`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
xgmCMlDBLPxWLVaGuZ7HLhr95fphlB03gpJe/evJT2dbj4ClNun4eANtutaK9IiVxYuMg6kmeOrp
60EfS4/r5Qcxn3dzDBZx+OFIy/LUNOu72+Vft/McI51r9SVQboCFixHXlXrZotiA5U11Q3jwH+23
k1cVF1NKg5JPHceu32yghvnY5VhK5dKrw82i3ZV9h5o0OF0fVrkCzUF1B3wWVXX1OMGnYr4WBkMG
ABqz3z4gOk6vYpZmyrYjkm0wXbZZEdENdV0UqRGZwmD+zv1hdSVDzCOT6IGfmbZsCoEfSUZYovnx
AyxlEitSlvx8T64Gjl5Q6AZph3gWXaDb/7SJZg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="l3po92ZmnO0pLgEjD+e8dDrGcXfglD7vJriM8tQEKDg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77968)
`protect data_block
9i9Bm6sV69d4xyOJWhFqAq02uWp4N7yMfSOa/jaeeG/M3la3VKKbV6ekHX1R3U3e5YPb7hloGwNR
AjHcTdYPbTyGK4pmvem9HBpGx6PLwDci0w2yy+tnvbXLRcfav23QpwDpzBgVDOmPR2vEg0U++imj
e65ggnGZ1P5wc/ps18aWSkyHUJZBQmieCONgmIshTK9iSgxf0B9KQ4SIhYz0vRf1Hz61z118Zx4I
t3JMBTu/zW+lM2BItR7xmQq01GtfPlhGFrKXoaj3IrnnOB/af87Nldt5iuInnFZ3zhUSDYKAMnEe
U+ckUZHTuX/s8tjdRK1HEwcANGfoTTO+HOyExbLDrYbYsTuokMakWwjgpWm0tJhH9a8OW9XQ/Wgq
KuivJyE2NkjQR9RRv1bUwSTjv+Trn3WSa+ip3jIhc10lr8W0vubhOEXLBYYypAc3C4h9NyEy85S/
E6PxSTk5bB6gaVz/K+3YSpBNoUIxdnADMnr1mhiOvyw5isF2WGHwmL6/z95w5tJVEJyS+vGFQtf+
SNfB1hMEXJo0Bd8f1aUQdGY3e9QiEYPmYzyKFS/bXzjVXeN3kqgdb8NxXsdZVRw11IzrL5sV2YuU
+tvjnVZ9iWiWKPGhEuJNZRh9KFcjzGVGGxxE+UDK0gOCVAMZH+pUOc977rRbjSlcw8JTpqbWMB7B
CI4KZzl5q3YW9OmGWPMtBROXc1ttZIDGOxBuz/BV5GsVpeGBT3wxw4nhE/JtesOs0bPVb5b8KLHY
mLFGxRS84EKcu4dCuWmcOoiAZ0x0DeiCJa3DmxObXMxMk5F1oRxNoM9L4trFgpWq8HD1vJX8nqI8
nPstYV+rH0j7nF3C+q2r/Z+fdKHZMPauDPRZQC49aNmviRfD0u/PXtaC1ApFHpxvQkiprbg6G66U
6VCG/Pf4TOlSbyeindptoE376rZtud37jOfm53TiQCRry82LfITnRBgGdQZWIA0z7iLkG9cfezNY
gedrW6tSNqyW4xBrLpAp63he/K2KV4eNiS1cG7XkmZ/0xnQXwZCrz5BkKjnM+W79Q3OohYY/orRo
c+g9W61y6nCndacAFUWOKqKs+1urf4fwUeqcMN56mK0LK5vsmrDOAqBfcmR/TAButD7gRNIzcASp
1/XZsqmV3VyjIc1APh2Pi6WKqkWRHiRkeJY86ssiDAhp+w5lE9CRUWU6PMfeAEMc0QOebxmu0Jgv
+M5tVlnFCeSBUBE/7oAHu5GDc6AkO9FPh6EoXLa0j9MzXEJRoqgDTF57rwYZi3e2rp4SyzlXT6We
kOrjtkj46nd45STVx8TKA+Djoj3SFoSdu1U19kPJe2MAWQaWt/rEs7H/JQklTfI+8ovdOPPSejLO
u1bLenpgI26UcxiZhhC/o2bHPV9Y2UQkDt5Mx4KBd+eu0RJfedekqYuckDL2GAp0IV+WgFF6nsof
dsO6PIU35tQ6svRfSUmaO/CJtlTu5br4vTzbRftE+JySiGDuVjGp3m3MMOaA2VGgKfW18Xp8WDa6
ddsi33oKI6lxiezf1TlANpuOfin6jx6s4fmZmDsot84gXfyinRq+5D2j9ZJZhUav1eUPoWzfjk4x
IkSq1NFP8jhxL+6KYD+3ysjSdJ9NlaEL9kq7rfq8KxsCO2oOCNNsp4zHd0UbEVLP1/spLM7qrSmw
+xc+LL7a9W31z6E6fjdnSgU94Hnw/2/7fL2eVbXZMpfjFWhozP+HCMIgbmq4omqVYzu5f/urlx4v
xtczwXjEIownRuH3H7u78Zlkpiw8xC6iaMgkpPnIHkzepLZvYZ5xvH2iz1WAoEbmf3sF3iv/prWs
wwFCkw3+Yz/fCB8nQXdl+nwo9gZqeXZvUdk96C01sz1p5kTdhfZg3U5kBskGWIxC2HNXHFDlHU+6
+n6h4T+ADqGxpzloJfinbItVC7uYz1Q6YYzykHELngPnfmNvZ4J+B9WJpHxeILpjOnZyVByWbvaA
wR3KeKGGK3qliw8FUidsbwr9IuMeFL6UfZiLJrMMMeGQwYYzqTtLMJpyDcAa+rzz77YxRedItXZy
GnR9WpqElRLPbMGo0ilKhTYuYnSGTt882oYvT5475gXtfrx5mBp2dvMqrsXvufZ/u6S2ON7rjhrN
1TV2kEBm2Ad7EXcugE4/9UCCQ4dsv3O0Iw7QNON3lxah6xIRlhHXfYDU/rOCgqi0NfJogK9FiExW
O6PQ2BejIz5BDG2/yBHPBQgBnHfQpRLW+q7cc59Z28NP2QGfRQVGbdRnsr4NqLevHRAUelYi2hhJ
08SKF7kaVooOyzMMyFxm1JrhoZfL87MaDA4aBafXPOynm/1BRn4NkK3Xnhhd5Vd25Eu+yURJhi3I
fY12jd7Kcm3pOJshbCRWGNLAqbYXGEtpHbNruu4vGElCNLm8U1GiGm3eQ/xIaiIBqPwCmw+5oEyG
NbWx995cSFlgjDHbkMPnMr0I2qA74GxPInxuFP+jD2PoHry/mLyOvSuuaYR2Rw36iDD5jc9Q5nn0
ezWeZ1ldBTDA+OkRsj/KZSvgOTVLED1LmccB0bvO9W3s+rmRyYRWdrKaTAkPt5rhIN3vjFaH7LeW
2qS7FWqwKM5a8pYBRxMB1RGcp4NLZBxzsdbbrnw2FaBUS/SE+BxZq5ttfhOohvlXRG8Xh7QIyQf8
EsH//OjGq8UvPf8kjXt4NtjcWE8kvE2NGnDB4efDzRLjvLNJ18xRu/EU8SnKYGoY+oLi6jWKgwjW
q6+dbvdmpGJSeH06NqSCaFTRnab9919KzpYLGvDEdx2sVlakeMITU9e6uBRFi95fQR0Mtqtvxn0B
0Nx2eH1RtOMMMMNeoE3+z6jdsj+P1815h2E+4cC36fLAls/KyI0vwT3ZMHahVW74k0eIGFm7fUen
2IZids0lZEdgvk1FCWNATnucTTh7IZTuUBBUrQ+Fmrj/tp4MSSiOeU0Zaa6X+8Iio52/YaDtSpXY
V8GZcrl4h+HbJ2hyBms8Nd0U7I8Y7Rkqv8kBdY77Ev6z/6kWY7V/mBMbdxpP28xhy7D0U+JpUDQs
QlENvS4iUIPPGvSEbE1NsUOVrg0mp2Wst8hkdXn0S2NEPgEdtgf8eU303aSzEZe0HZgmO+IH4lzH
7/ssY9BsMw3z2MWCtvX/gL0yhdzfy0dsJf5qrHL+X2tNoU/dWutPH/SuCCis1TOMgRoUx+XAu4wY
YtMhDeM37jBvvUKmgNQ/2uEHsZ/xFT56uC8OeB8lI1at7jsYk0cL6x8LsVr98dgI+mT1G46S6mfc
nMsu7TshL7OfNO7NC8ch/nzDMoycFFYljZIDcj9RMy/aiCrupsF4JoPvBGyMgDtqug1JuFHqE8+H
dnPoOKqBLHgLhKJwZVatoRcpoOAobi7T3HAiuYcDRjUYET2V+EwXf4cNX3qQPoSmSrjDMkm7qgOj
W6jS/zsaOM9myCxpkG2jYQo7rZ+lpkkYt2GWhOLdZlN3sZt5dfQTrdcbRu6sH87qrbIXrfZchyDr
p4ty8DM/mFOEe7X65ErUjjs2V5gsYRTzaknls+i7ZxkSNHBLsIVskaUQcRUc0fwixgBAOTXYq1Gc
SJYt6GJ5XGcvUUi0mp+0IwM77xkY9fQLqxsqncv9Pl+OwcF4BW1gtNMnq4B8ATFVEDaf0Rk36dza
0dyKyp80dsLY5XNaAG61UXrnlOs6X1M2pKKw5p4zZPwZ49/wFQY+zfI7c35nuZ5VwusGcTVPd3PL
R+442D24W62qJB4KMpC8s8h0pQUlZLgJ/+f1PTXjX4BFdPTB1WyaCrg1jd/RqO2AIk0vQgK6TaVl
SRIyL1nm4C70cRgrzRgLnIG4zEB/8VaFXWmZmr0ydH6pUl/BHD9soLYzahZ33b9vALv6ZV3e2eYd
lKKw2bDkHU/6/orY59jDGEw+VUwil3z+XAawHWO6deF0Udco8jKBRjuDjny8w3mU+Sv1ot9Yrt9y
cNRh49MWGm2Sar8gvqxoI+ZNMhWcVx9XezB73pUsh1kCogcrPoL//2OyUcymE2zu0EpszEXQL2Ku
dNwrbyy4j+ow54i/WfftLdfpTUWRerucE5G40N56IsOJUXCILde/D5y8jtuER87TFiz1/z4LUwcj
5GL+ib+MaaBH9BfeEqXbzQZ7XewYZZqve+wmYnKqAC27fR7fQn30+GetzvTf2eMxlsLKbEaQoKxu
lRwsSzygSpVWauYclyv+3OEb51DRZVsTkrPinKkV/R+WWAJKYHQKE2faaV4tDIn18JnzaNjAa17E
3OI7hXGT/qMKZwyBKRiU+xdn3hkxenJOAnaMO7xZXELFORvtL5xmuNufjSvFiYw8gKzntkHGupFu
ZS7cFblIJ9CxD9S3lX2358Sba4zfNH8UtlqFB4vCtkc4TkSaq837xgUZwgGNXi7P9yOncCtjpfTk
SSNnSrFVyBu+SsygLP6MhfBJqSxcSA7zAbgGhTA9hpVTIXxq2nShCtDN/PR2iSwNkJE78VMrqH22
HtEtpjzy3nDbmU9Vjt5OYWTRnhnCNW7fUYNTItauJFVaN43jFfi+xSLwGM3T0H9kBl8EB+JEjLWu
iSi8KIUxH60dIZZwC/cOmfOlPQiNDXkEdf4Co7yuW46LOTzhqpzOlfWEQd3i5PemJzN0FZqhz/cR
RdBXBCQ8tWeIIA0YgNFaXjZDQRISNS27oGIYfiMeqyDegEtQnkskL6sTwdSlPfo27eNgmqf7ZBaP
4o7QQLtknQVtaWFUsiDuLmJ1GFkEhm9/RTUo6qMGrpRuLw4HsIp0r6e9Heps2/ktp9jjgASVuf59
aXPJrldBpxOj5zF4gRZMevB/qdrHaNtmYEVZgytaQ8cVpH43wNy6QYy1+rV+D5kW0o+fWTXx3xI7
KM+aZVFFgK0LV0afBZ+LaDCq8wPluRL+7MqtFp1Yl4KcKMy0oUaGAxMYY+20wa8SmQ8ob3eLIsDi
u5R0PIv84U/btCTtCrCKLExpvvcO0t1aU6ptKEb41NC06M3rJIKS5QeQElI5Rd8cmW885KW8kgLh
XOnYGdF9cKKDgEJD2FKxFYLsZa7TroUiiiLHL5krJ6LprmM4NiStayK3T4/jD6CImjP+V1xG4miu
n/839x8hjBfMjO+ZuvSQqWm92CeqiUZz7hd6F6ocOKd5rBZGr7JB9usalxG44vhy7cGbJ/YsqAzt
Y2RmEmY5j4ezOXhYuUk2d/2LKGiEolj3tfOvBkOLlgbMwxp/IJYZZRE4NYtwcn532rTy6ImbXHkG
KXXaRj3xVAhtNl+Ap826sh3yUbCdcu8upviIjx2iXtLTgZY7/h7BGJ55U/r3qLpC2sRxho0Ye+YW
1q1jLcMyFDPfjQxmRVNR+TRe7utI6fr+U0IVU/Jwv3nqtZdSioCrQT2IhKdOe3rFEcqWoqhih8Wv
daShGoCsMtBGI3JEwa/nKwhyjimj4qfNaWpBTWAs2qWSxl08G5jDgLkiqgNJ6lxiZx6brS781Aly
PA9kLKWBM3819WDarN6kGNamb3kTtnPrKCvxXRke7RZi4vXO1xaUQ9hqsvoK/18lvl/WwRrPxOcd
UonPYEVhtiBDt8Nrlr67MadOoEOH66CCaNual0ICyiYge8hu/QOpjP7ChFdAXcCxEtPpF+ejhpYK
B1tuZBaDeB0xKHeLh0Ks+PlgJhm8F/TDcm4vs0sEC8LK4PCcYRjbgczJRTm5a7H6d7e/bPjxKgc8
2/bFlKEOra4wW9doTtYS9jI1YimJp6yuo140YPfqoh4eqxy1cwVZ+d9Z8BOiYpNztaWho2L+ukgO
tZ48eFt8op2ilQhwmQmRhVuViPdGMu8q3pcflj4Tsy8p7E9V9hye1FHyydIZoFee/Ihd2Aw7QQNI
gPXfHuS4Uoccv3LP0UMzNoDNF19cTTCoM3xGV3pTkLIbc/Zk096V0RqxLkLQitXcE+1C3IpBBptC
QlQr1CAIft8mRODMNv8mLaZauTphuSCbrIyHHip2CTXenCvNskNzQ78MFNnqn/C53WlUGpIl8TWh
f55+tqG1yTykBSOHXhO6UlwMeOlUeJR63YwUOC6zcZ/SqaagCc6AZuhN90NIUxb7s7pO9+TbQ+i2
5+yYREqfqyj74c8whMrrdfo5K7m+JdZb+p083PVhzT9seULxOXUnav/RLOeJClnj9G/BI2ESqYRi
ecVzwr1rffNxYMtPiDp0HvKOkxBygdqnbuGf+8V9tmsQNkTipMWqvrb/9kdffVvEbc3cgQzLG130
nkAo37iO8Rml9S9lBdfNfnqvezihXpDNIG8QfF5vgKeQwWECvbHHuePjITVb9MD5cCzyNYuNLIWx
es0TSf07CTRcqcIJDEMxfV5YgFomdTYSZ4wzFyoSQ3QJyWzgPTrXBvQAFDHm0ObmE+xP28puokwC
+LRcstO17vuaCcpX/S2B8t30G2Zux40x8skjxvQlv/VzeW0rt5ti55Lr7nZw3yS9Juf/pl6tm6yV
ej9W+ceSGLI5+iRItuQjD9My/cgR01fgB89/yZK0U/dkSxsmgh9EdR1MC4hAuKgqHZSJYOww6FTb
og2rf5vDM/riwBp466VDQF0Qx8kyPClYzeiLb/JWiG9Cn2IwyVqdlCAU039IRY6gyJO5xuzy+maW
peMNX7rfQ51iK1FF1zKWKfgotXWIYQZOKAKOV4ok6OiRMf0AfxheNZBJsMAWJ1WDqGp/ZuEfUe5G
0hVlKznqRjxf8vt4hjJx/QFebYO4FCJjCvnlTSRwfF9wPFFA3kp8E8sVbeFSK20klmjzEWn2vy6E
CncoXP+odY3ryyRW3d9JHi8LBlANdZbf4d9MLTuDZMy3x5NZChd8i7dTUeDqhul30a4C9i06ff7x
wFH5OcVwuJXy3Gi7nlR4BLsAzNt7w5H0x4sQHGl2fuWK60sD0UmOhGusgR+DLuVnEkEFcECi2ERj
zAdy1Tyrn7Wuhsb8VLHLoWBELllRPjuga5kefHaSMJe/sY7a72C0ntzSNvInFrj6h44Loop9BSOa
oLZd5XqitluQZaH7KYXyNLfu2KnHh1vD65uEqFh5tkTNKvVM1Fj6c5e0q8hydjbzO3VrVHUk9TFI
fR/HbTPVS6IbYTti3bQP41vaKcodMkngYXPBIccWzYFUCgTfAh/69MqrLf3+3QNysvQAEX2OY4US
kpp9C7W/Q6hT8VjHUPB9cSCnyyVZp1UVh62Bf0DKTSs9pglV2dkeSXNfFCZIyAMaifXSub2BtNAs
g2DTQVNZuTnoXrowE4S8rqA7DyvO0C2NPIuwJSrBhku57vZuEy/3+InJ6vhgYgtnQ91xlcrX01OH
p9qYNCeKctO5/G41fWHYIhcsTNec/4l/5oeeLpsDE3cuZ2aYRvfKv4YUxalM/+GUuZJBPsEPpRSx
CY9TKfa8i/Q6IhV/LURqN6U2Ki+bPF9x7mAKNvI2A7PA+1uN8+1gnqIRUA3rmXlLoiNWUGSfCIun
BvaGEq2fBicbUCoCJcENqQalsUEy/JnJSqb4RtgG45PwSJw2QlLKIMQVIobsdweudYNZjTYZcG/C
D7gNa5lHD6GonTMi8EZ0F/tIhIyqTvY531gPmHtzHTZBHCYV8/NIAr2nFWoWNSRuGHxL5p0tLmFv
iesIAl0TaIeMb3cWqetHwkC8cr8KNDr1oE5KFmgdivp8AjDIKqyScgO9bNCTsMCpn2b/aO69PAo7
5aEe+dQrCgJU3o8FbrGIyTHWvIzkOXFeM35f0d7c6dmJoclrfhcl/XLIet0a4novztOSX3DhyxoR
9d5qKQSAOZWziuYSxuKZx01pAjGvJX3/WyGCENrDJPvdfGtqeChx29P3oXv6lUrJpHXNXPemKDwh
yrsnaMKKpvMwy6A5b8lerBibjbmV3d7ZZzB17i1rBisArquvT8hfpMUxiMHW9XXxzfQRA6ZEKZig
FOz8nPXlTZbvCXSvNLeiJO6B1OHs+h6lCpEXRn28Hl1irTHiGZcQ8TmEf1272XmxKksAx1eZxBoX
nRKCbW9M9mPLpuJ5YFiL8yUBYnd5ES/1XCCJ0gUFFoZ9uq5QDWTFXKyyOvQSPlFhzXXrzLVPb3fC
syPXvnhsbvjTe6ktd5cIFYtjyIjmyIr2ge6YOTCR7Lfmcnqk5dPuNmNajQqU7QKQV3Am9IrSFixb
pvZNSmTgwOOi8/fmkRYuBpNCgR2NwyVuHaUxvkZaJkPrqV92ZmTjKKDN+RIDe5Ipw+fYXBt/4CP8
ux2I1pIanuiV+R3UmkZ/JlTKAhyhLKEBJN4n/TS0Y1AbPpL2M7hYaPmv65MMel46nLT0t3ucN5Kt
DeDfUF5B+zjc4CDX6R5sHSfSr9w6T0//zlBCIEateOaMHIq2YvEf+woRU7Zl60WrPB8YcewamlEO
op7euE6TYSJQtwwoSai4vp8AS/8duV8qi8pbSwkKnvAn51UwWK3SSyD75bRZJH0DXQFkMTdJqR9M
5ATtzX2vsbkofW+yJL7VMz7GnIXPMJMdzE3V5vg2oSwW1i/EOeXGIBfJCwtFtK81qxyT/B4FVy67
IkVJl3SlTyjYs4oXl7E57n+m0Xti/QCHqeJaXGLV27y+GzXJ9jw/rlQcFImhagxlL9qIzRjPmEgm
k0hv4AP2zuyyRH4b4w6Sl949CbLkmXbso61i3vXw/cYQ7leJmcdFN6GOIsCP0+JKW1JEQElrar0c
nz8ydo4A6jNhHonKaWa+1Fl1yKoKArfek4qn/Z8R8I+dPQFkTJAnLJ1swye23udPS8/lUI0eIArs
UhoZMmaYp/RPmeDBLYA/5BV8ToLkUI021bjRSi+ZRzyeJH5rJ0gFxylQnKTZyVWM891QFJlDrHVM
fw/bKVgg6Ztk0c2S7aJbnSb/dzb2zWBR0ukWyhAudvA0EI9RmDbMSeq2A7zkWbkuelTr3GgiN9Kz
coy2klQhNQA7YlDjLwBGJUKyo4qe0ICJhCSPUu9/Aj8/BFgCa1QgcBtYsBhOefXQAsfCLqYBmyii
hShVfZ+5rBTbdZMAqjf+bWRFIOgWxvx3S7uf1Yv9nHVWi+mqGGw/C2YAF2d1pE5Ovmyw10A3e84A
MIZ/41/6pnpPMCZPbalZTeqiMynaV7akWirBh9YTUmA5jPYISq175GxpmiysjgorKLPGt2drXwTk
Lh7wxVSEz0zLt0GTfhi1vqkKCFF51NVh5sxSM4MboTfHRL8JSIvfp9HQ2Ql1F1D6eK9544DZIa5Q
206IG8RRglyI12JFAgTFzCbvwcSQJJKOlNyv64s+xXIzUSsl8M00J1PlIOqVUpkZ9RNCkdVQB120
MslZd4zldxxj2qBaN3lYXXKZVbc5/KhTapMXdZxSufULSNAmOUAokuVw4AaisztH51gnRttcK45M
It0mFgyMuq4nZJxp0yLBVRDyz106mfEk7Ph/aL/5Rpua15vEgJDVD2LXH1DlvBWHhM8BBiHKJsiq
4KgNdTPUUT/smFw+8CUiTKFeyn4y2JzjAFS14RW1bnBNkPsSXLGnzyGQibgNTsSFbvtqoNN9D6gI
BI1uznNI1G1FEfdS2wrIlVnp4r2sFBBrQdtSsNeYOR7zpjroIv+ybbBDB9+k4UAPhBdLiZNXE6g6
A57Bu5ZyQpVZi/wVe6hZ/FF5JvefMeI7IOMMED1AEMVOhB6OJiI0FY23NQzw2Lw3MUms38weZnZm
0BHwvXnXyo8gn6rotMfrNVtA5RM3wldkOULa9pdUpO3m4Reh3ZMGAFneId7MieMzTTAvZ9q5aOFS
9Z5Wv6G39Mu2MuJcvdFdtoJmCYV6iz/hKhdjCHGFJMRTCpqR1RxxSnSFzvj6JwMnDGAB8BI2m7Wn
zuJcdCeXO8ksYKg+HbWsyqVJdCMdOKbWsDVlzlwzpp36AFpr29esQclR/xy76+x0/JaMBEM47G9d
OMIQauc/jsjjZV6TmXUA+55OEPtW49z3vgCiBkLoQ27wRLRGwBZsiRlGccSS5zzGgD/cd1Fntt+/
m6Z4oCE+SXWMc4D+w2uTWC6xcwGYUJXbc34x6OQew5jpHjlk8iCmayGprp1Ou30e1K5vJnQCDkWZ
UQdUK7PLlLyB7Ezl2R5rks184QBBfjkmtjisRFK34SRr6zKV2n5vhTBIupBzU+R38fywslYPJje6
3+eJlLL1mrB7fOK9mb7/niAl+21jcV9s9tt5vtjGEVY12q8Z+v9IxFYBsDWdG+MNrCw6pdU2q79T
jubBrMInY9WEjNyeSSMBaAcmvkzDduxec9qhNGYUKtOVbgtRgYaEyRpg7uVCquyu0oDyQYB33UXy
kQKWzlLOFfmWRjOZTKpyL+UVgDk/Cf4oNCmLVvzrpxd9Q8pV6MsIVZshYtvKqhdYZ0UNvrjb692j
s7nIVQFMgyHrD9hLe0RhSAROVv6qYBCEO28uOgSc+SdnfApd5CXpTV4W2qRX0h5atlaikOSa1JpO
c5hk61lXwER485dx0T7io64kKNE+jHHDOJGvEk2ueBCpVOkC+tR94msJfF7nG9mC76ncQPG+9N0D
EOPWTBpn+5uzTSH8iatX4dNqYWsbGybHuEIcgxBfD2sr4uhJOR0i6p71yzNIQgv16ZaWbydgZTqj
/yP5hlNeUxIyBQErOemBvM6mFOUv5oLncYgphps8PlaZgpyNHlraQBbQHiqP2+pFD2+MSAy6nXbP
yutI5TdLmvSewvKi7pABshoajvfHnukvHxP206FShGVMKLgsex4oZ588lZVO9+2j7a7w/hGlmn6T
YW719gINSxVg/CKgAPpevNE2LnJmvYrV9rYjqlc6JVhbi8Q1kbn82agpH2FAUD8v3aiebhTm8NsV
2n8Mc/3TdGDFrjcl2VTjrTNZNNFGNbM4HwT1I3duFC747YoEk3DgF3iJ1rnlOY7FguLApO717tQi
DUkAxX/tO8RM616ZrNHif4pmfeAnd3dk6hj3PJKyO2N+ZR0rb9ymv3brGhwHefGmTg20NJVJdrkX
uNHprLhQ+Mt9zruPiLFDiDykomtc6nK+ImvuYmHslIzF4CARccyh6R/5khP/wHqctBUykM8zHjxy
pntslHZwDLWM19wVbq2T30w15aJkoM/RLRanm92/OqX4h5Vcq+hOj3YXRWR6JZP3GUO6y5HnWqeT
+x1dZP7WQB+KCM4ul6afw7uOVnW2R7KAibNjg8XmT5am6ecj5c2dDapWvuyDad/aid7VYrdbIdG0
AShXODThdjJnLqIPv1j7oClEz0UsZtZ0rq/2JN7aRDP16Uv/9+VW4yHKLwcfscttdd530DbgjVxI
2ExMpptf86CPFPjo+IlU0iD+Hoo1A6DCL1hdpuESkvfFBf/HIjBW/WYiTLjl7foN7ZPeUCTn2FgA
XiGvGNYY1rKfZu9gUW6Q/1cZTdDhGvpQ54JG5d/Q9Oq+SkBK3PqLpZvAs9jWDYCQIM2i6IZqu8tY
8vdG62fhOPgXeoT7kwpgLClT1EpbFgvxNGPn9t+5Gd29W+fnAz/ePxIfSuMVNIRcYt3+YMf3jKIg
XkGONwHyjonO7ShVfpUHUvCFlvJN1jgPOmTxZeKQpRpxw5f+Qnsg1H9fk925QlDiL796Ktt1mrAJ
I6AzZqfhgTdJlkcRTzX2+63mXtDkC6g7thnIs0j8Z40Y+td4wKN7RY9p1VDVrdABCErCb1PN/TUR
l9SlIXoNaaWH0PXWixbtyUFgipmCe5x8Uspunit0hyPZ15eDlB8ojivREJ/FCAXfrndObzslkoA0
f+IrbPePMSsQnuWdBVB7c8SbV1t9RmLJ61bm9+T1lhw+ysg/GRyxWU3x740OvSaWMRSQDF3Dv1c7
xwzN+ISz2KzVB/zuMMg+rrlI0yl1MzZwYkQ0bJivO7WpsIVO/8cF5sXxjNateH/rHshsem4F3VZz
EGkWGfUeUXHHmYCbI+pRDrZmD0lmzygeIvmZSo+ywnCdIM7itF8G1f8jqepkA05HAmVG17iOL4Yt
0pYhc3LXEJe08AqCa8ZVYPacAf1lN5OVd6YZP5JwBvZeXINqVCST5JouMXLwYqJjMiT/PJdLlTPx
FqyIPHNB7YyPsjUI3Iulmp6HZlMt4UAy8ZlNqAzQ1+nr7Uj4P2Lkk83vxw+DYsj4YfodzAVoIRKQ
LUcKVJlGG8+uYs8k42pRHZkUWEl+Boe46F0jH1hUsg6q70BjXM36RP7cZiQR9lX22RXwboLRqBl+
EmFk/HMMJoDMQvHJiEgU5HIN6cHugJoM/55hgSRKCH/fUXRmrpre0reSWIbBHHdjsLkjy3KiavQx
zAF8HI8C9AKIybHUPxmJ/lbiR+TK513aQ3JHjnCZI2z24jpEcVVI1/KDNQIxHWhnqanMzSaXTNuu
7BWOR1g+/hMHbNCFPbdIEZ2qPfkGpET2+rT6S/b7+RvTDw3cFYUyTLui61j7/ogtBOjCDoVagFiX
AQ4DX7F07ftJrcybo7/ZVxMENTvogXzIxbCw+jbSzLp08/HThwLY3aKABXhBgDGMXB7xyus9t1F6
4qC/NMF0TScspY2CO5OZVDyR7elkoi0Nxdv34/jFLDQ4ecoAZYfPEqspKTfdUrj5tvz7H+UfVrb9
ODBGWZ42KKZoXgQZZX4qytr5pYOj3k91wmwnjCFy6cpnckaR9lHNZhsvGGqovmb4z7emLSzuIFBd
0NKDVJWRdA7lJaaTGHcFM2LGoxgMLTVkSd7sWjGpHCNMiSh0Cm/gkrFRyT2moTc28R2r/Udwf0wS
HqwOdv8MG5L5R1HwqAJvz83wmwe7EoL2bgqdFeQ2sw7n/K4NZxxYUNV6KLH2X+uqsiMedogmrT6p
mNuu/inW3qh22zgdHsSVAhybCJnx3A9fmUMWqMkh3xkJfYXDy/V/k3/DZwQY65RKNSVDgqtd0Nkv
Wb+X+VGn0wP4Tqxp+o9WFnINSGkABF6eKfHL5I8xwsimuBCwl8Nk/hvDPv3IMsRtaLg2oKtLbq8J
E+GWbeWwMDXP4gNImFWd6p8IChtclhRoLq9ow0N65+0WNu99oyAX99GTNwaQP41tUnnZtqvc4ELP
bWXua92mBBNq7uCrZYD+S2UKFTX12TkM8Rb+rv/rVHI3yr+KO/hFwrBwYu9O8CxA9veTFLdsIPQD
PWCwap0acC/APMMkCYpsM+bSWm7QlgP73pTlZlEgMz8ZU+qptN0o4a6Zmjr9EcMHRXczWw0T51T3
wQxvXKhHnlSH/XxBfP8UEC3K4BBqn9sIjp6ITxWNfdBR9iPmpBTp381VitYswxeMwaJ1LeJ/mfub
ec/o7fZjvLRNFdM/4xXePpy0awqkUAO1/McIRDrd51/P0KqQV0sZDXH5PzMwH0YW+Akr+3yykADc
kITYuYhdwiwp4UaDJIqsfBU7NxNLxnHvaf05LVG3w2idXZU/W4iFew4RRTL3AdrnG3CD2aH3teTS
mgnXJRmTfkH7r8P3uXU0dDpHn12A7/CXjLC6McEJ6aRaEUJze0urIYwAIzbrHgF2GWOybVqd8r8/
5JPbHmvW8QrRAYx/VT1dwHIADI8rp+k+5STbelS6zTOhIos2hQgg1MJ4JmJQY0OS3Ek76irG+7CO
+2buKGqZJPTkQBea7kdhMxqGrwh/YYuWRsFQrKD0ovDOKvGMDORSzkwEi2cizSN0EKwjj7ohTU8u
e4o6xZY9eKRQjAvz+s0XhTgD28a9D0PnWbHs48XbUoTMaqEvQJhJKpE2D6zzynwqlTIBtmi1bUmZ
Awf3MNf7K/JlP67ouz5p2ruzpRPFCoC+Kz+RkUte1rFV9/Z8YONKqCT7Swh/29SQgvtzXgmtQCY+
3vXTewkGR4gioeF0kQms8C0bWXtPtAVPtCNkEkfID/XEi/x67Y2hgBQg+05niZhLWS973CYa8Hhx
m9Fp+o2z9rBFw+PPkWvcA0vCo6TF27O5EzYtGbnp7giQjip9PKb7d2jXJp1p1kGYs+yz4J+FflAR
ed9rhDzUhDHvFAVj1u3j43UsKdqlN0NGhr8/Fhbzfl1uZ9TqReEyWU7xuRlefCzctS26xQ3ESAMW
CmpaatK9XLFTw+hUz2QdF1HPR/05N1Atujps/vUDkJ7ghTkJlN/y8hpn8QrBoVoLzNLvC2cNlbkt
pegLnAximZzCn8bED7P6FJ3TbqYNee23WY0rL3qxquOMTQqgaUFlmqwwhMJin5gNZF39qtcfe7XQ
OoUlviIYdGkK9WMj86+jSpA1ixIRkGI1hu+lfuiLN5SzedVzQwbHtTgL6jyzkxiNDLNjxqU6M7YR
NLHSUKgpUowEnhXqQJBWn9R6I+xIOiJz2s1I9vuMhdsXfN7zgRy9a3zxVsIpzRbVDA4BA8ycxxda
OmYJP+yqXEveCrtHwn/WGs2Wl6TE4aQ8Eze8U1HHI+JeLu4AKe5eqwSHIRujeVaww4kECWsdbul2
J2xcYzmNXvAVwVT5Wkn6ctICJIxTF8CMJ2K2LfGnpNXp9QASMfBjACGLhCrZzZ/thp8gvgHAJ+rs
BFVoCxm6eE3T8cd6JmvuWTs02fcxiGNoRCUt143YL4N07wn6j76VSofllCu3BP5C589S8e4heyRy
Qi9fxC+m7b17VC4aha5PdTUPMG3iCcNTKZSmD0ZoOLLmkKqU1TlJsGQG3d3qkDqQFfkjH29zvNeA
awlVhfcDLuwHIDmM7KJhCk+CWpFb2VDQ0ePgfhfcPGUKV/8aCQ+GxE3UvUeO5zevOWEfYZ1kBiGE
ONBvBjPF4hoewxs2dKn7d0GEQ2wTaF4iyBcrNnpsAClH6BT6D13jCXXCbJ7lMg7KIkyNazoCJknX
AmzJHxxQZjLDVqS1S3XO6MChIDITOMb6a0kZ/fsqKv3DFW3cxy8CwrHKA7mDeRUPGvlx/m/nMmNJ
6Hgzg34WV49RIaIBEYx8njaau5e/2kecXAKMhcT0AuozoLyK9aHbY7qOi19BoTu/J4XdNMxeQMvS
v4Jl1ZAUPmsC6b6wadSJWgFIIPSo5Y0Ay7NV2rsiCuOyilFqL+nuK/dIm4eMFoYo2IglBOBYaCWT
gGjcMLa+VaUV7fK2n6b1/nq1T9KZwVzUMiSGKkiZ4e3e3mub/7sKfKaZrJGtAMAq68+L2N5aJ2fB
Avji2jbeqTsO4GS0Xexd4HB0LSnotpA11artBRtIRuWzs8hr8Nk6Qo8N1IwxXPTVZS5d6r2jF8kq
XhrxA74Yt5nO4VO6agQSNtrYPaRa8VMkIooN03eYPpTgWpBa+r3yN3NzU4lMFI7zRBeqoef20QPx
vwXXmwnXfIzdA77zk+4sqihacJrvfK1dMkbF3rh40IL7kl6nUHP5T8EefnB4Y81LVuKPlJStQ8Dy
FGNNy+4FeiJYa0xJjPh+dSKKPO5ZApIpXoIVgjq54V2b9qrC9ANB3d+ut8DX5j5s2o27XAEDTazk
arh/pCBsulL9ehEP1MQUfeCkOx5Lsbs7ScB2Hr9f0qdADfGG2SksYrAk5k5DwGQ9LuZbjiUmrzs0
ch6gAVLeKdz9+2SckRr7Jz2B8gwyzAEPCKG4VMh5DtHoLi0hZCJNnysxHZR20ILbMj2xK1arwtjd
cLr8FjW4OoHbmuXN4kXe2azxyS9iIG/wnKJ+PiRbcifm7ZUbMnE7o5qGZvdk7puLgj4eR4pfDOev
T4qaR/a1rS2+cn6YqIoPPQVvPw8OIcfO/M0NbI4+GXe/AhMwrXqPrEU2CoxiX01Gpr/eIZzcWbdF
//LkKM+EugLwEGf5P5pg+ktPrnmabtXxzA0iPxvcK/pjhOnhXe5vzaSF85XdLuaKY4fNR2gSyl+e
VPJgDaQhRaVVv7OUWIUuAlXIvTZktFIENC6SvhIpiirmOW2dsmevKBdsqZtZa2nXxbAp7d0OjHA+
rOQRHWhaLMvdQ1pOdZv90DUlIsZbUM7Fw0NZl/lZCV/4v2HUEa2+iD5G6BngNwG8LKWz+DUTLSvp
Fw6Ga4k1oSUDaGvwGkDMqFQSsr0ETjH/opTIwDmEGPW8Zj96ZAKoCmRTNoVTMm+M/rHx1FQyk4c3
75vKWI1UyBjroEc94+777hbebwbNTddzopV/Ro++yPQ4c888Eq7QlCSq+VhPYf5YN/NU7TK5XMhm
lqs/TQ/9hrNMcD7jmwPTupsFQAfqS7cXJ4j5VLBHY1A6Fkgo5ZfsxSrlKRdwWnKJlJ1KM494af+I
aJdziDisWugZybUAX5FCdIHvAgqlimmDYG7suqOlQ9TRiLnwyIWq9pep5QHOzgpDg6ulTwOPzvLO
5GG2ZtOc7S7j2R/3xQ6AfDLeXxLZqF/anIEYCtLBm9yyPPk/prQXPDwsXCzubCdGewlHV6J+XLau
cEBFdJJGJcrXzLgcM8hD0HfuAxdyGz7vzoATCMWrpJveGyU20vrHTN6bFWgjgavbRN1rAbdkZ2xk
BuG8TnW/1ZuW9oIOGiV74xHoIHCBE7ihDFBLgXCBms1Pf4begFRJjEF3e0dfbu3Wq+6S63YlUUhP
OCyt+XcRXCGnRbAlG0GZXMryerAt8EPei/EpKv04Nh6I2xpuNySkGnSFQXn/CuVbRCCyWA8J32ny
lN+aCD12wybiGrSBvBE0JFYrBWc2vEt0Bc83w3TsYCShcvCeVMRfLFj0RL+u/0rSka2shnCJtGip
CrqifEYfIpJ6OOg2kMrPL+MKZm3Y4SXl2HFC+CxgkJJpYi2UC1dF2uFv8UMU0TQMxxg0lbl8d8Mk
ty2B025B819DVPU8t8f+IAQ+pUFRFUNRu9oZCG9yjs1etQ30ge/Xv/ywFEhzKR0VawHDGwoNrOwP
uWOgCwn6udcNatXVZNfz3mDeQiJUheCxwxaykeuJPy/QkaQsrvO4IluczBeJJeM9yCFYHg7FoDGE
O/3kCMUZSEzaAbksxuv2xMyClhQJa1g6lZsCblmn0KLv42Ll+KGszWewhCxXLvXsPYkTcYnu2OkN
I2QwHka3HvF0HgA2YQyceXzZMmfBZ9dG8tpKA8SJoQmsYWrwODq4dCnkf4foJ3KEJEoWOvWTawdm
X3j1HH+ySbzehrfOtq1vG948bKclsxlhvV2TGYfwYFuv8RHiyhwqu31JADt2rg9ybxDUXdLs656k
VdGdb2TLcYeM8fL1nEGCBcdkZtBAvcgriPuP2N+P1YKtOuDiv7m36hJ6wzmch/+CyjXxZCwbTi1L
SwXie5OyYovPeVEOZEIae4AhfctBw9Pc/xmku/XguQ8YtBmn0Br3SQAJxRMuQ+8s+qpw0c7pq1CC
FzISdnmM2Jl1M8t5iCI+I3z3Q4M/m3jg2KB9Prvkn+QzA0rnMtABKOxYHboWcaPnzKnJI/NfDVha
dOq+fNxa14vzPwJYgOid0R7H9MvRe+je0AUfZFQRBuc0JJOQCwpAPy4CpkAS9gY+bcvU80O/Ww9O
/UT222MDcXcxCpzSU4y6nSwTPBBqGoiiJtwP5GcLwaUkhyb9y5VXNK6xQM5fhSq1x2orfkmdHKKk
sbs5VrdnP4E/XTF04zxwsRZJcbYNurbBLVU2/31d6Qt2z96GqRxySu5q+Wc9wgY5XbKSeYdmh8YU
FZRgE5/H1imK9KISuK84OAabdfI7NjNzQ2wVhMNLe0naSn9vT6Iscqe/ppMtOYxA0krw0rM6Os+O
/kEYCEZRNIe5Rcw4zx4eLwmRVtCF1M3ej1hInZ/DWzGU48DMiFt0V3DcT47l9N5wLVED9foMaHlm
dSHYcgIv3pz3SYXvDKeaBdXnRqGQkb7lznce2tuoalwa+0LVjVlACT1maXpa2g8jMV+sJMoioIDQ
44SkH9x7vXXyM+02aMfLOzrA9SOzaFumqEHfgVUatHkJOCF0iVpMX1rhlLSb0adrieIR0L4Tlk+v
oVHjUM7dYDt9rRZ9KwC8zPcSpkHSxxMBH+RjUwoINLRgu7iyBB/iu2JwL1ZwVTXm92et7cdlhpYA
EcgIL3s+O2mbiB3W7FoY1xsn3wQt7vMbuofacE3i7+ysyBvtVJcqH1YEXK1shn0UMRq7Zrk0IL09
a6+coOzBUdDym9XtoJbKAvYB4ACRhVP/MGgf3em+ohXsIyr+nyYjGs+7EhEf89PsMc7GgllgyiYb
mHacBiIHhYVpNcJISvZv0nQgJOSMQRa4VPNdslmt7dmnyPNyYVCNq+RRT34VQImYxA/S5w6HzZ7y
u9zzZcLYeroyTZirc1yGr1fb5UwTlBzfhRNd5KXMM8y+Mdzl3q6SgMBGGz4HOllv+kcgdsuAc/QO
YSaay0F54eMB7XkKMjxOklKo4T/D2TJA30y5FMfVINsfrPgOx0YE366k9/j6G21tE7dBdzNkdaPJ
B0oUMwViL1N1fUwmSM9YPICG6LeDvHuz2fFAB0CbkwOgFcUyB62bihL1MZbLkB8GBAwc20ZrdLFF
tGRxVugEjvfO10JFSE49NwpKWLBox5h4l2UXgInq7yv9NVpYiZGhg9CBJGVnIiDsJvuHeApFsS/C
kUMfSt8aGm6NLkiNlaZBUYv2++KOHYaZn22sDWHjXaIHixds37K7Cjs+R641UBQAdDnFqymynx4B
weBxqCFFSqkB3epY1kJj/RZb8G8gZ1+ohMiDCS3MRayPVKtMk1WGRxTnZXKbkor3Mos1RETMJRtf
YQqvV80fEkHluB8No7rkpFfYPMzZ9qnX2xPh+4wN9K0vjDnme5vey4Co6DdVVG+KT3qJ7fm5lE4e
I4oPxo+x/maK755W6vIXbyZwlWmkSytacmo9FIWlBgUfiIjcjrhVmjlsj+8cpV2TgmX7YEedPjC9
dr6WCXFVNo8f1mjS6mvz5brGsmznkQA9edMEr1ccjjSpjSQ4Wmg63aiWS7zVND0677IG5mKDGrvz
xs4NpCRuAaqXFG2p0q0ZN6oFFBZ+qe3UYth1dSs56i41rN0vsBHBInHk2Es4Bub91ZP0Uri4fQkk
KIJuaclrGh60Z1RO3F1a8p92DPS9KngLQatQaotz7PRGYFxHaMUM4oCdn7989+mK/43FDTAfnq9P
zezB7R603GLxO94v78a/2+iOk6XUpuvQqQmqCmePuEvHKK+mpiTCsKK3VUU5VQj1WQgBvCh9j5yr
FmBFbrXOdXtPjDp5hE5hcGWQNE4Upp/VxSGRJnqC4TZE2bqRgFOB2fqLRT4zgaPYCoLPp7Z0aXwM
JHqMy/ffmHjffdEHR3Co/lXlQwSzxbwmFPHgzMxRhLUL2yQWeDEfG6gDeF+PNiNx4Kp9pgBO3EYq
W+CxD2QL8B6SWZ3izNzkA3uE94l1e0u9sIuRXDDGnOyeyleV6IBgKO+IOAmA9AO5U0m4i3RYNilU
Mh5XOeqtHqm7bhc7lM3aEl2gt0g3l4naOj141a766+X0K5J0hQ8xa9J4pJRQ8T8c0qNyYfmAOroU
7j2Lsx8vOSINp9h4YVJPfOiXI1T9iDvppJBg5oEVBk4tYGkNSeBhB/WP1dpZK53EG4MUZOGxLied
62zUiVZ8GXsztKv9r97HCqrbN5ol+IB+Rr+LUDe1K+ASl7nRmlISCWfuVvFZtJu/6lCknrN0UPWt
wOeNnjJRNiWJ+MDqmQ1o3HFgsxnFO99EZgJzj+9kkDIVg17Guivn8rm2gCLP9fAjx/tmWLFB+6Gl
7tlYnt31frFBxUHLJLswFGUvPiS6m0JnrH2jcUOPoybpsHatSw5x3NIhoMfdDg+x8ze23K5pb2wd
j6nY8q0FwPKt5OlYwX7nda//OGdntGN+RuTyJvNXYo/l7k0DKfLuIYh+8OLZ0NNih+pKH0SzYog4
LywJj784o2FTKnVZo42LND0CmOsXK8kLW4OGSv9WSKK78EbZdjUx0vnu5n+rkahZ/eb+R+EAhwaD
uP+kk2qDsmh8N5ui87/BighXkHXkOP6F50hXVcuOyuc6ynm7158/03qhIQPAiImcGsfmyTlCUK73
vRcNTQG+RxMhEXB8nPoJ3vegTNQIxAgVjcOf2w4CLGHhCL+ZqatoCG5PxCc4GW/ta4ZZych16cYF
rTVkRy7+ZGv/+YEvL6d9Gd2mNZON5hZQxB8+w5w16HRN4WVgvWF+4QUE3jnUEDqbUubm0GN2dCXU
/V0G4qkzp0OVni0W7G++b/fjWT4xCPnFeps4SKr9yK+Wilz5vGrd0vPX21OXCOWD32yfbjSvCNdn
6swhd/Tvo08ZmD5aWEgTwqiJ3ZofqfI6xTYiMaO8+G3R1aPQztqY3Q/Won+7jr5Gv/wY5RYZEt6q
yQDdoS6dopJCR9e130LENfXQw7LLcUYJ/a/XvkDKaMbt4K67+Op+a8rnQ1KMRTDGVkA5NY8n4VPd
uWAW0DQmu90WCTV5gWBybiXlGIYf7m77sBNT70MtJMivSMjoXLJw4gd/IPO/ncLhP51wQkSDdHLA
z2vJIWRp31YiVFr0dTRBoqeYR4J+jHMLABVg/inPoe9TGcKfHTbgAjy+/3fAx/QdPOaLf757GQgu
F09DS4SoVnOfeID9jS6d9drEoixS4M+mIIBuqTscm0+yq8pbcZeZg2382xBjRzUeQF1hkcqT9aRj
aB/UjPBRSrA6xsFRhvT6gyjf3zveS6aCnc3jb23l2L0bgafgh+ibYnNDH9oZLlp14noCx5h3o8n6
KWrE2h/3LDg3oSSx6g7Bk60tYjuF46iTTUEKXdj+Ij2becZTO/6CgqiHL7fJmjf5AL71IYR4vnQQ
GVLetO9Nxe1HrqXmVJFSDWNhJ7znbMiq5b07lR4ts1UcgnsC7Z/y+wFI/iBcIiDS837vvURV4t50
LshmuHZIDGHo3bw9xGBeEIJb7Ic+n2sQ8C1JmCb92d/xPmVDAeQ/FTm4xpVqQsmxruuQb3RVDOvD
oPgnBd1ytdpSvF+iyEwmARnsHiw7vljy5doO7ZieUJus1O52idIzepV9cSLNYupXqEJ8VQHTKaEf
0EiAnKP70aZSyaXeXZo5I5PnZSikrTo8URaYMKcGyQGO022cExqYz6Mq7UeEQeMyWh17xibwbZ19
nq/LJ3fAcTsPySzF3Axdh6Z9wOrKupzTVU3xj+GcnhElCw4ED74e7PhxtLfK+LfPK8iSVEClJSEf
SO4kjlttb+Ec1jzpJiOUouoVqbR6H8/4XvZVkWgEPfOIw9wvHkyI7iJ5g1anWJEt/OfLRfZY8qsk
8yp4UWnvYxbHXtW8OPrX4W64H8xNRJ3lqflZr09WLO64+MtW2QhVdKKA3WXt1dAHeuhkVzJswx7z
mMps4XoZ/BGYn981Oq7xZI5/epi8e+etd5GM2wInsWDIa0TJGPtPruca+VHfaLElsFPeHGB2CJDO
CFGxlg8O8HDQfoV5u8rRf+5K0TFeHu0otOWqYr+slLIXY3OWxw3Ko1P8bmOSIua34bAfnMpEI9dl
ma6XxUVHA0RKUexB3paLsQ14y72tZkqS0XKrU+KZ4PV5oChWd3zvkWL2UvYqDHztlHSFtTWqjX2u
gMC0IqIS7hjHXk+zLXGupwBNCib6KlvSVoLJBTl0l5qdPFL8Pf87xb9AX40JmnKLVwZcxC5c5DOZ
ESowxR1oQrmWlTfCtt57z8H5wW4pT6iSFRo+nxBh/5vrnbOXmE8AIywrlHPu0SA7RXssmZSLS0u1
qtsi3b6NLIEG/YMJecLj/gsc2eGwIJJSbwNyDKpP0VLVrMXhMNZVOXcNEIJpsmJD3VT2A2QS1GZv
4xDkDRit0IqfQoYqc3e44Zude61ykhH2TyT52beWyk90iPELG8puuCVBL4ePLvKuGQMzQ2mXK4Im
kSUW83qCEZa34ms7/8+XUoeFCOsIDAiHjzOGj1VGUtZPRQAKzowARX2EXZwl8MSZk92m5Co/vevv
WzBYuhl1zn74NWfbAd+4U6qX5x0jSn3OsBtzGh5mgnzQd5Nki1FydSWqk62ViveacVEU4zU5+Rsm
dfOK5QNh0Or5pz8qGobn/72G5X6IXvUCw4WO+eW1GipL9xOJQHUlFiTA9BfSBiMoaRsc3lwaaHYi
ocVMqPTyEJZOEBMywSwsgUfP60Wz8ixw1G26oTBgxsKrJPfg0gQSbYmxfei9pjCXB8qGWeA10djK
4XVTnL7e8ECm2vie9YvsgjCyZJYx2amq01KUKvt6baLl9D9WRvfRFBtg2xQ5VEN2S67YueVqTtpB
z/eleTKtDtTPgvdrwDGKnGXmDUxYEJue1cfuIwSAniu0VGR9vAcuPn3eFXb+MYieiSfTxFQjwHxy
+8uDjQQp9tvDWgY17tOuLJTnHiKiKQXnvD5vjvBFigN5vcGidWyySLQsc6KMEiFjoz9Gt/rhZ/MT
LvinZaNLHnrH/cEM1sZyJ4mLfvf/9osK8eSvGrK9D7GO6tBaAgC2XWG/yKd4b2iiA5ZRdcaSfNiB
YEiFlfg/e+EBavPyZkBpMKhxPnMY+j0bZE9pi166QXuHh4heOeLIG1+Mv8mYmp+DVz46347UDgKZ
d1ThkcaHl8NZ4bgwEJSWFaMDslfOeLfHpuJTpBUy2wxaXlMOY+bXWd8NOaTJl93cf7bn2aQIjXKC
RoTsR9Eqa4eW2kxSUfoHR5aKmATYwa2turgWaynPS0Zact8r5mq3Ed3zpi+7c/g+UCqz4RSQeAW/
FbfDijePElTHWT5u6kRlnshHj4KQg8HeeW65pRfxR2FO4y8jEbn882SBVhXNeeTiH5bUSHZr7pUE
O6Qp2F7MQoik4eW4u0jvjT+xz/n6+MUi/DfLfOCNstba0dPr6kv0bFIOESG5mI9FHL+icefcl96+
QG4AwWj3xuhymXji5AyvkAAgK/Dxiy1JPHy/Drz7OaDHGo933GWFV6m6oeeFxQa8/2cBMYKuBwmo
tzxlTbqlGDVzWHa9SfzC3RtH9w1K9MQ8UGzhEeIrZ/qtHAvZWUJuPY+rlzOs6P2C8eovMpQMA+xp
Rp1r8fEma+7hkK0bY3KWpeKrALGPUVE2sp0HGTMcqteoEBxmcKCfOkIAZkagJavqGZLB6GM4GPjo
u80dh1OOGdS159Zx5TzREzh54MJkBps3jzc87EcWTrU/IlLYfmECIfNqqdcvULNyMyQw1DZeSp4E
/tf6RowZBrD4Kbd+FSL2poj04HgRF5N1tEsmxgg06YJ9yyWyEFrB/C46v5GlGOC7sBtjjdRYnsP/
QZCI7eDoXUoKNTkk9uZakc1TyLYqQndIUw2pS7ekG9kewqOpVGZ71ARSloWy6Eqezwz8Inu/22Dk
YfgFOfPuourZ5TQzjyUf+C201ERmw5iSYpFzSL3gtWylAE0Bmt1haQr0LysWh4uhrHbfXK/BYfd9
GY756phJ4NSzDrqHMH/wPinbx+IycMhbVZpAwUTkOOCDuZ9WulfjpJonfQl4vlf26n65rrR3Edkh
SisIOF3U0CjEEH0tL+EwlTqZgA8K9Umo9zrv6+DIG8UGbCfuHXxQWmT5ORgoxXhnmr65vnVGckw9
OcgPfVYv7ne61bgz09ahsDR2kITuf8XZUxaUzBhpZkO0jVy8fCpXmhGpbSQtqxBwMqrzCtznk8TW
TqBbAA8Yxl4CzozgCMR00/FB9B+OWcLFZtitq7pN1hxNxXEsf36OWomu5Q8T7SxjSh3nV9ivyhH4
JJSMM7gEruqJlN//aOm7GhC22IMm6It+PZ+EhHpcTKn56M1Iick/TAwZlXqa69CicY463EJn1oCZ
tca0EHakt92uI87Xy5KsO/9tA5vokE9NTCXEaeUALlAGcuqIXC5pbGP0j7TPAW1OsbOULt9JRDUB
9KY2i/IjWPhuNqzDn/J0ITz9F3TUm0TZMt78dkyv53HQ8KOcraPyAvjz0LZZy+/7REG9pexzyQcd
d/prGpZlDyrnOc2VYeb2I/pgkoXBcLP4YT0iqgocAjsR911wUiLWFvz0rfZRGAbFh/yIeNOZBFGK
WYmMmMXcoqwBK51ky6OJnje/oje1cFKPOQNmtSi4E7+O7KKRGBGHhGojb6f5KBJ1rM7NvgCib1eL
mDZdtrQrx80/Q/usV8bVJA6jk7BeAT9+re6IbE7zYPo/xsU8ru0K/Dj8QZWKRo5ox5Rb3EpeLEJ6
vBwVC/hqvqVYtResvVetgWrrVYSCVyk2MPIHOy+UxoriUwEEixVohSuhoLUoL9fr5b/6EK6VqY+D
HXhR+hoCviIeY7k8tnrzwGxE8Cm1ltPjqvDdJjdrz4Fg2vfjymniDdAuuf6ehJLw6aQTkCcB74K5
iv6hMTx8G2+YbCYxX3efrdJCoeBYsCCwyipiRyrx63IEURRukIxm2u7AUW1zVEQhguxbptqXZ5Mt
brgbRiRj9MAGTY2hoKLvbgJZSQba2iiWh5WHciBzLusAmMvKo8sNv245g85FKbd5yCqQq+hbLv9U
aWV1S67vPrUI/Vw1rqcjo+TPvBpACmqJmZKBk/k9R9iUKB78shYceQ25j1QjU0R5NLZ1UEnKRDyH
7PKq0CqWf1Jc7jEZj9NfxcR3CfuY3emM6XlPQtofiZBJMgnmpy3HtfRADASdVklXx4ZhwGEYw2ad
zUvyu+OdzQOShQD6nFtx2AUCtKbLTheM8vBoMDypDwOs/OLyyyNLxstLBWWVgt19ZBgKsRF6oleE
K3iBqGQPyXY7IBGvYb/G7GmPnPiXqqFlQ+RFhf1lI+GV99lMui7r0zSa+4BjK2XR3OugufLd0sBK
+cXYxFvLmdGRVelDMQOiRqEHsIKOl8yDSlRy6RptH7m9gy6D4m4vLEEmLWKNIjQH9Y1wj0ithEln
8U1JP4slhfu8ka7zOb/LnuAmA3zg2lVpK+vQh9cm33Vliz9oQSZGjs1pI8nH5sEcEeu7zx5OrbDP
c+lUlM8j0wxMCCmMVpZhStLbnCEDmk2eGoepvaBeBsDwTg043h/JzfRM5uRM8dbudIDizX24vKmj
X96hAAeDUB9uDdRIOPmiNUUaHgApuYE0CvnKJMHQgTyWOWLTUJN1xAmh7yomETC9+O2H7iV5ffma
XOcvb6KAPoOsGvCG9kzE3xGjr9A40wq9ISOD7cRglf9XnfXlMOOZA2oP61DqKzk6qANtv/WPPQo5
+VaSyHgSkqWRUkxMQ9R9GAgzFmR7TcW2gu/kYdD9VuviLV8B5ocFny8238f0GEIJIOTY6AU+dnCA
2JGlhy9S0SDtEW6JyNLm1uu+p0QqVu9a3iYj9CfA86SzvTlT58ydfDyf5fLHdqoYFj/Ajeodhk4w
/ibDfYvuADSHo8Pu1Ul/gPKZy3e5PbGflH4PVmj/g2xHIbZU08EXFJCsN4M9ROwA3O5iA3gs9xPD
wQh8Wwv/11cHsoWfm+iDwc4lXErvUzw3lFerKiHWcpBTmYsBj9pMbZnM572V8M3KOg9rhLPJqtJb
xbWMDNmcs7JwvKWDqmpOyi5KgzY8M04H8u7I3TNhb/ULc2cqc+KjB4WZE6kyt/1dE6qdQK55fyUC
DlBJ5jvRlKoW37UqP7PrOcZDObNVncCZGYqZ6eJXv0PtU8GpXiWjOuz13C+Sgir56Ir2Zd7pnKdI
0jdu7eKvG8GDblbs1nnc5jdsykpekq342Mj0Htgd/M6Xn8rTfWMzh+r80uX8LbJRupvF6A+ZkMXq
66RuOoq2SHt3kHPKSNXAuEpPkZBg1JSC3fIJRGp1l9Qjvi72IUVX0t2lwLqWFzOygwgzhE3lgY6t
E+CElO/kXtLbOLggDgNae//h/4G/Y8NUV6Gf5SnMrv2deRCp9NPubokOhX8maLipLkA/Zj/Z8RMI
bRRPIkEz5W4Im+9/Frti4TA03Z9YCRfRP+4aRvgEsUGOtb8FAaHKLbfFB3zBicqlMbAVASSyj0ln
hHgaf+2efxRtt6Inpdvk6FvoFPgzfGZO5SdbvzWZeTRg1aIW6Kli/cat142ED4fAykWMAC3hjWyj
LetzvpiNLjSmsJU3GIOjnAzyVXmXkTQsHTeho5bRqfUA/8ggdN8JjkoozDohBTztXWTgSMULti0l
Rr47z2F380KsxG6lT/KBB44NSiSwjqKF2Rdf3p6nsFa42Q2YcA7RmtYfFN/tVqatpKVXQoMYMThx
iCZD6KCJ6yrwIzf+mxvmRDJ2BYr8y62hjHo17Lnn874KHBa87dksxsjz9RTsO9JNuBauZJWjoY9V
iug98MVdnyy54rqx9d0AU2e7bQ6mC/BwykGZ+gOKfqjWSZFXpR9FC9/DSy+KURfXqEkJJiKOYIO5
Gn5OQXa5gKE2cQhmNWBjPb4VymRiH6k6qi+WA89ORku31kH+hVKwL6yOia1jCY6KOj75IGIRy0TX
xEWl4LlSLSseQJVEgH7a0a054i37Ml6T1oTgOOhyuNV11SZ0Zdy5bqPV7Qs3lFakn0O6TCcEC5vd
rgeJcEAOL8CObMKxh78inTeClE1CFyU5QUoi6nU8C+0a/6T/3Wh9gBkMYiXTDpPWm1Gz8erwvHpp
EvHqWmo3TQ8MbjXmef9bFENOBgp6gUxiCDFTtUgt/zIhcU/0T8tUrMLiEc+/XkoQ1RMH4QvakHVl
wOtpcg0evi3vamXzDgaLDzdzSffF6C/ILuj2Ns4xuAf8HciOjlX1imYRudzeIHi1g/ZY9IZS0scU
jK4GUa9dhtVyMw/43glgOwbwQly26Rvw5FcF5juns3dl1WwDF4mL4q8x7n7GXBNa9Owi7MuA/pbj
UzbKlJ0ctry1hp/qiX0KHdXem0up/F8JmOhkBjNBgG6377QHlX447HsB5mSlx53uhAVt6735PrEc
DHxcvFYNsxBqeRddMpiwRd2nOgJ8SNj+swIwpn3a8GNPOSrMGrNhQ/ruNMj16jXb0+VM/iNvTEiJ
1IwZS/KLCabAKBTG3QeKoF/yxs+89N428XaqV9stWx+ZhgXJXKsBhSjaBVYsF0pr+LN6cbSt36ru
BI67jrkGvir19teY0+Advy3bLarLZzUozPysym+wGAFj+WBYr3Qo6DcVHcAPPO2qZoHfN8gKCAIM
7c5FWpBT6zLzXF8iC4m1n6zB2K49gKwvcvJBQUYxh7WmMfk2GgHeThLVvLBmsmq2Hv3W4TRBzImj
K4hKfU8fuR8PE5Ta8TKBkJH/+QKiiS+wjUnbeaBsJAHyu1BmH9IiTEOEDF88M1ycWP8rp2BDS54p
544usAkksdtyLnnAVTsRgRiMhAYZS/Ik7RiEYoyMAhcDFLITH+fPTT+djVaMuTrvsdSX56j3g49h
GTU3q4tLdFemlMV0N/XPric5lu4mxBSYoemIWA0gC3v7viDHy9KcMX8peBDc7s87CJe9I1yuU4Dm
C7fcMS10ERWqJwSK/O0G7/AL6V0Ax/pestQQPJfjRJPIkv1Yrv45HTLRlbkn/EZnscj9qiiqwkdh
seIjnbjh3GBBiLtfEwjKP2vvwW1fmAkiXBXp0IBZb9Tx2IZJFFD5uKCG9U1uOiU/T8MDt5W9o9k5
IYU+npwtjQzIUo7fy+bxzZYgQZ/tkCbHRcsRfrRI7Yk069AePFBO9SK7ymfAroJoilnyjIqChbuC
4qvGIT8pJCuCa2XIiYix8orayqL4+38fxh4U5SpmjadV1NpHyPwnKFc0z61yWk520JYEAt8AZj59
+7MboTCo+JFi4tlY4AT4zKRIZRneNK6XRrtC2syB0IAS5nRIvsu2DKFKuDHBf/NH3V9jh6xu/isC
AiLTXR8sYaQPt8xdx9Pvhgb0Svd+CwEDziwTml08lLk/+nUHck/r5Utvu+Eq94a1wEeIXdvoh5yq
oeNjdIn0g+V35JHTYVQVRFuAvPN1Bb9UDEofZHPHYeDmNJG5xQ7qrirxeCfTWtm2iNkq5E0wsARm
gyN2SaScdFEMA+bbqd6+9/G9rpXPlxbhf2oObRTW6eItK76MU0vd+b1BGD8/NnY5wE5z6adDOCyg
6ongppNvBaDFFz1P072p45c+I6nPlAdzlUggzo1KQoywBqH1M3GgWNFGu3iblw9lckVevZOaDO+8
Ms4VGSiKm6WzIWSy0OA0RlRCOPFnTY15FP2ryvXGEglfhK67DZMa/B8oQ/o8MRUp5waDBCCLCCCb
y/z+uu3OfHtSx7T2iFI+/upOlglT3FGonFaWm/77GwMPxDYJV6JlDGbyeuB7DWP8N3F2ow/iOdFc
XimSh0rTZDsLt3KPo0Nk4i0WPAHEtOdUcWbrbYN6Fy+4opEi6/frDS7P86IxEhq0HQjdPMuIB4se
Dhovqz+OGadQK5vNHPGsqJNiO2v0jqmu/uHIeh6lyRBwqH7/pUQzbuDIqZ+R7DtkHrykde1Lui8L
4LtV8fRYdSppl6F6YE21sddblGxSQowdE0DCrW3svuiGdmWgzYye28SK1pocSHRY0ebJjDSngNFO
hgviigp27NnSObay+pW0QtmCGLdB4LEnfLzY5l112235JC9qhXeryTAcWcuZJKgf72cWDGWLQX+a
KlQk/uR2q2MN1sI4En4OnQ42K8DZCNqb8kclbKFbGZpfPW2Sc30zusNh4dm37ES6Bad8eM/btDbp
S8h8OZnYhHKlZGz+DI0lwDj7B+eHeySO1XOEZuTCXEaWMVCY4RyoDWVP2QFSTo5derukPX80W+pC
LdTNM9bVcQZEMq8iRhCihvYLBzq3gjO2KiyJK2dbdP2hQYz0c1SPzQ+zM/zJPiobdEO8GoP1c4Kp
j6IRZCiDsg75W7vPuHhDPFzZasiTKahIUQ+O8Zz9+7fMtZ4vqOX4imNk/AqZdYH1E+PCicaCA+1r
XWVyQ2XTixVGvUv/rn2gLqFiPo6uyQJTAKEAtxMoPfCFGbeFdr1iUk9IR1WvQSimsCx7IsW9Q8Jw
sY6R7pTGn4eg6sQgpr+7MPEozLY63d/0bp4A9Ez9y8dDhxJKSimYeaCnT/i33ONBMWSxFf0o+6k/
+lJmloxuFRoXLrvpoj1DVU02AJtwj+MNitDP5OqNpC/RCkBPehCsirsWg5jkFouKBdz835NTA+Wa
ov5/RRTVtlo2c8l+lAk8XCMS0H/ViQLpBDdXj0QpUketqFIwXWckNmoaR5CcoKAj/ATEFFc60lWp
Sauhn6R5XWL7oALIyeJlVNTocRhkA8qMZOy1m+eYDu5djgSoZ6MJqO4Ovh2v7J1sfBUDO7B6orwW
5AcKXeAH0ZTHuc5j77ASO+g1cnteJB34ftRxLzUBtLj0RfIKv+6e+KRBXA3ZYjMO/KgjlhgL9aq7
PbZtbUsI4DQYSNIhPMWGlEeXm5D7wC1g/Nctb/Rs+6N8ebgwaTUoUvYDs/mo+1b8OBYKyWm9+NDN
XOcjssDhazZclTyFeHIpl7nf34tATLTNT4hFeUhC9Qp9IgvWMBhPhJGjGpWsY45CBhstcea6IRWC
wlxnncNMEXpfaQGfNoUgh14lA2JTXA3COoh+BP1sTtoO5GezC9Efw7OA1PLm3UsAZcR/Pc5Gup+i
eTWgQ8ecsxcuh5nsQ/lskWIjxr3nPCdEpVG66heJUz8c4uny1EYMwmqYtDHaul7uv/O2fk/P9gzx
kcrGYvJFeGdtH0UCk8/51amppHrVGYMtyeIuGjXAlKeqsxiTT+BRbWZJV7D6HUg1XK823fdJ4ioy
DTSLyH7yvLtUsfnZyvveqjlB78Ew+5MGeRNgdrnoSLLVdHKcguOyr7KdZbaQHAIfDBMn5ly/pKrR
CwvNyvXsKwxQGUTqPaWeLy7MOTwsNjwUVJPTYyiwJTL+5Lu0TnqEFfotXFethJK41zdnaXtLMxP7
sHo/K9cJHMg7pUfCrMLd9XYKaejbPkYnuzyV9RM2HSPmroUjh1SYtqWksmjM+tKrXbAj7zC40hAJ
dttWUE78bklQF3CpzIBGZizFou6IX7EHTO1CopkK8n1Hs6vWPNrPaMqc0n+OsqgisRRleUFlAr3e
kZjGwFhsDy6Vxag+NzADNpIQDG2CQg7LD1+wT6E23gVIWn8E6GKiW4HArXxaYPKfLHWPuO0OTXaS
jFr3WUG5pQv4kAw37hvmj47AzCHcF5DMSkixVZ2avTjaSPk4qKVH/Yr0lrMvXLGs+EGqjhsPsK6/
niMupu+yWCZVPpiivGzVfQ23as1fQJ9Lu0kUZo1nC1LrOWAOqNS/jppID/tg7L/pjVgiQSV93mFT
jC8r8ofdVzPlyrfyXeory0fIDMFfa1d3XyxGSiP6rgwd/EpYSJ2+Vz/9pvammo0726B8xlf7wpX9
JQGBwuk+dd3wdNrKbewWlUOEyBWfD2HmV1+xQKnOf0YsPUJvZoxBLAhaATSlSkYTkCYF/WW7FyKB
nx7X2JRfrbvJog2E+71lnGPh+4j3iRPoqIIW9+r4hBKHIFs4Z+2WUyWIRt3J0RC12oZkutdNQFAY
ihCyTQHdMb4PL52W8d1b6TNmLDk/kLxf9i2zG5cc34qkC9y9kh4ZGr37D23Hy1n1bCpV0qX9HTE4
kzklElHx9x2T8pCD1uJTrTZpfcdU1LsqnWmBA4nVoZ73u+DPZ4Tnd0UNPaF2si5nGyfk85P9UMSp
D8zkHPJnQuWonESmzl2QZ+lNTq6+GFGQKcCbT/VoRv3TBi5oVCHZdsQZO5MEn0bWNWABIgMSf8Ni
uN4QAvoLEzgXGC2llzbvOmVobKCSdsrfPeh2D78aYmPAw+xUhEhTs/YjWCBOJoNmHXZo7k6HgLrE
XFR7aLDcTr7OsT0g1VNYJRCehrTamGrpsKV99DPCmYmOfJxEW6IeXJLRaTX0pqPWzO4451lWBgh1
+/KRf4TKQayWRJDKqXWN/1nxAY+VyMt6U17uUWxhn3wFcAF2Um6wxQBJaysAgFWAZulDrACp16pt
NQl2nDLQ5gvcc361UOG1XES/aVGmzekycyEWf3BUsv6BbmS34WhBtZXbOYAZUTN6QKAbG0d2osxh
5FA5zKkrOc/hDU1G60qLP0EVugbkZlYnOcqSbNWswFePkGyskRZCWc0owGgE1uxMos/WsijaqgqF
1ySzGV3TDgsKtIPPygftnlAZhV6HrV/5blqgZs428UINYehXJ2GS1FonElj7VFSMGz3czsKxAFvh
kqXB7EqRBP+HfKcxQIkbPw+wZDqss0B7+Al9jjEJZKlUKThA6n7+lLpBTN6GcYEg4xZaZ9p5sqV3
ou8sRPwTb9n1I72p/VMLRpryV8XucCFggGjjLUEjtz81vgQomLjkBDnI0N2xYSo+0pD2TYTCEVHg
LmyLqgo8k75fCp4z1vy2V0xzB+vRKVZHtK1rs486XIjUo6Qs3U/S51+sUwovfQgOvWSOb5jHrJ9c
8nJZ+qj+32XASpPDLloGoYLmKyvBRk+jtKmj+4Llk89fcqMNNEF+AtpGclT+asS8EXihcgkugBzK
xGVh+tq0YjWJ9WqSkm92HRUy8btVURHUN2CfKJiGsZh7pgaz5EnKuAAtFwnqRUQPIMDPaXrTJs4U
suWxFGlEjmLUADLjT/rD1WNemnoOYZHKO5jr0G/IKbAE6S/m9HBn46XCDGuUN9KISQntptOF4dzc
ld6dSrviwX46edpO16wXz0D7nORrLL+yJCAcAk4MEEBafoZsx6j5vj7XJ9s211t+H8A4VMT4BO6A
cGcPW+JImkTerN1CP7tYaauE0zLdcvFDscnae3Al+6hYAMdK6WT5n5qqzFmBmooVmRkc3nGwX5qg
whOEzA31z6k2CyfozmG0oCvsMurcwZKUFMdIsBQ7W7Z/Lsbt466cHtiqPPkxlDxA4Hn27mhczgIE
5nhbrfq6JmPnUx3vApY3Y3xL9Mexn7itCeyEnscCLjxk3F7YOBDEJgfpb6GSOXX5OYRA/pYzyti2
UCdi2bOTHlHyY1Gh5TksY7kBR0okjYafU46Xf3vlKsJbPTcaeNEX2iMdtVP4BL80iSvWNoBBndNN
aRyZDiKcvadxhFcmRgyW7zNSNHRjn7JquTaGCfFrkJAhqiSe83f4su8c0p+A3Dqef2m+noxX/HYx
Q0dorgSATv+ZjjKxw3VWukL/Amr0bpu1xH0VH/MRUQFwJry6dG/vhVbg5t8NBHk7d9AMdmK+LPhW
Pfh6dCq8nML0PnpW6Pr4h4hd5EKzaJafNjfIXD92A/T1IGUyyLQXBpNVeslhzz9fv4asIqeW5Fco
flHL2ZMSeFppmLuP+xw7hvSka94cKPgw9BM5UC1Cfj9jFpa+d3BDhFoPR4AoEeYtjeDvPuv/n3EY
kzb7gxIU9/cp3lZvs3W1FbLyTp5/R1nLEGSaoqAYYYlA2ObHK/YYsdTBZHT1kQgjTELo0rCOEAlx
ctfWBUGZZtjeInoriDAMAwrW8GWEPVmmF02f8YvWNRloa1XGqO+lBtWixEWfW9xkypUXn5HW4UVJ
8AbeGZ0KAhEOK84Sf3Mj1hSBVM/tBCUK09binxcJKz82rAIxUV3cN2Mw4/OXTSTkTGZzNgJPpE9R
GqizjiTjEVtv3FW13etkYGRei0zks9PUfVOh4HkGtEsq5ExuRAfThj2LGCddDLSwFbm7wpw9X2N8
rV0P4j93gH7bAycHMrTAqyce4EcPIZ65hhP+oanchug22CH7gZ+l8ohYWpxZ3vjf9DklVI4xtcME
H3ON8/orE7CsZrCEkpgq9hOi40hXVKXNiPlEHrUZyuqFEOHk0m2Ngk7n/n/5iJonwLcx+FsHgFxo
1qnOArkK5CReN7jZlVa+HqLk6NTeQx7HLSoIulL/Ko/qxDpBYxU6mJB4rJUbewqZ3tGPQMVhClqX
u9xk96Mc+6Xd8CT+sY+dkaagJ1+QZWP0CUJRSQsVOWBSEckzbOmNSJZZbF4+45aZkcIgdmCIaW4X
/VaaCZAkfJuhJkP9QKE5600WYPdDV0q7pV7XjX80dTJWFdXROWr3JuTdl27f4IF1P0yLilhNsqeU
03isnujhk4NG+ENS9I3pjN9v/hfeP1VuYHw4J0eZbxBHZ2cTojt1eRJkWJVJ58YNWixq/IUnm1nu
1rIJgtQrkW6JSwBnlPLHGn9fbYl69z1O+WH2gYfZWRwK3YutGPjBE4FwEAgOLo9KKeafcXn1mhQy
45i5vE4RTLzqM+65Fl6SBILf0NxohOupd3nd9uvHSGCCznHvrocg9JpkrGuI9LJsKW4J7aM7hqMf
iY8SXPMftX0wqKYE64QCuC1rMzRFzlVECOdQjMrc7vXxiWmYL9zhCXwhdYewmdhpI0mGC/l/Uaxs
NrC1sbDgGiMso9XujuaKw/92w0z+gpseCe6ukQO3zSbmB/VUB+nsB8XCKwMGxpooznQl93HLbsxO
i2Bn1P3RB1pMEKIiEF1+uKGZtnK8eaTK6tuoRAP9flCmvyYsRgEz8l9pfFuy/egf+SxixTFUYMrz
jBWL+8EgYz5R0oFY0z3YnDLjdNu05P0vlnu0AZhkXbeuxh3JVO1V2ZuN9Dj2LCbGmQqYhw6EqlmM
mwIvhmxjWwvrb2VFckxqkKFYx6V81g4Kr3hyE0gZt2c26009V2znhGU8kW2LbeHw+3JxdLPEVZiU
F6q7OGIWxSVRmODi4d+vDUMrg6UQeojX+Cng2Wgvo0vs+7n7IVUCZivUFduS02OTsnEytnHLH7Dv
Fo2WWEGqGH3zlZwzPacvn2L9FQCibWAGBmKX+u3TRtypTLLUOPSeoXSCH2YVJUiiy65vFUZFh5Eu
mHMOIommpqL3yJxbU7VHgjd8bFnso3IOJZxU8QXj5lAYqz2qpJnP7jo5PQcRfqDlp3k4kyYufuS5
a3ApWBoMS9ic/zW+SXpF0tPd//+IDN2C7np8Dypj5W6qSx8N9Jq4sRILZDx2JQ1NfN1C2zc+UKUr
AtXGCSarPWC2XkvW567erHuN579ZYTdxqNq5zlCWUK7WzTrxOnSabw6BPECzKpYuDwC/V9hBmKqJ
8DLqykgtnihXAfhe2Q1sFdQ7TfokFoFmVxn/sNsTri9qVaV3g2aSy11i3uY3oiongdh31pZYtmZ6
rGKqRUlAH5gQPLohn2qbsEyWpunC4jLYVfwoE06OM19xnrPHjwlvBrk/xxzDoBOVlqO0mzCG3yAo
s2rnviakYfdV7ZYi21dJ/0xOM1COkeGvfkrqwlku/psr1dMjxLaKAlkapzEGbiM2FE6CiDgG0v0J
+1WXp8OIgEjZhiXHcvzda1ybXLNdu65o75eunyjZPHTxkkQ8iTACbH12lQvf3w6oxrRc2UjeuM5T
dMpK3FWHE1jUpSDpZeBRWyfsQEt3BeqXlMQRZy2F54PTQpj4rYvrwmiu5+FILjAETZ0fNY6miMlg
BR/++VvLsnUle27t4qBfx88wNOqRXh/A+1N8VpodjGtGu2fkq1JvZ6P5ndeJzORe77I8agjcMDw/
SBt3Y0UaILFykb0XlQKyPsa2IaMwvMs8AROXjCPpq99fRXdiZLXDcL1V8M60vZWD11l3TweO5kph
fWt2M92SNG54azv1qbCMJCcZIQyyWIgNbdZtQl1w9AMj5hBfXuq57eZIVQQXKLarkK++wETrpTaQ
wiXNSgfw1nlmeWTQlwDmiakiJmp58VcONAm0ulnl5bM+wjyEufKs3fic1KQK7w+imc+tc+h0YwCL
dXVFNjIvjdfDBHfPwy12YEjVFki0pj78VQBFTGR/ADL/oot0GSM2HV4UcFIdhrwlURKwx6bAruD7
kXCcvdyYxkH3Z08rACdcsX+aIMdK6WErSOaBj6nzVxg+n1K5fPlBZma/umuaTra9RPh0kKj3gY0t
BK22JV4WfUUemDTbktNkfaIcREsQP4vl3DsfqOJH48tmW355+qPAYHOgIgPCrANWll/n3+DqhQ+3
4TJy7YWosTasQDh2/7dOgxfD30meX/0CWCdLFXXxCxVnAKCab3Js6j2jeZzEIQM5eqsXELde+L2B
LmSagaFSppXjhZLEh2cJeS7kfjA8x9jQXmP+CxIIIAgj5/pJyd+4RA7gG22ZhLShNUTccHIR30pH
RFZmm1i/aNWY9OhOtXoMlef28AfIQqRQxu6Dr55ki8F6XBVE5wJxWYdpGSSKVZzavynvb4mURU0E
jXUKZUKl5ScTeq1yED2sXnx0ndnBrVX2uz48CSJDffSowECafnitckgedDd5j2v+h+j0Zgx2laVr
wGQfIV5qOMpF0ke0QPprnrbUuufMAplmRfmr+MP1QbshQocBrwtHNQzrah0/nK+i7U0wjglG0obl
8Y3IiDjipCdgv5dPv9j3weYG03S2b27eQ0G7M8ftXmGYVXzSGOQxNsvyBBiDz22AzW0Vl1a8eS29
KIDO1QCIDkjlgoWKGs8Ti4G8Rw4ci5kp3NZ6rk8oREa3xjFJRwpd8RHFwm1FJxxIZIs/2k7NNbJM
+0aruXBnQtI4ETz741RurziDclZ/69r4Q6OQUN6QS5R9EdZy7QIUWIXfaIGuM6oukZVlqp/Gxfz1
dEbyoFVnN2C0poMJ4mbOjkEiNC2sr17iZRx47xb+ji2gTLO6tthq28Y6VCRdttMvvn5dUY0RGZgY
mRvHasEMdTzYJ1qWXJF0ipLZvQ34wnfAM9g5kiQrt+ugZhEqFyKCt1wRu+/IAWnjgpQRwrDLMQq3
ScQf6qttqX6OlkoPt1WD1QTyZhE33GTI1Tpw34Rew267+kqnGWD98SgBCCOIn/WXhuv+mDSCXLFN
7T9//KVNAc3N+9lsktE41yzeUeagr/FWHCTS2ICjhraw/q1ZErTQukC541du9pOcBhzg7fqXBgjM
V/n8g0bKT/Xpu5NLsuD0Xr6/a1jNwkvWKvUTrGNChiRoTsJ0wjTgTDoMZRmIOcF1gSTh3bryWXTE
u/Km/GiXBCQV00EkDMkX6GeDOhsEPmkFXiDnzJFmY3iP0vpDZFSdbnxnoltKpcHWqf/N56UZ90x5
5FRxHZfJFFn2cSTd/e7VFWFNqHu3b4ed4JiYyc6te3xKODbNLgRN5YzBFSsWpQeCASV3yGZb1jzz
yM5SPjA9ghEz0O6/nGlZJhruj1x9QDdFr8VAnsm0dFfBF1a/q5RG+tr8h6//u1YjeIghK2bFCi2l
JNrCCqWW5mZ7srAUzSIMW1lOimqG4VC7ZTqd+KGE4XpQdfYoT9TR8/el9QSjorEaCAG3X4jq2hB1
PqJwkfeIo0ryYdsGmGHtjg1nmsPGF1sSNJ9/tX/A1EiNi44ut1HV8rrPPJ3134hEJGI1Tdklv+2m
VyrO+UsHgifH9GDhS4ey/h4yNRC/2Nl0noE6OYJwrtdeAvfzPIAz3DV3EMnAw63XnhSKWXHENLNR
7MgWvayCYyJegC6DKvSWbU8c22+ws1KJf10o3KKpqBXLTFqFpD6QflXt2+e7V5MydecBMe29/8l8
IZ7Msw5gneDlS190VTgj//+osMlrMaJwlmNgGHy5DjOoEbYZfoNOSBVk/SpLpc9rUecLT9VXqzPq
u0YN1eb5wFQye7cIpE9LErxV0wpzuO19j1qDtlzjZXPtLEH9wjlramZNxzlVFQQ50PalPO087HJm
dIK9YdPgQMt6V0KNMX/Gto+fYiU0uPZF+BSNzA2NEbAoZYkglh4WAmU+oWQ3+yvKLz46DQTEIw71
LoyKL0X/OOIjY6iQ+uyz2adRU+HQdPXvM7tyQUHhKo1rOLQw2l8I+XBKwN0P28YZH9C9Y1iNSHJa
OaY7a9lvy/ItvrnpEVl6DWTt0B5Xi+MpFkrO2WyTdcQrcNYP5MMacJYJa0n8DD38fiy16svxtR1b
JTU/uxlIdbIMui7BKMmH1MhKcJ6EB5WlDhZM1n7/OCojh778LGx7L6lb3QIzh6Q1vPZxdBm6Y0tx
sEeLZ3Kpo7TwccKbHbj3PutRtjsrh32SQ4cdMNZfSpXpa18WPBIDgV9XPr3gT4MLYL7VynuCv1re
y9aTON3hqvN3ancVAQ3bWW8y3/9IjbkzfA5fagecl6nY7o9/aWB4TM5RNAG7wS9MJWlTLCoPEFMG
HxbhtxEFDwuHqWXz891umosdBPuiVmmlM5Fe9rak8aFX9Zn1AsUFoDNjekzSPx22INbAkxUQWuLS
M4QlG59io8XWgXLn3cw9YEMjSdE1InKK09a/gJMGnjwKynotNaztJLbIV3YXUhEHFfslOsOeMMSU
OeA0Nk/bMCSMW+DaBxl98mj4iE48ZnDw7Fojy00n6NLPTXXJgtKaAg8XtguV3Ow4Kn6EnL1obKTX
QahH8rw/HWkuQeg75a/1bw7ZZ8sNFC2xQu50qOvhwl+SFgMHUEFw8VL9WbnvCEoZ1PYVsBbd8G7R
PoX7XHFhz050fciGMGC4QQ0zjTAryFDIr6fXnyZ6609SAOed1IJ3a+CxTyIuLdw3va0lbS2zab2r
f16lFbApgvKiNmg2DSF35r89OBdey5Sm1S0v9PttX9qtw5P6QDi3RJROCt1HBhIDHWoHeynFT4lR
fAi8aWpAiYPCaeCeLoUwti9gF+eEZTpgF53iHtZtGYyaxEjcv6DWXZMItaKdBuEQmZZ4qVxipXeZ
4fUo84lB0c1eLbOFXcHWKAhzUZ16e/xG3V18Snw02Nhk3LSsVil0g5oKCTB52yBm4ztk3vRV+gQp
Z7DqZkE7Xs1jLp5YuS0Qts/h+i8/0tjPL/PkogCM5mqoMKmzRBPvnJI73IK+F0JISeCtidFY6+sM
lEXUIxSgFPD/ieHZ0KdFkAGSESmgRp/lKkNyb+8R+v+PE9wk+LBhT7Zs8Wz2FuHNC0GTy6mOFdBw
muI9rtpUXWkS684kNQiGWNln5Nt2StrNvt40anxbdkTyDZro2xDZGuNQn1CBMfLVLN12AX9Cd677
vnRjQT2kxhANdoUkFPt9MAX5gEXp7+4K8hFER2VaaKrw3ykRJryePzXK1SLWzTRdxnlnlD7sjK1i
JXC7UkeQQapFJ/EsfMd4GR6EtBJJbfPLWSOwxiNJhM5UbvDNYYapAbYhl+w1Nu6TUKkE+K61BDmr
bgNUj1dw3eJIIk/fFtA7fKWUWhc2TRhpjv/qsVWIFdfpoNYaX1JLfRDghoFlIM4LyGXTXBnhXCqs
zpJ/dhYtqutsV5zlKS8KWv6/ifdugUeAdMrKaay/neA0Sq4+EdfmVLPRysvObecPjuMo06GQomV1
xB1QmxtP/DGlL0Fhxjs5NaWh2TjICdqjuKQOiGWwlEr01kdWpMULUh4Uvif/PbuJuO6PfwBqUIBn
5dgP+01OEPu5oxDAgLG7Ns31X0KFauYKJv2L3L+WmDNhejrgEwTxfm9NgR9OMpvhtXvntyieagai
73tjkPZYmbwtZPyqO16kDu7UkQTIb51/31t+O5oRjH8PiTp9mEpYsvnTa3HR/Hi0VIBOKO7Vl56Y
U+G1Mvw39D55SX/wnOWrjBb0UPHvNu9aqvdXbFfLmyzO1F11pim/2XAJGNkw6bEduyA9D4SjRieh
to3wHVZFQRehM0ZoM2X5NHAd1wEhyP96hvxJHoEfhzJiVULjNMFOvpcsOcYQ/rdKvE/VRBI+w/Vd
3YtZmQamJFyWESgtbnaQk0ElkE923R2JMf4cdcFkaSJETsx00NZNyGrWdtzJuQ3kA1JFS5xgORQp
oebu9zVJV/LrmpSpStlfBbT1rPTSPYeeTNuCW4reSPhxdVHHabiBFGXlJLSZh2O0cGT030p+9unT
CJfmWIjSQ0n/Oxl5qqXG5yqiwDKzZWdOXfxjoI5KRjjgngjCWhuJFdYGdj5TSNRipEwbONzwryzi
TvEitrNVqWJI0A3X4rD1pypSXRtoFOyJvOWo4oj85llqpjrAGkH8kVDK82mYDPj0aAOuk7ZxG9D/
hggvwD2qIOPGLwWXajd8Zng8CW8YXbn6zk9CZXQe7RzpcBAU4Tz4SStpuik+3r2GFMmLgBIxIISF
rZ6SAAJbK0tJru/7EBv2PTU5S1CAXgiJt9Fr6XY8N1G/9M++cZthvZpz58RNYdUGvDlt9MrVSmjQ
tQrkDHxrQmfPS6b45mtsnWbLq9xTcoZVcPImmaiq61Uae4BojXROcT5p4PyvUUI8d+dXhg1G9g+f
BP0uIG4mKj47VP/A43C2PVDmSOLp2+Hl/fHhRU3FFHXQLFXqcVwwtubxOFZuQAHuzjFmuC6AHWU9
F2QY+GvHNd2Z5OsKLi0+qEMlTv8gB5Uo6Atxb40nttC7VQbyHHjFKEVt7Aw0USUQbqzopW9XnMIV
fN0daotlDtF90k2Ysu79LuHbt2Z2i6TxaOjfCQb2JzM/yS+spvBr9c0HsPRKBtuEKiElTxBIbOjJ
ympzkVWwHNMyW3/f8LEg5w/hmjeQVeJ16lm2PsTMNFG6t5ZF5N0+8l6D5EO1WK5tWSToJ27Z4I/T
SkCeTC/ZfFqCQowbNdkSwl7jVEknjlTKsgRf54oLVkJsHP6oC7mbeRJ07zfjRo8TCNB7vAAqeXG2
QPi3L3w4W9cdx3es081u66jHKFD/sLdHpMI5FvGwCoVTAvLotfcXBE3n+7rN58WtefYI0zVWac04
AqktoKM9AKsMMKZc7izQR3afCa9iaAUY08+K+tmwthoCFmZzvAqxlZlhb4TB6rYB9/B8L/mJW60k
Aby0zWupo+QY0GRb3VEqM12gzm2dYfMfCSdqrJJmJyHAat6rj5QAqpbIEwLL7rJ36jWwjhGwlfhL
+7zW9TL1GNRsKkNu9uj/P/S46j/euVn2LQkz6FPwuZGfWB+IQNw+GTBsMYvHVd7E08KseBmiAjz9
c45uRleLVcCAsXy3UKoyBhFCUeI/r8tsbL9Q8o8d1wmb7LFlMcjTjiupBXzb8CrJTeLW46cP6Rqp
MfcCXRjXHHbqLwSKHhjp0jTPgmYwGaWcC/REcfE2wnWG8hB8ogKbbngBSFRK8tBcRVh5xgLe6kgl
Rlr/uq+/ZDuUjaPH0H4e5RMuTX9/DvHOdaNy9x9qHpaUtE2rxaYTHIXlte9ClA9TYSpagDd/8dOZ
mI39S3mAjfE0QnH7zdP8dNtAT8/vEvvSQGwsNLBaVlbzLj0IdF7sNno6KubHiTQbsNoeo3dshUfj
OZiFLKYIYlR6RIroYx16ZC8psNz8XufkHHTtxQNsTEo9uDZCKn9xOwe0WO9O7tbmAaCp3Hmc7ieQ
zyHzp7SLedwrgTbJVcWGqtJ9fFZtDfgagGRieZVaKf210TOoequU4poIpcxmBo8pNzWLo0lNVw6z
VNo+NU4a2N2Ee9YxLRVyuZBz/j8M698h33x28nPMBnhccT8ZvHItFmkNDsCuZ9GJ93OhCuGSCbr1
rRh52SBpHzIu4Yc9MWGmkl4mTizG5j3dvnbgQJpfaz0r/DK2ShBoCTXoZP3XvVJI/8AUbuvqyJKA
BN+Oq46DGpPIvDUeivZkyKTKEBdIk4X9rTwDFUmtGQEWSJzP6Uw6ph3JOZ7vaQeD0borRm1ZDPSx
UyIdIcZhgTwzH5cNAdfjswug8kUxUv9z5YlzbpRp60YhqtUn+ACQ0b1vWj0Pv4hiOWcHgfHqk7aH
eIJDZSE9S2johZLz33cMJtFHmPoZr7iwry9/LxhIU+Q7zEmg3VvlUZZDoKHLRmsIr6y4+8gDb0JN
uCdJjzeqFcZYY7uRyOjW+IBA6kRDJysjS/MkGV1caozAzlENbGdqPr5hx9lzTxmoIJtxrznQEJas
/dBaEYzlah5NtRgDPi7XayubeQNPhkekvyBOP1KKaM44ubzfTa9d95SZ7LOM7Qyr7ypXc/zaLpSJ
fHEHWX4vqc856BOYO2wJfCJM2WVEkuzIQj33XDK83ZwiKq8SWalPdqEANhKUcI/8c+nwuKqaIXQG
gEKqZeCZeMfz+jU7pjNDT/lRHm2yZU4gOhC0kO1FIw9RJekmqJNDkQYP+CIW/1uOxEWI8jR2Ch1u
xPlStVz33KCSuXHRNBYWCrhp7IwqqUVvWXgkOQ7aydVkqAfALkixHhjTxhF1WrVRE2/CggDg3EQA
zZ0HLW5iU/NJVDTS0GO9mLLkTzdkK574ErmD6YIBSx4sha4tbjchKi9De+Bg0slOzkVUr/tddaDP
Rf8A4TBW33B6TuvJ8ufcFHBXMAUMnACKpDN5ObfE7hEW1nYfRYzWB5bBl6giHJ2fbfxBOxibN0AR
cEJHO5E0dBtjINLm+y+a7gW3/S/RCV8W+L8FS6N9cfJbi9XcY4ucx3+RaftXvhU0NUxVSuEcDx8i
96VhWCIfWAQDlAcUjrEcjK8ia6fLMQrrvG0s4CTzU6I2tBIcqMKEeK2DBvxzwS5JaC7coALKLtdo
+rfOpCaBpWaXeEPXD/3frKzVemhf1kOc89OOl3MnaHLbxt3WOBX7atI8ZzuxAdumFWqsnjuXX4Jp
iEIeyQd18jWfW+IWHpd3CyEOc+APMRxjICMWwvKDRZPScL8RMeZTfvbYmsjHo2e7wThlivJ6O8xn
z5ccQW+oS8DpaMRpED9azMiCJhPTsV2/IhKiQc7kpvEv14Fw+Db0uhDzhtbKkER+MT28N9qWfPkj
h/c37NSq1F7KArzK2g6aGHtSTkytEHxQwPy8NVRkBtxV3opsHMNrw7xnv1teEgLy3QhK+I5VnTB8
yxHRlpJslzXRKHRL060/k5qCn5tKbE9+gIMFsBdzX5bMIlXzpnwoEmjgoaIO2JevWG3EhkK+hPAI
k2cpe8YL0RTWiyenc+JyMclC63y2UxN8+q8nrlmNB2XgCbNyIlOF39s1T0bEdOybk5lBLDbj3V/B
Thk8qXOuZWsfySjPz4rmpwOWFmvw8KqU54v+A8+kadPMiQnHcGL/OPtLBCOowSndE8nzJgO5c4ci
yDbsoIFr0AhjLIp06PeX1irawNLuYlIpiRcEGI3VDj2+GGIo2i/rhc3tqH2kz6GoZLzA/3nPu41z
0hGUJGYM8OFZuK6nBahysnk17ww+oBesu83VRru1ZUVAQF6mxk1DnOkktNv4bLfuLHMgwgjT7D/s
jw2nqGRNiZv+htW7HhYxKAF872poeNYUhNbPA7rS7+wbChthExPitPZ5/5Fe1bbsHhEQXaCEM2qD
ajF2jESC9TuETBg4WPMB5+zhQcFpbGlzwo2kk9R//1v9BBpOdnSfWom+AG0LBkHuAPFzaMNSOQ0i
T3hRoZ9jq1o1VIBMTPwdq6NnfHhpjwzLBCXro9eT3tMKenczBjFCHGXE02/lvNRd1uFOySm3DHmm
kg2CexSDhj0MMOJpyBvTAanJvF3q2kVbNFkWAiPLpqReHfFzz8rAgxIdDKJ4/4VHF2paK0GTj/rh
S9mI0UVvFrbOwSNck0wYA3MmBsWLiywUjvCOcqo3Z3MewRyl3YXauEfDeTphVPIqM8lybwMfg8d5
lQ/VvSs4cbENPMoKfxJf9PGcvuD0JAQT+bfZWoZNqRuQ11D0SjNdUPfHRuYwL8usSXk7XX9KumSf
XWvfTy5xAHfQRipXnpnpSlmfll001tRXwwzAWVxiZmjXqY3UGLKhxjgBxiedhQf0P1NOLuhorT1R
Y6iDEjLo85LfFZuPOzRBAq2DoSxvtdvF54Oz9be9dCFLlhChd6xOOVt45pWBntPTeF6APBprVWEb
JODwT+4YDQmLSVLH6YN6avsYM5A6oI+JvrFZJfGawOS79R4gdf8iAaV8zQi6Sw8DePLpDw7wreUe
YfYpWzAD/6Ln/nzICSAcfnHCk3ndqT3s5SsB9g52DfSrY+GX0r8jetnMhCGtl9khlVYuyxRg2V5i
o6f/Lm8ww3ojexSzqIR9bNzErjQz+u27FMiPBFAiDqgNXvtQSe9RDu3OkRUH0yE2kWpWencC/qGV
7dr2ykpAP91P62JDiTtnixZwMSTxGmo+aVWTvJbvHC+uWkI0UNxmjI3FZvm9t/7JXaBtdwioVoZ8
LYp+BujtYN4S0xQM7vOS5iS5V8xwpFwgmgpxyMoxZNmhcU4qmoVZxndoKGuqv4HHD2r0HuU/77jo
AMEFqyD0tJ1O/gWIU6XJw/oSTpl6NRGZrm2+bIsbo3WrXBszS7q/q4zmgdbolYEB0kXpZtkWsZnj
3jv57A8k5yfa5zOsotD6ZTsunrPCdsA/Uk5Hfbr6cXEYAT5c3B/0luzYGpD3O05PPm5237sERJsv
H9HrBSHqrWdO8Es9fUFm/7TIIfHjv0iaTJ03RYFCKCLG4LTB7pAH+J1tMq8+2A7eGBZbDzfDnUUo
ivJNmPj5KQ09O7az+2FiQQNEOF+EGsC1hWtFWneijMrxeQRchlPoAxtO0QdTIV5J0hAHOISd/f61
/FQeJ9aCeK3bYywmaJh+pDyIpMk6bynWt0S5SVxe+mwjyVvxC6tgpDaKLFd+0dFeOJk2UwYIep/6
x85IHeGjg64H4RhU9lpF6Lz1xKLYsF6PaM94H3/QOLIMhnjC/kQmyLNrDXeWxCGu+0z29HlBytrU
uSMKZeRCggRmTgRoCGiOnKdkHJ77JeDNVTCCgnE/80yY1SHbmbrAaRmkmserX6mPtCI3NtY4sndJ
D5UYTWgAEqB0dzh3m9IMXf6tTQOG6wGRxAqQT2nAa6hibriiQixLwHFXeQ2YxZbnA2wuAuNtvr1m
XHNl7AzYOPloJqRKNFGHTJdKdBIyWyD5MI2x+vv4jpLo8NK/xlNu9m7EhBVwpZg7uPteHNcI7O26
xoQuM/TQyxNI1OxVVl22PtJ5OMc3nztHWv9+7UGhxV8HDW9hZwlc/X4XM2DLWU5ZV4ZfUpB4CJE/
AMGT5LZ4Nkdi5uM4Z5juiDuKssnaItLJPJHTtKbPrOa0Jf0+PxPE7jPao0DtO5qgRfVCCWpok9UI
AeYRj/WCibVBBZfcir0MFkUM0ou2+9PkKpMne4muqCfTM2kKK4QmSTV3IMhIOfKGPcJYob0+TM98
NX0/FHjkJtoHamfV1V1IwCIkLDHXJWBekkFJLZ3o6heHK+A/D+vGbBwmRlF0oer6xJiJ9G+UCMpg
ZBsofPMjNTis3KxdR7tXOEOYNAP8R6nHIY4wNrrneiNjkTBKD+a3+yWxvICH2T4PMvT+59aZQbQ3
NVrirjUNMnQ2D1INYnU5tMG0isoKcmsoy41iDiFVl+mpMILey5PD3zyc1oyRDIIX3QJe4XUWTvD3
kZJh8JiCgQtqMkDSUIM67wboeH49dUozMZlL834vXDwgmJh8u5EplwYaciuVRxRNM/7U4fwVVeeW
xkJlyGbKZgXnm+8sLHk/9x5FrlMV8vDoFQFR44ARooMHgNC7ml2nLAiMyFOboLRb6ZFQnohpKGJp
q0esfxUxqB7ILt/t0decFRINu7y1TaWg4wXxFPOhbdsMfaW07ALjQ8ufPD2F85NuhmDO2LfX7e8k
PNPihW6IwXmYZxvuY3qj+PjYV7ic2tO6QHs4EoZ19XUeJQqa6SFvHx6IIycN1Cg3bTYCcmQB9WU3
YMyhLGEzl4Mo7vrMxQNG7NZ64uCeQRrIFlJbA0vkVo8W4LZypsqLUINv+bqI3uzVsH53JoKyjD1n
3kGvP6P/qJ7Xvovc3UQy7bCZQzEDPanhmU6JL/6qBmWbJVbvCbL7IfcvgR9MWG5jqzlItl9DPKMX
6c+L1FUigGJLVY4UMlrtbgnaonvwdkPyXfYmP5ocsLMk4U/QNbQyX2UuT5bl9Enhh5emNxTXPJFR
j3li+ek2iDjtfITfGHBAx8eXxjpbcAzqHwWz60Ox36m1uixqfgQD0g2rDz6lWWCjRNwVSYGc8avr
lqwXsf1t3PT3GE51oHHi2D38b6752zGQ+86mPWlAD3bLKJTD8r/lrZpWyK9TsLeTnD8jkJ1sJ4pG
F/wcQAvmZDyBO75RERbrLwBZDolxjUfcPSJ3CuJ/CMnK9XZZyXo52APm/3AOtVaglcN0Pto7gR03
jeP66vVCMqEuVMAowK68AbBIYx/gu1ChjxdA/4MHpcfihbtgyBoE48dZLMQlA33grgDimqmAUXxe
VkXuCB+ONV5xTZuWyGDVpQVA2t7dXnfdODvs3vjpzkxQeuycDFXGUrDArARAwTzQw0ttOjlNG0G6
a+6Rl0mnv3UpfG7dRSIVfj82hOWQwlTHDQLyPH+uusKszGaKO1aDTImouyi7+z5DGjXaSsSyL8t8
RvTeUEhsXKtR2F82gaqQ42XqzMlCEZr2HULbwplMS7LoTuw683K0WoxwoQj8mFse7iN5mxTqmsWe
Vt4Mpk6miZy9lLjQ40PMwRWHWBHNt3bJ07ANwsy6nxlXl+F2NUaFpc1H/lSvartH9NkZHKaKz9vR
wATFxEqhU1YOzlh5Zb2eAGAMIj3JPn1IGh+g3iUGnNWfiqSJOY8O19vCcWdLYG2x3BFEtqzgLzgC
58OZFoiPYirRGiKvvz+auVmcEptifBIXE6/Z6f81Pn+/j3TSK8WBJgzWTvHai9JYNy/wtt3gfsPR
ou5tt89r1JzMFsHyYl40+acup04Fg2wE9I5jTRwsqZ48Jb5PpIhBWpAWWbATA+NrsRTxqNt2vAx5
x6O0XMnyUahpM7eIQQmaHMLCPV2LVo6IKDIVFkF0K+5Aw+bdXNHcV237846WVkE3jOm/UnfRmQ/x
NKBF1UnjbOD0l9IJY0SoQGE9FlXNu2c7qFU5h+txjZSgQDxJdtLoLceA/sRSFX/e71wZhrjjMNMP
ZRPY9fD9qgM6h2uPf85G5cmj0ZT5xpF6gG21NI7Jdv/j2cNkQEjWO5dkuzXBmtvopOz3RGAIVGtE
V1UBSBh/t9pjKx6lyfXOZ2Kg7E5gqnFcs71C/jIagvxnrJtMqvcWmT86QYAYGOlPXHB575JDZKQi
4eyViBTnb907GuBQ/gs3DHNRN01BCPXQazt2xFXJk5CBqRJ3wjqA8L6SE3UTFenpY4IDs6ystlaL
ah1FFomgnFFJOiWdSev1eR4ZgN6eTc0687ER12sdp1GHESq6RJjjLS8aHRWFd/nb5Pv0tCN9E7XF
r+ALO3ILYUR3yuFgevyaX1llNs58Jjq/yluVE4vui64UFvBEz5LUXEefY5fZTdkInO/SpQCsLghE
R5TnhEuEk4+As9BUC8beviZqloG2Is3JeQZndbuykno5H0X6BjNlr0vZ8G8IVhD4r1+nbeTIMtjp
5tXzYlMGrNVsCz7mAr2Mm05gUsv6zkER74VEwYsYZnknyavoLtx/lslP3zz7oCeBmacUTUSM4WZB
7b4S953vKQ767ro5DEh/3Vew6N1Vv9jlt1hgNXeCi2162giYyaQvEJlAfjQVDp7+2QskitGf2SF2
lelP108VcYg+ytcfnmK1+UYB5xyoJD1wSsPpZu5THotX0AtqpS4aqyVPc+UwStZi4Er8xnTffhtm
fX/5goHhHJDupfKLGX5wwUkXr/I1/w8q2FTRXB4MzIeDegFOaTIVGuTecAiiHCbAAz1Uj4kT1DLe
/hPb5MygEuKP+ozPpt+rVw+OkU+hlZoOtw5uOzKAjy/P4CzWfxvD7hSYcthWfIZ+r190me7+uepq
S0l+3Jv26sJTyKcg3dozI4u+bmJoIvJhdXBZzoM38JKfuG147uNf6ezlri1SSBQev4aGNa843f5P
OY/k+/hSBtakZZLXywGOYiiwLMbOV8wTSqpHM23D/8EvbATcd7JkupagxEkwaRKNYLZUPrx3zrYC
iEUp2gDqGOEOAnv4DMbNOMeTfi6b2YmDbU3Fe1XJ489Abx6Ojzks8nPcO14fBCyWCpVKW4nByK+w
0rTQSge7L/jb1RaAkpAaTl3ZgF58+jaQd3PEmi3bdc/AN3AQNBprYY8ToWDp4vYoA4Vi1c8RbWEv
cGTTywlT9Qp2NfUcFP8iyIJzj/FgpIRoz1HhJbG/Uao8FSVacPUVaQhbjSRve54xQdG1uQon8sZ0
M1/JpQr57RdHvcp/Srp9bUxAK+IOsQc6QI6M0oruAX7xtnsvwWVWNW0xoTSqypeJLQgOuaXhtx8a
LNttjaA9JeIgesU4so/PpEYbp5WOrWT10FQle0ok02Efr0o8S4mC1cT0NLPG2aK+v4149KxLIYZC
YPxEWZIuWx2Oxz8H81evJmFdLu+dLBLuKfl3LY3wwK2Z8iZ0L4Uo7N6JRhyBXJdB8Cw4b3CrdtGo
DS4d+we77RcmCY2ZBz1v3k1tpbHMx7uEPSLLHwAEc/UmYfYYkNbArRtzNzB+7uVYjUGkCDchoVTk
JGHEA1yzWZtqvuRLYm0eryguR6t5sdFOyMHHESgs0WWWv+Op9Chd1CZozFjWkhb4+J3wBGuOywTJ
Fcvd4DWE92Wf/F6yH7nfPmY/p710Qb639jp0RoAhvN4BbiKperoEAcljdke4c3SoPDlUSMOCQmQt
iZKvGkpGcqiQXwcxeQJkhCTN8NhSHcDiEYQqD1KDMWI735CoguxJD29stYOalXfDHDmUaI4u6zz8
hROZIoT5RsfR35H29OBtCszCKZ+VfLKE1Yii8Lgjo0WgcGkmqRT7AC8wT4wOCau7YelXcIMRZLsx
OEt0YV9RWOQFeDtHmQhkB4FS7cIvwucLW7RiCHdpura9yJla/cpL6526RkHamvv6Mgy+oaGWI7Qq
V6xJZDQc44x9QhRv6UFaSDxSLz5zg0t+KnvVM0o8DPhRVTkbB0BIC0xqOgkxPRKOxu9NCHzoR2Ml
nc36RGhb88UtevXrCpKie76qabkvbS/AGlvEU/PE/W2cXfucNNn6Q7ravv4ZDvEqQeQ5Jm92THUK
u61I28cakP4SnxS1aIuPIs+OtdSHRvj/h3H5ajPGB/iakC4LlNWmNrd9KyJ6d7cqYYaUfI/l+8JN
DkJOan8u/kl6S1ZLhP6TzGTHXhaxXd+4CttoZUDitsym3xsNqg+qTSBih20Jo78hvUVEVPL8OrcM
nSoqKqNI24mCfF74m6ub2eL+2/LNmg7oBEAwCZxkL/5w5gS0iA8F6tyNtQ4Sviv+mSird7y5pLj8
txpq7apcxvS1KHm4ddUNg0gG8ONQpWntKDQAEoRmD4AQXWMRf/9O3QzUioZrwWhxuh4rFwMp+fgk
EKO8AagcpC7OBVwWWDtyUUQM2ZEAMtglwyeD4eTCevzIIa8sGZGAT76+zKfYxeevpyo24hCOKLLA
D4zMzOjrf0+rOrqQ/6vA69+18nrYupLaAxJGRBbuWEoWd8F/F1ina9NPraoCvRl9pZ/zPLS4Hm5k
jrLHqjTfzYqoZoV2cwIPxFpHWRYdt+FXqecXAT9/Uj5Eiz30FdjIlys1gi4hF9/R1pH3p/867Oq2
/v7xrDsGqvJGlEWmoILTKza5ekUkbpMoGVR+HDjkcieyo6qhfWxYZhk+5G7evidgX76AI5U8pW72
QMGa5H+Y+f5PpYyJH74vDkZ0j54HAfrq9cfs8qx7UuUchT8fK28FiMUztMSZCEmNOvaCZKg9PDfi
teQPJ6LDuxlnO2P14s0BpKYWBaS/vrkncSat8lQ6WFKt3QwRGhSH0GR62AcuQelVvdvCMUXN8iLv
FU9lvvxR9PZw16xUO3SII0bBhviXqbs1h9jgJ7VMY99l4UuyiBck85Uf570VASkIgvqpWLQQr14E
WjkeutFRhMHzOtyh+Q0uRAPKfLlqivdCHeG8HNU7HL9Y7tsCfkHLhhThDvuXTE+dYgUpw60rZWRk
K2XJxoMOuYDKUjAV1wzY+I01cVPnP9O2N9vJ/+2KZ4QJscjo2inJrq6RNw5MfXbt75Qd7Nsq/SkU
3rZaxgj+BDWkLH8EvUjcKzON9s9cbHJQIYvyWo6qyBiCeKtlIWFA+Okz2m2kumYlskE1lOyY+Fth
NQ/GigYOyawont/XeUVptad2ejpCQVxvhmy+ZsaslzjwoGyoJK9oJWQrWgsO+90erhXZxjggPIul
eIxhF6fxaY9isUZkTecENycX+nw6nTjnhoPUxEWhYLtI0NGBE8zd75CQ8/QOATZ5gDCQjnBlViqy
vHgvYyFygeenCxvYh6LC4WMCKGvcNQC0zxLanorRssy2ARWYsph5NPUGgoC0AFBpy9Tt36GHihJS
EitVYkXN1CRTXClvdB0X2bdxZ3TGPX7TZ8HCs0K/tLSfnV0Rmm2hmcsx84tIUPA2rCBBzbcKU9gm
f6P8rcqXrTFCFNqJIZdVt9BAjz1w99FYc/PFqwLXxna1p7VpsNHdbs71eg0XGqjhkboY/y3lyMY4
W6/aEaSQqDRvhM5mTyaHf4iDZTnfIJcmFhWQf10fxcSMdkN0x6qjeMjkj88sfXvR2/T7UdUbZlYH
RfDflhVEpiap8jdjbJPbYycR4x/TpGvxSuMTlTnWplWI91hTX1ikL23wk/4jm7xTRITPZY4fuTeR
nrRrbVU6tN0VLoIWooflom3SNVIFOUxxpkrbR9BI6iIJYbL5Rj9yEsOv0o7wSN9nJRZFyo5Rkavp
HjSsmLRuvjSWGTCd9eAV9xB1m9yFQ2JBBqIvUnZwz2nE/ChDMSGnxC24W9BfIsv61evFWAUOuaXV
tMizW2UJbSeaaKO7+F7ay2BziOjRrXeCYtwanC4MXYIuIdERZOAPloQbsSw/cw0/vPbImULNRErc
6Wp17kBJeC+Vh88ZUX6fqdM00Vscg6ygkEQIJfr9Biq7yHlKxRaQWotDcf1h3Icg9P6wVs8LUHpK
AB5/OA6v8tbnsTJsfoF00QFM6BjxtWlTghIUcW8ScSquoDQYebKhJCQ0G6f8Caz9AyH7goOCwV69
8pumtuNwDes9tB37dGiJ2dcIQXk99xozes2ENHxujNMOARy+vFncf5SuR+YQ4K0xx2YvQ5dmXs5f
5USTYFPMSMstYmnKC/EE6FCd5T2kgfQjDqQSpFfeKTLWIrSln7jGsfhKGyopnHSMZP55LPsMfozm
x+1Im90Av3DLT04eWJPjivnaZ7umLngUFlNfzpY4F999X48jfBv9SDIq+zzuaXqgNG/IPq612xzn
hneBmOJWOGey783LLKg41AA2644uGmr1JM8KMGK5DlveedVKAskOKd0YveLbXxrH9fFRM8CSNWwE
5K3j281mR06FCJfGZwNIxHTCY+5W1VQuEjqYu7mlyWfpG0THsFKk7va4+ix7QJOVTdf+dIZ1kiE1
VQxYFAIUSovdpyC8bISRbckIRlPx+O/akqqBk1bJTwFBFSQSdZoOzQfpBobrxL/GdcgkkctmtbvB
Cs41DAvM3YDQUMeK8MJg5DdgK985qgpsgY/N0cBbrzkhyQYJZ0FBjnCfpr/wlojf3vuuVaSAvctW
XLrUXopkTS89/oEVTK6uuCBpUFzcpJos/BwQGym1lGjmZP26bHpzU5hDF1MeqLZTsdeWfcEQgfES
RCiDAymXiSyw8ay2gEgZjhLbZEiQ4S8wVBefPB8vM3vNYbKHJs5VmbXnWtzHjTUggQ0zHOxOc8Ln
nHD9BFR9V0q2p0ypfOLhlVlKZfO2+/jMoTyvUPmkfLVXvsFGaUc5RdpRSNKEmgwmtt+trA4+amwF
Wm45oueaPeDSTIpdNFzM5PwysI4nanDc1snaD16oZFIXbAiem7kztpfYZu7TvLrMJCFrsllcDszR
APDkABqR5/uUKXRmmUbgpDOSX7KemW1UKREQUhzLmL5/Z1KDdS7NP73BWQkDFjtJu+IdoPT5jIvE
mrqdwV5105k4S4Gw/zVdJJpJt/3F82fpZToDxeno+bkZ36W4AxXFR+GV7CL02CQ6cQqbd/S5trJt
0Q1Gx7TAHstjv4JvGuKBT3rMv2aBOus66YSByeJJiejZtaCUcKFDnG+IQuM8qjYwkiXVoFCxvlk+
v1/BGtpjIreLNZWRgJDOt2Ji81fpsjEJnSygyeJ1x99RMauR9DJ+j8rwlEoxapJuP4I/l5SB5e0i
mmt3JG5U7apX9Jo9n6vjLUrL3sw6Tt7CffYK21zx6hiyICoAK8Fg2+UApKQGcIa2uwKQxRvCvhTZ
r/Et+wj754sewTAb4yFmcEuTzRzZhbxCjIM8+gEm2NOzd/em1/SswjxXNqUq4n7ycoxqx1MoN0+h
caflLLCl+64BwVLiCS2qrMDp/t2LexQGkP2natPcW0+/R7AS7cmXmwSPoNY7myujBy9FvWnrR9Gq
jFIuzG5YfhWTHYCSvco5/UJZkCGGYdxRLorL9eGazdeI1vWOzDyw/N/RaHFuGO6VzyW3Mhxi1Ds0
pUgTjC46FV+SGRguBRUwAz9gnVVIdrghP1JYTSbl5s4zOBgr3sVcCK13kmPeM4c3kJ8GDml+E6ut
tzSkGMbkWKC8aTgUEWip81rOOOh24fHdBZ2w7ONRiG7q5fL5w19Qlj/PvgNZ2YFY7u7JdV1ztRx/
tu6h6lL/L3wiFjTpQM5WKNw2vc4Oc438c4mirblVn5vV7ercnWPkNTFzLoSK1J4X9jnnRn2e58bt
neZ5Tsyx78H6nn7fEps1nCsumiFTXICwVR5URFUsTuVxxepI0P8P+ffVKU15GiqcXHYyFECivci3
XmCLKOvnXCtY/AND5u7DZarKJkcuazEfHjtcQR6ROO8AiMrZW8hM/qRbudHI374w1icb1efjAblY
EqapjR6igGg7ful6dB3dwadcD/0BB6absJ0t64ZfpEXuwbEODFsUb2hJZEaZaT+nRuTbkCJlXPTj
lVS33GIw7buB3vX0VHTO1iEu/pMZ/YzZuxCUiyzsAKvNI1LDTsDi110R07/uYci1DX8MA3PdrtVT
+Tt+BkZE61JhCb2igY5QWIiESLHkD/TBM14iLfDw9DSYUir1+BM4Hw/eONWdZi75GeOEawh74G0R
mSKuTvBLeaQa6XyHS2tv6paC97OnJwzdOORPoFNt/gFsCCNBA3c0pymTNzLZrO7N6iyKdTDWomF6
ARLxCEvajjfYEVRV8dbFvaRQ6FrEp7NAoD/78rLXuQMAauEUlIUrfC8Kq35emQ+0sZm017IpniU6
BTRMaP3jt2QF1d3c3W7q/Ro0kF/VQ1OOuRbtGCQOIHc/4ZjhszAF0q7oUAP/3z1QEy0M2SVVByIe
Q5ITqz1Qz/yQJ9uf8ZKhVxjMHSC877HC0P3swKL/RT0f8nhP/fELiRA0dtux8woNLEqDqLTBSFSJ
IDMkgwBrSxQvTPHXj7m4MAD0UaOVYVIQgxZwjb2/RJzFANExlSRq6sBciBdjfeCUpduZNXqKmkxQ
59uK2NMmR6et7TnjiuzwQx0HIONCPl+T1UPe87Lj02Oj/HuA8jSaDIikCmJCyHlXjT53PNZGGiYB
7psUbZ4iEethfyf9QTtjT4nd/kWsr4cKKk/LF1101rsLGFOreIM0JfaM4upynXLdFei8DNxKHKrr
zJt4IwvJEaoofxYgMbLZKJe739GDjh5l5J2CCtlINy09jdXlb+Nen1YaWay0i3g1KcPCBYXSsSJv
fnuXhXakKAZLP1wvGtBlosgM7a592cuczxzygOjhiSN932+zkDkVDCzQNcJeg5Lo8L3tglmS6r8K
/mgdAiTmrAeBoaY9rAk/9B5sIZKdoFv8qroJ+rVdtKRx2W6C5I0ZApChKXF8F1Lbe2SdcacQNj1A
kx/vO3CVZRsz4ITxI4YCqEmtNgwHYLjii2fUHv7G6CN6VMN6GFJh68aq7kyspHthQatbs76gxpR1
A+31h5i3c7NaHVOKAlDhcnQe58Ty1i/Ry8pejylYNz0a9nsHxYn0icfeT86wNP6VVcxJfYxk1puk
Kn6EyZlCJEFRmqpqXUWXK0SitiG0PrG+Mb/lC8rFdJZSer2AGBpePiTAmRHoWHSkgmCQd/PkSW1e
KzLsFviPiO92Z/9Nku2Eh6gYZbBiJlxanphbkBU0dq/SIDFE8vNv/0fxLcnVCXhgdj52DcfF5/Ak
7JV4TI0ZutoV4wf23fp1+KWAxXxefEPvxd8UvM2ULQ3mAVjeTrbuzXOqisw6KqDIu5J5TwLL1tmc
J+rZolUqgDbJ0aqJ/DjjEUQcDQ7eloR314v/IbAz56RHb4dtKpVBtTb6DaDEvTxndtqVxWo7OxNX
5TWgtMo0ER9fvaiXrBvYkPkhjmR65a2LeIEqmCqiy9DeXLFQcn6MnRjGLarOXN5nCDEoDQzbGfD+
BNaoccsP0JaDyemoeo6zoWUaLcngy059tzjMb3tZb1wb7Z3avSVCLkFt5ndcCDxRDX0NyBRPwB9E
RoEEsYL0qCQ1nHq5uqIi/BkFW63h+1y8tJfFWGJydySjqGTjC0RnxU6faDRdcO9UfZpzX6aYgBPF
02Dlp0PqZ/12+bLfULeksVJYbEm8EbjNlhfXNDwsJpIccxhUwWH2vHNsl0CJU2ZcARk4mUX4raaq
V/IxqTC6tRLawE9wO+KtJkZjwt0Pv8BoNzAlK6tZJTqxzrm7MQm0iup4lg2eX03GEKepThfqCZPo
k//sNUyjAleMFPNhhc9AWrXJ+igMRmoE8D4l66t6vVT55P8T5B2KBzitoGWve+70CnSaqYyD7zXk
eSiTIQufD3VxQcK74K2CRpkNSAV704hAWGyf/APOblRlvxIZeo6FyXwLAB4QR5IVlqQhfHZV3HzT
fH+329cq1r9pH7zfaazNbTBlewowE3Gsf8BKyue8d5BnoBklbutq69JIswZqTaO6zPlkzS24+f06
ip1nZakNY1rC1qAQSdby+fvU1v5Pc0EEdE6v6GI8Ex0EpZnfSTMZ3967IEHKJoALHmIwNXllRY6j
RHYMlPVaRn0ZvmGQ7nKOEGo7hrj+yn3jc77UiWFZIksEm67GO8HRsrqhEaFooL9x/oUz5tV8hWnH
8AaItyxrnDH+d041Q68vzeQYt0OU04p/RZ2VyzTbVtM0wefjM/fUi59PXhaqwgr6w2vzJLxWetPw
NWCR/GWo6PrFa4MgeJlsV4YNKQzyE6yxg++v0+aTUZiIunRW92OtQEqzcH+UEHHOuDSzQbMfXqUO
TncVk2IL9ky/7HW6DsrKB+PU/OsYsQoEPSb3ac9FBVRJFPrr6U2MyYbWMX8Szsf3WGgjwoVR16Nt
dJB540ltXtCIgx76OMygkHIgihqtUnZtEHDcd58rzEpH1pDObk6cWfFYSl242spalkrlIGQ3McNw
AvfOqmsjSYrcB1/1t3mBu54FLLsGXqxrA9TEnU/wurytL3Fy5VEYPwk3lpjfGgrGOsNAfFX1v5ko
Gltfjj0BbLfNFZ8GJtDCZzIgb/fmN0cspnHjfhCrXU2L/wnKn2IDyAHuQ0TahIEQk74zF2rCDNwD
2NL/HTf6VB9YoPA0wUjGGgft6gSm0HOyRyZHfXMye6cl+3EF0u5rUC8U2geWGCYreHVlr9AZZqLx
SK7mtD6WSFHYQWAYImdxy9CLS55HobLJp/YeKhuy/b8NT8c8Ir31HiDHhBntn2w88EnitNFGvXFZ
wDlN8OhZmnnhS7sfBO+mssxY2b3esIN2YPgtgirthxODMr71PAlqw2PQqvMp50N02WLxkULEdZWv
7Kw+ayodlvTDAuQrGWo/wz9b7e7yEGAza212q2YW1ZrvDbtGbXiSIK9Tlw+ocR649ymPbhMfMFyN
qbYOHM3lijWj1NCBnanuoHHZBQX7zYbNwIG0xD/9xQkXk7+ZUhVWMktcFGH6hEgQ7sQWerkopJif
KMRrmvx+HmrggDhFpwqyUtwAgzchwfjGdfH7uk9heID9UdvCOD7ZSdUeZN9ftiMj1MRkJdmO5yQr
yfH5nQoK7LP/wu23ORXLtUqfDWNybxMa0uapOIeq9tDtr49q7JpzSvvqdm0myoRGZWuENczcfb8B
/JYqB1y6keHl7tOsjlPXR5heCgKoFgCnV3Wdvil80UbyfUb5XNVf1lTDEqw3hxsjP+f5kBXOj1Sp
bcYs0T3TRFyFOSh4GyM+THCq7VxnEVqwDMQfEVWIBJZHULAe7gJNBFvKCbN3/xL28Jw+S0t80Qhz
9B8/JD+wYWLZmgJpRQ9kqW8p+4lBcyzDwIb961zdjk5QsSreYjzAfni/w6Nd3+AgTzp2pjeYAIie
TwLAaGjE/X1eusZBnA9kk9eMDo04odqCnXPbr/QvqBM8vcyMG4qdmjUZkHTSostb/PMqsMPnvY9U
69wsckQu0mXppm2zSyXX0461wfo6TLMniRi05+e3PAQ7dhvFTvlYLqGZCUGOGxCvyA4E/yufiC3j
mYuos2vsswMJ9fPCAMkbqrd0htyG86fku0KMxdnHIxKeoSxyNiw15+ppSfPq+ct30P95TdNa3jvS
jOAvcTWDHPl3kOtpE5p74i7d8Sow/65gVgvviIbi+lsaYsSmC4Q6JK3gPkEKTzsXe4MLNz3wgenc
h2gz0GuD47+pCQ1lmX1/SZAeIfm1IOpszpB1lB2VolDoq+OPEQdv9PGt8AdXhp1hkWiOdnCTpoOn
5mHyqwAa2b13dN87FFp0TXycI51GNwLouoMC/s2hICtgvw2iBuVrHXso/wUmiuXg12cZqhOld1bp
FRcGC2FXWJ9MgYwflNN7cqwz079pXMfUIfhFHhu2rzVgFKzz+eQjrPvEjShf4KL6U9CIvBC+gaJc
sO/FhubJEI8muLGIx9M2s7ueG7yT6RWjuj/7VdlJIe0Q2W5/A698L3X67mnWAUR97bYMGyWIuYiL
4Uc5gSA3KnqeeSsGZvJ0JBCdF7LvpJSyWfWTeiyD0SFqPfhIIW8WEkdie2TWQ8GqtWO6qX3w2Wwm
ZkwyQgRkRyzaXcQLEWZNe1tUcozpioaZSZxvsmWJeXJTi0q2TGPESZ2au9zo2Kzn7NZpQxkxetFj
XGyxuy6HYu3VoTZ99VGPHRuQPff/uxoWsqLkNSlXgXHC0HBGpOZq5ZWilKW6kcxRrTttaVTUVZjZ
aZnPPcbzm3ZpDb5CO7K1mCSA0EMnkQse7uB/6FPMIFbyXqp0hXhZdzcrQLScJNDFlt8qfXDftspE
4DGANm9i76JK8ajgxs2sX3JRDZrjy3NkUwcAMU1935YiuypmpohaGlcxdBr2uRzzmOJQ81vY25J9
kz2TxJsol4FIzIMGFBsboXyT5xNBsdvRx0Pn3roqOAKBZeiesFjfXqEjCWpCfu99yt8mHTDvtESB
QAp6ETPdL1p1/0T9A/2e28zsL43mzIbPjhLyiVDVq0gSGDJKnJ8qYX3M/mbODWclERLM+ZEvQgll
nS5yu/+cgCjeEB8uhOSWfTMWxwvBfTcm3+8DQEvBYmo6IYAveNcyM3b0jjvDTWpUEFRjmppN/Gbf
jhfjFzK01CZh6GmKyVlQgGibHyMI9JMpeKK+PfIkGmrJ57qGgRWOaU1ZjBtAeGXpdnRD6H55A6ZY
b8Z1CA3TmPVJmDpqDSCA+G+53sZwzQZlr4cuoWXbcOnUeA4uYWBuEmI49DDDqPxjgT6ZzKnQJOAy
8kLDDdTK8hjevdw6jFUWPuVHCjY9m6JL3l6nGmptuND49ay8kZbPLB1d9dqTlskH7kTvk31tc0pU
1zUIX02nhpzMq+WfSXwPfCyAOpckHNbI0Tm3naXQtXYyKm3TsC5KLqYnVmI7xdrJDiKun6k0NHiO
RF1Ka6R/FR7e5jy7XabsPmnXjs0XBzBTdWcqQ6GyGDOH+mEBv41/EyFTt4AL5kiUnOhFn0fJL/Lg
1ydUw/NqiSJA9jHdomE3i4O0qR1Y0dFaSYGRNVbWKP1llMmIBnQ7OPmWD6PM4B1KGx2TVJa5UDpt
qKu5Bjp+w7BhtRTqtBx5ov9Q/dRbqPnLq96qJnCfmdLZABMg/Wnv8iAm+kux4ule8L+durpZqRXC
jjll7zorFnppPvxT7t/6pQiiPJjg75TesGHO75f+XI3VeqjFHoUuuf4Z/nyWE5RGdf9VvTeVd4vU
C2suQqn5G3/2gR7YN9S2yroh+EQGfw/cXnjd/xdZy3VmMwamvspulL2f7Hy5l3zhl5hgb9Ky8KNy
exOUooqsgD4ycIhLpZp/lRwGEoiN+k03tXYRjX69BEi0/tfIDTzD7MyNBB39qiV1ebgp42db96n6
ApL9OVHgQdUw8peRBqCHkfe0o6hUoL/HEbJs6N5WYw9aaDybQQAdKCiLHPtzcQFvfifxVGMyJvsC
Uv4CNAa52Y/JH/o+iFdUQ1FJiJVj+Ruz6c4lp0VgDmOplPyxhTNc7UqsLtCbW4/LjsfFT52pzw0r
dbqvTvX8gOQaFNMMof7o/XTxDJuGfHbbfPThKIPFJzwyMn/zrjU+h8hlwWnIQQljKIrfeLQbBG0O
zmvqJu8w2KFlDeH0/n5WXqqJtYqiweskA1YOot/5SdXaeB/IZg6PNRyNriAMDTo7IVCfm48u4i5Z
fzCuETFaoxIpB+udi7wl2jUeK9POqFtYqqmjfYOHr/ug818JFsDIJOQqZeAtCf2wEsMmNbjTT7HV
TGB2DJwdbCI1ouDk7qODEOXPjC/mVu23k+EWOPP34VadIfiLqyfB/lKW5dVhoTM7BTPKCZqPsBvg
eA4euj039E6X3/4T/O9nZjkrdHPOLyVAv8DFgLkWcvH/L8ixwE+Jw0I6C3wHZnFfLNoIDfD0MyX8
kvKpV7c8iSGmqX1c37EUid1PZytk1q6uN3zyaRxNTiz1McbVTiVziZR31SCOA6BOn0K64xo3jIvz
MDPDGrNnZ0k0xZxFLCI1pWCj30FLA5ebe9EOoTtyw6NOxip3zCafImGG1Vj7bh6CrxyszlFNQKWi
Ix6T6w9KQM2L7XBdQyzBUJM9VxwVy8E1tT5rBk1dLFMQ/PbLBVG+88+uYgIg7phm2+GMcLMShXed
ywokbnU30mm5EWUi8b9qxEGQf0x/TdIqFMj2xrotssLNaUJFZBNTlEwilpooLefwZMivkDGfGrZm
PkhLwAMPJjj0ieo3g2l8oB3KTClDT0Tusn+2owi/fTqAJwgepXTiqH3v0EsHThfXxGvH7uiNvr2W
Kz4mklDviFw2FffgH6YpAw/AK3BthP7buJORl+70EecF7rCUQORbqyXCblavvERZaPw3+QQXpyM+
j0efz5BwFyDmuV+968Xhgvg3piB4+iGMiusIxvwDzJxiFhqtG8oURIC/R0cb8sLzRJ1Puh4yiMw9
3rkEvZsFAMprGr+CXCUSxzwyAb+16l5Tsnl8TS6ZMyN/XsF9MjPym5J47uaa0TgKxoPUt24vO6ki
lYQqdorSqkRJzUCnLNM7yOurQRaJz7qz9eGM2NsB8jAV8V2YtL9SNbmAt3GahFZ7BI4d6wiY0WEa
jgViPjHLvxaFUxdVql0kkdyiE0R88WJ/Wo6oyO7/AqMc+ankvyb5tc16OkzLJ/nAm/MDWgy9OYD7
Mw/Of+R36Uil9rh1aOHecJ3yWlnY+M3XFXBMTXT7KD5p/dBCBBcsPSyxgao7viCmtpIfpOIFMOVJ
4UbFpmINvw0+sq/hVCyk7UdT/K1AOBMd6F90sDcqEvhFklmRCUU0mBRiV9QYfMklQG7zJs0gUBJF
HWp3weRea2xEb67mTDqNqH+F16prgfECx/52GqIFVBCCVfRaV3hVAfw3QK4cW329CMQmyO+0W+3V
DV9YJ475XKdzBJ7PHmr1tAzDEOnsLgKTIR5rTEtYPmaQ0F/Q25vnKBysv3xblsocspjAp3cILV1O
qQZj5veqBZbWgP5fLxAGWNLlYEmlK0qhdNLiOM97RJnecPk0i26KbrgMIR+HGzN3y40qAm8dQTfO
YpCHvnkd1Xjp8lIl94UMM8RtaQjQgCQnQJPFMqWpFAgAQ7UkIO6+daY6+uWipWh2SN/EFU2eLVBt
iG7f64UaAgNDGHOj6YtmMmf0fuoAnhi9M8tDC5vRz576trsFe+5wDAxoKwFb7ZFR6bPkztJHXK3B
38YK/u//6T+gNNdDAdjT+Dw3T7UJNEpQtOHG/5PwztCz544xnesVuBjeOfcytblZty8Pa584zTwY
awZezHI4mO8D3LQ7IgxHtFXFmUTppQAErN/tvGF04lKISVBQhJ0t6XCjOOQ6wuadwjXsFqmuDS29
7Bo4L06QxtFGy7N3mEmBL11wSlu493BrJkLnQWHKbEYNNRmTspUCu+MEYfW0xotBKwNqtZGmpQYM
LlyRQUcinBbMkgMJ7dsLS7ZcOOQu7TXygIg1/aYAwkJ1g0/HjANunk0Jky5d7+iQAyfrlc5ZaSOK
le8v8535HOEDFFQ/57qfBoaJETHu83XJPd2e9Iyieen7wITdm7HePQyveWmeTRRvP1Gq/ViEMIHp
KXuwIC0hRA9SL5j4r5bLzQ0dmq6B6s2ccg6yOzUNW6hGwhaXYRSdHAgnJCBfl302Qt+Aw8GDKgU3
BP8ZghFgg/JnpLNGtDusRRP4TK3tLGVUvY28oFRP4NcdKmM82U5L1S8TVWIzYEINOlWROYNiigFW
SXtbI0GYvyk1jhEadX7bDcStNNvco0NSoe22q9MyhChvmE4kS0WHhvL5FaYPapPXUVJj8TuzqaXk
A+FqP17Iuw+Sj3Ef9wpT4sgukMgyKJ2gI7gr2NsciZ/7aLKmxbtCSKxnofLWT4RzmtWmEGtBOCox
vhUIj/9Fb6qLklT+3hKu0Q+DJBTJdWRsFu4Y7INg3stlitETdnJWudK3GVcJBsfYA9Y1shOi2rUf
xMyQmt76DF1qFPTjgUlufM7o7SoCVoDvAbDGgzyco9NftkPoFkoh8EbOwjt1qVz5v7/LXpo+F8U3
9yaMQVkJsY2jMFlVKjWGuagVSQ3NpexIcw3DjOCtZ/KMRsF/YKdquTTMhffs8iWn7o4zYoW8kaca
Mc0IROti08j3xD1Z8Ti/j3WFH5GjmVX6uGETItzvFixQIRH6R5mItlQsKQ/tL6vMK8GXV5bRwH7u
rFCmWNTVygpk0y2lTByi08oQeLGvuB+fd5s7LjGcns2lN6JHjmz/ixJqesgc2KOzWWNyapMmGXXu
N+nEn3DrxtNfrEHY5LaTvUaxNZb/xm0Wef0MKhQV4T3KrIHQR9ZTvnhPR/nAhTzVwNtxfCy2P0ij
J5gMYWf9ye1Y1n8ZEvDBcSZIP5D0pfUPpJcsHGXICNxfmIJfCIch6792QgPGiSbPaa0Qu9gzM1+t
nkpLDrVnWt5Mq+A1jV7wkKxZ+zQAf6D+ZthtBIe8Vzl/DqPWRU6OtG/XPb/SWCmUe2YWP0Pki5l6
EujSAIHEHALtC1JNlZVS5DE//yu4mQmsorQcT10Imr5N6DeYC/pl4KF0eKFWV9zZY/vwBLUhqrAk
uhw3I9RV1VNoh1NZ0Dsfp3k346ADQJqanvcddqWqEgi6Wtqp9b3RgeSHGWS515wRwjsy4dcmhVX9
wKWpj1JOLXJP3MLvxODqNnNAE/kf/9wFtDaYXxIvWneN1bd+bPoR2RNFficBcfSkaLZ3K8H5FQdG
k1qPMjTKGWi5CJXGkPC6qn2gu/QWd3iEDnpK9gXifNXy6mAkUQ527bjguUi9g0GHt05mv6A5BaTk
qxnW2SiSPt7Gp3nV0jx2YjkzIqB7UX6hqOdTJ7oQD1f/Guvu9AkQmzQHTi3PtkSL4L2Sz+aISFwO
ZIDnO5ipXV+lBzzMCMBcA5YJc0u4+iS+Lsq1JTRTkq43jLNKMlYMAzS+V5VOSPaq3siNmu0B6vjU
4swN2JFJFTmoqI5XWcXaFYmKLVlK0vnkWN07KYCl3aPfmMeqfk5N19CmVavXAw0YIrnvTZJxY/pw
9wfBFGgBy94gQHliYamxTlBzPox55PY682M8idQawNsPLvP2rYrtcmqdLiAL6NBIlPYa4C+9JGU3
pXq8ChrYz8Sws7lgxfHjcHuiqZVTrq9JGno1oOzZBkzmMO+nmk2bQ0KmVRrV6m0n1wldh3pb80+D
J1GsqAfGrt8iuyGZIRD2IizQAgCn7adTitUdiQnyBnLL7W3TM5TYofLebtDjxKQzKfsc1NVkbz0C
apZtVIjpj1uhUMTaY0DDTFdAMAoJ4EwB0D+UZNvqQN9mx6raYRsaSBFFj+i+zTLLfRwVWGiQ215D
zugyQs/Wb8Xkbx6HFjl5n5ZzQiWnZujnuKQIZpYeJYJdzbfDWz7ZYSgpdgDM6ZTrIhzynHxHa7zR
GemRevw9eeX8QJN3/fQeAIUleuFjTBHF92ZEVB3ZH9LDztWa0BL1Gqbca+wuaGHBLv79A8kc1kr4
YJWeQuOD8qBMMi00xfyv/vbYlY5YJm28CLU3r+a7Y5KTGbrsdHUwQqWNkiarUfXQif2hFUxNIaqm
7C8JzyPX1wIkaFqx8G+MZi0uNQGwAubLiG9U7g1MFBz0jFKSlU9hFaE0rQ/UNDz8SIZXCYxElZqb
DdAt2FShtih8r7r8qd3yrVBl53FmrHY2tofJNOt2GQV5477n1bcdtORFbHFzMzZRzgBi+AFO5BSU
BRJOk6C2I5yH9gM6kpqZ+bXUZwyDRHEdc7XlP0p42lZRKD1OohhAPbSA5NIBY/GUHVUWjZyLU8qD
5u4aEFYBDFutSbHwEbsO1QXvQ34z2PeYfXABw6hAOFbm8o2M53CDDzcBYElkQSgff+vSFmpgRnDn
0qaJuZQ/7167kup/yEKnsFsXC/rHZonEZhfTz+wpap65XnQ46+dhUkuOy2anpNCiCSrl58aeK93B
EcHzA7IngVAGlKmWlwT06WjjOmws28kBRDQTbQEDcWawgtfPXOfrEABAWhq2tIAgQXz+b6HXSTyC
zC6JonnzL3Eo2LNRBWrE9JOR0WLl0dYCb1bTTDQgEgoxhvlehWEdw+nLkr+Mq4eq3p0zN56aK88k
szBieMydVhw5Vw9wJhRRWvyrGwFK+tcdPmsztijqIXkX7lM3tYd69YsdqDYVC9D6Ke9dMhS7ld9f
avCUxWmBmKNT87/sm66qzjcmrEnuWFoWbEC//HKSP4p1PH91yQOuYRWIuLzMy84jsdB6B6ivAjpB
vWzQeReB2DNb/iewSQccC/9z6C+QbOgXv3te1HzUZD2clTbKJRDeMejNGFUvMXHc6Weq4hJxgge2
8AiHCSNGHE/NEVOMds69LZNbsFZYvOtDxojFOV5PzIosj1LRer89V6ZcYho1PwhSz/aiZb9TIDkW
rBCInNIgyt8ElTQz6KN2oGpjLoyKhSsqzEg9iu5x24TGBm0tep5C1adY6mmEc51zSU8Ft5yf2sXD
wp+3ZE0wLEWh7yTQhoFSjO4rvaOduevTGErq7fRe8gnA4dqvT12Ny5ogtv0pET+/N52Av7fup9x1
kNgPe0xMns6pe5E2xBJqufRbPStrFJGeuNI+0wUrCLO86Eo6ScnT9IT1cbsDbRKZK0f8McDwvQ1K
F0sqiw1j/wKZ4rcvAmyBR1yV3r5xUXGgcWEnZZcuQUL8XwUagbik3LISqRTXslt2nEIrYMK+Ktlp
wONpNXXYu8W+HVmRxwUJyUmcHqXaFFCtL7h3/3CrZ8/VPvgsmvQG9Oqax/jjrGo3kh/ISMsUkuc3
HH3aeiKAx//sl1T9NW4Zt00utwHWGaDInoMCjDHG5ZHh5FKQ7PVTJqJMK2aNHpHXqw1r5VLnItX+
js/eLXAv6RmYfgsLn2sNNagmJJr35fN3YO3QX+PE46g9tdpQnSE1I7hjxiNkQWsovC80ABdJU1sB
sKbKTlfbvguf1laF1f2g520X40VQm/QmmHBDXs33xV8EaSl/xHk/c2hhTdSG2/J3u6JTNSnyaMKj
8fP/HXX6Ww+HgoJJd5wZjmdoYElSMTnVFs03Pvkrd364mDY1+lb46Kf8mSLybuCx4jqfqguC7EAA
ZNHETcDCcIKt0an1koLhVCIltI+4luYaTkHQhCHla3GWTUXg49kRyd89wIefZikKU5ydbxM1nYd1
bWy76s2KFop0jMVwOOC0eCpprK4cvFhfXxR9e/Wlxs5FZ97WmiexQl/4ltsN1dx0K/wdzpNiUuJw
wPD+Ixm3igS1VU141qPPB4khOy6LvUB3INO2aX91zRLMXfzW1fQ6Q4o4Jue+LdkDBTEyUNF1j+V/
qbzvLFHBgrSRrQ8VZbca/R0IHNEhEV27vk9I7zV39ptXKM1awA6kw9eG+r0xSW/+hZh3b0eXahRD
3HVtUUuzFPq+4F5FMAE6mcWzpikZFpr7sLpY4CIrq3PHD31PczVCKd2qQV6UKiyXhShrYoRRJabv
6fo1L4pTO/LysQbJw6pxIIUfHVqEeKFXWbK8MaLl9bMddG7uyS9lwvI3COVpAMTb+HJ2007Ql13J
qRgEghQBCTg+GFmlS/xpPCoz/9C0EvYSmUs8uklkinnDrKOpX3OTFNXyTMoWUZfIf1UDjAGlkqmA
aEb/Qy6JR7WDMIgl6IobuZOX9CZOKDdiWMfn/6MgKCcA5fVVbTH2pIqIn/8d9tND92wZXxhAShlR
Qo788/8WTAX4wqhx7Pfm59Yl/s3ltKXyucj3QkDclEggI5jND1vDPoN6AUoeU48eKArJaFNz5T9O
A0y0+dUSaNJZWEZ8oAu0dI/Zli6veuGZfYY96bjrG2nzv7E9tjnw95WSC1a2kqHJc9yD+p5uPzU/
8kR2cq8g3SXbB98kTHWsWT+FV2fqn4z3SwxqAjschHWi+sfkk+r5skEFbpVOBlNnqeo6dYMuTDik
6mel5VvVCECwYpE00e38PkMa4ZDL6VKtLEma413KNusRhX2Mi4onug1KsAX3A0I0n83Zlc0O/frN
z2T2AKjTSPRezdQ0GFEWSabFnu+M0FLpUQprSU00sEVfikdpOhX0c+dDGbz2JUKLWAtgrmEcj6cp
uKljDuM9J2Y9dCz714LbfaR27uTjdsBKNncFwRPAQ8LLUJiL28BZ8bMbn+s3wx3UlOrME+aCO5qu
wZ+ELKikBDdlrTxbXtz2thAGypBBnhm1OKu/WQ24PAecEOVCDml7tsawz0MoipHPZvOdCqDQcNDm
UhHl4ck9fVXjfULDd3hpU8atyysKspTglVDKTdp0kJ9Xpt03p0gpS4udcYLmDvrtOWmKWpJ0DDS+
b74TkCjQxms4gQeyOnkFD+WJ8WI+Kg5OVibHT+YahyudV7ZUx+7DOSf25BXLyvXdjE34LTxzbKaB
yyM7Y37XW1AthqUxUvQcL6eooyOcHaIMFaYon7d3ni0CPWcuy5EEKAWsdyeE9DT6jopEoqNDIRYw
Pw2GDjmtvpjFS7tNC+hniS9qFMXkvyo2QXUdXmXk3e53j0Br8svJFz/8Xk69tpN3i2HyIzEPP8gW
q2UxUSgqcCPlw5EUPcsYdefibG/NZdFY/nEoPVYZNPD9/1ZfHPmScB0WxhUt3OgbW6+QDS/7uxUD
A0RJRcntAVH9O/6XWwK5NTdZLlIMhiif9UfK8viLdqOlOEWmE/+UaDwsWinxu7LzeCYOQ3ErcxL5
0UUaX5gO2/RdPWu+dQiTPPp9YxtyBdm2k1H5xUVMBeVU1/gukOzxRbOJdjEBdq9qXv9ENZ8pv1De
TEuC+t55/vWXdFeCCmrvr040qSNdAV4cw6xwqjPpmQy6teQZ0SpvPnBtuLZmnW2JAaE6CBPAerSA
f5Gr0oka1zo7Iu6xcrSR3j3XOyVIFhKNi5gU3nnQK1ksQeYJ6kx5EFFPVOa3HZP8h0z0sPYtmVWs
wdcWqF9xsZS+UlSx5XdPRkhqQYcsqgkc53AT1GpdHhkNu4rjSyilEj6TGw9vG/rzm33pLC4uP84n
CUkvBTsniZsEuAj7+KVAyr4aWR6X/RydTJPAE2ekU+S6BSDAsJJTje4WGOl3nsFI8lQYZ+ZI4wkW
dXgs64l1Igpb7mhnqjZjCCax5aTgq65EuL3e8GeDa5ZC+zYpsUK6A6wuRhdS69gobHWyIs18yg70
fFskRPXpX1wC9lUwiBErJx7np+CyUWzFnTX8OYgW7p1e8Eqj0Cn69TmyCqz7T+4bxyNminGAChP9
zFe14RMW8+rup0zPhnIH6DsEjz7SIjXbjyEMO5d1pZPU3uCJTeqX0ZnL23XDQtb7HnXHCUL6SjvA
IDIT4rSXuWOHkxZdKom7tTpePClqADKkzcoVluglVrNdTtblecyK04ig15A3SLQm85PuV5S6uzXf
sPt7kTXCXurKMWSKpen4rJOf6qRHXIx/ptP50jLBTFrUdjxypashcJ8NNi3vvz6G5zFfP7TuU00x
gQceCkHvrm+EJRqKR41DtnHRM9uiMH8lPIP4o9XPYP1IJNI5oXNeccueNMOSeFQpoqVqYgdwHqRv
j23pLmuTKGjq5MDsCBR2XG/sf2ftFvT7ss5vN6uyriqaHJBiiCWpVrANYMX27oOjaTml6IAhUbCg
87uCq2xm4PBViPvOpfCYu39vXDCuWE6B2AcZOWSaksqus6XBZdMIK2EM8ySYFsvRLtXyn5rofe/B
wfU52g3sqgxJ8Ksn1jmMCTqe5XRuuzV4Yc1px8k3W1I7Cywexs9jZXvYn2eXOsHie4NNPZJ2CiUx
eDphksG0XQBUGveFgsetRqiRKtRaNVTIrj8F6LIt7I5lH2WlnuANjAKsIUxzbVEszVwkkvrMKQYL
suqAMlLc3+8CMokJRMOoSwoyBr3t/4nDlFBh6yDQ6NKb5DyKZkwskMYU0O8kABdKATIsf/uGgFpS
w93sLWeXY9j2/xrU2VjIqTQgnnpjQ+aaQ0JbXErm/Vr07b9CaTAYWf4XL3wiAt6jxo2ThZWw5B5E
ppt0anGc3TR/OK6bGPxTa4cEkGxdIkHdIXVo8xPNIpuAbrOWUUSs/rN56a7kSVMP8Ceff68wjTfH
DoFPjw9wLaMOLoCdnJAQK8MQ4aZydKB7elfRritutCJHwtSEmTxYFWxHlaTveV+0BpCXbmNd6QCx
UbtBTc3U4vYT4RBbH8QLXfj4pwm7k8vp27YMjgORPRl3VvNuPowXSTELpRdNVM0PUdtHav9tdqyX
V73ZyXbWHwPfIC5u+gn/NudeUN1Iacfp17xIGNw7pviujasGapU2Lgb09PLmGZTwAWLpJ0IQjtQ+
gxYozaRdhmAqzFcB9+fJejhE8oeiJ0h1G4r3ak5Yx0Da0AlfoUC9lEBZX5savKv23b49nW0oTv2P
j620j93FN2sT/z2RwYcRkLkCRtyaRzvH03tQQs/ZKqYBjKKcBbZDtmgp+157rYOsUP6Zp5akp5mU
aeQihIhlcjMuz7iH5fS7FoHMwHiizfafdYA+AThPIIiVLww1M/UgSJ3hoHe+R/Rp/XE8MdEjI8f4
2Y0S51N1sFyU/uq9mSD+TO25R11Kw0cZ8VVwpq3yuXQs8QWKzzv4XeJb/Noe4FjU7D2YlDaXkzo3
UTr5Y/t7acUmzlah8274kWlCbKgMwJXBD27hIBUZjOw3cZqMpgKoCYss5I/WFPRLJGgRmPlIaWN1
kpEedCXFfX0HGktd4OxXtC0mbptMkNqu91PTyO/8lFyJrJPPEOGQYxdh3wWAt9xZZ7sItPlGcQwa
fvVVHJZdD2qAXk/OlygkPSHmiUeU+qn995Hvldxk9yAfD1GVDghV/Yn8JcpgZJtYDXL5Yz10eCFL
PhOt1pgFsPZpSlXKTXvSRQiWMlslL/XaCucccaiXE3Qbb6/0FPcEUqCPDDjtTZxxv6ZM64oTsS+V
ul4elb1mc+NMKxiJL4EPewhXeXAoEfAPMhglj7INPiwqUL8XfeYqX/JHZpl0A+IU9zqTOmt/ta2K
N0HV3WXrufw+kP4R3k4Jh/Q4aRm8fBUgdaulwolPr1Xra3Tjb3IM40UD6zD+p01wG7t1MrMQnkEW
kU43QLdLf1P3+dvQdCQa4y/ktd+egRkFeaQUgAwr5QDqLLHwNRdRwfRAygNxfuJrwsku8u9j4USA
d1Ah1daaeQFUWFYJUUtBpuYtF1Lv13qAqMgWhsZhyth1xEubOIJh533WEYAhfKuj2TyGoeGTjYhn
6DbnceJ2x/NGFrQatm0Ah4AWVKwYFT3ORVQfwyndckr6yhZI8h48jUwbYdUAFYtcbXz646yxYudG
1N/kQBV/+hle/2etiPvWGcm8OLsu2LB6XgNdpiC9yxBbU0o2qTHK7kh7Vi3mgy+vVCgauxEmiO/8
BpcpK6Ywef73g/PmxBclC+IJ7hd4aaPxQguVW4QnixRbXtVW/0n6VHA2TZU6+rapGfkp1dqT8wiz
SX4XtEJ9nROkJIUgwOzl6UEFbVhplYAtxW641iZz91yOvCQjgJQ/vsBXB8W8wNaIxDIvK457JTHA
OmfgDkEt0KDCAscWPhdji76TzWf8nJBip64yuSRcSRsBDYF0HlapOcny8aMiqYQLaqav2yTJIL5x
mc3D1GRt4jpw6SMNBqzgcPcMhuePgYsFnjl5ZG0zfKRGyq40BgI76mhpu1FM9qRTBM9M1NddAIZ7
+xzno1yLTbdHyezmVxDt6WJ6wdhCJHC4EyfIgmV/E6R+9fgI2VNFwvVyinuc8C+z2r2+02FNctL+
G+9D6mwqbVKPi0iHPVKMvkkphotCNL8oCMin80ttWJlUvrHA9SEwE/AJpL1aYMdX8JrGxSfyknUc
Xbhmjd4SAcJJkfpbE+M/q6vIqymajGfp8WXfp5pU8m1NHV2aaMteR2BqMntx0dRHfOh54lUElZEq
36K/y/9BhlRAkK3WMee6kjk7GVjA2747Gv5h85IePGFekOBBngp9VVnvvTPHyFs4B7Okf2mI9RbG
JpDFyJZQC6Tc14VRqS6xRPw8U1KPsjQH1rWFgW5rxhAeT9mZOEikMeS+vQAGWqMtzChNUetyDEkv
2B2MTskhhHU8irjGmw6SxJ2uEFpvfOca9p5E7yMO4cF2N/EZ6uufJVSWD4v8BcaE3bURXfQWXY+M
djplB+jB3NnvJP4JwWTHDqVsru8xe2+r0HpKR76dhwXz9mYvS60ZXmXAXW47EgTyg/bWjJ4utpvg
m2y4bkc2Tnwhd2N3wilrMJRYHgOItQjnujfOIJY4bfTH9BVRMKfzYSx9nTr13eqM+BpZJYwhQyLm
sK/pTf2PlldLOz7VUzA1/+zNuRZowQTOp9bwq2nxmNNR6cVLyWwe2GIT9O9Wq5myFCWNZdX4cND9
zsqDpSo0KyNYp9iHX0pv4tcN7mRv6KXqHUfRhtnzxPIUMfN1PcF+qTP1yy/UPM4qibIxBvwKMkDa
9KsC1+/xNOY6gjvlLIA33vx96z+353kYhl1bg3/buiMyNIH25VoP4uFccSIEfBnesqT+YaJAsrIp
SMBz4SLyuVQ/g8Y05GwE6vRH6b4TxDNYS1KFduYZaXSz6oa1PBXqLCI6zgsCb4Z08zRJnnG9QT7f
3NJSl0zGIdBpXdNCJWbKQok0g0OtRVdT2Qk0nBK3wOUITKPQSZOgfBeWRkBG0A7/N27vdWRiceIF
3s1LaF+qSz7JeAki54x5BW7BZkWxZnOeol3QH63TTbgP7/X6nOyTNRj/P6sJNoPuAU1TmSU3G37G
nHgpQi2g9m383Lg+GjpJecRDm++KwWvCK2Dk3AnC03fXvpP7ZjF15xBiYPr0cDSmbYuhulKNwmz4
DJ9m3GuT4jIn9f+MicatzAN3DymNJzGJmcAZnhb1Kqc29uNOaS3GaMCCGaw7p9SBxfEXWGw/T5kd
ExFJYzEmLP4lHSLY8XcSL2LGuyTFVzO/plqN2M5c2rCguO3MQozP2mH5Y0Cajnu4jG5IwoCvRtck
JBPKSGy8UInBwNuADQEx0IARjkNYj2Byu/XWbpcrSqE+RNcZUttF+lGEzCc9DuXzq3Zwh55Zv87y
Cv79ARPZXWwG7eVJ2WpIPChBXepLor6cS6WyTZAGMBjeT44xeSummWLyStTSYvb3A14nPPgWYFew
g2OqqWzbRIiEw1cS9Aeacv+W3O5jcIztBYzH7jtjcqpITerBhH9E41ulBUAaFJ+0aFP9I/AsIsNt
Z/UtiqbVZuJ4ESkP95ezMalCacNnvr4RYo/Mwc47klQTUr/acric/rofnClODONqn5uAX7t7Nbcq
cttLqMvw7asNecueoo1J3lxorgGY56cBWcm8QylG1wMiJUZPCuwNPVhWmddtUaM3kWQ/ciAjBwn/
MxkbtXnYxF2npw5Xw8eVX3YgYopKrCLmPIVnizuHQvVc13c5rwNAV/k2r0V+IpsDALhoJWrU4Vio
lRDPFMTUuFVZ97fq3QXef3NxmWJ7Q0iFShMU3H09lw13zEpYf/SLFw4iKeJ/vg1qQ3zTq8yHivWx
FCS3ZobFIvHCEUZ4ZgKLFg4oMH5V4+5tyOk7aOinU6jIgzhTvE9beXsC06llhf6kytabWDKOWWwG
jm2P1rsYosL61OWxpVcJjBdfGiKLXxErlf9n56PkVCC14y7Eu/WBZMLSFWpwyXQrJS4mvlEFZ2uY
qZk8woiI4aUsHwYvyS0OiYpkfeqZyAgtfNFSa2kKmDC3txy1kLAC+1rwFBOkClF96jM1P/fbawzK
fuEY5DRrpPzbn1GNfp6m1fAzsgUnnN3J1S6Nckozbyloude2t/Hay974XGhoS9aJCtLhRqoHLM4Y
1+xty+ksSHAzRzbdGtP90+N8L4sZGAC9lkNCJ9uaFPBpoYjicwSFcxCoUyPuwvt4n6uzNgVNehxG
HOeFy3PBdtlyi+EHIJo9tyOjbF7CXTzfWd5kelW8/Tqtj1rFAqihu6w4nRXiCPXmQy3EJxLTutzJ
GFqP77X6rmgoEFSyBG+uLsk1YugtmNKdVuxoZHuE/wNSPlCwbsod9oRx9QNoBy4NCbw3iUplp0D9
lxE/kpeXOG1pChUBjCysPXrUvq7p9EckqXVnnVvjXIVw952ehOp4sXB2OOFJKMbPQyIipVaIIFUv
3DSd9tWbpZelOcxEoaCcaY7LB+TE1zZMr8qlCJUs6SeE9lCJIE0mSDF38CNlPnI46bfhDwqGliMr
o4ZVbOWbBfWDodUxgP3kQAJrf8/ULFDnHfqNqTxW58uxqdUw9+YcLMEMDK+ACqbVK5mu78of1UG3
oE5mytAr+WOt3ePuNKIBihot10EewC2qlDejsq2i1nlY0RU7su+HJTghUOCu5qP4yl03/YG5/v1W
Kgz6cy5+sfKecUjNLPprhKRpjNfHzrbFAZmU4zK1ga/fLkn8wHTJz6121KSk7HCjHj5LQyL/P3r8
3pBZl/6igNJc2pDai12J7GxWh0zrQYzuiceWGttKomBcrMn/fL4V7tYI2tckfbzLpY/jJAWybQ87
/4//KgfEuz5tOA5UJQY1o/jK+ykwm7id/MHVC3CD0+036B+hlW4crBZcoXL42TKNDcXshuJ3Yd8w
cL6cSzs+d1ZKWmBjY7GbGJ7FWCQ0iMcEQjE8IKn4x+7t9g5dYhrR0OV8J9oDl1qxD2oJlheAa9Sg
1aVxb9kKKOfB2CGUwQ2v+Z6qQp3mo+TSGc5fegGUbMO/M2c6uIkCVPyH+c98uoJIZX0ASPWHn1cd
8KrJ0OXd6oqso3vIKLax8Yt7ekpTfQ3nzsfSuxJ74+vxxkKFhxEunapcAK7+2Cus2oxUEpj8t1dI
visJs2bZLDsmTSgRF/ZLxBautMTb6M6uLjdV+In1RAnNsH4z5Z+NGihMXf3BiKJow0qDrg7o/cgV
1QPAsY2A/Cclh3M4H8mzEIa9rNNNUT7EC266jX/a679tBqiNWkP1QZSrwoH/2EHtkrIbExvIU2EG
1YhJUvxHOQIfecbFVcLzXEzR+3PuebAA4hd7pwGpqk/8exEgBb4wcbWve3X5uMJkA/dz0ttbIoVS
VYwwnqgxws3w2OATe4Ns98YIy5us3aNphlOYUi+YSb/4D0b9l5nIh3bVdDHObG2I081/3zI3HyyU
w/7TJFW1UioOA44KjuzhcvwcQ5yaqbMZlUTC3rFUUdje7iZrb81OdYvt8J+I+jXKBzD+AQrH3D7j
3rzIvArEyo39XF5xGXmtdHzjbo4z46La4GR+QArbBvTkvnIvZQ0/13iJrVdHLX6jUybElssM002h
aebvB+cCv7Fj6rFHcvlSEQzhmAoRSjWyPK/0/b3S4LcR/4VikIeakpmOlfA+yx3dJVHJtysSApSQ
SQQUbAdUCfpoHmGMmWl84d9jzp1ziV+BF4PYgNnAuIGwcA6+fgldAS01NI9nwGVXN68C5hrpOG+e
UJfSco82PnLEFyNVWePCfbdKBk1DdC/oukdjoSkLyiLGnsNwbTyZUxNZQV8AE7FnAnCfulBt0jCc
YgI4kuLz6AlDk0n4IdWZLSMmDHTmSrU/4ltoRQrh8HgSIKcHS/RKthPCIom2OdQ2udClESdw/mja
dZqTSc8CacWiMobbo7d7OYudumlULdbBHHZ3PEhIBZFrqNonp985xlvhMAtMdtDvz6SCscbyiq2c
ux9QCwzqRGYjoACg+9uQ5a8512s5F7hz133xL1nrg4k7FrjHOhc0E1iFzAGaGRj47l828lh0KRsK
woUKUPhftdAqsBenPGGnLMeuECds62TtMWmh+uvaRA4JD23aUJWL4b2hHQOCmQRd1FOg1GeJmh0/
rWsMluNkA1HzlHAiAPBxbcCJhpVd38RGFRuklgmhvxRt4YlnpwhQw8DiwuI0M3ezinMuc4eJs8Vk
V+FR5HBhDtLx3ZJRehNBj234tbdfYITy0dZQgUJfLJeESrJ0jH0rAJ26OLrW2CMZWsaMf5c3QMsx
SJEcu+PSko7JeOMLhaznchTMEl7oKZMpxdz441jHsTviP+isn2Q1ynXdpFUHMTlq7ToDbU0VnlvN
Hh2SAxxFNqPL9lX04BAr9DlNILqa8dM+uWD0+JQyMbSEP7ZyhKIrdOBK0XN0JWvczn8MkA5QjB8e
iz7nCASzbDcC0mBIQNRMMo6+QkIDYhOIZnlekNVNrVVM8i6tZjsP4HA5nXFGSrynwFbh/Rl5C25H
mJh82vfHL20QA+WqmDGGA1EO9rPPvKwSmGwZ9WgX3wXMWzplR3nK+S+DIOdX3p2cSxlO8RpkSiXq
Ux33HW5U0aSQmmPP3rjjGiSXPlzFL3KMYBEygMU5+hbtkkrwC13Rxjnffvd2hGIbe+nxjOo8MrWB
IwMQ6Ghc6rjYcsoYrm6feoUtdegwCiHYKXGX3Dib3gUaTt7Zua5Zl1Rij6FilZNFhHD6mqPKx2/3
Sht7SuvI15XRL8dmCya7eMFyONPj6UZ15ClEAntFshAoYtZYURzHhNCtf+GbqfzJavP5J9cXkpJh
kO5yynevw6bshJiUfDLv6WrHmlgRuJmqLf2Cz/74yDGRW8W76dF0YsDYqn8qoR92SWocWyLVI7q1
FdJfrArk5Z6092J2sAZGQKJgg4lIjv9q1V+T7cwLE97Kylt50WgvTvFx19Rkz3+5zY2Z0LJN2Dab
z7QBtGr4mqUdcnoH+p4ZYFyd8GGcgrj0r4uCpoGkpUMjtEyiJn5/ATIsb6MBZfZw/SEsvYW75Az3
Jwv0n9jxsMshN/+2wx4q9p6lQneDFt3guQS6PjkEDyooSkULlVVgzeNVHkB+WeaO63cl38Lt2Y+u
eNO+HRawApMjlJzJdflxdSRMORgefhdltgi03dzNqOmCvWcBh0r7aCXRZ6K3uci5ntTpP6fB31Ge
IrQQejtUEPZ36V36Qsde191XwRsAdblIR7LSxfYSMfuVZtvbXl38C5FW7Qa3zprLM5tJNfJOa6Oe
da2NgwLFgtZmqyUhjiTT24id5u2yAdXxppS4yCqbTa6m67dZDhU9o3ZdMJKMWhQPKmRShO5ql/EJ
DZ5O61gm173Ug4OMoVvGtg/xndXYQHKXTRfALaO8XZLUUavvPmVuyrEA+Bmls0jWjZ9Jj2QkGUdS
40SNpLA1DxJUBaVDtrb/IUpMlnSiTN8c/Y1swQo0DFVDT922amBjifvyMfKVDD7Usi1zmM458S6a
SuJXjl2XmRI2VqY53rhdDhCBPVMR2VZxSltVKwfG1VQXxjwGknLMBvfCcBJi8r/vgt+vkyvF8Lm3
ZwbRcemiHwBWhppHkowWdcEaKe2Jn8WPYO6eiQJ78Ncu9mpBqHkw6pwb8OakcyodLK54xuMNMGWR
F7T92+RIEke3tBxDn2SugLjGBKxp69VkxSDgZ2U+fOkrnM94RWAD2OHeoqKiSH4mpJEji4GMT2gu
XnD2yiV3nSuagNsZrB6usyL6LAcFAyV9A+Qyc+MpRGz0UH5gxZJy0P6cLLJLk+7/ogi/d2Q2V9H5
7z1C0BuxrxenD8cSR/T2byUrqLgUNHbzv5FV7a2FjsOlTaPsSoRv5c1WJhExwPyPvc/9KESZeENi
lmaVur6g39m9z0C7IjjPcgyy8SCjlxUR6ThYLA1Q3mw7YBmxyW4uO5xcNmmFDLc+iCZVBK/zeUBP
fAfba6sssMOcE5GwUIu9B8bj/NkZ8ztr8koP5mA8YYrx4hRPS/hzXaJzHCHidQEBUQYfmxJ/I/hD
sQxFKhUW2DuZZEhm/Q6QBBSYSJ2ydQrS+Po9d/mQd0FeBKrZ+tMxjKbEcUDy57wyqmgVNXcAjtwX
2nUyocP8nf7hUn782ughcpjucvYlvCTYErtk3YN2OJfoglRWkfmlhgDvytTZ4JcJCMFK9Fy84jvs
axE+BDGUQh/Gjwn0/MVcMp3TniCGZQ9IlJZpW5Jti0Fq+RMfpB7OjdE/V5jfiQpXkFx/vtYzlP4y
5eJmspzU3/EizhyV9FRpDlwioW++srxVoJuEHD9z82RXShUs+g4bXNeViPBY5IVJT2G+AkOa+fex
QijBA2B8w0iKPgzN4ya9+5MKVlznWmaMeSA4LoFlkKpkD3Gvlg4IBsj0Uj/nBY4kuGoo5mm5iHtf
xSrD7+bA6qUA0RWgMjTy5Uq+lXVIoo5Wb5rw9atC2VSMSKitRAw2SgBRxVmycWjBaWGkGyjsCVqt
fAogKf1Ru+rYSenP/qE+tBc76Hs4BoeB2Xm38BUO2srIxBkaZwpoAxcheGQKfbBlYjTJ1KqqktPi
Qh8wmED60npQtj2fEBiWJaiHVO0/k5wVmmuXL2k/L/3gWeccBXnQy97+DB0RYCVXN19XcDV8xu1O
HwxP2JNplnlo5Fp1X0OKmuZeNwKKKYuV6+E4XroBRoPwhnsk08XkCIexLv7zKIPQqUIm+QB1kggU
odQyruShgElMjTVQiyZ3qtPNIgznUgtFxopDbMB9vgpPzekP4++z7K3gC2UhkQBk0ePXUqEnjixs
hAfV94I3vLHOcZXFCqZmpwKmj8FfQFv14Zo4urJLfkJoeUQ0ENL1Ob0w3iahL/D2mgw/YHdHxJhJ
cPktKrc6hrjUIaTzAARmWiKFjgHuQZIAyix3gh8A3x4qe4J5mHOmWaLHnlhuUIjiepMokvOGIY0p
6sAOvQDQqVrH2Y78PzMvlixhC6+r/OR8jzW+aCix1VHQ6JBXEn5zm9SndnsUVm4YGjO4fpdy9eFG
Sp0OeOvURjytqObiPzdCU7wAV4bSe8N/TvtxOVmZQrGvZWgipd2c11+N2FXtTWNX3uwMg55w4Oaa
446NsTLuvYikBnRCJhuVjW7G6fP3NGYUehfC/rWeTu0UGSStOUWIVJ6jyA/CZ/K5ZetCqFtMNk+b
MkDNfmjqUo+TrNMwdTUepdE/UViNp4nKwhuZdRLLQRQZSSry45sDNew8o/810LooGS6C7OC8RtmZ
rae6p63xQO1UyrOgmPK3J2VznKFgek/EbCPXfdw6ESpeVIHOELDDsLxHJHwliGXQhLnqHbKr7QCc
wQ68jNSjIUREx+cyJp8jU5u9GAMpAzzHS8IuIJYC1h9JreZhh2O7vNHb2hYkYPRHTrX9tWGiCrk8
T8ayr01DZnj4bYqsvXeRVdCAj/YP7Ku7rMOxMap55iiefy/D8Li9CqJbvVXs/ZFVa+u9CvdlMWQD
ql1kbsW4bgQcnMsPBE0tlIJUnAwanFGdPpFAjWeWsgUpFPj9O44TGCL58fOQ+BMcrFBFHJ3ofWCo
kwoB2mc9L69UFv1ssadwgsfPaAh6XOxBTmeDkl6FhZ0a/r3XjnIdNj7jOFUJvglHVKHexbGiftcc
XEDnmOBjAH+9S5PHWC6QlTf93/l/di8EulBARd4kDh3M/zWjIFx0iEI/0ClGuYIYPXzRwHDFG60f
HywndnBWphIG9L9wDd/bXaZAAs+GTWaWDr29JJh/p9oly/NlcXdxzTDXhVIA3Kq0ROJs1WdbLX/P
0ElQikGvbtaWWHyta0otaJOxlOmyLRETiJ7WTR0YDNF9+d8CM43r6dXxL0EZjI6M6m/HYvGljE6p
Q1qizx9Tdqi2feH3l3vmLSu8sA6/No7MFCmEah4K+ndnGzbnVPiee2XbWL9DwFA90rS5dAsEYzJ9
vxFB1nXcqwEGd6BAlWEMnCoNfgg5ep8VT57fL9bey1nirSW/X/Pok43ZoCP34dSFgsc9DMBLBbCb
jCZodYp9EYnbOQJvq8gzv7MxaWxWl//Y8wUYXv+n/QIHTY+LTGZYzTn43mBMUzMHLdlQu8oB1t9Y
5+lHXsHwFAO8mc7Zn+j0eNKHYJdFOoOWBmls6bWSAWxoje+KzSqSi76j1+JXwC122IRBSCA8WnhF
PX6AiLRhTE+qmR8SMYdBEVWeaJrm2G38wOdb+Hc5c7sWmm6kwAL/8MrDk4MleUMT9n/AxcxoneMW
DuEBcABaG51lpf3nuLfjMYEgpywOnFYNMKrhW6Q5jFb4eKCEIvuN8Jtyj5dqdJw3pV19l++RhXKp
O7t+guJwyzjyd4cbgEu04fCBDs+m3wGfYh5/k6Pc0HIQmaOHsYgT2FOCnI91DU8cV/x3vL53W4Ms
m6aLB8jBPZ9Yk7WoI5TCWx0EjOGJWkq3zo3Gwyj+xsCF/RKqLKTevuWZTXCqfC8wwt5z7TJ8wP3x
VMCSTM7FdWzBSgB+AyR1seCKdAjRMLnZ4pzleyru2wS650P0EEv98wx+kbQ/XUij6HAEDrFKFP6i
zvI3q0D9xjB4EqMSgwMTrrD1nvpaWg4VINk7cp82UH4taNr0Jubqm0NqMrtTDyAlv6eb2K7Rq2v4
py8QfcHxDPcewkIwLMIk3Jf0BYxsheHHcd3ka935fwlWlhPfbjrJbSfN0HNnDvzvX/fe6a7P8xA5
x8xQ0Y2IwAk1jbJNwHuJOgwcrbHE3RCj9e3WsImYWsNeLmAvkBLRTZlRZHDJ91gXDn4Nz1VNf9w7
L8KwuuNWw22adGiY2VuYuEXIv62eWPcfL3NAWe458fAsBazmpJP98FR7/KZ4Klb15MvhSvAGiuP6
jXkxV/GzQeuqghHhozTU4YdFycxBxXXghUaJHXNPPCxRRBGxFGdul4YEWoYJ3YD3/yvd1CpE+/dc
jLbuPygXTD5BtALKI3qyjV4VDxAOP542l//tD7czScZBQo419SU4c7iqiZjHBSNT5IZNKEtUg7f1
Do+oX9IVDCIExNWntFazozgLVhXIPGeLMqn2J4n5Ax6wbom5YzjguZXrbdJDniasq6nEr21od0A3
R6xsTVqANLyaaDiFImPsJCW7NsbBqgS5hcHC9bmS37NL9hWBiCxozy0EbXjdvbsR99Trt3NVpFw6
rI8M3d5hn1m5+9PRg9+Fb+pc6dBb4pFVULwI0PuRrn2rJN450Hv0WoI6iU44GRvZ/4DiP57P5r3j
94Io0fT9UxXZgzqZly9SYhXq0Wv1O8HNJYO9okEle+TTESE5eFvareAWn7J+oEpcwMB439D+OQ3L
DUo3cYqik+WxISnrncy2IZQA3EWlzF/IIEFByjrltnMYDy6p3HLj/jnr4PGh4V+3y02ttDHzNnSi
BeBUpsse0xPtvPO1P1TUBW8cmLmIXU1FVcZIXEcgHj4CPKAV6ICMdKVMKZEZT+W8T8no5W734ORK
Axzn+t8MuV9D3+HBfXCW1hMt8G7HTOoEiyssmGMxsJ+9zDzwhlDB3clQccxLNAEby4W7RPD658KU
QxHzKBzpHswf3ftddK8ETzZDcBQeCVD5aOU/HxIsxNhM2PAxvZkhx71xsf3HAjO84CF2VOUKbTOx
+mc8iHGnBTkPpsa+k/5idP6sH1zCtLJR7HA/XbbiGcFUKvKglmyxFzj1wvp/uKlY8JvpfdOK1W1u
eSddjAuIUsgk2MLk500fd7BGrSlMB90GS1CUD4eoFWbs76fqUcUCCr0lGQO5fTCFu8psB75ySOba
/tzCNbOebFF1lITGKVS7gAu2QhlI/xXRytwiqn+haVYisc5Z2/gST8Gn6b6Oho8DHjFGbVze+Tt6
I3Rl7dBlgWkmwNErE1RLcwAdfPuej+A50ApdESeod3Dk5QHre3WMQyvrlZV7yEsEweOxjtgAxFbp
wtvOinaVOxQgvuuGJmlizRs1Nh3BBZ3TaaxxW7bu8AvE9mKQprKRnzF0z6oy+nHFTgce2jpUbZxH
pn6VmvHVUvzJWysomtJILY1fxdm/8DZi/COhZayCISMpm/vWIUQNnL6w/y6GvV4RBeQAtEA74Y32
q9hgTEgPnizpMy6Go/mLGNtA9RDHRZYmKOZpA98tVahNTPcthzskJuegX8lxYCTgKfq1MwdB0Nss
TMjMSA0aCCl0Kx/NkIDp7T6GwKmVKZzOdz45oJ0Yiq2Cp3+46YrSDbtxIiK2pc7wtlMiJZeSIdzj
KtkArhblRPekCJp2IIJVr8vbr33zXbNYfCNBJ1W/cfqsgTPod/w9y70g5GUhD2N83jrN6qmUolT3
Me+6PPCAebhKXhz3njRO5Po5U9/M4uaJJorzaiWGGw8CnVYDpEDsfvx5R/8a1BkLNH/1+PXk2lZ3
FFu/4AymwtRheiqGDPC7aIHyl7tZk21CuXMDYB11yXm3xUanKWzXC7LLjT/3vhv7HSGKFuT0b6IR
anHYJ7IzDcNq8TBqrf70thD2MNJnioqgVwm8pyMaqnsypXEgg+VKobYtb2P9/NITlioz1OO9RXQb
ZSWReKw/RwVzNp5MuuwxZKQHbZ77/yHlKAbgYgHbMb8GSUqpI6F1zUw9ZwJflpONnuOHlsNmth0r
2JYZTFDRlQgBZx9+r9hrzZUzK8oS//v5dQvVYp5JMTG372TnsiDRHxdd9pJSbmXKUeqs8mr+RDPC
mkAH5v0Lz4Mb9L2MAgAlv9IZEqMtS8kJEOsUIhMtR4TfqxYcpXqssPX8Z+dyrr+lYax9MnG4ODr6
YNYIVB/dagwF5DG6ZM9B1cgsAWw5UsVOzgfP7U4I95Rzv7ArP+VpfvbHVMsXtkrzHH/hCM/uabze
sCqBRjBVW2gGAWYnmFH+C7gpfKJFVSTDyzjYXElYTLGmpn0jZEPYeR7glR5wl7YIz3Frye+By33Z
0j2TZFOf5++ew/kBEueF0thjzDUBzitKl8Iopze9AivZDE/C3pKUfc1gw9Lj3rCZGEbhfElLCGFt
rS3RFjDh4iqwNSRdDSbPBXD5HO1I8TFGAXUhamoCjdb/rzdoxYSlYkl5718AK/jRoDKwuhTxE2IC
RVGAswiP0nSoJchL9NSmDbBDUtye3gvp7mphln5NmIETQwUlHGagQKnhxtWLzAkV4r7HujpDe/3J
532iRhwiVkGp0MvThsl2iuYQhVRYWgxysgOPkRoNRUfoouqBLMG5EFuc7VaRQdEfYqM9lLbzqrxH
l+h19KRLVF0WZkUsQP+ehY0VR1XLZM+KhoaJOtFEwTXneVQ64T2ClR0IBxy/wy7FUxQw3wb+4BZZ
M7iGgPTfOczcN/mrEzLUr0plmxppwj3lEf2bGaWHLAX2UimuQeizgweCLZFlQI5K+n2yi89taQRH
B6+0h1cNdyW0DBDC+cb495WKj8MfO5bR/xh705ftLHFmGM7OMA8xhlv13VF3MKKGWPuRfywkfXIT
puYwH3HdULZ3rgWby53jKGlTWAqx59YugM1v2nz+H1ieb68XXXu6E/+eqBtMH7P8GMeRUDrVO9Ja
oWpJf89BW5gLEtmYChkqZEYF3p/RERxap5/qkZnJ1+2ItvLBWQ5B4KjFGAbcUXF60G01rPMLjgn4
dMeJr64NKq7mIcBYGkK58BMxvBIusK7UMNCgib0Tuxsdh2DvT88pwlui30AohVzKUDhF1BXEy4ok
MBdA6aAKeCKsC1NObLEN4aDA+W1uWQ/SGU9S1qW3bdLRCUE3yF+hKa0FgnYTn4+nUt41E9Nertqb
RBSSwMZc4YpqeSrsysgBjJbsOBJMyoWUj1L8v/09sOvGZYozQihIR6QqpA7U7CDdos9hyKb0AlZS
2kYTkLuGAzHnj/jOu552GElZ4hVv9zMWN+GWUxXZ2O9vNxpRusU2Xk3cjj6hKa1wlpJfTx9oT5nr
L1fHALDAlqx0TfRxb8gItr22D2cwQDDjj60NYSzUENleLT/s2QVho+VRhjZVMDFIAhy2FQr82Sdf
FFcdQ7TUpkVS5wICdeVKpaE4RwbGMOMCwM61stICoBOKvVma4kSvPez4SEuimmuu5+LrJ6d/rixK
pYYUDeywO+U8lbqH00Ef5ueWM6qxtMBYt0Cq5zqg4jyh5W4ygRP9jn+i/jGBajlHJER0pyOv47D1
IXVR2yFvRufKJj+f+Mz8hTMVTNpNzEaaOohTeZqY2kCgQpZoYIRFJpKc/a3LwaGKyKVvg+eZqU5D
ttC8iDfTOLa3CwCDfHQ3mAPtgVxWpXF7cX/xQ9NuSOvRCDDQ+0ujbtJTAV+lEZ3HkbiVp24GCvQi
b2eAgPUCa211tQ83mhueb/FZC308sTLo4RAIWUKrEAgyzARExAHLUzpoibL4YsVD945HcTMKbJWO
BqM7ePOODWojT6eE+nVlVN6knJ4kYRbgUtMCakjSLGiMH1jsbLiR9W+mKlKrOWLFt333HwbncWZ7
ctYzed86tmsYQW/QRli0XlxjD8THKJmQtfvwyQn8W33H8uNIjLBErhTEmnXTXov5ngKKvRIqln/w
o+ewyIa3IIWvGBnURN5/MPlorO8qnq1iPndIK9wYJUno419BId6difsIA2Et8bc4gv/bxtj9d5Or
GjI9E8hkRKFax6mXGdJ20DxxZKexaTFmeQurGLdBui0CAOd1XvuVhhtFT6lNVX0V4Ty//2OHJiHU
yNLH06hk5/ccTUNwnoaMrJLxQ0yx9R8YmwQQ7nPyNC9Tk3fl0HQEybzgCSb8mWwsLgFDlT9sOX4B
9vkpXtfdI9I2RjKzjAF/tJu3OVq3lnBl7ljQrygS7pdIacslTWBiCVgi8v3GZKfkGGGOSsxgXmFQ
ovZ+PQX2XRvmUgPF4/wUvpRSqKmT2fACmOJUr7TCV76oShPlyO4TTmUZUk8GSo0zWCOjFFLSWNkZ
NBrMSxGQ+J7WKfB9ZMxt26HgMeOWKfTULDqgmpDmkNxQZgQrfTdaHI4czuEz9jLObTFx6C/1jFei
8SSQtg5BEWtC7CadR8lh+IKtBiNFHzjgOy3z/u+OwNxtfWsCXZpKs0f+m8+0c4Ko839B9MryCrV0
l4tqC/ZfoTO9HG7kmDRMVyT0+D5BK3EVjSATHmITQc35F4Z/XeKPB3DwbiGsK+qNVo1CMnEG/bE6
Vl5bY9I1LuYzoc7nZj78JdWVmdJgUxnNV6AESrgs8WBRgYKrd9bl9P9RC0Ed4ijcxGWjZHZmqnyg
+5oKvUXo/VNI7LtDO6fpM6lesi0+zoxz9svaYkU7o8gTds7yGre2TPPqmBHV3K8guqmPGNEbwuem
X/GCqMNl7i6mi6yibcsg1Z7u2+XWC7eU4ugpaMAWbwI2aBl6DOIxjcTBmfJ/f/M5oHNorf+VB/Pi
yS+JFWYMFMwLBVg7uzxUtq0xQH/5Zgf2RzuTS/eekll7gVHHnyPMp4HWQseSyqhVIVL9iIp900bD
PIpZuTHeS500CTTsJfVOAtPXE68ws6lXK8oqwoRrwa4KwfW68U/5SW5d2xg7PUVRapKlVKjbIpYD
NADrOEc7A5DhOcWmQd52poCVDk+jZPj6Kcdq5Ds2n7tRpjevZi57xolJvmYCiEiPgX2CSWI7wP/p
pU8x02tSp98520QMOpDct0tFBsJdZQgE3L+ZSzrIKxvVZnTKt8aru7DwNF7I5UNk27AYVrHo9L6P
hrCO1qeK6hhi7k1s+YRFFSh80c1F5O6YOdGkyeXNqthApOB4AXQhF/YaeEG28jE6BY3uhlyGP0iW
lX9xYdPzf1FMMRTY5TpGvcjxsQu7WI1CuGqdMTtVLsj+oiDM8hyzovnB/0jB1RZoTE9iGfTQeGwm
Aq+mX1YOjHf+GcaDsxKtmEhyw7cvT/6LJ9dup42KE6JJQLhBzJ3tlOHSOw0hoBuLZZs9+Ea/LhPk
tme+Yq0h12ofe2DPxbcp9DlmmP+aGTn0adaZe0vsKI0G2QA223EJH0fOcD7z/5CHV+PWXjO3t66V
ItWj7WiUSq2xfdt8T4K9RP/UWvaM3s2kJEKFRv90keRgzPZMsZOTccwwz/KOMWZIv2W7ihQ+XVEU
BOxwDI165v0nHOeBAIgRnEZIRu2Jf+lZDZaXB5cGV+ENkeU4dGHFx7FBCJRli5h6bRCcAi1LmZXb
InAGeDcmc4lj+Bj1foNplEfiLf1Og3lBEl8ZhLplByqDEh6z9lXaXi1ZDM4ETpIHj32P+wcPZ6/j
QVHDwE/dwkQYAMa0C3FUdqjvlerFc0JBz8fnDwjENtutej2U92CbzYS2WuHpKquQV0+flhSMnV0/
u41wtLi9lIcP22rXQzZXe29xB48qB5Q4GMQJxLoG6+umqi11oGN+8h7uFk6NoWeZfwuxXS85frJy
uOGt1yDUPr2mwekWV8vXlbsClC3x2rR3yPk2AiepHAAWtQzr7GwDEGb/8jZ+dUKNf33YDoRW9IS+
cpYdVMs0DI/x6TiCzolAZXfaNZD1Yq4+Rnd/pRGNWpXjix4M7mJ3pciPcHplYRvLj4cKHqQJMBRo
pU24gJsnw5gSxk7ADQMfaNcI6dJJ1L6IbPVUQKAGmdpZvW2i6/8GVmNIAnUONf7x6tdL/AgWi/57
zU+88AZSHnBPBnpaA2yRjtobSq5KbP1teQEcWrFRZYyen4a8iExam7HPVb1KMoipSuQu3o1ZxGNE
kRdWxWUPe0Ppb3RS3WTagLOARr3L5hzWVb2IwQt/3WS2R5R2ykDWjUGuSOz2YssnLNiDY/a4ZU/3
je1npopfqMO9qi1nOLkxkbnazdPlHf3yD1/eYEsYPAfj/mWsrb6orNYC9uAujkZ/VIehPKdrdKiY
J3IFbJ4HoXpbT+6AJalrS4bZWu87AWnC217W/9iX9NoRN9wMpw3f1ReSXKNw8IYvxD1UV5UIVaTi
VHl3BCBUEjgYDEosKZgxDEaHHW6qIUTih1U3BTcTX0TG6f6+V1MJON4Mo5A6gqKoR5VZ6TBfNV7g
z910zL6hl97ix4qLKAuBG5IWk8xNRfutems2n64v4fewUbLnCZM0n8afxt3DeczTYx7iK9EA1Ab7
lrLca9lGzq3IlQubwdF39pRwVUaA9tjxN/JofH6Is9Tlk50zIiq1cSEr7ZcpbQj5dAl2BVufcwpf
SRJ8te1GRfyyE8/w7Wm/+O1ytd7Qzm8fn2tsLIqiC7G+VxrI4unnyAV74L3//aiVnxCPkXcBdyna
kULy6cfN1MQW3ZZ3z9hFoyTabv3xms0lleH1obAVUrbvKC8yjEcf9I4sKRA2J6bArBcmUM2DGhZB
Z1AeKsg+e0xPIMsuuDUosNBcIaQ7SMCPMbhIXss3e67/etmxdPI9yKI+qD7sXntE8sBCZU4mqt0u
1yypJP/bdSwBaFlG8vFAQpR0WvaEvRZ+qJlKxngliYSnib39fkUBWm92/hetLxrQKOLe6bSBm1NF
GwpA4NBj2m6KW3foh9/Zkha9P7DghvzmN3XEl3LOaaUx/hIM0aOngM1sTudK9rM7SOVzdJqLn9nB
J9SLkjWLiIf0tqhi8KZp9WKw6nnLJ9GaoirTDA5KhSXdYh4hqNTGDPGOUxY1bKqidWGUdhNt33ei
1VxBZ7TcjqXYS95sKdj6pGDk1E+Gh+t35TKmNumOo2JVquqV2o37kHgFzacn+1CkNT1ny2bPMN13
zSzzqdalyhHjSdjoGzH9cPm1wdoHV9PYrPNT6ujDwaMdmLhLRLN6DB7C4VSCDOh7qEpRh92maTT0
6xvKFxjrpxRzDyUOlV6hFTdR8omLJ5HmpnqQafz8BKR/ZMsD8QSU7/+Dfh63F7NsYP0ErDF3oI4K
zp+KwJTjLPlApyM3IIA7DGKSqfQD1Occ7tTjpmgEfB9QFeQ79vYBq2Bc/iYTQDFz7PeCLpUHQs8K
TbjqpYQQgNHfHqhsZAWRfy/zQXfxur9/bowQtl/IRGsEtHN+SSEp0k/s+NiskraisxO9hT/vkQm3
umME0I/1XmgVGLbObELUxEEgg6lbfPWXIZy+LcaiHdepyUNgj9KNSPbyciQLnQJLSABMk8NwSTLn
c1GRSbexPSgf3SWw7TWYZ0Q6I/075kMVWa2mBiEJ/63rx7SL+4PLch8rSkufRIYGjsx31L1GwAAZ
8zCm9hLOilrOr37X/ApsZ4Uw3ckDwGpa9e9U92Wpyqfsp8v4U7ctYB0rgT0E4MU8xp0d29n7MhZR
clndJM2mqCK/+9HjhYs6bOAfExCkNQRHnJUo8StZ0rECcfyvht5R7q64SSKY36WtpS8ahBTP/jYo
w2f8yz5V14BAap79l2D3rnGIBLGYMwqFnVFwxDyXEEm7ahuD0RfQMNMcpYvNU47xyBNi4w9jiQKC
2g1HSVWMVuNRIlC8Fdf4vCAXmBb4WF1ldWF/W85HQXF8VZA4VcNEMK0BgcIFLBvlmloHbYtZD1gc
g+YMNVTWgOUehnR845pIR/isq0VEdpLhAM25EwfWVNDu7Y+aCY35SsGVM4Wk9JiD2FcoUSohKnVt
NaBfP52pOn9gjz0vIcsaMgfB7WQIZneRapq8BDnLuKyubNAFQ/n2IirJNXMpoUuBkMdZ82w+Np3G
wlTMW3+SUeN/Ly+QuhPF69M5/UpLgu7HOkM60milpvASEyndb1/nhZoqIynimMbGz2ikD4svDkUk
P8weXwrN4O4wzlS7uFxSCCB+8YvkoqeNw6tWBuu//6namxRyHgi1+GZDu/0vXWVif9IyLYk5TOUb
MKyQ1MNTpxqch2TtK5RUWAJQ6/y3LBNzCWYE/eJdfF9pF76Zi5qrKJXd9bUe/w3lgvVbXNgMHlmA
mJ2JrOtoUNJRNsMFYgnFvIm+2MD4h2idzB5XuoI34uDpYqAjPdDjRPTX0s3EE/QDKWFR9+ISumdh
o8cZSJ8sAyV0hBe8PlftHbcYtb2jx4cj4033GAksHdG0jPNepMIxsLgH9cPs00T/Qrq1b5XuUUw7
xrjVBKhLR5pdDQjRONLhjtxlLmzgGatd49UjcnEdVKXCOFG4RKDrierDRpiTFpw07ayyDEfUytIQ
nk9aIxc1rGjKjRal2q8hWU0G4FkBmJRGOpD4QFNX1PqXnHHjlBKaYqIVQyOJZhq8JsnepI+N6H8z
pIOxIwkIUe458IbcPmzpWa9LeMNm1NKDlhWRyYpe+YxJvsuplCXnD/qB+5S4PrGdfJwA5gR09VwZ
vbGvvlUSCMA0vOY+FUg20n1PoSEkQXbZGhJbyG+2OsVeMW4pPz8OXPU5ou4Rz3qRtKoK/CIsDXyR
9yRlaayZu/eUdQ7oCf3iSHojz9NaHloRyJRSkHuOWoyjytWfTcN0ZqjPddyTMMFObDn3Y3bWYwm8
AAFhpH2QzTwEajNRE7HYlRr9c/ls7pxOSlXqjlnDgpT//Hd9cYUaiYLKfFsV3mI9S6NnQ3uJAY9S
phZMmExh0VOfRviUn3rbfKbreFnFl8OCWLB+kkKarc2TD6SOCm50yg7u55VwgWBnmRZYDLkiVQAo
3XWNwIp0Mql28lQvN3UvKK9SlzicJRPiKGUMU9p1YBiO69XKOxuhGlFkMDJ+kuIC9GarHvf7zo8F
c7gWuQ79tsfMsbGWIZdlaot+T2uE67buGWvmE5JKuwkK5Kxw+3jvZlp+2OWJeTxPRqZEdKSWXQLd
TQk3WEo0xckKkdHrpKIi1WQqSs1rXxi5xcXHRST/ASWxIY7LdsmhU+G+Yz55wgdGqK6abC0EOt/D
Y7rCZoXaY9RCDQtXxBZyRyz0Ma2RaZuKISKpuwA9u1Zfx3rc8WZ/7jrJtF/y1pg2YVW873ynO7fA
zH2e3COfrrKCQ/DnHpZX9dePE/IDCK8/BZKIbN1Eujra/R0KdQII1oNloZZxX7+niyDeNb6gBHeW
6+AcdKrSZhs7nGUR/Ml8nTiv3It5uRR33WxC/NkFAm6Hl7qSRkbo5GebeY857K7mBvJ/fqrE+MF4
l26BWFGp8UKP+e5McOUxIz2GGCIBu766svd+RWXSbdyCCmpxfaDPp9O8LcGaRDl0Q8828t7Quxbe
opZ3OnqQk/xsiaajP1X+bybzqzY3942iuAiHpp4SpPI+kLP+bw+8fUJHH/j4bTJKlm7ErvGDp+Vq
CXOKTxTLCB2T9h0OwMsVplkD8VuCmG8jVs4JGZzWjhTsMSI7SLnydUVSl4+caPDpGkh84e//4r6e
ZxX/audG6ncprf7e2tsOILtEF/brwXXBdsX6L7X1JOJFw2EiBu6OvqEN84UhU8tYzDpim+5S4iia
S0kUHMKFB6pEprdkdyflDrnrKG+3W44cVOzm8xAXvvOkqG4OZiYcETtyWqywehdpV6/79tDniiqj
6x+Xv1A9Jfl1WbeWUa2R4nQTRTYkb1+xD61ILgMf4Cv7vDGcJr/qP14FgPyZttP5spBbWJZZHCyn
D3+iff8S6pF2vJCylKYbGec+M6NM1sbdKB9fQDzUmJic5aKfNJqAs+iT6GBW67gXCd4nXa3YBRie
rhzlStdb2K474jsIAXJRf0NCnhvsvODCXw7ccVd6OpDYQHFg1yal6cmWxIkUqG+MQN4zlTdHVHPY
Hapf7EZWCl0091xl6nbLwJ3FwRVikPTZTmtDG+t6dxFF7OhdDCbfrcML1y30bHNhlGKVfn6pLdIJ
QSE4WQHyxypWveb1IQwXax4H2aqKdjDtBAjiVd88OQbYe4Kml8ycStry/w3ocAzeOQ9Z6zJucnb9
5C4/wOJ15byOW6flPv7qqaIRAfIdwV9CdLypsDJ23przVR/g8RnL2fVjTrNU7k/oy0HuOSiIXMYr
lZnBei7dxk+EObCTjd908FrKouoeFiQhB4Vh3oBkn9CnU45SzGQ823KjtMLcEnkvZHFBP1r9cZ4W
LgglLbQ+FIyMryXvsMPhTnjazIMhypvAxu9kzP0Y5yiYSWtVTltBRCqNLlsMJgCHt8VLHUgWse8l
bhk9W/rQO6pKXTZ55kLv7Ose6Rq4iMIu+LCvQjPyIfzrzejvYOrlVDAA7IhVQjGZBxeHFKM58SuD
Wi+RzxQLuJfqJFcsWmC1CxVJqKWT42Po8Aa81mCAJcN6F7p8HsguWORPnWuQ/Nnt6Gpwo+eb9qL0
vAANn6ZeMyh6UHrB5WKfDUEoZ6EelAfn4O7BYkF5LXgN84xTSFHHRK7VnCDh7tyD1I+BKu4KUYVz
2qVSlHxPZLwN0VGLHP9X+7Apx08Wa8/a2HAB/4Np8INndxf5TfkKs3kOWa4X0k0j/lk0k5dIuiI6
ZLYpQikXJD66tFgjLwm4I6Vs9Z5puc+/LSQ3j1WKFvTYJF/7GXIaDRUFwe4AVw9BnT2MVO3PYgfH
sTctJlGZitMjbMJ9DP13lDX5Z9j6XIqpop9C7UoyEBABWo5VCRw1ojgIsit4GrxXTSgDyVAriKZd
WChuLrHCn4uFqPiixYj7kXO545ggvhyVEUJAyLX51wecdiQFGnLh6i+N66HBQSFxoxxscOgPssRF
Btv08gb801R+vjCH9Xit01ck7v6Er/HWi3hw426iYM5iNw0HqlKnjhBfOYRVI77fSgrjfP+lhYOi
gAsplvA8r6vVQaPuzLgnRUbj5lEue/csEYK+qODNI8btD/z+QEnZlkbk4bLmgCkzbybBQ7hGLzcr
TcML/zf+KUqcf76oaXYwO1O1NSQErypeCXd6VIs21PWX+Z9iyXGU59DltZyuFccyhLlw0Yb9G5yI
eqcWRWA7BDlb79yGUc5MwRaQe0stNtnpfPMp5dra+YuHarPajZFxkox8onTl8sIeNw0mWD/7+3Ln
hDDACZOvxt9q456RrHrIqpUlG5S4t8ui7o71/tV5xnLshaQbL2hUtrZ7jqS1J9+yJFi+BJfqeFWB
m2S13dfYmOlwJ+IRhkwyJURABClH45mBQC0wEL+b1S4BX46YQKy0STaJQpQI93yACBcUH1Weistk
8cvuxI7kQu0CNfNr1lKE3pi+VhiZnfRRylhqQfjIB1bFkwm9wdVpelelb+9iLwoZNVvi9bSA0F15
i8hlF8JCeJaxxiOl0folJTlZyhUz9yVP35qlZxvT04C25+SCLiy1MetrWn6XHEmndvceibwnrnNb
TPY81yHY+fEbUgep54k6ZhzMk9VgrgSLh96DfxUBPdhj4ohpj6ralQUaeMJxfyFmwiD3UTyAFmzv
vb2ng6kfv/MPexnoLXl4pyoBoQcSoAf2+I08AZaSw6lUic18Q/cA4sZGO9m+0xvnh499XVVwzu7Z
4cK4NRMcrMv9Nv+JgPmqdjtC7meMd9Qwfyak3+SHWsHaxTX563y89LeXVfp4b1lLpuntK0BrM/0C
QIBRevsdRvQi112aLMxTbDYjDaSU8KkES4DQ9rsO+BVeeyfnUvbuplGBQIxvxeiTZ3lWFPvgMsWs
fNVlNCl5MF7SfEoiO0Ayl/M1E5ZAaZTVAFIdSldIPYDgkWJhc3nvedLcHuNSv8wHC+noMswBldAd
l+Tm0kiaIS43nnkltYVtSkQBNGBwRDrFkGPPXBim1MCTu6I2kcnmL23XlbZk/y485nfBTIo09PnG
Ogef882Qcq/bHVpeRemdnroZDYmxCq6GxgEcrW7256nusC+c+XSqx39MtVfbkTArglgQ70nk1J6r
zXaW7KtqG7yNqjYuIa0/mG5Xh6jykUQZEAVnbOc8zF5vNitw8JUniq7KVQurb6LPp8UZeNZY9ntz
uKuO1GF73010vzWvcsqBJtkK9aNi16MkkFjO1lHrwtybqcjd0BfR9l8FxJS2B4ZQA44ZkvvOM/y8
jPjWTvOdkR+hKOzfMkbVj021OQnADs4Cl21xwj8ZILNFMeszDFFWCdlUOtgkP+wHTgT6iEWNjsbr
O4rsCoJfemuT44UlvNiNbeYp5ppsRIpAUHgnEvf0Mj6PgAgeasu9QGjFfIo7WA8zvLO2LUNhAShy
t45LXciMTIiycoPLX/mnMLDPi1SoEta/eDeUoGiSQIf8/jE7E+Zy4k+iRf1NZaeUa0DsRp4s922p
SB7xeqHDLPtlSm6BjKnKeO8AFSmtz0/JttfAkiOItWgj4Fy028bBByuqloXDsNwvcBfG1qIzKha7
eY1E/C/w/UoyctxrJ8AARTUmRFxl9hz94sS+EV3jEsWjBFvieAehMb8x3oJj98XZmD7FPv2IIDbV
ehFHSzrrvIjA31uQ+QK3Xnbbocibi4h52Z7cN+B4FCtL0syu/F75cRUpoKNNpl4sPPIHAzEDZaCz
3CuK9IIA+n/k5/TGqUZWb/GOTof7anrOET4iyvkrxYb/ea5Imv9p5R0OILKV8r7D9piv6e1+b7Zl
451/z0v42+gZTrkl8nJ8XNYUPShzil4vzOeXv4KUHEDTtrIkcBmuxyPMoe2UkP/nhqMGWBd0H1qr
iR93QBaGBgs5/ylfSKCBH88JHji5DKKEQPvezCYPOvx0xRCZ7GiwgWXktVlMb9nWuMQJIZu9RNqt
agx2ub0GfZBVYZN6bqkVd908ALitGOp90VPVABySu2qrLyraxfuB2G2Z70rXComOH//pFyjDIMk9
klxxk7YQ/pqXuQMJr7qxo6oaXbX/zrXVDEWD03ouJGy0xl7ADejpNA06rSWSrwQRzvysEdewitz+
iIyK5FhoR3dihQYRtXkbMLZHYwd5/BKnTJUbOKFmhrHD9MbkEm74Jtltd39XXYNUoEWUbTaZ2OSY
hs1yLg7rBzrKKD9EsO4kTvoZLe6NV6njufelg3T5PuhzKx0UqFYdzodNrxEqrZolhQ+j553n5NBK
dJF6TeVZ5iXuRkeVvXkjUyQe3kP7HfUnuno4NaZeXjDsNC3K3PnZasm9Tl+bRa0ICd8GpqZt09t+
LDcAO0U2OHN076MAj63iAVE/agHjHjPbs1FdQ5upEcE0MlTFgPFGPq9Dpx/JNu2S3l4rQJL6cZ3E
z+spoVFcHYDMcwBi//2MqsLiY4sddkzeO46LgbmGQ/MLCtVgpDIJD3o5aAu5FxfR5gW8gVx+X0Vg
SCEd95e5n5SITz7FIBa6gSK1Ny2CDequ3rmv0TnrCbZL/GTDQJUVRCvCwwr1gWj8KFAFVNlOk7M6
fTImpSv2ivUma2KowaC5/5o39mYk3NtaPHro5/xMaTMnGaTrj3a0NfqblU8H8332ER+lBSFG8zqI
I+mW3GUFI92STndIRSnyVdlIsbHq/8Lg7+46dcdEfDL5HvbPYI7gKKH2FIUQsCIn9Bi9cFrk/ur8
/sU6tOvqCoXDBN2jB18hAvR/gaEJ3MpOClOwi3C3YVURxmpg5VEKqlyo4zU4G9XPm1ioLlP/8Bay
iQOZbe6arPQ1TtVoFGpd8R5BFZVSTSmobW93QkHGOwSZG3MF5l0rwEX9u6WtTk5II44iDGKbRp/a
SNQbFk148eaM4E2VHwn5X49DszeWpI6+geM0+lupQKE2kNp3sIU22s647x7Wa3Tx7mzxvvINNI+s
c4Bo3ZEgBNdLznEKB7g1CbKZBJcjPjjn/CmLHLzKZylWG62Q7EO7TKbO2bktmJP+31cPYsvBL8yH
KRmlitEBBTsxlZkvm+JccVeKp7sSIXtbqna2AZWFivkFGkrAuD2H0Y2eoM5i8hz0qeErORchK2WB
PmBC3YKstNDyqKfdVvcukfo+dpzc7s1EaVXB+cLr2svA7rZuJNMG1pEnpAIMJz5yPVpHDWaLh2Ke
J7WMQRHXNUBLw+R8P98HyDgZqEc4gduMHqTrMlUD7oIiDnJFebJi7JIE6kx355A5qngP5Cfitc1T
Atjj6TYFl487FfvOMEQ4LtUlnBeTqrIoArWItQaYBC6DBQiQbGtS6SYyOOmjt180zEbECG9EP7+W
hUpQw5oNXIW/ax+xnRA58eRdx4D4GEdcH79yvOTuQYtX2IROdvD1b22r8z279GaN2aBjdJgj4dJv
3//Vpb+A/VzVWvuQ6oaahgXGe/AyFsLpWlIZuvrxw/2ROB/nGqkHaBG84mLbWfamYigqzwrY9JRc
NbSw8BicQCCKCdgkxGZoIHuaNVvjhua1pqgIAhL/YFkiEGbH2aqiOcIDzdS9Q5cExbt/0SeIG0Ei
qRRpvCxyT1Fz06oTW/eFGQJugY0T4KzxfYCdf3rccG0AtO21/crb+d7z+nSRqZpomUA7W8lsJzvW
XpOyDzIhwR9hPl0ZoY1VcWcBhXQQhq37jfvwQzZ8KpmBlKPKtkTMo0J5FxRXVrhHN1ZTxKJicr1i
Ibz6B8tMvtHpX7Uy7fExoCM9qmEBk9dL4Kp+7q7j/8H7YP3ip+rCRLGXZ9qPLkT/6hYVpYq7VNdV
iOUIlpSY2SGtMzgf88SyJsy4sGcwD6HkYyRzp87QRhGgwj/r+Mf+ugxkuCHgdKL5b4LNCyszkfXY
Nme97L6VGXfB1iRSS8Iri77JDd9pxzr1zSEhg0c1zxsBEpq5qsZ9SF7eXB5Glx1f3o5Zq2HolNrl
8PlgmNK27hvDM2WDETIlKaAkos5t7bF6GocDTmtpSsr+T9/b/8BecLrhWfAUe8aDfwC5zYqhlbTQ
K1hQhH3FiA3Yp7Q+0Pcz2hffrtW0Gb++lpoM+yaAL+UpSPSZZ7WnG27k5mzzgXBVS/SLoweGN3t5
ORKPD+2w3aQrqhf4jeKT7vmnTbHsFMTa48TnaffZNcKj9k03bVKHOMw+QoaeaEy7UyFuSEMxPb6o
J9HShJ5xTqLl2nyr+fGvVqa8QkLC8CAR4CKgsemt2hudzf6aGLtnKgFLUe7sMZoEMbCmEbDN4xZn
Ueq3Oy4m/JvsqzLHQ32VYBaqkB5C+BFJe+7fRfzSa6LRbrW+gqG9XcMv840/IZIbU5ugrs6BSXwx
3bXvzzXcqWUGpf2if7x21W/T84aE7ULp/t02Gx9jKKdbhlVMX76ZrJsqogsqL7YzdPQNO8AXb+8S
FR04qlgwmGbSjAnHFL0HFIY0sH9iTitmoWOrVXP3GlvQ5evIr60h+TzhzLUnYlPLOPKLoStoQCkT
gT8LhhO9onHm8tPUmlUuHsD66u44CS6QZjlK/44Y6ZZSSyZbjyx84/k7lxLN8rwm7KD9kAp/IdpP
XRIL7VJaQSCWg5JkfF5cubhqDNMakWc1KivcqSQXilwt05XGH+pMjhAgTNQAmZr5uW3zgLvPeK/9
JYJ9xSSHMDQLmJN6M3p+PjtRorMleF+py/k8z59YUdk951jBoHKtwmE0FDHN6VF9wclLSIHxWFN2
y6kFlpkIBDdV+uGlLC075ArloO7eNABYkvcSFs2svnuDVt0iV9IRkJv8YVKhOUGA38waEULI8W7G
bcYz8TQWq/8412xX2o1gDPfL1bhpe3KDdqN2bJipKyTEX5deEkhETxR79rKpcBOtRhv7fSUpdqaO
MACRhx5h08P2dOCk0M2K6xbtvKjd1q38TJkdbB+qJTgB+kMKR+oLYFGGd1YDRiCCYUYMXzyL1e0X
eOayXVh89qXmCzmHeyjHRR3z5BucweATR8nHKm/M8pCVhqFzknFpRaYEQ0R5Vc+YUGz3SVdqzTA0
wHsdADhZ2x+qvzYEpEDVQMXRXqdqsJDqmNrGmuAwmRnvnuq/IMkiE3DqCGsf2SDNWlMpC5DJGoVJ
WFIRWqmfMjbBnqIDAzjD6dNJffcpukSVwyE3ZL2oRN3RPtK2VX09i5sz6x3DwjGEA157pE0gUmZS
ix2XT/AYLZwSvTPjd8S2SbmSkC3KyGFEku+fo4jO4XomxTB+XYRL0k6T+X5rWAwpuvHPfTi0MqHF
1lTorfr39zFwkEAJ2De/F8P/krBMw02HM2Dj86b58QwOAqJBxM0PeqOpjfoA/HvF8B3aZ/f6d6hf
CDJqnU6cbeZLwin9YhC2DlsIlqtcGZeYKpXDHyDYg+a9gKXgkQ/qhRzpbksWFznZ9v4V2Z2DG7Su
6SWkjgrB0NQlSGeiWxTiI3WVRXwkyNIp3XVf3xYVZvA1yNc3+EYlQDF7BnE71kdeqSDtwZE3Ai8v
X9OakLzSWt4pmo4hwqpwmBN1+68GwgoREs+PJ9VdmKx8HtsNyAjR/68ws5n3TqVVyClsgEO8C5A+
IXfgtOwow630NufFSn0aDJLvNc71DjjN5OHpW2n99KtkGklnJxZJkEAIQUZWA1NxXEd15wp3XrOj
h1AvzOd0E6XCl8USzVf1uPfhMYA+gvZTPsx1gnuXI68An16YV2hewqSzlhJt+ngWLm+a7sUru5Ni
Q87EUAfec47aW+REs5Fsan1Fk4ztcQ+HS5QerMGmyLSbcCQi/lIx2XjPASKjPa5i5mEKrkajeZh+
UwYfFx9rwsTCM4hYNZPmyOVOKjuQ4IUJUMIHUBZC7gWQNq9T+/Z2pRBzpmdpxvDePFxFwJRl4SyK
DcYYk9nCvChRL9ho2ayqoPGNbLHjfDD+xDiaT+vnsYbGcJfzkr8XJvYWVQhC31UB1krqlRdGndsn
EESajlX+1Y2jy7OoGjfu+4HleFvjJQVH8ZB5ZrJMnnmoEGFv6k2/6Srx6iJR7PBTZUeRNd1boShU
D8lz3plirhhCkscOMh7ml7Ot1TUrf/FdGc4jh7jd00f8zjwFE+dLa6ZnYEIZ38UP853yTOeUVn2V
DdZzPr7R6H/ShP+pyp39Rks7PiXzJbEWMUE2Bk2jWF33EZt1PF5X0C0AKUXUjvhYv6+NjJOgkR0R
4ZEC8w7oVo19ZX9OthK1c7xT2+7GhzuSt2Ar7Fi3aWWk0538mRE/U4J3R59vCgobEDivk1EuqiEf
qRXnqdRINEnzQhO/MuqmE74sJ5LdV2sbSumcg+RfPPX55TxGMZQiAOOMB8V7uG/dz1nelNaByFiq
EVVT37rZWZF9eBr1TVq8rm5SChmlU4S1m/T8zr3meZLPEfQsLmscZBAa25MlcOwe900noHnulGzI
HCJzndp3upk529i+pJTaZ+qveA1TBC8R/AvN685WUjWp4Nl1EyAh5cA6Mf8J1bhLweTGCtLQAXJU
UeT9AZBZsO2bf0usFL7C6eCt6mG/s3a02Ui1ZfZII1TQLjfeRyJjL210V3RKOLetavS/BwBmOvwp
JnFuGZ3fSeqhvMJtXLdyIAl/yxNhM8GDFw4eq8Nn3bKFcgrEqXXmarQlaExYbDQNwtkvPrzqkBmJ
TD9KoBMUIQMG83Tl+6fT4+doM2FuiPmLQnxnlJseVxbmv7Hvljl0bkd6BOosC5BvwLLsef5mBpCI
5LoKnW7kk/OBdFJj2+EORGLKvhi8xIxmsSpsWSmERxQFg1cRHbc+r+FV0Edj5byTMRmU4bQLcAYC
ETBIZYvh/Bst8VOaZvu/G/qIcNFtKRlCcZueTX1UV/YnUjO7z1BgRfZ9NffpgeIz8uAsu9Zaxyah
ONGWXVKCwfG+soTGQfPixnnBDf5kEhJKy4jPLLf/Ds0G/bfG03GjSVshaR0STrHXOvwGchr1AVbV
TKXIR5vojsolHrGdJDucQTHiYw1oWSm4X/Tc9HZ4DgaeLvY1/lxSUaSfcfj7+UuDbSXgHq8eOG+u
wKoLYFo+2WF7eSe7XEZc7V7WbBIemXvmE9gZj1Hq/UdcwT5DXRX2Jw9Mu8MvpFkfYENwdg2tQm9C
hKkJ12qn4yuiGCrCHvgZ0fkZfWncyhrIhm9Ief88/z16frZQK1nZnFGJNs0TYLi6rH/GYXkyLdbS
iXk/3qsU645gL67hBMKMzbIPXC/3/v/n6ExrvcIa0v1f8d1ZNvEb3gs0XHZRDS4POLJvZpe6/atR
FCuhbzLHlIvFwRaX9oKB3lHxDLiCaPYqbkdBgwg3bHVY54UCO/+wuLAvEvTt5C4UhceTdUoXYU8x
c5z/5Zbg9613X42afDnmIQ2z2G9s49atdtyHNvonPCp9k1+kvJZR7Er2nrdO1k54e5ZqZ4O2WlAu
dkvsMbj8OTIzhPS8QU6w6iUbNHW+uv4gaLDyhcL1lLGK1UQrwYJNEKqi8iD4kLg5gzS8jZPsHuXc
m9qE7+/00HHM5vsR+BS1JE3g20y6fem3uI90ULY+mygDBThn7brVuZaTOjKxa/teV85qjMszYI1R
urS8r/t5lN9pFqKAanb613l+04zcqmuxNI2fnm2SL36fW4DMVkcMHvqne8XGB0BNpaebUjnBx/Da
nJd70Vq9nDCHwkgTFT5PlD81dqsPH3xyh5s+3W2Mci0r8TX+d3vAFkBON8S/BPHDVTkeuJGdal2L
3CTVS5C7tDjuuaMIMijFwCb30wx8thJI/MXvUhKkKs7ilGvWhf52MOgMK7mVSpYmKw4MdmzeHlLi
mECvfflejzzJ1WdXvmBNVlpst7hZgreKtoseE7rLE2l76/pqlCizzH27YOfmndOVqnaohDGWKJFL
pFX4XQmt5qOIn5UhSwEjxdlBc+Ct6wzUyj0K5XaUULif/900MhJDTUUAd1IWjcaM7iIaEmQXfKKi
sdivlPFZt4DyFGZBkUN8mYjjwQievm0sWRWTow2Gcq5hHYVCsr5DtEXp5BOjZmr8dteTTOxMcgpZ
8IuYU3ncgO0mB0uDBsuzIw+Ov39Ikk2tWymAxeqVGUyOezgKtT/jVhtnzHXqIeV1RzzN5oIAtmPk
ftMTeVvxK3pO2JbRbHQJ1HP6ewGNCnI9PR4U+hjlFJMlWR6iacUBPfo3avyx6XlFObWcK7k80mK3
Z81TsIloLgZ6kLm5zx8LqYNLUVKdiUU7tV3iTiPUlqPxS6lVqqgZ96TjlXOY0cyVtULXIfkuwB82
LaJhtXWd5RlQxbCp1osJFEvnD5O8bzlwo2+Dzor9OZ51p1t3+HXE4bXjaxbq9o9utqd3YDEqg2lE
8XxK+Eabb23DnlV/+uy6cT8KeLuLPmwOTnFwWpkye8AEBTOWzwt0UgihYJkojItksuW8rlnS2nEu
55wzbtlnl70Ue9WIAXbLQ4be3/7MkqRSi7Ii7um4hBvgDE1hkE/q0CiNk0aFslRaoxH4GSw6i02S
rLySMnaKBqbyv+335CCOVTjJh0aP9nYyIsNlrYm4OIsUpTetZ3s6IBsvnqHJJxblUhW+yGYOcLTx
bikmOKCrVJYPeWXS/zFLpqqd1LFVGxQOthgLYunJkYgF2v5TDpO518ZQUvjZqEtlirpbSxP2V3Od
sX5dqrKJALOap/FcZJ6y67vgs5tyyCBGy6auqRfLIEBh+OTIl5HaWi4cAWdk3zHmhivj0W+41Dfe
SLCQn17rtW0oGCfAR5I3a6dGXyHMsjvq9+EoRZaNUfQl3WONQOVpLhJ+/8xg2FK1vzTMQ6mGscCL
uRSt4TXPwC6iYYYtomrmIbWjJsbQV8i5+gv6pSDIOI9qQkPKVrpgNN+ItKWDEegkE7PFNDrm3kUw
2HIwBde8Hl5AeVaIOgz2X06BGAfNtjfo1cq/knCfcDYI2mTklDpbHXJpyBfmlS6T6362cxq/9d2z
O5x72URwA8eb2fwceBa9qMGC/qVgWi+o6DkKihQhqF80STeFziQShj6qJ2eic/nDir5DjgRce+MW
wdYh3hmLX1Tv3zxFdtYRpLyHYK5r1xLW2ABpzHHl9iVDL5j5RwW96S+W5T/WMA7u4/qB5iGQdKK2
SDE3LD2ZT4Bd8pbSKF0KI08Qw/3xsE9u57y6D3LahB3KUSan/ztSpYIT2LDAfSthp5FTsYBy/sBT
geLvsgVs/JyNtvAa05WPFM0Dof9OCVdmURIKGHZnk2rN2mzL5r+FqHJvMjMPNEHTONmT1gqVCeEY
TNr+Q3atx0SwXiv64YxL3F56QVaGOxB48ONItKpPKm9iWXduNYdLaWGeD+BjiAyf6Z3RiqKa7rh5
zkDsTEkokKem5kLTOuWQ3oFzJLU/4E6HvOg4C6Eu/gf7pnMyc3FtI2RWI7oxnECV4UsVTSwYJrKt
NtUIYRYUEh+tH8zN3bK2SF+1RVNMwEVocDDWN30irwSyCGus44ePw9Mdpzc2/OYBRbX5s8CJf126
CqafjZrm8FxibkF+hE3ypdr42fMsEfdmxi33nmV3c826Zl3EfSUBdKCirVD5fcRFqj51LKQGyS/n
bUmOQskxMfEMn4d7/QdascJk/wh/jcwrD3lUyHIhMjiFWA7rlRh23UWEFXle2I/zloUAFJhmrIkk
siPUANeBd5asnnjCyUvvn/mR96Ie8HAPupqYcQFMKkTYTXWJ7NmZ1fhOG3S3Zsq4vzeRujZ1XVN3
E8eeoZ8ZpNMwaNQd3MzApHAfOzt2kEvssKcShAjO5wPGH4DxN3Wk6OTq9FvLjP9ttjaarJR/CFqn
K4JRNgQ5M0UzXUbJKoDRCcQiir6MA7r6cpyz7avnBTYmwSS4PXMeOM8t9tkyE8EV3Tg6/tA65HH5
9gwNj0EocsHFDP/iKHrbyZwPw6uFxE8HyHHbg0UFIGXzf3UZZO+7qxnOLTKk6sCHgzcRLo3JpQRs
MKohbVCcub6H3i7DMzgVYkwCJQyJ5tqWk21IHYLDPf2uqdao9SMHtZwfz3UhozqMaVAgxDCQvi94
xl3RJJ5i0Fs+tXDKWwn41TQ+CGczv2EdG9rVxx1S6A8djZ3YXA9GzXmnutSoAmQyxGBAUS5Za1aD
oX5zUNpbdnwhPyArL7N5brsV9FEA9VPV9DT7CKHauPagZwOKOIFaiAPCG0WaQSHcnBG6Zhn6umDE
ltfha6REc5SNgjEBvwlAfkIdsf7ZQVwmDeEPb+pFxk3SVkRIMfMR/Jw+YYnfEsqX/YYsrSYXA42b
LQbCwidhwPf2ReUyZr5NhNP5rsi4Nf5DuYPwfkk4vgnO3JPWaKVfHEAHxzjSSYcSGfzgaZHwVccb
qacmxSBCHlOXz8VdrWdXaoUTyHqBztVsod3GacIypYsOmHfNC5sZQdR7RxA6GTba6aIO8nyQB3Qw
NSw4rZ4eoaHjKWgs2SNly2KW1yJ23RaFOkeX1/P2frpX1N5VnJbgSrKFD1oMOKugeIcch6nO9gVV
SSxekGO0FgeuQJeERk3ae+W6h7WHRZo4WiM5YACVUXjX8wkShAeMF6441nRfWkakdqd0rWcPRakw
VO9zvWrPGfU8lfEySMgqwXKGUdv/QcGO7W0ofsFOvK6ZvvOg2bf4zxlVv7XshdBYk59xVt5OszG6
vKkK6NfMhK+bYWdud1SR1NfbhTg+MuwAoPeH1oLAFdPql2cm859UNz5Cvp0lb0mbvnbaZNiP3mnm
XmYevwqY9FXnyU+ATcNGHAA4Zfq6KFwL/AmnI7eHgzU+nbjNZsBemviriUnN0ckOX+SaOr1Zqb2B
lv/oqybcWX1MBX1wfMExKUslZW15pHWaeCxxKJCzpZeA4Fms68DotfuEX2Z1GysriPdTHfjJcNya
bJpLYueWjjfnl6twCbSRnoLWYEkddkqu83kYLYzZB3O1PfGYulv/sjc46ceaB5FbOpVYvCRHZilQ
D1yR+HD+nczFnQ7NzBYiVwVAUmdaJOgogL/gGYZpdsZFoyJq/+fIVQ+PQXU3Wb3SjT+eTh712x6h
NBAcH+t7VFgyk8p7JLMKyQblV+vRpH8uBICLozszjDMOaZ1ZS79EzfFxP7UwWG+1E8IpezEs+x5J
nxrbdoA7pWTxow4RpPzK/tlVmuGFOWpQM402ElCsL9MyJUsfUQdOzz6J4uujvCR16P/CCaD44uYh
DHzMHE4jqxy7bKnlqm5hFqK6lEqoQX/w+/XXSVcEHTJH9DPC++YukYRQ8xP4weW47g50TES4OX6j
GDLXUiedXqtJvVPsKEJO+Ed1TzIX48iNkHsHQhZdxddauJPa42DQ7Z720/YJtRPh8XpIt102T0En
M71fb4APoudpedQVL0fb4+BuMC1Qk4MiVY8BZbxKKhKWkawh47oCe3tKwLHwayY4jVY0nkoVYHJj
Z7iPPSIfswa2vgc0p+2XpVyA7phBDTITP2bZWXzXwuPYQ8v0BHMEVl0ZJeSO70fhMs0ZDcD5Sgde
StriSSFC4HhbA72AN/K0LMiRXoJ3ZTXQHVzkvjWZvuwNv8CaylSit16wobxSK8515716j8rOMQcm
SJlhHe+do3BiKjcEFn4qc1xXmMiu36jrXz2R3YRzbkUY9uMaXTA2tsQwUCLCBMDfPmxaBmqovzf8
Lmcg0X8aMHLJFMN7NWaG+NUmqLZk4UUh5R6W7tk2ycSyHC9ghyPZA0tsIrm3lW/KzO63MyiN/yy2
dyxFXDBYKria0/n7E27KDf3umNH4/NLX48V3mPqNFcWrDojAGivK6NQ3yEWSLn3unzqGByJA3Wu5
WQE+G1gxRjR5QVcf2vMhZ5ad/Edontq8h9IeLz/RkrXb6TD2FmnYpMwmYCHU/iwpgO9k1SXRlFoQ
L9nvpbpMcRYZytWMK+C0JX4ldBYXK1D4Qhj30gGk2/Yn8Au5GDCt/7AHlsab/HiMRJw08VJYDf1T
+uazsWh/xEuH9QVTaqNC+Bx58kw9Z3SZ2sTrQgG2KqyeYN/yr4/mZq/RdVq5xuDWztjTE09irVmN
5jwZngqAOSio+WYAn/RiLJvnD9SSn1nqN9QpU03LIH7K7P6Uwu3GyeZ9o8srbDXw+Kg4aToqsaCO
MF7JDczmam0tG+IC7b095KYg8r7jijz2rHnmuM2vorfJIvG7dADmPGd6hN/v9PEmVtNg90oCslrX
apTfh1bnnH0dsl9iF+iaHBDOE1sbHnjTcQImCC+Ywo/gYeYBbNPBMChTJbxKiTYPzE+srA1xHg5j
wKbHJgHqYZFL6MN8/wu5eko4zFcnVdhxijze3h9yHeUtbcKgR9ZgDGmh3JNp1qsyOPwkISZXRn5t
DzmjrNA5igR5+iBXiqrrHi1s/dZr/arPiAdRs640EQ3PGHXhCi4Q5WEXbR6nVwwjcvHKbRBOR81A
cwOu0nyYtCSmTzJPMGyt7/aiom9iddTlCLxerDLUTFhVpEnwUVxsX6rOZOSH1ArgsY79wYsHg4A0
dC+q6D2Z2QeBIN+TS/rZH90IL7L2ALe6wRaanhPUmALl5AQKtymJwFH4mZfUQnI28f+ZCi1YNo7y
Xa1X6N9rs5gRe554NaDWg8dSTfeJpHpCMCdh6b8lmHrrWXxn1kU5eRemktyPUZXw5phAmIxaQ6Sq
mc1Qwo95i0/MX+ZtCYKR3lvesgBH7CrNlOUOfU75sOf/2UBTCqV0lxQH6eU0ZdAPo9kbw/mSqpTY
Da0eGymHCSugmu2je6klIs4a8+YD4I/CINE4VNuXttj7m9ZjBN9YsU1AvrQt5RBthW9GWt2oacGV
xaMAmimpc4WgvBqGcJUrSbFva9gT11J+khfMaZ1VN/cmGY+QqKeAHRUL9qVoPY8c8LcN30gBBbkq
zY8vUoPSA63DHtF0VEZvSnViCUzKDimHr0GnkgXyfSWEnh6rENcmc2vFxPuIDKsrRZwbYS4jSXUE
roKQKyS5siENEELb03FgHuaFwJd/bnMMZ98gz+DaQo1PK5deGaV0m8DLSVn8xxF/aVJ2hKNpPviV
CEZ03+iK1JRlT4nHF3NdJUW4l8eM7a/CtfS4yk0LL2mkjC5YFcMNuT1nKyFtK5Nk9u+olhfMHre6
yWKiirm0OW3kGOPLbKxCZ0Q+X9ReW4QkAnLTjQWIsRU3D8gbUF82ejHLzUwsZs6ccu2Xxg2GaDdk
9bjL/jnNcXMi/3UXxtYqLb2iyzmD5wtaHkdOmddfHw35h9PwooFJfRTgBWkuRS9oQLC1+Rg7Bkyu
YibbbCMkGxCXekKsTXYCN4Q5qKBcrrPDuc409XZkOYoNIBPGOyMhTwtsO13IvgPLjB4B91Yy7LCj
DW2mI0qo1Mj7t3mb5k0pUresZDquF4JnrTmUz6qxdpP55BWoCHglPTWsFSeWCsZITNzS91Zw54Jt
fZF3/o8KEO5bGMZV937AAPkl1yvK3PbcNgefs3cgscOPHs1jI39FEZmGEocHCaH0qbKAFRrv6yMP
6CqCTEYw9cX7qAdAgnBLTFtW0pPnqsRM8SrQ4qrsAFd0YslQygQF5TQ5zLlik1Y8QO/hOBXw6qvh
2CHE4EJopB/Dwjji+5fEiBYYs9btVe46uI1xklsbnE/YpGUw+/Md5kleI+cPWpdL8ZumbwlGAWeV
tfMuV5N3bErp3LM7CvGS7LgywVihDdL/r3BCjlN1+M4/yHLsfTJOZeeoGhDuYy8ftuH2EiumpxYi
I77Q1Ehh/euzra2PQqmjFpmDeGjc5LkswUp8BwxqPUn9Il0quBc91Slk3YPXAwhOh4zjSC5ysWvJ
in2VfGBznWAbRBRXmwxZ7l61m1nIN1IeWXHsPnYmH7PRPe6twelQPTXbxzIV45PmqQkLHeUK5211
cYEBc3z4nzO05H/M1j9I8WB3Sje8UjBEdnHtWcWK+JY8lpQ47e1v05razyyuMM/nGGbalUCR05W1
O5JABCG1uEF0qlFbTNdJh+91YSPpOtypb2Z94qmk6IB7eQ4NBd7UO2CZsst5cVi77Z38g9kTsnyZ
e9kOqATOWmEx6ZTekImegwvCvSApuChJ4odeLXk3zXJxF/CGjXgs9Ii74gDwRKd2Q5fApWkJQ/71
j4+wewsGKZ6MbwnRJcCZ5OGWq4HzqB94UQsc5oCxJ9GWzr+uhg4N8o3qxfmTIdX26GlHwX9jJ6Et
l7sMQ59qcElkF6LPM62Hw6hlP1I/Ri2SvWxw2B3P9hPjXVmD3ndpWZH10GS1FYBYMWb+Gl718F5s
gvdoyDLydcyJlfkRpBzJyaA11LNeaTLUkgpqCKzPZhgoHzP+my6a9w92KORSgjmVfZ4AqV2t+F8U
V9dFe7Y69mgZVIxlmwecU9XY8uni1IgD+cxvBJ5zJNRPN8r3fA3pxTgmNpxCKVu08SpGStHzaQnW
23LnS9ne0Wyx4qZI1a2bJe9Bh6VdIG4UCkPTjNFAO/wQ1KkOu5zpV94rCte3IBM3j4fh2IHE4oFQ
fVtufq5L1xBcFSkCm1k0m2ZQ1JLBKeI9f6ukLsyOyW7AZp3dclvp/xWEGALbJUyVLnZhj8VbRPbH
n/WbaGO9Ixhdz1xLaw7Dk1d9YgXgLQ3FPl+Ej+3sCcACF2HiGBh7OqJooO3cJatzr+6ems848848
gEfBa4XLo2swEW7bc8TJpbH4DMVxhF2M8IJM0C9PR92wGJI4e9ll0Hvb/aajNvtKbGuAlsraXbRh
Xckdu9SzxzsPcLeT5iqx9SjNhtKdUNrSGzWatywTilhe8dIwrIpK2+/GVNPzzZDix4D00RTnJ/mz
tcvIZmwuW4RWMYvUR29deYlnfnZC+3B6tH9XvoNA02xDGMqOTAbeNEFfrtqINb40RZ83xk9BrQSB
zgTQhvzswirXK/DX3tved52HBlRbt5MWn6VDvH2kG7LgRR3+G0C+NE2Jf7HzZhRgLQQcASQLvpiZ
BCMGsCZIDg8h96+5NiBpEGmzAzwXOHU2UXKsRgIPqy8p5BP0xQ9urNFCvqsjQSkSHpN2WBXbUUky
A7zCo4gNqkXGuPfqDLmhrLi/23fCWbsVlm7YfGoGZfWkaaJJLZfbjDTyMc5F/Sn+5Hbd0zlzCSa3
lZ3G+iT3tNJLU4RIXQF66x/XDzUtmKHjkgBmtZnK91mnBCtozJDg3Zw4tniKrqlktmBq8UNOBFPn
7hsd3mJDe88zi2miBoRG6zhZCkz+bd76CR3B2L7bWqVbhLx/PpeJzIkRP2Hpzv/Ci/VcaRFqRGET
i/rFsiYY09fFWGOc9e4++dfTK3tseSVUt/155Y5z+gVu/b/ns4jNJCKeTATfsgmxQTl1o8r1NLTC
SBHw02MKdziMEFygKNrEgOLLPQi+D2KTGLsibPDc0suVxRexq5WjRaVRgJUd94XL1zUeLuNKtAnS
xp1+T02JQtaT5HmHhokT2t8z4Y+VbvHwRQ8vbmgGfNL/ZklMUE4O+jjgVavom3GHC7GuJ9z6HJ8Y
FvGnBCa1IRSECfRshcDyHr5dgEid7a6P+bP37CGnh804cu8/zz/6q2DwwSqnycTeDJzqEqSHKSsn
8qcAWzrLH5WsQ/3Pu8Izm9r8Qp41YxtNv4OL+ub93YTdwlfG+s04nkQv8frvRLVFQS5OQmBiAaS4
cYwuDV+X+b7GTQp4+JKQetdj2JOZrK9jVtHD0f7IVSOlhAjl847aoyGBQJlcF5tZmSVAb4Otad1D
X4hGrTYNNECMzuSoYLPLZIi/Y+DCgirLM5MLpppBAwRJZYv1sEtHwQa6B02ILv4OelTfPhdIMbzR
+42C7sbkPMxd4f8biXvAZZUgfcjZvl8Zy71YXIDxM1l6hoiuALhQ1MmDvyGIGa5h4zZ5imXDtw2z
mIkSHhTL5Bp5mo4ZcMlR4BA7BWJEueNSNkIG4x9jpgUldRKOlJE0pBFgzSuLQqSH6odelGyTbTDj
4JTgHiYxXrlzYe9bGyL05hTCD+WohwsrxqsXgrcSRia2VJRgZNXs1nER26lEWfqJXenWz49zWKzm
DVQgdFTRv6CAILa5WmTAl2gLyh45Ee1f8EDbbBXSE/8a7+/PJSzJESd7i5AQzihlCyM84jgNjm+t
bH6eAE5dB4jRnY3EfYUlWcszaSvv64etVF6meotEXeSh8gnKDjiN7keGxAP+mLwfUKoDYc2nVbGD
riied86RU7cbywoP14h1jZ6M3pOw/RR6FuYtmugWKN4WjJrcWBfXtNqcfVry58VWxvINaylOJLSc
YQrxT+COM6DnNPqfi+/7M61Zj8ih7RcxX29+KiPQJMA88QV+UNRp+lyoyCbaZGUrSUj25VvmXLJf
RdON5sRMjMTwnqyU6e+9Vo6RsfgFufU5jx+7i2QFWjJvUTkkH62kaWcCxvr+fUCipCiR2GKjggun
1i1kddEFvbohzrN9aR2uaeVuWEoTnQXNGzBid5Pb9vBjCYVmVzrtvfxZBkDkRRElY67r8yz99ocp
hVwLJpiYBvlG4YrN/Iqg0GlVFDcc8evilQ1GObN4bGruyIgE3BPyON+/RxoFSIVa0Kh3beBf3OyU
CAXJn3s2nPQRhJ7Fgbb3GO7B9mikHBuqSsPil4xAM4SnlBBoaTZo0Ou4Z8TnmgO99/LIUmtd6JLV
Qt0jf00+mJ/pzNX3DivubtcHm6mz8fTDabuMO6WGksB7hk269Kyb0gYXgYdiVHidleuSJzaxec6X
/p22EK9Dv/Lq2bjtJWys1Y3RCMIv6374z377ycehOi2ahfD/XKV7RzAcGpj6ljl0V3G2GMAiXjsN
v78D/Q2IOx0+ZTXqphmLRbh0ZXIt7QTzS3Sz7jeJ6BHEfE1nS/yIrPHLgZJO4+tf5j/G+i0kyvKW
rHvHQPwXaHqlN/WhstNbAu0Zt4uvilc4zmX+XHxZ0R7xTpJEtPb1T0veBNq4hXmOkT+wwZVMevgr
BBzWFLaW7eK4ncKE5jRTVTaeDohGAyGP/tIZNhETk/Ozy30IW9XUQ9lN/Zy6QtcZejyuFkrVbKXW
w3AZe0hMBhkKo74qPRz1rw5Z14SiHM3IZXUUroTz3K3rGwF9Gpld4zLQtoE2/0k/Y94HpTalu/cR
LNsTdU0/Cg/99BBAhrA+0bHYJSu4bwMwHJhJtmQgAYo6LzvAPdytDgMK9ppch841/v5lXtOWPq+k
u7v2dliGZuYMbmwlVm7Fa2Y/9KM0F7rjV53iLksRg9wp/roCozseFv4P9+eE2FQZ/7ONPMmS1bTm
j7j+jkdWcAxNfK6A1eHVDodMhPlr7BziqzBhei35Hz3MfxRrWq6ACBf7FfAiUBqSTXhhEhL0ZzqJ
cMy6KqLKEoKnQW/ao3/XZxdRjSC8alpW4TftNWM8TRdQLNi2OEJUeB16CV7Bqcg9xyU+geV5y3yR
iA7B9RJOEqISNma1Is51mG46nI7zczn5CgNK32s0oJ0JpAqNxs5bW1iz9pYsdEgz7gN6h9ECXVbA
pZbWp/3LNyTbJskyPJCNzFOycOigdAV3qJdQXRUfEtUv8k37/XXurCZF4JxBb11j0FLJT0dDtdLH
cCmZie7wnOcZfZykEOyON65cAcg9kIHwXrjO2w0L3dl7hEeSDUuwj/N/llfqk4ixLUspL7nHWwJ5
y/YLIQs+ZbWdT8P5kMiBQpatT4Lnv+XfbC4+UW5U8pteYyJqiBbji/udwkNINn9sSh97TY1UW71u
paUbZI7bu4FQkDvK3cUWSRb9z1vBjwe0NfLzX1uJ9pAApMEXLvZH/gKhOHcGrfDjpxtfBEgXniOV
4PvvB76wEH3zlZSesCrpM/NoQ6mFGX6jBTEezHyMDaxE7dV5vf1WmzWxAlAkPTg8kp5tWVMuzMQg
wNqmhAlUyLbpw5unxqcE3q+bYYN+HfjX940Wz/C8UiofHmMdysLcn4Uf9t6ZKc5uJQ==
`protect end_protected
