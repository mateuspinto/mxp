XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� Z>� ɟ;� 5%��G�=H�eg�沒n������a�ͬ�+[�
(;1���YK����j�23=�=�BҚ)p b�!��^�#"�1�]�&f�ؓ���m~��4R���)���K���G��Oc��|���ud�����y������HqRԎ���H��K�ED
�{׽�v	<Ұ���N�������ޤi:VF��f����a�mG_~��<��Y:O�ؼ"��������[� L�5���T`�7�&�AӁ�Wՠ���E�0�l�?�Q���q�3-��f�?l|�s���k3�{�����jr�@�[��`�D�	ZU�ȃe��9����3j�s��j{��k�f��v:R9���Ҥz�����<����6�q\�(������u)�o�!��()��6��C�#},����X+�L��h^�K��xV�������+�rt8/cH�G�~��牁N�}�Q�i��+֬�����;p��=m����?O��T��i�ު����l^D�<{GN�GYp��}6��B��E�̨��?����g�F~Pk��p�=���E����0��Q���9�.Ga����Y��������r�*�1�o�����f���˳&*�"Me��8�Ӣ]��>r��C��`�B��_LE��	"�S��.����M��,��G���3�����H7~�^� ����"fh;r���y�;a��ǶぴJ�D�8H��}��ni�(?�i�B|�B�C��[1+���s�XlxVHYEB     400     1f0w:{��L:��2�����\��c-�	+�-;f}�&�F��:`�����(��~��r\�p)��K1���a@�\�ǿN���T��f,U+�����?cnӱ�9�����Ȇ�?����͆nd��>TB�����(B8��g�~y��
	+m�N���*Z�����O.e)��$ȆJq���Y�ԫ_2�]s��[��{Go�0h��,��#Bͮz�+0?�'�5g�f�˽,���,C�X�����8L����0 
������ �LJ���@��4��Bc��b��Kf?��HR:&1���z"� �ݴM��Xs0$</ln"���}z�T-���}��ÅU��c�U:��p����{��L����J�"|�c'���5�wۤ�9}0��l��U%�Uq���@��0���	�@uf����7���9��Ꞽ�����W���{&����N�cu�A��76G�[SR_U���(�K���Ҧ���Ʒ��XlxVHYEB     400     130E����gd�c��/ml�x���$�����c�=�ԗ��u����q_Ж-yƌc,&F+q\Bԁ��&�F�FB}��q�͔�؉�"�QH��y�7����"��mwԅ��5�����6$]���1X�"�̔��L��Oӷ&T.����,�Xqu����2�>43�+B�\�ᝩo(�U(wSp얅��c�])�T�\Ruj�Exy�R 5����̶S�4	
 7"� �t�`{��1M����1����;�4���Le��b�F5�MyX��܆��%�_�N7|�U� ?XlxVHYEB     400     120�_뜢nh����yh9�!|d�&�n�:N�`��*�$�e���%@6��{��R�'��C�m���4ȑ���h�)I>=�%��}"C������}�"�dڐN[
L8e(�۰�j
g஦�e��
�BM�����xڹ���^��S��j7�������;!ԼR��>�y}����b�$���#�R����<5�1k!'2�x4J�$doІ�CB&���0�H��>�&gI�\e!A��|�\�pb�����Hrg{]��Y��y{��'&�V��'��2���`�W����5h,�XlxVHYEB     400     130��II�V�"],Xs��0����3|��C�:��R�]�"��h5����cH�b�AN�����ܐ����	�������(�����y�����xspԪ�3�y͌2P�CY"�&Y�S�w��E6]��Pٮ��#�Ӆ���y�4�f��S}Y6�YB�6g�0��t<��Db�<����3?�W�����P�.i'
A�ԑᩨU��2�,.=?̆0@������@4�L�QD���Ha�:@��
��7x���Sfd���1��ܧS_xʊq��(�w��^�\�2tB�S��7�l%���b&XlxVHYEB     400     140�ZR�ŨvL��M�����O���k�HOa�����6�$烞Ѓ
�֐�l�Xd^*���\�-����=���p}��`�8#%��VKKf��J���	��W`\�V���*�1~�/ҵ�|�z��T�^�=6�,G����J�H_��1Te���bE�D�%)�A�.�^JXq�G"�=��ᾶ@5}0�d2�w`&�+;n4ES�_�B�#�N���������f��w���%9KX�Е�`����?��ۊ�{�3�Ӻ�)�jh��:�$���H��Yv�[���Y�i`�0`�»�hi1,�%[�XlxVHYEB     400     180��G42]e�8�w$��_�%�+�(%��U�w�P�e�(v2�,�>���G��^�5���4��{P�Z*�M�!\����,�눳�\����9�%��?�g��@�����
�,�r����uЊ^�N�SAOuQ��M���Y_�� ����o�z;�����亵{gm�B��}��[b{��9��[_��ڎ�$�ֶ��&�Uk����V��
T��u`t��kU�a�m�}\��S��ڼ1�'�/��غ��������[>p�D�`�&d�"��>9��0�!��)���3J*�[z?B�]]��J�rL+C����^|=d�?2F苋�uX/c�TC�׷/���v�S�;[�1b+|N�R�k�(M0��E!�/.�]TV/5XlxVHYEB     400      f0�j	����h��6�~DO �y����[K�VwD?�ul?�/GX胿�nD'U����>��K��vo�.�����n=���@�"�
�-Ӵ�KK٢5��n�E�V�ai�]k�Aq�x��@�٠ D��]�h�>7z�X�P����PG��(T
�H��U!K��tj��|���!��1 _�焴�{`K�sp�a`�X�ñBe���)��{�[~�P\ƫE��Jb�Ǌ3�#q;����[�sXlxVHYEB     400     150���^�BmH���h*�w��L�&�f���b��2մ,%�uB��Oh�@�܌(qr	�kw��n%�i��u��P��������C�����yl�V6�[�:Yjy�Z��Rq���$I�����Te���m�K:� oіU4�&�"��;�Mp�����F�e�?��L���+q��9,-*3�mJ�KLn��,�#�wq�����*��y�=�W>���<u���i�Akn|�I��4w�3P��m��Xf;�Є���`9pڷ�TL�'s'�f! Ox�ʍP���3}oXw�.W��_̂��kT���l���ӇK*K��:]]�Ԏ [���˘)�weXlxVHYEB      b5      70�� ��Tc���R|�Iq3��D��p�j���G��䟰����=#2Y�lB��)\���_��c K������S:���@*�[�����:����܊��2�|��