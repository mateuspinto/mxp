`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
xQho9hpoS6LUpIHEXhyA+Gf1fv0W1GYPBAf9Q1YORXId3qSysj1+iWBZajc69CttRgXIET9H0agO
pugkicu7FLIxu6hzZq2F19aEJ1/H9rqWKsqXVUwv8V44MCtLCpBC6BDizwW8UYd4uOfBPJur70vm
TFLfWvhmaUOPdSlzRS8qrGHmN/vPj5lvWXJ2u/DJ9MPxjSJXBKzH0Miz2YRxLGj2cUi/zINWhTh9
yq5X5ftGvSsjeYMrlDlPTsMaEl6ZyYR9n1fLpW2F4u8bpwN2OC7/yap1Wpmpb43oa8/i7ddu/ZDr
BW92EMCDyH9xHY39FoqF6d3iehmbksPdHoPmG+d7GxRdpmqhigQjMF5sjzm3VkDsF/01vkVWruYu
uvwR0a2jAIe9gHmq9KiBR+qspA51c/1gm/sGzD24NDLZ/EFX4I2PX7sj5DhCwF9MA9sMp9FT6l3r
/h6Zv8XcGDgHdE1XQ8twuT4oW3u+U0EC54r2tKGqnGMeJGpf5s/FGBCFjFcJ/TDJHibwQYJmm0KM
GzXPY9dqdipqoHGBkBWsv0xRTRIJFpZqHCXZG5mSBbdn3yaXybcLpZ4iuAf1dPDZpEcq2906Q6F5
lM14CsSGLBoKgtxchcalhBPCXTPNaTshbvyMLH2MjKX6m3POmw+sfZaTn2wGBxHNZbqVqLnZIywz
IY+gEINFuQ2TXPu9X4cf3npNs2kHf+PZIuxrdMEyUJC3DzUewPJVXKBP4S7Z8nLvi9I4AJhcohnG
DyLX9H1x0tWuzGCg/fLEEWgvI6n+XZ8nET9jGc019MUB/nSNFkFxL6lnv33HrfkHuEpvF4C/pJrK
M5QCtoRKEOyBWRinsqNv9NSQ10KciXQAXcbfQ9G1HfXYnWKRXugXjDbLiJ7uPJWl/XxqQWk5P6zf
inl8M/ol6IRW/Axw6RA2Gqv4/Bg5j3Kn8jGQz/KpC0NCc+2W5WYdQHWzKvsBIpoj1xCDaRJzssTi
ve6AMiYrOxsMkf+2CnP4Ls5KZYQRCXWnU9c9yrTGc911LK62Gog71WT/avnksY49aYKOyTKW9GAq
DF78mZXXbFX9O/UmqnAL/WFVsGH/zkalxoBwnwjKxvOL/vAfQ+WH4iVQ4NkRKwFnK3emAEtLcnIR
0sEJGAiMW6HdaQqKq3zl8lgAeTnaLtjR0PsynfBFDCNwvyJpQWPBBqzlIHh7Y0jgyqhbgA3oSzHt
bSLRf/UND8oBycBKcDyYqvSGbA8a1lOsFRjtkY/zCWXIT/Pkxnu3H4MgoMhzRV3tpmopiB7avBuE
OVBBGFDgPDSArrb8SnYofE3EerakancQQEr+mW79Gty7VTcu4/7Rs3LG8SO1YLcTbPUig+itsumQ
zMXUBvnc30RO/OCPuHJSS3u/z0STMeJTyeBOb1br1JTnFAW1cdnH17u1NRzd17zCt0kSL6cWB4LS
mWOioyNQUl5cwm1llqY3hPAJ+KBE/wxl3e2/a0UnID8QKRRfxkLxHqW9n6DPamzNQypQ9UtxNTKT
7LbnHOTt2BvVMkE9JXWxmUoKBm9q/b0AYlVp2fhjprRfh0+DOvDxDRDJ98ElBISMZneFJ6GFoP01
RBsibITf6g45vP1zFSOgJjK88t35dbYULh/sN2LQCFTHEfWtHsX0ff3cIWjC2VtYEHdaAzoGjLYd
QwTys63g+SpvRdMBsMNeDXvI2EyjAL/NwdT97iWfVrZLQ0v0nV+wgqb4L4i/Epc1Qc/Cv3FmhXNi
e6TKPKRhBTt04rix+p5/lstevGWSpotrA4BgBQr4Qyhnd0NdmAFJZbuRxXtwQKUydinBD8Z3jENQ
q+CNn7OUf0coKwu55H3pY5kTDW6HQ5Pg7s5wOe07xA+pWnOqjEPzVBbcQCbYUm/hlrUD1ZGkxCyR
TOG1+X7j7Zzy22j/oGmnF5brc5Bf835ntgEiirhgHRMNdSMaj1lgmttDQQNnlkqDgIGxR1nfw9kC
5UPfhd07PTQMUVc15zLQk6knUc1m5ZIuOQ61Nrq2UE9GP+TdqmZRQbPbSgBn04DBM9lEsIwcqJ0B
Xp6Cq7UnmBM8PW7y6jXhshtsZ1tgt21XLxn1LFyHW98kRggCH01cvY3IRxdY6PgXypGGx66fkMSV
Z9kflnFsH1IwRlypGFa18DbZvt7U4i7uCqGi09A6LuIszlbTPGHBlTcqFjR+PMqokD18qJJxKFZy
f4nxxsHgBjJ2+PfeqGZS7ohgsIcWgi2fLgotg4xPCkCSwABX9w6BXkNzd9kug7swbAWRGQtO7k7i
d4vYJaTE92s/v0UeOVkW8GbyrRE4RDDrqUa02T09KDenvgXf0Kvb9vY3U2b1j3v0ns0Y0/NzdmD9
IUPKbEJUnd+VQ2CHl2RnQTmrYWyqc6MMXNfl+OTcOqzXSGCW5JeDCT7Re8Cu0rDYlfP4V7qgefZD
BpLoldM5Qo37aHXU7nLUMYKLeztWFwJZjnN7Ci9/0+GS8iyqSvfHn81CkFucHpZ9cgmGUs8Ic8PN
NjwhtjQVre6OHpIYvpbzgTjmg8PWqN96KCLmQEDncggO9nEId/zoEX7b36cv6Q0cpGGiAhRrtkdb
jPKGsxfltcTLocrgwi/HULTLuBsiILkR1fvZbw+/jL45wxzllviOovQFU8WZfJnFCayuao3yfw9E
L2RMfBmUxT0UEjr0qdDIM51YgY0afsPw942x3rzO0iO4s5+Qs1tKIBWgVF0Mnbeo10PpqeHTIWbO
cWeVtWnfaed0aC2BSPg8cQq1ZAjACxxOC5sBM7cYAHpQzMP5ZcjIp/ScVNHGpmL9ioJDik3rj6ix
U6KDCWZ3pIdsS83rs83jQjlDpLkPoLA/YWkNzXkzJWOp7Zy+Jwg5QaoVhOuFOTETzhXgc6A6R+tR
DeLyCDTS3HdASXYMkm5BZQe1BrznxpRY4Lxy8VkoQfBap3SzLUT2oYIfZIqrnF0xtR9jpf828NxL
CO7K658swkTZvjmZAnWoWuwSCRphW4s6q79TT56tO32YOi4m+yXnUZlfB6qIntdnDf0THIXTKNQX
rOj+zj/k+ZP3+Kd+ioHw9F5UeFOIwV9v57u+zdeDauQTqsf5uhuf1BY09znDnsGfJxYm43qaHpeA
7MdNsTCUF7AVIuB46HiEYAdAo8QmBuizo2RsVov74VT+GABpYTEI+dTBQ0MBO2x4D3BWN1JXKxWB
SrcM3GnmjMIMtr1zRtKu8DZIhajx/+RpH09zOXWsECG6e8ORyvgxmiJ0KTtnw9mA01rBdoD+duIS
fYMiZJT0ChcoCFvKrSVpm5VuwRwOcYQPyEC4H0DCRZpZKrPYVxmyj5EIaYkMsAxdz6yLkR5vuT9p
+oCVgxZ49zapCht4BWLaTn3OMRYhTO1mdOhbcyMCcltOemSinOVs/h5w5H50YiKBjzfYZeO99fMz
dAbxW62WlaI/nvBzkIW4YCmYeBH7d6an1eNoqWBzff5PdiyhGXrgYm1FqBZB92F+ibE/EPBuMtnJ
gRq/5iglc9o7G3F9JFK08XY+Mdng5Vil5ldkHpInjM0sZtZaxydj09dJeBZFF/RJcUsWvan5zE0G
1Uc89o+HkVuxCHOiYi9OwXtjq5Uz4gnTha1ue+KrRTf2+tlELkAYyiz9OPIzoGumpwSZ+aKo/DMX
ts9XRin08RzdohEZvz0IkZlp8yzLVtnByCLLnv4WhvbyIGiLSDswifwhBxK24o/6I0tSmFzJP6oV
rfZOfnHrguZUqTpx3AQma0sLcQv7psW2yYhJ39Tel7W2lthhYaxkNimmzAsvb6ZIDN5yBYCazx8n
R8xCi6EhlGEQBFuZArrFUIDoyL+1YhpG7iTKgZ1mvrxaPqc9FWrN+J2pizS2ZdqGKcF2Az11jqCv
hLBatvzntYzSMZJ7MUEiiU4d2hCIIyUBeL43QXyj0XPZKsIJeAjQ/J32QeV6r5pGCuSP4M5tCuJc
iNCr/PPkgl06S2T+9Z6F+n8Y3u9IyPwAbqOFX0vG3hRNVkBJ9Bqgkt51+Uthr59yt6cWGda+Tl7Q
G3BOsVWmGb6aX4AaFnQXsuCp0oYdXgIqDOKPCGI3lT8lcqlru1bLR2jOREVIW9Bnb0F3qEcVqNKM
fVPW3GWyxsxREw24CZv9Uo3x0+1XyfVUn6hPKvL1m09SZfZfuIScWOgD2T87fyyxxxt09n/jwud4
YIl13qpUO6CT+RLG26jFGSm3e1xZDbzRhkpdhTkfT2qOAXtk0JSrb5HmskuLf8MoSyW+MiOarQEc
n8AdymiUPAwbuDAUB8WIR4wh+vBhOf7HAPJnZyC5pHN6xxbRhhFMdhfIOOWdaPZ7vh9Gzxx9SHmF
lllEi/Hy4yy5YLkAbn0Q2dtyQNw8O+GsU9yBIxic7i7EZDO/6jOtEVSXiFpF2paZ7WwSrJBuRfOY
BL1MEQ5dYQZk9WUb/xjNQCgAeZ2MwnLf+JT0SPsGehuhvOIJ5+VseDmlmGh6SoT/IMU4fiUe+WFV
ETpAp6ep2KLSPZhJanejyKZyrzxXAjnCwNi5l0ljcosFhfb26J3FnIFuP0UTKf3L97ny63AklIDm
t1Je1FmAimUm1FJ6CEISs7SDZ05T96+NQ36TiqA0pfNBKjOR3I/7nGSFX7mbDzQWe5ThiypPhkKn
sxjRyzMm9MZkpCvG/mLoZKoma1kDCYXhTTA35czo5+WDrpbqGOgJyfXhsWeo5+0bcUTIGHvSfM/q
Q6XYR0yxIkxnCVvPS2+eLeoIbztAyagGev6cNizJRcuPHRoi1/Sk8qibCHsS1Iwk+ZLi0I3ixb/p
/d6GKpJx0jrGSqpwTN213JLAUhBCtQkxoTFHqrQaYJg5dc9KmHVx0My4YjGj0MF70w3ZmKJORLNj
VtRyGoBht+TptxkyBD1P6+etGClzWDGzVj4omJEYH6MUCO4LnDwpazLOOI/fLBwnVjS0rcSa1eBY
5G/x28mFLwQkgZbUPsmlN4wZi07nrK9/1Udv7ZxnlAWH5Ze8cBL6MsUCJA2vLC5oBGLoP9yLWQQ2
H5z73p/9wrgfJJNUETrWT8DLZQ11nn6b+buORRHwYH1SZDNhefMIs23xxBSkCdvveg+BcjBnUBDf
pmiQSC9kaac9vxdSTX3IBg5hObaqVKAXktYY5r7gjdU4SEH+bNyYXtm7QA441I1PDbvXI3jey6l+
BqJo/4zCV1nmof6CIqH8qTQNdDcBJU0N3AAz8J4pW6MeS16AjDDFeRahaU7hMEM8FbwXKEBGkMQy
aKcGsyuQsbASQp+RnODLxVOZK+3XOJMD4pjc344NzDe8/1fmMDdBLNL41sVeXVYg7x13cyZk2w1Q
MiAH49S+cPA+ni2cXlBvdBsulZVpPx6oC5mQAz5RIxWaQK+0ba3mz/kqaD+r6izvOz/L/+O/nDEJ
1jti8UyPBG6j4wjBRfTYssTd1v3PNxJix5zcZYrW6VGRUSqfx6HU7XXagTavkqm0tGXG22vI5tgQ
FFLVIrcsWAIdJfNL7xkaS+rSUVAd3VXdS1H/5EFZRjBEFRrYDdu+PaadmHxsxy5dw02mEtaTDmVZ
u8J/UKAs0cDZL/4caRuBEim1qOC8XZ0eHpI0LaBVT8sjbkMXsPAkRUiaHBip8LAnJktvfF18v/Ny
kRBpEM40+LQap0suyP+TEM8gG9sZuljaj1VhU8w4t+7pb2uIslvGiQ3qZQXy6YrVlByWBpYGx/O9
oJKSaN8US+5p+F2fyhrnr+SiJLcM3MqmBWrc5SRLgDzgVBhbSlwimddgi381MF7bLi+HmlZ3IArD
yJE2kwFKUXbs0vc75NysoB2uqNS8F7o89j86NBtVL1uggFlrVWLU3OGPIABIUAqSh0XLtDciQsGv
onz3C7eecKpfq8kyLqroJpbLbe+MN8KSdBGXZazCQayCGQdA+9xHNoNRL0DHJUgsXYD4YUj41pqh
1QbOb54vg1Eb0e7gDaqPrWgv9UCwQtmlAf63vaDjQoT2q2IZf/aw4sXK/gdYtTKEL5PzYU/tLamh
DJw6DSa0UTX1gZO49gskqPIdcrQKoFS3oO7SwxG2+mmtAvKERz3CHf9CSuOdS9hD3X8lKwKgJFKy
QI02WINaFkGI11gRafs+Ush8wwpZOjnffJ6Ic4HgDGNv6/Mew4bY/aXZDTF1436qmDIgzX0bFkdG
oXousxjhckU9M1KjQuoCD95B9/f4gHD/TtdgSs6Ug9A2+dZiZuKOVD65ZJcgnyhaOJFehSaWC7x8
H0mlOYc3kH0NGLZYv+ju+poVdEn0QUiR4pVvcxP6OOq3UvZ3DZEa21pYH/I5WqA09rZEH9Q6hD6F
LqYV/b1ZIKNxEMVbFbmjeL9ljljPu9XumwJBNR3fFqNnAOFTrGYPgu8GDFkc4NgZOPRMP5YVbLsv
2vlsDsfQjEy9UcF3BJbqR4UlcR1aKn1DM3beWOn7M/GDC82LhT8qbu5v+GtnPhWce5tqDpz+kkio
o+L5tvzD2gmM4KMY9GFbGns/vAdg9PCM9960i805xRqzxfXm8wsUNc9q7lUymBAloxwJTiufgSPZ
sHzkmUDceNvK65Y5mHdjdqlmcr5OAMHMqEN5QSsA4/d/NuLv/xwZhtfZBtUhPaRBRnlBsF+0LT9n
8lO8oLA6s7z9BRH17VpTcwo2Q5J7KVSfu5JNlxVjH2FoW+8WgNcz2XtP5QnH4Uu1YVHClFI0jw4B
WtgXCqDKfnwPizXDRsjjl4wPsAtrTR7V+Z0HKDsYIfO3iSnNBWwv77Y6Bm2OvdYguz1QMYmhkWrc
WteJOup3yBVa+dldWlbuuuWqmZET/L+WYG1OjVWDCL5HyKZHpUVw4Abzmr5Vlbe/4iBXqvgAYLOd
RdvFI93Hpgeqbp4/GJoPFXbeQFR+SXd3m24zLzR/sgY0YwtzldJ24eBedM1L02fZAgrgcAFFUR78
RM6OCVIidS59M1fNcbMSRsLG9h+U+s3wYQXV9oiNQ/01D93it/ef2QLf3d+IOhdJshKgWrwGYHe9
udnXLOfMU+d1s4kl5vwAACGdRR+GFd4mLP6cvSHUWVvbWjEaT6c36yyOHsx/n52MMF0eO0ViUgj2
OZRYY/9DHDUcGz0v26vXNSxz8yVTW9wXeLceR9p2ze2/E4YiFukhF/q/7QgsdNcWg/oW85gfwvRv
G7QyDG5Om2bzmRRpZjU4dSziV3dmyfnwS78x9gFBO9Q/tzIO+x2ehS2+bDERx+RFBAy7KAunBF54
1LCUNJdUf1tCSdzMukKkWBSrLG4INN/7KxekSSMaHyMDcX5WzH0I41i3ILT8WaFQz7zDP+gpYwgT
a76JGejBrS4kZ27W8d8QlM5W6B/3xbiRTycVksLfjLycVxGGWiB/HJfdPyLpT665MeI4s1vvwt+b
2jnnp4+kz5Mx41B6+pLsMNoM4yNjhnW8ZNIig8W6IxR+Qz5fHsa2C/KHASnZ3+5VueAlv62/Ktkq
55T3/ZQPjVsnt5jyoY8+wwFHevaa3dmB+zTxLi/NVUHrKJjIdQEX5YfgjWidkaMu8etAW30nkXS4
6oIuJTQKe5DtUqaXR1eKRE91D4gka3zSIbnge+Vba5w/vJO8FLqVxWamx3CmlDaP81y/bBwA7EDP
b1JT05f1gLArBj4mNps1KkKfaMfGDShOPRCMUA0tQn87oniRChvtqE/tUdSXZfIZv41E2pBdxKMb
W/mZNcnUVoPhI4CYDUPxnivzkTQp1HjdcrSgYa0xhq6xqMHEPci4W4uzDQ/SLOaF/k8FUBi7Rw/z
jZnaWi5ZIQIi2GW4HKSwTLA+mzdgJH4d7J33Pc9OTIn+r0bkgjozKRovY/CsTwFtlJCMXckj6zGE
XvYsn5dh5aq1oWjkl3yUs8F0fDGqDXFFxerYrftiaOeCu9ZK2FmIQ52F6a15hs3MOnxK1+YxGyjV
mCo/MMHpQ4X1THSbqIOjyRvoffdlnrv7W4kLL7doCzvelK2qmUtu/eNUMgQl2FyDF8v5VeNXN6HV
cSKnPSwgdYU6ssuuWuTyfE5vcJZqIfN8cQ8bAB52wnppweHYgHkprVIqvXE8JCIec8gWZSbJ2zAS
WUJLk0iHC7LBA/yecW8Ex9k0OY4sU43RhWJ8IiC+1ZVW3WRmcph1dyBofm8msxiy9FQ7WbWRQ9fv
CvtpuMAxAAOGanymLf3hxOHeONkzS+bvWzFAL2qnAVT6lv14bYobWS4Xk1R13D2azmHfd8imUOPZ
3BzFBYmwoDN8OuVhKV0nIrwMAUyrqlTbJG6lfaFf0Fhnmxvoolor+KP1m2APFmhuUkiSlcpMSzkr
qjnwPBc19vYPhd3Y1Tz1+yKkxqI2Zl+l40+ze8bZLFN06g0Sm4TPHxTrRPLGMiV6cnAhWFVytLk6
5oiahWFtMM8M/l2OTUqIaZDDiAZ+14OyFWhyhTJoaygX1URvSZg3n5jvbShk4AdvPLJNxQX9/D1J
PSMO+1daIrhlWxLb7RIOOMefsq/je7xcPFq1Dh7rvRDaEabWju9yXpQ6O5znU4dV8eVSbdfVY24b
BrovU4TcjpbZcooyErAvsPDyE5jdA/OJKz0jsfZ12csAbSiHQO03wWx0FgpTyPhoFqpCYm1y4UQ/
rOyW9ckhnlMPlx2yIkvEZhyQ7jTgTfsTr4/fZlHmaDq7R8VXSLY04btRNwuL1RJt1R0EFbZwoQt2
iqK1YSFFKyF8b0+FI9YefIuJ17KTm/OXwd3/uuDMOxsUV8RTGTcBTpn8d8mTDTIZejIbN/GdXa3a
eSw4jEHMm7bVVIhNaHR7KLDuQC/NNUcKWrdVLEaUHphVOW1F7I7hpodKVL3wUMjB/TZ7u7Mdpl1a
MwJUJXCi91iYMzKGM1krT4lBgrCUTXzvwhlEfcHiErzITsbepiaN1CENig93dnHfLkY1UyGvYnSJ
qQm58Fj5Nr64T57td912kNXXf9AzVmvTEXvnFEvh2HFrTS4EBEoNT2F8AgKcA5pXwpnvGX/q1zvt
XMCaUAS4TjOEpgEppoxKxFdkLK+rSP/q3CR/bZHml3Xzq8XZScbNFFZMHuwTS9S/nW5Ywk3t0JjV
GzWmF1UuQ3AVq7R9Pt7n3faMGCPAfIaOz8YuYyRkaHhN8ncQJxZxmnTpG3zkN9SkzqlqB2YwI0S1
2xQPRT4qh4oqDwyS15mpu7kwiVqdGQ7CyuR+zYQpKQyYOHpLFmxXOy609d/tKwG1tKdg4KNpvURv
IsZ7iV7SxrPcidaTgtRzmzxevDhyNivW6onJdH3Lnkw9dhe1UXmDevUcXPIpL0fg2tQjo+SOtVAI
gaE6KYUh5Sj97RC6vLXMHu61YNnv/Z0xf5mxRlOBd1BE70dT0GmJLuYdEFCpFQpRm19feldz74EF
7R24dpq6yBgq9Z0XqUk6u+FGfnciEzWAnNyf76qTydLTHbuDTbjsUDcqPCCtQiJe11at3/5vCmIX
6O2DULteTPSZQPLgvROA5tMKJSWCypAID0OY6qheAVsj5iim9ygURddf1Qslmn9bcacV64ocgk9x
wNiSusuaIo6uGV7kqRqUMiVYrAs347e6FJMKBH4pNN8GxgFADcpo0NOu7KWF2V7jVu9KwNEtq//H
sIPUOIk+4vSVRG2kibNHiM9ukmlIl1HIxeW2AfjgBoIQ38Htd5OA//lv5RIiI+HrDU0oJEKGlywh
u1wK0r42hJz4XMVZw4uRuJoPnLuI/jJBZaUWSNucBcEgJVQmGyO0V3+DtWSOy3IYxniH3uDSX/sf
rwVVbSngTG7kCYrq71gSK/zLE0s3Hs/eU9/kDuithicXzuYYt/UbbJAmKTbxbBmv+Izzu2rC3vM0
nUIJa2Cbs8ywgi5ZWdBFXxY5xnO+7msMYMDVCaUQp5yn39SPyu9MHXHqoNQzddljyT192ueLjKwO
tZ+mAzW9cKr8oqpDUy/fbee6SVs/Q3fSApp/lgKWFAeHX7uxdCH7Z7gpkWwD9M4S42WuHHWO7ehi
tKZg0+H6UdoSyAOYoPFx2/AHWR4ouRJ1A/UtYExHapywsanXR0Ux3u+KvVUf0nGtRAqm7/DDbVWX
EuqhsEKWkgbTnAKwKLNTQ+RaG/z6JNlw1wLx3nyOkSEfAs7Qsbs+0Hc3RQoRAUJ14owYbczI8fPH
IOfP6/Fybf/0nx9v4YK2jgW/wyt/UQ1QMQc4sRwG16glSPqhxhj3aKIPVtYn3tA7QnQXtrHPoSqm
AsG74LWpTI7aPGhhq0cKcj1Pr/e8szg+CoU1jVmqdO0S3+Aq7+kC9PtsltBDIqeOEx7WR3ZXYt8E
gdHOJ+9aJkkAbCucHOSvgl4/L7WX0jPXXSmDcV47KjSADuAj9HbpxApXIgeAtf3oxQHl57tY5FWn
K0L59dSFi8EU0y2i7F7azw+8nwCSweuOnRa4e+BwxrHSkpydE99xvjNqo9NsBL+KmYsEOIAOYRll
GaHQky37xAenh17b1PnGvNueFFmUX2XOxO72oLCLU7oUtUBwEqEJY75LJGiMlqgkP0Jx9S+DPMlU
HiFZn6cpqjRClIrrlyhNSstBBD9h2D39/fXnY+j+9zZk7OujtYbn1Sb5O6t7ak0kgt8laLJStctL
zJJKY9VLQ2mVyNKQT5FP9pvaLVRX7rlzyKtmRssPQ76nab4hq4JtKCO2vZx0fz7S94zPiBLePFvo
aFe1vSs0RmuTApmRdKC+GdG5/iqAtM7TKS9qjiHw/HNxiHIg9302KIVSCGasr3S9nnRGCrTUugIM
PNgVOWDGOwBlNDfwyf8ioenfG16eaDeysEZGrymN5ZbLcPlid+JKbvqtUySn8WffiBjhaY/EzbCk
/MllLaw/M1QbNAneBPzha+nYeqU+Amfy6X+fwK+hyjtjthK43xf74lBBy84ylAujCXwceZ+i+G+C
VShRwwU472CYq4xxm7CNRUMI7D8dSnZIWmxUvJlcF5nFd0iZrgZtiqE4Gbyx1YOWY+hu0kb94IHd
O1BIx6ZPwUPMO41BhOithMDzwk2zxXpFE5bX+sgRYhKQmZP4v+fjCWAncUZ3ESwA/2x6l8N7Bnha
0Mk0BRAE9a2yPZaAwbzW3h0Z/dJCW8j+ADj2l49hJ2H62igHtLlZ7nhcqA6nEKQQgxhSuCcMJVQj
F71yaIKUNFfQUg9xrG11RAUw9C0anfx1xftVNgsl3I/ZAK4ozoCSQGZZdWJ4gJctfxB4uxlX5knO
11+qDdMMpsmNTyjx9zN2wwgH5jIEVDJHZImR7V8sHHwrHm6pXbNUSE4yqQ5S7O151nxf5fycYHaw
hZBTgzsth0FE7jYrrQ6OIdSewtP2OmZsTiQuCyXAhKn3AnjQQwP0YS6ilpAqXiMCcVaf26vYat2q
nvqbFvY9E1vKEEoTdUEPR2HliF8qxffbkaCS7sLlwF1UUf9WooYQh/x8WoD+l+PCllDkkBwLKTeY
iuuUQ6iR57D0J37G72vYpmMMdIhU371MntTO8mmCXLJ7IbkuyWlr3TwYMP7J3AmfyleN45UZv1kH
hJVBCzsKGrRxBxPp+Z9VtuQRZi8hB2vs/uNc8e/PDLUjcv+0ZyNC4ipLUiyKjYHA5UGJG1vE0CIn
bIjWCbQitOAXq79U9OyhuWGTtyooJ48A+5QmHkLG4Ty0NI8bDS46l6uCU046PewL2dp0h5WORIYf
QvNFWLcvELc5LAK/pt+3SDQ7gVPbavetS9B/3ePgDUe53VRYM9H/sn9wYu+UQA5JGiKAxzXBHPp/
ESNx5WFgjf4hWF5GIu1jgMxm4iKHQwWF6cld4o/11koGOkgtOwHioJ6A1yRQn8Y9wHWND4lKH+LB
Yr4IgnxetttM7QFdpyM3owW/uqDJhNdCoKLb841Y5QB7XffJZlBEnSH3OxpYHwoBXNzcDVesqSf6
2cTnL5/J+U2vrUuEm49RXqmZcSo9JS7gUkbrC0aR5ka2ITKKnHlWqntOI+pvfX209jJSjlahkYVN
yOQgM7ARzI4HEmBuG06aCIYJKBft6wfW6rROXbDJhfWlQWUH30ZS7HtAOq7RQBEltg/+HlXltmp9
cpAD1Vp9yY/IrJFgmnc4wLjx6K/WqMW29ukxGeYXPnOS2QaT2vBWNLo+kImN/5KPwdsilGLZULuk
gl6TnlDOn3HeMzbxQfaDI9mx6m1hT8aLd8FirQbPrsXDmSs7fQODnPietS0cemNTSnDp8/f5rD3N
5B6og2nTUAuPVDR22Pc/GctoBpEF+9T1+fgA6LLIbmVOkhWkTgaYzDWxBTnwGGqrfb4i6OqggNzT
ySFam4t5wAu5RJmTHw6hgji6fyAYbwNSD2yf9NN66rtz8LDXK146OGtKkCHdRbshUYw/vwi2Qu4t
9972acbwy7M6eXicAtNTOljoofYYF2u9itzuQWbELX3tbrjSSW5IR408d6MKhFhD+eL7iGeiSkKJ
xud1gXhfmROMMYVkqY9gYC30S/HWAOsvozNkb5QVO7wYHH6NZtDlE/yEcqOogArWbiXc3AT/gIt/
wnkXMR+rDrGewJ1AjtlJIEQKK9kJrl8wNEWtRaHJ8PkNum22PlQ0VoRHRr1CKSvvMdyKmF8d3MaA
o+YnOp7pB3XoVPuQFEQuRhEccJhZFf1pbXOYOanFiXfwXi4zWC/1leYY0AjMMm12RTdvVnSGWBFe
oJsrvBMzQJhdFXmC00SD+Xk2/9+qVSnDswKTMAiO5N1BmyFi11x3YutFJXWSIJOa00EoHdS47J6H
odXKaOe1dCoPJCa+KEX3YqcBVfCV1vNtxntwxEGQoFJpGf0gLlMiaXnajszjeiSWbQxBzYdFfFgi
zCpigFsZ9j6viR7rfh4c6xV+xCJ1Ph94uoNmw08JX0hVDdAVdqIQEOMY1BB7JxHMDXe/fNfNi3tH
wbdHpscJmjxMNX2tfnL/ue1m2Zwc/50/gjMlKBWcagHboJaN1KYWzBI429QdpajHaxJX4cavnOn+
l1vSlz26XocRClP2MeEVi+wndh+YyQzae8NqUZP3uOjupbHyZ3H3FbT+g9C+C3x+zhC0s6xrDVMj
vxCbeXwF6MfJYiuSk7OLk8oPOuScDBVahREnZcb4xuPJNQTSquxiW/oS0rVPthfmgiWgW3W20yWa
rQQRuIDQDN3AZ6qEZdHG1ugpMimrVCarM4AO5lbumLt17rJF5JLnW1IhGV2wPZEB2zw56ZTToiYx
GqCM0cR7Vym08tGywEQQNWmobafRHcU3taY7W6kOD0FxNjx0jtXQBpA8TvzuE9QqIHOqTpskYYVj
tyeScebt29yjL3Rq9i6wiIkQV67pHKegUgV21IEMyLulQQqdnzZNT1CwEmcePH6WfbZAmEnu3d9/
LrAbA2RS72VuHK2P2KGzv/LEkmZbE6CN96lJ6zFhlc8e+FzoCjJLzDZJsghUdOTPw4Jjxh0x/ZgT
/f2IPPZikJTMuuiux0ddiAjsxVDYjZ5uR/aBPBXTEu3I931DHidNIjraqvrt4d/S0Y1XsLQB1BLq
JheYHdlQvmvFO4OODODA65hkcAzSxfbagOpQZQhtYOB7Hfk3cTYIB7eyrtzEQkGXsJShCScgBnSB
PEQDzjJmYcKaOfJjz4qNHrek1c9AqdhroHufB8ZfxqZSIkjZ37WyejsT9JrAjdVdsB0l6+GXNtfd
hb9j6oask3TthpMHxr/PLfn92Zh7zzYXlvF+Gvo6GOPCbyngCQ83cpFECeiEXSl8uaadmUKGuHLg
O8imkQy6IFLvREx+b3ZO39pDrOB6GeIQy665xTcfuDQLYkLan9zvA14krgZi1dnX3R421sVqEgT8
MaTsJCmqPzmyKSRZOyN75vIAfLArc/b68PphHsfWp5ZLJGm0PvHoSGIpAXfbiAMQdvdySTiWJrvU
Ty+nlSTE+LJ6NdcdnvacJfCruudMR2tNes19jTZJpCf9wU7UEeAyOcvfuG6Z//PzYdXNMS0h3ZDO
pXSPzNvuh5diuiNVpYKkeEJxJ3N8LopHRKW6G9KDh5Q9Z0u80X9C4JGaFjA6OUhcUR0KGwEKzj0A
wbA3RhPWdA8e037/zNSid+GhI7a+GnMr6jQK5wv3Fw+SWB0z7lJauh6wM3Y9V0tD4aku8NJklTrt
4oH5Kn6iSon/t5j0L0LGHL5sQkrVN51pGFX01xH22T05lFqS/Ju+REhr3MkBkaazzpO2nKsV/Xse
BWsanrJuTe6aGgvHs1A2/sIQ0TJU/W1EMBlCrpOs+4o8C3grg/Rp9U4KcTv6H5KOrvIADLtfEtEm
hhcnZ2YmBxAuPHkA1TL1vlSnqEzyBQJAd3BXRGwz0Zd+9afW5Z2DKYbAF49LTSuahIT/GPCKDGwc
D0Yp3BJXZ8YkpT4Wrm4cxqYoCyvRjfUR7YhGpgJgERTptTzBYCZypLHtjsrdfGOovL2YznsQ0VG/
LHyS6D+dWrkSvn5EY54UCuQdZL9DzDEvWKdV3p0s72jeW8OC2vi/FUXPa0ojHY11qv8F0W4C3BCC
ezdxQjyUXi4/kS/Wywni37PBirouS/2N3S2tEBgAZ4O6hM+/d4+l/RANxJClrIAoAEmtaqyXJVMK
xTmUz+WZj5nwBDn2MxETtANm2yQgZjdFY2D9l8AZBm+MDoPxM4UHbTXMYdh7dSXgI3vUZ05qtVs2
HUKRke+qawLiFmEPppp1IpZzywJonKqGjWroZm6MSSkbTQxd1yw9scCUVV9HetZGzbwMJtq7xNek
IpiLhJhHA8AqghWiQjaHGP5Ff5+ZFyEwwNRwvimjlixlEPgZDetUzO1ES+XFL1f9h7bfug3Syh9o
qqsDBUz8T2zHyir++kKdbpg4GNoY9Gardhew3w1UrdmjiO5uoU2kRlSBQ1FUaPqiAL+X61h2hZB9
v851x2SxzeYPYi0Genkbx83UyA51wyhAKITgeFgww9j7mjw/dQL8a2l1jwcQMgP33L4BojXQrD5p
iBDvHsTi2uB3YX/3A39O32ZN09acGYWGbQ0IFiIxCufd4BGuJYFfQ5lh96E1u1w4KCf/v8RoQwV2
ei01vMAVf8ABMT7MUFuMEPYDLFKT2tfLWqaCFgdwiLW+Lq/2jhkJTN+7mAmsaanWiWiaO1nD04Um
+irgGZSXBT0h86xV5qk2bZkL8cqPxXrchJt8DSJ4y6GygWXE0wQpXz1Q3I23g6ITgh0m0K78KKva
rJCJ3E/KtmlCtbh8RJ0ex0lpUyAxR9r63c8pdueHruwCTcHFWJMJL5VgV5jTuU+7HxfmH5y9v+OI
SnvrKvcLtA5sizVilliEL2eTp5cmizChQFTvWu1sKbgeh1dNdRjeQ4xmH733UbTMxtCplgVJtoQy
5F9Qjb7b6NvCtdjVTDqEFIDO5a6BB0FNsyF/4XFuIDjiwOzelRBp1jTYJbg1aey7LO68X0IYQVOl
UkoNqHONnrUevYYZoS+1dCHrXPOVoO5b3MWJRE/8PD9UqFfBHity8DdyxAE4KGFQlpgicEddlApl
NW4pDX+qG0FdhV7u7qdM1KMihGKj2v2U/ETNjYlfklYNkump98RxX5nS1DRr61kYOPoUoJ9LGGvY
M0a3BWitiYLLm2N9Q5m3LBKqw0c8l8C0EUostHn/XjsBxQ2iEC3QR06xR4kqQl6UKIep+EQBnP3p
G6IlfNJ+bRix4peaU2zBhGSjZbkiyDj1knzOXw3cjVgzlR7sWwbaBDcXqyU2yUEc7n5dIhk16KWN
ultJ23q118jlTUILucQE5VsitFyEEW9mXnYdmn7jQ1NNYEWjOU5s+og/oGYNcwX2cwWmIhEmj/6Z
txMH3lYVZJyNvSlNjUO2C9iNFf5oXoM6pen/AfPCVuUIC0o3IvCtGoOM4CY/6+F+iil29zTS8jwX
Zg8oUx+KIKP+ImblDU+vaOwHODIVvi4WNEorrQMQeD0YHJOA/x4y989mh1KvGp1ufJ2gJP/3k5MG
h4JoU+Tzson756Z2zFFbrYefsy7ZwcCrDIbnWj0+Z4+flKLv94V4z0ShF4Gdvbu18H54Y1j9Jm+g
GNeN9hEarv0Q/ddG6ws8Z6ji3zYVGvMrMYpnMEdUUiubKQnju87nZdLVAF5r1XXzv1haOMGoxFzt
FRYWVGLE4ujt1/bxPLtgrl+gZgIQ57Y+cWIDij5JpgjcjptQKFYnX8lz45FKpEhqm22zIc3zh6VA
QEQb5rN5LtukDPMRy5Oz8QsTzbwHVPxI510JthpQJ/efSrw5dhpeFaVFlDu5zs/iEOoj7l1UKuPA
LP9P3LpW4XnCt2pH8VXXoQuA5JKY5TE02tPgcrJfN0MyuFY=
`protect end_protected
