��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ЦT��q�e����6m/��p1��(����F��'��1� @����Gb[@���"]$���Џ�2&��<���(8#��^�qw�\�H��%�rI/k�͕m��-�ԗ�^��� O��t%�zKI\�����#1l|�"^B�꽘���Co��J�{vx]���3�w��A�*HxK$��x�T��`�\Rue��;x�wnȜ��;O���w���Gf��ʛʛ}B����� �ۖ[D7?��$��mt=��βҢ*�a|j���<tR[��˟�,�9L
9
Pq��l��2[&�w_��GWQ�Ci��.�B�n #����p��%�U��s>��v+ �Y�x��;��>p�,���E�'0��cF��H�^�1kiO	Q�Gg�M?!�=�TE�q���S������d_ck�h �Nю����Ϥp��3�ON�Vi�_�F1��%�"�''�!�A�af�������g��k#�z��/Ѩ�}YxK�-��L����,�g��y���J�x�s�����!�];v��~���P��\Yo���#���f�'�?�֥ppFw^������ї����O�Y-7"w�4a�f���Gw6f�#\M����z�M��f�|H�`�	�Ǐ���Il\a�� �����F��Y��:}����E�á]�%������~z�&=i.�Ai�73"@�ܴ&܅~��?q&V�D����M�#�?s=FN i(f$�b�44kv�K�P�Ɣ��]ZFVE47���[����KZ�܌l��!�,���$��V{�)iGf0<YO~�FsԊ\�Sp��켠��r�[fT�c�~<�W�"�U��H;ӂ�`�x�����tF+_�{�X�˶��m��g��"h͸��ˌ�AvY�/
�vNG%x)7-�Lȅ�j�O5*Op��/͜���L�<��x9\7QQ����yj�S�y����4��@�y�v��j.������=��}C8�uˀH�mw:g޷�IЖ�}���O	��{+-�A���mc��4�H-]>�DsrŐ�/Fs%���qUM�K*��K����z*o��m>��#nA�ʉ#����7Q�4���{.��Om����Eo�0r��eB��b>
���N˦� ��L�|�r����F�m�3��bC�e�c�g���=d���+�7o��(�y�hM��2uݜ?�)SN��vF1k7DT��K㕊��=�^��E&��y�Jx�\�R���u�<�H�#�����Y����+8"�B��T�R��Zo��$C"��Hp�<��l>r��x۲P��F��#�̩�*�����b\�Ϣ,�{�eU!` ��^�!Κ��$IC�-;�������� AZ,����6;H����%s(3�z�QI��E��o�r���mޚ}�[.K/� ���ݔ8�{_��+�/͠_@����p9�В�{9odXa�\��`�Ы���������׍:2��qa�p������m�C�ڪ���y�m�I�z�%c#m �_V �Q�b�߯:�w��GJێ�8D���Ýv�.�����H4���Q�9�_�$�����Z��v#B%=�]e=�D�&2�mqbSzo�|<s�1i�Z��d�T��掻��1�*�F�&K_�&�>82��:n��X��#�9`(�A#�SʐU�.��Q�n�u��cwɋ�	�b��<��K3c��I�
�V��v%����L2�*�Rm��A��,B��Z����Xa�������H�o)����ޠyj�3�����^�gX�d9*>�L� g���
R����k���\'u^���#i��Z�wY���ˀ�N�x�{����cB_u�a�Sw�"�J]���?3�N�xQU��]��2�j��k/)b`U����ty�������7 Ô1<�Dr[�5%������T����_��#�U&���Q/<>5v��km�<d���H��a-��
_{B��9��j�P�E�Be��q�x�x[���v	�]Ag�ý������Ňe�VsJ :x���D��{ �%��?� �V`����XS:�4�W!� ����۪�S��,�F��0ΟC[u������b�D7 � &m�a�2a��U"�{>��h�[��</y���%�����b)*;�@SmĎ\���̢ �~���)'KWD��)�$B\�ogMT�9�Бg��e����U��n[f��� {R~y�0��B����Ym 7���vYp%7Ms�z�˪,E>�=�
��Kn�Qx�LH�+�xW:�8�X�� o���{���E�Y�L��[��?���ST7�Ճ�T�#�K��$U�i��T� �Er������+���i����m�ω�>�^�մ�n��K�G�Oԏ�t�Τ_�^����C |�$�n
n�G�.u�货�E!���c���J���S~�89��R���0B��Um��ɪ�~.����Z�=2M�"�?�(W����\���B����A�����\�O����$���{i��%|*�J7Y�Z}�l��8 �0����`՘��qd����!z'��*!�d��1�޽�������h���H\�]��y�'��h̓�+yאl}�.���X�Z����jG�ӥ�X�F�3�# a��)iQ@�'�3	����p��$��u�F {�;v@݋¡ܗ���]��'B����R�Ȇ�A[^��7d�j5�x+��O�I�o��뗢T)�@S�����nO8<�yv�m�����������Y3oA�G+"�n�6�f�J$�I9kx�����u4e%7��"���4���y4���F;b��l��~aL�G�M�=�B�:�fT#�FLÁfb�b�@���\����vD�T�}ܿ��@�"i�s�z���Aȳ^'ګ(�)pF$��)p,o�6�\�QU�k9��PFˢ�Aaj���~�z�;�#�z���Ӏ�[������c������G���]#�Or�B�Ȕ��T��<�ǉ������B�r8�Q�38/,�I]P�(���
=��Ȅس����H�U����~y1-��lV���K��^t���5��P#�o>r 4��-Cw���R�}��Y걞�M�@F9�N��^�CϮ�$l��ɀ�T�!��8��C��l)BBs���S��_d���/������а�&=���?z�<�:������i�v�]����n ~<܄����<�������S�&�
J���{;삧��U��c9Ɇ��|�l���J���㫯T��hM�%�s�u|�5;�ӢV?.ƶ]�e�Y���3z���5I/?f���B��l�_���d,)ܤoԼ����u\Z�e�IH�T,su��Q����;cCޡnw �1@s���k.E١�!q���&��	�j@�:�@
I�iOG?�Pj^a��3gXZB���x�0�_�l���sc��|+�+��b�%B�(�`�2z�よ�x���Ҭ�o.I��`A7�r6���`Sa5��J�S0��jz����`p�:�X���q'���u6RGHCn������9�D�p�>׋���^S��\Ѹ��H��QQ�C����0�?�I�[	&Pb��~z�[a=0��@P^��X�u����Α۠�M7�)��X.���x1{(�w6�����~�.(|��g�SY��յ(㏄夐��	��)�!9��A}�! v+j&���5��Tu�������~f]
�2�H�����"<$!�~�a�(�6G�43)~�Lt�Y��a2#FŌ�|gϭێi�Ɯ����050	���jb\�<��`�נo�Z�1L,bJ�K%mw�!Hч���̉�yȭ_0�Aj��5F;i,j'�g�pc�;m|O;&��1�ƽ{��|�Ϗ�w9���E�G�>�VBc8��*k�"k�t���g%�_��}�J ��>�2F_:5�t��]��	�a�X�q�Y�!�n����g����Z"����>��	�~��@��~�G����L��9�����c����yg�?t�92ٳ6Wy( Z��8�z-�25��6��XL���,_t%<��j��S�2;�ܶIh"-~D���U�D�G��5bG����l�t[�7���	�*����m!0K�!l��_�]liEg@�wIβlh߶��7n������	��#��~���w�6��K�FN�~����)Ԓ��Ek�W��s������H�/��Ot�cb���s?�ئ�M$Q�5<?�p����F�:b!N�<�
��Dʱ�da]:m�˸X�]�~��\��������ߺ׵ouf"UC֎�y��L�!����]��F!8&����8G��H���z.�  �Eg�|�����ǿ;���y��o�2�X�:�a=3�(����a�A{�
�^�kU�� �J"ĕ�]o���O�S[
��OoR��1�P�Z�Cې�%�e`\S�X�@j�ʣ�4����]?s@�1�1�#����l
� H�sm��mڮIΓ|��	��M��,�9z8u��(���9������]쩋�Iw5�g�&um�a\<rm�h�s+�i�v�}G����}o�����41����J��<q��XlTw�?%�iE�"�H_K@{��R��y��ŤŔ�H�(bB����3�Fr\�"��l3�ˢ�DN�[LCU�wS�#>��S9	�����vC}�HIueyf�,�~��� �د���(�k�,�w]�X��|��>L�p��������j:���Гŉp���i7�_ċ��S�mTK��kh*o*��IUAr條���q�>3�VI��+�����P�ܸRn����ۘ��oMO�W���U?K�4#�A���(3�,�8��R����ό�{�[���,F�t{mM$�H!��+��"��5?�\����5$BK�d��]·Wa8�f��ݻ��f�+z"K�O/�u땍᧦!t�U��+\Z�a%���s�/���6B1��eK�zT���z��q���h��w��\=	5�!I�sL��l�J��L3�[5)�¨2�#;��k]"DW����$zbor����;���_��~�����3������'{Tw^sm�ظ[�����{��r�@W�	� [<;����5�2M�Q��q�2]+j�I���i�V�#��2����6�.�>�0�N<f�Y	5���� �UJ�-6z���Y���\�Q�s�LMOvi@�ݤ#�2��$Z<��z��r�R$UE�0�|B�j0Ӭb���L�pt?IP�LH����{�jo��hwZ6䲏4 ��4�L�������R��׷�c�
�ժ���Z��&�-Uoѵ�����N\�	��Gan+0�_uް^o�)Z6�8�n�J0��+�A,�2���~a]K����+@�c)4Z�^NA���Zm�j�[K��~ ��y�$RpF݆1м���qC{��/���p2�^ �*��06|���b+G�jj�{�G�2�l�(n�+~:��<�\�D'�� Z���8N�uݴ��-�My�#�*����O�x�iw�o�x�z_��\7���W)�����ъ�j����"ZX���3A��~.�����h�aU�'=�f��[a�q_0��.��Q��[��>{q��+*�"���Ĭ2h�5�Y����Z���@>b���e��}��aw=������.��%dh�M��s݂�㛍l�)I���i8|Lve� �DX���1PQ�av�FJ���G?��Qg9�#�e|=4D?���.1�+�v����v����_&��Ӵ=-]K�RJ�D��<��x�Gn��R��A0$��[&�U���	e$��0�����ȅ�&��2%�&M5	85� �3Se�����eS;1��7-�[R��S���&ˠgôt����b�q�}�QBJ�;��75|+=3��!�ߕ?
,l>li���q��d�m}�K���Z�XO`h::/��FŜ�W��C11eh@:�XC��ْ��/���N~E��xF����p[D�kq*vܞW<�5�Ḣp���`���9�����mL���n���MSڗy6���คI=�C�*ОU<���B�T�L����{�p4rs���#}��&���4[��Inw�_���EЧlQ^�eSw�ec_�n��,L����u��Ϧ3���!h9��O�y�����C��4�cc��pE:���WFr��9ݚ��M��:��\~��+)hjas�F8�[).Rgv:�0��0�a�5S%Ny���%V]��"@����x���=�#�2�g!��"Q����O�z��ɣD��z����O�:ř�5ԧG�9�������a�R]DW� v�哏��2Q�ᝌ��j�9v��m�%���ϩo�(��刎�G�rG{������		px+��x��Y��ha��(ڟ�V(�ܵ8�xָRJ5�՘��ϐ:|s�֔B��RC�,�S�����1��g��k��[�C��[��2IY���>����U��!�aY�y�&�\��S���$]�̀r� ��N5��6����p��d:��7��m�#qb}|p��x�G��(�lڌ;n�MZ��N9�l���!��<��@PR�*�y���G[7\�G