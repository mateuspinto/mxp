XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Tx���a�e�l�� ['D�/�ü�I�=`��gm��0��c��Փ��7dqǶ��8�B�Ȋ�;��&��hw�<(+ݙ��T'�u-����/2��J�Qswѣ0����5��zօ��l�\:`�)>���P�D����|h�|;�љ�����s=��&c�jЉ��8{iq<(g��qpU8�����}��9��t4�U�biΐ�/��l�\A!OҜ������H�jq�d�Ml<�8^�$k�����8_L=�z�6y�tZ/ͬ�ǉr2���01)s�G:XjA�.[���v�������N�V�l��+��v in9����_x�,X�ZW%�A~>;��a
��77$�=�i��K̍�О6�z�/�ËR6���Ir�FKm�1z	��t	�N���Kl;��Y�
/��22տ���:��_�kwo���~�˿�9�����w����5������^63�z��2��d�]n��ihh����{Cq�u�����C�5�W}�z9HQ��Il!�3H�Ӑ@���4_A�t"/�M92_�W%��������J�)B�B�X�I���~�~��k��1c)"0���O�.����� hF0�l���P�IR�_l��W�>8y_4:���둈�t���>�kj�\���#n�%s��`lj� �Ǩp9��GI�!�`}0�t�"Ӑå��bަ�d�	-f��)��|�b��qG�h��ڐ�?Dٗ��mf[���}�x|�Gi߀8��f�2ȿ5�����0�Ƴg0�vXlxVHYEB     400     1b0C�`<,�-I��T
e��d��~�>��gЊE0_�/3)�hf���DY�8�� �
E��/tNX23���ժ�4%��aV�H�'2�"$nq�'_$w9n+��gy|��c����4]�1B$�T�H�Rn�9`�n��|ҕ�c��f�5���O4_���	�矐î�^A0U��K���s�F
a�e�ȻC�8v��3�f�i�DѢ�d@��Ao�)5�=7��Y���i3 ���ޛ�=9�e=��ާ�i,���� �H!���A��ʒ��P>S%���Oˍ.����7��))�E����J|+(G���Wj�{�$��L�'�6�`[W�y�&���ʌ�E��y�g#��&�WQ��JR�XFG��5�F�>r��c�w��S@�}��g���>q�tȻR"��i��B�����(�� ��"XlxVHYEB     400     170Gc�O��?��ķ�u�x#�|e�w��8R��W����
�jRh�<�d���XU��š��ޭ�iSr �r�Ќ��1�$��Π"ę�UcX�9����;�T[v�nFu��xvC�e�%��8!UVٝ�jv�~x��.tuei�����?�f�OG���y���Zvu&"�Ur�i0��dk�m7i��4��!�@Ҕ��nȽ��e�lKo��M�!M����f�v���0�C������������fUs݂�5��m�^� *���[f�� r\�w�;������ؕ%��[�V����w��`��a��2�A����gPܔ�v����!���}��׆�����|xP�t*�ۏ�?{H��ٝ;lL;[�clg�XlxVHYEB     17b      f0��뛴��$�9�b{ɸ���w���4�w��|��Tr�d��3,L��C0�Pb"g߻�B0�W���nЅYh���Rp�7?mg<����������$�x0x�>������ޓ!�����E��k%�h�;��IJѻ�#�5����NT0f���k�����{�n�m�U�e`��H����Z��Fa{�Y#�VC0gKd`9��M
�����R$�˨��9+x�D�)/~��(#