`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
pRCqdBXtNxkf4COeI8hkvD0sKEMxczTsY3SsGAk+Kpj81tmFlcdLXTG8Q001t3eq6gEdhMTLJyFS
3q0RPsDeA/67VBHN1bnv7kDCH6lb1QEyKidzkgE6WASp7f78HzrFFoXtdTPg1EgdwJUQqaDO1Cx+
Ry+oKguBgsiuLDAxuEvcP6SamuvJqP/1SYZwmGMsCZd61zCLyaar9n6saMfjcqOHGvUamJhvNqt4
o0GkHMeAgz1bMn6KgSdJcO9H20+kBgzQ/EwzRBcTMsrKwIPrx7nZAMc4PbVtdObFIpSlByZvCdg9
Ch7dc4jQtmNMSDJx7vNX/4CamxKYYDdC1S76IQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="sjcWQngevlFpF8T4gCfqoNE9ds0M0Ush8+OrO3nKdYA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7232)
`protect data_block
PeFHc71Aquo1U5m3U6/EQZQs6TuKMdF7/qPXqHGUwbAuDX7J+SQXXXgB9GSKlD0iebxLLrWfoqmb
axfgVJHFX7MqABJL6EjEQRm5U91MRphjpds6cEe31Gv97pndHIee8QZEu1bHFEsV2Z6tk1Z0046x
wyzSg0ykQomoJcmrHzpo5Fc3HhX6TgVpEfu2uA8aam93CibZKcmQXv+2yoS6Td0ljGzvJnCQTzdf
dsiBPGcvLtPv/Dl3xH+bK3bsu6lMfOHnhU+AqPk5XTHXzigNzJ89Tmve0Ebs2WvlbJAlMKifcCgH
UTlnaoZos2uP501n6PFTWl2Z3oUw9whi6AKiB4p1lmSwiU6qWWLTt2aH4SrVqktnuyuMwknH6y4S
ryQuGziIJLvybv59ry36LioEAmHRa1IusbKcLtK+JVf0UguitJRTPqm3sDeGjCTM7hVb2SAr26eP
DwcLhU4H6+/z5Cu5N4qL769cgtqnbNgLv+6SCwH66g35dZWlgOI6hvsS/k2NOmB276ZheXypk0NS
dNzdugJPoFVFLGIjVE4A4QFRFiEm2HLobg+Q8MutvYN7/uBhREMuliAqd3DRkhi3zpF0R+QM3JoT
Hj4JtdpyhbRC/TiTIofBesyBqvuoVVCIUUhFLih833IhU0/HBKWp38lV8txrCDT2EXXdeSIItxex
bRY1NnBaWSKSv2V9SH9PpCZzRTInginBQCxRT8flVwZJD4aBmwDJ276uw60YxsFrO1GV7KKc3+M3
ofg7nrFURyyZdL4QCSdaSqnV8oxotxCRRqDEXP6X1PzWQU7v3RImK6GqLBWtzEqpeN/QMljXm5Ue
VS/+fNd6chIjmHkABg/Iqs1xX62Xfl1iy0AXXj1DufJbtX0Lc29ZufTURTkHdLUApIfiZo32Jd51
qzaMxpHKAwa4YCOmGN3ENgYJs80Z0EYAZDYFA6JKZO4vvSE900z/sEo/dZlFeS2NmG8mn58P8fO9
qA4VWtwNzqKvhYUpA6zEnHWp02ZHJeUz3dXa+vXaV5H21rX3qKqkPaYNB8w8DNQhp3Ynv+B3e0TD
bHmH7gIglT/WgeB6mEIaQn2ulggtkRd9oNgdcm1vVODG09uYiGRZo1DvAUdxyZtSNUTdD+Q9vfct
ybJwMvAN1/qHl/+5otuIDg0Y32tYQXDaHfzCPDy9lKKgKlI2sFv7+rr+pTgPYzBoO/OBqypfH3yq
DB6fud97Uhx/pf4jd0sPeesMNxX4POAymZFB27wOp/xvIaCfWKwAfDbV5BCtS+DE9Z2GI27CXHP4
xMbLuUJu6tGJ2aBH7OFOLX8FxcCcoXwwiiLnXjo57pcZfX7kRY8Cq88fqdLl5UrkKW9Hiz1BRfP6
wZJCgTp07n43keGLlsbSgvZEsPpeiugJqMvx2BQnwwPtihCvftTg8RHetXvUWa+3hoMREgGNpTUf
auarkLpXgZIUjArkz2Dz1vSPQlCbMOG3j21Vmevzt999Ngj8dKassx3HvgIuN/yBlCiu/AORmWdP
cMN8SClhxgC2GwVTft0CgnXGgAnncattZkJx3OL8+/rFnHpQ7eTAfHZm4vVXAKYyy1r7dQ/8A9EF
ydQSIRm8DM8NMAnXit4xBE89WvVzC2rKt3D4FQ8jP5P0CmEzlMUck/Tcc49L4SizGkZWNDcVBwF6
rtnogqcqqmFOYCyDmQC8xn0MwYKiLXFImHQAX8fmZwjFtt0Ewk+FxOSfNZKU4/Dr2Wr06scrpDiW
5/cAUkbmjpQGzfwJShd7csMUutc3DzMTv+nPjYNgSSbl0awzChYhydD2xpiHJJ+KRgouLHv6QZ4z
R4zsAYpWXZ3X/sNM3jKTMNnSMitVkwK3yl4y2IfbibwkpC2Xiv+RICf4LeHRg4D0zIGts1LV2AY7
DXhicpzROIuas4ZDasNF2k8r0MU+G+BvDbU7cpkNzPYxtS0KHcI759goOcEl+oosawrZZ+PSjMQa
FTMijJ0JbB33tW/amwlH0uZyG2gC+KCfuP/DQ+/MnF3cK3iTUQI6NFWB82wIhyoj7Uf/oAPbGGA6
aCBMyfsp+tM3HYS1HFybtPAdtZxE1f7oK940ZcJWJI6jHvH9oFzb3YlEdNLuZqtV8pMdIioRYekz
W4QW7N5VlC3Q2q4HPVqkDLRNGO5sfi8O4P+PEns1cmK6FvDUBnGEs1uPshzuF11t3FB/vXD5VCly
LjQuN/iDYyYai42/MYb7z7cNod6Nr0xj8f98svHEwhjAy1EWUZIKxNtJ8zNw/a/mEmxPJq3hTMC/
0S3RuDW2ZqZ0HknYjoqafd8nC5CsE4BDAi9PisSl97PVL6UwUZ4jDZ7mBhIwOpRwyftrNSZ29EBP
TBUrMqOyrqKOdhNbmmUh2hnmGNCYmtCTbV7IbqkfjAvaEntstlsLrNN+R5TDLVNpyuaKaTraLdNZ
9Uwe2K4oD80SLm5LMtkv/Jx5Ss5kTIBueOS9JVEKlG1fLnjjM5v/oy7M7bDqpynoHJn2Y7w0x7VF
7cz7egiLwIPTolFQjwCLF6TuyHi6oQ1qkniVhWnddK5Vv3ud63Qu0MOx0TSLR+cpivHxp/aDc9Da
tXEUetaiPyXoN/wa+S2DrJXgZNQxxvyqC/eoH6raW8BTC+LrHatTwaM8rl29yoEV7hentWrS/N0+
anuxXX9Q+SiFyrJOK4lBous/mozSvVqJxEI1LdATCo1wkOruu27v8tJNPb0YSSZbflGeQfEmoBMK
0ID3uEeYwg7/QSHJ0U/8nqBwmyRI9/hZXmM7nRk1lGgiEnL7AyzWCapL2A2fB5oPi1FKn9pFW2t0
Fd6pxruQFkFuhT9I78DjQ36KhqqDyP+q3M2+ABbACv/jb8dn+4OkiEFPMrXtvhzGEeO0hGlZFbbB
FXaFV5T0PxZ/Am/nwhtYMA4/XkuUzIw4Nh6EbaB31vbEf4TYg8v8Bs9b7+5yFFCNUYNon7eveUFK
ZO0kP0FHzKTpMWMFdJ+RX91hWCxQ/wMiv/sWXJKHxdnwXA+nyHeARs6fH6kJ907ZJE/ruTylF1s+
cS10dTEp3RVOOQy4ubtHMzmVzB7a0it/tm+q69DlkKjVL/axNVJ9hHrw91GevDOxHZA0o2iGIx9j
RQ8gvXabejeotu7akIfNDLcLXZm+NDFqTDTd+gr1eMq+NWcpT3wAo9tZGHzOr+AGttKyzi2EB1rX
JyqYErxafAXK2H1CWDm1TVj6WQAoT/obw1isgTtkXaTRZix0xKokNayOBYFnNxDVCL02ISYdnQOk
9Kk7W7dwz1xsOkSs1SwgqDzQBcKD4AryzNTGmK755DobSB7Xyty0CGRZGLOzCsg0fdM/wxzx7XMQ
F/SrZgvgwZMy/Wpt8s/zhFHlAOMp4+whRPH/ZPMELVV3F1aY1rJ+rP08JZR7+AoxGYgaKlcfXwXQ
35ZCbHDeLWlyNmf5RfH6F3fmgySbPIvrNM7FbAgnPg/oYoOr2ludX3WW3GE/YhLislK3kXOJCfFr
n/rTULV139v1HH86ReQg087PA3c4T0wP7xJe/OG3cIDyuOxIC0TDJfzbtjMNVAAIC3ug51bY5jNX
/RvTdZXcePVisjorf5pCnJNQJ1FTEUEyJZn2zxOiWWszB+4Kxq1UYxFjN+j8pQjeMQE1BGdCkPRc
HqqaHNL65ECiRZ7cIUdw6ITmVjP53YUwRfGaGM6H10TJrW0DWECrZ43TyyMpPgnjvWJzG9DNSa4q
4MKRnVEALyjPc5xxJiZCFEkQUKoHTdPAIrLQsdlaJmh43x6Vh+AeAm1KZyZ/MjqP+cPeDDW2r0wV
Qg7NH+Ctuw7R+Q8dTMomiivSBJ6rJSCn/9htfZ4aBsFYkzUd2JCrj8wubNoe+8C5a35rQgRogBw+
NTPSd47wx/5R1HAgnVEKMPmXSkPC9g1gIjJ5+HSlgWbJWSA7Hri50CgTMBGR416aUWoBglD81Exv
EICli69D6r87aryII8SzRv6jndSGtJzVKiVMYSwikPLZi1HJlEWMSIMc34s5uKnamud2+RN22tUp
6+MVqSSJWndIN7fDmKz38nVtQ4Y+DLGvG2j0dW4D3pzk7SRtTU1qKrjoih0Dx+eIQFs1gXn5+wjJ
gVs4H7fijWrfQ/UFhOnc4DR9SQFmpkTNKjyCGg8sayRhMlPYLuoKIX6JJjUMC459JRu/NBFxpXFO
b+Wlai9dRqvyLzSJIF3i/TgjYpJVhMUFSwyd71NqFZKLTnlzuQaG9dGwnQsku17Y1a0clF80SeL9
YgbgIrFaUhk0MlJNKZV2WkN18UsazZXu1+YP5+2RYis/8/pDz5lrC8EBY0LuxkMYVCbRzSzEQ86E
syHFmnW4d4xQcx1JvJIIos578QjBefdqD+AVkgGn03MseYRaeJfHMf6vquFWbz5E/PRxK6L8yVH9
4/Ace5ap5OX47Sc2+j0oO1Eb83TFs6qiO6khzZyZ32TeeXDlZUwtLJYbsMz9CAoL6DBGrL9adWwI
InnmmsYqVdEWf7sIcGw5jABPR+viQ3SeeXZqDMoT4x0uxlv7QbpuRrEk3ON29mEo3IfQ0N+dveYM
Kl0/4FoS4BqrAf+VrZKFfwC7qH9sVLcZSnlMG+Ey080h5v9iFL+3yWLdwPwWS/qvdZohxdyB7oaC
xNuwiDJ/4MOC5KnEaDSJTVHnkWCCMxmMVU3RayhxeoZKjvqzKB1k3cbUHRkZKzzfcwe5i40Fbu/5
1LaSXojpqjpLeqbFyStGqvBuuBtqf0SFVHtYVopotsDYIYgW7ZtcaaOI8kGbmg+r0EKQDejzkg+Y
9znYJA5U63h5P3YdxTf/PtOfapPmqv518Dl9/KP45G3q0+XpdDOV9xLSiSPtSnJXYTTQY1Ww1D4l
tnhWaXggnb5HQXxbzWOctsnHHZnQDK2ObOSCJxcHA2fGUN623o8CpEUNboGEC6UnwLxWJBrtOmJ7
Yo6Bv2D2OzPWGdVE0gbXW6wsGrhwpztEY7Vsv9OBpgSPEhvOXxUX4icYoqTHF+ot39K/iNcrD8Hu
MyTkJNaC8OXBxzYCEOkuojOnf54cxM3fCVJi3JQTSKDmSgO9jASKuFuviVtMa0UrBzglq4R7qCUe
U8Lauy5/l/wBfK0LgaOzjwtKAziO+nDMld9yY54e0GeAm8Ta89hnsXgPny5gbxG3OUA0lvcviTaP
ObAtwnhnei5K4daTDWOZZsxOojKZI1p0/ZmwFA+Iz7SEGzgUkt+FFGgDcksuZBsUNV0j5fGzb0Q2
Qyx2HNRDBL5p/DWxfzj107xJr6p6ZvF7Ee9/iXhIjeEfJs4c28K6nihbxd0pdX/BR5rGCZs/sikj
Jt+JsksluWEqNLqyHLjwtUxyC8xpm+WulWuP+6wg9e9GXxoFIHB9xb4QVk+dMG4O0Hx7r/Jh+Umd
wih/7ZmiaYLCiTAGnltPSIl38b1kjTed3IH39v0NfFh03g66FkHVcF8LavqixFTe1rJN6Y7/A97x
LFuV2jnkm/72win3woKyRU2oPULhInPi7IXS4bFTgZZJaQYpt8yIx8Vu7no/EzC3Y+v6Sg8eI+bT
R71McY9ICYWhDANEe9uaZGWvoMN1E+vZIEOMNIrtaX0YxNPS3uRomVxvbARt8hoBNXjFAZTVDhsx
Z3gK+InWIAlRrazYf3lK3zdtLXncwHMhBOMO1U81+LiTWGqLlYyp4rosWRmkct3/20osOtsR2u/u
qWy0ARlrF4zZt+OdUETnwKdf66j3ZKxjDep6eEQJlKUbCP4xtB9DywgQFIFxjgYtLW9tLiH2KCvY
8HOEsaIulX/RQbjXBge+U+YJDYIKMyUeVTKL9ztbHvG5x5o3aqhVsWw63ESHw8Vo4dydccgZeJMR
I3XCUFtm8nNIdAAomeGLwibEMl1GFN2v0hrQeOFdTHhySJuciamuda6OvcMMptjwS9KhfUkf598C
rzEiG9wDh2WzYf/5Hr8F1GYYDX5+SAPmxG+3nVZYIZL6ei10ilG4wo2wu1Av2p7t995aZFZ51CPj
tjyUsnpKMKxxUOuOvM0jFRlJCB8hrYiy+PP1IKnvDRiO3qDYTnYxbKBBXHrwloX4DvrfYesvvdcx
+7Ler6/JCuKFPycSt/b8CHbXOpQwVSeG+HRuMZUdCB/gBChP1rUWG/gPKfGOaZjJBK5sPEQHwxhw
J42Id348nB7wB0+gsN9dzBiVNuJoWrjjLdz75lAYUzalzXclvH1KIGrPVJlwJVdjiMITNL1IQuij
pCQws28rgUJ5q2ugYqR0NPiWkgGWyipGrjXwmJWR1+UnFxP6ZLBRSL9e65hP4GTIUeLwc9lXhU8d
fl9C1+TSKd0HMiILBNS6iYxoW896+YZB1wAhKUlfYWxjtoxRWN4MseOVLn2P66wMSsx32rnzCjyc
r0Wap2Zkpk34t8og0/wC5QtvdyXggq+jySoO1j1KyfRvVHyGcIQDA3jzjv21Sk3DYOnbVo/Qe0S1
8Q7wjAiak6Te752oWlJu5yGsOW+Qw6fkzrt7gRwrxepXAuV1e0xTGz9Cdl8SAzw/mGYt/McKcprg
T66jhaEQUAWfw5AE99nxcBTAFXgunm5AeS12MwJXZ8FZa3uRhDRTdueYBoHZ7DIjZDrENmC5DBrq
R9OOgwGs/4B/tD/oCajOkiB3GUsdys86A9wV3bDfrNd2ErXdHO5C3RZ17AkOG3/2Oc57NcUTTWfp
r3P5G7u2jhwHbw0xRbh4U/rcTq+UeeCntdgS91oUhtrSF2dPk2IVOPPZCGxMjETTKnQIj4yaCIiz
VfONbXFA2tcEI0U2ktC6F/C+DyWZC7VMwJ/ppgyczByUQX6lGz+WfN2zE67En+4EuX4IaFEFS/fv
ku7mBA1VN9vkCGg6cWfM79ruviRrGZYZ/MJGzEMjod7lalpBh4k8Mszii/m89YzXBVZW5bBldorb
LCoNpI6Q3oo3wa5kjY5qfrb9aWBhmP5C/mI5z1BFAgOlcOUC9iqauBY0md41xmJaFUjbSOti1CXo
LueFGx6XsHrxGwB/7t3LEiYK8QVPCglcUaW1hCIgn+rKNdzkCGBga19dIW2HnVo2mOwaVwdJAxkS
Styt0Z0RDLqYG3QIdkhn0uJZisF4LKgxNR4DTXCqE0o7yOF4GU03qUBUW5NehEwXT6oCm5pwt3ju
BvPRtogSi45SbUIZQZmDNRrfcOoxGlIvKz5yiu//G2fFpsE6q28gxAugP0qlyUc5nVTCjbM9EMkN
6x6PR0kB7iHd/swD6Z7DNdwLCTwfhVyg0vX9pZpGYLcEEMFcbJRKIi4hPH64a85bT43E/C9fVMGX
XobqoQf41/XIEhlsbBHrdwocIpx7RBxU6cz4k0b8ug7ZdWyRmLvKjxbyCvQ2aFDUa0oXgUZPOxDc
puenRH/n6Lx1ogu8btMwLuSp5qww4c/vwugDfGXzY+0RXJUEFDbrZC+tCo59NU36/F+NhJoy7y6F
3LEeCfGt/7el+rikpCY8QNi1XJvLHhwfxOqOTDtISpQ0HCmVXiYL+/YV4n06RyfTKgzlF9oNi/AM
6VxbLCgaVk3ddDyuHZ2o42nIIbrtboxG+XNb6SRmwBxCDZOc3z1Qtj4M/+YgUL2ZEv3oDCQu4xh3
wkS/+/ZKOE0jU9Z1oHtA2BKaaB1bnIXTdbm7l9vjWDFtYrKXJfz9l2Wny/0VOOHd7Y8Cu9j5z+rP
vee05yVSqrgQH/q+Q3NvowZHAfNwxSLlzrd2Rxa7mYvOKccso4Qu97WdoVoCU8XXFGIX+u093KXv
FkwWDXy8eDFTxalbS5pSGDR7dGvALYzeva+AlmLk8rptMZtEIl8DP2SX5RXYzVekc3v1S+kXetRa
Pb59k/gBfbfqjDoiGC/Lh8Z9E3aN4ZH4XlH5bMpdSI2dzgAzfuf24e2YQmrzTNpsNNkHY3WRqxa8
lKKYI6WRdBxxYUqtlB1fc9BElQI/MDgw+HIhXUYPQFSJzfvPdCBOlYuksS4N1DGJWznzE2fTFvUF
dbgk2RAuDBhnAucHBtCPv430VVKgHCoPIXQxWnBVkJJC0GTc4XvxesUqslMrPZ5ygJikid7exHfl
YhpjG/QVvLng8u078Evr8JZqqy2m1v7jExfYwtLeEZqFgrXVWAsbgF/XMo0hb7ypYlHwBKfGZlrW
daLq9Nb9vJD4Fw8xu2ovMmGXrAtlKW0UdBG4YNLVk1lZiI4RUU90XGOccN9xRkEed32FlBSX3lqo
gjf+ApCzsTmt4ZwAAtCqftyXtldDv8thRAV5w4EIZ2PImr8eTIJZQUNSx5YlWLjxqjTbEvwksPqF
kQvcGmUQBE0ue7ydiOnkaOSnHZjgVJlytt8AlFP/OFiRieI/QU9BAJLIQgYKpZCMkKhUxy4lR1hC
b+S5ba2iDjCHW8v/yyHNlgE3Ch5njt6Txw9OPQm/i6R6ne+i5xKKfQF1PDSkEdOpwXzwaZJlvv2p
XZs6A0LTf/gm3D1jT4/vZtGS3mwkpC4Ankk4LDkebh4mjhU8J9W5H1P1o4ZLZ4f9EqFNEmctlndT
1qURaw/9LLml4KILAzDT7mVvlaVuuvl9Hy803X4EWx3+bun04Rzag6nxFnUGg2YjL5yIopF0vTHa
mQFvrm9ug5FVF7GxxcVz2f/B+G3h6XLnQMFId7zjKfZ4K/1SLivzWfaNGVKA2wNLEQQ71Kn3aE7l
XKoWGnL6YMDJTDU85VhkGeV0LYAIGmubS1QV+BvzyWmYNBtaLq7/0aktuO2V/hGbBiHXIuoDkQ/t
9iQzTuS1gfqq2YTFqgKQUvycaxsq7Qbs1XpQY3Qh7nmDrO5x9IsLZyHoHkHoskoFcmAp/WtaalR4
8uVSTbYMPm+zoCZ477SIVWLcImY+0wNwQFvW8ZWr3JEt40YbkCqT1RaVueoye7yKilGKF24UYbMC
t7bXuKxie3OukCtQa4HlEUXg83KPH3GvvJ8sbqr9w7LgHqbqAk3OBcfrnWBgKKH/JjmkAUPz3oTm
VeVphsN2aBMNuDPpOKpElaoMEsafiAT86wGeGlbTnEU6g7qXAfYwP1LKQTtBE0zGcwbRIgHzOL9m
SDzROHxhDAbEllORfWQrcev1Cpv+Io/RcKadi0tw844LtFsObRiXJgTskHewY/41C46tnEfvuSFG
DipkIcbt48e2HVCNzZ86AflDKvu2cl2gTbCc9iVJA2y6f6O6rF/yjNbnavN195GRJ6w0oi4YnZTd
rbk9+D9vQzK0Agem4aaNNUmTXXX6oyyXyhIX9dPBJuu2W31tAyKB1wwBlUeX2rbVSGuEXuZv50/A
GxJO7z5WPZu24sNryS+XjeRJMMKA8/W5ErwImq0AlwVBWc31o7X5r2OyOIdgmaklkC0kg/vLPPqd
L8ssjDmhhCwfDA8suvrwENadiTXQUkFNX8qgvIEw8ZGxxHsAfv8HSxO2KNlvRA3/p/bypcdieYM+
xcfQWgVT3xxq7LSaqVbgHn8jbsNUlnlf1HOYn7rYqRahdUrXJBev+KgSH6g4yO3lWhe4BjwtYabr
tk1M9KRBezykU+qOx49F9k/CBxxt/ozTkfICm5KzDgM8FhKdpDH20YsnL6SuL1hUvn/+ua/ZSqIj
7LFiwJPlV1/RQUHEyq6ZcFe9EzbUwSP+5PpZ/549mJlC8ExkViAyyo26oG7zaW198YI=
`protect end_protected
