`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
cPEWnEN0uTCRSI9me06oq5eGzOyzImLro+30j1n25ABwSXKBVMWJMlof6NbdKEJNp02vEvQLgP0l
gdVzSBs/lxsztN3ec6AOlStYcLTQ1gmbZ6zlukRAmuhx5JbSKQPumnKSyopQ5U0FhklELPNeT2c+
BX1BNOOvtGTZ5wN4fYBp0tDHvyUoHO+9IdyhCeziYPqBAVYQTRmXmIknHhAfhw6hzDv23Maum4EE
V5nzXD53gJS6ik9UnH9R0oTpyjtilS8aotKsjARtrf6xD55tTtwQno/rF5ADfkNt4hrsgqQ7FQ3j
D3oQO9sa7l3UE66cC1XkazBo/LqADiE+ztDT6ra78bBn4GRaS4+GpkV0ldUKvA33E40ZV4fbDivA
rbzoHPG8tLK7yy/vjmapQnHp1ehOpJMB10zuRGvWNRGFGR0zN2Q7eW7/XTygkUd6Sr2/yBU9mcmk
mU6VNen6IdP5GBAcNhnGcY/u81Y02QGIcqaBcCdJZkmbEaCz5f/xmNDjtk0cXaO9bYZN1qrQC1i3
nNAQ4X5oENxUaQDOsAwykIClmm+Rbq5IgactcalnVZPrbmlMfdhcUadAjPD3CEhhbDJj/5AsDheu
31jJ50U+s9wdiwqW+/UVJlTMpjSsvxsd2P5jpXbkKXk3GlpS61mTbtYz+m6z2G5yyemrDPt2iOlo
6IemNDGucSzC/K7K97//nmwebkhKHquQQwzK9oozUBvNNosU/CY+AruEDYZHp78T5A1lBEIMCntf
+PQdq9I+YeK512vzbh5mNgiQoaPzY/QMRyxjlxKD3YXAdjkeKmaFLWW3PuUj31JjMOetLyQrCJjZ
lCBD/yHmviNjj9YUSDNJwI06vUrzckbabaU9Dgf9QzHSIveYeHuG4NNbLQoBUWfj97ZU/PeQJqEV
CcEfDhAjdSNVExbgJTAgJx8ec78SV3Cdgsu+bobnrq5YxGQSH9R8suHwrtau0hDO+hWv+gRYfoL4
D4SAfeBtX3T5yPnFIxP/H+kcossLpf+HqSxjEU5zNHitV4ZG0vFuik060sa9zCq0YhtaZ+r3ddW7
thJSi9xC9lTObRZfUWtfGHANrMTgN2g47XWArf45qEAXV44VwEApz46bv5J/uRL7hm9E3KvJAE/z
s2MQG2IpxydW0kTUfaAeFNk/GZfvaUsskjbJ+1glGdaX56qs8nzX3mTy8bhqdcQtnR4BKjTs3H/l
y8/k5kaXGauMl8f/Gx2VToTwXbx6Z1tpCLPxlo1zuXpsVkvgPd/hYd7SV41U4bD0LyJ1EDpkANbq
KaT35WZ7Ygr0xXUxU6NapjOdGb+dVw9Yz9OhAlnW8pZ9eib6Y3jkzgW7nEXQCCy5gKmAUI7eHx5g
H1vtgAoJ7F6IFOvyzkW+xZMooAv3V22zeCMOV6iArY9ifk9v6vX1bW4ke6NRyBKAuGrO/B1kCWBZ
phXzbccA7ulKbmipUxl8U87EvFCOKFFU/dGvPOKUm3CDNxiS77fzUbmOZWb8Zzmj6hcXEL+Oxdn1
LfJZHQCquYeM7BCEq36CCB7myj99L7YEbJeljm9jNnwdpewZfNqetmPMGseJoTLwDtu2Wjnf7j+7
uWrUOidDnvpKeOfLzHkrTboO6XhjgNbK51aphr30a1YVqj4tHCO6VyWsAL9xGVTXHhf/SjZwCeaf
Y3UegJKEXNw8QL2bqodkyCX5Wtc9GyAjq5CO5PDQOdkyu4PMIiFtUYE829yDJKL7QZjmGB7fc29s
hLrGNe9GnRRGRhVZ1vutFAvDBGGvYk56xGc3RR0Y/liURW44cVB8auhxbPQdYoX8Ro2Bwc5SoJd2
sWFSVD4RvTKSMviuzagI8P6Pe2ffwBh4mVl9hRw+w/FlE8S6pcPbv1FRleIrNjfO6jw52ahuPdTr
sZzLU/CxOgBqD+hWDwTFj2MBV2mHn3w42bA2KZhAMMqUmv/9te9pSm2NLE98XpeY2g2tk7dKUZTW
XU5VGMkvoWyPa1eITV0E2ppDqOYD5tBQ1p87Wc0kSZ5sb3IUS1gm6DUyUcC0PnVjMCvbmgPxMbNS
4L9WV0Qm35LphTO2rF6AWGtuHO21gNK4H2pbUd1hxHmnfpBQdVX0I+88XebyvOREoGqHTdRcdxy3
HjUDzmTWwBNIXaHXrGB1h6O+mfPHCYZQMtN5YrTnIlVMBzljokZpQdTtVuSBwgW2vUpL6EVG5AvI
lpLfAqa2HFqMFBJHU66XyEUBzNqyqPfNzWTdK+HIMRhH2z53YfvgPyFjJRLQre7CrnoY6oqpbB96
AN7Kr90ek/65/LPLN+sDF4sGWmX7Qw1hQdIAz6GjhsNx6XD0EIs0Xq99gfUTk1aGp4QD6k921/b/
LhlSf4dYHvAK2rcPQLMqC0hhafH0xCfkdC8H1KNXbo+P6wASllbVwGqgzFeR1wT/XzRh760u093/
vkY8itAcXEklST2+jturtQ26SByOqiGODZRDJlpbYeLH+cITEpZsYM+yhu/k7eCYpiXcz66BnHqs
Ps9oPenqVz5tkKA4jfPG/RHcTpQHfJ4O3ikEdRFkyOogLUvUsqwrOJjJoKbO5Z8KwrLcUtfbiIog
fuV3HcEhD9IBhqoErK2qN2wWBuXoZLrWfdjtWsVnElXlJyl+EIbj3FRR5ZvsnPpgx4srJ+NeCU+D
XaZ/7J/8cPIOoZJOzinoPPR5Vuq6sRKTBqnGH3DDc95kMhDTtYluwH9NdKYz7Cq6TnTNBVh2JD4l
lxhrq5sGxKvX0r+A/iIIXw8wZVl6UXJQYbBfsr5sE1q+9bJhotpqAPRl3zDfDqOlb76ZXi3EpEsv
8Xx+frtOcNGGLZePEU8Whqi0Q3HDpzfI8np9VP0avpejs9JDMkQzgzCNn0J+3XdbUTAY6arRlN7G
IwMK728AvE4A5bcMBu/8oC18xmBois2qCgf2YJqphLphbu7F93ZX+dYz9N6wBRvVm6x/DDiwgcEz
JwZlkrn5jD9fFYutZkY897CWKD6AaITfGuWKAGf2jQs132wExIYRgtam1FbJdxZ7IzArfhBde307
fXeKYMDsDEnWPm5G+dgFyLMo1zCOO1KyzUHgBKzW+fZjzlLUdFba0kMnhERDxtnIMT1qUekdUWup
AHzp5zknDggZrfWrCDpqcCDIKpellnQVvpzWilqZz39p3f/oMsk6ubUtkUTTrT15mBD5CaWfrqg9
Gp5/Uy3aFwCT/gQNvyAdzb0SXXjfOLx0TnDTBe6dduRGDTJ7mkoDikhkSlEJLU3r04oqwFBwlLO6
CYkFEol0OMJGL+wllYT2cSSKDKMhMVTYUaTdgMnh+GAeo6msqqX8Q0p9DPoG1SQici3EffxFsq5j
pfk6qvWuMBa41bSjwV6hVwtckuK9c30IkOCxJTOR/+qgjNWtM+gu3/+XpIZ8Dl0vRrqCo8D0UuFF
j+d1W4oaK8LcmRCjINJ1acz1Ve99iKsh7npVBRGKcpyeuPfQfj9KuoZGZg+9gOg0K7Tav4hQ9Fyu
GhXtWZd+p4Y5B+UcGPc4SPMxsMmeNEh4imwD+0FJrr4KtoQWnQjtXup5YfWgobINNhdH58DFztry
LhCieWIM6k1bUrXHjwwK0gUVedFEhVA1mZOlipYT9AwQkmcCKPpFfF3YSU6aMGVK4a80CjoK5mwm
/7FBrHZNV19NJWnGTaxqeokpj3OxJJ+Pgl+ZKqDyFNeZEGtkjFJhTLUJOjUXWcAQcaaL6n4Y5fdP
oB59KS2M0ICwCfQP4qkFeWQ7yKFDlyr5O5gA346b3Wet2DPUbd1L1jq41GeL0Ph85GseFJsPRIT2
f+h0qzIFfRq5Kq/PPmSkSkWh13lD5LDv1yk6RD6xOkZjJ5FmfDBJyBRoQdEQZA+slpFgDMltRcgo
ExlkelnHp2NYZoQPwJMx2zJIqK6hRdZYcFGSHwgeaDhqENhnrD2KDUjPNLbDipViyHqdWG6HDyO1
VRA9tnkrQoM/d9uM+zo/kASSnQ9X7WhNnM0izUvcQjo85c6jvyE/ZQoQDr3bKrYp6WES4AiOWpfI
rY86ePOQXgyoSNq3+TyRJI7zQkCHODLfl18GNSkAlk6pbi7dTrxrftOllWY40qYAiPrRyD/pDruL
3MD866Jvp4xHMhfmJFLgwHYAj6ejn2jx+6j5+aafjaJRV6nmm8yigGqTmCaNCjRjMq2GrdxKnYuv
h6Y9FMMdxp9flEKCWfyWMPysYxSVXggahBdkUGtrH77yQIv43EtdolVVgQsi6ZU2i3v+JMxdcaS0
AmQ9ZxgtsMRWVkxHBXectXfIu/OkTDsZ08PI+b9wrD7WHsoJahz26Hm1weOh2GhyETzGdzzjqOcr
sXAjWvIbla4v9QbwQ65wYYE8la+M4VyIExZYTxwM6icel/kVVrZyRV2tO1RC25cQPDTah+bWQvJW
XVL0BVCCRYV21sXC/75aaeVaUx7kyK5ms/P10TRlHklx9Rdqc34wl8u7L4h25/LlYN/vLREw0Bnn
zv7nlZXQoWD0nFouhxrEWMUxALuKHgbaGBkn2YDzz+UcKHfknOZvXxflKR1LcpFFmPdmj27g3kRH
0y007/Pp0xnQupSsnQC2bbE5k29e6yvcbYD8nGg7PkhTpGBxJcFkbdSAqYu8onuKVUeVYqj8+/LU
COFU8Wj9/4dF1Ph72K6rP9bKjI+rYlnJuyeHLeig2GS/32BrFCSziCsswV/65/Fw/hqn6H4Vgf2j
QGSW4h90qSVhvTGygvD7CMT07sne/yvcgYgZ4MwkhH5DSgspni6ooD3f2Le80zaFW9y27GlqJELO
/mbp3lglGjEAzRDTgXx2SwxDcAQX/RPwwZABU46diysj+nqO/UcbUOLztY6T61o3kZUd4DY5cRqs
NJTea5jr1L04bsCa0QRZ0oi8yKuwcE2f8/ysiP+DhZ1ThaTaW3RX8DmWy6T4kFdDccm++AczDwUL
iK8xn5hOb3se7+UDqWeEOc4X+cS/Ij52x3riCPblS73HtPb3syvxd1j4eChUtTles+oZxA1Q8KOm
GsSXg7oGSdg7Ugjq0K/aaac+RfI421Q1jardrMdeNVKJQA3r3aMcDznoILI8UDbPKJ42Zg6jwXfv
JsBwuuw3DnVEFbfOT7+9YaOGumnl9M8tZ20LHznJUylOaka4t0sXIlEFl0qhzB4RXT1OQibqfvw+
UHUXHAX4mLqehfaZBIXur5jBgt/uhKNHDz10FqRNN/CBQYLxiG88pwOb3b07j/ZIEZLu3HCp07ox
ZSeU71dN3n6rg0bqt+K4+RqK3WwvzVLKrtHJzdNaaMZJ7nUJEOC1HxEgdz1koG7E3+Vy1CLbquvw
uiGrFM/z8rzo0cpMSEMWg645rNhNqVeXBKccmSMjh1gnXLNzNEcn4vnBBguk4F1OU3GzKZlNZlCD
+sr3uisgc6bJ2fFTlOZII68IpuwvvR7TCUDcz1ftmmfakQdOdkZ4nMIangBasP/dAxD8Z9uJgnGg
q4oXgkr7mIBcwm78eFZjv+drNvcLXnuGTkv5JIp2jjwApgeqCcdstnQA8JbJ52faYzvNZfaKZ4iG
8SAerhE1+sZSiEQ5oSP68zsLCsWdXptO1ZtBGizFMuay35oPranrmd5PExj6p+1fkNndJLwCxsg2
ANItOBF9ZYsM5F7E3krbi1ljLrARcw7Q9TslB/ma/tK2eTf12WkRsQvH+q0u9360PNIu3vIFjshF
Mw5zL5JnLzxIS5YBUYmARmQpx+W0TBYmOIgJk2yfKgGasfBQ+I3pgr9CwANNpKE6tEKEAA2lKpHk
DWYL1ccPWftpmasQu8+zxxwaQstMYeh5qES3a/Koj8WuxlEHLAtsrX2O+07+Rm4Zia4D9YE60245
4qdCg44d0Y3azyiwR6ci9aUmtAXfOMR9/RM81S4yCsiIg+Hqw7insrU+Zr4HQStoEMo0Jx74abIs
zElJBl2Je+CT9dGIFgizU5Dvs0MCZoPD24VhC1o8CPfjg4UfHjvByYNTNyQ8H102IzqOAXGt+6Eg
0AElr4YvOFAPInjtzuogQSmxY9y5Jya0f/E/ivM0mMdZHLQGwYq6eFhqle5apRejae+rF1VF+ude
cTlQ22RUAeAYNeIPsvUQ9oPgdLGH2vXCy3aCBYAutapw0Iewau90arnaRx9dsqahJSUl4n6Us3zl
R9VcYzg08GUCeg+NVWJbZyMaJn4/XTfJIebcRUNj45DJWQObPxjc9PAtkOAiPUI0u/Tp0BRY6TRO
BDG6zQFUEm0ImSlV0rwaPdLZJzZkRjPfjL0BKoC1Fx4L5gZ8QMA5UXQ5CUk14O82YLOHiF1znj3t
5gEXWemp1uaX3lpjDEn0+Vcaz1QDSF/fNgSSg2jfFj/ngBDNKH9+os885pbpKvpYySUxyi6tz/RG
sL4jiVn6oYhTAi3s3eZpcIN2ZF0BvMjRa6VxxiaM0yiktWdStlfEM8tExsDOtfKDkdWNowSBLoHH
VDK+XSbFC2gSsSk9HhcHbZrTNBddCC3TefOILki6Ng75yi8mKbQ1sz5Gtd9Utz6QBrFLvd2S562s
Am8aom1skD7a8m6tH4V0z2Sut1XDabteNIbLA20GHKTWyhodZElCDR25KTJEf5RsNLU5M+6SOKql
fjoatKrgE6+Qd6LSSfO5/+aGTbbMZvW1Ihc0NpcTM2p2fwWrXo7xI8doek91E9DyOEiWjHRn+vlS
2hOKQHl7mX87XZiq5qFD2TqTn0qRA1zfEJF+cHO2VIqxYD4OLFCwQ4+85M+BdxWkMao8MQF/rTQS
fSTk7UqBp3jrR36K0jqdfYa4cjcCxXb/9UKv3dW1VY8n2HpyKiIrSajEWtMM7cT0ywtyepQkN4YN
EtgGZE8Q4MbBSp53awtBOepGrnhhcEEx+2ClsohxUDxkI6CfjUEZ7nauxxSUL7K5LU9OJHSJ154A
+q2SsUAzeK1p2HLZUHR0cKw6tjuIwC4ezPgj9cBN/aNK3aOx9+a0zQoSfPALfZFMKenhoj0n0cOL
CrzeNPGd0diAnuvpgfux8z2epPbCw/EV13Tz7Ah7OKuw4snY2GE3+tN05a8m1QYmb0fOYt+O3fBB
T6JhOTuDOvuSxsVoC73GhCAmE99LSEqSypn3wcOpcPcympUcuITgXHs8X7H0bTJXaulZ5ZtrOll5
Sbj7nahOTUB9YQCd60qQ3LdUXDhHtSDxyElzXCVXcmr5uMTtPKl4F5raQKspARzc/v94lpxCa8aZ
qJM1QFSwyk7eRXADqZVxkdB1zxL+DiwKzxe86/9Xdf2++7MbIJDNLSEAVTucYHUUu8UgtOADF9ne
TPjitldRzxu7g5iZpts9wpxeF4S2E1I8F9h2oZdAAqxF1Tr/kcA8zCIz7nXq7n2DSby55ADGu+zx
YP9V1ViWL/OWHhUdSFJwslEGaH4h3QsYTod7+2nQcz6Q6bJV8xcOYI2A8DbGQ/CiexZgUfj2m+kF
JJ7+RIVb1E8MgkRmrpimx6g36X3w9J408ECXYDpxYMl3ruCJBrmP/pTW+bmWyg5zRVuWM3OZ6irE
mhQig5WwcLuMne6swQR1dZEBM0ly/6tiSFvH7SCMJfp1Whdzh5pAve5DGoG/EbbNcAmW4YlLEZZr
C06zakOR+M3PE2pIC9GUBmObFS7GanQ+PluatJtFT03tXSSwIFZGWtk/oF1x0aChtvnbMpkz447h
3soLPLEuU/X36XmGBQyPF858nO6+PrABh8eaZ4to0nS3wQuvIBjlsWZOenOLFytJFPyeue4vImsF
5SCh7rk4jrN1NDFHwPd/HnWN1d6wbFBKJEllpUZAfU/g8mGTNO9EtcJP5IJiOdlTnj9VHcfyamKa
31PX0BwHyWGC4HyL/sQnAEP2Jp7UebEwx5hfaBhTngxK0QZyCHRxGogkaxyhvE+Tr2MrTh7Vqo/W
ZjHORAOeD3zlT3PSPpSbcYssmnSd5jlYkkhMX8fJoJVeBqocIJze5l30fDQMGNxxasMIFEUTw6Oy
LcpJ+dvAaQzZv8jNHtmZTQ1hlFz+OTb/qW4fQ8tTuulmUTnV1lx5r+a0foIPj4lmOQFk9ETisjvY
BIg7ss9/8C3SDUKE7J9yDIgsE8wtr65QqHB6qtSXIKqDUCJ82WcIn4U8EEPpDv20xfZFy7Aj2dH4
iaKHzcLjymKAMZEmVZASNYRKK6urAcNpJBaYdCDAbn+56c8BnRbfJXfYBlFIyeFqcXh0WUau4HjS
LcJGTyFvu3CHuAq6hoVRlg881lPMdaKUNwnRS8wyJgM7bRa1vNiolWrXp/4f7z5x1gcUQttBnaSb
fKV/3VhawDMGzTKEdjLvZRJ88B9Js9/hvenztmp+4LIw1ILGwnqBpuA6TebAA9bYF5dxgFd2qTCY
iaJF5+cXXP2lqYZ4GCc1m+Xe/+GUA7gPO956WF9Pfhi5uX4fbn+OGXrwPZD1eaKvzhgFjrgbUhiw
gfnt7O0Mx51urYOXMafAM0YkSU7loWPUKZImyA60E2+Cp8w1ZiEMwC+5rfQvBivOXZE+FN5jcv0b
qYJL6V17N9qdeJ//0UCCElb0bp3CgeLV2/IBEPovFhw5eXIgFHZSPVHpATtc2wMg5sAVqGXmpQlX
amYjL+iY/4YQ6Ig505/Jyf6BBjeDHMPPnI7fPlUe5hUhpAjdxusOLPhNNOQFhVLYNtnK+4fsHpOC
Kq76XvNfAdhioQ0HYgVBfvgKRzk2mJOOFLvdR8uI8Ik+V1t2WoMdjFx6uO54b/qqV4zh9OJ4WNg/
HmE3m1NGQvqXK+ZlboBvqhtfKFm42osWiycjkRJJoIQv0OtmS+vIFRlYqs55SUNvL4ryuuPd3FTT
wVMdXQyhC8sycEkQr29l4cvAYpD8si5UB0UfTYZVxuNk+r0J8CP5KE2Jzg3jRK+beTpRMFrAXKH8
Q6Fm/PHnlxIryUwVJ83Hi7BKtev12ktiXAq16n6SfPawzdhvK6lBUJdGauorufaguurgElC1/Mlr
lRKqwplJMu3m/ng/XY11MvXkTbla0vIWP/jUKmODgI471TJZxv0xS8Gog2FK2A83zbt2TzmwkcW1
MSJLOKFQ5mW1INZURce8RDYCyv1rgTTogDfAjEdQ5zon/3P8KqlxPiNTPQv+hjul8JJQL5s7QTXw
NwrqBYz1iJbu8fzcl2XQXmC/6FvcBw5CR5YjaZ58yPz88e48hsTwuDf5iCYCcfqnVdeJ1841AZ2u
WPgdTAHHmZpVyVVUi8QakCZtPFcJzDp6Erwo9xrC9PxyGOi69GgZZ+zsqJbepHWczDiRyosFmeaF
JONaHYQhPDQeiwxycvOb2jQ/HkUBMq+ZHkRlURD6OmIECW4ByKqWn0vClFiBX9rtJVFELwiT7sYs
z/Q1joUvM8B1NdYy9SK0//+GpA/WivfKFKelSgcryspAGZ3xIkroDih4Xmthk7fILt/NYuUu76vC
CrCAPYMaq9feS8oHyY3IRGFiChZ6RNCvpJ1hMdUX/KDPuCsCk5/TwGFpiiNR+ixCemgu30MjUGbM
RnDLxqHMv3s/ntEVlL2BMyfkpnauigK7PF0quiKUEnQXoMC1lpWgQMhwvkpMowjsJW81gyzAuiHp
cmxlQPeYuTGEybxSWzBoDoHyMyFzqf0goIg1le7elDcv7fuASYEJB8sRp5Pnn3dOwWGBTzjDhucw
Iok9K0dZSQwpWHqrYbEtXwlRXxFOABnx/VXv1nG0tO2Ea4hB9pG/ucPlN5imPg92+n75lAxcA52x
xV7TpIlLn+XAs+zb/8odMQ4zCOM2BnjP68ZvDh8FBmvhwlWOAvI87JT4y/KLxJywjZFpYrh5ajuI
gE60bYoQmC/LOWjA5xGtEc8qjVRnaELN3/kjnkRvRUGohbVvzScjd6ZKayzrwk08iR7QDtuNUonH
T7J9ZLEOdmN2y4Jac9DlwNvsoaP0k1FiJn0EqMW4gdU5LbdKNaSqP9hdxTvws7VeHjKyp3F2mOur
eNDGKiba24F6GoEk70/23ios5OCq1zdZJ7SgOUWBFOvnT2X2+KIyGu2PqoFKwBEx1xpcF8Md4JGH
6rb0uEeAbHE2ck1iRSuQ9m0DHFxgl5ZxE5ZwtepNma1i2uBPDzjtxmUIlkZAxIfPGhgFAU5espdj
2xumk0e9hbchVbAdBym9C7T+bXI6oOYRDAVTEz99L4tA4xoizUYzCpM9tPt+xSmlZwCnu6pqHvTu
YRVaqSjVq35k3VJcY/Uh0c1QohWbArO4V+KI+zsa/QV/j13eEz/VZbnkKOnBH0IGY54diVOsPHuZ
6S6oJQJbFsj0Dtys2n330Dd2q4J2Lpp2cz07HfsZATyWsYiFIRyDSNsIFPYeJq8/REl7GVjbzoUs
fAWJRTIQDuANjUy/8piNBlcF1qzFJi6UZ/I8nTHM0P6g23MH23sgvWTlPnGdXdFxRHgn8H1/3sxV
KO5hrynxJFAn8XPCthg5QLJH9Vifqtlhza1djKE0nb4ktJTsZSwHX6ItF7/Sdf31Rm+KugeRfF26
Ya3ifFxPmIvLBB7BTmTP+welZ/irNTgjnyNHGYuEnE+41IdrU68fgjfRXThasw08D7UqBhwp+n+V
1nyitPXslMXwkjwDTLxNlzFlyPx42wB+W4ghVLZXj5MNd/UgNImQlefF7Cj9KAC6N4SYG77k6beb
firgEsXBE2nt6GroTqDXYCRhd0niFKJHRuA9H6XK2P3l6WoxtMSeYm5SfW9rD80sJjrtkqglWuS0
5vNw19oU7Kc2lKIDg5WUo/6wY1ZuRXi0hsD8IlPU1Z5Mj39G/vg+EQCdkfZb8dvmifXrKNff+9Mv
pCjDT61vQUuKwRpMtW+eQPRXSepPLNkAxDhuQg82h2RHZrsqEzw39a3LZi8Mz4RV8hGHG29iIIX9
32N3X9opPMhlLjujXGgeknFs3Y2zFDm1vyGiUDqEnDRnQH9LGciKCm14HE9vkcfXwfboMi5lWDBT
QdeHYs58X30qjwB+aLlPTxHi1d+8PJeXHUa3t5a3iocvrlYU/R6XlHnOge+F2BDpJ6XRGxdbKwM1
WExISKyFR/++6ZaAFrEjpucH8LLymkmMx7j606WxyC819ZBfmmKu2TkF/DfpLQ8s9m8ICZlnWYQq
+sXLsekHu8U3KpNAfM0VV0gBGUl/p3j6INw9Lc3eZAezxwE+6N6mTCbpgpFTigfmDmk4sZIJ3XoH
f8A1Z/vk5qcOhRu+OdQ6VGmdYEiTMcuSBrdIw9uWpXVGbIUwo1dso6oCjL43QEhs7fr0+OLnvYGG
DWvkrzxoqdnEc2RI7Q7nb+cQxWt/2shyKhwCwbNNn+tb0BklPxhBkrWQUTT1xuNk122Aq5m7WlXA
4dN8FmqgZH1e4sW8e+6iW0XJv9XBVqBx6WpWBAZcB+8lvNpw+TrC9AXiZc6SR16Epdnc/lkLy+kF
VRS3xA/8AK5HlwUHZGfaF9BFl17nppOZDpn3o7C+Ol4xUsMyVFTyov+5KMa5mkio28RmqZTyrkna
x03mK6LtQ7f8CnYVonHFl/meBIXfqBg3zIL4N5/0YsrY28I6ik5qSK8QPO/nj4aSWXrPcH1ADcn9
09C4vzzijvfpKkumct951sO4JyTsf5HVOiv7V610q0Jt90CoWJz57jxrJaghi43fOSM+7tmAVtH6
5j7v5YNOcx/XGy30yv26f41Az2YRFpFzf4SLVgGH3dNxKTeplHS2H0yMqcyllDD1EEQl23SfoD+E
zB35s05DPGEsgjRpvajoacbb0I9BqbXmkOx5NZOG1yDM1eZELCkl37a8T2CsWAQ2Z4zl8kYuUOsq
Cq48hmwd/N/1f+UgJUGC9PAR4niZ/n3Vwul7oveZ3n0Elqr3EZsi0khIj5Qk4Qkj2idiTr8AyNnT
HpblmA2z773m+mTVImAwVKdcuuUgSk1TEGwxU5Klldj9WshtnT7684+GK+Nuh0iiocLSde7dy0PF
rVoaRAVll57mUA8wfs3yeOVZ7aS/KTys5Wj4OJcd7zb7jwruL4bD68fAKIgkl5QcKW/XyFdxya0w
+yajsHDp1jDdAIOGQJlGltBpNwbLcIG9LTwtHI1eTfDsR4HbFJApKYyLdzXj2Ie3WddHcRBj17/I
lrJ0ZiTZtzisRR1wD7UsIBRjNAjQfOhJnuG915SxXGAN3mdlcQPBVQgF0mgvxTOJIk1IlvhvpuVh
eVhVbdKs3RYWQVIxpgG2rmVq1rUBZtGOPX93Kyferzczj5jXTnoNsnquJlHQ/FTYH2LJCkZPEff7
iPqf3LU8TdbM6O1YFxqZBTg6VnK0QWvjluXGvlM/fcGN6QWvY/1zlXoQtNmSbxzLCXpCFMqRxvma
BqyNzC63BmsWaQDCukZ1q+9Iqj/2lln6EigEFFskrI/J7DKWNwYsEYzrajpUlvZiMxAkcZongvT0
2NZYGAE7pkzTGdA+otP7S1ylI2uJQSUED2UPCJ9lsODuXO9mm0NuoTp9dvUgF8TVxCd7/JkagImf
pus6Vzcyl0DPhrZIaSl3NnrQsGDg+om6wBZqWlRInt7vdzVDkQ7qaIVCNzOk7V9I+/QPPkKTQWr9
7qK0V2oFl5nknukoNU+HPIfLX3O1pON8aEc3M1KaIRnKH/VULP0F9jSzfuIfaLxV3FdnuXiZmIEV
djVaYEmxr1/9yAzVCEzD7TxmcT5UmbdmQ/nEZg4qCZD0qLIocvU9hczW0mnNTFEcZAig4FKzWiPv
qU41NmUkw7uv/SNxRrPxLGhZz2Ii9/iK3g8e206WdAqs22pWXsGQ4k5u2OTSGpYmcrkt8WwEsC+i
ldZuMiMG/eDFYDediuQNQfSg2WUf3EDlOy8UzoYBYjYpcDmtVlALCK+oUXggaPRpfqpj3pDgd9mB
+IXB79jCUyMy3bLfXHb04xMpfwRkWvZBCr2qHRfuyteZUaUoiWBOimsJL4qlKKCB1rlGwQCh9EIt
9Qh0pSQbrrjaO+q1wZAZBBkUVYy/Kv8shXnwSA93+AOfWrAZ9HBvhpWTrfP0wZhQrHbYyBFGMf4E
1fOipLSLaeQ93jYqBK1ufMf145QjE+LaPDmce0KTeXlBNhkCAD01nrHM/M+xEgkCKLLpIY2KjmKb
KmZYuOnKnP2DcMCu/yGt2Q3V+W87p4Um5Vg577yL1VzqcKALnNZUXn4qG7bpH2jQ/q38oN85VgsS
vdLmYlegWTYTXbV1rV2e/FoSzifs6DITGXWJX90DiBD70t3sJfG5WtN2TB9eKSfWAmIU3+LvIjZk
503NZ8YSPMWVyodEyH/AGTxWgaUnNWVdJBwaUHKzZiZp5yfMN2lv/xUvDBJpND3t/hOi6CxUOvvg
Oj0CZUCGTiEWvZFGNZuPan+J+bSn3nXQh5RPEadWnBN9pNWxqvV5oCJ7Zh/qtcwacgBFJzpTuz9u
ot8ybdGkFpVxJfDd1PeElHfsRjd94g5Ecn/eAEyZhXWFVX2HsT1fvJFXmNp2fVATVCskfPJsZJ6L
RwrZjoyTtxxrwsUD0UJ+yGdcqE4q+CR389gcdkMNMa5IiA/DMFkGhtoSgl6TS7dnV+t8KiMSHTVQ
seTxa9eW4HlaVzc9OrCS0MqKIdM2NsIMDL8P+ZwfqpOTpgh4HsJBV8U7jtPvRdCZSLv7rxr2dfMg
eZ9wZWB2aQE6IzF71dt0yOUiAWsHhqpBaanhI/wvz2P8ya8k1RjvRl6ezche2K+AmOUiOmYteTFW
DRweq6gx1ML/8ZLi/pzaYTHoltfleo7fvlK++AWsF0zRjovbcLUFglrB8AcH3M3wlp7y1zcy+3CL
HTo2jGRxdhLf5wprFsTCuBbxICXrZR/t75Qk03sow2RNoVmKguUGFHd+4B1RuDZz1wXCbO3VKzDw
KULjl6zMeOX+291LKY9Vbf0lCHCu0e4YIuo1ryDxBnxf5ureZdBTzFCanrKNlXEXWiddNS50bEum
O77JZxLPMH4Osy19hqXDTtpF9hbmH2dyFe6I31Ak8IEzwsTVd/FyK6+A0nIjt2ASMlKXXpNeW9Lu
yIkYMFrCo46a82cVcUoUoxy9G3uWi376rKbY2DkoiC/7WhhaLXibPGxyvWeiSlSdPWWqW+Ee7NM/
fXnk6FD2JpzDB+pyLO2hJGMG2J3LyxF0QVut+EsUAFAJ5Gou7TP6tUa2laeHH27mYxhfb8MAoUbz
mhX8WSTIt+10lKXDc0U3AbPawuHHnkRjkwdmSpeCU0pjWsxiKDCMzf9xvEZoF03e7uNTRArFz3In
+TeiFDcGcGnRxZ+hI0bkKdtlzAPh0m6hMwCIt/x3S1DJTXCTJcZOJZ9fXrmTtyrwBVmyKP8D8xQr
FoWyMkqQo57xmDa10s+45zHDw6Gq9QYPraAaSv4RAecpSZYcOhnBo0ienSGMr+Z0o+5FYIdfzsgu
RlYVcAbbzTxdUD6obsdu92drVfrtS52AxIaoA8OCmsX5bogrd6fOSYzyswRI3gQmqJyjDoCk3S9I
2ens/CeBBZxAd+aYhlY9pKDUeKkhlkrHGo34oJ29UfnL+kfcvzrV7KPc8LPY08HPPjTxgByBha0q
JepFN0KpGkUNoqjbTnOEeIYcW0ynjh0u2GSccV0RHT/6TWrbXgv9AOTK1RXxkDADMWhUstGWoGcV
Zkh+tJmPnca7v8lDkp/NwVCbcsQP4kedCJU5Yuc0SmfUk1bZHr55bLw9/ewBakjsK/Ktzt6KgAKP
ZAoLbeI+DmKtj36uzCRkJI6RVmYmC5/tlgiSTCRdeKxipPAQdmArzAz/dcO8CVpzq3qpUFwZyYE0
mCEPQseRv3JUP1hOR+udZAW8Z04hrYojOp3+50jaGgpcCazjrGVJofXOhmIFU4Fw/yf2TfLKi0v1
vDcEkZqWc24cxmA7YbL7wfqR0cqdJVihiX7r3B0v8FmFRhoceks2SLOFTbw061TNEkXnSIhJw/ye
cyAiQoxSwyivo4MmIj8KZQOV23NOex1SadAVpQ+6wyV3g5TMWvXcjwqWC1+HjS00zKfIgDZDi95S
HBNkLroYS36zXZPlA3UrJJUG7hAkAh5OQTlwhlIbNOa885QJbBluqvZVefVvzC+XzaOSyOlMjGLz
bBH1l+2otWfrZpftUKkOs6V6EP2gAh2NcEhrBkmxIJiHBf8QEDMMCSLsyzKe9OkY9IA2fh9J5aOZ
8llzfowYUbCx/VJ/hRPIrDdWREddlQ/agvBQw0zqpK0+lCLtZU3bdKi25ufBdvokgqXLeGO/lKmx
+FjgqDAV/nGkvbqzDBEMv9Gl+mf5cm+QGkgYMzU8UVcsGJyRL8x+u3Oq6ydJdvMQaTAPWRh7S4nE
S/CfSi/eL3JedDgWx+E12/KwTJDqXRk24SuvFsoCzb70sqTnGzSPB+30L6jzVhtvrKS7gtp+jOAU
G5XWmuKyhTu7iDnhAHPGgvz/+u97pEqVm8RS6z9rRNsqRpgqUNBfOZE2ZtDjybB7xUXsO+OFosu2
oZlrH5BkRcIzU4zsL75jsotUR/LNJstnMKmfIfSArSsUlJl6qU1NaoYZZ/lgcIVR+rxo5Hn5jIty
QsAjlZi5XzD/35ZFMBL1Rc30kHii1NTFe+Tez/RaO95hTgWX5REOtODUSvEUbe8ciAFhJ/9HdwsZ
OLKC8xLfLG+ILO7cufup0Tkbw3gFBO78/GZU9Yr9SS0seL9gLEn59nEVpC4b1pfly5UyJBp4YW08
mXR/0KbSu1+9oMsxC6JY0OCUNVZrvIiHkECuz9iouIF5EUBDj6r8NE7oW+ZZZ9asFJ4cchLTG1Xf
/epDsSFOFw268JuGRfaeUPnOLfVvG01lbw==
`protect end_protected
