`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
gGE0LEARv3arppTyDOrehnuYE+VByRdAR12tUhZN6TDzxj5/W+PE2qoxQu8aQEQ5QjL8dgL2rI3n
8G/d8DIPNzm6cBgVc4BHiWKMcQDm7buLg2OfpY+ecrTwHVYVgUJc6weSVY4jqOvhxSdkENeqMvBm
c2jVExJ1fE+aO815/W0Dgh+dt+eeacls5xvYW6R5SvNz3lRER/SRZfzAwfksGQIqOfkFBnxKMHV4
aHWk3+HR7tAhdXtu/DUgMcil+h54lDZjwPbFPZvsAmWEf4ykblAKTPHDt9AW8lKAYnIDJeMORqaV
RWBEDsX5Dxc5gIhHUIySEl8h5LVjE4fXnW+AQT/TI6ib8N+Y4S1aYQdgMWq16DPOTu01j/bdNG14
7xMio0PTAuXSp7Z0B+10NRx7r7BFH6l+LcpjIZQhWNEd3ct+xIQ7jsllNgBeTh91FJFumiUE/wPD
yoEgD1kCrr8QmWHhFguVkAppKkwJCOVFPY1zSHX4YmVUUF4MM2Xf1W3SIzM6NXKG6DEDU6DPsdc2
Tqk2TUVevvlToqed/PAOzXYYGQ//NtXFPaI6z8DBLTX+GmlkDcZ2f+23+/FJbtqTSg1zdhP+vxNd
m+N/lnNI4NY2onYSIzuJsH4yN/AhYdoViDn1MhV3npYihWd3FmSINGR2dqGbfJ3WnSDjzsDBmVLD
IDtyyPgaI4mhUp4EiahYTH7uS31sJ0HTNZarxV7zLrPoegD+ia0cuYzQHpC4e54ha8OUiTO5tHHW
kbssBxXPdJnK1fB/pYjcp0vK4nhrK8gypTobdQB7+aI+puGSL/k/LqAAS1uHTLqlbH2lowH2SQk4
+1wBRwuHnobN4Qc63nfBcTAQCIET4V+OBIWGKdOcBNUlTZllvvpWfxBbLFlHbYVnpSbCTpokmCZj
vixBgJLAs7ms0uz+0WQRwuokHrBRWLE/hkzPElnyByTiC4WMkMQsK3MaaBU1++Ts2FK1H5zK770z
Q0SiGHMfXOsO9PQmOSB62VZ+IPLioCw2c3RSisgNuZYbJsDREVtWfRRNcJ+cpGpX+9yz59JwDy/K
rylmsteMZvAJXJr3PcYuJkWi7IyqYUNEMWFFTTxQQ/4bLg9tJBMqkvAy1YnqQxr3bXb7x4a0vEV6
z28nXTsSAS17rlwKCBNEzpiUTZ6rnxr1/C224he1RwjGy2/BOPuDn3RjCmco6ubY+J/NAIPVOeNp
mZxONYK9iDoQ5znsv+XYP3P19zKo4JwxS0KUcUuYtg+Z67RQBtyFk99dlHhy4filaA2JHTQL14zg
uWSb8o3Wu4SOqWy58b0zd5ILt7vHALqYMGjUSoKnlj3BS6y1FNGLH9OVDHGWUygr4BI0737nTdjJ
uUScGPQGx/ReMRwTofJw+b+uvTZ9U4k+9XbDgAsgWD3nlwXFbHjftbuy6YLANCmIq0yF7sID69k9
FqWOUc8QIEt+GFbZh93b4aiygc3zCqKkezt4QvZMxEqGP+BB7LHcLZA44AM5LJ5jjKJLOxbqc6EV
qviPe9SpBSxLjbfUY+gtHiO8WY54/FTdO+jgwGfgELrMqODztkdnnLafGVknVT+zpkBoQ70OqrTm
xIK7xQfLdBJIzmJhtwdZVxExcyNK44/zOK68qxFRq1EKGu6JZ2TYeBNdCAR3O2q+Nnni5CXByhVR
ty1ujd+mxWfq/VCBc9a+6M0j5Zci1/LVmJNfIAlEc2JnLXN3rfCrMTqwUwbrnmIuEyfYtbuZOSNd
18uujEFNHuI58MwJhftxU4edmtuVP0/d1U1eOW0np0gYdORUProwJpVUz2q7pwjQQ4C8N7M0f/N7
XUZ9z1UcH68lZEw6mm00vVMMJ3w4Cb5Z+M2efdipU9f7QnO5ciHH7ZpfnBcoZWfphY0WSv1nu8m2
t1jFgznEMD7QWuqjAI4DfxFToW8THer933S1ywsPT5c03QQsHXDKQXEEjYJlN19D9IIsB12sv6R2
WdVnsQxS83rDh9x5VxUxV7G4S/qkfxGpI1SYQ4oNXbcaerJAXZ4bhTj5sl2EPHfygfxUVrcy0YkC
71+K0VWzljQehFp3RMok+05z2oo5U6G4JOZs2HVeOfig6B/0qg2B9seudUw4n1aANkrbIMOklCUJ
13ITcl6PfFlLgI4J/xZeKrav+Ki6KOKtUTAc2zEw3FO6RN9jh7XNf1ne5cHUKV9bLegAlvtEI9lc
lZySIc+TWKdVDfRUedp9YILAxlBw+rdcMgotoJh0OO9z/jHH+XyqG4ixwPCX4K0xZS3J/BW20itS
Yx8bGJSBHVKQt/HbBw+yNF9OJTYWFYAQZubCYVWEW1vcxA2S9/c0Auw4lOj0NmNLRmxxA/XHt9Rg
MS+BTn5bLdkJArkfpArT+RE2JglGIm8LY11GSQwUmFWnjYYwnubuBKcXwPN67Au3Uh5PEDZ83tOp
YVuzy1wH+PXrTYzW4HnspYn6P9V9MoWKz83CCcAgK/aVuBB3YFi9jYeMgwCSgrVvBuEXJdKeIXNo
J0ah6v82gp+h0d7NFUnqnZi7KZ/wmyqT+GZnIndoMMk3e7O58Hl+dadQTpk27bwn6ByqXhP/YWbO
G/u3+RkpGyrYtDz1WChpk9E9QN2kMGhQV+hu06kDt9BckdjqYatmoShg+9t2shHQIBJ9nG7cKu6g
SvS0iWAbhM5jxj90pmJzRJ/k40jmmhjjSe5wlwKSsO3GYklJ41QdVcNeq66wNU4qT3JtBM+aQSTH
g7qAeGRDuAE1Z6hXfZgfVZJiLoNGJbaUPPGIB+NqrOhcpJ8EpbijO+w4c+MhxZ6w2uroH/wG/8Ns
o3YK7MRowpsdZDuQsBsxtDa6R4aOh3LF+iVHmdjZIQOxLLmY1BAeahTJcU+ptSPsZLtQX7vr3osX
AWlqQ2wuYtsq2IkBcNVcQhRHsDC7hxIG26H/J1RzxZyS34ylnN4fqzoFZklRht/pCQlwxy8ilLdL
Ol6WQQCwHyCyPhl7RGCPFoIb+0fdhQjYvmCN2oN0fTnXGD559skNs10G6OFEq82XF4urYsNj4Izb
79XDhsCD75qIm/MF0MdGyihwJtpuntC34cARW1uY+9PqBLOrL6krB072b9pf8CJqQoUD8ZwyX6pL
6ctWXi8ERyqIBbAfRf2IfHBuIkOMgGfd+DCW8H2itKcsXv1MrTP9VbhUZFnSUniFZJ+oZFaVQYfM
Aw8+QFgSABYu2NO+1Wm0PNDwghDCOf4W5GVnvUxiC+i0yXH1U6NPumK/WZOJtWrikBtOIbMNzYA0
uJsRVzmjG3U9eOHvEmPduKHRm8h1/X/+l+q17nWUg0FuoPElLy3YPe0az9RrPD6slUDKx6RnHcWC
ixrln/35FLKxvvoVWSpi5T7XglIGpqR3lz+I5yr+S8SEcUF+Nv4PgM2/Zlm8t7dV49L+Jf5sbhrn
pJhee+iQqSGCzsHDs+5a9i/Oc8NNkDP5ffTSGpfMC4feG95aKU9ZfLBfe5bJSKfQvQliVsoiZ0rb
DKiyn4/bbveLCJvQpjItpOB8EjcjZ/b7qLEOIVviJLcWRek3sHzlG0XTi3yNb5qrFBtDCWRl7Y7l
9KrEqI1ksQINGM1PauaiE+jYKFC0Dw+mUJa5J08HYhPQGwX/Sy+dPuflCiyHS8AFhBL38hXuz41a
2iZ1Yh1kAuHdbv3SlxCvKb36OKYW/WREnS+RoZ72N1MJM5aY6k0XkPF+QBsnElx9VZufP7A7UdRI
wgJO/4mDKe9rvxoolos1/oc6dbQPiTLTsWJYwf/PFG9yU+yiGY09sq9WLzcnuoIQJfyfdCyKWlyi
4lFpz7Fd6h7gJCCrNwbpZF2WVXAn9QNK7a7VV4sE8IvCfhpNPqL/Hga0bXjG70WNIvv3XktSlJSB
2MHGR9/843UW532pdt196BhgC2wGHN07w9NXm+sU6h/V2uy2b/3xorJYgia2ncPJMQMJuRGTQYDH
vJpInhf8SVzNxCc08sWNSHK5byt15OLxNO92hVFmgUlvBjjSJwnXeDJeY/WPsj4fWJrOP2NXSFVu
WoJsGaEbxKtOw2W399WV35fyTcNiuJL0O2ch8n6ZKacMA7m+O4QV5VjXlWxQIV/t73VLT6GJAxhZ
CARSWrzo2ELdwzr2UuhiR4rVlVz1GzasKKpUO6KZM+BrqfhPesYJ3JWMs/aifpMLSiocVTTXOCpH
ZQEYDcZWaFKXKNYIK6xCY9rWiTvJ8L0iNuNf5ylvuA64RQIkh3g+xWaQPU5+ugUa1sMshmGm6KJW
EvVC9CINS9P+3Y8uHOa6g/IgZXpjbU1Gw1afNX/9TdsCQOLmNDI/6YxuMACfqP2SI+2NqeLrd/DP
anOjq65WvLl37qc7M9OENeo01MT1aiUw8vbuFRdWkbbLZt/9Um2AltZNBEEvTMTjRTGXO+CYtEom
SUJwQhoNvD6lWuWjtm9iAElfqgZaymQRf4fKQ+kAAF+OiOkFUMSoMPHtBB8gcJsvTQVcnutKfTuX
yMc7lJlO45bnsBjIqPhH1BS138U9bH11El5w/H5huTNdLTUW7KXOeyfV3/fvkL5DPv8AIWIcW4ww
Bsih7jXz62BmJqZ3HNe3lQqbzAuJhiK80Gb/oGDcLqCwJCdnBfCwu517kcu1rqxlv/XZaxEY7O4q
WuaF21f5+Lx5sq3l1+ldljqq2yrKU0UiWU1lexPwIMsrj2pgB4fiB/89Wrh0KGw++Thmoy6uIWnq
ht6rlKM+N6BR8QsYH0T3OrTQRxyToSXhIAr8O9TrQ6xKQa+svPPS3e5+ZoUvW5DpytVMXDM6F3Ug
MpEwiJ6eIrc9M4ajBfsdh9s3WA2RxjpGheSyO8lrHkHVwjuEJI0LSIw3CerabN2SY/dte5WTfkl/
5yZmXMQJ/rJPt8bQ48ktDcI+zfJtbZKu5HeXMdA1QsnguhmKDAZqJAS0iyK8vKl0QMn3ya1gmpKQ
RYA1KtlBnZOghvL+9zpryquoxUwJSKBL245D/1wDCc2YSv5Bd72YxEuA2PhIL6cIjjZ9wFok9/Lr
y6hvsDWpJURglXtXTSHS0UbR8ZAY5gJ9dkzVzJ7bET4G3+ij1hB3jb+Z3+Aq2RbBcjsTbV1RnXfM
uxbO04cEccnNzoJQdxYI+E4RTa9fN1B9pYnb4NGEKrSSkhhvZDDmGAxX/ZZGIcQQasp8zm208IpV
jFRJumTJCC1mQ0kOzvAbBLBiIxoJRpDwVtPLeogLIimuIK7rY6M/nyKTUuGOX4CakpK7ioQy2bG9
NtrDcg1YkqSUR4Ose92DMIs1CycZ05QXteF+Hzbr8eBGyUsiqWaykffNtPsoF+UjSPRhX66Qhli7
5VQZ7KKQlZhmOggCt7OWdgOLq2OmTbncvbp5HixR5F94NM6bSZIutqO6qme0PhohNnM9J1sNcxyc
FQtWXB0HJCKO7snIMf+dzZzWTDi0AWTr+evkNwiA4zHc7Lf6SiO5ffo0M84+MQ8k3K70L0G3QxnF
bsVk6jXU1TmNxzAS6Vtegt35pVM2Iq7AtRbtDJ/Lk61dp42yPgxw8btOUSjUVCvLZdA7EM/onVgI
lCEXtypPYpmiE3LQj9VT5I2JWbxY0r7A/7vRI/lg2ZV5tboBZuLQzQoP1fu0FPgzcX//hR3Y50uE
lSg8TZApbPkotLsEEQcsKgtI67tI/AZRv5wzyVh5egbzJsHFoQj9eHmLjzMaAB3192zbjKj9GqyR
jinIYYklqYRLdCgewEwX5nTdIUgINC7vHFJRY7KQLKkjyaI8lOvglqCV3gHqbrvb0up72Zv1e6OZ
UtxuzTbjwyc5vEjB4xhM1vYqnu8TS491TXsQBrIMq8IVHS/jKIvXdSL3mPESTDD09Z1daASxzjOM
lE8IHozgR5RJqFN5+1nfosIqVCVTQ5Gi8idkmXxoRoz7FIZ/cfx9UK2A0mGWRhH5A1bAAoEr2c2a
ZQcKJl0vmBJbSis56EXOGu6vX8VM9Qw4hQSwpeAvKZjE9p6APJqHtw2iwkTnaQUmUCFgq7uPKfZj
DsBGRE6A323c7qNyqrBPfIPvukDl1eBx2p+dkIcJIUVW6dVpeGw5JOD6PWESzz6EbpJJGWqsRboB
nVwpgKQREAF+15vq2giq9/UrQTffRkm0DgcKF3rl4aR5+7P9yZq5e6aLLAmRIBWaH4CJmiQhc/YG
DPylr4w682FnRT3GgE0zuudiBU9WOC+k1oYmwHjljwL9sR2ZZozkYOej3OrOJs83DeX50mj1m6ti
uNAlt7KoHwzGFNWkhxJW2qM5gdYPLrZPgjwisSUxRhjzBjdMP7S5HsIjDDYxugwltTnMXwpH/o0I
aGPeTfjmvfY2+HOxL0g3tWM8S7Iinam7+8YxIjnyyhea6vyGOmJCS9mhQnp4GJlxhKkEIINtMLZQ
iGkC/DTeZeUfFm4Vs8gG7ULhrpdW25YxgL1/S7hBDLpZzVlMHNJ6oczWKTCV/6jbt3f64mpM1h2Y
rdiEkKFFIg3IlkIV40eLzXKZMArh/Ad9AJ5sHlvu/0JM/ZKHDaCl8lfsTcdsIgjfdzXtYrAI5KJK
FZQi4D0hayxEWoMOVtkgDKuDAxk/yolwNKL7MCQcjc/pcurf2lWV60yFLj8PHhmksrirFCdkN2U/
LJjuMs8OHNaH9sYIu5UPKGJ4HHxqKTfsLdAL/ph1Z9mqLmjjPaYNPJBByb85oxgfwctMDg6vMMmi
o7DHv7AppC/Rz+l66UnzLOYQ/uF/4qzi2dH3niSggqsCHCB2buFQfcRh66TBA9+RS0T9ys6xEuMr
lT/LqeGheLROAdwjLHDQ8ak70YIit78lwnXfzr6aH45ady8X4yeLmD3xWKrNwzkDg2sFxGJaKz6/
0LheKQMsdUcChWxQ7aFml55aceB/z6rVnxYGsF1mCF0ApdS9aqIhrKGe2jE/5BvOMEd4j9K/YpwD
e+ZKAAY+6zWS0QqNI2FPVG26TSqBeRzdVNNqcLvkdqxA1aJO0B6QhzrfkwxwtCjTJ/qscnDhX6W/
FvSNM76m0zhBPo1fokN7Ts6NXhkaHNkv8Ult0PfD8GP5dV68S99uIGRlYaGAIy9avHcHye7KJi83
1qy+vTAR/yBFtznmVJBS3HWU9ys3v658GFFe6cSvutkFDXZlgHjcvjNimmTt1tDVr/FaNPrOesuJ
YalKFhjwchdqfVuNMU+wbXSfBawSIoey4Wz4Y39YKVsDZPHOpw7y0T1FfetNHEC/QjiABDhUoGlA
57wdSQjVC3J5Gb01sIiWvtf4j+V4NnCtByq/xHF6zfaxR1iY3uqxYAEyDaLHAvg1ekMCcwMtupxQ
XFlW9skQTbJ/ihtxKJSmk+aaXhlMzE8mfGm7mdWhpChR4d0m7zq/AjUHKwtZ1u0Sy7VdRapxxBnr
D/hsWl/NYY2J2sebkIfXsrEFIG/9gJ7SKT5mxYnMmWjTxNHvQ3MuE6tnG708eS3mwLwAJkbO5fdo
yE3CHCfpCIE/T0LmfIAqb/BmJsczqcN3BR8MbmMWtC9iL93zBeXSoNhiBhmsTBYDXtPgKd9ehCiF
TiNhYETHfQzn7hrPpnitjser0qlvnKc2NHnrx8wXYzB941jtBLssLqUtfG8no11BtXw0SIr8/Hqg
pxSgZg3UELZuhC+vEQgQEuA7sOaxZHzigliS7deaA1hM9p0tn7vPo4DjODjyoNghLNxCgJ+Apygn
GTwnMX4YOXzj4NJxysrIxQcyOjv2uHQP1LM7QLB9dV4LyivfDYxk7dJHIyY2uwvqV9qVTGleqhSi
y6DLFurzQJ3eDjmOmtN3gRKKU8P/SqzJFxC2GNyRcouhBI5CMw7wqcbX1PGGoOSByInGxXo2amd+
prBkNroCurFeaKIILqPvdpM5Be6eyTxgTuA/Sdw4ywsjnOCEV99I65mSmOF3jYar6MJykE284sU3
eBU7owp0nuT7p1TW7IIr8l3y1u7VeNQF9Qn6C9BoR0wnr77xlzmDrci7fyUOpeS3QGTtV3IHWazS
1Awp0clnAyCSARPqOVbxz5OD6J0UwGhRvhkK4cT7NYY/vutdG1ubWa+OAWl+KimAkMZDJVkI1rKv
Hh8sZSXL+FZKAdhFrHM6mV212JfjYCSvjY2Mi/4JLfADVdZGCaU4JLhMyoCx4kHMpYDlsqyoFwRD
8Bb1ctHPRnkM6uBmaOrj5W5r6qOR+HXHPR19V5TqVjg8O3vLrIj7DAokra7MeED9+rL7wo35CjYu
uKENBUtZlaain2fFIbfXfiDavYV7eWem9WCfRXJr9vAUTcl5c5wTFXWK1Td8HajcWm5Hzwy0aEgJ
kevDVBJ2AvgcotTBAvK58NC58Pz0lrjWNE4iVu1+RjJiF/qw5QwGIQ551bgf95G7Lczr0BhBROLO
HhAHqbWdiD65MG6tO2FIZTZ0jjeAEohgQFf3nPU8NgdHL0Jj29rDUnJsJ2Azd6xqig0T5KRyqRPO
h/S+pVoyCKxZN6p07AH62kTK0kr7qtgQLJi3aJrjleLlgyg2B7yVAoeliTVWLzXyq61sfVy5RRhM
/i/rmU3QyY5wM+m7te5RyjsaP+BLYI1tEmp3mGzNE/cHUXu+U90mkED4t4TZdiQgBqeAqYW/0Do0
gx5jdIzTF6WL8GCq69nFe2f9JyEKfmoJgmxKBDQ2JeUqFDyckVbx8xT4gDohfUUOtxnvgGehwH0y
iry0wn+aJEmTnrztkxzXxAAJX+mXHzXVcss53baQY9d4nkVzPk5dohclW1D3GIXsBYE2RGg2mGmc
ec+wGYH/KXjlIM2Ptny1XdJrmme8MErAyIBCB0jh6oYzMeUoolF15fCEpjeCOONZ03UkCm4g1Kl1
i6/dK+AGmUbo2BWHQZeMw55VjxD/9+NqDbrqBaupuWj2T/QK9Nz7RRwkeSSqH6eI1J4ZodJzTMOT
y7MCte/nyDtAQ+ayU3lOPEo5KT/slomxsKzLbYQz78l6gl6Cmb8CU7GuoYIBwVaKUyjlqgz9GhJq
ldWHq/qEipaV1hAPVHcwqfUS0NtvLgFy+WsFF/QSGDKJFmP8EIZzjQNLgwBN/4wO4jZo89o5hX0U
V5XXQnE2c7TuvACfY7ccz/h5SsX+1bUKYbODrvyQRmoaudF+rs283+Ujhgux+LEfU8/nKRh0FS3s
nONrD3Z0uANKQ4gXhAl2FUPSfWRuq4QX9vfl7/2yh/YYtu0M7tRKFQiWBjUrEr8zAyJFceksMeku
voYWEzRpszvT3GWC8XEOFgY4JoOUgeT+rNRvKe5qfxJlYr3RukuyK3C5O87IpAaTLhTryoNBeJFH
WFQ/9uCgUCkDFDOHbp7ozy1w5G+acYEjfGAc2lztBSCY7Wmq7xAn64v+UnBDAKJi5HQqDWUokr4Y
AiDNfs+P7RSAlEm3xdZm23r0flkqt3VbBQSk3LZTTZdIbp36/KMfHjVZVqzJ6MLijMF7FiyjrNna
KzG5Eadhgh9KrpC273Z79xgVj50qNYqOPTenK0dTwiyw7Lf8kh05qNuCgl2o0jAl7axGRy6dk+jc
E0r0rpApNn/xlNs9m3a1WSjvovj5KtW7d2N108KG/H7JgUsq/Ki+zjytloscsuQTYRQQ2FVuZaVH
JOfjPBWBoGgx+XwwikTnCy0mEk6HmQ/Fbf18t78fMW8I83g9e3cpMI2oJW1hQBC5AmSjs1tCkm/4
PDuxjUs3Erj3l1hjU3fk4SLrCm3cYFrteJQO1idfZAxHR8Tqzueb5WCpwwzqMw5JfVqJtJ7j7GQt
4uQRc5fsYIndJJ2scLK491InPTwevHzokZRa0yLKBzXrtraFehtYfBYNSb01dHkq+RTgQAsVqA84
U4ugWC8kKqj05CA781G0kzWZtFjqeYMe8fYPo+dDedWAmvRr37S0UVn47EB6dM8s7n8r4bbXdiEC
edFy9fVuCjRC8DQuyrVMhE77b0Y7LerdKQONBk7tp77pWtIt4WdAXiZ5cMpQVcfJW/8nDERhbh85
eqiwhUbFtW5fG2Xmus3sG9r0lATdE7gKW2NaqXkCc5Fn2pUyaqOEamhJiJyZOALAw8xYB6WmbuUc
TwHbFTr8Y9mtz62OZ9ho9NzsoolN3qzv2Gzw8L2Xdjui8w3qaBr/yML1dmyQT4o64gQydvn6s4xj
ZfxPRNkBIJICnuTK2hpC1l98J825QPcn4IzzghxMwYHaNmfuagEH0d5VrsMKkt2DmbQjO9yRcs2H
rh3zOELL9pxBSSFQQi7ntlJCMAVa0UCDvXYHxSskDenitx4Tmy3sL3Ehukp26kz1wDdYPylFUaiu
UAp9yy+uZbHDOKQM8SSTJpc0eUAggSd6R6IkKGB5U33atn81RTPqOgLx5Qln4MOhO7Oc+B1peJGW
IJMhiN+35EBHnQbyDsibnx4R0cbxJvfuPb3ADdql87U9YwKbomzH+KEft61gxUUNTybshTWdnRlW
L97GVyAmC+kFzU5LFHatfeb52kPK5hhnGex/8SBihz2mjtXXPKJCKcfsjkLT/2Wm2MgfO3JlNoya
36PVThBddMzH574Pr7kWzthr0PFcVbtsYmzoYjTQmvZ/4LoFfV59wpyG7EzMFeUb8DP6ulwa7Wb/
tZjogbp1YXHLTVzhVanrF3FL1qEmb0SMwa5LQwYaVwzMkNrr43oxOolMC8FFCUnC8DcA+0t96tSE
nUMY1aKjPdMHhZMq++zr0H71ZVHWjN69zkPsYTdSfyXpwgT18GlfdVhZjC0sohbnTTgf7cRrOhg5
lrYpBah8gwxrfj42nmcwSGCA08fyIdPtqudXF8Ut+eiTTzxUrQUWVRKdDxi6ujPBKDaXDvj5ho4p
Ujw5ZcGELk3eE6GqMC7WBd/oizOfMCCfu9lc01EFRF3IRnCSJQ218slriwjixc41p5LY+zujKWLs
BUWTvzMnkLf9wEmEcHDOHaxe4MbA4NtpxAvpnSMWCEkOsNXAJ1MZpUO0CpiCqUgHyx4gqI9ZeipY
Mg3qq5EhRlUkF2IsUFTRV4IgghavjWeBG2HdT8k5umn+ADzhXGEt4Kt+rlXR3Jx1iAXU1PDJnYNR
Bccx2gkTzsEfbL89b0EZ9XS4L/Hrf90Gbq194uu3zRKZt/5Lhqs7VlDSTVh18QdgaQew62bmvNM9
rYQqxxqCVfk1O2hwuM9kJIRIUW0A01uODNUX5dqkh5l5ZzzuV/uPfOEfpCNt34+jyq4h/N9j2i0c
FvsRIe+ZObnD8P0jKiPQupkw4IIyF5DkazCBeBYGjBUgGot3kHX7pA3UoXj33EOBIwTPp4Z3AWel
ldS7v4ZDoqNQ99A2v0LOGnTz1DoVuwWoDUxigTDyeCiitrteYfP/vxgsr2/ME1Vir+jgCZfSclgq
R35MenvugKIL4yvfh8Atf2I0o/wNd4DNKb/zMQZ93k5K+fGeZkWY+kbgfow5lwXvRxNRa6b4dAJl
r+7Q2ii5rNCfQtThMdXaAAnHuPFlMH72CMZXM9AdEXhBYUgYuiyjaHtBZ37mi1cEJWGsGMgRG0eX
kasZeXBePYsosf2NcVfmn8c9/ktJSNR3Em+jozCvWz2DGPwAF3nUW6KN/aAauPiKwqvRaEmv/esP
2RI8QOJ1mN9OBB6RW/8M6cdnzx796rpu9h0PDOlz6kYgwPpJdKZTIQCVwWoW/vwwqAXbnm1aGT4s
LwGjt4+K7yR8ITWwllwVkNFQHal/TCKBaXRhmWVJGL4OqXu8A/ZrHT86YIM/yfGY3LMd2LccXWGs
TOJeGdgcH5/hVgWKl/vm6bga5MiqLp8b3OxY+ebSj4SlvvCm85w0Nzn2vjBye/5pR7DZ2W3ij3at
lxdGO1927LlTqtla1jrQa+6mRqDNm75KO9JHAns7QEcabE/5wL7PIWGMfW5FlFJqTKvF623Tc9s+
drN22Aer1B/huoaykeFGZ0grNW+N3h9Qcji0ZbXiuJ8PhQFZlY1NcJoi8dqqZFpiOoLmO+Q5wCpS
vMzqQWt4If/N0rimOkQ8HI6Yl6Snfp4y3NCQyadAbX+T8so5zGl8aSL5aLoxygdxAR0CLSsPwlCV
XbTxQa8UOhkl/9gMH0hu6GCheiWDeGCsx/38fqWi20nmfwy/pb4H55I2kcu9VH7IEu1jneYlaN8B
+cTNbPrjUU5G1YUbeCa0WEr885Wd97QJZPDsgtGuWHVyAkpaUBEiJA86jSjEMq3j4PgPTzRnUBRo
abuOhRAaH2RsQG7ILLFZGEryfcDe+MlSZO+fBdvzvJsJgBmRD2dHhLc8ef0bHboSP9ecQNAk6JiD
k2fNyqXzR6J4rWjt0I3kRgYHt063ni0820orekkA0fEJGZ1fmBO+G9o9yIQogVExfffatzOFWy1z
f9/A7OJ8axOMRRjrXD4UBynYqmIQJIqPp2jOomhJI8bX0VYOEP2KSGHkvlbpXsEkuXjctAYQivJh
c5RKB0UfcmNGHAhgYtpT36Ke2qo2xFM74gV4U93erSSlAy8P+L+i9C5w1SUbMFSKOLbXSVLRnTgY
Z2jnZ29f0AzBhVmOxKdepmFFv6VVGRmsF6/PVXqn3Vs7Gg5DYuvHs2RtLClTmPgX1gOXHv8txj07
Hko/G92+gPbKoKfwOtd8E84mFMtpBK3o79ZmMJibSOwaWlC+5wtFNR4ZGvJI+4vi5AfaIzKwB6FV
a+ycy7RQg1kj2Q8y+dS+zpjEdQmjfyynRarh4MpiulLJDniDGGVR4PEqOc0SVQWT1bNqSoWVn56k
5k4HRBoiu7jaR6L6mIX7cYPoDO6iFgxo9lllLJxAlA//Pc8YmqgNxSakl6mrxAYZcSQQo1XT0j/T
kR2Ef7Waa4GPZVmRFRA3R9hKdZ9hXLftKepOUv1biuOc0BrVFKjNuJHHW4H1AEAg5vzrTTi+T5AC
Ub64ncKedDYNS6MRC5JJuFmdPIJyph4iZnlsUfPvjPEhBj06JrCLvGjLky/+VKw6FKkKTXqYQb58
KHQKlY4v4k8Sg/5NCIAoqyZC+rMAuF/UKavbT0H7wkF5fkSgH4OcXQlEi4IG5UR0tmapLgxXAMaV
SNJjOm3qhcGD5LvYFMXW3xKE0dcHGNdMCeWs1A+WlmRaIlIOOisSM15anRSXKTOD4uga/BqAEmy1
GaJUO2TTZ4r3CFSnw3M/ZEXB4vWfswb5zAlVZm+Hjq53lirmIHJVDviiW1IctneiHSEOtJxIRFiq
VbKinmaM4W1M0o0QZF5OHvmjanvmhn5AF55lmTSrPNT2kNRIuQgwZJDsyVvzuYPfqiwWPHIr9SdN
vK7ift69q+tBanaE9MmZVVqlk4hEh6EVp4hqyooDlT1ZPOlJVTC3fXKtBpv2R5hMJdoJ2lt4MpET
9VhWXOxevzCXTNgWxbykutt0TeGjzrgacgkGoy3+fWHjazKI9X78xLYB4/UD07UKtlV+W7Sto9+J
I3tJnX0wMKz+AaKl6qpIb71it8kxJzxAKASfWRNbg8+ron+Ha0i5qdMFT7tz8s9Kd45scQc8rMDk
j3PlMw2BNCTaR9tSDgVDJKaVMREY+nwR8hg75/aV73AtP+tV3mci+JYJbIZ/1/73xOD3XHuoyvJb
YfU0T4VjMmyGsu5bITxh7gGB+hgNpZIsstIZ7XiR2Y0aQANAMiQua5+CX7r/Bt/DSXxxYwJx3Wg7
o0hOpXHvOZ2ZauvuclOszJMDFSPX1Umr47BsZK0XtKBU/sZQXN7gxs5wMs6E9+gKVbEPF0EsHACM
R+dGkiuLPs3y0BsgODYIaMQE5iloMHzgzaEgv/VCG3tS9DO532zKXy0+lX0WQUaE/bChSEZ/Y8rE
WACrCktr0jORmUMgAW/BfrGN4LZTexKfkYQW+ctNGavkicrbzjHBVgpDaGcUSHU6S/3qlIbX6Q9P
Eqfi47FOWLzzjxAnYKVH0yZpbCmEtungaV8HKxCG+O8RMrRin9ZICPT6U4nMFFHa1iGop+dQtHHR
bHls7rAxcgU4vGhb/Q+8KDXAGrZm2rJZwyxqkcLRwo3IzIRkYUwELc8ulMg546EtzvxQdlQKBKxQ
jp6mJcpe0391UHACgk/DRqsnwb4OPfGJF16djt3PooahYRwpRqp2202pe9nQpczP+FhAhcIsinYA
8PieiV4B9xzIoOU+wx1OMruLFuWcoq9h3/eIlBloX9fY4C+JnoJQahqF2pQWG8S5xLdkQjSrMNJK
u5E14fwnoza7oA8SzXji532UtMPk09AmbfQ6pvCELuGNXgXhlFWc+j8Tz+DfAK09CU+L1cQLNzWi
IelXNAyjCBxf0BOzo9EwyQWfToi0dWj8zPlU5Kmg8xavNimSEg4l7+d+Pq8V82yJfIikV688hzCt
ceZbsBj784S6wMNBDuGoxFYoslhY8BqFWr5/5hAlIG9ESNeN4vda6AlcpwfuTeay/HtFoi2wqyWv
trmTASYErCsuitIxj7JSLRuBrq5em5oxricmbA6gXb6pd797p+IjmEPo92THIq6UmMXfMBHiw6Ix
WlqJ/ZqNqIrfuGLBtz8aQ1FSs6LPJf1bTT8rpkSL+542LJ3+0HqpML2CvsWaeawTyGTIIQFfQURL
0rOVSoC98rAPWYTNBflnkmKuXXITfz3ReG4k4EvxnidmLpUEIr0DIQ39R6yiduIL0iDY9g96uy3h
g2Yb+a0e3f41aLZsCqH+0y7XoyptfkWWG9buXBwd5NCvupFag3dnD6LYL2JiKju0D2SqJYewJFx+
Khmu2gzI1jCnSRbZm+el1rWf83mxc8OtOAilRktQ1nZuAkA7vHQV8CkpW+U0RcG8rNVdLBLX0dK7
bOti49SiNxHL5gSrQemWHqtOv0UEOqOutv4oeJWSJhehaJ4vshtaYIkU6ycgWmoHExZCM9rZzNn5
9JgEBKtQQfqA2CLpCUUYh5knhDmsh179uzFwbtLHvzrU4LmwZ28ukCdHoNVJbiOxniSD7e+2UccS
a7W/t06kMEnIQWZuYqUQxckVRq4+uBdxiS3cQthHRtsnkFDrnaPlQPF5gziwPQi2ynr3My9MsLE1
A4b9zotVvqguL35j3GU8Sdmo5p4ddL2J2OntTJ7H2v2zVg0iC8q46PVVQeOT+HhGqXaBErfmtVus
JX7VqeQAJL5/lmCDxuACb/TiarUKNsv9buunPE2u0vBqwNzs4h9j4mbi4HPLr+r+sTu62TX3KWL3
MteAPwWz9Va/HdiURtJtMki4sV5exV4G2YZG5nQAuYl8DcXOu9kMPegHt0mFB9dlWS2VWb+e+c1B
cghiHjtg6rq3hX2BWiDARYrZjISRxqGj8SMYjzo+L/rKB5FxKanvkPa6M9ChugQ9OcnLkPV9Vx/i
VHlzQYkMGL7fe/YwFj74akAKV3b98OhxJM/ftnwQriDJYneuXDc9v4PZjeba0TlpTJSMkoS9lIc0
gAO5t2Xyq2kZPcgjMiwMrydReNtqPyhfXahUvalU1R/U+KOIq913gYNrNvlPQMtIGdxcbNK6UaWl
KkD2aMCl7VinTBAfOPbbYE82qkYu6ALXIU6XFLlPcRlYqcF3S74ozZQVP2+pRfyTEHhukyPoXswn
JD61Xle0CyCxMS7Ez4w9pCcVUOXsHvT76j1m0g/1JRNEmvnl6aoRl7jd8fVoRw1pez7FxIt02jT3
9zVtp5ikQDwNUa+RjRgRKGg7FJ00c414KPPQHrovMi9e1XIAQ24K7hzIb8HLmrBXHezgLmOv4ahX
vrVzY+EGREBTnK6iooU1xyIdt6ALHHoN0u3evta6eFFGR0660Og7rW/bzN5b0fZxf1tjiOf8P+4M
rJqvChiufyCHI2NrnuIMcm0ysL0wO/ZoJaIfhaadfO4EkgYcAyG6WoXgxnMH6li9jsyppdii6XAQ
DYIVZYiaumtIqTucleyd1h1Tw4o45hNcT9wnzjWhpTs59twWJcmxFT/9rGH29brwRTxcORFnXVdd
yPpzEOMZRb2uw+PL1DJngNXcd3HvAN+nL4Nw2YcA//c1bpja5Kb1zmGxwVezt72Db4Ot6BN4GcyV
FURRpsFqZQCnTI9G5MmHAMgc8xMImg4u/R+d9yJzEUtE4hp6o66F3aJoC1zvW0v/T5Av1jGgSFCj
FtnWfVmp2yrsdIAwDXHVnISWEB210jcVCBsW/3E6jX5H9cP4cVeaKiQro4xEg3IsNvD1D29iOzBG
zjX0QxKpzGJxN7+t97tvTPupuKSTVyJ9fCwtcngayVpmc2eC6nd3L0Vc5NtWU4Rx43eulCDmyM6o
jW0FMFsUjU45/44zY+QcMoHcFtMgVDgZyV4doi44Uh4dh3Cgq1uhE9k43xKx2dUk3PopljZGsjSg
hUkeuZsFv3Kgo6f0SRnf94Pkfs+D0KRNexwT1o+LZWc48Z1aMGtcpwbv1DlzlIA1wycvGKEvOUqG
RHuS2rTZrzp8uOAeLnQsyxqvyZMGGcP3vzxaGmLyySJCnKaAPQYejHHXoN5Ig/oXDwjbsuBZFhGK
tYOLgXDGJ1iS8X30QT+iYVJm2EvAJNIRqnAso4iZFfWzarXNBcWrBYBB+fowel3h4XWcWIcjzyo/
rhfzKxU37XlrnwItPl97ga4ds92Vb6oN8+NSEJpsUqyXCwIa7f0OZY3f4Dogf1IFdJZ7/nmDYz0Z
6n3q5bSpSUFGIBla7LIRqviIT7rBSutSHfJfc/bo768brl9JiFbkRJXrL+NpNo5OOlM4NiJGOpMD
83gBPW085rVcqTQYphbCeOssYQAikZv5s2qMeJRlqlI1JPTxpZlxrGwiLLKActmN1dKH5ybSsAQ6
ffFIhab5S56JE53rpwtNBTETQYG4vM0/vDKka2KAQlR9A2pBcZZtPfuSyjQICw3Pr1diZvos2h4s
2F2tY6VSU9a9yxUXRcd1P5TTJevAFxl5idfO3sr/I6pZHT3oiB+c77DFeRIOgmaegqASFvIiI865
g+GvxUHOXz4jVR0o8D8S9B8Tig+kaOh0KdJEn+c0N/xSOtXx8CZhiLOKxH3HXcFZt/6YQaL4H1IG
7HLW94wd8O+X+q8NCpRVR21dX1++TOKZTVIP/zTDnL2IWCAnH9flf+UxHZv7X7SW8j4MFISfAMlw
zIN2vVb1J+7mov2eCUX4VNgS79ZSmkw87e/31v8Tiqz0HEHYmT9ep/7uWAXXYJzRGjv2GEQvvICy
KIsqQPTut2Tbd0yTY2hjm1SdH0RCo4J2nGnWZFLY+KHDyFIxVwFzIniokwXVr5yjySyhdHO5sKTq
FVjj5lm8lJHqmdTSt1rL2KaRw2kEZhcfCegY3ULzrl2LaMEUERhDKzDn2gExnFUQctFdctXFKZgA
XNPbSIWz1CkbipRMWQk0zDUsNYCBQrLB/vweqvTUzrB7dBZVaGaxOPb1x+NNXyKDlLGPcov9rWpP
j5jyLRKIRJ3uphB3/BltLPS3LNXNhFGpM+y14jyfLX0YJfC7OI9nBl1C+ENcddJ1luGH1WlLQwKY
SFRctlaOZ2GrAlQia3gUyInQhc5m8cnWpiehJ6SUnYWHHe9EQanwA1ACM1JCIF93uD/u/a/DEJ6c
KAufjRJMSxAf/JJHb2VDIP6lgo4FcbYEp/McFkCDQlhpszj82X31Yq/Ox59Rw9nKsTB3WwBXYwl7
Q3dl35U31OO5PzAHnAbP2qLvRcWMZUIEjyDty+zjNyqdyFwZ3NxVnaDLdL76CYAueUbK2zJbC+qD
1GDS0vUzSkyFSqRVbShEh12ArdeTGhs6WvFVMs/oKx3jXoUNSR7PV+9cHbfdjS90fYBsHH1ixoOa
Kl+G4aEavmcKsPNfPjT1jWs8Vy1hiBEWBJ+ngy0EEXY4i8DgkVPxopu+E46FeNyAX1+sSrsXcrqN
F8gdUXeUrD13UMLPY9hIwNmL1U3FQc5cIvZDUZUwgJvAl5L1QNuoo4LLZMZYDvvC1Rkuu/HhXpDI
Nps1nLu6Wdmm6p1hyrX2FWIR4XfnF2x5PrEHAD60VbqFRAib8cqlsmuewHEbVVKZkiucRQCi7dQj
A48Z14ONkP0a39yaujsx+GXkoMPnbv6OFpZQq4g6xllUCJNtSRUL+pX87nC6yObitKSF7zK/3oYw
I1x9v1cvjHM/bVatDtU0jq1vdq120hvvoqtxDN8I42N0U2hUpeZvGwwrTyQ3sAD6GdL49y7pHHTD
oGpKlczMkNpb4CtiRVtXioeYplp7AYs+QLmWLrTt5rwjG2Ki8DFc/QZUofvSx+Q6gmHylgHyTaK6
b4zCQ2LjLysTVRdYAke6a+K05mlNhXfAdMBW/jjJfxTM3WL7rr5elRTPO57r8FjeJTIh/+0r69Ag
SNgHhFoobZzH932HlLb9QAkoPePs0BOZuNmDAQfInH3QHoJHHlFw90huWnvJ/VdoV+jzdJq69UkR
G/Lf00AKyml3CZZS6oISxfF9ufTDHxO3u+JeQumh5QMmFWDe0MSswlJKLE0aNwSMmzGfg4AcdYa+
NJdBCxtixbot1b7n/1bZ3jfhcEYWv8DnOoMeltbquW5GeaId0Kk4qwXB7QHWsxtl62yTptza7V5t
48ifqsx0CMVexg0qq3c5Xvv/qzBLcGeq/xSl1MLCTEjLmzTxESPrVlc9Qx8bju9ib5utp28Ax9cc
c4AsF/Ti0dZ9fhWtZg72laDeDoYxwQ0s9XA3V63FfXkCCZgiGwMhaKShxZT9jAJ5aH7M2MJajfS9
OE6I1CBBbwL7gkQvYy7cZME2+hbd++tcj1cHJmlR63UlSlr45ld74YSoVbQ9OseYukR8foakNQEx
d5He3agMOiuKzatOX3+4JyXYwpkGqoI0mIKFrqk+Ew36YALYbs3cNXQv1XjJjwpICPkF84V6Dfmv
0bfG46Y/cuQUnaTUhBNGrUiUyriHwCXTRGx9F7ioPa3craZTQ2XrxJD5AzR7sPrc+i8CXHzL6BSa
8IFho/GmrBGjgalOttPPxxBpByMTNN5QzQH1KvWJq8tmmvZQrnNGRXiqfrjEqOwVj1QBLUH8bulE
7r3j+t5DsNMMuXl5Z9MmWLGj4ZPTgx8PWimyZ5gHqT72eJYcFy3JnhvbFBu0UDigGO5yO4l21FbV
iJuBoILQ3hiqXiX4GfgrnCWl7Wi4NBc29Pz8WXJv8+RaEEEspMMGHfn+IZZKmaQh2Pm4XmK2mtjT
ADC/J/q3G9YghpBU66/iP7OxwHagTuhrdTQAQAm5uwwQ9hk2s59TcUo8Yy1EmjajR7fTrv0yfzpl
fQSOYXoSfbKYpv6D46f9JyY+hE88Cbw3UBEcKwphHv47bg/8PwGJFTrR2Bjc0mEDD5WK/WGzO26U
bwESfPNt2n6nk9uZN2egEXVAtuxs/9KS/VEEgjoGi6elM6XP6m2jk/EMCA9KroEaeTZ35V7Wpbbv
QPtk03wEQ6A6rUIsAQ+t4L+f2WJ1hgcUtut5xddftnhgVb6Ap0CyVQAvNQi5vww6Du3I49bWcLoM
8dATE0lFEfLjy6Kdijf7wcgA+NgbgzEVy1rBli5S3gZMfEa6QObkFuZkTIWgbbSaa8Ar6N4oY+75
UnJ7G4BaV7YTJNCogW57hEgKKvHwflz6X8ll7DxR5DokLWEevXJeygGOsDxNU+ZGe8N6OcTvpZNx
aBpuRbZP6vOZ1m/LRwdf/C1rpIFet1aS+yNUPHHSFX+vdVKevWZPsg/4/tQGFgkwiJS/Cm3+NFE6
fFGPNmDBvJ/nDqm3/B9o+sK5XDvZ7HdEXOSwLm1bxnVYTjh5q0ObMkeiyNjmcODVgvpYtyZx9Co5
PgQnzwcJoAEvqvi8OrwRiAuwfAYledkSZCrUaLGdmuCGLMn6iZ8EQPamzn22kEZTNg9s3vML1sH4
sYsuAV4j1dP0s1ocjxWeMb/oeJZKoBvt4zcqR+VuKhmFHWH5D+RpZK8b1vSxfs3+QJTEpvEs1wSM
MHkHgauwUBWknGdFewhH3cEggIm9pZS96HzqR2+8zIDpbFo3gtUR5snVhuqoQO7RvLyuz7KEp/NM
wM/xZ+64jE0InspIG1Zppr01xOzm4iD0+bZWQVO88ZmFcxa/Z06CamG037eEWg6bVDC31voZ3diY
qRdZBVvh6X2uR9TJT6ok1JF+WKjyyn7Pzj2u1fmwdWJxo+poo2hRZbYyDUbTFypYonjv7YfzjoSI
1c564xqEJtjzsXpSZ74S9swd08wdDupyqYn6HtKaYJZczwq1G9Kz3TrCeGORdRFB6f2X/BxzCOQd
3WQ8/Rfg5VlAWl/nSUCBCTJdXgpQanGn4T+c4PmhRBz61VjnaL9HgDQzFVDkuChpAZFVQXNnYj48
q7V+5vtMY58UJCY7rfys5kROYFmySKnKmpCdDfiaXBeS5xa9vWWrb8yY8DafnnXxMEeZ2diZkbMW
uSlCW9Lu/hsDy+bRMbovVsGlyRLEgI7O8aQUST2usgAX1udY/W2d2EU0zpfzNZNirXcfpETYi229
nMrH0KOil2cFFHD6MJKgZRr9Htv48FvCji7Cy+19bsl0xlS/wfJlrMQpCoFjzfGhrzDfA6VKaUAe
AGLK/oBaf5R74uGIBq681hXdmD4karTO5OIRf5la7KdQzANuzH6DScf8FV7JDDRJ0zdXV7TetjWV
WSvK2HgsUSwO1n3W7YjQ4/yuQo64cLcbn+QXcfIZ6OddjT2vhs9V0jhxBw5P53S3A5pT0YhpMZVf
ubhr8nHp42bcqGb2BqyvtA0W9WBF0/FmUCkWhwA4KzwRVHLSL6sNH/bUyPzrrz7nxiaypbCH9aWO
MzzLfJFD0J37ExAbKD4qrJLFAhn5MN9GNro2s7bOZtuUTA54zh2XvPH9DKVbbeYp7IPFIuRtRkLY
u3f6QHujrdXswvwZxwA0hhdaPW4dqVc0B/Ez40EVkbTbY1veCXG/6CMqWzF86n/J5Yy2GtPELqg8
NvYT/rBNvkb8YXOyQsXWjcddeWiH4hEILYRnixySNluHiBrjJ2oOvpd8IMrgLMUeB7LoO1x6peIM
cuLhkrkge9qxqu2zIY0AR38d6jLhIXo2joEe3ElbtoTJ1wtq9wmOYmFYGt/cw3n8TLJZvLtVqzOn
JYNLxknrqmIDPTvemh5mqU694LHh6/5b/G1Gcm7x8gDdQql1fB9Oi46o8mFF/bT/p+dV3Aoh9DvJ
oX/V0ZDgnZF2Je7dP5FuO5Av+Y5BQWtz3n2KyeHGIzeOS1CbEHSVHyxYHy/nB1IKjnzQNOUrz8MX
NI3eFLPzlRAiFDlM7Fzk6Ls/GY2AViYtpKsi1JChoq64w7ZOUINU8Sf7nmOFHDmU/bh67b3Y1Wvr
3q7jiQcJV6X/to/w0QW9fOx/YTXbS7WRTOxCm1tqWJJ7wJvQGx4XyBrYRJD3E2wsGaTuQO3vJSJd
k98fQyf8uhYFJhFVLbXGDlDrYI01yaygybzMStzAv34N7SrdRWYrNruoVbQ+qW7xkQ92yZi8XzQs
ACqIPfgwlwaFenuBiitbY83tPAixVt/l4WeDpqUgjqcNY9XuB1OIth+Og74Mi80VYfJbmxwlaTQx
hS1v74H/99oFkqhw4ySSEm4gFiAZ7Xs5T/Uam84XLS3+bZNdkh573JqkXFloW3hSehg4j3nj6vsL
nBWzsWJrdG5kADsMniRWcuPLVlXKLLQtinitIyeI7twZ8O64PxEqV5Y7OXfDVmUt5oioK+MORwzY
aJoioRT/mRsOxr7NsdGLz1MSX+NsVisczemH6zVhleUAZlEf01ulrH0aShSar0re/GIJtRVVfEG4
Zhks2oncQnQtn463vu8Ivn7zdks+2QX7AloAY1L0i5BTl+mycWXAoxfDxWOdQRZZSJ2IHKeaE3Cm
zJmCDQISoOcMnIMSknzlg/LomFKED0Dr2RLpBIvRj5QMDzKnukXpRxuJo2IoT+2pFEIgvFXhlFFb
6UgZz6NTRqQJ57qKpdhYCd/SBB5ZvLbDBIiHPFI1g7Ypth0kDb9E/W2EFAtZV1SnKVG+Z36Y1pbP
sSg95+b+IjF1LdW4lymuIjFYmJrJaMW2AsLoyz8jvaoNwyedAC5x6rPVtN5bBChiBSPTmeEZxmnn
61kvkGFPF2OoqcthZmFxVfkEKoncYVglfveh2EMBtslDb+MKe8m/ysf3RqTizpICV6RgxhvXxUWW
VQZAueGpLXCDm8kchQLtMudQGuOYJmN6qnGgyU5l7MxtMe9tUplMjkD5VfDc2sTXKeSpgkLD7XWH
ojisw7lbLnJ5BpvGwNCUJ/j2liWVomxG7IN9aNEEIReijl9V8n65Rt5UCtIM6cwznRBaydLzqUwK
+D5KXnJPGLbt9PANNRGU+7uWcP5XN4ueXBlQjIH3lyGxLlodwn3b/XRZD9lqvQZACqgrgMTZyF4/
4jEXH/29VuJxy0AyNYHGdCLe+FHQu5fJmNAz3tSTQMrN3DFujFaRnEqy417NA2xShhyMBwRzdlIc
eWNWbq9i++LX9h+ESvj4pb++RJG7l+ExiJI1rlVQpgfYGfrDue0RxOHi2l2ruUghYe9dW1L9cd7y
F1n7JnrFicTWNzm9+TD7aG6qhToV5XEojlq8W6lw12MA6Fh4fbZjqsVTl19f2ZySOp1mXzVUTSux
Sm950N+24mVWGhwpY4VKq1eefz2eU1ayCgmr/RQMbMwGMi5cSx2Soafr9raCrCf+31jOtqySQMUD
O2y8JGcMRW+t84M6mzZ8ALoic+9H3UJN5W4LU0fq2EAfcVuAz51LIcbPhZsKh52YC7B1578CN4h6
Hja8wQHN9udMmaDV9/zW97qDd2Rj1UAo7ITJDPga9gxpX3UUT0HCeULHZZO/9bWFsbN1v3aowwKp
lmegf3KtSz2lMf9BEwAYf7SktXG2N5np08nR7JA1+8vDWDVrOgQ6I5DwJJT1wOYCJE+q1z2oDDex
rFzQALiogRssNtRENkx3kiVC+aPo+6twx9feCZZXHcbUvvOXSVPMNjD2bHYSSPApSc+uRfoipcLa
uBWNroQ1DKMpxvU+VnOQXnIRgvPiAbYI+xB7R1wNRkUqSVrYbelp8fDUlLxjJ2AgA1biRw9aEEdC
Iap/oRhgF1+RPWFvQyuwIVRlH3AsAAqVf2eEpyaljWRx0jc1FmSJW27X/HaHnO8iHdmczXBHhSRY
tINtkqzub3QCorNKsackNR1qiB+27bJUFOEd2Ouw33RJmgUK3DiiVGEJEqKoK6p8YmryNfe0Peo+
lmSzhxeVv1PROhC3YHGAfYY2MMvkYStxVAitOq4ZgnfnQ32MDxFt6ODjAew7sRr3mbTqVyUQ9q2E
783ALZg6z3ZXkAQQkIWlCY0nTkjnyarNvWk4M7gkk5GEJNMXp7mlt5ZZx8O/oEvwalBsc0PZkXpH
F0/yB4y1DH60LDfw7zey5faC5XspjVHBnewzOTu4EHnuisWJ+g8q/l/LfXZj4j6NUiJWD0t9kYBv
vyaNQfSyHFiZyomtuDwHaF5xIm6cxG3Aul/NtQkabhIb65HyAPNcclCUn+V9cCwD3QkgpkPechY6
sAAqajLYWjomWBRqUdbx8OdeGUXTFWRqPQz+5uNMxKnYPUbP48x4iZ+dFAOb8cANUCRvIhexc42K
WWdDSHhNvpxPiB8BHWfYRmSfSHmFBFWzHNhNQ5f4l6iVq+L5BjqG+TNVRTELMGYk5X6WvjhQHY9o
IW9CcYLrLXzGDSBf/b0VFwcnxhgXvvkR0mxpHerkHVJBrG49KpEvufNvt4j3F7pTFZdWi6bCKohx
K8Prdn1DosAhGu1bkYIN17uwf9prrXV1IKOe1Vv55/DQnurUP6CrinAlO8uy9zRmmokMppiTbHFJ
MTFw9bd7VkozpMZHsyTK1pwmMz4OWyfxuaqJusuW6mEQ6MiHJMMq6aIOHva6IE8R7e+rRwuPFdFQ
9EV06Q/nTPIVqAQVElRxtH1anvoOEwAkRruvrM+RX7hWycTdoWWXa+/FfLsxSVe642++9sd+A5ig
iTXNGdKGEaOIBJHNDqFyrJft6neFaOozEnqxkVClJIqaA/fl3CdYa5GeyZyF14cYUr/gcIFEupUn
fvUJsgWIXvJtWe2Qh+QiWrdbTYnYcK198OvnnOPQ54UUwbTvffYbuFM8YTPcPIBWSPNHK6XiJvbX
lDtfxTLREYqtuOu9KPQSn/W+UnJawv9LCdE9X9TVA5EvBlQM77XPw5yELFCNUZFI3MVYrJzwU+Mg
2Ut2ObCDROxGJisk8y64i5FEYb4OvcH8b06MNz1kczvrV/8B6NLbp2MVzuJMS8v3lJipt/DEFubu
HggKvNHQ3lu1dvS2sqlS94bkSxGbCxR/N9OeewtqQ+dKT3/xzU/1YWhdWtjuEpQSVh90aEB+ECRa
MzbyEfaAZXN13FRU8/dsLA3sojQr7DMJySgTdYb3mKyZVm2UAZawfZSBpiC+gEgHebCbdRB4uaRM
gbNdYlr9G+e7oJ7Zg/kIl059qc79pvJhdaqMS70adNQgRCW8HMpNrnNo4zRuKjM5bmD8ILgBLujb
UREgouIlVtUNaJqfKJyTYuQGcUeuGb81i3jlBjUXy2YbsOL6g3dKiDEP1Bg2YwwFlSC1uETuqs5w
14NeXsg+HzCIKqjm9XtdC8XKvM+ELY7IZuOSyTt3Un1WW9bRCb7NAzqYAuUGdR+aKtDNTgakwC5O
zVO3oaMTMxaz9xIETYJXeRdb3MGL+hV6sK/Nar2WBTYg923VH4rEQSyo/fcH3/3xZnHfQLvqR35F
FNtbtOC04NQy64HyAFb1xV3SZ9+p+bEMKT9TpJFqvGj4poCs+Za8ldF4JVNKjjwU1EEM1nP5XUiO
iemM/8iEHXxhV5DjnegfZ84JXsyXRCyFL8qnhHo9PyCODIyS5aoaVTU49kLTakfXRSqTRdslmLSx
wpOQE88qucFZuy5okXBET0CyGEZ19c1oS9dHX5MEffbd+fiKBUT/mYAUHJR596kn6mxNFOeGZzf6
mTuako2zhZVw1lg3DYV8eIz9m8ViuTjAyGEiKjjn1+9iZnAEbmMY0khZeZw5KUzjYggaE6RQSw6a
iEXRe8+I7AkOVcuQ1PdHdX/ewMKK+Nv4h2ZT4HYvBDtLTbVJXOL+HvyCeSb/+Pa/zWy46XM4GZai
zKveaJVGX88RUvu45t9EpGoj0byrXy7inNUFN8h6WW5ChlKXSG2HIJHrqBkWImJZsfLBuPSNyNZM
rL5PhnCxhGsdo8weSg65JDBbhG1dMrmfPxUA1g91nOMuPJcQZ6N/Gw8YuaaTOzJ6Me5g1ovKHl4J
bBvMegR5ZFlIaWju52K/A6OohCfyr7XbSGNTvM7JU+x3vJHZ5D+lil1wXeYIRs/tXJ/nkmky4Ahm
jCxZL77PVfBArtN8L1Z/9A9H5qBTMJ1vHaMfeY3SaDq5NrgbMdxUT2cgAE8wMtz3vhfFAa4JXL+a
PY03HNyyo7C5y9xikbbRDes0PizdP+TSGDxcsKMGja5bjz8LYJBk+y/brWfImFdZj7H8WySzfvoK
fJKB3g/Qhz+fg4AYcYzBtGpMP4cCWw4tyRw/9u8hH8Xsix6l17+L4Noo9NpsRZQywLxeRM0PeYDq
lDCXoslChwbKPnZVQ/UGyqriZlZrncsc8OK5ad/zwh9Bp1FGmPZkHEyYJjp0A2NX4XE7vkKPr7Bc
GpQfmzt7WOIfjMq+KNxmpbjiUKWx3+tD/Igg2zttIQYRXAEKhtcTPbNnMtPL0IBbmFJ1pk5Df1vo
N9VxZdg9dh7cukC+yKkD3Y130OvfwseR30ay5jyG64wNOjri/AKG2cUlSvB74Um6TNiqnivefNhE
J//LEKEWu9RQvyU5HM4WzGdp2fOi72VluFlUC8uZ4eKUtYxf9OzT5laVM5d61G/q0VsobLqE2UWn
X2Mo8OBUsO/sN9ary8XQbAtSk938nnjUjJD//cK3evaSdVFzRGwCjhCfg+jnd+8QkwoaNKAS/InD
eUAaYCOj1hrftF9yffl/gVBgKu8S05/5qiD9zIoHZUaZtO65vJPJ8WKeCnQB06L/qBuG7GCHRrLC
FvBhFqW5fbN9m+5ahejIZyPG1PGLSX+fBbaUfMY6w47j1879gg+OaU0qKxuysVNfct6K16TaKiXd
LZttvrMWZdUv7ubQqEkVJ4Kv93mOcYZFzB2U04ayjyIpHNezGDphBbwxo8xKK0XHMLhKU8Mp+HUQ
PpT2sQn6i9IMgrSIX3oVPzvK1FQRX1Fldo01nTt2C7sBY/avbtxfErWMMzxybE9enwzFrX4P/MOt
ptR8GdysBC6uZhgG1whnk6i5B7evCbQQKvRcjDKJ6m8I40zr8LMe3UOwCKCQF6LYEwQHLq7c5/7A
wnj0Y5lVxpu46jD52FCM2lmdkBSIHrJJJDWE8qI2/MjMcBmBW7twi6p4iuoLjnLLSdIxOjK9Y9Fv
akPV2RaEz6Ymj6lM8kQutZtV3+aRxC2Bsf6/IYCzdPm2IojmaN8t9UVH5qa4WJibhKymZMQgNSVF
tr+nfhC6OKJ3x2crmnxWifJrpExa7iJkex0szwghX2maZ/8SDn5qxLco4TcdqRXfQ6rnhxvwEzKK
2JbTX27Yit59iPzelIFZ2wrpHNAKftw1VvwnRR16C6gTIbAOszmi26RBj3MSfFL72bxv7IA316UO
2ILP3a224Cqd5l/We6UtMIZ3DU7HFY6H7/q2BV8RqFxhNVA+Mq9aBTqSL89gKBtrA3S3eO0sH6/j
XkjLeSM/ScwGzsSHJkoMuV0kks0Y3hbxrDci/lkuI4cCR3iWfPax+7nMoSsRsQ4eFNwE1mmv+uUP
lnhMJj0AbWPi2ArNySN2i3AP/Wy89zNUds6Tsun19bgm9ibBj8C+MOL/vST1hCAl6+7d41qtlIu2
eJqvnjei3ms4jUl2YJzJGv+1zh17Yl/72jZglpU2XjxHGG0g7QccwIIdxDRfFXlAYEWrYADCu6p0
EmTK51TcgDNxa+Qa9tvaY4wGQRkCx9huDWWgzQOM1wOi3aziJ3hrngSP1irj5zoiku1EM7hc6zlQ
6sspUoNtb6oMunmDYAh/tjyerL/MGSNvtOTNs7rs3R8H5QpqVv126JNmSjoNf+4Pu91MulU884qf
OQ1mJ2vO9rhqvOxJD9T5Pu+YJYJdC9Bz5bdznzOdXHdgfGVI2lURR+qWl6CONnffBala0e03MsQ+
55ZOvSmblZhPKDiB+1rHH51gg6OACTvfjjUitYxiNv7+YL9fhwvDNTr1+0nJAQzyaQaih+S1XRtb
IK1OoqrXUAiqsdjqcxCvGAzjrOAWrh6ouqbec23Y+RO4mej9Xh+uP57lNk8VfLGjaefxiWNxc9AE
pO3a3K6/hke72ZSD1Pqo5dK8bcFy4Dhjd4+Zksr6mD82wLY6N7xPtMfGxpfFffloueavNz0k1faj
jCfNqJXEre79ESCUJ7YXOJsFQ0AFsF98fL6fPAqWrI4s2zH1XdO9w4XeYfwp3biTp0GxVmuO5eYY
ZJEv2IxIn95lp6obizRsHeL8Gpual7AF0scfe1DPbesFTyrZBLn7oKppS45Ejc+HTTiv+oKro23Z
m0/8F1GVQpohZb60nJqHzx+iNwS1uxgv7hpld4w+Wo0ibWa5PZBU5jHmkSocLTvNKqCzt+cpyH3t
BcREGnlZoyDJi5l0/Yc3EZ2uaPWzJx6t/SKfqfxd27nJAl1eadB5nE5BBO+RljsxOXmsU1vr3sHD
O+QguVJic5VFp27aUqB3z0Vs4MZBh93CgXMSVY7lkKik5VCM8Y+p4limPUI5bRZ5kkIvLYc9F8i6
GRvHdJBrTPawc7AzdYQQMLtfLWvpXEwyKeYmIJcNRxmxYWYeYpWcQO55AP9bOqLS4Bp3hH8f75Rw
btuuPfSlfEwJTgRzGhTlFnbMxQewGpF4URSCXdeXN+dq3rCja2hru3h/BONUd/Zh/4WqHYnWpfAA
1+zO05ib1HHG/yKb0rD24a7WoE8bWLGPUYKwwbsfjxUJMP2KKD1Gthp9ZQBYa3Q6Z4m4IVUUKJ3B
3rOKBuuCUrrFbHRctDNYx0JViQcN2z07Zn7bNNhzmmSlkMbscnHJogom05uwY/1mtLBZQsC0aN4z
WUay5x3iSkDZeE6PP+5WyUJ8WiKBJ/P5/iOhXWxZnWeyFXDdIZDG+45W3EofC5RVVTvuRrLhSiVq
IhYnJJgGBsU2pCHMs4ZfRCDVEju/0z7ML/iuO1sBWD+9S09ePcd5/IqGvs57/AZKpJzA1p1CFyiZ
8o8K0O+uNkQFNSPNlS50x4mgzU0qodDUODLNN5zjiehond/nWT/GqpDcV0S+RajHkDyysZB8lxia
wCcMJALX0s2DbfkgPogjIxWFGeoeJYnlUpPEaVUKS9t1rPK6HpYMtDwDeNObGlg2KGuBEkOduaV2
Fw9ZY3ZPUxE/hDkCYNs+61A804vQcDqfSdzWvbGEqbO/rKB1QEhqYMdlYZr0Gl+O1Nd1DLBFRgmM
rpHlLpy2iQhmIFJP6b4uiXKeOIvHY6LMFJIxrFlH4rOxXV3dTw/zfZjWp540K8PEi0K0CGoENcRx
7WObSgGz8e1ktnvdrfI8uFZ7xhA/dH5XdwzIhDtTugpPreoeynwWZChFFpjsZyksQCfyoT3IVUPo
xZD3DWqmbbNB3snMi8Ep3pABK58GnvjcotIvlNyjzxTVH+R4dxQsJPdwqykUx3/2IW1UQFsqHSvZ
ea3MzrCXJHg9AfVeEdoe5NfOlTbVUxLPaCae3ro7Xr3srr/ybZyiYsvdo1QGspLux+PQkK6h5vYZ
dj8+WvQoHeuJWh0NoNvqkjOooOBHudwrvZ1EVasvLHB4Ikzp0A/nS29Ov8WEPSJsYZn2ABHSqGXv
6XAQFTuJPnXLIIYSWdIBhzHZyXSRjXygRWmRNJjMfUS0we7uaIjYFWZcbquhoSpjqJyb5lT8uXUT
q2xdAzTMrzoXmTKnSpCvEBLXZxW85riK+qp/VNYvNnUG8AJZynaoPCm2tHNxHABAmn7BanfH7AVJ
A22UbVtfkTlFfsADJCFi8f6qf8B7b+UJrVJXcQoP4mhpDzMELl09gWN62hS/P2f9zef5iS6UFhk3
Mpjlc1yqHYRLmYjbfoQos2d+Wk1y7p0TXZV32ld7ecU0tcMfsoSuLEmG0sZTycHGOt2ZVw/vsnM6
ZPKEgdTPHGYJD/8Kk2mKDsbdbJ9ij/YZr3bQla/Sn8MA9RC52B3aSPY5VBNFaGc+14+dkL41EPQn
/aGwz4DcTSgoPrG7v630pfDNBJ24RzS02onNhrlT4ubg6mDYKqZyjyPXhZWQBwj+ov1/A45YRhZ9
MThgeDyH85z7HBXzZqjCP1YFJ4/A1BPL0GBQu7qlnPNcSrvmCsNpndJgYTynrD9bQnlgmAdyPtls
jTb50ZwAMD3hmRO2FFVDWOSVDdQ+8uTCjsMArfohcxlraXHCW/MEUdyjUELHAwCJuRHXd3R2rIou
4MFQMY5M/Z6XuCblE4tjWurVdCjGJ/fkg5aAxGOiqEAbduuq0YV3vIpD9WG/HBFzbPvAdEI9U5s1
r576YmIMdMC3IADtAPZwjZbNkVQ9cbdaHSxU0U7fQ2C8/KAKxfAmoI4JqenAoVwOpPSea1g7yz31
hSqh0hwndGGjTYMw8JSMUjONAi49Hp+PiLkfFnEB6sK4vHxDtObLnAODh5ah8s0NbEVE6iMGA12G
uFYRhDvX+A+HGJidS7ToLhx/veoozDCwjo0GzyuXaMdx6RdxXOIjQ+wfV+B0HeWBuZ+ef/blptGf
hw/WHkCRRTc0jsoA/zByuOWx0UJtZw9N7vMSL8JvWyr9SccEAQHg23W2P4/X+GOr1QDrfqjWnAaP
7vz15O+csps4mBRcWAb9rW9NcpylxnTleX3u26uar0TC4OY3zvFk76U0b27zHN/LJvAiOfeLi4BW
RBIcuT7Y876xzwMrrPhZHAnQd2SJkus1Cvj8BZvJy7LYJFPShLFsLaj9PMjb7qiFKOgbquvLP6Vf
UabygMD1tlKil8apd8n14NCJpsWBc6Uh85glzslasHorUJ3cWNgKLNAKDVHMcvVWliYnibvK+7ju
Si8ayFn1Ug6ZGcRtlSJ/en2diwRpYCC/FeqTv2kSK+19YF2tZ7BMkpjnCy+b+8UGaFm4aqpeZSrp
iq6GGo7vQb/3TD1iqVXBXedIZLduMQ1qn3/MBn8Vg/K9/DOwk6fKXXob2f7+3xM+LBPMaKn3tuv6
DQPJBZ5pXtUarqwebHoP/JaMzEmTpeIlKQeDkq99obdVy6iRcPjUHUvvswlrhFYJFSfrT63/yA5a
eg+SmImPylVUaiLrQwlvT+iqRiBgdy9jKxJb7OqkPo9jSlGrD4Nm6dku/3qFiwy5dRG7/Uz9Y0mm
S67qYDLG1PaFHGV+5eLXXWY51weIAMW36fjYt5owQafGQo8xoIjWbaB8TL7MwMb0CBALbpSr571o
Mutk1CU02nhPal29H2jNurWYH6hQTCe9bCBrC91hFNOP5LW+8iG2z4e8Ps1tECHVTzMLIsGuFF8u
O4Hg9svo5L8H5uNB6uPqMNbLPZ7oqV1xS9Zw7efjhPFG8nOfN6ArwUuOtFZA9mG0hOwUSjWgRPHJ
cHqtZSvKV0OeOm3ejz4UZlkjhYcXXKzqsi5rvoPqR9WcAX+Ku9cVshcrIu7Wig/6pJMlzOx9/eko
cTGMV3SJp7G5+tU0DbHr+6QQE0cxVx0TPSx/cUC48+bJnr85LkB0/wNjvE/tYGft9ozJkNP8cZy+
OtBb63s5pM+0JVbDUqR+JEjyXuotL9Fiqu/YX/BgO7kUswDRgV2ptpIukpdZdNeD+cbzvd7cwZXn
0iGuY1vimQ7U0FaD1usSOpIdGdg8gGcjIN4IXvNocLy1tXCXHwQduNn+AWtuwi3UsUPXtgcdNJD0
bVVrWFBoLKmlnNYFV2TlBuh8iOdwAl8gzPqKjjmikqv44pj1NHsNt9uP5bvuPr6M4ut6cGznQ7Kk
Uqgoa29f5z/FgPT4uQ/F925hSGkLp/GKdYfxOWrzZ8nooM8coO18HJ3qGX3+7Nobq9XgW95rsHTI
tMuuo5GxsP7uk0jeR+rq3t7CEA/iSd2pqG2SI5yNj0xUkpZU/8gcthUNmQmG4ldyivHxdOtZj229
9PT06fbNtd3insF0GE+1v+TQDoxiCa+MikMIgo/5u280EcXJaXWH3XCm5AAdYhoFllk0P8I0jZD1
pkU5WZpwtLHcHtFa/Er2cYvOX/poHxosc81cManuOajXrCoD/oOZhwdrvLd8m9Te9wrf+LcmafNf
BPRiSMKUEm8WM33DPz6gJxwUgiRjf5Bu7CKMslLPZ0vY/Y3UBx6Nsia2eG+SgZyunawgW00900gs
OLVohhLw05AjvIT8abPyaflXIdcRKnuo1/7MEgAmeGKyFjCVLRj4aG+gJmcPhRpm6kj2gdZ2pskw
tDXFDM4oOO41R0jTve7Q4/utKTJ3vg3ajuTkNIruQgy31B8UckKi0PtHFlAdalGk/XMLPHWSWM1H
uc2krxO9ms0+e3ethp9ayY9wgNnbzRJaDsO7mwXcLOMguHbidZFIKTKJGKdBPftn9RzjZaB1nHjK
QcYa8bcZM8Vn7lBBDpNTmQZcZuw3bUrcf2GNvob2TPWA8g0HitA6A0bNQzbCXp90yoXokVwqjIvO
x0kqYFS7Y+LNIQq3kSoMkkcw+MramiDvdqovWyN3qD7W3WCNbb/XvDmka61qRcSC2H3lwq6fVpDA
HmLYzaJIoR77bAgksFLVt9gZfIjQbS3Zzou2Gb3FCm7z9N/G9S6QbMibmblxM+zzzrKvtWlG04XG
d/98H157bVIpG8cllEagYR+tAhtdNrRzmHMY+s9YUxzQ8yfKJCe3BdaSOSzOYv/wKjJifbvm9Uqn
Vx6AAGzF0/UPNkRiRjKnU78Bm01nU87522moqwXoFWpYJxROx9B/fhRTf6TtbyCqHbVZ2K8OZ0av
YOKbGvJiO1WHNAeB7mXJlxpe5QWoYWejR0JXbZaJt378Q9Cyv9KXJjDe7bNtpzUQkijpTlldzDtN
S035oMYnP441xMmsJgAcj0VPux14fac9m1GWY5sHoQBkAb1F3xw2tGV0zsra+xUIN8/bwGgx/ea7
LvPHXDAy5zwNWm8GRUJNMbKMpG2DgDViSubH45Ns7nPR3oFz6cCRXX8vpo2smQcCNBmz7sQOTDbR
8GCHpwNeIysKiectB95WNbzy04lFLyvMssjV2GmlqrNc2WvH37QFlRx96N8aHjokjdfU5cKQi9g6
I9fC7Mi0XssqAJ1wSAmc36D4Pc9n5pH7gF+qErUgrzdhscttGMfzB7JUM5+F1TGNl1aJvN72i3Uc
8vCBLNPFrtRHP47Mk7tfsJg5fmdMNR8+VlrwDMB562/WRMdix2ADPGi43WfoOkafCcTaxuCslcGU
3dhQ+VarF1EY38B/ax26dNc4j0gNJym+sfEKwPUrePipjUgt2WBVVdZidWE5w51FJkKHRBmu2vC5
IXuoVnhNyUy069IHT5ygqSwXhkp/s8VGVZOQEtMKUFGqKsQnYEASxQDTrJs/bXcPtCtm2MfG0ZIL
dwXeso14KflElwKYOYOuA9aXDJ1Yad6d9n/vSqLjSF9Duv/jK1AcuANjoR9otiNdYeYv346mZUpe
V85/RfFvolBRaI2UKZXPU1AOzIaJaQA4cg5VMT5a1do83hBlWsEiQyHKvRRfaOGH9TuCtmEo0qAH
aB9ZDSO6KAh7X0A9ke7z58K4Sdd/CY+kQD+Y2IGDdd7IoCLCg6RzGpQCTGVe5TrBkj3XQ37QdoMX
ViXzYdY6qZNudxMyRLceowX8CPaOg4jtYk7cJbLQcIW/cFMxFyn4nMm+h+hgubYIGgbQ9uXZgxJI
GFcm1klL/C6Jgkb4p/y7FlBDe5aFZ+kFdiPhKYaPXlEvEc4XdefBceDWm89RwMS8qCV+ZW39qnJQ
Z9DMKq+r468yFeYPsRWIZbFKde+XOXaR8KA7g4upaYPDrX9oUMQikKdXCmveqijxQtDTbEGnxgZs
JKqp/NJGApv+wF8SXSrTENaTKGfSG4SW4ojVII4a1cAQiE1qCHpU4qu6Sj8YIhA0RBwrbVL9CngL
yWqod5QGFiq6l2PCvObFN1KA1j2HE0wKUuux0z31U8jSijJFxvWqPNQhv89xBTtxL/NbypTTMC2g
8NuRItRgLhBLctQJBpb6+byqWIOLXw2cQw7uluJ0bb0Whd1mNcDoQKRRi9uvl9FU5aFWNGce2sqM
uFkIR3xycSm5TQh/ZFekUj0yTtgyprA9vl2KZ63OkZ3bK9QXBo3p3Gm367AKXXD8ZKLN1++sGxIL
UH/aIr98OHlMU/DgG/5KCWiwUEMuJKHYL0KWBNIAVW0hTf8NDCrMs22FmDuXp6RyrYumS/glT9zI
JMeGdlNsMVyFnG4e6Bu9lXVP6DbXlA+dVcsZDsplaZvFtmXiCdKNW1Bk81rx0UvXqLRuLw/dt7Gz
uJz70IQHsJ3POXP7uoGjUdA8wb1cXpJKuknWCBRKStt12IaIgdcjOVVXuy7v+wEh0lJGmcrT0Ror
uDofU+Wra5WnlfHXbxJRvZfqAEF3nYFYxN2VQz60pxQOJ4+uXvQqbu4Ht9loj4zvqkgGgVWyqWMs
d0OLgEZjVu1IcL6jiP6Ay1zB6CdhuHhMPkiyfbUKCCCkNhRbhJAYPWP9NT2m/XI=
`protect end_protected
