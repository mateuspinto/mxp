`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
H5fpvTr3AjVCMZZ+0yR2R5DCjf7BeAIOUQ3V8BG3xkt10Me6/6iJkHHTKnlH/UmX+awTUepalV55
1sPkX/cgxG/9hITwXg/9rvvGh7DbWzAevTj+49vDJSphjZCznZyW4uPGCHn2VEepkSDI4XcNI6wI
13xyZfIiM3FcCEahb9MN3pPaLKaTyWVvSSl7RrDxhY0qwk6VRrRj/ZifBVt8+w6WJjEPwqNMQwdp
HjvBmbUBKkWsHFmhTy7Cf926TxVpFiZiUsWD3s9HwX5ZbhZvxZ+Gp4RUZeavjabVyx43P3ATVbNN
Zqhze3RSXOu8HkhE1sEzNNTuZwYyyZbwmL95GQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="5AZ+8wliMKKrQHGqfJLZUUdNp3917h1h2C/+0x28GaI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13808)
`protect data_block
7V567nPoVcDpQPLwqbyN3mb0EQOZuPKf494n+83f0/Vp60xVejqarXIylSDQjrXZC2XUVOTbW+w+
mc7TPfz7oubvFMbnlsf0OsxeaIKvLzGdKJyBACqYxicUiFrrBlaIewDc//LYd7IBFbVT2e4UFXYY
7J/kLmqCZOU3TsUn5O2d45JcJkKgRJK88SyZFrZOe6ExLpqIFKG1srgdn5SdO/cdnPAdyxrGl0ls
y275f2gTHCT19NJ38ewuCl24vLEH5z7hPsemkib/GQPe7DwMR3TU3rMelcX5ZpRnyHxfTZgC6w2J
EtoG7iI2BVydeqdpTw6FBB5QmG7mw4gfvKExTxk7BllrslBRpHkQybMwVN+aeoHWNoCRKP2PHxp/
GCFp5W7f9ywbRz2Ul6MxE3l4Iunqp73+aYyOTxPfax3G8/vCMEVh8Ctdup0T/N5EozcBbpqGxnmR
fBZqKtg4THoLOXcf0WXdq/jJNAUEqaEMnvC96rcBQRIHd3mq0U3JMDnB8rB5V9x+Jtz9UgEgBNdB
sr6fpat+dBiIpuQhZwH0ZY/VoFbBh5tT9RlX0/q85gi331m2mQWzq+U/BxXWQwA2mgsGRE6XVvib
V+UXemVmfoGzSHnKYw6lizc1nub5Eu4FifsQ6PDzqFUPI7KWbjmWZ77Ylk6eGSIX4pvViCrgw/u/
w3PYWIQPWwfT/gX9JQCPfnbbWvWJbArq4zzlz4rKa/bS0I0lE9NU1Isg/W18htTGNioUepSFukRL
nnK7vI7djFmmzSqbYZYvXAYQUNejGcvRrtV0L5fZOawijJWXHzZwnrgoKuALI3GTI69gbbZdh5Wx
Nz9oZLyjJjA7ClVAytBJgIdW7F9AvhZEqcYa/8aTcKRMt/qsB25tkL9WtxEEDeFgBzWkW0QpjE97
rOZbYxbwZsn9wAehiNOI7//Xc6msFWH5atKEruXUukxSX7baL6BzVajzYbZxNpUrWOHTB0kQ9nrb
OGGOh8Rz437+ieqEAbpzHkoPUaSh8EhzoOK+X6C3l+ROw4eOzp3iRHRIpjvwOIHS3GE5HFNAIRAi
uzSbFEwMiOykHkBddixoRUD9jp4Ye6SNVwxj7Gr+h8g9IQXVsvnzTiec+40mpG1mEHJQgp+mYBnK
YG8BRAYsB+BXPHSgPO0hHYkwOklCBLMKgpkLwFw1jbiPDf7mH2De4bCcjLzK24Idw1sxPKrLjH41
M//mAuFxa7VbuPgMW4qst/LywVAslrVu2nkZw9B3INr6GU7hvhNgTP+SSl2cTeg1bVz3LrZ6x0Fr
rWssQckyOzp4d0OBo8mFEPVfiRXW74gFJFLRE/9tFizng5MRg2LeFZYGtySiBTlmq2XcgDDZlGgh
Sl7vH/Kk4WBKhZGd90AkwreEOjbPQRqYRx5IDgqp9cg4s/qUWcovov//PULogMe9PqInd86jqutZ
jJOMopDC5Pypdlu5zMtGC1Hi9CSeA2Ackf/LSCpDlyev++ciIsDoLqdm75qIAHR2NkLZ72ukLJn7
TugFTA96O9kpGcGb/iJkIkz24fIJ7IyTi5zws2b1QIp4Vi/b0wWrJcIV6JTBdmiFC5LRQDk3Em9t
ye2PNkEJ66A2Lx8T69+ES2lH9pk/XT7dj86Kxpu80367Q8JSjgkH8R29vy/VkpbG9rY782s9F2VG
I0vlZ21KVLjrWHn12PYfCjlh5lg74Mor+nMyGLlCSFPx6u5CMToQPKJQImZecVVQ68MQNtWqF7eD
3icLk8Ib1forxx/xlvdhtLuU/rbF/GrjAkFFNEQ2IbjASsZtqsmIiq38bKu1XJQfw8DoIGbQBx7h
TKgS/OMiKEPSHo0q94ry5TnKsgcXAx6H3vS1UyehRftn//bEjASynIlgk5m+ZvU6ly3XewbUlaxt
Nr5zNCMInLN3r6bA3YzzZvGkGu+i9Pe+iU903UkjC7VPiSBehwr+wU4mbtkumfktc7RSS1hMbfor
qNEPMsqrfPLi8eg64ZPomydd4OD6H+b8mXM7SxJe4KYe1UmTCowBvJ0cXyDy+fp1zM2sqOkqFE0b
E2g766HNilVgXyPjGbPXow+dhaMbg7Id2bwRwelx3GzTEqVLLMKZpxf3lfKXa2JXGeVv5lb1IHaW
PUZVTHQnlXvNXehZCABt+FS3gE80je6mhGjpM2wdCT5IETGxQoPGsopbwuYkklrjSEGqjbT28ZEP
WUNkmwsjhUFy17edYf/oo5YS8C6h8dVfzb5aACAgs3yDarThxZlkcVFxf34vInJ2K6yBmE+FNheU
yhKRi5f447niyN4qRpWdQpBdLo0Znj1TTkv6Zj64VC8GD8hs6n/WH4hQRbsLdNqRxCGmLH1yKrDi
N+slUwF12YZqwTYHDIbSmPQkYK15XxJWknIRPu0syrmydw4cLzTWi1/NIykSOkVvgLZlDu0/inHi
6HslpkPOet/mwV3I5eHeDrPh8+Gtmmlp7YSCkUr06fEVou6KoEHQddXyF9IgVccIzJSB/KU//AnD
oW5qo3QBEldzh2Ehymu13lWj5I/rtDp2ezAowLMA5pLeABZq7I0535KLRPr8vtSZ/PwpRRo68JAt
ctMAmAHRpClxuIjIjZ6kG369xj436E+CxIgpzmPyhjNgx9wZJJlYHVDqWHP0chc9fhub3Nc5i8WB
XzuUpueBzzJVKr2vkmCuZinyoYNCNcYXpr0+wKT1SFy/BHUqljrNdwsbxAoZSxQZ3h0+DfTuWuyS
c4q27xClmRK+xETt76QfXtjQW551dXsm2RloeZZDjRbK7ytl10fOdqGoXOctp1tjXXOvMlCECdaO
zk6waDuN0+xXx888WQ/dPzcqdM3IF1XeNp/+e+RkQ7Z/xkH7nYVX2pKH5uC1kPgsorn2zhjEOSUd
aJcPui11YNh8bET/hicFpcF19/1MRgdvH/yABc9RMWnrUvv845Q6P90wXcPfEKnnFFXro4pMH0ig
h2EtGTy4lXgYKmSkkNRBNIV0N6QNgMVH1UjQfs9wtkCYsUXNYlWPi2An6zsVAgCpjcLbO+ZnW0AV
SaguvE7UsfRv/5ZMYjn2sWuBYd5lLYKAMDd9dLUq+sb1ip7i/6Vyp6OJxC3IBaloSIckG0udXPkg
WGt11yXUYIMvvdTgeeEghjJypagmuLcd82oXUROvfK8d/Vifft6VwL2vYfzHptgavvg3sgynm9Fz
P+GrR5OJOkO8mcrRSihZL4/YYcuoZDjjvoBnfBJFWFwkupWp0uw+Y3T5axfL4YMUnguZGwlMKNRK
Q/0QitEDrHJqoS+qcid3ALskX+EGufNdAKAWw8vmNqau0b323pd9yO+P/43Wn8YsXkJYxUKC6wxQ
PeNzgDTTXy5j5Db5PQfwzAKi8sRn+0+wMmaIbDrPRWIbl0sMLehkUuZdPobCAzpVYsZlmQCDTmfM
KVGinRNncdmFhmTvgcWZ5eWnlGimBOPhRDOhyr3moEmI+RXukIBzGCDqzEwkFWE2nILS0j27d2Wj
EfCdG2iXCsraGEzxLQS3M7crgOUh+8NfgjN7MvVu/uM04YFlT9GeE0AIazy0XKkuorA/ttXsMdwa
/m4UekhN3AF9l7OaoAvHkVzazm9B13K90HVwyFszBmIDkH5wVu3sNJNdkagLOplXGB3m32Om8lhS
17JnSWmgmjf83rCzmTj9/ZabBiLmSygdE8PVWEs+UGAsePOcStJZEs1fn/d7zQlZcCAThZjbnHu1
r1fYaqLS9VW/Kf1qSO6VnW51jZLkjl+yH+ykv77M/zMy+29IJSpqtosgjHJC82Cu0pm2d40u/6gZ
sjJdPaZGDcdflU0hRUMEy9KNP4TSw93yjapF1Gxp11WrE5MqOp5SK2m7B07XCzcAv4pEAQV1iWy3
YHjO8jjmn74O6EgXE67vTYJxt4OxnpU2esyVzIL8679qQeiCMjvXULGT7yjpK3Rtzr7eL7AqNXx8
mrSG8qeNIWi+Ufc091Q4KW3G34civas9NAhR6stlJLHYEZACxirfneu8ynuy96lkauOIX79wTXBS
iMm0t667gEH2dT9hEZ26rGTRd5iBvELFAe8esbxsfTOQJKirNKOwBdLT+ezysqnJW42gwwebN1gm
pxBmDpgwlPyKQ0xP0/qBxjK8HRhvr6qf51LKE/AxK6iQmldKINXyL34c8sA/g3Xxi5HlKqy5yipa
jy6lnFPh792n4JtzVPDL9rFRjc84Vx4fo2xO4GPlEPd/Pzw+EWyug0eKx3oXJRIipzF79mgPSu+F
3CPm+/mYnDY5MD8gQ/3dgJu/PLjQ+t5rb8GCyND7iD6CwuMFjAVQWfnnGjAEqH4Xu8Dwvr9KnexE
nBQGGcQxE2m5r7py4tj+MbYoXTY0IgSu7ezPbGz2lXi8KYqkjwvYzRS9HvGH7ne1IZ0B2zrgb2dJ
XGLKdLz8ZvfzQ0T97HVMcG4iGB36Ty18Ecc0xhkMplvjKPul21h+i8KMNEW6kAj/7jtHGulVOZmA
C4yccrgIWjJYxQabHDfLgkeCBqPUylr6ni9Tiw015S8ofMVfNrsKJsyxmU6WAp2cxGBseSSOCafY
hlIcIasPdDrdVbrb3QrpmthuL8WyWm1W6ZCMfQLgBF47e01aHbrprnmAt4GAw0iprAZccjwa0P9Y
B6DDXVInKO4ct8IwopCByyEtfb3Hn2Ym06blJLF7mRJZ6wtiF+tCbNVBpOUIeItIEuL2ZD8HDlSk
NcB5b02aJj+fmmsQeojTsORVsnU/MXB+Zcw3RW+ozoLfWBtQpzjfOb7glLg4wpSRqnCCxch4p82P
PNrGHLI/hjQcbos6GxA/ZRqHP4/gXFRdddPOi0QjzMGuEpOIZvi8wCTWut/1TvIaQs87TRv5flU+
hSj3aqwUs1smzTccpQP6W400LC7ooJLRWm7TCsgmeFokXB2+whAwcSTBW2B8nlXzsFj5TvsUTq7K
iLhrtdEy8hjQy9AYAS+tpURbhb+D1BzWc6CwRMX4m5wzEIIjIvAzB9hQ5QCUAFsiIjRvNqkgxKec
Nf/GCNHlxhbbKdXnhzEwvBJEoAGTaENb5FkIvE3ENbqdGTs49QnJgdZRxJFGOLiHy+rYNphctXYY
ajR41LMAG4iv5Vjh/ysn/CPWzwK45yRILvEmrJaUzjGv1zKm6UT9NgNKGF6Y03Akp2Nvf2mncyGu
XgTZcKUGSz69YZhS+LzEniAPec8n0fglFhTCRGOj8tF3KQF/xEZsjXuGaRsPH03O4J2qvZXcVgLY
mtqk8iDKtScgeoMzWdPGb+/q6p1SZybZ0tvcGCGJJ9xd5TaU6HiyNI1dfAr0pdqjA4w0QMx1t7pf
76xMrZ9+MnvFMEK/AHlf0wjlSJgilxfkzzt7jbey0TmU5gVLL94qds8iME8NJHVKvWu6RtnCOfR/
8eu8nOWFfTKkCmZK9+9wPzZg/YKQNvsDEPePEOtqbZR914l5xTeNQZgED6PIntOLZjo+vuH+iTGw
0TUxD3v8UzBcaAhVjnWrCXobgsOI07u0KqCuB95npNF14Q2vwynjUkUdqrfwkh8g0d3/ZggbRVho
u4nMZvljBuOm4h9SSxmJQ6NKRpBcnN/pDpg5/fI//TBpU7rCs+4O3rZpDupNep2ElZGkrHVovVQ5
Ua/R/AyrlhauBKUdJ7RZDxpPHQN4tF2t/RwBuh1X1vlOZuJ7Eu//ZCpy3QRcLq+avERhDILVR0TT
e5c8omTBDGJBsDxG+ku6CeP2MjebPNp0WItctcaJoc6j2Q2cs8Ow9qPJ2rbfiwIFUFnsvoIrMPnc
Ora+TIXLGxLHLwhzFlZNpxbxmF65IsusP1TRq1irNWcGC77GavdkyH/XeS5tpC3AWBLqoXBpQvOH
Cuq4LNqmOkRqp4Ka/Er9E0Tp/WjNKBJnCBWRuygQeUws0tBvbIWd5OUVKJ1YswMeF7b0ZS3/4nig
Zds4K3oVqwf5FcqmeH0HO/Yn456GvmA7EC/fsyKBV46YNNVzl28kz8t3ivgIMb95b8f2rvXTlPJZ
kwJzSYZKqAys1m/2LdlbW2PEslnK/HzOuQSmosueeejun9WHTr0fAfu4WAGHb4M8TDQUHpm9PfSb
fE002veSZC8Rq25LkFhjjVU1ohh6DC7D6QJBls9TK0E4l31OoZyJAwCdHzD3/Rlbq4l0E7B8rPG6
uYv127tnU4Eu6Mt2c0TdRCclxr9ScTD7YL5CWPiojCNRU480EO+4vcueoMx0OrLEWWy4G0hXEjFb
izdO1zJ4LO6bCdmqiYjK2lCKfkJnkvdLGF6OWnl35Lqa4Mf99XVbSwLXzZD8X1/mb+Zf67mxsHxN
oSaTY9dZzKYwT6LdnOGFje04yweNhms6erxmRu3vIQUu6Dqrx1exfSj4wzmeAjMKtqTRgIpf/mWA
E74U923yPd59T9HqZPJQKE5W3LhzBE5Iq7msj3bYB7b5ZGOb+t101H4JMvm0hdZCCNgn0EBQW1Op
0hg8sHxLE7aceYQV9/aLkuPo+33tBv/hU9JkQNbnKalPBn3Te0wAt1xHxJUFal291EK/w+bd2OQX
L8gd0JeH85cbOmkUoQdt50eECpXBTjzvUbKpqqHhWBxBH56aqZSRImMQcdsfwNRoD7BBVFWxIm+g
KccoVcs/8DkQcMUZlb6Eozr2lS9hPTAzopXUDXUO0OqRfL8B3D3OTBOqNSFRwmVjItb0R2sLKf5Z
CdUM4Ml+RvWDfsXfhTvvZF1Ai9sUVB7+anmdsBcl8EaxBR6qXTBsCIqA+l0NIBL70nJm+kUft6/4
G/oKnkmdqbN0KGYx0VG5Qi4JktNuHm18n/WVFx18lV80RFHdDfX+YSlrZC2sZuJ2xivANnrql/3/
NqIYZSc7Jents4lHqf8fwKZ4Galt3HbSYgm61ni71k5vwbgblbtNxE+K0lHCvVj91Jt/RBtEiRaG
D84EJ8hufm0oLBx/ph36jI+ab4UaG8G3ARTfajQyjVKgM48jnjlbVCz6eEv6i8mvmZRGOWM5icce
nLuPwWN9aIdqcE+8X6K5ikeBWzRazo88SxVftuGE9kPWOBR2doW/3Sei+ddCWQ7L2I8JoszsMHsb
Y5qnX8bs50tF9hjhPAH+5U77zRFBmWYhLYYiJMLIq6J3d9H1BGhWFPNi70uKgywNk2XnFhiW/rlq
831RPlfiTztenMXpdq/+2kLVxsAINwNM6vZBNrkmefR77WpCfDKPtPaz9J39Xzm9JwSfDf5Zv4fE
zbhN06W/Y2twf1sMd4819to1lBke2ranrtrzXCFvKzFA2gA+I3XZiqR+vA6MHaATSzsxD1wAmin9
uoX7kfqogbqGV65FEPM8mm7oLeUW6KJJ68YUOgXGqXusWyYvmvqLBPnL4Mbg1+oaw9vk5U0cmo7q
z3lASea4JasvVXZG4CgB4BlKbQDi0oxKCwQS+VE9GuwhyDxr4ZwN1ZKdgxrWod+E+4lFxx3+WTRM
ec2hYgWPQVXtYpSTpcJ3nVwny9vgBI2w+sV0C/hFSzumI98723xNnO9E1cFX+0YY5/g6CdIl8J5Q
sPpVF/w8bh+4sbzasGYmGfRlw3SnxJ2SdPr+I+7YcVSmREKCfrT3bT4+SaUqiR146sNmFsh2e0SY
YosShj1CMv02VG+O//I56Btr8q3ucnB3x/bi5HvLMmvYrlNtXLVvJtgSXw3DL1f1+A4rQ44i8ZYc
wamzszDVQ0lo2qtz2V9AKfeQnABQkeCmmRh7cdodSceprO4G5q7fn35iLLo50uSrKfPoD2Ulpuol
M2Ha3yc3WQslijXLtdKF1/XlSInhKhkr0hUUCPX2EMcdAZpKiFoWb1S1eDccpLFj5nuJGxq0PO0w
lEWP0IuCRikWhfHoMJybUacJ+W3doFLIA+3WNO4jEvHUSeYkL/N7+KeAry/pmFyblSal0mLTdoob
LEQdezGqx+1spPoLORNsI6jvrXfETeKADzz36e+DxllCmHKTiZwwTcCdTK3MV4OtPtuOGv5Fra3z
sH0wOLU8b3jZlZyz8XaoxLPrYkpRHA+fLRCFODgJNbv2zj45mvUSMhtOSH9E+q1PdvpohrgIxZHD
XHvfI8rNpGOO1wk6bBNTKm0pAL2/V4U2zCJGJtrEhEfa/7Yjui+wIfOSSI9xvig7PciUBlzQ+JA2
lP/WgR/H+bnhE59LT2llEN5p0dONnzxO58S9D4lBkm5mJaKcPcPidkzhKRnF4oaNRRApZM4DFa1b
XQzEmtD8doTJtWeQKliNMIqxsMxIgU2kB/G88JcJHBubSM2c8hvTvt5j6jQHgWNw+r53jnKe1nOO
Gdi6vK/BIG0YbLtumOU2w2lhDNBz9+bmQ1n+bwTEF9hiHcjkbT+RLYJnMDBo0AvJtDGj1jd3+NhX
xkoDkJHcKmI0VbRn2iUAPqrJa4SpXE5ohxi0jzw02I+PCyH2fWUfUMwyhITHQdI9URgIC11ZG7/R
wb6NH5S5h83TqRTcEf3sszrjwOqL8WIHroI5o48RWS5JyJnH6jE31G/PJY0+1fJGWNZmE7uBalr3
3bujGWLiuc/6QRIHtlwR+xWDXAriiXsOtuOP6AI/B6fA/q06SksI2nGy1G5AhGUFDYGB7lTDd0QM
NXLP42GWsDSnIIWaok2tYRmni0lJGWQZ0za01LOhTyqsnyXinPbeoxaXSGMdwLfkhELtz5LtLh8X
KquEdAQYI/OqR4u7FsMxPsRKUFlnZhXgCi1UK2oohDonWZX+uW116Iwq4MJs0aMTFWb8zEHDxGin
lZpF83Gn9ef3SOMhW2Dc+TJtHhz76vPqNRXLSZmXpQ8/jrmDhn8X5Mk0UtQILgpJeuLDbWrNWJQz
BQPWVz+4bu5apaLpcWfv2jn4bkjg54rPEq8FuZ8vzm0bwtXBHVqJtcVJWTsbJnFQHaWVlmILR8fx
AdhSwh4DBdxhkrDKEXmVCC5mBJGKqRxv8QIDUU+MhVTgnQYzeey7STdb3JXJFMlH3h2h9X2XRY0I
DTztJd2QKwXqaRHItU1jCu8BAfAyP5m+U/9MMYUzB6X1W/rR5Vx+6/9+Vqf1qnZTToKhOsmnIPU/
KqL2P7mws0Eztx8IoOGaaTDxgIrK/gVlqYZnYYu2zVL1apftypsuzjqxOW0XHtsebC6KQKYKzqm2
m3B7ziXb37pPOivV7BAqe1S5hNwnbueja1cmh7atzkeVzbktY5SjwX77dUi03Hh58UdV1K8ghm2K
tBnzTib+pZ20uBcINL7bcM/EB7tSuVAoMRSPh0S3mn2sKSvuZSz6GNZFuwtGpHHUcw/HxcftOOBW
W+kZ/1f6RUCEAOK5GBW0s24Vn7NdQ7C5TAOP2OuZw03k0H3Hm+RMsbPFXRGwNX2cEvtZ12BO89YG
fGNa5ECTLVFKPFvZfh5wxM/6BeWcCEtEX+CBTlcfV3zgeHdeLTV+6uOt8B3/z6dyV2fy+lXMmK3d
yf3nKtSy/AxzixM9KcD3EPxRJkw+u1ZZhAKIVuEDSvLaiNF9x0I4VASgOl0F9mBoYS3S2eWfuicR
h9GgqYT1XcovtVUKArhAb1/L+AtUx4Itn5Z014JrwdNxtp6CL+kmGlBkXc5uEiZeTIlZ8QcCaNiV
PNmodykKvAIB2HzYIpoRoAMFD44fpGjTJQyaQ8J+zNM2SHARWfHx+4MFC/rvtcoPZGclTszMRLd9
q9YuzmX3Aal7I0R00kRMP/8+QjJk6HTpOZIG+UPscuixDczvMEz65fKONsPkA7vD4d7galfPLmgQ
qiqqye2WNIbvvVgknWomAFW8O0uPSqa6bQ1aOA93+QTLPvpzVQvra+L12RAGwSbKpZAO0uHWTL0g
467ktmAnfZWjJvuG/86zbMaVr5Xy4E4lpcpqp3G0knPaoC2scZnLnfyd62k0RN3WrAibLCP7Rc5X
qxBA7aoRSJn9yXgURzl3N0+dQwMz8TF/ozW41ZhOhxJTiaYKpk+nMoHhrxA/wNRbJy8zTa5agtim
bZ9H9MIICGZRUA0BA9AfQjTg/zzqZm3qGZbtlXH/B/i2RchChsCCXUk1FdQYS1ibAAB3l1U/N8IO
KHuVxtQsewmKSMRGL+qRVQJesmlvEpXG/IeqEZzPUjlg5MUm+sNC15hOT92y8ah9pqThTPPylkkw
QooZm23e24cglhln0lovIPYTvGdliZy+W7GcMimEw0fpyZJj/o49Toek9VuJIDlI5zQBjw27lPTM
xJaVzGOW3W2oVEzAenyyFbbhKO45lPUJDYsyYMr/P7chyGV7g4Z4ZGrdBq7VerE9pQ88+/u44WOr
QPGdOPPF+qwwnl13vinO7p+MMnqz4GzokOYfkYmTQc9dE3DbzmamLHDUekfLAg6jas1/8BYDxewT
qGJYVuzDzmJzryb50MR9yTF8XvgMclvfuSx1Y0tuGDxPA0HF5GlIVxhTXGDHoIIpiMWWru8Sc3Ao
6KVwNBKPo2WvNTj95kDY/R8NmNbtH5PBYX2gcIyCISF1wEL6tilfaxQMgwYoM1F4tVtnSEn2PzT0
9mXI+OTUCy6b+QeHV14FKq/XmYJNrnupuYcmQQbBIGPoNisJrfmS7+vx3dViQTff0llE+gMktNnN
a1chkPaS0LBeCqwUkDFlpx4GLfy0a2X61jEDBYNjbRbmWL51POFvKwnY2qd9vzUPZxQFXIacKoOU
SXhvasmmtg+PTsONPhlc+vxAfWz/tVPkJDQwDBhzhlxgQa2Jruha9MriB9r/5J5+5g0U5L5N+n0Z
FOOFJyicS76xc3ePBOxhpwYpkkYUaBxzXV3KAfI3Tlc14lfhNBrXDQwHthZROOnJdLur/2MnSTHD
7nimUJyLy1zRIC1ex1AW4SIEgLp4LU/F/wRNSw1lY4V6tL59+aCLPrYBASNYGYEILfldTY36OUSn
CuxIhEpC3SpCTAV1T/eNDL/hqEyltP6Jg8GWd91M+plLrIbNAtsQDt4SogTii8hxENruMmviupHY
Mb1fufR9SdlFn26fkLHV5Ep12KH4BanSbGWVYUvJtu19LqA5dlyoUAwvbMTEo3KmUojCqoHhCPxH
HlBHDpqA+sBzff1nlgW1QMyZNAiJWK7eLhrNshBn7T+pLDGFtH+gQpDJjft3fCHDadxtq380k2zg
JpUt1r5GTV3XFwAjLE1PIgUlgj2qHA15Q90Jjm0c7ks6Pg7MlJ/Wo1OGkRHXJr102yqJmb5E5eZS
OzoPPR6YYHUJEEbs5YvFtztT7orjM+wuFM6XU/R4qg83i8b+Ef53+qGb0BJfIawD5FW6ODa5+wdw
4I/CskoGIzcfq9z8vCgP8ruI6fozUR2bRjCacQXbms26drxINOqtRp7LIoGs3O53qdWQCrN63Vnf
2786YiP/FcjbuYOymzDWf5kzCMGKhcnseTsPoM09jq5vdZNfmp1V1bR8j/A6bJb74ova5FG4fVEw
lgO70ICXDrf3aUtFCTZa2f/RurvQy/PKswlAR0+06k5rVEIQR54f5ybflDqvNi9vnZJZS35zjcm2
0cMFCMq/25oEQa9lKlwOWWfCInzykdN9bPS2Ew47j+2guCq45Dg5s0yLQmsKi5EKOfd+VRH2pOXh
a9x1kNxSzy+K7nAXEPA1Am5Z8pdabTl2c9nBNtrlTGh3ivlUzIAi5JaTYmJGm2M+gLyLOjByhQ3I
+dafN7GHIx/P0d2Pn6pJk+KjMoIc+hHX5q/wUwm1QLLqEkjyEW7qe7Fg8ftFTbkkha8KuLtBN6ny
7+646omAVFd1v707WAEvvIoq2BL62TQUhL5JDJGkbj9HzBcyybHmLCFB3mfwi/0bKXTaZtEFZZT4
1R09Vg1MpupIIWNSl8lbz3UqNBR7a22sg7HsDk1osLio1dHF7+i7jt86f1tSX/AJUq7bdZYpn/Pg
d0lkUUQxnBNcei0TVTmanbOE2myxhHbQ2pCpLj5kP20Xjz5MaNIGJQmsXvcPJhNw4eb9h84OV7d7
EQXpc5WTakXofF4SQCaNCDrB3zyTMZp3fCD+gkxmmxIUeuq+/N7UDk3+JZWBIliStw5WdDl5j4s+
5IrxNm56DxynSWQaqvVhKMFuApZLdsMSArTQI2wY7DmXVjyCjLCFdHI8LHu/YmSdTAEVj4eMutC8
W8Vgfk0mlB/cgPp3uvaQNKjApYR85LAPfwMs9ZPTXzeHSxN+8eWJ2yv2KKGYkZ83gP5mnWOjV+Ew
1lZWDF/trH6N6L/g8lnNRRzi8Tk6rA/YVNOI0M0zZyUTQ7izH5rj54TaNA7VqwdNdFc5k5yX4x8m
q7gMFYnzLrCI0sQh2JsashvDUPuEWmJxzEeld9KtTqBjWRgG7xcnLZm5WdFnloKeeeehkhGJm0TX
ZC8Ur4+paFh066emLkLZQe/LQd4zpCFBAneRwVFuvplObGTZmD2CFUsI38qal7ychZqIrVPDdFOA
368M97dAo7+/6kF8WwZW9aEmnvnG/Qes0LQlakJZ5627eoH0lgBtsc4ntdVB/ufktamiCjKo6hvz
UrI9acddvR2P66bJ1/UGvmxTLEEelfdiQoIojO1dObNAcHrhw4mg8ReBbUM5VJbtoI0ajVeDscr6
a1GgUb+jYClqAT0wbm4LIWK058VNlGoqYkSmcm6c48AoHZgOap4HAtnol2miniEwk4PP39s45RTJ
6wDUaZjQv73IhCCpW1dFdj4OnfEAr1b6QOARfT5nqxk3IT7ShdQnT/jVwnOudhxoD0V7txInkZ0j
wq/Dk/9WEP+MmAqRdeDCEsRGyKh0NaQUYPkLiTYRPD6q+vBZX+DOVr3N6cUo8qR5j8EfLwAPqjv1
5Jzwfw5t+5cN2VR6XWPKGH321BC4x37jONI72gUkH72fcSwhWri0Wce5amLtGyaxudgtaOJW0ZV+
9cZmXXXELGOaHYdPJByU37Iewg/HfC7it/Pfe1HlnQUPr+yWgKPOIc4258cPdciJI/i3S9/b+8z1
aSKu2zSpioHwndb1+OkJZyt0KbtTFrCBu5oZGl90xtSxRrvzGDka+2Cies437f2N8+ToCzD+/kGD
YGXD0HQ8jowjh3qK8tBWJ0kL2WNpAJtwznbdN43DK9a+EA2GHU3O3kIWESjCEhbr8CSm8SQ9grUW
TTP1oDQt+EaaIQqIBevsBVH7Rdgu4qoK/bwfpF6KynRKnbkC5IpJCo9D7nAMqH2dTCkSJT45oja/
xoos2pcOVSAgHGiVoniSkB+aRLw/jOTPQhmelCAicB4Vd3WVTtAoG6U4UqUnqXYYnJTRWhz+MBrt
HsUYps5/M95iNbXsRDlDSzCcT3lqDj9yCltB32Ta9DeAKJgDMe/HSDB1U1HuBYV4UrjuaKL7xs+5
0QAJTysLQUfC4L/Cee8j9tYbfz9JWYiGaRmWnVVjjl2frGRNXJGEYZbSKAw6fK4jn181swhi9BUW
TYmFhcB9TlGqlUVGcd/p5Y4p+LjUdpcy/hoRYlfORsfXrh1aLiUd85ffmjBAnWHtC9jI7PnIlikT
0Y5SiAYJtEBVhccIp3yE4ec/ql3tfWPthUzDNnrL46UgreY3yHIbqfQymGcAu7vwvHJQt1kRbw2s
tlqXmLDLiBAJ64fASfKo7FJ1e1mmhAOWzZBUoAD2CGtJq1zG2FKhm4Upcu1sfjwzY2clF5lw8vjk
QMubFtBSQ0+NwAZ5fLGj2KKkE8nN6Ahsi5Mqg51IAPFuetEBqJckMHj7L3YL7Qvxt2rj4oAw1jpS
2MxnOg6U8pMft0hcItEPFFE/bawp/bSrfAG0zAOsZKMnfHIRvCAZqzieDghqm5NIWh6oL3e8enRs
uVOQVy0ZJR3rLSQKXinMwAGzl2ci2H8Sb2JvowlK52s8FRY4EMDNv6fiFGARgQTFDjL0OL4il+K7
4Lz+E8NGrAMwGiqDyxxVi1wecTv8Qo97rYvhsmszi0E9vvJzDGFyndKJP7/TeDS1wcVttdNY94gA
2tn5fDgWCEpzvr0LKHxunAGnwW8rBSnc9DB0G3/KKpAuQxP94ciQb85i6gX42ZO5SyCSKnXVz1da
QgiBgSqh913UlOkAxLcLpXil5emy8A8bb6pXdeXXQ+/s9OwFA7TY25Ceu2UjiSdTf7a7LZm9qjQX
/Qdo3wIDVJmeBuwF+pGlllqC6OLkBfw94gUbXhDfjHAHqxkfXvbsb8bCGg2gmyXbeP+WWm7Gbf8e
nHbs3jNyN0T+w2kd5otcYd0+0+kG+G92m4YGEsVoOIKfUgvVYSK4K+yUTEPeXEe9bHt9dnlDLmwB
whgaBnMLhmTm5nwIwpf9K+Y3ImcFWjo8HQznIfa1eTydoa4VciHQMXJPRnJuip0rq0mnSv1ZHZ7D
ZnkJiUWoef8z++9UlgeRcZ7dcuUYHN3d27PEqHxKVtb02c8v22enhcy27PVJu1wuo+Bt3imK/2PB
dQF2VZ5NgEyN4MzbJ/IGiB7JY8LUHMiq4QUKXE3STEfcfmDQ2GvznC3JvewM7j7j7d5xBo3jE9i1
aIWaREDo3ugio3BbAMzRl+lGF56h0rXFwL/QRSratSf7uy73OtfSYS/6HtcSlq8tijNSQzopZUKa
CcZbeR2D+WAklivvFdIX7G5SKrqIBKxLdCSfSwHQxnhkqt24MR2DsJEBd6gUM1LG6/oXaJ3Ridvw
AX3EUGZpoAvFPCkyc03CS0yUYB81qU9Ett3z2ywLeOVUAIfoSEzN8BTcgNwYAlwLjpUj+SdE8g18
jcpn/0UFOOJ0I8fmQ5jCisSbRqi0g5tiNiP20ZR7TjcbWM089vnpCwIYNF4hpT6nu17Vh5jKaCYP
ZKjl1ORGanhi1Q3LWFnMcQplpoockFeW5FuB5xzGB9mDE9nGhrnp315MiTvb0wUw5cZB4Qv5kLHX
H5LG+s5uOH/VAwySbXWQTgJc8ykozM/jR9U87DFENKm/lDb8bkeyML4njsbPuFL5pjK+L0Ydgckm
xhQIYlPPyiupgjb7rwP8uH4HqcTjvWUrxetSoU8wvl77ARcTvrIseeiCD9GiYwl/kLVnBk5cLi00
qXJHCWqZmRJE2mD9Cme1T0ZmRsDZc0DaaiF9IjA/8+lb2F03zZFdqy6FL0Izqs97JQUezOVu6WHY
Vx8d9AUb41Ov+6MMveicC+B2AzgA+l0UvAQHdPP9/9qAC8HoUkv/9bIhVoj/G16NH7Hrr7H0pDTO
xNnuQ9BNCekdrgXjiI5+E0ErxHbDNS72UK+g3nZ4QCU0TyoZLvuGClCnkEAH0MLa9tH60k+6Uw4o
2xnpSFsnyvZYpdDfo8NiKp3fJO/TrHUmAGnuqNippgkKxEvJa2Khok5frHTjR5SgmYhrWvLrF4Bd
kQlhZ6jj8oto1LYcFK1dcV2YcgVIcdxFCtqCR74SabV/T0UnxjnudXIGtJbqLv6IuKMzieCXe221
p2fNNlMXIZo9HG/O3UxkKpe2/MR//EEPV7LGEzXxvnPV+Rq2lC1RsEHU311ASrcyAFVtyE5HWvjn
9y11bZZvFcTKB4/CWGAjTaGkiVNb36HwL6oTy93wY2+aGdPz6b/KrQ+t6LQxGofanAlpBuqAjP0y
M7Klzyv1yBWcbNovxm7EnOSSlcYGQnDPt5HgCrEtKe6vbZae39Tp+Tr14SiPRzFHqa5ZmEXWa9YX
SdpDKEy4P/9ZRjJQKP4as0e/xHuCGT87MTkObXJJAtrHxHDkiFp8sVNHaltX8opiM90mFfYZlYMg
0xaXDNVdfWch7Ae5f307rQaEI37kW9CecnRd6ySa2U6mWrJx0prkZprbMYicM6oRpl6KvpaEFHBS
IArkPu+Tf/5YZT9hnNB9P6OXs2Ki2YTSDiLppDxY5sxDptUjV8cLBrCg5k040kKiL5oF5pkI1Sjr
CkIg8KzEO096UlJP240qzLPllONLn1y2HmWzlxxT7QAzk0zC7WhcWEPO1qZMYN+JgYC/2rUSkZ/l
EH4/p+WvmF++CdPkXqFJlm9WsP9Bh4yhvaCbpxoOUhpdzvBWjpPBGyoLNo0+UrVfOzqufaJlDuCT
CzuaK58bHKVoKK7+/54+0hTkMtIYW7ty8rsNsXA+PNaWhz7V7JOrf+V94QrBeptk06eV2do+3VQw
ujU8zuelAzHsd1iI5a71wE2ffgS+ib7Nfu3PhR0+Ua+O8fK4cUdo6m1bhANdvWERgINHOWW0mnrv
fn1BTP6I0wF3NL/du/qt4e/NefN5IElOJiWzOiv80xU9CKkuwMVSh2s8zG/gl7u4ozr5b+KidTLC
xuYteziLQrV9I40ESWDxsk6C6cywov5aydlRvwLU+iK/qu/+57XogOQYfz03fRfrLXsVtdVNrpO9
Y5ODjoQFQ/QEdeHDegi4CyqJps7/VjA8JgBhR3S8FuYR7VcUxImqFS3t7L8dJepEfW1s6qcxKpbI
AORamdZiJaysFRdLquIMs33d0Usb7M4rT7uUlThqInYqox3VeNIEYk++9uwsHB6OCs2ft9QqWNl9
FWcHq5ho5LOunNwsanjiMs5+pXU2OO4q0fw2O8aVjYX2kE1KeTBKtLyOWPTPTUxag/qM6hKuEGxx
9DhB4HwfD3d8PTHdP36A/x28N4GU1qhyvzw1u5f+C+PcYSzuew9koQK8VxS6TA2qnlJZTFpQU7Lo
Fnyxd2jb7wzNm6+62SmP/e4w/Ln3RaonXYn2xHzI+7YZLQlYZsUChHx+7OvbKCexravSlWw/z1Gi
bPIX59kbSK/1TujlkW8siKV3JkE73I0gT7tZVFDT5FNaOlmY9G/5mCZLaicpWUWDsf8WvI01XhLn
71PGUzdsT6nB1rHWDdFAqoSIwi0rJOcPo7w410Dmhuv/k2TNTfUryLutBjDB2ZbMJkzhWJ2j+4Mm
CQrwFj3cAwMRHtHiRLPYb1LQQ6+0GhGrW5l3zw//OSV1L4+RpUOjkYVKw2IIZe94xDiv2C/0JiQz
TRNmYnTrbhfu9ZQWExVEEBBe7qrw9YrF+y2jW0LxFU25ie7UwKXuwaba0bLJA/gUEMpUhYGwcfil
vgxEStofqIR5/SuI9O/pwWVCfettbMCwJxmvYsRqxLZcKeQUoN7SAm5jUmIik8mSEi/6YwOcWQQI
vHghJG+SJnPcG8MSo6ZSO4/8KGZ8OxMxVXxhokjA1Npn9TcmUymO7/NOaUyw/Ey8G/7PMVqo4fkG
tjuhgeI6dWKkYWuXN64ajL4JDk5JOewT3C3z7MYGpceNehNcu/wT3XMAzTs6atVzwWYyrhEWuBpI
nXCkTjTCYx0JuEJ3JOk6VyDvZyHxLeCbrH41ER7y9PcpsVpnjD2qLKcFpgY/DxnwrqDRmGLEUsJK
Guvhe0K5eiUcDso0EdKyMoXphjgRmna7Bs0IMrHchDPVqkuALCT9XLeRfAw9A5mxfrbdukgQ5WT6
qje20UVkLNn+4xc/JkfEE8OWKMzWg4BQhW4gQAPnh4x4FcyFplVV2B13TMlzpuM2O6ksh7rhiqH/
wh8FBDpt0LwhqybOyhmv2KbXIaXDquW2tBxWxW9xnUbPefHK+9S1fx0mshmBaUg2fSqoWjLo41Hr
RT+KtnldcpNATPwGxuqtTOz8wcYF7CO2491uetlkl7oIhUxdswwS4oNgAhmma90bRAyMGp/EtQCF
jLZW78kh5WH8PtvT8D7p0j5XMcTPHhXViEzsSuTWOBQjuJLDnrdrglChP3Yfi5EDbGQqIL2AKqC6
A1o/5VZ0LFgFfzaRW+UpCnF4oiCHTdhBSDxFyIk+67qsdsghhOoyD41RFzYi4XW3HloroU0VdRPs
pwxdhS6Ow9AIX93HjDN3sp0Yt6J+dbvFHUhmWjUkYt1weAtQd+hrncvmAMBGsAfcyi/TRPl9JiK5
H4D9qyWw7xbP1EZhYrbR+FlYmLP74hkWf5SU2IcO9UxBIElePk/ZezbuuctdVjcGoMNTth4IGvD7
55kr/SpccOHX4JGrrngsYMThvDNRhFBhiMEUw0/JKTi6f5oYtsJb5GxfiEyAgBR5eChfZz9E6Kei
b/ao/zYXMsFIcp1NyphgJZqzg5FnB5iu0S38X4bBtGtsOuH816Pjh0Fvb1NpUAQDoEzZWYrSh8EM
fq5j+kxNFJtudxEgJX+nSA8W5EiziU4DBEoF/qvU7XXUkNq9ld1jUPAR56iHMENMpy+QWPfjUQZl
8cFywmTr3hnsmbtSBPxCFUSgdxe3qoS64edZbF12nMYmDIISkC/xX82FNzmX8IrhnlKXuOTv2CLA
8uFkCYk0xEAhhIaz1YArUM5Bz9cULerMP54c/MzJV3kSmTeFAMaXu95tLQVNFkujoP24gWv38SVI
vQvfX1rE8P/YgGu9pOemDJHD26XQZOWG15rrZkJCJEqnVlQ+3Bj2GqhqTeirIdXdFjZkI9pSZ7kj
bj1ervIqILcxsOuzdeuRfLFz4veDT9d1G8ZUqtPCPjqWsorAMMQ+84YIKEBTTmzow3MkU8gp32QM
O9RKPqKTQTKjvRKQ3XE=
`protect end_protected
