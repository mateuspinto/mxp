`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
r4ClqoQrkU53dtVF1k8aM14MDBumTSTcvLRtxlsY+wTZqTqE6dTVPzPIHsUF3CV9gekZtBxUxb7j
sEXwIDqIsFnWhzls1VptOdK1kcrRf/CfGwDyF3noMY4ViyNv/bGi3/ZIUx1XrihO5OOb3q4edFr8
NWew6h6rUtJOw3uxt2bl/LGJ+tAi0+E+6zh/NLBpcWABZwRUNCpN4WDGOEL2eSaOyLy410kiwmbG
uM8CQmesiXRx2ZIxyemSIcVoT/Lo9S0iQ1enYMREQOEpSuyjc5PiZoKn6eIEuMDSkX8cuxURLvVS
piL6qGb83yya+VRKx1IWtDe+MCEEHsOuiphXHQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="iuKwMJSzpLX9hPp1WH/8LTQTwRQIkorMckuP9+B4wyM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
/jBv7s0E7hrduQ259Ug2Jsd0K2hqt6jup6/1PcTPSAZGbUp+WvFXe3rz4rJ62GAB5zDxhx3XH7Jg
0EacSItS6NSsAaTyRcl/F8a4Z6QHmw28Wq7tQq8rmRLNdqbOQiNl3mSkgnBCch3XTVmjap4M0NTE
WrcrP+DmRG+g+qVos3xiGJrB4Bzm3FULADTae59dp2QuTIkr+ZKJjoybjqk0pl83c76+PZ22kiGE
ptjET982JNkoMgSODHnX2xM/KAuuOaJ+xvIH7klGyiCip02rhs4hIIO7C/ImV4Te3N/A3M4WJ8LB
zybUWcGUbEOl1Q2KzAazctJKZuvq+2GrkaQfrgC3UnmrISwRwFu9VXQfWNeKZxhkK2dB9JRMg+ws
pB77D9e49XnAXx2eZMP9vcTev9k8bLVp/Uw0Xlh5HAAcSAE9/hFNkDVtT7kdIWxFPRMG0Da4Jlau
CEHLdWTx1/mMWk5JcmWOJ9bRzK7mVG4Wcsebstqbf6WaHMeo9mSRsbP+2kOlbtapWxbXIvFlRB/Y
3dzToCnROHduGV+ZyRtTY1hQmMWm+Ia58vb0e/bVuBv2CYzhJxxzS97iH0CkUSJ4Q/vdW+AjQi1S
aArc6BzYelqrCNuRdrtlWq4eq9PQ/xIXN8gaGe1z8pXo4D72pWUaJtgDU5kfNdIqQLxCk6bw1Lw5
U8tBQx8CVm70I5qeIyN0JPTOv/eamGBC6WR22H4gOTqj5kWAp8qMJhxabzAp2GIlreF7dYbnuG5Y
AccTlS0Vf6uwFnMgpJY/nD3p02F0tOIXw7ED2eYI3UErNGE5z+AljEpH95BAO3VdkJo9qeAWoWee
yjK2+2jpkSxhGVJRdp4LOVQ1mehNrFI69lc+6bjh/mrEaBHIBMY+kKCRWC9s28HdaX1X7//mZl4i
bMXbrnWPo1vIr2FLmLEm+yBoS6GGou4qu+QlkgCDqiqW5Q8iRGu5TQ8XoP0Xr5lwbSUgp4FnOo39
Z3k2Zbwi6X59my+FuGTu0V8NClyTBS0a62sqquAw9CDMMnUcA3jDo/hvxZuyGhQreU0TLWvfC4on
4xFLEU6X7cfuGk69TES2XZVMPR7XR2pEBGe0TH3RSmktGtdCwc/wiMCf6lVEPMMOnniW73uAK+RG
uV9qdoTlWdHHHXkJTTSmwq6gUZmw2k62UuOrm2tOpfqJvPIVzWhxaoJf1IsiM8jHR+aPDThL82ko
bKGTSdKyCwfPeAEbVyixws5JWd9xSoHrvYoo2CmVrXv9wqG+e4jgoy6tnEKXxPl+gLxwYkEA3JAO
XFFufoSQy8xLm376nqjWxsIqp+fFNptvQUjqlbxXY1fJ84aUNuBWxYBlTuInNQPIp+M7u1c4eRm7
bqYURc6/uJENHohPpIdit6LdEfmmjmluBvCR0hB0vYfoHtgCqsn/CrmNy5TlnZpjO93tFbTpGcaO
Xi+1ZJu0I8L71PJRir8k4NFDI1OVD/4WmMv7JTA/cigm/0Maug==
`protect end_protected
