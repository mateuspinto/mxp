XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���'��q��������������}�ڬ�e�G� ���\ ���DI���\�.���!x� c���$K"�L�6z�
���B��k�U"թAli�a$���G�Ǫ]Z��=��Sb�b��ŷ+�M��pL��.�F�z�-`���3��%M�����|'���-�r���}g%(�D�r�S�}aX�f2����D�
�?������%*�P�;L,NP4�����Q&X7���z�$��W�/L&����{��}�3���=\)�}��p�P�S�4E�%�!u�R���]����y��:�ȜaH�9���%�6c\Cp��p[?�ƳN����V�}]��af'��3s�������a�ڝ�Ol�L��|�����p���p�E��]uս#�L�5���<|�������Y^��N�^d~�ߔog*��@�Gz�[���RD!�M���%K�{ٌ^W�j庳��-�N
�@*%����%�j���=��N=�!<�]4��ò�T��gM,ȃ�v�w���`HT��k3�-�f=ܣ�5>+�G���Ri��k��bdV0�@������z�dOZ��w})����Q�[����QB���������6>��Q�0��E�}㳦[}�<���0,sa�֗P�4�tW ����M�R�%V��@	�h� �?���:���\�w�W`l7�z��h�ô���c�R�D�>=���ҝ(3�@��b��"󕟄}��A�el����#*�RO���K-T�e
��JčM��{��SXlxVHYEB     400     1d0���c����M=9D�h��^8 g����W�L��Z�v��U����T����S�Xd�+\���-0���Q)��DRe��Eh��\fC=�����eC�y�g�	�?��q��m��i���xd�o^i$n��M�Ǟ#�P��Ѩ�o={%�����/@�C\o�я�n��h�����E�\S�^�ᨿ�Y�� �n�:Yak�O4�Y���}q��E�.;9���>I�1��U(�C��;�<�O����4�-����fw�Suڟ�⑯H���1���-.����C*�Z�� PE��ҏ�ש�9pJ,���,K�����]���0��&���{��/����wH�3✠r�HA��74��R�L�ә`'�N'���	��^�$2	�#o��1(`7m�pym1֏�1��a<�3V��k�-O)Fo��oE�#���z�t�e���[����x���$C�n�^iXlxVHYEB     400     130O��A2�L���ژe�q����J���ehƪ
d��/k��-@�n=6<��@���x&x���~&eN�4�O��f,�W�7bN��IG��s�q&����>Z�X)nj�+��j����0�Y���
ox�q�
�W���7���W������10Ad>L�;���`�P�����6.u�
���Bn��T4*��7�d��x�ȹƺ��^��?gy����+�����S��)�8�%S}nE��E�T_�f�Y�FRncB E�Q�_��1V�6p��t�?~6Q��t@�>]���̯��`XlxVHYEB     121      90��߷��5�X�Δ���A�̗�}�X��ϋoż�Zq�`{�cm�s< ���[��p�˒�T8Z�Dρ�.�[�
:�a�j��l.2��ǂ�W�X���&ȹC���G(��t!���t�\ޡ��J�Y�k!����˷v�;z3�