XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q$D�j.�}������$��+��&P�!v!���qUv�c�{Gm%��ZM�2���EZ�H=:�c3wFP"f�0�1l*�GǓy����RhoB��������\��;Ԗ����ސ�"�&�j�����.4��K��;�N��X�I���H�el��K I&b�����i��2|e6*~7�=���x�gwm��nAm��#m[�K^�xz�nʆ��F�娔�~˞H�  �?j�}&�<��$���!�Yj5��Q��d3l@k|$�L���`ŭ�]��Fz׫oZ_������:�������s/ʈ�x,�8c[D��6���[6M�>��'?uH�����>�`t��e^�Y@��ڪb_K����������� ���
��M:/N��km�L����@�G*׸#Q����
��&�>�|N�	��i�tX����� c�qw�g���[)2x=F����|�!����C��3�Lt8N��t�:�%�N�	���5��a�򠜹�[��^�;�U���O�_I����?�}�kA{�;��\�7E���u��hɹ�ߖ�ɉ���|D�[v���{1ڈŹs꧶
��'��^��v��@r��F@W{[�R�#�qp�䡾4�y���B[�/��eF��q%C���7��Q�t�o]����B又��0�3OLaw�raY���;(d�\�u���'�mc�?���?YlQ=ż �<���,4��K�Ǔ1�Ԧ)�c@>ɐ������̆���o4��3_�2��XlxVHYEB     400     1c0��$z����ϕ��0{�wC�=����X�D�[Q�b#���2Nsѳ�!"�J�#$�u�s;ɨ�C�� Œ�Z��=_>H�v،Ӣx�*5ˎ�м(�wk(����b�olY�a�MA!�JY`Š�<1o��]7���JR*�۶ߒ*��i�,�[��۲���}D2�R�[�_ppe�T6���ȼ����\;�d�� ���t闔�L ^vp��T��H��C��6��\����%����4:W��5��n���"�o��WOt�\y����7E)����L�9IW�Qn�i��~hQY����*���0O����G$XՈz�6<N�f-�Tz��Ň��G����d��
�v�n)�j�@�{���V��
U"�eYr�~�Ȟ<���/��E��7�`��쐵��P>�`j�b�$|I�gn &��s�[�7�j�n�&_&��ӠXlxVHYEB     400     180�� ^SINZ�^�Q�X�b��Gq���HtbP��M��E�K���qwH����E��d�%�pl=1�j����4r%��ㄖs�B�%��De~�˞���9.���,׍mǣ��Hj�	�I�4˪fh��=����:Vc��\�xa�#ߣ}8�9�u�m��*�w��K��85o\�����ڍ��\◚�1��V�#Ā��zL�ӄ�鍣��WNJ�>U�%5JM�yŘ���ѕ�B<��Z^�&<�r�y���4ܜ�R��TQu�+�6�#F��{J�.m��ח�[�-�,z�������l����I����ڽ�ߥ��c�H�jGV�^T�<�3+o�n�d�T>��P$Ǟ�r�E؉���p��7��1*�g��4�̲�XlxVHYEB     400     1500g�:�&��B���9R�	����V����0�;I峅�D� Ă��i&;/��'QDZ�����^�k`��?w �/�|�4�'�h=��-�O�$��sN���K��T��H�S�G	^EdS��p'�SR��QsD�� Z>)�XBt��h
n���G
Sl�*��2�8˲��!��DQ�d�����:��A�%�o�[�y"��~_k������&�f�s&|V.�H��O�)��T�W�'o��͒���j���0�K���D�BڞC]�����L}!B⩵�O�[����[;�sT�c��O���6�Ɔ�1 @36�n\ᳪ�y�XlxVHYEB     400     1b0�
��D�B�i!#Fɲ�:�{(�ƶ�%$_-�ɝ�x����ٽ�6 �r�3�0��;嚐hd�1(L�?�1*�>�e�Q��Q{��#*���}�E�m��f�0�M���ʝ1)/�VQKt����kGMي4p}�H|b����J�ZZ�N������O�<���B������-󂜑� �6�1���[��Ya9�T�y�,g�3u���^b�m�9� ��ܽG"�G��h?Ε�5$)�?x��(��:�mI0������m�`i6Us��p0��V7hX�����	�߱��[x�(��j3�?i,Ka�|��9=J}���IE�+Ɨ{M�'���¯��f�fJ�t ���4���=un3f�"6��N���Di�r�)8g聏��le�8I��؍QBmVېGB�KD�=B#��b`�XlxVHYEB     400     100="�^CbU8J"���PvGW�-����l����ַƯ�BG� ���7r9ϥe�Y���P�0^���ԓy�X"�f�U9�j�&�7�4��Me%WuL@µ�nQX;�#�Cq�C�<5�>�;��c��1T�ȽUI�A�s]/^9��,�)����5�b���;Ų����9^�����p7"��6���%���Ҕ�.Џ٨�ب�u%b8��	�N�e�*�	�|����/���})���kl�ɹ
��HoXlxVHYEB     400     1202���)�G��O~��	���4ߧ@�{}N(>�4:�.�^�g)�S���	�� $��E�B����
z�A��K�i�wL�%��[r;8�����Q�S��xV��!���<��ǲ��X���;��+W�ٵv2�yw��G�������sD�u�\�$�b�-�FS���q�����|�|6��`��#�
v˒u���o���߈�t0���H��y�"O�� ^,jΈ�Ezj�1//Y�����D����Н���4XIIc3ad�w��1ߏ�ƍ��˯��)���q�-u�6Y%7���XlxVHYEB     400     160�U5�4�A@}q]>���A�0�Ŷk�|������r	�P�� �׿N�]�n�gx>���1�윙>n��+�J`G'ǒ�
�������9�%ǔ�8h�*"M����F��?%O�'y���JA}rȐ�t�y���q��9�2�)�� �RPo�"!����n1��ܔ��?�}6���7�#�Yͨ��s�:ؘ�b� ��0�R�A���Dx�4ޫ��$�B����T"5m�jbc2��t�Q��)YŢ>�9� ���G�΂E����?[��Eqè���uؼ5o+����%�Ø��%2w�G�^�幖?�n*�Fj�R&+nMD�Id�z.Z���}�.�q�H�傗�XlxVHYEB     400     110��k�rt�3G���z��N�&�k:~�Ή^�}mW=I��k������uRkr(���)'���{V�鼙�0���-�L�������/�DZ�;I�����Y��=Q��B�&]��%ݨ��_=�ch������0�ȷ��d=0H��w��6����%
���?�׺�]{����� ^�U4��c1<��P�O@�=�%��� @� ����=J�@�\�]�vU��������%zl�J��a��R����?�c����Q���3w��R�qXlxVHYEB     400     100���	\8TF�XO]���6d>��U���/���[0�J٧�͜��aߴ�>y(߆y��2�{%Ԍ�e����G��ArY?��a�kb
����G:�3�������� o�3�N�O7���F�ZyE��-��D<z�~q�oeXv�E��9%a�����n_K�!n~���4�����W+�q��~����k	�@���B+3��j�dm��y��I�����T�²�������;��S<��rm'����l6XlxVHYEB     400      d0��Ҟ�9��?�M��-��MtᕼC[���țP�]@2-+�.ۛ�$����6�G5[wkcL���ycڵ���}��0I�K�t`�ȘQY>~�ff��2��]ĿY���E֤	R��V�D�#�<İd��ה �.� ��(O�+ u�����`���%aW��օ4搿�\9
��B�u�;`o����~Zq�����`��͹��5WXlxVHYEB     400      d0f��C��� Qc�Ȱ����X�zgTe��ac�&����"|�2g��7e��˵�ު�Z��ɫ
��ryɅ�ֲ��k����F�,HRZ���lW�?c�B0��+И;HC��ڣ(˨�6��"(����XF�����Q�����䲑�R�fjy�z.v��n�BR�����,��d|�c��h�\�#�<�c:�
��'6Y� �
��)�vXlxVHYEB     400     130"�l���{!�� ���\�re:�*��U��3'�[a�˄o��<Q?���ܾ�p<	�\���x��@��@r��ں(�'��c-�@[#{ -��[\ Z�br�]�â�/5��9%+
_�:>��qgC�K0 
{le�.�'y3bh����A\/�Jɡ�˒
4h���9�b�B�͈��)�S_��Ng6��������۟)�鏴����$�$Do����\���RN�J�W�
��P��pn�R�N%�@�=L���rza�b�Z��Q��[%�̶��k�6�J�5�Oā��$^�@XlxVHYEB     400     150
.��bـ<���\#O�D�1�t�n���E��!��?�K�d�@�ms�,P_�_�j`$9����bB�#����M�D� �)�Y�9��u��{%������6�β�h��6ma�_�f�pH�톧bu�p�r6�g���a)P[�Θ+v�mK�l�qu��󢳁��dNFN]�W��+�!rf�u��GK%*L�71b�&����'�/�p�'��w���aF��j�Y���_��qg˱_�����Z�f�@`-U7dH��;�LM)�~��γ��Ba�r���L�V�l��ЃTZFB�~�������v{4�>�)G�aD��<�XlxVHYEB     400     170����WVԮ��S)�s����IL;�;��h�x�V��t[���Vû%7��x>oj�$�MB�ͫ&]����_��O�����S�쑄�K�o��n�j��.4������N�hyЖ8�9��V��7��$���v�r���LgT����YF�-?���'ߢ�Jg0��w�=N�V����I��]����1��y�,��:Os�g�f�](�|1��N�g�����?���9+�;��
��Q�& s�|�� 4q�N+T�,~���r�/�]���r��S6�;<ѿ��b�R�oҦy�B��F��=<�6W��^�9[U��P�\K,��-7�g;�4����;�xq-��麛�� B� -�i�9�����XlxVHYEB     400     190p�hK�+�as�l0�2�(K�?x���||H���-��`|&�H������
L�78�(��y�Y����7���;�7Zx��"Р����h��Z!O�;!f��.q���%k���*W�K�A�S��9��m�����[���O�vŨ	yu�J_pc{��E	�I&Ϳ�wr���v_i��bջJ�)iy�A�(8-O\����n
��17��\Z⍿^�<�Y~��>�g�՚k��ñ�#0�4>7yg�f��p=ku����FQIY2�$�rM�~��U3=O�D�`G��x��C��G8��v�%Ͳ�GJ��N(r�?�y��=\b ���pP�+��z^[��T� \_H��7p]�F���x�f�	��R���!��wl� Լ+XlxVHYEB     400     180��y0���m#��� ��VQ���bjR=���w��I�mZ��f@d�cT�]d����������e���<�<E�m���i�5�M���&G������R�(�	�<6s�l�L�������"�i# ��Ð
o��8m�D{�Q��Yzƥ>�=�:AT�)��J�xֱŨ.N;H���Z*����LC\Z��ڴu�X���}Y�:[��ېջh���)�8)%ʵ�lt�n״/�ѽ����?���Tn6il}���P3��Bpr�`�����YA�x��[��sOe�M��4��/0�AQ&S���I�"�~�``�%���֔�E~�`��n��+e��r����a	wyǋY�Nس���U�lI���2�b��
�wXlxVHYEB     400     140)��%�9�ɖ����\�$�{�Dsf0�`�#�H�����0�� �c�.z��@��������]ɫ���c����ᅡ��J�t����$���"n��C��i��ї�,���8���9�?��Q�t��uFtgeo�����)�Q�m�>�%G�I���5�bKxim��h��?��E&�+�2���B���䆔SZ����)cy�Y��U�I~h���`������o�h�gL�14l�j(F��3-���6Q��7ҹ!o��\@�Pt!Q�J��'�#L�,eA����Lqi֢R%߲��.Tp�p��XlxVHYEB     400     130��oj�j:4^^��j��y{4i:���G�C�cյ�U%*>�p\�ki�:������₵'����e|"\�����_2\a�VЪT�Q��EbZ��}�	eU�d�@'�D-�8K8���5����ۖ8��9q���rUd�v(_X���׋4�����#[L��7s�b��q�d*����a�����g��|�@�@�]���ᘘl�]8����#�9R��;�O��'�b����5��؞%~���TW0�[��_�f��v����l8��m��j����VM�Q-�f�q�Z�:���iwXlxVHYEB     400     170ϊF_���eI�)��+e�gq��3-E�Ԍ����y%2.�;Ft�=h���J�>H.���hF��m��t�=�_�1M��V����!�������$S�[��q��Z������V�+FX��
V�?"�4�tS[Ÿ�q�iM�z,F�k]�&�)���o&p�U��#9KN��	��Fٿ<b��,�9p�S�C@��S�̓M�̟G!-�V��B'Q|ё�6��V��;:W�``��嗓�Z"}����<Y�#�(�?Wh����.��կ�VA������\��w��ŧ祾��b�6�\��}6�r��ǟ8d<�8�eB<�UB�zS?e£�U�̐�_��1���}H�8�w��6]N�N�=B��dXlxVHYEB     400     120ʀ����Ш��#�OQ�e6��������xI+iM^	�r��������}L�fY���Ю��@�Ӽ"8>�7�z�7�^���G�E:[8��)��(N�'���)#�|#��aF�sS;�i9�#'�Cwh��v�Ms��a"-R�}()f��ck����tEl�C�g��Ds���&+��X�ʕD��u��eJ#bgd_���GF�M�k{���&���GN�";.pI��'�潊�H=��ݽ�1HЕ��w�L�N�Wu�ٱ:�����Q^��Ýi�MUXlxVHYEB     400     130��BxT~%�*g�����K�Ȥ��j��։5�a+B�j���vټ���'�^�W����ۻ1J%����iJ)�l�}#"�5P>N���7���"�}3�EB����W�g�"[��EO�������(�nO���1ө�y��?	�B*�:�-��Q9$3�9� �GΖB�'���f� O[6%���zK�%/:�XC|�؇ͬc%�F ����E�*���Ha�j9 �<�]?!���U�72)U���k���a|������~&7>4�٬�C�`4�_�q�϶lAd�]��ߗ�qu��Z>�XlxVHYEB     400     1403��+;8K��g�b�L��������O�4۲t���G�l\�vk]�/􈆆���G���
mv>��V�%�lE&d8�8���[
F�Y�-�v�d�8Y_�0���\�b�#��Y����p�zٌ�SYp���aZ��;`����w���σ�TF�������{z�u@�p�C+>1���:�evP�{�H$��"G*I�B��1�D������x�
�7��1í>�vjx���%;_EE�x�Q Υ�?X�Xv4PK�����n�����~�Y�r�(���D���\��L�H�H�~��W���� rwXlxVHYEB     400     1a0��&G�7�fvݩ
�I�{��!1�
v������̉B�n�вQv�g�zT�GV7��6��8��fD��\I\���F2hV����i�[���c//�rT`E���^p�YIˣgv;L���4@8�u��7/�sm�)a�8H�/94�^�G<y%#Myy{v�A�s�dS�]�*�0�7�Zg����O�Iht�'�ak�on�uY�s�S��9���l�	c�kheV`|K�Ex�7�gY�*�6�)QĒk��"����a'ed_]9��?��jj
����XV8�g����������C���B�ٳ1�7���g:>(����V�1�/���������Rz��rX г�-��r��& l���5���,�d ����b�x]R��B����瑪�VE��<	Pd�0��NXlxVHYEB     400     180Qz�&��{"�(�����y�#ӍKu$�7ߏ>����#l��6#�a���M\R_�~XA�*ኋ�d�ބ_6����b�����\����U͎���A�>�n�l���ř����y�u�:d
���\\pf��}�AJ0�ca}$���p�w/�;W��S)�tu4��K|����$S	��4�"�ݤ:��+g�H�p������y��/E7��	Ud�w�e@�!�fU6_[	�m�C�ȗ��������{`$���,a=fQ�"&9�'?�#��k/�J3;�e�`O)#9��G)-p��E�|V����@.��e��ނhI�d�:�H�FwA�q��a=��y�/$\�7�!�3�s�����L1ެצ����~�W?C?�XlxVHYEB     400     1707��?.��Tf�m&���'oݽ�Dj�A�V�I�E����)�AF~�Nw���#O�9�3��a�sN�W���jI⏿"���X����sϖ���e�+dwx�-�}h�?�l"@b��qG5m��c��-\>�1V��M�J����-�_f;���{��s�s��9�����_����a�{�&�.��v�j�ũ�	OC��g>]�d\�j��,��1��������d@*^��C�P3����ck+�1�e؃�S�&�Y-�lF��9�i���#T�_�X��h`/gꜣJ�.Q�P���|�E������3��b����^�U�X�}Yc�~�w��*O��7�P ���eW8��	��T庋L���XlxVHYEB     400     1e0[���'�ׄ�U�QJ.������Ƕ��:2CbsY@�Nj81�'T`eh�l5Lf��OD�}t������3�&�����o	?�]��s���tE�.��4`�p�V��ЛE�^����m�#ZK=b�`Bٮ�5�ec2=�{��M�tb���1�n\����X _4 ��w����'bO9xۍe�y�F���P(��y1{�u���"w�������lb�Ц~�&ie�Y��9O#�e���g;Mڻ*�'�3���D���S�F�f��;|����&xG����ީ���cx��IC��1�Y�.�5�?�	��sh�>3�ȭG��9�)��M��˷_\�/��|�A��{��9��y�`ؽ]�U5��obU
j�S�4��#�]J|��bR�Ո�S܃���i���11�}�O	1�n��Z�m	��I��x�AW��7�ss���� �/���hG��\�e�O�W����#%���q=�	����XlxVHYEB     400     1b0�r����l�Z�M��n�E��l�AŐ��b}�-c���3,��=�1f��6�֭}�z?�r�Il���Ó�"�@�!������������Q�"����Fq���k�4�G_WA�J)NW�-�[|Ӻ廥J��er���Q�a�>�9����g1��u�;�cx�N��I^��b�QY�Ľ�_�A?g��}�s�Rk:�˨Q猻E�*����C�l��� VX�_7JN��|Q�b_؏R{��Y��>bb�J�`h�UP���DMn��}�?G�6*��njh�
��24�x�_���-�$v/�W���!}7�jg ���De*�_�[G��g�-ES�G_$6�; �� ����94}'������[$nO�K��Z�2ͬ>���`�7؍���Y�L�ef���e'�bB0SQ�g�R�N�d����Z�ݾ7�XlxVHYEB     400     160x�	]����=��_Pag���ϭ�l'�w����"xӕ�4�S�&���ƽj�r�ç�?�(�C����X��y����WAh���~"�� �Dlѕ*�V��t�(�i������O0�\T|�J�3���Q�*3%�ɺ��ѹ�Ʃ�H�7�:X�;gy��P>VE&r��Kt���^�߀�0� Jo�x�/js�w�E�hq��m;�3�h�Y�O�Z[p�"��F�axHO���4tm+�sW�w�q|#Rqo�Y��ɲ�H:�÷L2�FmxJtr�0��&IXu�އA��Me�"���/�#׾s����=1GE��ٽ�~H��Seb8��λ��w�:pE�XlxVHYEB     400     150r�W�-��;�]sڤ���1�J�����n�Fv�/������>���.���zj�dю���6�T��ʟ�9!��Mv��껄�P�k ���B�aUf���om�.��1>�����*�sa���a!�I��1����`WcD\������\���ty�d�QfG�$E�A搰�˽J�95��s�3�~�2n��Y���% t}����Smq�%)�}�es$�����ڜ�o��)�����a�����I�(��F���(�9�X3�� qX��RF$Z3�@����Q��1�H����/�⣊�ԝ�{an���%XlxVHYEB     400     1a0��X�)���^�!����8�i^tĖ�`þ^Rȵ�@?����Y�|�:~VT�y�ƿ��O�J�nH-�b�D�$������AH��;� ���P���?���9(�? ���x�y^e
սY�ZY����/#�k'��@�1U���<=�$�u���O�+��[.��*g�z��R�H��EF@�W_�wq-}�u�(ty˒�)?�~"� ���+����������&\�@�����wp�8�D�/�\�����9�e�`�D>�.łIt� 8���)nd]�H�3��*ysF�����3���I̎�FSj��Fa ȶ�reebjg��3��6h�s�/�ۡ�\a�fp��I��g�K�X�N�0�ǔDBĄ|��NA�,�mډ"��$IS�\]h�Up���XlxVHYEB     400     150�\�{�"B�[v\ 9�{:� �a�xוSmhz5]�PON�:g��̮�NY�<����C2�+�]̕JT��{ʹ9�+�y���5�$1�@bE�j�_;���o�G���=R9�\~�Xxۤ�(<6��䷩㚾t����N�Z�\�L�#}�LC���� �pnCd�D.פ���x��Zu¦���`ۜ�b�@�V�._	�ր)O���b�bzu�@O���#��r��F������:	pTc��0k��Ȥ��o�X'�y15}�Q�p�A�@q�lAa��A���պ �EMA!�o ���Ů�m����o�L�\@H�l+ :M��� XlxVHYEB     400      e0pH�y$21��,��)��?=���,�gf��r޽���A���?�::>lg�8�M��#h�a �� ؛ 6�����,�P�-�I3E��>o�ũ���)y�C�m�	��������A�q�E� RMW���8�8�OUoI&�����\$ �l~G��HI2U�*�(ԮPi�b�h�����4*���ˀ�j��OFs�;E��ɋwד3�LV�}�[��h��iXXlxVHYEB     400      e0vC�m����g)	��zY�%���Jm��&P;.P�T��ψ��Z;�g�g�n��e9��j�b�25Le��%$V�Z;������;>�f�����~9Y�׸��L'�9�pBB1
P<9�'B�Ѿ D�7�8��Fz��'�Ho�Ջ���W���;��'�j��I��5NӜ0������Z^���{~N�Z�,k ��SP��y�;xU�ַ;Ő@w%��w�9XlxVHYEB     400      f0�����q�'fB=X+rZL^�Lp����z!0`k���4	Cc������V{��1�r��ۺ�.�  %pK����Us��nP9��g��zF��;Bo��s��÷�<ߠU�Wa$�yj�4Ai�q��T]?AP��y�.���sF0�]�U�����uV�(�8��ȱeձ�r^�"�1��,A�������h_�%uL��.ӓ�C���5�D����źQ�Ͼ�̤ �ڤ@����XlxVHYEB     400      f01iN��ӹ� (�^�*w�L��������!h����㪎G����XT��,��$I\��T���5��Í�L�1�>��Y*���w��ь�}��>.�M:���fB\;��1�]�
F��CPr�l-�(,��Z��YE���;k·,fLœ�ֳ�Z|��[&�TH�����sL�Q��҆�(�O�0f7F�'�6Xi����(ڛ��O��j���.��(��ؑX4S�D҅�A�n��#XlxVHYEB     400     110�J2�U�ND��'�>]��"�P&�A�ZnG�,�r���<�Iրб_T<�2`�:m��	8��ms�T���zn��j�� _�J��1O4�s9�d֍� �ʢ�C݋�[����(����˲���@i+j <[��*\��O[�UFx�B��^>���DN�1C��2�l9o��>W.��T��h"�G\k��,��������$�Sd������:M�^#?�;:m��#C*{d�� ��&�R.qkK]tf��ȈcIr�����@aq�`#mXlxVHYEB     400     1b0�fBW�Ng�9�����U:�3�ҍ�J�|�����y0
�ݝ��?������a�f�H�m$�)��9��]-[�m���"��S�K�o�)�\�D�������7(�
2�p�P��~  TqM�Cq^�KX��eJ��BSkk\l9����gѺ�"q"�$Fo��2@zl��Q�8����<9X���%p�2�2��m�(/x�������q��!�<��T�6v�qeb���+a�7�B�)�|!���E�Rh�2�V����'��y�R=�6��@���fQ�1C�`�O#��{�r���[ؼM6�Q1��	al�n{a6�^|���=��aUט#_D����z��\��.�eJ~HԎ��` !���Ē\b�`��¸��q��끳At
i�_�X����/̯e�� y�=��׬ ��XlxVHYEB     400     140�� �����D� W�����I�E2c	�M��A���?�����o�����%�Lk{`$B���N�JD#�ϩ#���YĆ��X5A�~f����QJy��R���>����,o����"A���3�E*�'�ַ[���[D,��TZ(D�y�Yb�o�Z��Mw�3式y�i�k@(F�+�
�}.��$˫H�VHB&4�U���>�/Y�9Z��� �G�}QP�d���' �8d���Ӡ��R�c�E�Gi\YG��.�k	��f��[dH%tɄ���>�5q�m�{*Gi�+-iL1%lpr�ZP���1�"�(�XlxVHYEB     400     160٥���)ԖŰ�`6���)�ԧ/����8�F���OK�
��*ś�"qe�����Nm�L��������d��4C����D��+�J��ꔀ\�����B��hx�ϸ���l�v��F���0օ�H޲�T�'#��d�U���b>!�Vg������x���2Ncs���k��[��F�3�B�@�a��N�������׼[��������|�Ƽ�j+�[)��ͬ�������2���#f+��A=��W������u����.�[�F<~�G6��LŏK�zOS�+��������,��.YTp�yL�]��N@z�m�y-��Ŵ����?fӍ��@@�"�k]4-XlxVHYEB     400     140�ɥ����wHudN�Ήi�͗�}!�C����5��� Xف�A���w��F���k8�cG)=�ڜQ���B��`�����/P���=���	 ��2�җW�Ӡ;�l�C�H(pЦ��ɠ\%�\4�t�+.��<��ss�׌��\!~A���-�	��=�hES"�6���`	��3\�f0O
z�;���ߟ���@�?ۅ
,9�R.�i9W_O�-�|��7�sS�w~a.�I���l��?�N�!��J�4y����;���#Z��Qu�r��{.�jI�H� ��j q�Vu)��M굇�Fs�/M�E���n��!�1Z#XlxVHYEB     400     180�bJ�Qg`�ׂ>'}��������e\���X�ۀG��_M��<g9{i���k»�oת��o��h�fv/]��<>��V�l�M^��NNo�[ha�������8����˅/�v9t\�N�~n6��e��M�V>����rR�e޾���V�;����^�(����4����A��QV�%"ϖ�Ω~�3}�xO�5��.�3��� ����I/��KuR��ɋ]b���GK��ʫp�}1�#$�O�d���F��݉<3���-"�R�|z����ku���XʏO��!@W����p6{��`^b��^n>'��Ν9C`�@�'��Y�\�p���I|�&��(�o�x&e�^���gOTs�M.n�XlxVHYEB     400     190�~���.���[�����C_W�et�Ԟ��٤mcʼ��dh<v6�hV{��7c5�d�(���s���k�h�Qy�9)���q���6�̀Mj�Rae�ׂ�?�/Ag�/?����I0H�u��n�@��;�]�i�L�-��/".�����u��>��t��b����g#��jL۱JJ��\a���0>HerÌtM-F����3���8����Q��#�������޹�6�R�=����hF~�E��qk�����p���^Ecu6#�.	r�R�z�0Ĳ�ߟX/ J�n�tu���lD&rP�}�|�B]ϼȰ�&�Y!�d�8a�O'k��=�lH�Ύ}ϜY�ٽ����YBH��z���Rw�����>�c����i'��b�/��V��d�)w�'XlxVHYEB     400     150�ʠ0J�>x�ʇ��L�0�H��s�Hu�j�W�?nJ0ȾEL5;��1E��cc�����>+��c��0�4�M����QAr@ ̘�?󒬢�y�-��״���Ɏ0�
���'4���)X0�Ot5d�/F����a!��Ve/���I{�,ny�$�U�oG����?(YNWZ`�c!��]KX�}N�������(�,�>=a����ƣr0,`4�{.,8�2 �h�JDސ�3�z�#�:�!����F�"rM.F��{������~���%��~}�Z

�N�|8�vD�c:���v��(:���-�D,ϡ��:��U��MMDK~m	`��SXlxVHYEB     400     1a0�{�y�e2���=PO���P���{�E+9��y��E�ս�O9�?E�P��aA�x;��a� ��~�e�n"r�gB�l:uG�򃜢x
�\�mB�v��On�+9��&�Й�n��b�板�m�{���+U���tu"-3��6�\S�н>Z�s]@F���&��!��W�e6T��/���H��A����T�N*0�K����Un����&R:�ȟKo�8(��c���9;ěB�ְ��bEq�������w�o�9��ȫ�"q�<�Uz��b��~�����~��Ӝ$1*S���1pC�h�r�+D'��^����+���K)Z���\jG�J�	7N�WPR�!(0���࢙3}�^������%͒�R�����'�3��5&�/z͈&D�PG:]�f�P<<Y�@^c����],XlxVHYEB     400      f0�����WLs?[��E�� M������Z�������*��dva�y[�.�ڄ��c�wԅ�vKi�:�6���=��LE���r��,��{tS��1�ac@����Q���ǔA���w��Y�� $�����e,i��]$����_����N�
�r�&����x�� ��f:�� ��y]R�b�;ݟ
	یu��zt
�������v�}��O�Yr2��)w9X'?����*)���fXlxVHYEB     400     100����*�[���f\ؾ�b���228â�lϟ�S;N5�r�=s"�L.��:u�*�0���$�eU����{����鯨�NW�q�^���!���X^�;���_Zwk����c���"p�`���@7ۗˊ�g����ۦ��}�29��o�F]'e��Q�3� �? ~������h%vl�&{�6s����I�JAͰ���ζ�|��p��Y\+� 1�11�W{��Y�Ms��d/�^��� 0��XlxVHYEB     400      f0�n<k����PYe�Qp̦&ԩ����9�:��%����J�_0�e?��eql~�mp�h��B3�F��������5d�Q����Qb�S �'띦G
6���J0�ӂj��v8&c���O��� ��gd5u�.�>�nꚱ�5QuCHN�n}Cv~����{�<�cv��ܺ.=Ƅ�-�s].�1����b��%͟:��~�ŵ�۫�F6J6��Re#�1��4���G���XlxVHYEB     400     120���'huq�G��;����@ķ;��7Q#0�̥�kn�}����'~��̊8k���d�%���K���sf}k�O��Lo��i�tjH�R��5sd`G�&$&Ё�wd#@����Gb��5�y��q�`r#bڙ\�䦾�6�bdSP�}<����
4"�1U���r���p�)�1�.-�����O�����s�yFh��5��ȉ��� �ɬkƂȫ%QK�R�К��6	Z9*>���� �J�X̦���S����8�ɯ����Ot�h�\�4j�.QMXlxVHYEB     400      c0�6V�*6�����D�e��p��8>��ʒ	�m��RD;0]9���&s8���{���R���H$,���!�㕻d��}]�X�5C���H��~p�1�'�o�U�:Tv��m�b&R���S�To��;�{����/�P�Իӄ㟟�M1�����	D�S��b݅�4��KN ]Aݞ+���A�eݡG)�N�XlxVHYEB     400     150��ZWG�U����"������"lz���D���$z��/P^SD�Л"d�N�UY��a�\L�醻�}��j�=�����t�ۨrk��IM��J'zT's�zO�f�%����p�2&(7��$m4���<1�6��"��j���F��5�;�x%����C��ޮ]������>�4?�,�u*�`��5�X��9"3���T��4��=������Eܔ�I�Km+���S�#����'�d\C����Ku���m"Gݡ	Cѣ���rJ��I�6���b�ґV�;�c!��>6Ҭ��@�:#�-aI��Zڦ������8h{ҎѮ4��C��XlxVHYEB     400     130[䉥/S���#�����X"bToh^Pj�k���4�r�HH�����Ǎ|��Fc�\,KRȗ3S��)f#�fc��8ذ��itU�� H���#�ŕ9:35?��,(���� S҅�#��D���Z�1q� ��d�D��݄Ŋ �����t��]�=/���p9�&�,�g0�(L|
�����!����4����ʽ#�C )��s��"ϴz�vi���e^]�E%�9
$1L�P�So��.,W��|����븁OɛD?�S�M��i�>�?��n�_������5kMsgXlxVHYEB     353     160�OQb���.��z�����D_�u �^p��%RƀZ?L�f|�%�,��X1Ic7gK �to�5���B���h��հRnI����;l>��c��ʁ�k�L�`U�o����26&t�Y%������4��8n<�J6���U�o���'9�E<�=֗1(�>�QC0s����]�i�Zj���Y��<'�K�o�BI|i�`��lC��[��"��	�j�y�Lݎ;��t��sR-y12���92lm/@��w�K�T�0�̧����x����e�ާ�e����fo���<~
^�̂J3T�n��?�0��v�"nER���k�m�OG���~47L�(�_N� �*��\a?�"���j��