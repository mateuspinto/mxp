��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����$B'���1�5�i������~�S�$�L%TE�Z%ց�i;��	9�Wc�=jg�"��>��8J��
���HV��,^E��TlR`:ck���/����~LE.��#/o�'�����H+�iѸ�H���V(���,ͤh	尞d3�o��9yɕ�Č\t�o��ߴ�\¶�$(v��2�>Y勻�Al��&��}�r�~}��sq�1�9��a�B���1�K�0�2/��u�ͬɱ��s���l�����`��7'�9'd��H����͋9v�J�g�_�ZK�4�D��%���5���9�՚^E<�'tFV�� �7��o)�LV.�R�3X_�s�*�X5jz^Bٕ��ɩ��4SȪ�D�m⡌�q��"TP#���s�s��g�q��k�h��Rh2e��	JFĸ�ވ��<'2uH.��?4vE�Dz�S�5�h�������P��Uܠmb��9����ڋ��R~9�[۷�_HP�l�bw�!��	1�F���_%����zE�W��s�O��
��;8�י��H�!�XB�H��bŊ�Z��r���h��@����e�@2�ߙ:�?r��	����`p^�5��֟��)��C����8b�Lk��
jsso�+z�����>��7�;���ѻ�G�!A���B��]�}�Ћo_��E��gՃ]���[\x��=�0��}�V���w��ʥ�1�Ҍ���/dC���"�a^��:��61a��N�@@@��2��a*;�H�W�(t�����ʴ\m%(&oL��_��o2�=_����:�?��@�{'���#�Vg�������)6�D19�~l^L�Y���EKn��p��9�H�4�!=�A�*�D.��;"5�#�B����p ��>%���C�	��Y��@��
�{hD,�]'���[��Q�Ҟ�q�n����%ai��r����a�W'��ʶo��'����	���0N�S���\c�W�&�:��M�>_��������MXN��n9��l( �U�h �F�wx�5h�,�N��@�0G[Ĺf�qM�QJ�99�'�|啞�����e�骖�\�y� ��b;��)A,�N��Ϙ�g��Q蝰�)��n��"`�8&�������hu����I~�6h�%F��2�����/����e�}H�ҋYE���O�?\tp�{�wW<�'J���@��aR��yO$LY��������S���j�M+�����o�1��<�`����=7�F��`�<r�g���2�J��u%��A�*]��U�1�f�|]ZB��e�@��Z����A�E^�����!9��D�~𦼬�����P.242����lgj'Jdo$+���.�rqm������#㜠/H��jS�q�pFV����m�ӳK
���C[nJ����l�FЪ[�|
�kR@KA��Ǯ�f4�F�H�?���]Y�Ҡ;��}(g�>kCjM��)������s=sMj��Blu`,��%
d7��͜U�M:/k���F\^!�|�h�4�c+����D�E�muW��P����X�6m^"4���l[�;�zC׺5婭1�S#}�F�f������SP�I��;�R�"Y{W�|;��=*u�瀻#Eg*�O�R�t��N���%(�FMi�;�z1�?4%M�����~ֵ[�"�i&7�Q,��Ng��j�t��.i!�"��;���m.tg���|U�&�ȗ��oFu�դ,���r$�J�����m�L�=9=aOS�8B��V�g���@f�S�-7H���Dt^�S�$;c��<lI�ڌ�N��d��c��W���㿤>v��	#���c�~]��T�;-g@�Bsa�d��&6��l��� ;?����!����<�SD�ن�(��%���M�~��c �6x���ŷ;L}�����F]ɫ�%����$�	SdM��0��u�tM�q���8dM�'젡E�|����P�J6v���IM�T�9�u�����|V����[ƪ��][C��)�w1�&tY�3����p��ީW}�047&xu��q%&��)�9�T�Kpc-�Z�`�~xx�vu���1�	�Kݼ%
v�^�����i����d���ۙ����8�8���6�@]ۭI��6�줎ᐃ"Ѯ�p%4�~�<��Ej1�c|�"�H��ˊ��A���Wz��	���{		_X�aZ��ru��`����CC�hr#��9�y�+Ԝ�h��w$�x��80��I�'q�V�&�b�~I2x�X��R�Z��]�4�iO��Zq��	�w��c{ޮ �DV�����W���(o�.�O�dX���F8�ߧi�dB ��\�d�ʲ��.��W0�w��y>��=�^�b���`�sp7�O�������Ԫ�X��D�]M$quG���ॣ�E@Ʉ�����6�"RH����?;�G��3�@��Pԭ�ܧ��� F8'�1IpK����uPկDT	�9#�T	�}D��|W��h��F[����7�|5[`e���s�{�<w��&7�$��!�Cu�-�>�f�r�:�Դ�����GHy�̀����!�U��z!���c�5��8�>�>PRC(�:8��~MBM#9���:έ� Y�(a3��A�)ŰMc������s� l@]�0���u�x�B�bp{��7C$�B3��@��t���bWMnI�۷YNSU\/�T��?�r�(fq�#_%����i��{F�)*r"�+����h�ߚ*lªq#�U�eX��v�l�u)jb�ji���D��ֺ8T��É�(5ArΕU�T7��'�� �E�G�!m;[h����	G��������/�L`vw���� �úo��:�/� '��d@|#�D�^����ϕ��˪�Z�M�}7^M�l8�gw�d	rQ^^�Wqz[�)�Y�r'����B��:C����da�~m����� Tu���L\��S�D�����pʨ&Q�d(F:�V1��t�s��՝�]/�-�	�z�n�F�97�r�/����D�0K�"3�l6���8%���~���Ȫm���Ad��Z��`C��Tyل\ז�U\��>��w��t�cM\�P#�x��9�Jq����.������(�k��j=�ݞ&��N_�+�G�hk\�����{8��o��=�x2���
�<R���E�(�Q ���R��L�ht~?&=�[�u��ʬQ<�*��A��� hO��B�[�W�8/�Xv^�Qم�'���:�pYTAt�n��2{�W��*�����q���j�����<���y���Ru�A~p܋8�	=�m�t]��̶D��<�T/@����{�*��3Ƅ���W���ֱ�0�^���=��>���!v~�k
�[&�#�&|? �j�6�>]ZX�o)�W��[��5��z��F�{	�|��L�G߸��Zq=q���[�T	l���O���3)���m:���v�
���N[Č�ł�H�ڃ�<���Ѡ�:z��^F^���X>�'1���