��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���6��=&!��EK��`������H	�ʍ��^��-���<:��L�7炙-g"� @ג�3�CS�
��Y�g*��Mo0��#δ5��:cpPu��L�c2��� j5Ӻ*� h����~����-YS����R����. QC������l0+F1��pL4U�(����� 6;�a���?�3HI�%͘d�$]'��G����"5�v1�f�ǻ��1����DT+��H�6��H4�`��^C�\��I:�"5���3����x���^=A189i�	�v�ޮ#0��e�;��C뀉ǚ�_��*���k�}����Ub[� 3��$`>A4�xH#YP:u3V8)�)^�#7B-9����Fs��>z�s�.��FT���;��H��+;�/3c+\�,�Ď|2,� |k�<�������qV�1�#���o	�y�cg6��� ���iWW����̛���<�,L��-�ZV�@F6�P}���ϔ7�g�rM&�Q~d���d�"'1x<$��^�4Ǯ���E�eG�,1B��R
i��V����)h��+y�h��޵�/�C���㦝�z0z�fO��U]|�p����f�F�_�T�0���A6+ˑ����ԗ<\A����o
�(�t�� d��G��p���1��� i�[�Vu�y�t�����P�epfk�ͬW̩����d�'�6���آ�5���aCy:�����r�FnS,�ds�d���xn����b�
����膡����.|�\�
���	%r���rX�yxQG�Ri&���@����3���� qw�e�w,�'���c��k�a&u\���?���z(ȫ�q
O���OC9�����'��*�#�u�����N�����������F�ƭN����J�� ����b�X�x(���� &� �E���$��?�7��ɵ<x�VL���ײ�M]z�_,j��ՠn�8��o�ϲr��Ec��*�T`�b^vx�������f� ���p��c��C�-T�ɺ��U
Y'#��_n|`��d?t�5������\��tT�_�2 ��W*�f���~���t��ϰv$�W�����
xß̞*Iwį�#T��o�ST���_��Z���yFQ"X��S���� �{^�C���=�H��Γ�.8x��}�5��v�V�O� �hd2R����[I�~�G䮲�]c��|ew�d���26�2#�67j�t���UNt
���bԪ����w
�@~����5�u���(!}w�V^��9�o<��^η�k���C��ֵ -��)��( m삨sK_Fl8�t���#�)C�X��Z�0(8��
{�U�
M�~��MBX�?Ԃ�Ǻ�㐮���s̖8jEI�b�Gz�&"Øi�z"��ÿ�?MY��C�K���",n���nS�%;T���+n�t�Ƣv+3��H.�g�
��ь+�#� c{{��m���Q�^�����	��R`ġdɂ^��Mr�Lwh�_�T�<�=b�v�V ;?����D�Bj�ϸN���2-@��M��f�)�+������%�]������+�/��ڥ��ms�p����cC��~�=���:_�=Sn��m�"���J�ƈ���S~�|�	L�4Az�HX��)2k�y%�ҏ����Ž֮����65C����aQ�]@!���ȅد���6�t�x���r�M���^o_v7Y�}�qtv[l%�~��\�h�n�EO�{���/��ӗՍ��s��d���jbJd<�-56hG�'�2�^�������P�[Ҝ�-���<{sʨe>�/{�8��օ�����>h�l�/�"��s�������w�ᥔ10����Ƈpf��o$ !}a@�!�^������%���n�?�9�1����T`�w@2[�j��@\��o���Q�����^����2��/�AѣZ%S�A�|v���?�']_2����!��G����U�k����^��Mh�(�U��g��>y������4���P���n"���$�_w+��)V���F�,�07�.:CKJ�s�q9�;G�*!�?�S�SK+���V#֏�hҨZZ�_��4"�Ѝ��n�"hrˬsRͨ�U;��s�%5�����g_.ohV�����REw��Տ�	�]U�9���cS>3�\ryL������L����+2Z��lK��s~?���k�ww�l�1Wqw�!K�������P^�W���SKV�Փ]��k�L�O��r�=�n����p�g��1vy�09�$xy��"X����e{!D3�E���b�7�.e�F_P�a�C��ųü��?���Rᒫ�!z�4�� G���̆�\��UQPrap{�L�g,����:c�;�g�m��\�Ѫ�~�=q�i�\V�1���$��5�1IS>�=Ǉ�Ƶ���遨R�^����Z]�Z�ɠ��ֿ&���r��o������z� �ڃ�/.��5�L��zu�%�g��;���S`o���������/S֢ȿ'���?p KC�� ��K�C�,	J1 q��ylC�0�9�;hj�ў�乬`���ʄ�5ʦ�!G���A���$ء�/��{���%���O��KC4�e.�[堝`n��"��^(����� `f\��{��E~Z<� S*�{8�e�Ϊcc{��������e$/�
�|�LH���nz���5��J�5z7B�ߝɈ�fN�t��@�L� �RK(�@��a
�G���y���k�^߆|��J��ĒK7ף��QyFK8+ؙ���o����?�`��Г:5�wVPtl���Q��I�*����4�$G�V�5�!e�j&6:��P��.�bLt���9�7qO6��g^���\oW��"��s�[�� �0�u�	���l/�#�����[����N�b���F�(v����(��A$�)�3�������4U�0'l�p��7�5�)��S0�rw��H��֠Ҵ�<�-#���e(Ag��܈��d�[3�K����ș��P�ޕ[�(}��� �i�J�T�I��8p��נ�����r��4X��?�+a���A^�T��匆a���Ue�l:)��Nf.�O{1�&�U��`�)a��ڠUA�������5K G\[6%�u��� �za��|��F1�̡q�MhЉu��*}��H�7x�^����xI4��z)W]D�����8&	�3o�f�G��>��'�5�çYխh�Z[,����F˚PA)6ݿ�x�����Mn��)��X�c�@㧾$×SO�˫�EVVWNBnnyfe���� a�!���ê� L��{�r��[ᙸ[u�Jh3��������%��vR�� p��v\ue_qs8r�;�}}u�w����ɻ�m8tp�k`ʹ��=�x�Ss4�������pЉ�������r�~u�+[���Ko�T�G1T��>J0��|�L�'��o|����o���,�O
i���\͒��ʵ��]�>!��䜥\��crnVQ>��m%fl_���b�3_)'���У"����a,4�L�h.�D~״<���J��v�hF��˺ܐ��<5��M�>����.88~��5rT\�zP�0Z�`x���#S`��ȭ����<g���ߡ{�̚�i<ޟ����U��Ƅ-u�F�҈�.�S�zr��
� R���B|�{q�� �~�XJn܅���C��B�<^s��7��*�{�xg�k/��Q{��2�X�^}��
�C����L�9��m[o�4S�+�%"���߾�Ir�P�;�Ⱥ���D	/��x���[|��?�h���]�{S��6���a�����$B߈��C�>�f>E�~^E�V����~��RE�C�H�P/���`����<�K#,�W �Y6�җꌾvI"������b2�+�_�	�((�Q��E>���u��xԫ��Pًl;��K����i�jш�L�)�(�fDJ��yS�C� Ry��[6w��U�?�|0A&s�i�����50��d�є��������+�aoH&��~2c K�9�/k��[���r-&r����w���~�;��� dS�Ď�N6�1R-�7�G�{"|vϤ*�_
nxV���"��\�_w�ן]�_���r��ظ��F����{L�O=��h!C*z�'�ͷ�������T��k�;}�U��)�Z,s������K�q��a=̠��=2�,�K�f|]�{�A�Lq�J^��糩>�q�.)^,҄�j� �,D��#��d�y��s�}�8ﬨx'�F��ë�UW��u�����ZJiw�xYQ�h7�Cd~��$��?���}B&�6� G�Q�Z,/Tc�9~���J�P���
j]�r��#4M��*��>���I�Iu� 9���W�ϑ�����-�2�(�`�7���
#�l?W����D�@��-���4������-"P��Y�9���~��C��L܊���&Ә��˴
�Z�B-��ۓ-�MV-�qϸ�����jN��7��B.�S�8ɍd�6�ڰɈ��z�_�S�v�W��&�^J|!�	a���#P�U��L�k����R� {�$i�u�P�9�4I�
B~lN��w"~8/�r����M~�mR��d�����J��}�����DfPQ�d+7�zꌐ�	���a#4���-����f`��jl����[  ƤSUi�b����X�-X
2��0����7��w���h������ R�R�Ux,o��O�6q���4�ZN��s��ɭKi�ɘ������e�Һt ptX��瞀�P2����A�}������!�`�@)#Jy4�߆� _qE�JVD�gҀC�_0y���Lq�|�5Zp[��l�JB�%�0��ih��y� * =e�J_ZC����)ڻ_݇�K�N��Ѻ��݃���w������S�8$�` 8���v/�[,*NQ��aǉ��_��bK��`��:���6���Z�0�����Y�"]8(W�(t
u��X�������.��me�1�t{�ˠ�'��x�eR�4�3��O��<q��%�}E?T�hB��Ǵu�<�5�1����d��lb���b��#��khCh�wt�!�%������Ku����UΖ�$��|e
ᦗ�_-�ͶC}���d[�sԈP�����:b��+&v#�m�:����n�1��U�:���g�K�u"}�^��^��P�/o��)�OӃ��.�:G����}���;"q���-�����m�z�D;/y7)�f4�S@�I҇�L��k�����`O5��-h��e�P`����}���9�������ߑ�[�6�-"N[))����3p��\)�Pm�z���Ҷ*�7,6�`�����T]xX�ײ7y�i@~qit�:��b�B���8.y���ѥ9��V��x]�rB� L�KfOuc�;:��]�{YAw�P��E!O�V~�b�:4P�y��q��f�J�wK�c����/ǩ��+nќ�-�UZ8`!9:5������#�;hE��h�y	�DAf��зe� _Q�-���lh�s�&��B�w��!��7h���@ ,�/;$�[$UL	s�X�6�S;�v�����ډ\k�r��6ʯ,��[S@\����P��q��?v���ˏ}�ύ�~ԁ �z�ڣ�x�p+W�m��OҤ��>?�Y�|�hZ� �0���#W�Ee̊��o�y^�ƈz�r�,3�^(���Sr��eq�\��С9��BUZlqt~�u���5Zi۽S�:<S�5uvŴn�,��0�ۺ)oLk5�s����of�v���>�0�����k��'k�����0�zio_��і�ePZ�>����l�oݠYd�_�7PLa0�w�޽��-%+<6>\10H�m�=5#�-�|��[x+g�k�8~�����ݴ1C�gT1,ы]>�r3������U+�&曐>�Z�V��Z������ꋛ*�� ����z�g�LyR�\p�i��[�P��K1G1vy����-.�=��H����fʇV�&R�{󕭏oĻΔ���p�}C�ٻ���A~�Upw�}|�Pѽy��	�L����FN���[�䃮޺3���\��[&��;T��εQ�a}�l�B=9��?q�q�PK�}�Z�:t#e΄U�}�\��۫]v���S��0����vck��e/����wxi\@�js0q�:��IdU^��PP��\�`a4�O��8�p����.C�$>���E$��+����Ž4�g������S|8.�\ISu�l��� �b�7�+��W�
Ume�ٞ_����S�)(,�i��#���M읝6\�8�u�e1�����E&�	�q�O�an�)���?O�b��j���N���Y����޸(���9?V�<Q�JBs?����se@{슩�L�K���S}�S#�!���mY�at}��V'B�U�|K�F���*p��-�\[�p@�E�Z4�r��t�}e��>������'���k�s�KlC`��dv��"ou��g��^(�h�_�8Kw] Kŷ�v�s�c���gL0�?�օزZ[f��O�S5���c�ut�/��1�f�9�`���3�]��ـ�*ɿ���>�-ST?�I.(f:���cޚ��2��G�k�;2�� ���}Ǽ�HF�g��ť� ����G��zT�u�h� |��x �}A�}�����+�m�"�~��{7�R�\�eCTM_�P�5�M�-PY�a;��l�73w�N��֩r��q���P�a���Nq�5�9l�Kz����5˭o�+���R�3���p�% A��EP��]���P����	D �"^�ssP#V�C� F[����;��ճJ8�p3~���}�v���(Y~}�3E~2$��p3�'ģ5zgv\�Ğ����O{[�5��Q�W�(���Ը6��6O%S#ޯ�w`�@���([ؚ�� @���o��hV�O���k���h���U5X"�/.��\����'��4��{sbEg�6m*��b<��r��t��ٮ�1w8}K�Q�Ϙ>���	G�f��%f����ك�����6�0��r��:�T���U���`��.$ؐ��΀N�H�v��S�w𣏕�� �΍��Ի��7LN��]��l��j��
��������h3z�G�Q� J�����䘾8�^�E�5?R��_�Xޠ-Z��DC'?F[i�����G��K8��O]g���>�#�[�{�8Щ(cr����Fr��e2��{1�N�9iŖP�w��1G&�c�|�� ����);�,\�3�������un�*���1���^6f=�)n�$M'g�}���Y-o�c�H��i���U�^,�Ԕ8�zx^?T~��%�mb�Z������?Ǒ�������,#(���`N�T��A�}g�W-��g���4W�p� �eT���%��ߢӴ�׭M9 �"�?`��m�9|�p��s`��nz�ջ���H���Y�^��.wQ�KET|`�9-N��q�ﾾ��D����S��/� <aś~���AS�k,uЍ@������A���%�@��9r-�PLW�@�UNC\��~����i��UΑj?5���F��e�Lo��3]�Ʒ`�h�weo��-`~��}ܢ�L�"�X@F�~f�}UE��������b$���LΦ��AOg�f�����D��/����b豊u�^8M����R����,�5��fN��:[3��AOֺq1�5���ڃ?*y���O�\b��#�|����H�̃�$�`M���	
J2�xi��۷���2g�e5z���*�Bst,�B��"EW�x�xޣ^Ä���'L��$���hT�s_����r�U}�R��k�řw��Y,�􊙲�%^���L��q����J(`�za�a6�}�
�f�_K��")�k���fE0j~ `����V�S�e�֖�����P�{x[�Gw�*��Sjpdk3O}�p����?0����Sq5Dk���D&���f���D���|9�k��s�G<����81(�|����%�Zȅ޳���
8�!����ȆQN�wV�'֒�A�8��M��۹J��x�̡�%��i����l�q����fd���r4�NӰYƄH`����%����Y�7}��g0����>��U-����?�����.�O��vR�����|��id9�`��
>W�]
�f��,/�����'�];J�� F��̪jr
#l���C`Zé��7��3�ВQB�=BM�E
�9�Vx�����ڴ�'/L������TFٿ+q\���+(�1�Y��(���yF��}&�Bê�4��V��E�M	%4Ql@yj�*�zY�̌.��m���Y�(�*�R����	w�H��3�4m	63�?�>^	�P>|�����>��-dR*��X��1�|J8��h�� MY
y~���GEp�+�����op	x�S�tD1fC�M�������
ͻ�^:��=�o��hHż��/Y`��A����7�&�Jpu�;�#�g��@;|��-~��*�s�t4�-�e9W�-��ý���?]P���$��ʞ���j�/���[Vu�9 �g؞c�#[W
^��8-��x�W�6�'2�@��d���ӡ�5pN,�"�N��$��_�M}��D��L�Wt]�e�����)\*�˟�� ,��&��a�:�����5��ޔ�݄�6�m����9�[?��epǤB��'���%;Z|����?�V�����4���OoĨo��E��7�-����Hn���RЙ�5sid3`��1=�k���mk
�KaF��k��W<��硹�Cz	�*��~��D�C���"�^�&����J|��[�x��ul�'��f-ZI���Qb��z��G�O7����c����6H�d
4˴*�G�ȷ�/�� .��#�.<�ۥ*v13ޢ/��M��O�O����M�H���?��Vdl1�L�L� ���&^�ό��u:O	��jG	�_Jh�$�j�T<��oC�n 2�����|t��F>K�%p$������C�[m���Q���[|���k�"ҽϙS�ޔ2'�\ܶ���na��~`|��������R[�**�H=����P�#��nA;ǳ@��F�;�Ϭ]H��o��q�����Y+TO���b:�JJ���;�,�n&̅��L�u��{�}d�����T��q���[��=�C���Y��?Ig��D]����K(_�ܮ�ɞ��(%O�=���f���6�}`i߳\�D��p�;ݦ&�DC�����4q�,[_��>͔��^�Vg� �et�0��bB�,5�,� �<�}3Rp���ε6Z��c�W�t�NȝY�)�9�3�ڮW���D¡)e��:�3�[]����ߓ�N������dA������F&7i)�7����la膆س[4c�����G��Z�{ãн�*ܾ�񥳩-������.�ǃ�aй$~"�ڧ ���!3�.�=�V�Iqm>�P�T�X'Gh�MBm1	4x�����#�1^�B�K<A��	��ځ����r羜���µ*N�<eB����po��_��.jгoB���򝫧A�~ī/S�3��l�WǟU���4�j['FG���D�4���[6�/�l��wN 7X�~�.˩�i#����L�[�6��e�s��1A���I��x�b[�� �!+�Q��'��1�2XH�I��K�A\K��@+!.��W��!E�d���|��E|K�CvJ���Y�+Nv~�K����2��DԎGyͷW��)�n�K�ʊ�m���-)�J(����&%K2�*� ����&ʂ���O�6�G��C���9`g�Dvh�Y�}U����{��B���\FZmn_#Y��R��v�%c$b����m]���o�(����zh�{j�+V ��8vP����u �`vJ�]���Ϟ�:���Aܴ�h��	�m�e�
Ieq���]K��#v����lsK�)چi��"��$�PGzɬ��#�)� ݔ��`�c��&�$�5+8X��v�@<Y�O�q���������o�GO|�k���%(�r�a�:�^`�h�������^� �	�r����0�J��������]15�J���e���dܘ�VI+�ozbh	���D�f͚�D���: �
�WM\�V�񷴐��h$�/,c���E��5~��MY3�6��k�Ix���Bn�ι��������탮5$���U\/Ɉ�M\�;,6~�m/u"�FRR��ۤX	G�ח�܊ �G�?
/�ܠ)�K���"����`qN��9�쨸�so�
�O}�|��0�noИQ�};�Z^
�Bv�J��ZF��#�F�\K�!���>c#-<ښJ�샋���#p�� ߼"�.V�6f�)�7�����?���I(����X[ �a��v��KC�u���3M��
�_$�]H���Jʈ�K�82�����f� /�(��\7��N�s�}�DkȈ���(���ؾ�w9����6��"����^.�h�5�V�2����d�#N���ެ_��S�~��o\����B�j�A7b�G���9t����0��~�IOи}_�	�c<('�� ޠ>Gx�Itv����:�T:�\���������4��&�����g�k�i�w�z��� G��W��;�#8��#t��?�y�'����x�&>l��d�d��tj1\���N�j�Q���MD��SI�M��d0�j���AI/wQq��i�1��2&�e3�9�@V�^@��-���}��
�W(ޚq�8�L��(�^q?���c�pd��Fe���(��[���Aԁ���F$�����	&��>7����G�����<C��a?ma �e�ޜP��*Ֆ	]�q��MWxcnQ�@�u�wn)#>��мC5(��$��!���j�}��W�pmho�LB�D�'%��p<<\����G�V��3��?�YW$M��\���`x'ͮ�]�?�~�£�y�o�.����x�IN�gF�i�k�x�.�It}nr�,��s

���L��I�TQ�<�G�)���y���z:~�<�߲����SQo؋������\�����0G�5����l6d���$2���0PI�n�\�}Z�7�efw�H��
5��=��4�)w��}��F����F���[�ο��^`sT��bb��#\5�Fʢ�Ę*��}��y6�u��"��?�wU����*���|jthW���)]��Z��Мu!8��kQ�;�����7dr�&d'\~��M�5w@w�w�34M������`�8���{X@�e�W�����\`�G+"�����&������r��ɴ���OD����d�a	�!%���=ln2�[��m���U��7qu���W>�G�����|Sߖ�A��.`G���k�_11*}8sI���:<����~�wpy�
��FWWg�4�(܀��p�*sz���U�V��x������ �v6�@�hY����E��LrQ������~�)ӭ�|j�a�"�e����*u^
��AV$O��|`������WuDum$�`d.����������ۛ�nK���=ig����v;:�Dܷ�V���`$l_W�{{c����6i3�Y�zl`_���K$ dwDT<.�"yoe����/���菟����-,M@Bļ89l"K���V��ׅc��:D��!�t�sB� �L�x��_�"����8?�G�K|�[���9��WZⲬ�8A��M�fև�^"��^�9��E%(���>����Cz�[Pb�����A�y���^h�]=Ay'Ѹ�Z�?���Q�����1.��3��8������&�����F�F���Y��6v�_���Ei	��G��k¿(����|-*�ϼ�K�Xߕ¨��jt�OIC�p���uz6kkc6iU�sׄ��3E��k���y��wc�ND�JdB��4@�6��V!՗�.���x�����q���@�5�?��V�騜��.��V<|���:�-��8m=���4�EQ����XE{�-�ҽ̹j��s1a;LMQ��m4�O
#�[׬L��~��&��7��H�������N#��R�ɸ��ƌ)yc{#����{F8\���GR��nu�^�W�.����_Bԅ�6�<O��^s��χ�u�ePGdA��ű��ՊṒ�,���K�v�M������D��x��>��(e�����\Ll�2`�@5]���k��q�����G
�_�wlZy�;X9�+�\��R��<t��n��C�6��c>�K��أU����Iq7Vk%��%�fGyw-�I���y��K|�H�K�j:��e2T�p����y�@z(���,/ l=o��L��ꪌ�gՍ�Z�d��ܐ���b�(f�%�7�����@X����{�Nܦ�~'�A�N��Ol�9�zu_M�[n��2�d����&/s
�Ku�4��ts�R��pԅqJ 6��?�ϑ���;���"��D\ (�YB�m9�^5��ĠF���=_����y�18r�H���b���� Ջ��HHډ#�!�z�6_�;��p7�=���n�Rw��8D:��QdJ�P6�í���o���v[ӂJN��v!�x��&E)�Ni�g�#����q��Ɉ1r����2���̓��,?��X����M���U�Gs�T��e������E����vb�.�dS�ǡ�P�0��cGIE=$\���;=ȓ�5k_�m����4��Y��g�*���Y�(Y|+g�b!�.��x
��Sr� �Q��g".�	�͗���΢�)ѐ����w���G+�y�[�я�3lB�f)��&s���F�E�'�dW����]��U�Hߡt��!���3��I�ww�F
���w&ң[��0~�+i�'Z�v�:���Ճ�U9IP����Q�5ܓ�6�
V�a��8�4�~�0�v�Z��_%�k�дס�$�%�a��olc�j�FN{_W+[<�/2l3��i���&w�Rj��"�Є� �?̽�i����M ���`(U�0%玁�n;dc�?'&��"U&Q5�s�=g@�Ʋ]0��fɊ�*�K'f��:F3���cd�fQT�wT�:�%�OO���<���蟩5:_��p,��CZ����`/�!����xEwHFTOWw�tDU��T�N��yv�� �|WC��э}�6�Ww�*�d��b�i��o�v �]-pmYs��N�"����[ps�ʤi~V?X��T�����Ι��Сo�}�����S�mn��6e�&1��!�w�w��X�{P'�s.�GS�>�p&ɠ�@�~wA������G�M��Q�`;a�p��)L��펾	Ť`����*�)I33聋���.��	�F7H���t�o�"�YӒ��v�]X�[�S<c4�=�1<q��� b�-��LU�O���k�:�U�V�'�RT�1NV��~
�>> /��H0��I���N���RUùne�9��!G2y�d�.�|�kB�Ϡ�oNW���G$�4P��(��R@�%Å/�=�����?K�Mi�s/��X����8Gt��9����������]� i��yN#	��+V���ᇭ{n�C��=ml;x���E�Ȅʾ�����2��+�lC\(��n���/�8�S�$o8ۄ˭G�ɝ�uA�Q Ŵ�����?��`Bt1��>�jS[�lE�#|�wV ����a�CQ~}�Z��A�Q��+�DN���:����:�:M�^��1�6*Y� J����U
��*�,�gV�2����a���)�bK
]����|+V���P�"e���<Zlm����e)��B�R�{y�C`i�)��;,�=t<�撕C�X!���9��)�@��a�B/��.-Z/3M��J��벀�ҡ�T�Яk����e��I�a<���ś!K��"$a��ۍ=;n'�f;��z�at���E�H4w\�Z����T�?�2j�|�o�A�� -Kz�>�$[��K�RjA/���j�~�I�C�F-�!�ǐ c.ʭ�N5	�!�=5����9ͺEFF�x�b�L��$x�y���whDD9�-- � ^�;�)G1�Ч�|KH����[�A���0������4ʧ�cP߀V8_U��(,�VX��o"&�㯕�%�R�n��1�; ��Tv.Q���{D��=�T6m{�I��(�jlN����R�G��A�'Hzo��&0�H�`Mܑ|j�X5S"o���W��7UC)�
�q'�/W�mP3��	o���N�Nű�K��.M�4I�@��pP1�e�}d�o��:�$i��<B�6z��
�͢6�"|IT���S.�=�ֺ�����8�%��G��/�A�^dS��9�܇F)�W+ ��f�`$�h�����"�n�P�xR��D�-%�I\dP��T�
߽B,%����M�s�"#Ҫ��58�����	��=]B��9��U1����u��f{�|��Ybw�{`���d�F���&���_Q���m�7�X�=U���7`I�A'��:`�x\����Y��E"�q"���?r0i;�ea�Vώ,��甸1)X�ڨ{��Dhώ<i~�W�{�S�I˲���щ�׍���]M��inՑ��K��%+�Z�U��R��.N�����o�QF��������`��t�F����"��Mƽ$`sEf�2#��,Ė�1Ѝs�����/�J|�H~���;-��ن�c�v�O�������k�Yǝ*��ġ9��b�����bd���۷�w��!�p�b]�4���U�W�3� ��.b���]wj{V�6�8����C+��6�4�~0)K�t�{��k��Gw���e;��{���U߾�ʯ ��B�rQe1����2�V�_<O��)'RL�몢�|wt6�c?3�e����O���KHiU5K��3�١�i��>����0����Wm'\[de�\4C��]��a.h^F�:-v��_�q%/�Ȃ��nQ�U�Gn�'v�i8�*< &+23���b�k�lCʺA	RS��e�Q!=�B,f���Ft�W��<��2���V��۟�	�$N!v���z$�@VZ��1GI�Q��;G�9н�tQ��A+,�2̛��V��\U��fq���Q�[�O!�E �{/?nB��GW�"K$�Ĺ�,�d�;VOG7*k�U�2Jp�/�21 G����YF�FW'~��ق^�2_�/ �[��y�*�Я�*m���[z�CfSu����ә8��d�S�,��}erDe}n!��1�|6�jk��Y{�<+F��[�� ��ʲ�V��}��
�_�\��r6��ec}��Eg�`
�J#�l	OiE�d=�
lW"�o�C��,���uz��WOg E���	aQ:�'`�mA�rȲD���K�Q��}�]��� ���
L�����=����̬q��뀔dM�
08&	'��bK�B}U�k��XG`3����W�D͎��:E�|`�=Z�n|"H��s���2����H���WRD9�4W�kBh�r���庴|���h�N6��"J53�;��
�?���\�QL�C�	��l�DCH�v��d��|A���&Sy�����R�X���O&���2�i�3� Q�l�p��e߼}'�u&Lmg���pv�����pO�|jĒ�=�)"�j�.���z[[�;.v�@��R�X�"6KʮwA:��;{k?�Jj��w%��^{;�/2(AeJ�ɇ��C<�ߠa��Ul����"�C�0�0G=ē�(⾜�>I�\ ����2k�r�'V��h����C�;ǁ�9�28�w�n�Oe�P�M��i¶T����:��$��^W�������#��m�ݱ�L��+W��%d�,���C�k$����_������ ����!R�c&�ݳ�W��Kl'�_U_kg�e�(��Sr��:��oǵjĹ�ï�=��WwW�s��;mp��f°� �ɥ�(�67�ߡ��$Z��:f�\�HDͤ;L�C}H
��Y0)�E*�ꃗ�S��.��ݑ��5�,^(!��[�8��Gt��y�w�b�*��B����uMѢo�Q��Fz@�OS�1Qn�)�&gH˶F��^�iP�M$�w@�������ꂝ�&.�|$�W��\X��DnD�%���73�Θ�|l3�R�.uק�O����Ճ�S�34د��ݮ����Iş��eET��%�]s��?��</�g�M?�Ȑ$��`�U^�{�J�F���G��L~��s�FH�
��T�#�=�c�"Z-�:���3S���ϯP��Ԫf.ro(�A9iU�x
�y<D��3�������PN�$����T\����6 ��	�[,��	����|>�I`���5��ҧ��F0�j�JBFRR��l���֋{�:d������0A]M�̉YYs��d��A��|dMRӯ�`�8��
{�t���(SS^��Ԩ��E� �7�5x��F�(TL1��? ����d:����:���F��c%RPF�x����-�K���l+扭����g�>����ao�����(c:xB1��Yŏ���uc,�I(��a$�hO�s��Y�Zxj�[�m�u9�{X�
�U�t��$N�m�����\1�L�n����#�F&60;�������*kKJ��'����;V
��]&T�(�y��������#���>-�'%��Ɖ
�U�*t������e8*Vfh�	���Dz�"K�&#����A�t�x��Y������B�nMD���A��fEܨ���!�(�һa!�U����L�gJ?
]
j����ߡ����{ò	ړtV�|-��ahI���~_��nF#s��4m/0��p*�f� �h"	��v�XL��eF��Zw0��WQ&��Bc�+��ɟ�k��Ik����!L�$ig;m&�ȳ�t7�fUs�Wq�P�b��{ f�܉�R&�����UP��EI8���;r�(g<�P���%$��S��ڕVq��D��	P��&K�C:���n���3EnyE���*�@bO 
t�$���5�K�o�k0sW!Z���h�>e�2�]���c3H#?R�	 ^U'"�2y;���QO=h�E����c����j�f�4��P�Yw"��8�D�vHc�s��\��;�n9���"�`��Y���	�)����̖L�/`F�<q.q�u���?�F�t����x��Šѭ�|D�#EC��lo˻V��9�J�!�BƌN8���fv/���]
iXUĊ'���0��[�K�9�Ԡ2Z�$��4�!f�C#߭P�$zH)�i�"jb h�Dm|j�y���
�x�+��J>�D�2޺�{��	����mO��;k'W��v=.>�!*	���6�7$D�?^Q�K�j���\|�+L:{#-�o:��� 2�w�R��ё]\���x#��,��d8��e�s�g���'���7�d�|��@��d5�"��e	��
"�
~�y�� �x�ߑ�Fv�D^<a���2��x�4ԭ�g�sa�9��-uR�ga,ou ���Y��|"m�/ѶA8����o���������i�9���Y�6#�h�D�.0������bWjn�uS�o�?���TDD�vR����4�:��Le��c���X�G�޷�j�C,f� �����6��>Rk5����r���r��T\�q�e�<���t�"\��G��9���=_q��-Z1����|R��(?��u�j'��b*���``_+���5T*���b�Ó�'�K��:):D��	���.���|HH��]�if��#U�Ή�c�J�7M��������8}�&A�3��Uf=]�@5ş��)9f#F}y:�:�Wӆr_tz���.��b-�dN~NS�&|bccx,�/�*���ҩԥ�,2���p���_z_ �v�|�a���	�=������B㡒v"��G�v���TՒ�+���S^3ȞO9�T�|��=����#I�ne����v �=W�M��.E$=���R�A��/�H�*9���벵�e^g0��}d��Xvu_�Ro��ǲ���{�t`�?��O�
�� V�HAV_�M Zaϙ{�"-&��A9˩���t�3Le���l��j�|��-�C�TsJ��H_
i\|�v�7�O��s��M�-έ!/g�2�q�G���ۆ6�w�����Z.�sA����u_�<����g�rB�}�s3C�����N?�Jt��M	- RQZ��W!pH���S�e ��t�9#�fH
7��jׄq\����e�'\�|x��e6@�K�t>S����֡�\���9l.�@���uG[]�A�9vX����G�WW��ҿCn�fB�A���C���+bC�g��X"̖�ZJ!�ڽ�_�S���#��}��6Gه�u��,7�|3Z!$��=�+K�����4����s��>�l�.Ƶ	��S��D�$��t���0�8��&��9�����-��El?Z������=*W�t�b���e3��r�9@��8��"����ƥ���B���	#������(�-�g'C�_��Dx��ZqAѪ�7R)[��d{ #���BОf�{��4�<��=9��`�&O��O��e�����%~��A�d�cu�H�xTw����Fa��߲���5J��B�����)�^��;�n���Z����[��-�f\$�.�Վv��:�2J�Ƒn��y!׹��Pc;&SH�	��Z�7L,�g+=VE��f(p��Xڨ�KE���#�28@��G�>2{,�3��pM��dɒ���o*������V9No�C�����v\/IXn3$B��bU����eU����)��,d���' +�ػ�Z���1d�Dz��xU�'V��6�t,8h9�#^�P�����q�Hj�����cL����k�Dd`*5<�����	XG�e�5�^������ER�1�Ϙ<t������O�K��V�}O�@�s�P٧�͠f}2�X��hF+gѺI��(��QI�O���Vg_�/r�wFQ���I�T�w옴1�o���1�����4y�7Č	C����}쥩ΑFW捣7����� O>���h��z�|��n%��=�,Iֆ�U}����"�u/��o7�	I�F��6�:�c�}������oנ^���A�%O�OB6�TWN�y�#77��K����R4dǴS-��f��`k`'��W���YˍU2.�{j�L�u��["f�T+KP2I1�̬0F�v�!���9�YAGʫ����'rv25cx�x�3[)����|S���OXoޝ��:���~�˺R�l&��׷��z*����eSθh3�Nq��N���5gչMϷ�	3���E9�%�� �Q�C��9,�HK���¿�3k>�s=�.�~���S9s0ޙ5���[���S�����")��Puw*(�Yg�|��ȡ�ژ�Vp �I�>�[�H�O��$����d��?L�c��1WsT]%��H�U�*k{��劵!��eT�̈́�`���|_�3�ׁ���J���ጝ���5���wɡ�4�FZ3�'��fr�2�	)q�*�J����c�5�)o� ��*n��>�.�oJ�+��@}�VqlQ��P ����ℽO�%y���gX��M"���)�MS��M�L���ln�wl�-�%A�DV�af5�J��-�±�zܱ�G|˥S8���1d�'M)y~���^�zZs(�rb�����e�{���~TS�;a��k����C��Cή��zh�~�ڳƒl.����t
5X�P<~�b��֦d'_}7M��g�Lb����9���j��E2I�«��ۜ7H*��d�w\�*�mn�e>b�����4Ĕ��=�^���
Jq�zKb�ҏ'�\+�\�0X֝����o��?�b��{1��`u�{���RR,g[�>��e����A�0���,�$�;U�y�mPy���@2�&�tn2o}�R*�}�j\!K4l?� ��{�b���䍌ѕ�{��b�۸<��H�ukI7��o������@%N&����@u䧵Wyd@�񧢟�1��n�"*�3D0�z�w9c�������J\�Ww�R:A�e�t�̹3��vq4K�֫�RL�),�Z�gG��L��?��
t�n�;������s�8h��"�'�;�PS�t-��6LMK &ܝ�%Q7�=�O���꫋�S�=
���C�R�������C�Zj`���"�,�9�$�
���ϊ@��K��|��Xh��l�u�%�	��$���č_���U%_Z)�$4��u�(�D�](��"�L \G_k����h4z?��y-m�n�d���>��Lj;�k&(W�u�"��
�\5	F�v.!��H@��^h���'� ��Da�j݀����-��1S�9����ߤ���S+nB��E#�h ��sE'�.V�/�-��U9���&­We$s�FA��R[2׆2���]`�"�)g9��:���$e"�!�`�-%p�q�$L��L�<#�c��˂��ܼ�g�2����3��'��G;�Jim�� LF��t�]G1neo=�	��.����v` 8��{&��F�w#��ܮ�r�U�
uP�9f릻��a���}�.�by;���
��M�b�D.�MDҸӑQ��9�n]TA����@��	��؍�s6�Z�S�8��)����Sk�4��xɴ)�g"{���D�����- 
�[��a9�-�(�T��},�hOA�>��T/����¹A��x�k���Ƽ���nu���n-�0Ǖ����&�=(��bd N�O����]�r �r��3��a5������r�!�˛��j ߤ#��d��Xɘc	h�ܠH6}�b7[a����GU��t��Ci7�_�;�އ�Rd�w�X�wR�L���{?�F��<0�����{޾W��
0"ω���ue|�G�`ؙ��^�����&H�����SȀl�45���U�T�p��:u���Zڬր��8�����G�Ҝ�"���d��_�L1�)�ϰ�43Ks_���إ����6�sZ�m£'$���U�2��n+�#(�!�^�}"*�M ��y)d)7�\�1�S�?��$%��RP�H?L�NU{>����~ F�E2����۩Y�W��凉��~ቢ��ü�P�Z��� �IZ�˅�Du(��ﯬ݂QC8�}v��{.'���A��D�s�G���t����0��M��m)A]�ߗCW���Dg�Dz��5�1���ߓԼ��5��w�Ĭjӹ�d��]_u݀8�[+��.?�iޠ������?�����Y����ٷ���"c��a�].��9�ޏ'A'=>�q��җQ4<'c���d�lS����C�Y`�L����}�Ն�I'��g��D޶8�j�e�'��1;=��a����� y�\Qk�RA�3��D*�U�#�)gb�JO��_KoӇs�!���a�c���Q�ŧ����#d���+�M�u&�G޳(V&�� 1�� �ٮ���nA&:VT��l8=K�o���<4'T����&���^̾1�E������6�*�Oa#M_����JَcI
�$�5�Ko�a����҅�зi8>.b�62�o�x
z�P2�{oN��V�b��_K�
U=O�2��(��lj�m�D"�6��*�C�w��>��%��{����
��Y��W�{!��j)@��~� �_<ߌ�P�jvn� 3e�G� �N�:S2��+��(G>,�l�?��2�H�諪�A����InRu����ej�p,��2�OV��OX?��XHƸɐg�^|Pj"-ִW�:''r��R촺'�Ǚ�	{ژ��d�@���y��ZpluQ���.1��L3��Ǧ�fG��'I���E��������g}eu�ge�F�7c�A�
>o�P�cD�_�fi�3��?���e�f&?��_����}��RKtGj~f� O��Mp�'��=G8�K������Al9Q�\kԬ�o�K�_�����a�Me�	z���~�{��e���x	Ptn��a�M %ܔjdL7R|e�y����eb_s�`Tb��_��9Qe¾9��;7��v�77��Q[[��g����ŷ���Р�^��v��H�����ۤ����k�Q�v)�,w�����U�mF�F e�@����S���]%�@����&�{�9����д�D]P1��VΨִ�1��"nrX�;�Qr��
�!��0�P�&���!�6)��+Xs��ƈh�X8e��~C.��`� }s1����9�[nE��N��<&Ԑ2�И��|i�"ֿ��@}�VV��M��u��gޙ��}M(����:nK`���������~i�����0GŹ-?�OCdc$N�I�A��8���O��ʈ�vN$��l�����.���`C�����X��#ό�ىÄ �/�����>�d�����=S	j��	s~���<B���D�+B����լ�*9tE���Bb�a|�~�:�	U�F�k�dU� 7a�`r_�v�?�
(�bb����ş�t9.�̣����Ԉť�:f8�7 TB�%����`�JD�׺.D�:�ߑ�'T%��5�XjP�aD�݈x(�/sy�h����_{Txcu�o;>�Eo��M_wY�����6��F�4�1��s���y)2�l�����V�ڂe�'F�r��Ƌ��t��*���p���t��]yyD�V�ڟ��]��8u%�k7y�w+! 8�9Ѻ [�,F�B�*��aK���󂊠���n
%�ʓ�)�+��=�R5�!������)C_X���Oո�,�h<�.��Xp�V<J ���'JE���.���~��OG�~1��L�x�o+#-6�i�k� �<�h�%�4y��e8V>��i��//��^9��6�#A�K����K�u�54����H�E�wh˄���v��T����2t�!/���ROja�#<2�<^��<MtJ�>c��<�� �(�m�;�S�5���Ӆ�eD��ce�S�R����?�����Ϙ~ZO��������� �2�T*�t��~�E����H�D~7�0���^ �<Y����\�A��Fd+�%�-�s_��IQ�N��d��Z�Rk�ǔ����Ƨ�zY�����?42�Yף'����ZB@���F�	s˺^e4|2��+�	�~S����W�<5^��ͅ��i�䇨*p�GPz��E}�_�S�Xb�$�D����e�+�Z�aW�A;lC(��'�e�55���1���ױ���ǿ['q�~��5��+*ȧ�X{� ER�w�V�s��/�;�<if�y� ,,m�̨�D�4D����H@��v�O\mw5��z��k.N��\w�G~E�H��-G�I��	Ӿٹ�$�i��zl��x���U��P,Zry.M�t�5��!W,VL�*F��&�'�A'�4��.�9��K&3/)�;����F�%�Y� ��N˩�JE@��+aT�il ���r����ji���<�̌�֠��$Ӿa�F<}��U�mPivo&�酝\M��槃��Q�@�+L`��;�����-�=u-�����
��9���)'n���kH�����unPBS�ZxJע(k30��"�c��Q�A�JQ}�ry���澵��B����E�{�ݸ���Wz+�K��W$Nl�K�Ix�u>�/Z���QU�Qg̷��|9$��3M,i�ؽ�y�:���a+�H\��G�d�xp�[���${Sb����:2N��5-�y�iĮ�x�;��L�6z��e��e�εyx��at��M�g�WAZ�	arp���|]��	uS��MP%���?�d-?�ƄŮ�����k��0N��I�NM�x[�}�w��S�'��G}h߫B
�f�P�teQ�*s�*�IH
�|l %PD!'vIl��$LK"��K~ȅ^��u��76�~O�|L)&���߇<�tI��Q*WɧE��aQ#W�V�Zr��>�Ъh��YwM���9�l�Xo�w�:�d��E�i��4�Z�Mp���bQ�q���(���('�A뵈$��J�Ja�,��}J��:xz�����c�<���1�p�>�W�n���Z��1�����	��ـx�Nc��3�!�FS�_V�狥e�Ѹ�yޟ��o��>M��@�H����߱��Hv�zU~�J���z��ni��$�&ݬ����x{��Y-)J�L .���J~�'�6`%������>�"��kx��Ҟ��>�x�@M�:t��"ͦz���(�v���<j����3�Q�$2)1Q�ݮ�V*m/t&%y�8
i�����&%�8��X���U�,��ӊ�@��<e5��E �G<Ӧ<�	��OX����+Sm�PlIl�t�������4s����#���ҧ��n93�oS����� &�8��OX���߾	��v��HCޠ��%�Q?W�g�����z#|I~t��fڋoKA < �~�k�:H3|q����h8���#�%�+mP�Q��Y��^}	5ēNo��}�-��aC]�)�#�����d)Vs��ѐk�[q^N��>0SB}��_Q���L.�Y�=�vՆ -Zd�ᮬG�%@6�N3�2�b�
�m���X��٠ς�~��s��6�ژ�;<���ʺa���r���]���;Уv�a8�у��yg/�A\��۾�?'1�@� ����ά�3v3��L���d��P�M�)���*��+E'�+�7���Ղ�9a��I�cZ��u���'��ar/ܐ��Mc<���^VZ�2)hc��p���(Vj���"��`��q�x���NŎ���_6��kq��nL��F朴��'��R�դ #��E ��G�� ܔo�4[��"���x����5sZ�_�V^�{��T�x��0���-=�����:T�����>y�[)ߣz���-T���8�&���0��R���ܻhtr���5_���[�ҙ?�������k\�FEKY���iR��1��0���������XkwX�S��k���o���<�s�wi&c�}�X	h���a�53/�����S;���`�0�@���^=�8�Ŝ��i&Q�e��j$m�c�t�E�hJ+���4������i

��`��Z=�����IVE�V���F�=��S6�XD���˫U��imH���k����������r�l��"����;�$✫W�b���V���rqq���0��@�є����ƭۭF4a��:cd{D�[��&�[��L=]z�s#����߅$!nW���ҟUB��X ~��x���\bṂAs��Ya�`X#R�ၳ/۔����Wx�s0�?��$]gL�!�MB�XNub�LYBƂ��G)��Dĥ~W�z�� '�[STf�*��	��u"U�Ut��ѱ��}F������W0߲^�٦V�Ég����w��9��a|WK��o!�#u.�7�xpG�bΜ��N����m)M[*Q�Ʈ����2��b#[�%Ã�����,���{P;��ڲ���&��,�e���6����;l䉹��m`�NL�<}�!�z͗��KM.�@��~�%ߐ�j�e�BPn뇠!"�w,K���K�	~�O�:i�$tB"K��8����?	s`��f�<�9���{�}^3W��_[�y%�l�,�v�%�&�lA��+�]��-+�5�:p�2�n�
�q8�z���L��P�]�:ǁ�\�q��;�THu �
c��|i���я@��i(
��4\t�~�A��d��QtqR�w�\A��=���\=�5�č���6�����*E)8��Tbvw��jy�G�\�4)_����r����n���=Ƴ����nj���;�B&9Φ������� �B�K�)�{���\�k%N[	&L�N�����'r��nL��˔�djEg�^�0�!�.v�4�BB�L�XO�XY�U�t��*��C 0D5��B�8r�|M3�'8�g����c�¦c֤��
۞��p�U������_���:)r�q���^?Y��;8��%߱ �"�S�*�TS�L,IƟO�q_&~[g<B���c@�,�(�1�^Ϟ�"r<gC���Aq�z���$�Ul0�Ȟ+��Aq�&�������E�a���Xo��ԅ#LՔ�T���&�mv?q�||�".����ArAy[J��A2��Z4o�m��D*%(_K�n����̃_�:���`����}�'�R��r������^�R�d�l��0�G_�$1�P�1.z�gZ��k+�
�~;N+ak��KFQ 7.�ǃ���;O���B����f�@����%Y�q��aI���g�:(��qUT�<	�HuxE��Z�zN�p��n���7ć�7�g{Vr�zr^���vO��QW^Fa��Ȇ${��
T���A��HQ�sx�ߪ�ܑzDqç���QF�U��d���&/��s�-�� U�Z� ЖbBwW�(#��~�mph�k���^iE�������dp
�0p��!{BY\h��v䴛a����/{�$�0��uwl��5�^$�"P�a(2������ƹ'��d�	�N%���ϒx�ɷγ��e�펊vu���-��}®��oX#̝&;1��W��)��C�a~��/V4/�CI�d�c������G����[A��`Y޲�� NT�V��K1Y3+�E^�g֬`Y�fp�}D@�`�0�����f�D�e���=�0%4!��z��V�>�oY�r��x�FzMZ�QɉU��yt��Nw;��dg���}/��,�����S>�N@�M����D����Ե��p:�Y����R� ����f�jS�����"����c����tB�j�萺۵߮++]��r��i��͖{o)���n�n�5�s��E�>&�M_�\2שޱP���#yOS��+F�cK���'�a��܌3�Wz�H��Z�qj�[�ea&��C��#��I�n��/c-����3HE��S���H����F�1�d�W\�ݵ*D鳁���Q�u�E�W`��F�;-��B����X�:�f��~�:5p�=���K��?b� ����Ak,��ؿh^�$Y�Gqe�$��{�jW�i*�C<ä��=�zxj����M�tɑ6~�W9�0J��� T���B��63k�y�+�GJx�n#$�.4 nǋ���2�)��D�f!T8�/s�4� �;K�~���o�k�у�7t~p�ġ���h�6��'.F	n�P�X]�7�w�����eI��G���B*CK!�6�Y�a�%'&�*X��Q[YD���1�%�>9X�{��Fl���/���>���~c1M�:+ �57��ؼ���{^*�7m�=]gd��Si�_�I�H��#K��Sv��]�X+���ﳊ���(|���Րl����n�;��WExVn��qqψ?�r}���O���[YF}(��0�ie_�k��� �����ٛ�$���M
�y���$M���	���6>W�U�a��� b^���R�@�g;p�� ^;�g)9!6�~%$�I����k��+��yf�.ҿrހIl~:Tд�k�myR`�S�	�7_ӈ�������{�@h�R��l�OxD_!Ô9!���)r��bG�5����"�-N�JFV��>��9@��2-?ԭ�u}��[;P�-(�쌨XZW���������}�]��6���Ȭt׷��Yޫ��~[����O?u�L��9���8M�NE��g��[�+ӟ9 :-�dx����*9k�=uN;���U�]TϨA���$rU�c�:+Ĳ�w�*cz�	Y �?�`����kF�t�1%�Dӕ"#g�苵����02�4�,8��=�4ק� �ҁ��!��ygYG�64_(�90\o
N9�bo���vQ�n��!Ge�g4P^ȏ�y�x��CP�����V��}JG�f:ԠÙj6�ZX*�C�j�k��w��C�'�e��z�j�<[�u
:༢"�D*EQ�K�<mU-�(��g��E���-7O�g�F3cM�hׄ����g��R�&�j�f�)k���5���X����L�t�'��[�~�H}� -��'X7p(�Y#k��%R�Fg�N���py����ֶ�O�"��=��,1K~4D���9�-��"3h@fS4S�7����xy�X�n����X�Y���lf)�ʇ��p@��0������,����TR@ߪd�%i�J�Rrn
.�0�]g&�h29!HI��B��]_�9���
3���GS�ȅ����B��i����-$�U��b���D���S橗ǧ��)H��
���4��Zټ����<��y<zj�D��x5�5�Ӽog���nou<�᧛�vI�B���%fg�L���Tp��,�<��f$վ��7@�Kr�L�Z�����ʔ�d0�n����U:�^ڃe,8��U���E�=�B�b����λ>]�7�7�}̮��A�7�z�O�v�Ih�^��Nk:��rT�t���K��rt��"G��k�W" c�Ÿ���^�b�ic������"+]<�q�����

��1dqL����i�po�	-I��8�܈��|��h�.�'�UV�cr_�~!z��Oa-$Ա�!�m�7Ź}��KE6��JNq����W��Ph#�a��`[q���H�^np���.��,�i�je85�^��"�|�u�1r�.��3��q��`'U�d$�L������*uͰM�3�',�s*E�|�]krx���l���81>��~Ϲ��E��>�3��_����	�%K�NM'�?p�঄�Q�v,ɧ�j-��ڛLH��u4�n����d���}��B���g�U�.�D���$Wf��V�)�+�3���n��FN4��gk&ĺ"�%�_Zo	h� r�G����sH����B�f F) z{��i�P��db����i���
C
����7{��^ ��F7�@��/,����'� p�_��*|P��c�,�0|��Dӎ����������Ǚ���X]i�j��6Fb��2�3/�7$���B� ����PYΥF�x��b����5V��f�R�� �
��a���C��C9�7YiI��]��e�U^���=<�qz�)^�\v���=�Q���J�h�wT�������e�09�a��m"��f���h����h#�$���t�Νr��#y��v����a�4T�*1�݈3�Xq̓-d���pg���`h�\���l(6��X������pԨ�q����c��CjEOH���>��L�4"�}FS��v8�Nh�����D�uA8�O���^�ql����5Uh�p�3x��F̣������� (��I��,���2���'�f�/\�L
2���Η[tNN����n�#��(�S���tn�AtQ�h�\Y)��G�吏�z\$vh�?���{2�$�{�a�b}-Rv.w%�9�x!+�ϘŁ�)����@�KV�>S�>aRe�$���iz�y�Y�'C,������yt\wɹޢE�A�a8�w]�"M2��i�lyan}����Z�7wr�-jf`E;�:�LhZ���D
��?A�&�䍠ٚ;sn�K��X�:S\�[)��
�M��M�ڃ�-Ot�0�%͜v��{����z0%���2[ fD1B�U�B/Y��Q����nyVX!M��фTٻ7�4�j����i��-Cbrie��e�N�mKE��8=�-]�|�O�	��> C&V����Ց����5��k2�G��|�rr�-��h���� >�B>�@]6'srM�z���V2�C�^pc�T'�S6�Rv�	}�W�V��}��<�t���_�����GAs��v%]��X�/���f��0g�i�����������9���-��	W�f�b0�e�6�d��e-��?7���^%~1��wnN]br��|Ny�)63ڠ�L�}�t��>�u�(T��k����pd�0��Vւy4Ba>j�Tq��j�v�G���p�F�I(*��7忌���B� !�9���`�(�#�:�п�D"����3v�yq�e16I4��$MMN���:63ݷWk�[��ͅ⹴�2@5���&BCg�p�p���V�XL��uc/��ʊ�NL_�TU@D�z��<��T=��$�'�xH�ݶ&��=��E@'�g��
@���z�[��vP���G};b[�?�-��q�>DA��hM��+(n�����	�Q� �$�u�3J�{��]����=��.Հ����l�Dsh��W��B�|6�v�D�ھ�`��S���S�����(�H�?��r'8I�2r��P��Tا��?W
�RD�-g�_�2)�G'��i���]�dP��F��� �{�>�g��A���髲|͠��Q���ɲ�"Վ�P���ԧ�u�\��l����� ��3M�����ثÓ|�,b:V��H�̮_�6���ё�I�J9}�$<k��|���{�`�h�P��])�8B��m�\�56�\螘�{���~z���P���r>����~����~��}y�vVIq��ǰq�i@�;�icz�sbc�_��ng�כ�jW�s>������Z-��NcT�� �B���1+>���z��,d������R�[��p��rlOvl\�*c�$���+�Bo���:���}��Ip���Y(EmEᴝ�yԮ��3��
�<���������-��c�Nh���ˬ\N�pVʺ�}��MFt��hS�]�g�~R�%�Q�D��:�zގgȇ}(^�3�1[CF��AX0�v��]ùP~��'+.�+��N[]b2A{�ERUl�
%�I�6�wa�фEn�÷��)�������qm�d���:���O3���6���*g��.��>DTЖ��x�s�3�O�B�O�G�*MT{FK�r%å�	y�{ۘ�8���;����`X�T���=uPGg8)��>�]?pKJE��g�i�]=ޑkPa6�&Z5��4j�����7W{�ċFA ��HU�އf��z��x6l�o5V��'/��>8<��^&�{ M�b��=�m�E�]� �?��ˇsM":uF�O�Nn�y.^ަC0�# V��I��L˝�h��^�6�WO�G���z<��_
���������hc�;��ֻv�����I��*/�`ݾ�Bt(Tw�fk�i��^W~Eט�5����`ǒ�H ���T����9^�2�;2�_�y�*���-=�B�
����ʎ{F�L�+sl�mz?x�-�hQ��"z�vv|v/�;�{���Nё������H+,e��~�}� "�4>&&zdz�z���C?C�p�ؒ��0������Tt����T��*p���([�n
��������Vp�J\6�r�/&H��(�H\�+�����|cG��}䲐����i����ؔ���$�{��:e gAF?��G�A���Bz�T�3��Jeϭo���CL�S��	9!����$N����	���T(h�E���#wPl9�J-�b�Afd�hi�tl|�FHI�n��Ḥ�6�c;��&>.���%��ȼ���A�f~5���/�*+(�~7�c��F�	)�+6"����Mv#��T�xY�\բ����o�D����܄M`+��.6/���\�+�U�n���L�@JАՐ'`�{L7D���W<�{���O6}L����N��㌗�ʑ���D}���=�y�lv�j��"��s�s��l�>E-���M������gӷ.��2��W.����,��ˋ��bs��E�������U���0�k��o��Ż�q�8y��@�~T/,�t���p$"�����;O��V��@"9m���}]�(1� �����	��C�,�g�*b�
�F�s���8���Sf����!J�����4@y�ǰ���Z��®x��.�m����A���g�D��֤�#M�Q�P���c	7�w��J�[]��/�G���N�wrU�N���;�)�O�������I0I�����o�j1pڞ45� EV��@�%����J��:��/-�B6����ͱ@���t�[p/uI�x#�m��J��q݊;&^*5`�ՎqmȠx�Uj��� "(d��k/
�i.�;k/�F�+X��#�ζJ�����^{�*���hq�|L	��w}D��^���l��[4N���`��=Oؗ�+ƒ��������RY���L?}�.r�DHKD� �S�@�!u�tV���'h'#���W^�n�ao����_���uy1z����3�7��`�4��]�ȽE�4�p��BC2ԁ�N�Ң���l�=���e�E���v�Z�V݆Z}(Iu��p�v$��̙P���D5W$P�3�^�G�:L�\7^��rN�y��U"2�k����,�,���]��F�%�1�M��hc�x�Ҁ���*�\5�����$4&����:�w��E��=�y<�.��'v?��9� � jU�������j��F�w����[o]�Dץ���U���jmXۊ8�m��?�oN���+9'�2�D8 z�x��.7�99�Lԋz���æ���ł�'�!=e1�L\َ
�ne�s&'��s� �%��e���bH�С��$�SK��P�J�����1�y(v�L��1�9ĉ"*#Q!�k������L�r��آ�B�V�Ԫ�p��Nh����-�]�⿫#Ł�P��!�G{�ύ�N���r;̾��:�޲Wt 2�{l2���A�@�s3;iG6�,,2�eGQ$�	�ϰn���c�~��l�H%�l�x[{��{	�������8a<��$�)Pn�zU����/�J�=�X^�63�0gV5�Zk��WN9�K�y�S�?[�Iț;7h5`��x�#.:X�@s���*�30��k��_ihL�t��zGc��;�G˫��, zJ1?���Y���:r�mw��-E͘������$k�q��x��ZX,��/u=��{���Wz)����<��d��L�L,L1G?�p!ۡL$8�i���4�H;���Ϯ�� ��7�ƳO����N*M*�4�s,�JU� �(+芜���m}���`-�i��en�T���$x�^��XhͬĶoM�}Z\w�<o�Z�����_�<_#�®�ØZ0��n�,��i�D��v�	V �δ��c42�;h����T�sr���L��8 D��eMu����y`��5�f���
�+��,ߏ�o?޶�L����Q�ـ���F�m���~����T�i}	ک5��=�=���ƵX�N,}o�C��0Ѽ#���fċF���r����-�ţWK�2��_�-�[X-�{�x�8/L���ә:M�^p�aN�� �l�nWW�A���gD,-�d�C�>�5d�	 �
�0�ܔ�0o��I��}!��`P�4%�m��Μ���}�1���K|ħ��?2�4�`P��498B�_R�-��J���R��v��xm���-��A�B��T���Y��n��"X�������H���~>-���*�y�>��k�X7����`�=h:������*	uq�j����/�������E���g���4ͺ�GЅ-ǣ8\�qΤ�J�
�ַ�vd8�Ғ��,q�^��P�<��B�'�eW�ɛ�L.ۙ�bm���m_b�#[(���5��]uF�ķa(?�5�f��O�_�Bx3zͻ���T��_n��=Ny<��η|`�m-�N���T����4�	������	��mj+��e�$㪁9`�D�.Ǽ"�V� ��OyT������a�M҆/$�{��x��=����4�I3�Fs�
9����raD0P��\GK��ڞt�~q'~4K:���/�_���1ܡ�C���{H5����ʈ��yq�;����|L�N�K����B}T�䘧�#�nU�G������1Ԓʵ�(��!��
Lوw�"QP������gd�8]!�X�S�N��Xf�7����)��P�}f�t��m-��9����k`����x�<}��z�}����:
�Ƴ_�s���f7��i�`���C�E)R��e3���Bq�[->��H�'���� �EG��U�#(
�`E)�5�E1��%�h:ﯫ�i�Ur�"� 5��h�T�@�"X� �H��R�j{q�7;)��g��Z*��O-m�w�ľ;^-m&�䡞MX�^��>'ɇ���m��N����(P����E�sK�>I�|�R�W\O�����!\�$ut�>%b�L|�#�*߭1�I�CI��
��K
�VLٖ����7���Tӓ��Q��f�>+1�!��;
;�fɍ��@4��T�G5�`�k�}�I��Y���ˉ����e����e��'w1�y$zˎ;[�#X���]6>����?���i���\?7h������s`�g�:�&�_�9�8EoΓfO��)��ljy_� �jrlm}���l��,ީY�UE�4��k�l�<BvҐ&!\]{Nit8�r帢����'8�9\�JF+.��I)v�lrhX:"��f�u/FT��h��H�-l;˘MԀ�������)u|:}��'����7�n�������q�"�<�dd��`� ��(a@�����R�})��M&A���t���3	�x�M�� (q[���3�:"B�7�������ގ���RôjP�`i%�Ʃ}K��w)���2�dA'_���\ݿ{�q�%�#Xn��d�=˪���r���ƾ�y4�6c\�5�(������I���ǽ����P�*1V9�]f��t[� ~�-�� }�����L�,L�Ρ5&HMK>@�����Z.��.*�NB[����hx �J�g�_��+"�$�qi��*��9QG|����۴)!_w�nw�e�s�� h)2 ��v>ږ�Y ���A��%����ו�*[k�HbYp  �0P�-�v��8���Y:����1���*i�V�+�G��|u�7(f�/0{���nOeu96J�@��[�yoԺ'i�Y�9J���ŀ%�[�pwyMǃ�v������|�M߸z>�N���^�% �{u�V�_��8���W�C�J}�
�$u�+���^<P�����ӧHc빝��1��pGc ,���'�j֌S�-Ʉ�����x\(VB�72�k�ߡ%_Ŗ�Lm���6;�z�$�ah<V��gE�W�	r����3�W�4:Upͬ�8H>d�;�;���Y��J�"X��c1�g�b�\�%��J��~^9��s���^2���l-lPñGSE�2��n	��@/�7>Wxo���ն2^�����/oؙ����N��O�1+L����Q��W����|$��Ա���ݚ�m���U�G���^��p�� ������&4�Z}O��սƱ�G���6��cՇ���t�⢗8����� o��>��x"�f)�Ը�(M��WPg/��xJ�s�N��~�	r�O*C;"��J���}n����_u���m��I���p��@?��l���HS�EBи�q����h�"5�"���\�'�_}=OQr�v�����]�+c�R�/LE~y�H��u� Jg�*>u�[�u6ȹZ�Ȥ�	'��8+,/<��-����YG�6�si��#���?ȇv��$G�2f�d,����,O����T�F��_���rR7�F��p�����g�w" �x���-[��"�L�#�~'�;E�M£�>z��/����M���?�f���ż����S�;�x�`����޺g�����Y��/4�zn�6�x����ǽ8��0B �!��Ҙ������p5���|�M��n*F�#�0+)]��?�$���l���xXK�Ey�:4�A�6(lm�q��L FB��gj'2�2_$X<���z@��8~�
&��JҲ���тΣB"��#�'����2��ܨS1�~��\[�W��h%�2/ë^G�x���T,�E�����<����9'5����	�V �������i�'GKP��eTPQ3{����ZE�Y�@��3��S3�S8�g��?�L��_�m۷0��F ����כ��ؚ4�i�r9:�2�;Sm=t.�q����-{�R��IL��,f��Rw��|J"u���3�3�-��O�؄�n�^���}>^�>@�������"��y�LCK�)Nj`�"E�	i
�~��Lr5c��Q�)��ǟ^� J�jS�ۻ�d�k^9/إ�!���Hx��뼖~��/��r+���`�Y�e�I�+�	ҧ_�� �q��A��.�nݺ.�_���H��t�ō�L�K�C���V�e�b���64�Z.PG,�����#b�v��v>e�P�&2���7Bx2әx�G�>݆�O���}��fž:i�t������S��ao<��X�~���;������U�vUC�p��0�ڴ�w��eF����k��&����u3�,�q��~�q˞�!7#��\A3f�v�)�~��]./Y%h.�����o vW�
��7?���V���O��¡�]�wm���7����� @����j�.4��z�����@%���l.�U.;�ae	oO�Ӿ�o���Si���k��H�p�˛��T*|ج�O	yΑ~�&�ڍV��*e���ؤ�4��@V�rq$T;�+	���q6X@qΊW�D��ٰ��āzeȍ|�,i7* �i)wO=U��g���ӳ<�����{A��L�� d~�?4K(��(6
G�yV��ZV�9�Cι��/��4�Z�ۍ@v�KY��h�NC��������=ٍ��C��!)�Kt�柛Ό�Хl�Z�B͚>��x@��)���I�(�j!l	�߳�V1��Ax9>n�$��@�f��9�OOg��XʂE�T���YMa��R8����>����h�Ƃ�F �f�lư4�6��
��|���,��ѥq,,`T���.�O�����������M�q`����g��}�`���k����:��0�v��ti����Z:<��%v�9فl�]��j;��E���BS�l�д#�p�V$Q��Œ����~�*�<uk9Y��#�B4��m����~J�:?��������B�B���
��eGE[T��t�5��Γ��TfpR�(,n�3'X�C&+���v��VL�Q��AgZ�ay����[s��� <0��jO6��uMx|�v���ݞ�Yr���ڐW�%F��p��Wӹ��N���\��hv��9S�(�Jө�2�ƞn9����Ķ���b�M$vx��{%��)�2�&(��ԗ�厅Ѐ�Rfyta��ʸ�f$�t{(�T�S���O+�q�I<���i��@Y�w��z��������È��/)���� �4������dCyί[��]���[�)�Ӿ@o�++�P%j����s�$E8�~;�T ml%q�Ӷ��Q���cv�ՇZ�u�N�4����B�$�{�F����N)�]�GdI�h�r���4Ir�,h��n^r�~��:E5���	6O*ǳ�O�5[��ӵ*C1�e�A�z`�>�)k���DN�Ձ��B�����	��F�%���h#Yѥz����YRA�#��fLt6g��~�D�y���Zh�~�3ʼ�/�ǭ���W5���W�b�Ѣ�vE�*4�����Y�%����aF�����c_���*���O'͘�1
��S�05�')��^%e��oXvP\���<���Ӻ���e���0䶊�=oh{�$��D]5���H��>d�����7
�fox�&��\�� ��4�Urٚ{z�1k� �+nGx�6��'�Lk�C*EGƳ$�`��-�v���@��Vtk�,8�ط��UŴV!ޥ��C���`^G�+w�z����N��}�ҹ�2�Ǹ|%p�S��`�v��[(w����};˭$t��ITh,]r�.#�_��Db�>�t�Kۻ2��C���e�4s�I`͆�S߄�A@�Y.;F��i53Hk���S:�p������
Ɍ�B��,���D��C�|m}Mt�r�B*����18(kF�h?�;?��R`����g����/��S^>�X�*��9�⧲=��)�w�{*P�=���?��-Eox��#�)I�� s��<������Xa24�Y]¼����#��y����
P��w�8Rk�Ādp$�$H��=�2_
�RG7��N����W$|l���Ǣ�T�p�ǜ�AI��rZۢ��oP�"�~M�n�1�'�� ^�r�� ��x5�S�4��l��ܙ��䦚d���NW͹��j��Q]��q.XR���n8��AWZɝa4w����Sn���K�W"��u��[���ii�>&U����]6�ӊ�%#�,���J=%Lgz|�`>0{�λIX�b	��+��5R� ��H�� q]?����1xm�������B՗��k�G�V�;�LL�u�����)� 6��[txF}�O�>�Q2�KP���S�8��FQ���0*S������Ḽ�0V3U�����[�<���&�D�O����*�xf!����)��>+v)��I����|�|�X�"����w�Ud�4G�P��чk}��� ������<�x��̃�_1�s�Jyc"�il�>��v����u�z��G�et��c���s=���W��������P��mM�w\���,_C��N0����Xf����z��j�}��_�������8+>� ��1��h���2����S+'�þ_@�����Ukc�S��?�g2������\����A�$R:���9�A��R��=�x7`����y�� 0��e�9 (��W�5�|�_Wv�>���vïb9	&�Qzs^��_�%��.�X��Ygｩ�a�yc�g��t!����o�\�,��4����/x,�����D�Wl�4T,Tem����d�ä]�X�8���X݌7�Aݏ��hD8?Wq̍�r7�
 i�i���]�}3�/�Pm�����_0�<�����l �����x2��V�`��Y��#�]�� �X?a�Fnlf��d��P�jנk��ᜉ쀬��|��E���=�������R���+�S[��^?�T�Z��k ��Q���:�K���P:��G��Ff;�6��N�"�ِۜeJ��>Yj�ؓ$U��������=͕UVɀB����4)m5a��4�����ةc�
��g��X� A#����pC�Z�~��0�ը�Ԉܽ���}�摯���sP� 8�C��ƭh2���	A�tz����T&~�e�S�����_*Yrԫ�W��ĥw��>~�X��֐�a��m�2���o�N4u/�l�j���IFf�+�va�������OX�Nɔ:�2�Ko�I7錋>A��A�_�y
(Z"S-�̷��G2>�q�T��e���;av-����G+.:���E;f4c�y��!���w�n�e�y��!��@nm?�n��򉠦ғ�u_�����@ȶ~�������ֆ�	�d{ُ�N�\�3�2;/�t�p8cM,WIl
0�X�P'�{�&���@!�P�ͱ���_y[r9O
�q3�;�1��
I�l�Е��B�~����X���Yֹ͛��(�9@���H&s+SS������Z�M��$�	�me����]��� ڬ��-Љb��9rjAZ���<6̚^T�gq(��t�^+_m�}�I����5�B�#I�/�������t�6�(�5a%�:F�H`�b��f��&��yulb;�|��|�k�F˅9��Z�p1��W�L��%��_i�l���E�Z{�va������Ǡ�W� 1�GDER�0�Gܥ9�:�h����}d'P!~n��;YU�����3��i�$=�-��8Cž�M4p0�^1��T��/3��y�W�Ips��2� ������o �w�:����Qb|���p%,aF��LCT2&8GɄ��6�D�		h̠R�<�$rE�x}+��Ho�$�7�	��Ɉ���d�Δ���e�XNE'Ƿ7QC���"u'm�w�31C�P>��C�)�wM��w�����������21}i��P?�(L	�Ki���h�W�P@��~_����[��=��`����BN��3��L��tSQ�����v�qМЩs�q�l��٪	�<�&���uö^�%k^	7��P�d�P3��\�*���
]�65$uE���@Ãv�0E�ʎH8��#��LRnґ�5���OJ2 I��)�ި�
�\r`2L��� ��G��Iz��ޯ�xM9�1���ʁ�^�RT׀w`{����\�V�gVy÷l�_M1��W�_蕕��y��@oHygc��48bg!�$�)S�U���'�����?�e�!t:<� Y�W4O؎:���s��3n���$���T�e���Ϊd��(�L7��OQ�m�g>��"��P!��N�F'#y�Y�FX�E2Ǥ���\�w�(����������SԤq�s.yOP7��k�4�(]\n7v֟�z<*�^�����B�ZA�8��.tnC��v6d7!��~�7��R?^ ;	���Rk�h|�_��/Plm�Rq����M�M���ɂ��Kduڏ�(3�!)<^#�ż1���H��t0��fd�ƛ]]K��Xb�ٮ�)��g-Q@*s�J玎�V)��i��<��l���BH�I~��dSO��3bw��qȤ��f2K�U��U�*��pKh0�n��o5�3X�yD�D�Y�,�n��<М,D�g�7k<��64+�i `��R<}�:��^�]2#�5tP���P%�|��WOɬ��+��BE���]j���j@-�o!'d]���b�b�8  �v?ƿA-R 9����J������ّ�OWm̾��n�ӎ���6�U��2+��LG�4�L&py*���A�d_����Y��H/�V�+G�FuvMP�Қ:W~��j��j����_O�^ @�&��[{�ړ�$���$��M��\HW��Ͽ_�m���\����n����Y��^P>F�i�F�� ��l�p�Q�]���a�	����r:�ZӚ�'q$���l�kޛ0��]�����@J�ze�C��b�0U�:��px������9�ö��o��;��nx�ڥ;l�	�\�Y|g]����;)%��a]���c�;��9�l�M9�""ic�}�+%J1��ؤC�Ⴀ��Gi��Q�Ԡ�{��x��_��I��+���V��e ��h��.�[�C	,�ۂ���]=��l�y��?�Wa[�^��etU0�s��5��#(˨urVN�O)��؋�m
�����[kFR(S=X<nG[���j��	^<7$MY2_����S����-��8��"�[M�#����>���������)6+��0����<lSx}���|@Q��{�&�'F���GJ��^9a�XH�/�W�P�W@����[��pj>@# �/�F�=��@����r?o�x�!T�Z&0JY�L�<�J��NEbN�j�STMԼ��T�ͪޏ���؈8���	��Q��:�B�ON�|XP����u�&>�^^>1��'~�}��#D�ߑF�NsT�<��||��Mcx���+H<}�@��]Zy��c���x�6k�?e�>bv�M�W,⩀���<)lT��sS ��rZ�B�����;����l!D��nTj�Y����3��/\"�����gX��5�:_�q�C�
����uп��4����o�K;�e����m��l�'�S[�oŠ��!�}���Y��w|U43�><ŷl�H|@�'&)�"��f�_�B4�-B`�5�zF��9�ۤ�_R+Ү��пa�TEx}9eu�ɦB�SV@Gj�����ߋ�M�-#�<
-ճ�x>��Ud1-*j5�$�!���KS�9����E/�7f[��G!ޗQ�A�_��a�'����Ye�T��Ui\ M^]��;Ȑ�D���!����N^��+ܙ�2<e\@ܼ��S��"5�pA��Y}�ǻ+� ��K`�5T��4V����c�5�m['\�Q|��܍����R {x��x��]�P҃�\�BN�t�eh�/WDE�W�6"U��#��4 �5��~�.��ђ`��ִYLS�X��L�m��w��<	��_*��(��?�!+"�l�\%�×���@b�N��l>��	��15�L��5�r�	^��{X�\�c`�Pd�B�	HkP���Ȃ�0�|!�^�ߊ�̉`�V�-)s`�Q�	C�<*��'���4���ީKj$��Z��P��7]��/󮷆����bC���C����ll4i	 ����!p�D��آ>\g����5w��\;u�*��9x1��}��4���Y2'�|8��zO��+��'����oAVT�����0�c[�œ��rN8��M�T����2��Ƒ���v���ģ��%��Ar%̷���R�m��h�L�Is�P`ܣ���(�pK��:���1��'GN�AW�NQ�{�LU���\;tE�g��h,��~��f�I�h���x\9Dv�<$���lҟ+x1i�l��v���7�G���-��ָe�����t3�/����p5�P�cvΏIS�s/0�� �F�n�My�@W2^0�0�6.u�y�#��	��wqd6��:#�/� �`p��Z����#0R<s���L�6����'� ��q�}(��iez�����y��!R*}3�X6���cX_οk6Q�~G��IF�	]�gm�S%���K���wČ��O��=�T��@ ~�Y�xz����3��JSO����oz��:lN�㔍^Z�C��:����6У�sS��r�����R|E�b�L��P
#���9&ד}�p�+c>dN�m%<N~�@����z,HZ�$�涉�t��^�	�G��O-��SN H���X�;�e�G�@��A�Q��e�ߍ�*v:�m���*�ڣ���0B3|4~o��r �����jʛ��cܮR�y�n<��������xK)�
��	`:�)̺u�OU�wu�o�W��E�3�s�2�J^d��2�36r��_��hzعc��D�w��`��4Y'v���#��-�v��啕lj��6�*�t���RS����ĴI8���U�c~X�'h�rH����<G%S�Ca$��p�<�LOJ!.G�[M��$��~�%�� Q)��+;��I�̠���\�[��e�_~+��1���fu_b�,����u�uv����?[�Ê�и-[Lp(h�7��c��f���J�9�9 ��~#ue��b=4 ��G�
:P��+;37oD��@��H>�!ܱ]s;Ni
�r�� 1bp��(	JO�]�'{�I̩�HI$�r��	�	�T�/��<lڎQ��e�FBGԃ$Iۣ����
�8@����^�g�T����/n�qa�i��Y�����(����i��0�b�0X����������c��y��#J��`�61 ��q��'˟ɵ��pӁ�zV0���A�S���8(�����G�w��2$/;yc2-N��F�[�{�T��e��,����|�_�W���I;�V�g�bDj1A�m`���P��á��t{>�������1[��`{c͋ ���$�k�Z�͊�κ�h����|�N$,;�W����~���~��6����ɯ���p�Ӿ��,�����s����v���(���>쉍u,�o���GC���aMJ���z�O�O��!F>�l��`��q8&�>Z�z>�`n�%��PdOo�L3���I�x��4��\���D���nJ%]�F��\�l��pNT�o�<`/A6xv��q�)cb4u �vG����[,����.���F�;?��M���R��\Z�F�Dy���M�3�_8���ͽ2�؇q)��M׏��:A���^c���'3!	P� #��������j֭m��k}/2v\Od!ی9�e� ����p��� �6b����[	� ���&�1UqH��6	�L�h߱�`e��!�PF�9�Aq��p��^r�(g �Ó�}�Kh:N*�4�X�4��t=��Ѯ�\�{b
�Gta�H�8O۱e�/�BC��8b���0�GA��},��b$��e��,'���(Ukp��x�\D�R��[<G��C̐|&Jn�h!��iS�{X���6�h��İȢ;�"|�<W���_I�_��a�.	��d[ߣ�_�P� <�֤ݺ�#&o��Ŭ���ƳVo��P�nL��X���Gi�bC]�1P�P�ݡDpr�|���u�I73����ǔԝl_E#-��dNHʣYm��r��ݚz�՞gJ�SL���iDMm�ᯟ�E\��@UR��.?.ǎ��(�OR�R&�A�q�DF
�zt��c�S�����K80�k����o�a�5����v��`�]����^S�.����l�&�{��"*
����xf�I�'B�`Ķ�m� ��?��w��d�$	$Dl��Y�po:O$�h�B�l�E!pڮ�]Ub��|����^"�Q�,)��/���&���w󠏒�:�"X\͞G�K�("[&-
UrB�BU��i�xC8�݀��jy�s=	�Wf�)�_��a ��)p����L�Sb�	g-���_��j��0���'�-�<���� �K\����jn	ͦ��hb@��p��E�����v�4>�J�''����&���@�l�*��hD�p�liy������qs�C��7�S�8�h���P>m�s}2�E&����U��:=]b�Ma���<���%��g⁚��/b���=c�f���Մ��1o}sy:]g����u�����7���)ÎFV�����L�f|���[k�����yKiէ@���	p������⤋!�8#�[b�]=���Y���+`�3P7�ǆ0FRN�l�d&�$vF}���滰��706x������{/��U���1�����?A�� =��
��)�X��a����K�L�1���#ܪ��1M��[4P�
�G��*��7c������Tw�8y*�_{9rZ=����M<�+�nx��L��L�/�L��?�?!V����;�'[5��N/��r��0䎱���Bƪ�%.�.j~Rϒr����[u�ӥ��R�E(��мhu�'w0��a�Z�A���o3�"�J|ߒ�.OZg��u#�|��� f�1��و�� ��{�K8��Fn_���W�i(�<W���\�U�(ls�|�j V�����v����nɏp*��(��(��I�v� _�1�M~>D}`�Gwʮ��W�<�}���ŝxK8���q���^��m�}�쾙c�2���Aa"��J#����OC�o2m�¢p�Ӛ�{��{�x?�i��^��_���OWnl�,t��T~j��[2���n�Nx��!J��TY��j��q�~����$�����$��W�4��馡�1D�y�ȶM`�Awl$zإ��-ϟs�\�6;�cjk��W��^��D�GV�0�T�nL��ǰB�8�׷T����0Ԥ�����#YU5e�S*�n��s�?�J����	�~Li+�pK[�E\xז��-fշ�4œ�&�)[T/��$CeJ�X�vþ[a\<T	o���xT�.���Y���n�]��-�5bj����ύ�f���g ���q������{Խ�^�,B@��L��<��9]���)Bv�KrP��"Ta���AgQ-�Z�ם�[��e7�v��t���C��<$E�4&���1���̠J��)N���O�ZP},A��Ftz�UGu�tR�`4�0�Y2m+��o�o4eiV��xLm������kv�h�{��=y�$���w�O=2��s(�o)��������p阮P�?�η�W+~ɴ߅¡Pܮ��p��!=��B��r�ǔ7l�P�h��3H!`:�p@�������ȡ$DB{��#���*`ڕFk�YP�ځ �:[�a��wT\����m�����m�'�ɻ��!��]�d�l�`�y<I �B_X��w^8�e�bз>�/��d�:.��L\��]��r)�8P· ���B�7�D�~��]�8�u�G�O��^ݲ {E1��z8�� �dj�t�xx���nZ�qԄ��zL0Ǜ�V�a�(@�,
s�8�~�M���q��Y���jB�~�ca��x��mR4��V��HutV��.W���!�OV�:��iЌ=�2��@2I|���,���",���5���^Y�D��5
.��}1��q�j�.��FՒ���Ə�P�!�K��4I�D��$(�~^�ަ��~��l� �%�
����.����f�A^�����|
�|Ϩ *��.	QF�����|�_�=@&:�g�E��"���h� �j&��r�ռ����2�Z�����M4n����Hs�<���Y:�+_�<Qs�~xƮc�l����ؖ���r��D�q<:To�읺�f���Hv�%�e�<�y�#�3�����)�iK��ՆH��
g֣��-jhL �jc��I�سV��o���?�㑨B�3�F{��̵�Q���9״��v��B9F�YW������X��X�|wj�>�ւl)�V�+8�O�?X�.E8:��;'���i���������H����n0M|-��e�r6�N~G�����6�>��{�}�w[��9��K,�Y���%hi=v"x�J������LL��<]��~)҅:�$�D<hDG��A�ƄS4���w�?����7J|i	.r9����J@[����q��`����C�XI�t�"2�S���pB���R�^.�uq�Z�Ϙp�L纅;�0�$�N �
n��S9�A�"ݺ
�����GD�#��~r�|�?׽I��4��E�ȴ� ������>�';-�������iwj��4�)
��ڜ�	���Y����G�i.D�6/o������f(�3%['_"ή5��S׷��O^�_���h5(H����	я����h%��?&j}ΰ��ʀ��W84�UU�hT1n�y�,�?�秔��Գ{y6w�1�:�B2�~���8�w�@lh��^�H��x�
�=(����YqBٝ�|KkJM-}�C�������n��Vs�H ��[^bn����L��,h��]M�����x'��F�v�3Ҍ[�F�R���k��5�Z�[��ݰ����|S�AN<Ex������į�sS˷�۟���L�#~��e@�2��}��3���t�;�3��S#����&� ���)��
6hB)���[����\ +L�U77Vخ����B��EXo� �;��'F��ɲ�3�W����t~}*��j��P�HB��s�b��t�H�)Lv���[��c��N�JI*m�u�.X�	��`S��G�J�p�T��7/F?�lE��^�;Y�M�MQ<�&+V�#��%%��,�ob8�2��E��#��o�!
$�q���y�����܏�>
r՛���$��P6��}���,n�o��dN8���4�J�J@>.�gmZY=4�kf�Kr�ULp����ۋ"B+�3��1XS
m��Lr��R��>'�eų��E���k(�I&��P�:�4�-�;�|�p,G����K��L�glsL�.��Q�H3���+�� ���E���N��߽m�m0>�e��>�1�� D4��3S��?��u�p�O��NQ��@� ��	������=�mJ J��T�z���񆰥*$��͝�O�����5�
�c�0�<vz���c^�[赀��gb����?����[�> &u�K��7�j����2���'���5�K�n�4?J�fǟ7���Ā
"�Nc}=�|�Ac�#�4�|�F(��`B�Pz����*��sa�&fĂ������W�[���#A��ّ��U�7��p���!l�w|;�j��=���v��c��m�lMŷ��;e'K�a4���I-��_E"��s�j���:����;�Q��ay�fA;
�
h�O�o�9�0FSZM����%󷲒1[�i?Ȯ�zqy�X�k�S|Y������W��Z�S�'Ė�i�	.$4W��F������$HnY����1�06���>�;�e���X��j�~
?�5��~�uc�x�3K�w���o��{
���(���ڌ���.]fġ�'+�����@���/M��� {c��qL������n���zDq�<6H���F0�"MqD��W;�zRjM�0p ����;lL�zG�·f�k����`{��N�ud���ϼ��Vc/�8j�7���Ʀێ�Iր�4Z�~Jh=�=��k
����[>s� ^UerА��"����!�3�Vr�K�Kh1�]�U6��t��z)(����
nbQ���ɡ �{��nV�5Hv�\a0��},^�P���x�|z�psF��ڌfS�����M�Uݔ8�O��7}�%���54�ϽJD�p���W�6���;������E�c@bףQڃ�B�
%+�٠�{��^y6��&6�n�q%7H�����si�N�X�'*z���Z�ɦ��v�4y��PcV`aѼ�E��5��� ��׺P�Ma��]�U^������լ�mW/���8j��B�6?�UReMa���o�5EQ��fyK�J�XW��6x�XS��9�oĽ����j&�;"��_%	
n1U~�=�:��t*ak%i3F��;f��?H*P�6_>4ç����f�mY=��T��� �LDB�+������l�.Mt����}�dߎW_���#e��PC~X��ou%GN')��(XgkK�$9�4��� G�C����pGu&U e)x�}UɌ~ܢp�c�e@t���}0��:���&Z�A]�=1	|��d�8�V��8�1���\1���ϥ����D�P��'BZR��5Md�]t�������.w�RJj纶[Q�X7ͥ�T��y�g�ꓙ���!�J"$���Fx�Zv��f��;�����������U���� !��6��;-�۵o1�J�֙���BĄ��Q��V��߻!�J����5uϳ�c��J�b)�+�g�:"��I��Š]��*;�F�#[�	?u�����Y�e����Ka��:\�S��1�t��
~�_����i�i�@�������:��2X�w#8���\Ԝ���gΌ����ʁF2Zِ�h��ZÌ���Z7 �dM���m������s*���<��VA�qL�]�9b�����	�������W����2�[+�Ԟ�-�IN`�K��1ZaM,�����h38��+�Eh�mmzQ�E�"F�T�X��ձN6�#�ZQ?	>Sl�)�ҝ=ֶ3]j��!F-�VU�ƹP���0@y!�c=<m'�^�q�_���r��ӊƂ�S�`���XΉ>5l���3>���ߑ��2�=$����*�4���L;���u��w)d����Ag�M��c��׮,�+�l݀ƥ �3��5�`.�[m�7W�<çS��"�EW亖	���H��2�����53�G�*� ��0�w*�`md���NUL��/詭���Web�DV����<��H��.t	?�E�x�����,e���j�l�ztN�zg�#U��5��a�@'Cm	D�V��oqj~�=2Q�_P�a��Uq�#l�=�X��c}$����k���q�U����l���v�t$�������&���¯��j���v�IG$�su�sX�/���*��z�TH�9w�@3q�$�QE S9��71W�ޥ�Z�iS��s_X6I�,Ft��\-T��5�Ej�"�>�
|�,Jo��q��,4/S���9���o:�J��B�vZr�q���0'�+X�C�Ns������_�7���."'��>�	��G:;�\�����7�9���P&�*P/P� �4l�(bЯk5��j��1L<���N]z����0x&P(�mjP#-�p����Q���/-�^1�O�����p��n����2���:)sV�G'{x��/& �������:y��5<y�&�V�'�8��&��ۃ�x3s�j}6Ӿ$ټ><������|ɜw�'ҘQ�Z����+��������{��p��F��vr����rbm�z��0:��?E-��Zѽ��&8v2�9h雪�a���v��Xq��Q���FFR`��0��]b~KP[v�B�����g�����#�~��,��ϸ+N�;�s�V����C"���������-������^�3�@��Q腰�C	����^3�n�/|L9=�
��[/�6��;U�������s�V��|,������� ��V����#�I�%���Ʈ��r��w�,��k� G
�� W>{'[5U�FB��ڳ��Z+��n������߭�F�Õ	뵑Ѥ/�S�I���.��0�l�@�g  U�xv��"��5�*�8�A�72kr��jnr����PW�3�Lt/�z�C;���B��lQ� jV-6�(�gba#[�0��6�>�6W���E���B^�4n�R�������!F@�ͽ��֣~7�ڡ*[@&LR�כ ���Du�z��^��_1r���nu��S�����Y�w^0O�:x����-���Q��\Zn`�GQ��o#�r}��� ǒ���z��l&�eI.�"���jX��Ą�,�f�*��A�/�����V�����噾�'�UP#�k�F\u|��"�8�g��D�'�ogF����S�l��)�Y�kX��j�8��,��1�~X���/�c�wgs.8U�e�U ���<Jj���K����SN9���Z3V�_�B"���#>eW���Yk�2���ԒK)A\%��<�/�N�h������ؘmb[���(/'�϶<b���E���D܁6Ʀ`J��Eq�>UɻB�=��Z�����kϙ\{YQr�WN2�� Z��A�=�Y)GzǛL�N�Ӄ��V�>������,h|ݧ�k�����V�'�ّ֙���w���;w�i�{��"F�v=�To�41�!�dIK�,�C�8��o!K�{J�c��0-.b�5	��S�-�X��;�}�)m�����ݷ�v��ܣ���\�5�i<5ڬ�G�e8x/�,@f�l�@*|�||�d�+!�|�b��3{���vO���$�h[ҟ�P�7=ϔ�+r������ ����=2�%��l�Y:w�v���6)� ��\��#�7l,���M�Z]�)��	6�O0������D�^χ4f|A|"�jӎ��|�.w�߾�G��O�y��.�޶�vu�?i���]l��������rU��򽗶��g:��BA�:� $t���K1�o������Mmߗu�7*��ژ+��x���;��qFq�x��͓�ew|BHͩ9�F-]y{���S��#�F���h�Uk3��PX�d�r`{a'�i�d��eC��d�t	�j�_��Zv컥hK����f3Z�5���co�mN��F����yQ#�;˰�)��Mu(�t��S��wͧ����ӵ�X�&�]�,�E���;��pF���/�E`��T`1���ƳI�킍U����3<�N��I�@*J�$u����e�����)�:�����_�y��ӂzU�w{�#
 ���b4�6{Ɯ�O���ۀe�p��2łnY,Ixq�|Y�J��vg���=c����Uj����"B�z;�wpz��<���ť� ~�3��u<U�}�ל��l��L0Y1a���ZjM�c"��ǝ��h��(��lHBd��2z�+@��ր���EN�ëM�2L4�t0���؃����iڄ�^Ŵ~�A��ŭ+^C�MC���X�|��wB�'��to?�N8���8���������O��f���p���I����N,�QM���>�^��;��"d�g�䰥l�D09���`7Oo߄�w��%���n�g>0(0c�fMĮ	bH��RC�T@r��{���*~pr�+*��r)�x��jg�nM�t؈i�H�cWO��K�bw�#�*�&EkR�߽R��
ӯ(�N8.���oaa��pN�	T����~;>�/����9�?A��%��B�+0-x0�Y��3�
����4}���(�fH���%���!-Ϙ�8)x�n�ð�� �si��WC��r�7c��%�a�}��WI�=�ݤU��WI�[�a�70"Đ3
�2k"� �\�D�5��Mr�'���z�����C{h�(���Bx�D���d�Bo�&�Tw�my� 6�;1(��1�Y#(s���Y=0�a�xn(#������=��xl񋘿��E�s�pQ\�i�����f�k}��z���Կ�)�������N�a>�B���Y]Q�Se�D�pvĬ���17��[�E2Q,�.�rcy��1��֫,m��(����"4xd{9O��Z��������}�(KJWY9\�d�g���� �?�M�ֈ���������� )�N<�����jH�����(\#%u�«���6ؽ���&m9I|c?`�1e�����`��	�;WJ�wq�:��EQ���q1��[+.�jWy5A�k�-OM\\�&Ϗ�d3s���f����ı���.�\ni0�ya���h��|b��_^�g�5(��[�Xc�E|$�ap�w
o|�>����|4R�Utՙr/��;��g�	��k
T9��T�r[_f1���>��]*��O�LQ����"T�
�NsN8H�J�vK�b�Z��j zQ�G�:�:��]�zx���m9��P��V��^l}רpB�=8��`Eex���+J��+p{V�ڲe�d���WDT�w����G���(�Kʫ1��@���k'�腠�d�bN ��m�P�8�?�4��Z�3�~!��_��W*�D�T�PZt��2�N��+��(?'E�\e&X����v��L��ܑT,L�v��I>�i�ͪqf��Jd�=���]��4�A�d����w=sx1?���HQ�q}&qD�z���Rh�Z%	`�{A�%�`P��;��_��⤛^:��^�K����0��Z�p�1$c~��Z�wiqS�=�H��o��s��|��1� �3�̜_��Ƽ�hp���&I����8fM��2��=L'�W��g�+^�@�$�'���u�������'��m����] �،�BB,?��
�I|7<5䄝���s��[43E�Ҙ���D?߅�3bQ�Å=�ǰ���I�8�A����d1�2r7�D�<��Q[fC�s��MQj�ҽ����*�n3�<�4F9�')ֽ��OUp��� �n�_Kˀ橦W������N���^d߶m�S	�̤����dxi7��_�z�{���}�=�g��a�՛"��X�|`�_�JW��=)N�����>�d��[��_to&���A�J�@T(�b�'E�Hǝ=Eܜ�+{xj����S`�e��Ae��F�~����/��)�o�N��J'<=8���k��llV���Y5}���mHp��T���n�F���~V
�ܞ����AR�V��}�a���pl�