`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
qyebNVje4eZUP7kvnGUaiY6/k1hSK7SS3mOjazPRi51vpVPf89uk88kkRK66ROSEHnnBFC+qdHox
UOvc2pRLQO32Yui5KGY0dKXOf+3aYV+AF0Hsv35S11alduFy/u/VBJvENRsuJb5W5u9qIK0yqDij
dJCYKFXIafPY3rYNBpiJn640SmDpo7ba17a++qT7LSgbGUeRObanQYcf+Q3dm+C7CPRLkT0WZuPJ
KaW6XriiZ/m1BHIJMqJqtfmAkR8LiT95Tml+XQBrsjvKuQajVw5fnSkavi6umVKEu8+XTKbj/s3+
tgdJbvdhxXyzqDeCgvt9LT+r6s35ZoI+ZCuemJqNyrCCbDTcUjfnh6QsbdvejJd/e1BzW2nirixX
OkttxNwSbs3UOv5PJjrn9IHP2JIwNOHC8z4hYN2KOEVzyDAGjxLV6aSBkW4gMqOirjciSDtSncK2
J1ASYeO0mHTuhRSP5hal2xxDQiBPseajhWjTgHhS2jfsh8LEX/yFhBChWMIHH0y/ecT4cilqGOBv
W9w48KyWAoK/iDN0+e1NQ65Ty22XoB/F9/db5xjANryfNe13YCwxCa2p7UwQdiF3/A7idzzAUGMl
H5tCvent8XVk93DCKkIzUBJmnuIhuy27GDp/HzEo606cFCmb864uZZxpZ6yLJ2irCTuBRCgn01Dr
UlLT2CRIoaM/eWCTAx3niCd5rYiI7W+saumPYmgqP18XmO7By6eXrFVX5XQkoKwNgClta5Rcbglq
t9ZfZgoxDE7Q+w4nhOQu1juzgHT1iIE4bBPsyg+7DZWsphmHn7jg4utJzrnN8Fbr3hGDlFCAqmb7
oeop0O0+bHdOD8PwIOL1f+5FJjXrb6dI+a3SCTvcJxKcaIIqKZojxuvjgzAipNhXTpkjmP/6I/ra
C/EBIlGxM3gM+e+3jEM9gSqjvLWs3UT33gQly3jFfCp18RMmJffWF/VuWJsd/C39Vg21HJn4BIVl
d+RipHdidD+ggY39XjBP8L4DFADk80iSpZWTPV+Aevhkhe1BrmID2IKs5f7kWxINsHH8XA+cbIHn
5VJbA2Ojn9RGxolppi8jOHlukziZUfwDGe8s8TuKHu/E4+hcVaqle1rsJtpRoMQDG4BUW+XXBCeu
FZ4XKhmcInAHiHITgo2LPPPBz8Bn5GCBVrrlm324c8Hc2dVYnbDzFe1G5M+oZ/sNJ4etH45NG3OS
DPCBUaS+NzkH3iYtG2wZQVAv/1012+0Il64IGO8QAnnneFsMb1mvoeHr4zTfrGVkHVYYC8IVYGMA
07PF6SWpcxv9eIHCR12cuEAUsnPbv0G+b/L0DJ4ShC4vbN34xqXIVXvcb3zhNf4oA1mpmn0LL8Oc
HIbmky1nw9QFuS9i4+DMjnNffzugZoH9aWh/QNFKpcq/+DRFuCIFEzsq3eASrBWV/RD/o/dNfyII
4sa7m5Cvs9l/gTNBU0DHGEYO9aGsnU5zkNvwV3xlrXJjIIHO5MMaeVEt/pOVykcAlO3eBEyby/hX
oiyPS+rEV7GFQhvbD2aFbb0J85Dn5AetbP7mnDdCa7WYjqc+ITArlk8+2VFkV0GrdDx65+VIX6wp
Xyh6CAmTEKYxvX5MtBpvnHgRADF+c+Ri6rtJJnAOZBL9wdxcHS0MgqMCNQ9pffav/dbvZzQKmVfJ
c1lQCc9TgxR+czX7C4EPyN5WuCj2oU/newrEEvMvR9CAb13uQwy+jwWoEy4h7yptfi39NbU1kvfb
ITMugxPL1PR203Lx7V+oj5ZJDaksTESjDeXc+G91VZQpvgG5qaL+DlWcbW9K1OccHWeiuh5qrrIy
X8nTmcdzuaQWIITgD6sLSv4Vk82jrHx+33/y35OlTUWW1BdXe1GcwoDBnqzhXgtt1o4pSGJrF9wF
qIcJOqU9Br+SnRfqfcTLoO9XoloPeaqgZWL3jZbB0//IZ4a9Yy8FbYeixRatpDWTqmna6bUarboK
VOoR0Z/AZ4VsIfTl3u7O4SGhaFD/PeiBqtjEoYKKlNBplXEFngV2DdP/E2DLNfLh146x4LiNLAVO
ES6RMF+W9mSBKNm6pg0syjQz1NKJMk+89IKrQZRyAmkaExziJERG4wr3K3pJRVQ9icSR9fLOlHrf
2PGTx06HUjXvC5mtSwr642aMGFRHr1XAjOx1JdWR4Xsa9XJc8yBmp0fiCe3lCghs85jV/FyvJ66c
A2C+W00guCHVbPENGrx3qObfyhDk7B7YdZWO4NlijpuwIdOiXFka2QV1jWNbVjyGVmmxijQPFxgO
cd8uvrcgkNu42bXoWCOTyMNVasUbw99lNt/vBCHn4V+l7rEf7pEOyR59KIIlViX5OgAnpzHDEyAp
wkK+qpH7QwwKM5OqHKK1V41GAQisg51thHscJNSgcr5BYNkF4HMKKFNo83JGITjZ5dorqA5fortr
BjIhG5fK88L/G9vP0O9Tjs6lyFNJ/FyeYlAPTnyJUBZ3lkKTMXqxwu/CxBbrsxxjuYa0C5wP22fL
BbucXpBhJe3fdWjbnH5m/ziS7vdjSYz/KCgzuQN8UyM/py6qhjMIbdbOVGb0LQWmBuLIAGeGrav6
UJ4TBrDcv61fa8NuDv7J6+QBeel9IflK+FXQ1tgpWozIfrnjQFkax/uiceQQFMTHhl90281l3t2x
YHP0qPOyHeRbVuav7u2DlhpBq7OFUYVCOLJ+veIYRHO9qnzaaXmJntnzp0wlnrS1dZtQXALzIExk
QApAGLSz4sgYVLW1SH+fCf8Syr84hFNA9vEmZHhPS5KSE94LUfghHtUi1O9RPa3RlM/r/80kBhi8
5USmwFFKY6/S/lf4dwzz5Fq5qZtttXnqCQfAk1+i0XqNzCGeeUKo5jex8wNRn4UFd/r9UQbSRwlv
sJPIDdoHz9whPSMtgcZDQJbOY+rl3fNGDnAam10gPaV01we6fNegGobYXCtO3K39Eg+/Q0CPzSkA
LQQO3RtliOprNqt+vdxvmNWBnFFV3Zvh+iG9Hj4OjuHpTf40vnN2P0/u3ttitv40H33AwjlNNvFt
K5tA5PigblboXdHNRs+rUZLWOmVj1cBjuNvSRKa3vPoSt6H9o73oJsbygP19gfilG6tuWVSIN6mh
SiFkTcNFup3rq6ZM3CpWcdOrp5V+ArK2TPOC51thSTA48dcCrDF1azZH5XmSNCbKn6NiKli/cnlL
ZfxFbcmqeltF5viwLqlrpMXE7jOCTXIQ1EnbzYUqejmCAQlIa6H7E0Anbi6IhCLwVaR1sY45
`protect end_protected
