XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>a�'�ߚ�4�J
&ѡ�)*ὐ!X*X� �/��)���ǔZ�9YP'?���o�Ƽ\������e��βӜ��c��N�ca&���P�����$S���mj�څ5����O06g����B�����I���p���	��j�G���`82+�"�_�I����=c��.C��f[�'a�ǥ$�Ӓf�/MU*}��G�{m8%�x�&��4E�2A#�nDQhX� =0JUW�W�]��b��)_���0��	M��ǯ�C������s$�0B���G-߈�ਦ��:7�-cش�Z̎H/]my_o���.����yVL��3���v�����s�Ǘ�b��J���|kI�����R�i��XmOS�n����gQ$��d,*�y%��]ĺ��.ko�� ��@ԈE{lM�'������0�����[��	qFD$�M���oFy��_�0�3.+"5wC���>J���Q?�p/%����H���3���������n+��R��P��`�e��&r٨���Ttǟ�G9F�-���|U�9����O�ߍ-Z'Xп�b���F�r@�p�ʿ���%r���]�ͱ�'�cY�G2�Rr�Bn�K�1w����r�k�n�7�����Eb���:�`i-�y�cG���C�&�����*�L��]1M�)�	���p~�kT%�A��7_�zTܱ٪G�d�ET���-���G���ҋJ�ԝ��1���&Lڣ�8(��}�m�VǀB�[z0^��XlxVHYEB     400     1904Nv�����DqGJ��(���rKy�Z&o	�C�lT��Xc�����|i���p"�X��(`�t�o�����=��g�$eӧ�:�eb�saE�VT�Ό�)�8zlȴm�}5Di�B�®��82����Hv�� ���x��O�S�Q�p��m�$��%��[[x��풋4.J�`�����@|Ǐs�n���g;f����f��� ���ˈ�rS�*�%��]:��ѱ��N�bnY���;�q6�x.�Ğ@Y�^vwR����Ʋ��:K=�V���qC�
5]�8��5��g�rއv��2Ъ�CqmpH�͌xG>��Š�/g��8���pyl� ����~�o�eTj����
�R�^��!I�R������iXw���&�x|D�XlxVHYEB     400     170=C?�Ȕ>�ۡ��okHO�%*�ݗ��{�LJ�Z���QTv��߳m�ژ1���N�	�'�6�j8�	H^J�X���d��}��B�����K|`�����v��L
>�sk0�6:ca�[���ZD`�HL��� O���F�^)�H���a6ɚ�]�`��3�\!w�=�c	�_.W��xS��Ws�P�x�Nr�Z��$�yIF���z	),���'V�l�w���G4���ț��e�����Gk�Rc`�H՗�o+ ����x9F24�������'��R���6�ش�v͚M�����u�ȓ�{G���0@Ck�@\9е�#���{���a�q��]�� �����XlxVHYEB     400     180�'�O��Ulܓ�L�HZ\�$U��ív�Inꑓn��2A�C�K-��|��,�؜.�A(,�B����X�S8�1�	�4���:���Nl�;����?zM�[�_����Z���F�o�Z���0��*��Rvf:��*e�E��x������5�d$Agӷ�+�ĵBD1۫2e0*'a��ַȓ�W�^O�^�D/�5ݿ��zP	�.�"�V��k��Yӕ������D���1�;��1K��7���G�O���WPG�:�96�h���E@�2nЗ�����8م|�q��a�����\Zi�#ƒ�ޠF$c�:�����nfc�8�*�$��-pk���c���sΦ1�ڂ�mm�%9XlxVHYEB     400     150�.�ղ�i_��3!����<�-i[}]�X�Il1�	�G�y����OF��0���C��d��Yc�N������(�"��e��K�w#B�p�PUYy����*C1��4Sd����V�-�a����!Kwj#�w����
���h�A�X�A��y��e�+���
[E�,��+�\
�)�4�[�Lu���dGD���xo�gb�}�]�}@�1>ksЯ!#7�����_q�M��,!��a�G[�5�R��(x��-nq�,YX���I��V@p���T�R[ ��f�`��%�֜?����i[���%�P����^�4gj�D�8?[���?bXlxVHYEB     400     170@��>��-�M>ʱ���T�)�.T� @̎��pb��|���3�/<���=��C����:���	��2���'?ĭ��t���#UO��S��{^Ȗ�lI��#?.[��dk��^�6BKG+����8T�mX(�M�F\�S��ҥ�=c�>d�^e� H7A��2���B7 ��ף�	�<��#ݳ���zFqp�AQ��L�r����47N�	oeIg>���t�5�7��t���?��e&�֘[3&8x`����7
o��K-��������"����������
��9K���αV�LQ��E����L�n�_D��aND^�s���*�W�iC��"&�p�+������!7W�oҚ���XlxVHYEB     400     1b0hkS�h�6���1����GnYkó���{D���� �b�_c���AF��q��+OV^�De]:��n�'�6��l����d���##=��p1�O��i��Qr��.$t��uS�e�أ݊��� 6f�	��������^�K��M&|i������<)� D�75ϣ4�[-�����F�(,��I+ܑ���ӡ`ݼ�!nq�+`d����btiF�҅�xÎ䂞����GI0���n��Y�¢my�)]G���.yU���K��`��i�@��4�
RV��/�#��<< ֟�jv^:�7N�ұ�fƷ�9��G6���|�=������x������Ŕ�4�R.�,r�3�Q ��⯒m6�`�I�����(��X��hYeQ���ꞃEM_^�L�O<�3�dsrBN����[��XlxVHYEB      e0      a0�=숤��8Q+�g�v-/I�ȼ;7�ᩕBԒII^}�.���r������o8�T�<���:z�! ����<>�_a�c�y5h�ߎ:��V�Ȏ� ��܄�5�X��i4s&�d�m>��,��~��Ǩ��M��baB�3�jA�
��[>�I�y{��3xG��#�