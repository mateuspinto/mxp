`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
UzkdOxJzYewJlo4zf9sJx9P8N6J8YaVZWcHnBfOSg8WYgR0qd5dg2oCXq3LCfD/jh5nehs85A0sb
dSOzN93IlX9MHkZqSN4fOidCVp5WoaYPVo4TuiU1j3MOnp2c1w1/9OtEH9mTZZTpPAVjeAfmT4aZ
Zulytrpk/oXuPZ8oUOiawpmE9mEWvgMeMxkw+Xn7JkwdLb1Sw8SlR89aY2flsE0LiojkOZwvN/XP
NfCiF63C4tmmD4ieQIl5xsKD8Q+0HrtJcuE3HJvnPM1f4ZyLMkNL/u6htAV0gBS3sHls/jJb8LrC
VLNBHkiubrRhaniXKUix5DGB10K5OszlK3OKSvmrhjyuhQ9dRJXYgVp8p//Rm84YDSErHNQjuOrJ
dN3vXB1X0JIACGO+Am7sVMDNuBgP3wYwlyGlqNywXJkrC05Gt03ffFiQfFviN+AWjZ+luyPMALAo
g0pTk3mJmmWp1vtl9CqpLO7wjHMjQu5P0HG9GKM+nLCFdk3n4XgpQRbzkYmnVBDysOyqPu65vh8I
fpkuJtWs54saeWlbkfSrXdosd95m2vg8/G3NjAJgPET1smxHYnSQbOrX/sIDlDHoGHyl+BWpmyDf
nnAGkkdq6hgPP4tPL5kDrJ45+YbTKKc2MsTFlwrmxoK/J1cDZts5Gl/nDZelIwvzH/xJXLxv5deG
usDnkvbMcLPSn93cVr9QDlv4bOm76DOvz01+UHP4HyB0B07AfkV+FO68m2Ka9DFvBcvHFYixkJpq
DzP/Hwo6/0PTfZ1fVu8Bf9UBlJ/qNvHlWh7o9Wr3FWeXKgMwSQamILEI9fbBtD3i6KqaTgEewkxa
q21YgomV/1E3ia0rhLNuUOZ3CNTjJZ9tX6kdkExIlQvdhEnXM1ekGFOAdMCLZHBOusokaVsSHmDs
WoMCnrYfvc5ku0cY10jPAmSn0SOM251ldcvDO6hbgWbnaZYXXbfodEQHz/9M6545TdWHkrjKTERr
gIIMS3hLK3KiEKkSMSLGe0sm96ia1/n1p1ziYVIDnyWk1YqWZRtKE01DUBxEHdPsPgGBjAcrxXwN
MufQaYF43waRC56yVGdLWaGGhA9XUWgSTt1OQqF2dw4xSGbkPEnYRi8zjJDjrzn+tpa5pyKwOQHQ
Xdq67zvpfvsVj+Cow3AW3DMBNT7OpW/t2/iooGKhpTHFudGWOqrCcfrUuXSuB4zM6CpsCp2JsMEH
yDeMENprj4QKrnbSmhe3zahSt49CTtxZhLcEosqCffjlGYEIhxPW9mg+Scp9tUr0we3UPlzh0xY0
xWM5SzPoSpJn3oEqM9SB8ihdy42HEov87TvC963QX9aIUBbc7C++PP2YXwN4G20LO+s//cqJDjwd
j5dlN39b10QP46ULyoDDa9T2nj4G0R7M2BVVoEwgGsiaWlbsuNtqPt/jiVzYZWVbCDg3oNxegtEV
gmXo7rcCT7Zd7mgSmqTAASiKLz1aJrGpesIBzd3mxT5Jm04C4ascRy/AorHeaLTZX321ML5vyOJI
CGP2tCPNRenVouibqrnqA12hzc80EKPukS88NK5TS7SK74lo3VP4tmtBSEswSFcgry0iwFbtc+Fw
Pd4w/CFisLlau3sphEZELgH7wM814Omm3Fz9XqrJfwd7Jg6osHKfr+7B//1pkYcpXHrzBGxAFp9A
4KKAnsgzmGk/fxYSVBmgKS9zXgUmmLVLW12qmJ0RuVuAEflHzsT1oIy1T793JscKOhfxaQFsu+j7
imTWYnYSugaX9t5B73zH/HPFYUeiS1VvxgA56LXQo75AjTFwCAkTOTGYWo0WE+Er84sdRZlNpI4n
UN0SzXvKUioT4uW9hpFXRRZn82peK/M5wpbqxVJJ1458LkS5jRASwO9P9VIFxbjkrXSiT/RDOUbz
66CuTIj7gCrWPMQ4tIpFvUscKTYRw9i9yvt4yRLbP3fsB+/S9YmbNCtib9hBMaTyCKGKsnP1tR8q
N0KjOKcAA73lyM9xP59AGGytXuohOio6/7PzECUM2Tr6lRA2Gil1uLVGV6gOAJbOHvx/HQE6ySnT
nqyISprpB3lELG+LLm6IzQJdDfm+4dw19NN+85/q6G77Ngf2Vkj4YlCIsL6HUVw8UHo/9VF97Pra
sO52sJ4eSg4hjxQP630FtREefMMqNl+EfxilP1tb+0dC75PG6ULQ4pONYTnvr2bUzdohF1k7N2ps
h1o/Exkr2fxPMjVnYeWH25czHd2C/mlscOZ3LGYqT28gRMixCLSQU5AWf8h+tPlVLvCQifjefVY3
BT+Lw59wB+kPYqGwicFHYuDcQ0ebPVeSAkxViIGFzXnA/RhgD1HdRCoEfnN1oH02TSUqwTQ7Pf8Z
a5X7E7IqTck7mRfmRtkQ2VCHWIUFGH0MXVClbcMVYQZtf2NDXTgUwqZLPGJXi5cJhFSae2xdQv64
WJG347uH/djA47fwl/ekx7JBbWj5Kq5CtUjiFKlVVgqeySbJbDf4nabWc7Sz1XOJH8mld93a/7zQ
zjOr1J/kYvdieMsEyI9o91CPYd6I3zuP6VvkFD4q8nY7/x4y+obAzeUjMOPRH9krKXKhpe7wIRdO
kgKE7uQM/I1oJ3MaFWAjOfrDVihS+U50GDuK4SmtHOnDPLkLVvT0Kg9RkX8yuAWQcgaE11al8MYy
PGjEcrfWcQhM+RNX3gkqck+4sv+de5wW/rXxRj4YrhRBowoSB6bIuTlWjFe9MJ06hYZpNobWD02G
M/HmFTnJFOdioGQy/9xm8jvj3QCKO/WpaTsKefJvr33nVWNAVlqwqHNmQldyQZvIjXo4hy5eFRiB
j9fZeR703N7qDBUcZWSgi2Xr3ZZqE71HgygcWY7lGPBZ2Yf6v1wPpM5Xbf+wzuii6tgtKBHxN23r
TCdnpUKhSZY84F6c/GXtixQcU8FH6+YaoJ+PBO7qGITf/GG6XOKHFCdrBT1JkxeStBU6T9a/MFzI
ryWhsrpi7pSQwNPEqZxmPK17NEolE5++uOkKvLvyv6hugbb8/g0V3VGgTpDBobn8re6NoQr0HIXL
9T7BZO3GZP8GyBB6Lt5+vE232QAGAvUDLi4a8e1ZvDyMYy6B3vjW/JS7RgtiWga4127/YRqev2CU
gT0r+FSHR6+FepUesoFGp7xTlYyxSZJj+V/jE0/mhpRFq2kCq2KAfwgw/rx4pZHEZwPEQVkosGbv
W4nUAw/F8q8U+CJEoDcaNu2rP1ZV6EbjfDVAGctjmDPLBPJhfT+1RytnkjUV7O15iCR9yMSnNoyF
Wosi2+7vAxlbpiwUA/bjxuxnLfbkBw692mtorsRlMzgEgyUUWbgG6MWd7WZ0ix4r6VsBDMIk0lfK
4Ix03eVIi5jQyWTRW4SNR0UXI41/tdvDflyWXdRQRIP7LR07QZDbAirPbGfRTSva+Yc0Cg9zEJp/
lFnQBAsVFCxB/9V/M6gTqovSV6GouaQgTumE066+Eza+nn60rm0hrkPCBrkqK2WDdAzsm1j4i60K
W3ARpmEsEe4IDB+MyiDOofT+J90I/0yrPvHCLUVe1xHcnLo+11F4cuZ00Gt9G3I2JuL+qcVkL7Jm
qIHdqbOpNI0V6c70dq1illGC4G0DvBZKK3g1N2NyRMdCqWEdL2zOGMAO4ibIQDxDocKYrnC8OuoO
QDeJCeFYlQFJ6ztIJG9EXVYl1/nq5WElPhWY0PM6sr0X0DZNIU/4MzwSBTzkEUwPH5mP7FDm93Yv
JAkGMbUFnwuazoOy+MB4rbFCj9Yuu75ukmK6IlkYTibkFzUYmhky+oLyfJG+BZfZpQX6iQo+GY1N
AH7MnOONkLwunoUp9tliOH5Pe2zIjURJ08dDAmcWadjpY7luLjiwCq8dJ42eIvs7Zk+cf+60QyJz
+35URnCqhAGsvBIGP3C1ylYrU18Xp0SNYfdRYYbm6kbLhgFZ8+nJ/eVEvfsJ4hiQO+1SmLX5pm84
WT8EyJMYeZs9EhKf+trIMYEr1p4IEO3LEDnQtMhaUuZveoeSC+yFWOvQpIyhFFQvUugrgCpiIdw2
u5VelonaWmMAnd7TuSToTVydfDh831bkrpXyyRvDEN43Q6QvCXd11mR2mDsS+rahKzo0oAjeYC4s
plCsSS+03njRpbSQz4At0LoWk4UqW6JYxXvhTp8ZiH/EpDrCMlN9Viea4ZmjEdakLMf5zCdVxwdL
XF4+w2Q+HRVy8dCqBmZ/c5aIzmPjXaNoUFHhxx4wayyku3SNoyImrVqpd06dJ7DnatARoEVkaSJV
kXYTttzQ2yUkAUm0QDt2Ld7dn4md68qvKOFT25IAUrbXqiwEAQOeUparBzDwe204CK4F6zGZp7Cy
xgPVgpgREeFb/KmIIB+lLmJDwiFcDgoPxcUgAuMfKOC6WB9uGcz465kIFzqHKqIzYeDGgwM9FyGr
yHvp2/UqefXxJe1UuuYDuQ8vtHzeYOVd8Twpsv4Y7zUcwPgFFtvC1qvR9UJUsFmocVsvJAyHwZrO
znNLK9BdpgjA0ey9bJrc91D79ySi4zPwai9ebbedPHDTxPKOjLiNVfKPmb1ouDh/aZoo09ErsLfH
9jPXqXTOdc13bS3n/8qbAXNrmtEojvwW+cklFs9pUqbpiS81r0KhPwO1yD+u15CUwHYjYIB+9jJO
LOykBW/1FQWFlvz35b1FPU7lxsZYXdc1y5ratem8tGa1FRBBj4hmY82WiZsaXZpEbwtozvtYB0ww
jt54+KqyiMOXts0VFG/oKACm+yCDNKbXbFsAAELjTdy6q6Jtx15GpamuwHUK9s4YCPpAKvshyiJ3
/2gEbH+Of0ynVCdslX3xT0+6NttFSkqFwpgTMfl9wLt+8UEzeuamXyO102bC9+YjyjXnh4hNoQUD
x6k/SikPW2/uaXPHG4NaxKEx7zsbSJtVaRbcCTya3jutbDf6T6f8+VM9Sz3GZ+EeT8RotMicsqep
7869MDVhOwAofEqT3lewu+84vTHaaUkyooNWlFozTdHLccdGv8229OGdIrIvV6SPEA1qRVq+crUt
NDjnw8AMdlA+ROJZPUPV063CVlUmty69QR5gstC9sy5lyHD6n9cSbTeOEy+Rw0pLjncSw+VitLW5
UFuPJkA8Z10lY66ZtU97JQmkY/bv
`protect end_protected
