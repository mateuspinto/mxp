`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PbVQoWD+pN27mQ1tjKbwlJaSn7DbFJfjk5sksJlnHArxxzPjBMtGKI+lSBmLN9srdyOzDeCS2J9g
yOKKC3/jXLSic7HCH9t36FIU2AUkoAJGolQuExvLyfObV8x97a2Ofr6McEQp6u3dYhcxBRk0K+el
62UbYnlrHgYV+LRWRPRGHsdNSwYyh8aPRQOwBKmzyQk4ZJaAtfvvGgg2oxbIbGvBZAwjqMbyCrn1
wmhhi79KdXk4fO6c69TAcX7MxbbEbt2yRHLfo1a6q5yYC16TFEUsp+E7Abm2cGiWN/jkF39Yg70P
+Rnyi+FfX17k+2x1OqBXlzw70u7zGwd3i8ydFg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="LxoDx+IGH/SjxUXlWzLe4+UTfHH4Q3cj2QxJBWhJyBE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
jZXMihkHvya3v5Aee3bgHto1/3airJPH2GrYob+cFcNLTXvOprTJldGWvGIIkmxrJ9u1OframGab
GbPUqIJOIasnNy5YvXdWVb5btTMRMpbMT9uh/r7EanmwyAZsOe4MGM46oKLN4GWHlq0pbJtnAJ9c
//tIpIyZdJqeCgdlcpVaUqbeLFQCkt2qJFqgQGLTZ86+H4yYwg1oxXPbVTmczZlRI84mmjC5aocl
KTd7lm/D/SXsugtoAudZtMZ5p4JBl1fN7ksHFhmPQ2hnwSjQaG8mNbYVcsWgoSndzv1LoKiNljvc
0lnZ/2xHPhTlq3TsSRgokvLI7x1oik6J47hllMyy6/VUEnbzL5aBr7jw3sPG6MdAg4HlYJVsAkKv
B9r3tcq+uBsQILhW5Lu2g3ClMOuWGP2G7cYZooxUvaee3aBivhl17QF5o5D811+CQ6o/geWpjZlB
t7N2udpBvRaVUNEpX/G7v4g5ZuBRSSrWEIT7PNKcUk9sshF0wUUu2zi76O7JE3HwxlOZOFgP4yXl
mpeOHYkF63fSV1NCdt89AvelumIthM9R4O6SP7PG2xbwftnUyW6gJHpLOvrDsr8KyK0S+ABSmYVk
osUVIIZFlZPggky9H2hjBskAtQ6sB6eP3j7FL8KYJi+6+gOFFMErj2Ok0aYLbbZaR0oIo7VCwogN
UT0c6gV4zJw+a1+JC/qc7IkaDtDZtCY8oRSo+JUwvxAYQHI5lbg61zDsbqS1/ZtOWYGp9pSLAOsh
s0jpEbt6dcO0rnaEhMOyn8YWqQrYgpb2TSCa5NxcdKQdE5N7dPKLNADzjY2quDFskTn+Oov6Mj48
7LsPeFUP9nQR57n7yiy1UDYsbTUTU3pMozwx++gZLAwCZQ+rhFwKzXzxuJ3F6DHnZZWrrCxUnr+v
qN1DX7NjgqqiuEP+75GLC/hNajrSF9hYNjMbz2tf9u1x46KqawsCls+gDGrFv2AVRxBbYiod1Nzp
66bU9/ok9FgOsX5H8FALWi2PLeLjR+5fDEExjlpcbYgm45NXas8MWLNbE2wvGmRgtKw+kPOmeD9x
IOdTf0Y9ARa4MFFSQO9Nv9LzFS+iyCn6QP2Ca70B9WXC5pGsa1ZfJ8G2ys64tziV29baC8NhLhbh
zMrbwhjTrXo074UvG2EI660G0YuOGmQ5kg0mPLbPmWZhLqM4LAknUlej0Kv82NeSiXBmLnB3uLVd
WtN0OSYIvVAW7u2ThYe98WvSmQXHVqXRpOjQIXnBorLujWXCH/dFedWZYLggXLv9hEjIl+JeN6ts
2hAe04BRgGA6Bz332Qqiiab9GEXNH1MxPbLXPFt2RtiidxmoHcZcwL02ukj6Lp+lBE3gPKrpGti/
2NDSflkFijdQRK6I895QOik2MPpUVRB+2SPfekQ2RD1tplVlwEWjX6LY1UdflLwo4Scn03f6lECL
DbzYKiCfeBIF4vT04cfgPqNSpd3UxNukTdtRBnSrFMjvhrhzWTnJy2axxPlY2ng1YuFsuXlajXWc
0W1XVldvlcpBz9JG9++lr3P19+0g9TFsC9xVYx+VJR6ozjxK/ud6Q1cJfucTXYt1cAOoiy9Pjv3q
ZDIp1I4rCvWsdIZjhbB5gDtlSlz2cBqwjF2xOqYjVO9e3jlLxNkpqf/VmZqLf5Zz4U+xdm6cGMaV
SK1osqJ4jTzZJZrnm32IrtkWUS9lJZWWHcKzPL0AsiomAecxHZbrejvIolrsF6mfstp4w1RVyoai
kG+hHpm67Q1BI8nlRkrj0IBLi5B1Hp8H+S3pO7yZv7ZnjnWuCmMk1Lq7wl6IDKs97LIGdGPrsBP9
5TKgIa42Rd6aHOd8TDTWD7+OW4pcMQFX7Qj/pSVnD/MMl07OVxQ3vzcfEvcnzz22Lx754ILKQVaa
QfOTAXXyXyQ9f9Vv9K/NfXc3/z4dmWEbu5Wek79wRi6DkNLbsMdQEw7NDEJgBvucZczdIk3vCDlM
YU+URLMgTFcloo2B8fR0b9/W8ctsD4TRusrZMZ1YKyIcj9VcbgK3Tmcqe2QOjcOHUmq/Sab2yc2p
vQXrvzENnndb4ZSLTPoN4Fayn2Q+iV87ple9dZimbrdla7ous86+D47YvsvJqYFMlxT37iuEOY9J
SbWXgGTkOtgmOnFPTft+WB++/uzJcQsr0WnGDSFdqSI53UR0Fj8RKo5GrtMxsN4v6znRXZDSEva9
IQ3Ekk3ott+VdXKUYtlgsG29WOVSO1safc+pAgKtdcIdv9C0SWP4ZA/wYCe1ez2zD1qPYrrMVu+u
SO0h6o3gyODE01BtlEL6KWFMfin4oFD0iwcfU4E9VNqOOXOy5DEegFq1G7/0fG/lWT828nQcfdjt
HaHJpee0o0LSbU26AB5MKu4kNqJCwHfcC3jX4wEMh5Mclsl8yilCYlA0ROrEDudbYPDso5SrOlop
yonRFppd7ziFWJFjmHcz0RcY0T8+FJbmfwhWD63eN8afa2fyJ6cq2mkip30T788ptiEtBUaNEO2v
M74KbuUDPJ7Me0TIWQoidbKrwvWDTMQ2sj/G5LmucZkesq+xO7B7zkFQBvzk1VU2fY+QNl1Lglxc
XCPQcoeew6jUQ3NLe7RKrDqc6yBh1q584FRkzEKSKebLHuuqb9WCko3X8AmMej50laYAgnwWuJ58
JSvk90yyBBwVIuqki8YMijBkKUmbqI6/xgOS/1h45Scc6/LIuoKwfrfGlsedYwgkLSkM3TNLxuaB
KFK5Vehsjm+Ea7Tq3qDaxDFizSrqr0HP44j0hOEs47+EfPKPVl6z1gQWOkIaWIr/lQCB3W18N5zk
Cs2o/AJduyT9cO2YQBZLM05wyuOddMUDhab5ber7T09/3lAUuAKIvjgMNq2Hb58E4Iqz9eEKgOH5
jYKIpUaFIExBGy1IluKfvMQVnVQYTIoKyk0nqP1PQNjABKzjluVcQias83NJgwm/NnYoauHUIELF
2uK2jb/J2rzosoE3thlTvG1VrYH633jNq8luDD3yohIAKfIErXJX0AWl1umDWbo4TogMr7xo/EtH
HK7t4YTOs0M/LtATix5IoYJ6LVtGNhLaHqMeurh9c1w5vAQZZwB0Ckhr0YKVBk9VhKrOR0GQgU9c
qZvbaQap0s8YVHTLnkox3hEtlsGWOuDmimlVP1668RnpF91ufDeaee3lnZXf4XZV/GqY74ExCYwH
uLDz79oVMgILDV9o33tie4on37njghqzUJ3zzU6kfjrTNx85LIsU+UHQNJSn1Mb8bXgjMfwb3M2U
yoG9ukztNB9buNIcTK2HJGHX+EVUPWrLgI/3YpwEaqgkZalqDwrVPXpck3TntY/LuVxi2B8HMaCz
2/H9glVB8ErZR1VxyPhE96QV6Qd8Jd/1xYttmYIZOkk0BWthcSP0NmXFV+36QfLm/nQlZk0wEMXA
6T3aA2q6Oa1naGpuPKfREsb/I75bwXXfLpXmiT4Ai3FqKPkm/oOodk/G1arcILYb/eTuOvCizum3
BywBcLIielxUvQ0KD+3lDaXQZ4Jv0sX4ItwJsABYraO436ft31PZ1LXCmm/32WdqmIToNBGzt9N+
qAonlXAqJin3P5PvL/hEq2WHGsG+P48/FmuGYQ4nq0ZQX7RFRO9q2l1qS8OfIA0hYqjQgDsOr6kY
rsVSwac7tKfqCb0NA1i/ArnlJBoSQv5BsDHUsGsmfzCEx1mmE9xFL6RiIVTgjNXF/t3LgwpKVvag
Qj04OASFiPVdqstR6N0ptSVT2KiUiCydX1oZ8BMTO1dk5bE47tKSOh1WnASGYzZI+l4INElim+qI
FoFmMA71Kr9lk/OwK1ooJGU+h0OOCl26yxm+EcWBbdduQ9WzABfNFQLIeCjzH8W+uUYvCyuSNR3I
rNLOirfKYfdqE5/jy24HfxOLJcuktKsEYQ1pVA8004PXFIfyNUaLQYVo6fIaNLTfM9MD3mbJ6QNZ
LAUKoEkCx6/lR6Rb4jrU0jz9KUkmELCaLRXYhgYnfYkP4beYOnEXqm4OKQ8/mpTl0Frq2t22bf9w
c7JKWBcWi5emVo7gYE7/KlTw8z3B9F2wSah+NFt6a0jYXGG3gatmXEHBnFYn8Xq0OKq3kLtoYX2f
JW76dnLWNuZKNNQrwovoPlmSNwxx6O+leSk2UCU06Nk3H8ghnM/UxuEThGal5QDROoFWDUyrAX9S
iFknACKAv5XPW3jTuxGEo3dgh8MtgZNAiajZAB3k/QQ0tZasvjW8WnHOoz30soqxz40c8EdMWk84
ZZdfopghIq7nF6L4QjvGIGTqnGTtO/QUeUFFTsmeovw42fVbZJ9BcunIxJC5+INh3vcMK0ZEOzO8
DUQu2cLyKqR4Hq+V5Ai/6F+hM1OPYQ647DUMXVqKrzxrzqafWC2QpffD22dawJ+syHqvhEgpZ7FH
0RqS4m6tu0Y+niK+OBg65DlLwMtA9whvS/HMD/jCzgMFFd+w16QcD9OBiH0ZJTkb8sss0ImFnYlw
cuJaj5J1wXRw6/NI499bezGFBR17Al9jB6DsRWQ5rfCipiZFUE/GwrmUiBtQlFuU6/dzsFqUCA2o
A4EY+dHwiM0LqFssfecS/wqjrMkXjZabYQmN5HjZeTJ6kKIBXhQ0nk570cPZbrj2IvCGGlwcyzPl
0usJZnqqNP3xeQMwCTwGskEEYS/d4ZcGFskNxtMEog14HL3BhUWlFwhIqQCrEXn81jkJKmKktFMT
ZcqKdL/m59tqta4l27YmadH091k2zQIgACbuz+Bhuboxa7lFAmJz8JiZ7Y9jhuEKIG/eBEBa0z5O
X204tRsM/64moHIrUbFJ9JPUZPHNoV1TWHSoiVcbsexcjidmSy1IVT0J1BdU69Z9ZwLMuN9gUPS3
GADUQ7XnPxBBX4DAPoVEvideaAPekFINRGGFHSqMhALJXYMu5LlsSuKfgptEzl2kRocd8h7QzdMR
beEEo9glQYa+YQUYHB9sfHR/mh/PZVgd3Wwj+eOEUTarDqYdckGFhdnk7xnIiUZOJBA/8A3sNKkA
prFuLXZqgS7tXszB+iEkCKzhXk/4T4wp3E9wvKxUaXHH3Z/SbwKNwU2EF/fjCTsYqOh43NksHU40
BuNq4VnVuq2gAOIq+mcRTF7TmieG2T+Z6hF+wO8lLAE/5ylOTxRtC5VW5D8+U1bWbDgULmEuYr7q
L1H+QUuJZLS7/TgsAXYqVOH7i45Ki0tUemGlwu7pbVH6y53/aQMiJbocYn+8+QEMfAf11ibOrZbV
U1EIURvXOzZxSsbyL9Myvm5V+brxCZdDwObsb+26IfrlMMj39tAFjMzQhj6zbpNUcgAkfFAjgaUd
wtP+hA4V7kEl5nSPUVxmuyXTTapfjzWhm898flRcvi3l4t45mDLaiAiVNk1UI9KHFOJcNNdaIPaa
q2NVJVLzQHsVfwtvATcAd5Yh10EvEfNkan/na+/Mnxnz890LRnYgM5o/yjGzP2w+2fl/58qYr/46
3sWeEnOW50piFaBIjcfbEIeeztvrdaG+y5X8EI7lFc+6T7hQK2/DnaTK8/CQ5yppeCH3ZFXO+muD
VYRwvxz341KhHLNkXywfwayn1OIfS2t8nIMl8m3UP+q9k2x2k+Mx3cRIzD6jUYyuidhRmTEAegfI
MmfIW7oQ14jGdSB6YzSSMczrGPyDR3QHBffKw24WRZLFfkpWsVokEKfDJha5NIOPus9NbQQcvalR
m/BmbmSZ61spI2lo5qb9aV+L+U8/CAezA/59OIorbFNHxXigrbrHqLLPh4PIJO3WUqN5NtshLvZM
zPbB2pl1TpUd9Ax4tVcQ0ivI6K3/qOFwaaSoilhRBzx862zgSGT4P6/8gjH8qreiX9w6WtVkD2Rk
bHjsta2wJF04yN2b6DYiAMJWI+2I8hAaTAneZfOTT4SROwvOp13fh8OTVJJQgOEiQl/ZcRoNQvdw
BHXMBba1R3h4TZut3dlI5hrMjLMtftM84M8MVsm1rcDvWwDZpz0qe1ttxulSXi8SsV5sgqCZ/NFw
7SgiH2IFAzJW+IUDwi8NYvWKwNBgZPzu1OMqLaOw7APXsTNDXqtYkcJUahXSPw+hFJ/ziT85HwAH
bnzDnBRKvhFV6dC+CgMOzSV6h1IZntlSkRl0H09blG2eRTdZEiXbBK9PSbjKUSGOhaRHYtZWRV9u
LWU8u+BFb/KVYlQt3vRni46ov6Pwf2tLuUFIjxXz7ioDnt4GkfcQF/YoYZEFDshy7/z99WvjEyTE
5BOm7xQ8x/otH0SOjBgK2Yn8dD0kROCe4ximt4HcWEoJA0Eone1WGERS2BuW+DTI1MHYNMurkyPf
z4jNhtZj75X8R1zoddvXaOS1DYj5Qk2s6AtP0n+XUBvx4vwf9TruY//Furlx3PLSfStFHiQ9dc29
LQFjUw/Ki16c7coSqnWstDMEMn4NDMfmtuZswvj21r0tK/X2APyJcs5V+tJv6rV9iwDhpBqG05bx
TK7unYU9MrlJ9mDWy4OCE0kwbyib/znCaxJD8FG0zJuHk1f1BpIpGdNJdgKnFyXmaBt+HuIgzQs1
nDHN8lhI+OKxNQQ/W7+6aZqo8CP9VkR7tstqgfm0zzW1lwpKABFfS/Shi44SHApRXxivFLaNevgM
16B9vq1ZJaId5+vwv9DB1/Pn13cOVRfgd/QZY+JME68kc2elwpNe9hQANb+QZUGlssnliT4mjTyg
Pbzhh0HWa/bbQhCvKNLjjRfBKyBlxWujzZpiE5fRPgh9RHQsVBymAUPqGNjND+LfIbQXecGjkmKs
KkNUApycZueKvlxw7k8koqOzDUkLo78DqhA5U3ui5oZ3inmJjuUwcuhec1ZjDMKUah+jMlar+rgR
tUJIhQEEg6IBFdlRcjj7vBKGaaS9swcWKCBDmEHGeMc7kjE5fPdredz7Vdp1KUYna6VPjd+skyx0
W1Ymqf6zr32wrNAAWQIMTSLrp6F89atqTsh8II63fu/Ydh1xEa5p2oNRm2sKUk8ttJLv6RH2fbBE
Tw4jo3sUnIVAhNXlBxkpxYZFbDPJB78QvhBQFTLsKChu74M5OCDTom+5h7bJ5CiYqnkF/X/1otch
k5+DSqZcGmZnghjzZ78xF1zwVl2bKEQ3aTM6tIiABtt81mL5FtydAmh6qSvEHFKcCD1FQ1KV9Q77
sgqhPIGCwUP1CJlxf2j0HPYzpU1vO+Ane7rH1JjttCs8g4WCmUZcqVKqbXKP7mXhkYjlPtF9T8Dz
HGwlmjR1PxOInqEx4Imt9SIxTpsq0/VxMmVe69r165c7vrQuBvim5bwJV3HrCHhbPiH6ZRDZpbDX
9F9ZMlOBfuP/NkVZNcaWBTYhvkqFsEUS14/lW83LtZNlgeB18iixBVtyse7dA+muNT5SrpnpGGcg
knlQ8MsbrlfuotAxi93052vtgwVeB3P8t2UH10CUEC2jul5uu8fzbEAp3lZJJCAuRKi96qKkSdnO
3b1n1eYdncoLqk20gJ/yQxzWSKpBMKIWBydgZtMFdgPPnXfrqt8i+Sm8o1qh+sAfl4Y8GzTXanDm
UAJ+10iRgJdUzwRc2OVoA/R65GXVpAub4BojKh8wKytcBC+1isyUZTJvvMntD+x6lUi6SKeqEH3L
kxDpH56f5HNfEpLEgPKW1H5wNWhmN0E7lQLj98V0vPTyoz313UIvrsQdnVU+R6p2nvbJAM4tUgob
t+VKrs1Lf4aKS1RcsylhxYfyFuYlu49tfsapxgx0V8Qne9phyvl3k2KFnr0SocpB8FL11gAfVT4H
V99QVpk5Lwyqwgoyoey0oLV8OZSF1PIqSGtW/QADup6BWzM3a00s2K0X/iInNOiqSneL9tlugkXw
BZt7/fpMls0nzfKiPv+TSusyY6E8ALakEuiFG5cY79vXEMy8T93vIFqghfoUCTGe4MzVJl6RRe7K
a28z4uvyon0888AsZLPG9dCHwdSQAkl+NoH/LOyp7q+7qArCdj6Mdbt2JxVX9wIhqgtBU4s3iuNK
c0mSN7mhE7HWfCwBE2k7yhkrf+I8ulOWbmJackd5KCv/DL59yZtzySFESnrOZXnoSJWSA2uFC/+W
9nzpe74PKFwthlRvb/mUp3VEFOMbdaR9MfjFfl3jeoeNsemAJecPUyca1cpilYu4TChL8baHBLts
hJWatD57ofobL6S+H2HBMv+EtsC89NmzNPVi3/4vxKnxe9ajoZdlw/udQC2jh0o34xvVKwS2SEGk
Vje2cX8KB8hWClj/2sp0c052fD6rpT138RyQpsZu1cSgOLABwCwhGbzL1yFH8BBXufo1o8ErLb9Q
buQe6Q3o2+Vovl7HatkWvtDnX+YseM5XvMCyDTaGDdtDwDQk4nZkQfqoBaAStrPNCrtWsbVkb9Z+
XZrGiLqPUkokFUNAUokU52INhel5u04QvTgP2taQS3QfgPnX8/dRVt3bFwKBYMHRrt1m+V+eKVnq
ZxxpCTefdH04MqTT4b/ntf3d0XAejC0JxoTeiW62N5S/jFH7hLPpuZGo0P+afv1wSsohkvW4Bfcn
5n7kNspQFhehrFbXq/p4pnfOcdV0mJ+NFq2bUxbEoHQTHfj2GfXQ8Ultvp0XfVen4Q4hhSqXV/R/
PwXFs7FAQZqhKiHgakOmyWgdXveJxJcA0sNSn6CtO8ah3JFa17EdEh45SbDdYkwG1HliyiRFVrUQ
BLItxwqIcbHoG2ms2XuVLZVC7CJnZ2k0oUK+ubMWWzQGM+fXG4aBVdS2/lWd17CHUSeFXJBtY3D4
9lesmwzcG0fZEIDo0fZIvJYQdbw+gVZyL/TvVJKHewGNqmIOlWxWpdJG8d1llwWy336WFjZiqfQ3
8/w0s2+0RLxLgFhFnaEILfkwCCb9jvF6M79dkU7aLqEHRckxH0N+R8OU35ybCpMUkj8gV+GC0JOJ
jwo3tpr2DVbGxwkhw64aA9NDYaJ03zsjzkVGRrMPJ2rGhS117ADCIhi3PvQHEQelwXRQeDyWxNwK
9dZNg1iuA0/GLVJagQcZ59c7rUssakBowSgPtfgdsyhYl+202Lc+K4FpfzZw5KO7l5BN9Ylm6CMX
Y/KSUewMKd6lZJTq2gLmaqXUdbTiOKwofzqvE0wSgcivgRetr+iLYbR01n2H6Y2JdLlTKN46PL9I
AMoDC1+O1pgrl4gX/82diDEu80xMb+h8WEzNkYmDJ4lEaOs3mXwFGzPOT+2DiSbdDqcCuR14XeKL
hM4CiD8mQA4WTVPu0t8EEReMjFH6FxD2ieUQHr0GjNWiI7jJdpkjxdyu+rP40bEEbTofY5r2UPW6
FyuJuqxqarEdO1i4mB2UJgfyC/6FvM7ebvAK6lksbWolV5soPjGMNhPgzMzjepi+KLL8O4N6NgsB
e/CHCY/3GLT5cIBziCo6/H2o9a7gh4YmgeldaJP84d4J4RiX/1aTz3c37cHrrH/OAtqmhY80qq1X
BV2tPD36hkaLAaUCoAEe25WMTcWoYHJlqN1VGMhcQhLUCUMTJXWF9nk7klaqGNkElVO8rPrWronb
6S6+KlmUr1uCBasPP0by/P3jBvs6ipx3NCRwQhDJLEcI20nA6l+mVImJxs0q/G2N2hAA92ypJ/Hh
snGV9p3uYWiZQ0uqsvF3Qlm7cv5F/eUuZgtcvo3bxabGxd1HMJK87XLPj8oozMXbmdB4eMkvBN9o
ZGpET8XwfU+l+/BIEJukfQ1xTvdqTjF9Q23sabFjJ68cVWsHuPIAlPSov+nF0L08T/752pt8to3U
DSzPUOZrpWCmnKCaOv+DegmB2XcPeaa4Aeg38BA9RvT9k3vljKdtxcpNx43xzdvuzlsGsnPK9GCw
QyQTe4d3Wp/xNuqgmTYA72t6hBr21j+++Ckh8ISyfmqDsxqggaL5tHbuclWcIfxQyohA1TZWypfH
ShRnOMJ9wwAxmikwH3oHFzKsuqZn5vEaNwG5Ib3gQvZDcnt/IE5Z9DQzSjXpjiY+30S1y9X/Gdjt
xdd/W4ZqFAoF672SddoJqJG000T4GrFF3l3Xic1gvTrWFlltj4pLZ7KD7IU5lRt7h4FX+qMp2ijs
QFZkxdXB1pyBd8jG0ucHy6jA+NbDjAyeKizlzsIdv+boUGNP7g5WSdt5GOHS5+fw4DsGfJLKeAa5
EpzfWACqwkOcYokjT7x0OppwaX4yzY8dvu63BEQA8pKa6L9k4uOl8PcWNV5FJygKMB5CNvuIRbHx
sghe0Fwp/m8Itid54NLW55l3cYB0x/8fpUwQn3nzgZTURA3WOD3tEuUy8bO247fubS7wTjmxw8AL
1qOro9G4CXDllOpish4qLHQygjHGHHOaVXyFdrHwp0XYiUCQxuPhjHU+Fvcvz+j+s4bhI09mPHNW
pRuc5sgxwxOwdOwBTsQOEXpd5iM1ZvEYJFOjEaJhT8IC1FUVXo+D0ChcSQZF7Tqjt6ylgwVLXB4v
LM4v//CGAYdR01F/OvRvymKIjhSJ05YOk7CiIV7rSvrHrQEwGYlCWOHZPuJwzGT28QFyCBBY5CVg
yPGpCo1d5pieunBvz9Pa8a7z0liSQHr5w50YE83l4977tCDHcBADe2wFKBqR+6eaTNJMthlU5fuQ
xbtwlgrqCTOC674sCEiqEGiagysrDK4bMT50dYcoAfU1xMWTl5paCrHpzHnBe1eeaYQjScGNxuuy
sgcqY6d2pzXGG9/3bLpJXzi6CxzfuG1QqNgiRUlzTltHYNNBMO/dh7EurIEDLuaPPFS9JR9RvMY9
H1vsm2j4GvLzWokpIcOHVHt+qWf87cziAjEXPj2G8tsTNBbnO6sfyxprzgdEj8pInczlgfxjpoAN
cjPUdua+BlXQ8j4n8rMSm896uY3FN7Yd/GjvO4zBKSsOZNmmcBEtwjD94sP6EBLpr0gVq0ZqD221
dVE31R65sk4HWifkoHIo1G93l/9MOdqilROYR2758WL7oaCD+lDviymwJpaKNWUz+XqcyVlW3Srb
jzKrKwLPJ2OOG1pwkQVtI8TwpclPq2TL45xG5kyEM1TsetdyAKbfLLsWR/2ML5U4lu/DhqRJmVrz
29Zr7QyJVuCEjd3D5DBUH3PGSP9oZq44W9w/0Y1NO/p35VgPHmKZnblltyJaBLvoyvFU6g6bHhuG
JcjjMhmo9p7zaNNLa7dwFH4Wo0cFKMaqaD/GfNBfKAqrLWwN5IlHmvr8yhu6/jnpU5GR94goJVLZ
FZvE+sTMgtFDZeSQpSmPMG55vz5td5SmebuaztPSmM3HJPMR2Fz2VSyWcM8r+rbVWYMQ95nKQXzp
W4kwcajr+EcKSQ5JK1fdVWbq0Kv3D10umW+ZeSMWDiojqS0hClJ0wZs+butGTI/QpxBE2PKI2V2m
zWFhZZLPAWBZzw7jgnaeSTF3TQlleNxfNJBD6KQAb6tybyuak5o9BmpftRJa54fsaB2A77sipnev
K8gelTdshaORZZ8aKH1qf8t45/rm5eZ1KNJLVeBE7Bok2hT6uEZHa7bAm313HQsvnk+xGXSt4vL8
9NIVkLD+UKEm1+0raAAS2aOq/SdYtgoh2qFom3rps1bYiYxMrz9noF/LOpzLuuvC8FoJ1zIWr28U
vQWx9AaFGxlbl18dUVypmdnDDPxxS3XGbOuOLJGysE/2cT4xS6v4c08lUgdq20zbC27naZq956aM
bOhyQn/qL8uFviWumzlh6rMsAtBHHEM2oS+XVye6bJ6EGYKa0mvtokeKZVeZPAnI1+/j3csXJJWq
ClP/ltbveqRNOAA0ZMS5jzU+b9mDajdx4Dskw5iKVymhLay194HK2lVUN98x2lJdgg6mABkm7c1C
fT4ff6RJkrefb6cNYrh+ABULTbec9W0Q2HbGwWxPC921EDh38sv4DJPw3K4spJQpZsYBHFyl5jZi
Bsd4cKsMUZzGMCSgJRmlgIOUg34zBsiSuBIGUFhBmOEhBMEsf76s2OQonpfLG+HxHxzsz0/rY88c
2gT1MQPb0eoMMu0nVWRgS/aV+6Wai60aoz+cE5k7RoMLhOrb2Yk51HsGr+WyEww/xxfklt+SEPxo
LvrGHh8pvFhbAzSG4ZVtVuSNqr6QOKNNsAaobMe5K2qZuteWSlnS9ZwS1a9OciX/wZi69QJCqRe4
hKsZ1+lZEOe3CjW3PoQ4YguBJVZNsRFhAPlotEUC1tKJRcRO0NsHkTx1MWypwAZ5sheJpIHajhqQ
xQyADtm5b95kdh5cL47eDHwCY21PVkUdeWt/pB6iXbw1J2mpi0C+rHKGWY23I/aNa5lwbL+LCeAo
lKjEzS+MWYGpwGdYWlZvfRQudN3XB2tIj9eHsYnXFHXfdWmSsMQT3qZ/xAFptSIJ3kofPg7Zr74O
hhYtR+Bg2YJMdZIzA30wPBQIMT2mJ9jZ7AS+Mgb3fYebWVyJW7dsUg9k3cbmZfO4oK8HFJrFGGv6
ib0qsGCK3USe68SgT/cwY3YCfxdLZ0gv+ZMZRQ/OlafMZdtXw9wWJnOlwGuK4PccyvPDMlvWOMPP
Re53D9zv06Hyuw9+EbdyK4Nkiz4WPKTBocphgNkdR9TedupdsKiSerI/xS1nNbH8GMB1EcC0Zy05
96jVa0fHHpm2KcVkBw8GXAdqIKyNaMAwFuKK/df027bBO9PagFLGmDQ7diGnd6XlHcnBAIKYou+o
bGyFxeoqqcDbbprqHNlGwi3WtazqOQu6qyb27aSZ/u6xaxIJoX3rIdMZp8w5tZcgVanXuP1xQEom
AH0MS2ym9eSGl+F30bKZYW6wLuoaCE2FiELrOHoEdWEvvNw0jOR3e2sAfwCjZ7Gf3uvpo54bbSGC
0jMIWgd1QDsVARAiDQXcWLo+294tgIAt+UQMHNVBfLUntlEYhwyDnysps1lQbEaTYckuqZ4CaNXU
Jsb6bVpsI5Sj5ZkomKffGMpi04aLec5KkIs4VUahmQl5GQfB+eUepH1Otyvfv0okWgeq0bdv/1mn
AEyXWVZWOF17Zf3QIiGe39llhDRuisfSuyvtGRhlbqZ4wV9v1XNO/dOM0gwtBgZhg69fDBAMYcBg
b9yX9zr2F3xomlQKsvjtOO0NSq4mV9oVct9/5g7LmKUhBtwccVx9x/TAaFNoJHhYZY+qtESD3Fzo
HiQPSYyfCa4JfmPN7vkHErTRxC5Zpt720UU9QYKYxVyAklpCvqzS64M1jV7stKFHfC0bxU/5FGrn
QyPC00UTVG1Qqy71jJuR0Ve8B0P9LMoCFS7FjWrRzrBwd5nOdnauiWmNxmSgqmfqQoB36cAcD3iS
fsNOInmm+jy4L2KNqnCGhRX2thZ4ynbRLzlpSOSwDX7lqEPb9WUBNUuDwUOKQh90b+bdKqLUqjAf
fKHN+4r9bKkBaap0Pd5XPJXzVaBh3FEdJ0wAZowmD0lcBLkIJ+CM4TducPeNP7K6sWipqmnOkn8N
9cd8q15kcLPiJZzH/g5I46zHP67vTTwVOGlgkJEsDBId2O3XiOqxYWVPUqnRi96o7fZqs29AKej3
hd5SnPLx1fjHbDkjqlp3VdToVm4570klCymOXKpDEjWAECAm+pSZEPY3Nz9v3k764uZGyPLFyoe+
aA9WBAEuH3dE3BX+cF8TxA6FX8qOtR9tdiRrPQR50RNbASgoyaROMge64HuHJ1hpVHYBH+uGn93r
HvOJ7KDALv7f1NDnoG1QkK3AJCpCi1Xsb5WSp/3rRumCLwvHNIuh+tvH+PiaFgWJ6oejzkSSolf6
s1rWkZtxXHb0DM6jygIgDSQQ/6qoqMWWM7kVK7LAtS986pL0oVL93dyD4IPkF8RaqSGvJa3vJ9uo
QXZMaLQOmMpBru9Y5gUoxUV/y8/YS4nTsp2iC2UnyAENR8lUFkrU0l4EaU5ix9EUOIj7InFVldj1
Mxx4XzXYUWqmTnF64jzueZiNokPayhCSOq/W8zD1L5VlbwJJOBDVq/tzXVwD72BbO+/AFqhFlW6a
44OV4jb5k2Ogg02ZUq9bKpSvQ3IlmEP11ezcCAxap0/RhdMXuSLMaXzss1of0bVRbV2IXFLAMo9j
x7hx7T3LjCapvmouwstkXtQLuNrkZsF8bzqFaiUM5l9o4dk5Kwy6in9qEycFU/UOvWhGSDpQTPDq
6YW7Gy9f8ljKEWFu0I/oxiGLFgoHVTYhxV0/1wREi1SqkFKo+M2HV2gYlq0r62tif/MwrUoI4wqu
FdLd6rgsj35Ab/TwjJAG74tjaQdEVB0fO8ccGE+vitjP3cubbvdJZInFQt2sPH0XPm9xyfhV6Qbp
2+KnRnWOKONQ1mD8ptwTEJcpd8FlF9gZv1VHLjH8X2hZMi2eJrC9N0oMUul0Ygcneh8rUXUKPUS7
lc6f/pVFtRnVnVD9Vk6M1K+juZopOUH2SltHEQAQ6mLukcZZoqke3/c0JQ5osqJzLqzl8KOa4lLJ
HVnqAxilLjzagdFD1EUi3XYkMqJtAV4WX6M278NK50Jj/L6uiopexIDTRqfAZU+oo+0BxdiSS2CZ
6IanWS3swRKAsCaAnCIjqAY8afn/1dtrWSgDE9R/5GWJcv+Jjlc5FYYkaW3nLzjubsL+8i5p+Pl5
LMYohkMIivE1StkDjntQIz8Btmah2yzs1xWB49KraQiEAmg/lV5GU8R+zaBtx8DQDRkD94CXxL14
wkgPhpJGPOzAPa1uvv3d0c4WDxpQMo7ry0jbBC3HwcAqHL2UzWw2JDYafp9gLunOpwMQ7aWcLHBj
Q0gi12p8FisA34l1tq5E+xztknmfvKuAeo5U9NsI6RF0Dkp9rp8yguHOdoiKbIPsBJsM+VFMGIat
nl/SZXFzul1FjQmRpZZu72inDG4Qi9M65Jom449hS0XbuEQStWqglX0ir9/t8C+Qvlr9Cayu8DBT
U2/gHX5WRLclipL8d54qnMeTpqPsJwx1BDDEs799pYYyUPhD797/AckdCVFxvmm435k9r27d5YR3
bKJmLJTxdxcHDlrRk/CN+pzACUJXxa2JMZXjUgiA2jSGRIXuyZxxCNjnCqYEvO4rpi7e9Ji/RZGz
7ZB+UVit3x0oOwDrkDeechN5jS5Ls570T5YhBa6SMsEyBV0JX3VF0lC4kpX4GstRS5dVmNJpKX4C
tTsZ+1RqbUqHinsZJi48kemVsFbTE9MIA78/vwB/cF0U3HN/PaVOO/KkFM3qzft+E5B1IX02pshC
heTKDqw8W2ILqsEsbtzf0fpfSrc08fKoLGZBVFGwQmnkZJyngpo4rU1xz5GOJcKhVuyaeZNqo1LK
vlzh6mDkKEdNu3FFFB9Erofq0aMYoXKHAOazb5K0FcRnVxs+1COMu3AaFwy9F2WXKjjcurDqECgT
Yk000+EqusxWlnDL4uFfcANC61kmBDYpUNWxmhfXHeEIs52gbuO4UH5utMJ7Bym0ZZ0pGwrVJPg0
q+TG7UB8EYYlE9BRe8m5ZgUnXobAbvhCK6MT1cL6qUaTMzPxaE6At11RWkNVuXGXlTcM2mAku6lt
SUVJl3e1En9a5d5r0kdRP1Sqy4O/p23O9zNZ2WTRiUlmJCbUK5yE1xQC82RFJ1SEc95fG+xdHUsp
eBzhkpY3DrxYVP1QEvdzM+GtOEXvoQ0r9U98x+m4xkJN8f/5eBtoUD05AUPt82v79YQ4+jzg57cG
+OBi2BW2ORjRW1lot9EARv6U207vAYrF1RD2qqN+LHv5ldSC2USjCpO7d22ChJBUYmhkeUC4L2mt
BWu4pz7ctG0hB1ItuYp13wa91iN5odIEEhMdymDp2SXV8VSurTqRx/HOzRLC6tQlmp3Lz+yHA71l
fryADzbCLWqCxDSExNmXVoJKhBy071sNwigFdJUXy7PTpYRWkYn9CF8aloq1ffD86CFNtB+6wTVH
RarDwWnGMjkAGSKu5lfLXG4HnM2gDmGSIVo1Ywy4s3jxHBh4joGCI8ZN4EO0T3j1+vHeBwYQ3ABV
TvWTfhXccCEQS4UVyQrH0w4A17Fqa/wVOXZmY+XmP1t9Ew5dCkH6ARxgx2akTcegjKcjI1LfoGIj
cDK9kVnbjRvFEgqrx7GDPPmSeKb4o4mXNuwewbl/HcQS1raHUZjLH0jm7JlU9D6CY1wrUQ9gcwfQ
1k2a/7HBJ8JlxLVHZN1v6W2tQOZaiF+Plf0NNTMYiQEWpsvjA9JcQUsLvbzJzzKLpUyFnHW1UeWA
69PyinTPQTI1VUKk9OXlToiWZ9PvzWI87vVycZcDWDVs9LKCBG1vJot928TkMyQMk/FTyEmD9Byl
URnplr4Oj3u+l2FAQpG4sG8LeXOa0C3iw53F+GpuXJga2olZMA5SpBg9HbW9aaHr+0dY1Y9p9XhJ
AMFt263ofUTpoqg8FHqrSZtRkFHKHaPdd4Z8PWCSN1V/LU369rO2JbXEcXjBeuKagH9r54nU3OC0
lkwNQHrU7ZxUvpwj+mCjB1/lp+Og5HSMUOv1aj0TLH3ZMvphbpDsereViibeJIdZhK0rkbBjvg8f
+sbXi9faqzJd5IyPiDltzz9MZsAqC1tj7gGYsgwmQFPYNPg/0/1IVLmLj4Nn8oSQdbbo0RBC9LFG
H0hMUM+8+5V9+HavZgkr/KjCKcop/OiNXs/onZukt11TKIu51ZcACyLUA4l5nRZvgoksfFMYPpdv
OJ2AGlBTawpzTLHYgc7WPj4AffZVFBHX9S8AfKZU3wUBvlI6swt5jnvfccXRgs13H7qBBhqQLkyX
lMMum27z5nfkKHuq4QhNM29HdoLAw7cmNEdxjlwekt5XwhT5cqTPkMZtD2ExtncsHAh0NlkL9G08
XYPa34S8EjhsDq2Pjo+7L9/l2FaqSc6m4JYbiyxuVxLs1Futht134ZPvkroLZ934fFN+tVQ5ey8/
s7Pe7WN6MMzhwIjomn2B1/jSY4fgjMSsKVmziktpQwJEKx+LBeQ++yRxImI4DA889t3hS+WBN7RD
uaOyfB0yZvbQn47XPPYcW4fNNfCcq3M+tBvvneV3AGmmaSR2d5NCN+XHUCFAcm0xt6Mtp62YW1Qo
w8wRlKVvZ0upiBrd65VJ1c/UAiAI9vKrOQ+npK9N3xILXofYvyojCqcwhhE9Zo/sRIkdoMxEaPnh
45aEYShbLMmuKarYNAlD3eqOM7aMxcaO+hTNCM1FrWcgsfzyzG+tulv422R1x5VXrWdmAWApQ8ra
080a/KuhRFYXThcY2SgeL9LWv+TlDez4YM7HlvIQYHujYdGQCTaVObVCwiwBqPIwdt8gAAiqyp3Y
aQ45qqjFkmQYeKOnDOU3P1askHNyTKiHuYlJIfSITEFMqpmfUTQXXXctmmzfFmy12Tbf7xpt8j+/
7HCglHKDOrYmLWsNNjfY+kGsVwFZwRQnwfZaeLSFUksBsJtvqVA10skxRYJ4MlAOL2gsdyxI1bEP
tPLBHYKk4IbMqZqbOVzG/D43LCatE7FOzonCBpTZKrCNfr9aNWYL5V0ZHH6jAFscTl5rePN1yULf
2Lb/h5Pn6stePBHzitAOdgaBxOc7OoB+NyVQMnss+y7WyeMLjdkGQczktJFV6Qt4P1eT8eieyqVC
HpvD3yLjt5lbCrY12Rg1j55AlLdJ+EMmnMTgh4Xy2zJJeOSPEwdaVwHLBwKRQG78tx8gYLBX1FiP
PzjYOqE9DH7x8nnqNkjex1VOsIQ6i9hSHzJGnXCxsydeE2HYeAfcG4fG1rS7RbQPD0ae2mGB1v/O
dyG5412qs8oMoUBLeuVU6ky1VhJuygSD2dxoSvwuKMUw3B9hILwhhmpNlYPVpHEyO8SbVI9jVgHC
KlfuZaIv8xXp6DJs5Ip1wmJNex/CECzIobuARRUU6u2CjViO8+mFv+uMOUTMSd73i4wEynKSG5Wh
h6/ZMzbKWa3BGnOAo/Rv4JxvbdLIqwPFp52wKBYsNfgYuCT4n5vwaGMY1knc1jxUu09T3a/dL27o
3JyLM5nedsbd2EmcFTVdvyTTZ/pcZoxW0BSJo9wi39K5yjP3BMWo7zdXYHCK9i29/UP4zbGIC9MK
fW+FuKC//Q5nozsgmg7V6TGn/FJRqg7mj7X/iZRwX9WAjrn99NWfOTuk8+fNzzS8OEvZTQ3E8G5y
nHyKwktnENlVUaZPucNC9+bOk9Haf7xQjsdQQvjk/icPJ36mftimZzMI78ywN6u1QPUM0FVFQQ6F
2L1cROf0csJwKDN+eb+yKmf73wD/nHQuAJ3ElhZr1NS5TP4J3s5mqtETpC+UzatbtvWZhzNvoUhm
tKH442V6+N5epp/CgXWtV/iFW8nlgO8Agy+/pFQI+sNoVaFLXKRKf4GMxwmJVr7uf4uKU3QBgloo
Xjv01/jdNfe5mbaWTjnIlx5G7ViEx96V5dH/3FzVlBj0CDtWjUm7tgEDCQwuHP2TAG8ITcwXp8Nk
ekk7vjCgUJjhy0YS2XDiC21dNZij1Snf+z85rPi/vUsZfqcJ2RUHQFkukf47VnAOmwUr7PCdL1Ir
So2txFRCW79w6smmXKyzH12aeMu4viwrMIEyl+KWL4ELnPR01q02H52rc0bkClAefZ6wfRDaCHc4
B2M7pSTwGbHy6+/T6rKxPjeMs7Il+H/Y9uEJzBnFk4nlNUcjKYOjSWTHXW7oHo6j/nQXK1LdSA3b
6ZMk+7JTfE41IjNSSMVl1akM8rOlvtYsUu7SVP1kv5mGcLRAp7U2lICwHUCG9P1B44IsJMnW5dak
3J3vJB7UTlRNdk1XA+J5OsKwehkwue/F94U007BfwmVqzB0PbrlSEaPFf77sAX7g0tzXNLWtWupC
8kNdsEHh5cSiOd7hX+TVduiyQuepZu79jeuyBLGL/EPZMKRharvysookBlIy/haW4i5WVeIx9pAX
cgHvX2UBTYfByC+kKDn3xafd9tJ2GxWzErj06qhrqMvYTXSbYEvNrB1gfJK33v0N9iiNDTW3m1n2
t+t4NjIx52rCqBZlhE0ph0e/hY+lmnkpwZrcQGp+XhC+pOPJEIN1NFpHr7xIXg0Z3AHnXYCI8njC
JlL3kOiU0C+JgDAPC1wcSrQbnqPDlt+2E64Cifl8rleymiU3gnrjFZhAvIwKmyhkj7LTSoBmj2BX
eL2I0+foPAdwJpxX2ml9aiQhECSbjPX0Y/KJxxQVxoSxtWZqjN2Bfz41gpi+Nqq7VBHZK590rP5f
JyDrkipZHiFlWFWDAx6jOcUkXH/ba6wCH2BogxuFWCiVgIDLH6l1+XJnPjiYjVGsde5B3fFeNvZ+
TyS17KJxmmzivLlPOI7cMn9QPOlI70jik8ez2869S//kJtc8LYA0ojQDvsFhojVIdIZsrGfouBCO
kidn3RWq25r9rc+nA++cq24SLNVbjkVeg9JY0WbUZVO50xmKwMXX2qkdBTh8CTxz9t00Y2OAjrI2
TRPU0YRvvd+P6PhRmOyosu9ZP3gT1aCIL+RYC4IILWV5aIa1tK1HTTdBIthvrj3DPxV4JeQAAl3r
LcgaVeqvmWOwXuVdYSKGRbFpAJOmyx2N0ToXRYdQlaI/YZTanypxDsC6qv2x7WaM3DjFoJzEEjJw
T6VXjieRGtfuCxjIo7pm8DHtvXvr9HteRrIHD8atmIgitYTNIreQORmllml4XrPo+yPwiSpnSrLS
XnZ6IU3WqsOn4pz0YGUpCdhIQmgsMPDWjRaBzyRFo2dj2fovuUhM6ai/iXxl2wl73ja/xH/okGeO
MilIquAJ2qaKIXjg5HNvtzKt51sbuVrolqCM81lstQpnF4ahtySpBgnE39HTKi72mrFpvqKAb1Bv
mmXFl0lStldjkr1qqIBSJ0BwcmxzX2qHGXhzGJsyFh0wlpu2bMOQsEZteKEqAfIJ86XvKpyBQTWm
UrDYD14voSPhWrnLXPNQ6JYngX+g4Gy/PfKzxUEIF20gpR5H8vn4ZGpwOOxlDSGIbHEj+zIEDQsY
n/F2nVZFENOkktN9KC3Jeant2a8oyp0CdwfsiqVeFetB0kcimAZMxrQYUkmMoX1v1wTGfCyJctc6
9Vvqqe40ilpsJfX9YdkcmM4IA+I7rTuboL/CDfqqYncPQ7pjFEVEBVmPAYuy2DPS7wD9fxLVQEoL
JRx3Idnm21lRbnv/jh7blHaVEORxjbiEv4KzDY6vmmKIfTsO9GDPp/6k6QRyi9RQmW1EQ1oLcJwL
6a573CLcpCygZwBEv40fAFa4fmow/g7LNegGsJWpjvrhHvr78cT35+oh4E++EByQVQQwkyDjswZh
ZQx3dZ+M7Sa+ac6xJN2iImen5Fvs5ctJOf524Ad9X1X3y0bxd9BE2Sedy+2ioOuWo85NexCT7s4W
UubGS0eP9CLJeXHX05cDTZ+VGDV5I7pOOAaa5uIHp145FeUTi0Zn2Mg7FRbk4Mxtm1cxouE1a8ID
JHCG0PzESg5ZXtZfxgJN/Vm3HhqyTpCyNREf+fsUhaYsiAWx+uWZft1kGXLS/abVMarExVeTb6zW
IA1zLkdtqDrtZj7kXUosD2GxNZJRSXlqqawIz4usB/THzeJ468oCrkxSJD8V6NcNFu3D0yhK71p+
VBmCSqfExCvC4OTRI1rnglQ9Nd+01uYBxHXtwIsZJErEYkhqV25RoEC7Jf4IaEKoA5vGD1h3P/0K
D9e0HA+DBcDPx4qL0NenBblwRWDz7pqLHXt7/w5b/SE4BngndaBv/hMb3fzbt8XFVn1eYJG9vCLa
yxLTQOZtbL3+zjezXGK6bb2dY5sY2q6dBV4OSVzpZ48nRDrfDltaEOkXxd88w4pz4wAG946XV5ep
aVwgocB7ajhuOuVX/zDEqI0uL0rkGIk5kRGKrFgH4XNgCOi0k62H5MiOMK/hNeRTciZlqYWnGMrn
GPfU6opL6ch1U5HLkJcRP0cIwFhGr4PqfvFNRRCjkebVXxwJM2YFsGscqbft16UjL3MbNCfVc9lW
QshxG3GPocKfz5NkOeSGNAFsifBthovvBm1q2rd5JboG+PwVjOqzUnouu2m9aB1Y7mXLBw33XBrS
Zy792f/hbTHtBGRHwK2G4oRI/G827xicezW9eeijkNJkQILObpkTB2UG4uE9Qch9uwNxHfepellG
AdHTRFN1V7pHTKZrkkxhhz9bxNfNcpfTrJEkpM1mWlxHrs6Vyc9HAtPlMI5LEncbpbTvhaVEH2hM
a2mF++s/2PvM95x7wTiGpb17gPq++9b6I+Va9wk86KdR1RVcYyZ2pGWzR1kSPtM80M7ykjOZcJNw
4kdZEQT5kkUNncGsVzo1T328rxSWEAgKb+54dhYgdwOInw6UMPUWnzMZaZfGOktqG+1ZCVq6oD+N
+Hkq51AjLEUF54VM0Z3fepSvYPfg+p1JNZQ2BY/CNB6YgVYlQSgYOcqhVqe5ZVfvFGhJ+RZhPQ6g
wnO83gQQXLoMj7FZ1NNrhZRSQ439AnWrxJlXlp1jnvu8x3XScwz+OeSwS10aYQrUS/PnMD4cKTJW
HzVDnOVwocumg2MA4Rn3u4IQ0qhbUU5iAwa8QTz9jZhosBvbLrOo6gfsHV1p+ghi8W9XCGpsYfaO
C3KgQ2G3KTWlAbCxaYqBJh1dHmJeN5xKPqwmc4AcrVpHKJuQJztdsaP6ypTp94A9PAqGLAhjm19Z
qOMV0/DhUsHgCB1y5bTpNTv7/P1yeLwlqMcqMmOHsmdIFJ2bSxguW3Unln/uODLTfvMThjjGPEdl
WwM+uN3SWunyrCQepxRoE1R+05IWzBgsFHFPs+mNHarz9XLX9Cc+cnae8n6b0+3k6lw9w46JBO9R
jFLXrj8DUnUSX2r1hSJPRstsPRKVJVCY99I5xwCRWtPDoh2xYLZDnLUrmgtavK6VQ562OMYxOeDb
8Eq2I4GH2lUbZTjANUyJEclSZVPbVoVDMonM51dkMwDLhtumV1sNuJe09wW17k+xAHRtHweHTHKx
V19PR+R8QMDfvU6gCgkK1Ij+GJJzdGJDZxs5DNlhrZq6vjcaBBRY/r6wyISchVQuNu4/pYOMeGou
ga7w4394FXffMyaIsaeM2FvwC2fdtUk7B8WhJyQmRS7iHb6WuReQ1b+TGtJc57D6qnnG3AAwQ9do
MAGiAa5dfINYwUJoYHenU+sTJbPnVGpYY/Hd5K5x/Bpu1oKhuqvUHIG+q/75db1WGytYrYmr6Gd9
dyHeHzR+w9mAHKfBBu8KfQvWMpvJM+y/lMEm5IiUkDHgjlENXfY5zVH/B6ZjQL4+Kh/fSuD2tu8s
3PFHuQGjojpZCsEhaiyx3aZkkZxXcfJTeD1omplMq6XG5Q9IyYJrTRpf+NaD3zX/PfTGZHArB7OU
Yvq1eUKKQyvVma7tuIuI6rdJT8nXCn+Xm7uqa1S3zJByrTryWAyfbEGeJ7KLsOlTjZ6TG3QNRQB2
0v8NymP8lDgbC1gguhG/hv46HI9LWwTYwMloj3Y4Jm2J+2QQXTHkz/K51KWj8rDIHhoJ8DtEJPwu
GON2RdPW131OZ8pxlUN1xnpJBALeTVNde0dNk6paWvNupCKQDrLXUoBzUobAKDkkabckooxofyJD
hmBVwSN9upIDvi6CZPG6uRVdRugG1X4Ua9oq+uuaD5TN++6Qxe/smdTeh4L1obWhjdy+t+F8VQzT
Z2ymQJiBSIXtTp0nzQRRw9VG24t0SwLSeStsFPlgjzCSxmdwzNZqUVgIzAVHtKAk6qXyHsy7879j
T3Db/67/1uaamqWLlLC3GH3n/3LihNPiUVgdz0WMPfEjxuCVFp3+xgubwwKY8IgXbSR/vGnIc72g
1U1TgacsFzZPJHfLwjpXkXgacJHC0agNT5K/ALhXdXt7xfEyMNQ4CXTYxBY2+DrMeUV2tfrTsN04
WvtQzTmkhPKTKnjZiGHeVg2jPrnPwcGSlMa1mhZvui5bmy781x12ewHUfNOy+fOXV+hQCcSCf7Vc
v9L9aNunFZMfH+8x/7bcKWCfO61ePmYriWrGQpngV8RL2N2JUW++R8fE8CQtEW9aBy7nxtg9O0Zb
+DWXtZbWQo6ZcXONTDyIz7LlQtxaQzeT3c7MGEKQD0UnOAevExmi+U/B69wyaFYAFKtFkyg1lcU4
OcAYWuWTkAUMHLjP5nimIeFu1Tf53I0PAjR4lfd6VyEeT06l/VyHzI8SdsP/mfAlOwCkPIHvU+Zj
UEXz4Sv8quA+hM4kSXaRqzC4Gmf4lx16blhGx2KkPYrRRCxB30SgXw9C8BdBjaEEFWt4ssdkMazg
iS50zvjDX0PxE+Qt4TkPK+yVdIg6VgfXBupAoyd4kQ25If9zojWUx001LRRcdYE3JOHp5UABNWQ6
yOqesa9UXZYDOWOTkfCKXiJYdYKCy5hvAOWXXCGxMoU/2cu+P+FaPkId5fraDsth8QA0B3dBTjJG
8e2r4JJa78IP1yHmf0T5LNFgVeYHyvQT/YX0jYP0qtkVwwmG12sNDHhM6sOSckKgKA1sLtsfv4uh
oLm3WpfLutkYdVnwi/qQCm/za846P6Jr+0DqlA0rTT8Ued9GkignHx+uJRIXDO7sIZTX8UrDiqkb
hx5GSwqmzyI4sqwjXW7GTcfFYQEFl/pLRNvVHEYZD1LVslKF0opq9Emrzhu/N+0mWCe8OXDOMSQP
hNY94AQXn+xsy7f37Qfn/QPsXJcc6e83JSQQTb6s1YRAQUhChiV142fi0Tpf7iRR8PzEjdaqnYDH
GLDIqjax55FE+1nX9VQeg0QCV9DaoszSzN54gCqeWLyDP/FqDLkeXlEDU6g9S/mVObppgis5NTvt
BlvBWR36dWCFnn90I6+M9leuTSQDoReqLNXwtHM2XX0ch6q35zb0MP+/P9nfSQZLRTex44L0UnZH
uJ65l6XYktX4yN/2kYf3u0OJh++ouAYXqaeybyXXYebtG8Vr/JTaUrYVv3i9m5RnT2rc0DI+ubd0
abwYPODQdRZWw/zV+w7AvvVN9r1w6Fo19XaYUfwx5vxN9K3vK+zfEtEAzjti8Mx4YDsv0axAM5W1
1o2LjuwZgve1Wx/cQOIMWWRFHPwZksfv/yDBo8FUG4FSa1Xgh2d6bR6sS2rQE1SR1RTmZtOAXALF
RqL4oJRf0BMKwEOTudCb8+IESJnaUma8Y0RVSguQ4FD+RVZXlY7EniiB3hy5hHl/kdQEVc9GIca+
QsJTNMqokbmiQIF7Fr1FImOtFG5CRXtoALcZOlhYD158Li8yJN3vc6i5l3rdxH7aUubnc9sSx6aU
uIJypbT7ZBXF28BKPnbtXuKV98gahponMY1pND2ujtVUaGXN9wOySRlbWJ6Gpk/hZo4fygKNgHr6
aXmX9vFdNhskUR9jtD+Qr35zzl5Pf288CzMf3RjkNAHoattKsaT2HDpBNOTO5MlgEYZglqBJ44vy
HGvhqh8FW0eHLRuddWZD6OdwcvlaST/K9zc7yLmfUe7vs1Rjl2JqBrzDGwmP7rRrpa0usKcXXeES
RMyLChfLyqjaUk9FJAU619mRPllBkikjw2N13ruZ05ykfHucxll8cervGt61XjUwRxERCwR2c0we
bzXCES3MQPDCczayb306iZc3ZhnV04/7wyDqWenbK9sIIkvra/JMHZS/Jku4KgRMLoGOvhKJ0LSz
NI9NrmLWDi39p7/9ji7WiDd93zFiCHNtDl9ojF19hU1ZuKwXP0TdezhHcVH6gmO5yBvBcU/qW4U5
DXSzbHrS7y9od6sWmbf3i2rbECt5iUn2l6VJCGhj+p/1U+RgC8SRq8bRcbhZG0wJMF0T8XyraUGo
QXLaJHA6++gnKMfpoSu4Z6vrXdtgrRoS5OY2zHm90gN9oIonsyLEs1f5tTSClKLzH1G3riUgcOmh
sa31eOcvbb0PyiMxAcqfbPd6Uwod1jDc71v76D+jyugJBwDr1GBvLie+/qiV0wVaSdjuJYCVQd7O
X8G5Z2dC4efLa9LU2JFFqNw4o9MtPvuYn4i8jf4wDXxGka51v09Kc/j7pFG/BwzgOskowKhFtW+D
7kOtTp1BKOTYZhZhUV09xAqNzWWuz5a2vgLUqvfWLRwVwM6AI+3smuJGcKyvs2PZWexMhQu7msTP
zS8GWYun4/CYN0MvtnFzHYibmIlfPqBrVtM0XvWPIGT2Pxoc07cA5vdMcGU/5bZTysVtyxVGdgFl
8rDNttmzvhhaODctbLle1QFPa214SnFkGU2ZxYfPmHDwR2kmqKOSnOxRWQPE+3abtoLMtklSHL0Z
wCd9YzrnEUBKy81ciKO8RrBpwSu5ch+gCvlJR83bdICWJiTe2U9PlSCuyxPQUStg7ubHGO16KTFF
grd6vlAh+ucbDlerJglVD9Eea9YN1RFqHlR/IlaV5fAH9qrqfWwSFyQIr4zfdXzy+yxonOIoLo2I
trINA/vamWBASPE+S9vZjBxUfMMc5qqtX8nSPoQp0gdZqI2N7XKLCT18JxFB7XHfpQHXQYOb4ahf
H3HqDx4f8tkDEmlIX26Bvyw9CpqfZxc6puwgpk5PoKcQTWR65C8uv9xOUln+Od4DfwnvshXFRDVt
mrtpjGWzGyZXwF2QE7txioOInsckk33rJkMQpldR7VwRRLT8l9/5far6z+1IeRGSjZf8/zLRhr1C
6g/C4VrG0fC5NgVM+K0hAcUCxdati4STWxYR+/R6D2DVb7PQWI831ILuYYBH+FexwK8u2B6wkYtb
O6w7NA15vYz+++n5lUluQ14ls7vGgidOLHaAtxZGqhnZtFXV9/eXl68ZBJKxBhbdI22s6+E4LKN9
Y9dz5QW3iZ+d8Ubutnd9bvJfql8a13dfLsfNf/9bK2OhnYwMzFiKgJ26gbm+aejzpHbXgHZW+Pq9
83i9n1X5YR9fIzZbDG09cDH2hjtiTjfpExJsnaMneXUYxu/Yr8FF+oZKLjlimqHfiNO8Ju3G+oDd
/DUOWQqkfma+nvB6hnCJwkSUUAqMhemO2gvD8x66BkmX9+0JHRPoykZ6SJL8akTuIJkkYLLKpfAV
jVfEaad7t3CEcqOf2hj5Vjsga3Y/WWpatyKJXDSNn3kUPtx3sKJHOcJ4HOTnYW2EncpL/ZS/1zOH
Lt5SQxQ3kof9gF0r0ZxWjL5tVfiKi4VdyvhmL1lwH84snxshQwjtEy+GRuIKCOXvMy9nMseEpe9C
ul7fSaDS1FePbPmr5o0uktrixC4/+oU61SFqVUbmm/rxXYofWqRBvsgzcsoTJ+ktSRh7Atd3vP6m
awUoZyPv+Wf5r29waXtB3Bptb8rEnv49Wwn+iKBHszQJUyobOZqb+bE6rvPs4R/T88eCdZanAM1p
1a8mgyku7JzWJgBwHQq70E5aYJUXCsHoOxedVYjG+JFkcojuYGU5oHkaB4g5/DwSbpeSjT0l6Aet
6AB6frJJ0eAc3MdMqCqC4vZQqqW2TVtOOW71p4V7YztJE/5q/d8hgR4mra7sARt01xM6Er3vWooY
NfbjGYIcVkKg9stUe/iF90HcQrYkSj3pze8qifFAkoJZycj+EixOF11PhI3Ebv7kyWOrrC/vV3U2
BJonPEKk3g+W5C5WNmQCgZuM/H+mbKvdCiXz+TirVNKw/7K+VPC8z0w654sGwynWQrM5qFHGUoWt
Xme7/RyXOMGQo0Cj8BKo7XyLD3JGJydjge4/+2MSOTtOt1cfz6+0VzwxU+fosmxs8Tbx3RSz/Fnv
qDk7yyhd55VBbDQz7GPeGxWg09bD0q9jw+qOSmEgaH+rkUBzPW6G7Aa/uRxpiBayKcUka+e3Jen3
MToyuGU6Ahj+3wNYNVZ+/PX2FUyEhqTKYpiukShqf1utOEH4o1yI29ltZ45gBb6wjBc/O3BYJ8Ab
IdjxjDS5PPSCPEBf0OYfSj4+xmQLYnyFHxK2bnVb+ghmA3MdyzhRPUE+GOSFFIQ0bKLzC+8SaWHh
xKEAMIRVba/dXrTDbL34yKpWePGLe9Ke55X0fX8sB25tiRcRWqQnxSSO9USE/wwUTGnzxWilzPZn
mvelgaNDcv+3cRVz2bO1NlAMoJaHFr3aCsv2nETB/KyT5GAcEU93ZppEbpFnGK6eI78QoXw3PmMr
YJu+9bup/AktQPD62IuMEge8e00iE1XoeJMj4OSCHiT93Y0h2+L0aQizLDItewKdk6MGbbqa3O6G
Ub6jmM2+NM0gK+0R9AorYOheKtD1eHChjlQ1Fd2YbivXsg4DlySYQ55s07oftktG+nnvzdgmF8Se
rMw3bYYcccLXCckkosk5Cimujvic4krLRvm54cdyMwvQk/iGg4AmyACo3SnvlFGKZPduwYfZOKLD
68YUYHtbt7UhPJApDVlf1V7a3g0ImF3FZcs2ovh9ZuZl3dTzuKOFpr43J4gndPOIlU0MojwsffHN
7v2kiUAiNVeVhauxmhVlAVf3QO+Q/RiGEj8pNgLp2mBzQQNJnPRPGSrKvhHMB91/br0CDf5An0Js
9be9V8aN9dMIBDtl0MCDwde0MVXuKAhB/zIp19oW6dSJsBHlOtCpmf/1HG99rC0AXkU4E1Lq5nIO
V039zrgm4wfIvG5GdXYQPwD0wv2o9twnsE3zikoJp4LYo9zZ2onessjCuj4MQj9YaIV5G1aNavwl
puydyjuuZFVIGQtq/WKEvUXPnEnCjk9OzlIR+2RUorDRCHCAqw2t/CCLpy+GiJ9sEteeIEGblZFQ
QZqFYj2UDHLKvw2kfwjUNi20tQPfsCVpeI1R0Pfl+MAMYipX5p3k5+oE/bIIeG+QHYcmmhvtCMDY
BmcpgnWezyfhADQ4aSbrEcxs3H0aCo5frgCqj1C1ERE9a1nJy82l3iLeGqt6FnU+pQtc9Tdoit6r
6r1G7ATnCHVXXm2KDIfSaeqTgKbKF/GNFGYreXG8cvMAnLdPJb3c3JBmBV8Wj7ienfZDXqiApfEB
gmciq57rcEUYxBd0DR20+cJZDbSTRyDu5yAmmLLBpMqQDR0kgOME5pbDKMN5TbHua+30tCHQYeX2
DrFkgJTOa3WAYD8JkXg68fJwnGmJs0m9jtjbfIruYpLHoszSz6Fzc9antBRpfEvHmHHN9ro3ddTZ
ZuLs6lxezvIdMBUMqDtK34gemc1V1VF2AjkqKrMJY135oV5h3CU2LBpZDqmc2LBzW9qKPj0nvN3L
RHs7gpUkHgBmcLoqIhKO8sTGycV+NBM6SBLAuuBqo6gMJrM+JR5QNRcjKv6tk83d3EK+mH6SNeP4
7O4itWaBQsdNW9JfRwCyWl/jhnwpVSl8JR6eGQXrZ0LX591//Fy2+/i4JERWQ+o8pFHWNte/Ssq2
h7M8v0RSy9cBVfgQhJTaXOshDYtucVngV1nbTRh6zLjSnKP+bV1U46igql24NnnQXER1s7x6VG5k
B111R6zO3ontPLjXw1FQhVxYxrceAezAJ7KCHT3XBs6dhdiD28aKpYlxKzJLnxRE7M414XSbx2Pz
nxT2kg/S5WoxLqG0hALaSg/dZ8/3C5q+kfmNBffs9jrLRVdwRHpE16oIuzMKHB8eS068yk7AypKb
avXngM2zMXM82Mhs/gUnuH/EcFcacXBwL/4Gw7i9MkqjXadMzbhwTP7VI/jhVm/h3Nvy0xfbdT3l
0PfKphgFQlAmRYJoNhrIUdt7FWLcdKsIrvhGj5poNqwd6/GcIhDCI+XJhmoXXlLtTraMGWxniMS8
cid7BHh4i/bv6wJzXG1teUplEAwhFTVo6OoqjeMhoB8TfKdVFeLaoCUXOIUzGnVXVv8iBMSsrdIl
5nAQ2fK3BqPx/UWGog6CgitQhuLvF9g0epdCiduDKFltAp3JnZJjYR6ZGIlLH7Ew+83yoCrG/h7E
DXnOz/qoQYWi4sDkMEBX2A+gclUWcWp2AJIlQVOo++dUN0XfSevh1F5IOJGw9QoyvTqJANDecWuQ
QGga21cwHHfryyCCMeQwZTJuyjiE2K6f3NiZ5qWoLgWgSvuVHSm5Z8HSR+M+x5JLmMZeSAdYPGiI
kLnKESecP2fNbkp229195tJRhx2YHGbqyg46FmR7k5WyKJebvvQCtnSyqRP9lICHL/0kJzL3HtvS
eZXnGTk8SXBhZ87Ay3yv2Pk4uivnffszih3ms66Ho3cXR+ah4ZoA7AahVO9T2E9PbB8B79ajPLfE
+NMYXAEC+MDjwqRbtXJELMhBkXmpBzvfMSEjzk/Zgoua4dJ2EJqck3+cGNxs4/Xkg+tAzPNaeEr0
zipnlnDQj8Jp9PsekO1zUf4ZDaeBcW66+VfopsmR7RRfj5/SJEalMTgdm1+GGJiR16ex1KIjAOUH
q+CUyg+DJTJsnCm1ZwGTCAPPomTrg4En+roHFVD/H8cAMnMjk3wkZpaX1czg+wI/ZkyfD9bIRFTI
AOSIBW+BIEMLpq4E+MfmBbCVV8Fdwx6nCmAo5oQJm7JlFPkEejW2pAl/T2a1EpEg6tkwuI/NViIo
zC6D2aGsoL9R0vTgArkztNpHH6ViTCjEWJ8AibsJL1jMsRdwdwzeIpiNXdQiHp3WGNk2ZHI+dgad
hniXCPTSFN11CBVZmpRXSUIiI6YiTKPviZO0etDOTFNcdrdMIEwPxr1zybVhRS76zKSalRlXwiLk
WAFU24P/pVmSaysttrxsgtCHw3tlt3ai1N0n6zyAb1UNNsQV7/OzC8BRKT3oQLf7+26aWuLdgEca
vHFNR7/0sEBiwz6Hh5mVGqXGLi287TQWUiIAqlHDZythhsOXqPCuKeCKL33HInx5tCogp4BQm5bR
5rPhHhwG3+n/gOeikggGTpmuuW1x1rq4RSbZvZiX9TuHBqB12TLNIHXPxRPZWviibUvi10UXvFjV
BpEPL6xGSmdb79O0ZUVO+jExLuDvCxulznZZ5QucYOKBEVgTEdZRCRW0wXJvwBUZxgLHg3Aw98QV
0Y5m2mWqPz4UYAg8H38dSsTQg/uvCDfWZ/QF+js+dGiaF3BUwy597gLcy6pOP+w9ljqQhCcpOHlD
wEKgQ4oFT39WYKDMULoQH/BUIder4MlHEiF2Nw7woqF1M2CB1mJwxw+9cUc9u+7ziPqlYvMscwsv
4m4Duf4DtEpWHRn/o89yMHwCcl4rDPI9acN5M0689Q/QFAs6Ih9bWxjgxbpJrQkm3uDdnJYLIBMC
QMWFevcScyqgJt5wFjV+2NDApbIEGWmzHXYsgVP4E7OpI9Vqs0rojVoVFJtkmz+90RbVJN/10XdX
ewnMoCknaG1mWPg01D6jqs7qDAsZFTrAoFryUJJtRznuwxl4wpxJTIZWBSAk/QssRUzHXHv/4WTW
KY8S0saPDHdGUuraC0ImDRxMP9dcGYWD2nks0uEerSij1FLECYn2pdG/IwE0efgI0dYiuyEytSno
6wKaoooM6p+6AB9pzGm2iCsMBEcf8IcMcayN+BtBxssa5YhF6dgGJS66QSlSJyV0b1YpgG083fGG
erSjv9TsABi7Z9g6IE5SQGmqpMRbSpbI+Zi/zCbZG8Ze6ZJ4DSzTxcwsJoW9SupXm8rtQK7KAYrI
tHXpHxwfr9W8PKfGRPKlAC4fV+p5EWiMdR2UKrqjhPqG2O13qhDTQLZC3kfwwArjTIAqMoSfInjo
cizaPkpqL9ibgTmEQGCsNTpPFNJzp9nj4FPIoALhTqL7luWCoHjV3qXvWcULr//X4hbc/Qa88GMF
S5wO0yy0faRmB/LtFjjm9bmuqBjrxntGBEC3WZNkuI2pZqb7ujbGi/gIfDRdMNAyHrd/eYutzPSE
69th/eYUbuAZq51jLHsu8TVhyEiJ6qnvKL1dF8Ug/QXQbM+aH+Fi1xQmIACKd6h8tGDQN/xGMLtM
puB2f72m14KYW3mrum323RqLJXqYlHauQqVUetTNxYVd1NO8cCnTBZu4jnlwxdGusaLL/phs0hfv
v0gRpC2xOuebRjxqyjVBrGJG5futEIAcSWrXcLNlrhgtEUfgr8dcU2Vb1XFNF06LyuLddN9s8nTC
NWAi7QLM7ke55bryLT8o0m4lUGfeehLD6hkDRp1J/ROayzyPLIr+30oFqyHqzT1dUwbUBGMMAEuS
IjirD6OcmIGeCSDIuK88kKDp+oGML0vmglRYb9uEyUZfjs0cZneh1bDa0DX2TfkE3tzzI7mz8Mi5
sZf9Pn/QmXNZZLdF/TSDeArspoS9dtHwvd0FhFCpkoxqV57C7GPrgyhpj3Vjo1Z5NjPRLEl2PHrM
ur+1XT6gI0rnUmxE1Gzibspy3rEpeCPfTRlyqVEhownaU/Ho8FjD969PoAKLOBMwLGLdsB/ChNuw
dme/UZyhe5jbAim+JVPVmWxExbs83GPMzggmit/h1RTNbkckFpAf9EIu4Go88lm+UNNg6q39DCYz
pVMs+CFrv3rxOfP2JLOTfcPv+jy7EpEKE7FBuVzcGlBcp4+Bkh8f5NDkdAaU7XyLcKoUYfM0u9O+
dztf77xQLABKXEyFQd0cQOZm0AyPK36OiH0z0q6AdGpnnUmDccbm/JbR01/+Tbm/Ub59ahbY13ib
k2sddgej7tF6oXw5zmO9T1NUetkpFXFYn2/u10b37zyGVxFIqEZnODmEtzAiI6n6+tDiGTmf8htc
kojvNmcTXmJnMyZMREEZsGrwPkGDftHiEVNN6Z88/Zl4S08SQN+mYgnRcJZcEAV7roZBMOLP9ktr
a3FJJijll4LbokXp+onN0eiJrshzO38TEBCb6ip1JLVYJXCYoniNNNDsYHDKEySKrS42oRLTTrkC
KpoMXt2vvyw7GHQVc+TsfOZIMDV/+C0pVgKkPKmUhZis7rkfGXKMPgR7nBbXbBCHpMh1yjoS4fls
0QaRshr4HrIOQiMmsv1NESG9V6v3zRCnotp+21cusQWjix+GwWeeXi+cy+hScjQCvsgwEqqxlL36
KDSnF2F/6hdY9b8pRMumiprsrz4ZVEn5pG+Vq7drBrkHsxjTFiLb7WH1HeWG7RaJHQxWm3wdTw2C
DEYyW20CQi981IMQM8ohuAdGUvrvBl56zrL3uMLXgax1EJDYiEeC0kv6wzL/Mi3tvRXxsGRV0k4N
MjPZZdrYPXRBTrbNtQY+cFEnAf0GTQ+ekhwN0TO1yYBwDTmUEjGaLJB3iF3N0EEp54fCvf3mvYwr
6lixKRpIlMqBaoDaaADFbdMBee+qcrpZHYBV/V86nW3jZfcQ0lEI33nwKWFLr8XBFJklsIlcpJBC
huylHBlFWtGTZrYkzLfJBKM9QvVMWvtw4gZk76gFA+gGERcI/mCp4i3qJB6vkZxa6YPKBHSHp3C+
D0dUdmjCPI676GtoKDFOUaMou7HRD0E4B6yVMOS9ODj1aUIcb83dxVzDwmdNFTB/lO+/kOKN80X8
82uM79u1lL24inEneaOwmcHW5OUY0Ny7yx6IKzTwrFszT2ey7OhzSuJy6yNkCpUsbT3Ew52XXJji
ANBFXgAHLaVdhVjoS1RZMh1aYwHuLfbChQlmNA6IPp/+wPEm5Qg0xw/VdbugCdKinHZhfiiatYB+
OAccGKcKtq1zzhN6T/fYuJBEMKxnGzNWcmkomjshnkEOMhD+phMwf8YOjsH4YlrEDycPCU+nxFJM
8CzeIJwscRDYPnas0PKG3IXWaUt05sDMlFaAdf/kFqx9OncpSRXB7bBvk98hsuSQ10JiTERgrngQ
dCkYFBY9XokBrDSko8AnhuwR2kqEbUsxsSLDsCCewbxuR71m6foFUVSiCnw1gkIytGS2/fH5NBlA
ePSDswY9CbQZ3s5ViDXbyiW9TOzZPeD9rLV3fHurScO1rlcrXy2wlGv8eXxA1txjVSIJaxgZE2nP
EIlsr49moMRSMVxlmqyeK2+71HAifpIm918MAzYdXMjLuMgohWLqQfGmbEYtjHNo7WdwDnHFm4YW
1sDYU/wSAgnNcRckVNieh33fU9fzVET3jrxpo5UjH1ljZ+HZpc0+VF305shSZmtEXnmZvUEFXMAJ
Ug71IZcA6v2k84tZtjr7ezs7Mer08tONJJeTD6twyrf5gdXuVqdx9f140/cHHdWBv93kmbLGNazO
0fIonk5vTNEOF+a8q2lvNYFj2ebPx7BGyUzkEA896fbLLavGlrDY5A1u0n2yM3lE5c7LM/amjh71
yZkYYrKK0/fRawz9Z7rktD3lIYnk3I4klyApGHFvXgJMPtjm/IMfmyqykH58LPRplsHj5r8UDQzB
AAbEVJT255PLoYyZPgcG+FLsWgJOGWTF12RMxcKfgHlAlJnOkdC+GjHK1A9jTML7kgeYlHPNsiox
y9oi37TjoX2t8pMteggDbMjV97g1miHT9X+GWDpTV2EBgpo8Ad9sG+bogWf+7AHLYm6Q5QmjMIQl
UQSIl52d6tAMT+i28stnoDtEatx/kuniujhg0b/uRwD/FgzrFysLacdUVL6p37lc+AVWlyEOrQmi
gvdhhQhYPfLYlMzocIvILRpYwAptWcsMBN9cCsm7SUudONRX9sBjVB/dh7pAbRW9ahpiGeAGHGPa
jornPtrVSCvELiOjgvvoOaXGSkYH60kzst60rVaqGhgjZMeJtr4//4HM3jQ06H8DGcw0g8rsmPHp
FtgG6Jxh72XjunOzjp4KDR9aWBNmSMJrZVgrRCgNtDmdC7eHnS4P2uEL5ZIwDTCeKyvjYCqaXzHL
btzsm5SsGEFlVLFMdwASCgYJ/KDi6T7IJQ+VHG+w4j8oCfgCNjNKfPR9GVDBFsAx8n9KIxC0hHB3
xSccJi5YKLLuaA4+rVkMMiKar3OpH390//L7eQzoRD2TEuVkBKHsuhres0Hi93B8121ERtnPAWdg
eJGX0pxGawmjEF/NV4BaE+TUvT1EGVDM5jIQFmf7JFnSDnZtL38j+rqBveQMpM41rhKfeWy90Sas
pS35YBZQfx2aVr1qRrGK7ix91P+5zio+WOsxGkHRIcU7zZRu8IQm5PSqbtkxWOS/8kokraHwUd25
2oXqseO4bgCLcohYQsWsg4Q2rGOkJOtbY/lIIcKmp6eYbuH3UZA7kH9tVClTizH82YxatNhTDP7p
PWk5UH6hZYdGBhuyjI1uctjLyPpEBYutJ1ldo9+guTwOwecLx7BIxg4zw0Ii79JDDeu+WYBmSNnx
Q6z2UwWSPa/sqFTxoP9sk2BRfztLT0SzdQ0mkmcsfyLNwVyCtzfk+5qnGH5ymamojFN/SSoxL3xJ
OvZdNS5qVi0hChlsAfs/J+QFjW2qHwVWhbboLB9rAspduPclasaEpyHUDioUwT7rQYof5+UTFqXg
VPggB9dzCnXzYKsnHi4eIZfbsaKeSfY/jvRVoyYpODY3ujP97duVIV61n+1ISMOJNTfJBgOhbgeE
WvnpYbyCG68MtW2GU4Ca4SMjJB74c5yh4clB6xMF08FRmVemXaFApxdR4peY91eVvi9zZ4T8nVgV
e9GjgAjV6tuu5L/Faa6vqqqgCcWJhjm83HX4/0/cwjAZhfYRY0ZcTsxH9UiZ3FSEY0PiwUotvw6u
Xh+p8f407h6U+mJWPgIMLmBTTYQVl73GXh84Kgs+O58LcNDruoZPWn3Hi4sor8xf8u4zXdkGOT+7
sdmCN785XtyKhxvtKXb144LvAoZliEpU83zZaaLcGHAuA/XLoY+Nj4cAhgP0j3/E1y3V7ALZUIVs
B7iXMhUya8OnyIS1vfVXUiOKCWdfq/kyyi0++k/rR06b0d6a4HFE1HwdkuriGeUEEjB3EjsQbvLj
NeE3I7wvNk/R1+X20a/rNSnZI9ZsMJh51/zbnO3Fep+17/owkOdxb6ck+LpysMI62vojjgix4iC5
9Kl3AHtMqVbUe5kFyqbqYagV3hB1LCJ/Q7mp4WvRtM+K4V0c2CP129sksNqqHQB/MP89XRIiGYtg
Hc9nOsCXKRtEzE4y2VFhbZmxvyvn/OMsYU3NVKDBlJs+Sx+b6cBcbH7SQUGDdeFOvjxa82y+UDP/
zQLHq13T34rZDDrFLNdYR+tjnqu7wezfJVPnQySuIiSs1a3RYNu+pefZzgBvRptSHQkytDypSbJX
5VfcR6lkQdfzIyvbgtpZnzxSeJZ9E8J4vuC1FJVIqdu0PtRganbBgLV06qEeXwP3HsPpwUJ2EhYY
/uJiQ7WsJdlo8QWqVDZjF9fiEDjrn4jthP0Kuv/trZNJlstlZAAZ5DkKhHNnn93Wcz3rKYGo7MeZ
dxC8MqRLDkn26NZHNyxZR0LyitE+0wuvBmQ5ECIE+5i/puYs59Z7fOEFfOCiwfbWMx+f0YC8TGkT
uTLFX8OdIoQkOyUZ+5Pr0zCKZkGIQ62lPpaXm6WdV3FUYVj68uemhnmF9kCfwxQNkYBg5QvjWBdM
9poCiqCiHycbs9KPtzoNebFgSG7eDg4avcHhgjO3LoceM2S5xrihjclpt0GZY0E8DaE6QUIM/Do7
8F+F6R9/BmBT/hhon8YsV9Lp9ECnc94PRsTeqdm6EN6QyBXMJu7twrMtE44Ts8J0WhJneziw7n7J
iBIZk5ZdtHGPrcxFV0cC6W3RwGFKGGt74KyuB6r469VYOvmXKLZZhHmCgML5qt2YI5va1NKaMpEl
UfSnvyvQ4+GcG338KWlrx7H9f9CAdiUnZXQy9a020YvnbSLRF5UyWrQpWMPcgjJ0y9cUjCRX25gU
e5RH6ByXfVS7BlRr92Z1OMNJ88l2VhkYGew7kJeApEtQ9u4FGcWWSt0Dfx2pGrOZiactPxZAaA3c
tv8DKP3NzlvqhbyQgIQrZni+9x2QYLA3QOPx0+DiWUp+R1Li9xgGo2gjDcQuxmtWscjDaLDZWAR8
Tasbbxv/qUUVrdAeBw9jcLEPvDl0nytkwdNgu/95A435DDAOxAHVLJY/KcR6daW20+6gG5DYH8DA
NH6Yb7f+MDdR9iobBvSozwZg3cmAPT4k62ljq0ylG/+JPusN/U2DnGEjkSGj4i1cbTZytnzRhOVN
pl3Wm837RSH/+T1cepd1Z7Hytn8PsgxWQeXSP69C6WJ1/nDaO0l1ZLP19XBWbBKmEiRjRuFRy1Si
xP4OgxtO5aOWTuff49VfiYWcrWZF1z/WvZtU2OafxlQ/Tsu0gMjo6yu4urvFhglOF13On2UezsRd
UHa+sKKXzvii1B3jBrc3eOCZCx+PxOTDUc7chLGTNBB2OzgBCLpIUj+t5DGJtPk480GuERkhr68+
baWWJruFLqr4Q7hYaFRS91A+ArcFvaSesUlKeCxBF3n9U04F6y6yGqPR5NstCzbxKsRN+MmgMrxL
Z8ft+d3alcMIBiUR1OxuufXTKFmmSgRMjfdqa7rJ/gQlccEFtvhDAlltWEq2bQ0X29cvT29ZuhLs
WckRrmvELKHM/OrfafeHegGHKqStXz50TKw8XWl/tkW5oFGa9vQUMt5aqwfuPGps00S8wRyIUmcJ
zytRTG9til+xTTGPeJRbuk9qL6rjTI+zmg/WTdGEPZgmeSMdo9kSCaPEyAyAVrTz92EdeHDwsl+u
K51qwfMIXbR6Ai0xiQrcMIJhYZaYOLwkfHaFZfgfnT279aSOs+14wJHyD2cJC9zILJXkPJgWNT2m
5cq/iDf4t1v/udyBWPDJiHZ+rTWDPYkQ66n0xA0+ud1TkTAxpFc3idR9lMtsleLRV0MyB+BSU03w
VNXwZ998CI8H9V9fQDbmVYnxO4rnq7lTYuZgJxqVs+ArEEANcb5z6YNE9+IEVXgUZZnrE4oN/2iU
yD8BSS7X3ktoiwe5Sx6oSSjjK22uMSrg78423XuU8UjRpDgkqYOXaX2x8qAOiLvod5aCoy+fOPVo
bYyZdp7fZTMv9ZqjR4kreTh0P59RaqgPEqRAjgqGg49ACIiw5a/lDubUYVmXmL+ozMDIKguoNsGL
gY278G5h4iDdx9XeONxEvVo6gXk4KTOHtR7VzrqmQj8gLxxfXr1laAhKOe+KZW77ZLVO0RPdVK1P
NZyY5V72gW5UsE8QRRW8RIGJdyNyOHPtE6rSFULu2/SM7/+GckZskiE9gJB+fgLV8nbGS/1x4zAk
2sMB1vdzAUeko70Sc37OXg/hsLd7KIMI+qlNpWRbeoorem87WK0lt21Wujto8NwYw4TQ+dN7vGz0
ykd0IBhkGWhXOa0Va9b6Vwq2aDV9CUOsf5nEbZfiILirRLJPQMGhts8Vlh2pEizf68T7Bm2bDLgM
EkMqIpOk9kA1Al0U/EgDMMdJwUvkJSr+V86PtERz6Tv9Bu5mNg6mHaWdieadyrRRKQ2D7W9mwNmw
hry4SPW4KqNTjjw87tDxbQk5SjeE5cdPJX5mcK/Xayrqz7UQOmfehTxwfP5iA033ruEpWpZJOzcb
CRQchJR/pTN+okq1PAj55BC3XTxm23sfpbwOWvgR6DHnmvUSpXgf+k4GTzN6HIty3JT9p3iimxj+
q9Dw115sJK3kvC9IhQ+AdVZ42WUOhoOaAu/sNriyPvF9aAbRJ0l/4uAa1yy1e8OysgIrurWG/v7m
XmBFd1r/BqQpLRzl881YJhQkzr84zp8uFc3S8cCzD4iCcDV+wz9r6mBp5kSAUSUkbmdbZSks0X6R
4eTPjhniUmrPt2ke03DdJ8ZdBH0rpXfMzi1s3CvEOI6ReMTQMurhKv5dbfcYuNrT6flCIXKhLkWD
nSgYY2IVOQYQV7XXTyEJavDV6+GIKYMMsWphnBVy2TwfQkaCYueIQDH3Hh3ID00wC0AfZ50+SXyR
K/S5q6us1+dOCSA037TveoAZsmGJfifwu44KxtLjTHD0jYFZQgl5GJ7X7z2A2/fbmobAqdwm/Ls6
qu5+xT3nFXKkVoEqFanCEzlxAXNK8vbjGVoifnOQr/o3U0Kh29YW4X8ewErgH+//UGwPsJtHQcZD
RVKd7p3EBMOn9e/oAjKl3Y9iXxmTu+Uv0fwiDz3KqB3jRbY8dgNPxAzM05ZGC/gzMFrsB+Edaz3l
3pcM93+TPtlTcEx9fg2UvnSIUNouPaarh6+d6tyGCI71uZxNI1TjxrpYnt1UxVt0UyfZOiI9rVR7
m230yDSEi7UOyA0yASgSefs3RBx7/5/b53nCnH0BKf5zDMLB3t+Hp77PkOrd9Lt3fsGhJTCaHsaL
7jXRXnsCekAn8iSDWBFMpDoyzBVqCXEH2ESBB4KNPtJT+oypnGx49O4LsDr0mp1cUQLBc+4tKfop
PJk2J0QHLS95YOe8Qe4tmKyC7NHgzM65tdhclHjstHJhENk0Y4X+DjFlo2Twz045GvGJALR+EZoW
W5nrDUE1Nz/O45n7kiEHHMY/PPQOMeh2UBqt/Rgeg23dy+4tNsNP6XkKoLD9Xy9f7eJK7q83E6Sm
pbGWVtT0IXlUHlc/pLIpiuVgMhVBPEiNxpQ5shh6o2zct6K9Hq3zjuwNGuE7EQwDdQLaAsOItWXY
oNL944GWp2d81FNg6CpShFhJc7oFDPV+Eokr+W+iOaYjN6nZcREkcl/chjjqzu0/MBWqS0s7wCHU
uhIRx3kgG4yF66ENs9Zmjpsc/DKaOI0+5SYgGkDMYGenMCGgaLwF/P/E7gtNhqLdA8pvGFFzLgjp
rIuprhwwtQHV/QTKp9SJVrMnhkJ3+XPcQ4u2o+eH7ojWp9PodwIHuJPi+vYNUXWsWeoTDbw0R+TP
aCTB6mYCSlDPuD+RIE+u5u1Jzaj+6eF0OaGTQS+sHaxpipqCubVYjUX6w/0Gbo4EAp0/6LObEGAw
xrRuhMHEMxjwHn4LesgYwGvBozmArG1sxqnIM+U9NYFcD7U+rtbCV4xtloUvIK/W7VZgi129ApC3
9N5qc4Rez0t6GZ4Djuj5XKfHp2qL2920+ZebBJBGOI2vFwjR5ksMnaZg8lsdFhrizkrL0yKVQmAQ
fTpG8V44S9CPbix+rl4jnx/YS7aYn0IVCUI2Jy4os2mWNJo5f8IbCOmHKXwjFsOGyIoY8gl3rpOd
bTTMVGtklQ3ZVQy1TbdsrM7cHl1rtY6tAv94sWrR+DOuMLAI+gXlWNbDJhK1uf+R3kC/pyjhg6Ig
pThY5zGmrDc3Np+Gmm6kcZ7XPtmonr4Wc29eq3co79cEHoBGCy+y71/pJcbscelnu5In4DOdpPK3
SxNjWHzuYhh3AS6lXJ/vzneo3c27uHn+a5zQHZZcWsviRYDFi/ZqZ0oPhXiwQH/4Cl8ndVLfyVrx
IG3zt+R4479O6BaKQTVklAl9BfS2LgfAGjS+3wa6otUM8TgAFLPHaTLF6xVQeivaRKzFYLv22GQz
0lSo1GGLEMuknwe8zFr9N7zCrIgvJSgRDC79ddGA8vhscu6opDVt/BZ9Z6kv4KqCKPBfwaiXKGa5
hG9ArPel1qrhj7rACaZfFVAaX0xegE7zsZk82gwR70ta4NVTaTGDm80wN3iW+RM1mirI2E6calQv
7nlSQ/UBUSZQigz1nrhllIRaR6gUFBnW1XfDZXSkC1bHbI331xuJZ9OPDGlX8CkCpOaQ5SZkjumt
HKKIERQ8FqXzYRBfZ+Hkl0I8ytGpB0n+ybr37gBQZLwgZ36WolEo/IbTOMzbRZIuwDacMTU7FClP
3QFkKRVmPnxqrT26HwpbQW/vnA9wQUYBb0zlvtN6ujh+tEhhav9Rz1rxcJzbwi0RKrWKiIFNNelB
Z2q8IixmjGz/phx0xy+eEqcQFmKrmNRLFr3Ck3ItjrVfqjGWkNGK7kX3/nYXr1R+09qdeJkVzILN
m3b2UB1RUB4R4ToBCt+zElRQmHEDYGZUl4s9n0R6vjNVJLR74av3P4J297ExU2lRKyY0yA8V/gXl
fSMaOUscBI4kkZLqLYWEBwP+9iwNFeFMykZNEJ8d9Z5U2EM8cUl9DiUU9+JlMyAIGgPz2DCm+UWD
a2rxMAWvJcDAmBpXwWJO79jaxc6rI2FWR/32YCQcITSMuZyEglITY5ccDJdtbcY4edF9Q0xWaujo
1StKwD8nMBJlqzgIgnu0QiPR1WgJvy7cgCScF6reyHoWtX5INnpnurMDPwi703UjCNjbnUlrPNve
2yCvro4WDsrY/s6iD5iA64kBha0acJ0/RfQV+RG3GuXK/w2YFU2lnnUlF6L+MZsYI+B3cfN4LG5A
K5E/AAWhV/2gp6X5Soq44GjyvirLprhewIcpf8glmsuUD1Jez2MwNMx59lRxejfemUouHsNENql9
D64+PVxJe8tRSY7R4xzZ7c/Pt42v3Yhkc3a1TcHuYkoRwB276DsiP5W3EBLOObUel/WP+eZif3Vd
cRbgIVFuJC6ie+fzioljCdavW556ZyIc/KUa2FonihGYxE/HatjfrqMV5kVdZeEj4CTr46NcmKUy
07DlJa+3K07U5o92s9fG7wGnT38aIEgZIA3JOUvxmmfwrOaF9wshcLJJDWYZDfCIcWPaWS6OEOM1
ZBt/pd3aUIauQIekIseS4hN+70eP2AeiGzCpP3yxBOEtRmJej7zCDTBd2uy/hqaWpKVydDGhxo1g
J4nfu0rhUlGfWWxZ+/Janzxd4vRbrqhRueTq6d4bn0OgecnnoqIsqdGpd+eLhQryqOQa+6WIEvN+
JdAv/nl3cX3Ddu/1N+6VX5Hi/ImwapuP83LZHtx9jPKu/t1VFKddN2ch0dNt89i2huZQpl9fJTVi
Cv0DD84i+T5nG9kMZ6IEHC4DizKAk6nem7a1k6KY2Rux99sorRXu2l8DMr1nrLBTNRG4pOtVBdDc
tcUjroQu+bN2NUKTkBvYyMUgR54sKEzFgXQsYglBwRuKh1qWVftk/PcIBx7hNHRCfw6grud/iKT1
bumd9sMW3Bdt0Dt//k7Tv36WM930Wp8fxhz8h5RdJbglF+TKkaAzGv4rAy55Kz5dcSTZK9ShoSvG
s78Ga/4jWj7si8go5AmFySqI1lPFhVNDhXWR4Pe8DMGNxqiSzb5U2xlc72/JeoIKIIOrclzjy4Zd
dXOtsMdvJuCUOLqNLadOPpf8cNHYZT7iPjRlEg26L8fUtcnTS3FXTAXEPS7rjdrPENSdFB6+FKjy
5tPImCLANXAjOHiOfpaQEIKaIl5FlyrYrTtZVSUBMs/bf5XbwifyJt5Vu+WAHwn5pKLXg+ulTwuA
Y0ZW/Jnh3rN2tstLzvTzqVNOiStjWz6gcwaBuzrxLJSFmomBNctH1xQp/dgNA49hxQf7tKzB1zIw
qxsyvfhIfvBjjrV4xbrtlaCngkCWa1LgWYiToc3QeXNLu1VSfhS+3yx3m/gWIDucxL7NgOd6kl0A
Q286q3s/B+wlF1/vgQZL5vvKeyc9B9/W19b3oUo7hb6qtpSi57SsTkIN6A5SgMP4RsLbjLkJ/aQX
RJE48GEvrjB/97HqLIICSExR9p8IpnFDWpCr5gZ0kdXFFVUxSxZ91pw8xyJf52rWH/2f9h7w9+TO
DKEqjiQLMD+hBIos7yLcAZn7zjRP9VI/BRiOdGtYp5PoNAIWVxvP05Z5+SUD3fUoXQYU5eJc5dwm
XndQziNbw9w271Q6fzoR6kFH8QJfEeDbwQM2dVK5m2vHi8kml7sUM1DAA4nYeE/LYs+kZ0cdJ7Si
LIKcgWFZcJTdeIwx7dAi1sRqvaQsYiNNeWR0o1vxM8jq+Fvk1Z7KWFPCcE0Keww5AYuWUScarRqi
MY18epwojsfcqD3IrDFuYvfV4IROz2BlwZtJODgwF3QBLExbPvlathvFslB0TtNeMYKRAB0z67x6
pTlozUpEOEG27STos9PUrucc8MVvxn4BWXpGf8vUjePBvGjB3lCEzE9JGMv9iLnpAYW/x40wLMmG
Dw4AR/CmrcKW9GJncORnviP6Bg8UafpGVERLjl97g5aQiun33zDaqOhPqsrNkHaHwCRmTPdC+VsA
fSDhJf/x0FBGbbK6OQVqKl5kINy2Ty6s5id35ltGkqxMDxGxakMyq5SuJ0vVXbVFbmgIUWJH871y
KzK0VrhEqJydtf+/12gMSoXbrBzF8xWcFjkcC6P5Zg1Pm17o808GuORuUdBpD2mTlsPHpMeXSqDE
uTHnF8sYgPOXUfkILmADVr9x8gigxzGcs4RRW+ejqGgHzC2HwhemHnlpEAjWPZf47FBSldkiugmT
XP88Opeefn4LyTpNdkusUwhml89UZ6hdueODpMQi4ajP23536Oo78mbC7jTCyMcrnH29zx2+Yvcj
1GZjaAep+Y1EPhao7LzPgYgAqsmB4x4hh+d5S8rahYOXiuRq6HfU+TnvSR7nziG6v5puqaa8zv1e
m8RhHgySEaFsfF8Xx341DT9mFc8Op0xveIIyR5bPMhD4i7FJ6nMHvr3ALEhHfOwEl+lSiYtwbnsN
C9CrDTHN+1WwGkcbVZepPwugdi3OtwB2Si8LXhnS84r6sBGWxIXxCKHn0cfN/YBb2DwQwj+M16Ly
YxlkHSyl+K/MFKUHqNtoC/aVbGIqLl7bhe9bQs790Scg6M1hgRZy7jS6i13KWuSmiQ9wBuWijvSy
4uj3pmMXYCqMWLOZ3/hbjbR/TG/oQRVYsPy6gvxwYEiYkWU47pHbvbVf9gO7ywOwtj6HI2ow7lf1
FpC2hmtPfWDQetpOB8EsqG7bsMEV7hsM0dsJJQraUrL+spDwWAimnWdwN2O9rQ6aqLalF0Ew1dGw
niWs/UCGYxRIhYZeLb1IQtcbXjUSSRTxRZWejbyLR94fkvASpF/Wh7CzVf1qBiNwYUnPp5l5oQ2B
XA+44x7R9voxFsP0U5V8lKgi2X9uSyQksxhStlp/4nTWU+WHOgTrRKNWjVUPvlpZZQaKb25iPXyZ
FrnOkl3gHAb7tnX29INYlQ9038ot6qi5wGpbD4Pd/Y5aCmTSOLXlapjgABCpU9T1Tja+ar3+hzCb
jksLCyx0cogQmVZftLrc40xjmgWM2JRRtq9I0wFbTsGATGFqkUKhCIuB1UsmoxO4mvoszbOaoFZm
NCry7lGqgDU3rbRSzLk2Ub3p4q1MghT4wqtxl1Wv7rzu9dLEqHnYA8Qq+uARqQKGjxGF8BerGjvQ
n87JQbRPrprppc0zZI7LQ0wkPJsJbXK+8c1tdN/i03Z79rQGH0MYTirfNrIvLpXSq13qd7kKUJm9
uuhr1yjhSvDBEmL2ctXHpAD0aMflKq5Uil6pLVa9XGn9Y1ydEfcS+scqECgk2f9GN2sITxbnaBER
y96AmMhGOnkvrCDc3U4aY7D9kaTs+Fo60UklqLDDlulIXaeeCDNbe8EhF1cmK8G26xf9nogmTLEe
BfxbUyY8jyIxRjuukK9lw5P1sVIURlOsPlMpXSuT/K1TlSKHqatNar2RlEN5o9x12krHlQ/aLXP3
tVq/L59/2FT9EFwZdBOYAuWldWIKE1oWePtiggHMOAAmFPT/d8YuzSHAFfGk0cOBZAIShJKQplBV
ACrAx+EyPdL53QOYGX99vM76U8p679sEl+GpAdlrbOfzQrbj/z+8iCp4ovNR6o3Sapznezg2sL+s
irig4+fBNxWLybv4V0hD1LV1zPzjIEsaZ9GZ/FOYalnk85pvjHHuGTCLSPBRRW0jjcKSduC0yfZ+
0v2489g1ZehECR+zOD/crBSPOxJaRFvh+5+USoVQQ92hGWgDeU8aqTeOZXMcWs4KH2PuX7CQ++Br
Igbhy/BOggiHWZQCkB0T/2lJhZAmDkxXM0Vk+p//5mC9Yoa584E+NCGfGxxrJmwqazqZkVIgRDmw
DbBiQlLPlSmh0gYJ1d2ytK7y46DpC4Mq3leUnBO1Zt1kTen4KjA88WxDGAbLyptJzr/i+b+Jk3M+
GB1QwBtfrHBruwetB3zOurAmsNNdYJkn+jkThl/Kk0J7lvxo9odpYUGZXyJVIPy16RqhsfImaTW/
1KuJGophtgOtyn7H1rzve/RbfGrFfHyxvDgrZzmKlNaygvTlaZa2Wqf8oxRqYta9vpdTDyvlbgsc
Aii8y6yMAatquPdO6Qao2SQaGr8mKSdGmCU6jrRmhpF3O957JA1/z+kwZEUbt5I7Ng1Wdn+x7hZn
fMerkokXxQHBkqATx3MmJ0gRCjcDtyJ+vyrLlGch4WX/PcyuHAR+9J0W6xF8zHITqWuMqN6u9JZY
qnaXjF5U7VtUD5HhAJz1K5OhOKmCLDzeHpe9RmZbuNO7s+RQrSWk9DN2tRwOA5CN1rMHkjGJs/kN
njkQZJvkIUJL6WEpIqxfCyJjR6UUYmM6tf1qJU5d/Ofp9qB4BYEou0off7SF6oAjr/ozFrw39UNr
AUWGbpjc4ldRoOYgW0GiSIxqM3JwrRFWqsv+FZGKuAaJiItcY4vQVuXIAgRuF6AnLnHj0lByvu2O
EK77HDGSIeaZGNlYv99OmFlq5yGwLhTHAbLaT5TKRQCfg4GgxyAhb2BCJNwK0Nj2qQh1l1wdaays
4Yhb/PO7L0i3gL5LrQWuyjslEp7icWv5eD24Qo+Rp8VpAMA03TcBxSmVCAjSJOPVa9t72F1pWh2B
E6WRG0CDUgZVwMF6c64WDV+4Vbe9C3OCLJHOBrutXijDteM94VlVks806B7KwJn61Mu0vS6kzG3N
CQL61NKY0rPPIiSLKpLWQ50E/G1lB5gyXnUysqC64AvDjnMQ0MSqr++r6lqppro4dbN66nAzeLUL
FqzLGbmWbFHBe41AF67rIphcorLoO4p7P6g+Kv0XnZ66eGHv5EweBOzxIyKJyk3TVn0x7/CL2vHb
sobZKPa6YGBP4AKQFiIraFt0iAuthZK8y4idF50Km7a8kp3xU6hxHNm/AZmDUe0v384M8tCRY5Li
CMSey1bE3Ge9xCPNLYAAmrs1V117MDKZ///ucZyu5EjaayaLjBRAcsiqK3XCq7shCF8F5bEhZzLQ
55FeGqdMEPpv0/v/qEOep6IKWGg8mEqqIUQMjpyuFttglITTu0XB7O5nNnaFdU/EcqUez1gGuDT2
c2BGZ9OHiOAr4y0vfIvQv7CnDbJT9ubdDbMkbepoTketmrSDNdjWWKO1Ls1J/lOu1hOkN0LK8D40
4xZS07J4N12f/IaZtD/dpGfO785b60zxH+xj568D/OzvUfwhs1FIh1I7XCQcUps6yBBLto2ivCEM
ej/0aOOgojZP8Oj0kPdy9AtYyab35X4NU6/CocYeu36sOUeROcyKbwTxQLNLDQiDh1O9x8Cuup1k
/AHD0zRb8tMURYdpYTgyhCAMq3bGyTHHZEDXXh28Oc6eFoKJHjPmVVItoAknaMUCyw7/meHDjsSv
5a6QPvA1MtM2/l4Vj9dqMB3Nfa61Gu4KKMjvK/UFbJl7W+dPn8pYYedw/h69g/R2z7nQI6h5VYV5
ITHldCjIY6i9EDnVYU/VkwpgY6vBCNn0fnPDEauFIMQin+ZBKTmInhXDQCRCWy0Fth7lRxoHa8H8
Wppy2JHdHZeNUGZVSHkERAzJOmoPYlxiyR9Z3A6oAdza/JBRRVfdAoFv3KwXgRPVgdNrI2BRzZX6
Ogk15HezXF7wepqRFehF7jg46FGv3QLYiEjUArTAQ37iOrda4dico774dKsMMrIXFpkcyFvJn8pL
I0PTVa/dOY5YK69CfyiSn/YmMJ9AiJCNWvaAe6HtBJGIw9v1vmBI/kQERMqwG1T0UMwlFHHZxyv3
QVtaZIfE/3JEHuA0fhRn5dlCeHzUg3jzFkahvQR3I303ZecZyvM3Q3km0WSYHRdHMQvwq29O+Ys0
fRjMUoJYGoaNuPoAEv5BV+1RKfPPrL5MUs6xPMlqmONmTJlkAmTiitfpsFrhXIZdoGlmWNhyTX9S
zhqqh+E15aOoG97WWUpDNn2zjJCnRi6YfrzhZOFkqHhPDSsXmP84qWCByEd9Lem4mWw9AS2O/mr7
l7uS3HLixjaRfN8HCSm7wXQXx/QqnpwTqgzpBuGGGXOx41VtEwiH0xrVShDEn8L28k4o69YCncXw
mKdgJDJpywSWoMylN3p3Vr46uvsXPwli4WKVeUFJRL5h/JXfI21kBz05h8n1hXLMiUYbTYfXvVBV
p7G5Zce/iDqHDa3hi7bfdmpeDJ0Ld2IrRkXTwwUa2tMCzQedUGInEQc6qbZMSZJQNAAhYezgtvA3
0jirTYLhHGEce3FzVym/wikbixL4RCKNewgbzTjOmePV1lNt/6kfAUwzUZwp0wVyb4N6+rS38qka
4oO1QAeqNzVvgZBAbn4B/HI081aUzgVlfqd/SyMwntHhkSypYGfrz8Dcp4QOg5cqZrAnrtIi0Z9r
8V6xLAVHGoGAzo925MxBI4E6+/zCiD8xRiMh0B4fxAs5zWPVNduojyN3dIM38A3Kbq47BFh5xSIM
jk5+jroXG8JhjLtzvwiuZllsOWoaqQh7uVpjCHr2MtZdOv38jj87fk7ERRCQi7Gzfxa/5a4PNBF6
70Wa1b1PlDQ6H5V/bpYXx0E58WHZDbJHxKaaP2ila2jpeBZLkhVCokBGMmvMnAfGtXXMZ5NfR6m7
i4GFoTewivgTTw8CyjpX4lg4Mwh0Ie/dEr3Q1WyVKy0AQ6XuHlZ9ogmYX8lG/tyEmn2QLsRPmmwX
luq6QZ5WJGgqeeLibjNXKYfCZnspqOjr0n9jKYYCx7IVo75OjB+Xr08stETUvBph5sk7IOxdmHqr
Qdf5GKRw+hXJYIDDUq/dcp/Ck9NScDWbr3/VZD3YlBM1e651GAHl10T4Vf8MhFYvoAzie916WHbV
LGTh25cnrlRE3v0x2ka3gX2YTU3x5iZV7chyGF6qAdYqnZyEMncVNcyCAwQqwMaEBjLgJBHQM7mR
kA6f2SedwNpyqK6xtDalzYNUwI0GL2FTdVzWxjApEZZYIaQ85jGRHasgS6lDfP4+8A46gVakeOeE
PL/CSb0c0srgEQXzSyubsWxGuHgVHKhuFKEKCryzIvTvIOT201LC6Gv1/ocKOpAFvrnx9oGkN6z7
z+PVaQRZdapn0q2qz5vt3m/S0WSZCEi7L8gMM7kUKRMg0g/KEoM84XfG093fDmxLQIfaq5so2tKf
fkk8eglHRxX8j02zPIJdSRFpD7pYNKtSeqI86gSXLPYAqAkNI/St4tcN8vMw3jpWWwKBE4AICj7G
FXIsooZTvdTZy1b7A1S7178VjRfAfhn4d3T96PhRzn1gP5yxxx7LNFFBMkPWTdfJA+6t3u1RwMz6
K/thvLGELs9CdaL3r9B7iiAU6kx1yRpFB9Z031ufLbhOBGEPIwCQqrDVvxnoop0XNppHW5aOjFKc
A2s96uDa/CjY9aEyjHtqHb3vjCChmE1LvpikGQe6qhkOkQOoGDVTvTNUo0Th59rzXj6d41TjCgyi
dm7fzKpzJZgThC1OehEtSNWvPWH+b/DT/jOSiQFcOPBSac6bmZqynBwxYUX66J+ivlsTWUWtUOQU
uNCR+9BGWhKuQwf4he1z7x+N3NfIF9DQVEz14LLpBdZAW9mYxIQBh9N3CTYQOfZSkWRMpulQ7pp1
Irsy6zn1xflCSEbcMFLkK0HXj0pg9bFoWXqnOxqbbqGJZ52LjqXi6xso07sXu4H1s+hlrwopvlXY
udHDeX9+Q1ll2krR92N9RcUKn+wSPfTqzaqhJPiuAC40QVvYS3xBjnACpQwaJDje6kYlZ+0gpwcb
a4HzgoRERNnYg/1Yzn36IA0TQf7tpE2rpfTT36YvTqQaxfw9YUJUgeVLd+VKhGivfG/Y6pyQwJCI
lrnsW+jNnXXhyed4b42TbZBZP7LzAZ5hIulp5UitqZBCRfkD8O3P1MPfSwr98xxPk0Iuw/keKkVP
AaId/75myKCgQdXQDMvq/zf5nVZz0CbVFfLPx7XeYBQJJDc1eRGo1jxNvRUrKLgYRcwqvwLVy1v1
VClKwvtRc0rjuuY9XrqjYbo3uufbBHvfSHPrsdojFhrL3GiazqyaHcP0csj/H/icyZNiDR2K6VdZ
DWQmlpq/rddPPMwcnPKvL+8uob465YT0veejqjDaoI7sGZ/klnY5lt4dnK2m8i2BjYWaOstq5VcC
xSGoQiUiswMMrudHFGp668iC1TeUV2RjPVf/IbmbDCYiRbRJma4pfPfD7cZmqvJyPzbogE1I2w/f
OLa9YBLBki6p0STZXrFDtdVU/jTUhupKtT/iKZyxm+4g7qU7YS8lGCXtOCCfI7LM3W3jR86usf0s
XCyx290bZGP1tn///lJHykCFzHIf+cYdhFnigvDAYCyyvXgyDWQ+8R5+tKV31amqFtAs9r3k4ipK
tzHcXZtVtO2Y0zujQiqwk+V2tSWf4jOmDjN55lC9Pjx5IGU/rkg6GxpxaAhTmSpcXYK3P2HnmTCi
SYGBgtIObdINaKlpcWhnAXfkLjJSKPzDb2ug0FxMiFYsniuOx89RFtFKeMbwqRo+4uwU5o2OP58R
f1svhAIxLeQdBpOYOaFZARRB5d8+DVTLwLLISNuNNJOfXjCTh7l0tLXWSwZ6xEYKbN6EkekV8chp
9cxVH/HAMmI35832NNth9gg2VoHAMrV5poD1SNfj6XsIngLt/wx+U+DGKNmSGkE4LwZH2F0JjN3q
WkR3TX+hYOWBhv+L9UNhTdA5hqaDqqoG0JS/hTY6oG7gDJzdwjoB7DzVASjhG7VmzaYvG+cXMn5L
49r3EWIeaU/P3CCxG0InLjRph8h3PqeBmzGJu6E04DPUML4Gd++xvlImRLTP+VpvbbOsJ/8jdS/w
1x3yfYajfn3cDhEIKKJTPEE4jMzAPeWiePsuj72BjDgdsPBAJhe+8aAxn0jgzCkJh2IGx+lCfl3c
PWwMXMQEkF/rd/x7LXRow4cTzU//SZdSQMQWKFG6sS0C67f4wiuyArcV7pj14fJZRURAVXBqQHin
ERB2iXncqdE9UcwcaVIdKcdSVwx3Jc3lmG7GhoF1baAHOQmaONebTB/YLvqxv+WhhfhHY8YfJz1s
QaQv18+Sk4/oiNeIz1mRqplSNrQyJ5y3TtNxXR0XoEAwAm5Zy0p+CExoj2L8LpBXYmBlFM3niN1D
oW7TJpGecF5x7CdxmC/VOPYMKjY4FdMjP4TIms4qtLs+LdrU1FuPwKnPiwzw5e7jDngEehXFXvoZ
WO+g8oHg0c1GTrzxSCy7VvokX/tsC2tXnpLUMK/m4YQxO+yfIXQO+2iGlNFtThsZmByETGgj7B2M
xQdLmvTUpcZp1EE0CGw8K2tBGmnmmrI/QmgbMkIp+0u897jAjUn+zzklabIUBxdAVCibS/x8ptUB
Z6QeZqjkzGhr4DVl8LCFGFyEWldBy6ICDVlQhySpCs90ENGgvB1a4a6ySBuJvumecNzRcaOYcZ4+
R3EetqCqCTT29qUhCspA/MuTdXTrv9iGm/TsAWY1TiURnhrEPawfKIF59L7L/giufcHNACow9uEo
Js7CyGYrwn3TOm9buJX2hJyZE3egZNhCloRCFULbg5bz7JAz4InYOp7dlmhiRdUIQzKbRK5O+SJL
84BaZwcFlbBHxyBX+rBFgnudmS+BKR3eyxGMDDP7VCDjtIumJ+FRqq7hhZ9nM/XJEJ38pDXdM7kg
NkOQFe4V2imwOPT1zEiaakcLDOg3rTOQp9Dbm/2acPJIsztxn4nMlT5f4NDYSi6cT0q+nXJflFer
PsYG468WuEorupRfM2S0EH2A54LJ3c5+NV06nxU1B6sWynT51YjzEZQ5euqi1xKsSFXxjWDMj40E
YIYoRjIOUPwDpoEk2/1vtO+y5ShKO7LJCfoyPL5W5KT62ukuXrKOlah6nX9u8nUvKXHMv7hGfTMN
rvByG8ep5QfaiWo/0QoWxvPBiN4MEUQ0tpqLdTXHwAkIP724IyIQBTBkqUtdDVqoglMwvVsr5HQo
AoH+NjeiliMS4TGSKrGaYhsOYlo3cr6SD+VIblLKrByVMn60nfZ7sOj4M2AbVxIWS3e0+ywIYkXz
NsaRM9pc5PrWsBN+kzBDX6Ruu5vwyFQc1WRx215zNyn9KSCzukiodvypAVMdZxBh67e/E3lEPoH/
nD4rFiBuROzYk3qYiREG+v0BDtsFilzPm2kC3bFowIPktlubYvxM4r531qMDBGCYlTkL570O+qb4
eEaVs/vNtlZjcfNiqP0HWKhxLt2Sf8R8I7hm1Ke2OrJitq6p1SzYGI9Lk85DE4is1P8WFNVDlkUv
TDYeoODWxKP2pgHqy8z9/P6grxluTVVzFYoXJJaxm4zodLWWuu6FubUfNnqhEsotIuCoS6pihtjB
RmI0A93yZsCi8C7gxHQ/j3SAcWl9qt00WBX7/8n5qWCoTtbmrlK4ysgVWbq9TCZFbPvuZbW8YmSk
2oBJ3yMBQlNDD2zUEBja14eZBOrDHzBp1TITrMSAanQsG0jW8hpvRJzlHwPzoof1ncX7Y6Ur9NmE
oS2LNZxrPWRBgwiA0X1w1TDY3IGuHGkA9LfUk5ypS66TlwRvM7sJdX1mo+VHsJvUN8TLnNbjuF/u
j6ob8g5VeRlVP7QUF2lToekiIN810qY/XyLDeHXr16eOxR/etA/IQ8qziWQbo2Vh55Sovfpe/aSY
BFJk6lzp0fp99/qgWPtIESUEZkFWzUJnUWJcqHn9P0V8v7zK+Y8aV3sV9h2WcndK0ao659ShcbMW
XS5AQs7aSrE6RjdjIkRcRglEQ3IkpJxZ45BRdq7HTv1qFdmtGPy8VxC6iySwAJKZ09z2yDdX28Oi
4uX1VMcCK+frM8koUQdHMzVwwXEmAOTpVZJ9D98rTkWMJD7ES+e7yk+5VRuVkW9VoOm2hiN5O/8W
eBbafMjPYWVYiUvPeEa7UG44UJacRCcBWBXRar51XanEzPhMy3Zf7UvnjOcIGTbReldaHtB9ICXA
5+TcVkxedwz9CF5XX/0mTBeeiLonvt3+68I8ub3p4IgL0r3gpZiG+3eQn4yWHaYE0TBH4BTlxPpq
MrF4NnxHc9joAHFG5Nz8zrwvG9AYwlGkL3PXl/jb+L7jWbF2n6xpucl9e3bVhny1Em9fb7t1GNcu
o/9tJirnoIF+x+wNe5jgdMo/7GMwTbLzJ7qA70k/kcZR3KGmSG8QuVM4bAhWcuJzCULM4E2fqV4d
tPq5Msr0vEpDKcRlopmjrexkqhdPyrEBroJmUX0rANa8urxFMd2nyJmf7hjZ7riGjgDIknXO/wK1
QObFVsI7FrXInyrIfcos4CxXfn3I6x7z7nJawm0hr0loOaXe9BmL+i2Tqv3xEV5m4qwdZ6seEYMd
CYGm0pf8YreHsh4l3Y23ko/Ohn0IcQbK35wHzsRYWU8CDChj4CL/C8kDGBVVoPjM2YZReFx1GQYb
joCTbMoystAjOEFi4Fd+ptsBBPullXgW+GB7cKUpAhMpBYzVz/jkHcVdYmsl0vnLQdUujxfW2pjf
HQMRXxFax5jRphOdjgn/EL2y83Glua3TP3aqAWLaYwXLg5b7zcE6O6vWvi25dw1MlCukIleUM4sx
ihv9JyDuLEAJ3q5PmHDUSXur7goOabj8J3Of/ldOxg67vfhhXxV5oYHc3KucEXfmcS4n/9QC3gkD
lwR0CFlp+UfjyT7AnQg9RLYWkLY+VVaSSlbMyzFKEeWrWtp6qe1XzUUBfZQRCMGdTjS3IoKpqyN6
crI+VPyA52pt5Qo49Ba+RheWfRVh6mc+CaCho723lmZ1nmH7a99+0YN3gcpopOUHMHTV0TQ/xq+v
HIPrwUFUe3iCidFyMB2+JEMBjE8JMwNIvXlvRggUcuGDpYdWJS4uYv6099Iy+Onz2kKTWKzwf0My
ThtCZaI/DEMx54IXNMMyoV42+D2uwcmx9S0Z/Mvm7WF2+igKDU5hdeayvd+3qUltN6fEl1kPheQV
CMZd2+yDA+pdlK3FUQdATszzWbWIxRb4W6SW2E2Owc3dEK92AV72UWAVmDTSD7uaiOgSP5CrNa/a
4VB/QPd+LNy8z87qIX83vjXxpF/Qi7tRGzMe2EZIWupQlk6vyG82tnFspwMHxDDS0QumJuWJjlJa
TODdg3p3ZNLIUJSh/+GyYZ0jGD9glntngzQhnLjs1ByIpAMCKRhEX+mecx/ZJ7WEubj2MsBrIfCG
xzxdg0FeJY+zPzqlOXyYZPLXfKleWcvOXbgW7Pso+PxRGU4HpkpO0QFt0KRqXE0tmyx2FDa93ExS
xIkU7Nr/rj93HbHhR/QxCkGXBhh98Oqb6/KJAAh1vytQSh62R8Oy4oGmV0Kxgkz4xu0yQOeYsRwd
ev99nSt9q1z5jmYhve1eY9hzQCiwIfrNEIdZbA5LbqtF7tCr7L5nJHRy2FyLOYgLYRvCJHNATGGb
i8FF1p9SoCkNqPz5PAqBpbM+neOhVnXWsUZu16DkEfemYo8eCuXD8QbENt9R2sZIlB4w7TrusqCc
/TxfQ9BwIDQHEf3kYG8ylpUfBShdHxvNSa1XWJ0p61cQpw+jQvw67MgmgMHLyzNL2EYLnkfoHeNL
SYlZMXVUeWu1tFaliVTjUGm/YxRyWYrjuXGK/k8qGJBT0EKuyERb1hEZp5m8izL8qXUHdXYhjiRK
5iKMSb64IKoVAPOFTUJO04j9dQLAXncx8sOTLr1uROcmayR54HGSnaJ3MK0pYR4F+N9U9EOWDi68
zTuITTFWnXwUDIaCmhXzpq/EdlsqYrQbeMaVof5Lp0YMg6QJqUDfx7/xc0BVO5K8hv0FbW7IYu9S
YFfXEbcAhKvSXkVEN6rKc3Znv3t7b1i3i/o4+Cm3lUaYjXH0dPAnUli18o/vpU7OUtezVf0AM8Ld
+5Lwsqgu0VIN8xtLg9VrBMz9gwMpM3yDk4ZrzlkwcyZRUtLiq4CQbJt5Xz1E6/mxqyVJvMGUb/yZ
vtT89EOsA9ycMMpqMJayjUVFyTah8zhxnNdvUX9uB2G7vFk69rf6dp/WcbfGk9RWbAnI+bT7/q/d
CTBE09+fD/qznUmmAW+0UdtOQY2Q7LXc2wrRxykflwFGxj+OmA+MsTgpr9bcLeja2qP2b6/w6foF
9pzYLh2Xc6LedxbpGkqN2OmUiEDDxaJUw6DxTKH+zSJYW5P3D8aB8ZJL2hOdn77H7vvDZb62Kb4s
G6+a5BZMG3H3rdHvQ/33E1FdnetTxkF1V323gSA9hhdTbsHHz8KLww6k1vVV+iG+JYPCaCPU40rT
LuD8rX9KhHBsSWjMiyuQP6IldJhWLvJdTz9/lLdnseN2uW9MnpNJHzgzUMOaY31ok6ccSt/hDxQV
YA5vPwe0xtHkRwzUAfFHsevtgW6oe/7Vp7k+tJ1OiET5IY2APdNI7eqQahgPytQQKHhWBFzI2sEf
JRyvI4mqg0wctqfyXDP3SHU6P/iTl9igSfvLpUm8KNfW0jWZtC3noB8TG4M7Epdlf4ujsQUSRY80
HuHxKLb3eTj7pYtrQT9t6qby/rEhSlKGc0gIRSnv/4Y/lpK455IWtbLXumobM26FjzMgPCExWiYS
+Yzra0o/RFtgPRun/ovYkZono9Wrx2DeRTaA7bbwpTpCHHuJhA74wYkfPqAyWrfOtwdjhQWxQNlg
FFk7/4LLgV1nS+uEgfwGeGMT4k+lJqA964GuwKgcF1EtamkJ4A1AcJyNSMVn73uNLwEdRYEB+EHo
N8WCnuuOAMmd+XLrOcdtT56BHo8m8HHlkF0VBosEcmQ/nCb6hIbJwcn4TMJebTXPD7MVjDtwU0Rf
r3iTSUj/O8ctDd+JCXqqPLnxgmsFTGmpcepRA1bIuv0N69ha5i13Itqj6pJKYVIotLiEI/C9C924
SrbUqWZvKDubBdNSNJvSFEDAk6FL8dU6Je0u8FiBvwO9MYej5c2I4fb1KIxwzCYrTft/SumWqfAC
yvEges7kbH4Ci9XedaCYVSWV2BWx9fbm3efmkbn+4NYuBw2UQLJp6IkmumWFZzm+F4GbMdVVXxgR
iKql+aJv+2VqUyqN1RCRnnL/yLsFOrz3hc7956w7bgDJF/UTKH02tvdgxMQ8kvWqM53u+m/Jhg8G
XoCVKnJJZzCnFOMpVaag/qecVb+zikci3KtDV6hwjAW07ZvAxvojplwWiCCsdZiAW7i++6PZhD0z
0+axdCvLcz2wE1Nl1PBPOXDvQq2qgs7ERZJ0Mtwebd11We2xM/+4KrbcZ1XVOw5VUA+uHmn4fmdS
l1LDPXENewS8GrL3xNvw6owyaMk4ZNsncqKhiEk3gdQXlsqaiBS07slvvQ5W1IkrFgZrw5D+EhLz
eFmh3E1V0D5tpG1xhC86SyDRKhnW5yjIeG+9Zo8mIqPIyyKHyGjj3E29irLJGkohKhsvrLezWiwi
JgHWUkweqG7FvyTDowA4tyqAog0QlCTsack2MrVQFticeEUX9sQpIY+9ef3/6KMFI+xRSHKmahy4
o+TD2kUML8Pyms0C4+C3HipGKKVkgHYleqajfuf7DhEPY1Zz4ndoO5hPg2kIyDx2wrABZvz6xtyG
VDn1MZ8D+WK3gUV77ZIgL/JCuLf0/6dYkVRlXdHY12986mgXY6Fc8WhzXzvMmlOxoXudFAlI+w7M
kS9zQYMNMZlmfwupTruUUi2B28m5Wz+F2q1SvcrLYL9c5WWBhoPvCh3Hc6QO0xzrfG4fAf0jshI1
hRO7hZv+CkEFaUNsBETcYD5/iESku92S1FulX7FS9BnIh16ICxgSMsMW4F558r0jQOBvUbogqwbg
AYu0Kjp97Rk8T9Yu+qgfY7v3mi5xaSBpvH0zEcrpheZvj2s9rUECGFvIJo1v67bifgmwy+qFY9eq
J1xB00+OdjmZzByqWnsX7MeVhrz8kKt587QTFscrKxtEcbIdGuazfER+sQMLU8QNFheORi9E8qcZ
wbIaVTpKKlJBCaZXMvF4Ovp2htkNNhM5rVax0/yEbLustC6qKy7m5/1Q+Eknj9dBx9bCDuYQaEMO
aLj1ovJI+tRi0dGceaaxwiax+x87iiwhPpU1HfMdcu0sUe7LPMJF6GvOSHGxePsjRkFqGc7WpBpy
fM6NEVEdpngxAXz4jcwVchMfes0v5SMQlXvsQBRhzv9UsMXaoPrF7P0n7ostaNXkJD9hsXk/I5h9
0JWxUJwABp2x6s9yzhXX0f1BkIvmopOenjeRAEtFfuhL8E+v9PBocU3Bzpg9aSefmcggWbCfWOt0
JRZdPZvmR0U6GWpt31zyMk2CZX6yhYNj8kbM+EzSJTk+y3H1DlPIrDnV+OlT/vX6WIHqNurWOjwm
MyGzbSvnCb5nCmu9d4pG8cMzjLzrOTYWXQ0TvD3uCTizX1KP07b2UJ4WviZ6Cip53D39y1MjOSHy
pR0cU/kLqlf97BG1XucF6r4+DBmo+yP9q/9nGqX4hivhwosZVx7ybwaLB+o4FTrHSQYtwHH0c4r2
O22jb3gYZ5hku3H+KzglLHJxoqUCNoaP+i0zEGH6YzMxucsXzPAtVbQ9Gr5YVzBPVKP4X8+wKvFT
2cchuYE6zoBwtfTyn/EVpf14tMjZGdZCJBXEsKPBH2OdVOIF60Qk4U0GEJNMxkyllcgPs6TGKM3c
7N2LeRjEnRdn7RPqJ70rIni4639QKavTtRkgxGvGb+6L4BDhTzoUVl70irKiRoXvNiPSApNz/mF6
ce+uXr9wzI4T2wUWk15CYqXwGU8/NPmpYSpXKGwi2NTw2urL5Cfj0E5223lw99Ke1ZyGNrGQYTtY
fBLYugjuy6AySg9VpAo46sTaoxLEOIlR1U5GIMYXi7bqF1JrmfeW+C9vSJSgnuqmAqZ3aghjMDum
8cxJwmxTcfgyl8/vLNdchB1+CWjF6Imc2/Y1FfH+kdFdTiZCylrDWws/jVlUJ/FzAEvAFLQGUdQ6
72BKbHQfW4QGHyQePS8r4ZAQIzn3ohQcaA7lsrOQv5yYGL4DXJziX0KsGXH5DIE3igvXyVpo7D+B
NMKjwUVOjVNsW+nKK2cMrN+RxKQkCrha3eUb7UUsrq7U2OJc/yT8jgsTsbmuxgWSpnFCZCFldp6g
u5MlSBOADa8KBHA6y7pt4okFOcWTJtgaI1DakmXMU2w7/ctZDT1aN+/cTdGetMX6trxOjYi53uMZ
OQ7eqh5Z5AN0ItCyg0ek8zeknpYXlW4sELKnflxO84nIfEwwqPQ5F1TzldLGT89t3xAUL6px9Mjt
W6Kqb6LUV2OSnWVc1u7Xx2KCNtWdjaPEFD/cVlZpoZGDZZdZEf/GsproRqT7jdBWVnhsBjzXRedn
7li9Q8EUz1xfSxuWv2R0Bx6cleONq0++slUrqlZBPlQro8rNDjr8Xnbq+SH4Si2CCZM+sqzYK+W9
Ltp0qsdwMwS88Ve90lM+jf3SO/B74+qr1ksYP6QlJZB3ddVF30N6Lx6n4r4d3JEYynWwJ+rX/9CO
ZzWT6MW2ab2qjpMDttKxSHY8yzUWt7mxrNkR94g4+1LASrRTl5M3VR4q3h/Aw4+ZvHl/K6AtRfvz
A4aw3TZsbDPkAEd9ZS7PajBsTzYoK6QaLiENo2DFJvbZYGXuTPv4KAPNd+OO6VZZc59cS0UhhBgE
0DefDxAphEdz60mudHVDaXLAuHB7D0iaXX0IFdkSnKJbkLYtqI7gBUfdJd4Pl48rtY9WvSxn6IbG
2cnuf9lVP3YA4OajKNpD+aXfrPEQjCWpYGxbl/yhypyh4iHwBnMZI5COLysOm1AOQUUj9JEY14zf
Oxb89ExR81w1wCjKAMuKCpkHAYA+qA/rHv5RgUOL8f+SWETncdSgmAvCB80/zSdMRq/D1rQX3Mol
gIm4aXrFUBiMpFDiij8nMOJW7G23BDLqiWuv6MZTiDaaw8U6ktLafYihQpr0ZfavznnqyYmuqxJ1
z+UUNI7bOtvId8zpVJVtm5k1vynMiyIvfdFGVN/LRFPdv8PpmWA3U4q4czP7w+8jUkOCtJm4kdU1
r9hBOX9yIW5rl+GF413NKrm32TcxNEPTxnMpcRzZ/p/c1m+bgJEKSICepeOvG/ExgOI8BoLtAvYn
K1XTrGsHI5F+W71rlw1xve895V6sy6fYVQiu7FvcxQvvdVd5yti53KdOyj3KMxHYUp2JvOZ5zkjZ
cvnJp8wgURFjN0osI9Eul/hF56Xt3p8fryZnfLV6uW/APTVLTAAOxp4TFGDx/iofZrcRgBXsKhkT
hdfDE1C20rDUsIbT5msuqrX+iVp8e2Du+mBgO9WMe3zJeErX7BYQsesqqTkz/TnEfhuZsHg2W3Rc
tGMdTurJL+rabNHQNWv895BqKcu3OTWeqbTJWc9Vco9yFa1EgiQVfh66TnJDxa7if+9UmmUY1jja
c2vdTLSUku/SQk/Flt3IT/PoH9Txg+CIAxb57k9EjulH/LMWtNWaBK2K8PijZnIo81bGVYDo9vDt
zoeHFEo3j8n1rCuOYQr9XjpVnduY4zYBGhrF/vSQJUaqRpG32mkwdbIOv11+Z2Yn+T8WhJmHcx0Q
fP2cnDD/S+AZleXthA8/+iqh8ID/GlpDrxQITxqIL3L5Vykp8dDIAxr3VIeGXxrJ+bmtVp9JA/3O
c6uwwa7uTg8L2/btPRwZN657JaTU3pyIRltmeLk9MIB+vTFl4/BYdEeX0avY4kpS7+2HUEGsHUY0
fBVs6mkV+sZj5C2OJ5argbnzN+Tcfrif6UcdgibKyyn0i/f9y4uudNbTHy/1XO0dP+fO0cmsPTw5
tlnHX+mOvRhHd46ChuRJLp/9GD1NtES8+Ya6S+BN4y+ew6dUoPpbiCh0eHEP3fR8Xfl956Ti2qSV
eRZA0IAD6BqP1nSPp3alOnQcajVpO86z0J+FtxrJC9D5tW9ZNZP0mGeZEIr0dAi1TEWOWiL47BxG
yhFcWukC65POt2aF8gsjUF1gjFE9NolnJb/RlNrtPLzrcVmpdXXke6rhVeNdA73+QVAbMrpVzol7
94umieJfE2fMNDqOlofZFxWdNvMNJmvFMXyLrxs/zwXpMZTHIJLZtEItMxOvvGWSTSMI5vf9adgF
noZnzdsw9dwKuRO86Lype39ZetsXxvzjoywVZxp9u5CvxYZtyns4Hscf2Eit/1LILgKmEdrTlDW4
mJrsEXmOwi5g74pGVYonGjNmY0Rk/hBrPLzlCo4vPw1ScnlLyMRhQrYbQ65ptO1hC4JgnOdQ5Bwk
mBBfu4whjWbzAPkAkgnxRu/tjJdNUTAixVKo3VjUlxvxS2VPhqi4YbBmbyeGThd2vDf/novmjBJI
UjUvmfHt3piIH6wQxtgim8l0QWBLyint3KmRJ0swu6uDuCj18O8w2MXqIu+YWRkHWX3SmFulbYwM
p2Ps6eIO+Bb53AK7EFjiFtH0bFI3bLnkgcUiuHC8l+lL/ilsGEQVQGIJGF7SC9Djoh6pnwB3CbXd
YUUqmtKnpThjmInO+iaAbRAXyk7MHNoVHQ+aYjk7JtD8q3+qMioFM+aZD8swvAyzVxBvZbG1EbLJ
uwdu9CnNNBcofDeb7c0iHlQ7BhV8JqHjA4+L93e7RgnVDw1MbZrHLNmdZGRxsWnGjrwfhn5kkphj
bBAmHb+6vB00DKPpE2fpy+k9BVKU9xSpaLJ0QuSqubHETelamF/chIDSg5jlO/px958tlo382sfH
5jdMrVo9XkWrAJqFJUlQLi5MAx9rNsaHbshCZNHtP3kSqs0Td3LjSVa6n64HbyjiKZwJ/ayPqdaz
fgAhvoS526DB7W1PTTDv3LIkmPwTd6CibuvhdpgK0jQtIPb0gmsJ4fazbz+s7Yfgzwhbp/Ftqrlb
T04XMY9IoAEq4OK4H59qprHVWzDCopbpjRyAESNwbpAUqHBjMj19YzowriMb7Qrb+1Xi3tySSrbh
eXPoIeX83JXS4eNXiSyiOlMHV3+AIaWOjkoCO+c4ERj9ZFldoNuJTxH+xOhCWd9i51sqwQ5T52TR
dgIQtMjdKkBdyEaaoWCzhO4PwErXawi0BkaHCeQQUw/k9+5sIATTyi+2x60S25o7DZmdL1KtbsSf
CYS5TKwHlNCIrHF2czIZcHrT87Zxd5C/B0XUCd7J5Ail8mQs5mEAOrrM38kSyNIolWIX7cyjh1ij
QY7dYqscNkDQSJtp6VdctscymDQZVNaEMSNqeZn92P/G6ysQcgsCrTC5T1fIHtXxEyQax6o6hQIJ
O09yq9+cDlR/cDiR1XgUYmg4Dhut+8p8hjDOFu+zUN2H4wZWj6/bT6ScREuip/h9E/hFXLoF8m66
gUv0wLWnWKhK/vCZ67yFvXAWVw0tOW/ToVqVF+e0Acs6kLdUXqWysaB+B6Ipk7wh4297nFm74Xo0
9R3Ly4MZVatsvYNcLd273We6UGmD5y1AndNCY63MYvawMbVSAXwCBv0OCKfmQQnRgoVaw+FtGmph
U92Ti+wRcqi4DtO09lO4YBrqO+PnANiLJnOot9R6rw2vQX+a7iJPLNvHFpHln5LAXbaFrN4+eksk
QYMHdy/2fXWlqtJQToFVRZwVTdqKawzl8AOhtQBoGIl7+J7+oCHiDOb/t+DoSwMN/KkIh14fhuf0
5YbCzL+TPLvr49RlIoTACZ9/cxyFzg1Atry4/YlpBjOeYqx7r7ULzwDwH8qk20ZoBkSC8oHdmetg
S5sk1o3w+Xek668TKyrvA8XVazFma8fhUr/T5FScpLeNHcs+pI7floh4tCfALiYFM1Mfqs1gC8fm
CbdAfVSXQmHuRN1SX49fxlyPxzvNzxbemqxHDvzNJtomdtTsEGtlwICrojN80QFUhw7f+It+pIvo
oMYf6qOV4rumjOr6/ju5uRhGcRSJh6lI2gPKoWRv4ymBrM1nW2N2OM2nv+w2XYgUFJpi70ytwXi3
BfnRaS6iEMnKmZqdWEt3K+62TjbBhqJRKOW98eeVyUSxlQyjMuLsfAfUZetiOdXCQ+z/ezGZKkhb
IEtpbf81rYQlwo0TFbikL0b0R0cn3dNqkXfZwSZTLEw8dMDKrAmxDy1fdha6tilMUKA2GGc1yyHB
I8fftdqaE5i4to4J0XBrmi7f7LBunZ6uGqSAKFkiqUrPVQIsBNiRea7mEXKjgDKPLauQ+za3hA6a
7MH5HHshRW1hiSbgQ39PPM7P8Ed8SqYIFWeLmPEnJRzXfoAMYHT9UiSnGrpQi4IlpwC7o3T3m06M
Q82Hno4FqLYLQqI0ou1u2ko5iMdhTY23rPKVIDxHt9H8o4N0EW6+FdgEOLIOQiJrMv/WgRx0cEO8
rReIb1N74RA7D+r0RVIJiIEe5GMa7mJ25Bi/MmRXzG/KW76M97SVr87qIAweuld/xqgJc5aEJIfo
4fgtBWkI0TUeJmvg3Nkxgt3+XE/GZTLhDMwxn1j25nlVVAsi4ne4PC+eSQYQ7sB/gJERzgRsaSZv
EppxpXOaj1D9oVxE0YJLvIzPYvn5Z1ppui2iUArrJkVrqYI4/dQuvkujz4pbUnugfyeAITXqJM5q
/rjFrEeVcVoEG+RSBXSjMTgtk6MffYpUY15Hub1NUhXd00h2BC+kbfPXgwrHgbK5FhVm5I10Nyvp
oGuMTKb7hAjTUnkdeP4xclM968bE3jkZfbiNBbxm0i//J3XusjZOHuELsKNmnTkFxbp4Aq+qEZLt
EQa1fcllTC7naCwfcW/DXf7Ik1aJIVOEoh1EPHVFrdBXRcX3Dj4XCKhnCNjo3x9qin2Z/eliHFxB
hiSCMXoZc2br9R/pAVJ+SVo8k6CqWnZ8zDuDFcSlZwtkGLKAdnpeOeXu5OZWwVDQb78rgQvqv+Ia
zECG/1DK68hZrHhgWEH+1dT3XDul9SbnKC9YVjGXxhjcdmsEg1uUACnzRXsEW3F0Nv1jAHnwPi+j
Xp+Lyfy60N+cr+2WC8w+qObLm2kJfCWMx/Vd/cngAxRKW2WusINWu2wqdc8O9YxnIsDHecCQo5KD
R4mpT+iMo8MStFZ1nYAf+2MZ1mYtWxqr0Z2MEO93AnRyGjaUxqwiqcQypWBLvBdGuYle2bZyRb3P
NPuS6G+qVLSNp/ZCoguvzwcVNJdtQQUZJ2hmwEI6FP1b1LKLtP9qAGBWjSYylotxOD8PSupjV5BH
vap8NSGCBSIDfifjphK3RbYjKJc5uom2VzHy8h20guHAjsc5WzRRx3sQhvmbV3NRbBpUlmVoQ6Pi
CxIKN8hdFkh7NXr81CpP612dgKe6gVOrJ8DE6YuKlKiOy7b2ZleS+jrB5AeCaaIWM2vw09pNNLiZ
1n0BeZimyAwhXu5S5SaG2eOvFMnwuiTexyhD87hDUmkm3ehUwxrlC3wXDeIfqIYMjCBM2WrHJSxH
zWpkE/5pi8qQTziCE6Y4UyZydNXoshM5zJ+IZMrA+t8CdIBfRxIrSWoj9MpkhPtOaS8lk6OnrD3p
JZo492xG5qNdSfDGDMGgrqKBdlkeDMl0v1QfRucJCyHWyOF3lJELS8Umf98l27UeUBuaxErpqys5
oxSjaBpzvjQBfUCtbRbKOoiHyZYUPsBHAftK5E//GwvaBC9bDNavSXxTRA6BurYXe+8d4Cu9OuuT
zh9UT6Q9C9UF7eFRGUJqXjafBm1gVKMmPGkgfAtV7Tb9KZKJVogSuU1oNTXbx1tb2TOAjyoRjukO
X6Bnb8ZdcqLf2PLffKSuB+Vl0azQidH+NeouCfiMbsUa+n8mtzf7z03q4Yj/wkTwZy3uit8GjlyV
UjBdIjiuh+8FxlBFpxOBIVeKbUJ3YMeRwWi6wd25JqLHz8LpTNeu0CdWUiJAFtIn+/2/27yG1Zx6
wDfEHTMEUNiiTGnAJAwCNqgleEY5ScezOhE1qlcSipfkrreWDjueTsGtlJIL+4oXQLvghtbRNrtl
vsldaG4T8Rs42TiUSDzbvN6vWCx3X0NeKLv1DNJx6spafkKAUYHDktlkFLPyBfQJDsioCw0nVlsE
G67zpX7Z+IddUz5Jz+dR3XZUVkzYud+qGYu1kKKF/xTvpWzpHtJFQslFJUW/YN11wdTCYy2rUwQK
ud88bwZmzXY+1JKkCK8iICBtw39m+NpEcS0crrJLSa9PYzmNQ+LT0HUp99Sj6ng5ZXE1k4MJ6MQ7
UbmK//BOGovQR4p9myoQuS1kDcmcW+gV8d0pdfzMH2fBlUeX7K72KklWIj3obTicSUJf4W6utiti
LE1F2zGR5T5afp+1S/IuPIHY+Eihl45c4mo85vjshmObz1toVbWhuZhuHQiiJD8zKSD4riIgceIz
RHck3a/Y906Coa/b5cCvJ32JQqYncWbOwn5lGThpFSi+WwL5sbWpSrDSduhM0hKwPQpNECUcqjpd
x20r+zRiNrV6cKDWLSHCkjzfQGq888fB4iVJjdWgFxodat+AQx0O3N/VXJB29crJOSEL7QBQ9bIg
LC9Dux/YGn5a2RZQq+yFglCTlqIJ9KaMMLX5+eNpOZ7+jdbVbnEZ2C8pzXa2wVsr1KiVPIZv/sbe
eiAgGSjH36YC2KbKvnT0HfvdrKJbu9RRtKotO7yBhYs9yveLw7uKu9uVk6PV1rD58UgMGDVWPa6y
SP+xrhkvJqkEir2XICkAufbhNGWq1oa85djtuQNL90boTcKcHUnqVrr2dewKLSIupetbmqu2f9Qv
0YgfgYkRiA9+7N0INoVLsrfIucDsaozFo25+4q90AFcRUMog5OU/C8VXlnhhoEl2u2cisSvmugHH
Ix5KYugdP2qgIc69CDhpRITeO2XyzZHKcrznNEdfnjzv/vRb4BkU4SZK9mdkS7LUpKKJNnydP3d0
HUL6wL8kzZ60cvTtpLAHWDIZjwkSC8F6f+62VERDG04Y6t67Z2b0v9epIxj6xp6iHRHcr5/a30na
8P9DXFGKOi+LFWd/LfBauwT3LvYvMweBq9gA8PzF64NmjFn8Z6zXYoubqv3tXN1cputuQTnlF2/5
ynCnKdjb3Oo1Mz7FRGKO3hdrJdf1ktPuKebmkzVdPRlDuz4WNMEr4Rv4eIhDRgx1GqTU4yLKpiqk
ujvrFTVmE9sUSiOefwBf9WMlHRH+qF5615PwBfpiMiGSNIarKR1xk1dJGbyb4er890XqenBJytuI
r+HAWCO5KLQ6UIGoRtn8RZN/Id/1+6VPdryQXoTTGjqjAiSt+PhMUU7bebi82ZysmKxmLsR4uRNC
ouWRMw9THpnRi03HbavNYp6fXiB877wHSyFqjOgr5EFLsFm3ZNeTT6bWKhLwphzYzRZWPABSQJeE
wR85+uR6saFeKW8VV/MIH6m4Gpjgj8PvzJs0tEDO0P7IFjbqzysYb5SWjVP1lUBU/Bb65oIGwYDz
xw+x+3MusgzE5H88pb8etAPLQuEDIFCw+MPTLWmTvtXIgNszGMEqalYu9jTW36sxKqd8wRw6Dqin
8vqVs+cLp5rWW0yKc++D9czMXY276dwcuQql6m19AJcTPv5erVhoda8f2PIIs/fUuQRV/rHxFiYb
Kabfnn//Ap8AsmxUV65DpWl5uSJQVe2TuKyIrwNbro55YlsxOhZVmtYv5cimQo54bEUWtNoHY6/N
HfXaLsuqbpDjogbCvJeIwhTlzUis+j3Ltf8S/s6gOMOXy1fFnZiMkTnQPHqdy7KZhUzZySpwlXF5
mAgKBXrZgjy/O40RUWvgWw5MEo9V/u5mbMR4t4crJzd7ikbOeCCCCAPaAt3xCHGVmlnRxSKdy+ct
NehdqSMq0W5yvd3zgMckRnQa2viKrzkMeZeRZnKpZFJeacJMozfYZ21YmMIiIgWEYkZ3EJdZO15P
EUdME5E8KT2lQ2+8NFl3Si/mnbjpF9UZEJ1e53ANRnyLNDtEyqXTfhbUowLJJAhG4gZlYKzRPY1m
kiSmUR5xtb7LdXzmRQEwYFEClQ3PR0JnHzrcXasSzKIAbugBHOCqJT3ZhTNahig+2LsnBmMIcY58
69Bsk5Ul2rzOJuQetA7aP2ikN0jKYjxNjZnQcNDAXcX+FQhdE+8OJJxikukgGs9LURwlggUaC73p
e1FcptlPEsKsVnqptyfDx+pRgkmS586MgEDWEdaXwtj2infPx2TK07W9fwyN3H2odwtQ82c7d0LN
gNEfvIjlKLWRsxconacAgS03r4ocuhSn1E4g72IPX6oYZx03scgnEAWnnbEdWPB30eKuGWFF+IMT
dYDMsc9nR7CugPO0XMhd6giQXc2xEaHRuX48MXFVWCxVsC3KJ34uG7lsxw7LgLpnQ3X2ipdcWxpl
3VRBMlZfBBHjDlSFOXbu95WTuKRTC7NWnhrjwDNRcI07YGuYezNinTccB2EwI+EVcXmZSkBAeljv
BtroXlddv08EYlL8OWD79SfwMTT+KQoQ2rGRRhOeR2C15PiAwE+t5we1FmAgxeTgEiwKfGxbTIgE
ik+pgwaOp4kvPJNKNhcUg34rsWyuk1lrKgBjMs5nzw6knrB8tgJxbh+a4vQDH4m00eKQjrHVKwUx
6SirChvhmSBaElXSrVV+aiIs1fregX1Lz6yFRrtAC/aM4J9uYIZuE3R3BPA39dGsH7BXYLQrcqvr
K/1QeYNR4aUEjVT7wCxNZg/JmbOsdvkwgxatuoFHBRop7oLtcsh4qBPVj3BnGaf7rfNnIuzwDxUr
QGsRq53hwSw+al53r7vH5hCdVEScg3xB4W0cmnrHvTANqGX0oNZdwM/nsJfdgTtop0xaWeih5moP
4/nKaa+DTkY1nMxDIe378bvxbId/vP1lT/np+2qyNNXl8rnKlFyo4nEo/PLtZcxYzvhOXbS9qyLV
qpf0Dh4YnDIO98X5Wky8aD/9qnfpm+FFDsWIfr4uQFGjBjOUtXKa8S0L4gq/Alj7nBsY+/hbt+k4
+gF9RGskXUtYtIOAgcHdvxngDgbt9am2zYe7P1PnBU1uchyh9khp+CFcY9Ntz9VpgD+infDyyAgR
YyRv8ZDcGQi9Q6tkleT6RV5giEDnhBEtvFFIFNopT085rqexfJt0ytuxYnpg+7QhzVSp9blBPbvb
oWXdDGdhIwm+QlgPRWLzxbws3NsjDGgcRGK2Arpiv2RuyytYLQA77qUaGIuwxFDn6Ofzb1RGaAqq
RyvFTreSDXADkx2E0DJGJTTtX4rSjiAOVy2+BRbZNT+99zL1/nytHKvJr66dnaiy9+7hNDAh8QAM
uuf0QIbX0DnZggAyXk8kW60NXO+ZoAy6P65oCzWQcRVxtjIU8EKTStUD0ox3T8mXyIcifcVZvKAK
ZKGTJQX0hbL0YuF7wwEq8QbUtgzZpXKaVRqY/X6DWM7IGNcTIRsS8DCw8i1Ji7UzxS1bJAhJ/7lo
23l3hjZ8sGyTQyApTMSlXqbKF7HJNXGF4aCa3CxOeFCEeW/knmQ5DOh0YBLgXyapM2OQ/6TuMEtP
5rBh0yH36U7DWlQcx3zilM2rB7OmOeUxEPcuB0XmEyiPFXv2pUOr/45ubvr0i6HYAeL2nUnBWqEX
gP5QcbM8sAu+mUb4KqE04DVpoqiCf4DKJkIP/AvPEAt8lZLjRDEEfih5ZA1XfOrAuqaHDi+iA5lJ
zshj4ytz7cPsyv3grmL4x4VEMWkIlTjC2oYsyZIkkwrQlJwouANSCxGQyiBgY1fqqAqVKyyTPvN/
uoZF/XGaYRqs5xdW+44aiWV2+0Getv7VhaIcx/m7Axv+p/2jUG0YEA/Fqxj2x0OBmtIQd8/A/Y1A
nG2n2YpUu0DMdVQOi85EdZ/ePDbxjVXVSyWIrSq9gqpHr1x23EVUOyUX45LmjwgrJLZmx3FsLm3/
ucRQ5Yn2KW4ujLEuwSOTtJMUtcbcCWhgqO197Xlc5GGCnvsOFtGwELhsXpU0IP1sNs7vSNVJWj+p
yVVONX4EmNS7e5HP6PoIy01RL1ma44OAyFHtSfTFopUkd+ZtgKIWt+BB6Os8aVKoEti+DYfC+mAk
I3byKBfCdxB2qbXeiO7+IhPenJCXWjcUx0XepqY68xXCbUKo+yAkgurrRmbRF54w2Xlfq7CTVi1x
oPSGpB16slxEgz9trZlNQIJKP82oUgRglnqZ4tAHVjV+V2Y1mskbJekp3WPk/TVYWbvn74lJIhp+
E/fTNtKVb+jKSgOoNVZiAZjkS46ik60oN7CbHzAtHJ2UdLAtWS8RPOF5Kq7GWvCGglTqOZ/GKJkA
0R3u3kEgyvvbbx0jCFmHhKoMceBxuJzswb6kPJuLbAauR7GJF2I5KhXpz2R5m+S/CeqmpsIxWKwP
aaSF0q5p4ZYM8xDMDbOi2PFe7kiMtncWG8jmloMIlz6j/z/Pd9NrjT3z5Z1YjweJRcL2qkVm9bP8
Mc3Qn5EebqHChoZ0/Sb8eRFUSchdP2Hk78TBpFvdPdSXiRkxFPcCtGg2ifKtHzj3DBjrs3BA9Vzk
2TW6t7uN24lLB2pYCxTE8AjsXgMrirMao8Aq8TK+tw4ed03c7zaZZW3J401DPnx/9v0b8F/YT5r0
E/iWnoJ2K1LYjcaaF+7AXLIhQPKEwW+igpphbnDglbtogChjAHgET8cjZnW1pJ0qIa8FygxF36z8
lyTZynFs2542bB07gL7VfF77k3HJc+mxTjTsdt9f2Q8czpWyb7S0lTxveAeTGq4HH0fiyzccNCwV
kWHTfovrsZIkc2Do6DBN3M/lSBgJ/gRMOHZKZZgG+lOITcOWiQvKlky8c86FybNhDUk3+67ajIbN
UtUvJyo07b+oEa4QlwpkBiUUJcXIssb13szHnEBdmk15j8p84ioC/5OAKQMMJ6MRAZkQwoMBCyUk
PGzkCgzfGGsfM51071Onl14kg803QUbrPnBBfFwNPpG0zkVfaroLvwzcmA1cegH0MDseNen6HQU/
BtVtBPs/vFlSVJ6bd98YjM45A2vKkuB8Uly/6VE5sb6hC3lUAupT1PpZi+gVXQ+bRHTFqcXnF4CB
1J8ISHQWuxTd7NK+IPni7eSbTbkUmq7v86kZK9/PI90QGORetRewsmEZBkW+Ofxm6CGVLA+XwS35
n3DlePFc6nBEMEFaY15XepigUeHx8Qa5iNl8KVT5/ztEpzFpPW7v1zG2LBQWeTm2Xs9lveOfkx5Z
aKGpMTosqW6D/B1mogaIAp9WqE9FkG9IBC3KiImnHub+0Gjd20QpOqZ07ppIIs94tOrfnmaOh8ZJ
u6+Q3jgYjb20qssDMmFMXafqlep+OGN7utcl5QPUxB8iJdivI9wI+P2qg9VbQC2buS2AvmPTuqaG
dlncU7KfSgr7ArVQEpSYHiu1G5JJE+DDBe/w7/HHttF+kNszXOpOpQZK0+WRUzytIgAHb5AZBmYA
lislD3miwkHAfCgbEbePFyLLp0Qh7H735SgtvNJh0Lo0ibK20rc03efRhvt42g5ZgdvYJr+7R9il
uauDggQrJumQ09gGbJPUsR3kLYyBGjSS3cbIO1iqG/xSp0FiQNhpHhYB2St14PkV6SLL4dh3B6wW
zoiKLE9VzXhmLiZ/MTwPHLD8vbFcNHRnDi8t+c7IqV9+2Zzs5DIQHZXMmBXDSTF292Vw4gwaSz6Q
5aKUshOJyWmxj/YleB36+EfL5fTBeaP0SCx0wx6jbWu8nmyei542PpLgVpPANzPRMf3n9RLMxNF4
48JZwxilE5LNfC4gZNbtgAaxVAasGaH3rZ51HXhWWlqBsUkSibW9mmvyl16VqrIffPQT0/kFzDa2
amXXFDoCjJ/kJt5JhQUIJJZdyqprKhzsMVlRuUbXAl4l9fZyfrJq2ds3FK973aEW5UlMCR+ttJV0
gfPymFglklpnIrs9jFs9OEv8UGcPKybTKWddkSYCFbMe3rNnEsNDxUwYqDtupQJge9TNpVDU2gd2
6jbmtOeX9p0egyztW2pmVT1CpzI1VvmCJCRzep69Kra8X6iQpZVoifWXGG93g2h1YMj8L1APIJro
zztkHSv6iLn0MEhYTZL++CGAPBocBzdVgafhzlTsoAG9YtFXj5glJ9kKQhneZq+eftBS4Czs6TXN
waAHYOxaXWl0/NZ23OObKMyzdQxIu5tCLoM8B3Lo1d1ryNLpjd4qDsbtFdYBeiOqXFJJj+Xahoak
PRBjwb3CQZl21UY3e+K4m+QSlnnVheHStJ0X5DIDmQrfnWuIuSFzCm2A2WazOQ0O2Vher8RE8jll
V6rbDlB60GMyvDE4RZwanfNu0WArIXXVo4hWQs3rSmZG0WbsW+mHpMe6K5/9veHLFjEnkhXJ08mn
evQmVD7MeA39QNNAClM/QAgdolfLrIR9FpeND9A4FNwgu8LbEQhoUnT5JAmW+GWds6ivDk67wxu8
08R2t/eXc26C59C195ES5QD15r75kmBMuq3zWtFVoq5JSXg3XC2McfYyFBYVgbCdK86NvOmr+DGa
WspOgwv1M30oqs6bzOQxppcVIIy3bvsXbSTg5LmZkX9/g4RGo/Y7R66Q2i+o3jl35arQBkC4ROLZ
AgN+fjm9g8cC4LNFfks+L0ayLgQ6bNFPYmHrgdRxXVqkQzQHDBAnc352CChs7UUnL73FvAF5tRPc
C1hcZGQ1aBf4KSgR5dW6n2m9UWN3vJx//sWZTqswtrc3qg+wGwjbL2Qr7F7iQeTBgPy3nHNxuRYY
i+UvRWDtxaHi+x7YrrSIoNn3mddl0Ul54AoZQXyRZeaCJjdlVDCZb6axmYoSWlVYyLUouSVYgLbO
VN6ynhIgJZmreIt8y3UUoP0lA/4u5IJ28ptkunQ728U2ML6vbRWvgBke+wC0nbigoF3PJ+b10tzu
L/cl89jHUDWFCEDciF8/F4rN5HLXF98ALfX8ZSIa8hWuw8eAOlKNJmmHj8PnrRg5aw1Hx9LHs2iq
H92vflsk1tD984hOZ2ou3TEr1Mod32T8Ch/SBT9bgGIKPDIpIBsyYtapoy6ANiukZsN0UikFbYRL
gdPFC6aOJlYWS0mT/D05EXrQEy+B5UyO7Uq1RTJC4okpVT0g+56TMs3v3UEkAGNAQGfbxHmX4WF4
8y/OC17H4mx8iwO7dx58swQrlSKvMb+F/jhIweuXi2TYALIrVJARuW0GQpf29B9WGUwnWodmdJBv
GRfAkdWc3o6osfYAWPGmS9DSW9KkMX0vhiO3CEDlM2wzbeRvFvnWYGQN7j4lSrS4XcIRV4PkEelC
FJY9zTwI0s51HbFRjfREITARSapNbp3FWd3braTr2FBc/PBFzhvii+uPy6GtJ4q13eXykX1xgozq
8PbrG+8a/LEr276Uf5gh1IqONDvNZ70uHsrvwr3KxnHtzwiZm9QEH8M5LH+utjSMZStPWUIjn8Ir
NErON7eES22hcKjiMOA3eMMCDJo8PyDdqfWc1fX8ih2Y8pojovDJXvnfyeiaJMGeh79qxFmhbmJC
8n2TKzhIctxsUYWXhD/OeDHfiKVl26R1yiqxrmv/nT2uvAl8X3q8Su/CjFeibTwojmr7cX0qZlLj
usOZGDff/MW8Ppmqx0/nKKeOT3eGnWkxpvyZbuZdz52Kkq4uy17VL+svxmxUM9TOydVZaVDmLOzQ
zNu9iRW07esoLHj/sSJHLjYDlO+7QssfeSi2WWxXhY+J9Amil2WBXQk1MTdWdEUaFbOFdofN1Vcb
emd6e8L0rT5iF0DGe68rsKrGmDSpEY75EYEbxsVbF/TlXoQK0v0f0wp8SCl9Ja9dR9txpRS2q8Rp
eT2uuvW68UW7y+5ykcutVGSxAxSG7QsDs0ZAuAXW0HgjYhrtJXf7Fdw7QhfmD7O/KazDyz16zEG3
sh+Ocz31MtPRRYvM9CFg6K9PP0bXHBUGqv3J0fMGcOwVv3jl3b/JGVeAYlsEwM/6+DC1QT5tcAGD
JHccMVh40mzdHxGnDPjbVQdnqrXY9LV6tygcZPZBKD5Kj+zPQOEJvfv54iUtjaLt3wcJO0VHBLag
+9seUzGtpmKYUQ8MiWI4k0Q78FHoITZet2HvP3uNfoJxGZXn15mEIFeAqvCak0sMfOPgv18m1TM+
2FC6NhVWOsBKXYKkKYSOFRRv8fEasgIVFXnp+SJf4rRCVHannKN8zD+Bn5J2TyAP40wOti9yiJfn
5Lc7csGvS1zuTg9i2tBMk1YW7hvzRvXAropSzotYnh0AMHzaBZbWNrYh+FdQ+oX8I+XzTA8SfpyA
Q58OHYE2zlyZ6P8veFtz4QM6YXX1KlrMRxqjOG4pefPx7Ot92lvJc9tJmt92KfRa6hLUNtVAhTDD
7UHiWzgI7KVZ8CTH0rB0CojZ6rsodWPC/XNShwWAhhs7S2nt/zyP4j75I1LVOpjSqJvGHDhvNSdK
xAbr1OOun6i1TTOrciPuAaCegy2i5jZnyfOtwDBFmSLkcsGtOm5XiTFoaPfmSG/XT7Q/UU1UfG/O
FdTh9ow9k2EkIKbS22h9WrvOY6O4b9Sa1EtoUoNTLZQGXFJv3TagmPeDzrBnOjSKYp0Zc8xpXHm9
tOVXe9x9VHpx6tIi2HWOTLGw6pj7jGG+qwv71p/M6MdYbUqGZdbTr33rYj2t/YwHcPm3BTPKbtKZ
h31fJjr0mzH1DrrKUsqwCJp1GFufKAzuJ0KeK6pKrmLwAhrsaTiCpalfLdRQ6R45hT0XzWw1KOJ+
xyC/yTab59vTZzl6CREtu7HkjuFqIBBJBLfae4SZ/1msd1f6tqW23suTDKoiCejUaPzEwhieIxGK
LUdmPNmX65GLltFbRB+SOA3GqA/3MNTOOHqBylsznMZayEwO4UUem6SWB0EhUrTXBxhqgMcMerTl
eXmmAWJxT9kQWVa16W35V1L6ewEz9wdsvHdC2A8Uy0MLUly1N4zhcVV03ntamiKOueVRdi36zdYY
msUqMocH3g+6icizbe96PF08RqR6OrILcg2ZyYTuu12rfaN0P0jkL4q7NmM4BetU/1hAPFltJ28P
GjUrhPbQl8dB5NUrh70saIkiPAxK5kNY5b62z+B06OcZMqX0xY74KGTL1pyRb13Hwndd3CFFX1EL
QIfCzD5Sfb2jKFppNtJMCHhHjxywBYC6BaiXmrF+Nxi3IelgZIXPWtwe83goUHVaJ2jKt7u2bS3v
RQovRWBfPjDgizpgnzQXiF4+McaSHo7rBnqb/vUsXpDxFC2j3QD5CqnIVkwSpAq2hHxCTgjldbZX
kj0NfK5s460I5Y/YVL/HANUKdeDKO0xV+Bxvx5yWvf4SLlfaHK08IOeKoRRvE6KGz4rT89e+7Poe
30qHBmrUd3TAubcsryC61P8HZSkOtIwLY6eU3JDpRYw08zVdP7CRhk37eYAO5PHWyEl4Xx5KKf8L
acVVPo3rmmu8HJRq83HPaxtoWSvbIH9+vwPbWKuPlN7sOiKkS5EhLQFpKLRu+ogU4FnbjVeyGMpv
ZhruXscLbR5UvN/t97kam/hY29DwwDqHs5XL5NOcmPSKkJfqNbmU7IdSzxeaoMiqliLHkBWyFVvL
tpFCb7iJetmWxUepw2OsXgr25xAkr1FB1X49V4c/tAciceVjdD3eOVTQsozYhgkmMHFMnzYNUKAE
AWDUVXI5tKE0kFmtHWj8SK0l3sGvlcJxXxzSI94QWLwsx+vqszHs36l69Gba71YiTMTBDOQcx0xR
MNb2TyRGnD+sRGzwSeDG0NPTkjkTAdDxnVEqACZzAK5tjI06IWPe6g0CbtsVZhF3V1gZidbKYSQ1
CHxCrCuxNpV+6iJmh0t6g7EFopN8p84EDvlNDgq/8MSIS8hLOhZQgkZKAWPPwsTi3vvgcM6vuEdZ
ueLCfCfqzM4tkJsuJN59/mH2FmaRnsQl3ElKUbi/a0dmjSMry3832IglP6IED8RagdPwD73DQFz+
88xkkoEKO6UNv849aCWWAXondm10drRJsl7zL/BakxO5pib3gT16zjO79tx7cPxcoB+nD1QHXA/8
6ggNLxnQbnENtxus1vMWASWtGcvXpkenju+WU3aSfKB3KNjiK1JmaB+mOED3VYfyudNwlIMP3sEe
wa9F4c4lmsHmQoFAt4vYwKtPSCeI+JVb6V3xnrBtrAKmIM73PJIF8kc3yO83h+jEKuvfXS09u6vZ
uySjKW9G/8yKhdj+IqeJmClREBoJGoGzEJpxlnQ/8qCBMzUDmDxJndncQDUpQvBDmvYB/sufLMJ8
t6a645jrTRnzBAdDz0lASb0kQA4KjRek5KvsQxMguvX9OZey+zUw8lvNruUp+THuygntruwB8FjE
jGYY4qOfjCo3yghNNA0MqzIUJU51PALSUr5syV2YLenUI/7rZtECby1ekSh9OkXIH1FI6rOI8YPm
ayp79ngPpp3WJBMwI6Wsm0n5Y9HdtKVYcrgmGhZPlIkHN8zEqnXVmF+hZf6n1QU6HtJL7Ik4GdJQ
5izQzPHM/gQWg0i0OnsnsjWIkECo2YaRgCo01qtjHqU98RWHuQevRLe4DoCn59fT/X89PPrWnlci
vvDRDB854/UKLINONFCGBEQ8tQCvJmVwW88vT69tmebhjdkmIlY6VeraoO4MVfVD68mVmkVTUnyz
0cCUMpVFEOnkBupIV1Slmyi/AQ7YVftMvvtGcvUK6rgwVzT/cdP5RJB8WnIobTo6QFqeaVyNzSqm
GdPkdcmV7sZ69ecBpu3amYScHt7ZyHN3Kr+mf+4t7etzQR27zGVBkaKY8G1+Vr3FKi+7cStfQCFq
/AgyrlmAaMP8iHFed/1dmj245QzsGbUkMLbS+x1OWvRKwpNZ8jeQ8sb1wCqxejdNQyZg9huWCpIc
mhiMe7hn/BYSEDk8hbSlLzqw1FitHqvEg7zPR9+uCSR7ChO4SUJK1C7BQ/bPAtEOp5OX+uqQGf0V
heYCMknktdnn81JyxYoDV9gYU4VPnZB6C9SY+ysiDETDHfsjl/tA93Fo+zB28yy+EtJ6OhhZYgfi
oI4rqaZYypk1NbmSwkGvuAsnTYj1QlASW3gpCMZt8S/6Ui8hKZe1hci2jhXgg1bjThltb5KW8iPA
et3guySahqw2w4RSWPIDihwlgqVO0H91YaTRRLwomWKYVY3MsQq/gzGE7P1fIbeuL5dYFrYXi2du
pt0e74NZhG3b2PlfqQki9SaFUuc+RZT9mwWCsh2CpSzcdTjbZ+YazT2Wf04gJYJSBq7GZCWlqoVZ
2KMWO8zo+aj0vHk2bUVxYpFaUBW9btv3bgJ7vQ/bsCMEo+xXrHGdbdgBDK3bDRSC+3+7039yqoq+
7NGe9TVTsH3icu4qWOCCzZg+xI9IZz+tXv428cdHlnpuyCOY8inhxSGhSnMxoqZiJegK7UhvcDqq
AizaRggvBeA9MSJQowP0jLSvI8gfWmf6Wpihy4Qh9CKfNfwohSiNgxgj6IvsdNj7evkADFaRxUPQ
IddbFHdRQyYpV+Y5VZc111xveLdrQtSErx1ZtuqBqY5k1wwxhiROBL0NRmrIsbSTU7ayUcdoRfyd
+S3TyeBULzrTeY/in3wxVnMfydF8wCQLnxBgo9hx/rrCLbx46WrfXaso2b6bB7+mHwVR5vAX8gwK
ZEZ/zeWidelBtK76MVMjfreb5wGJH3GN8Nbfi+3+/VJtb8qlaej/EFrmkVhi2JFgEBFJW36ySQR1
1/DU0jgZOBYcBZ3QfnJURRUgt28QpOyLkOTvvrGkxwKVCZYHEwgBirr2yqWPlYhVrii6kCcUVjLq
0hdrU5tYHPEgP4c9ATJfzsrabqsXsEFi3jrKXhej66y68RpZhNh/KKZMLbijnEEGolYLe65jYC1g
wC2+qJJKHEMW5j5b0KkFtXlv29ejD0xsYhiw7+HT5AyfAQyoYOsqVvdQkbiRThrfXZCfyUkvkhEg
DsNYlleLum/tCYX5nITMW8gneXYTeIYSLoU49OabPwXBOJXga1RyEdPF9CMzeWBxAWei79j0o4ly
hkXmRqQjDh1J/v1/HiF4OvNGG9Kp3+KPVmD5hh79LggdPdqnWPvSXoHCiW2sTKEIOQWyHcc7o+Xc
lLtSCymvHSbtxQ1XhQ8Mbg51lkDFTQk4hPazg1LX10ILKNXpiNnVZyzm1HyyqWmRnVZ35bW2xnw1
uXfeagx78xUHZxYpO/Run2wQ6h/BG9qX3wvoeT1qXFb2rCjJ0LJhNOgbb0Ly4tV5QRw6bsWjcIXF
hqcnDDMu7P/VSpIZKylAO0vWlJt8RYPOH6OosfwVzvmQrSrEflp6dNYBZSPyjAnqax5VcqbhdCnK
0JU0irliuuE2kHfNh41o+m8hIe8BgjUxg3h1CWP+VtWKCrFz3c0oPPYcz4poALv7r4y2FGfqYSB8
3AcImR7aViIxxh8GB+JE993Q+y0M4hQm5BInS5F7suEfz2W0eCCgwnLj5WB3t2VbUnWxgzSzR2cy
2NfRH7HIC1QsHgkR5awmb6p7HfokeKAjgDQKI10aC8RhgPl1sBNFPMGgSBP5ddjKtFyFFQ5W4B9u
BYt7F6x4laoIK6MfGqPKeU9DbctYLqc18XogiKc0DSk8py0a9SnemxX8GDLkLNsn2K2Q3kfO+VwL
05270D8dbpNYZ5YYkC4wJp14PyUrml/nB7fi8l8XBM4S7K7uVIJJ6rv2lutBvvpPkHZzkUEMMulT
6HzHg9fr4w3QRuAxIzGKJXTHo62C/c4gYyB0Ttxv9XDuraVbo48HC0BjgeVohoOIl0bYraTgpw80
eM39BHAESWZ840RHCACLMeeRtf9B/nTPUFw0M9KFbzjw74O9mh6paTNBqdH8jsirM9sT2W25rqaW
PE+TkJ+NeRz6bEuQlU7KnHm99kGxEDY/wiq1/HYTA7qBpox0fTFfETdZo+st5PJR1eXhDrtHygw3
CK3sW0QFdA9beTvZJDehFZ9yhxg6aCRnDmf6F3ma5+62M8KkTxUqogJQwPzULonnM6zYIXZ0axIG
6LSnHyDtLn8+LIzDb8rMAULq3jlppqLTVsdWCO+21EvhnkyE7i3Dyx6fuGIFJ1+RIwrCsufMS5WM
Y6Aux+nae7Up1TvaznGOPKJ9ORECDbwQrFBrGdu2PZE7BwLGoBPy3od403z9SzhZfBqsYvZQG/kk
ItO4oYOReevtl6r4X6hL0/jL16V6u/YqrH/eSQZUBqKoZ1JQTrNj/o+PKjt/csvS1Wd0vdVIHeKo
FfkhM3LA+dumr6c/6jP9sjVEj8+5YWU+FYYv+hThnjn74n75Gekz49ehwOoADl5l7Ijw/4uFeEzw
iBlQ9slLESBhNfusoxqCvqOV680drYX/YhSrFxUoX3AEqvAXRysht8oWXsTKApdDhylNAUjmH42B
JhcR5LoX7V/fcVaaJRntI7LQZZGFquCK/uGQa0H0yBMPoGp0CyA/ILuPdWG3yi0K7fYsYlQ4r0Uc
wFZh1uTm0L+YBZOio7JwX7FwCvNNgweX+m3dzLtbEAuhZIb4J7e93ilvAaKKT5m+xasF5oGw16bK
FTF2omRCI4Rkvg9iJ9N3cc7//XzDp1uKdBFMEtwL6aX61Ex5sdUx+sQdWjEM7pQFwfsQ63eJe8MZ
ISMfozSZ6OmHYkMci4ESfzua+MKxyVl/JeWyn2PsOIakHtqgYg+Om5EL2CkeAHS+qKJJzRtEUMG4
MUnoUixgELPCjchkIXgVI8kH05pqM4M7pmTqY3Zjyh/NMmZgyWCZSpvRFQK5svWeuWCtX0BKQb6Y
gOnNbPnfmb1bI522dPMbI3+4f8+x7mF9lrnePRxv0RNx3AKuCxmVkdqm18UJ1KQ5UGSisscRHsNt
V8fWxbCjIu/vsRN4Y8k7ycxlDu5sehyQpwEm7/CGj6LeqN2d+V3dmsg1VvWmpVGagDIs+yspOUfQ
/pDEdlXf4OjfYqBT+dSYHQE50OheArnHrEeJj6bVB99ZY74ReJ1aotfVuYnzOm65GlZQcJvMRjuF
TC7I8kS1BonAhQ/qBzTX3srTTTNr8LDKpCBs787rad8Pd/+dg3tsg0hQS5uNVeLPB85xxPQSY+/I
16yZBipcZy9flDmGM8/dG2HmJBPaSd5G45jqK43xfZpF0LKwsoIYpduXFjKADuEsmLPLlB0F1226
LC6LNLyfb5Bl7NWQNzmiyJi5BSc10oLGCYWB5hfsGDwBDI2iF/cA6Xxdq2eudJvVGk2izRVznnNe
+jHGyV/1CMHaX69UmxSTYUaGXxTTDhfImx7Ai//pDLAQmOqFcxryUsyYOA1uETX7ihbHrxvZozOC
P2q4rpGQZP3xHeAyhl6CLEEqcDrRSC2BGFbEix3LdtgjO2e5eKQkPuhdSlRFCs5ngXT32EnGL40O
Pa0121HAMXLBG+xdGp5ccWYeoh4ti2qPIpiJR78MNZ06LbZIuzpieZJoBqLQH6QtU5MEVC6DRoXa
F4tpgr3Q2GrwDFrWoyvuLCNYVwRMsNtR+wfRVFcDvSdkUbTCEl65OAAwf8mAGmkit0olKz7JMrv3
p5Yx4gFC11lEHg52CyjBQJnZqD1hInFLuXSaLn17coKJwV2liHnZm9cntGgSmJqyX4d/8b3sAx8g
UCys7VZVqlI3A0clC0ZceySTgzmu7THhfIc9rOTdcL5nsPoQr1YZGFixV/yx/fVj3jUkGQnqpW/p
/GCf4ulGcbbXH1oAgJhU4CmBTFfGKvG0A6QTkWJNxEGDFd3dXxu5RXDJ5RPS7nLJw22IwnIUAlkI
dTU8ZvbQy5xynganLRcwIZqWfEZ1xKPSTgibUTb6LQDUKYdWrZrFRe/BozdjAiddChJP2/2nvnYo
/r/R6FUvii2Ufgl055aud50q3KFE07mO4l3dmqGJKD617nU78E4MZcDurfTsIOLEKqoLow1wwxVk
VWAp9aeCDswoOB04ryC8KDgGjw2sl/XHqBhRyhstVJfGdKfCuRG4rM+NUksL0g6XYbAFR437QD03
he5wnNxQyejlTHXRhNgTCZGronVT4T889c+4+InWQHrJb5dMMXYtr7GPFbn6XVlZl9xhqMyYhDpC
cYsYsz/t05SMJqWm//IkdH9/5uDDK6RIvm7TEhQYpBXzdJtaWowRsqjhTbaiFsFKqMxLzm16Mg/q
mFxI3cYB5AW+Ti77u0rtUAnL+HXBPuc7ObXXUJEINrRKrLI0387rH6p+l8wM04h9KsT+dwGBaNun
40uaLyWprYURjeUpGk8lHDotyUXhx1UefJt7PFau9u/hGJpAsj83LtP8SE+EvOl2UYqlQHP3xcZq
S42N5mT+0QHOHJf5DPHVJR74I5GxObrnAihOlFni50TN88kyWUnQx5dys2DHLGYthIx+TP0A3og7
MPESPaCuo4HgYd6YAbvaH8HjVb1fZpjjI12wQ7YtaBj7vHb3qdtohnhtcYDUrWml1YkQbrN8buWJ
rD062yLwNXLzAeK4AFquMhwZ9fnZDI4AYTtRXnT3bXdJggKv3SLdS3o2a3S6hDVwmQ0q5YqHPsvK
AE/J2zuzEHqzvlfDPYxwez/hMEZJrpBjuJBDjWZmJXIP6N8yGPlKY6z2futn6uY/c/QT+MPAgZat
xmSncAlDM3idZvZWap2xcTGmP7b3wRqd0m/8lzhBlKJs0J+NRqce/EyDvDvNLKnWAF9QAmAWO4lR
SzPbks08j3qPhrEFM0WceugIeyIGDB874ROXsIGOlTa+AbXo1YZKDMj/jgA31rqFHuv9fqkOxh5K
i/uexkmrHbtia8VSgp3y2jkigqchdu8i3tK/AUG+5mHbsUqZJ/4G1iyPmpcwfRsMJD7gGN+PFbyw
zizXaMEmORnq+uKlfobzKr8p2cfqRiaGEypADMa9doiQEFBQOo5z9JYNwO3fluAgcx0wctgBcr0L
ae/+aLbrcu00i11gG9wEgLg0iSxSROkCfFg0QDJaOYLJaPySwqshm+GBCpxdnRuonMa9Eg/vWm21
jieWHUfHwFBklqLDH9s61tjnBmchT2zoXy+CENSMyYQ0I+GEVNOneAsmdOv7/sBKRd9ODGZzzxo+
iZh6y4r3/rRF7cnS2jfZjAPbNDl3VqmZ7gBQO1ejEsC2cnJYeGplw5utZAoEx2F1xDdfQk0QRGM4
klEQflH0YI1IEpRJQwoEQAbNt7d2yP4cBQ6iNjExia6CongtUU4Z/uGJ5I9NU+HaQO/ifUYItmm1
sZ9NWeGn3Es3gnYJ87EcxK3dyxh24gtYecomqk3ucL8FKP4vqYM/T8SzHycWmkd7A6KJDFFda/j5
jFelcb72HznAtU48tXH6TCR0Fc/9GZrz97IcOGx2JCWGPKteP/mHbQp6NMfKcG1fgufJmug81Zyv
CXKVsBuQFBkbdmI/k9Id1EhWXgJhhhqnW9bxepfFrE/9cI053pWfdQdK1/ontb5A1ds6UA2OkTsy
i/R/oRlK5ZG2G2/NhbA/H6ayX7f3lE1vaMUXWQYl0K0eVUZTtVDRTRGSbUc9laqOfFHguEKBWIYX
cpdr5WFZdk6YxCoSkZmkNiSa8BWpCs9TS375Gbu4B7J/74CoiNEgU+iSGuZ6CUGVemPyvoh+sUjt
kZ3a7WQijUNa60I85Qoob3b6fcfBeHSTvlBJ7YaSC0MocZPtvBZjAZrZcHMOooLa+/TeofZA6U/N
b4La8O8re0T5c4BmVlsig4Rybxq7TUsB9dkmdUpapS6Uxkp7EjyvUUymSh+CnTHNAKFjhPFODes8
NLhhH2L5URu115JhpajCUVlwKPJRC+rPqwSKIFOLw6xnZ7wCsCL1iTanqYbVESVLB1E2PHJzr9tv
rooe6ZKLUFFQABl48/k2hz+pyJ8OF0R0HsdDh7UUSMsZhLdkd0BXuF6ts846eGcJVX6o94rO34+c
cjqKuKgUfKM/HhJi27qfKnAezYUArAyX5vIJjH0AiLIVFFH4pfi/hQbkcmQma+wv3AhCrScyYE2C
a/Pkg494IGZ3QM5fpvDy3nsQBctC+jzvB9qr6uzEL33SVcH1wmW/jJYlFmxfena9hTZkE0SEpw8D
Ts75lh9aYN9U+f/mESozWf+dqsb9n6ynbdzbNX7TYUrWZEznjGB9E7mHH/LOZf3T/khDPeg43QSq
P3xPjTDp0IOW4xTjGEeo4bJ85HP/j3nh56gwuGAfOgWSqGJiiOE/IU7UoZalMNCek0lfljIfK7nj
Cf/tfTgs/lAU38dthqZoO3CUmUktjZv97VjbnQScYqY1oeLyb6uL/fwcK6x8MjzqqLY1OA0T0Zy/
/fZoIftQUnW/oE5P1C7OCgIPw3JVEeDdOZHf08JD+mSByL0QkdO3wzkkWpwJhD6XB3jTp1QdXZoA
AAElxw/z1M9Otcr083+zzlmH16cQGCbjpa46JLRCBbmtcnxIOTFLQNgPpAaj3Rok35NM7rq1TFfN
zAf79JyChczG+MPwoBxmvcqBOFfGAifnDYgEUTfHeuor3n61aBTtLSr8MDSidZ5dLXG1iCqtzPE9
94/OaE9NZae/rIbAgHStKeELQM/8CkqlXuKfXVLvecacUdTupE3xRWwrsO8vatrzNNioIYQvHiHn
FS1e2J8QyjjTofC+e7SW3fyAkG54iVUXb/hGrLv1BDDsExqWWdMe/+B3ho1FepJknNpmAdGAFrv+
sTSmlVZ1HsKYGIZVREMiDA03bqojEsWcycz0icppL9ZFMOqdJm8IShGoG6TNx118ZtW90CvH3Fzc
c61FfJZdD8idvx6BMyeb+RvEDtHA3loixwzb095GQYhZy7oDeSQC7QWCGzODXa7T03Y9pfyoU6gY
h/uryJQJthkz9u8U5YFvi+HDP2PXsR9lcWHbXNkVNF1WmnnCyLmqFCk0LMgFHhTdXUgrk+VtI+Ku
Xo2Jt1XNdmQsEzGiNskQPN+Q4MFuPA+Qsk08ZvblUwFRy1ba9u26wxUfsftsYI2g+rlVcZp91zo6
LiLD8z6RyveYA892NY1DreuLqmGkuUfITwJ3zmNLpqbeIc5ny1DFQ1ktskigO9loUr7CZVYy+Eyo
FasxSBwcz1nBFH4AoAiK42NiOwuu8+Nn8uSH7i6++QzQQDxc1VRnJst0RlnssMhqZ+Gru3mJBmqK
VkYObK63bXWOjdNzAW9yxYnBYe4hNY2QDl3grXybsySXvVNm4t/7KWMVMH7SaJG4d2iQlChfhwtY
hDm/FP4glyfk0t19sBiupCPcOPlFn0J0y0xr7wJAa/mj5f9RcLB6NmRDuablnK7XshPNAhvMH9/Z
yUkVYWY7oyCNei9sQ5ri2pcI4TNq3vwvKinBwNJyvgTWZ3Js5VT03int3U4iZx6t2+8AsJogov0X
BZ4Y4v/GjoPqUPKrEcIgmA9u4Gd8JVfn0Yw4ba5wmR5vpknt9yvg1eN+ZwW0Rcyan5pTbdW92j7Z
CFyKn9a1pufGnGJphodQGFFaamS4tgCwAPrVU0OxfkZoag+uPs6kM6PHCCm39MDWUbWaM/Jt9lNm
O1TtQ+ZcWOR6RmDSwHj7a8rqz5WyLszoWsliowAJLMV8yKsMcCMVwuWeUw5T0huaY8Det/BgnFMv
IymsraHhDUs2cU1en4WZ1sT1xK1kd9kabcjwqdK2QfD5h750uRTzmJLHvW++juVooji+ZE4Hecpn
73StlJEK/l6fD/VE/qvTux167rKfD89HmvwgrvPpRCqAz7exyfz+V9nWsc9cZ0qjXOAcekP2x2zB
8zytdUd6hDXH48FAc6JZllhDxhP1vtqkXXiIBr9D9tCSkPOCkjcLbcRumYSc5gK+IZJg5VioG3Kc
rQQZ395yftN6lPn37/JB9zLKrK3p1blHJBMOLvHuayptqf9uCiX0SXCD0hwCZO7Kub8PMm7plwMn
gAX0MFnfA5+EgtX3K2gailj2OH79PSYiCGj0WRFnZj3w8iHgKziCgFi0J16K43iiJI02Jkev7qcB
RueaDVxnCn1Zib/oqHK8SQrLINylk5+Wo9VOdrERljWboo6RtxITRhJB207+LvdUZRVzvkkKnco7
Fv53tG5JLpVE6bmJc2AeZiZLfqfUgRsjwGLGgUR+RDGESnP3YDzt7eoneqgugRPK+MNT3PNkcmqZ
yLexP9cOUQcjRM5ZF6BmurRMqsGPpPw3qjHFXiZjBNFex2uyStUXkwAUFT017/wA3PFpH+mEGdgG
sAenan5tIxQTBLW1GNxrVasqn7vcc8i1LJ2ZZg2qiKWYij1hx3kU7famrln6dyUEk5xehq+i7XAC
ErnyMzOcd5Ij19S4i0IyEaj5/AoY35utpRnKy3GQCK9tvSQqVIGaJfZJwCC/VePgHW2bA/FZpemx
uLXedMmwZG6nKOBbnM/Lj8udlV+itrK4viZvMwSbuWsx1pBiEfpe/3UaTKgFuaFkmJnK1Ssu7yyQ
ypWLdU142FSCESFff/sxz5CacYIpKQZc8Msv41mx7P8dZGKusA/DVMTdBU0jSFDEU3d+4mDo+1dw
8+1y1sY8IqMv6UyT/5f3vJFevzHOLnilWgCuu87uNjakXI1QXjppUW1oRSgAXN+mBJY8m/KthxdN
GK/qzWbPmic2moqn/RE503nt6vKox4c7YUmjVdjFLgOeZ1/BeLfRiLocw/6CwfEkrV4gyCaNjR9q
DzyZNW5mTyhUqxi58WAUuDFTQSb60P3ZjMd7bHjglHKUGWMhb/K3+4d1Hssitmz1n25BmJgmLTbi
++qn+DysTIe8n4xHF60xV2pAeNja77e5nmTAHPCOZphhsntGDL7Vljs/kmifzxf9gKziLcOUGAKx
Wk8Tb3C/F98IZ7PypwJRA9Yhcv/Nj357b9rTdPX40yMl22hBKL8EabV8/fjNPI0dZSiipYaXXDuJ
tpG/eGSyWGsfvju/jcYmHZ47bGkWCAhDEIyzWAawKz4G+/csQHyRHrqaPrjJMF+WaMyb2uVK9sXA
Bfq2FFlTaIdfelwZ1YerRlIDCS66CHra3xHgbZYiy3NSHujTLGoeTG2b/zsQj681ytIA066ivIQN
u3LOwfdTO5aG5fy5Rx07Ve/Z9cvVwd3Q3bDwWNHHVJiKUVWgj96FzJjHhc/pUNlt7dXwyWj6XNZy
GCVXp5iPHlSv1qIH2LZu/LSeCVFP6q8PjwcstD9j6CDKhPuOuIuO3jV6hA6DawEiR4/MXSnjz+/a
Yx8IarfRGv8OhYSDQOQHnrVQGSmq3msu5CXJxTPvcQ5mpyzbJQmXGgEaXvErGmgnNTXKiKiHkfvH
3NAe0AFOb3b04dcyregezeft4x9dHtrSS7wCwll67vxFh0H1NPJ22xMTE/Aeb7iMQzrNAtev/10W
TxmTxljWZQN9MftW/QmRELIYkA9fr7YRBQLQVZpuYe2ggUxGYyjfjXVjxNaVhRSyC3CrjHFvR5Ns
9c4Pp65skZDPAVQl2pafFZSU06y998q9BMe8fdufXRH0HAlLMU+GiV2Id2pERmjpV2iuen8Rly2h
I8HD/YAaQNod7VEk14F+aHAlX4Wf2YewcyTqp3NHwIKrHsYdD+An3TY4mx5sI4y3fWcgrB+W4Eo+
TH1MOXVidF/DmnetJWLF3H9SDH9BHhaID8Ch1KzoE/z5+U9nj4JSE03DAV4/kGB4Mp5W1cbSiwal
5XRwojmN8i+DJz3zKdZm7ncxt7N61bkfjyIKiSczasfexe5dfc7xbIMffS5VI8Vz6dxHz1g1P2yy
n0o2RgT+sYPoGdMXbPFNxW5n/telxide0fXWSoXdXTgWl1uWmjBVe4zv7Bew/BtiWHRyqIs0jO8R
h005I48webQKOCeRckAkBWo58UKRFQju2ZckLGD4VZZTVKZDgfCx5Ef54KVfEdiwF+f6nG6P4PqX
qEXPJ8kG6bhAPcjUlV1bBnWKHlSRVBb79IYVFJn8bspvi+UXTx/qjjfiDuLk8JjFCyXTgl1B0wa3
9TLpPFEaiaq0nxI4sNTHYb29FApg4HpT01j9oWEsOHzhXy7x6q4ZHgfW8kqDJWLy1CtRuwcXAcQg
LfzqsEITGGujPF6JKrRbWf3oIgyBjVpZjjQd0WNXZThJ/FNKljh4eunDXi+RzqcoH6Kvt99JXRl9
oqEXV0tAA7inb/ma+Tjsicn/AEisku9GUyGNYRprYeW1RTBReP17kq7vuve6j5mQ5J4Qe9hfGp2E
T1kPVQod8dkS9b4eXrfT1Unl6M7ZVAOLjSt2u4z5VQhcGNa95xDDaMkS5pJ15V95b5xcHHTMbuMW
yfMWo4DG7trrBWG/yfkGFr4A5/U/Q4mwQwAmE5dVey8SsQ+SfN1Dk46jKmvwZBh8sjDMdrCoA183
8fF70gQxHP9L7KhcvSxL0WTM8O8rVBrRvm5Muai3gKT4Wue9b5IQ1OhDClLPCu9trWNDjlEqLc2s
2ERvSZBmTRyXJN6ItLjcpgXo7nebXABWoGtYv/Md89mZgy8sKbWdjL9TnVJRKyIkVA4i6wgsF1t5
d2+t3YbNhZIjNpxKesK2HfV07SFcAB3xopu5ofT4fDs16h1IBPkd54Vm4CEkgQZeWv0WdYi4IBlW
97gsE0AzV8E1xncstfeEfb6BqftQu3jpneDFzv2eJcHWpzW4D8eY5tB35AHCy55IVZKT0dINrzN+
DL8Gfe8d6Vu7aQ1t+AjotOZ0DcZtxMQbSa2oGyUAu4pkqrhOCwqdZQJU97lVQsaCkAbOypfs5Yn7
9zIA30YngWF7UpUlCncgthkKCsnp5nyqAy91UtQXR50zQZbTm33RDjWP6qpiMY6DBQdiKHCmTFSP
lis/Xn5IiUvnX5e+G5b7nv/C7CyqdT1jFr9+hK32G0TwRdl/Vf1nLmiTLb+fHczQwY8HYbPigxtY
/TxcK3bXyk4DoCk3x6RT56ZqQWqnAZTsMjlSdc89wGuPNqfs+XhnUl/iOFcqos2WM2JT/ABUTH0b
LoJUnvwUuc1FLXlcZg1KEnldWlSX395SOFMMyLwPjSkRrPrNZTeLrTdpJbpOL+7JFS1ICHPvyrh+
OLtRvpHds7rKmFfzMF6dJXp8bs0MZveMjSzaL3noRronnqtgnAXrSVQgvs8Rg4+m3loFrIyCqEF9
zSN8Ece6gFkXXv4lcYjjZZUAKQ5tKJFFvFLnxhQ5mvvqHVThNimFf+2gqXRxf2LxSJpyHFSgYpzT
xZu3WAS+lOtVDHrFVlqLM11BbtQGD+RKQSKEEn3GPgJGwJPhzCasuI8jPDnVq8HN8vsi/fAngAbg
eTAtP852iEQGiXA1pdpcFv4Uc+TJS3wpkrtTmYPmrkD+J9bzbcVx4ZMakzyv6HSyRHIrDc8uvLHZ
AxRvXuilypt2yIU2Rh3g7eO7BpK6skPFMBQwgJtMIeoNoDtBZOiErYc+U0Sy8jFu1A0OMjl2G99g
IA7g+XBLxN8vNMpaPAo4TKEpPkyfE4VuxYMbeCUcGQyuYdZeHYOTsx493ZK19oEJPYIxlh6IXf+v
jUhRhFhgCzxrj1jY3fXl9n7dQXnmsWvB5iKaiMApJulm7bMMogIPlkERfDjk92QX31XPgQQ3gsW+
HQStyTINoT8axFMq9Wf18kptc3ZabgWiA6iCn7UTtWhw8Ek7FvPN2bPTlGCfMK6vSLNQIxAksJWn
P9uKdfRU2coxo1st9pZCtin+2BR9ff1Nihm+7wkgZpMyLAhl239wVcUh01EPUkJZqE8ZATmMVWKI
Sa43oyKip6NtSNfHNjIRIhBue5RLHIXm2HE/zGdaYfx3sKYBwti1T07QFuuKAIHuH6QY/55WWrD4
cXOVq9ZznmOC8MyCPuAb3fUknNJI79XSNc9OuLd0+gBVt1tTYQ7CCNp8qoWiPFAAObhPgzuSRigj
BMUYSJc+0m/iGEq9yvmELhb4lcxAcRcSqgm7SRuRiexFSzOMsAudL9iHg+EPQETHUhU7CJ7oeuL1
TuSIxCtids0OzdTXy57hbBagYQ0odaeHAy02XOkokAOAtqryhwgVshAbmRGmcKMvPkSjHYRtkW3x
LebNrPonyeXupC/cwp3X932LZU+mLG3SKZ9qc5ttdcQ5Ezvf948lB3CsXl17qzvWfkggc546cqMc
7zOoQ00RXMe4E5ZQ+SQMq7dpkJbYHSh4qfya+J+iFRMhlmE/NR/RtqByhLvIs3JfHVO7u0hq4OXV
ZRVkJU6btXg3HJ16D4KNfqVWcge7oRAlqwtee2Z0LINEv6PX/Wmn8xFk5rdjoMX/i2tPBRHdBuCl
jmfhK/Et+EDYEGxFCehWtje+rO40BT6VfQmH7buw5+DuwLieaflHyERoOE9ypioYfj6Eoy7DBDym
+Y5ucg9ERfnfZkL1gApAbAT6Rdb4BewqzS+9YY7isqBM39tmxKHvkjSEHE3RKLxO82wPo5CClUAb
aJGjYcJ3+5LNWUMyrrtnjmxE8x3/Xj5/QEhXQxCXoOypoyGiDnfH+z6R2N16e6ZWrkzxk6eWy8hJ
wfW5/ZAvwfhGMriwTS8fT1Mg1Ob7qtbUJuDXHekd4qKOMc3RGCLWhNBCYVEYOxehrmTdvsUv9dGY
jgq1OROb4LTE8imTb0xZetI0o3dGhLIFXTVWeratMMeALTblAy+oEBKRJHhhyjzxG31TclnZnRwl
e9NxPYDvjB5sp9FZ03JZdQBVkgH7u1jdmWQ4NLNzg3AFWB4a/qSd3+Ll8Ts0dkMWiw4sEVHyMhCl
NIzh5wlchukercqH9IF0IJwwqEM+rzpEaVkbMsWQ05OyXbPG53pqVMkWP/tnDV75IN6X485fto8a
Oa58lczg9SrQP9gOFQ52aIhBfeDmVXOwBvqHFrNOZU/KDUdYGEg1L+psEQU2sfSrJTZLdynUYbyf
26sJXllDW8xuCEva9wez6Ym1+N/qVdz+yA9teHZ6ZjpfBLnI37d+ZRUM0ss+1ZGdrsIE08yLgNrr
9AMppDPyZ07cf58p5rD+Sg6ZpJ3pjdhekesX7B5dVH2G1WGsnmloeZJv45ihutyHPbSyEgWTq3LT
AGR3Rn3H29aVjY5pQU+8XivCszBbiWHbBTvtl7WqixvSgiKiBR0jdlvTS3yb57W6mLElIGbpDX2F
dJUCe8SGeIWILyDkber7sJr0Pj0Huk4DgC2Cls3B52XdV6hWM3Bo84QibIzNmpDD+yIlrkmCSwbm
WUoMi+mh3N3vpft8BaIMuVEl8qKiA1EdNVp1ycd5cgX3DEYzUi2A1eLsQQFSEJIWo7aoUlBMhkDL
cwSQzbSwIEMIXzmtQHQ5iedxmV9DTICOlUGZiVlcltjXDcg5OrPmE4pfs9fXgkumPc/GgiddUdH0
gNKo6UoeSBYpAD6uV6CzaUkRxXKh7tg9GiHXITDhvAKWyaDaE/rP0T19psq+Fz3eg2uOQu5WTR2W
0esf1WDTe9VmARgWJT85EOLTORTL4gDIXtl3K93HKJEWX5RLuStFc7p4qXeb8c00OWRetRsDcb1W
153U4W1I1ii5+9TUwfr1pzCbiUVF26GvuIjQcuUzDd/dJZMZ71Uy7Kn6+E8euL/mlGTnm9A2IEXh
GGTs+k+MFuz/9Z2z0J3peX1r8bIQqIyS4dQBNv4Pl5ExFZCNWVIQkb3HAcRu4RrQbJCvtTm+sYhi
k5stoeU9ZuCIyVp6gqrHxLIgK1VEWrihU7olvrvIEHOCf8dcE0tRN7oCP0mL8mpaJF/4tmd75l9K
weubJmZMB3Pr11hhaMIfAMqWp7gmVy6lDe+Dh5HYAn8Rhr6qObh04BO3sVHFj9JC+wv48k1IP/j5
ZZnceMxqtayU0VffJxGrfINE3JlsImF7J8RLEAWtHxMBUo1Y1b4XE7ZIRynzb90zo/oSmsa2Uq2M
L67D4cgVI8y26dJAN/g9UDVC7wdDsFXvrnugZiDuOVX4WW/fHFr6tUoWRc6NzgqFuz/l/3xgcJ7e
QGWswX1TKFpQ97nKdycRVvzDli6G0/azTu+Mcs3bcKEVQAY6k4iBaK84DfaBYtx0MCZbmyitlGH5
L8Gz1F6qnG0gjbV77pwQ+itdCiJcMAkALZRfK6QEaej1FDPUVd9OBTQsGENM5uFYTeE5b9A+d8lS
mh1Gw6V4+YflisA94YsdHbhihnelvODIt92ZRGDG10U4GuPR477hLFNzRpOsHr127fQr2dlwq9xe
ftmWv25rPmurbpG71G7HQmWYj56WCCmu2MtavnOsgwwWs4y8PBCrekrFF9sVA9+an3AwcNL/mtzX
o4bzTkNewN4Mq3H1LRpO7BuIt8jWsywV/GTf5NnLZCPc5zEOsV9GAJ0qWBIgH0ztGgkdLtd7OnBP
tbfdpf+B1L8jxc53/UB6AY2MpT+7EtwSddOIVZHW2eMjv83xYrX45UVEIv7KeweL3ovGIwIry3d4
oTXPe9/jPXVH8cBOzGG7xksSEtdDQukyfL5WNQeFwsCjzdeJPZiy3jj1OQjr4IfVZS3xi0Gu6UH1
WC6mrP453/HiaAgmG42DXyyKYMVEPUzD03veIL/NrxcF0kh2lPSO5hRAajzEent6LTsu+Zuu6FHB
0IhL07ZG6WhhYhMYe10FZja0eCHzzrATr83gsg0wfY3RcLZOhnXE8dmdam1yEU3wMtIeoJQ9Y42f
s/f2JZSTwE4VfWn1ryFSTVPhQAuV0gEOou3vJhtNptSbQ12/QBfoyqh5bxmbgD4g/69JGyQb5cqj
+8S5YIEDRBd7TDR8CSEHXBy534eyI6J36ZIrRFlEKvKo83wr+KBknujBZpB6C6lcXiOVyYkawiAK
nr2Kp+jEknEQniwzO5H9ud6e23hM+vohs6z/vbxtCTL2KgOtvhahCTEgC8FlvDzlfzcTGPHr1aM/
DTLX7Z50onNRot4QZBcwQXZmITBD9n8ftXIbtHHVw1Ucb2o3sqGHIhDCMb8iT+/n4iNKJ0e1Q46Y
y1mSgA/QW5HzMSQkqYODlSy9sRFia5Wt5rcs7jdwuUNZu/YWCYD59l7ePVtXh33mn9mUDr129aXF
F6QAq4rZqa91t5L7aNosag+dfE3ZgJBph0JjZVfKAhtocjBy7FOI4DaIFuDLi7boWBt3cfmjAv6/
U33L5ELyUYHzEW/r7nMVr9Bp/Fbbn8EHfDll6F/UyXI4AjuyKkcgSb5eUCv8YsV+q/Q2jqzugeWq
QYWoFwP7ErstyReYXpJqhyYpeLSNoH1YQN7fAd3kAgaSPt8V2NXhAnIyelekGK8A+3X0tPjd0SyJ
uB8yWjFz/MGNk8ohqMtW4XPUvrQtHbenyXxaSFCb5yK1uYupHmgXXfuH2zcNtA9uvwdIHr9V4Guj
kxTsTOeupoHSYvPE5wiwoyUyv7+TPpScZ37wB5RER43lPp83LQO34NNN6MXxsAQmeVz2HSVOyiGl
e2f4Rvp8IFfQK6vB1+61tBQB+zXBh8m2/rdgKexD1DDUQWnmHAqtfM8NmXoGjhGJsZW6MqSn559y
mGnbf3B3W4tm4gp5JKPjVlKBlg+7aINMvtI0nj/SGgBye7J5UGVUp0WdAk7DujsyoVwTIjs7ZPsC
Z31Iim/2js1iwkw07vlCXZ8RtohoVkLuj4SUy6PP1xLxn1uz7qbkqBpwZYhS9qql9y5LwzYDII9q
qmHyLhLhlyUJzpUyhT7irrwj+FlhWYmNXmeSTQ8ikK/qS8zI/galnug+Dkt5vV5GEH/GYPyMdO5c
cfdMBR99whuYyHEaVU7Y6Lh3cHqCH4tQBuOyrBDtpErx28C2a441cKNCrEjm+AeZWECr7hqzauBL
qpQXW1JrDTdjbE78CjVhjwJOzesnZnm5I5CFGisJslRrlPvhiNWCOr34lMv8+q1qvO46G/5aHJuO
TklKIVmvEqBhYQz1pHNfyYoDv3zliAnMdRr1yXHWmPz4uXLugxReDKUMaQhnFAmJLfJo9N5OQyY8
77jNoePZg2rx9QQg1FZ3bKFfw+62ZMiVwnXZiNfYZ38/FAsa7WFaowP50xRbpDpp0AB7k6SOTunK
sKo//mOSx5L6VNo7UqbOoHM+BLiXRY2gwDtm4fwMh1gk3yPH90kOO+4gf25naJTe3Do3TvN7214k
FIqHrdkUekMsw8EzH3YUD+QEwBnjJv4g1FVA7bmLzcSEAW6Up2ziRtaP+Eh3PLnDz3UVvPUBvutN
UT3bWoiarmU5qqcC4fnkveg0IOV6vrhEwzyJhXgpIxAWycRaZLrxbQSmw8aavg9yPRZCOaeDA9pb
CTMQjh+uFaHv8QSOJxcSSZ77VfKP4y+ei5DZplWb7Dhf0f1mVWvorTkM5sf8PW16L15M8HR4jwsd
JDGxyWKmsbe8fCLi2KosIzkhvCHkS6btBGp6QAGUSSJBnPx5uIjt/UgFsTaV5o4F5SsfcAhdV0t+
0RZdHB1fo6OTknKuVL4IsXJ9dSVLKcnG3EgQ7plMpyUXp00PJjlTTw5ITHHL2C4+WAM8X8wKdFmD
rUN29vgKkJNWQ2Yz/aVhU/htMNxIjCScx+CIvNObuPCoz5ohcpqsZIfY2uAbpVAU7W7z6yL1lbxo
bTuKYf+GQ7trlviOoXUDRD/HqoX6MVk7SEKEMCbG47HOTCcehMSwSJrwv+Wn8RDiKD0KErigoYcs
8pnuWGl4MkbTgJ+JvUzL1kcuxdufnxW71hKbtGyP107WeB5Odg3176iXjmudzEbp8Nvy5RS1ieEL
aOzgHDLqCK8JqZUiQswV8p7NokGqlczpwQR1CasnJaZWzUGNDhkTbwxxDAW2UUjDNlFAg4cHq1PY
hA8EL2Ha2ZSsRUuTGmKXhyx/QPyyPwzjjpa43KF3f+OFfG2gtXTLfdLr4dh4iVxnTne2Wb/mHqBo
15DHFQiBf766Qm3UdPaW+4TJYSCEE8SI27NXhcSb5ZadE6tijwqA6tQheHY+sS2CWCnV7KpvrAFM
DksISCX7lwe7y+BjkCsmCaf2hSYYUE4awqCPcMkKwUgYA6fgIfOxMWkgDov8Tk+77FpjeIR5BV53
E1KeHfO6O549eIdsS/T0wsXrTaQGywFbre4DQ7HmeP+MWRMBaVHATk30FyiayUMSzfgHcqVfFc/C
VdHnQpfh8Pm5tbjWgCCVzL8IHodVG3Cns0GIw6wBYCBZexxhqGSW+BVZWVLp+IXQbQHvyQbju/H0
J4RICOLNu4uBmboZU1bed3ClaM+Rc0++1O7rNBeZpT2QeaZ0wgenXm+SUhim0w8vE9dvFD0zNoTr
c9m/Ne5AATvPN1RSvv1EYndz0BtB4QMCSdn0EgS3fyxcdwedrEUKopifR0njW3fsJqJKIoy7a+bi
+vF+I3KnXpnkpDdeiDq/RIifnVHljcqoE1eK0jvpHsQsqrY2VwO+Xv2WA3hRmL4C6eEnq9Yd6NjY
L5XB46XB2Q9WH0o6OFDZt8HrvCfPiN0eRSoziOrnOj4YVKiWLwDVtxkvQEHDxrmpkd/+VslvY81l
5HKVd6X48TP6VrPPs1+/6qPJeIku+J/6w6UCDG0tx7/OMju6qVmSqheLfjHAvRpu1hk9anjTirMM
3cOjmPbU4XsyfjZ77YpwaGTnWexDO/VpdGPm5DUm1clNarN9AzBPN77LXz38NQD+LiNjTuEQlgc6
rPQxjYZqThHEOsOcui4zU633yxS8bTaW9TujKK2S95nSB7tXwfmqlx0pI2JTGxwkk2d8c+QF7xtf
lZhIBkhUymAV1McMnZgF0DwukehJkiR3YUqJH2LRiMhUKp4dO6jkURTtQLkcGnJhucXIhkB/7rFz
Vcz0b2vTk6hYMA6y/3Pa25MbYWSoeIrYhbMzSZFTaj+ILmPeOUl+mDrWBPTjqDBxdyP0rFHIywDc
N+XOLZ+XiUqycpxKlVqRbbwEYqa415EDDMdEUhAkkT7nJ6nRMyA2mnFN9fsrP50vQrXwrbKktTyD
1LhmxBhkPRVq/QkSRsiQcP+pqOHin9yf7sX8LzbhXbEYP3937th5y6P5JsgNROkFoVt2rItoXRtY
L7e9/jQv/gEp4sqgMkK1Eo3IjHkhwHUg9YjMUOSTlJPjsSenXziVLTKpr+laSKxPEZ+wMwrnwPw5
OPr9/r+FobC7l9SnqR5dtXplczhQ3ecVigMXoPJ2qWbA4sGL+XiDzxwAUlnLZVUsBPd8+ZUQ5omq
TepmFrdAgXQ/H7EgGuz0e8HCxkHS80tYy6tfsEpxf7DL30wRxg1XYnhgWQBkPFWNjw94nS7zr6iK
HOuhUTIgoCtAs8/GLkXkP17u/tY9sbJkkKPVKaz+NEn8JcXAYjUCQl9FbezMAhgHKpYsaQXcog71
2ni8NwqNtb3kOLgFu4lVJ89oJGhbUdDdSu8UYkPSyjWZmFba3ngqJYwf0gMotT272QLrx4u9CrVC
B6WY/id+IwJoCdvJo8oc04X9ysVYpGnUOZNzY1XTHgCdGq25zCgVOid7msqLf8cu0A51BQzxN/fh
PxWMJzoeTi7EOf+vPuYDjkQCqMx4ZHZQDD9HpVuZLARcDMdK6xLtP3xrItWgX2eeOxUxM6jWVfuS
4ZRugNk/ZAIcBlbq6VYNUUALFICnISikUAD52j/pzAK27y2aR0D7UnNfLPl6Zrem2Vs6GKJ2990K
yO9pxkIaJtyN3H81aNlsT7EKX6EDOhLDH63ccusqZq7pjJx0rZUCC29AzbXgdmew03VQkpVeBeOr
+LJBgJbkLDxwM0piBAOLM0RFgUNXABLMnRnSCaqLdYilaqfu3CDHh3euqscCA7tplYzt3InvWpYe
g3oWriC6UDldn0iWpRxcORNBk92UaM09eJ96IyxkAl4KnPOFbwzbnYla+w6QorMCFBIwbrYALhPz
gpQ3nGr4vRJORO/SW0wLF9aVg1b5ZVXWCEJ8GvhJkKcVYvyYI+x/JOuyCw7lAH5lyIGY3Q7mfJtK
vAbgehz9ZNTdlhkjc/IKnneqnRIy15LEHq105zx9bWTmNpTcKyOrrtOfES/0iYZIN0C4dcPoQf8o
U4+0FM2f7psWOcqGeUavvY2ZoG5n/zKlCW9NdIl80Qwz72duhVlxa1rEgv5OjZucNF9HcrKDjZwI
C4NVF0ueMnVwxX0Y+AunKzG3iDQbmcKzjUgnXNhSCIOROZaLSYCz+3GWTsvBzXz6eR25hel8fJJR
b3zLHtQLrjxNAYwJFjI3b/52AUUTQoJuNmeFLX/rFUThofRqwsVQLHxmmEmCiJVwX2gaX1yydMIL
F8HFHByqfIA22RikhhzZvR9goDQ1rkn2DHOo+JtQefyZBYIORQQuRUXRr9O4B2ZVQ2VeVbq4nteR
F1aJ/KRzOgVGRzgf8snMZDixfo80VSorwyKj8yhkStekmGaILD0vsxU6QHI8JIznS3ckUcqcAMge
GKSLJtFZcQ/N021oa7LAas5ElqAVGMCjQBMf2uygMg4JhxX+6CUOWcgS1iSeEVE+TY6uKMYBE5MC
P55OunbEJFjguCM/jpMyWpd509LOTqz0+xjTwkCB2Okg3JF/hlq8Oywm7ilpWWVbpXx56LBV91/X
U+CiIS3eakj3L/gRFDCZCZw56wbTwY3RyfuuumjMw7UeSp+b6f80w3BnhLKQlyKLdX0J89MO+AS8
3SJh7AIhWnbHX+7cQjKpjhSXmolkTZa9QqpHjaJ1tnzyXAesk2d/kTHLqPlhwq1pugNawVW4yVpb
jqlbgm3XySIwSTyXy4RE9slVqewqsGe/24abBSc80+Tt7RTw8NF2ZSup25asMnMVHbYoC5JtjLf5
x/BOsuyOlgyH9WDpBwV0ASDqmmCD6bTVQXOD3Io4l1zO/VRRX/NQSFsJIbaA0TQTRKRZ17wIfyXW
rlx68HQEvhiYh8EPWRLtBUlYKsmBFjdbDzyXLc60/6hUa3atTFX0amjN0c5Z6AgGQWP/h2Ur9Rzb
gMnoL2DvdZWhE8nj4Mw5B878g77wAmNG+l2n/5oe8SbNkM1vFUVIltxH5ciyMol/mij+sXsOSvsD
5YPoZ1u7GtsRiP6Co4/wI3FpK3eGEEYKB+Jq2zP8jZEHM5cMvPnBb6nsoB8HayPRHv9BjNCa4tar
Ge4fmsCu1AX4htRYlvVQ/P0NfqiBKVBMhmCd7eDTXlfKl0m/wZ1EbiQXe1XkgKTetZtM+0x7YQ2u
32eIO4N6A1ZvfUsF66PMUAnXb6lY6G15sM/aRGM/pRkB3RpTQfruXlDlDNHTkLfuvPt8izUnEBpC
wvNOvDKN4iXTWClXnSVU7u1CkLcNtSBDVdU3027iUWYBzG1NM3LiMQGD5WmiraUXST3b7xkyf0mD
uPTfmB/+nPwLEkem+FY2WLr5pjqCJWN07hXu5tlSBSWD3BwIBZvTZsSTdLWLSbkiayW3ypjlN8gV
FTUYZbYDA+Gxng9z9n7eytXhFHunaUYuxhLW8fLD1l5bFv2/oWYz57Cr77ivNgxakybPhTF8zKc4
RfkkgXgNea3WSJab4GQsTHFKci36J0oD7Zh/t1rjXaMrPhH/k5+RZHLO0973CmMbtaHMaPmuKfT5
+isF/5rWojqCzJ3+bKqf1iWlJHXgLUhkp3jDI/8k/Rl1e0KJF4dziOIx6ecUgLLsjnTEWggmcJTz
dF3eYVKJrGlY7t5vMBPKn+apFZBcmBHFK6Bm2OYpn96igHX+/hPGPfy/yU3IZcG2ZUlSi9OY/QWo
amj37stA6XJYdNcHqoo96fJPPcpH0iPKGniXEogCvzAF1dMx3LjAFopFXSCGTp/XBHuFm916aklK
rYzyEcHy/R8+kEN9IYWij3dJOybK8xI2YWx5EbIlhohrITr1yuapwMNh54Kte77TBKreEuxVl0fB
2BdoBiZckSp6FVJ8sqsunsW7ouZBTlborB0mjbMCrwNK7/WhJcjhOQmVRGhlOsOzZ/DtKGZFvd7z
nOu71hqfqsQs6p71a997L9cq+boaD3Uu4n4aY7ZmhZRfBgUqHRwj3zX3Bk96vxU3LGGTVhVu4FAn
yMN/K84yxjT+SZE1m0q9WkQa0IHlwlSpznrh/oY8ZAVzXUx3GgQg0FBKL6TKCG7Pj/Hs6qlT/lYx
SlVbJuWq3wVFhC80fLchgQkBuJkrxu4Y/czYpQtYCL3953fOSaNaBWkEFip+wKccNysFLwGGY0BE
JdI+UXXmIUn9IMw/69hok6rD7TaOaTP43b09yUNQ7rIzurbGD80KjJUj85tUt8NYX7fM0h2hNqYn
Kcpd7V9L9g6TtgN+8GbYf57MZ5qcWWJjr/K9AQucpDA6/ODneEgIs4W+hCSG3XEa265p5WrG9gnD
nuv3pyHr2rsXpItWticQsuHdQ2QMfWiC+6ZaoirmHfgmwN5EZpqqtlLUNF8Ss476zta03l+s26ve
gkBas3nEyDwIVGQepvbNh6JxhSz54HDN18fi3iB+LvXK2ci23kwyg2I9ZBZLVSVovR+SXR0m2Jfu
efL/nhAxxFappYijy+UkEPfY5ZqVBSyeKO9cXslB4RdGuWw3AyJHjMe0lWsSfQid6o/ONgWyzHJj
mGLczlzr65HxuwC2kYurnwNWZAU8g0JpSgDUYaZkAeJ2OY9W8AW1EvYKk/0VVfye1ARAMIadoqBF
M2mHJPid4opnJiiEVKT7pqTkKhnFfYssaW7I7JaNqVcThiUDgJyIjytMx5SYNN2QdLNTsr9vbGqT
XtEx1s7hNxcRAvLuf/GyTi8yO+sURHielpZf45d5SaQiBOAQyxmxjgNe1tXiXNQr/y5lJQyvjwqb
I8C5dVkSMuRqsahk8Q8WNXJFwHtJ7joyGM5PCBuIVSo/0nP+HDYuuLbP+08kOIM5nS4jWV77k3bG
j5H4gsNukvudman6VA973ze75SN/ecaMFzEKk1aK4Px8QDGldZXmOqY9EBJsH2D55FUz886pALp2
s2j+HqMualA5zvIfEe4zDF42hoNCTpSROB7QoEVWWU6OvvMEyZM8GoEaf0oMHAzNsJ+6gMGDvkKD
uYqUymdQLe0bcCOcOFB8xtXc0w69+LD8cbMz89j7J7lxvDprh5ftF9Nfp8W9kfl6v893UHnwe33z
759WjPrnnmOXWKPck0jVOncGWRB/pUNtIKTuVPmbZGs+ds7zN7aACGm0u9DF6169Ugit5JtKTu3A
0cBCgogtU0YysyS0Pm6i2FzJYihD4LGnmH7JQKWYVtdIdnLfhzyJ0wv4LkrCv2aofu/dBcKI4+dg
aRnUfIMSzn56m+wVRRpm4YrMHV2u2PzTXk3R6+a/87ET9G+dM8Sk6XM0j70bv2y5q+JI7Xoa9lve
aij+skXsaosfLgHg2xTdzS94+/cV8dROIxDLd1WzdlZP9ZzCwl5Z2U1SQpM0vHxrEqlBf/DN6hvq
+uc1haAq/bXqc7F5axmIBZFxRETBKdLcUZ1VjiVZe8iBInn2QvOVHbeGSvCiebndbahowHJrneaG
pl2daZT3NTtRP9tyNoYjufsLlPPqpHijEf6/HMUygxcLs49vBdXwz52MtmcW8STTjXdaWsUVCDST
4OO6rX7o8NlpPfsdWbEDwCzSIhKB7kgzddgwNoHQbzjrh8JCYy9rqE9JWlzApUVxDcEXhz5U2y6L
EjKC0zisbC3habtQXyCPhVK3xNPQQaZFwzs8XCntF+OzBIyRd9K/g3dI/r9DlV7hPFrcIqKEOLOH
lHhPNoIn6Ft3cuEDIr1UQ4uE6Rm9Ppaqn0FJynON5TeK9vRkEH9x4UawTHRpdWMbo0mSe4ZnNnsn
MZO+i6RB8UxjcBrVt8tabHdZfrxVx3oHGd+m+C0bhVx0b1HudZh8t+Y6aEFbOCds2x9hA69DD+d4
Z9FcjfvzgeVDqxb5Rr5cOkNF4o1w1v+4bbirylJQE3to/y6qEfkN30+sVxdelSKC/FszQR/9Cyd9
P4xiSWOq4rgPCeWDf6Oa41nE7xmumXcA9zs7lzsm6LtDpeUf1ZTB2CowPc5cQo83MAYubXVcsGia
5blOYM01ii5S9ArMl1XmABrvU9e4jGBR/SfGpxOGHIrt9ewMi9tVpz9vbHAZGgS2ncx8LPgp4NuL
mqz9mMTQaRQG0WuaeS3D4s/mnXjudomCV6dazH+Kmmt7cLOS3GFVhvnEXCS3duK4wdWW1CP6CPnZ
Oqa9DgiuPwA4fT+ivESCAS1ZzKL34gu0Vzx7sqQTlIMYBmnoVPZcQMykCEols1seE4z0+W7FzOL1
VqrutZe8TbBHwRAk1waVQPUVYmPYYbj7769yXaPsmbtDCeSMOls9VJeP8BKv6+OHiLZ3n0hXgDKK
Xww7eq58ZGynQs56Ht5Rcr36FbImymUPtBI4WqW/zEJXft1opubRr15UGpOncfi0LLHVcM9IYsbA
UcDmgiP5G3nyaLbdhDzWWHBG5S3ySC6dDD5AK/rRzzFEjJ9sT/BEXmTQ8QhPOnS8x1vdEF30Dlrv
n6MWW+hdnlNEWHBdnxTF+K5gOicj7i9AIS4n19fkwP6CL5rKeRyik5DcXfPn0IvB6JpieW3Oidbd
8ZLFfZVVksVwQGdIY7wrXAOYB/9tlfcyXOxZAEsUxiOS0jR4w83TxlRf+74A9qJtSYq14j4wWpwD
qiWpHMx4yKxb15miRWL3uBukL4r+O2xuVgbKzZwCIIW7zS5TmqexPXaX7bsqFhGT1cfKu263Vm80
ef19P1Aac8ISA+pHJ3xqN1GTHRqKkB1RVFIsnEzSDUGXToZIKoSgIJlWU54KFTf6HpGzfCLnbR3t
hyTCTwo39XpV0tModDBcxC67Fp0BCIRT3QLSP9tntWAhvLDIuMNKuaDM5Dw7FfxJ6A8KudWEx65i
OCorJL9I56+pNDrJ8pii4jdTBqTNI4YW2kMK5VR+jwUXu09fYcxAf/IdgAQRcCpcJGcKJZx/cv7o
BNvct5jCKVr2T9F606ZSftsFDmIRfSPSj6pVzhfXaq3SBxtrGnEaADUuvr4oJgD2b1hQAwPyWG0o
WKBOATqt0ZmNIi1iTHbRa6MKNKvduX4b4v3oar9TnF+jJoAF9K2isUVbiVFPWozVht2NmxuF1BXe
ERBePaX2WezOck1oEqsrBs7oDCPohPo0U1nmDumBJAG8h2ljd8IOF48YXjYK58O6gU9CAXubSIBE
ckaAoK+EI4w9QwLPS/dyX2Lfcpu/j7Opu6DC1f8wpJPlYbA/Dc4jE3lukhxkQM9alMctzPKoE+PK
diuaN63mYK3oYvZgTYq6S8+qLcGxq97EJW1S7zB/giC0c1jbz4ZiYpS5TKuqnbOKR/1vOOK8duSm
DvZp2/RtuIh1rmNgUauxvMNLt8T44SkDClZAMZ/1PTYgTnVsxq760kJKX2ySMvWiWLAmxU1MYbVe
4Zz/fbO//updGNk5JIeedOO7hZGYIEDA/Q0/tDsYV8f8scau55bjBig19A4ZGBOC4W/6R70lysge
2iLZ26EDPN+RWCfw/f4xZ1Hu5F4XAQoe9johiqHcbrJhtRuLX3fXWWQLrl7k/wrL9tiGRaINB31C
qCnBgw+euwTO7TDBlO8PBP8pTNR5z07HLqhUngoTKLW/B7SFSj1qDKLZqZca1qqthNJt0eGA3RmQ
cPskJikWcqMHUb3cN54nUZexh88mpF/x5/TXEJmWZCf/jdUksZGOrZmRU619IOZ7rtbrBX7L6+Qo
g8uFk0HqH3ZN+jIUBgmNk+zvoyiI1MX9EUEVOkooldrIaf3eJ+KqnhV+2RPsIwKsdcnNN5MYTa41
tGOmttqIR/q6MfvN/31z7+vldsmdgdSQqhjBAZYK7wqAM2dQNKNjcgGQorJrPo1EFGU5Ee8rJhGB
AfNujfo+YJ7DZVn0lCHFUhoA9E5FymkbzGC1p3c7XO0gw8yCWMpuPSBJmNU7ZnAlNF0s4oCrPpKp
P5KJ8j/kYYz05wG4+dnCh0RDgAYvwGzt6C/RidpIMLcji1dgKKH7OU5um0DqKmWjTzRcLhPN+R4C
PBS3koZrL9cMkLDgORdEmbiueOTTJWQDQJpGjVB/JSk9PyI884TL8gqnOoMbbFiY9KhieBOHWkgy
Lns2izQ1TLIb3GsLOASjLMSSZ8u8eqc7G1nBfuztYVT1iBUZr5wCXmZF5oILA9MsoGyYXG4wSh5c
HuXReuA/RaBfbqHFAJvIRt3Awh2ksL4QMhFqOA2A77jxhLE64QoL7i0vTXt4VF3sA95d8uq120fK
Ve1sb8l0Xuv7OYF6hw+m661lGCGhslqGRthObiTraUJ0QhWI82wDEDo7B0Nwu9ueoQOQREVDgur3
fjTd1d7Xjw0KMzkD4XM7hmwDB2cvJtPBncz36JqLCTOM3k7Z6FyShctgLuBkqvlNzsQeTw4VCbvV
5EGgHEMWlGuhSSUVwezStLkkmjcUGZYGZF8ZyyvVcL1vjR8T+3Wh8sGaudmh/ZcJoHWluFG5v+d3
2YpuJOoZ/9YKadhxxjCWzHkiTB0JKE1DlRxJOa2t9FsA1jtvNYO5510J30I5/3gmxjw2e/F49JM8
r6K1rXfHaDnKi1kfSqivbFwmiaVg5dqeH9RM7bdjC7iKxwoLqt+c+CkBxFFWVQNxw6EBVXbKBQ3m
1LY4gFQfs2IPfdLuCkPePW2e9q3c/ne9Jtckt3cYeSHP2/pJ3K9b6OCmHMtEufN85NbjENDQJwBq
kcdFruBjb+i2hMBN+jT3xK1nFcSWkuwedeq/TX2JmTJKMPx78iER/KfpLPHWbUBwO/5mbixfk/lO
wnQw70kD2Y24dJzz1N0IrXZGEotysppBY1cQQRXB6XVqHrYTA3dA2MJ48DK9wH63rWr1dT5uMB+h
JM6pdvAMr2FCF9Js8fSUutxlA03rtL0bE2xuriQpOI7dPomazUlEqi47KQ2UUrXMvgXxNC9hpf7k
lqLuNrVw0SjnkAuZfM9ndjJREVI/HEs3M53xYiZNaAKCp/BLeyqBqnVA0vzndjLdjbLWSE2zgaCe
BrZRxSL60aMLwN2PpQ6R5QtyTww0lg9NaKshC/xFJlJjsh+Jg3UJgqOSICEM98VufR0DPmvr3ifI
KG+fPR23HWvLowJ1TZhgFPVnfsevQKEW/eN82EEb6b9q85+2OjfICk217jfMAN4xljJ0Fy52iuTz
Hbua42c2gCaEwHFbXzh5SRPXXYq0mtsNus55mQ5wHAPskUbmjOt4IaHrsDoZRiNb00iu/OuNohui
wbnCM2GDN9pP/LWZKDb+fSklNCRVSoaiuRpOHBPo3ahZ/gAuF9FqaRWlfYNGraDZoNqidoqsNXsJ
mqLJIQaCm/3efctP5VhBGfnvLvLzd0+0tbX19lRhtR6CfvpUJ1JBEpRTJl1z5qTT29sDLWLCjCRk
DYDLEnpRQ2CCfuI8xrS6ZwfoEXxkXWYmS+HMWS66rgIt36VSPKwhOTh7ZfKx7fEDlBBLywN166Fw
/s85rf40xtenEitKfBkoIJrTlhbN4KwP27Zij8pK4q4=
`protect end_protected
