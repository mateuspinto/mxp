XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%l��@��jv���eٹe��3�a8�ߡ�5��pq��)�4
b`���"���� ,�<X���Cv>�E0�ut=� ��HG`�dl3E�N�C�?�/�.�8��O��l(Ҭ�u=���1�"?�2ZR[4�j�ۼ�����TD���`�	n��O��4�>�����=���{t�'rH7�Lޟ�E����Q.� �M�_%��.� 4��9J_�E���ɇ%
�|�mOV-0�������9�<��k�θ.�=��i��ȫ��k���]BC����d݆j�!]�K�Y#�4�z@ǵ�D�A�z�P}&�Xx�d�̼,7�Azw��"��-ڒw7_|7�r���W�i�]�n���H9���׸X�H�3���&$e��-�}��v��@x�6��G�qAU�$��iϏ�A��d�� aY�o�>��������h�T8'��-ԃ����F�D$�Tx=�o!�����%��K��8��HmԷ�vk:u�{�|�kg�4�f�'4b&8������n�L��^&���k0��u�����F�(ńuQEs6�wcBꁍ��<�x���{c������ħ�[�S{��RPn���a�,9�*.�3�9I:[ٹ�e8���g� b�������.�!�����_�~f$�duJ���8G�k.E�:��K���|yP���
�v����n}C��0���.@A?m� ށ�n-���.�qo��Ynt��x���h�E/��XlxVHYEB     400     180*�voޔP��P8���k`� ���DU��H�{o>'-�!��,˨񇕾'+�Ԑ����w�BF�Z�y�|���[`5���./��4"m]���0���ul
3��mh�!푇�zRRe�k�f�W(���E�X�?���A����d����i�b�w�	��:�-��sE�j�/�Щ?8�T��Ι-�}Z,�$u�df�xq�n�UGbP�t��hOP>���q�?����\8�VԢ���ށ�4a�#�ߗ�u3X���-�/�n[�"��V�q���6I��&�?\C�{I�G4��~)dI�tDm<��A�X=�gf���s,�"����V@�cȪ�+o�6}!�ۆcg� 0W��h����D�갛3����tm���XXlxVHYEB     400     160NL�z@��o>�Z�xi��N2��Z�]��hOË �b�����`�X�� �}���1~���;f�����
�`Y����~�^�4��^��}�g!�̂���;W�����ޡ+����fڞi9��}����ɶp�&)�f���M�����Y�ѕV��N�?r�$���p��b�!n#�d�:)�~�"Z3�v6�b�k����Vv�����+#oPja�K��C&�+v��jzj u
���V�%�H�P�ˈ7(Ң����E�~ی���v��Dx��٦HB�a�d�w�E��C]��m��۪�HX\}x��B�����8O?g>���M��'�ry�K*+\6��:�XlxVHYEB     400      a0�QNH��4%S���
�B_q�E�no��^y����{��=2�%�jX"�f&x�G]E��1���9�L�С?֟d��ϓ�D{i����F��-N��lĕ����>�o] ��m�3�ߘn1h��z��$���Bj����s��N��y+4���u��v��6XlxVHYEB     400     120� S��"�����)	�1�+�5��*x�f���
f�`W{5��@��)�R�M�7t��?�h�s��ԣ�[�Ӂ��䰅;�X�Z��Qy�5?�b�i�N��d��t��������L{����"go�i��EE�{'�g[��1�)"L�"��S�jRJ;���9a�'>UR�B�@P]�0a�A���<�^�A��RW�߳�:l#з�������p5��|b���r�ק#�w�*�y�r-�;���C��1}�;)%U/�Ә�L� �7M/���M�|`XlxVHYEB     400     110����7@GϺ��_��p�:��#����m�����K}�v�I�����w$Ӌ�>I���8�W�~���T���*��UcT���,�P{ b�6�Ֆ��l�`��<��z���ts$z&_!��nI9�91�@�
.�7�F��\L�g0g��pu2]|_�+xK�N��/����)�i����øj��mD���׵��h'Y �VBvܗƀX*���-l�Tn����{�@���v�˞<kQc�y~���>A��KMmv��[���XlxVHYEB     400     130yOM�ἁB��sIJe�b�� �F*�֯:���nD�Z�JA��	�9mx1�0{a(g�����e�/��6�aԌ�_��-��G;p���pݘ�D�N��ı��_i$T����˕��}d�f�u�Ad�?|C,�	�ѰJ�'ޗ�P�����,3?�������o{<��JM��Q!f�mQ��J��!¥Bo�`��Vz�|�En����\B�!Q\YG�{�&@��ؿA�+M�_�C�2�)�6^/Sd[Q<aT��v{0{}TF1H/��XTJ�*���#]�H������;�Rt.�zZ7ҁXlxVHYEB     400     130���Na�)�_�]V���B��U�=`�Xy�M�x�1N�������e�nK�"�DL�@�mD5�v�V��.�X5c^ ��"�WK�����i	��C�$����~ j�6��ú���|hA�g�Rj;zx�� H��z�5$G���懽ڄ-��UIx�a ��N�<`c�;��ӂu��B��_��iuB�LN���>pl�_c�qm�J��g���4B:����Fy�2�lu>�+֞��n��� ��y�3a~i'Wd=FJi�Rc�� ��qw������̯	C���XlxVHYEB     400     120�b��"%�$ s��#�V����c4�쬏�r�OK7*O��(q����B�(p�}�U�*��[5��1ڒ�7w=������{NM�o�[
���( �G�#���cW^�b։��"�\�OIח��^������J=Y*�Z�(]�Is����e��T(YK�m��l�T����46���X��E1x^J=T�������9� 0Yؿ�xx'�n63ȑH�k��%�s��^-]G�����t�p��_
�x:ֺe�}��O��2H9�no��]h�޻U�`�jz�;��XlxVHYEB     3a6     180������܇�� ��;�Ю��DYI�V��Y`}Q��YVr�u!���z�,rYo.�}�;����&6�P��w�'�N�<<�E*����������m4:�X.b���.�4��Y�q����w>��<A
Ϊ��*��|�_NA���m�t	�|�I�Y��R�׷1q��9}&�l�A�=�B��N��R���ϙEٓ��-�$�����gM/���t��wǆ5����1���t�q����GB�,���nuS�G���7_�]r�P�J�G�,�(�����{1��HF����*�"�Q�J��g��I����)0Or��Hp_е<�u?���<���Fq��gzI;|?�܉��a9����XZ3d��ϱ���X���c���