XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����V(�a����DwS��6��x�ٕ�S����K[i�l�
Fj�Wah��}��ns.zg����dy�k­G!6�E�&�~�b�C����)���|$�8 t���	�kB�4������L6�^�d�DVf��ܘhTP���0���grA�=�k����$t����o����j�-'з�sT�,�;R����	�#Y�C�A߳�������$�T�)��&SZ��a���P�;ι0T'�GfKn�8�O�yIQ߳���H2�~ڶP�FeG0�o�:W�YVd�2��Y�Q���_Cy��S &'��2�}�T��EQ��K�}���%Sf83V��_0�&�;�������`��y!�ONw�� M��y�.�^C2�+%׺�������S廎N>_-|�k=F��P�UVz�Q��Z@���կ�x��_`��p���B
0��iG^��D2O]N�6p�u�r2zS' ��G�7t�̒?�js�g�j�հĿ�����n>N�~�{���~�-�C�#�ȃ�<����ʒ�P�Ҵ<�]�	���ydf��]�m!�@7�g
2~��#��j�5]�x���=����.�K���K9�U��O�QQ#'~����n�P��,�ڰe���V����_,ri�8�k)�?d����-�ػI��m�F�X�Z����=�l�rb�T����$��OO3QXyx`���7s����8��T�xō���R¬�z`�x��'S�)"�a{���*VM�l��A���)2�K�XlxVHYEB     400     230���K�~�ƻ���(�nPO�d �CK�"�8���b�ۥ������3����	��g'��"���ݕ�z'�R�5u��*��	Ha�ɥ��1[������ԩ�%P��b� &��lXvH�4��v{�)�q3�`�Y~���c��X@��>����r��Z:Q4p-�9�G�h͸��x��N0�wGl��ӛ�
Z~=��\���N����K��b�%���̡��r��UɾC���tԌ�DP��S���]���� ��#����
s\F.A\��q�otV'Xh�,���������a#���^#Å��%��rK��q0�ƴ�*|� F���R���9��N��U������B��42g�,}U�b�Aݞ�0>�B�1��2Tr����n���/�t��!ɚ� �Jg�N�z�oui1%[w�/����M���=��d"Q��l7��W!���ܦ����>#��2��f�O>����
x���q��5}�m��W7��կ�� �qA�'��~���v�#!�đv0Z��tPm��r�<���:�mXlxVHYEB     400     1f0��ԣE��J�,���xLK��A��T���[��\\���8�k��IN�T��2�L*.�b��!	�X2�m62��6����2+#����@ݘ��&@�B<Hjg>��0��a��Y��;�qi���9>�2:�ɓ��4�*m�3��W�!����'῾�߹���3��F����)q��4[�Y�Q9Hk��䱀��|�S��!�qAd�4�gG8�QӃ��M��M�m�Q��]�����M��D��hb.ܽ���¶�� QF$����`-]��4�����e�i���[ÅШtܲ"��/y+m��+����0~�J)����~�d�T#�5�����ot��R���Ql|�N��I��=�mVO�����$�p��6�����0uT/��5l�R��X�f���"ꅔ��,��n�B#�<vY	�bA���~��n!捗��
s"�w��i��\����X���J���I>XlxVHYEB     400     1b0�>{��5��֖�,�=����c+J�h�y���h�'f�*0DW~�;�h�I��	��@��F�Һ/�a�w�=�jjEh6%��<s9a[T��ƽ�{5s
"�[��aZp�r�R@�2�;h�:�����,c]
V��+���[ߴv�s�R��Au��7�
��ؾO�7Ry�d�+\v�A��ά��D$:��S��?ɤ���m!˦N_�'Y=:a�HF�x��rm��_u��!XO��
5�Υ��sS�Y>�ϫPE�`�	�[S��ńh�T!
����Hr��8l��[���.*�qOH�O��g������`"7�鹁!������Q����ݭ2kl�[�B��L���)�9����cVh�D�:�0��|�(����C�}���Yg2-@��(=Q�{��Ⳑ��α ���0>[�Ҧ �;���΂��XlxVHYEB     186      b0��������b%�":�G]&Ӈ��i�f�I��+V"�j�ӂ�X�eR���V:�;܊���d>��f�(7������<Bb��D栳����@��!����XB"m�|��gN�yu��#��(�9
09
���PtލdI"�}Rz��5҅G4v�J�@�v�`X�{����R�pT�#*2