XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4��a]�4^����j�OP����ʣ�گ|���,����lӵ�������Jx�{t*5��ou�d���i}�q��s,�����V��z3����T&<��0�5I*�����r-w	f�f:�kOE� �i�)����W�s\�$���a�R����Q&_��y�q��0�G��YeZ�q3*�0�ݐ�@���U̓�K'E��� /�B?���7���xHM���Z���c�Z��(!޲�F����
&�\-���@G�jhˑ	��Pܤ1"���8�1�D�/|�FL����p�ʭ?�E��Š�0p��A�{�\���Ӻ��9�<#��ӻԑ��6>��4���ů�g
�
�d�ޒ@�����@߿B��%��	�|�n�u��C>b���[��a0���D5�������y��@:����K�&���D%ENZ��ŋ�Ė��<ݕ1�%t�5f��?����R�����a;�� P�D������b[��w+a�9U�����z*Aا|C�]�<ݬ�lҞQH�XB�<�0�}:�KE2��O�`��sS�O�W��M�4����`k������!��[�+�e�h˶�rd� ^�j��(���t�մ%��?�ye������k�-����]F�ڙ��" "��N}����<o���+sq���'��0�q�2;!�Jeh�m���^�{!P/}�7A'!ro��&�y����H �zgP�O1 ���WS$b�3�M���1I|XlxVHYEB     400     190X���ХPx�u�q��.���k����2��
�A:�\�4/�i�r�n;��R΂>�u�o�9	5(�u�<	-��[���-���<�$���A_��J�X�<ǳy,\����iG�ax�����S����>K��7�3�UH�/�w5��\��2���=|#����@�4�Q������ �|Bm�{���2M���l+:�L���៴1��	�W	c?k��/S�$Յ*���S
^�s�%#9"���U�\s`�����<0<*�/���?������Jx��E�B�H�/꿷< ,�O�t�Kdщh�'��V�OC!�ձ�5�*@c��Ma1�.�\�΢Zc�Э�g<�"�s�`��	�c7$m��֕Ѣ����3u�XlxVHYEB     400      b0)=��]�O)����21��/�W��(���!Ǳ���N���S�(��U��w*7C�q�'�2�!�,Ny�M�ܟ����i�
�&�V�6΂zd��˗���uJ��OjF[2/L�9ӮS󲷱B,i"a��k8/�6�dgi���c�Z��a4<����ש�	��ԅ5���XlxVHYEB     400      f0��Ϫ�,�uy:����(m�L���a^~ϕ�V��I���� .��1�z�"K2�:�1���+zA��������}Ke��V�⬒�}/�z��gx�+"��l@��)��o���$�	��X���/F�t�Zzj��<ߨg��'Яw,�{�}1���,s}[#`�Ka�mʿ/�0�b�q�m�KH�Az����4w/"h�)1ON��eZ���0��+��YS�vK%9ϯ/XlxVHYEB     400     150�=�z(pY3]Y��5�d~�#p���gzW"R�l�� j~�T$�%0��$j�칕_�[p�����zӧ�Ot�`�X$|[�Q:��V��M�[�I80T�g@P*Rę���5��B(��|ygH��3�y	gPM<-N��Y\W����R��:�����J����K ե����\M1�໗�Z�+X5cd�F���cF��i ���Q%�g�J��4|[���O��v�DL�c K�T��~�)8�2m?9\vXl��{߄��1|�O������<yk���||�+�#v�J������m'�](jDf���2xD�p�:[&7��u�tf�Q�$"c:�<l�XlxVHYEB     400     160���Dd1MGKu�q�O�����֮�Yz���+�d)��y��ޙJ#�&�I(�����*�E{�3˛�.�����4�k���B�� Q�А��6D�ev�J�v{Z|U�\䈋�q��>��G�L�~>
+WzjA���rg�H����PPuW	f'˷���#�͓�f�J�����8UE�)1A�L��ax��䛓��g��-�il�q4����)t�4�lH���������ǙL�D�U�*Yl\�zzRS�����1��`v�ys5hj�Y�TM�!A^`8�����KӛQ��O�ZiQx��a<�����,�:PY��<�i��Q�M�����B��XlxVHYEB     400     120�}5<ӧ1 ���]\I�h�*osW£��0pe9J�Ǆ�İ������#V[��w%ˉ5�y:`�>v�.J.�1��~!���-�� �Y�\2�|өޚF'� V��{<���2i%��A�s�K+%��D�����q i�
��v AL����%t��[Ο��͓�fWs���v_����A��%<��o� b@����,���{�i���s��=�t����oư����D�i�?�1Ta*!�;�^�Uk*MX��"�d���jeu$&��#��9E����JXlxVHYEB     400     110�Ϻ�������H�?$iSs}�����G�*E�v� �����:�q{ti�Ņu�|d��n�U��B�� C�U���?���C�׹<����=w�w'��M�/�y������'դ�FX�o�ֱ�_�tT��;�aq=_JZsIb�M�5�A{R�.g{����ʣ�������1EH�I@�d�]��(����D:"Ă����k�)��[��9��3��lڀ7���^F�Vqa��W��۷��}H�� �˹P�ѡ�GA�������׼k�n_$XlxVHYEB     400     110�?A���P�aTs�P6!�k�7��W]W9
أcu'R�D�B,�r�EM��ɩզ�_�E���@�^�@,�1�����(��M�bkk�M�fkN�Y�������g�������N��	)`��Sc�3S� A��kT/��+��6��]+`��k����)<��:6�/���U$&��bP����)�{`�|Ƣ\�,Z��bHy�*q����Y�q�=��	
M��K]��.�b�L��T]:�e
ܠt
�����*�XlxVHYEB     400     130�b��72=��>n��l��t;xh{�ؽ�;��~!�{J�<&��l������Hf3�X-�"��rf|��͇xRm�5��d�\ip(��ԓ�~]kq��	�x��WhW�XN�R�#�vؙ� 	.=�6I�Eά��=e�cCf��I*����p���T����1����U�����z3��Vk� �5Q���}M�ˑ���'���D\,�?n�z. ���λ�f��A�>,k���篣�]����̐�
l�%WK��S�#V��l�sė?�3��*wc�!*w�8қ��f�.:=��XlxVHYEB     400     140
��ejpL}�I?c���g(.z�4Vf�Tk���4N�9�՚��{�yXe\�[��I�^�2�+��F"5m�E��M�������0�c���ÆȆ��zf'o���p�{�i0���34�0;���?�{O�c��x��[Ȇr���5�Dˎ����Rک�%����Ω��)�����Ha���zl�Ֆ��2:���C��N)�c�za�OfEW��!����G�a�.:�q���Қ��S�u�k�ћ��QeM����õ&ٶ�7xjEl�����1�ax���,z��謁ץ;�!"|�z̟�8�pXlxVHYEB     400     100͓~����z�08H�8�ݿ���-�R8�TpX.�Af��&N�=+ͫ�����$p��%C�������� ��,*���SHe±�R�����N�p[�MK�2�(H�%.(���[���oˌ�%�9E���#+T3�=?S��%������kWl�D�/�Xlr8�6����~H�,�]����	FY\�W�a{V���i^v���Ab[�w<$2��%�[p Eb	�%2���;���$Hu v��}�XlxVHYEB     37b     140���Nծ�V��)EQW磼WA}N|�O���NL�jO7��q��-J�@��J��S�g��V���~��������J�J�6��.`�K��87=C�"��gdt����u�/DU����9M��� �{�?%C�,��vn��sR��[s;7��.Ozo���J�Qk���nN�"j���7=��D�F?�XP<)5}�0N�hB��F��{��Շb�M�Pk�ɯ�ET��ӈ��#%3!�
�&�c,��``�Z}br�"�ө�>�e���)t7�+����cmA��$�����a\��/�![{;K�@