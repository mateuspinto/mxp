`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
NzJPAaa648jC4SrqFtY074/cmM1mxZlXrL96sgVeeWWlj1ge8zvBSkil8enADxNhaZQ4gzCxgXT3
cwoVlBNE6TRhu92LEpqpwRd9cEOPNsUn+TuySZX6Xg1oC2Sy24ho3tvY8fmf1gsPs3GVV+ghyIKN
FIFaHUctlUE6n4tnKOlKK4ILg1WK3Qz1UYfrUdsNaxmAMiDqyKLzJy2XEWSBGOlwdI22yY/V+fGz
t3iMmehbS/Pk2yG7vjUrQE7fuS43bgZTpBfy1iguwOovorgpF6ORFQCCfs7WMeShzHtyDILrRf8v
KkXjvUns/RTqQT+29AuJ8/jHNVzZGb7mUn4wdZuKZQqu6aVI2gehL6tgDNBLQflyBhd9e+i2G5Dw
yFP7pvBjR32mQQXFgRn8Jvd+TCCWU1wnbkXQUpQMbPBOHaNaYQrl40g3Co+oiEXRPY/91UnpBSml
NPh0O8vWBr4SMy1HmXYfmnNziI6k3/PaD9SnN/UK/pAJgTGZROqYppNB9h9RI4DKRDfwrwSBPMTS
Lh8y4S9vewITJ9gduMHSC45XLTjakEnhgON7ynuysb1g6sh81gxSwzC/Fp5noJS2C1xiZYBpM+2Y
PIyEGaH9ifBGUyC0dq9DCaWN0lhiWwpAiE1S5MlGdfER6eWWVnm6ccVBByCWf8XILHvzRhq0ofZ/
N9x+V4+3p8M/FitA5a9P6N+Pyu9GZpK8knPpkMeh6MR/lbsY+QaR/xNYx9yFcCzHDkdxXUehiPQU
esHscR3gmAExsHR4hnxH4aeUpL9QGbdYThqJ8Nxv27mY6mymO1cNuSrg2MAzJvnKBpgUvdSamtH9
4zFvhQOQrVM9x1Fytk3+w1OZWmz/ZygXxNqpwnxtvz4uCnrxqgwSWpLwC+8vpPrMCBVCF/3xWn1X
DqfJJsimpMSQK0m2F5RiteQiouEThPZ4EuN4ckgL2lgfzUjRb4sVaB7yzw4tTfOJnjfAkQU+VOdU
hN2E867UdhOF3KV9ODY0ZSAW3XInhodMjMiX0WWdlNtB9K5fFyOJSO5AEeSFPVMC85hi0GDl8pWx
WlQ1XhKF68cBV0I06dNyaGpUemMxewTlZFBBveFvtRr11KGshsx6WIlwUlCV0oD6a8g7GTz3QK7Z
KoJTK88Gvf9QH6kJTVehPp2HUgZ9xgMtkIi1I1Bhq1NKUc4i3lp1VSwwtB2q2NVcuwZ6dHT3JVMi
Wf4kvnwzbyVwR7sDrBfUZ1JVWG477m4Gr+GdHUCRq7fWkmPS/rVzqHy3oIavN6/H8fbyipD/fusG
ntSTxlMwSY3Ku4lfCDgl98/i6iA8dGRaVL5iNA/H0zFknkhRDZOQK9b5V8YF7c/pVMHrnipf405y
d/MjkiD7QS9iYwNX82fcrZQJlPYbYa6CCUuP+43q/Hrc2tVWWXk6B99vUnPOtFqvmjZmV9wq/VoJ
KAov69ic7VGaQ/fBQKM08vxQgJjjlsD7GVQGRAG8J7J+WiVPIfPKNIO/TX6MtWSSK3AAou+L40u1
HV9hMfQNdfxbfu/iNXkdI1C8CWrP70db0hXIeHAo9CivIL1JLK2QDfFKTODe7WnrkMK+iUUbAXt6
O9KTFOKj21RbdkZmYl2StUec+9BjspwBzh7mK7G3sLoZwupCh4Q1IdiqV2z/DECbAeH6x1dbh26f
XUkfDIJxj5ijnplEm7zFpj4nV8UYZWACjFCHP19R895+KVzJUt5fvRaxaUxB6hQsATdd+mrRPZhx
JRMssuhPS4zcTmu4kiBcbAxPq8E+1COP4RBPDVIuEIybu+Y5rdrEaFXn7tBR32PexepLW/8sDX3P
oEvwGZTqBr9l3WwbtgR7gB3qQfrMwO1Iiixs1Hn1xV7XM6YWqVj+zT25PovosIUmj5CS4mWhDbkW
xMipBnk/DpUb0cl1VAPdNYwLzH3tceyI8y4A6SvH6NCsyP/kPV1YYgv5kJddH4pj8kPyLiGnjjE7
4LynuAGdGQv7uxfp+rVv83FeKnTkr/h+jQ/Vsgiyk+9QUxvB4/KCzAHWJEWAvZN3+7ANYz2cz12I
r0debGTem5fCAkFhiCY0Qzwf3tjmMLAmqafpQHdU6/BDhbGyaR1Xrz2mNsy2YHLogXeJQ172KJxn
LAjNpl7PqpfTV/3QU+FpYvtZE4C1RNX1F9xeLki8KAKWI5lXVlbDRoDYJ31EHeSN48hbW5Kg8jmT
uWYGjVglpGXGmj3dDPehAh9ONjBhrFZEjDX615Px3OyauKaAiE9XChEtHRhrDUmDks+znPp+sZqk
1fTPbYSLon7bNclHeF2xZBqEb30i6bvmX6ppN4+fnQRnjF3SgiL84YdAblUo9uAzlnjC9z0sCT4y
k5qMqG/x7YUlHyc1EN9fyYIHrk2ynNRr9lVRlRUFrDayiScv1i6MY2LPG0CAyAwVsl8+G41rbtXt
aTSCicK/cevwUsJTabctqXuITwEOvRAD4AUnNwyJZLGjnrTi+zYcbvi8zT6OyJhyTnsyOO9OXFxf
UIyn6Dg7286YU2NKByIg5X5RmcryGffLd6TtupmbR5P47C6K+Ilc95TlOC7RHa6N4RdbjN31lqLD
D9VsaUpUQKIIc5z/9wjKP6zuO1wTScNJtpH/8h3TM8ghbyxQk3QvBNgPLlMeXGfqUJLJmqWuMB7K
+LsEqlcM6mhl5HiUL1AR0ngQG1leS54paH1A27Yn5rSf0yYOM1GC4w80ncDH7GWata1D/y2lus8L
9IxTBGzFweGVxDGdnjDMEWbmiE4yLHzKPBRGGKV4H4pHTOfTziIYoc7R+GUNqorkAnkc/camW1qH
3EBhEnlEgKkaM83ctSfRxBDGksnBmZYroHKRxEKH6El7Cu8XvBa6v2Jhwie7Lj5IcyUzAj0LhivY
4UjswDEcPoTgcw+G9UxtRgmoLYwRVQ5V/mo1ekBrBtakgkbo64bxfLcH3HvEnEDFyv/WiQjg9n4f
OjOtkmKsFtePvUNQyJv+zLM4QMwkHuQtWZ84CUm/EWufGxdmBBDfTcGY+bdbGagigl74/6OR56vb
iAA/5bSbK7gvzU8SK09rxI3faTZaXPz3Lz1ESL6IxpNWFkl+D9ox6ZnXIm+uvWNUWE1slOWqgme2
PakTBJOqiHlIWIus+Ys33IbYsuN4Me7h/0YIxShiXB1etMmWcYDkw7RT1Og8fj/1ycBCEcZ+fkFi
RQref1iw4XOMvVxqHtMl2oSCb95NWp/qfPE7GxNUprcWF+H6zs1syQweqihNujwdVeXQzExkl5eB
esW9mSuLtzG5t95TVuyBg3FTRchKo2yuqUh3RFe6nJljj8+Kzpe6pJumCI8SBN3in9mqZ2tLvpZd
7QBeb/peRnPqmyqo2LKcii6q5EczAgCXBAxbMWtTBjKieVEfyaSl4yDTY4fRedvKFsJR6bKKVKEB
N2D0mzkbcy2p1GmqUBxpE6qgLtWnoZeDlyJbAhKXq6G+nnVMIddc+TBYRP6G1d22FoucD5E5Dt+z
PVREKHeY1x+FIRfHYQTE5GYob3q0LTJMzPSPtKLzSQ5YbE+vYWhGj9hxKuaCt0hD3zV4+W5DP2br
OHOqLFTgMKnV4mIKlnvEHKiBkdU7ukeiNDEz/LCiCpT8Kn+xx6LipMeTL7TpkmhoH7wo1TLN+rP+
vgaDF1ukJ++cKSe6ghB2aeOYcv9/zqFD+duuQPDgHCxPxkiO+h7TGFxhX+hwNpyYyhM3aRCAZkFX
2e1epDH3oDEfBXYWqvvHNxcFvhyyMAxOeawNbT5IIPHlc5Nq3AKHrDout+qWzSK1SkMNfDWtct9j
sn8N+tGfq9cvXuuJia4odReAh1y4OhPxZlQZcX0bVYHWlxSGPibwKYvntA2SNrkGk7Ulgp8lFZox
VfsBGyz2HVlTd6eDM7xFn9XJ8shbisCGo3JE9BkhAfl7SLJGXUe/jn0xtJO3XmnRWGAorazsmAFc
jV0KNjllzhKPVzCQPIJENQi//0uwANwZgYx1vsR/GvH6mtlghG+TbR8e+WArEpxmIswrG7Wrys4s
BIiFgfLPauZ1/VKRcYpG4eu346DySIdtrPQ2LgbbNDeacaUIeap65TC66MsSgS1xxRStxT31BHoV
bz0r0kSNzRL5F0IjsiK1HRMRYqUpdeBoNjEW5AnEAQdDRbLEHwP7rTZYsGowGeWzAsr63eCXP24P
w+SxxVIx5MnYLTVRCMZjZFmpiuGV9p+oIQGX7S6N0Ouk4iYoTWDFot1JqWT8L6+3B61Pi1UHT+iJ
+vS5IpigIii8G/fQJa8aqhK4QMTsQ3y3TU7Czn1mz3lxhlrFoOg0wcKSuo8OouZlbQZj8KrcHzIB
Y861RmnwjDs/sjYgOHvUU2PR0h7bKJxroi3OpYcym1BqORxZWPp1x4oaYj/I2t7cVA5eVw1RZ/Ea
zDjPRAGBqFsDZPzSsxh2wM5/vIYygYSJ3yA2Qrm+EeEdXnVja9LnE4mAmnQu4Z1Fh0QuTd0KxY4o
cBdd8KdfyqyXlkue9UZk8zTuna3Yt+rehvqPjB5ExEN52wR9yGiilW7yuYbvQgtIkozIU9UoEchJ
bmsKZos6d4KeVyrFTMBloucFaJTDjPAwaU07w6phBVtNM9ATBPtoU9sGRAy54xiwHmhjlT0gj5iy
ZxSkdKQxIhOzbUS3apMHduuRoXEpUk8kzxdGhypt8BceZ8OEtCX8MtOy2YT+9YrZqkI+ehIauK9d
vztfcMc8az0bJhhg8JOV5aUKBiOevG9VbiD9WPD1Ut0m21XIbssrh3pxk6azhK7hZquxE4Z1CyAt
BSh/Mg8Gnfh4Qo11eplp6zaiwNRgdUZJkufcwln0eXkm30OSBq+VZKmiIAqXK+RSfLxtyAPqwUH4
ez+EJBvMq2UocTX86k8HwXbeazIOb4piS8bhXaxKv1xDbqc29ikwYah/JWH5YzcKKYS61XwoXu91
fodXqD+lZS6lXG/bWtqgKN7ua/jjEIRxfK+aK6Hkg0EyFO1+dVH9zivoL8igIPd5UuJq5R3gUC8L
Th8+SZ7/ghmtsPzHOiilqd5u74lJPhARf5RPEkJSLnYCRQCCNbMYjOx0FyjB5hymerX2Waag5NiA
smm+IPGunVJkr92zWXp0yVzPK8nJlyR9IrMlPbQ3nNveWvicMJ6Aw96p7JS7gIrqXsu5hxyvI/v4
vif9GzJRQti94DOuWKjY4Sh4HNDxIBGFs/bN8XDRrfx8fuKLJN8LPEign2OUjdlonJtr6zaSB5xd
F43DAsUrzhZF+myHWlDBYWq+5H6hxqFEmiRevxKTPynP64ygBgKUiwkhmBwJgSenJK4qydLzmOUK
a4QIg1mGQ9MSvHamwwPeIbS6cD2jt1Ty+q4v0Vn+kpXtavwvXNpnlbb9NgGh0aqlvrfFd5XWa/Ux
b8f3tiGv5D8dd78JezHc+o85x1DIBX9GSelKyfA52BLpQG37aVWyVc6FNuTZevzHLDueZXm//3qW
KNk9jE+ZAIJM5j1Wce040qDBjteA0yIF6USWpaAKhanIIvKWAT81paigHui0S/471YmyFHNIphsF
WOP+eakOb8mnXmq4A3oO6iePgvHwIit06yhglCI/KvP/PP9gODaz+dYp4ePRWq+4lBSdJk9SLcN5
9CPbwolBY19dmcJqnJBStVTFd26FLss8i00tfVN0Yhd+ba+ItXGjFV6qcnPKCYOoDcrMOZfFGVRQ
kOVGPb9lx0OVYenA2DFmbpPQYLehPojlUAwpIG81YxcuDwVEHQBuKJ3py07LizqHxkEuCUH7uSaF
xlIL8Tyir5Kq8hlNTlUatQ2beLvxaZDMh94T4dFY6SWt2iBVfnUksR6mPLBRM/51u15N4+q3ypC1
dFfSZotwGU01bQBfghqOPa1EUIXt4TXcHqjO+r2HIdg+6xVjPfSt4XBiIRWEqNWwDubC2A1dzFk+
oXC4sdX3Sa/DvniIjEYvXBMIwyJ4D6dQ16X3R4oPXjXvuL4l5QrOwKXAUCTV5tnGNvGm2/y4/CMr
S3SDnmSSYgX8t2GHxY2L5e6rRTn4NDtevVrlZQr672rXZKl5ExCNQLl0JI/Ep3D4uneiM1cEua1Z
M7sXjIymFRYm5zoGi0OWWrd+XdnAsMszHajRlBH/6bEdvhXroE6oPuKa3GGJSBwigunPLHVl/vuN
IxspNtmMeb83doY1kgjphbaW2sVvhxS2tjQmyVf9zEBGBhLk86IbYa+dbnn264Zh9E4X7KaEfEd0
Km3Rh1GAMzsv+ex/bHvU710XQCAqFiA/nOwr+8vW4GWZaa7lIS3n5A6x1++k+aIB8ihYHoTzrTIN
WznF55efbaQtkQbAOOTMrdkVHbviGRqA7YeEgCHwxKnd0Uqe5yLlseT4CS1fbK+QNSbOVZei7X6N
ib02+JzXYft1WJdy59I3yUMh8RgOuL9Ja5WV+zRssxnPN0hCbgU+2ZQCLXFZ8++Y+85Hd583/Gx0
St8oRgc13DctT+o+Jnt8FMk2vY0RlAxiW61aX5GCLxdBnzfJNQhe0LLkBFCNCy6UOyRGiJmRIcfv
RZPLdudsalCItgC9TOT7LOPoURU4SJ7jWFoctDqqJV4GVNzWUuv929jutlBj+MMz68WFa4nooMHy
V++SxqBlQ27gNdiRaZuuZtCr79z/IN0oir3ujXT39HuFbtDTayJy6qcjXjMed0ATlcGwDpBc/zee
9p9dGE9CxBOgfC4qz6EWtGzD1q9pu+BM5KIavN9IZ6nOH5ajK6RiTbZRqxfoLjCPCOzDNE5rVMXc
29k8i9uK7FQik47tvaONnJdO6DFl/t9s6yHUcDaxA0HrGKPl3srzJzRvRxgRTe8HiE0WiO/wUJ80
FcSQRw/zZCoOchxHIrZE9ebcIfDgR8ji8kSogjOlYxixqKo71srvGR7ZZCBwVPVEJJf89X4nvPk/
cES5nSPOPcCO3N90RRwyIglOC/tU9CZrKzb6lqWc7EMoIHZvslABF2oY5YFB1NKIs5M3JeEOwbX/
KJBOrmYOs7XPtmGEXVM6cvc+yENFYzkBo6e672/1Dpp1z6rK0oQMvpadYgWvil+7fMh83rKgXkiB
vOykwHOKDEcq1J8aAcyALiR4R2CaTfRDEKHjn7LhZwTDvoeSoa1EihQYb6cEq8By5PHnnbxyoiO8
S/F9TaBXg4Tw7sMFrFwNomR7HjhoRl7nKyZokYMPI3eloqRq7v+CVrtWtUakDnBAkunDufTqpgau
ZyrI22PglRg3xfULGAMGID8DBbt9/JurmfZPz7/pv9iw0tuMq9/xTfjAMMC4DnU3QS3jqqZ+eRg7
BTtiVJrIkYqTZ70ICv1NiDr4AKZ7yx3bApaE6uwTjcD68HhowP1QIPIX5/qclt66BFLHgnX9MmNV
LWTw60jFApRgj+xD5ynXpGLLgb2nSP3CW4dO6NedZsiEnUUV4wmknw+ydiAjTj9tcRK6PR8U9fuH
kO+SJLNRaUgpgRIvcmTusFORvHAx3HLphzqrdVI4fD3KRnrfrTEqg2h6SG8kqFP+5qj0lmDQO0b4
yAbA4j06Jl0KKHs4qceLn9AebZK/NKD3HPhlE9wq3Te1Ppym2hgHstdm8H/1XZxs9VT5WNkjimTS
p2Wv+adArTrYoM6vvoP907yAQ4ekX39m8sgdjkMLcaEnlKCvFdCpf8oIWQS9MiQsf1cJQcc+VUoo
f1hGkvXqjJGUxlSbyZarBUk2BEerX+eN6xQ0BZiDitTIJQ4Gu1p4PLhIV3WjMwcyquvsj48IUP7f
x8pFZCMN+8yFVQ4mrEg/Ilz2jnFgb6WpEg+BUO+PfeLDK+bm2+6cOn/cxZHaFom/eVVqLXGnc2Hq
IHK+peORv4WUMAG6JJPdUk7rApLkPXwgbHFEmcssg8D5cPP3uwWVH71y8bbyyQqw50hZzpRh5fud
ADTeFZZHvj5cjHdcLW0Tz6qJiZj28Z6VGwUipJBauULwfQbS5taNB0/KnPK78Pzjd2l/I5ImbCAm
ArIEA2DyHvaj9H5F93x0iX9MievJyl38AjESgH8q8i6LVvL4duB1oXAXAvaXauoCaV2WVADTyy3L
er5IGvdvI2XkQ9GQJmUAk/LuPt41JdMpngAdrsNa4SlnjPlMN/zXYTsCyokODSnNsLUS4oCUEvrW
noPCScDbqubCaX//IYXZE4vtiGnBPQPre1i0eG0D8f2rdfjPPPRs+Nohxpcc99D+cjOfsZ1bm/aH
S4+qP+Vqb2EUKlYj2norC8m/DmAVz5aL8gT8r4yIAmWZxcY9mxA/1KuBVN1D8JZV+iN1cmXmKe0j
BsCFaYcXpqPcbGhxtaOjV1xp6thTAnXZnlnTZMn3z4igxRlS9T+Ml3QAg3e7FPLdx2Fm14Nnw3tY
iBMksgL6KmJmEzjfvaVy5I9CFf9sZ3lgoSmHYlFuRtpdClkGhcRFId1UCStJZiKC/uabKPJpbJ+P
KL0ebjJMDdzHxJNcpc22t/jVSwA63NjB9lthQQjlOj0v8EdNEtALd4kOH1GU6eEImOGdvS3tGsx1
do0c0vrPMMTGC/Cy/iWEf0F0+POMZQoM2ssZmnGrjsYfMV5VHHd+107zom7cc8Tq0Os/YReTNHki
uVYHQRsF06fiv+udGX8u4HnUFAls7cqA9NFGz2HLbDdiL/cKrCUE1xk0AbNJ4sh12D1ptSfHQd2L
11Wwk69kL8xvv1z8vs+yAzsg8U7SsXyjhmJ+7CClDb2gQy72EJ1I0ePK9F2LsoT5b7+NydifDZhT
n6qjYfTd2XaSub61A/EVfGy0Peu6YIrm2xoQLsFxaMRpUue5ym6jjEEdmckcz+wZ/ijMulCnmrhp
ZkDSIRe3salcF4eONj62cxpeGFHCV1AN0k+oRbM0d1CtYFFB4zQqSnpn1aWVv6hyEady5aBkJysF
OpMmomVOK1rHQD/OV9cPWyJUrFirGKAForJ8bpXuLOOIprCxWqAe5yK/5Q6qaE8dy1aJu76IYkVE
puVwY+lm9eFZBg3rFFG98HHo5Ha4ku1JptygXunhM6RlofcjG8283FeKFg+CXNbB2cknKYX34TTh
pspGdbp1OICMlw2vH0x79uMSlK1bS4ObBfOf3vEpBhg9/ttd1KNJj+nFvpzqm/t/PYwWBiZsz95d
rf/KyJ0fjdBu3Q0t7k/y/t5qMAPlCz9vtl0/LD32bLID5q+Q6pDfeCNtofrVxZoQGHVi9GGLIK5J
D1DoNf524b/Ce22IKG1BDZ/DvZIQ6xSL4dW1mnTVVl4xmurn9d0iDTT5o55F/OC1qJzL4DpD1LAD
2K3V28zgqWaf9gycScGkBly4iDStl+Xr5L2QJjJPbIdeVXgHUi2wlZFAFetHKm8K7XmanZkXlpNT
yEfhgp2/6cCE3MxOQp6pn7f7TnGJFHK0+1bIQxbfY7DMCizyE3xVk4yo8tD6uSjZnCBxYiSHkwxV
zIZ+G9gdBEYFrLsXTpkJPbQ5lR+92De9QIBy7Wq7SPl9HZ4RWMU9ykUhlcT/lv5D+tR/gPQlL/tX
eWggrvM4D18l4vqu6ORHnWBaQmj0nfhW4fzJg/NFWQ+UnmrXjwGhObjm+u87KQhCXDS0KZvNUTzK
9mw2wYeyi7+QPWtWkxx1IDQWM2N91NZEZjTKItGhFuFRl0cw2PvtiZk99Iv17gXQUgLS3qNPZxm5
vuSOKWTmdfKhm7t9xd/+ZbzD1e1CC6CwpWbMQjxUHRHtBtePFpwN5YeJHScdcbvKyp5IiJV1YbRv
F+gc65kjXJc5cvmzm6c1sDd2pQlFAQxPouZNYiDuKNzF6hKfywLNFnqyhAG5RrJR2UzajPnl5irz
xAh91u5c7V9s9lzLE3ooBlCRLxKbEo+aNIbEZDL1VF+VGo8bbHz9WcAH9cCT6P41BFJxrTXbTTg0
djVA8Qn7JID2r3a9v1utSXEbDcoWYwilLNF1+VV2bEBcI+H/gCa+9vQjqFi89THlitDLTlFLly2l
7I+CS+7tqaS/BvCz1ZR3tuGZfxtfnGvQf1YS1dZCVDNxSHQ8Gm7msoNVBEos32cCKUa03Xlc6qSs
IYymA3VKJPdzPEQmhpIQZgeF8ZIlpdfA3ljAbJGbFcRFnKyMdKC/UIU8ORxiZoiS7bNxoXJGHo6M
kVVlhq+oJOpWs6Njd0iypnWll1K8aYHjKmJLqUTniPuMrZIvHqflZjB2P5TObjg9EmYBIheOOT9I
AxoPsL7lg/KcS++yg/W8WDAyg2Cobn4Xr4kFnhPKa6WL5u8AlRHqdO+lboqYtbUEOfNyVUTlsJl1
0Nvv4uiRx9ADj7osteRVjwLoU4rpdsnxW4i2G5CQJ+QEGLsfzknLqgwGKZ4Pd17yUGHK5Tzm/a7P
1F0RoJQJZ88s/hm5fAL6/VS9la52JLnoMwa9mrPlNWoJ4GLYpAtK0X/VV8fe8bIdCnL2QS/dD2Qm
aaI88qL41XW+Qb2Qo3TN67yDMgneblKRBCzRd5RO51Mcql5RQOvnp7RojgacmB4s9sWQIjCV39nu
g65NIZG5ZU396hzjjvbMMoP40SVNZRYfrR/6eKvqDFjkDdijEq3QBjZwVzCJr5wCuI+qys6GIMP7
u/epIdiVdxUGjVCNklYRzs3sB2J6QaNiQ2f6aqRPl6E148WGiiju5G5HtX5o46AVQ80dju5EafeJ
aOB1/qdQwcBoJB4c8oNWGj4a1r9pfakJpqw0fjSJjVRoZjvxMN1q5igFgv54jILzh5z8zCVS5yVc
90K9/PmskvaIpJYfuQQVGbppvt5mSiSblgeDaiZBq70VTyPbBRlSEWB+PejBZCAl9fQ92j8axatu
lwv6y0LEh2yh+GMAjt9eQSFk77+9S0Ft1hd6V1uNXb/cQ0Gni2/q9VeZaAmS3NvU89QmOUkkwEVN
gOQkCH6qBiJ8kwtNwBTN/5lsdqZGdFmIanM8Dm4t1oYoM8aNsxO8Vxz4FHlt9A51ks/4Q2asawXx
pS3EyTHklUuITaJv5vzRfm+o9UqLl47XnJ9KkJ0aFGVgNpslinLIQdykPTrys3BWAc701MJ9rDrR
68Veay7NzViobZur3inheDviqZRlfNE6hTuVWnM4RMuYA0vHl3fbaGV9JjD7mQizZHuH7gJquF35
qj2iqT9E1mZlySCZXZg625QPfWrvZ3oEAo2k5QINKJoNnd+MrSfZQyRatNbhJumlJV/F4SYdqXSX
jaziabM4sq03vkJHzejX8IUeiUUKpcczmlSCelix6gKpQ7fvpmXCSry4mGGjxSqCym5dyaAlJ99a
e9JMgodZg0hKOedSpq6xCGBcLSN9wfm7Sv4MbRn/rpi3+rCdQ8Cc0hNneoA6K/Ycdswz9e3JOeza
ZNUAw8/c5NHjb7Wn9lNcjK2vIXi/OmvpZ3VSakskn0VssltWHLPoiXeskty6zPpOf0bFRSMuN+Ij
61xyeFoI8xjAhlxChFyqYilk8WkOxYsa1+vIAdz7Zqg7D1WE0j0HVScoag6fa5YAOn3ssFDBrJVd
PUQe8zDnNZomN0gwskoJo+GjLWjVFeRsUVXHJ3q1zTQZ5NW7iU58HUQZUPA/4PBE9e+pCzwKRzge
JPLkc+bg7DYsYskk4XR8X3/WRxXoiGIr48Pc7SuCCle+rDY9uhSmZutB4A4X50Om5BAEvHFpIk91
3VmKGEs7bdk8gkHOSvLSIzq5G8G3dGxYq9kFZuTJ9QbvYqFUxT8FOR4GRJk0v8vHnO3bY5h2wiOW
L8xcwDHda6O7spBKxol8muFHdSAYpgYqwrQqbPvrOc5znRrZYAjkzDG2yQWNwM6RGUGyaEHEuDB6
8XcAIaC4BcZCLNrccZeTg1Zz54LoCLwflT8Ha9ILlz9OavYeZ+PUiGjBA8Nwf9DdSt8+i3Ei/JWs
ASz4i7kIdOvimAVKGF3e88C9nXnpLlP5jsYU1vOF3rTRN2K20PznOIId3+p0OVbEO8OwDGiJYBz7
bdwrZYH7Wa0nwx8aBZZrbjUun7Q5dtTzOGvYwBZg2vVFuAMW4+C327FjNtIG7fTvo6lQbtbAzqjR
vNC24aoNz3tpx60Az8tUIYHyWbb0oK4cXZM7J08zZBWl6efH07feSB2/gFZO8IdOXtG7K2dLSD2S
jD0TEfvj6C/MnydRDfWAWIoLtvhuvUAYb9w6uXsBWE/773srorzQScg3F2qXMLZHEALpBFMB5lKU
IGmezPeug4Q5+dom0cNMilJHP39g4LRkQDOLJUdSeUmLhW1LRYy+hLVraLAJPR+VmILq7R40bCxz
z4r2Cg6XjxbhSQ2spdUEkrDKBb7tWi+11QBnk24rgoNKU/AWdiwolBRpH38B+dhFmFDa79atjMVY
C4BQUh03vTGY1ij3PKGs74fZq5VM45r93NFym6mivnD4YrP3sz1vLPBgbGruXb9Al22t5KFn9l3n
iZ3BkAD28Hx7ThHlLN4JUJSrrSLzjtj0b1RiX0R1rJf1jCWSy8/Sr7azHurN0UcnAk4L/7m1ngb/
du0xmF07UG3Z1J01scBFJzVMJcTsLgGpKitQQHQtBWnMIJylZrBfZH1Rdf532Y7W07SMighDPyIg
SLG3vwBARNUSYyAOnHOXNON6W4Cobv0GvgtpJ3QmwU1r/s2U6VoAREygwYwXzh9981NQwrrrjQNA
Mq2E0aSoja4dj2MSsJGK8+h6d/xxRcU9VsfPvQ+gVq5S3cHtapgXuILs/aGrmtXLYDraroHSOWzx
LHHJp9fHif+BrzjloRK59FXMEi3XWSPoKI6hX6jgvndAXYiw9ILvBKsXYf9p0b71LsKomCbueXam
t1OdwUaNDYmx8j0F6CvvtuknHoTq4wSUZuprv/4BNSk64TFN+vL2c/J3G7yc3i56VZ5pQNeln/wY
uJDYCTTuDyB2S5HD/D4DZt4jfHtdhvFJT7LUSSFXXs2hO/6u2sZIFHa+hlilLTj0i12OqkejZAlV
DY8U2gjro4P66ZPamlkuYyrsludOdCEfxkS9x4LWJJdv5SqNQVSs8Bz5jwZoRf05zk2D2sjjKdaT
eoTNz3LZyMIW2KnrmZplSlcd9pjV11ZwQCpDNviIK6UPd0HeJBubGFbnBDYK7r3ancwtGDZM4uLI
il5a+XQ8OKuKgVVynJd/3Ok4I/CPqmHcj8053yfmm1cOpqjxdWPPa/Qxro/CzVhLohm2y1Q4vm26
XZQ6NdU9FLVcrx+zxc24N4jiy8yEuhNQxUNmhz8CKVTPI+Jk6TznoPfzqjMesZCjDS8Mz0RYrtY/
BOxayr5S205lBCtUxx2aAap3yBXValJvy34QYhsACuSSgwFG61cSSGj1Y+Cbk2prve00ANwcsh2V
0lH/oMl1iTeTJya4mEH5TL2+dfkKAC9MAXoMAJ20BUb8xyCFWmUUv5QMlp9dJVLgCzlsZ99mTNIj
FGM6KKvK+D+LLvuFdqGyWwooCrGEPtIuJ6iMzeRYE5RV2Aq6DSDaiitG1WlvJ0dhFsdgoqXWcpDe
qWGAmI8k7zFQ9YLq/iw2KX4Pi1Rri//lHb0dCRlqZGv5Swk+DEOqK8Lyhqk4zv0Ng4VpLeIa+AW4
ZXGBB25mTycw3HTpt0rzkmnv+hhtt6ACwwY+aftSfu0IMnL8p0DpIMlsno1KMEbwuGFdpKjSIW8B
2P0s897qCHf82+YXuTW52pzsWSpQ7DQDd6VEvpRHWQE7l7V+VJ+4CAufTqwwp9JSobbV0Ygq4WEN
9aPvZcNtRoNTKmM4vIT0PnE963pMCtabKZ1m69cyg9JWHy+jk/CQxQX1fYJC3Ue6kPc/HS12KSL3
apvFisFr1njzUhuTl/YJ3K6zhSCASY/qtlClwwV6qhQ6WQW7S18mlekJyHWPgJXX6jMgMLAPWjnH
3DgyyCGaAmvOysAHV8D3CeVa+19KPNjVPInu9ejCOD28WU/RDpxAnXVQxJoBgGy0Mmn/qekScP4M
nbUH2q6AeE9KjCX9ptb37Zp6AiBNJFseuu7RDTUAHC0js51qYkhyXIzeAUOk3yHW6cn7kbRvskHh
s5/sipewXLbBhJeZQQpFtBLXNKMfURMBU2p/U2LLk/YEd/D3sgw5QnyMNzi5zEviTodcaSMEoIn3
aP0Cvfi+cztRo3wMFDXVe/vPiq9szJ05gs52wE4Ft9n7A3NgJ1qBN2AELqhcGuonqZeXa7KyjsBY
wxj8/Ou77bUIpbsusSE0OAz5LeuCpYHtXDfHKN/BUZsRWBrXlLfeuJ5pNTKnim/zQH+gFLqHW5Z7
akyMvJA218ckuGfeBaoh/Vk/SSua4A73a3Fnx0UxZuuTbFZoO22LCSTFuK70UIzefRf3rFS9WSTr
GCPqIeFNb2pcxovwFxprRrkdjDwj5x2cfQPeE5yLX4zOzidegswntR+sUuxpCddL9v1zQM0H5mbe
kSQCxKoeXqktKgSWbObqEgybm0ohr3ifsyxlHWtgg2K80/dKqnfpugkAYQPNCPoUagg+PX7ZUu1U
nemQh8MbKk0AM+NfUNyH2Hghnh93MeZotcNCUQzx6XijOLocqxCfrKHg23C1wLhPKOplW8Fv1596
9FqoGg3WytCviJkaIrAURNSLfKPx195XmcjO6T4+XBRA3MrULlDruUjOTKcqnFUMAaNsSFjyfe4T
9s4DmdYWun82wuef5JV45NpFL4iDSi0kZP5KnUiL9pEu2ViJ0LtxNG3S4ucJWwCbakqB0AvzTT3X
mBF4SQmrPZ25WGUQvNTNyVWhxg9fio0HfYpXYM3kWSOnzfKZyZExprK4sOB3sJ/ThNhtDwZSrBQA
zsW+oS/Zyi/eW0R0gug283K6vOpCxC7CUa3J05cZ8poAnY7F7MPwFb+O//G5JSM6Q4NujRLUF+gv
Ca7HESEEg3P0gDVZdgOBG8EPDowgd+3YdzWP6mt6jrZq98odyTQTII7bGTuPMmVFogsrkb17++NR
KUwfZkQprwcU3+sTc+RXmNu4VjZShlEqMRSqG2m8xBzRNOUcehapSuWfpKv9xKMEo9ntvtV34s6x
+ao+Elb+lElunrfJJ7dayMtJh0wvPcPCEkCQeYzTlNrV7HqbxIoczjZXLxlomt0B6TFnGpn3pncC
iAmq+e4nWya56C+qMdRrW2imxS++d68CnH4DQKjvFrXI6hrkVcOjVgDcMowjHjL/7t4tf0GAXAKm
/zIZcu2ihZbBOnGGkmtsHWFPu3tB1gSVqkxsQ3gahfrcK1G9aXENo26emAvCFyduvjCRatBcQ8Cg
0Rau6zuYR/EmVC8AqihAKFIehbSmy5eNxlSHq/2kiogRUU8wmnbdtYuCEShvaCVoOZSDNVHDgBhB
/OiebVQfyyJayNMTcZZ4wOPUbhyULn23CVvOjhCEV6lLMxhjdao3KyDzm+dQbzZF9ug/WOpQsGtx
1knebrGBXfucELFcckQJp+vaa8rGLY6RiR7fXuX6YZlJOen8YU/FJ8OREJKvUQHUNSLhyCAyLmAI
QFOTq//hjKkhvqaZM21DYgV9orh3UK7q+6MpU3s9p+F1n/5tLZ0q2FvoKfglmAntzFs+wwwvFJBm
Hk1+W4qp2a0EBWbiJ5b2Mn/hJh3QNWPYUkRt5IZVTgQDsnP1t6cElSzv64gyt0feH67KqIeSDaur
rLux+S93FukUBw/tdOPhl+2hUzhG4g5GCFBMg+FY1FQNA3FIDH42BuNau41t9Qfhg6aRrOLe3VRM
6KfCMAx9I8DegGdYBD2rHcdUOm+w+Ki5aH8mv4gQfFOEUF5uRe3O+d3e0y3pLgZGo2VQpw8HBsO0
YuInvLCh0S1fwOK56hXYl3qWqdmj5wXI0A==
`protect end_protected
