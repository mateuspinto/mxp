`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
HI6bCReVuVDTLq6Ngbwrz7kF2afxJM3hSiCDawCMHjwGDBf/Dg8YEN5mh+/rBCota7KHBrsRWS6Z
02C9IbhtGmHpcV+Y+00q+LaYdtMAt8zspDgreVMSckfbK9MTBzYWi1p9oQTKd7BoPhdXYiaHuJRG
otNap2/6OU334afdYEMdiyzVieIAOORYkb/I7r91lM9jyo/jK1F2A8s85mdZMmci2Jn0yqenThIZ
g+S9Vj8VVYLtvspzIVQg3uKf49sF3dwqkbdE7AEzBpgx/DjsBscaKOxZPpLs5I2K0Ps5xdLPhzAJ
IMs5VzdfBfRMKFA4idTBIN9g2uAHkCMUCyx53w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="fDkDn7BlqUGf/mZWEqlB3dUBetDqf11dcp9ZvBS2NRY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2464)
`protect data_block
QYvyVMAmlVw8gXDsrkNEHwDsXHrJ90v9PK93u6sIGBpKqeQNTeW7LspAc/1l5WqzTvUmULWT4tt+
BAeZF7zfVk9J2QBmYqF7eTlWhphPEskxF1aEQ6KvKx6sQJfU4GAk5giNptdWdaWya8nIGF3XSkiw
TzCX7TkbZDmnvGrvWERvelP1HnNoX7kd2MKrRwvbrHEv5UpJvcT7PTP97LM9VLCc0G1DBHwBCc8D
sBMPZQb5u5HcHcokHGRYJk1fk4XHEkGrGnxjx5IK+kiUI2SiinEl38xVi4jI8cxxU0l42rhY5QpJ
sbAq3phZEJCxwKv+teacBPgEklJzQ0IRPa9L6BhZDgZe3eyzMQ3KU8eND4fLRp/j8T0utGV1Lg+w
iU9VOced2TwFcX0RrqrMBX6Bg7UE39og8m9Olf9xbCIRF/3aODz5V47WbNnjSg2sQfLNmWTT1XNq
xnHPHQR/OJBLk7UifKnT1qDrlZ5RdfYwFZjBSdmtll/kMnpg8gu+Xkh2Pfc7nKHYHFKb5JGwdinu
VAUbXxAQEOom6KCxfPYm3+lp3fkapPiV26hlA+GbxZYl9WLaO+00jPfRfASYRk9/+N0n1YjF/c0I
4fwjDVOMFgvCEGvwAFJYDmCvPrLs+6LK2U0ceMLWIUtwXmBwW+YMXcwUQXyb7MpWhoprlfQhqbQD
w8WL6Zz2xXRNIHBtQ6WFW2jXJz1jwhuoPLu5cYxbYNay3XrFv2krbQjDjR2Rw1kppIbwcu9ZfvaO
RcEhLGjvQTnB5W83+gNzm3l/qQHYUFwF3U0Zm1XyQlTcwZ+q1XFi+QhnAEEPJA7Q3iab/vNjIGLt
vf2aYUezIfbD5KcutL8IPIeb41oa6/edR95ZFgOMxmrw62+/B3qU/orNHTJ1FcdWJPX39UeZPGCD
4osBEr2HVANyDy5idOhFG0GzZNTn5wp7DBaWQ2/TbJHAqFQyAhY/Rd6hI2e1K7xFemW44SkIUFJh
JJakvmDcDIsmCUN2w+tKWzz1PbC+Fa7O5w586Z5z9NUwoL0Y2r0YkACAsmBQI7DLSsYtSMqyrigg
80anrqJN4d+ll+VzckPQe2Q68100oyAYIJ1xkVseK2sD7ZGHYeEWGVQeHPs/goXecOYx8N80Ytk+
ZwBt3VkY9YRMxklknIWYxdR3/E6QabbVOADRewEB0fwhZEuHMt/Qt3xIiRIy+nv41+Po1PpSAmMN
Ct5raF6cwT+i86PJQ6LDk6tH8IIfRLxs7JwHsDnh4EilVOq12l0Y+qMYMx7VuE9NPcS4J0CvjPRL
/ZJDn6TChsEw8IO6lR3e8U+8NtLWYOa5cl/9IXbBP04cJBYCrZklmxL37XvM3wMVxVZzfGk9QqyW
N6n6oVFv0n2Sd4hMLtJxSpJBMK4Sd1e5xvmofqCtgpxK/XzipoWxPEpWBC/ivKfSwtdXiCejTu5u
0GwHtPvpNHrId7umDaP6HGDTZGq0qhU9fnIW0HRT9JT9l02dRzL5dRnD99UwYW+XaTmQm+Qmiv1A
4kKjNYybp46/eARNWRqzcAGNdLTDPirc4QNgdxBPHD1y+qRIj9pPlzEuKKMcDkHFLfe8StLnZvCN
NCEd8k7uKtA30NZE+3pek4tUebN9WnwOUeRDNDeXSsddSdPV41mQzfL2YqOYHzNfzGZwMsiWMUtB
y+DJQsD+mwYJ1/9CflfAoGxlsXk61GQa19+g9sSBsZoKgm+OnHKi4fRdV0hUqYilK1AOQjLMuMGe
1lClvuuNzmR6dAlmMvNDnRjzJLLSMkMpfIr0jAVvP0oFmdyTiNg0jvmW1S9mMXQGf9kn2Dv1Re73
/Cv9xuY4T4VsSevCRarVEacgDvFGz7aH5O+W5hpk2vffgVXoCDqks8azLN2sTlpVs9rol7pFfEXT
Zv2J13fjm/Vl+VuxWJJ/KThhXVHW6wVIYMtwoQ692tbvUS/v9VdIEAHlWevEUupaYSes7uTWLibS
uh1GkQu7e/qkwAm3aJmXNLLqUqZ3ujpol4OB+KPLMIKoZlZOE/L5sG02uEbK64JdYrZwZCl4IAvR
2/DEi9OQXBq43SfuZpWCZxpozMdNji4fiTjb8Z+HGA+gOLcjIbkgAK2BQcEwkeMnE9nNWBjpYLht
a3wH5UuWUzEleD3/xn2XU5PLKis4RSKDPlM3mnM9SoIMXOIl9Wn4NNcTxlrukFwr4KN7Akp0JctM
9jXd5FpWaU1pX5qVVWn1mXMJXFryQbA4WVM6JyS4Pv7/QyczsF4j8Z/XBZuzVNSK0LYXY76MAbht
Vkn3i/WckBrYnAtKy7S+BslkkXemXVV/OPLT1sHun3wlFenHs7J7V3vZfoPe2nnvRce6JT+xCoY7
1VcukRgOTBadMkwolXQ458bkr6pVvr3a2iMbmjoKjylfFc9UqWLs92us7M6dUapvXlEICOi11vlR
bBnkGTl7Loy1rsuWDog1ecP3FPDmyD8VcXGYW7ugCKC0wcs93EZR65Pr1YCQ90YR8T/twwjk379Z
Frm53xj1gWNqr60+6yXt4XWA8zIMqf6gZUwTV9+b7PPYLHP+jweUr7STKcHwBIySsZ1/NPfTbJ/5
rvmonKeShoFIYyRmwn56eN9QtcWqLZcCeU/KqHVM9Xs6hxfZV8vDAC3qeS0ANdDlN7iLpi1Y8l4J
CtXJNtzOueqwuO+zQt0yaiFUKIK1QYDpE2V24/7SfH+7fRS2o6sRWEsbRDrFa3NdeULGDFecTq3H
KoMmwH/AdlyQPlDcx0xBk5R/l5+PBFz97Z2AoKHdyhh+5GcJh3NmvBQHqqJ6MhLrVI3774EcZ6zj
nvO88sMbHK/5RN0WX097dyV5BSjfnD5rCBbLNiSSp6RNisFhWtNH7fWntls92qpLhjgxt+NqJ2Ln
ylBfzDk02YJ8kRrDxHFxJoVWsZ2mfHWMZIUl58xbsd/sCOGQBO+HbOiLlST6j7L/daE13dfZ2UKm
ubuqUx2Z4woG7EfbRP8razg81QjvgP0HNXHXgU/hnJyMC3HaPZeM8HHCTMi+dklHZXXuyDrpOtlp
haPiiPZbFoofqu1Lha7+vCDaKPypR5T2rHAs9X1HJtmtQDCU0snB8XKBYr0kZt3GP3ulT2zf0Bbx
LpYtg9mCLBrPyf+eDEbm7gDk9rUSlLxMNE0lKJo9w5QswRx3bbttC+yhqVv2qpKmQH7qFAp7Jw6j
WxvpV/Vv914qAjbXtetpqdMun/pe7hjn8oPT6x8oLOxim4T/CQGklg9OtusiM2JAHUqPSAdA1A79
rWG8iaSYclspclGsNA==
`protect end_protected
