��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���/��J�EPz���b��	*��G����?���X��!�4�P�q������$%�]ƻ ���׃+��H��[��>M�.��S��v�4���~���䆧̹��(*�+"�a:�W>�"s��`D��� 2c��"���E�@���0��C�Ⱦ��̿�Q�@�/%+
�����8b���M��8r�[�<hՄ�{`�k�1��}���$&f���<���V�Y�\���"���B�_e�.��=�͟ �`�Q��ge?�}��
ri�Dod~������@R��[��g�b�Y}����:�����P5��U4|>8���G��G��ӭ�ƙiLm�TUTԡ�f�˹����X��{����~]���t
��� "���/�bQ9�d1j0����]��
��>�$>�I�{�=r -d0K�� F�t��0m0�u4���߄+u�2��z�vJ*���A�ϰW9�ĥ���Эc���վ,B{ٷ��y5��GH�FJ�#��O��'wm\^��:zc��x�S�{��mh�]ퟴ/��pY��m�eH�\��y[�Ɨ|;���I��i�Kts�х.%��_�\%«��a�6�bLɝ_���Wy��z�F���]��
�ֳѭ<��S;3SUr�m���m����H�ע���	��*�a����v뾒��-�b�,+�x�~+a����,=�xL�/�2u5c.���W�<�-��L��'Hm��NP$q��!P_VHc�����ҧ��)<��W'��a�ߚL:CN)C���<j�t�hȮ#_�y �5�z�>�C��ỳ������(Mc?*�D��[p���~O��Y���lݢMZ<��*�U$c�=���<%����	CF.�]t1�xՌ���Ǹ�Ԏ���y^�o㦱_]֍и4A�<m2˻�Û��p�Rr���$�ӧ��I�#ö���KׯaCj��Vs�Ŏ.��r@��CV{&(����z�-"��F�.��㕿��|�3K�v�5�'���=ق�~_bO�ܲ#_� [���)D	X���7�W����Gl"Z,�]YR�^�����<�))�ZN�'�w�V�4�>?&�������.��۫uQ#g\��>}��n��@em�s��g��;T������VU������E���X��0��6���<��Vn{+=��W���)����jΒ�&�����ौ��'���{an�����YTB���7+����MGS	P�P5��[ٴ+���<5	�"Wz�q��>ڊ�
 ��2��N_o��S�C+LKc����"p�Um�1���h��0�L ֣�:��B�q�u��)��"�>ȁ�J�sceY��9�V���!i9J?�*��R��w@9`��z�	�����Y�o�!�l[�m�)�w����ߛ��p�x5�8��w��|���uQ�I�f����h�uA�;�f��\"oo�XM���!{�w���|�ƞ�h*��������*��G�z�&�ڪ�(:Fw�J%�Q�Lr�]e0bxp~� �X�\��3@����@$ZO� �?�H�q���Ν'B���K��3�7���7��˗Ca;���?T���q6}L��y�7ƺE_b])H�[�::*�1}��5q����7� �nO��8�^�`=�[ʹ9t~��CB�@vL�c�����cV��w�ϳL���С,��tt�l��f�<w,[*��Ėެ�z�H(�5!-���$a�T�
���Z�3[n�#����L�kt9� �-�X쬯ps�����;�;g//�
�'��I�̘V���X��'����EV�I�p�$��G-S`�����rP�0����W)MZ8�"��Nv�Ǿ�BD4`Jׅ��'J��O���Y�MUh��п��ȱyr�R��{�$�`?������N8��t[_p3�S��!�C�{���A�yjU�T����TJ��0��לZA�G*��d�*�K����\>h�1���w�'���c" =��i4��X��E���	h�_R
�B�pU�L����g���]:}��d����2)N�n���;&.�4�F�yI^U��H���G���I�
*�cU�)�mfzc��T(��DA@W��z(��4��tE����)��B�m����0���J�{/Tk=����ȸ(u#u%Y��7ky�e�I�6����=����8��º�0�:��Ԛ����G���r�@?eQv�
&)��4�oqD�2�:'j�'Z���n�'51Ȅ�G�x%���pD�(m�O)�2���R�6�2�w����Q��jm~�����xe�Q�7/� 2���_��C{� P,��;��Y���?�k����T�ò��\?g4?� ���ť.�g�F_�N�
�F�.��ڥ�9#%��&L~��=�V2�+cE��Cx^-��b|]���Q=�1N�QJ�QӲ<�:X�@*&��$�C���q]���l/r �,^X}�uΨA�� P�z�U�`��H����u�)�m��Z����ĎZt�����x��̡�ҥ��$����@��K@R�����Z�ւ�H7/�[��D�?�s^���^�s?���V�b�(йG���;��~��+	�X�9S�~��J���<U���6���wn����ε~l96-q���v!MY����T�������	oK��	_�2QuI@�J~}�N\&J�W��GXt�j�5jI�Zi�Vn6��մo��%RS^ܕ��h00��r��ζ����W%.������n�MC�}��L��XW0�?]G"_F0?����;�RHBs7���g�Q��4�d��吾����{�RmJ/���tٌs�&i��XκĶ����&�<%_�l:B����Eγ?�
�]�H]�t��
?�/9�ԑ�e_g�����>ҩ����x@���Gc�("���Kם������B��%�fT������#�%-��V��/���Q
!�Vz#�'��/�u`�n����߱��]�ejs��i:���:J"Y����Z�C^dE�W����B���ʆf�,Ov��䟑�wdիz�����lc*I�<��>���Ft�"of]ZF.Ib�R-����=H��O�P!�{As�ؖ�tHA��Xf@{��"���V$ýT{/������0�F5T9�K���)qq�����37�<���bh��f֙2���D�
�u��	y�.W���g:�sƤm���W(o��hЪӛgdȜ���I�ү�E<��e2��SG�#A���D��~�~/ RՊ��P�U�����I�p��^w*��q�;$yb J�3W6�
�YC��
C�@.3x����^�%���y
���$�������Ǳ?3�{[�)��I��fk?�N��4z�j���n'J�t[jO����e��7�|�s��{Y������S�20aX�t:rs���7.�a�-?X�b�]�.[��j��:?�F[ K���B��_m��|+�������Iy���Be�^�E֙/��d
�8ჺ��|jMZ�F�X���5�?Fޠ���Z�hLb���
�	j�`i�o�k�)�c�;ڋ��W4���WH'����sO_ʱ�JG�5�����nq��~���?�rr�#�J%�s�����;�~��(�����;۫� r���D�G�YJ�����h@w3�|���u	����H+59�;�\?-1����6,l��g�Yܜ���xӖ9�j��[8q��p¹����>$�j���XT]�o�F����Q��]��t]����F�&��d���:���Q�9��)@Z��U�`�0H{�<t�0�~�q~���� u3G�f/f*���[�B�8���Y��2�b:���O�E�W�c��X|[B��N}pp^jL�0�%��-'�-�I�s�[�Vf9B+�mC��1mU��0�;�pW�p]�nɺ=e�y�ƦG���T�S���ȥ��F��Mi�����yb8���G#���݉��r�I���8B��#)f�X���Į5R��B�x��1vg����j�-��&Y�F}b�@�����g���,���;���^�9�P5�`�3$���}����`P�z�P�� �Tg���Պ`Q"$��)yl����:���:�cI׾z�$��g"xC�;Ҫ��u��h�J�������(��H��!=���r����5��]�� | �}u}�ٖ4��KnOY���9��4�s+g Hd��?�3��o��"sLm�x�&[(G��z�{�7޶��W<D�>"i��~1�k����4e�E���DH�[NAs 	2���vv9<珙�~�ҍn(�28��MxV{���������w��߯ �$p�e����X�@��(Ag�Y�-K����!�x��]3��<ne�"e�Y�Y=j��F�D�5I��l]��q��E�ޓo��9f���mDj���[�	��Я�v8�ғfbo�`'2�ѝw��_�jQo�|��ў���M�=��
W,\���O�Ӵ�#?
Ex�i��v�����ݧ��,@�?��~g���:wg)ͳ�PA�$&;��s9z.��ư\�R���%�dK5P]*�i�FNv��wF������{ez��\�������Ʈ<�[Bi*��H��M�A�O���'��F=SF��p�b[>������R�B�\p�{�S��a/��_��ԅ���r�٫�^bs9s8��dGafhzfo�����GI�;���W�����{��q��)-9Q#�^8#��yЭz��޿��&��D-JMX�+l�+��>��5Mq�Eˉњh,:~)����0눯���&�u�"r���.u�g�9γ.�G8`�Η�X���s����-���k@�����S�:w�]p�ߣm����wD���#tS�6�E�N�ׁE*N���"�W��ˌqK����'<
	[ũ�"��!��	��	�H(�X{��L��튯@��`��f��y��s�q�8q�Q��G��P����c����/�&�$9 i�8nK;m�{Ԑ�πO@I=,;MVJW�V��Z�ip@$�?�t�������(��UiV��}F�Ȇ�V�n��%������@��L���H����M��~S2h���A8��^��-����l�/۩�AM�[CS6��VΨx����V���u�b���duYt�3�8'� #4�O���6�-	�rdo�x��m�y0q���p�+���b����f�a�1!Z�`���u�Z�� �4�Jz�]�Vt<6 z܃;!q����e@�$?hgS̯��� �� @
} ȑg�R ل����3����K�<�	�Lz�hW���m�ꅃ��1�ػ0@�'�������B��'B(�)�l�G�ȏq����+6Q�F(Z�����ʇ�X��w_!$�VG��<���I���񮹥�;͛�-��]�-��Oq��D݉K���8`7���W�(�O:�46��I��\�F���X����A����i����"�&d,�
ì�F1��W����W���C�]�ODYU�D���8��Q)���m�3]m<4�J�(Y}i�����<dk�M����r^�,��+S��Ys���j� ��`	��+��Ax�Rw�@͚��2� �ٮ�������%��w{�� [�҉/�=�^�Bs�0�
qM������N\INn'���t�=Ɂ�`3�Q����m)A�A m��	�I�w9>;Tީ�?|zq1̍��_�ТB�j
ЈN���H`h;��mw�@\ofz�n8t�S�D��[X�]Gܴf����ˢX�?�,Im�Z~�g�:}9\��M3��尚��6�Kr��V�Mǲ�1,�������b���=#������$xR�[�cW��55J��-7�p��V�І�m:N���|�F��7���/�g[�� ��9;TyA��G�"&��etJ�
ӻ�����/�䯄%|���oS�`m�����,3�"���������Ѧ���"'�P� lw��5�튬 ��UM���	���8�*����5"�PasF�msM����ȟ_e�U3�#�s�S�������!��'=�\'FH�V�� f���F:���s������k�%��E��ZWK�çQ�����H���r�K ��>���Tk|�ٚ��š)]��e��k�r ��֫8��AY�p��T�ް��$�p"}��y�٘����=�b��:��x�oP��M���0c���W�+�c�����eb7�A�	���?��,���r���t�yꅮ�b[݈��y�I���;H��.�)c�w�(�9�5��Bm�NP�)�=�)���V㳯/g:��$�x��G�>w.�ٙ��
�ȋC(�]�B*H�Wa>,��d�ѭ�f%"j`�\��?�^
����0�#S�p�1?w( �9L#Y��������$T2��[��1�`x�������
z�Z\�X-T\ʊ	෎��)"'��]O7�?����-t4�"M��"Y��>��w��B���OP���7���I����_ì&��s�6Cf��C�c��~�@����� ��bJ��R �l�6���6:��'�CR�1?qLv_2�%$4۪��Q�^��ݏ/!2���>�L��S5�r�R�S8Ll��p��L�]p}k�������Y�}���7m�z��4-�����F+��/ǵW�C�]��r��Vx�u��\ہ4ES���P��)	gI˝:@�}��B��8=a�$���3�T�e�Ȣ����s[B~��U�2U�	Y��"�c�w�Xp�n!�3���r�-�Q٢|&9J��V�i�x��^Xvc\x�i�"̖�v���%p��d�W�?Z���h��]��[�f02�z�ɠ9��,_��y�X@GD����M����,���~\�p�|r~d���vX3�y"M8�-�Vx
�3sbw7u�n�#�&�+c(^&�ݣEU�Q�l�b`�6�3�m����ɖ=�0�=��ȨM�zD-�l�P5��O��D��kΐ%[U��Nt^|S���z���4�5M'�y R��iRY�٤�L!,l��h:���������O�~k�I�	A���{��!�����L{)jO�]/��`�;h�q�Y�������6����qx�+�6Ή�[�z�Q�3����ڪ���	������"�ȧm� i/=^O�]���Ƀ�>�גf48�H��
<�$G)"O&φ�&Ǐ���xQ_���g���YU9O��!���:1{O�y�����1�ta���J�7���~02�$����PO:��y�94��x�	�5��s6Ӝ�\ܸ�K�:�Ýe��Ҳ�;bWe=0��4nТNz�ĝ��KH��9�)?� }����v�(�ѷf�t���%z}�TdhXO�d\�^բo�4wN]�k8HI#��x@�,�j���k�+��xu���0p�{4��R�=����.��܏ʊ��Ŭ$z?.�9�l��W�����%2I�v͠��~����"��8��B����}���G}K-��l
1�T��R��||�����:JW��)��I(���G�{���o����؍]6ƀ �p᫜�ً�`��m���g�V��7�lǝ*�=���_�pɲ�8�QT.d��
erY�/!,M;
�X���k��6t���������	Q���Bx0IZ��G�|�P�{]�u�a��yƅb��Bi�B}q|T���܌�߉�a��u/���J���s�K�H�*�]�/�,ż��KMɘ��:|��#�tn����Ơ���*�p:�)��j.QPk�#P���䆝]Դ��8��j��&;M�^d�dT��ه��bcВ���
�,R_d���r	����E�z=�l�����[��$n����dCȧ�h���_	0Y<%��ŧ�{Lݹ[�J���*�WQ��ZÿF�npT�|��I�q��%Y�s\z���.�rG�~��1�w̆��b�~	��⻢�0U�2�������7�����gy�6d���G��;��k�kL!��8~��'{��$�y��i����=�-�UM$���tǪ�ݤ ���Wn[���!VU8��r�f+�i#˫���gHgAM��c�Ң���b����+eƼ�uX~�ұ��)�n�:B���>��)��-[=iE��R�A����)l���Uv<�X����19'��ӱ�/��/X��G�㌌"(>�&�x"��13Z�p���q�vԕF6���4z�N_G�3p^,����"���Q
��.b�Amt�t��%��=��O0C��8�ԭ�&t���Z�H�
�gQf�AE�iҔ���gK'���q��O�=�#�^��5�<%����t?�X^�&���^ )���@Q�r�a�e��\��}ռ=�dl������4����R� %`�dMS\ 5;�-�z�(��ء���Y��梴���]�������U�)��6c��NB�^+��T�C�^�*���Q�~���/ sf8A�!]Y�L��v�:AM(�*˷.t�}ߏ5����� �� 0��o��G/4���m�����NA*�좐��zH]>��E��;$��qt�� ����e~ȷ+W�A�-���T�B1�JN���-k2�ۗ�N��|���{nd�IX��*4��m�/��`����c%{+׎�|�h��Y���k�$��BG��K�%i)L+�^7��E��-��.�j���fk>��c��հ��T�c+4���;�v�8ү�*։�w���{G���藃P�K�A�����y��sh8%�l��u�4<�R��*��^"�xªbi�dZ��� ��HQQ��u�	�Ū�$>Ɍ���aE�U�O�8���n�`NZ&M�� ���AXƀ�8�\>�V(�Qj��.�R�I�u�[���x��m�+.�(���o�,���{��u��}8�v����*�SGR.f\:�!�_o�Lu��"mZ|��;��+&���~ַ��רa:�X�C���OL�W�2}V�lU��D�GA2�ގ"H
�cїˀHP�8�*
�݌��f��M�L2����0��v"*�s���;�k!���'�8�M�	c�r�ӹ�uW��ڮ�)4�Y�˙�Lc7�!K��W�.�h�_K8�{筢E4)�J/�ѩY����j��j��3Gh� )~&^���K�x��{~�C�M����q�%X��(nH��=9�O�XFRf��/¯ �9]`Y����"-2�������CvX�J����5NJ5�][e���`4}�	�J��+���9u���C�39w���P�������ț�B�rXM�+#�|��4H{�zF �.G��˵(�(R�����fz;�J��A+�
!w��Ebt %>�s���sad{3�T���y��#�0���N�$����j�<m��#Zy|c�R�P5�����5J#N7c�@�K�ܙ.�%�����p��U���� ���衅Ə��ԫ+uQ����V=$��q/Gn�S�/���p�_��*�P�8Y���?�R(���������ϻ�@ �2\/�L�6(I
���,�{��}L�QH����g����!A9��
�k�6�K}�Y��;�7�*���p���H	2�n�}%~\L���J򳇭Y����p��<�9#�� �%rb��o��7��{��8������N5vp��Ak��}�F����sݲ��J�+����ٕ�p��
�M�V�%r�Lɽ-!���������Q��i�T@]�0x�]�i1]�[\)�?=�֊EH���{רj���B-r���.���^����������V��r�'�_o>��8WVY7�#?����X���f�e|��v�3����
�_�B���);�<�/�!�A)=[�U�V0������қ��l�S�(Z��Pm�e��8Hgn�G��2�����h���d5�f;]��NQ���1��;^�������i5G �����;��o&~K�6�Q"k#�+8В�}v�#w�ȼ�[� ��������6\��,��"���p	2\=���Aތ�tG�c[R~�r��}C�_�4Ht�@*�W�U�cy��7(������T��F��r=�ԇ�b����,�յhj��ˇ��u3���B�J6��a����m����Ö�@f�ts�/�y�i�{�)�R�L$hJ��x2۩������ Z���|�,���"S�[�-�d4/�����x����0�V��|uE�f�3�����5��v��`n�l��9kh��x��-&'֜IY�_%xNqD�'�:��˒��� ��ݗbw��~w�?���y3,[ͳ����nj�s[�- �f䪑'�	!����,�����i��W���F��>(�5��m��ہ9�b�������BeNyV�2�n��=s���N��a�r�/�̽��] *n�K�-��d����%N&�R�{p[3b�;0�e�w-C(���Ǿ���t��H�J�5��)�k��j�D�}|���aꔜ��&b:����9�Dd��#�\�L�o9���. "��Y4{)/������dm��	�>��Z ],G ����O��X�yR?�`�rh������h7��q3��Ꜷ٘��+F�:$g��G!����y
n�=�a4D�$֕�yЁ����ۤ����b?T��0=8�I�p�J�ZsةpY� 'U���tvD估�h�<���ma�h7�e�䇀0�������R}�El��	�"�ܓ�:n�2�H�����t��i�F��J�d2_�_�%�����8��җ��e�֚ �N��f8K��2����L���#��輑�U���W~��[U���)vu�9J��P�ju�i��ŧR�p�u���R��n� \�H�K?������F�`���ZBOL�V�T�a�"E�s&�P>`zη%��R6�[���64z�{X�a \����ƽ^@����1G.��R_a�lm,:��T���L�W�#�vg�N��!lD����o�@5t9B؂N���	�| :k�^e�MqM�t~���g�o�A멫������k��~�� @k�9V��s,z��yҊh�Rt*@`|���Ğ�x%�
���ӅvkOEDd�N�Y�.�潸���j�h�]�7J�Ay�������mH �@dD��<`�7{�)ڀ&w�ɲ�ܒ�oI��&�� ��i��N�Ӑq�^ʽ�%I*�9�,�
��xM�d9mkr�}_��f��2��^=3:4��?��
g��qt��ׇ����%���]^
�0@��ž�4���4p-��7+�z�%)����8��X���3Bi\ˎ ��.*�%}�OH����]����Eu$i��/P������ug���[�gj�n��A;���B�ݕ������	*��0hY}j��r�~�I<�z����M�( Z����ӓ`.$iс�U�o9�^\?�U���[wN��q�7�mˆ1�Bs;xƼ�E�L��	]��@(�ћ:�B8RY�8P����2�[߉��D�5�J.��tJ"	��n�yF�G�(�ӊT����)%�'��u�'̺|O��qN�j��銘��o�qG����	�tzα	L�&\��,{�[�1��C�������eo�Q<���G��4�!6(�ՊC�5�s�'�+�I��>���?n�}@���ܧ8�]��a����
&Ʈ�'�������XT���`3"-4���\vF�T��Q(�Ѷ ���;�L
ǥ�l�vIh�j����5�Y �~��~�'��Y��E���v�M��ok�JV��-[$���,KGR�N6|�g��c���7��d_�c�{s����3_�3|��BJ�+�d��IU}q8�W8x�;�C��j��6wR����W"K`�W��+� �G�4��M]��Cwp+m��/�t�A��U#��of��7}�0�'rC 
�N?�m�()�Ç-����s[�B۷� ӳT�ޣ�N�:f�b�{��H�(��\�.�%����Bp���&M�)�;D�q"'�� ��T��I�V��i���g{��d�N�e�X�P�:~��
!�Z�q.��������PkNM�d��u�6��@�$�8�#�=��N�N�?�ܺGŤ�Ԍ\���d/�ȴ1X~�+���P�H��\u1��G/��|�kpC
�@b܏ldn���ԏ�Ïj��=�3UMr@��@�������$Oj�IE�T�������v/bF9��Of�nP=;4�����PW����u��b�c��]�i^�/��={�#o�K�?��F"�
��\$�C��$�r�� ��.G�C0�d�`�P�ypc�9Ŀ�_y��}�����z.����i�zO�Kb����P��p~�񺼄�o|�Us���9�d����e�F�9ڠ\F������b9�<�2>i0��bC�eRE�v�C�*lN6��%8p��-�ا�q��c��B�0<]��r_�+�:z- �Q(�}��@w��DF��j�_:5��M��kƘY6��)�J̊�oo���������)�h�Kt񢜺A˒�a�i�2����:�1� ���>��z,�a6e�9��.;��S\x7;[��a�N����c�nj/�lAB��>��*����p�}EP���6)v[��"� ��@�F�����ІS�ZT�÷{;G�r����,2�h�{�e�8Һu	�G��Q�[�GU�v�� 5�*�b�iSIEH7����I���Ƭd/��U�L��ה���(�~3&�"+ND-�K��̓�9Z$���st�׳��y��?����R��8k�L5,A"�=`cX��{I���o���Y�I!����f �^���\��;w� [�z�~p)���Lۓ�J.�	Հ�����ɂ:����^��r\JOJ2,g?�\%�2y�V�V�Pe�o�ɿ�	�V+Z���&vT�]����ȿǢ,-ͽf�v�6��:Ԙ#�L����̰��"z*q%ւ�Oٵj�!>�]g
�SQ�-��	m�@^�Ȕ����?�◑,!�Ӻ��2SOwX��G"k�$D�i@`��I�d�f�mT�Y\uST��'�	���{�n�!:nn��E��I������uϭ����ӏ:d���j�Dð�$�1��F�LG����pN��p)pH��J�,۶2��/������g4�ڶ%A�v8�}����:�j�8�0?�m��S[ֶQ�Z�mp'��y��|�Ŝu�dO�މ�I9Ƈ�Y0O�Μ+p�)��1`�l��8�%Q�����:�Po��R���O�lJKd��V�%�CKn,�p-^*Q�7O���4Hs��$��~n�:/t�qo@�{����H[7�(�4*:s�홼�|�
=�p�Go��S���@��������!KJpM��%��e 6�XA�G��E�?r��E�&@����m�-�>�f
dmr�TƚX�;��?��hD�|��^�<\U�����i�ץ6�.�p .� w䍖���)�Ƅf����õFa+wMԓ��x�$:��ד�a��r{�M�	ֱ-��F������ωۖ���^:��zY�S��~)q���5GQ������{�x�SH��N�)����|�Nz���TAf�8��~V�~q��
Q�MCwR����oHYk�sM��O�����[�e�W����z\�Ȧe(��в4a��қ6�� 'e~H����+s�����2�ʬmT�uM�=�Mpx���!q׿�e7���- O�M�{�W F��o����@�
"����7�4B�{�[v��.9��s޻>8�����̖^O��}=���Hˑgc&g�����C�8�k�X}�PEg�䗎:�?P�P�e�6������^_�{�j2��w���2)�:�ѧu���g$�w���¨�0��0���DvO��ޞI��JDDne׃�7��i������pw��,�X�'i��kULϤF�]7��~���Ϡ������1����^����d���h�y����4֟����|����;�s�	9a�td��ĵU�ͼ�"Y���萆l.��A�<����K������q�æQ���+��w8�F��|Ul?�U�RH�u�Q{�p���� c{{�P�Q�g~�>0��`ދ�����L�8#yUb���1������Y'R(R����,�Ȋ�ㇱJ�[el�,\V���5F�A���.�@/r=p'k�1G�$�Ab���Qp90�����9ѯ:�'��'�.��՞ANޘ�����QK���uc���؛�jg����I6�@��c`��KI���t�q�Y9
����h#�����Xtw����4246t�0��o���6�������hAU>s,t�_d>���vd�`e	|��%����_s�v�]{V�`W#�-��/Ir4�ak{5\��#;����Zl�y���dXM}'ޕ���GN�ĸ;�{r:�zR�z�*������g�Y$�k�(.i��:#-�	��#Rש�}r�9�x�-��zʀ_��G!$�g�t]���_��Z+-�z�V��?~]�m���#C���g�mr�O���[	�4[ڞ�(��Ů7h�'+�4�k��g+(.�����	L���IЂ� ��n�nv<h�qڿ���,&0��`��F��˾\0>}�m�佑 �R�9{ClG����=I����)�!�Qm���<l��^H>�}�ʏ�K�ifv�J�'Y�ܰ����r��K���X�z��b�{��8�:����n�1�v�����֐bdkƋ*Z��n�$Q6�K4���f��C��;+��c��jw���o%cE���M
Z��V��C�9�d*��&�u����Tu*��V2���V�T� ��W=�mN��<�5��*��P n^#���b�e�Bm*�)�g�c^�L`��<�q�r0��9��k����Ώ�U��5�Ƞ�8�3��u�kb�4v����ī��'و��J��!��	�����u��td���=�|f@R����f�ӥA|�L�>�,���z���e��-�[;ae��d�N���P�&�o��@����mG�e���w��8Sn�g�o��^f���r����/����.۞wN�+�1	��5�#�ie��!�<U-��m/7�D?�G�nSBH<��YkCe�k�6�\�����(EH���� $rV�ZGCY#/���y��E2E1�&>���I
[ �(��/��h�R�Qԙ%���r�lZ����x,�YܤK��6��P���V� k����[)�"C�55����⇀V� ���G�1�;�R?wE�^���n��>r4�� "4$��He� �A��(���_u
�F!";���ǃ��Mzۼ}y�T�*fX��y*=7���o� ���1����Y�P�Yx�:���0�K�I��ܐV�bb��5/6 �	D�V�Y���jd�N��BD������8�@$��px; ��ϐ�w�Avs8���~�I�Jp�n ��fxxc��-���~\0�9����\��c4	Qu�x�\�	�ߡ��2K�3��x\���$�l�*����3Z��ӓst��"�����
\�/#ĝ��>�A�e�w ��wsne�I��ֻc�<
W4&��5�ޏ�=^�3I��rCB�G9S�&?�=�R��:�.y�R�/�K��B��o���u��F���L�K������~�v\���^�r(�����JX�A�b��1��c��7NZ��Ѯ�S����(������FutZ�W'R����V�߂3%���_|T�͕�STвI$C�Q՛���ָL\D#���c����)�<�	ż��*T�k
��!+���ﰘ����*=Ѹ��Z�%���1�5�WΌL��s�����/h�6Lt����c����Pʑ�Ow�wF����@�V1<�2�P�fx)��5�� {pu�8i�q��U0߻O��F���n���$��e�[%��������WZ�V���}W!Fox^N�W�qK��~:�����
������^v�����H�:2�J<��Dy�����pe{��gy�2��"������y�CriU�\;E�qo�0(pEY��iA�ݺ�X����*��=E���GW�=�aA�{O4���B�<ntބl�l����y�s�(�q1���&��d!�j�j��ـ���Jp�M�`� �a؅����҈���KW�*�H�\�`]śȓ!ͅz��x���D�ox�(B�&����Q	��K�%t����s#�-����W�~R�l�����8,�-�3�/q����6ٹ��<����%�z�����7D���K�^o�䗰dw�4�z�|�g�R8x���]F�c�+�`��ug>J|��p���謫-�����t�H�.!��*l^�x�X�']��-S��w{c�d�%�EG�@>G]�r$�
f��5����#t�B%t���2���T���ϮL8EwAp-e�'����t.��4{� h���:լ��k���ݩ�qW1:|z3�0�i8<~`�\*g3��ݐ󈑉��
"Ԫ���:�c�$�G}��_�F�'�Ӑ"�I Y�+�ո����a5�Cy���k{�8�KCL�$x�`!#��&�E�c���� @��}@�=D���A*3�� 2,����I��-{�NK��3*e5�t������/!��ƙ��ft��}����R�8�J%�k6s�ff���"�)�a+p�u�F� +�C��dԬˍ�4�`\�C`R�[ėd��4��
O��E�\n�
��%�����H����j{/��	R�ÚRxE�
��B|d����;�8\۩��S�.�F 5��}R��Ʀ8�&�>eҳA����VV�k�!�����F���0������w�)C�?P���!�w��mQ]e�:��7����qF��ʳ�V�b��1���shPԶ��,~K�Q�,f�_mI�n�2�����(+�q*&��]ϻ4���u�\�B{��mJ�����*<�W "g�i�����k�̂E6n�W�zݸ�]��a�@������e_�*��[���T�q���&�+�~P��3��A�K>u�UC�P������)���t�H�4v�|%i�S�V��b9?��ya[
%=�]D�����뀜��$�k ���渉
'1"�"�&�b�@�5�.���yCW��AZQ�G�xY�
8���⺝��B 2�Gյ]C~��[Y�I�E�=�Gܸ��]�yӽ�Y[� p�S�>ǳ�(ۀ�W;�͏<�w��i���bԈ3>ʔ��Mm�t!��F*��G%��˝�#���ć�IcH&!�9��۠Ox���y��l�@����Qu
g��D)���$f�������h2�<��F���m��9�����A/���.{�K�>Q���ֳ=}����xQ�S�?�sy���6F���j"�'Xr�h8rm���?P���n����m�R�X1�~K��A��-l:U��V�x���1�}l` n�=�B*K��]h��ECɮ/�*�jwK����a!�¬�x���b��Au�4�A-�o��ę9�q��|G���a����ZJE���w�2A6e�Ҍ%���-H'�`f]�yݭӧ_��(s�:A|}�p(�>A+3�YD�&ޗA�N�4*F��JEP�Sb�|7SZėߨ��E��J��5�Զ�;��OHm�v�W���'�.O�X u󎕽�jkǡL��f��X�N�
��i�
�	A����X��@
D�"2y���hr��~-ֲ�}��/=d��މ�uw��O��Z�NVssQ����RsIDˈ�3S�k�)�_�`���a�^]?�1�n�3;���K[i���`�8�j��[�J��A��>���z*�G���%�C-��F����`_/�r��M����3C<��׶:i�'�A����BA��0>0�*�Fߞr�sD�
�k9�}�3�|TM]����?����F#�f|b��j7́��c$Аb�6��E�E���Z�3b��E��:�,�Uxz�V��)L~�=�]�Ѵ�w��\��E��t$�89ҪT��;ա��b:�5�J�)��m�s����*�0��Q
V' @d�DSY��aqU�{�He��NW����O�����1>�i�y)x�-P���2��.,*ByFW�%��`�����B%��HF��f8�����"dI]h&1u�(���˵�BQab�b׍^-Y��.,�)�O&3�]"/�Œ�`�c����4FL���kݻ�cu��,����I�Oxcƙ,�5�L�o�ǯ���o	�m�֕��t�)�3
̪bv��qo��M���d��H��%�*��?'���X�q@��'�gfO�
FW��t���Vi��٧�t|��.3���7��a�3-��j�D��Z�\:=i���>* rs���D�##�A�}���")E7V��K���%��v��P�l\�������R�t. k͜�)[������$�,|��]�@j��l�7�YI@���2���/�p&v�d�,������"��-ʹ���W��a�z�:�)�B6%��5)��_����� v������C�����N��2br(2>		_wV�Vt�Ds�3��.�/R{{s�b�kZّ��[��	D�BPR�l2� b������zMe�Ùe�>�y���i�����PRv�T�q����k��=M���Ԡ}P�l���L�П !Gv��`�;���v�\�6��)�#��\�*��S� ��E>��j���`O�����]�ٓ�z��<�$����Bb�HQ)�}+w=�"�?z�^����]J�Z1M"]h���/k���ţ�����8�Pw*ͼ^�8}��ا�N�b(��!��5�rm��1Ny��J�K%H��l{��Q�E͗Ҭ~�����(�!�fRʋ��Mq!�<���~��+� ��ތUWD�fR�ސi݋�����%�z�B��c7�`}DN�e�-8���|
��ŌP�3���`�m����N)��K����I�_�r�\����H�&y�^��{�����uA��|vh�)�1��Ǭ9��S��:�'��&����g��_�2���x
bQG6evc�[E�ǥ17QDTqi}��#6霥ݖ�l��v�y&J#K��E ޺��9��m^ܝ$1:��R��O4�R�1�Yf�I)�,�l-��	���ϡc��ڴ�[W�Fp�	���Տ�E��Uj�g��-�
��'�M�����I�L�|V��E����M�,���\��8F��'�8��$!�վ6.UKN'i/>g/z�h���2/�ۉ��yN3H�Eh�lԙ�0�1L���9���1��Nc�����L\�Հ����<R����c �cu��3�1h8����s�{�S���*��pf��2C���yO~�n�"�}v��yKV�ۆ�	`����εS2?~�C��]�N��P����+�����l�����k`�Ņ�zvy@�I}�;@+ˈ�h�=�!,p�Ծ>_�S$E�B���g�n^x2�7�,Z������.��� aA�/��8�5�{��Z�s�����������G���}���ZFGzgg�}�x�lMޛ���u����A]cFw�����z+4�?Gv����q�-�3�\�Ĉ4��}f��pW���5��Ϳ��]��ŋ���_3,ҵOfh�sgBV�	�y]S^��+)�̙cr�~;x���K�|Y9��s�	�=�E��uQ��n�&#�z����P���5�i��>����^��9^�î���*zR,�iv���Oކ�QSƝ��՟+�WL'�
��{/�f�Q�˪k�#��R\���5�8eS���I�m�)���tM0�B��[���B���WЕ�����&�\��Ch��H��^�7���k���k��B�v],����l$���y
��X���8}���XX4�P��o\�Yi�V�#	�<�?���#�WUk���0Ը?�������bM�o��[m!X�Yv5݀]i.S��/y�`�S�J#��R"�2�5���
��.�oi��K���i���l�~n�B_u=��
���:\z�#�K-���K(��\a���2��G* ��-�b��� ���U�5)G�a���t8D;q�?��Hos�\h�6��S|>K��R�ҮF>�ɢ,$���T��u���ڃ�iӽ�:r�v�q��3è{����RǑ�9̞�iG���O����f췶"���Ij{���(�F�8�r����H&�0���B�Q��RM�b
5aO�v�(x⹧8&l3 ,�J��SDT�R�9."e�Ab2{��<���v��W.ų@�9�wg��4���Vp���\�YN�~���ؙ#"R�c���$96�l�������0 ���j]���^�����G�]5u���8�����G���[�mTo��|��2�n�55�>�5"�t�I�O�孈��,�<m�Wvz���*�_fe�x�O�E�ZxegM�����2���%���2�"w�����`�IV�� ����=@���ǄyeL���C�|��"+�ۯ�/��$3�;bt�`���U���(��Np���wde7��,M��X��h�gt���_�x��K�0%���~'ֱ�ԡ2-͸;�˘j���|y�\wst�2����q���([�қ����MFq��T��t�T���_��Ad�!��аzE��G�V��ⶲ�M��
��ӐҺ���m[R�'�o��ᩝ(Y���1��5�k�8�6۞�5}�!�m������m`�_^4��澓���k���YA�(u�q2���"�J�t���]F���v���>oJLt�Q���2t04��m��cʣQ@�e̝�s1�`^�4�Ѹu!n~D U��_R]��}���C�B��$>G)�1(�����y��Vj2')b����!��>���p<�wg �9U�9O�L�m�����{>S��ܞ��C˕
ύi�].|p��&��Ɩ����&},|����ҩqm�#<�]%��ťz�1wnW��=~��v���������ʏ���Խ���*�aE�|��-������c��?a��Pp�"�!�s��Ƶd_:�+�l�j�$����XZh������M��)�޴'cW���NU��ZFewi�Al�����*��\؏��Aabpd�w3O�4��y�|O�1s���^���F%��m��
R�n?h�R��L��%�ڵ��ߝ�d����������?�A
A���Py�`�_��A��RJ}a��OY�F<�~��QH��g��&C\���Etw��k:,0�xl��1����ܨ�C����'��X�Hf{�֙����A��I�/�^�A�B�;��(��v���n�P�ʼ=�J��w�d?|���� ��H��"��c��#�����9�<��-F�gJd4��"��@��Jr�l�A�y��q{�s���-eQ�"`v��0gJ[ݬH�Iї.���s2�&����w"�G��OR��*WƑ���qzv�7��z/_h�W�h/��*� ie�l�@� {�FZQto�D������Xw��<#���Q�Ӧ�foҬ,K;��Ĺ]L�-���߳V��Mw�����[N����P(W+���ċ��d����
d��UO�->�R�3V�!��+��|��	�~��<]�@"oW�),�e^���ڃ�.��%�ZX��A(ca���[�&�<?,#�ᭂ"p�R���H�8^�CG�5;:k�8�)�����a��{5? D|��{<��pÛtf�O�1T*����#QanJ9/��B�cF�?���sWZ@ց��G(Sz1��'7��Q�=��6��@q�7*�UH��
�g���r^��A�g��zH�x�	����2�֒�� ��H��H'���P��w��M(�/O-��H��%�V�lsփ����G��Q�ʠ��$�<:<��ٱ1�d}�K����w968��)������]ʁݍ��>�I���	<u~�p�>�Z̐������jf������U A������S9C�}����ئ���R�!����ۋcs��@�i����D�d��e�iC�ib}bO% �cR<��Z��*�;m#FP�4R�?����<]s?�~�u����壟R�rM)b̰M���	�J���\�j�G}q����ȑ����ȓ�,,�a�r�1�̼A�������a( ��m�RG���g��!��cr�Q?rKu���M08]@��&�ȟ;s5���ޕq8�Iн}It��0�<HB/b"%ߌj�;���1�����>u�*�_d���4w�^���Zۣ�C�K"	j�dU5����Q�GĜ�.�|"=?B� ߶p~��C��$�������b���}թ� 9j��|��O?�5��5���=e��,`����Z���RMzi��y&��4O�D���������7�	��Lد"���FwS�r4��?��a /E%#B�$�J��	*E�~&_���y��8�mx�KٍxL�WG�����n ���W����?�Z.�����`U��PI4���Ռ�:>�Q��h������bI���z�ܡ�B0��S����'��,��jWM>$k���8G1����k{��m � xn�þ+�-�_�ScqU�����WR�x��~-�A�xp}�����~�La��`�̨�ӱZ���g�fY��Z�	�����r뢪��U�?p��������d۩�8��F���f�ă}٢�J�OĊ��� \P:�Ԉ4(*��Ӽ��w?�Iևe����>fpm�q����編9]��#q~��e(�~�&���x	eq&�:0�#��<���<�Jb�&y��^F4��]�Ƌ�����B��v�1fNB�>�[s-:�4�T|�t��-l`7����f�Rz� ��k��KŜ��宐y���+��圬0
�g/�e|E�
�q]b13�4,,�Y�����,a��/{Hp1`����ħ���t`P7����}V]6���ʄ���K�����z���:��Ar�N��%��,�Oq�t�^���.enVq�ޮ�;�C'qo
軇�	�_��wL�B������~y�^�ɲ'j�}*Ɲ�Q�=�����!���Z�Gr��u���$��*%:�b\��~1��L���~����x΃|i�ⶀ��@�gij!i?q�
2� �����̄��쌝`�2��*���M�|�+�r�	�ii�����o����bwl'.!I�]��I��}m�����fٟ�"�|�O�z$��;8��m�a�D�f��s9I$�>�*B<-��'_D�p��!cs.8�/�*`o��D���-��D"����/���W&���3�پ�A䋆u�w���a/�D�oYY ^�Q�������?��61n�{�%�K���N��j�%������q� �ۖ2o H͚ň�qD�騑�֢��e���6���XEU�5 ��Ϭr�䷑�-m�� � ݆:.��A#m>bݳZ��^`zM���	P��Q�@�����~#|�H�Cw)o�m(�]���p���q�qSli`��)iNVF����=�3�<Ǜx���:��,Ӌ�F�B �XnSTr-����J��g�Y.(I���8�P��cOkֻ�dt``�%��D!Z?S�Q߼v�Q�����t���"tu��ܣ�$4�QJ:����>gF@��ᵩ�.���w�=
ɯ�Ĉ�;�pE23q�&T�]>��Yy�F�N�jlD�٥�}�H��N�{U��<ka�y���C��Nx�`iܼL�E��4֯k"�9N��[�O�{�7s�%���~��7C�w�J����0�=-��_[kJ���ԮO���}Eb!l�	W�}��i�(A�*>�]=�N�E ]�[H)���t\-��������,	Csy��LV^�M/<`�SB���޴s�<�p ����FX��@(����D��|U��O���F��������i=d�9��Y�2k4�,dq���34��?���[�*؎f� �V��qQ�}������ @j���[�q�Xw85���s�*��Ph�qK��Rr���BJ2i��$F���g���[�=�	�X�U��j�+�ա��,�i��8o���"�ӳǤ����b�4O�ko�}X�>a����$���'�q��N.�L���u�T��+f���%�)�m%O���͂g��n[4zjo#��������}�9��BZY�g8����k��Ȩ��e�]�'
����p�����&��*�����A;����אgA��� ��kA�c�1����L%?����O���_lck�wj�E�rQ���U��w�`����T����Gn�x�k-�R{��UZi�lD� �/�>ˏ�<�{4��hu��/Ꮙ^@�t�")���Ց:#����nlcN���E�~%*(��"�:1
��hw^?`7L�C���ngP�9g�F�L��>�vs�)9�L��iB��x�i�,M_ɖ�>���V���*a�dH3�pB�b�Τ�v�M�{�;��ۢ>hz,i	� �Ş[���g�������
�SA�7�҅�#���/��1������s����{Z�˲��n�ERC�MqS��̃5�U'�	�Q7�~��e���K2W�Ȼ���){���Xv�˟T�[��L��������}<��DY�ʟh�@[��
#j���-I���e��O�y"��Җ��Ԭ��?�����aNܠ�9"��L��!|��:E���삭���_�)��a�i���P ��)W��:�:��c	jDya�x�����F�:ڟ���'-򰃶�cZ}�z�'Yq8=�z�҂�������]>���ڛ��RH��Di�N���C�y�aBki��N�~P�y^2���H��
�t�U?j=ibT�ѲV�GF�܍DM{��Îp�y��)��R4�Kʂ�ˮ�-�I:Ȁ6�����A7���u��T Zށ�V.��U��7ŰF�;{�YH��;����3��;L�m맪�mi|��3��|*g�9[tv�]}�`�sIɃT��@??[-�'�V�N�@8��I�'t+� %�/w��K�E�*�|di�lHTP����	�9ʊI\  L	�`�4���� �Ы�Ĭ�	K=/�B2�ԽہM�[��Zn@Gp�D�A�c4�L�e�?�[�D6�P�N�o��{E
ɽ���0á${�Ê?/��6���r��B�'�X'"����}"�e3���ˆt.��>����h���+2�p� `GV�@V�;��|k헀�8���>B��I��H��ꥺ�%�AC۾�0��#�#�2�'+�!��O<A�6�$^�7�9B.u�8�l_��
Lj%ڳ>��epX��vJ���;52�5����>�Ԭ�P�4�fmI�P�׉���D�:sE� �R"�nU[����*V�d*��Fz<�	�F��7�a��kF?*k`%��l��Z��:s�����V&�>�La5m���gr/� [?C���pttü�j��#��W�mO�~���7�Muj�ݒs��B~��tD3�V�\�+��?�~H��L[�J��>�w��x���s`H�t��&T�!�+�ĐT u]��a>���pъ�� =�t�m\'�7��p�QR"��٠�����o����[�]@��x��s�Ƀ?�S����J��Sa����L(��2��Wm��Y���!>���Z�L���ŉx���;����q��`����s�F���Q��!C��GWE��;�Ç��f�])zx�����˫�y�.��l&�:m|�8e��]k�,IQNʆ���ƻ�KϞ6��Q���81mg���o�}���qP7h_���$�}�ml�(�~�#f�fW�Ȭ�ٰ��Ha�����3�e�+z���!�2F��s|n&�������{w�v�G���g5gg`u��'�'*��B\���8����`}2NB&m0ΞK��=P����"/`�{N��������0��].����E ��%U��� ߈�y:`�ZŹ+�E�����Q��S!�	JT��;Н�(���a���آ�~U{�P�qaݰ��9�gu�;�j܌�ģ|��	��P[E���,FT�$5��_-V��K:�zl  �5�p�d�8��-�
�6t�D0֓�&Э�
�_�M?7-�h'��� �+O�<.|[��B]C�q()5~���m-�|���ϖqɘ�1�Ӳ�5-m~nR����f_Ӹ˖�7:1�Z��ܟ��\
��9�E��_:���7\:FDbv�Î�Vv������O���C�c*e�/&h�cJ�Q!�nXnb�4���u�S-ɨ��x˴x"A��
Zp�E+A#�
�Y# �%�������b��Z_�ɬ7��#��z��d�~2�L/ޯ��S�T��sM�l+�&��P"Z�m��I�p������ǈZ�T���E˞����4�z�)2�r�S��|��/n��{�#��d�Wg/0����s�<�*i�I�b�6Vʍ 7���# ��,���$v
��hD��A��;���/1��l���mʎ�Ub����]^�Ѡ�z�IMA�po�5}e��n�}jɷ[.Eo��y��}����L�~=����-�U{����7��"F���
��pF�V���uWp��)�țqyZK6{��P����e4{e*�8
xHy�[�lV��0�:�����Y)B&�Ke[z� �@�7QB�l��|�8�{�
�ۋ*f�,j#'3J-[JE��6Z߾*dE�����+���k�PƊ�����6Ȇ1;3k=�K���?��f�����9Hye��G�[�81��4>ĒX��@�a�*:�� �'��*1�7]s盜T�K'!Z�n#&M!�]!wVLH�YBf��ݔ%ɨ
s��k1�8�&K����r�ihyjr�eչ��B����Kc+�t��#��Z���w�������]k`�U�8��
c+�3��J�TYӅ'�O�[�hàff?f�$w�"��]�&�&D�!�	����>2�nc�6�T�gh���e��瘀��5�&��T!mvJp�����|�y�@/�*sU�`��W�Cς8�Ba�!�z&�I7g9��[1|��$������/�jo&8�'
��uE�Di`ANܲc�XO�^���٨�u+H�����^:��B}��r�<E��꠰����H�I�	�w�n�� �D��i"�(H"�T��"m8�_�~��]�5�kӔ������� �^3٠��sMV3q�(k>��7�]
��8m��۔�I"�@ԭ��;���bX3avľ�e�[zv'�b��\:c1o��u�wT���>����!=W*��f1�G�#7`^�&��12�#��@e<�8�>�B�b��d���7v�)�2O؈q�O�����"��ߙ�;_�ȇ���'�� M�����Ueِ��H�z���:ڣ�������%XVa6�|]�U���v	��(
n�z�n3�,?j˦���a�������oceq���<�o-d��k��Jv�]�胐	��<9�*Ҏ:��:�J�A-����^T7�MK��f<�٣`%��u	Υ��D�Gl��|����Z����	�hDb��'Iz�C��IC"��9c>6V�+>�]� �?a�9#ܮ����zBݥQ~a��݈ZI��
"�Ѐ�Y�:=�_DL	o�By�O
;������J���)f�V$��6w�[�M���>} ہf�N�����tm �Ʊ��p#���ׁ�!IpQpy�|���־�a�`(�H�9$6P���Y��������/?<cJ�QSh���b�$	ܵ@�ud��2>�~,�K�5�n�;8���a�#�������&�];.�	���o�@:���x0>��!��X���*}�	���m����t6)+��p�������#��r��k�<�)���( �J>����(�.c�Zه&[��o�M<�=�Ó�b���c�������6�6���H�Y�j�u!R?�e�6�KzWW�;���ȣ��h�a�.B� �9G�υo}��M4�<�7�X���kُ*�ajj<o�{]4�#Ӭ��<-=�XY?��'FbT����Y��;��Xٻ��J�q�;�cB*���)*��8�RS�5�6�Y=��l�G�H'���c��{�4����/ƟE���S4伩(2��1̋@`*aE��d���Y�ʇk�i���o�`Ŕ��\DP���A���Z��vm�M������J,�5obg�F��Sr��ޭb�=/uO�(�g|�HWT�ڦlNk=�{�����"�<��)e�W��s�7!s��))vq���030B��8?e�o^u��|{���z"p��K^�~�e:�6��묮0�q�ڀ֊���=c̭Z`w���m����'�rC���A��R�bz�
�G�da,̮���L�HGk�@����]�j/
Q��m<2l������q`���꓌��Tю��B�c.�_x����j~�ҩ�� ��l�ߍ+�p�X�_�/ʑys�*�lܞh�Q���zn�����
���¶YX�(���1G���;�i}J��(v�b>�`��u���^M��/�I�uj���e#"�H�S���w8m%D�Og��Ĳռ�{����nV�SMLM1Ю�f��|.P�ؐ�d�XuH�p�:7gj���n������C'С��ڟ]=+�LDy7���r�D�v[ۂ�M�Uc��/�$"Q4-\ܲ�9)N��C��(�$��5��s%9��}�uq�>c�î}��T�l��v��<��U%�G�bZ��݇xkCh�:$s� 4#��Fq��#݉��N������a�n��'i��~U����d���?�Λ	�-66��u,�եUT�}Tn���8�"HOڮ�6K�!��Y�7������#K�k�FZ9P�X:�����B��������4����s#<_2ځ��z-���!{V/��!�|�sl���	�LoD�Ӎ�����f�����@Cz����{�Z���m)��W�Ur/acO|A#s�4e%�c:;����F�~K�K��PE����_���|׃�%�'�!D�����>Θ��?�lA0>Xm=t�J��k�;����J{�oQ>��Z����rF5�tV�������(������d��5����l��R+�g����f(�h���
�y��s#��vU��᧡\N�)l�{֩������տ��O&,��u��s7��K�c@��#�"[�Ɨ����h�ͱko\H�.�ρtR�\^ﱀ�9{-�u(޸-�X�نI��X�0����q
���P�S�۶	�ńw#hG%�P��̇��.r{�nZg)��h�So|��L��<.-��pX����y�1��2���	�*%��n�?Ъ}o⍦3+$84���{*I�x�$�J���s�q�sZE@;��0�'!��z�F�f�\ĠZ�! ��������C�4�����߳����$�s%��Ni;��
^%�8�ֹ~Io��{��y
:�S3�!�Lu )Ԩ���£���� �0��Z՟p���Q�<aG�gtG����r���:��K^+����hH�\����N�ZN#%<�e>J�<��e�r�~�vQ�#``���Y��Y����ޫ7}�Z~ �Є��?�J��V�r8cRI��Q�� Q�jj���7�W��;`a,�����_���umمv�6#~�܏�Yc�1R�Q��
���K�͙��&�>�-���
��vS_�L��X�k�+��B&������j:�U�:~����G��� �n�!�L[�@����}\����1�j�i�����Ԥ=�[��Lˌ�V��nM�gx���.G{z�u��Q0�X��%Wd$V�&��et]��H�P!�����P�Y�p��:Ê r�����7\p1��͓���O���s�Q��DB�}��l�N{���X�,��7�R+��LB=!�"�.\W@������5�*ʰ�i:y�E�i��2/F��{V��vb��#��QN�¦� 5i\�7�h�����b�xj�64�5X�u��ZS4f0���7:~dn�9-�ԃ	��C.�D�<Qi��$�XK|��o�	<E���N��J�3�#;H�ץ�dx9�S�꡹�[��1L�8�g���l�>G�o�����2�Z�z*<�7�YO�S-$c+χk.U�����A�%�O/��8ɡ��a�s���������Ϩ]������c#�1��H��D�y�`��q^W�"!�pME֭�ƚ�Ҍ�n1�3��+��7̙D�&����;8�!CK��ɶ��o��v��d

K9a�����n�h˄_��~��`��侧Oy{��=�2T��D��io[�@Ӟ├$@�x��Μ�`���<��[����6}<�s�����d�2����Ǔj6"+M�T͍�s�d��)��X,S�c�/��ݫgfDv��G�ῼ<���g����Փ��p�����DE�V<�U�k�y�/����U���o�,_ӪY/8w	,b����i$�fb�Rbh������C�����x�F�:5���P��N�Ok��� uGU����n���~�BP�������0U�^-�� N5�)T���V2�N��zv�����]�"?��sUi�F����g:����1�c���U�h@�{���4�Ot�T?΢[ྊlD���ڦS,^�{�PH ��t*u<��ִV¸��<�ALFS�F_�M�<�8W�r����k5BcK����؜��f��<w�����6���<}��
��o \�ɆG؎�\�Z�8�	�#���u��DP��<��+q�<�&ʨ�̩�h�H��~gS�	Ǚ�|J8r�FG�νb� 	�	�'zo$���t�z�����^�%݃�.=.�`J)ԖDz+�Ҝ�T�(����*�-0ˤ9+G�/Yj8���aL;�C���SbPx+�.O�-LU��b�`�ѵě��E�aB�L�.&{�����ΐ\�">U)jr����3�R�yz!��כ�i��0d�n^��3ox=NZ�A}�R}�<y��*�'�xNW�������	���_��1G&�E؅�~ߚ�㷁T�<�N�m���o�(�Y��RPUt6�<F�ʩp-��R�x_F�����ح30a DX3z/��������F#�S�k�|"�~J�e�I80P{�j$Wz��|:.�_o���VDK�)�Q�RW��s�!���o��4�j�K��23�u0`1��v��=	�*y.o��?�����:D"��"�lN�j_�t�l��١��{à99�ȑ���߶~�kt���u��=�JI��ģ�{���E=	B1o��5��p��=�'��ƕ�`6���t7e�2���0�IG��3CB�C�l+)�k�&�@AZp�&Slz���_�\��&>�E�e7ӗx	>��`vI(���/�o����eN�s� w�*b �~I6bY�����]F�H�����"	ja_m�y�P:���d;���`QV��7����O��W��.�h�����(�.��ḍ�D��v�s����[0PA����t	D 8�*j!M��tT�Z�;Ng�C��3���5ZS?(�j:����M���g�BK� x4ٷ����A�@���ق{z`i��he�&�efh����T��$���뭪n��H'E��
�Z�4n���2w�j�1��Yf��#��c�z�
]�&u�i\oe����^1~���]�U_'�
C�X�B���9pƬ0��ˎEڟ��ZQn��� �� �6��̱x���s��@u�*���[��u]���Yx�_
�b/�'�|�vϕjki�o��-ut�%T`ڃ�ֻ�O��P�L�^T�*��&+^�`�;�s��
�|1 8o��?,��\v�0c�Q�tT��֝%>���?���R�A��%�͍��@����YKD�0~�jn��6
�h2_͊�	���g���B:0�kc�ɥ���:A|�sB\�x�����%{�g֔׃Y.,~.��+&�� 9�#��A���a0� u��������&/F��1B�Q^s|����E`��'�?,��g��?,�>,MuLN�ěPK���ڝ5��hH�o �����s,0~�X�!�ֻ�k�o��FmS-1�@�ͻ�4;|6�����02����1������0++\d6�kȉ�T��[�E�q5
-�L����l�H�t��KuI�xH�z�W8���JF+3�ʂ����s�N,uV�}�Ճ�s�u9�2���,�t��B�ݤv�D�쭧�@�p�֞��>x����Z�Dj�v��~}.�w�ewӝ�����C�X�j���F�|��GVD�\��Q�R��疋�a�%Z��OKa�k��x�u�ħd�@�G"]V4�k͜%�E��C=~C<��dL��#��>~_Ӏ)�n&��ma�惒M/�`����ߧ�8��KH� !�(���/���zx�N
����5��\�� f��_�^���F�D�#�
9�fv�Ð!\K�=�b�!���ϫm��#qkf��b� GJ�FsN����7v�)�����Z���kn���KSR��9W��b�om[���QI��Y�v�(�O��|}F)��`6�z�` �-��sih�h�Q�\?l�u�QJ�2C�>�=:�)fd���x�b��-�����@�P���+K(D[�M�A��6��Iӯ5����={P4��_<q\����{'z*��3\���1f��AL�V8�Rm����y�N�p+����={Z���5; H�1��ҷ^��F��]��E�b�t�P�p��	F%V�|Faȹ;"�qdA��@�b��)zr���8���:�ɔ�@�.�:+��[N.<!-9_lX(��8��;&u�R��)`]={Ӹ4����k�h�B��I�r�@mJ7���x��w��7�g��r�`�eI.{��m0|����v��	$��Փ��]?f��w1��~�SH|�!���h�V�W�-�Կ���^���<|����^{��-PƯ���j�����X�~w��*��w'�7�Sf���/���Tm>%������y� ��?��t�$��j
=����8�͠nb?m&�}�`�~��Fh��9͘C��~äұ4��f��ߒ�^�f,�W���d���,ᣉUg�N���j�9�%�Sֈ���;wF�\dE�F���,j���3s搾�
	�{�غv> >V����.*��)qw��:	�Ed�K�za�ז SK�s�;ZH��Ђs129�j�F *�˩n11M�Q��Յ�f
�A�1�&j��	�_���#e�X����f��0�PȘ#��*�z̂^h �@9o��Oy��n��RN�,��@(!�O�Rȏ��x���@^�xs9~�|�,²����<`�9��1����ù�O���N*����0�j�������sy�L��%ر0H��5�3{�!���kq�]q���	�-]�Z���K���}�"�^H��~{X��:�Ng* ib���l���m��?�@<#��`|�(�Z���-����D��9j�# Ѧ��M{c��Y���&.����޹�n6=�3	�] �T����m���<g�0XpF�w-e}�;$}��B��Y�?%��2ӥ�}n������x�x��C>g\s��'��:� ����X#8zPu�nȂ�yH-$�[_��l��%���S�� /�/¾�@CRS�iA�:��o~}��o����\� �A�<'�-L���I���Sٻ�[E�^U���Qm�䃯�����,,���$�,��P�&v�uk�B5�����2��G��Q�Tqy��G��d��
V�_�� !
��i 2g����rF�f�|f�ӏ�vL�3օ�ZN��h*J�#��5ip�6H5�"n�W vq-�z��ל�Ct��yu���Mq>�b���j�d�����{{5�$�9'0^�m,�v���c�bM��^<ZiNϦ-<�m������@Ve)�r?�v�ϳ⢕ 8�3M|RrA��Qz�|�:K�]\~��G.$��h
���`kc\O4ڗi�Й�j���%n�694�PD����d�:�j��*�Gc�H1�h���?jb}k�h����ϊ�_�HH �i)�C�f%���w)
��OD��2P֌�.�z����J 9���F������ZK"c�ʈ)���6o"�F�Q�m
��r�m��+�I|��u�E��eOH9��@����_�r:`��2пI�U�� �/e&�Z��ܳ�ȵE��zzT�a� "�.�zw�J�Iu��V�x���
qO� �����͎T���{�֓&6վ��}W}@[zvJµ�9����(���l"K�	�U�O�k�ˈ$�]�z�4.�> _��
�C{�E�T�Qbg�#*�N��7�GJ)��,b.�	�����3Ϸ�m,�~lQQ2qdkr)TD��%�@f�����)����+33C��tc(�,�qsq���wF	+H�@Q�SNP��孧�n��3_�e�֒繚 r�z�W�OS�|�to�D�J���`�l&O.��	��=�u篰��tKU8�����+U@ͲO�����W����tҶ�׌\�"]^)�/ɂ7ϩ�|�-��`07k�b;��t��
Gn�j����SD��L��H�e�]iό$��O���ñ�e��v0�S�K���Q���N�Mdb�]8P�0����i���NK�,��A�qa��a�;Y~����dV=DU����EVv���~dS�n&���"h��j��y�_m�>���N�9WZ5���
��>=�e�qњ�!4�g�к]��M����o2W�C�?�SK^�e2�j�R%��)�q(��Q֒m���C�q\���L�Ҳ��8���g���QF�t8vN��n�������U�xcO��S�4��@[Ğ#��gR��#*�P��9�P���	U�p��9��7�@S4W�Q�N�����WB.ohK�1Y)9�$����E�i�_���m���L'��⣓���L��vN��П�+���X4H�a)��6	*r�.����:��j@�q4�ӌQ�w?L�O=1i�ꏊ�)��� �'�!߽�Y�X%��#�d;�jD]������P���>���a��l��-�;ֶ#�az�ʭ�HI"�����e�V�^����$m��,UɯN��}�?��޺�g`%:�)%-�.l��Qy�����M�Q�QP�V��vg)D��F<E�77K�5��D���~D�`�������/Fj�(��_�]�w�sj�L
Ф O�@X� "\��{*�p̽�=�1�bͻH��!�OhW�"�<!L����wgT�^R4�}�绵i��:�zZs2�s�-Z�$�ϭ�#�t�T����!�P�D�q�a_4P#�t�oo
|���ؔl�1�>wBz�FX�3�x1-�όyFw������?�{�Y	�.��hB��+6>�m8m�?mB3�R}�$�Q��?S�':�HyP�7�٧w�v��b��@V�\���,66+N���?8M3�M���o��p坢>K���٘"���<���V�p=�kGݢ�1��f�k���ɜ�9~#Se��V�7�,M/)/DF�QJ]��������)wn��v|�/(��=�P�c|��k��NL����Z�h���Wػ�2b&>�O.7"���')���0d�B�W+*YC}.�qX=���6L���@&�L$$E��hb����QU�p�hM����߷%���I�GĬ��9Eͤ���\m6�"�[^.��_D�:���iR_� ��!"�$'F�����ཀ��g�G	F޴R���'��E��A�o���$0�{"X��(�@vq��l�{���]֞��4�Ů��d<��V�+fɃ��=�t�t�5��lKRl���5a�R�44���&��o����B91<�C�\r�c����S|moB�ֺ�ɑ�_�a�EW��y6�8r�z�)��ᮬ�4�����<t�=��@~��1��H+�j��!M��Cz�����m�V{dx�8��ԋ�����;0L�d���������>�#j��)�`�M;��ZN��1>��Mt����m���r> ��u����[�{�//=�P��%Ê�U
��g���JU�}q��m5T�q�@�ڇnq^K�\:&z��L.7�`VH�.G~����Ս�4���z�8*�����@��V�b&}����v���X�/�d�|-���סG#����r
��*˕m�Zm�T�����9�E������ ʩ�P	w���t��*#R�>^k<ϻD�&x0XD���7mR�G;}�J\W+���h������WQ���S�M1͇"�4	8z?�D���+V�!h���O S-aYJqR\*q�� �7<(Y�=*%1<��`#J<#�����Q95_��%�E$�sP�{W7b��������N�G��ME����9J�e�\��­��{:#�ܿܝpK�J+1 :�o6�쫄�#���}ۘrwAf��=����(Pbd����	)�毖�)�BA�tЖ	���a����lX�j��IZ�(��L#"� �6� �7�W����)�0����a�ԿZ��:1�Vp x�:����6:爐��l����t�mEq[n��  I���m�����t����|����M@��ѷ�����/��:^�T�S�5���W������L�*"7Qt��&�"��`�
t,��	���;Z����W�Azm�@�9��*b�*�h��y��h R��5=>�0�8�U��ɫ����m����>"fJ��ӌ��Dz6]���$?������T$�P��r@����f�{�0^�P��6訽�Y���]C��Myk���_H�8L�[4���?L����D� 9#)�u��L�`�����o�o1x#�����������"斱������s��Y�,@'_w�D��q	�'��*���MPκ����+��>˙ש�܇خ��dM��չ�q"Gu/�a�F��K�'�Q�Pb*־��Hq��9��ې�=m%�@�D��2�������:�� ���&�@�������,9�2N�{�W�yMU���{���BYC����W��v�Hd}.����lvf�CҔ�����^Բ��Ѝh��D��Q�u9���i�ʛN�Ʃ���	O�(�i��rڍKtS�Jj¸eط���I�G�!�!�̣������C�V��_&<�:E��� 0^][r}{�\�w6�trfw����#@���aQ��M��N�S ����8/�_�|�'B�V�A�GUl�� 3����!e��V:�ϳr�e��Κ�z�A�����o]	�u~��X�/�B���W3o�z�?^���jR��K��u���>	�I2�Tm����8��f��S�3*���*�z8��)s��p��]��Ws��B�����V�9��W��	�J")���-�!���b����6�lu�X�{v[\��H@���L��a̠O�/��H�$���t8�$w�	��,�Pa8',���hh�2�ɵ]��([����O$��Ya (����M�8� O��[�\�0ġ�1��V���s�@p;�=3��Ss(�ڞ�( u�����7y+�,`��pc��f����L�(��4�#%���;���Dl@f��N�R��w��)(^6{#4 �D�����t��vt�|i��[>��y&p2�-}�\��/����B�b`~�Ť�b�4/��oEE�>{M�^@���
 )�'0��M�Ucϋd�'�3�%���غDR	&}�>����?-��igI��hm3u�?ZG�?�����R�y|S�<�5�if?#�u�˓pO�o���}���W��P[�{~��K��6��ơ����[Og��������-��M��)���|�'��Ђ*�N�+�ЫŨ����֠��A���6u)�ȋ)b׃8T{Oq��/Đ)�����	�˕�F
j|)_k"�E&��0e)��
��ū��GlC�{u�]�1���z^4wz��f����{�EtyF|�l��!���R��#�V��u���Ic�)u/£��׃u���f�� ,�3�=�֛�r���Uc�47�4myu)#��	�.���Gz��,��v�mG�.pk^e�Ĕ�|��L<S@58R�t�oy�h>�Rۓ)v�	rC���%�6����bf�A�$�����Ac��ģf�#g���LB_Z(K娂�gU��
>(k���	����fI�
���<���0�+ �n�&����<�[7*!?��h�+�ц�X�w�l�5n�g���J��m��G+����s��麎�s�rD�}P��k�#j�gt3{�
&�c��1���Ά��A^sAU$O�Q��^��k��A���ܖ��1/�@�欄��>m�r��sE#`�,;��3+��)���S�I�Z�ZV�\��2ķ��ڹ��D��l�)�*�&O��<7k��'�8��p3���/��� )� �Q�qY��,�v���M;+f��ݤ D�H�����1.Xe�ا²o��Z�8��j3<d�����@��I���F�PG���d�f�6@�����	Ùi�ۋP�������Ƨ9���Ch�N� �m��K��ǥ�������OaA�t��L3���;z��\OYRs�&A�1c��&��>�������ŸA���(�$5r�T�}y -�,�֥�]�"F��֛;�s��Ay���"�u���(�R��h��T#\���)���!+pƮ5��j��PC9\���G�E�ک�W��Ӯ �����gT(r���h?���*�.�4��ƞ�HSHF���n��5.�[�+���:O��|����ӷ��^����Ǿ`P��(c�h��p����h�h�	>��-�N|�qaUxk	?���*�:
s����x��`�Ŝ���M��u>����Tӷ���Y>XX��"i<DL�n%d����u�U�B��U�t�G^U����j�'�f_�_����l�Z��uҨwL���!p�M���E�Z�k7
v�9Lq��ĥ��$q�W�����h�+3�:	e�gy�}��=���5��j��an5q�2a�p�FB���AY]A�R}.km�2(���؁��a.	�J�F��ܪja�������6J�Z�=��JA'#�8S)"HƐ��&Ao��\Đ?�џæ�r�&�D��w��- �J��N!1@0�-Q����<K��uQ�����J������7�6H'e�Z�:A�a�E��JS�$��ٚ����G�/�!Wt�� ���<�v��!��/����0)ʆ-%��	�(#��V�ߞ�E\�������.�ND���卋���L���h�%F=L�-()�g�8��N���eX�dfTRQ����5�!�)!=��{:B#*��L'-n֛%���t�x�]����V�x�`�!�ozH �0�IO
b���ʫ��%����v�;������a�.ϒ�n$g��<C�߂�4����n�Ҫz%�ɞ&�A|������~t��|�ң?���(���;:_�Q����/cqa��az1sF�9٠ ��ڏV��9�/�m��9���>>�x}��bt�<Z��g�S������JS�'g��}m��,��{�y�x�q��?�gOd� ^_�%�h��gqh�ž�w�4%��F�P�\�|�ITe6xu֍_sT��?<�x��8u����"]���D�*�,��)O��?ĥw�vv�r(Y�l���٭8�F�g��Y�K� ;�<�ʎ�I5rB�(�A��V ���|q2D��N�����1nA����'��SU[�\J��/�F:���v�ȣSC	�Z���)۾�74��{	�[R����?8��lS 8cg�k���|�������"m�L�q�GdJH�'L�	���*��#*��$6�QA]�oS��Oxu4��F��ńȂ�s�Ľ�M��Bw�yD_�`r��o�k�KG� ����0����ٳu������?3+g�Ǝb%t؝Q����H�?2��s����Y��0�'egC��wM���w�±82A��r�l��������)���͕C�;1g��E���D��I��}�JsL
m59�@�%����ӱ�s��O��QO���+ �^��*�̩��T< �~�e(:KG>�eX#�m�O��F��^{p�]B�hTm#3I��\N��2�g�=�wO)(�>v��N����L�ӱ�{
:����!�7�S���AxV{4�jb�x'u}qY��j�p5T9d���lF�_���U#������F~�t�9���&n��V����Ę���Q(�����5��N�z�Ȼ�@��3��?�7���R�Ey�:����-q�G`�	�_��xU%xf�A$ͧ�a��m�h�G83��%����!�P7�q���'�x1k�`�/=5���O	�IC�g���*cԴ$��2���eo�@l؈]|	��$"׈2٥�~Z��-��V0�*�c�����f���!����fT��
��ߢ�Y�*�E��'�<-�	�L��)����<_44e�\Q ���u�ē�!��4��t�z��� ��~�YԈ���.��Bq�Em^ l%{�����Q�u-@�s�eQS
v����p��axK�ͳ��f�u��]i��r`�q_X�1z�.�4�?Ǵ���<��I��WK�s���%���CBp���E�R�k$�Dᨍ��~�6��O)�a)�exx�V��ùVIR�K�%6i
95��1�5��4K��b���ˍA���|�T����¶�9K�{�O_�p�tM}|���&(Qǅ>F`y��=�:���34]L4�m��h^�u�=�1@z|�D�)�4����A��˭������Φ*6���u
z���J�7� J���<ǥ�X�n�.�h��)�=bl�tU��T$����8�I�C�!_��Ar!~����)5���[4O�]�@�B�h���b
����)�V]{��}n��t�Frߋp�����#�
�	i���W;�},T��_^?�y4Ri�r���Vd���7��h�@��޵A0����M�LZ�
��z+)1�+~_tj�h��G��Ɣ7�䭯"�M[��F~��Һ˻���}U��B-�]&�yxXI�k�t/󯢸5A��\������O9R���8�y�Ζ��t���&�@Z����$�����淿YM�=�^�fpx�՜%U�Il
��CF�{{��]�4m��3	�7�a�<R�����K^A=�P�s��+Ln��Mz�fF�9�uF�w�i�r��	�`�አT�����˼�Q�)9� ,��[����q�`��������iɰ;=� ��w�LS�e'�r���7��"�D�$xA�~=/��oE���)
L9^o�z=o�f�h�]V�w?���5C�d
!f}g�ܥ\�hH�\]�pQ�,]U6�ݥh ����*�a�baa �;4�)�{��X5ݗ���Vk]rι�%��H�g G1��<�v�������i�OQ):w[�z.݊����ܮu*�=ה�,��+��.H�'�����?�P����KB��0ǐ<fd�}
�л�a�Su��n�������P,�4������W�u���|3\!��Z�b��0�6�О���w����jU�X)�%��z�/ǻ�6$b���f'����{�W��j��k�fX��0��d${��j�ZY_k�Ph�
'��������C�=�Iouyzֱ���P�p~�i3 R!��e���u�; �_��d��E�?�����?�U$XC��n�[q!J���0��g�"�ў&�OD����Z�Z��=t=Q��tcz�f���#8#��a��N}�M̭���_J����[O��4{��2	���t��m��ͤ�i��!�D����2��!!y�i��Sp�$��Ɉ�Gf�r�5q����F�Q�g����fH�6�h	�G�ѧN�0�����]��+T����]�y����h�Y�ҏi�|�3i�t8l�:l�a���'�w�kM�b�H�?�$�K�5B�x?aW��o7.��#�Nϼ�I�O:�1s�����-)�3��F?$�&
�a���laz��M�3%!�'�_g���M,:�����.A;����)��:�f{�`���TT��XÝ:f9z�ȅ�}�A{��J%��\�I3]%�e�1��K K�_�^(1 O�������:[n��p�ĥ�����ɀ.1a2�h*����1��>��\b�D㹌us�4�g;�� ��<�b{/�L������(��5E?9�Z���r~\���K�@OE��+L�����dN�w~f�۵\��I�x��d�+ ��SQeg����/��"�����g!����p����%}�d�UIs����j�.��H��V��n���B�I��p�|N2*��rx�$����T��}��h�椀�wA���)��o6j�~���5Ϳ?9��_z��-��0�p �r�R���}i�-���@^�[Ol��|R=����Rv`�JN�M�g�Q��$��cE���aF6�J��x��u`+k�Fg�kfMB�j����T5�j5Qq	���[x�W�ە5��
��B�viZ(]��_�m����R��V�SM���S5��W�/+�ۂ���]��<VNS͗���Լ2e%)����5�^X����B�\%������|`L������R�."����
�����S#�V�A���`k��8]Ź�B�q��x�ɖ�,iZ�����-@6A���c�a���i�$e%}1�(o�7�@A%�'�uo�Q�{�m����7+� �Vt`.�'�@b��*��~`X�!�+S��l\���h�A'�SI��<�f��'�~�ؼ���k���@a��b���e��|<~�MI���x�� e�oX�2K�5�'�浤,+_��F��~M���ߢ'����V��f#�uـys!0�5���_��*��7eq�rB}X۷�`�k���r�"��n�G�*�gB�|2�`����\��B��'�w@������ѓ���,��IvX����"r�og�+�w�(Xe&<��{�*X@I;�^�
��83�D�w�U	�-����"���FIyb\��W%k�-���6V������(H��Z�!o'l��-`����.���+����J�k0�ΔE��U��+*`�� 6z0��ZI��X]˶��K�?�"�k�;�ylZ�]�Y��TKE,�)y�wq�:t|�aֈx́�W��-���T��6�gm�I����Q)�A�����f�a�ٳ!��˟h��͗���h��'��K2���������*�*x-q�	Ǔ���'�.��bI���R�)r�{�f��0��ɀR�{�xNXEv�4��x�Eu��qĠ�v�u�\~\�K��n��_¡Ai��K��A�zBk!��p������-�U0�H�ڽw{���M�;ZI����g�9��8`�q6�?��,�ZqMe���SP���I�iМ�2�.�9�
���5��'|�_�r �T����=� �p��/!,6�b_"�e�	~ḑ[�b2�ӥZ�^�o�$k+�M��y���5b��2`-M�ᖪ�����\�?�)4�Dy��&Lg
�wKH)ԇS.��\�F�0�	;g�=����*y/CΞ*f��K\��0pѸ��设�RKq��ߥ��:�?��S��m���6KZq�� |�
݄65���Ae�S,l���kU��-�� ��D��>��\�%�,����[[���-:&b�ct8e�ݖU�hȽ#�o'�=�&wI�`�r.� �=�����<�)&�!����*{��֧N�/g�Y��5T>�غ�	Gm�}��d>4�~k�\ h\´؏�d�>)�֮.'����� w��:i��%��|��Z�8����]57n�&�t���|�7�1Z�y3U�����u`}:�9�O�[���#�r!����H v褟�I�3��J���@P��-�7D�����xBa�p�����d�b�Y)K��^�i���S_�},�������s��I�w~�,�;�ڕWa��Qq���r
����\o��w(/u�q}WY�fFb�zQ3EG|�EIe����|�f��q��+��Yh ��B���[��4� ���c$�ЋcL�DP�#d$n���K)�m����l�Y�ca�zfD���u����V�+�ؖ�4�e�xz
�q����ĥ+��0�����B�)�d>R6|��9����j*�[n�%d}?Պ�r��E������	�M!q��M����u�A���)�6L% �I��rJ�ߌÃ�"^i�a�0ǈ���*���GVm�w��V�tf�,?��ɛ�c�F��7y�d�d�&���UO!��|E���B@��9"����<��z$�5�]�Z4�AKc�����aM&��m�񡬕��fV\+��u��m�w��1-��(��SG���T_]v��4�B��~���u4�'��,�H8�m�8����yuQ�.�%�=.ݟ2�;fgj�Z�(�BAw��uސw���a6����GwaP��4�:��ȮЋ�XԦ�	cgA��v�� zە���mKL�����~�����oԛ|=�����T�e�y:A̫�c���aD{���qI���K�骼�E���)����zХ0F�)2�|��n�2��X�8��s����w����O�p�pPgM�o��m����O�oK�#������oR�ђ��3��/��l_�Te�:#��;���83:Y�tE��@7�����
F�0>���y/�o�ً���Zي����`�Ns���j%4����/�8��M�=�:�&!|qF�b̒�Ք)�왅ђ� ���5��o��-.K�Q�|��[zӹ����0O��;4-̄
�U�N=w���*0�S�i������q��	㹋�h��jy��&叜��f���+�v<v3xG�Z�KT�f�N�MPk`OR�mvtx��r"��Qe��X>�<Vn���&��3ʇ�i��.S����6am�=P|.���9�|�c���A�E���4��Ou��D��-��	��h!B:+����c�t�Z�p���#M���4����-ڟ���~Ng�JF|{*��:��f��g��ܖ-
h$��gc�7�6��9��<#�i�Єp'!��:�$7~�A�$����eL�Z@A>N���r�..WWT����%J@,��g��-��˫*�s�Z�Eu�q>�}O�/ N�z��v�������O�)=3�r�r��v��D8M	_֥�K'SU��(���]j��k��»:A�T��S_Z�Ӛ8�N�ɀ~�wP�I �4��]�C�c���[����@|��Т�E��_F�h�#�)���0�����EҶ���e������LHs%9�Q;_�N�n�d�eh���Ge:xc5ˍf�.#dS�/�� [J`���^~�jD9w�sj/,SK�&�=���	}6~>im�����g�dC� 5`�=�6�{��˿���Tn���#n]}]����ã@���[�#�ܰ���{`�ۻ����S.T}�/hsSĵ���l�,���.MR"ib���O��H��i�\inzk0k�+�����u@�T��lO�:6A %��6s2��`G�(���a��Y��}��E[�}����b�fb)��3M���F�5T�E˞�	���6��q+I㣊�Nd���<[P��}��R��v�>=(��c���2�$���+�7�p�� ����I�}���8�-�f��#v*�^���҇�����Ů7N������:�� � V�����?��xD���>=@��NV���ۭG_]-���e��G�"����n!,�aZ6�֯�D�4��p�+�F�G�t
�.0��#0�e��LA��Y�d��GtQB��>#zK�2Ѻ@M��{���6iؤ����r��
�c��}@"�S,��4����a=K9��_�G-I�~aᴟ���M�~��A8V��=殚P�!��Л����l�B7V(MUK��D���kz@}��ٮoL��IT�rP̣Β>(�+�Y$|���}Bb��1�Ҭ�	A�J�@x��|%T�?�{�[��o�44?����g����@�P��r33�ɓ��<�f�U�o�aD�ǋ�FL������{5�z�'y�H2'��f�$P �	t������u#ٮq8�zvq`w�3l�כx��ނ�q�yb,(?(��%z%��H^:s�1�u��>�^�5v&����9�w�5"2,-����aTD;��#��.��[�+�A]zy��u~z#��dt{�!���$��M�a�ç�,��?�0�U|lE!�Gd�Ӄ�����eYd#G��릩?A���%hC��p���s�+w�tL�a��ʳ(����v�ߢw��_��PZ�1F���U��Z�Oii���ek,�6�z6X�rd�m�����YF4M�xSO��\�q����D3�]��`�M=mli��_�R�{U8B�a��or#��cK>�A5��M�9,q��%�&���O`A6ա���w^��m�a&��CF�X-�,^��uv�	c����~)�ߧ9Hz1j�h��8l�j�	tɂN���_���$��vS����
QL�l!�m���F�(_9}	>N=b,[�S�F"w�|�p�bF���'W��)cWYl�3�{J��V�e��1�w�bR>RŅM�Ck,r�쯑z�Љ�oq�d�D2��icwT8x���s.���=l�4)���j P�3�A!����Cw3;�Ok��a/�7�ʟ��T�I�����}Y=+�z�<R�ޭA��~���R�;b��T,�]���e�حE��{�	7x��j��5zJ+�R+Q7���R��p>��ie�a�0Y��T�d,�^��`���⫁���zQ���k�܅̿�"z
H!�P�����[w���a��u2�ܵK�z�TG�W���8R줸As��]���EĀ>�>��=S r��}0�t�5�\�l��O@#�O��fQf Ԅy�A3��iϏXk��<�I��\��E�G��M����hxO¨3g�	Q��7��<'�q!xL�,`R�6[�7���|��»ꂋ�p��ڑ�֫M��O�h[�>G��Eӝ.�.���(c,'S#;��IV�����_��d{��|[t�3�f���t���rf0~�b�oM�N$�#�Gq�Y#�T�ԣs�qQ�r* ��u}0�>���V�f��'Z�z[�j�K`m��e�4N��b,m������ƪm���hC�w� �6�Ѽ���Ζ��W��;���/9n!x��;ǆ�룵v��� ((ؿ��ɯL�7��+{l|޶>���Te0�������.<󧁴���{A�J�Mȟ�pW!|cr���d�[�,�3�|�CP{��@w��\պ.�b�Q�F��ț����l��$8T>���wz=Vs\1y�)��G$HF+����ɣ��O�
�u㢶��Bm���?�Y��r��B�Z��\9���f�Jɠ��@�'ާ��f����m{�6 h��O�[?�Y�3��2Ľgb*I�H�,�m@��r���rD�,�t_���E@ҡΟ*�N��ݚH�mVG��,B��9�)�*�N�I����n�1�޸�ۼ	.�)I]@S�-� ]�ړ�Њb "^���r볫
�wa�F
�>Y�_c7ܤ�Ռ+]���2���"X��4���#C�*���kW���[�?c��]�~'�L��*��� X@ߒ��� ���pj39��㈤��x��q]�2�ۚ��2����.��-?j?Z]u6PF8m!3�� ����tS���8�=U+"�Ip�r%�.]��0���"����'��#w�ur-mY+��D��I�)�Ai�FYޥ�09�/�黹�C�<<M���R �) ���I**-�
%��~��ܾ<Of%=v�����%�M�觤qEf�n��l����"�Lb^ԅ�Ҹ�eO�dvܒ��}C|��LCĉ�M:��FGF�����vi������upN������+&���ݞ����k
���ܵ�� ٝm�J�}�{������x�	��.h��AZ�Ui�*�x��D	!	�V�RR�r��@����	r�ǘ3U��f�=e�r|��{g�r�pF�Sr�t�Nz�cS�z޵g�ѹu/��$�����ab�(�#��b�՘�g+vd��~��3#/�[5�)�{2�:�Q	 �v�/������y9]� �N���΍/o��q�zN�}���i�P����֝�N�=��C]|e����@���s㛰IR夑^���bƦ�h�\j