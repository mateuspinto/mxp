XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��vTy��]U1�'/�\���
��o�H��9*'=�t-��	~���ث�ʸ��6J�3�s�@������$� �z�u�X[�B?���̔(Kn�Au�=q��Rh9�j_��������7��a^��JeM��0YǑ~���(���O�
٢��2�ֺ�o=0� 8)��f�U5x�S�82�:�t��JT���0�"4QI��i桶,n_��_�<�{t?8��fY5����d=��X�p�86jЦ�|���L�2Ǿ�����7r�B�r�^��@!
��6�+GJ�Jn�@ES�
�Ѯ����D?f�B�EZ��s)+��/q�M�=�I]C�����o��`�]E���Oɣx5n�Yu�~��%� �����E��*[9�Y`�z��V�7w�VG�M}| Oλ�~G���(��%V�3����C|AȜ�|�e�$�U�X���j☼ J,���Fҕ?��P��F�Q�yQ�&�]�mF�z�ѓ��˂�����­eKO�m7�oJҺMR�ʡ�@�!g��֜"��l���?��]7N='zC��B8����j|f1�'�~��̾��,���)�Y��LKal}ʨ��?`-�O�X��O�\���9�]�]H־�	��a�:�N}a��e���Omi�(,�za")��e���.��<���J1�����+Ⱦ"�a�YW�[3�{Bec0y�B��Ɯ�����Y�7*�^��Ƞ�r,J��]��b��S�x}�`H�XlxVHYEB     400     150��L�4� ŵh_���xX���祺�tM5�f��sɢ��� ��݁�g��/���DN�8�615���X�mX��+I�?��{؜��� ^,�7�]�}3��HA�I��B.�X��q�fݷ��8�w�ޡ&U2Q��߽qwL��Q��
%+����i&���U��"�Rs'c���l�d~#��[��V΂�R�&B>Gi��_;�k�?(H&Kb�s_==RR��p,c�|�)���&���d�^nK���&�7��УmT0��E�幬�`<T	�a ���Q�����$W�[X� �3�0���p��g��2�Q��E7�^|?�K���H��G42�!K��XlxVHYEB     400     160�~��x%tS�O9yB8��M����fS�"�,��(}�B��L$R;��y��g�gUv�	�&�D�]�^®!@�_�A f���D��ng&�s�F��%�^�:��ln/=f�ia�.N�m�a׷\.D
�. ��&�\Q�6X�o����Տ�4���6�В�i�{�3��P�-�,��5�4��?:�r	P&�F���H��s��`i&1�T�DoN��Tr��?,Ƿ�+eX�%ƙ5Tl�ӳU����n��[�CA��]
j��J�����|Z��B��V�y��R��{�po�q �_������n��l s�������k�a�}��/\��PU���`zӦ��GXlxVHYEB     400     140�'
���N�ثN'��Qw��֏�പ5M�P�3��B�O��X�7U�n�\x1���O����Z�7��y%b� �͂�vE�V�?��χ �q�o��c(Y�O�#L�ydV�F-���)�����f�f%��/�)�t��<G���9��`�~V�F/KkH[�c-�UK1��Za���dq�Lp�E��!�ӟk�)�p����apy۾�C5��pѿ���V�Ͱ��1��y�m����b�4ic�
�&uyߪ.�޿5��L��p�r�?��<o���I�����&b?����]�oBT�Њ7M<uf�j����XlxVHYEB     400      f0��!|j��+�LN'N|K�98|_3S�����w����U�?�w���M��(bӱ��܆�[��uC��|�%|���H	�� |x~����ZǙiH�=M����2�B�yPeUj:�8v���WY��E# X	��m��y�GI�}����ڇD�ӝ�+kzE3�mWX��غ�d,�L?./����Lo��2 �p��$��O1M�)�uГ"������EI3��5�T���m��tvgXlxVHYEB     400      f0n���k��$����f=�h��R��c|Ÿ�5E��
�[�B�B��2�,�����9;�1����_�e��1��@l��6q�57�⏴��D�>�Y���VR�a�����qf�"]�3���H�r:c7�!�]&�-T|��/k'��������hIݢj̠K����C��4Ǡc#���OT]���H'�<r��Կ�$$����,���ENg~����ҍɢ��� H"�ʥ��#�j�Q���%P�z�XlxVHYEB     400      b0v���m��DZ����;�#m��1_��/T����Ǆ=�'`�gl�_G��y��3V��dg�����ú�kqs�ǯm��!��c�|<d��� t��Oz�D|�%�w�؍�*�a4`Qk�W�vyF-T~��)�Ձ��K��̆��`�^.�_�p�< <yh��Ϋ���8/c0&��XlxVHYEB     400     150���@L�}coL���?���e���Ӊ�V�hӜZA"ɶ�)���=��R~M��@.�S]�Vч�|T�Y0�%��]��ǰ�D�8»c�z�����M}� 3�4�C�U��oj� �|�q'Ӯ�(�
���֖�@Q�Re����b>Y�S�Z_<����A��5���,��w��vR�

��+�dq�M��񥃢Q�$\�nk�dێ�Kܯ���R�S]+�X<��(�L����*u����\�ko���-��U	���K��]��b�K��Js��͉�4�Je�)�%�7���S�C&������nZe�e��7������!?jZveXlxVHYEB     400     180n`pk�L�V���� ���9�>�ON�q�0��#6xݤ�\����ہ������Y%Ϥe�K�*S����"�'��*�,��0�uG�������{s(��TԱ܈i�\�Z�� ڿxT_�6�g��h_�ΚF��:��-w �I8���#0��X�SO��^���"���o,�{�i6P�H���q4���?�2M�y2�Y��zH�`,�Ib��x�lC�$�}!���{��(�SF��-.bhtA(��'=t�~�_m7�ܜ݉-q8AƲ��=���7豂~`(�� B�Ý��3�HL]���ȸ)��s�ҥT���bo�מ�N�ы�	!�s��8BEi�M�o��()�mA2lrlUṣs��,e��XlxVHYEB     400     140ፇd1��Ö�)�]v-�����PK Ώ����V�<$��FO`��%!���S��ɼ���_�����a~æ
�}�G�X$o�#��s@5c'�����1�߷���Z�0󀒨<�t@�� cvj)�t%��	l�qj�j=P3��qmy+ ��'��: �'��$�Wbvp,މe��jow�E�y!-ض��iN�U�VJ�I*͛H���4`��.jʸ��<�>
������>ïc&��#�Auo�z;Ds���M8�#Hi��*8~g�ed�*G%$d��dB|�k��*�Z�����m�~G'XlxVHYEB     400     170!)Z'aWNgA�u��Z"IK,��~Gi�J��ۊ��f���S:���j���\����9��FjXYpxvm��(���0��S7
�����f���R�]Z���^v���!���QTl�p��{��w��"��W����l��|X�Ƥ��=e��tC����:�d�G�O[����F�ī�Œ����$�
����`&����^'2VV���v^���g��&_��g�Q}�"dM���R�]��bDh.�b��{�OɎQ
�5Խ}
 3R��UH���{ϯ ���#�^���$3�V>����8x�g|�znh��R�Q̑�ί�_���W�WЫqXlxVHYEB     400     170q��ܺu�P��o�ȱw��� �:Du�S�g>���e����B�U��'�p�S��YG��#�Y�4]���yQ��JuZŜ,y�r��B��w	�K�(@�`�	y�;��-�������� G1|Sf]��]]�:��Nq�?֢ܷ���#����=��̢=��� ���&�%������h�Vx�_�����$M���M}w�
v���Q"(3����iŶ�Ҝ���5��b#�p���'h�������p��~���y��u�Tt��o�o3�]k+��[X�ӧc�i�4�m��lo���L�+e>gjǤa�_��vYnj�|����^D�E9lX����ᙞ�X�%�����3w�Z�XlxVHYEB     15b      c0񯆥��x����4m%�J|�w�N3�|�i\���ݘ�Sn�~��̚��%r|-=���Hz����*���X���f�P.Vz�|HјG��|p���I:���`��*��L<9�4�Q��1k��Ry�h�@�G���M�p�TX�XO�"�i_ƹ*��~&I���>�0�.������.D���R��m��WA)�&