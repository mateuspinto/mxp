`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
hDhzwfjoAEQHppHYzGTqHiB3ETYAsYkvPTrO30sPa0COEhUkXFUfhXd/gduvlFvgCTADcAyI02+p
3EK6CsLvKOoAQs/yRs+Hql7AyDpiJTLXHcjxUPNp1cgLGyvuDcjtOXpHrbxZWDaKrb7ZDNLSvD3u
gYVB9HsBsqPnbpZKMGp3MHmbZ9yjxpyDQFf8tu2tOCnro7TKs4nl0J5PTKuTo7qTpp3PmaOR2ZiA
+U1LSjCn0llKMkEFVtmVv8IzyCUfJzqPL+rY0ualH7mwWRZG6zGeMXq9B/uh7JUwaYCiIc5h0dST
2Kogg8On4Al/aXNWo6t23zie+XL88rR34NGxhQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="+WflggqmWQAcIP4l6G/XPpuI2VpryR/aM3lrySjZ9TY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5792)
`protect data_block
5XFFAPT3M/SxqydMTINIqswy0zqBWq3NXh9z8+T0ibWdgqj127bfXZ3SeqUvrT0jAhb+RJ/b8iTE
gcjt2tnQoorTtQTsFtVy1isUVt7Pt4yu0d6KZ4mO0J7ebUh7BLhjOjX1Y5TLcMAN/loV2AXcjRyT
PEjYWRj0Dn3hLU/XIF24BABJkuH7M0XNRa8VoX4C+RVhKfn/j2m3OFmdSEjuP3xbnt+N5gtg0HCN
q1pwj23EtcvpOryGXwtHXwrUJqPKNsrh+8lJOrAVfe0eMjtgooPjP7Fi6GUNCIC1qFYgAZ1nQ4jq
AjS1ufmcNS7bCGo5drNgmNguxUSD5H/Rb9oBtR6TDrCCF1WHRfbJLRwEv5LrkYG91DsIu1nMHZ70
lo8wyGqEscwi5ekdsyEJgRN+sbTeM/5fTXaJeidGcbaBkSk5lTY0vCzlKxYjQWT4Q/LtPwVxNB0Q
pilZArUsIg1CITpTcEMdEd4q8cOdk4KZ95N85uGGdtMTbT/sypztgJ9SV0HvK2xLEzU+iCDzS03N
q9/Zrsyz13LUPiozdjS1MN/r49o60FimaXTQaX0OWrOmWpKr+j2epmjzwUksfqWbAaApiOZDGHcB
OIwpYT1a8m4gAmiqTQjaFwoSPHCR3c66RRz8tgzvm8uhHbOyzQIY/UgWCaDPC4tNodDIN4MXaEnA
d+KXqIkhrAok0IxIN8HciySY8FhJjYtBrx1MYIHKaD9GUlHEtKz/wPY8I3W03QzfxcyQmioi9YuT
jYRpEh463AwfgM410uYDK9wQ48sLNoXE7sU5KSzUWR71hHXMbvNVbnKPSxSr1cz0pZM+TOTz2KHA
J6RRbHlsWm3qSDqnmBCdZCv/8PQa6dy2ol4e3We52+PaGedRGWr2MJQoO1vwUD70Cp939JFSAC8U
NhPxNrEKiO0jrl74/QFD9eZ3W+D0Nf0+HjEwYjdKmnsjc1DwJbqawF1lQeBc4UcpkA6bWYgBkQOc
gB2SqjZNIRmcl03OSxndejlC1rd5K2MN+Bcs4Uvr6nBZkbE7EB09dhrtvDLSTm29m3hABxLsrNI3
w+Lcaw4PXAYAgKFbVCO9DhsDTXy/+kVUSJASfYXZSZyUiH8EqtXsRFWcZTYYi8yH0AXhdhCVuGq2
I8IlYVXHfezYSWLSDfUxkAMYOlvKm8MX/Nt1YfgxAl1V+AkSaagigf7g34RJZ8La/+5sfDu65Fr7
mmraZsS9MpvY80teOEXSBBka83BR+mhIuscvar3Ur3bmX+WylmuZd2UMmvYE2p2W/K/pTykso76u
7NM7TqT3DG5jc3EeuKhfLeDpBBCB6CqefQMWi6UYpBAuqrvF8OY1QsuswTrkw86bWu3op+GEPCkF
XtBBep1qF+dQ+2n2+abZUk3TecvIDgLhCAgo5PoLTq6XjvO7wVqlX6JnHEhIAxNyfESWWQwbvVEL
8tDwAlGiTX8XXXrVTn07Nhkx72f5jyouV/SW7NxplWp5RScr0xO0fBoFrK+tgdBthPIb1OjyIvxD
z5scPC18dkr9LAvvwd7msCq/iTMU9kyXIg69A/LUyjYWyKjUfIGZd7nUur3TG8UWVh9322pIv7ut
0fBqoNP5t2K+MMeEBpqUa34WDEuYAXR0ZbCooquePVsCPRg2l3n+8/+57LPMCwZ/rJA9ItyfdeeO
BfvYOTlNcvK3eKRuEqJYqTg1anbF7tko9w8YqLnTFE1vQuHyoeK0rOs/3TkHe/hSlx7fZyC2hMfj
GZ9dJjSWlS9QQuNMGEfqIcffhS1nBperdAjDliEf9XoRelrpDnmUxY3N+rfczfOIdzXu5uuaBIud
tIaSh14/yuj9G4WrOPm9FUWjVI7DJrbP/FFB99Eh9M/BpnZ8F/hlorCWZqnHKtetEOP4GLGpmCSn
lEsOiHYwOdHCBGDS5ZW8tPM6PoZuqQbHd7JsMUQvSo+OvyaYhfSy/q3WeZKIH3ood/p84CWT4HFW
4YgZfYF6wkP3aMDku0X7s9T+0f0k9twTanCXcDcjqIcv7ynkBcD9bfvfVVHowF4RvvVxJqtLulI8
shYhJJecT2tOWeTwPr8u4jELgcpCRYfMEmWEdKTh/cypY0kbTMsF3bbaTmrHpoSMfVynPKrdJLoL
6BNc5Q1RpqBPzTD/Ky+Jt2ahx1bD0nfLrJsNne6/h9c9Stsx/x7Av5BTJn8NT5rXHf+qtziyQkZa
ukryjTc++I9ugT0SAzF5cSWd0Y1DAtjqIKCotz4ss+4y9DbpRSNKWCM0oiezh6QEhQcfoTWPnVPT
alGPH9O7Ok7Tdb8KzEbeMcLieVKL4zto8+kcvn2jRWh88+LnWxm36llpKx4I49cTspAfnYIF6N0n
A2xbqu2TNgZ1BGaucjM66XVxeEEn6j2GASjo5KbrBLFc4uEF2OrV0Wjl+YZWwPkrztbHQI+JP+GT
v1np5w14TeNYmDb4eiblFHlpQqaVCYBnvturJiFGSX8Xl4OBWa/ar6P+SpLW3DGQOz+DjjiUVcgv
IdDFV7YJVChQDKmCdxbf71bjm4DO4noqbsLbhWVzUGGme4DvKJtdcr8YCq4J/pnNHxkUnaD7USDG
N7RMiBPIcP17EcTxgUlGm2A+W3CpZqDzYMui8DBXhErgMXK0vNksMxRreRIdoN0oDyjnDlDRK2n2
A+Zi5VUsJAplS07EuzLMZnRcwfJSWTGPdeJRVy/1p5iPvOqL0VERaviysSEoVO8/dlUCXJ/OGwSX
263XloT7zsxAF6uO+2cZn/0WZZybta18lKrYjK641C6eJUOia9yL9tzREqa9O6EvA2JpEqCfd46d
yRW3m8UuH0yiyQQ35IdI2RKVuOMoMAXiH90YxCaExS86qAHiZ1XGTzR5qYEoktMXI3Jp5gF9XiRc
DXKvnPDywh2EBZs1S2LNLD5ijZ8Pgb/YQ8716iPbgK8kvmJ1ywNb3EvXWCPH+2LZc3Fd/RmO8Mwy
RE+Cy79ZHUTC1EdVz5aurv3uX6jB9feZBdn/FavkXDBHJufO6R8JR7dyLUrYKg4bOOW8r0VOHA/1
cKbbOxXzx7pWrDfAZ3PFDWPAtPo2zipvl88W0Qt5MnWNKaX7XRfLyaCKMUoeeOqZPPNvxS6aQ1qq
a1mLkb7AdwTULoNarxooGtfOjzoTwYU4CneQ4jbyTgNt1iRu0iey5s+XEqwt7JDuqQnvCFnGDGX8
rVpCtEqle/6hVLjD9xS3ae9l10ZC0HUGGElaaBqox51bZzZQ2/7aD/mXkvtO8D3h7O9HT2mVoBKR
DJvqibupTIZo1N5oq9xQG3PmDFTNQcyz/tUoz5CWXMB8EihHD7+nl+LRzMCBcEE/xRGozIIo11Je
ctm9vJn/KJzSBEdi1BwCeFQ3PiMXao+qX1nfWvWz6X/O/gqAHeDTqOi9+yPoqX7vJE9qjL7nimIZ
5mtTqCSOoKapEv7+OB6qu341+KeQXa0X/VSAWVAEraot7kDdcxBFz6YjKqDf+Ulw9Ys596eIvE+N
klaIWEB5ZmLgkqjlnolMiP1UXv543nN6do8h27iTVE4eiO7NOpldoZCS/fQXg5vEOutGIlkY7dSE
SfM1KqHkv9QWzJpdrOGdxSbryKY59vUrZz/mhcDdwXWWDrz4ym0KDfAAIdplQBv0mfQoGcvSZl2q
gxwbnyjcop1DJpxyv5+saT+bfeC+8j2T/9hHItvnVugtwA3OF8ZGV/zytmjypagXMSudiBbCnDvy
A7pzD76Pf6BMikUiSGOWrmVfAuNErPcyDhxf32E3+G/dgyMgATrg0DLZoncfLMESKLeulE1xO8Vy
w3d0n2b2QEslZZgHcuNKk/s8Gvr3TQe3AoFeMQ3Bb0kRzK6wSi7qlRGjK85yyIHmO3DdDtxjHyRK
pOUgTrIdMtRrGqvZZ+0gwnv27BuhgBT5TLTs+44mwXbtiwBRXCrnas8ChOfqTupUsZVm1EUArTMO
5ycenCriqkvTIt8npGoWZUz+Sv1SgoZZ+YWFvx6e2EmUa4oYniw4Dy5s1A/5ZfGdmyT8HDUEblsY
U9younr14jlcHKxYBgt0VYLKxvZmNcrsMdeexcbN77tbF0Qrjwmm8gx/3HMaPoTxviwqat3a6Dya
VF1y7OceaeJkrSEM+skF0by6YCxBkBE59M35JhqK5Gll6/QtoUhwc1c/HkMDkT8JLUd69/E061T6
3ZmB5pKIZPwOewTFHgI4ZKsJhGDE0CzigHn0ZpKPEzxGR4+pRFcc9zi1zE3BRJ4bilAh3KerU1QR
4fDcYZdSEzRYEse6rlwbJSjE+S1jhuxfMCJhw/ehOvoDoF4aE0WQb4Kr5988EnB7lD6afWKfy9bK
NqyM+Px19xS1EC7ALBaEm2AJX9ggz5FgSfCpUsApUbJE6uPnIcamDbygA0SlWqW2UcpVWG+X7gMW
CDrBsaSk/PWtA5hC8EUXUCRvY5mxsD5ZceeFkhdYTvgXHoAiPXD82ycqMeU7QV5gI7pkskifPDWp
UFtGBBY4XeoTu64PlHgwsM4tb8lREjiexoYdfCyzzGLCcdKgecv6BeqUig6RZJ+J1bAXH6cS6/sD
gM+1nLBFqZ6NICt2e0XcAySZ80Fz/PRuqD8xjPmzWecYphEIAJLMFwgfShUkLXVY6ANzBSWjN3tU
JnaFTVN2wnuBbzP6aFyoM+En2RSjLyDKsD1xJaA1eub9rGx6WGY75xDsay0VK1QGc9RVbjKB5X6z
oDZlXNaw7nLPHKoaZ6ecMMyCFsRbYoT2Bk/sbX3a9e2xfH+5HBkSmMySsICcIWvGl7xn2i6s82U1
HkFC8vuu44jU8P4842KPSkUP6fgd8NX+2GBNV6CRmU6BAVUHvSaryJnvDCpsCv4RQZbD1R9aeGY/
33knPuNYcjSGa28sv1864jAkQdApPr/7TMmOt9YEA3G5Gr427qltRTFhC4d0PtWSJzuCSAvbD9nk
bQ6bKqFsY0oodxQyui3AFdoW02VPFUj0f9Tv7DYMm1I+PM7r/xUC6SOIY7xC25dVBIuI+ZNRQFD3
vuyJbexyLykuCeBdQnydo4ngpXOOACO/KbeDUMGRR+dBXxHVX4MalQKN+ZKbGywfMnvKOAviWTpQ
fOYi3l8rb1H9IYUss6n+a654PEHGtAGiZeUCj7yMB/x6oHi4h4tX8ChUwzJNB4a5F5O8Ld+/3x5P
NYJYS6YBtm4ZMvtlaKxpMjmEtG84pbAVEruQU1+VvfwgTgPvbR9gkx4qLiFwDyYmsOySMs4qbOtt
ik4ZeBW5N4QT1VokMBFOHie4y4uvNwu2E3Dy2Ujey4AX28dHOlLWekaeNC2AWxNf4M2J2eH3HbE9
xEfsZsHvr5aVLbxzE+33jOhWbO70+lMiGDOAlxIMU9EmnIRxUBo862UBMMEv67isjtgd7bHvnxHZ
p9vX9hzUl+NC1Ovd6wwkSE3U8LBFt2lUyxBz/gnn7MxzDpoyiZDeiGVnGAgv9A+vDAkqSH5QOgqz
T45f8KARncz59yv0mDmtz8w63YTl0kKfHYLAyfWWMEvZjaq9GLd+YCYLNeohHiNlgSg89EqvB1Te
nEMZIbEOKPdwzdECLIIv5CD8mLhuIpep4Mb8NRNz9Tx/mo5gH1yQuN0JDTbTyaP2U8rjS5/pcG6g
ePgqRhTgocEo5TSTSW3GJ7It5bxW22t2/CHm7BfiChcy3CurGaJqKu4BnPqSOxlsGgXnSinh3zbS
aK0iyfMphaToOzMpyfdmvt5Ye1fMsCB+juG6wnL3VZiK5H0GlbT4JPNoJdLOVPgSQQbDGkORCucR
nPn1t/rONi5wUJMpkCcy7+UE0sOjHxqvm7vHLGI5RTVZBjpc1ud6nEKaGaN49T+yxnliextpZRIm
BJkj2NF/22MKpboN1T6Pl5UTtQ17uy/S4OLrHf+n+3J3rwWFuvAEArOszoyMnDUZ9K/ln3huVoPr
DbNd2pTDwNvB/6uLGGn9tLqKR5UyXJfY0JI3oCHgFvVBoSuJ3v0Fo+L+IiSCVciiQqyM1pwHsaAP
DFp1C9P9aFytxQavPvcJneyGjGitjjVqP4yWwOv0sEkSG4NFYJViu2B7J2UgXX9E/7Qeyy+XLpNd
35c1xYmksu4Zd4t1MFqr3dfKLQsj3Nqd80gwOjvw1V65hQkvocImQKp5HSOIUQOqRV1W31baA3WL
E9cgG5k+koLWsROQvyntzCn71JhCbGZWBM62u92q+fs3Il4v4DG0Y98y2rInNsqpacJpLn6rFn0e
Fb34QMJ3KDJO6y6aKLyxCyVkcMxUme00y5Ncp+1UTZBYJPcquV73R1RX/nqYlz2p2bZ9/uX+oAjL
12wDch7buKsunqBF4iZYn7aLTJN//VYjmGQ4bO6sB2AbhonR209M7zt/FvK/bPIJ0A1J9M0ejT3N
q7TV2GGMUnBd8HB5oGKSFF/cQ1B0IiRaQpDKfjouqvI/8uEnbIzdBoUzs/IXgmxLpTEJNQK/+vFr
JQZkxLHFrD+dYp9DTP6T+ySS48QmnKU7spK2r5hWT27hzxoicmU8+FvWemNg8+ZezCsdfDvgbpAV
MJ120zaSKry3IwmZoJt5yL2mHcJr0DF/qjD6EQ6KCP9PNpyekNeluK927yCquqUCtqHZGQ/BpVJb
bcb08clWh4KcLqocCjyRhckZSLiaNB9uC3OUGBViRq7L7/xczjJ6Hv98WI5fHPtZNtWvZLRxGZ+p
y+6ZC3kBrdRwO6pXIIuofbPf3JfF0fnkhmXrAS+pt5Dkw7VL8vnupsPXc6aGdtO6ad5QpouiR3s2
NxG/Edc97aFVgpOBm1WVez3LrjusqvFCN07F/k7QhEgfVcjZmrYwnEccCQSgekTalik0GTuWWrL6
CSs8MDecCi1ogGTj246MljSgJPUCixUAuhouatIXMdPT7pW1LKUbb4gPUoFM6mquG3pOJdFhQhyL
2Zx2Nxlyp0VKiCIEgS9LtiBA/Dh19LZI2aG1DMSXAVmWLrgRebYhB0803txblmXQUQgzq7oyTv95
LjZs446dAwuCfgZq66WrPURYtSrOGKOdKad6Ap/ll0mM3EH0goTfMv4o/VH+mxv8hHvNlXTk0I9H
PegOzZwhWgEPOLeRqu9ZlGDZSd2QkHklXCxO7xcDJaiRSc3bVo96ELvoW5IzTMPdjoDNRwY587vb
QeGXXWF5JJ6T95OZsg5uAj7X8i7fZ1JdJMzC5Z31IlyQI8ffNVE7F3PCJ0xhPdp09CdEUZ4865nH
VT6b+tfhFddAxD/yd+hXaLAelFqQGqa6UBFty0wawWWKyAhJMreTYhvTC0AAErtEMEit3iu8iWFm
7lmH7nIauqTKCSqyw3tXd0HwNct8SNtb3U7zQWlXB5v7DqpuzkaCbM/eU0yb9SyCTJu/Qse88AhD
8Y49jwPqLuTbb9JKRVypxj0FjyH/fF2klrPHF6po6MB0KDi32CZwvQzkj+vPzafSBi0LtIMet9fM
y3s6gCx77SJkNS5F3UrHWe88U0fs6WRvwQvgU6ZfWIpA9wZr6xxr5fy3jYROb41+T4QL3fmg1Bot
C8QGeWY/Rb3oePuSJJOpvXedFTo1ttSVvvFEHX1G7OcvUeBmt0bI21qrfuLVYxnthiGGwh7PW7i1
rT/lVnx1N58wtta4B8HNGgMd0K2PKOLTrrCDWFq7K3VUKklgnm3T6/g7ax8k2SJShcEaVsKI9pqC
Nlcq353JHWGsiHfK4///lBwJ4b6l1zCLlBqhZhthXCS3E8Q=
`protect end_protected
