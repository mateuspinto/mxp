`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
avjSuA9PaVqtXZTQwB6sx5P2oJ5wWYSDZYlziZG/ahchOpii2d6JBjUjodARTS6TcA+s90KiH4eN
pLQC+CDiyd/zd6HRdcPjb5/bxCinrx4WuRlBR0KnMvdEe51RU2NV7z36jVai31QjFJP4YlSuLerz
fUukYzeug+HSvFoPLppHy0hjtxQ/RatDuzmCGuRMI8mzw7PNhXtYoQS/A0CKTy9ZU2fILeLgqorD
hJv6J4qAoJbPSTDrGh4J/mYfEtLX2jb4qWHAKsDD65zM8UJ/myXK24zI+YkHa3ulefXO2hENIgcs
qcfnh9AnTFj2MMknmnevsMVxjswGGXvgqlJhtA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="98PwS0xB2VXMAXj27O7Go/WsUTcMdtEAXgQd/rHFgYo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48960)
`protect data_block
OTw4f697IAupU6U/qxUD0jHB0RbqgiEBOr2UzomOWJGGfx0m0/DaNxj83Gl1GoIXezQED4YIwSn6
y7SyEgSLYt4ayy/ZTnRudGe9xyD+lRfwPQvPFYF6ha3y5H+wWCm/3tXKzmlcwwGOpiFO3jA402CE
G017xtKC8F0Qpo0LfbFme42osnhqVohoL9XToxW3gS2IHmMoL88GrjNRns9Sg9+uNCTkiUayUKy9
jOR8jysGf/hVoVxtomAY2adL/iafxIpNcHXZzWAkzNGuOkdAHYiR0lgUXCOIms/cS7JVEWJCvahc
F0vNuvWS9Xc36o8TmsaLNgqipuRSrF2DOlOHZmlsOnKVyMbbvc47Xl0YodRh41mGu0t5qkEO+S3w
o1fzWPh8llL5ZfeJfh6Z+Wx/L4xIvYHU1V1JMix0qsOfyQFaMmsE0Msoit+dRSoCN0F35zoKV7AW
7TMtfu6/yZl3a09xLtamAA+2RGW5/aWq6OrGqItzFqUh/JtGcIZ/uYbIclH8fxZNi2BsqocZ55fq
YnSgKV8iXO2LvG8M2qe+C/UAtbeudw3uHNESyfc8/t8uNL8zYrVF/tgyqm4TsGM+HmkISiVVNsmO
T4IUrSntQif7l+4Oagc+FrEL9yqscSRE4ip1VINmQj8n8fwiz5ryUSb8HR9M94ya8aTScIh6ej3W
LN6LiqWG2oT+nnyD+PPdtaPPlnzJwbso7uRMia+8C1BJeoPDp2ctMoUHMImEv72YC35+aan98yKD
jzt68D9p3a/HtBlqxQqVlAbZmC9/ZxQqt42Ml6yNTMVo+wU72zGVEgIvkNxRL1VScoWE5ItZA6oW
jlztjZ6FT1EXO4ZAVLD9oAtPyQo1hM5JpqdBL57xFafndkADibnsX3+Uy4Zmw85+ME/ppSeJgPiv
fRwnkn0Akij9KssmjlmosFo/i5bnDc8fTN4r3dD/HghFdFSJqkScAX4memeX7d+Q5WW3lnEFOuK9
N3SKuoJPF2a0PpyJvYJMJxNUnOV2rauKyThVEJmLsW+aEhrYErMSW1w82RUDUEkxh58I+JwqDuCd
yfiRSSWJ2ZyEOA6wyNW6OlMxPKKuBN3RK/UoaRwB7zLt4a+576NLjJ20lCVOeZyDjXGg1oUS3vMJ
BcnGgm/Rgy6B1Zp1Bg+O6t05ITdcqHwaJWCiawBaXHs2+OiIPiJxhF1eGVCaz3M2c4Mx+iSKxdLv
csL9G0a6X8M7Ruog+Yur6qYBG/mkQ1DZZe6xTaAdvRxofJgYyg5wxuJxy88WRtOk+wJfQx5MThGS
bSTaBi68daN/0MjRO6UW3Y6Vgf6O+xWXLUpLnqWmV878Z2jNdjULbNMqcdhLxarNnUpJxKSwBYdt
a9fqIHAl1R5rLrDbGOdcZkNGfQCaNZQ+SUtUwMQ8RdnRqgvFmjHLtikOqjS+QurfTeQRDK0sacPr
DK68ctJM8NLcI4rSwjWRKzg7blq3C2v0LuJTJc7apIMIh3cDRXBEIoZg+TpUxa86QPtZkUY3kUWT
GgC+pasw9+4oqIuGqWEdjd005kdfqiPvfPr0wYMumu6RFBeRjdG+s312yOsCKShW0cYOUy1du266
sehmvHw+Namkf5Cp0qilhFOapXhPSnPzVJcT3AwdVNK00paEsgGUVTVh+do0YrLfREYuQvKDwWYS
K+LZ98D/6Ls2J0kB+wjrQ9+0O61YfdhL2lAJVGQa9ghK+VarbCrTKDF1WUqVjjZ8LAqUln3d5aUU
doAiTa/ATd+woUHy2pKfQme5qdbTTUj/sWjS0ZzdUC0NUGemAItx+uVxokB5xWU06heTAfxv+VV2
D32KQSEQfGpfaHeufO/HUc4RNBGzV1uV6u0UAC8eJKYJ3LuATxEZNAvCQNOJkY1l6mICiwzPKZrR
TuSeZknYTC+6r1vFBzKPUOaSdt+SRNIWbl15QT3hAQJY4MsKEXcUi/AW8l5HBI/KHrXRr4+Bp3aS
aScXhfXJ38+t1UtIneFTJUxclRKypR85zgkck3u4d+8pMGcViBGe9Gj0YySKh790qY+CGSXJn1Sx
/XziGOS6JTtJmmd4VrocuijZ8EDwlUj/NgWdAKJB22syPUPVo9RPwdJslPBQT36mwNHLnfk/A+t6
n/oYecs/nzqiFo7QrtsKDtLb8TP3ekpXEhWdKqw6sC/lxLU7Km/MYoQV5JO2TgSCkCWHA20GcXl1
9HXISC6pw/MAQTjQPGnZMrmccic5h4kaEExs2oBlIeg5EvCZbDRH5X+kOq+efF7vI7QhI9u5itsX
+4m9BK/W7ZGe55GAkfSTSDJoUsrZLfkxZUFyqZwRfKV9gMnf08ymeatfzOpFb6BitQdQ2pkJbSKl
7eMi8duWY45RH0TeVY2PdBrv/jPjAKbZqK1r4MNMY6kNTIh/SOrDA++Ib01s5GEHSADZR8b0Xims
B7Bdfw2eh3DgCfB1JwAen8sQnFwxlN48hEWQVkN8IWojQ4pCtftHRV/N6kVwmOkxj1bqfTih3k1L
US6CmFoWnodbLH6vaapLE/7KuvS1hO0CB9YfiVFDiMBvnjTdgavzbkW/lVY+TdH6rf0QcYe9fMml
YlOeaWA+phrI625YIAJWC+delMj6APYYeNEfNmIDUn7qySpFP880Ewtk6m6EfAZmpkDcxb3fxYmc
TaSVILy9ebfVpb6PxpqHU3X1ynq5hvGQzq8oGsaVu8JRyBwUy+ngxBRQV2X4DS7huc7HSSW5JRJP
qz8z/L2z0RgrfsDSwVjGn9r/kZHpYPa+bkqPS2Fj7Bgpd49vXO2meK/I47OjEYONpO/gpTKtpuul
C+9rFEiwW1GgR6IQaikDt5vgJKPQn8XrmMuE7FwWfjZX4CVXBNGhwjqkA/aUJICmNAU2k8EYLSAo
iSE+OPchlwDRssq/I7pvHxBbx4mgRP7B6+cMK6X1M8BYZA6WMfxTX6vgVnAa2MaZxFTBeJe+Hh+M
XiuqZEiKrNFp/o5RkcKC7YZDe8rztiENO5frMfCRyZpX7c7lU8CIKNvg/E5Ox99dnoHbWR2IKebc
e6lrKaGCFARmRLGgX66afWY9maQWl5g2/JOSC/gUGi9Wo45Fpluf1Jlq9sGys7R5gq7iNQcRnJZw
KziPpx2a38VqVou6caXD+l059zYsTl0nvRMXPIxt5tRUhZNxuJvCLsLYL0dZQaBVbkJzp4r/2OKn
ZiPCBpy2zQbMGVDpXeGbBSbhleP4Z/hMHPxv3y8Dk4VGBVlr5Hvnb83hcLyAbZEFE1i1ZPkD+2QV
0aE9ezwyEqytrc7fzsf938NzRpCCP2ea05PfiNibUW0AYT5KDFYM7HRo2azSHN5ev7C3068IZdw5
/UnCVgFIr1SJGULNVVuh/073Yxo6lspSf7V5VjewFECRiadHxKt3nmyYHktDXLIwkfrjlVX7ybuA
oFZ1gjVun7GWT4sQCgUUD2fhfDiOiXDm0Rd3UkJbnVIHKA9MtvECyV6cbgasjtXACw0AlmarKA1o
3J+WM2PZFCOA7608Z6sRXD2uQAwd35t2q5W45Sschd1mAflmUIrxI1TusEwlak/yXqy+4/Oy+Uo0
gbaof44pkeZOPPXq5MOI9XtaKHFsXFn6trZ8+q7ktdQfYEkeLwXCaM6BeeGRz97rORIoLddF+mf/
nof9qWuHT74u3BOaVYWVYDxNQVvUqvKEhyx4604Z0k31hbkvMYstU00nIkc2LZgLG+zqCtxXbRJQ
motX5+DHm0hZI/K+0DrBJsxsDuvAzfPbK+obwfKcHLoQ6nKE1Dkaf0WymquvUw40Ahe/QjlDLQ97
q82GR+lhTLW6DrmS7oclH9enqiLCMJQ8Uz2pbJPK8XrKAomLvrV4Y1F+0IYBfwSS8B1T9s++Xcd5
hc1Gqez6D+4npqX0mtlbpulvPoEFt5UK5g09/0dAq4MXzxZ3GYp6FmQKac2Hak/zCvhn2fE96y+2
ZYDUesoY/SzCMrWtQ2m4H5MfV15EgEyzV1LAm8M5rJoBD2qWNHujqYokkPuS6Cdxi3VXDexRRgG8
ozER4inffR2Tdi5cW8p5BB8wMhwgdUpWRns0uAtwB4QRZWqS2xVb4qfvAFS5Cnu8ycZSD56uA5/f
6naysl9nmee+HowFSWNn9wUqPaTiVYIvyb1IHfJ1HiwzryVgrUUQYpfv8kvMgX+RBhJRVacCAuAz
YCL8wEN1CB82jAtaE4SxC/QdJhEHqL0yNy2OwDoVxkAStuBJaaUO14sA5jd7vyPwwXLYEqtI32kd
8sqn9K5FcAEJI+IIIuYEMP1h6MUDVBuE9KGaCCWzXqDCr9/jB+4Eb/yME7B/1kSPfcn1UBaN9O6B
9nbY6A6nqfRtGxmjbNCdvoJ+FVzsl9xbCOwrlShtcZwEwrDiyhtedOLX1d08DZ+GkboZvSsYZnT6
nUMrDqc5zh83ETz+ezYuW0MHuvSGpZ6F73mcGQlPdBZZ22cyoYNNpj44Df3nlrf227S0zlzduvMQ
/J6nMJ3NDfRi1wsus3iby36LOCYsSgiGkZXPP69v/LIfVvqTEGd3Wuo+PCDpXU+tKt4bINeHw0Lh
nBbZ2ruZkA4z8pUVHdffNpXvVJfQV5twM4+GsXwRpCHe+afc4HEmDVHdxyRu9rDlSrSPSCk+OdqO
dlfFGvoSZM18E5St3aCxh7ifkFcDUWx3TduQVb1OMp8GW6NxVlZPtrV6wlEekb6lTht+cM6ao/TZ
7GHiuXPpGWPpLPN15/fgCcFqYR+RIRAukNvhz1+iXpWSVXHFGXkW6Jq9z2IJx+TUNtu3BvLReyqt
gKq+l++PPyGyP+Zm5a0rYYBxperbzMJrN5MoeGyNhFq5N33i4UfiDR1UP4CWSdwu+l+VvCn+XLHQ
rBLs9AmoDUt4nci2dEiXAw9NGujbxflXq5kXykWh5EUY0ObjRpi7vusBQKzjnBGOPtw6N+VBgJAw
RNDR4DYMuiBabgmcel3+TozyhY0TIphUjPl8EjgB87ye98sSeW0DlXrN6BfVxRL1KnI2uNzaIRIm
QpMgxaWrOZns9YkKvNQCRhDmQTaSF3mQtbIw0WZzuvO28E06NI8HpfcdUHleIbFprCVUbM2mZBWO
dTqplF4iJ8jwhTF/Z+c5JXeagIMA+zc0Yt+eveNojPJkcrAMXS2P7Kejm9KiIvvhlpQPUNBhAS2q
xgvdqWUABssGgaZtEaaATR4PpRHSRwcDxm7YghfUHL1ST1dQqGfTasLr2p1AEqadbnVVSL01rT/T
dkv45O1Pgw5WL2Xk1037I/14RX/jeZc+gPBb9jNgVedkTKLu2jcMQT1chCiTh08fpR4ovmyLtQUX
R9KxzAPPKOSWtHIuzgFWXL8FgsxX5GUAlOZWiGjKR2BUN00Ym93cHdVcVGHaI2Q0FSJ0wxn7t6d+
aSkTBBBGJnC0y6Cf5z5qFqRatBbILxOiCkJuqjhSKcpX9ydM5T393LHLTn/9/mHzqDSz7gVObyOs
zUD5P2zd0icc/sx7XBHEqB18iOB0mswOeAn65Yrd+St0iYZbjL8bOjvEq6HqAe2lzF5Hf5tXrvrQ
BJTW7QWKqASbvOg0M6vG2c6dLn6C1eGm0/Gcp6RTKDq3l5V0AmGH21JJnhXXnmtaGHlsM4LlpN85
tZuWWd96RyVJakzdJnry9WvF42CGLxJxhxqKOhqXES0mAP8nwbEgBOgFh4SOwbH5PBFoniC1vApv
0OYaisE9wlMqgNesZrhw8QCBddbH3cg4HpETfNJ/lhnabDqzM9y4wGNrq+P5W9hN7Sbk/Vhy7lRl
olFeNDf+Xyc+0SgrsPrb5u6oIi4kQbwpOAofU8TkmhmaTq1NU5HSuA7NN3AcQVx5zpEG+6PJBXFv
HspDEpdgSgQVEx3ZM1bjTEVk3BKrfkjn9rofcjyWOcl3XMTqyal6/onr4yeNb/aGPLSKfmPCn8mc
kR5Sut0cj1oChkqIUXldZ4opVP5PeEfcVnaeYtfvg69uR5Qjx9/PJLTwMaTwR7Hm1//QPHrcKnAB
1Hw8ciAUsEtNB5Lpf7GbMLsve0288AaSd4pFGQbToexGbEp3kzfgSyCu3c+qW+6pYBC16GVoRkwa
/B3FPasv+8p1LmEz3+YcsF1+8oPoQ3LEj4w5GbR5vkWsN19BrnVoCeVp+S0sHUMdiMnXYUPrnjRh
D08KHRNimdV70Unb0t/vtdGUAOeYclbj3MGWp6cuB5EvquP/WXV/CZtIn7E5sBhGlkMwGn/1Kkno
F8bq0BvDj4mCpNqUB1doiqYVk0+PGVWIiwKyBBPBv664a8ofktN/EilX8dE5GNAIctgW/4N/Ilhe
kHuCt6hWx2/6O6YiW9xFrbDF+4pglORYQlS2+fNX9HwFSWPw4vnXHJsvc43k+xVOQ8lJYz/sv8a2
6B1J6GAkhXQbWDxy4DgWzwJjCVAAz4i/VBaYYts7rVgNSxasWbIlvw2PDrnRq4SCt9eyK9xa0GKN
zvzs5mI4Eub2PN3znsvEqcsM4yKHHmzJ3OfoAVROjs3pxG502OrjOccqVBgdBPZts5YjDY9cT/G9
CpGWhAi8VuPPNlBF7qlTpxmpHDEWg1/dygJtPO2AveoUKzkGhIS436XZnRGR1+113YWKnTRQurSR
yYbeMbI2eLhgQTcFKYmFYpadlRC3F8aT3BUJKXbVn9eX0OFAyjRafEkC7g/pv5h+NanssHmMNWvw
8CZetguYtx3vZgS8Pfu2UU6Q2h1PLydE/csHRUrVpepCcEGYcvZ/Iq5NmLEYYEJYw4piQZxosWY6
vmJMnnGcnnhSOdeUM5/8XfRIOffTjI9EIdZYO04uVjI6xm3VbNZDl8JdK8EBB0iA4P71bc/BoTQY
hqM/qxoUwoe81HrjmNi3xdyodD+8PnpnocBg7yb7PmFnsAPKLYAchfN1ODQoB/8xZrBffYGWLBX6
GyHlHa3BNUNE6nyYH/wbmeVB1FLaMf/rDf5XfA4iuVsnoeI3ABl84AXl1C7m72phdf861F1wODI+
ezVdsIjatHyzhY3X6ilLc57SUNhg3Vkmermkm4+CETecPDbTO50S7LFzYrksk6eLSxwmTHuqBLIy
52cnqTqEF1dcHthimHIuTKGNGwN9+8kFoMaE60dTRhGOo5jofgT8i5F8/GtEKEgoCnfJP2eSNPJB
qNZy2DTgGhkFMk4JuvFzUktMD8NUoZZ8tNbrIJSV7lNJlT185P9HaVSrYtB7IMpCSV/T5G/0nMZ6
r1jNmIk3Dz6RSxAbObGYpb+iNj9c7vAJKz6cL4I7k4xXUm+M9JEDo4497Q815M8XR9m+Rt+UhJ4N
xgSQDw4mBxq7mfM0guEv7Bfeiqldjst2dqULdfUs4tQGevt73rg58Ci1O4KJV911kVW+m0iaa0SM
X/4E5eattlr3YLN6nWkrXDu214Eyzuc6z17PEgbMiFOYTmaWzlCoGw4OacdImPsTR8acFiO+0qTg
srO9MV+HknwZc9ipPUVjxAMpxmKYRAta3fJnsE8VJMxpCVTQq+njCxgmbph5kjijk8gPFtzs2TZo
vZn/rcrzkteGit8XJtu/ey+KoSIfdP6xD5APvEeOwg6o87cMfyjTg1HA9vNxOqnEkPwZS332uJjF
AwPNneAvUt15Dt9TK4+I7M9Plt7vbq9LBZ9180SUgCq8SRTRIa1L71LhzoojYPSNVIUuiS+XMwcE
gex6pXyUNl/u4ZpXVfXpTaOj+wTlZntUmXMwrywQX1wlp+MYPr1ANGY7e6XSS/5/Rot9wR2a3HbE
I/u78mgxhBNgCSuWgCnfAmIdN2XzxiV7kbQk/fILcex/tzr/JwHaA04RyW947V/HTWHAfcST9A8p
Bw0YGOi8Oaf2Jes+zSCQmSJmS/E0yrd9Rd4I/jHl+jWD/livc692/deBXp3RszTwYDwATqYpI6hJ
HNRt9YKi6UeMgJODCkJ6wkCoXt0Y6WVfA8rbnyJ8LBObdxJvNTBxMTqBDtwX1MsXwlK/grdRloLl
pxtkduL+HmfqH487r1XnFm1SOLJ/RypmIYm6Voe0R0ffOo+RmJaUFW+CVM64WEQ2mAHmDx27fJ9F
c8ubb0rxJOqeD38vW07FafJ0jk6wBwzZ86tS5W2rzKc6+LnzOFdjHYNYsYFOa9pc3aVvTAmxluFw
WyrnWo+rbMoAfWgNKoahH2Rbo9Xy1b1qq7iiVsgZXH19KfCyrxFQdvtQHTL8m+7ZAt3E4GXXXQc8
uxVwz6hNf2A5pcSOWC3J+gEtVrvfiPhOJNAdIXRcbhiZdIgoE1y1djNNbStiMWyW5FYT7+xJ20XN
sEH1gc93k16dhFha9trwyAGNxDNBywpzJqZhRi/yyit0RWb+raaYzB+sIdrKelDUww9Z4hGZs5/s
l69H/7IOtvXQ2OU72rKb3CA0iHTQepWl11bpZzjeRibICsZWc/CLg4P7L5/L0z5IgL06Prwkyfbt
tKi2y+5aO8suwOigHtd6TaV9zulDZkW/D94CSG01AtXz2czrtFWgOLkHrzvbox4D07ClJw/UMXEt
1SjhiIHIMtOCEGzCrkqhSmfKeEsXCecP6XE9YI+GpL+n/KT6J0uEyrKnKrRLp51JasEntWorFyfn
NdW1B61t9o8oTS35jm2HDo5+45E9xeLHv274P1hKwalmFhtPe7iCEi7jcaSiQxRjnun4tDM6Pafr
Ik3DkVjTu1v0pj0W4RJ9fh5p1kE+fHG7kT9oE2MyQCG++6j8VoAgQo27zOA7PMnH1Ia8bba548dF
TdLruUJIaHS/Pz+gSktQfmX4XdMoq96qBCsHgOqGpOyYf9c8WKrb9G6WBEpBXNepPSYpBy5Kbvm9
eJgMV7BAPhbckh/GQcXcnpjzrbriv0rjXj/ovu0f8RwLM/s4T4lPDRZsIAhaep6BftCeD/ROVtgp
+OauiuiVj2z/sAqablHh/xHZ8rQfCSXrHcPvutWhPfaFLNSk3Haf7Fa3VddXKPt9WkXj5pWa732H
is1pUyhnRPXd2HNDLFaN1rOeuZWJka+EjpHr7K2tMw3mORAYL6jCHqsqdS+ac9Qvj2yu1t+zJHO4
ey3DC/WYYjwJnh3FQexNX6q3qpxcK5nZH4F29iAv3ZizyZ8xqRs99ZNxZf2VoIb8keFQiUdTAzMn
n6W3PMEbp7Plqc5+UMl1RW1Nf4gYGyXdYs0EMsC2mK/ck7+F2Jh84PH94tgXuzbmCIyCxAcHH2ZZ
v4sG8sMEobB8StgrAPH46bUO6K0PPyDaK6eesI/LeeaedwvqosNeTClFSxX5nPeqRpSCLWqr6l+5
x3oQNCxyaXfN/9FsUfh+/daSUkwWtgn40vAC5Rj2JBjOH3EJ/GsOwKxt+dID3PkQNbKM1FzYHZLG
4T09b61zjYrsyNcJoX/5xhy/3YouadQyTf45M3jsdZyfmzcE2DUVp6yYdgGdkbgTfJw7gowD4Qyc
3JkyGkR3QJsip4GTtjM4t0lvsDXsA6bsNPix3wsY5NN6nO0qP61A1v0dtzRS4ofhfVdV1GZrZBJE
NA4kYmMAdU5VLf1CV7UxtgXoHB5z7jbcJuQkVwJCJtSTB1XLmOMVSaW/7xzFBpjuBKf1sbDiwCuR
hFB1ytPDTX1Y3kKIlj+yr8qmWkmIUdEKPT9vVDXNAS4Gl7byY0DLOoQlCEzZ93RehuL4qhlD35vh
jUxN3w82jRcE6GdiMcLTauu1BxzFlZFximshpYL5oUmRDhVZ5rMjp5MNywJdTDrblRF3unGwNF31
g48vRZSg+nJquAfzCwia1gvgW3zYSQo1A9VbODd8XfGQwr/nRtI8swy5klMVUQl2dJMuXGrX2cve
/6tamZ+H5bFwJ02bpa0d3LIGs0vgPJC3OuQ64gZzFUUfz8y8GYbNMDzrTi1VV+Mn1DAcFv1WThj2
eZWz2tNoHyMo9tNX+KzB9isAG5ECghmwFTYZ8xdDJ9zyte1St3VsxxMJwJyVr/xtnh698V83xGay
Lxofk17TC6O3uaLG3+ZfRiz3B+gDESSHvECgL8JVjqB7l8yEdGN1k202GLuGZlynxv/MXVmg8Pzb
vNL3rW3tSpwxOYCQlqwOYFVjJPrXTpwmsRP2/dNm+NDvKToELbl9NMheesIX8vCrhKArH/Tl2tKv
YMyUUKV/l1FjkWgcj5/Z/VT6TTnkLijwp8QPD2wdQa3kdwcGu35OXR8W8LRJ0vHeDFvvgc+bQ77q
mEgrmpEwm774i8gYyvfRj9QlN64+NsWpl/x+YHikqtznI0E4x9/yPmdfllM312Nlnij/O+kDz2Jc
I2E0yAlWwEtgh42xUJ5R1sFDi0yJ2+8ePGtsMiWRzuobjDBN4HuJG5tQXUw3Qe8mk7Ux3EfOuH5E
NeqPM2eZ6fVnBW6KAXLRk/YbEtvgI8votn8z/WFr+xvzr5W8cKZ+HDFlsdrl3ZZhYgGrsotdDGto
HlMNeI58EvF36kd83J7umpi1PGRfJnebjUaEBRfETi8XiqgtTc9bsysW2qW0ThHDNz1kIDwUygff
Gsit7suTOI5lEROivKDQLu6480WrdRjc+ncqic/XPGafyNs8e4HghzbXMyiWE0f+LH+K6yBFYUCG
RVz7GsVwa84HGrgPFyrczxDLEfcmRcaMGjuw6MFkRZeq6rF7QLENotrRF5LDmRYYGiuIpXdSGXbQ
Nns4q7VryyFgROy6LASYw7JqPF9tDvC1j1kOCnGwb7H5zB0ZLAGQUJslqHJArwRuLvnPScgd0rNd
Q90MUYG9lGOYAiuP40BHJlQ1r1L2Av32zG7L77F1PynDzPrhx7qk6hR8CnHZLOkXHw3+qFRAr12U
XWBsuZq7cVUtijtMwuHv7uTj1JQ4KP7TYqEo/4QwbOZPRz3PQ6vsPC8axbXol97WuOL8AE4oCTXV
iXAjLk8nvAR+C6FNx3GG9yqXzZMacmyR4sKNZt/9dQGXYGpTVU/xnrnatFN1pgEGM6Ayil1HJz2h
gw6LrBPHs0SbOHklpPyS9JVINJhJRn2/X6iCerWVvbUGTbExCk3Gn+MxofXX4jzeyqpn7ekqP9ZR
tFkwFM55pEmOpAmHAZ1cuZ4DJ1Z6ueSYmK86jqaHdLS1+uDvIZqMY5CpfLn6l/K2ET/Yw2bmLdWD
LpJVB2n2le+ePNXI+IB9fJGVrEhHXpV0LYW+SySMYISq90Pku25biIvMVb7s4O4lpwWHMKVMltWW
6CFdStBIU3kcFNvoRfVOnhKvUZPot/gxDYKU7B80wUHfki1GGwCud2NTHKnxTlHOQq6j/Pwup1XC
UAyeNEMJZQcwULZlkFIynthAtD0yVZx2MJ/GXpPM8RhT9zMw4a4OIiPVFfKItUqTrgj51IXVbM3f
vClJpi8zvApvNpaUKv7azMwJKaa7DrqBiTR3OsqhSsc3FiNoXmgQN1NBzRiuA9UquP4DiLgK/5Lp
NeFz7D7enUilAyEKd2/3GjB5ORvD2aOC8LiYIA1RRiYpqmdpPsNC5Yinq/tl/qSzMnQ4BuKvFzse
WrBF8+pRgQ16YzMPgXalRLZ+MCTL3Vr8MlxdcA52AGo/5Lf2dqpfglwT+7UwnD9CxY4i/jOUYM0E
RBRiycLjF3W065Vpy2Pk7TdiuXku8TfFw7Ai1QklObu8SRIvwJ7WrbeWAtxJsDpc/vDzVPTtRiaA
UdCn0bex/e1yE02bYhy0drSGvGr3iysdP36/YhTnqCtKQcv6ef/rIZi49xNpJbDYWNTybl+enF++
571SJlfq8TWNXGUebzxVy1l2a/bWcfQMZcIvbSB4rvXUowgzxxTs/vA+J60StnXR9gpENYWXkctX
EcCywF7O8+5HmhIGKdxSDQI1II1iUapQlh7imvMpPMiMwrd7nDo22w0DcyYgqSsz1gai5hwrfPpQ
gVD1DoMcfTKr/cVhYn9oMz3abmNr+LVJcMI9pnPubPUsYQGqc/bK7cfW+ns9apNu30B9M4JUE+tY
9LOS7ECgX1w3Fu+v9uR1APhTo2oC1gOcAOh0iprGWeqTUe8qNYn9itiJZvreXmtKGiVUpCp1p2QJ
/dhuqn3pJmJZErzi2I+jpGK4M1tQswOPkg6NB11GRhvEX1yJ/udXpKJryAO5h7lzAvskVOqEAtN5
nocpFzhWjccP9s6TnspUNZiWrvi6rH3dL7X7uewFl8/5l3UVwQDRDpbQU3EHExM0OvIh86bHZsaE
piwdIrLD2Nr3m4Pd0rNCfwPOvObxKyhtt7WU9p69pl9Oa4apip8fLHewIVAKxHtgNoXU4yMum8dY
oKpgI7p39P06RggN7CYlhDXr2AWdUxUnJydiiGrSrJqMXHYLvQhsevqk393l/ibUBw0MKDDvWt+D
dgupulqoQfE6K4B2qVqev6aIl1Qx8lC6P14VwbhN7wV72CnUkE3JTQBupoEqGwbKCU7rdNenyAGI
byEOeJgxVjhCy4qBnkn8Z1lcBsHS+k6/r3HO9QUUUv2yTerUeKNf1OM3K/9fhC6E/NChyeHuPs/B
eTvUEZ0gNpO897wlxmcTC7icejsqQ7G1oUSwMhtJOTN/mu8/l6M5i3Io2zY1P6bZcqoMkYWRoYnD
nOtm4lkQBN5ywMVtCearmRstbSdJ4WhYP2boKtXSc4gG3XUlhR07A8jOj+LQ6TqfkamQ3+M64WHy
/lMkNUP/enKBdTh9siP4qysRRfcXOimUx1CksmgUcQLO9CEEvAlLYwZpiH8mroYsjMaEu6YnOk//
69pIa1b14KD7j46T2azNbSLLiSgw7O+Z+H4qxqSyek61V2CVOfldK3O7ppc7QfYoQ4RjONbX+EXY
4eyrxeiN6b/eBsU1rGamHgpigdQ20hDFcfTZH+3Oypb7O1nuIB56Kq6z4tZaSwapsO+0OiSbNc81
MzJGSCSjwtYtBvMAglLfu1QwJa78IqkcD6rfuBtUkaoctPoR/3cCjjWPo49wqnzZYLdCKwr3E3+Q
hE9He5ZRFfR1wyKUaOLoKYEcDx5dYbIuXcbka+3Rla8Rw9xbgbWMHI8GvTj5RFU2EialcbZ75QYb
XvHca8aLjy1bCBBXxWr/A8Qbk+NuZOeCRP/bL8BxysGl2Z2PjDBIk+06h47picPOLpzkqAZyeTUp
F/2pKR3swFZIIvTXIs7F8hLB5akfdNhuwVvy6AlfpJ7tcZPtECcEjCnbJJRQ7UxFDw12wieSfKvV
fgccfD8qCtPRK0e/ys9X8S2XlmL2yOKhpPacTy1Zt5hdi1OLyGs2otwoO96GL75pnA86mm8bjl5A
hc0FXI5UzI8+hQwsbqDZUYPFlexSo8FriQP2hE9Gw7vt9y5j3a4jJjLSmS6oBABOFgVhNgmDom3S
IjFSy6fx4MYc3KYC3uwhTS+YU3hwternI6Yn7qOVMbsw8oNWpABL0abqRgPT7rcHRBOQpO8sgqs0
c5MDugN6R4UAhSASorLgVhI5U4pkBJPeaEXO79F1z/rG4DyxyjEQ0v1+qIQdNhL5jpwqaYNN3aGl
nZMEbgvG1y/CvaX+iUsj8dgnarBW7OaHycvnNNB9lLlqoiGF/mYNsARq3Jk7UaEpQ3t3jhhKUFzO
Py3sAz85M9APnHL43zysCqh00G3Ix0yzUtNXE4jAUYhTvqvnQAT661qiCfxqeEIwgi3pTsajM9Yw
wYyoveIqCFSYJvAkEOh0czTfNynCrvAzjo19A5qXu+eJi/WsjJQDnVzO/sU1M8k1wWEYe/R5eP4W
RfB3XYoFX1gIcL8M6/pxvPv+jsc8L/mhNYnv8HV0f4805JPylNhNxLTodMw6enWxCBK8ceKrJfGH
6+BAXQNqqoaT1vxFSuXTAJJQImMZx2NfD3gbs7T5kjGAbn7PdkRbkUazLMRxQ2+DvTuiAG+jYSyv
3kHrLLLJmCHv6DmYdwiOorQWtqeTZiW6hQER1Uq5t6CMXR6eLl5lh4BvKV5Zd+k947Go379HHVy7
hk6AaIaBB1WxC2uHxf0gUev9O/2ptNppnvQ59uZQi5Z7iW3+9LHx6UfG/wPz2RnWj8ZngUbg2rgT
PD5DDJEPdeGBcIavkBROvH/XDvU8qKQYhCCv10jusGm4hLNfWXwHXK4+3wKG3JujLrACSo3ZkGww
E9YQ3vIH+1ZWsASIFhwyzaM1XLjNuLntZ6UFCFD0XV8jdscXFVe5IqtLfwNJw6vnKee3pweSpcOb
wF7UCkDXEIuOXo1IjtXQvgMdaR4vuwxZwPV2BXmbqIbmHJ861u5fkAnI8BEWXBgH5arBUt8TsDjQ
QXxx60jE6LV+LqPGlWT+3eQ4C+wfZ+s9DJGiEQkfUUoGJ1YDvwf/tw1deBXsHxp5XmQ7O7Gqdw9b
Mo2eO7OFC3gYijkAzf/lYeia9oZ5WaNJv+rUDbfcQ2I+5aAd0QlLaUBBA+Pqfy7PNVkojsT1B3Zn
OObiZ8g210p0r2JKU60FEfzdDT8EJF7ZF1DT4L+tIZUqJX141/4GOKC6dTpGP248XmUOVodVDIMn
fXJM/ZmDjxj7ldRn2yO9myJ8NvmwxYLvKJiODlVGfBFCvXqLlQ/+Sio63Lo8sBVyT+jDwliK+Rij
0wQ7OHCaYdVcgWd901sRhha5QJ7iVMy5+v0yMbslM2cynGUQJVx9WVYJf9TdwgA8KuWBgWyYpB4O
oHBv6Bah9wbznvScBBijvrmwiGuWM9pLd1dkUZviajrQcmJ4gfZtnydANklagZi4lvWfRbR6J4SB
rs8ao+Gx3U2b0ITlYaxZOx2UYS5vme8WucW1cOKEJvYqZkQvnO0OkyzVsd7rzw4bW4HakzsiEqwa
Ro5gaP+l3Bjp9HQNshgj0BW7Woi7CLPxbAqYNVh4VCq/EOE/Hc7Yf8C5nXzEmn6usrbbFsdwzJGz
xnnsZ9mGtdNAAcIRKfvRqOm5usIQv1RQ7jElwtBmgR2++ig/MhKwj/6mbd9DepkQv8AHTjcBu4Ot
Y3OsvX8Nrr1NyX62icgdrI5vqfCg3sk3GVWSf/nanVnTzSWIjoRqB89n757JduBNTNR4z9N1562P
dlSsew/9dFaTfCD7xTv4Tb0gSwkF7ayPZewMIXId+48hL944OPdgmekaliQquxM6sbpnkrQiYSf4
9NhzXintflEFUyej6hmiE+fZeii8r6wP8Q7CCz44/BDiIRtKqRlZ4ieZ/H6XbOS7XIswMUBcX5t/
N0zaMhmx0t9ZVOIQhV20OcvMAelfiyXw4TDTmggMo3YLEexdI9P/B6Rl2hHBOOCAwR/nFYoLNUv3
bGo5owmc8QQ859gizIcdpa8hkP+g9ArS0g8UwPJEFChn3oa7jibYyV3Yaer216ot62Re7mppSlfz
S/RJ0HYrhIPhwVTZYghrQLnXZSvimgXqNNU+Gy0JfOgovST9iFhWbpzjwrZs/ppj3M08mI9NHism
NdzRT70Fr3ERtLcGY1CMeeX30i9P3t0tW0xPrL08lB0W1TXcPU5DGdrUpUQE1Om+PWIwpoLJV7Mc
pG3SM3IHwewaxs8WoSiejA7fVChPmL8Z1gqxRAWMGUakv5qqbFYOj7GyfITc4LBZ9UlB7N/JNbYX
c8azQXISZafU6kXkLWgDv4EIPNstNya8NAaIhHqH5V6Q5Ng5wRmDFV/U3dxN4UXAM4+W0pOhEG0/
SZwa/PQIvSZMoXlQ38atlEdqBbz1Bdke/CSV/A8Y/x2HGQCdok7ZWaDrjQZm4q+DEU7Igdo17t/s
bLpU4Z0CWqrWB8xXME4yCZbHoNUi6Jgxcans4vdUVGdooQxbKpNk+BdTfRYnUn/pAwvKIkXFQzmo
pbvWR280mx18O4EMFYTrp5u+FgQ+ZZmYtDXaUnG/29qxxvxi3Hsszn7FhjCrWHyG9h+XLYYxhej2
cvNvhRXfGIDvD3dWct3z7vpLGt4OJPH8bbuJwsB1/xh18423Pbl1lH7QxVA/MVBFTwAIU3YOMG0S
et8sjxcS8UVA/lklB8UioZh94PxeXN9pBRyXt+kB9kij7mpknM3yrBFxoRVD5/nL9Mvy8siriBeq
uFyqlVt1sdbFOm7prWvZx8ZVeZvisl2Sea8Ubw6s3vhqiOwBC7ux3NiqMyUTPzqoJHHXitSbymY/
ipsJsRFWNI7zmsdDRaaKlEWVgNz1zBk0BKNA0oao6r0O3xPuEZyiDpQwZhBuxfYy+j3j9Hcr6Vus
Pt8aXYPDx5zlbhgt+Ulb5vOeFPwzqBZx7rsPlm1Vvurzq1eVkq02ma2MzttmHf3DiJVLLHW+EulD
0LUNsGqU5IR0nAdF9L/1/hfTibukU+JtmZOABr8oe05nvNDy7G8C69rxUskYxPAqtCnUkfub/L9A
6onn0jlcFx3PFTOPNT5mhhT8+pEBKgkJ2duiS8epuHBYM1FUmM5AtMoXHhj68WwtruPy7LjtrqNr
0f1Chn/7lTuNwD11Dm2nwAkJbdg06oNZ6Mb1DxrCm0zBXbS4LZ9Aan6tJLhtJICtAYtyq0+yXa8y
GD7WI1j8c5YRlhFwHX6JPv9hAtSAcF0Tg+QfARFYi0WIp7m0KjuwsztsfoOkqQ2L2OKqdTFkpVUb
c53ITBBw4b/71dk5hJ0prcbHAGPLbjpYY/a7aZEMRQEQ2hFx+ELc/7ijlhbPtHRnOgeCTzww9PO7
Ual2eKOrNphrlGJYFKfx2fh9XQuh5e35I2Q9SGDlHgCqvaULpvDuCnMnCvMe8aT5d9uaa3c5YaEt
04CuTH45heBSk3DytKLFBMBaqy8oeiWVaQZHh/UdAjGcPT9rs03oz72foxAKBGbs7PXVyy+4WrD9
UtIAQ4NCE5fyPzDyMmr6I2+2KAvuF/lJRpHOFKa7qc5AgYAQZMDSqRV6GRPMaEyopNbTS2QZpltM
kOqalW90i/BV26lJniNarEybIWXacEpUiTPCeGh33kMYDr18gXVRYbmrO3yY1bUJsO548kwJZpOP
6k0HyOl/3cgUAynEdRfC2kWe+W2wMp3ngVt5PFJKC+TH7lxxygY39aYvMyENFo4Cl6LJwvfHgzT2
bEbU/s0sWxHp4Daky39BQ0BYMIaMRMwdSYf1UFNognHrLs57NyL4Cje5oPFuEZWolTGwhllIU1jY
nKQQE3yRF2cM8ZZO2l0p15YrPe6Ub0C+I6uCct6+WlGBJ1VTmPZXeAR/mwzUKRDp/YHikOUnoXy6
qWkX2GGX8to+rxXZQj0WKoZhjHaFqzvbbz9r/CMKwmtr7v+NeYfyU/Gk0FE7H5fd+6stIkeOPFUJ
WTABD6s1SatljP9Tef54C2T0hjtMBiS8//C46DoaqskOHhgISGgzj0bIieoOV/reyyBA8Nr1Crg/
Ss47RNAXu8CLOCTMQJL5015W96uWo/EAa94CssF97O7xykCDMht51N6soCieIblyH5OYYQdL/LHj
THfih2uanPa6Mtc6qdkS+rsao9qEKDNvN1xhdHjzswRPIQi8wDPYQZ62DhOBNmkLa+c4+CR/+wQC
OC6dsJuAMYjSq5oGxaxCbiFHlu9sRCzSDIlsR3TYb1jo8Q+JMYzGN44Gt6WslvqgclsBoFZ8/Vs3
XuL1fIi8tenADB86BjHTvvb7o9do+/lgoVGqsNXcHJq6afNwAbqQ6ocYiPZ5a6Nd0Gh2e8WXTs5G
AWzge8/LRAzmHwBdqX7Gf5FzXPI5NeLICVMM9A0qqfyjkV3Y5FgfrhfR8bW57LcJ0yGyHdMOMpgY
U1s+sadfj2x7Dc6WCZupIAb85JK03eNzYtsBepQGiKjvrL/mD02odyO51nXHfn8GKbD4GylLNADl
X/wYjzdVLjyx0d2QfpaNKNxM4CDe7Sb2rXXI7PQYPWiMOF9UWZjmWi6GalEBocBPCUwu9Ou/tzB7
0vWLUAAmTF5KE0XlaH5pFfa5bEhDanGV5YezABYH4Uf8txCthXGm96QWVe6dARSpuhU8M3LiKsIn
KfHLN3ZDMRpbjnP8Tspdi14w2fAFZxIt98DIsfeE2A0TIx2YA6qrWKgWxBss3dDCyNhencHWYcYM
ImUssB3FJnZyqgDE8w1zZu/b/nAP/jSBP9JVkDpb8/le/EZNx8p7174e/I8CZWxXlRV6o6NGn7LZ
Ke6+NAXDyy2TjMc3SMzoasDyMPuJKW7j3pmu1WSJbvPMImGcj7m07eEdhNep8JbEQqTHp+P6vsKx
4QgZR/8zKRp+4WXSjgNAz7fyldBlwa9aZhqOZrDqRPuTdq06dmyR5rkesMnLd6w5uUYrBqys6BTv
Qi6DP0TVdRN+vvPSytLR/9wpzQDwVxCQbUKKCptlJIv1e8o5w8ntHqITwWOzTpIlXwwRkELSBxnX
ra70L9mNFWE8bK5snJg3/Cwo7v8n6j7pypAumiiHVLkw/qEnOSL2CQQevXU5Vf6YbUjqD7wlajya
edDF1s4pEAOm9DFx2gOT5qyFgHUnNMob7pFX3q/8rJOfkKh/22YPakxG2xV89GEohhjisLzDISQw
dOVVI570da4UFDQLkY9Z83jWDLd8hcshKOE7C4m1/WmjuAeVmBQd0RLgo5oj3QQtt/ua70bKw+xv
18h3WEiZvvlGZmzpFVP3ZoiXzMF5+C3WJjF0J7HgOV9+GtE+HOMr5O2+qcAPeZh9UIX3JnJT1DFA
FHZv0U3zBqFRYRP+vVgMszlRTUAqjXQRLcOaYzCsEhbElEcTsvwmctgS+cEGaYZ2WObd+kXv2IPH
vPNRTMySXg3/rMsoPkvnDrMIeMylZKQ3ZqSIKMac8PtnOvH6fEwXFASmNmoJRNp4OzUynmfxGfdU
zZpcDfxy9gCHovJgR9spPcQuOym2jgeAc2mIfe4EEg9CcpleBrZvxE9hDrSHVZ/xQ5IeHwJnHE2K
waSl3KMnTzbl5UJ7n1FZDj74TD40keZ+tPOBnWIFS49NWo2sV5Erd/iO+FanYAdj05zKfDUjj+6r
qz0fq/iU+YZkNNpbrc/b3sPLIuTI9GcRnSQ777lYm7EPuABrOg4D725xppXeVwJGNGA9PA6ZgFzM
0xSFLthcgsH4OZ75G4l0jcKL1dKRfdtrke1HFJ3TzZtFodvEGXA76z5kXWOLNh8A4+d8iB8jjrO8
jt6jJKC6fYBL3voNupGXXR66fha6fv9KULHcSLvkAnY1x9Zqgw7UzraxsX3RYuWYj2lsQKWSadk+
skhPROxEyyTdLkX+1HmJX0SNk92zjm4gal0fOqCwaiV+BrRCTeDdL4GNAAAiVWcAeDJZY1Bp5IqF
IEcRMX8g8tOrVOETDGNDZcwAHcS7TMLwU8OFcntcv0d7fMs102jD27yVqnhbEmdTTqa8ebebpLpr
82g5WFEwPaL4kMpmzAXvK2siqnkgAKbDtpiTA+jifEfXYor+WcJflFH4/JqJqZ6B0kbNxLj+hv88
pUOCXxbxIT24c22fzXK5oGTjcUEBKaGsAHNyGgV7BB7AIRgT1KCxE6KiS4/he8K68umgdk02QKbr
Lwbi1ylp9qMlBf4VFgCHFFB4u1xvG5qe3C6D3QZkdQ++BFJRXxZWD4m6RdJi9MbosppxeHEe7lj3
ndubmt4oj1MREOlzFwJ0VvrWQ4NyLJ5e9Wuh5pFU/fryTMqNnmH6oVtzbabu6W3Gn2bDCQwsf1sr
kS/WXsh8d/pW0Dn3/64i7H4VEmNMfvCH6m7aFurjhUtVRIGi/t37qGsk6Tlpda7DSKWXhdb6F+5d
adZMf6ljinBKJxiWGIyf7Zn6V+TUATEdG+4li/RQt7AxYTA6Xq7xPj1QktuFmvva5XO5XlMZ+hx7
cwH6pytcF8n/q4YFV93ZrMPfYM06hMaD8itZSyXCWjKoTF4eZV8kDvsdMnNRMCgBrk68S69+bamt
jJDLFIe8JSxQwsaZ1DSC4TcgkNmocfenN4UMiCutAjVr+NbioZmBZlpt9DVKwV15cHF+IGXsKu0L
VEHgNG4TAcgnkXIg83bBMP5CBjpYRgnP8LpcuIakPAXYgeNUPlMqoPl7/F5ju7h+7q5vVBssgJrS
hMSmIMIf2XcRNOYTj7snSPL53ZV361zo2SVFQDfLqCMYe2Mlb0LcJx0HY0BxODhw3WEW77KZxxJF
hhJfW0/cgIKc6VJywRT/utM3WTByOhB1trQWDz63HP30fTAEgSEwoFdsDAsszs12KotXdda3jT7j
WE7k+CZPXhI/c0FkK5AYRjmRmZJThpaN+jh/DIC53lgG1orXrhbWoFhIb+i1QhDS0g9xrRvmMK7o
7VExWawzSCPTEYfJhGcJJv9iMG3K0LqrBjR+m23dASIPRTnipcbph0i9FDur7JplIIILC6w4Es5Z
MgHUYI15r9NanTWBeudquMXRc3WvzCZE14fMewoWcAZROTh9njP2g7GDouVqypXYMC0tYwKl8DnB
GjnOMC9TYAb8wt3HyB2/oMRNFaDW3MIHTxZ5enwPNPBeKLH2BqdfeDpftXo43RppcfmYxUzAwNO0
cZsi0GOgvCXOL3VUKNQeYrxP/gNYFEPgO2iecdmPWmYIcVll8LJ7n09vQESQSn5KGwLR61u3Xp88
2+tijcInA0JiewL6KcRxN1m4RwTTE1fZDEBC1TDUKI3/tvLG2qgjfKk8fHeix6B1RgaDh1s/h3M2
SHnISzj00fGq+/zdA4XZ4e7GUSpeqVMVbpGnk0iKh6kXeg1MoFdy5jipYIFN9gGhqydE4F9gIZEU
RV/nZ99INtChOBbOz2NxcgapfQATk2f4miCWdY6dVfTF8Dn/+7xWsrf/9E9VQ1/TJZVYSmVLg2L0
bAFWZ1G3LXhS1ysGPV7v7+ZNZ6ic8HlYKmYMaR6y8cGJUjyEf5fVHxBnoOH4UbsQN9M+DJUc9JMT
6NAaGHm2N9guYJiv/McLCQ/wipjHLszZII4OT1Lfs7i+LKm45sdC7+yhRZEmJTnY47XxLxyca5gs
7+EczKKkS3J9dEQxbmUAorAjm6Vogr7xNCaq/wkFGAV6daVrSw/Vv0NQiJVIBJgfNe+fpsax1ZTT
t1SiegnVHozASuHV7RggkqI5ipDa6y19ZQ16gK7RPP7CiSKIy8RK8s1WeKplJTyu/A+z0m3Om/uT
i5kUhVAyMSoDzVktRR/mUpbuA6yVtCCScdFTNnhR91ro+vUlZFlyzIrdMaHF70OunxtOL4VRX9EQ
Zs3QY0xeq8PtJ+7NjNrfeZB8jaPB1CnrU1PRDFEk+OOREbgm1qTBl0G/FSR7EQSWX+UAxM7IvEg8
vaE0benmFHWx6YXoFW25LYxNoPvcrpbTaEWVadf8TkJ8COqmH8h2fFFuJZAC2H1YX4QRcxUhAodT
ixkX/KLFnYbH0LWtCI3kLF0s0O/oczavvn+0Sa3yLZpmDk+zm+nU6AMX1HEIag8VzT+8d3J9g1/1
9xndiWm49Tb1giEL3RVyQkFHGlcTvnakWFKcjTwh+PvT3WSjkEERewDtFmSRLaONDRIxM/gl/dWm
e0jyzLxdt5Iqf5kAenHCiL4PaU1uaxIMR09lUEgdBxEgIGBPUuOB6fgfCQFN+FshXNPhZsXU0Qkv
SDiFpgMzwKZInz6Id+BFm9dOm+KoXDahbO+CnRzTX0L9REOsgkZICTCeJa7mjtGZSP/zWnPfVNx+
3hGveZ8Ht8RrfylHX8ZA/RMr6r+MTIrhzY5DSkdrPpESaCA8zLsUSQVkja1cFlyUZpBfAr2PFLhW
CYB++64PttQj0EKqYefzSkWmPorNJBb61ig5m970b9C+prPHL9Rq17hj6pZqmgz4Kg1ZS9NWBE4N
pIiYn6oKVl1NOrBZCURHTgcclXwmwl2EFyd8fVEygiJpPvSBOncEqlz041YDRWHJu9od2TxEWLa4
CRUMqpc/a9HfiS5/mpe5ugiegXaueXxbWkIjJ68EPnkOzzrrIJRXCfrYUS47kKgglTV245kcRdPL
UD8sq/IsrYL7Dzb/hLaZg7dlZrXergCAxnBudWEIEFyufHIad+PGecOcyyVmZ89wfxOq+UkshIMI
AKNd4Vs60dVfi/8Mmq5CEt/Jo/MmpWkNmvQZal1xJXXEUZ1K+cEjnxTGatmopNxAOQK50hPLWHFV
eN/MOiTEp7LGteS1bjhCwXI2NGW7Mu5tLCSp/RC0TrdhU5kLm8Yqsh47vEa5WpH4hwetZkdM/icp
MycjdHZrPePktEd6pcUZJ5f/H/Al2yLawKODE8s6kX9urzkK8wiXA9VGQESet5SKBn+FiDZLjvWl
G9APRWVVVfwTN0s9/31XtlH/q0kX2gRp/8GDtgG/ohBXWo25Q8apQk5tfmB6pcVpye+z72ZO0kR3
L5D5orPPR+FQjtBgpe/IThLuu4xYi1k9jDAnDN/W7qQIAod+g+jmp1B2PuI/BxSj8hnPBbDDoPt9
381nMZ0qK//ex2UWwtSP36sOm5HR1XLg7sX8c47z98x8KXJWDGZEXkVjpnI5D+UgQPeq4MVOqjUY
H6o7lxAMHGgNgTYI3yurnskhyOYsQ+DvtZOYYKdQWKtGYJmvzzaGG/pn5qfe5b1PP26bR2FBTW7+
CdBDYnFK5Ph5XZBrlYrHhkzbKqfYIVT3wMlZbT/CfIDPjlh657vRt0wIfIcHb7HvpBl9S5DnjgIu
vL6dN1l2QmLBYenhydcN362NeSahpDoCoHWMABejRsgJwIp30iQ52cnRvKptx5j7IGrQ+oBSdn9b
6Kud+AGnL/Y+CI+E+IINt1NQ9HeST/13r7OGVOnVjws672pXbvb8mIaNRSAruxyub5swrX2PCeTo
93vSyJfQ/XzVY7xzMRxFAc37DeC0LqrpQgnjSNM0pvImb9X+nzY89l+UDfylblxIvqxfnF2Rklsm
ms5f+RgHJ3+MRBPjATvNqkd0dwxg+bxKGmx38eX1a244Krwu9dDojJI4KUj/VsKOMsNCAmTUtXQm
PVhUjvlN3DeKvdXawIAEDtGAeUFLy3UGGVf/FKLh/9hmI/523WxAJz1l5pCh3nrvFhkdUgEHf0QB
Pqpgy9gczKaI5gHKXMGc69hVfvZd5b4flfYKzINqziYFGB0cf5Sl4r3xpOe6gwz4pAv4zv3z8kfP
M94AsFiIg18kJyExpNJveZ23NjLqfyehmA8l35CclJ1kplLVEk8BPg276m8Whak4gbA4T9eHeYw/
xzHCDIl5PniSU69mA6JsLUP6gN1BEYi7aLCXOSal3Djrxo2OiagJDZliaa3BsUGNQritNHGwSfqB
k+6yCtgeJKGGMITRlkqSK27yqHyVEtQ9jGMO8SGAyvvC/mTyojqbGBOPzLBi0FCFwMG6+OBQTUGP
XXq/Gp+8kdIwHONMBP4Bw3ehYupvL+0/9t9gc7MeP3sn/FLRpDxe+rLVkQ51DLdeJFmp4p9wGxgC
7WOrMnsFHF2gIM0HEdDgX0LCnz2uxQ1f4Q+OC6HwbpPzCdD/W0T8YWMdlNoeo5gqn5X3tnaZC7aL
EM47cWn7fuOfBSB1FvV9tO3FPC8RKBsFR3MplmOhg2sIuffQHRSuvne7muHH3f360OX8kvn3yfnd
6jB5eyH62pbuBCwe2l2zPp8kMlpS6xhpIdUZcZwZvbo7MsSLUhZpRpJvw6lTweR8jLxN4SSZufbu
0N7yBaVwchuMUl9IZm1RLwxTdHmqHy3LaQOSUorrAoHwUC+Wa218xnuyyjpDfI5zPPmKDZMJlpZP
tFvbcwyioAw0GFo/6Gqi5Pe20z/oh70eUJNbq+AtHKOww6UWgl4RrGJdPaaShMaArGZ4AoLuCO8U
aavF2zyjcnK2ki7y4pYZ47Ozc+b4vHNEbk4XqD92jgkTeUNvHOhHSG6YUX6CsjjfnLiXB/K2U50l
XUNmcFd3sqvcC6fi+U06qNPI3AN1JVCWnnSFT7VsJxq8c/d61pPqtA4dxCiKDbiyEl5lfvJ/B710
0TCsRea8ItxNM2FBAxtgPjSrFbfecuW0h4gg0zlwkIZfcTtHLpRVJe1w6e8M4rrC38b3SxBSUAwH
uQHCgKqlPOZrQRtKh3CkNH893ReuazPRhqJ7V7D4mcbUVqZbXAQG2csjHODv7oFle1o3DhwVBibm
3eXl8l5D1I0uYZa01C4fX0rbVyeLThCh2bDV2VEgNfcCXUqRSZ8X6psKHVscPlJi/mIx0BwJJCVT
U4Hqebi80bxvP5w3BjY2LvSIJWxRLRpcGqBDgkT7uX/ftiCCV4tzUKpvs2Nvu+zL1nmX5twTMgDL
Jyw+KR9nJRnIFR0lNC/FLzRtAAax3OY2dcgN8YfXrg66zLGrXDZwmxjr3fEtrDiA5ixzbBCcfc6f
RRL49N9L0BBbLZVPpsvz1nwfdp4w+Ad0nujQ5U0mrV/8ChU8RRvb1vqmUjE31ThUxZgDxJawIi99
oJbAagOoau8rNSudt/9osQyaqF5fslitiP3V5mWQ6UVjUhCS3yKNMOxZvw89sb2XU0j1HJNsdYJU
EmpTCtLvwikKY5esAxWLGqC/A/rjsBwdz8bgi+fQf9dp24AxbL9udHe+K7QVpXBRQ18LrhMZlOg0
3MeClKvLR5iLdBW8IvMzeTmnfgQsSMhxDUcRErsIXZbZq2+RQMqljfkk2DzoyppRs1mc+SdpcNkd
QZh0ruyRb539EW8KEdD6/QPg061JYw9VTI1Ll7KTIlWbzFf2BRCXRBrSkuf4vx6SfUVh1q9Ph7qu
giNn/PlnNHeJwBdBM4GMUWOMpA0x9WopNvM8WAPk/Z/zDDXux2nzy+mJzy81mKePsmAfo+07SMGE
xXxCrieL+R+ubZZwoOBpLGO5sETmrvm1RIvf44H1rlkStOKPpvxt4KKdqLxEpiPkWdAQXSA1OXTt
uXKrrNfEEebuty5CwgX4XYDqD1oWlzQcNhxpW8Nh1ckWJziaYsHGocaOhr/11gygEc1nTsNrP59r
R/RwgKdNu0IsHmCo1+xGsICXlPLbZ9u0UPzWZGscLA5wF9xqpaViarjVj/bXZtpdlqgHwFhoa4S3
TxkczsjThN7LKaxiacsotvRI23cSnEocGh4mqR1wjypA3K12mqnjHPXBZrrFmQ5hhyLWdWZ4o9Sy
vR6R7ZkBp9BGdmnKlJP30WOwF01TZIwUKWaPFuEp48sdoNVeblYeGQw7EHUoPADX2KuXxWciNf4S
d2xw5cwmRzvOQEs/BVaoENGqRMFVNumF6c85Lg7A8EP+lc2UGTIyGoQWIIekgpT0mvkdzOU9pG4S
m/wfjg1d4C+8sMQCBIpidAQ05sEil3JDRZ7qfepIKOgMFayW6zFmSUESBO3mIvVgkhnXsYURahgA
pyM/AfiTLv3lqyHeIAMkNoxZR8AzA/I797mBSlCJQflEp7/OBCdbPSoNfFWZOcWZpxwRyhUAlrsz
IkymEjiNVg5xNVmtrTAkFJJjm2IvsHwEZnhoBZOuRYcVnIGTNmbCzG0SRj2BR8MbgTwhngLHHVfH
74QOqllZfd5q6yNLU0Mo1ZrvArmFKrQAtHz3TJZ9u/KZck71jTwlbjhtqbqlBKdX5qGizNjZ88NW
pe0H4hw2hAmzKGXHOwFbDPb2svKYpcMK2I8kLeWF/3rKR0gB5NPCqZB/QVAqOVH2FlIRk3aDOPvP
JSPxvdIgy8oLvYfBNDf/d10C/KsPKGpNGHnxXUuuKSXoktPIS527PJeFuNrsNraq6StNEGIASb+E
3MmRDdmAn4+InHCz6B9BIEgqecXArvkIStcXy58kU1JMeC5zigEKckh/cMJ43QCNEr6M5YHzSYZS
+UjpJF+wN2r3krx1DBBwlbgVzruQRnj/WaQmOI2G1VFadOO5WibmAdrBNXx0zb0sZVbfNw1kt8rB
IjoxPF8LZC/NlDewuwsoSoBMosqfM38O+15KGfQDdSA5jWlNvZXTt1u4pvoxNeuJPdvIuY2eFnlV
6Yayln7QBsGo1NBzzLVOzDroQaLjJoNKN1eKvUAiXBHVDl9sPJU4bzn+eDpyGiGk2wXmbQsjw6LI
Q5fRxagyAQKRhClq5nciEAHrVVBumUbDEi13UpOWNeQ86XLltTdtNk8/n+R7J+Enal7J1ZYAHTra
3QVancCoEHoXqUbWQ1k0ukSmGD/J5j8r5GkL7hdROdLLbs2XSR7F6i7YJ813rIcVdQK7ydYgPI7f
M3XJEPfNjMFW9GJfCJXu1CIeJ6IlsXFlOF6NYWqmoRTp3hUYoFR+hUd0E0dIqxhr5+o+bHYvnIf5
izxwbPAhH8k556ANqXrJi67GaRg6sVQ4eBR20YfH5eAf2fiiW1wWHdnxkbfGoRWllIpp1xTfjwqm
1DkZ3Lzj9/o/lfI3VlYeFrjSiIvv1OadSPsUhuWB9m7CptC3wiKApk7Q35zypE1AhCxLh2UwGmZS
TvUnpvb4iqE7U+juRNb49JnxnV5qvAYUgX81gtyveAM5sI/DwycDLgn2rFiCklnTKnGg84NPqb7+
oDdVpi0oqyZJeCRhQW6ND6v5dBY4WnWVGs0JZX4a1bPMHGkOrNBhCupe8DmLI4YUPoHnKpe1pVRY
zBb2W70RnMolSXtBdd/uUNPJsY9vBDaM9nIkGcqABiDJ0PfdRy0IN9M7n2VS5gopv0d94kDuTyxR
eF3Q38HwnHBMEgbvYyiZf9eXWAPzMGsmSBVhhLqqsMQNaZ214qlTMWYYL+gTWkaGSKrcD8+pdbWw
y+i60ZwNbILM/5PFr2Ffm5rAcsScFXUyjZZkRyFX5xAgj+oda/78shS2JUagJDknfsGKChkTrwak
6jUsewlId4egP66VxinUn0/V/5EyO0VeXMC/UofTawW4IV2xFqlZbXrIxb2iWay4HHFfBwemf4mE
i+2mBvxnaCZ4Ee44khsAUdFq/5x8aX8+SgLg+zkPVDAp27GCFFvVtgcO7WKewvykjHj4dzH6oPob
eCGMhEjcGKfx49dQGwi1u4nfOKaN352hRcpDQTKdFvNKyUdDn7TIGMschNPjD69ebNmLn9tMgG0o
LPhI8/kGYSzYC6mjkYZXtziSJ73OWMzz4EOc//j9CXR8DtDovL63/itCBYMZKGJn+dE6agAOwypX
WFcr2C355Ba1UHhshyS98OD04Ts8jtFqg8YOqU2gGNzKW/JaAlpRGZzNltBo9qEK8XYBg+z609sj
7zE532fPNltrpTA4oqhDkU9BOLD4h73pzbzkd843yZpO5RE+i4cl+K1k3/SuuznYwz2h+gBgjw30
Yc5A4CCiGymW1mbTvQg1145aiY0HMUmUs83S4XiXcGq9VwXFk+IjiqbnEAROo6oAAXOHjVtItxld
YlE7DyYOexOQIAqfOGUDLGg7piIflSwpOcSnkGZ80CjvZ1D3aDCDGeIUS+xVKNQIMq/4n4vKO7AH
MBLbGoYFecwrUv7REqmtA5Zbl1/4vMNfqGWgiF0TVLhiA4Ai5GntkUAQ6A6PybWca3CMUTSXaPZh
RrmBN3GWSc0rcSgqgOpRIBaq9g8tm7ISTESU4R/bO+GTXQr0kpuJy3ec+c1CCkJoxB3NDzAd2tdT
cNxusZrbkKKqxpcuWzuP59Mt4rcLwlHAX3WHrtSxMKZizj2uGXYzIWRXj1vIumT9rpmQQbZshsoU
LkVi8L2YlYSa2yvqbczaFk4ln/xi5fSjrEfQyTYE/iyoYuTUvOBr3jJO6WR1f7bWQsXfptQE4QSz
cxZ9EmMm/cTHnlCXDwGj4KxNxNdWVQINhSQtW7YKd3GWPT+C0h3aSZG59aqvZKI2qU4bgJmlcHp3
OX7ep5ZykQFqrwbURdsuj05T7wncwlrJjD2kkO5FdpKzxPEKR1tOH1m8q+uJvXLeXJuTGNN6LOfL
58rp8KMCHuYgBS6xuv8Cmrgbw0DDMooldF+FT4GuGbooIxAahB6jZJeUeLQcioq+sbsVz59qtqDS
FJolv5Fz06R0GeXLiYTElLtP4yz7wfwZV3iiuh6QWxhfk6tHktqlV4yLsu5vtQT4LqNBA9WVnp1P
Q+xfem+gMBjVx454NByihKmWMNEiGcKlf/XNS8t3Pdbg0gT1oRBE50oImXVhqxdhRCUwFIPbKwpD
QyyWvWMBIY0N7dOa8HOUz2QawbGUMPF8k5VmXLiv3FG0a1U1DQtVt4XsdyQuHLjdRATXtpXusJDF
0Wu00E4MTdwGatP2v6mP7fOuqIBjHaTKe/FzDdOlNJnz3PNbRTxk9dhb0195iOwVIs00al3oT4/6
vKKvHzMJkcQXoiFE/GfNGW5l0A2QKFKbsHziIyZE4yJY9uY8/Wy9uHW+TZYf9nI7aXzo8IVv3ED1
zcsozYD/ffgQkD8RZSLQxXpbAzNS7wZ36vWVciGBcDXqfj71b4D70/KzgRPUoFgMiVD0cK9YEwi4
bnInS4rGtzEbIToc5x7s31UwjX0ypXR+sk1TBeMhVWvEnGQ403RpqAdgCba2r+p49pQb1KvDSe0I
smXSSmndJyg97d2N7jcRPe6XVpexBmamuarXnEeEPlLPX3yW/+h3SP/rRWwV8ucjJ7Mbtl8NnFJg
dlmwW3LtNcKQJ8jAEa3UuMiHUPYroOsZobXIQOnb6mcLQC2znqxLhM1imbxDLzE/MPP+iobKzB5y
ElyzBM7FxuxkxSw1scFHAQLHEPwJI5B0b3x2cdKiBDYLD9/A/WYLY3rR+4vjlIWVvF5MPCUxaMH6
KdgBuSQWiNEQwGzI9vaM5I+FnmUtji90I7EQMPkudA5XbJIknMcZlb6fg/Ky7O5121xTWeXSOjJ2
Y6mE2nDv/+HNRzFgPM1ZdezgI6U0bv6OhBOrB0RSvLgyRsYw3Grwj1jIxwa/Cw6QUFqa6hkQ8saI
D61my38sPBtOXrrV+JEezpUfUxX0+ZVCjGdWorMfU9bDBdeaHJC9WEA7ydZNm3/MX5SXOJ/sv9CU
qbUKfbnqD79/lSHvIQaACoW6cFeSloq9ul1qgGoXYbrf4yjqo5Y2lJg9XYrpyU/cTXG+qdvKSwJA
GUs4ssSVqtcnX8KLDamvJ5VhrmMmgsSTfxRhWO8epQu+OLgNtKKI4RPkTXC3qgEInz0WkAaxZ99R
k+dvAuHYxvWiuU5EvPpdOOyJIboL+7ZNtIIo8WfbNz0tqRaDkFb01GUdhvA1Dqu0vS0XoBWZbKvb
hrI5bgaRq6LR75XWZWy2MGoDrL7+N6FzymDkoN3vllfPAj4ls2SJs5hObsysZ4JEacX8qJxGoJu4
E7pNzWdXPMJnwhD+zjZ/BnqBKPzhX8kIQCdl50MUq/88dTJWuSHwW5F7TLrKuXhoYBdzrlHuF68V
kNNYOj+MtMU/zISyQUcuDPXu51UrzEvTDb9wWAIMn3aPPdHzfOpauxa1bJrYewKeU/G2h4z62W78
qpKQ+aitsgyHXRbVYt1cpiLPb/bNgu0+vnGmWJ1xZn5HxjkwAAviBgGthKMIhoj0QiwgLKRqVh3u
w4nxys3gDCM+8sKYn7GIxrWgF4dTXnokMBT4U/Mdw/uBEazR/jCVeBcGX97v5kyJVSJWeiEnq7v1
EMrTlDZT/ItUEA0krIwLC6O6DNDfF6uSkzQzRreWf4u75apzvtt4K796Cg6zQQu5v0PmpZWnHIIF
IERZA6258OOYF7ltIMT5EXMbTodX/qrQNhyK6IZYtSU70iF96sCFBZgWbcDcFZ+saPcfTFTsfbZv
1SxIk5wIj/lcvqzKqlbI2ErIaK14thbzuUPHnDRKUDmJczbsdcUSFLSIxAGUJhmod1LAVwE0zBdv
aRGxVtG+0giYOKgK0Uf29Jh7Ccr0UpytPTyIatbdTNEAhtxIWjspErYk8TZuhUL0Cy7HFnynx/qv
ol5rmqsAFngutxkpitCiDYJ1KbMX0s+5jM7PFEMR4xgZAC400hgBqDvaEFhpz1/nZ1ZXeVBF/iRu
nkGK9v8lPccxJo+/0J7GfYPg4vAlplMyiCxG6NT3qzhp4BQ5ATo2SQu4cpy9qP2pvfiqUJKicFPf
sxOlAmBR87IMX4ocRjVlW/na39jFUKAwXpM2I9tJ3SKjfr1zyZT7k63KnMdkoC2fOedx/zAGdFu+
gGYRMBNfD7NIgEW/ZVekhOPrqHqVUQX2YsZFLvkzbhlbnNmwO2TFsIms7q/9+SnK+/EL4e2HooFX
Z7jSuVdv1US/1HDkhUrBGxlDv/igVAumvpV6GIikpD7OmZxYH0T7OrTGeG5bpUq0PbdzzZ8ou4Ju
6nKe6KCVvwQzpkIF1N0IujfXPaz3kwjy+9mZyyhvr0B1xpROmh2DiX6K3/0xpW16dpGP+nxbSTvx
GrUU2OzlyiYcCPajo7wYhwmU9eXOTdoOO80hzn7W23qsLzl2noZm89F2AGkIbNSPgz5FQY7FC3ID
e6Q25k0SDjG0VvCOHwkjcN/VmLOIiY+JfqVTnWHvrxN/9PCt6ZzxEMScbrwErQCYLx2WH0oqsxMs
lKG+Wv0nckQqIPaZ/kbQ8oznDU21s0tfxE/0IkZF26wuMNpOXvRAjp/TG0FFcFIwfKPOjSYPGT+4
Tr832sjUaB0ug+/JttDVF7obZtxkvupU1XdK+zJOf8aKIGDdotU3v8O1serWVTHIYYTglhH6ZVwp
URC1xp2AScw0gmmOj+JCdcoJP7NzVnIzvl1VVu6s4DnZhr8V6Lu0np6iskqkz3T0jhscrUIeVzVc
ANb58JYPLPtjUukiSQ1IGIiz7F0tdN26z6WjODSGqBC+TJ4jIu0j66UVhe/BnmhmzaRnKORLYR9h
0IDeHDfaiNXQa2/8p5xqjgxv/tWO5mRB4KuUY/t9oyTOszzOAFC3E3PgIzGNrv//s/1jC2dItwaB
YXU/kMOrQlhcYEy4Fi33bzitZV0ao4WQt1+14W0RBHn4dnLJR0216TkP7/WDb6dd1E0dTaa7GFXS
EnMd72c1+wWBMExRrodPDZ0kcqdKF5nKgny0pvqU02fD4cGSL3vHxo4p4y1+/4kG6mSA+IPi3JOa
fTHOaVuoXZBqFrdNW50+mvPJYnrLM7J2iE5BsKrCrrM2f09j/8BRQLHBaYr3YFOgvxHFQ1AG235j
MFM9o8v0Y9SCa54mT2BqbtyQtXBrVoRMb1aWWM0vqoAXYeXebPNW9cOSQrapbfCBgRvx7W2k7Z4W
Nij8/flog9KkkEyxiLkgZTrPIsMGmJbE84/A996W+Oz+14Y435U9J4ZVkyuyZLbxaPQuQ5rBmSUo
HgCdVtXaIq7GQXgGfhUXfzFdUn/07S+FAbxmyneLrFmWiAl+l37S8fwRL7U4OQkT3vK/cVvw56oj
ovXw295wVUj+DNqCsI+RCUiqNW8JAJvEBkB99ikB48mWtc+DXiMOzJN9elhTHUHTgLPTu5QhEKt4
bI7qO07APZx3RPbbWYO9ViMBvg2gEnjcE0PY6CAq2GcnErLXA2VZfr8ChH9vGXc1u3+xb5fdiH2l
chfZJdGT22Fu+xYui5gTzlmS6wpbnT0LoN4OIr4qdK9hyzdz2orMNX6DFr6QifF5Zetia1JsKJqZ
QHKvEU0uAAZFudRf0jCqOkQpOuNLhTuxZ8RVtx+dogrreaUJsK+dg/CNEbgOjMpMNc26Q53TcOXk
0s12SFzXJhxtdnZZAHMLNl5l9Hzpt41gZEvlWxp+5pCaHGo2TrnHZERM1jPlx3jM+xp+qITksXFh
ONeiLwTVahKMhrNoraC4thzpOzhqVmjfl03CKG4iiauYp9/4mpjHPHHYCsR2/ejJe8qz3fL6WcG9
rSDRB6MQO+5hWWZh+ybnwibl4L4PD6YU8MCubcI6SlaEKFBySYUriPlZm18MxuiyFxJxRfFFJXC+
tIMdzCOe0wyqRVei67iw2K3OJim3Qez5hcV7MHETk2GFO7zOxvX3hKKtec8/sZi/XQbQZqOw+HGb
IKYDWmoMS3dptd7+GPm1TH1QFFydse/i643JyN18zaD6SnpTxpTAfG7OK3C3imJ2uc6r5IXnI4A4
Qj/lzqXAxU3slgOYoLIyQU56aS0ubQpi/0Oxhilv9gtagFPrFHUy55Uv+/W3LtaJH0C53NLocF6Y
GXVqJVI+7jAefiPg81w5hhOCspTGL/b4myXRxj1FYm1cszu+k8IjeAf1vhNPGB8//cIEhu8PZVlK
Koaig949qzLZhN6BnfLucu7qsXWcAixasObcdDAp83S+wHktiMW5GmtbvZ718ql2cg5JJ/JqE6IW
UtMy0HNuZWpoNI6nERVBr2Gf9kirbKEZQlKRsl59Wf4crAlN/PZ8G1R2GwCdP8mtzaT8tp6sorMB
cQwcoziUF+TtRW+DRJAhxbw4FqqQXyPoM+eilxkNLTqmrIongsEPorZ27hteqgnbiatASN60I2rO
ug5yThmkjXnTBKQEboUOOu5ng+k8oHUe8SFI37cY/yYbYCYD497KL8bXGV2k20GL9xDl5tLJgRYt
OwyqoziKom8UoGCdvgU6nmd7zCSLgGJKUR25CAzN8xcXsyU44I0aNK4ME83AiMDwOkKPeRgnbqA3
rNpnabmnZs99XN/kouz3lp1QWWo3znFHTvv1VNkOmuEolvxsCe+Pnfczu3NsBv8Ur7j4FF8aRSAZ
jKB7VrvOICA6SPZHv+PS1CbdqoIFOPzEvPyigFeuUI8ZHnGH+YaQa8pKDz5erv1dIlDwDayxhiNi
wLtSphe2bUd227lIzNZ75H4tFKPmhC2+DrdEyGCzSvtCxiUDBO7NVMdUul5qCccRZOrFwYi8xIqr
u6dJvBqQ0J+09vk5VQyEj/ROrk/XEc06HUPXY8JR2Y02TJCf8er1yl47kQG+WXSm6emqbDYwfzmc
Dj5WW6t2BRPd1COaDZYclGT1fi5ht/QNkbtzqNVbTEbl+S6tQd1YaPPYjk7UpOk61a6vaQZ1MxYx
LxaiwRJYIjcqV3Vy65wGa3G/uRBAd871LFcBzPfOv2GXsJSXfaSIQVDyoF/jUY9rURc4gKav0IhU
Qu5To02UL9YC9r/OxUfSM4VchWlmbgOCjGz51NPRgK4oIX9M7WNrQQENifNw664nhCidaXxY0Ikf
MRl6KKGABjTcQU0NNxEf1Z7NUjI0Wk+JJBiv5WmD5hQfxTiNnNou8Kxzn7vmWy9AyaAzYnNx54ky
xEAOnT//eyJ+2R6vS0v+YuEhV6iCksfX2hY7/i7TsTV5lu7Mn1eKdzf6Vmdo/x7+kHDVi7VLAtcA
t/8yJsH7/UoutrGy1zCmREcxvfbKRdQEHB4vxK01kbxw9wDpCUryFOkqzSMqVpEeExoJQdWaH1Tk
386fRjbJ89E6WROXp4MdPNU8PtKgE7hD4ujs7U6wl3bIBK1PG6AWx2hSlV1gG6gFs1/9BzhgITKC
Ifhc4Cy/YtlWlEXERo4MI4JB14oDjEguv+u9TcEuYGlyJliKT5iDWrGVmEq1nKQibB9FM/Hwbi5t
bQwz0e458LO/X4tv0pycdQ5arE99Ju05yinnLta1SZTPmjnXGX7nga8JeKinqgRm2gPjyd4fnXY0
7vIRDhjH9/LbZfS8hXRPGTJQGgNAMV+w2InlVETvS+QbIVMHXGFmurRInvyuBBRttbKGsCIKrdqG
t71zPecRrTHp7UYrlM3mfwaq7lkRGzVX34+f/629iBTOoVedBomkW+L8ejs9GLTpGsZ42eB2+cw3
JTtVmmptyclEOt3vVEAIULFMoOYN6TPPG2eeruzC4QDylnDWve9YPLKuVbeRPGZ7Kfop1ajn24B6
MelfZi99yltmkQmvSATm48tyvQ9NARcoYUcx50T30vcb27fncnRblOAG6yG8JdlloHI/F/rbWrRq
qLBmDcR9o6+PvMZkTX+5u13yO7WvlZiLujMc2bVZXswYLLytNHy7y3j3moWcDRmbLjSb8zfNfhzh
DaXI9TdHWco6yvO55WV6KvfDTfDwLQGPBx3JoYV769AkjEWkF5ach5AvTFi5rY/bxTpMzbijmaz+
CyS6BreqpBEJvhFdj8Wrxm1a/QQQPj/+B5ueXZBXB5mTXc217E5U1nSDNj3zxij3Tt4rDqwF9ax0
fQmqTzTj/tVU6UiGz5DKv/ZxTERaqs30DtThr3vClM1v9l432w159Slgt5WYSsywOe2ISVmXpL4w
/MHxKalVx4d4OS4271YE7JbSMyRI2rqHKOpU4C91vXV8yCB3EvP0kCsI9+KvG2OWlCfs5tnHcHYf
KS8RN/Jgg0Ma8EeAIUhSnpNw6R3s4xSuB2I6dbxF/hwnKSOvoJ0AhUqHUZ1RW87ln0Fce0PgIQfl
qcA76nos/j+XHUjZQdOud/0XCeb32IuC2U7bBNVB1KdStUV6dZioFeZUpkkpFCSQn0qoVTp/keQ+
3EzmzzyaP6ukFXJu/F4lftweuLxqSGHyvVBwr47cnLELc78OlYSHocdM5+AaCvNHodCEyu0hpxiE
BGUtePDEdnpxL4pV7EJ3vQqZkwtjwBXPl8MuhJd00cyKu6JbeXv8ZxolHfi51BIXZD9cnNoI3qXH
348yuFZTNNMInZb/X6nqYh0H19J/aAx2MGryLFrpBuPBk2tv/hFQLWNzLbLZDkQO4ka9+PGQ7XGQ
DeVxa8vsyAcex3/huHzjuXpzZzbzvxj4Wzr7ixvZFMsiNhnXbuPgVhdSxRYneusfzzcYBK4n8JhS
HBmlwUM4IcU1IyhdOHQxDEDVGAjpG/w8LHhEIDOv+U7NrJHZeaxAL03bhVxZCqarkMlytdjdBsQR
BTF99RvrykoDOl2uWP9ATc/l3WvGNVkpGDqoNpEfGw7nlNM2pV23MWpC+CcqkjHSDmdTDPqia5eq
wkTjiK1QvB42qRpKcYccsCWExHWJZchJGtHJz2ZzyEavZM7epmKWf4cCwPvpLm9/Y/4EpboK85Wu
BhhQzZ1B9EY5PrjOFVbZewIfYoagEZhsihQlh7jF8HJG5egZHqHKfHflXAwMdFmq7nfnHvkFcC59
JTSORBUywQyPCfHsZQRkd4uF+pIV+eK3Efz+WfwN+2MvzAUZIM7ds+rdLPuDCQNwbGq0RTpLh3iN
TjZ+GWYMdWhQgtTuW7b2Ej6IUomIC5LQKJE3JAATGjr47M+w0ymjqyM6EAFWQ1XK6sZFvIHjIiu+
gPVvgzPdlrxPMoL7b757rah+iUdiHbyTqjUNNrvD1o4naYYEtx1RSR9gch7Vnu+x9t3p+v4VVIZI
2OD8US4DqtdTxASR/DiLwnwbJRKMXCnRSB+PfGM5/utzSM309O6HP736Ga0KTaRWhKmKbzRQGxAp
WF1ap7zZoXDm2GlcMsWi23JWxYZ2ndz7ult7rZ0H0A8LY4G3K0BpLc01YSmk0V/6sxRiWE+PDQbb
I9/FsUffB3MHv8YD1z3gtHBG81gN7q2nN2u8QuZfJ3iC/i5fFQycN9mYyUhu3s2UGYItT5RNqTtm
6slu/ZiZB+d4ptYWR6Mml3ynFmVfCm9qYXZQuiwL1sqai3P4T6exIYuoPza/skYbPQPPghXXfD2m
ksrlCB5qjvpOTJHSeHVX5HLtsYXcL4UKVQ8KTC4gFTXMji4MGxU7t7COOJxxJSUXlLgbashb+9uN
YLcrkHxaP8XSXTAGxyEeh64Q7Zr5dkbBlsDH4o4h9MOVxdxZxPGxOY7fe9YYwzbavGdA13yCkRl+
ioE+cjJzznD82OxB0eTx0teTTGKRsvmDC+4Bal0TiIklLZC6gcu2AYvnVfKGuTR6vS1opi+spjFA
OA/5gnCmeU40PZZRCF8PD8mcKoKYTZUVHYd1isiQkXgItEbzJerdGzrPIqsx1o6N7QfN9ehnJS2x
Yh8Bgl9AsnUeasnzkeYUji/FceonDjVgmM4zdGo9/U9vjkB2ew2r1LC8GEUDX0ThdKsYsJ7nUZEo
L873nkZlw9O6q8Xn7AwIKBp3ijW6Wa/Im5HkCbOf+pOYLZhcJvWjAWR66SjN88PkYATC7I19fnu/
UfZzEvQpwNIfCz+u2SCZnD/pdkjRIteKCOKU0anjPjVhb1Ew0xlHIn1sQgI7cOa8hBtJctbE6xr+
WzA1SStZFQT4UG3O6ogEabkoPjgz3WpFRb36/yJCVQyr5B5KHRQmPLzwx8GvBOKxQysgCP+yh6Xz
pob5D208lZpsJOj9lHoGv8Dzpdj84uVX24uISmjlYeampo3VorzkeB3VWIaVfwcb8ILQsGLCMeF9
YGLdGAUgjWUoRasNWg6JkfhOT9FyEdhdWjQZMVTyUJRzWv02Mu+8HPhdpsTD5R/G3MvaEJZFadRM
bb+xjmY8pbtrLefVLvuksoy1PH8C9VixbC3Sg4Sp0P7Yqpf4zNTftYbdivI9pwQIa6Xs7cMa5uh6
NoVltJABuguBtjD2vPFBIRDVoPyIOdMGIeriND0GFqdFdGpLjIj6ZtV7oxlufZc1vS3Hap+1M04i
JUXI9O+SS56ii8UPkeWhuQxkQ1xCFuInAKEDyHiz+g4OAnUvPV5NQcVQjqSgOvsfWkONWVhcO7r9
XS48ni5yOFAnuyVO1DfEvLprdFFFgFKbx794RJy/ECDTqtkvOTJDiASMbr+xZ/Fzc8dkfIfMmR9c
8VZk/346y7YIhsdMYVaXXzVXs6GFObIN5tUR822hVxXigIRb9kfkzxtXRTBfZBFr01rlDREYgoS2
RsDTyduDIXFdkTRM6He9TKwIi1whj12wHVbDeViZW1G0hiQu4S88MvEcq+tUv9NKTfhRjcVtqmrL
Ds21g1kpCvEOkgY473n9A3/8s8wWFnfUpFzDtAnsjJLRcRbc2GznQL+06dM7tN2aK13wvI0++uIi
Wus2FcAgUvn+IQGJXS4ZM1zh9pluUij4ickiOqlfJEUm2lo1HLfhMBDLPYcclyZ0o+rI9V3AjSwh
CZihzkT542TtnFhD1+edZ3ER3Wk19MJZuGq0dnmk/5s8AU7hbSfh2CHF+/dca1PMB98tGpzIf259
aoUcQIQxjlCrT8YELotHpwOs8G6wZLm5POQd/uUPLPEE1Defw0F38h3qPXEPUdWJiCe9ZyQtpSVT
eHEtDuHsAOMFWSfYwRP1uW8PS01UB3+Vs2oNrLuDHHzSLgFelEHPPizv1Z1dhLjNwvfa6Q1gNDiA
L/cmBeq0s3AzMK0W2z+WoMJPeoVZmuM3XdSWcrvFfao1mH9Ag9aVjVGPLD16eydFXVNwebv7TLzX
/kT8JxnxCUGeFhrxK+AgZFep2cIsR3veDDJteT0BM+vX+D82HH91Of0y69LJUSWxx00qnp7kuE9s
dpfasc5ZjyUezQGBjPhSfRI9IbfusyZ49AIzJkbqNlh4ravmKhAGahWKA4WaJKxOkAhRqcxcJTVq
3cGkHxu3/CcMx8Cpl9OhCKvuyY4LD0ni29mCO97dr6FG7drdvjM2PITKNJm5mLSZzWP9jpT+drgL
bt2KWAj9/qFNuE8KEGtApwrpFyFhVwi+xggeLBjVlzxHZ+LXNtO8aLKtXcpXu4QToVztUvdJ9Xt1
OwCnzBTUYNynOJwJkSp+q+G/0V7qnU4sdDW+wg90n/xs+4E0ff/qNxgJb7eY+sdYBKmiGal+20Jz
yb4x9hWj4PmY4jwnOsqLSPR0TnC+atmZboz6Qx7bh+yQGsoQMU93w73Kw7GWWmi/ntvNVBX1BH61
06Goy0YJe7tQh4+ZukExhzI/hgKPVhUJVi/jdqLomLqa1chgLBK+wvsQPR6sZMBbLxrnExcYN+/j
h6VFyarxxEZQuEMp+R7F4X7Xqaj3s8BTGnkJzYYAFmCohxPF+DDb0lALhguRgSMVwRO6/wy5inIs
jdTVnXNCEYT0iIZkLOYgdjwDwgqlWKxvuNsnqBHp/1nCze+tC08MVpNKz8R5WuuPoi6Zm0oK4Vkb
IqoA1zkjgCbvvHVYHngYUPrYszYvgto42E7lkcXVINHYWNclxJ3/UzV3HzW+QBcYBdW/tZaWVX9x
DdpZ2MORaqrdNYjerOrd8nrhUE7+16gJNiN1/lOZQeQCvhQUsMU9v+pozczlVgZlsUh1tZnub1cD
/FAWL39VsWiGAiiQnWNWsCGnJwN6Jp1KgaJXg43sBA7XM9Tv6iZA7tnbV7ubSCWLZUEjKbzZAOQL
fJXa0fsRE3/j/EQy8uGtMOFHXG/xnac3eK9u5BuIJBlNGDna4aJdJGsOeJPs8FtdjmL3gi1fKdn4
cASjYnq0H2YLhZ2fFuu/hDyny4DmNaWAnDu8MjOYY6ScgtvUVjYoRcM7A4hTvi2a5Uvif5gGibsr
XLnejDZ8R1cvcip06xTirFEMKNgCWbRsC8O7z+JIYzfQLYREcDzPNn4naXZ0OhOaMbLIiU5di0fE
OUgo7rM+bV2dEJsIzSRI7SVLgRal+Zr5BpiG25wE7w4UU1+BI+oSl0MswhcK6v3cjdGiliV6F4W8
OeKoVhr3YdKyqc1AbjliBYyKRkeERrGsPYMkvYKUWlCBicTXMJxKzyHwfV9WVmhZid74dGsQ/beU
BcsG8dcK9r4sFBcGfv4Rcq6t963/kpf+xrK4xcgB+8glHGoa7eZ+X1lhpdKlGrNhLNjE6Q/omtAP
DcKNY12GI0wsa0l3x6AwqxVUla9a/V2yMHEw9834a1lV0vHIPUwS4wX0h5ukiPKC1c6pPJoOlpj2
ka4Xs7eDEeEA7RJLFLFFQgswGVLR664ZH80xTBf21L3CMAPL2i5i8fENn5pwLPmgXk0LL4rY3706
etsxWfBa+lPAXxOS5jFc5CZ5EQ0uXbGUeS6uco3urXiP+4K7euNSqTwz8ppb8dBXs6rdgBoO9WIp
dTKZoPvWII4jjRs0+F/c7+iO4AQplqih8mHxEbwDJKD5ZkPLuQvO6oqgNU7D1WAZdjaFT1fR3/CA
57Ep9IWiRHUNkHk9Q1n1dgLv1G5fYeOK7GX19oIoV/5ra/WZtrSvUBz/Cy8E+TkEDxtAqDyT/O34
4w7gz4xMQXnnKEm61fTiGCkNlxBMd//Vv3BCwdya647jNAn8iW/fNi7HNPq6IVU3t0p/h+aKfF/7
yMCPG/5E6eJ4LyEbOHvOzzi9tETLzKS2zvawu0VMQrJggd78H49z9rM/MFxYPp+AUApYbYufzGtT
cukIE6EXMW/OGP2F1tktOeas7kKCjq/tLcWvYps8u+QbVY6qbtpDiGDuZv+jfXhRW3yeWKmJtCgU
K7BbO3x4OVLP7xaLRl+pB2SZgPXoanUd5JRPZiGMrkwgqZ0yw2gUmUUClCf6DIde4+ZrTvqNSBZ9
PduZp9o1dmTc2UlROoxGZnJU8DHuQI7PPVfDmGTbRaX3yS/X5BI7I/LNxmdWZ+B9ns5YlDmd5uYo
HdwU/NJkeKaDPeb/cgUessWIdbj+DWOW3VPvoB/21KRKGW+gWpP8JvO2BvllIvsLbUPGHCaZFBkt
reYZRK8oI2JZo+YQsWi1ovDCaZ3jjmCa0TQ/PEHb4ez0k3GDODqEhVo0E8rii6cJImcjEEDNThIo
ejNYRA5FWTGSlEybqHOSGtxWq+OR6MuLbf3I7f2hnCQB7j/mbl8Rc23Y0Esvat7KeV8BxVpAZI7n
1kwwM9AN4nNKwLcrWg4TmcJDvcK47Ta+z4Cl2QJpVxmsofjSBajgjxJoKbAEDtK3oKSJeE8aklTL
sP20VifcU7LSQ+tPQwJGM51Jt7ZmphexQoFV/UwWJFNPW2VgQ+4WuwuwgC4Xx3MCF5lXBgrvJyHh
3QqD+fSCTscCmLh2b9Om2mSfDU8IW48hS/NHiJ6ctq23ir4BJhN0TkaSKs5IztwGuC0tUwMT6M0H
7KVaXIG1t2Eedu5xZCaVXOMt8dcnKDNPOCiSMCAWuyXVQC4v89PkP9fg4ojrBePLdI2EIqBvyl4r
Hndz6sFYidwGH7HafkPk3Ug56Xh+1wDu/wDZxGCQNDdUBSfJSiVlfcMEgOoL8c0vlQkBv+Efni+V
zuhHdDJjmYhjRTiUk8kc3IfwMh8/6igwXIh4L+SBYzWmd5NBj8ta75LoS6oO7LC4/NJ4cN3umxns
AsXbt1S82Dr1ay9z3IkOk32M4Bw1PtfK7vJ2JJ1SGmYqmH/4M7cN4gv71wmBr3y4yfmwagwUrF4G
KpPZ/zWtd5EMXlvJ6JspRgxA9Pd+gHm53Bszm1TCy3XH43niuBfllEmhmLiN/eSC/qUGcepXTG1K
mmBqP3Eebj/BDeJ6B/HJeDj4Ll4ltWRT9MQ/ok9NsnSg1Hccc7nuZ+zpCAfoPnVcUGDpfOUXmFCE
d9npCrfqpr8Wr8mc6oVauyCcjQNRZAGQeVJiB88pGfkIExktsAj43rl2zaQOQHO4D2a/eMBFNtVq
s3IIu29zu6J6+7ZJ8THBOWEn9ef4X/WiioQeAiIDHKvwu9JrFicdDBnmeIt015BkJBU95ma+vBs+
Ql7J3SWSG+Thk9MmWzikVIhzII6fDr4YePlRTFXHOfg5XDTvyGh54PRfUwp7erpYgGCTsI1QJarz
OF0XQcc3S9kY+s9ZySVFYYNFwEJcBVv+JeTfjX4UqQoNH3VfTs2HnNQEt7EtoGRfDT2S7A/GCQov
+Fb7DhIDFXcjm8ddP8vjQAJ9wC3qgHSvvI+GfDE+9qqPWyoshNzEiqXUttfVnhTRg9mXaDrkgPIy
0fAjaXXeFLM59noND/m1praAT4wiulIkqGjc2IGYh1DYEjJCi6AxUt0kBk5KFKPkiLYT5fmLAq8z
rW6RDVEuPiK1HdUQiqmr44aYEJqOV0RhTv5ygz1IcjbKZvMKE2YBpHvJmjx8x/TweBSP7hnmulfG
Y3n8xtHP+gyN6FpNOG1apFlxc9xUYnkBhdYnbjUt4mDXo4B6r26G+E20kPiTPsz+4Bh8OWUJnLjb
a1P3Jm8beeu4W06xqXur+HvUyEekQKHGpX5/xOaRPnG2LdFJEaaHq6Xhge7u2W1Sf0U1st/fe7r+
qCCwyZ3czLmBw5XLpWl4dkkGXmfyTLdvtXvLPHWu5V5O7t9MHpEvtuBW9q/dV8gTKMoimlZpjpZe
qI7cccZQJIKfsa2O2we4cAm9JrYLg3BjKehW5t5ByIfDBv5oXJbDl/UGdIeznUuNaL8Npr1W6OP7
dNFtO8nBzSFkGd79M4RLwezx2sXQk/6yIlAQJ90XBcXejQMQ6jGvnPJRsxMlMgQINFojafqBPt2z
qNVR0usEVnRc175wIT5pBqXTOawjoZi9qxfwiYSsPfmY56j1gmWUDJSplRCstVcG0ghojLTYPred
FAL4HNa5n/Mot5HamlQqT2OkKB0IJmJ8UYr1fHxX8yJGcQbkqlosWfscQceHzTDcnCJs1cUhZw0D
du9Rd36aYmGzO+rsbbZB7p5Q9sAIn/DcZmkZXK5/0A6E3OfdeMX+DDYeFSBwXlBkccB4KsI6MW4z
MAE7WqxyCR6FrtJNTzMlMyr8XmPEQMZy0nLxxiRC+23/VAl9pd/SGfkrviqjq626JyeDOEk+G6CH
ncdJ/aHIu/kbhSKUb0PMRazV1GxymtN9h38bBkenmMa6B1fgyeYjhDn5mKu3HVBsut7eKZv7PPs/
/SnjVlI/vlPAHRZo0GMpcoCdVrta5ieoD8/Y92XoGyzbWweTB6WN53qVdxjsg3jlZLZxZndcU06J
VpU7/Rbyzrf5FC/J+SdffBA4yJdwo+Pbo9KqPbIOpWe2PqafSXK0YV6v48bUUXI7o+XanEc05ohb
7kotga6SHqaRUDAevFvopq6Wrib+RGx8WwVnyskkbNLedhI/r0CBAPo2iCb490ZK4zqZT73m/aeT
mPEkAJvcZCNFMDbf3Z2NMAQ78EIoDJGNRL9VxYCMFnA5NOVgnwBFy4G93nmpYJUdmV2q19R6DLu+
CX5XHOdBEe7lyHCwJqrhicB244I8CTpNDAjiP8Di4EVOB/5Ny9q3aWUUqJt0xWG2UBAV/SaSonVG
S+OV9T+CaYkKZ2mdu7TQzmNTyMHwS42Vl8HVMZlRYsh+DTxgY5k3TzrqAZBeTzVae4yB3fEJGeLf
MezLBWKUfMhJx6K0bdyfJL3FbWgLHdshPnJDELnIyKis+JG2bkeZ2e/7V42202sAxwdCcvi086AF
842BZPQnJfT8NRPmFefCwFwLSRBdAKA817Whf3jqEDhQUcN4hY4umO+zGeWT6gXQ9UdyIo3Mejb0
mA0zWdSn/A520SOQI7kVFUV+8kjjdessJLx6z2nSvbNX43v9jmrNQ9k7OkAaDDjpieJKBgUuNGNe
ITN5iuSNRDO5uWiabsjh2cIC5pBdLeQ3SX6zlVE6zp+bTucOOulzTofE6Sx+WMAAeMnFm7DIWa+E
WrBAHFctF4quUHAnPMvVMk47/nf6O+E8LVQe11eojRQpPo5Lm+mw//siigWKqMpaTLI/cij6GHUx
fvWvspxKmj/kVq2uYNZZTb+EeHcKqbqlpyCkuV+96d3Ot5in5jHcezbXruS4xUYez+WaguzRKN6d
vOP457t/le3L6obrsM6EzpAEqzuqmJkMi5HobPZcEKxCY2Jjoasml2AsWiCTk/USsu3DnW4OFI6/
YjY5O4wynNbLcL1cj5A5keq8yK7wge5J3Gp1gJb5JTYYbh23GgnksXjBejm8OT2MtlR6qCKHfa6O
q91ebN8CBI0N0PxQYeZhkk3XWUAVLtJ9R1DNlq6TyMEEfOgjjDR2ZE74p6ejb/V2WlC8wYYOeDQx
UZEk+OvDDAATPMeZ5HwABtwfpR/QErkmV52XCNO6wiPSJvJU64oCS1MLMotWWQiaZVLtbYlPcGmF
NcJukpCcPfH0SlmCnfDz7WVTRjT+Fygiw+9v9TEuh2mkS493BIPNh5H2yg1NIaOZSgAhn9ItTLMq
dc+RvDCthemuSP5YDXNQHaMdLJN63tFEWhQQW6youZ6bIb46Zlil2hpHmTLeyk2RzCOR88bLVr8d
ivjFaKs5cqdLH+r+IoeN7bqik09jfsiAar5DzJSC3FbKrZQhCJyEnHE2XqdRX/PNCSliy6T927Di
4bCnUVhGqhmFOtsKI5PMh0IcVPtSNeLVFoCBFuLpQMX9ptVSi7si0ycfXTklSw16psX0zUpHHPkh
yg9Kkkth/X4nRefHZ/btJxYJw9d8v0UqkwtnsGEVRP7U14kGrtM+A82YUFsxYKY08K546uXZ24Al
r09OY09Bhd2MbBImV3m8aaNBizvYOL8XNfP53YxyTHijL73shXYxlgDKkPpWEGvhvDIWAMiiZnbr
tnqMvFSlWULLPgcZ3AG86apvp+BTxTAZoQcLjNhKrRkW1Lr7IQKXAxtSUPrSghrngm6mo7jDe6uW
gl+QBwvAV3F7gjWatfc0eoqK9yQ55W8msS5PybY+FQr+EHBMeUC/5DpTvcnhAo8+z8oL6q1yxuht
TiQJ2CRSMBO3bJJ17megJp96CraYD9PKrOGnYsl1RtVdsq8PqiJNiQJQgvW+6lySHpn+kuqXnYa8
1FNci9JUQWc3obEAjCgp8PyvrX/KAXGlm2FuP/z1BqdgApIZD4cCjvbbomhUpIgwY2EPxeoKl0NQ
qsRwWtSh5V5oe5K/sFb95RpFCYTcT2WYHRoOYharMk5+VrrCkiWJ0qAn6WDJOr4StSThh1I+LW9q
idjm60zA+cMnfi3GoKfPoIFyA8tso1vm1gJYEma0JsUy7eio/AY4TzY0To6hK3p2+CJtwWi0Zr8C
dSv8zZnnAkBS6CBc7fNnv0Vol51AqZVV8ScK45hFbdkav92PnCR0cj4Lr5MQFwhYLXPhFIsyEd+i
uujkuyY9stYe+a5G2zg2jNFwiIBCM/RrtK12bELVNfep+UPhiTmHSLB0nezKewraxHfUDGtWT02T
qUGErjJSrTKoH1fGo3JhragusHxdi14vKD4G1kTI6RsSpp0FLhN3rQeUy4eiHz1HdnAFXexQ3xWa
05Q8rtWWSGuOq+XeZkrSRh0R5HpNut2usFAdXTDoPZmuCPLt6vsbUmYE7Jp9l/WIbL1mkZUfRoq7
15YxmbYnPNxSndoFirHkqu0VNlG0wkvvtb0gnTkkmsNkIbuoULc9nQ1XMQ1cfFCgVvCdSZPgoIxi
8TiEB9rz0t6/nMwpFEGc8Hx7e1LAaoXYxJVhkl0Fng+KiYCtsDOImWUD8WFGEy16Rj0HN5s4KcWX
zQOWalryx2IZgFkvxDaNNCJON1QLxZRQZwcTohDyVMuY8yek5VLO2Tl1uo1Eiryw/x4JEYnyAGpa
z+HxFsmIN7ntjz7Etb7JuIpgAW4TjCbEqQxtwKhMdcDbw7hRzrwC6xbXazEQV7zkfbSCiRywASI2
1LxGDGht60vun1MpNy3ET/bsG/MRt3dql+j3PD10pyN1Mdoruml5cd+AlEIheoO7Ziku25+PWKbJ
l2XAFVsCDrf8xTGm2QWx+uWrjBJyYbfCzcs2tQ6TtXYeAILN9o86Fmw3d7jwEj91Y+3QwOeD5nSI
io4SgzrnMYcx1IA6l86Pw6WYQRsxd50wfQUFLbiFRsk76yB0dBBYeSnG7jcgFpOdO3PhSEAZlDMA
oaym4dofVphZuE2a1D7MpEQEtPCx3zA0MM80j1g9xhKYZXOu29ojKgHc/WdlKJcUAcXPX0+0nrAX
K9WBB6UoEAy5YADpHD+WAM/VWlMQutoPlZz+FlzOaIvLOtP9Ncdf5llr5QKLt5MXgCNkhUOyF7z/
ZYMIY4wVteBuVV/vlyKUt01TVztDGzZVnzFJyNOXI5hoTDkLdRS/atk+Nw5Bjkbqm3vy2AfzK040
PRfrRcb1+eLBooeSEsOwlylToiDrPje7aBKAG7tRWq1x7T78fGhdp8e2YCxl+taCOkKZruCWDfM6
mtqTMAIrA5esPp3Xh8Myr7FBCuYOlHgrBLrnL/rD2e0lClFLg3CGQp38kgGsnD51f+rxkK4v3iM1
to+zl05V7H9Ojt+Ufue9FaMDpZjhLJ3l1OL91n2q8PS/XfTCHJn4e/wDT6BVHH7GoE7FztB4FUUD
2hKLEglANOmtaVrxjd2QQDii+ZXwqtzWjWnXMETHCdBqw67QFS9VQ/R4HNxpVYpj7COTO8m1yCHj
cUvbaVYBb1OuKX5XGdcKPy0nrUJjDqCphwj02VxDdY0WfQhb0Nx3wdk30+wNUquVPKj4oqQj++9N
OWcFTLBji8Yppiq2GMYdfAbEq5xNK+TlFJNO+pKnU85d3tUqyih8PhJBz0aKLxSPTJ+8qle82zQ4
S58QIavHyBpTXcG3e+cIJfz4+hTYVNH40YYri44YsZzLi9OqRG0G5y4LxdHws1UBhZLBtqaiULy8
jdZzBfxKqMJI21j4XxVyivwefNhx03lLpe3RcFRXP129ygS0YXTRN8zGuvVZhN8AL4oJckeMp0bG
OEmGP8/irzwVjwHVlkcSP2oIECZR0CLShVaINxRpWSDWNrzb13oNzUk9iHCm8mtcNZtIbBTzyINb
bIs4sgN9IPNBwXaKGYTPOKQaEjwrm5Cw6yk2AWf1iRTKYwVgFuKR44mSiUEVrCrwuB9ekPfXi3XD
7Y6P8ma/2Lt9jJTq6l0PfcDFvxCG/EeyQU3vg6lux7F249Ji/sx002nSM3tauNxIZf7pBUaSyoeL
JT0XAlue9R3+YX9r40vwfgnl7r0YYt2VWtMLal+SnUEqhkTPeyHUDQGkIgOskQMzDZNifW4ucQ5g
/CTg0MWJIE7xwBycGTPlMKUd8r1Guz0aJprKzZZWH2HOQa42Znk3+WWmrageZh/WovGW5P6sFs+X
dmf6k0xfz94D0fW2Wyeo7wz+NrjcD+U9+8sPqOUoV2dJS9Dc4BrdXSygeyymcggvcUU3yedTy3Hy
YHcgqeyK+Tx54J++MuUEAMsAIkuKUbhugCZE5C0vF14buS63V9/K8dYfAxpPr9DQ8FTp8lMbfMMo
ig64gYgDKuOAcdfDZYhrUwsLVIGRUTve+J+b4+f+CfFANlLTPGwWfJSXjb06HHmDY+0GwAu5mM13
wEh+1SlFeUyDWO8eu53K52jgPmHRwj5v0Ut8oPBXimVzlt3NP0XZ+H3WMIIls/oh5TkoulDkKjGT
fi6JoDdwEIi9kXlq8HEOb5IYaV81I3vRDjsYNxE3/x0zmDznbOpL7P52gfvgakWPQBsB6Azlf8BQ
0IegYzYXz4UXxMUIkWLlE2FWvkN15wButJhN4Zo0spw0zjos05nSUNtifKONjFUbvWbomtsOVXtJ
nhZIw0GCe2bkKn0HwqfLVuOYtnuZr2KNI1jR390+Qs81xyWKflw0bX0wGXSWHcdnmHOThDkBK7fm
XEOxH6ApY2Ty4mAJPV3VjsL/1n6jTPkyfcRLQgVXNPCCIJp19kAsXWVTRNXhNs7MX3xagIXo95Hd
AmuK9AcYTdTGrh33zn1gS3RMXAaGmexTiMR+N0ExWryfdO/Cy0re8rpI6v7jaH4xKxXDV/w5NWq4
MDO4rUKpBoNjkN6VgAtzOoTD33n6foOB+cRlywcb8GLEwEzQOZYlC7SPa+/JnT45wHRvrE5e55vi
SAGd7WKHOG58VCMlFpXoM8eZYXqo1dRVW88LVcuspdUHok3sDl8PkiewUFuvIqwc4FkPEqSeRUck
xRMW2mG98zUQNT43W3ifA2Vxv1/AAwLjMUVnhQBUuumcqFXTS4wRWNzcxVQVSOj+yQdkOIeK84/W
rx5/23yHoiRqAQSbqKlrIOMv2fV/K0OSikIISuSJIxjVVDNrDVQPBzzTRTa/U6q9ysSlauwuG0rz
0dQ42yOyNqRV7k+VJ+dyhJIxKIwK3nmEn6mlztk2ImNyq7keh2wTELgAf9IK1u597Ij4YCw29FPG
73U6R4MVNmZ+u06rg9xD5PmCBLa7sZFDL6O+sfcZm4kgvmuIkxrYIuHg5JURX2oc9WV7/ym+ntBZ
iYk1rqXrDBV0UP5hGI+uk7E+KsCFOkSKFFzfECCJpSKK1ae7Ac6pgBtBqYyfiPi/6P9YMiq8bD71
BhwUcnmeHaEgIZFGd+Y2q4kLQ9TshPxnVZbT5luFQSO9CoFVvsCFaJ46rBExuQyTvebs8CEoXgkx
uSiDOLTJHXgBKjIgaUmfSy9FvShAHhk22XUI2BTvmOZhe0y0uiINdrSx+TFeZ3lAaPNC4yyuo98y
MQpblxWC8+TKD8yb2COz0XGp9s39A8az4Gli/QgoldpW/BSp2enrk10NnlBqgEc/5P3m3oEkPHrA
TAIfJqJZYlLPPWQTbAi1lHZIadOlO5TucSyVqddyQLiNbQcNmeZtAq91hE0RhuSn369va3KEXIup
OilY61QFCECOV31NGgOqzdl8MOJINhlM7dfzblG/Zqfgy4khOkkQV8iOghVomPHWGfe8YIMcmdTS
dN3/0j8voCXpIyFZCi07y4HbVb+/357BNFA3kX85Ms7KZs/zGb7B/SkQ/A8Flp5y7ujXDmCA1HTD
4XKSHFvepJRAoo9vE2/7o6a/0txZfYDiptw4/44Dog2NJGTfSzCnWcqADVs/wjtFvxJwvFzYXzlS
WN9DSd5YxZDiFiO9oyrHoSxRiunlXY/dOd8Oh9DRYLGjNfvSZu9y0XvWP01AVQrVhWkQGk+hRkIF
nQ8/Pvz2br/8zK4mrknSfPaJ5PkajuAoqzxvzHhqxlcxPVgX9qS3i1InM1NFEJkq8s3ZGwpYd/64
Fytqh4E8tpc6iBz2bRj1JDYSd28Gna8xk20oZw6QuETXtYQIolIbMbzyFo0jqlWtdPIdW+S2+bvf
s7V9PRnQ8qL4q0SHwWZRF7RVhYyaJ06l2laawL1dnqSAG9eUyy1gobhwMKW3PzPyXpovHUe46zb2
u4Aj0gD20CRbd5fkpfTv3W+J3GRcJmgErOHuE03QN1btNpRIdz+5/7/rSCOVTxELfIyxA4LCYArB
yPmhZNJBDCoOi0GTVk3bWIqCaCH0UeGQS9Pj+wEG8f5LX4pBopPVWMUR4RZNOSMhcaxqfod++icC
0dR8rhYpehFtWh+U1Lh/XlXskrACdJ6SRMwnMIIQC0HmQyi/knNJeN75js+TnP7Ti7deMIxEPO8c
jlOmZKxHN0dQu/iWPsGwoEyxoXveq9z7EYZ2QS9JPDS1As87+my67evdg4k3uXXgutNsCW13ll7x
mS97sr+c3EDTzh8ZMeYhSCt3co+ight72mD4N06SuGYIIxC8WXQ5o6k09h2/JJWB8VIX3atORa9Y
jmcNY1Tz2jIHJdLrp+sA4tYPue8wMvypn5i2XFM7al+yhqMpEyUNkRNT1eFX+1XTzKGnjtKcDjh8
NmrwGhlIHWZQhDeFXu+PQLtinLIxkg+AR9p9ckeEY0iSyjsCyMl5ok4+4eyejo8uJxz92A+S67JU
IExj4OqxAHM3dPVfNPHOA3Eo26tOgNKIDeiUHRkmo2AaZv9463avTtxRFKo0X9bHCSSFnxYKsFtV
FRr4lTg4SuLrMPgfKOWLwCSrSVuGpL1UMw1VCf27olfwxovqNglZhD7qf9MlKnXyEwNpC5Hkw7ld
vGsLVgdnuonjTaQXqIm3Vss0ut/SSzuQ9j1ePXHJ6qoI7UQ5M8Q0za1uuf1aBrgeQIr4mOKsgx5V
VooL3b5FU4mQ/x2hfDHh/zEHr3Ia7rCmlnUuFCkj6sTPwIps/zuqTXf0/xaksNuvF1ffAwvAPXRB
RY+2/1qsFqH3TQ/ymO7M4+od6cmA4O75XHvBXiYUaRnDLJDla1k0mz6LqsG8/NgBvh/kHj6CWNHL
zF/xEjQMVI69nY9ggpslwrKswgR+ytz4B3denN3lFxKxQs8jwWQccYVlvNRc0hl+6PEwJUP1C4Q7
wUWvQagH3Sjy7gaFZR8pu8Dhq/5tR2lddytGCqf6M8StI7BQVPMVNTqOf5Sw+AAfZoXJwC8MOYF1
E5dc4CEgeXXEhiCB0yOb7VjZRsC51c3YC6gUwj9lbwDsQdCVl9hxEoXHZ7iPNFf2qEZqAJlZRzHY
Alkja9YwREvUCVo87RFg0nfn+fBoHZMxkRTHBI8MoQ0+v3K36f6iPsb2zfg1rWtaid7/Bi3c04dS
wP3oEWiroRbeT9LNonGbGhRd6XTetjLoRxjDztmI2PmQzsNaEFHCOOjqWvuer19+NVFsFAvLmdjs
EnfKYnQ2dzRUA/7ek4DsLtNQRpSts3r8eUZjXE5I5SUc6AcTYG+w8maHV9F0IFHU0cJufcVcTm3b
nGvbqjtTqs1PNWDo9qcQfRqXWhfAOjeHrOdvqD7IGKvzDTK3VqF0Rul4MPty/SteROLzsvOQr+D4
snjp2GoIB6aja94Yz8astmGfb0cNh9d3sN9gWkrpib/Gy9aFz5cC96pSBYwujIbPKOqU425V7ZQ9
Hl8jUqQfaAp/Y0m4eIGD1J1BXVRCqSnNu5TwPQKo4zaHpyNSzl0//aRKEoeojdQ7nLOmbRwSJ/g6
eXNodgZWb805kRVs74JvfSWgtRHqYiOD2KxbaOfSSsZ+bCHxubq+hP9C30DdAjxUV7QAfp/5OLO0
I7DT5w0ELaMNv+3KxgZ7ZLPA6VxIujEmhn2GPOAAH+JfuzDy1LJ8H9hbaK6lx+TU6dxUz4ZpXdiD
XWUIMv7TpUZfwyh96GVBwWsTomnSxNAI8ZOyex+gdIXvm+6yDy2pOULPYDeVB+pYdA2w9vya2ffZ
TxmntBRRJ/MWkvvPkMF+DPKS65fv/pDtZ9XypXK0reEQBkxwJO+q+a/ADJ0GgaKWrOyQfowHZuJV
2Ilk2Q3L8w5FRaUJLaMF/C3AhXoMK1kg8tGIOCZw5qIOx1QulLknPiudskfGH1ZG2roiuv+SNfK1
xa6cMnaiI08KqQBaZqde9551or6hzwlIFRf/9jQe0tzLpoW+j6EoFWTX8cDqid6U98+lGd+qnI5v
MggtFg6qsm8eVIsh0N866TaOEByrEPEJ31HZ78HeJCQOnlNSzXEIlpILMlScHCmjmMk4seBDHoIf
NoXtLBeK0EAVyG7b/QCEyiIg7Sl956/d61gRxa440Cp004AZGc1PUstocq1paJlhA2kLOf5RUBoq
sdE9O71yhfQUr8ldpEg6GTKytWE2/rf1H+WN+tJe1vClej5VhOqmnglIpRLu/UvJGu3XV/zX46r9
B1SSNQk4cI/pOTpOZrbP+mGeHi4pNUHeDQ7EDXs4UIqWRV5MAt8+h59/ZUACReBpYDKaXBHKHve3
/XNQnyU7rufDNl7G+Rd4J6Eu0EzlJ9weqQQUz/ZPhoG7lI6foqmehCdrQ5islMn8i1+1Yz9zvJGn
rYCancLXYNsIVyzDHaM/zvj9xaistRxY0Ss1ae4NPTVKhOomxoQNnxZ+nwU/JTesympqDWUqJQs8
BTH2GMFR5RuqleTLhx3wp5GY8AC9AtBgteRUoTSslhL9EvV+S+5/I28/6EMIgyXOLXkrTqx7ZaDA
KndAg1e9PrxwpBiiYee02/fP1OrV3nzrjDQ1yg/qUoeeoBOAQ9lyK3Ymv0Amz4z8V/P5MKKHe4CO
AJxsVCNJBiJJ3qh/DetQaTh/RC7+gzSoO0U3Yf3YSWFzfI/YR2pRVa5RzkXNzAEtk2wREqr7GNB/
WTcCgtiDgCsEG4QuGuwfxEqldC+dk27VjItyFiZydkw56eM8/XLJeSwcNo+o3RozdVUHaSnq231Y
nzBbr/pI3qNv5tg4+JwVFEuKXhdShIfUVX55P3lTkQCtVl5rH50/9ND17gtiGffe4Xs209BmYQFb
YvT22F0mnxevLC4ztmjYUwgXEp1xDsAlCgTVHmRz9EOLilPNlUEoiJ0XChhbeAr1ZdIth+agLHbq
vcnpxC0sx4fDMVUBl+ezFjWKQSpsxi5zxQeP2DwWT/GASn3JwjEH0ay4BZQARlcc2exj7S+Z8g/T
O7/f23FP/iFS1JU2998PpQXPAh1bZZgZGIPri4xDBjpGB1OLCq8E62GAvZom+xBN3cpZpoUYXfxo
69dvSQAQDmai0vK343/gJJegkEYBibh/95h/O8PIYBL0Y+h526KYLuqfVyu8PwFE8eV/klj0rpe9
z6ICQSl8kUSLQ6G5ftzFoWm3GubfH6CZLJu3DhKZf/+7DTufvtEZoG8a6Kzi7jd+AOyUyZpG+YhD
vlDP+QOv9kRHZEcaL70ht4G+TXeCkqHqKC6KNOt4pQVnrSFvDxk/+s5wOpQKULabvvEMcNWqFQPU
0oUqStYJl8nbTpxtE95sm1OiWX7te8YdWhqLujvGOhbtSJhFXdgV5bQrscNujDTF3LyEVfEIDPiu
pL0+hcZah1CAZtzWqsNSx6uG4DR0GVbPGn/FAJAN8yZbkNobAmlpf6gv1Vue672trIs9AH0gGI1W
EKAie6pDWf5Mf4o7d8yFJuRuqW5BA6j4ZUjT7TODXNi6GFy643KLwSloWxHguJ8/qdqDwwAJfU/2
NvEsB1lyZ0t9rfQtS8Al1Z4vhjOz2KZJOYwEe9oPgoG7+Cp24LobXGTyYaWloS0eHGjGdnlI1t/N
KdPa3G2I4RonS//PFzE1XDiV6XFw3dzLuY87pkyozwH1ihK57x0NWQ8iT6ZVGUv70/cyy761vn5C
0bjDdHnrh5g1IZWQnrH+6LcvtaVc0F7WlcsH/GAVF26JtUgydHeXWbxt7Sdj5W8V20bpcltf0O4v
V29yiJAgbDS2MVZf1J6HuC5SvfBazSckV8A4dvjFiz18nz1lV60ZDDmXk5ZacLWwEfrj2Igyl52b
3WoqNoTvwMH/kYAH49ctjqgS/bjrPiWlBV2LbDbvYFC49V5V5KczRzsRNMC9H7rmheErcNGboem4
7lK/rulNa7TxlSUKFMEenufLxQ9ackH/wAoy6wlMUHg3hhr+SrjOQSj2mCuNsWWLEKS2RK1UZbol
iOsydALmrTEdjkKqMNTaxmhraeKTrNcENWmNS5L8CG2rmCHDt2HiDdX8J9skQQ0evf+nUZFnD52Q
RZ1Ts16ybM5EyhTeA5l5gxXaWIXAIn16dR/0QrAZpnY1ghPRTB2f5vfuUY8WCscmZn3hvmFXvfCu
K2cJT0zdGCdQTnU6yYY96UnoYVIfbuNi38Rd7YoZusE6uYpZpCgy5aNm461ZUxoz6u1RY02K1/Dm
LqS00wmST2QJ/L22rlF8DQDX78ZXQxwEyUjrC3FicgO92ZBg2zxU4taDHclTDXG3glaX2SsfK5Z8
3ASq73726Va46OiX6DqgM+x8yEUsLpCKFOOO0c2/EkrIrS7UN/UAbip2T2gZch2BGCsaMvsI9wCA
gF+Io3UHBqQEWLMg2nmCI/5ByFKXQl7jFTnEBnMgYWHsyrCyT3nIneFbtj+Rw8UWTTIm85WBeOtX
sfxtcXLqQy6oIKqInqW7y2+AO5YXBELFjYcwNhSDR17g3i0gqV9tUR+aB/x92uhvcvvFLb9UDNT5
jnrg0cGYPN4wOTAVubWYnkDw9NR94qHsS/48Fl/E29cRJr/H/RgQwAydRW6SQAiONPIoCBMDfbDs
H1W3y2w1dFEnpAFAjlD3tKhuqYtUPYeGmQ1Ntp/LYtBHeS5ko4ZGTnPwp7vLjp2szKZhs18PpsZk
S8rNE1ByqBbkEVhYWv4jVzTTiqXA8NsRLSBaBSr2SOw+uDwUz2upT6Cm5Toqtz7SWt4/ib7xzWxT
94/S+btklalRrQfQfTkxlFL1zycVgAWgS4qJc+8Y5btlgxLqo/HoO4ZL+eVcPi5kA4V0kKO8/DAb
lqh6gK3WEGJVTMnNBE7VZsCQurvaWVxGEKG5x3PyY/49AunmjVWkhyW8+JFiRamoqFWXGLjNxNB4
ocUBkSHaj7NnvSR/pOAI6R2C0G6x2iDZ1gU2FcQzzKrupGwoin253tooF/6vzhWWJE+hnRvN7rTx
MksMa4bj0UXWg0qcipwO9fMkDsrRyDJZ/0hlhXj2tGRSNJRbEUrax4Tf5cMXY8WL/Bj1Gf5d3cHs
M+8krAww+SB6qbBBy/dRvGa6Rcv0e/ux/x6kFhHTceQVZuaYl6V65SjeTtz+QECc3LTipoGa1RMG
f5EotMf1ycXZSsq1ollkwihW0qf4seXXolBgNcx3DbpYYAmJF/Y2S+OOiogFyMEJfF45JBv76u00
XrjlTSY7iwmZCAUqNWlU1pk3SaPyTwJMLN0mrG7V0Sqi3U+Rh748Q1p4rFXYGqHfmyjMX8vuZnWU
62auq1IJpemjiKBMcJIfUQ3vv6T/8FgvfNoW3Thh8hRsqc/4HKTR9Y/jOsez3KuOBYPOP071btkc
gdFvVJwsSmZKydE9+f67x9aN/18hmHujBIKae62wrXeAmNWU7fSPe9KW0S9kUWDsgkWQFdDam8Ze
tXsN8ybKNFBirT52sCnSbiaLq5lCZpJM7noLpYbdQTj5/sbx878v85fvBWeaGKY3bHjPZM7I/0SR
YUv0A+omz1wCipY3yiEv9qfv91gRpqHNlRNVjI1EoZUGEnxPQzj8/w471OgQUEvc9NqQQ3U3/oU3
von2Dl3VZELWxoytZyiUkyIyqkqXZ2TJLAm9hIh8VvBajtSWmiGBpm0NUQt+1njXwQSMyDONQyRv
1cE3plHMmK8nxXEDXM2k9cE4VdFaECIH0WRBchWxQbCHSMqrmugZBcvVEfKLRdAJ64c6P84dS/VC
qQYWRnsvarAkPJsP5bxIF/HNCqD0VT9dubIxKuo/pGF4p/KFFfGZeNS3M/14C8MrPfhx9BUq4EzF
2bAhfVHZL568fnwSXOMD3mwpSIREg4vROqR0dyr92iqzvenc9p4n/LaKpfNeAULAyG4QqKbSVXhC
Y3dh78gwGYCermsjmn1W2cK9nglFT1RrG1QCIl61ZGqhuq+GBdLoxwwovUZaL+4lzMnUV/liwbzN
BVsc6CvLhbHghta+HHyFJ7Lo6qX0QHYGPeWRpA4djBlUPr+nQM62LNs0R83VZvu9mXwuDxfND1Iz
LUlib7lBNfzZWJHKE3SNfov2mN+SCf6m654y60RKhWdA6cYPtpkISUv5i0uVq6kFrxWWab4hj0n0
VgCA8d3rK8JUXTRz0I/8q1VptoY8mQ4E0MfBNuXN86uQ/DMayU5J9MK6lWMRdkN7hJ8ss2tqHHq3
r7c3LV53dRu+HuHxMl3cSqJJhcCyYN006z6IWkEp257tmFmeAn7otQbzgT/8mGeNPSL78X77RkV4
MX7B9UG5Y9U6nOUczob7+/pXV5wC7qoOl2JsxJ3YvkbIyKOcxWegP+FskoWJSdFdj2He3lDDIw12
pO7vPyLOvrCJxBUp8625ONR5T0sP/BY2sxSITNfomhp3uNnWkmqMw0JH9STQkMc2pNy8b4kzDvQ0
nFkzyL/TDr/Jj0bAwGnKFbGwTAlMd4DG7/owtRKo1TyoOFeurJsnr4GNjoLGTBhl5GY5z7bc1uSi
aehsIysIJgumZHKpyZ1gBwitYOpjSe0WtMkRFlGzt8C8uAMctX3CMjXv9+h6BzsvpYSD+di80Jgs
z3UGr6CMgl6fsOq0eDwrgCq/QpLhoA+bVI5IFzRkT5FCDl1WHa3Qekqfgt1jWsyqHuIjr45WymSz
65hmvhuOeIJZ43puPZRDdhOwviTPnr98kmY73A9eQLPcZwn0l/raojO7quI2KdxnhsdTbEIsu45O
F9EEhsNUszXx1I7CgzoLp2hf/YCIdZ1YZeQWDzFgd6BrDAM1aEKobjl2PresKzVyG07fvBscTcEn
/827pQ2UdiwP+3k1nSWKsRVfi8euCeUG23IvbYBVDz4gOQ8RZ3dOTJwe4lLJxCGuXqy6/0cXHB1o
kLkWWWFDaMtM0qbngzSL53qBvpF663h/j85XOxHBjC4l5DtttGgRZ3aTFSKJ1tHwY1+95w3RsqDf
/B81IhsfqI+7B6jdIHR628wUgKebFYs5E4kqg3ZDsogJ3RDvxNULp4vCfekkTe11a0ux6/d8IKOq
uSYT7hjMS2IX2ZFxT4+KB0Hd7kyU4gudFAOt6w+fy4aYTU/rnZwVxW3IXcqhAlOim3k0LE2ZGssY
yXGpfB2VsQWFvKlqZ3Brm0puB/k0C9V+5TS5OuxZY/Q7aNRZJ7Q99TIfhfYryQC8sAEGe+/3vjXP
7eBN8BozKBKCEhYPYtT9o0r2StQqY2TeOcCJXeUccuXQtNECcypo5nIH4rtj3/qYe4mzGWlxkgXR
D7SnF0eOct1a+h1esgNa5YEaeWw682/V6gbV6CNwRKidOq76IY8pSoH4GAXVg0UM5Y2QxG/9zTkF
YuGtIODla0UF2kkVUEIIBDuyrn+9Uimkh0MUPj2bowtPgBEmUbZtgRgEsR+zfQL1K+Q80PEQM+ej
98IyQYSGJ/oBn9Hetn+x8vQZnbU9xPddsxEVWEtQ9SIOlQZMvpq+zmieNon6NM7nPYYKyn9QScT3
8Gpseg5dL9OJJdiWMqaKqayH/1xCkYI94eLJIEIAH0gsrH9MSA3KAYOXcu/WeDn7hRc8/H3ayuyF
f4aaFhfUoDnY5xgeBqBp9wD2MV4p8OQt5OWSrtJDZTdIqEV1Lt7W709tU+LolRg4zvBw0yLU9Osq
Rqx18V2aTKxWR0hNjr6NqfI1ELxGavMSZL5pw2VvSPuXDBKgDHg5xF+8IbRWFThwfrDiEepOjDrA
pAe7TSWscu7dZehaA0MvQPHHYZ8sN6dO0poBo597H4lDTAc/XtOzmhPcsHVd1x8rOTZV/XZvZc9i
rilHZ11egRbVquU9cbzF4i/wi52X7bLGTJ21fWllfHCKRB0flfusTuaI3mMa6muCq1roG4ZUUcLW
JvML2YVs4xvHDdREJjIXnqKXxkzYxLQHlvle3ah4givWJuVt4BzKRXoJMyYITlM1f1o3VS1+IiiU
hISRcBu2IBTYPEg5hFK5No2ePu5YxdJTURF4G0hM067jy4qwJBIFYV1qoS4l9KHoztpA4fYskDvY
z9UFDC7vrVYIcuXXwtS6AZJQqPDp8k3qGCrckDTAiJfd+af3QmSj129SWwHnuQZJLequRckskosU
dYRyOC4xT58hyev6yOezmhaBtzjlaAnpw1PiaHUp8h7628pOErhpk9R/+CXRNWv0usW5p1WaJFKL
NM6Q0nxOmQGXCu76CODNg/tY3aOkVLoR2fnf/Cof1JWpjqUUo8RcSQp52PtWrbcO8x69ZC3QbqyE
J8WD9SJsblv/ctMtuyWDcSEvqgpjnfvumtfMwPWSYAlQEaCFz9ZTGJCb1xP7C05IxGEfDOxxv5do
eOxNJHvWgH0XfzCTAqLK2n0LO9fQe2mR5rOMAW51LGzqJSNTzBrSc1jz3LouLyRHKxzin8cl4dva
si4YPl2OXz97nE48mcijT+/iAzzBkC5u0Q+zwtw5mZTHYVgw1aKDvoltFMVHGgs+vFAsobFAGzwR
5nbL6Zo2rBhl0hb+LeB/+RX0ntyCfrf+fGsDVE7jFBsa6339Jd+FgxIqXu5JS+ciKb1Tk8wun6lI
iiLj4q7H2rGIM7WTDVeAkrESzSapKaYnTo+ug6Kx2s0N4qneAJefAqsGE4J9DFukTN01Ag9DeZBw
0EexvEGdhEhflLwMKmQFoEqmfGV/0Oy34RiZNnRZGTFZ3BZLF0SOQFgWbnBGR5spnlRuVQ8uttI+
uMuxK0GNtqlxVsAhGPRnnxYqjj+9XB4reyGMjESGdqbQ+Dmzk3V4WcwSo0Udtt1OuYzFDrmfBjE2
T/QYQkUQPFa0g5BXWgEk7aCfzyy5HFp40YrYl+QX8KU11rIqpUd46qaDjP7PukK2WWQg+gztV7P7
ljFD4FaCBCNRiGIzGvgFpmj3N/LPXpKD0jnLzHatvifKaED60Z1QQ1bk3moYPWXefdl8/e2HrEt5
Ao3M9JvPkG+ALdmj1au75uMIpm4KN2KKQIGu9Zjj3Zn2sBz8qawQYfU/BeOiffgGv8k9zUU5wx79
et8yU8ZlDPDI1wGRRO+qrX1AIgauQok8Nb+uI4pITQzqzzIdrkLVwVT4qRLR1poTDGWnqp+aaCl3
9r0NEljzU7GiZiB/9JSNBS8YJ2KhksovpWNks4GaYLexMQSHAEjcJjIL3++MNvrvkmWNpPQ0oB0U
0cP8BmH5xCfkSxiE54rcrubEyEObkcQnrSQa49oRnyRVRPwMNo3WPLQd8t6D903s6t7fXcoMtlsj
KcfiQRSTTiYJqpJwklnUC1df17jYqp2pUs1XX7UgZnI0VGU1CMDilQQeTf0jrsLIE3YQSmgXr5Vo
UCBvZsN6BhBig1QXJ8czYyfBucDiIIC9rVBb1BqM33EcVNjTW7WFUZ2nCVilHbC6VCW/VWqJU4iG
Qr6bGWoNoU3Ljk9Dq4vMtK1rgnSOToIofISjUoUtkqvXaPYCuQJun5NRg3bWEn4SBGi1QWUsBSW6
pix0ZgVem0v8tn9/bMy0jpx3HsIAE9EjB63rjqHATkn1v44QpeX/3F9yPTaMvCK0NCfuubQf25Y+
GqcrgnvmzLgRNH2UXvpdxvycnaV1duqs7t1FkT46U5qlC1RxVxIGFvNCXaLkggZmx3D1znSiaEZx
+M/U0JhTkk3HP/n/n0E2Xb+OrB7x5FB87P39jtNx5YirLJQzy9jaA3cz17DlwPpwMmanKNui4/LP
OOZQTITEb5d3ZvB6fUAwEySMfrtw+UjK6IolWaYukLzI5jO6G9XesYDUZJqNGV3DerkEvXuCegnZ
Id6OOJO/Js21OD+vHYxSjtNiGZr4f1bePWG/LxUcgUW7cIXw6PdKyK+p2FZ4Jtjp6KAIXEx/jWRN
fzAMtHcbUW/mvc1KcYa+02de77xznD5uQmnSmjugsh0wlZ3PDgod6fhtI5oWA7Is8fRkg4q8bA/k
qo/6hSdBRsOfv0yAA+5kVTnO4S9lUlqsaucmg3S+gyRWWp1UdUKDX/AXsKa2n7vfdgLZXo0E5IiB
+4ufCEdZp9mlLf5W5pKDfGwYgYEYABdeH/4+yErFgGsaoXmf1esQv1bqjF6zDEWbC2RSGazOVKzV
ZyZGofgcMnmsSlYkbS8DCpNdxWTCCmo9i5/KT3rxcmn4aBzoR8Y4tNn0jwL1/1uUIqzbuZSQDiwK
5eVxkqYwutcc9l/WOf10XVV7N4CIeXAVCgELcBHflFQVnZ1UsX/n8CzX3yedkNb6qwyF58FPHNDk
9T0MF9TMFslbqSiCkQmy6t6u1abZy4KX3RvmmFz0JXALx2rvsI9zi76UqPF6amT5mQbaj2liUlh2
BjrJ00IfQs71GiFJVL9Yo14DLMpEfH5l9ANU2vzMm7dYQXgIJ7WEjVWMtdN8velCIumzQSaSSjL4
bRHyrAnayXiXG9d+PDnfTmH4ASAssVjdoXI0HauMejJn5Hgf9ze3w5dpXFnP15ODlixbED3L3RZV
jygkat7XHAyFg+PeJ26qznmZB4H0mJaXoArBMR50CNtT5ZkXjZioEG3ib7ZspnjEWn97SZ8JRRjW
eoMKFJrQv7tFmYgYkdcg3tx5Xfyd8wyWp7XopFyUDlA595HpU9XtpW5iJbgKdu/kN0Iox2MQfLwu
y3SKMBFJ8D77pOSbV0U/kT/5XT8Nhx6mBBOcsNBqiPAWFy34k/BY0gc97++we90+8+KVmBVgIG3n
UZuJq4KANs3adNDU2JWbMcjO+ljgnkAdRr5D/nc/r48NddBF9zPQzpiU+hWudLUAYqbahMgkHFIa
wSZQDIvTuPQLm27LCfkYrP5CM/jsuKYUSbMUthpAhloLAq9aj/uig0tHbpr9hBnzZ+skhnj0PHn6
fz2LPYx4UWAyehvH4Sx0+BtE901OgDzHEUtNktbcjK+R4ckc4OduqguDJrkq9PrKBnYWClgRmMgI
ZB9rcO/HWhMN6EJLG3d85qFTYBCt7HVcrtac4cqEYgoiVnEIj9bz5ZuAhYuIHUE8PpxnhozqJL/s
C96pI60v4bS45pa6gsI+CavVW0ti26mprcKhRLohLJVyZerFA3prsx138BCWZ67LXGAXAjD/iKTM
o4mdzhHaYL6wtncGa2jFzAN9CUNnorOtpJttXwewnkBlLOeuiIDTe+JA/5ZPnFUMjkndku0iUjsN
W+ql05tah/nugdzZDGUU3HftwEzDTSlRvkJD6mH4BHJcqMZ1VwU55SUOOKJMqCzCA8v26GbDeb30
eTl1/zqpEA3MlAsso8yKQVPklfyiufMkyqhOkTMX8CsALLZ1acYQ5D6NWxH23h7a6K7J0mL69wf7
6z7yMnggabHnUsezR8aN7Ep5mo5hdNdgrkthshumeZcvrHGSq/ut/R4Zvl6suiyYkJ38ZoPiIvR0
MHTOTcX0gxCBDMfcBYXH8S0kkytNp4hMVZ4K0/ohfwXh1rYBxmkId3x4URcQxVJ+wZgFF3g5+7qj
6GYqpy+PtVMeBM5YprCVUhwJuyvd0Tz/CQdKMTowv2etmspMX8qRg9C8KczbU49EaS30hniinR0Z
T0FsLL9e5Imo2NFAmdPmeGbdicSbPIyqK/UfF582ll9K3/J1VUEIVkJeses8uBQTtojwnX0FdmpJ
/IA2Uy8Pi9IR+4Nr5AksE0Wz+ysJYxx9BB37gw3HS5PYCcF5pZqOuCR0nZerxvMCTA+aG/kECjNi
21KfcDouBr7dUUlCANtkuAK/Yly6tzGJ+827XpeAGWEGL5D5PTG7FeH3eR3gJHvlb3OIRi1vd7NV
1fA6qy24vdWiHyf+PZcNtRO4LiET5PtYx+Do2hInegLBJmX6Nyu9qNmjAkzvu4H7ipgRUv0JXhTv
pMt2PhjrXlVqLbDpH93P/GsyCcgtch/refz6jlgg1QH4SXIxyXYQAopJpKIpqApeNiS0bcUzYUQG
P4Ko9TWCoZhRZ9xtXKWLGP3XhcLEThYobiXIIiAb81ZxAXNC8bJKh9ZSTz321oz7WjOfqZvBe9q0
7jgr8H4rEyccGijGFyUPo0tOBp8v/AbJiU0f0V1hG1vfqzl+G9N5LxuB0VNJBiAPvhomKTcSsEUo
pfhBxSJBLkbDFbElPg0qKjihCblMoIwjSFW0wbp9ec2fTtl2YB5FZnQIzfRfFYilSEAhsKN/Hf+f
/VhmZiGR4zplkI+VoXOaXpt6/MO7wdWUEnPV3Tl3G7lEODdrMW88qIDGxPPnQSZVQ2M3qPtchiGi
p50q5dKaTW/ti25an0RahRGBb02UkfX14nsBNJ4SIXUoVxMOyUzgw8W310OsLw8X5nQNCA+zEqri
w2zsatVilfTgfsecZG6aiacWiCamyoi5vTAG1/gqI1DaPWRzbwgd3dr2vfz5aYJyrPKhbYv2Xcbl
5ditbjcXS6R2ZJ28I416ka5sZ9tY2PmuH1eip2vVCENUpjwNimtRaGy27CnnDZr8tZLfKCVWu0QV
Wk8eP/oMqF6UjfKYQVwbRXcXNUOZmNF9mRZrJATkcDDqVH412pyIM5krqXciuxOvathIOhEzokuo
ud+DCQO/iNAM3ksKuQjnG2BDBo3ZCUOEKsm2k0kgUCW+CwQ0cYZUM1920Lv+tqnbXTK4cXT+dOYe
NYayIPgEP/o+aZc9moKizGZ+n3S04ZICWC/k27Ae7TBF/XAl0OYmQxW41aCbGeQJrbKSdCGgcFM7
eRPPUEBKXMKmclfdl0uiWFfgmS+dRAFFQUIuQgfqOvQFXEb+tDYmRbQvQu/z0VTJrShJM8fxBmxe
rVRgVYJOpym+uXFKIFbN+5QGI1lfh0XioCb9fjtT8V6Dyi7mREHuwEkklorGEFLp1UIxhDC/oI5h
Bb/rLev7rmcDl51HSF362UaB0gnb0eEAhRg/LyKOOPRSdfTwKySQSrnlUzgwFY8D8B2/XH3Hggxl
VGwSkO+1mfokFd1tNQYA56SHedSi5+g7y0pKPZFt8X5jJ/kcoG+GShPbz6nIQ+8hrN8Eq3LH4Qi3
8p1GISmjh1XJyUAmnRCE/xsABrEVDOiMtAzWYB5cZN/pxhZQX+VRYJbynQIOx/SnmeN1pEFcy161
z+YvPkFH1CoS4QSKkhPUc8ynZkExSESuw4I+d/tdGcGHVsrGbUn69tdFb7X34fr7pyWVn3gJnMWO
fAhR6CodkPiUlv7CMOVMK3TueDyobOCdouWun1fxBbBrW1aMfNjgj4SeVTcvb3T01osODn+mzuIV
fD+6a55Ibik6G2hf/iA+mVTmqW1EzqlRBjKezq7yIynzrdHmU/OVyu3neYfc+404XVBFBmPkFjLF
G6QeE8bqIKFszQroA4tO54AeCojgiSGny/lYoO9YHc3oGB4CSd228mrLRkPNBLQEaPZ/c7l1YDCC
EVkj0BmZW/zPDC8/tepATVQnYvYtWa2u/sTVKEZxkRu29CeklfCy4K1uufrNXGZkU3BNZDXVxZ/9
ESu+8fC5f1Dd1/9Thv6w/bfF6CnPdZuQT54xK5pXzK7Kt+KXgjcNb2LNYwI55PEBbZRYdXj090ds
Auftq0SRSqBBHqkmLUUKvdbx6CGI6F5Gq+AFpDDjl/2xjE7ZQsAH24UZLS+2duJ3eVkEMeHhI3ap
pUKWnXouV6qZacl5coEJyufnxZUsTF8O5gFB2oH81+YmCiw25R1eA0oRNU2e0cmaQLZImQCRolKv
Inhnzp6nxigk//9+AWFriqMFZ4rTspqDUY69NV87z/tnPlL51UVzTQtw52kUeFo/k8z0JGQPsP8I
bO8R3oZGYzTvXSMMCu7YaaieQaaGZaQIrf5TMY0Bm8TNGtI3di7bK2dOciSSWTpIqsSqsn8nAJAM
mK44fllS0AFkIEODNNI9CBoF9+09N8iKq5naUYu5QNL+WvQqbV4mp9QuMEQdSnZpxI4tUsG0/bRq
feQDnY2Yof9F1LDVFTrWDjvJPSEapdhSsZwWO3Lw9CPuEOLivNwJGcVZv2f5IPFMz/qSdatBovY0
zNhTK1L6kgu2ya5LX83yoorUeGqcGZQVAP69+rilmW34ynGV+/P86SYxqSMaEAed+eB8tEdzRm0Z
QTqP+3LdH5elZ2B3p4JxwoHJZ3OB3c2OMf7Dn9UqO0iKoXFt13hMBd0OAzKxM2g/XU1F9fg6z3Uj
XUs/G7k3RYwGJjHAlX+y/hPQKMNrAEQcWrFtooZMRzwBx0CFDLkgX0qK2Au5mSWg/003bsug2zG4
PpXA4EhzzOAD2S2j1FB5yF14jMxOTwNLx55AB+F4kS83+QhoUrNNZreirXQiB2apZIH7yYEmmY6F
GDEvPjbl1FvX91RP38lydJkjVDM+HiOebUUodg/dBsHVvSTjNpufRjpi4Exyi4v/43skqtdGFzX9
OdEvvhMNyufh0l8UF9nMPZllLE7X93Y32c/n3MHp2itkLneWM0FgySkoAj+Z5C/wILGdbZrH6blH
OA5csahkpa2i/Ih0CcXLFLsOOTUtvpdn+qiYJgFLMhzu51vvANjXeQhjPtAq1wmga33UH/akc4Xq
wvUTRSNqO3xfgsSSB5/Qms3Ah3j9AkIGCwXbTbw9xWWBemrlg2Qr44oX/KOkjdptqOjU9Z/R5jO2
oi2bE1cA3aHOTmmPBqnDefbxkpa5chL/2XCaakkxLgH4q4YGuNnjgL8U6LbXIzPYFFcsyfDocFeX
i0DTWeLS++qtSllFisiVGZzngcWenvyxeJbHh1XgT1zvORR7H9Ve2m8GZD0Vd5tgdw0f6sCSrlzG
c95nzP1I68HRvUOfNrIMEid6dMqEEqMyj6nnf+KIVP0/RO8fBOob8txaEH4ZrERHizv+g3AtSM68
pPePUj/KgVUN4NfeSg9ipMLdRTeH6zlISGwlg5TiHIytTW5OxlfJgcJdurEpfn2XmRhqJrnfrxFn
7ltZPyGGym2/1Qhws+sv4St2mM5/iRqjNDgMDt+eGjRZ2LSsymXGPsNTTIw1GsChvkWMQxZjdogu
dwJccaWTg5tkNM6IGGVj5z6FRQjzjU4DoCF4MtHzKRHXvYRubcIgx7luedoeD+VYotCXq2Os1rM5
CNzhdyT0/KCY2L4ssyEYqLyqQupBJDDfD+LxyJYtB7TgtIpeF3fupoM4SS2Tla/x0KJLYHATy141
hLhkAKOI6GRq2M5JEOHt5cW6JInGMWy6M9YVD48dLBBv6LLDvIjzdXb0KGzD02hPjfLjYMqWcQNk
siPVuFwroGsS/xhWqv5H1hwSwMk0uUxrC54LNXrwVnewq7I7Hw5YR7v7VygoRLYBQaYYZhOc8ham
3VNp22byuUFpbiMsydBq2pPIpLI1ldzetalnX9YLm3eB5B3xm5r0oavwCrZTuTm808rw9R10AFVm
YgX/pYesrAqCajzKqVY5UfFnbpIRIX5rTt3n0ae0BiOfmEVPC7wcGhPYKZJX5gM9d929hnxWMpZq
fdnif0E00kKJ/2uIlFFCwbU3AY3NG70UgWrEzLW97r2+J+x8xM/mXpcE6vJlen0rQWdd0P90qnxQ
K4fIOhSblBw43yFGqCecLVIq7wVW1PsyfXTiQcHjqRPM6CabCy4Qd9Wi9OzKISD7ADlUwYHCOOgO
xmZ+ePif4XEH+NPCfUPekZ88oKzngrqw9Iee9nwvHJSEpqv+My+xvyLCAZkEM74rZUsjy/XIZq4Y
CIcKFJsKMT4X/4oS84u3KJq54tsLau3cB7OkaZIbxWcxEP1Ln05e550nHqpv35rKAZzhCmbXMWS5
UvepnIrinVPoIhfJygsdy/EIEG87FB5NMXm370lvsd86hfK8r60Oevfrw3qb+my7VpEQjOyo0dck
9AfSsanl8vsPzuL4763uEpNhbn901ICMJ4MxnA8HZeW+BsabMQLq3bisZ0e32DXRUdt3rEpwBTpQ
55ifTEbsjNXut0vx5FZGg8svs2MWWUbJIxtnx2D4gooFAn7vQZ7mwa4Jkkp8T+x9KdWEtF3U6jtI
PElOCrpstkrNIR65EmGPWHXa9vriMACyuPi9RJkZhcuS5aDxq6xxTlv7+aivBlNdF8AA7o62gTQo
Q8d2KGCS/tqXu8ZpRP3jj9l9NNZJjnqrzkKErDBDDbF7G+rHo7WzyuBGB6Kido+RR07/53mV0sdS
bgos/ILIDbKWJGTWA6AO8nW6tHZG7Lj/yPDrL1W0En2Y9mZeW3dQ7etIhSfU8g9imvVyiLp500Wa
jobGg9mt3fz3uTZkDOd61a82vmTrTaAfGZBA7Fu90cwwUfd8Zvgf6WQSWXQxA941L/zgOAXv3PVn
7JUVRWiWcexvmNChvfGq5BcTHkATtXgXSjf3fE+cKc9FRIPu3ovzNPSq+kJaoMBb7uHwwBEmiUY8
8Hr2eHnq++XX4wiuGaaqskKEB4aUIe6r4bkw76087mNnkEBjP5jUWASRw2JsUyV2bH1kDYtrDu8m
W/8Z7Ygj8uFXM6FdgjWUys47FD0vOOJA4ErObM03x73aRHAU3ICRlqc1te5ZSgp4AvLBvK+qVrZC
TfyHP2Fwu19tP6HcrDJyzbmulj7uxW/eYmzpZbAs7oG83AWxve4x6GNcNNutJyrj9updki/HDMzi
d5tfKTwc/LWddhNncTgkpzylI1z9s95w2N97BXD2Qa4nyLGb1ejP7wuwrk53f6byqXA5H8r2rkOj
JXFNYBTn7K1KskWo3/Zhfa8AOuFIrFAmgky9zfSliNdgKpY2/+GFw9Ih0rO7yM+ROyqTJHpeKq/i
lqRb4gRCsJ08Vi2jFM+96PpWWOaEeCDmmy5hfIkjN1VFd3Sc9e8r667FYV0zHDAUrRRavKGLv8C2
qqNG1BOtxUcsLNnbX8P1qnQ/C+FGembVbuDgyLugnpkyzliYjajsRhPcXDu7bSyOmpQpDzPlTZMf
aTTiOiz/PC0jHxea7T1E6hNWR2T2BMO/RVcyNfUb7deRxvL49mlMOzIUGZW22wpAlJWuJbCF9+0K
1bEXVtGUADNQLEIXYE1QtUGE+FvzfVQV+Vf/bxry0vjh12pKloe7AFa+KuXWWQBkid5G8KT3fUxS
B4G9HU23UAxRAFfjDWwRtuxsFeLhSH8D0Ymo0XZRtiRVYuAarP2ax5xQeUcak/dw1N6HoKjGzASX
OP6cbxBIRx4O0b4ccZteesqmEHQ5jfo9ax/VyZIqi6rf+8oKjKEg/FVdQnFCxsjrjIBZ0+YEgLZl
/FQK7SP6C9fEnmprYqtR/MmQIl/fQtVMh2xKDbKEd6x5evs3ie5b8jgCjNmPRJhfAuDmZosZ9HXc
C5gfcA9u2gpFmCUTgSvkv8Vw4zvYC46r1YO0OL44hsRT9CWcDv9oF42h+ii/UGcYx5wEf6JMaw1m
RVk6/UjuUp1ZRwtvnDoZ33VzCcCEjF/wbhdkVaGmfxgJ4Z2Ncrs6TdfwZR5VLs5KVIYvoIFmfir3
6azIbK3f6fPw5BY9pTCfQt7Q82VesPqHq5Jo9pQS5nnCrV+UqZ3LcS2SExTqRPbLieqrLoFe0MpR
SMciQgdL1pz0WZpVjt7rpYsEzN3qrmPNtDPVk84uo3XR3yhd6Wt0Xlfr1Bd4CQ2VdrC4k7LZOMSU
7RfUJwaAeCkRzp/EMW/YdwiBRVUuKjJ4F4Y6ow3fpcVSIv+MeV4FXpJK7axTbGYVpkFutBRXdCzI
FvHRUVGqy1+OIsJT81yBTQ0O7fJIpi9F22phmG4YqS7J6X85rN3PSSqmMvgPCYaVIJ3STEHP2Lxt
mCnKfphjoavhthggE0BtlkC+KzJ3ukO6iE5/Wxk8rMg3IIuxQSer5tLv3+4O6lL4jPCwCdjQ
`protect end_protected
