��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ДėV�ކ6�>z��3>�\{���Ҕc��z�JT����p\��4>�1=�������b�����S�57<�@��J�\��SO�\��g��5jV9y��6&{r� �/�:�]�fG��2�E>�E4�<9o�uX;���ލ���9ɣ�K����Ɛ�׏܉��F�J}D4m�[�b�� ����h�Sh��1F�2:Eř���v:V�7a��ku�ۋҺL�ZZG{6)*!Xf+�z�S�z�� kP��~�0+�&�-?:Dk<�GE�� ��Y�[Nr�A8����ӈ
u��b۳Y����R��G�*C��ܹ�YGM	-�ʞ'u���>�^Oc:�l+�̉!�׭S�,Ni��.��)��}[��ˉSP(O���>�� �.貄ʬ	��u��|pշ��n
��ȩa4�i�f��]�����^k�o�Π^�u6Q³�>\���϶�,g���S�-�����X~��u-k���&3k�,@�MZe��Jy[P\_��J�RHq-�\U�lІ��OJ�P���P�82r�o�E���Z!S' Vʯ6R.�2#?�x"��<�\s�)�肻�٦��\�9؀���֮$"��j��0����=�g�ݓ�N��$0��e��vVR�h
��%�?��́�s�_�R����UX�Y�P���	:�l�<#��ܽ��+G9��e�R�H@������⣈�ε��]s>��֧������A8�p���E׀�[O=���Bd%SgY%íU$�$��B��cK&�	{C<F[�sT�!����|0�B������_3>�;���$Vm��.����4;p��G��f��to�x/�����yqJ��t������gZ>���D*�1�cH���T6jz>�'�=u�;�m����Z��+-�-�O��$��֩�1�r;K3�b������Bt1��-{i�*:�a�X��@��J1ٹ٣p _��{
x~�������^��-��p��bV7���'��\��=\�<b�Ő��*X����F6�G<J��Bv(��ׇT��Yz�94�x�T�h�!�Yh�P���-�H@�Yl�w�ͨ�8��fU���"z��PyF����f�~�J�EN�Ƣ��~b~K7`������_��[���'��O�Ȏ��~)�$�U��"J�C��ΰBHM/B�c�DuX��`��)a�Kn���r'���ϼ'����M�e����	bjofE8���4՜$��,����RG`�Zp�h�⊢���hS�E�%�@C��?��]G��P�d�^�x�ֹ�8n�}��G��:�FB��(��bb�Õn�mVGpdD�k���8��Q������q=
ĝ��`�P���T�{-v^�@��P���Y��͏�ȡ�ޤ*�l2�»
�V���8L��+�.w�B�	0�7��]A���p=ً�(�( t�UaqVd*d%�:��J���ލ����O��*us)��wd�(v
B�@T�I��:`��k�P�X�ͷ�a�"��Ӭԓط�O���#¯/^ŭ{@��Ӷv���c�p"��#%ȁ���b"�qU�� �� #&X>��e�w�|�����K�3�;[���\����~�&;Owٓ��V�4��.��2�J��L��͉�a(H��(f�l�D��s�.�Y�pAi�D�[��L�iU���ޒ�H��17�5�M�����bՕ��&Ը���4{g8�
'$Q9x46Uݟ9:��%�j6}ߎ��Ѽf�֓)p`~:�!Y���%
[8��ߍ��i[-ݶ-"�ϫ���s�\�K`_L�8r�5��0�-�0��z������Ε���h��˛h��3��FҩQ���G����E�% �)3_�C�c�ؿ��_Ԭk:o��� y����~��vό}}��"�>g7�1��6��`j� &R��b/��%OsIC(8�~Q^�	�i���RF�p���B�DU�� /-�d/���F ��7<tA<�o�O������P�b�M�,m�2;6�A��C{ZBE5��`�23X�S��!H�|f*�p�����ٹ�ٌ�"� f�d�z�����dDY�+����t�xiN��?�4��S�p_���9~�����Mt�%v�P�N)^��&�Fl���@��������d!��R��:/b�t6Ρ���&��W��4�J�	����pu|�Z��#�t�iC{��R�o���8FR{%(T�% ^�#����y��(����+�]����8���ބ�U��/"yk��h%�d�A�њ��[I�U��V�`�;9��1�ɸ.(����~2��1��F�1���4L�h�%�bx�+�3�L���γ��
����se����֭���0��������&p�l����~��R	�D��>�<^��kM�H���ڴ�;�K���j���,�]f�h�����6�Օ������Ni�z%��T�6Xu@'2i�[W����+YH���6�P#���Б<�c��u�x{�D]��C�o܇�5@@��B��8b�x݊'k��	����X	5�����3�aV� ��+�+h]r�=��H�Ӛ��)51�_�(��zr��zS	R�iA�3�.�"ke!��5kOP9w���_�#�xM&�G��mYU@��2���(�3*:'������ P�����e#�g������Ӵ����Ȩ���qA �==��тr�)�3�,�-kMh��NA�?Tۄrs�g#�x�m��&�qNs�]���?��Di|�E9#s�&d�$:+?�g#AU�� �,�������)SO���Q&2��E'�m�V̰�ǌd>���bQc���?��]ޅ��)7!��DP�UB�o�P.�����(2�B��)�L�3��_n-9@����_�3T�Oo�QkQ�U�x�{Q.�	҉��5?��i	��T͎�P�:a��7lz��\���}�V��(��}K��Ĵ7[|)�CIl8Q�<oQi�v��Q��Z�?=�j9�g�ef2�ʥ"�0��l̴�G��I֢K��#=Z�w,'	f�f@�%|ި�oN)������TSK��4v9�����������>u��& ��=b�k]�y�>��N&2�����EH�wm�i7�{��jN4��p�M�<᱘%�@�/�XT�.��%��̌��󀜡�{r��l(G ѐ[�D�3cXY��T�y�m�IFf�*���CC�a�s�Ebn��b��>fs�'[
M ��to������p�U���J��]���/���˱X�Y�]K>[-%����ǐ��T%1�Y�I��޶t/�Brp���v��(�[T��eK�\�b^H�*?���(+�t~�NOUa��!���.n sj�6���mn�z������Z�2�?��_��1;;���S�q'�m��:���7�F�1q���@�}�R'S�O����@�zXE[�d�x5yf{�l��&a�SNB��Q"<߱�w�&j�R�P��~��B�����X�3�r�?`,�N�f8�mGj���&��re0E���&�1�k�ek$V}�t�t.�*+��Q@�υuZi��v�{V��%EZ�r������r|܋ �\yVp��pla����m���w�T�}��Ҹ��M��2�-�f�m/L��:��߿��[��W�xU�-=pyU�·5I=,�k�gmE��	°>A�D�C����ȼ���42�}�-���7!�Y�^c��`�Y-6��
���1�w���N+�"'Nj圖�b�YD�y�Ľ}2� 0ڹ]�v����=lôFE��n�G�4��&PH�����pM8�4�d1=��s�f^@����m��B�`Sᗭ���E������8�Yl]�����.$�Ύ����I���2���5�����X3lo�ӽ���/W���;����D��A������LM���#t���D&��@Ga��\(95Y�۔b+`����!Hbv>t�b��b����_ѿ,���B�E����!	0��2O0(9��B�p�9�Yf��z8 .�!��=�>6�-�4�N���PD��� 8�1Ш��؟N���(K$}�|1��\��!6��3�(T������k^qm����Q�f�g�����-���;���3Q��jd^� Q:���Iy(LY��%q��^5ӓ��P��0�m�j`�B���ګ��l;F�D{����6"��?�"J�\#��a�i�8��1X�]�QS���J�-������<.��T��r?���ӊ�ӭ����B{�Ťm���n1K���%:,w���1⥮�*��X�X �]�CUEDє���P:e+&tMׁ��s����p�׎1�b� ~Q�n@�I�#�E��􏱠��|e�+������9�W�
�_�*�!h f�tr6ElKA)i��"�@� �������������:ȍ�O�Y�����>owx8B:����S{X{�p�NDrx^{2��S�ͨ ������
�/0��~і���~�O
S��=+cRd��i����k�H-!�P /�Ihu-:YH%��"#�@�6�sy{Z/�N�[{��)Xc�[q��r@$�_�bi�ڟ_�n�F<�G��.�c�]mN�k��o�k�g���:���i{8={wM�jt�8��`�./G�J�,��1ϗO��)3B�6�}�fYzn^'w2wY��R((ȵ�۽���T������(SBj��'���#_M�]�f�AI��L��.�;�d]m2����.�sUTk����U��+�*.p(�&$��^5�RJ�􁐒SOP����ᚺ��$���#`6���T��-]�<~&D�wM���x�m�9NΫy�A���=m�2��yO�s��^p�"��3[-	��Cj~NX�ݟen>�qM��SO��8�faq[������L��Ԓ��q� ����2���׳e|�=��i�x&#j�}L���1��}tъ�[w�ܐ�K������!�k������帔
�Ҏ�c�K7��F� �\9���OZ�3w$�4,��Q�M��gNw�r
�YOW�L%��h���Ό��gكO��.[���gf͍��;�iڻ�G��<̎e/�or���m���'��i�Yd��͵��]cH�U������撿	�d
�5S}"j�t�ٽe����!�-�o9��J��oV��;��V���B[�+(�{�ns��� Br�����7�o{�yJ0�I�*j�W<���$y����m23_z�rA�!��Q2�:��P�K��j���<�f���Ig�ß8wG�)ٽ�*��"97(��Uhz�t҉ˍon���~S����Ach6� �뉘�͹U�MС��ca�����9�^0�(5�i��%\��x�3Q���j�&��o�ќ��_��Q�2�ÿ�Y���Wɧ�<��:��m?Kn�V��Q&�`8�*���늛�n���V0��wԎ���|ʹv?a�>;Of���5���6sS�i��9��S��g����nH�H�̼1F��DP�Q�e�|��bx��{�R��zPԹ����������M#r4yw���"$D̻��E����xM,����n�J�Ƹ�ʍ���a��C�6*��Fާ��h��0g\�@�w`�ȧi�I1��Z��� mM����E?7���4���R9B͉m�e�X~G�%��?sL����:Y�o�?R%f5�ȳM��LbՐ�A4Q��O1���N��] ˛u|b�^��$�����
��ɧ��Ix�Ɣ���,�� w���\����R��C�dwM�������"*����ܸ�ж�I��9/�g�Xuҍ���R(7�j�z��Y'k�g��6�i����`��y΍*��Y�ݨ�^Pm�^�uoXaۭdwe��|c�������U�xe��9�gt%Z�
,��֨`���QV��NK��O�K�xyA�5S7�]�X���zz���kx%
��׏$Z̛���J1���?9�!�N����fʹ|��Sz�=Bo�0�%Z�RVw��$՞��l#����
��xF��l���������Uv�8|fJ��'=����Vo:,�h���vȎJ��)�<��(>�N��b�
��0t&i}���D�H#�*�C�>����S�p��6���{��-����_��I��'�Mh���&���e�1B�Bڴ�GR���Q��^����?��P @n��ؔ�pYu4� �1�{���8\q�,�3؉�|�	=IEV����p���c;WO�.}Y�����-�A��H���I�;Rb�JYt��/ԗ܏��N ����*�5w>U<��U�e|0F���*#Ǖ+&*"V�h�ss"yy%�W-�j��Y88��gՙM$'P��F��+�&",x�#"ힷ��A���:��]�v�������g/o��"��A����7&h|�c&M�曗~F��F�A3�W|��R��׿����i�[o�M�+���>�h+�?^�y$M`�] ���0��FtL4����kFc?ڍ�a.1{*�}���D�]a�o#�NѢ�F[� y�</�w� � ���wx/Ŋ��������v)xsM���`�z���3z,X9y��g=�sf�Ή�N �3=}e���~OBy�)��	��寏.}�ή
cN@��0u��t���!Y��L��M�/5D<͞HI@��$2n�U\+*�s~�Q�G�X�$w �x�����ϸ��^;-+�O�TW�-��t4rg�8DnN~4A ��D��W�I�L/n
�N�a"��&�qu�H�h��
�Q$Ms�e�t}��.o=�BJ�	���Ъ@M��ih��&-ڶ{㘦"�^�^��p�C��DD�q�[�n��h���N�J�[��X�Ӷ��Ó��]�;� ��b;@�� 
�&�I�c�f2��� �yQv`@v3�)�?��������D��f�Nb�6��������	"}�����Ε�Qî�@*��
��'�%�U8��DI�©�� 'd�2ӿ�����mЧ��_���U��O�2�"}�c#�˘���WX�W����LNс������.ծ8 �/�e�+�e_�L&��8y|��v�9�ͷCgRG����EJMm�DXt�u�^��TS�߂kx U?+�s�~�C��nj*����n��d�?�DR��5ax��n�r��� p��P�^')������ɜv��b�.�/��Y��i�G�U�9[~����S=u^
|�W�t�=":��h �r�����1����)������y1%Z3����B�L����R�Y*8.��Ȥ��o�'��e�R�$���` �&��}����"�Zr�K���P� U:9K����Җ��a3����,�}"B�3�#��$E�N+{".�����z����MȻ�'�
:h5*I���'�;H�l�Ġ*��N�<��4�0j���M �aN��7A�P9%�=��_���K�m���o�.�F3�z+n^�7D�S�y2kk�3a���o�g�Oq.x�	ʂƍ��J�<�,��}%��Ln&�jc��H Qk��tP*
OI�'ef=���<����s��6�=�B&���[Xԉ�A� P=��#���o�gc�����L�CB@͆�+�2�?}9�No��*-� ���)�8Lrd���ڇ8�������~�䶍ݲ��xƟag󺦨Z��_�Ɉ�����޼��G�Ϻ��W�f���φ6{�	"�ީ�5�m�6]p.4�����ߑ�<���I������Z	�`�-�B�Jq�����2�c���a0�"eR��S��'�=�(�D+��'�י-����xA�hZ�hk����RU+a�.3h��=e�� ��E��h�2���-�+v�)��+P���������(<���E:�U�爌1���<d wtg
���]�3�DL�VpEYI�4�ۣ�ZD"�t6�L����a�!���
x��jGaDr�TX�4|�71|_ u�5"%\��Bat9B庪��:EKw0v��QB���(��	/fQ�����A��A�g1N�,���9�K�'LW���t��u�eg��խIk04�R��s~I��fZ�b^v��7��:���6�#y��F������*:Ij�����&H'R�N{�<#uT��V���|'ܔhd�~��!��Ω/w=	 Axٔ�z۹���(.��l�П�x�i$�#����l�"�j$��c�k+#Oܪ��^tq=.��o�?�2��@T7���6�<+������C�.�d0�Um�_�#���D.`ux�8ڑ��Y�L���ɠ?k�R�����V6���D�j�둪��� �ʴ��{��}!�E�3�V��4�5z*}]-hٞ�7�����)8N�9���}_?�����§	q ��_]���dR��ی1�0rf/��o�&9�ZH>�ׇ<7�-�
����G���{�(�g+�6x���$T��W]���k�|�����؃��|��
pe���\�5�]`0���v��R��E|y�Y5M��zl&0�6$C�`1i�H����}��q�ݡ�5K<�������ߨWd�\���E�&�$;�f2$_C�m�Efǿ�s�c#��M]��S�y�
��X,[ާ�v�RZ��)�Ҝx��ü	����Y0�}=�!XΙ읧8�0��uV�WB�˂�|�X��Kի%^@ tD���	m2�\j��_���L�"o�Z����N,	NnB;�r���n�<ȿϯK�\�/�����G 9n73��ϲ�^9�O�24��	j�ʍ���2g��uM�Q��|�D��w�l�?�3W�����>e�@�*�)�;?���eڥR;���b%���4P]�4
�f���޸X�ɒK����E/���Zz�7F��u�vh�Y�Sc���y�]�� ��3>��/>�xK��,y�~�u\-�8T6^q�(�ţ���n����bI�y6���a Z��̷XS�h]�W��AJ5�����~Є�o��4?�@�O��Rĭ��Y��0�������Gc�q~V���&���������|�;��9�����kˎ"K(�Y:^�9y�<���l��@=i
5�ԯ�?/�����[��=̈́�b���L�Qu�h�|��֙+C�n���qL��AH<�8o^���ߕ9�&<�JjL��O�&o��?R�� �(Y�� �� �)��h���&�(8>�
P���#�$ԇkBL޼ibE��4a�КDU]Ӂ7$�3)�?�Xj�i0��(�����^��$�`�z�-��wф)-fh@�+������XS���H�ʝcQ���4u���a���p�I�Yω�F8�����`��)�1�A�%�7]�n�m r��>���b�C�����7t���=p���ݷ�J?��~\bH���B��+g�i�!ا��;4�-�2�T���/B�k�Sj������j�������
��M+��
�Է,��>�45��,�/,-ETp[�./_�zD|�9�ߘ hC@�	|&�!�������c�D���U��u	��9�]��ʋN��B�ux[��K�j��Ĉǹ����J��p��[�\l_ΦQ�*͌ԯ�j�t�� nK��Wl��6�?��]���魞"ڱ��~�w]�@z.̪��غ&O�C+��>\9��T��{ �Y�����������`��Gg�֩�;��ԉ���_r��yr��-b���t&]��N�zOSv����>��[=U�\���DN�W���*؏hBQi�-�5��Jd5@m���W>��?�ߤnGBi��^s�