XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S��_8)a�F�x-���w��x�O^tP�<c0@0LR�|�Y�L������|����΀6��L��Jv]T^���Z��eʴ��U�nJQ$\l_���{x
�m p��5:4�~��ʳ�EC�ܤ��u����i�1�[��>��>��� �s.��Ÿc�\If��Jܱ�Z�v�7y���a�u��	�^��݁�t+��`����X>��,ʋ������ �a׌u��1�?������'K�wg��r�=�&�%���>٠�.Ҭ$���~����Hl�/1w���E�ݒ؇
�M�pAЕKUQ^V��ks�_y��U�PF+���_�|a��\�G�ζ�H�[7�L����Dl"X��W�)��@��f.�4n"�U�BWM���bcq]z.a�t����)¤�;����6����]�C��N�����''�w��F�%tu.��|$/��I�n�O�?�ߤ��߾���R�� �q�F;~� M��2نZ>C1�!�I7���H�fE�e��@��f��昑ҭ�f���"? D� �`�Ow�T'CU�,�k�ԴK�v���UM��`��v�(�,�".�2vo��=&+����EE���\�/D��n�-�n�wD�W囀
�1���C�U-Z�<J�_�e�x�R�7VU�?vҎ֌�(0��aч� VW���u��y��V2�[zA�V"24;��0�۽D��XV�
���0m x�9#�:l��U��)����3׶{��ˑ�ZXlxVHYEB     400     240�6�y/�uW�@���\�U�a这@=rZ�ʀ��f��fHCoo�O4�M��sio`���q�L���Z~�?�6Xo�������
u�3!j��$EԕB�GTl)���f~�Ɨ���ww�;a����N����mz��LY ��#5���ΨAS����_'�ѯ�:URq���BZU�}K+�c��TO���]��BH����x|Kv_|�	٭Gt�6�/ݹ�ai(D{݃_�V�=�Cӱ��s�D���i�D����ҙ%\B8�����?] ����E���S�Ԃ��[��f�5B�;F��Vo�P�ξvﶁ�R�К�HB�&n��:��G�əa~�E������m��(�C�
�M<aG��%�Rp��k�^��s�lUd��b�p�z���|c�3-|�Md��J�]݊�Je�%3�M��	M��F.�| �#�J���
���\
�ݾ����2ʩI�"CNI�r}�F6���n���G�'&���J��!%q������H��[���1Ŝf�Y2	�>"��OBɪ0�����v"wK��TXlxVHYEB     400     210�>���6���Aq��
�}�z��J�6Z��Y� ?׈����gx����?
ZGC-7�ܑ�V#�P��yN����
�DEw��z8#��tN9n^�XD���zu
>�?t;E���ِC�����N+!��?���18L�0���	߸�MM�<J�2��Y�j[�D�#Y�4���2����	��W����%<UNL�ɏo]>�zR����{v���p�߃'�$f1�錗LRL����s������TS�>7������y~"#H��7l�Y�XR�
@Q"����э�Y��2i�/!<�����z��I�?�e%�w8h)��	l:�zf�$����=yL�+�y�O1��Э�C��>�Rk�Y��!�4���9ө�"w��A����'�r
mvji�Ȁ��V]L�\��e�,�3���B�%tP4R�t���Q� �Q՜L�#�5a������ +��F����(L�I,�x1+�7͜?��D�`gM@�lFۺ���'<XlxVHYEB     400     1f0L!^8�_�@���I숒��q���U�?y���b�sh/Q�~("�핎p,���B����W�*��AG�?�,�.g/9������W�V���P�S�L��M��H9�4�}/�^���'�On�ੂ:	�E�߲ZHӋ\�5�N4bΕ�[n�<�Yw�S�4��Z�"f���-'���1!�(mB�װ��Y)�y�U!�Ȱ���r $��-��S��G��gxn��9]��3�@������.v�
��'@>3_'����?���t�����7%��T��q�k��������Ե���l ݄ޙ�}ȴQ��:H�붝avFpu�gLw�׭�����&l�2�*�&1��R�Q�����7��w��*���Q��[�֬��eҐugk�c;��T^�!m��D�td���R�SC,:�#��
}A?Θ���+��Cԃh�f-�ڳ�~,��v$�8�����x�GG�Zj��Z9�-	�U��}�wV���ZXlxVHYEB     400     1c0Z�ֵ��Ջ��X]ڿU��ʒ�]��F&��*�tš���2�A���ˋ���a��R�6��Fl+_r%=7��ξ�����d���Y[����#��Dу<�'�s����E��}�|�@�,�
u���ӌ�9;$E�U�(�.,a���[��o����Z:��+؀�9t{源��D$%��6J5iI�����pN����=���WBB��;?#���/G�Nbfcv�n]#?�*�{Ǡ����"�U!8Fubj
���o�� �_���F�v�F�x<��pO����H�0����i�7X���#������Ҝ�C@�>�=�uX���-���j1�o�!ȟ�n>����)E��eI��<WGg�6�v���|*c���aɌ<,�!]���0��X��Cm���%�2�e�G��d��t���k��;x�5�^�ܥEi�]��:erQ'�w;�rIXlxVHYEB     400     200��1I�Z~�J	f|���?a��L$���z���:��!�,���ѓ�4H!N�G]ܝ`y��ѻ�	���
.�?�����َ"���Æ��q����u]<*f�V}ň�%��iV�X�!��� ڴ�HK������wέ�Ӱ����Uņv+\�`�%?=k&(��OM*pS��,�[�5Dgln��ax��s��"ZZ��C�{yos^�P�p����C��(�
�vMW�9�Ϋ�.��K~/�{`�����U�e� ԂM��z8j�!^4��3�Ye0/�x6w��j���P�� �U_��8�.x�d��>X��|��&)
۹���sq,��Cp0X��l���s6�X	\��0���"M>nL�yWA�j��#���m�4��dr�PT0eu���u�N�d�,�'[����2a�0����!��};��#K�0
��� �W��<~&�ۡ�ZWY�w� a���Qj���=�U�Q�C�����9��`���Շ�J;�ʺ�	��d�A�g��
�}h)XlxVHYEB     400     120N������@��y�^�(5����n�ا��8A��I?�ߐ�cՃB�vم�e1���٬Oڍ1@<�w 6�k���;4=N�����!��=�T\��K}Z1�ƞ�Ɨ�E�6�d�>Q���&�-̈[2�@�f�aX����#�n�^ M��F�9���ðo�ٳ��K_�.��C�ߴ��U����p���ߞ�_+�ȍ���2��_C.���q]!d�)YQ���Ӗ4n�TDH�q�u"��w�S�k�?��@����	;��̏
k���U�n{1ɰXlxVHYEB     400     1a0�V���Oa6D{I��8Å�7O)��}I3Ag$����y��5 Р���j9ֶ[<%���L��`�J�����Y$�j�����V����G{<�t�0��>w����]>����UѼ�C��=�-�T���W���5�}L�;ў-��`W�e�7���ոEy�F�m��#y����U��r��.�V^q���v��8nFz������G���S��X�0^����)���4��m$�|�pN����+���	 �"F�!����j"�a�S��96��L_�PhA
ٿ�w���7R���b�s����}F���jR9r�Q�&��PI�t �����i�PA��"���b��1�LZ�=Y	�*�(�3.�vۧ�:o:��ܱ%4 �ک����5o����ԫ�s2{2XlxVHYEB     400     110-
O8���vq����)omʊ��&i:q��6)��������4�6���O�\ׇ%9	$w�E��]�T�'i��̖c	aՅ�_۟_.�(��U����s���'U�8y�#���/��k����#��2�*
@^�N��C>�2����)��Đ�Hv>Lӡ�lY�K�|K>�C���uЪ�78�s{�^����H�W��������C�m��#��Hby#>8	����شֈ���!ÀA��$�SJDT�:w^2���r�J�;{�	XlxVHYEB     400      f0I����3����Z*�|�sտq3�NT7�P�9՝��1Nf׏ʥr��Ɗ����܁��h5d�$p!�:�ؗ���U��b���Ӯ� �i]�O�7v�Hx���g����3)IC���fg~��u�٠03 O�';�(���D�{�,�r�q����QؒRI6�݉����B�]_F{Ibf҂v�=�0@�~���zF��0/����D��~���$��c 9>I= �u<"� �XlxVHYEB     400     130�U��.���7�J\��ڤ~�W��
+H�FWW}4�hZ�c$q(ʯز�Dx�}�/"�7%�$�Num0��&��v�V�}N��r\^]�~qH�Bg}���� �nJ��#����I`��U�i�u�jW���?|d�sJv�F��E��*ge�]�s�̯���c|�H�KW��r{6��7F�ž�]0�D��b�UB�}ST'�d��i�a'ٌM�c��L3�I]�&��w�A&F	3��o0H޵������M�4�"�`�ur�R>�sy�9�
y5UA܊�"n�W����XlxVHYEB     400     130�m���T�4j���M��l�:Q��x0h�cP�F}d]���Qh#�nS�������ŭ������z"s,��"�����x9~�ͭx�W��_��{s ��-"��qQ�=ꓴ����ח�0.�?u�Ye~�M�)V�9�q7%��+"W��H���h};�K��H��t�n�Z���/ؕ��蝥z�z-h�$nX�H ��ޡ#8��^g����o�t���
E�wN�,tթ�5�a��G����F�'�fcoW�Y�jb;��J����D���V�p��z�=R� XlxVHYEB     400     130k7T]eT��l,V��Fa��@�����o���-�  ��L�����,�i�eQ���S�o*H��y������N�胞�3�g�bh�.h��}Y0ܜ��_(87Eo��[�#��WG-5'��γ�n����TB})�V�������o��T�[ӷȐ�V�>җ/\L��M���rCIT����hM�d��͛P�+��8	�b`qO�W)x[���nH�`!|A{V͖�	:��n�\!�� %�)�Om@_ c���N��ǯ�����Utۮ:�\���ǧ��cIcp�NIU����V����XlxVHYEB     400     190����f�&ӝ�*T߆2YJ�A��ӌ*	i�����9����]���mלڤOW�p�hP7�D����Gh3I��x�K��Tt��O�ۿ�ֿc95��|���(�I������2tX�|&&���*��ɏ�|�QCE�;d�\�2IG)���6���A��LG��2`�k�"�4�V	����xf�'�Pt��.E_���&'��C*�1S��I�����Ϧ���i���{cUNw�Z�����хx]�Iy^m����H������6sU��d�|E�Q6t�,Wty�غ�5K�r$���b]��O/������ʚ�Z{3J�z>��O�����`�I�l��L:�u��$^
n��N�'7�1�(�1nԺ�mR��BM�������$�ҎM\'+*XlxVHYEB     400     110�<&��Ş�9c�ºQ����6����y��9�����A�~~@�h�36��_?J+79��ˈ����uAf8�x�7���򳯥����x�������iޢ%gS>Iz>+���v�b	��K)�Nk�>[@y����\�}�ߩ��^\d�w�R�(��97�mz�l`�ETl@Dr�a��:(�;��F`��Q1� �
"h�u��3��wEP��smD��<���G�E:�0��,,�.��e�N?�*�Fof6Y�Æ�h�|�lOb���F�h6�XlxVHYEB     400     1b0��9� jhX��,]�H% ��K��;]�.�Gl�y��48w\���{K��or�n63�xq�P�hJ�+�Iޟ_�q���|�� ��� ;�,nO��2!�?��,��]��f&��X?���a�O+T��{�u�Hjjݰʉ����MF��+�s�>l�V�\�E��)�tdh,��:� ��� ��+����y��&MfeѢ��!���Mªܠ�Ȼ�(��~��Z���o�UU�1ߔ���}�B��s�C`2�<��z+f�WD�Q#�Ú\�� �z�FU��M�p�#3�M����^������R̪���x���6�/��<��3yA�����%!�Q���ˉ�6�j��qh&lV�	�Ɗ��b�λw72�|��6=������7G��1+Σ��Uv��(>��H����tBXٿ��EXlxVHYEB     400     190�W8�P%]�����h�Z 8��= ]�}?�M������w?cE��f׶���'c�a�L.�hjR�&d*8��`���P��'��+�9	�C�P���t���g�T�D��ϭQ�c����R���m�i�L��zYH�5�²�NJ=�<��� lT[DY�J��e���|ތ��]� b��*[1��Gn����B�����u�V醋�.�r�ߋ�ej��$F?ZM�c`���r8��L��/e��[�Okd��y�[����k�J�D�����E>�8R�	X��r~/4��*���40h���HL�Y-��N�@7�ث6�3�vUP��aݝ��^���&'@�QN.t�6аE09�NĐs�L_r�rq�3q�nG��"�D�~��6�r�t���.u��b���5�XlxVHYEB     400     120��?�Q9��x�k8�D��9Er�)Hn-�P�����RHC�Β�&�&-��د��,��;�U�%5�yu	�RWܶqB�d�e��K��o��R���Y-�j4�0��1���L�8�	��,&�!i�H�ӡ-�Q\ޑ����İ58�܌��	P��b��7[�=��2�'��xX)���1>����-*�ӚP�T��u��ϣ��������\���y�+f�Z���5�(�z�p�Mc���~��9���O>K��Ab�KA���MH��C���<z�5�*8XlxVHYEB     400     120b&�uH�N'[����j��7�� �q �B�78�`#�B� 2k6j�e��[�{���r�-@�o�o �a$��"⚴�ʣ�mE`���6��7��0�zV����w�
���B���0m��5*�R�zd��0HEGJ�0�c��;k�9�{�����:��Q�v20�NEE&�AV�[���B��?-��S��=
��?#ڽ�}��}�+2k�t�)�Y�,-+���_�Wa�s6��n�1�ќ���>��D���K�(.��CB��#
K~��Q����&XlxVHYEB     400     160��]����m@3����>o%�a�c�5�n�\�P���� ny\Na�r����OJ&J�w�B��4�����>��	ì2�Y��N�e�-@ZiȢ`����<J�B�x�4E[eJ�&.LB�<n9�Lt{����aܚ��쥶�;���b�b�:�dۅ&�`�<�Cu1��-�G�"z��s�Q�^�0��Yв,�R������]̢���K�=���^�L��5yۅB�s�C�P2P�5��og�&6��ޑ�0���8���\��CQ(�Ӛ?�E`��P�(?�lI�h-��g�z�F"��'�·�����ƚ�׌���|u��&����c���9BU����=LG�!%��HXlxVHYEB     400     150KJ^���sLl�"2FI��"���J��C	\�3!�݇[m�_giq�.,^�H��3<$N�ob	�B��V9����>����n�+������-�����II,�N3Ir2�.��r��;�: ����7*f��?SjU�����Ӕ���T��C�)__��GTi_�(�=�W�_��q4:%��M�������-Z��"lu:�L��dJRA	g�N�mjBbۡj��2��y�ԳcՌqR��2��ʃu���q�²�ҖԪ4յ!|b��[�h�Rd��1c��T|EUsq�ˍL�u&D��/�?L�����	���/
J�WF����zI��LC�#
XlxVHYEB     400      e0'm&�sETi�9�Rѫ�1|��F�Mb�=�ѿ��ʂr�B�����Ŋ������;��Fp���[,�f�g�і�M!=N�XG��)>~/`�r���[�W��&²���%\�͛\�
k3|K���AE���+t"l�T�����U�'ϴ�-�ڜI��r]��*J�2��FD�ӇH�'��?TV��8�X����e�եg�	��	n}�|����~[��_WsX�Y7�XlxVHYEB     400     130���47Q��r��ln��m򜵀=�@�ɬ�ųO+�&,�U��[�D�M(�bq(��lKS5ɟ��ه�
��Ev�2�Xb�a�s�����b��1��h��gϞ!*ز��s{�*G���ɀ��z�uS��5;�a,�S�~�
��R�̇)'j�P3�?3`ns�.�E��Ґ�ͥ�9%t��k��Bi(�C�/�Lx�Al���|���6\��)s5�IV���@�}j,|0�[�Rt+�)xw���]0h���/�o
*i� h�B/9�J"�x�ϫ<�e��Ae6O5��qq~�i��f�*XlxVHYEB     400     140��'�|�-��0����@�JH��cA��{M�Q3���˽`���T���Uo�$ڸ�Op�R~5r�ֿ�:�g�mE^)/*$�&�1O�7V/[�P����B>�V|IGi�â}v.�D�O
��/�{ﰞ�{S�l���^`J�Ⱥ텸.��%�s�x�U��+���a�<��E�Ok�M}�� ߭�v��`�c�P�x����âʔmE�U�T
w^�>B�Z��M
Y ��z���n�Q�&�Ys�j�G���lg˪�,�F�T��p?�<�	�_uC��9���ɓ@�ϬP�t]|��/�6��b�E �Pu��QjXlxVHYEB     400     15003T��}#�������ç;�U
��d5%��P�-�,09�![N�c"@X�j�]�'�HZ��|dP&����6t!�{H����Z��<H��ƾ�����7qB�����$�[�p�啵�6L�Z�-�Le97�U�� Wx�a��td���JX�^�l�W�yr,v? 
�g��R�i`%N.�i�Z~��֙��6�h.{�q#Ú��/��\b��TiA��;�^�	&b�&��kX�3��YI(�2�uy7��_�����'��A��c5�Jq��H�Uf���x�~/w�G��d.����W�on���;]!&��UdV��o+5�Y�XlxVHYEB     400     150I��4e?���E�	e�GsJ��;�E#�������?��E��%�Xu*'��v�SD��]�@ze;�@�OGA�y�u�(�l]�sbx�79;�CF"@\[��(�Jkc�O�`�̨Y&�~*�Α@5J˭�F�!h�<�$���4
���Þ�mI��Pa�y�R�>^��?y��̢��f�N��T��*�`�o���5c�֝@Q�K1����3��:l�"��~�0,R0V*���
/ȳ�Qa�D,��"$��{���!��},���	��|�c�*��RÒ����a��4~�t�ׁ�G���/x9�*���RG�'�jZ�.z��6�{XlxVHYEB     400     120Hj�K_�/�UGΧ�n��s�.�.v>u����:�����o4������5�u�����ڗhB���" �3B���3��t�Zn�n4o����/�WCNk�0uE*z�o�
p��Ë��A|�-�DJ}�̠h�Kf�[a`�X��t"�']�R�Ǉ��
 ��y��,�VB/3�Y}�T��!�\�����g3������<J� �,��V�,0�n�hcr^RG�q��C�ύG�e��$o�*s�§����.���p���/;���u����l��A�6����$�Lt|XlxVHYEB     400     130���D:�Q�w"�K��M�CuΨ�=_���w�9T#�P��(�0
�}
Ţk/"�e.�[46���Gn$�|�#ׇ$P�*���?e�����x/n��!���������3(8l�p�����ϘV���υ��~�`�ъ�*�O1�x
�k����+��XI26�����%��H��KE������WK��~3��N��Q��M�[>�R''��9�B��4��K�0%����j�����/;�P�<���`"���¥K�M��M_�����9�2�c��\k�W���3���:��wz��!+��y���t�zXlxVHYEB     400     140y�g�Q�@�����������,�6�Q�� >�\� �vk0�?0YK9T�;�v��߿��_�ܨ��)}�#/�Tkݔ����$l�m&�Y�J���Rhu��n�-h��h�D�u�S*�;e
C�gg��;�T��ͦ�H#f�R�)M�k��l_��J�^ءk;�d�DsA�^M�Āb4�|ObQ.k�S��n6��7X#�y�~_Y�(V�T4D���y���)KМ{�A�?+�T�D�G���T�F�41�[����ӊSgV@Gu�2�%��G�p��
�5�%!�X�X��n��ݷ/�@�H�7Rf%�3O?�Ԉo������̽� XlxVHYEB     400     120�NԳ)o�W�,�%�0�qy��ݩ��W���y��vw8�z��#�L�˨����EJ��d���� ��W���N��D	��O�k��7��.*�'_�Tc�f�^H%H��w�ղ�Ἵ*������!1��jC�����k`(�<V�k�Р�yP��S�^��&����'~}��O[�#=ٶ�7�>$�0��m�h�F_�j��s�:`�\X|}����Z��8z
�&7�#��� �#��M��u�jKq���m �P�u57ϒl\������v�劶��{x�u��XlxVHYEB     400     150H�Ȟ}{�Cw��PJ�m2".��h����/�����P��,-g1�;?��<���3��Ԕ3�E�>�;���?'���6�q�HF^�+O�[yy�����~�G�d�|��~�y�j/&�[����ǋ�4��N���p�X:vv��D��!����6�;����:�s��Vș�+1bI��~F�ի�Z�&q�+�{�t�q�����Q���{���@�ۺ�x<�+�I}�}lp��� �譙�"��f������)9ʣ��}�m�������$$n�D�||^~�]�[_�&���,8�d��G�.��Ѓ���+���XlxVHYEB     400     150���*�Uq��1���P� �r�P7���7EZ�.bA֦����z�`&�i �\�37?�?�޲J/_$��E8��q��+ߤH�qX� YaoIQ��cs�=\|��qY&�i�ZvN��yW��J���+q�o�7]�0秏��l{�ȑ�ù�/h�r�lK�0��$����,5z1�y������p���f��q]B�F����~�3�@��3���0�6EX�~���g`5u3��g� �R/�G��#l�j�W�ƨ��_�Nr`�h�&X�p�U"{�e2u"h�4�UZ�`��Zy�bҨ����Ϩ�!ז�Vh��g(����-�H�XlxVHYEB     400      c0)��k H�Ҹ�ji
g�u���K�~�÷�f�=��B�zL�Qx5�dɰ�( ��f�.��_�*�Sʈ$�2�fܘJ!��OYk E���Ӟ��:,�</�b�^�U^1��6��@�cϕJ��b�MƙQ	e�|P�^ҹ��5T	N����5��"��
^����2�� �K}b¬XlxVHYEB     400      c0oX['�6�胗/̃�-`rs��F)lL���a� C���{wj*��D���a��xP�33��l��`,Ҩ��%�Tm�50D	�YSq��*�)��������,Vuh��_�F��Z�(��#;����;�l�Wcγ�C=}�c�9Ò�<�/�',�:�0�,+���n˓rh^��	">btZ+Z��*5��s���hXlxVHYEB     400     130=lX�J�35�e�Y��h��P㜇F�&���ת���W����]�(��`��p��==�zP�5F�{�ǫ+��@��`OHKf+�����>W��ti�]���`�S/x2�u����u(7F�B��AF����`�%5�e��(�+\Dƴ6�O8�G��#0W��zM�.�s�]��
��^����)	�9��w� n��Ŗc9?j?��=�� �1��'�6�0�x�l��2�̆���}?=��̙���3��Ʈ35I1�����2����?F�f��F����Q������k����NXlxVHYEB     400     120��+�p�7����$��#���3ܲ��_�E7#��	�Ei]�14�Ă1#�1*5�G?^VU����ؒ��a���ŵgRy�v�fL=غа�3�q[x��	�P��U�)qH��z?���������k����Zw���:�-4���[�5%L+gWG��:�;a��^�Hw/{r�y�&j��y�v���&еx�kW�3k�Pv�3��T5+��/G�O�˒��+�T� W�h7ڭ̴K�g�B�����\�M�Ʃ
jb�n��b��T��۽I�Pk$����	���|�h�/XlxVHYEB     400     100\�i�p�\`u3��n�p`)�{��ʶ�n�0���J����F:�,�ET'�q�{*�!F�dB��̀�{j�kإ3�-�d�}� ;���^v�A��D���g8�4tG��=hA���~����H���A?H��z'2��E�z$[䃂��Jڅ%�/�R�^7h�0$��K�J�CM�M����.�s�7��P���9�ݺ���&�Y����{��w�ht5����F@[当��e��w/E|���C;����XlxVHYEB     400     160���V'E@M�f~��+�����e۔�KG5e�똽��Tu�;9/̣L�ɼȴ��|����vsD�[���:�U�����#3җ6*��7x$j�5:�ӵt�o�)[8�ϫ�)ƆGB$���⿄��nY�zݺ��A_�.���N�إ�R����$��$�*)DBiG.
N��9��0�|�x���1�?_1�F{��X;h�y�gO(+�2�� p�����r�����y�	�)`[�� ����@���"����(�K�2-o�9,!�����Ͻ=p��Y�D� ��(�Y��
F�'?#ĥ�R�FW(�Ur(���D�$�^/>U�����O��'��X��]��}XlxVHYEB     400     1c07���{�qT���U��2�"��-��(z\�|4?�}s�Dt\�'z�����bXoo�&:U�K{ӗ�&����o��X���o��ۚ�a�w{�ul2{�G�����%[�A5g�:6浬��w�M��n3^��Gk���,)cvh�y�xM��S�?�T$~U"�Fp�T�8_��#
�� t_q����ncS�
�A�����Fr�[Z��(ĺ�+��T�i���{V�q,X@!8ߑ;<>�b	Z��I2���GH*�fzݖ���(e7�]�-?����68'6R��`n��Ce��%��t\H�<*��~��[�>d8o��h�ko�.��k�Hh���{h���b�fBd�@�#˲�C�ˠF�}B�`�a����2��ttt���>t^5�=��GQOM��$57�{Ub[�DH�+=k�ե��,K�O͚�)��4�_����x����3oxXlxVHYEB     400     1d0bC�ٞQ�E��h ��lm'u/�q5�磡Y-ԏm�q����b��
'bp| (	K��]�3g!��qo�'�4+ A����f�.t��	��K֛{k��W5��Vx\���z�U]�.�}���D�d��0��ռ��ս�Wif'�%DPO��=�׽�+[��F�5G�d��0�X�#�V9��
�$�������ȔG:��N2�;�K�|�*vʇM��S8<�^����\��'���ͼ��q�'�F���ht��<��P�!z'��-�4�	�`��+��ި�4����T{��I`��ي�J�Ҟ�9$�g�bU8h��=�����i%Nْֆ�(�<v���i��	�!YL�����`0[���&����J]�ť]�ROJF�@e�
�@\�w�Ɇ�<�Hv�	v֊��}���ߗ`��M�lo ��ڏ�+M}ڶ�zW%��4e��Q�XlxVHYEB     400     1b0��vOh�|�ۋ/ �"q�Fin���xS�
�A}%Dp�g'�Aߦ'��H2C�K�%Kӣ���:\�ҭ8+KA�4�ufvZ<�sT���V^��	��h��������8H�[d�όh���\A�����8�{	(%,\�&@DGG��N���}��Z��}�+B�Hz����X�(()J ?Z�%a����o�2�I[�.�ַ!93b${ �*-�	Z�pڒ�V�]X����\���'Q�i�~�)���c�_���j�Gt~D�g	�q_�7�U|��WDZ:�
��ע�Ԓx�?�F܃����&��w̯֜���g�sK����*���	1{ހC|B�
cS�Q����t��4]��4��f�K������Ww�PQ2*V�}N���%Y��1��/�qF��Gn�	qx�_�e�+M�dcG-XlxVHYEB     400     1a0,_�F*�-��L�R/&2Z�5r,����v��6�G��$R����i�!�N�4w�If���qdV:�!��jlY~{a�Z(Z�|����H�n��a+�Q���u��P��4�/�'�S�_�'���w �F-�C)h�!{��<f��%��W.^o�ߟ~�x�.R�a���7��
E�{�x�d(�2e����F�>U�7�t�@{���Uպl����k��p�	��í��&c�s���:��%� ,�v�K
#�����p$_��2��uS�6v�ęd�#�G�9%��G��z�}�&�n��i���|��_5ܤ87�@��RuX���?Ų�'� Ŭ��Cu�YU8L�TA����ޜ�]�*nYtİ�3[<����j��m�q��w�6;g|���`X��6�Ν���zNh)EO��s�e�$mc��
�XlxVHYEB     400     160\�,��@Tb+�F/�x(�:�����%oݝ��?ͧ�N�?{��Hb0���Q{qɞ�谲&n1�c�3�߈��K����r�'�F�1���OGh*ll���7�Y�R/q]~�K�V�����)����.�]��S�c���<�[./���d�`�e��CUN�:�'��1cA������չ��39�����h&6h؊zpA��[����s�!��]o��E��潵������U��E��^�\"�|(�tL�+��W]@"x�1E�*]��t�2���pSm4�yt�U��C�[��/G���Y>|/M4���P� *!"�q:�L�B��]LrbFm&�C4�~� W�XlxVHYEB     400     160 W��
�W���8mЕ8�̒m��p�}�C��C]�|Ik��Z�U��4���o���8�}I�J	o��A���k.�DD���������|ή$~�p���8}\��ȞnEv�R�t��L��ni�UѻF�/�= �u|��fX`)"�Q�bV�$d��C���cJ3�q��,��z�m-:_�c��&���x��A:�ic�V�"_M�mež�6����Bo�)}��
1�������%�D+KEǓk,R�n��;s�#�g�rށ�ɗ�"�Ժ	�n�u"�}]����Æ�-7Ŗt�V�	�s(�L��Ô|L4�~>�r:h�k)��0^�E�I�ý��b�RV�w�)XlxVHYEB     400     180�%ȭk�F��=����XA<;y�޵��2�Px���Z��x+q���?5�h��eM&�]	n'��5p"
�k捾h�I���}��U`�L��=�w���A��U���VXy��v��X�+�4;e�-�����*`+}dP�u�@����t�>�V� 㜧��9�0�s<���(wWtǍ�4�,f0.�|�˙NF\L���c/�g��d+N���Ve�	]�x�s�N@���v���8qj ^AGf�|\h���� HW��8E��a������^���*����(�g�#nu(~{&1R�׼s��V猫 �+Ky+�EK�D̰�q��C³�����'�^��/O"m��Ԏ�IǍSQn�Wr����&|��O����Fm\A���XlxVHYEB     2ed     130�G�I��oy���C8؝�.�`�]%[̗������9�+'�	�o����}K1�T���n%���yɫ	��ݡ+n��*5��_|j�p\�}�V���S�v���4��lV:H�#|z�%	�/T0mP�	F&F|�R�=�M.r����Q+NWb�5e�$%d�j���N��by�0��?3H�
��s���5	��A)ڭV?ρ���w~�p9w#a�3)���l�cFH�dkb���l�>_�,�x�ʾwJ�\�2b���U���~�p,\�;˃�ȥ>��z��L-��4~f���ϊb~y�\�