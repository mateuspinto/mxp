XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$H�WA���쁾,*�QX�͆4��E��zR��P>R:����&���|?��όu#��7&B��5��l�j�CN�r����n���|C|t�=r�f|@�-��h0��:�V:W��D�sR�M�W�h������k �ѥo�#��X�5rNV�/���9H�F��a�rݸ��u��ކ*�i��EՑQ�%=&�35l�J�@L��U�P*��p��A�s�nz5rGS��XG�Z��e@$�����פ������}��rL/����O������.�����t�f���5䶤�/�C+��.	eTs���~g��9$����"��q[-y���)�
�0SNU��F�t�Y0�����ذH������Xfm�ŀgY�(DlXkʱ���5���dF�q��xjHNT�s�|�u��*\=`��x��[��5��Ayz���c���5)��"��:���ߏ�8H��Gn'R��L���%��q�7j�(�����#�~�PZe�㽿�Y��}RU�9�?M�� )I��0[B ��~
��Q�-U�X�a�B4F:�`e��GĂ�$|���QY�P:
.�@i�^/�13D�K���8����cPKlhE.�f;�[�D%�~��{��W�l���~d�rq�v�n3]R����q�ϝ�E6��6�!��NR皠�e����E}�F%SR�\�H����'�/�5Z����勳�Ď��y���8���⨽c�ʘ1rC�E�ǣ�#�D<�?Mŷ�s�����UXlxVHYEB     400     1a0έ �!euCg��]�:���+�R�H��)ѕ���N�AK�����mD��i�u�R&zBm*i2[�H^���k���()���g���Q_���O����(S��?�M�����A"Gۣs"QB%,n��V=6�̬:syK��+X�HI0j�I�at;��6�Z�@�J?�[ �$�b�X���wY�@z�|� %��Ku�`+�ؐ���6� J� ���4��d�y.>Q�/@,�����/e�� z2JE�<�ښj���������a ^�1Q�#)��N�i�X����vLx�b �;�������7�K����~����S���C'�+��O�h��rڀ�����.?� �O�B��?��0�'4si���P
����2�3����!�ш��U�����wm]m�T�\AW�8XlxVHYEB     400     1b0;��7�986���[��&�:���;�O2��G��sӲ��ؕ�R?S6�hm��+B��mQ�B+��k�p���~��'H_�'�g�q�tS��8o�ݪ]ff�������ETwwR�`�5Dt
u �����l&V'��'2�p�z����q�}�1F�����:.�NR���L3�,�`w��h��	�8�ب����|W�^1Г#!�~�	�Ѷa�����V��1��(�ȻlT����jtag>���d��\w���!������s�	������Z>OͧH8�OK�q�	�cІ2�!����F��||��	�2���$GF(AU��ٮ�����kb<n����Gy�Nb�!���җ�q��AtK%ʑ��ii��(�_��N^n�t��*Eٳc}������t�\�a��&?�K݊����OXlxVHYEB     3f6     130ڈ��֦��<��xP�v����P��,eܠ3��l��e�Kw�;GU��䥓,<��%R<~F���3���N*y����rms�Z�N2ݥ�Ѳ ����v5���^a6�/Z��Z�-2~X�pѥ>(�ߧ����_����	d0�tP(���(���r"��=M��cD���jO����l��
k5��ҕ�x �v��47��c�̣H�� |l;�9XV�7�l��|=~.��"��8����ZJ�Kw���g��L�D�����X���&�41X�u1���5�Q�h"o�W�CR�Z�G���