XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@k���.f��v�R��������p׍0���m�H�Z��[�~�<S�U�jR�)�B(�F�My����Bl^�ٸ�=��j�M�uñ����_մ�5��v��f���ɹ�����o�[�w6���d����/��(}��E�d��o`F�.��ҧo�3/��P�L�F�ƅ�x�M\H_���k`⨡T������n�`�^6��8P"O��v�|)n���i#(�"�F!�τ��a$ݖ��
c�!��V���Dk)��
�8E�薵;@�D?�h	=����RD�L}��k�g�����y[��_�^||�[x��R��p�FL�|�����B����x�Ńu^	����B�T����i2z�(��t|q���,&�=e�(�j���G:W�\N��]w^��E�Vt�\�0[���؅-���e9�Q#Nr�\Y���A�� ��O�z�����T~�*U���Ǐ��//ð$�A�'K�[4� ��,ɑf�Oζ��Ot���⫔8�Z�n/ٷJk��p �~�&�n��nWᔪu������m�.痺_�^oZm�ͫ��:S�� VɎ=��xdN�Ԗ��>�a�¾,n͜�%C+G����V
�CRE����)�К35:t��6�Y4��P���*T�^޵�=t�i���bR-�Ta�"�ԥ׻͉� ���:��K��+�eg����r�'���R�Α�q��}�rj$���n-Q�x��:��������X]�h�I��̥i�.��Xy�XlxVHYEB     400     190��i=|\�8,M���a��|q�L���e��N�2�������t�Aی[�K�*�
`��aau��0�������8��%��~-�9@}oG7�Y��c�UOL��=~E%9юO�pq���+H���.��rm\?d+�a\����? 	�׸�<�x}G���D�{�~��Y�&֕���LY�"��B����ȢN͢X>d��%�M��:c�.T��HY���k�P5�?�@ 36�����R��H
�-X%l�h9��`cQ�5'A�_�{U{yz�����ͧ���z�)������@0�jj^?]:������ZK���U��}R�[�b=�h�y�;L|��0a�S��h�{��<~�g�D��hl�ؓ%-��s;P �R�Lm-���s�ɿXlxVHYEB     400     150ȝ�Vܔ��l��R�D,@�j�cIS�9܈c&S��z#����@�p��Љ���A���
������_\92�4M���K�FI�L����އ�q!-�>�9��O+��;�.M�k�ΰ��fN��H�IEd��~�ɯ��Х��Bg1?��o�/q/x�
sW�9BM�0G�?�C; ȇ�]΁�����/?�Y�����mo�f���^wU-<#� �,c���C��!K�]�-��73�c�1n!�R�=�`�y��[K�nl'볾<o4�ݨ���6j�a��cVO�` ���I��$�?j�gL=G�j����^WǓ�r�V4a��t��XlxVHYEB     400     140og�P�l����V�!∣I�, �W�����{��%�))�c�:��g�s�/�h>Zi,J��M�}�k� �}�+18���d��XQ�Y��]�_և��E=F�1�Y�P��4�����U����Dܐt��8�*�j������"��� �R����A�t3�X{9�M��t84.������`*��T�$u�X{��]�M��ȷǏXD��`���חЎ��p�e�8s���	;Y Vg˟ZY
����_��=J�("+/����-�;]a�y��5�|���L�ϻp����Ua�MwV>��|P�QXlxVHYEB     400     180�(���:U�>D6���1��P1��v�cWPD���o������"]�%vE� ,��u�d+[	��E��t:����t�2uOG'I_d��Slƶ����7o�\7<[�4�vdN
������@Nn��W�>�US���r1t��YrԬ�{����=k3�l�4��T�0dX� 9C���G^J�ێA�J�F�`@eZ�D��'��$����WS d���a�󑆸�p�LS&S�=�(�/�)�X^�f��h�~+4���ǌ`͙�\k~Ӂk��!�XG�v����V�#
t}�ޏ��<��@uә�,"�Z�H�^��3q����*D�҉�޼���n��Au~@�`�����ۍ�ޜN\�{�֩���'x�S���|0��+G��mXlxVHYEB     400      f0؋����%G��}v�X�g�<t�W,�B����gK/["�:��y��_�?�3�p���z@�{F��O���=��;��V��\�{F�G�lق.���;�ޛ[yBjP��&fWcq����F�-S_���lt^��=2�<�Դ@�6�\�Х�4���=��$&�t�,i�2�V6�����F�#��d*
`v��@]��e_c�H����9��K*������v�Օ���XlxVHYEB     400     150�al[��6A��ӥU&%��Z��Y����3*o�ɯ9A�����F"cibOq��G��X�>�DL��W�i��n����W'�C��ɾ����R�����OT�Q���u�g0���鷕���z�����Y��A�O�{�ҷGP~u�-����9�=0$��5�O�5���1��M+��[��TӚ/p�����P��RU�һ���k��厬�	�]-D��]	�v7��K�� Z�r#��b���ć-���"���+���9����DYDdѪ)d����۫]XC�9(F�V	,A���R|�ɛ=�L�cxJ�ɻN����XlxVHYEB     400     150�Y��Vь�����~B��kP�Pv'��@���p�7/�zĐ�[>��;,s>Ӆ)���m�b4��z�����2�~	�Xz���:�1nq����F��|P���2�jLK��ܜMH�n1}�y�����,�L�M��Y�%{��` ѷi�����١`����f&��=υ�z�����m!ak�`h%SD(	)d�|�����ӹ��/�G�C5�,O�I�~'v_("3o��7�~)&SK��F�'J�Қ���+�&�$"��a+Z�:y�ǿS���?���b�2�E�5\�=���0G��e�e.�˩�<�|v��#��XlxVHYEB     400      e0� OϕN�6��[�Ⳛ���)�+�h�����{  R2m	3��1�J"�ޥ� Fx546>��RR���V�9#m�*Y�E��)�bҰfE�ʛ!Ē�#�K�p�)���lZ'h0O%ڀ+�h-E{1�d2�HC>Ec=��;i��2��hޤ���&Կk��^�CD��E~�˫�XJ��5�Q��5h	��镉��}K@��Kw���f,�E�i�S��:���R~�XlxVHYEB     400     180R3c'�Y�GF�l���S�}Ȯu_s�>���,�b�i�D�sO�{���4�8�����'���$۔�^��=zr)��%˘u��A�{�3�P��vF�iR�c�݉}�֚��J�)�������^7��)!T]�6�L��{O0����$qG�?�uF���
7:j���j��x`y��A~�> K�5��&Ķ���0F������d���^\7M�,��s�<k�Y+l���,;Z�@8�����W�|d�^��.�rq���K�ߟ�M:Ż@��D���z!�sr���^�:������Ё����ߋ9~�e��8�ϳ��M�+��?%��ja�8R�d��ft��7\O��e��+��K%Q�ptl7/yQ猣D���9�XlxVHYEB     2f4     100XT������c�4MjtH2�e/�� ��A-w���E\_c�9��"������]i��r��rPXݳ(:J��e�o���K
��/<r��NwL�p��Q8`�T�2��J�p�Y'�G?"�6iwRކ7�d��6�(��G�
vʰ��H��L&�^�1���&�]�R��]�\D�yg��֡]E���%+\-o�FX�A�Aь�˭E��zx�wSx�� /�f�kE�O2�)-(��������#�)qtm]y