`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
lqzed8lF/Gsywb5VIuusjccBiy5rXQYyDxvRKdqr3KOg9FVsFNXG0tCTKEPHzcwVx4qSVzlgJ6bp
rXToGGzTtfLPu6GsvPMGzQQl30I3PrORX/YXyBK2Xeh5QsAMprmequXOxbQau0gBriwqlpz4Iwk7
y+RVO/UMv7+DdhLpyzwMS1hZUVg4EQHEHStve69YjkEHjWcKJpPtZtGabJuf/GQXRu4DV5i9KX6l
E6QXy6tv6F+vGw/YaSdxDDxfnUEBL1MRX74IsvbvF61dfavgjTyheyrR6vjj3vuWiraB9lN+VOSS
aBqBZm3/zu5d7BSyWDZEGvXfWI0cem3NrDUj9A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Sgp1z38zqo6kO3vqDKA9e3VetaH3za1K6lQdszz8+c4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2960)
`protect data_block
53vJAPxo4orlmqQtVCX6TfVpJsL07GHKxtVesWexF2s/AAvps8OwPrMzJztY5Dmekw7FO73S9fJU
WkXbis2sk8jXXX7cMXykYUp5PiN7sGw9Wro6tnwPqpBKxOe/CR7chzyHoX20N5lpwq89Coi7OfGj
47Ae0e6Ke98MaDBl3d7g5wHjs63566+LRNWl7X2EgfQVDePR95cZ+9ssvsqULi0gknw2XvkhVTiT
Em5YgvWL1Irhjg6AWsgiCGPelsihDkP/777vbojA7cIfsxJK/mGluy7VZCk+zwfJ8R8G41mAVyq5
g8gmWGLuhheBXqEp3FERIWalm41WVsHgD3nQUmVJV2bpYso+ZBwAIded5Uxy9iZv3uJ6z9wKi7l+
uF4iipwCJGp9Du7Wnbp7KksHhRAEqvar5BxQAcH6sOiLy23y/omBlqqqS271W7TRwVnd/UAzOj2Q
Bo5L9B3V9ZZhY1yS5oNQZtMHGEchmX41/qUPFiNJ7ellJ0i7MnFIEHusZDVluMZ9MhEdRlHT/XNz
4F/Tpui8im0OfzCxmetWusdOm2oF9mnw18y706mDaArisLn/Q3YecDesWKWLpDoc9UL8+7P6YtJ8
zI5slWtCQlF2AeLH30TrEfaiGgS75FLWmm8ldKLOnwJCYWNmadIkwXZ3dp5cdbmfsIkcmfmX9Qd1
IlkukqixFEJhgZ45g04KbYgWp0Zjw9NjqVGrmTFtNffwoERar1WH/CgkgxDECI48hSNyprHiNqKI
DWG55Tl9lsz2DGwnZn/LRULTbnevSLRphCEYlReARU8CNI9VYBQ3oTPNxxsizc4NYqZoSC3m+5iF
K3bnrC9BcyjTl1KmLDd8cHqPhRXSrgIMW4NYBKMTBaOp2NzuPpDeyYZtIiUe4r74RgRvl5p2cxkB
ijJlkSaMSls+VH4q0yY2l5Hrxe2Sdbb0i5M8+Oslp5alvpVyjOmUP5PCTyX3KFepHdn35zVozZJM
hQRzCC3mpwlQtTOxt9wubGCVA9I6RRSz4sKgDuk5pjjQ+fJcvkiHfTZBU2tJdUAkFFuDi2slk3dq
jFMAqtkhlXMNJxzN97SZUIvPExFnqFyrisnKyzu0N803T1BmAvN8PqdYwU+o0mdf2/rLbqWulf6F
vu5ettd1DyqBzXJW8N15D2y92nP9hMaaYfOqzphQHCYt0ghwAKNfxCz2rdJ8+vTsEtQnavPq9ZMk
GPgUHJddemRCU470niSQ/yU7bV3gLkBY+oJm6Ebv73s0dats4TF7GQycBjEb52R/Z0etwf8g/Z+l
fH75Et64pJwiYF+4T5/AQYbdQoF9EAvuwyYuOg+ZyDiFAsq7KNZwdHcTUs3XPKbmgqyFaPpaW36S
lw1xSFPOKJK91mspktlS+cCp35J8vrD+wtTmtDuk37F0jHyBpkwG/QWA+TXSPEF+5+3QEIkNdwfB
/nGel/XWIEm9Ats2LvbUYB5BcQbPxOkqQ5PxRicMCsxTN0Vef95Tp4g+mfxdAXuMKAiiFOChoTU+
ToB+qN9FLBEnK912PfwuzDk0zyHJp+9r0O0TXDBAwriAZ6qsdFUwz+sjWTkAWiuhieoQ7wIO+YjL
YsI75wjoUsYVHLJa5Rru68XZ/rHWCmKwEOshCXSDEIdSWRzc3K6aKNqnVYDNgD2VGhFUBjpg0Ldw
tlDkTHnx5VSyemeGp4v8wO2qexn2OjobGZqpg6k/eDyZ1lcziZ40MZeYWyoRKvP/SeD3Txuxc7/u
YT9Jz5YayAWhYXDoFlsPqzfpQnasQ+EPbahV+XIjpCvANNYbsZN/uoFKlRP6AwV3W2jexjXCUsFF
bxlJU9Ni9G9msVCoMVM+i+Y/NlGfymx2FzdbiHeMvV8O4hnjdgA/yvSTLdmaGJHY9YzDFa2kXol3
rwNv2BCE01EWMV73iR608J6nK38zStQ14YdMWRW22Vd5AFPmUA4/0eFCAxpybD8uDZ/SdAvdHlnS
Jrpaz2RyFl2qPIo7VbCWY/TB7epK+AiVM6SGN4NB/untdO+axWmKVj2My3cXaBKzh8HtTC99RIVo
6+WHmWGbw+M9S3kKDa5PGd2BSDsYNwUxVLUZPy4HsoqL9g6QDyK+pJJdYCflpqtbGZ6pVJpRHcgQ
GZqhj4eVIWB8LdonCsPFFGHmCcR3pifQ3YtVs9vmFliw0yZueeUapGNiEmYg9/o3A6iGIidCUN7a
j7fmcGmT1zJitkmqbtcJCI8pV30F3J22oKH5KPa+I2k0QexEqqsSvxL+tQkfblycblCVBaUqJ8iY
Bs0zGxgfsk58sGneScs8qDAQ1py1HDo2cS+U/b0S5GZ5lQJhFp7Os9tREUbVTscfh66KaN4LFe6k
hmaG7TUE5is1P7v+RPDbC+V9YqKBNoGbxFkfLUovd5iY1my317K/Cwpuf48M7pXt+jnkp4G021bt
klerqAYKluG3K+8NjkPMADhdp9Oj31aD8LoZOK//QBYbVFOjFG2DoaGE05aRW1XyCai8Yf2CTKb/
SLwM16W1qLMsfDIMZ+ZcI0dfGkp3vFSeWYQBGocEFLJt3YwZ5ffWBYDclDN4UkOO9r+XzcCHfIIJ
FMXkPEd/fl24Ez59Ket9RYxUD11NzGmZaoLE0EKNzO7MUMIatlPZYfCCiuBG4if1H8fCnVrBXGJ1
9Hk2lVrNZPuVRz1rlZh4m5r7FJpJnvaXr3PuBH7pym7IJAZjjkOfU2vrz3RidoMcXNe3xLqSFmOW
u/A5xETXZhkwV5AubfuoAYAmaW+AqbJ7xdTf7sJHrzRlM1QzeKyoKODFcjtd0jEax+a0id/t/MWQ
LhJ50JLep2mjnuh47uJ1+hND7s1YtyKBvVrl7zjSaCRbB7W/Z5M9gOVOMmpeTM3nsAnkBZlkNFfk
46aoJgp65qZGSEYp51wx+bU1am8a+83FtK/upwGLl8cyq8oRI++oLN8UU/RAfWPdMjYqgPx9rieb
BeovC6ScwBXejZWutZ1y8Oph2dO0fQH2+mAiK2Qcn1x+zOEgrKFxNHAd2hnutQA7sqxuG4jRg4zU
aVlzqrpaQJlcrLfQOsZHR+Tj9kTWfv05u0OgD/LFnKCD2p/Lrpx7puGuiD2CukNQDCwOtU7PjK9b
MzAl5B78hKsR9fRzChbWD5rlt0+yTZz9jp1SvOXHXkzfau/NYDAJBwKQ+h8DuB0+Clz11+J+EJVe
YCPuz5NTHkTd1C6RqA2EOcScQUDUjEplYCn0R9dRJf+JkWjK4hze3TEUgdwAFacuQwPrNjswCOiv
dDl78zeQ5hdPxGUmfwQ3HlWPNUkfvYsgdRWUnkYP+bvd2kC1S3DuSSVFghSfvVpz8Yy/FOCWJr8R
yD1XhfB3gSPs0YiWL0Zndu4iAssXgqUhh0Hxm/LpUf59U2MpDtEGNbtUPE9/VGw487Tj9O2UHZKP
rHN6QcuQnrPW/8ZPE63gnuMTp6qZDruHgV5ZH8JP1QXpqSOVMg3KtA1lh0gGlmd7mnUxJBMWlHGw
RKAQ+QqmzMMMxeWdt5GJaBTGrBd+m5K3GbBtBGQ1XgHmzXP/JszKYbgws12nN0YdT/U4k4xd5oXK
JfUNAzFV9xC7zYRojPxfvX91Y3WeqiS3/qKYoWw+vwmU9Wat44FhTEZDIzpeJCwPsnrXCsrJ+X32
6YYqtPpZ64gqiGKds1EaTjTo2lr67GnORHrJVQa38+cJDz1v8jx2clfjVmdr2xFGTKArZiF6+dR4
qYBIvR5eOnfJnV5vEqb5/2f9KOsbiaY5FSY+Mb4e/A+piGd2IugC6fMgKpbTTN3TxKcMoFOzzGN1
pqvnvhlMH7xBn6Z7ivVism7GXNZ1ZB3044+SizR/UmwmOsyDMEV66ZUdmqf6NOs85tlULIuuBGjR
jqHgAFOlZoxsDqiTl4s7aaiSNRzfgjrXgLVaehwY8BPySy4f8QWzgCG4lxvGE9SxT/Evd6Q=
`protect end_protected
