XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#xa�����������R�I^�i�*��j��e����}��R�K۟)�jH=����
��q�U�"{���%y�Yl�Tܷi@g�;4��r���'2�P�䳁U�S6����el�q��}��K�.}�&�Lu��Y\��h�5f0'�#�����ǃ�%x]��g[#ײ�����n"lcH����5;W�=������t��}�LS��u�A�mЅ�:N���ç��Õ�f�A��.��Z��O�Ɂ����t�z�ôlZF�b|���w����0��gr�0���L���͔��}
�r٣�`���#�u���$|�W�^�/�i\��i���C	{�W��	��Eŀ���\�␝��GҠ�b�3��v��D`|������o����$ƛ$��S�}�&���]rF��<p~U#xv�H۫�<��k�W\|�5���6�;xۭۉAG͠jǳF�1엜o��
�A!�(���!�L/)�R��Hґ�t���z��ں��̓�Ȧ�͡��*�1](�弥���N�����k �"Nk�:�LhtS3K�]�?�gA�v�[�l����Bn��2�����i����8ƶO*�7!N.k8���&��\�Nv�����tc�ڻ�7:�0D��D_���oU��n�y�������l��ĩ�q�\�2!��<l=h���M\�V���F���K�5As@-��%�H��h���Q�rh��ߤez ��>�m��z*3����#U�p<=�v��,�f��� 9o��У�fXlxVHYEB     400     1b0�Гaɶцҏ��4�ܰ����EO�A��/:�8�񙊋|��V@�)=�
��{�E�y�Ր1ᆊ�5w��fDHL2�*����[!�ȣ�8�%�'����~FS@Ǿ����+�J�:��RR�=�	�[�h-\-�cs���Q/��K�ʞT����׊��1x��:��K$��2��G�d!T{��o2~A��J�p'%z0���p.N4��=fk}^]��W�/I�]���H�z�<~Ǐ^0���6�b�e��0��G���0a�cb����຿�|:#����p<��aB�ޣ*D5f�qk���f��U�Mr�Q8|����JVG���� �Xic��A��n�p�^V��䞒�P�?��֟�Y�M���:�k����������־��	��!ܫ����V����;sE��<Hyv`p>N���t56XlxVHYEB     400     170)B�i�����;� ���� �~��4�!-9=�Nۥ�^SjCg�0����c��`���
a�������od�+�G�NHI�j��۠�jOb}�0<]��ť�q��4�M�T��J�S��yl�$4�mV�������;���Jhl9p�fJ$�8S�s���.!k>�%p&�-Ȥ�Ѫ, �w��#�M_E�O�O0U͹�h.ji�V&����/��� �j���|�qq"� �zX�I[Ս�o����xs�x�۲����ٮЬy���Uc ��#'vJ,XvWK�G�.W��	+7b�C<�#g�rY9���n���eo,H��L�[�ۑ��+���i�AP�Mm�s"�w�9��j^��z�p���<XlxVHYEB     17b      f0W$�&̽E�dɻ�|k<�DE~g8u����Կt�V��jo �M��d��]�n�N�Y�%���&���*��������H/�'?>:�ے��ǽbN %B�)br6x���J�Ա9�u?�\J�ί����5� �dlZؕ�>F�9�� �L%� ���֮�,+�3���<���˫iiU̩�k�z5�eC��@#�m"��YA׿��	)}̀/ꊇ4����(1�o!q*�}��C�L�