`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
LIDqRdDZDvuWQrM3/ZsixhSHsnGb8TPqTSS70Wmxc9egfBCHY3vBuSa0in99izilbpZ3d4y+wuiC
9p/0OgT+F8kaO263esfuOcv0ynrzkRBmprmeJJgW3aMKOHsIUiKyK/HhYMC7UGAw4/ShNxBMhP2F
zThd6smxz9cDmM7ML9BwnHbH4CmEM50Jf1cTisYfUDMpurMQQu1xC1/Rx1D25SaaL6UuaXlhVOkQ
Zi8ox5vE2uTlANgKPrga+iRg9fiLz9zu+8Gc4AAzdbGGUjfTnZPJYdx21Alloi4AY+Kv19wBW4lp
eTZKUgPj1ET4FoCmMQYFjalUvy9z+bYY+xoQ4Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="C4fkhtH+V6uYtTS/wSPvbHoN9+xMPupaxAurK8tmux0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11952)
`protect data_block
SNJuecNSGniyc8urIlayy6iYn/ODn1cNhp+I8uLIkb3XaQfz3zr8EWq40w5pyTHJF2oV5bFGhr60
/vlBy3Y925agjETKH5wzzZz//YVp457ZGQmWlJZ/qIpDrU7e80af1MyhPA+eKqTQd1FOvlCM8Zg3
OBpZOY25/gxt8ee16u/h1wV5c6RnZAuIRcgOpG4iqplz99edGucxdLOdP+mmAmRTqBJfYTQ1AKX4
bdeoNqNuDO3kADiGEeDWLs46SXGrCzqVsd6VRKXTowf0jo1qVOYyhUr6C3vAEtj4mo5/TbntP5s7
sSgIoLFYbncRpjdenI1mFb2H7JPHOTagoBFtDIOrilvM+D2OcrG/d8At/Gg0qxRuy7c7z/Fh+Wzp
18sA4F492scAUgi7GrKPm0ZFSj5FbqsSE0oiTnCBSvykGAUbQgxqJwn/CFEsulgaAOuHRZWItBa7
y6rsZ1Q21N8/HCB4j13LM13/G/td5OcPfddFkZf4Ct3sKNtGBXwD+ipBhaccVnl6EI0K4rZOIxQa
xK8yWiUaFKf5nqerZpnRJmSfdezW1b3rW+okjf/FlpZF1k0ZWWsghx+ncpF1Xp5/GastLMjUH90O
oOZS5wrxVYjG9oY+nT1V1aLBX4W20mOnMHcYU5qTIaolZTRjrdaRdVjp7xZbNOzm6w13Mxu9HG82
Jxt0Gog1sjnM5KVRCmPB4BXz94O08WZduH9O/mf9Dw3xy/b5LSh+U2xt60Kov1UK1a4Sf8BVgq0E
2jP63mtf4rk6nJUpQqv6r9h6sYxBhU+GUxfupZlxDdKQaZseEoUfVoR6eWUXDomeLrcmloga1rhK
MMIW6pBdfBlseqZu8JJ0KCU1yAYr8dzVRBFBGJSksJ5/DfghJSSP8+VIyaoVFqaoh3wyShODcos2
Zr6t19FJLVJNj+jC8qfQMiVCr5FKPkHb3fSd61d0GJxCwlxjrdyvAP0n1ddJ07jQWHWIzyzj3nFT
7Q4aLdj2H4aw6KZQIWnckqHxRILJBmWXkHay2CbOD+GWDp38jhFTjawbt6WZH+6FiqkI+pzAAcsu
ozAGXD5yUg0q/JzPIg5+F0V0VIS9OPqG0g8vH/1dKqW76dOM2ASDkadcAEjAze9kIRPG5zwxmkFe
9HIK9Ez+j9RatRjahROYA0AqlFoTTEHvQiHyDtEm6e2PB6oSotvGtIAioKGpwgXKZyimJ3EurWCX
y6ojkEBPrGU4i+wqQbhzRqtsElc0NA6f2b7kqRG3GaJ1PLBaYuVc90lwBqPUHtTIFGA8jDRRWKYA
WXfqHly5BvMIq410gwxoHCG6VsDLmT03EBHFytZrSNCMvKchBoukq5XfANjLcbNCp3qmCjMDL5St
yBXKRLav3CAx0LEBMLPFiv1N7t6UZhJwJ1pI889yDmOnsqHRR39i6vQ3qeNJqtRWXKGq3nKJ/2yd
LgpCm3CFNMMIuZ3+ko1pQabbij2F3WVfMBGblY8vK+92RW2DC9JfpCIJYCvUqhCwfaArWgN/aaxo
5b1a25LV0bQTvRVK4dZ1Qms+U1IHNFxwC8/L4Sbu2nKp04FQJBzIp3nRJASgLew4Vwn3o0/NOWCE
GLRRCeiTeQarW0Nm5S/GpPMjNd97D41urb9QqOVzZn/PWGiZWCELT5UB+OEnqzOo2TAjZm62oYie
g/PBpNPA9Jku5RR0wcMHEGXw+jI6fTW/bVv0EZMA0A0rtrAdXvG6ZNl4k4LfQ2PeLXeeMZyK6euI
iUAwvhcPk79kjbRXAqs3zXmbedDrGQ1HVzunPQ9WXC0kVB7R2pS90+HVhmrmwdknci+svbOmlf9s
Lpu8exLVv5beRTcmfvcbkewpJYQ+p79hxKoNO9PQPzm3VI5Zah5+eBIGkyM9aNHaIUxoIr16zN3s
HNsJ5C+8dvYszSIHyfVpb77AivWz8AXDGzdUIlpFLLQ3evdw6e1jiSMOeQKt6iw+5OyPhHk+ci3G
outO56c3MOEoqfYq6y3BLYrvjbAkIQfQFZtD4DcTMaCnSpi0KnyW7+mxxUbap4fRQ5AknEfGsnJD
+1mkNevliZN8zTWRJZnaLpoz0qb2ESRI6K83vzSdykahABlU7CYzCKGTz3GD4aLQ0XRgQORbiRY/
T2VStdIcsKUVuf3cVNJip5EUM6vMqss7tgUgiPNDAnO7hn2SfqEr/F7ynivCXrZcBdYCdDdV/jwe
jxV+J3kKKO5XEcocly8rCVUo75JF7ghlsCqFmN7Gh6cBm0Z2aNSNcYiN1AD3JSjt3AqOR7Bv4bXL
QC+MvIw1nLsWOXdwLNE+SPzPwWT4N1Vfb24TQU32ljz0qgJBYlKEwwgZvw2EKXW1vcqMyeTTgaRG
V8xEqCQeY9mowQB0VfTy4Zv0ZdkZVfX2gsNe4coromae6Mat/G8fDJTpWL5wkjSvJe6S6TLUwaqH
YBbUODkSI3R/jrSN2BlsR2zLnk2geUo5LJVijaB4eCiYCKmoXgeu0kFBKHmqEHdCCdxEnI48Gu/V
pNFOqVbuL8uuFOB1h9JX4CMJ3YIKqO6RwiFIBxHE9EZsRQPHggJVLXlpdRTsUhJCPY9XkoJ6ullQ
sFPtxjzAmm9V6UDHQgNSTMhp1xh7EwPg1eNpl85sQyPqwOw01gkdrHxRvCB5Gom+GAz1oSqrLd7O
w/NDmDe20TEcX6/jie3toNZxbEJMka6W9eY4Dy0S7Q/2+cOuSAnHhXVXjxR4sQceuUe6xtVZQMyE
VxWdb1fxqNnLiGAPtF6J64ZgAaEYBDWcbvfnVmbzQjS+UMlkCDitk8aJFPPWRO9BcgUTTDBFgTD/
saPUt02Wc4hpdSssLf1PMUgyXP4IJANdtU7dfLSFhNScOvmEnc0Qk3Km9CfjIrT0uBv5ja2P2Ubc
H9G4QBR2FP62WlhsOjdJY/FXVFzuydrjuJfFpdmMlcHjqunGoGjZtV15VrKhFmZ5DwIQwX9F2DE9
HVPq34zkkX3yOumvR9gIHxRorUjYa0g1+1nDOKMGYnu+mcUUh06LQyHLs2D6mvP4RVT2SfZMaN/S
t3bW04Aop/gM4JplELZdyW+6kNWIZKBZ47Lc5YNNZwhoZELB06CX9a0HEUh6uHUKXFHr8OJtC5dW
qzsir6wiTLUviz6XrC3YS2iANNUMWyQklBTnt4VZ8gSmpBiJVtdohqD8DbvinqW3NnmEuBG2maqL
1Y9x1jUPpbwLB+//PKipKD813X14YT9KIvoHp3Ur6mL4vsHRv11jMBfoNHkHSJU4kONl7B0awiOS
ip0jj4+B4gbFdgx7DLiMfDh/viCj4VS9RutcgUn2q2xYnmaRt4xyciyzMFh3kLvBhwM+yHu/R1LI
mhr0OYKjuvtta34Irl2y6sx4CrfCI5ZZ3GedUxp7NrD6EXULJe7Qqh/7o4OIr5bJLAz+BtS4cJBn
UamOXJCf9vnDxbpHKCDvHCAlXoPDoly3ALspiCO6OliWuIrLm7r8z+WnX6qXcwl5Mj2YY9LxX6I3
BMKWUxqKeBwhhBHy9RjfS6UKIazeIdVH55SHe2KiqVVJdxWABIxss7TKB4MvbujAE9ES8lhHpqxC
Z+MB4KW3JilEaIJC3nrXWki/40MBG+gF/vfgSWIgCoItTlL+3R/dAaFyASjihVeCr0jzYfqG+daa
f2RAJ1lMBBELR2nQ1t3Dp3hpkpj/BBhWqgQAoCCBBV26NRtR1PFFmy8Ea29+gjU6IErp9t0uMSP/
agCwGZWyxhAhXjYfecPKYLokDh+jfnmpPkC5y6mMqoNbQRvT56t4D2RIDo1vosIvl2FVIJnZtVAD
Pe1kjypiU4RssS2iXzMDnzkPYGMMw6un5LQ97HLRhfH6Ylh++xR0CU0TVQVfp7YghYsWnNQRY2BV
m27ptiM1Otwk/g4FOTiaf5bhHxGFO+MK69UDzt9Yosj0F7kH+1hJJtJiAH3+v/JUKgeIk6WyoSm1
pz0J2/RU+cvEeOXbOb4n/gV199LuTh1XHBSkE6byKqOa42d4H8T8UD2PE+q7ixREsn4Sp9/Y0Rev
dDLUkBbH82CCSdF+3UmU5wYbKo1N/cR41RcP6OZxaMnyne1ERg1U4pjp+QqNs2GbueIvsppNX4mO
qBe21/kV5/FFFERTLiNBQI1f2I0MPF/DKTeyqW9At2urDBYzFvMrRgZOz+au6nR8R3Pq4RJegFff
DSYuOFxUPpKxAuXrnf7pjHRJHd/yBTcgxidErmUoiXUp5l2Wq3A5RG0iBu8209BBMtxVoVw6B9jG
00pzeAkk6k9YCtNgr81ap/v+FLMEG47x3EHjig9OIDVu+w8hpuRdFnw6ccklPhY2wSBR4baHVRaa
D2p/cRq/p66jo89ixljuafvO+ET+U47AO1ikhbBn3m5tVAoUgG37q2e4sPUKqGRD1SBOG4UT7d1j
Lxj0qTMXKGi9K2pCK9kE51xcGQ89bGcez6n4caPW1QwYUN6qxDPLXldXiGmEQawk9+PBqJykpq+6
6mlvAQpwDu/lO/iUmtXzBk9xeZ1WoTYq1IFhvSED0Q1e9Ym+Q2H4Rbn1iKv5p0C9SNEGnBQr9Z5+
eneFqHVhVoK+lhCm/uW5nLShFHoeaDOjDPOMCMT6SfAfWabP45RblouytNIgnrKSb70lcyefp2hu
8WaeYjBVlNd77Yhq10Td9P2ZDKKRoBGIvCd1RB92ZEvz+5eCrVPe49xBpxeHI01w5RFbYkkcETBO
Vy759ok/MAHdgs8NhuKprgh/awW6j81/67hoBscc93ttWxPnJW7NvQK6ogxtXlDmGNRJKIxGV/oa
dOzybH85mc5Q1k6f+PXl+2MvFtpYqbrUhfZ2FrQC7KYX6R/QNmsDZRWAHf7FteNt4YFnWIc5f0Oy
rt+uYOlJ5maIaNr0otBeUMHSNHxUZt3i8qZJgl/B3le14TBvDa2MOgopMWhsImySnXWLPwQGaOGi
R6e0xk5+nWYb3nXKtpo3/U1RP2rutBh+6r+LeAOhrJASjbQqbGIwBbR/nxIJECLPuTBAZ+a/RyRZ
BTvFAe6M3Sq5lU2yPXPvV+LgvKgf8cJhQHhXa25Ejfi+nnF1wpvsklayfSoGkONLniVocpZGoRKO
DbtWpDBRM15JI8jzA6C3wH+eA2myP9FLtvn1gxanYdpsqmm9lgfxAXrohebU+Qb4OePlqje7oiY1
MerCrzg5c6rEvKIPZbttjzIcPl+RssFsj9k1YhEeiB9iXV6/qB7kc8BjVW/mO3i2GgMmRW/v6Dvp
UonGY0U+ddTaQdoiaW3tLBEEAENbRCbp2yY9uVFEC+2nhVTMJMVWWV/TyXSs4U/4mMF9UhKGk2CR
Yu+ecUoh5xh0NS4Gh60EYFT+KgoOrUD7GdUjIT3XT207I2yTk+PRawVCBijQsLoVDa9TRt/Dc7Mm
Hv1lRu50Pn+XV3Noz7TkSeDM2tZvHECt/uNMJs7YyXAhszmRF90W00Gddv5MU5pI6OYgBlSxrVHy
COHqz93qtreqwqEHZULJM+i0841tLOCnsg/bxKyl5GUxmz3cOwoHR4Xwa0aoqFNm377mtHAg7zzi
N9Fnb2p2eriAdBBmnqBfabfb8qmLa2YLXC7/e7RC2deMJV1OJYfC+6cxFPGoHhZtYv7pq5VGEllr
XlgtARD+yFXnvWN+MOgsECEWDodKTHZwsjzaoWqyx0mOz1bL6GFLYsy9mhETVeOPcZstTk59x0RF
0hNbjVPd6n0A5B5+XVxR9y+C0xhF6eLvdt5FpZZkHidN5OgGjl+Y+WJ05mKs33XkayttcsqSHWGR
zpCGLgR5onNnjNKAdmU6sizPJqxtwLRiSPZUMEEWoiDoXPStcBpwQaDvc9rRDdwNVG9ZNDGQubHX
Qrq6/YgQIegznlT2z+9NJLBasBqkhA75zDiODcTYxUPl8Ta9oOKGFycSSBGFcBRKr2pwcPC5/AQJ
4PxVveEQ0CzNa0MN3Ln0TuIGF6nSlomlm0+g/3TVGYlHj0n3u71JIsRERpjmL12j0Mjy/yJQGQbP
8tZAtLFqi5P+ok/hmIyQ5EmkNBe3tuM3z4IojH1rJ60hXfGEYophGSV1mZTYR83LoP0O5zLIPSDa
bmRCNWqf5nob4fg/8iwh1PucTiuXQ2fnue/KS3zV0VG4sbvAu3mBkTJNT+RWKz4mj9Fr6e1Kn0as
h6ID6AuTwUlgu4rBP+ETF9C8WoYjpBTQYFOizaYebt0clHUAVZpCXsbYZktSWnPohHX34EuuFTvS
8RrLxJQn0RAHjE9avP7ei33PXuaFCfcIkHPjR5XfIXdNOCY76v8+f90qR2SQX7nIjLfQQBLsE102
LjStLNluKDzZADcyIEzoWucYUFd2QKlrpe0SyeOkJgGd1Cjbtt9DN64zH/+iCkvZeIienwL3CFUA
2Fmg0jnon3mzbtlMwhFOJubWfVUqhJVe3Nm8daE3+7J3Qd5R0ZdCHrN28uqFFqq+PrCMNwgQZQ8n
/cyBmy5pPkej3ZN4q/VnTczJG8z5oUoxgn1u79/LvmslbiqVvci6LjvhUt0c7DySvVM8z9xrcmqx
lRGM4M/V1eKjkxSA6BnBYz1wuXxa0wSgU/MMMWWsWxNFvrfJdVPUHjfpN28K8zeV8CiJ2HI4MNlE
s4XY+vZbxfDPmL1QEXgOCbZB1FgHUQ5TkEuVZZGDx2akCrD/58JmgGSctVb6glZwbNEOusAA1RrJ
paT+o0AcYgh5FORkgotnjiUvkK0zi+s4LVy1Cp3DibNH8OOochhBIzRaPkBUfIgCy5J05FI5+jNu
Bf/c8k7/M+F9JkllqO31BxbXmwatZrIHj/SSOp4c8zgKnLN2pcJ+LimBnNFmacMDExQuaxXBX8L3
wleHHtcBoP5EJngKWPQEfEyvLXa5SaMxbkjf/07eW8OgwiCcyPpI6WI33PNxUkEa/lPd+8ObR9Pv
K7lyzg/Y/g6uvFWc2j0xGRkMmhKEzBUAN6QixJAd+B2ajgSVlbHpB5SMRtAvyctlNfdPuPM3mmXg
Zk1xFazY3AjrSQ5oTE44BEyV2MhnNjh0FSA4LnwbAQFTQ+GvD8vB5/mAkWRSjTqDmyP6xuT2XlaH
ccK8dkvTll27pbq+/GTNzzBa0DCcqG4Z7k43ZpZjnxRxrmEhUS/DNBOQ8peKuRF/ihBt0LZoKJ40
1hLgWah2wYbO3ij5GwZ3q7pMsWmsRxuWNTpacLmj0Pc+J/0hAmCHTQpUG6T3/bHsCsMIsazyrETW
rjTvxRXt7bEgeFH7SsqixXDrdzb+Pg4IkKAvImKIctsp026GOav1RikVid0rDiH+0lEJNkHkLjkg
invT2qIxvVx7FccOLawchlxFeFpG32mM2r3hLuSRkuidJaDUf3IKBxmKeFZH6bI7bueLhUsRfV5V
6aZRnUXwRXGkLexLe4n2B3nM/HJ5W43yb0GCj31lZfRr/hiXjdf8yhSHwFaeSXMyZeKTyCIZ3sef
enq8RdF9CzGA2QV/qZBj60qc6jhljaMJX5VSMPIltnGfrYT1UbU/vT6hURcQkHlvaNOPzPsZuKS+
YRdWOJ1DDLvH5nPjATMEYEgNDb1wQTMMpVSrbUT97a9YMupfCXbsna2m7JdnWSZ6X8RRoFjBOHKN
2AwDruOPazLqNaqGMRwgJwtZupg1K8HbwvmeUIpp+m2q/LvyC7nh0+fXTTs4rpt3oIWoS74pgcOU
rA95JwBQSGhfAI2POsax1gZrnoEtsvtvcxjqvKDNnJsofvaJT7Gc+JRJZSDTBi3NqKaLMnORwsdI
zluQKumPK0HBJ89Pf+JlJj5kMGDJLLFoaYvTSVcld+YwQiiiN8Dc6fHO3MDiI72SjJWzScsFq9x7
vFG26B/4hm72Ff3MqWP2dSy5p+PFY7kIHeLFGwdxIjTzyRA+j7sMvB2Q4dDrGHoHVGHLeZupFukp
TXSa2TEOqBb2aCqpzMiqaHfu1WLNgsLY7oAN5KzXbhAM7CHuJGNCflaz0ZDOImO/Q2UPthejvCHG
ulL6qdn6udnIGZXrAait/OHLi71mcv7cpH4gpJyMX5k4QVd2OAYXmbpfxm9tGTMRCOI37eE0GD8y
3wWaePm940LHBZqf1QQocBWK52Nil9M/eORzoJ5QZccwEUe1XtIAsmNdIochT7E3kU0iABLQlX6L
SlquP4uGvWsKGSrb+7CLReauFYU4ANMSGOFDJEwv0PUpuBb7z/9aap31DsE19C2/SNWHIuHmAriM
97Kzb0ZBTgGnn2Bk2zamUFH8SxpwkGMaYkhL3n+WhWWH7MqPPu/ThroeO22fD7Q9ULeNbbVCMlXN
tbsfgej1/ddPh0n4FKrTEVU0uOxpoUwkUBodjJukW1ZTcV7wmHQRpx0oTz9kLZ2CYxOTep4XH1G2
jF2KyMjrugrOn8yx0zqrEpRT5d3HQtFW/oRpwJAWOUGzzC11o2pztLe+B0NkRc8hHxX7nbv4NIGr
lOCvQ0QizSZzK/KLcqS1j99PMFD+NScgdfzZ/dOE5KZVLbA4TBVym2Eo7gtAjr9kQB1nssIchZYb
WunU1EH3D0VrJLhdHz4f6qamP3ZnA5Hdxax490yLR6/zRuVPyX8Yixw6EmMIT/YuhBA1Vw3/6J6r
cEzuNZBCaR+Q4yxxu2JlISh7AvdnyycrEv6NpHYCK5gjBvSqRrPs6XXa9GEnNNf/+xbLtA/Np41p
agUlhCpUzHyhKDqiO7c4asca37tbxa/oTnvijur4BfC6s9hV6bBMNAlXsgI5WzTGNUTq+PqNp6hi
CIMYlK2CBa5mlEwOJEJMDLxSGyqyNhpego7dKs+1uFrgVkI2bYP4Crti/A6ysjtarm/mB1GTzPz6
+If1VVoZJIplKL9qGFXlJVpZXywH1Psh751Vlm3A4yrfR76BUu0N8l0XayL1tsD2ZvqaakPeFVdr
buy7Eo8PjUdEHf+Dh5/ZIuhJAjbev5VNTH5bmizS2Ammb7AzfULvTdc3Dyo9HMDuzuN0NfAC9g4X
kCxv/XgD+UIqHAtz9MKzW8dDaVOSYKe1O5rTQjPU+M4H8m+EWfWkExMTvi0+pWML7Fi3j36PSnFK
vXGUgi9aWY3P46gygzElwi1fC041A91S7e7ffXEL2KBu5/eRvgOXQQY8k92yWGJvLrZOWn/jGbPI
rXaGR8wNv7TnOlkdo9+gtjfu40X9kLNi6dR/n1jZj+su/pqcXSWrhqOi6RAEByu27wcZJMaaVKPd
g7D4SQb0A7ljhnG9WR7zNwX5M1mV3GJc9mXg60wLVrb4kOBKss5DaEE19peIeXwVlPEIIKIOM5HL
r9eMKRG0hPo4F+8iAtSBkF2r03sIDhhET1v4cOrZYqx7jBAo5QKK3aME4cYWBuNFLQlNPaQHIIGW
r9T/MeinvohDzwbQAc4CPOqoWH9HIyps7DZgINE3a+wrul7qhyRYNpzrnauLa4KOFtsQNKjiIVx8
W7w0NlTDuVbKVF4lJiGwNq23CYNxYCUazOV83hAP2KMaNBcmkdoX8scAmS6HWkJnI9MLjoLY67kJ
GnaBIY02RXXniGNeo1bkQzh/5KoCJGKs43xHW4UJrLMGRCnhokh45drjam7oCryb6W+Aie/iZ4t3
2FPw0P/ns2PpSfLSpUAdLVJUmnbioUGVkiMBxuBI6fw3tlc9RxA/8LY0zCiahaT2Y0Bsp20827iu
6vcCfzM2AZBXTxWSmHflLNAqzy9nDYe/IApbwA037B8o6LUVqtpIbRzc5AURv3W0ZLbbot3y5bvP
oziKwyLndn3fbikdyqfNPP/HMLXwPLwEQ6fCMLev6M3P+Qi1nCE1UrNQYqnntIMlBS4InL3WvQfh
ehCZ4HDBygTEqkpyk2bEuiyY0vwaTphOPckNWOzjuRh4+yQQ91SIWBU4efyiYsakoW0ZmIKruKxJ
+DH4gXy1t54X8AMv6eLFoZD9lt9+6XCR+dE0hAayo+vH8PVWR2zE7o6x/tAJmoSVn+bne+1g2gCJ
M1E39VJFIVapBgQ2q/iR53NuAd/GBuxUQNX918JAJXC7wEf4DFncNRB20UbvE8veDD2bt0ziZm+V
epFMSxqNp1rXPoihzLV7VL3UbSpJQw74TmPzAMN+3RXaDw+0ir9J9lglb0gMXB+YPGUSR8Vm0580
Jg7qLtOPk5izia6dE4j0qRGZLZQbG1dhbTCRqXb9wAC6yQT8r0q4TSqYezzIowKXDIJuWmGDef3O
j1BbiujanC07wh5l9758AHEClHyQ7EJRnP0711d0GrJ9K1MD5jigGB+zHA6Lchymlzk/CeWT80Hn
2zCZQ0l1mRP1f6pFBt7WOQKeb+Sv9me7wjQ1n11QnV8Kd5E+rxHfzu53MxBlvzjvM21cOK+sT0BW
CDb7+M11SXB0827GIP5p4OIDjrGxlnO/9PdVPUGAts4/fkqhG5MDTbmNIN74k86/j8yO0V3TULnf
hX9PVimTm4iBYsQ0tTF9vYzSB8/jpO3H6gITOV0c8+4ds1ce1k0LcpfDf0ViZGW66khaUPQmmBO8
dpKGT1isJL/NwZVzKO8HhoUlTI66sgyPCBsa5BJVRFB7kH2E1eF4/d49QWh/rTLGpkPjQSE08zTZ
XIaPlrs5qsWb3wmXP8WPIPCylmVnppHHjiw5Q+0pson/Qinf8MuFPD4V495a/tsnsGQqPoI+3bby
rQjmxziIocKrY/K7inbleSjEE5ZDxlWgpEdhe/LiCR/9Lgl/rP6U1MSwqxStiRZ6gIgBd6ZZTgxb
BdZFL2nZgzkLB6Xqfd3OJBrtFvCFz64UZiD4aqjXX6zZeDQIX6WexXKlZMWpesXRpmfmifwRLDhL
+WB+lLBBagE7QDoXb02TTzJ0rdznuRqTuuGoLFYkGdqKFjxNJIg1jknbaV11uGvQWJTGwluwaShR
wUNNASy67YThRgfGdp9VVHgSgMCuqi8Jv5uzFEy+X/fiXSzK0ZbcCijUJQk5JXfALyKxS9W03oze
boXXNkMzyMG3GuItVVU9XyH4b+xKAlKK7o6ZBf4H1UY4x8kbbafT/ScH9jvAp0Dr4T3z3wewukO5
LldkveeJoIrYqgaxu6ph3WDLy9qs6TudvOjbxImDf4QwjfrYaw49szi/zY4Iy2Cr0On8vuNWk4s6
hw/miviDlFtv21DaIOZ4UGfdi5FIkX/pYst7s3tRi7u0FFJeZr44b54ZCwnU0X+C+XH8RoIOzV9p
2a3w22nyVGOjlyxI9W6XH6gpOwMBcHHPHNLwWBzqVWvqI/qoNJrUOmnl9wFW1a99W4pv2ROJiEkZ
dgp+KuTxoeQwgbfAZ2kY7HP2/v2NxYT26geYqwYPT0EnIsBP834Wlse5qsWnIAAcKhScoqpJ3npu
7jUK/zHVtIzr5vdMs3FMC0BgToD6fJqHa9Gt0QkOfHJ8ZT1O2S97+ejNqEEAPambcrF53epaiyc2
J99B13FjAkSTLlTbXftynDuu7+MOAKwxUwv5NIum6MnsSLlKHCtOV66meDi0PBKK1efCaq9hDitK
rfVTUYF1cF6cC+Lyen8uXROEKbVoNCecckMDySVO3vyqEci6aSyM/jWcgQi+g8BABbO5gYYForFX
z/VZDwo1N7k62NKUEKo0AObHP6bqf27/JXS5vAv59Z547kpTBhDRnYId6CZ0571DvLVgDD7b1TXb
Qf0Xalr8wdJUM3rjAwWqZT2WV3R+T8pny+ar6daKFo7j6iHBaWPXkAjnQLR/4vpsigGtgKUmyuBk
1qo/rInBToNgEfDrVvMUjhiA5fKctATYE8LbBq6+1ESLqBog/NPIUk5YKJQjvjjXaBBiP/d9hx7d
RGe0Flm0xWQp+9J++Dd+dfikBE0GPBWQmrucNfgzuwbZbQmV39ygJBYAFrc+wvyWkgifURjjH16m
lRQjo3ck+JaRS/44CzJtYwoKv9cYHIPPz20DZVMaciFkXrEc8DAMWbZvhPNFY5SAr387BEsG7BH3
TVXWVUyieJ3oObo9pwyFzsQ1PBzkE6LiX4YVNJP2ssxva75zLn1AvnDrBnWqqaP4j5IZKvgtlvfX
sve9IqGg9Plo7wVN/9/bLhQhPoqUeCWvBRzhByKScYfy87eEN1V/2W0OhyINjeQzCQ1bXy/a3zWZ
ytIz5pbQ4lfap1pz/qApefHcujiIMKq3tAUsfUqxyqxKfnqdyQMCDv4WbSG4lwoJRYVRh/m7YQo8
V0ONepXKUeZaeiOzfbKZ36MX8cv87If5WoirXOdCkBqLXTYEOEW+BLjxutiacNu1dpoy3IfHY1Uo
B88MqNrfHquUx5f0Q/g7PU9l5WKFt923tEkjMLKBPtf2/jaEW97ZHj7iY4YGbNoRIIV131vMabKO
umTZFF+aXLnMxpB5SAufsDp/+M3caspa5pIElNhcSFdTL8Cm1PrDX9O9wZ5KVKudeymL1eZA1JnC
HOS/h7N/KEaXLd3dqLkRthvOQMoLfmeStlMnQt+W0bbgn0eRe/j1lJwWG973VLhm6K90tz2oioC8
ALt7UQzjhP6c4NJsooeB3pBR3oUHEVE8+CbvItf5RDMTyrY/YT3SunKKuzeh1I0H2XwWb4seNjMI
TAG077Q2eGvLOcpU2UtPcMTt1pxChdTIPwRnuFhppdyB/5vFIDhxJnkaUoPJDF4Y/BpiDg/6YEdk
CxK2MI+T21gO5MJXC/l3xAlgj9v+rZo9HcDxVEzzAre+dsQ+kLwWur3obSHAhplwCLz4tpkGd3Sk
dKnTuTg+vsDhJXYf4WGpiGP449tISAhNqc1CLHu2FeYU3cDcnomjUHX0ed9bsAUsFlqAv6RPKC36
MX97W05Q+bAmgFAY9i14fC56bLM31DxfGHCbqXV+MwdFO1b7o6F4VfFYNzRK/pCHLJZBi6+sLTI0
K78saKvCyHkWYio99Xg2sL3KwNBBbiLSQdG2WhNI5Dy6E07f9LL2YjeoQezBpWEM317WBE7zlHYS
C/7s/G8vc7mxCKsnCD7d5KJ5s9z9n8R1asm8g3ZYL9G+A/fTRMeBhmH52fq8brZ1GPm3EM5v0OyT
fmSAXMXfVIA5xQ+8rnuFezNImfuHxmNPM1P3jrRiI1gFvpsHV6C688YT8sY8G5URGFTuWCLjRSPQ
oZrzW63GPmvvPLNg9HDv5jnG4PgGAcold6WABxZbWVGHmjpZeWfE1Gw+ockR9/RzRJpv0gpdqupA
pGH6EDrol9hn/4UEOiPlBkFN8i/u/rbeaX/V/sh3V3QaoFX+mQbnyPUALk/xS/A9xg/Sh5Dn+2Uf
BuYUpYrQL56nEuKGUMgDBpjsTpbNYCAvEIZXnKbminBKFCrV9arff9OoGA7x4CIGymsUndVmyW9E
vsURXQs5AgDI77R42zCWrus0ItLVfvNEj2TC7VEYO88Yto0gDz0dNTUeyTaax2wMZf1mDAX11TS7
BjK1Vjsi3Tmo7vOO5EqO6XMekxtx2ySeYzn19yF8C99m3G8UcYAZhcGAhksPo6TB8Uuvcyct5qVQ
zZDi25ldaadfJp7ukXb/mEPLrAEOI5CVGGzoNRwYceYkR50mZe8/BOhlqN+W5SXOI9DLdI7P9TXt
USLhKBGtkFWLR0Df9z2xqE6YqVdtnoq8UT2bPWTwW5lxetRihl8l9/lrWyOdrCjzlowuoAShx1EU
bmweE4MRu62la3OpLF0EyKS5bJm/fbr9PiYX3wkovFZcHCdJpegZ3NPHBE4fU5g02uqugOCV5iRZ
97Z30p6I9ZX1q/Wt4AOKxBGCyYMUbfblps1C1993MQ7Zx8IBqxWKuyptr4tIW+6E9ive6pyUFm5E
PcHMT7lIDdTdH6JaBRVJ1HIz85zafpU2ZZHyJRCf62XP8UAgUtY643sH23Go6z+qRu9epSLCAEI6
rjNl+vC6MEpXHhfMZ4u7DwyFyrgSKicraVEZ1gFmF8SnN2c1dlsX8dJnhE/KbeYHkuvonX+Gdeov
Hxev1DKh2GM/lDoxcRyatNuJoGs4gunGNpEwWdr0nJEeCUJNxjdOqFZD8fROX/Lgjz1N4Ceuk1zD
OWp7cm9focimyBT29bgj/vbqI4Wr5/E+v3YfQM+vg86C+1R+DobrWn5ISSWOXLPdp1BY0jpAjTLL
pSOqm/QqW8HIFjAPn2oEPEi5KwbtwYwl3gn3kMUs9Xvu9JQpFJ87UUcbP1YnwyqN8Uv7O7uBbJLU
SyP9rlS2+hxSal10Kg/UE2/kwfE5YJNFv40REXTqAi/ywzxyEqWqv+REWX7ty4W2bkUXhkRRyUIP
inv2d3AeWyRbreUBSyxVDyOrfTIZIJhCAYiOzNmtPRFhg4CYmGx2e7BAwaGWT1ow4xfgf6nUkCAl
N6u3mcUGNsrDIYBWx9zapEenT4Vdy5P3JjzJcO6YwnLXRWZCPbg7QS5TZ3XQLB6xe4J1yBF+3SVx
MY7jI9tagxx2EOCrGrjCaD2PHuHo4avLFc641c3La6srKN28npkjtAuk4f9GY4zdC5niB3KGzBaR
ZvKhfxKVZ/rySJNcCwG110oKmpDoXSXyVwtrET6oltuIjTkar3t196O2KTykO/kvG9sTVAbOmil1
BBzAWRxoL5Px7FOJMd1CaUUTJOuiZFlidupE587uxptPsL2WkYN4e8Xs2wdgEuUmEpuyj2xymj8d
yzKogtMcGOZ2kNpjNhkq3Ahxk2VDznQZK8He9VoAnE8znlbfJDQCJI8sEhj6TSqA7OaAVH3bDGQJ
vMF/zlcwM45aYPPjwPvwvhT69r4C0ImJYtMWkCbVEKotMAPOymob9Q1TNWlqLJSiB0iUdJDTKX/1
uZAup7CqBcgkxlJe5iRvTDU3Vt2ne/7vspbMosmtaXccIght9+hKVqBFbznIpRF/PHa2KaRGNJZG
yTfxuCunAGBReFyrXUdotwF5t8Mp7lCKrcdVEtQ5GqdRABO8+McpMNnr55uKWKQs8FV7Opb6JVko
CZ7rILfiH4XcTt39sp06/1ZwOzRaQnzo2NWccsCCewxvxqqNV2uxi/Ze//2FlBgAvwqjPwFvROXB
Wo5+g/gYqDLSqcKP45a0QpS6hwuELedBi150tTip3wQficIvMA9dEaWSSP2D7JcVaoN/I3l1OHkU
lKlhkVl9jDoulsQolRMGpD/Z8KMOZTyzdct/zw0Gb+6xZo0ospZZJ8JvPKQ3kDkIUc0zhHkgUI29
EprcD5XVc6Ng+VlE/yuoGW2T26tlcPd8Y9fQfBdHqjGfd0dyqRfF+fxMSnVSMiyoVmwVTXzJ6MYs
7jdokZR5X1XdZCZjh/F1870tZzE+R/7iOtV4CRP0B8FZaTi7cWJYy4P/MrMrVuGBEeeIqlxHsuzT
4B00bAk5oEVoSp+HT70tuUCakFtTlpnvJuIcXLjFSDlFACJR+87fGZQfha/6sWAdqyXjn4lW1NMx
n53PD/2mwATTP+AcK2GIoPe7q6Cvg6fDHXcRi4a30jPHt0L1e5mBSuMTBhuJycIuuN/M/ZDNj/E7
G9VraKU3IQ0n8T84Kn6NFRfnK5cqPszg0A5ygKkZwHqIL2763N5LjD5/5rc6sM+ySJoysIMzCqSE
r7wKfeUjjr5a3LT6CN+/jn7wY8FaT3T+NHV1UYUlIl229eyS6qeOTli8vJq2G7G0aEwX8CrylN5a
M8oLQ8p+onsSPDFxIxaaE7/j/0XwJWVkUGqhx97eDJlUKJ1HWMyBghIUCBdljuAsmU//X0YYpCRU
JZkGn4lHfbEeJSUv6jx1/hJfwPJf5xQsKRro0Z8x1nBHdDORy52l9XBvMCm5DAEwa2fpHYlrqRaX
Xgr54cgJnKlol/NUTE42hdKvoqED1QSd4x6OKfkkaLc4o+hVKhR9u0bkTivuFkMG+7keBCyJSEqq
kn8LoA81fQIKlyhDRy/7o8dXRMnxWO16EI0YKm/TSrwIN3At92CeIogYCNC6J+Ff3tHD9LzD9WD8
TH90uKlBcOShAcV74bK7b/F0/i8SvgOaLCtFI34GpJvIPKyYxIjq
`protect end_protected
