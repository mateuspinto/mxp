`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
RIgk+idS4BlIFjk4mBzWG2rvseJznMuoL2PfzuWM61VBma1VcJ2oLjPxXVjOhJF6JCwMvC/2mhA9
V1OnVsAle1nTy4i45c7sujymS8deaoUGX0zTSh1ayZIy44MeP5uXEfdbpL7NUT0mu4uo+exSTULK
+dSty6J7UqmkSorCElenrpMmKsnIdq72bTtlEPJtwLDxQcF3Sz8XMvFy2eIkOEaIJqN3WgbYkRKB
ynooiRF7BH5ff89hsZeWq2jioJ7KdZiOrqUpeufMmzGQUIELkaF1I7OAaLi3/6DedpidCQ8chDMz
YI7Uo9DETgu39XiDb+P5E5jKG3t/+9eZUd7eFvLhRW11DY8vu/KpfbjixNMkxdQIjn3IfBEpReeC
LOpq8tlgHI27ir6t5x7/plWtjRq1SUj/wx7HZ+sBX5CysDc76/PcFs8pFeh7emgYO407kJRABRHe
dl1WOnpL0il33xNNo+eLryo1GhB7eG69bsJfVe1o2GCssgeDmdi7yTAdS/N2XZiKtH41R0b0Tax4
SaP/zrr1FKNDJkRdsZOBEAImEiGbvY8awfTKRjaKOLIKRRQmAWC81035PRAn3u01iJ0pIFr3fV8t
tikTXHr26+QFHcUZ/IS8Jm2J+3Dq2XwZNsmqR/+Xv1I1odddApS0tvZxt2Epqt3z5CE2RTVpfrMa
MS+IG3LrZHupbcSKISEZVIKBA1rMX4jk/9QYLz5xr6POmpQiBtRSm2uvefYeYBiDuCN4wF8XEOkS
5FBurg7OfJazdz7bvX/8pdDQ1tESQURJ3Me1519YF5Yg0/+cQacmUccWn6OutjocB+wPT8mhv1nV
pFHHUqN0yIFvfB6sp7RIViWhey8S+4LHkx//OTd2Mz9g2+41CvG29cID1f01pEAOKcRY+3EaAgsH
ZklX0rOsOMcN/1g+SouOqVlGA/25yu5TgG9+o0LI6cyBaILU6mP+CfDcWCvcR0dTk+fztRuD/svm
qzT18f2zWAcmuCXHrIFR5otSQ8gavdG9k2M5WGLXQwEVXT2jNEm9rp89gIbbVmJpuCGhm0FopKfW
mkkv0hPMTGY2iFfVfKPyMpit23euzdVK/sjp1cXCA7/vWfEKhnfAB95EfCFFU75caXLTzptXzaRX
o7ggTCAHfDPVBu0bWqVI1N6vQbjaGVrrpacp8H6bw4NfQ1xWsTVT+zmW1YiXoAINvnWY5WwJGPWc
tbnTSjpDJI3RlLCopP3D24IcDhbUu535oSI/vuGcdZNuy4Ea/4/fGahnwEKkMUntN2/mYVRfrja/
bXyFABMUb/Lj4bcfPE6FFz5+0tmVGRllXBo/+JjcRf6Sg59gBMZsK+9+z3/JEItyiAtIOV95QF4W
A5a+oy6Vi7+pAm7ibrmhj0XW67nUF7VLL1g33UVliPTp0ZpgatkaGukO6Gh8HuAB+Pf6VwPFMxeX
1Qb7GRdD5ywuw3r2yxJSGAksbI+N41H3sBukIHb8s1diB2pnvg==
`protect end_protected
