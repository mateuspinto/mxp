XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���yW40����=���ނ�ݪb�;[+)���]Ӫ\��P� �3AI��ˮ\y~a
�#cAf��	|Ǥ�$��^B<rm�DT)8Xm��P�aλ�}f?4�^������x�R�f�n�ss��\PM4�$ݤ���(�%뮅���9P�]F?�_����u�^�Ŕ������
���,�Sq���s�Z�����4�;1*�ua��2k�Ķ$m�� ~Ng:�5����f�h�&o�RG���4ʠ�収5"=�P!�M����'�Y�U�\��^�DS��t���OX0?΂|�mQp7� ���]���9\]@�ũ����Ցb�H��C&� B~
6���+�/�"��$m^��B�A��.���ð�׺��O��d��0R<��a�w�u�<x��7�^�.�K�Pk�@<ft��E[Z��>�v_��M��Z�"��8�:"��f�;z��o�ەM/������gs��[�T�:��G;��n����ha��HXat�#H��i�om�+�M@p���x;��c��!|_�V��Q�蠆�eG�5�@?(��$�yL�<��K����@�^,��>T�J�G_W#R�u�e$���	�.�
�|4.���XI�pG�D��P>����e�K6��3f�Se��asz�̭R䎤��CL�)��Y�4�o+�*���X�w4(�С}+ .U�Js4j����6��>H�2ˆ5.�����am�3ۏ�Ek���BWT:^Ap�"���k}E�����_W�84��_XlxVHYEB     400     190�\K�|rV�v}���L�F�4��<o��U<"��(�J^w4#���7��ϊ��a���)֔W=���o���>[��XS�Ď�bo1�D!����N���#�[�\Q2
׉PA�.	��.�<#�`��t*�׍�|� �<1�����å���J��1�FÇC"}+�q�j��O8��|p-76�}7,/��-�s��{�<�3t�q�BS1�^U5�v�
��5E�Ą�������cUG޳U�4q��ŉ��6�0�B��[��?dG��$VR=����HH1�%�s����]m��dj�B߳?��4��u�گ��!�1�Q�xG�{x���6��K;��FĦ��tf_!�GM�X!��5��v��ob�|�X� أ�%i�ۓ	J�Vo��T�ڐ�n���R��XlxVHYEB     400     140����"
�ڱ��d���(��O�j ��wy�/����zVOW.�
�D��|r�3��x�h1�?�1�����D�+?BU#0��\~!tْ殨X~v���4��%�t��r�k)��$��xD3Rh����b=:.�s�{��Ne������u�2] SUR#�+/^Y*?-����1F� Z逍82�G����>�驒�.s%��%\�Me����"��+um����&)��O��G���jwJ2�����s��2�n�v୞��>g!��*"��񅇢=��~W�J!59P){l����uD	V1d�޷QQ���Y)���͂�XlxVHYEB     400     130���9K�'��x�����y��4,Y1��d�n����9$6	��*�:�~�����0Cu
�H[�v� ��`d��/\Il�ͻ�2*��dh"Ii}���o|�Y�H� ��F�KХ�[�A
��g��-� ��cw�0Y�1�R�zn��\��p��������4DA>���c�P���&�rI	���i��Uo>Uo�R��P�(b"�E+;)�o���� �	��M��}
��s�#�]V~L�,�B<b�����t[�"�dC�e�
��9�sZ�>p�幰�|��L�+�k�;�W!��$���3U��CI9�ФXlxVHYEB     232     110;�x�!����J�$��F�}��UI����e�Ď��(cd8$~���1Uh����'��1L���N,��ᜈ���P�x}�I3��?ZYJɾ��<kNȋʨL�j�47ۏM�>p��P>P�/4�ㆁ�
�t0c�^�K%���.K��-��.��h�Qk{�h ����y��U8t�6�wo����S?>[���9���>�N�{q�"��[\'��/}�v@8�$��ۦѵ��h���}sϬ6_B@������Ѳ���d����U^(��rm 