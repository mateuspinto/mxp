`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
j5BFvzywpf2jBv6fzVuRhs5xfw8K4R0sMrjD+pUPvQykIvaSWNlVJLi0EVas+0No48j4uoqmNlOt
FPszTnipeRv1Og8II26xtxcWpRMIzR0KTMyqS/4a0UY4hm0oE7brFAX8E1q3OLG4zPunASr1inFl
y1NRlge40r+A6c4dBhWWIbwdUJmjoQaKIlmrspR6CXgE1yHF1oFeW4XbPoy3ODijgn6rijJEzabS
IGqEaxYI9zhubCuc0iM+iqgt4cCle4Fx1mOvCjQHixmvZE2/slJVdjbxMDJdnJOLBNHth8mRZqnk
/lfdX9pENcOu+Z8KNPeqfIhG8JfBduk2by6quw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="HVvroYff9pUmfvJPFWjJF5F8wxTd5/ftKby+bYXROpw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9456)
`protect data_block
7k17a7bTyxw7h1cvWdO0v99zxZv4rxhQFOW/89xPquMqfeLpa2qUBQ9xnSPecXW1JGAjA7+ZF09A
+9k0GsP/Szx924QiMLWlGjDzXH4kCCU6DoR2VgyYr4MMVxDuAiNWACo7od8NhbJS9xHazQUa0a0E
n/i/IhP1BMe3aSI8uARylflmg7dxwbyTYVQYkyE6x0olBRUvR/fYpknZCFYoddRiiKIAbOb4apqb
ydgUG5C6duMHOnV0xe4XGB2/Q9TGR6NsLgubq6yJDoPPB7WTuNKco5QYee0ATVa1I87Z8seSTqo3
ac3iHjvcAuw73NCJbe+nrUeA8v+67RYRFu+m1Cdk4GjOBsmLkok9zn70E7/VqCv9nX7hlOoxp1bV
B/tWZGnnuu68eP8a79mI5ElKA81Bx2s5g+ft/n4w9+0jBAhUV22XC1cDJDgt1K/kJFCxLmcblFW2
bLNgjnxPYRbxFpM8HqyGQq26IT8Z1YgI4QvnKektasqjxIaSacsbjcn2IgVBM0pnxc7+sSQ4R+Qp
SOeGbsEfnv33DB9kWbqGnCQ1uvg9WNSZEX09htBfvkq7bdu5H6TQZq0YIrYI1S6I8dCZcPZZc3bd
bxNyNh5LMLoZW0ivLpVkrNIkiwZY2BJEOrG1L6AxGdorc+l7C+BKw4ksd9YA/nsSKuR8Bsqf6G1G
9ijlF5pfekNpeyiTINOBgm58T9SI3kjBObhK9Fy8Hi7TLlhrERwTA8KDQ8X3Jajk+QOKlW4iw9Lt
OJO6e1SUA68suVzA0MJ0nOymyTXXZ720akWfpQtUhGFoER7stUQ6JVtBxEf+dCKVDVTi5L2C35uI
hvXDEJlJZiFzJTtKOwgGJL7roXFGVzSD2zsXhnIUtrWXyIVoz0MvrJnRKV6R5Lbrc9sOhgOBe8Ae
45MlEnQHKs5guWCNCGvv5FFrUK+CKMKFxJk2Kg27Y2PPYc25x8SCeDpWh1jP4aifGIrPig2ixxjv
GUcPmYZ70vZshSN1saMUqdqFxiLsDlS+5bVZ9lD2O0gjRN0+rTyvg62+uUQV8JJUxDfLf8ZEOVJI
JX9jbD9yJPdo4fpkM1ovbywwL+BqWlyFkV2uj5tCOI9UuZSrZ4i7hxgKwQqkH7kWaF4q8xOP7tRh
6qvpEwx9hir7ija7sgmGfoMMZxUZduzzWbogUOOQwPjMMKb399mrbzgAzZddSZyndQENyyzZ7Vr5
JO4QMROz7eHBsC4m7IYj4JrwSAxM2CN1XYBGT+yBHhVeIdUt2NzR5DTzlk8Hu7niJROfPy0QRgeF
sGQ/IUp91Xm8A7aARf12pZ/k8fzkDKTUx3LYD4eshmyz80uV+qbVAamOY56PIwDoQsgfAfznry+n
d5mwIK+VpSsWfQKyYYEHSRn5i5jiSzCuclp4UAe32iv1QJO0NZd9tCSag9yyWbSy3aYej5B0MUFk
Eivf95/RoD5zis2ddICLjiDokv6v1xv5dEsdTGZkIVOZkeVJ3GRHL3MmijpO6HZSWzB9OcOcUs6u
iJLcRJR1Kt2ohwwlnONL3O6rr4y9i10Byg0bpl0scmqpeb81U/qZHryNFoVVLJcsFNlmWGw6o9gh
wMxX6k6HsAVC6b5kdGel2bjRVCS14LVITPC3ljmlBRlK14A7GwekTXt2+DlokpU3aLpyEDjmdJmc
usD3o123GY3NUZT3yTwcPI5ZaHVKv5htxpxAPLP5blDDWF+2+3BrQXl5pQ3QF4ZeHKspr77mlz+3
6pTaEvUOHUZKhZFpaCXOx9MDSVyO+9/O088QlHbej7HDjUc7o534nMS/BesC84V3FEwGf3YKyHTM
Ykgq3l0vzvZxhAiEnBBz/2cwqzKmXg88JSDer14khLYR5yYyt8/Z3dvhvb89tv4S0ENZOMZFSdsY
Dz35AXwxR97eAflgB80SX0jX+yw+vbLztSghX5SuVWv0gpE6Js7iqPsGf+5EjLRWq9bxWD7tFdTE
dYPql9PPvyjV7eLuP8GiHHUgzOPGImN3jZfQpYlEJ7BBPoyS6rwE5nZmvSYsxUI5MxUpa/KwFq9Z
gw+77ZuZ20RReRRNFIn54xSUP5ddch24p5zVsfiO1/hb+XaOqsJEp7zVbu/b4uQJkIAtH6JZ43QZ
3EvQ4iBhhhJC4/PPaJhD/JhgkC+LOG983j0tbp0I/xjhrxWnZfnuNXXtPBDWEB55m8VOX9XHat/p
QFiU5qRgQ+sW1ZOpOOIfpiGPC9jByTmn0stEUHwbxCYewzvPm4rE9oa2Ixj7epLOZgNG+IRdenJW
vTLO+p18diuu416Nd/xB4fcwUbG4KrUhI7MxV+TRmUXnfcQEUA2Fj4xp83NKh/tZ0U81wJvKbrd8
kQYtGb/E+EC+HuHK4Z+NHYixrESsB5jIPFieUUMAzzpFpz9LNZBgPiIsjF8b1UJ+pmWpyuJHHCD8
P0JKQMBapj659K1HDeoi2te1J8k3ooRsWzrrvcoipQ/JysoBvvtJ45cF36dDB64D2LXMrtY02mm2
n1xxhrECNSSivrqwcimlc3hSi7rp9XRzLrGtzCwX+oTrEd2hW/hZkhXXbTz+MNOWkROpE7csHRT3
GFUBVK3kz4cRki10fEJ/p0Z3ro2X57fhq01r1ZwOy+O0ko6cViGnJBayGp8nbj2TrXvzY4FxRB+f
Nyoqomy2VXzRtUyzCnmtw0IfhZOLCgy95KNF4yb23z5l0pm2ZDKjrph1Z6ynWNXMUyS37fgzSYnW
vIl4KPQqpXyjLVT9Vo6LopvQWKj/kd+W3wZwzvMiiPo4K2qKOVdAS66waABk/dLhCa9tnSBEpfqc
9iDevuCYvmc9TCFbUtbgUtMquG0itl46mvUGI0FBC4arqkWiqVPDOTIqCEeNtLHd1uZeYUxe1pVW
jXZgIA1YwrWk5b9sS6BHkw3pjSlvUfPxPUbnfHOGXt9esL38Oqjkf2nbb6/4mNIVDsSj3VeVbHyK
xsVIOYheKtQlhAy8YYnva/vws13JXAuhnGz980dxRLX2XLfqpHya3PuzH3Z7CdbfPDYYWm0A9pgY
yhqIZyPi9tS/IaVOcc8vImW16ux1b8fgYfW/ZAb9QLN0Ydw0p2JK0ddGCHPeA8bczMIL4SutMZh9
ofOPhs30IGWcCi5H1BGwiceZlRGI6uiRJlpEaLWZaZnbQCklud//9lDL4aemo2gli5DXBnov+tl/
Q8VXa6Os5fd4/KMbMBsH/Ziz23qBHIA6EMywXax0/cYtV6QXcHDE37V24sLuppUfnZi9R4AA72UT
D9F7PiJN4HssUGDIMvseyzn7Rvq4hu63l+hc0kwo82gPl4Ce8UxXnSVxnr0QwdYfcIhALjvboAQp
ARLBX9EH34OBlEekbkVzZRBgA7vVk2BfB37wG7QjTC6qK4bf7R/i/f88nobXTGVG8kOTV2310KXB
/ikxlKag1bQ0fINmJ/yA1wkEdJqXHoVkpcUEF7gY0S6c1gJ6FByhtPcccqC9DdnNCGePwIM02OLZ
oHPvBYQp5UAV45WiBZ5YATlvsJMhzG1y0DrjmOS2+fXe6eAG2wfHQ/7OpkmmNRPyYLsTXDE0rwiq
aSg13HqV8z5Vo7nuBqSlgHW70rneJENdzTzg9J3wGCfk2+BTnAciOn4VMC4C/ePBG0njBHcJlY7j
vza4iuJnVbyPjG+0PIsafPAvcoJutf9ZwBk7XAuZ3WAK1EjT0Th4jfk93cJdnZiVLYzyEqbshRkn
XKamTdNBznQTHjX+l5PLldIuMRPoqOXbYOQUM5WAIYrC++AoS9ypFAxH/YdaNIOknt7zQVD612IM
RHsyJW4wPpCMOnoH8WDu+xcJy5dRCbhNYdOfIFDwIUrna5HfmwENuHZ33+w+br3GTKRH6AZQgef5
ABfi4GVx8Y2vptjq0vxzOEBeNtYHAtFs/83eJ93W9T7U/2/l5VCAzo7N/q9m8U4tyb/yJOWwzwZZ
LLIuPJAzapHWpGvgeTqbr+iBWC8B1eJ6QFi+O/FoEzT5Jfxu8fOm8P/wQTBJcta4GRYb6awVnyKP
FOrXp8TstudKaRzJLQbdMjAZaBzFAIImHFEfVMFzI2mhgdiwRrymDFUHefT6RVHn/7aKS1Tp/mq8
QyhB5AQUVRz3oh6F0XaB/RBLN5KRaPivczXlpyxVUxtJ66XSG5/YQEu5Chpm3Bj5XiYPKbSOVFu0
aLvjuMFSqvirNktVXDsaV4KGOJzIIIjrKnCPjCVwDbyoj7dyxSBahC7hRoKWdSAVvxM5j7ZEXVfZ
DDA8Iziht/WrQMipty4uELWrz0VcuQrv+MToJ3WqQcXrOUUpHtHGw8R1paCRsmONWSf2TE8x5QcQ
fqFCGZsWEpHnZnP42ETYz7yZWRC0nQSz+x65w4juVloYW6nU/7j78GnGVR0V8jIgb7lYykPr3IPk
715dLIA2PVFnSiaaSRhfxwQqHxYyYza+aqzKuuPvXJeAajISwBxrKQMqhk7ioj7UEp1ZwndJI14M
BN4c9qsOPKDG5A7lxC5bXUOoi3UujOUhkPfDEawfOscXUqJB1F1Sr4ONk0/VRgv0Cs0SezCyEZBc
qPGXNuuKDE4Dk4P3n0XERli1JrEhPgjTCCVeQO8z2rTzlECv76kE603TPcfHZ5rG8wPLn7DcWQei
pNM0KslpWXqoCIs/mFe6goWvK7tag9qx0k24JjIrR/pmoCyXT1RKxf8rdYd1+zAJxqivOYWX6e8O
DnR9PRtzIF7NxcvIem3Ga2wWxN+CXD+fuXrRAsSP0jkglrmes5nh4Otg4R+rwQDPB0vSUS3zw05J
NxJpv/KULdYkE4vVEmk2uDhQ02aM5YShLUWqrIxttWziiX1lB9NLWd4hrKq2FB57ZBupnhy15PMC
D29vIu0TZI/cwaHRGoH4q0pMxHRX8jUseLS3qZ+mdKmUOn58/uMUpeN4VNbAKzZAh/YI2xA5v0K0
lz7BFGowoGwVQNekFfMBUJjp9vFUcGfeDe8R0mxOhDEf7oIvQlS39kzuPlPl+2YkDZDpIp4hwnWm
WRReHkVROe4zRqOgdiLSeN6uesb0Nh8JixhgLF/btZQ7x6wK0TxEKqbnsO9Yr/9vcaN+umqRULu7
9RV8pbFR8ZvuUONmppfP/3hRbUuw9K3yO3qmkkq5/sq73VM9VwyX/8zXoD8BOmmxJdpqUJHrRKsX
/FqBXOUggeolBUwf935PT598UnEWvVTARAGFCyf13jlOhQ0h1oR0lV5yUpEi2GoNNP4exnLKdUDb
Hqkonk09bUQDlsxBMwDZ97u0yCTQzxRjZrKpUzLadK5XA9q8fXi4MGjiOt0VPKO2jNHSRPAo096a
3rsonQ/lU+7V8hmcv0R/+ClRaT9GNkuz/oFVNy3ouxl2oQb14L+RXe31ZXtNFZYg4zBlHV7XR2Xy
Zidhz7ssVYCjFNAz+p3CHUWuTOiGb4kwEYgwcZkxSq/Q7sy9vXsjsHyyWbvd1/IsUFpqPMhTapvU
44wtZb5kAGYAy40PF5EizCFdfE6QJ7O18079CVTGl9v9KtaGEHFYOM59sLYLSXQ+WJcxz/gewXBy
N2q1/4Qax7Y0mbO1Z0M337xXIzPmqyCnKQrgsGp/D1prZmQcx4qnFEBmreveo+/7htDTtlwWx/Ph
H2xWR6QKXOfQMyw7OF3sacivJtcgJuaE2VV8MlkXQQGkikk6xPDxx5wOvBZdlLDNW375FTX16pO8
Kc+cwPg6uAXIl5xDXIl3vKZYQrLc/VLPxeZzvVH17aKXnlcfQqMN3bTEKB6xydXs9B5xe1vrfYVU
M5G1nw0vjzLpxuI8qSKlDAYafBj0kIzRUa2nuJkyF12yzChBS0911Q0EAfeK9BbAcQJL1z7fFeDp
hTL7YrBXyk7g/D3CsC7F4SPOpfQgmN+a4TnUZVHAmydMsFifdrrhMDc/3AA3zZyH+u+kr+qeya0P
43Wgy89dxHymtFsHTzmxoJs3K5yRNrYyGX0bU+vwsBqinFpJ73VtAOPrSJ+gTAJnVMEYa4f+CScw
WDWm+ZsbRyySMSkPgm91ArKe5QCdm0Zl29KGoo6Gygkhami+Tf2IrKfdfU0IPB9uajlTTLH++zA4
8VIiGQnFUDW4wm68AQVU1Nikudk77MUQW6cCyhyJpSqDSORz9Xaf419wWaPfIVGBsWLjYJncLWe+
iGK2q6vJJH64slH5pwXjh8GB0GSYgts7PWKVB9bV2Osoc0fK30GxnJA4RQS26l1OFtWr1CAbXD4H
GOKOaQNpLPC0t/5kOsBn1AAoGpd60deC2mB+OSoVuV/iJqX9uXGtDnCi5JbRKqdm9QQ26sRuFIVM
Yr3EZMfdzwb2exLvGZfnR9cmNb0HzaC5OIz8wzoGny2alKIci2M6Gp2xY9V9QEYHKmbVfFOI//xy
VTot/vw+t9wAvzWjsSyzy4RJg6DXOMBSZF6QW90CO+Hlj/U47RxWbA86Yy133coybESjhS+nzBCj
/YgUxB+zSCqS5Gne23oOP99hTG6PTTmEFthOLaiCIhBO9L3W+r7zEjmtLJOD9HXs5HNrhoeyivdC
C2u/gmmFbZJOKdwQkY/swoU0GVCUKRLjriypZhxlQue/mshksqQao3E+UAP7vQKtYdutK/Ts0kWA
iX3pf/mrAzhrtca21aJxUq6xtByHmAli2ahorTE2iQ/jzCnCSR7O+aCgK0P1+LGidI+ysHW6Dfl8
0vWcHbRosPdyKTCqZUkGScHdnkoxfnLMU8Kxins6q8aAnPfKXVQDLlh7osXKBAwNLxTXqtR3LSYe
QT1AdeL6/hKe/4w0NNXWHu8Ku8NLW81YUAGj2+y7L4tQeAQ+ONWTAkPDeSS3oQqtNVPsJ1DeR2jZ
NDz9/7JqlGhMh4JpzBNMKnuXXh0X5706bAGC9oKagBXgmBf/XpbF7ws/0Zc+unb9jDGccEDSX+1Q
oLJINWuBi/sJD5Pd2sFSfWfIWFOs9SWhPjDpSS6vDarKj4QyKK4yhdDlQHIr333E4McsRJn0xhiE
dvIbkaoR5jB6pmTC11SE2OX99jCzApXTRKvhT/dsCsjlgGn/Gn7OJQX0lkbiiuZNIK7uqpBTtJ80
mf6+qoABnKAhDOb6lsgyvOQiMTrN/8PvASsggY3NVNyBLt/Vu+Swk4LJndrg8vEcgXEgqMnVJPO0
zETCucbcYG7/zcUW0PKeaexjAnajxi7xoKvRX7q8rtpR/J6HBMsQZyfvogaLF8ApWVnpHO3Te/52
/RRmIsZfmZnr6g4676DXQ2rsuvFOkCZWcK3K/X4Acq9lmMYa7HZV/vc5GZ1/wrLtGofhkEwmplNe
fuXU0bTrIH6xMx6Ut5pkycdznXGmfIm7PMIGFIIveZ+ZvZTt8jwO9Fxr1ub2gTHrbAueQ+ZQe2pV
Ctw11V2RCdYW+op9+7Nl4p7lgrgXutdbC1HbF5/N3SzKtdNVVG1kG6HsGxkZ2tB7MgzUowMz7ysT
rGeoI7+8TMSySO5kxpMuJoFQbr2anLMzNbUbR9Wum5K97aLhxB6GGlm9/mLQ/ZFWrMweyk0IMS/Y
LFPNJ47U4VlPI43uN3oSxzwLPcbGibRcUuPsIXgvqeChzXsGGJ+1krcU16g5dpmimIWRMt7ppPSS
eRkP7tskbon3Bd2V7d0j8ZADUhGSc9bI12de13dzrPP6pLNf/hsDdu8Wv4BYn+VT9nShss4DY7pf
MAkMZ0mErSOPNjxbJ+XfQCFHIzJn2sSuabsYuuNUColuJlJzzZKs1nduQjauo47hLk9X6m+okFyd
S2KaTlDcn9OQgbn6b6Ybo8I/wantYxpKtQyWuzM/Sd9UNEWpqn4qcRdf3DgUoAVgaZVaf2GeG5cp
bkVKJhXiTq2UbgNZDopRNglw1AdoT1fl8OwzAaYgMykdclP/ZOVeToFB5aJ1t4IgXqnEZ2S29kmY
USlnbiFBOKsXa1bJftdF35zZG42N5H8IjId3jMtAx6OVl+7M1kC0bO2bi6yx2HUfRWotr3CDg9yN
lR/X0dacF0+qaPQVF8uDfErG+NdE9NO6Ie4/7sesfXHz7zisgQlVuWbtoVswPRUqW+vXwy0xfHGA
voZ5gi/YDCqlgMOhn5KER1LqLByyR70NbaEz+a5YyDOSIcwKBSUL7SE2qyhZmbWHC6CSnYOGrW86
f21gidifjg7slZdZAnM+RQMW++dxFlNYHlfWWBPH9oC4VqwFuGx4HyflxxUo5NDQBfLjmkJkbQmq
5GFHk6CpwlXuDO/ATktGverGVH3rmvdrHIdV7ghChNKa5ewOI6JsdRZRMtzTHnkBEuh7mipkl6cc
zSndhqv6SsbAOGh10nf2ptgGOud9UnIuVUwRUzQnMJ3v/OwMPfpawxv+LenyAb+t+mAYnz37LqCb
bwZ4WE8TdYoEYi4DSFDnk9UO3T6qG0tp/O24xOO6E/2LHPBgrDiHZQBXS0Pl2VxjRATm0xMjOGab
DT1fUwWgGo0iC1ehi5CCXlWXBbHfIeEjuin1xrXu8AFiZvyjIFCzugmqyWeBLti2aaUbmCinvsHg
aw7CV6WhCtd0vsDFNEpYRTEfSrOnaKOJ3llOZomgbeKigv+ZDozJPEVJqv0JypW7dD8JoY+z9Map
TUwQW3h/HAtBLVDYbJIe4h9U0wdfwg9CjbvmnO2F0oV7JE+VR8dsHhJRPetEFCGiDR8+gegIN/Gw
4bxLUhICPDhGeUtHcyeXSN+ObjFUr4Jlyx2wbVHR2fdioApapOe3WJiK98zOdiGw6ZQa17eK4gCM
zCLAqyiwuJRTOSg7Iy700l6jNhhKUL76HPPWs23Tg36d6BKcGcZ3nM1matEokcDusRTU0JLGs8Tg
8d5khVkVYQ9uk7VKvFBbiSjdhEuIwIG8qexGmaPywbCthYgjL+e0C1X7w09+1jvLSy7eJxjuSNBs
RKQtMfMNTuTX5eJAgUpW84oM8yeYtRWvs0y3i72a2okE33Fl0U54EaxnaeMluLtomuGaVdyT4FqM
WMOG3apcQyAKCcx4yBZbhDmLmd5L0YuZzIHkfWf7CRAl4bXEE+aDT1JRbsbEp/z8aoqAEs4t6EdN
N9vKXvsQrom+Q33ZMEG96LC2azvdszztWUVzc35DxP9/GfCiuX+bY4f9JCrMDxuEumlC/MrP27R+
C4wHBOD90GsPHSAHAd+1vbDX729lsMIsbNTbCsjhkAF4nIxRjg/9LYiz+whzYSotpIEjf0TatKmx
0+DIMwQMMrdPbgBZA77s3KVZ/dhKvz7Knk++AVC+0KK36eOITFYSAs8QIIb4YlCiZOAVK1blQa2i
gfdRwQjmjec7LMrCfItA/KWKNGvqyItcOpCHyX9S4evH7t9eidVFLIjrp/cjoQItyp5xcHTmJLG2
krrMlTXbj8mTkT1PAr51o6K26AfTU9xuFFXdubSGvxIM54trifA+Fz52f2el4BkDy95TbH0dNrY/
vdwvRGBczdPOjhg/170s0p3XYsIO3TIG1lMRrVbBFA0/3ZFazFZNYyphPjeTD6HCCcwLJ2+FDWa9
qtguerN3rl08UJonObAydCluMpiHk56nl+ZZJrEDwdUarIrkJ6CaODB7UqeHCnHG8gMG5zJF5ey5
d3WWdKNBV7k55MMkTGCiPbOqLqH3bvMy+LAxpnKhmtv517ZZNdtgmZfxb4dy79imTXvQctb9xrcE
eu/ivlAaBw6llzD4hl9gXKYSIm9a9czXhktk5UyKle/d6JWa5BXc6QmCkLFQjStheUFypUfFyAjS
IKhbGrNEta32uiTh47Ucn16+nmMRzjrHHLqbWk1NooUzRtlFiKAdKKYWXmmCzP7beS70E/NTO8H1
HNt/JNi4cC3y7o5KbSK26sUwKfAsnxeK3AuXhfDtjmZ0VAIK6T0deTwXx8uRDjdJMu5e0J/cxxZP
gFsE9x8PL3C4rnHta3nmI9v285ZFXqF15eHMBNG/D9hsv+KMYIYH+atpzTAbi7V6xJ6pDkysNNER
cGd+MX4AkWWTGJEHPODKhY+Ydvkx0jJQAKU9bDZUNTKH+k+0f2NcNv0wdBpctxOpqyvywJlw8Umk
94cyelQNk3mdzDp2XuuTrBWwr9TgdjXkmd4qy9paEFnzOuL0d4IwRpEZGB0VYVRSxiGcZZdDXRd9
E8pAEWJO6oO+N0TA5kyDIby1pKZTF6vB+XAd+857f2zeSbX2Z1/EiRonRMsxplGRD0KCu1Im6o+6
GNoKgrlKWmIxqxZL9kJTIUeqGLLmQvRy/tDV6brBTx5fvVsOl43+9IXChRfowlwUucTbOqXFiOJP
NnzIR0X1pCEQh94vCxxmhLU65i50u1HNP/j8nAmPkv4DzaqQ/jIW3OVKuzSc0aV/WZA8nJF2D16D
erCSQML7yChs5f04NCyw6Ys1dD9NTyxdNBa4aX2F7udZO+VniLiUYNAfClufiMWLZYmlFEioQKX6
pHRD2DnxwfYSx8WsESm7veZp99TKbo+c1u2tDC1iy3J2K5CZIbDnJ/rP5ChXfnrSizX/GbukOGJW
54a3wsRKFZvEeINNwM6fRTf9k28wsuB9SPJb0F2SPIFahb6sH1Hm19ZNOqwq21KJMsZRK0qn0mF6
wp6im/lCnsizdujQjQzhnzFB3ZmggZ0FwiK2F1f9JWhDUjGUsk8gAAQWL+qTo27HvVFt2Xji1wO4
2ZqpamvXgN/1B/rPrSAbCayr8y/F/800k55hkvxQhOYOAtyYIqxsuQ/IATLdKTfs0Pb4cOFusqsw
qQoPoD4rfv7E1FfrdCcne29i46TJlk1EA5unXYmSLAd+JfIbUFdvDmZyGqkpGel13rguO4eIVFrN
l8RE7ofhUEwAb4KXpAZDmF6RHx8DIwyVQQVWRC5HZlcmbHPx67UqblQX9pWteYSgC3Xx85Qn1GAl
RZXDc4oqsalolDhe5dacTizl8CxE8zckt3NGmpLJNKkgr3Qd88TTebPLp9Bxn+obtVVRahASW2aX
IMW3p0BrDOCPxQayKtSOBSU+iK9m6djRcf7pGKuNhoQ7jkmuzuEzcg7sCvz1RorQiUD/xRPEOuZ4
MbT4rSyYIf5DBeCp+8wN7lXmPlNAeTn0yOloJehn32XXR7o57Y3oCI0teRoDLi08mnTKRASrOQsq
F+1WvjrEn1VgYnvSQN7l7aGedxVKsglZYRG3TgqJkX0UbdUCWE7IGRqY1nbua/Tfc06OckVtf7jk
9BYOqJQEiXfC9vf6jJYXdU83IumQOYjOx3PTMXseBFHlx7soQpVScgRny+vldYF1zB2vMVEO66qh
A0rK+ch25wYrPgn+x9qUTNcfP83f5vtUm/XEICM8GeVgQXI3i79i+4N9xoK3Uz1Sw1oPl7k1AFlL
k3dc/R0iqwdBSIFqiV5BY+FKU++SKiTpitci/Fs5XFuibANcPjelciiaTzCoD7VEtF0s5KMah3Fs
wH2vNeIAlDZ63rgITaWqE6J+hfqovGS6Ax6EzGtXFpkfcGB6FwZq7WDYSPgq6KxqAVmoKfZA3U6j
pHayIp9FxkEha3RKSAwYUK3YzxIds7IdR2QXNoMxLyH/NuTspw9qopNKjgrfvPaTILPA51Ke4oos
f1wzkNkJV2rS6iDQdb65faqeGispRkIbKyFm7WxafUbNT+PtzsA62L7cwUzHc6oOz7lE5QY9f7Kp
h58mugST7pwnh6kA7XfBksaMTzhRYB1beVY0uTP4OwBjyVvidk0re4R+ATbrxQjalkpQ4V+N4tGG
G/+rI8+dZGyI2wo8WHoouxiT8rQc69me8KpdQAxT7gjaMwmg2Sl9968hsKAQnBNEkAKrf5FC7RiZ
WsppNFbjPyITvAmCsts9ugxVQ1xrcWgXFI1k1l8gh/1BY53OrifEgwrwF/CuSTCizJq9DnWpcfmG
D07X9OjesDjiSJ3EPVgPK4zJdatPSJ4uKUIhg5SpNSBUFH1PGFw5uk0OoPL7CZAHk8b8E5YJ+O35
6dxQP2dqyhu2iPYTmb+RoRDWPj1zZtrWmPeS0FoJsUgE5Rl4m0t8m44MvRgeT22O+owVnj3fV61a
qdEUTOO2yEnikYq3H0SXIFfDeOwkS5Qbi1iReKhfIWYqKviBocRQq2sFItbjg+advFwYNlwYH/8Q
jtghZ8vNlKARJc/dy0Kp8ewDUqKJIWDNeINFQc2F9e1tkGNF96IX6kzL6SjW93vnmrp8sXd9/8vr
Fc+EyvBy71POONUen5dfRnQ+cwWZqsVh1YCfm/DPqnSw5+Mx6tzX80aH9EDYyfBvCObAf00hkg3w
7QvbR75b946bAxhKeUjezXZKvEXerTAxoUYCBbA1v8EXVrSfYXjq/lL9QgWyC0ET6Cv3jvKFs5dH
Ss411JHNIlsdyMhaeu4/vIQgdVfQJuvlCjCzt0SZhU0RXwV4KxyCzM0+AZN7dUg8YkKofN0EeFbB
yZvqcC2RrzRO5g+poYK5Q/RuPFsOR0Iv+qPOfyKozGUQjF0a02+p+Nd+C286ThaV22CUzltLZbio
WM7a8D6c4tXOqpgkVwaliU/gz7q75D842q3CXKWLljHmWQTWvR3+BNfKmz2NiJTPGu4psgpQKDad
6xrkROWPUBkKg88XqEs/Q1QEuCzYGGxwp8mep2rYXkvhfDNpJ6ppY6ApO9iX/x88JURB
`protect end_protected
