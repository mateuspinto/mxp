`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
T+vwlj/JQEeux1EeSgNq1gWS96H+kxA6UYasMOkz02RajI13zN4UHDcpsxWTETg/DrXc5G8DW1wk
40gnnItfTt6LWE8T6jy8tuUk1yGdWXsKb4RfUKmF0it5FlZLTYFrbBegKSZXVpBOjUD7y0zgeXyd
jG+GPoaa0vsXcuVaNVm9sOpXWZKYuFJJV/Ho4k85JlTodwfJecbWrp8yUVYNw8cBHqc5sMbH5efz
uj12wiv3Xj6adpdxH1l2/TP/V2qLwq95P3hWsneIlfmcpTxBMzM5IUWUC1QF14OtslrS06YMxai/
9jyQks8+Xu4iaDH+T2B0fTvax0AXDMh77OtCHA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="bFRlYGDozH3tQ5LWC6r/LlPLR191epyaQNfYdFArQNw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
XvY0J+/aWUWFQ7MerVZBpdowj3JHgpH/hfaP4HKndJlGfjrk4QBgQUjk9QrmvRgbMqGvZe0gM6MB
wSIDevh2HiNzYSsUCieBqd70Blx2y0I+GeZqGRWbxbQHWKozR6jTJcONPnu0bUD2MPoWTeGRLXqX
EoEHWaUu3AXnS/7e8jlYtmLMvuGtLUsfq3+Ilng3/JqMpBJ+mFq6dDCFDmHk/zT4r7Oev3Wcx/pw
QQhOGjrfL5rHu4zxS0RCdB0nbQSwjkEB1yXakgHwQqyzgTmCwnixOv04accYuiJvGSvpALsvjDOR
E7a1+C22y5G4LCcL9lbiR9uRoXxovRu9YEd1SZ17g6Z4VHTJ7qUqGtnKVDczGi5E7mEISF7QUCQt
Uk/++/sDtYSsoLCcvrUGYClqqwbrxqETLeQ8UKCH8fOsudfl8aqs7KsmARflA6dVfVY24vmYI4CH
/i06sizyOWF+DjEej3rTpbIzDT8mrrwz/CvgRQnpmmzcVBRuNptQegQmnkti4jUArzne3MT4QHTo
RkuCj1Iqm3mG5c01LbKnbtiicC54QuxUJ84gkQ6cxb+d7+t7DEzbPGg0w2Hbb7X12ZqctzzsPFyR
gE7XxeIhDY6d3wQMXdDaSUwcSym5OSuy+v9SSccoanj+lqtlZ9bW0uUrhDO70lw2vLdu1FkQoSyB
jD1L7OK1ULkQhJlnHDkZ7Dkhf7eOetrwtvbk6w1ctVI9v/cyN2btq4m98jasobDsBqpC19OQl8aK
REAIGdtwijUcl6IyBuIBbHPQ6hvDn829zCzyyOzzrlGF44OKuKnOmd6gqeRtmg1/EBj+v2Xqqm7n
D7QqVPK0zNuFfN7X+kkjCfS4KGHpt9R3AxVD7m6+Yhsp6s7DE4s3krK/SavEEqsysvRwRUvq4V+w
I4Ctral9yo4sktKPlJy36sHm37Fmi8O9o6r4YvN/M7rPA6l4L0um7JzjTkI91AMt9YiOg6Ee8w+u
OG3FZW4p4EikR8dB4q/wmw1/OsTT4XdmolSZz841drkvZIe8MSOO1KM8KL6MCyVxU7yvnPxypN2A
cUXVenmDmGYH6BnNXBApRjewWZzN53r5FXpmY4ALYWyorJAl2QKlQc2QeZBSwzx46Otd1xQZqhHZ
qpMSP65hSL5jaDufCdF/7oFmRvjf7Sl0ammBRoam4lUjRIQQiymYd3zX2Lp5JB17/Es2IDHkzbGB
t68wjkcDyszhBz7g497Ek5tQjuxlcF17vzKslZW3I2b5DbnHswlyXzU3B7xAbfYKLNhHxnBeoVvi
ysXHJBs4VRF5BFc/0oeEkDayI4EYp/6Eatc84dFd8U4LGwUUlWiGL3uMKyOpVfXce8ipFlmNW20G
zOCVmY6xMVchi+vNzJ013yOq7PiXsWuvfCQQWTEIxv9gNg/je6A3kGgee7SKYSk0i18J0Sa8noOD
sX3ZQpbFQHAhyfFzmBlysaE5Gy3993o+OqqI7dV0C9mPgD0+QJfu9c2a5NVuN5c6744a8zrUG81V
BreO7PkleIYQz5MEb5bpqNQysm4Bjdlr8MGxwc/lQEnq8vQqp6WGS5N0BSFRVDkPhTaqZ1+VPuN5
REvfbKjeIiRQYyONbbzRNthPbdyHCeB2SXRkIMfJaCb7MTn+x6U0R5YKwktmHpyF09fwGbnS7O5I
RbZtqPbEPl7qkriihH7wSM63PTZ3hPzHEGGrxlBjKqRx9gx4ChrNa6XlXj1eoLee63KI0+xPFT/a
/9EPYyylGN1opHmzxi/Uii0tPVd+HnlSMv+Edoi/paukoucsHhKh5Z7Ceb1AOCueEZ4xHfRZh+sO
9vY4iUnruZcrH/0aF1U0mWnzCAhN6BifZfJdTSbZs5oiqrRvD5+HgWAWepPFwxIh1446bqhDxKau
hF2I9FeV4NJU2Ayh/550eQirimekJxu4SFxIxl8eyZMPLTqA5ApA3WsbH8LTdf8IhnQ2ATCn6YYR
yM4w4U+t3ycrl7d+H17BZmW6JeVLgUiBKQ6Nb6E8a9Np6qjpWx47QnILHf/Oxfy6wBYXqUjlFTkY
4A71dTiHHWzBzqUmK/W9EIo70lm87UHwsXkltip86hOC06CCcukaaaizA/rU4KQ+PE4rgSkEQ7iS
RZ3JS3YvEbu1LdQx2MpaEzqmmJwQaeskM/Hboa/MIt5kICoKRYHCHvuT91yFc0klnGsGuvpnA6kq
YNP9JhvztWzghhgwV9PVRocqHBCDUKB5hlxTlCehHm68pfB0UgWCK9dQhPtORjjHiNHHmuQrEuHR
3p/6+7glAk+wVFvV8QvcJ6BAoeioZXMDxWzxxzNCm6Cjvqfc6EtU9BCpv912mlv2TmcpwZUBXHZl
mmIdUg2m8uZeCU/RbJifO1RYCQZWOoff203RgeeJ2+J9E31C/9hl6teDNa20OlNXAHXC1kDzNkcJ
CtUDOfZK93vQAav4a47viqd171pic6H4lMvS/F7IDPGu+FzQNSTjWnlLBKkXwTzJDWJ3UBMr++Hl
CLsGbI4gM+f7rTP33/sBcXCzzhB2dzNrAjZhSGMAc8wpyOSkYX1nCtqfMKhnYl7H29fFFdISMNBB
EAu8dQ+YxZKZtkXa0FFAC0XZGvfAc3venCE5iGpyN3hfzN41wh84t3b3Y2FhcMo3oNmZZT+HRQe5
2lQSrfE5tjDJiYBK54QjBX1doMGwFFAQrbtEZWP994bM+9cHzkZc4jo7d3jybLH6lPaXExbGLDaE
qMrQYn/tYMs1IawfVECZNHvdXkiD6sDiGO0k5Ibg9bsYzOacgLYxF5QwzT+96mevjb8kZnbX7ivJ
266XnrIpBsKQWMeOyWXdXnfGA68f1MkiD6PBU++9+A/3V5iktJR7obrESlra1PNUBPfwKCggZuF+
xx5Hsp6MMyVRqdcS34wMFfQUFSsFv0L6Y3FmyWxJ8ceqsGoUKi7mNWvzlD08zAwbBgOqNsqNZKIh
qPIpqkilQf47HFGXVf5XMP+VXaYN+91e4Dc4tIWWCE8QG1P0arjIs96TSJiE9R3zzuZOQm3GMOMl
7GOnLDxo94qCkI3ANBDS8gxs1Tr3SfZ8LGV6bmLJaFHwegz1ifA+GzAQBM+OlfYtv1cGTERcUbCB
o/oBB4OKOMLUvQtDZ9M6aZUhK905ci5OZ/usLMkwjLFRp1LPH1EQFjIwwyDm3Pl7l0slPbOkKJAJ
Rp7MI4JS/cs2/mFs/WZ+wZcZpOskyz/z+GoYJnWnOvMAZlh0hivHHea5RIsf18lSSVTLa2xPBVL4
70eIkWhDiIdyr70DOrj5UPEIiO14iSklBPj0YMXvNWpxDGnm41cYosAZ3PAu2AvfggtskUqjFqrV
a8mFfNoZu1JEaa/U03vqD6b9VYwucUjE5zLXykwpbYjFNZ87psnwF7qtYGhCcsDawUPgYDloCjYe
7K8DbCOj3QDprQUz/BKz8rZRNuQHU7uqnS+sh81mc+w2BcZ3A/jT/Z7EWoxbTGcGYSpwpQZ3uCAo
Nz2MZcU+0eu2dB/Kue7DsUIOGeJX6UoJtD6DzvQj9WF5FU8gUKwmo8vwpzWN4pKOHmzJeVSnD1Rw
YIt7QjbUl3RUoWJSMCoeZgGjBbqA1pjBmtoQsgCvdIyGupTXKe9GxI+rqIYB4jHRE/J0e0qLSmNz
UR38Ot4AFiYaXKfih/T5DNsKsywZHOo3B75uKVP3bqp+dF55ua8lcfL8E2rigJfe6za152cl6dcU
1b+m5UaT7OAsBUZvsjWvWVl5oRk2T7Ls4kQ8hkBlpNUCQp9B3y7CCuhKhqqsz3rQ6gA0CEk9UhE6
RIsUc5TQcVVyOi8+iRU0BggQ7bpAKuuQFjtlXSwW2snkTSXCiO2hKmSRD5WUFQ==
`protect end_protected
