XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�jْ�����1�t�S��*}-�?Wr2x������	XH�a�)�^�z���Y��҉��ae�咵�h&ɛ(�[b�_�h`Pt�F	�E��>ŒK��ȍ��>�r�~�樨ŧƂ�gz��TR�Ѿ��������:��be��C��f
��=L�nGv�mC���c��7��2�v��c50ӷ�j� �	V�����S/7?��d��A%4��̕9�b��F��(p:��m�I��d����67̊�ȋ$�
x4���&嘿b��ye��3���}z�9��>�>�DK5���;���^"t�E̽�J s,�yf����O\�v ��0j.�9O��|����E�W�3>@�W��Sb����Ci�Qc��D��Y�3	k���}FP٦Ԃ�W�^[%�i���I�eAZu�U
�Kx��y�jߒ�1%�2|UO����	��"g&����fR���X��6�-̢\� }mCU��ä���mO�0��i���X�w��^��"N�`�·u[1=y-0���w����L���j]����R�<�5w�ˌ:.��AS���m�ʚ�����+++=�m��ڿ��h��#�*p�����$�O������uc�u/���UV'Y��Hd�'���G��~�$�{#SR�Z�:"'&���=� 13�פ�)��=L�h��Z�&:
<?\��A��FRr����ղ���d>14x�y��=QO��'�0q�m"UP���p�L�ڏ���NgXlxVHYEB     400     220�\�t0㈢��ٷ�Q�6�@�sq��V5i�	a"��b̘	�����~�q(�y��҈a0jI}��?|k���a���UWl�2�\�XQ�O�12�V-�s9Q���}d�:1F�#����l��������M��[�s(xR*`
e�)fS]y�������r�"ܻw������Kv d'��֑��h��<�޵��I3.���J��˵�»��gG;r�#�I.#}[4~/�-|bO�q���_!��H:Zw�rI`Ԅ'�2�?�6)��E\L��Ox	���alSW���8��[U�a�e�(_h�(î���ḣx3; �	F���g#I7���uT`�F�{��+��Cܓo�}�)S+�	5^�UQ��j�4��'`'beB�m�R�	�G�]��Dț���(���������z�QB�t�x6�J�#�Փ����3f���/@����a'��]�83i�O��%[�w����P�C����n�*���7*�3n��j���!~�K��$Y��z���y���~�Z�A�XlxVHYEB     400     220�j�7VH���?��A�$�j�����J�,ZI ywq?�B���E@<(��S�wޏ��� T����n���I�w�h��f9�n��A���$f��>}��+��"�b^��lb�Fn���5c���kF���!4�XP�׫����0>�F�y�d���	��6I��n��w$[�D�g�����б(�g��W�xt�{��ie�l��Z��O�FGsOysx��l��JV�I�8l�N'��n�c���
�lAb*ڴ�߸�IM2�T�3�\��RN7R���|-�l6�C`M;S�4� �;��{$b#�{���D�Ξ��|�U��]��c��g4�v0��k���"�ǎ���V�x͝��K�\-9 ]\>]^��Ry�f�c�c�����`�E�`2�)r��� ���<�|k��!Zj�ܶ���?��# `���������U�U�\��F�@���QjQ-|_�_�#Ȍ��g��ݜ�=ÒNx
)ǣS.X\�4�MR�YL��!#���催�G2����[�m�'XlxVHYEB     400     1a0�"�hA�</��B���S4رC���#��nu�:�� p(;�q���Q����òAO�v��:��䁽3�f�H��$w_��Mp�͑���xD1amb Ɨ�����X�[�4Bt�����w�J���Ο_I=���ޤտ���ȇe�+������̠������~+1լu���(�t���bơot8��v@7��@L��KxX���.�<�;j�'�p�J�R�M���� (����2v2/ �"VAGؘ|��Y�I�8�&� &p������#�9IWAX�`	"zT���v2�E�Ѽ�ն�<���c������CX.U��UQ�/�{�>���[Ãx����i[S�=	lB��*�����0��A���)d3��I�;㷼��b�*�@�XlxVHYEB     400     130��l��*�zs:����Nf�C�*}���7���gK>�(X��V�D��B)/l28��o�K�ϡ��R��6����ơw�����,��"�$T`D�}�T�<������"=��-��X���1C
�vnE^��M��0M�Ϸ�
�.ԋqō��C�c�[@�C��N��9���%3P��PwN������3�1u��Ct2VIĊ*։�+j,իK1e�F���pĪ��c||1�{
�k��F�*�,��N���X�w3���r�3坣�^PW�����k:d2 z�+R��=_�?��R�.Eė��W�p0?XlxVHYEB     400     140��W�ɲ0�3Z��~���R�6W:��
��l�:��r�@꨽� ���z�i�`� �Q܊ܹ*��Qݵ2�Id#��g+*�$��qb�^������\��$3{s�u��
 ���A�ٶ���&��%�z-�rRn�Cp C�H�XY��c,�v`�x$�!�ƪ�8�V�N��7�oV|��=��z�?�)��|�u�փ49��Ƕ��Ϙ�����/|�?u��;��w�Mb�w�_&0��aѤ��Goo{��P@��u�C�7��h����}����P �A��F����Ts�mO�;@b>����`��*�V�XlxVHYEB     400     1c0����;���(g}l_�X��hT8A�;�ݪF�EE�tT-�=����Ux_rӐ�������Y����~W�m�����%�ﲡ?Դx��|��Փ��y�-��~T|�T��Q�Q�SM&����I��	��p8�g~=��:��7��euR��MZ������^Ƀo����N>���B��L�.�jq��}���m��~��4���B�?���}ag�*��A�SM���޷ۿ�!��C�S����t`&#�H��*�B����ʂ%ԅ����	t3��p�ߺZ8p��w�7�^Q^�a��fh9
U���zT=߄�.��9�B���c���t��N��ӛ�T|."$�։��O���.�T/�"�.H'�8�����5�Tz�07�j��&��R�����YL�:��M�*�Tb������ԾA�� �f�����Yb	��GGݍ�XlxVHYEB     400     200�y3��6��rK||d���Q��g�J�)���R����vTb8I�W2���ʷ�߀����[Ս���_��4�}�c�>�cZ��ką�L1�3���'7N)������62�3�)�2~A*��'���7-����Q��3גÖ�^�i=Ȏ�vY@� (�P�㦩�~#N�-,1�'"�[k1f�ٰ�Zd�@�{,j�Y1��,��'�yC�
�aGYcmW${�zgTG�G����*�]�:��Qy�C�q���H�:!�q 1p���\:�_\�R�)�gr*�c\ s
�gZE�vS�x��%4r���	
:� ��r�NZg\Y�� +�%��ӨO7��N��)�O��c~_�;�9���y,͑w�v�v#w�0.:_����Xפ �]}�[f����߉6P��vt��w%�X���u4��< ���C�4�[��jڦH]o�[��#�l�Ks{�}�l]�=��"�_�S�&�u[!1_�p��P._��M�AX�XlxVHYEB     400     1f0�CMY��7��w ��J_=��!6����=ͦ��98��ź)i�֔��%��]��e�eZ�tH��Ct���8"_��������mK|}�[��xDw�v�D n������_|\���ì����@!����S��<��D�j�hL�h�ֹM����&eZ��+��"7���Y� /�_�뢯'}�c�S����Լ�/�jG���S�衖� 1pkǦY���	�᫼�~�����R���wZ�m�����ĉ�Oy�p6
�͉ެ�'�����̹g�d������"�R��	�ˈBd�[Q�;q�m�l�Q���?^`�?|�X3�<�Q?d�I�<��ae��z�z�b��fH��_ʝ��*�]q�s�]oކ��A0���}�=��+��G� ò����_[�t�>\�����vAI�K�^�LL�Ss�0w���7�Y�7X+�c~It)XX,��M����~��{��4����v IJt#�7�xXlxVHYEB     400     1e0&��1>p��L�I ���,ՠ;8�qǺ����繛|@m4<����j�h[�nz���Q�R7"�yИ2�a��Y��u����\dh������1��[~h)ˊ%�O)��T=�'G���/,O_�QTX��+Gc�{tTC$ ����m���;Mc�x[k�vA<�x���@�BD�{,Aڡ�� h2�1x
�ƈ�0��#ztߛy��˂o��5e��I��Ptj�G����#d��q��+�WZ���h���YS��V�Y#�~̗`�.v��M3�!�:��M@�����ѓA\���XVܘH	}�X�ۗSV
Ͻ��Z?Ѹ��~]�Təs�|�[�񇃊 �e~r��k��Pp�j3ӹ���!S�	q�� @��[i�e)�'�q-d����/$E�����Nb���2/��k�-{�y���N>�&ʫ6*+:�T؂��uۘ>�.��W`�lM�tC�O����Z�
߹�߱�� �1k�G�vXlxVHYEB     400     1c0��7ŬCh�0�DZ��2�|hO����,4��:E�������ׁ���dH��,�8�VX����B�'c�)u�I8�鎓��9t4���7-%����i��m�zC�0������С�/���м�pm�ӝ�)��!���6M���'���oҠI��>=�9~���j���"��Vy炍�jl�39��PI�����Zt�F�p��L����O����e`E��eX'������|�&���gp����K7���\ڛǡ ���c��/�8�%X�I(��V��u�GPи^1��$(����;n�&����E�q�|X������8/m"s ��s4��@P�B:�YT���S+'4�w����Y�]fm����_�:	š���{1�+u��N��B�2"�?�۰j�c�s3oN.��"���.{*O���2fq�d2;XlxVHYEB     400     130Ӗզ�6e��V"���Z�1���&/�u��0�".%!YZ�hPf�!�,�5��C�H�mqR�+�/�\H�bo�e�=��0éc�ܟn0�Reh$==7��2A��'�ulZd�o�F�3�_'�؆+v��D��vz*�h
3�讑xr���N�9��{۠؁��[�����` vp ֟�w��=֥K��g\.L����ٔh�����)��G�H�n�`>��Z3P�m�j�L|lr�Έ$~{�H���_hN_��v>�N��{���͑�0Ɵq���^�T2�gN�'&BF�As��i��܁�ZXlxVHYEB     400     170��]�s�2	y�(���E;2������9�-�H�#�����JY����4M�\�&ד6y��8��� �1�6<�)̃��#@�˗@�;G �8>\b3�t�f�L�? �+�����Z�;�K� &�a0�%r���Nܚ�ܴ�`ۜt˗%oA�TQ�M5�B@zp2��'۟� �FA��L7�U�	;R��<w�/q��A�Mpzn,n��%j��-�C�6u��}m�rt�!9��Pܵ�o�`"8�a�s����8�8�1Z�2��{`!O7�#|���y�0�j���
)���5�� ��C N�f�yma��W$�,F�q�8��2F5y�ꤶގ�\�p�{�?v���
���b��=ַ�fXlxVHYEB     400     110��(�lzԭ��<_U��<)���"xI
ŇX.�i��N:E���}|�����E�y� ��gZ�X��,ɩL�5���������`Ģ�����_H.��5ua%!ӦZ�h��9TѾZ�W���(���2o�Z&,u��퇰�&�a����7����d'��ٷ� _-����D<UҮ���DQ��n�$�i&�?W\�HB#Ŷ����rq���6��ʊP&��a��,��n��9���B��f���
v^+W�,��`�@���?�ĮE��	�/K�XlxVHYEB     400     140�ʊ
�6|l��<t: 9oN���>�i.�n��1KZҧ�;!O�{�̊ނ8�!�!���^��#j��`x���~�}ׯ�wB���,_Q�˦@\�t��>//�!�}���h`��qٽ"��M/�;"�k�01²�! \[ۼ��t���߁Y,ee�9P胀��gW�TW�-�U�gr@�vj��#�J����"���5l�.�#��O&:��0�D!q�F0_�����nbTy����\����W��z4��&�2�������G�?`��н���b�Ws��\��D�q>4�p#��.Q-_����<��zXlxVHYEB     400     130��
����!��j�c�+B�B"A��T.��X�Ztǈ�	�GX��O����уA���{�s��8�B�]�<��s���-w ���8A�Gy���g9,�k�%�Rw���_��	d� @��_ ~2���Gj'��.�QS���yb�J���ŭA�V�_VT����ϰ$լ��a�w{I�%����i[������=���jJ-8�������e(�+6�Y��Y�܈˭*W�! ��~:u�����G�ّ`U��Gf��$
�7s �C��8	��&(���Y�R��DXlxVHYEB     400     130ex�`E���@h�+������
�/��$XT�C��-��c��8���a6�T�O�L�`2A��zL�Aof*����j��$Wg�1boȣ��{g�Og������ .�d�<٤I��[�����>v@���#�2/��P��](pv�|�'s>���o3`<B�N�7�8�m�5� �e	���ܝߌ;� K �4�]-��b��3"� R��b4�k�wqINC�� [�8fT�9���r��>H�\��q�p?L9e(�Y�c��W���}�6�uPT;�t��VEf5N5XlxVHYEB     400     1509&���rO&��Lh���V�҈غ����$���^,!_�}M����j�R_�v���wSH����[�)���}�ѳ0��?i�_\�>�E쓚ge|��z�P�C�!�
��m��`ڹ��}C�KE�w�^��H�h&���T�*��j�ꑋâ	��U�L]\�b��s���Ne������I��)܅R��װLQ[|8	vR��5��|i�EL���@Y��5&28��v�u�n��`?1]���D���j�Z'f��"pt(|' r��en���K�r�~�ߺO�� �z[.�6�C�,^{����E���;�o��l�9�<�1��XlxVHYEB     400     1801��kBab�Z`��u��j��-���<�l������ԋ�[���&BW �!|���jo��vv�W>�K?�+4LϾF`I�41\�k�g3�;��Y�_�_f�3�/L}�,䄅-͝��W^����]�6Y4���r*�I����n{[�����:���[�'�4���O�l.�T7D�uU��U��OC�}��#k�c�|Ut�FN�<�i�¹��=���$�]�Gq���=�R$K��?��N6X��H�@�Z�z���&��(�3����΋�v~,�OaO���/{X�2U{b��c�Ѽ����'�Qխz��w���R�8osFc��HҦ�"����X�F~J�C�3A8K�
<eE�)��)���gXlxVHYEB     400     1d0����S�-έޛZp!#6��fO<f:�S��<�xx�Ÿ�CQ$�tH�%(��5M;����n����a��5���G˽�d��S����:�|�0�">I����K����`�����Z��>;.�O
�ՔRWN�޴P4�>�㽙L{\~�����$����o��\߆��H�UJ�����QX$�+����=�gM�P׆]���{�=)�7�yu�dTe��q�(?����������i�A�� +���J�&9k�(r�8�I[�h��:�+�-	
�ɖ��?K�P��!u��G�{���}�c 4���&�pt��I#�
`q4�T1�O��;@�'/�������]�H3��(����?�8VM�N�a�������T���t�Ɓ���B�4ߖ�����ΒɦR��@Ȱ�=�hhmU��,>�W*���ͥp�� ���PV��+�������0��`�M>ֵ!)XlxVHYEB     400     180c��L�\Vc��3��a�o�����h=�/�^@�G��J�����-iH3@2�������蘿�F��>��
�Rوk�����4�*��,V�VV���R[���q�}����Od��<��vڱ�,��]�����ur�Ŭh���Z�O��� ��Zƞ�a�J&X�ؘae���-�ķxL}��T͕������\C��O8icI��o��Q����xv��\۠`��Y��	M���B��7|�_�O��O���+�K)�wo̩����U�.���ԇ��ۂg����"At��3�/��:�e'}�] ;�u{�g!���"��A�mŖ�ZA�%��5�Ŗ�jW�.O���U�1E !�[�����P"���������Qo����YXlxVHYEB     400     150]�<��� ���Oz��R���Q�m!���2!�٩�VG���,Nx�I�U��6/2W�� �ҳZ��a�6g�l��w(
� �]T��$SM���<��-6%rCG���o��*�j׹���
7��{��SFΫbC��մ������~��B[4��u��12V�*9)r��[�p>\�D�ح�>>�Ҡ�_��}z�p��o%�g�ˢD��صl���#���\:�����JI��
�8� ��gh�2�m����M�dXH=d1�q��#�vN
��=4�[��v�<;��}��Bb^��M�`{�dܺX���=]d)�W�I@��XlxVHYEB     400     1f0 sf��uI�L�A����c%�q��*2�z��ܐ�Z&��t��F	�_]Y�)���s�xr��!"Ӥ��W����ֲ��]du���d�Cml?��@~�t8��\���=ƴ�h�Ow��4��.G/�7nC�=qb�.gx�,�~�CW����W=�!x�ܗ���)���?˩�P�ʌ�м�����~ƽC6�<���ݘ_�n��c���3�~���\|X�=���H+|i�_�kg� y)�W��������;�7VO����b�y���a��Jf�.ͧM}s�>�*I{Ȥ�^�򿓷?�-6�.�9Q!�>I����|ŻX2Lc���(��*Ɏ:��f����j��~.�����q^�&�֙��wn*1��A�8x���ܪe���XL�˽aw8Ɩӛ�^�r��͞:vV�Leh��"r�,PC�HV�Y��o]�$�J��4�e�Ȏ�^�qJД�#]��x��߇Q%C����v��XlxVHYEB     400     190����r�&���n�y$�nt�%��Mؿ@��3>/q�7�id���=�Ye1�q�O����-}��A�/a׳�l���ApB�k(����B��#�`�$�6Ԩ��5@+G]'V��A����W���;�����g�<��=�����p�tnf��� �+�;L�OК��dL�y?M��&9��IP��$WBjI�:���JNa��6V�pw�����v,'k���`�f�z?��υ߱���=��Mc=�g>�@��\��a˞e `��fy��G~O�8�bz����Jz�Z�gm �ˣ���;�:3ZU������ybT�k&K��AZ�z�ރ~�}3"��R�;T3ڗ��Q�#r��P��*��ǅ���'��m3���d$�_X+�����{����T�kyNF>XlxVHYEB     400     170���VU���KvM� �e�'�JXޤ��$u�o�T{-�p���f6��u�ctc�H�NH��� �MAK��,�l
��ډ��C"�4H�L�o�4��|Rn���O������l��6�q��p��d� �����1^砎����ֹ�b�Ͻ�����i�?�����~��; �tβq��r�w�ۏ(�� UE��۫�ZR�/�b��(Y�ck��!�����n�O�1�#L������Ř���W�`��æ�-���-�^���"��M{0=?�,�K���d���uƾ�9G'��4�;��
L**eٔ���W��t�*�k�	�!�S�s�� ���~�eyQ�׌9���8w*J	�x�XlxVHYEB     400     170���,PF7×�K��֭��I���ѷ�ʛ'��	�
'����RU ��ml3KLHٛ{��AR;��{�#��)��"��
�r��lG�X��f�~����kÐ�O�D���_L��7N?n_��C#'�kgaD�c��!����n��}#~:_�C �pN���ݴ�6�ʛ.�>�U�J���7��е��9W�+;��?��ņ��6$z+����47M�k|�m �j���p��u���EN(���F���W��k���or�u�����O��ՕO{�VD���l�㉼�JA�y����k-D��MT��dGN�}`�jʂ#���g���ݬ��B4��0�m��^`m/���j in\�dg[	XlxVHYEB     400     110!)2��R�
@!��!�[��������Bf�%��{�s�3?hDِ��6Z�B�($�k�V��:��<��j��.��pL�a���\~J�O�n7W�ױv�kR�0����	�V,��-��s�K�Z��;�8խ���:�`�am.v6�uF\�"� �u���#ۘfO�_F��#��n��������颙�b�sё�M3�5��sz0�\��n]_����ŏ/Q)�z;S�O_��xz	{6�R��*����:�Μ�W��n�XlxVHYEB     400     120Aw�npcF]I�W�����$Ɉ>HU�,��4�D��+��u�T��ݗ0�,b[x89��Y2H�)�^ۛ;wOg��\��q�SP8w�\%[��SK�wk�჻0œ��+�k%~���:q%(���vm# xt�:U�ƚ���1HS"v֛�
Xn� ��f�dyPC�&O��?п��/�n�0��G��0�%ei���r�еo~�Rn�]%�eEe��W�>��������:**�MUG����W��F��7�(����W��	��6��;7_��l׀���JS�XlxVHYEB     400      d0��*�c��'}��6������c�z(�k��I�~�����y�����1l�B��uK̢�C�9�N� �M�):7c�����I��	ʹ��5��  �*t��S,Jw��0�\$ky�7���*=��~PF4U�����ae̐D�I���T+���:j�����3o�!����U��E�F�����L�' ��W�3���F�08dXlxVHYEB     400     140u�X�0ҵV�J�<�Z�u�v�,�P�8S*�`��㺕H�.�e&g�ʕ2��̒k4~4x7<8nS �f9T�$���.|�
gRjK��7!��xs��������v��Gv�h��dJV�f2��n49�YB)��DR�����E��l��u��BaU���X_��gδPqФ�c\�3�0�TҞ�C'��S�m�
XD�r�ۇa�Ţ7�L� xI;�;��?D��,o�v����ĭ�i�JZe�{dg�9��ښ�t�3;YM^j�q]qf`�����A�k��
T�2�F�����
�Ns`�Qɧ�XlxVHYEB     400     140j�d^Q���5DYUt��B�dD=�;`G�7!�,K[�4��Yy}b{h�y��R�Ț�{�B�ѝT�t.�QS�r� �����\�K�=�"�p�`m�r������.
��b�r�Y�9!�\���D9��!��^�(7<;��0��v��^߰�+�O�43���%��b�E�U�4S�(�.�q�{���$��H�v��j�AI7��7��OU�{�r�Y�ӺN�03�.�̚ΐ�h��:� G��2�ؖ�i_TM��b�EU��V���P�y��������d����J�Wc�B�/o����'�K+eHu�@v�B�uG��5�@�0��qqXlxVHYEB     400     120{Dkv��;���$��]�IlK���(�OLW��'p�<ʱ�,�[��o|Ѷ��p�;y�!�A��fm��0ԾW�Ώ�_��kM��z)��i���wFy��O���ch�@�
��&��E���PЬN��*�Sw�uE�Sr�e0�z�6�Y3�ñ�o��8�8�H�'��j�D��/�(c�h���z19ӓ�ૄ�����}I�7U	�u�&��v�-��f�t��zzվ6V"u�RR�{H��s
i��ͯP�L%��	R0����=L	n���\V��'�sXlxVHYEB     400     1a09壷<r�3#�n���<���G��,�j���)��Z�Rd���KU	�1�$���a_:�N���L��;�J��o�Q�V��>tw7�{���3��IP"��;'$ˍ�X\��Q���!3�~V�R����b�S,�������,�4L�(0V$�1��6ph��	?�E��#e��+����'��7�:!	"u[k��p�%:��x�"��F.�&�|�N�da#�6�Dǟ���o.E����=�c}������ϝ��$��=U�M���M��cu<�?�T����d�zgR��>��~'U�҃*���ۻ�����T�rB�)h�=P�.ܙ��𘀴j�㯻��?�b-/����q����|���,�=Cͺ��Mκ�>u �K����v��3{XlxVHYEB     400     120Z�d]���'�J��K���m��>Q��C�̾K�p���s��G�I�Z��M�@Z#z��N�b�Ql�x����IЎ����^���j�8�T�n����V�W��4eŊį����;� ���/��
����tҞD�V:7�y�Viv����x�NzJ�y�!9RjcfI�/0U�ur���
�d�Fz��9�Xec�&����c(�J�-5�M�mրb�i��gg/��1���V����HOx���S`D>p����޴sr*Oe����#M܍��J���L���d�䟦XlxVHYEB     400     180c����E�� �Y,�wwK�Fº�Ʈ���S�B�m������QQ�7w�9�:�=��[ۥ\�F(�Ȫ��(��~��ъ�.�-�(�X���.M'��'�ۏTzտ.-���I~�g����yi����SfѨ�d��Y��|�(Jk��
ռ��n7��15��q>��I�^Wi��nG����ZNʣM��S_t^���X��Y�0Dԛ�	��.~��6���Of����Xt�S�]b_�؋5���"Ea{����'.L#��<<���8���"��t����'�|��:��2��tSG$���/�LF�B�X�����\Q�De�Cv�B��x��f(���������嵣� 1�g� �-="y%X+y�����XlxVHYEB     400     170�j����Z�jz���j ����5L���7�O����6�K<�̿�
�s���^s�b��w��o�{��ǣMoj�ܿY�-f ȫś�=׀&h���?����co�:���S\�әU���l^�o��B�O�송69���i���8X+��*�L&���b��9�L��%�h�a�gi�-�M���B(؂�K��%/j�or��7�s�Nѹ -!>4���k �3bT$��z��T���7+�zޓ�/V�MoS5A��ͻ0��m������Ma��=��̞d����a
���\T�a�Bn�Q��2�:n�Ϭ�>���4���,�!XP�/�v��p��rޓ8�涏�\�c�M}(NXlxVHYEB     400     1c0G9�+�̲g�|1��q�cH�w�^������/G��������yk #���{�9�da�u/�Ǎ2K���.�m��Rq���f4��,(c.oГa��J1kU@����>�木�30��Ѹ0T˟D8�K������)�a�
~�].\�	3���%�uv�L��0
(H������6�.����iY�h�Ml���%�d�Q��{�PYuL���d3���XҺam��V��n�4�X"�ZE����g��?
��R)nN.u\3�����`��.͠��Q�Ҧ98X��]Ԕ���F��1�HI`̙��}�²]�m�D�b�}#=w� !T�R�^28�Y�d�Z�<��/qF��<Yx)EsrL�M�P(9: ����1������S�����Nן�.8bk��	BK��]иK�0�w���Z�렱�9=���
x����+<�UK3XlxVHYEB     400     110,=�� �I�D��J��ʊ�vY��]�#��z�A�Ⱦ�>�Pi|T\�&[���\g,gM=�����&�YF`�ѯ�J�9��[-�#}xRh;W^��|�G ���|���I]�.��<4�CZ�����Kv
���F��N�#�:m�9�0�{b0=m��ݸ�vM
���"�*s�� �Q0�϶[��A�cf���Rׯ�Q���%k����a��V��?0�
`��`� ��_�Hvx���̨�<d�*%�g*�@��*r1�vqo�XlxVHYEB     400     170!�@鲘`��/��#,�� *��\�-�*<�����B�wz	P�8䷓V\��mh���Ĕ���l*�;AΦ&TK����3i"��ju8�B<r��A:g�BW�"wz�h&�K�^���H�G%ރ���n��<�/�a�s-%���5�K
S�������[ڽ�T갖�؍��`@z󮁯q(�� |<f���첺X�΂���0�MԜH�j�Qw���4
i-N��y��������^sՖ@�߄Y��V8~��������K����O=ء��_B��9v<�T�B�p���P-/��}CL�/��DY�	�=I��߈V�*�V��g�(m�o��q��]�BW2����=����8dXlxVHYEB     400     170Y]�����ZPq<	� G,��Q�$�F"�*���YP:5�w���A��n�T�m�St�������+{4鏤��#=gYa�ؙ���)�W�G|�`t_��R��e5��������E���w���}�G�Vw�b����"T\���]�V߻�3�9d?��]��#A���dc�ӧ�_u�wg������YS̜�wEЩ�l�lc�/��щm�9N���Hd	����t���O�4V�����^�?�Mc�kS����� ���,�m*�K�E�l	�%�P�,*�k��K�-O�&���(�,��&�YP��bh�ưL��Ƚ�l��?�WMe�v�%�iu�^�O���m2���c���CXlxVHYEB     400     190�H,�iH|��G>�����$�O�;L��:�E�@{��b�_��'�#̼N�Y����R+�Oh������i��$y��0�`�cg ]��P"��2K��!K'�3�Wy4M��@�x�F|dZ��ּ=5��=9O��&lx�c��������Ξ��eŔ�V���x�K�v�m��}������!D\G
>Y����2SN������B�g �e����:yo����J�✩r!�2�NEJ�H��BN�)��ǭ��.��tR��+�FΝQw���H�K��=��C3-'�F�$\J�[���~B���^J@�mуɬ���&[��j�S��R�$��|�T�[Ԇ`ԃڜ���q���������P"*��aʞK4?��L&7�%�b�������>XlxVHYEB     400     1b0�젝�K�q,r)�3�fĥnũ�ۣ<�'�by��%�12�^���N���)�0��-Q����ţ�h���Ƴ:V�[
��Ύ�Fd�ED�7�p���)=�f�����OG����6g���Rua]fj�7.#���h�X�)���|�ޚL 	���St+�.G&a���h9c�P����:
�U���}�Wv	y��^FV$fEР,q�%
(p�C^H��w���'�������>Y
z��5��EN����E�Iq�h����l|㟂ˮ�}�z!���Q�Pm�/ u<N`(r}�̥:�aflAi���#.���f���7I�d�%ː������&�,v�@?����yW{��Y��%�*r�d͵�#�e2	^�M}�󉮔<�A^���
�@�ЗN�m2�.^Oz}�GA�ל�0�S���i�ОП��~XlxVHYEB     400     1b0��*���l��>���Q؍%����I�'�9n8D���v�<�1�q�nD�'���n��wX$�q�L�<_"�hX�^%�����H��*Yyj��#&���S&/�"�Q|@�۪i�z�?mE����ַvgx��l��nQ�o�߶T����yx��PG�]�o��}X,�=���%��U���,�{ ��$_�������6�����	�k�W���x�xsH��a��G�/+�n~��L/kq�^����F�O�*��.i2��Q�g�ɂ$��w��cғ=����R/T�P�][�s�-��l#o7��(B�}�Y@�����tg%Q�?@�FNo��pQ	O��������A�ᒟ;�A�4�{J��fk޷)�,��S�vo���( 
N��ka�֫^gc�]}Re���bt������O��p�i�%[�XlxVHYEB     400     1c0���E� ��<ʝ���,��z���Vg�g���N�	��
�,�B̉���#nqa9��N` `BP���/t��_����g��X]�}(��(p�ךl�=Y5�S�Qǜ�i���3�t��<�$�ٮ��4A�6oR:e��uA��~ur��Q���İG��B=�H"�_N��zivr���{4a��H5�Uo�2�@��V�c��d�����W�#�Z��Ԙp�_u�	l�.r$8%�\�����_z��kX�:>,�l�ˤ� !��}��=A��U�3+�í���'�2�3�`k���4]���m����r��t�K�3A��s�=��V�w��)#��d�M�R�&	/K^)��ȾϿ��e��@\�{��p�	6�k@[E#rՁp��dk󬷝fr��e^DN�C��m��¦���c�=Mu�ܜפ}ÅA�jqf�sԊXlxVHYEB     400     140���.��=��&h��>.y�q|��x|Eد���"�vW���OA��*�������GMH�u�(�:�i~��C����q�!��
��/�����p8W�5�KnR@�Ǳb��6�e��bwy�c]z?�ҌH7�3�嬍q�2_�R���Q[�F����x�L'!5_�bDdd�R,���? ���+!���;��R�l�';���E��l�
�U�W�B�L*�#(R�8��*U�9�:{��TDr�%�/��Gb���u�e���������Q�6��F.�F�	G9O����/TY�&��l�q��T�v�nB\7���Kʤ�hXlxVHYEB     400     190��2���h�D����Օ�ػ�4�WTڔL���(ϴ�ӈA�����I�ߞ�G��p�D�:��Y�/0�!�J���
p�v��2lK_)� �
�򬭜����>��D��ճ��ǜ4.��j0����^��y��=Ig�+;��]������͑i�����e��8R��or˱����k!2-yRdq��͈��Dv�V�����ͅ���4�?�pj�M-�1��4��ul�y
[c�K�� x�B�/��beiQ�I:�y2T�jz�p�=S�/�� @ n(������l��ȴ�Ў�n���P"~Wmm��G��ʰd)�R���%Y?. ��X|�g����T	Qvs���~����K�	a#�`�+]�R��h&�)��7*ᳬ����5��~�XlxVHYEB     400     130`�a��jt�o�wDr�N��!��Z7r������:�F����k�GUف��ro�����^ؽ���e?ۯ�'`�ƾuZMb�����B<�iu�%�[�}QZ����2���Z>[Bz��(ܾ��|�w�7��w7B�9��~ߧ �����Tf�
��Pb�/��k�5���!� o��m~%�X+�7��G�/�05W� 9�\�m9B�>�}�O�l��ҤY]P�R5�byf�~ӣ�y)���E���<����K+�̀�3���Ӌ�W�i	5K����nZ����\_@`QXlxVHYEB     400     150��AX�D��^��@��D!��;k�E�)�-"u���5MQ���9����ug*�b=\Y��7�XǤ5,�	�i �]�0��n�2��l7N]�������P��SÌ�w<)0�W#(ln9���2욞��B��iO��ēA�r�{��?s�`c���:e�2sza�Ԫ������u/PL�}��>[U�V�рtO36���5l�嫬���� ���F�A�}���J��EJ���(s��oMS�����!�Ȳ1"�sk+��I
jGm���c�:�{J�"q�Iږ̬Q~�Pl֟dCҮg��n ��32t�c�X^,���-��3��4��Y�[=�XlxVHYEB     400     190FLV��y�3�i\驪NΡD�bK�?�r=�%H�
	Է����{�o��#i�'d��
��o���&�ݟ��j�K^�7��T4���Z����>�yڄJ'U�IHqk������*�5��<�)�Jn	� ~����IQ$*���� �V�O�q�HS?�Y���8�Gw��QQ��#��2�N�b(�ϣ�J�E�7�/Ŀ�(#ݭ1%��c���x����"<���1f��C�Q^��ҭ>�Op�rR���t�����h�z���`kk_�z��mP�����%5����^�S�d_xW��z?i�j4va;��,���/�1'������;0���j����U�FBX��c$U�!�0�U ��Ӝ��|��\�����$4��d [gM4��	��h��̘�Z�XlxVHYEB     400     130��g����N���hd�{b��d�~�}��_4��ٟ�k�3+2ݛ�'��-���U�J�]��]|�i�����Q|V�|{�P�<5�T�ڽ���7�zA��-���������(/�����!68��l��-�ܫ�a�����\F�1�a�n�mS(�Y��r3d��Y1�p��U��gm���D�	T:Q#Ζ�������s���Ho�}��n-l�(Sp?��&w0��bӾ�N�:� �{�s��:� F����'A�;�n�w�=�˭C-��U�ťݥnA����XlxVHYEB     400     150u�#8���aJ�u�	vآ:z�_��)�P�6���޹w��U������ɋ�U1�l��r�:�!�[ٮ�����Ħ������+z��w�$ҕVs)�!�2m?o���It^ؕK{��q&��v�ݧ~"����e!F6`0j��x6-[F���G�"]��꭫�s��d3%�ZԔ�����$^L�bo���wCk�X-�3d|V����	έ>�	&��nU�W�����:a����F�ye������W�!�ʗ��|h�edm�խ�/&Jt�?�Q�w���(z��s���]�̔wN�?O+ǅ�0�qhv�ޏ�B��wf.�
�XlxVHYEB     400     1b0�rV���*7�a���V�9������X�.��p+K.&�7S��t�?�քѵ�ɨz�TkG�:�P�)o�,��߿�^����^6��,����߲���	ȕ$0�0�l�._�P������d�������u��ҸԂ���q�0��)2��B�`,���l.NG�{�d�Ϳ��.�3B(����_����~;�r�4U�)���v�݆�M�#��)p���ޓGrB��C���XH ��<A0x�N�9��9�P ����B~Cr%$>W�F8:Pc�ꖼh(�E(��:�Q\����|tM�`��\�q��eD5�"��~�t�Ƅ2'����3�ћ�����$��W:��.�A20�c��=f28��;����ƙ�S��hE; V`B����Xi<7PHR�j.O^°I�������@���S��XlxVHYEB     400     1b0f0��ٵ4:C*����������0x��g�3N"Z�����#Z�}]t$�)��oS.�7:?`:��R�����G���<��$���DU��$3�ol�q@�S�cX\ɹ�K��b|¼k �������wP��Y�� �rN2�5nmᣄq.;�s{��K�7A^�#b�0=���Dhic;�]�^�(2��/Ǉ1��L����4ݲ�+W�O�T�R��\a�V�ګo�i�;�Q�qg6�6r�A��3���T"�a(�T�4���p%4Ӥ�<�o�R�>��òQ�[�^@��޺����֮��R\�X;�6z��˾?m�+��a�9��գ˲ �,F� w
t9�˒"�>����[fj��_A_+/���4�1����k�[���c@R�Z�͊H�����H�&�1��[��T��b����(�e�mXlxVHYEB     400     170a0��S�u7)���_X��z�Ĵ�B)yA߂�e�y��;����L7Qŀ�jy&����	Ht���f����'��K��uc���iPx��Q,U�HgÐ����?�f��P$��'��0��H�?h |��XUhU��u�ȁ��T�e)2�Ҫؖћ�7D���XM�Da�ŋ�m�Eή��DSf���&cxBo M�ۆ*�u���"���D �����g��;����F����-Z ���^���v��{�8�y�v����|���	�����,����V�8�n��C��'֎۟���6�5a�Β`S4M~ك����L�}�`�����ħo�b�������aшx��f�*�9a�'["�`}XlxVHYEB     400     1f0w%c�x;U�[ �ص�e�逊cf�l]�X8cQ����-�n_^��		���)�?�rI�|�k[��ʅ)�C�w/#�lZrT9��ֵ�IC����=��1�1�F��?-��ԍ���77>�p��
-�l��#x��/�E��a��#o�
�=����f�p�Bb��e3n5�F�?�9����n6��"Ȥ⋇wa�s|��!��l���iJ��V3ہq�lˠ�$�Ơf^�7�W���x��
��k g���.,���+hyH��?����>g�U7��!���'�B=��4����by�*�o�/"
� �����~'
)5Qc�y�Q_}�}�{�u؜/��^��f�Z��vY��;� vz��q�@L�Cs�K�N�@�2��� j�3#?`��e���|^����8!XUgϻ�e��Q�(	�ʰ��+�0p&^�����E6E��(�3�d�Л�n&���^�����8.�Ƶ��o�6��XlxVHYEB     400     130e�\K��r�\[
)q�]�f�y͍;�����Rd��h��]G�]���@��俬f������5@�S���x0(f>�{���{�I�~_�-���:٘lfNn��/��f�a��l3%%N�Bv���] �.�n��H�F ���zx�s�M�ܜ\�z���	7`����Zڂɷ��@�F|K2��R��&��F����x��Ȫ�U��~d��>�nҪd���8w��_W�o��aV��#�T֢u��nX�$ W��_f�9�.��Գ4���# �C���b�$�5i�M'��%,�G�ϣ�px;�W��hZ�`ڴ�XlxVHYEB     400     190�w!��:4{Y��HN4H�~��5h���X�B�7�	���,2(k ]�qE�o)0���23�P�l�����.^�ՙ!A��`��hz6�[#굟�{������~�-U���0����������o��-@V�>0�.mEa��/�6y�V
}���%8�1���:m8��~�K�qZhl���bҸ)������%�Q�o��Ua�J���e�,����O'��!��]���fWV`���(�4o ��z��[_qVR��85�޾����A��3��=39ތ��(Z�B�ur��;J	Ъ��d�Q�)B#4�,I�xn��_�yAG��n���؁ƨ���=�cF��?Ѓ�����d��& !�4״۲�Aތ0��S�4*- g�(.�����5=�)�8�XlxVHYEB     400     190R&#�Q�u��Y����
Vnk��]������j`��t�	1�`�)c��\��^��]FB�&��v���%{*3a-�`���;k���w����5ƨG�NH_xڌ��rj�rb�8I$��r5��2p�k������:�4g����?�FY)�M������ؽ}��k	:�n���x,�ݹ�U���|�,˯��`8H�Q�g)�Ng���. ������͆���%���.0�0�+�g�2����F�m����߼9�ln�(�B����s��i�b��\�UNg���m��uq��K�m���YH%����s�*����}m�,�����Uk|�:�͌�u���Z��R�G���P��`��ld�A@�89����+�𔕷��MYݷXlxVHYEB     400     120��Ö���l?�tl��t>�;�#�t�h!W�赥Rw,� ��ڈ'ݽ��cϻ(b�Ĳ��� �m ��X�-�\��E1�fj�Ţ/�F�T
�)�Dw��s��+y��6x"X٥��\nl�l�[��1D�2ť� ��Y2��?�JI�5��,�-��s ��T��f%���İ����8��Y�2��W�}��QmI���S�HY�.���+5��۩��Y�+�R�x9H���Xr"2��{3▹Ij-0���Z@D�S�
�0��v�8|�"�Z��VaXlxVHYEB     400     170�	���F�חҘ)#����e�Li���o����+���wJw.��q�e~ T21i.?~�$��QY����e���o��v�õ95�Ri�s$GV9MU�9���b;E ѲA��I}Z<Z���E)u�U�����ݟz�fR�K�$�t�'cӝ��-�.66��˿I�.�y�#�v�֞���Ggc�~j\����t�| 8)���.D��2���E#Q�in�8D�M��P6���y���A�HĩG�}��	�rUm1�X���=д��L/dQ�'zpۘ'��ȁd���f���M���D��+"��*G����w����PƲ�`�0��C�'��[�#ӕ�V��X;7'�#(+�ƣq�pu�Ӯ����XlxVHYEB     400     170��������=%���#�؝y)����{O�z�S��V�5T�o�|��X]'�[+|u@��a	k��b�W�-'>��J؂O�)q���K�@�v���5#���o��r��s>�"��Х`S�6Nd6��
�˦38lQ��Se��]��K1E����Ƞ��s�K4������M��g���6�k������b�!�1�b�K��'�ٽ;#�̈y>���y���{��x�7��7���h�1B���^�P�[�4u�h6�����V���EE^ZOM�S�d�f�ￎ���u�Jx=W�k�|D�����>���L�~]MBY�G��)����ӑ�RN�Z'�����]嗞^���V���#�)��XlxVHYEB     400     180D���X���H��`>�����l��rLo�z�z��=�Bljw��zL�¥����_�*�M�|.Z%�NL��_oު)�V~Ϡ����@��W���j���{��Njx�JN���I�/^�u��ri��$r���,�N�k���U�����[��K�`��u��Pk� �q���-�����CYР�ZG<7����f��O���x��xn��ݞ���W��f`��M>?z�^���Ƞ6��P�&Bu⒦n}���
'@3Oy�( �	����A!q���e}B���(�l�e�
�݆Nқ7���L�ե���01-��!���p_O��C7�(D߁���eD����i՛B�S����1��z��N�4�H���&�r�XlxVHYEB     400     100��:�dtq	��������p:�u��@�E�� �Pd�q�h�z�凩l~��;sSx(��� P~�@�j�#��x�?D�He�=o��^o��u��O�G�0iH��}���g��	��Y֤?�p����I�?�4o%��>�X�@ty���'����������u���en͎�K��5��J���5�jK󫛞9��V�̂z�=������B�׋�q�7v��:�	�Wl�F"���WK���e������XlxVHYEB     400     150��YJ=�����5Q��y�1<!��*h8�NTq�5z�V�B�I��a�	M�]T��� �o�0�"�هN���B�c��v
 �bv�w+U�w
B=hn��t���_ʠ�HY� �ɲ[]F@���#�(��C)�PW��������9Y�$y#W済�ˌ��w@������k��n̄xj��?�@l�ɉ�� 7�2��g/}x#eꨒ#�V�_��Fr��D�U	��6q��O�s�Lx2aX4F[�ރ�*]���:fgE�梳Á��~]�4��Z�s��nӹ�i" ����6~�bk����t��:7x�:��I�y�AXlxVHYEB     400     150|N��Mms�HvF-���_����`���I3�逵x'�oxÙ��̀��0\�͊�s���C�6���3����\���!�t�f�	���c���f�Y���c�s��ϞU���=��޳hgZ�(�0����i�S���]�i:�ѭ�h�H�.�E����B������Bu��ȩ����{MK��Y���8;ݦ�̶�`�=Ѥ-��qN�&̣��;^�ͬ��J@��:�ީc���v|��)r:�)DP�? )��B*������T�`�N-G��k�v@X��r�jF�"e��iyV��b�(5%P�]q�����M���3���XlxVHYEB     400     150�e:�ь��K � 9�=��>J��dy� �V���hq�� R��8����a/T�B���Ő3m�����A�� �����oa2�.=P=" ��A���\�V�S���~)[����6�$׏Q�+�`?�r�������:DJ��uՒ՞��n�������O�1{Y��1%%��}�"f >����aLVϥ���H�.ý�6���Y@,n���?�¤m�i�Q��k�|ȴ\j%t����C���O�F��V�6�>s{S�F�_�:�z�ƥ��l�`�~7��2t[�w�v��⬝�#�?Tc�Ts`�ܥ}g�}�����37��)Y��@���8g���XlxVHYEB     400     180��ƅD
AĢ�]<h�IF�>��SοZ}Eٴ��$ü�_]A KH�sx�Ce��x���3��8��'F�,�a�BI~#!��J�0� �wj�{��QcGl<ؿdH��ա�g��,٣�>n��GW掛y�w���8]��&|���ooR��Z�Q�P������P�$~T�w�j��ͦ�)N��@ �+��$�J;x�ݕ�I��޹�f	����4P�&��㩫��=ؙ����h�l3秆�N�����H�������q��"��</���'�����b�Q�y���e�Y��g��x�4Ҕt��ǻ��S��1��;YK�y�_�Z������,��*DU���T��c˖���&�.��0`�Œ�����a��/��K���XlxVHYEB     400     160���bsw�P�ͳID}��R;�Rg+\:M�!8J��]�{d��*	k�a��w60Ӌ�5�QG^�\��4�E�w0B{��t	op˘<1H"�f��>�A"C���I��|��X�.Á�� �_鄶ma�1���i�VNp�Ա��e`�\����b����-q��tɲ��K�c�G2ԃ^0��nc�8������N�z_�k2�լ��oI̍�E#��!oC7�e>�'rrD;�1:NUB�h�9'Xe��w��6һە�Ûbq?������x�E*���[Q���L�	5��?b���Ր�OT�~%���k���>�:�fnmO������k��f�h��@7�XlxVHYEB     400     1a01p4t��)KQ���ͼ��z��Mh��8�0�E��V�ް�1Y�<4�!1����I��%��̿8 �u[�AT�A���vi�a�CC�!��0�"��i���� �Ŗ��&��6r��,62΄�LL\�Xr<"HL�LqKwt�6���9[�Ie�w�ϧq�j���N�R��k`�n��D~��	���ʠ$�_�ѻ+��2y�,R�<�P:_?筌S�����W���|}ٳNj0����6ti�c;�Af6�#_�+��Df���H��77wB��,٦�Me���Ш|��@��Y���n��^%�Sړ)ǋr�M#{%�Z3�E�iI�x,A�ܡ3��i�:C��m�� Ġ�~D���ܯeè�\�)״	C���v�r����A����9��n
r�tT�L/�XlxVHYEB     400     1f0�f��I)��l�\a6?]���}�G
"^���z��E�s�NL�gNᝤIËB8%�rk��Z��as�vr(rf*�9���͛�į����75MoHڑ�K��s|<m���ji翹�z���H4��0d!�m���lY��X�ZH�;l0M%¾}�F �j�ԡ��MX-��[�˦I�:MkO>���ye��3U�tӤ�u��1t����7A3�ɜS��G�U`z��u�MwhvK(�h�O:7���Vӷ��)ńblر޿!��`��@s��n����D m\P�j�s,4�����S?P�pP��%Dʺ�ch�/�T.��n�Ij���i-�x�#�!���N�E}��}�!$�ɦ���h�F�w��am���tH.��k��޻*��k��n�Z��!�3�u$rF�#{�l�Knu�2�?s�i�nߵFT	o�d���$�d��"%��(��eT�O��1���4���@��T�AOXlxVHYEB     400     140����mT�6!��I%Awo��U�-�֢���$wR ��踕?Z�3��De�ye�nc� ya]��s����^�����T�������rv�^^iC%��_j����;�����{�m$��p�Y:�Ӝ4�Q;qnK-0��g��k�U�?���i��F���Ӛn�o��PW�� c����������E����[�P0t�ޞ�c��V��%m�Is\#���Z�1mFG�,P�ϧ�Y��0���"��N��7;1��KH��^8��+gH���#ȉ�N�]�V��!�Te�����e� K����')$,��al���XlxVHYEB     400     140|�Be�`��]����kMr����ݫ����5������r&9�2H��E��)���K:�9�8� o}�������uw�a`�4	��s��dmw��KX���%�3�n�&d���~�@�)���m���.)'�4�	m�Wp$�F�O.�tďPtd�R��&c~=���ߝg�03���'��,���2�bocE3І��E�t���*v{n`��=S�R�}��ACQvw��\��Wo�O +轙�M�?�L]����\��I<J�7.5c���T�p0o9,[�^V�n�p�	�
�8V87�	���WDx�I����f�FuXlxVHYEB     400     1e0&�Kk$x��a�1I�П�q\�l\E�Ǚ�ct��V�A�_�>��B�� 1Vr>R�q*b��8k?=ʃ���X����[�=�d�
���7+�9jfYJ�(g��t�F�@�0IL��ݢh�)�����u!�he�DjM��Q3�s}�;��u0z��;��^��!F����s+���^��te����9U���Z��e���3�I���RM���K� B��P�G�^�H�FA���nk Ɖ*ϒ�K8ur�����h�d��s�@��=e�1F���W��1k���0�3?��ǜQ�)(��;���F��9ei�z/ղ_Ѭ,����	/k��3&�q4�`祯��"����SD��Q�|B��Uuӌ�3�J�J�,��=63�ٛ���k�}�7�;�FtJhBq���3��� ��J��6�f��m�f|#8,O�"Ȁ������y�nJr�:o�2R�/�4C���ݚAz�U���J�8XlxVHYEB      90      90�����|F�!�qLR����AIb�^�eV���q���E�����r"PK+qa{�H��lZ��5q�y^%��t�lK٢9�`�F�O'��"���3��05oUī���C�"�L���WhV1�c�Li���C��"cL�O��0