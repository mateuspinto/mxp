`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6384)
`protect data_block
0USWSUGxovGsyBJteYpEodgVN+9UzPM4xcWZnw3HLToETt/97kCsyXX5yUQR8fUVzT8H03WDX0jT
6MIEb8zN4Epnn/MovzxysUohy+FnHxjp3kR1s9R+Gn186PL0BsouyS6WWaGfzUZ9PWk6mu37C3O3
fUFHruZc5n754ZnjZQLQ0C9LzUzbEjYDU6kStpsEzjcq09B03/tw71hjNQsArqVR+uhGvaVcUcfO
88m+0FsisPV37ZcTTpDYS9ulvRQP6oyhh/taIX4mcKm4u+Y6boXNmhNJW+XTrQrntE0htVkOJGNm
QdFPaQ8foF02p0lp0Vg+x/KtI4crvuE1GqxGvWs0mRIm2GKHcgj1PT4CZwRnBXfykMjzQFhEPTdS
XlSemfgfcEfEUIxNz7/jiu6xvCLdAhuzIRZGNvHa0P+8Eql3qT1XhAonZ9Z5yRV1AilrR89RzsGu
MB7wj+7eFjdISCRERsc+RdUuQEuBvh6MOD7xcP6rnbp5DTD+JPyVtxnVi/DmPUWEGQQx3HFqvqP6
URGXkA4fK5t+ErjMjkZVYMAa8szvYlpi0eb0MmRldvo9Ka0s2iurga7XxN5hMbqgWUQ1nbxuP7BE
QNjSkqvk+G6d9KEetr/xUAbMANbcZjts+D6LCLnqJHuntfJ42esTVOChXAkFJYoNkBGzpq+3Tsf/
df3i53TQd6oWkU+QiJ/VueFtvNC1wPD0/igtBlGN+hO6gpbtJL7SLDANFf4GtQM531DzFNyCLj7B
wgQQkZAHytVz6K/NQg+GOqZ/KqM32HSnY4Uz/xbePZnADPVVgLQIJI8o38/aQeqwyPCrjQNlDSby
GhJGrcwPy5alzID/szTdjVqRPaYx03GKBwlANnQwu6gE6XjGHIy1CrNAxfKLO73JlJpF7xway2X6
yPB6ewtxH1aPcxYZfTaVA6tBBaYYQhA+fe8e/TMHkCToK9bqvKGmIVYlr6eiaVTXvm8MJac9htFx
c3rGihrjQvLF6R50sg2Yn/wmq0pVGY0aoIR6pgQ/yvFWlVWIh3I4fcjGPs8Bkf7l5puHhxE7o4Oc
nfKrRzIM4l+Av2sVO52Tw0bhjb+b57//bTbFa2VyGjEQehxg+oaH1k3mOqltym0obY1c04FXIF+f
K7y4LQJyuwVDCp3rvPa/6fN58nUHjooZTCXAgdIxWkQW9Hq8HId5WhJneOQrolrG29fgHseWFVZH
x3fw5cdEGVW4H0HF4vJb0YFr6QjDxXm7IFaJh1MiTIBkoIUgcIBbjIoFK6L2FqshRot/qp9EoMvv
g3UhPx55/lzgIYeYUBmxq1UQxg/OIcqUtsTLQmoLXx0unFRSp3p9vzSxJe7gw45mlDiZJoKQ/mVo
zYc3/c0UM27Uh/uWiU2apikPACAW6f/lwaQBtOOhHlgYYyrTiMjJQ8KBWrpqP0T97Npfco4EWmX2
XarQphQdaXVX2Xu/hgu6cwmaUzodb0SD9e1sdv/S89geeymuZ/2Kn4CR+Ib9rXCCfwjLKO035qfG
kmkklSXecW7wwn0sOQs4cZW84Lmkxl2hCv3T0Zlq9zmrDDzsEvsA4bGPVV+2cWrCHPN0tCO1/uhF
hg8AsaNjoQZn1Y5gzPokZRFEtJw8W+q7mOl0BSSfUB3cf1atv+AP5/wH0/A9VOv5lOEmn29L5JzU
ZnffdOnKVTh2Nyr9IqgFU2kLnMYYAVkQQgu/eRah6DxeJ9QZQ/BL4xmHFL7OIpRMjx2FBRDxzUUT
pL+VMD1rwKutEJbpzRLBucXQIiSPmWWZ931U+Zr41fDjJERtkV4to3zLcufLr2jliCfdaqKZ615F
199sOPIHbalHV8QFD3jq6bWy+tVQRiySbmIdsFsLtBTYOofkHHoRcc1oPeZBJLZFXEjvEaBwK5Ay
oi9NIk9zJRAwAHF9/EjKQ1iAhXKhk8pShrcc514GQmywRP/jZKoAonqx87xj6jZcZxhX1EgL684q
hb8QlQ9udvREfIUvMcEAxX8JpcaXaeYhnxVXlrl/8qeJSp8PHkUAzhwxTaLOu2p2pY8PyDlH6hLi
fp8PQkjmYiyOu/P+5EjAi9O0kRYcfUqAVWWnt7vUCRfOiZWgm84+J1FEvZB4WpqN5bMtfKAhqO+H
vm+VjH2bdQP+uNBZ+QNBiBcKxCHAXcb6QkTC6KBCcjrLuY6n9eWmzmBc9Ri3D9aFMM26+6QeqZNC
TChi457hnPZdqNZN9yVzqLelytzR0DbEl6imytBNsZ3YCziOOJbQbReOAkeDqq+k/PzVI117cSrz
96u9p3pq7B1FEVWmbR1NgwuML41GJoul/kL856tmuzRtd9OiOtRAM9Upij+X+o6O2iG336/o00ge
0PeLfwzw7olbZ4QqXqH4tzwbbsKsCe2gZc8Sg5uabd7IoYg46nFxkk52N5Bo1Z7SyCqgFUDsdNqz
1QbBWZTVKlHo29tzehY35WKW+xod9jwTHWacCn8GZvsySpVQHpmXyWoX0F6pMNuK/cY0y6pvMtir
1lMAgLcqlxyrmjcSmxNNhnApzS9IWJ1swxPTNtYbZHSBl5FczW0l1BwG/lpCfKIQN5v39lWogeut
iM3p4PJcelG1ecLmAwIaAVq/Owt0w3PCFCQZY1f6wRziSnUJ9yyl3mXNcyLOLZAYoBIfv/mpGtrJ
iS5RANIu0NRPFUILZxZx2hrcnYoJhC2TGP7x1mveuTnDgXdDjXu3AaQUwLWdGLVr1c34Nu7/gg3x
+7rnq2bwtGDfODH/8UDFcEfSn1rVU8vYsWxbsU3QkEM1yb9yQF5Yq+OjVn2ZxNsEyrWe34cU7rfN
+cQGJhklzwNrHDueymi106WMQD62oorPAUviaOAKMj9bdBhrMr+DZrTmShGApKcPK8D2Mw6gVobB
fQm09Wkz8r9XrX9Q4TL4tJSKxGqYO725yAruXvhcMHw0iPYV9jUbcRdZxvvSKHeoDExYg9ydt2Sj
IwesYlgmIaAoHFH3XvwVcisJaAPH9p+zOSibnLUopALYC3g3sZt0IPT4n/Q7PEPJRuLoen4JwnuS
gZa2KzaGizxICzqKM1W/TRWTbS9DLctuFL3Unljuo4lMNGdTA1TBNTVylsbS2AOsG604mhLw85tI
KnGiSquZYgh6tJSHytZYdkt7fs+j0Jt8qg02bSWaZ1Ns8JhncXDOao6uLWoXHXggIOdj7N3ypYcJ
rTae/1hRylHNHqheLsAdcDVpPQwpodxb/Jtv8Luwl1HzKgLfVjFPPbtYCy2z6eQiLyIuf4Jiynw/
tuBNBfaEgQruhIM0ILolFEl6DmIkgAURjYvSEo7HLEL+lDw8u0fuMIgYo5sKpEuVO/e+Jd0zVvL5
u9Ee+Z+EUtOxC8CdEjTYpc6Z+JTYaFEIQot/QVdxNn1qcVl8Xh2cLeCBSudHd6pjGIjVUoXG33aW
7jAhoZb43aE51tOKoyiBi/lF3u9lXKw95TotFuzBA4e0ZKs3MFonA42cbBBlpIYIT/yfCijw0xa6
Z/NmCAax28LnMcJHlamEZKEUz+WGm30bHk8nxztdbFEMM+c69Pbb2AEruBFe/MbXszsnXyPQrzkd
HN6tzMCCoORzf5vuAMo8zIa7oqzfIow7kjdOQtH3e783NTsB8XewmbAXu7X/MyeLIu5QVUYc53mn
sxm39ntYRXBGUWmc3UdC8qXsTo6Ct84QfmBYTT4+Hn6HfHFkG1RKMPxeZD/sYNlpuVVXwCSBnIIv
fcbNG3KpDit87TL0im3MpicP6KHf7OTOBBzJHFbm5ih+7neM7vPNNRCmb0tURrJpl9E/QX9rU72/
15pHzodVx+nRviOFR5XkOMM56vKV+fQHppwdCo6ZYhtujEw4hZR6VYSG+deTWODGm+TWUlnOHz1f
jMh1YETIvrhb56bTABmc9mtMU74GmKMAK1L05ZJDllI4rzN4nZeRqEnHBzDTUKO/xuwXmpH2dw3T
K4ZGQP0JPZCFOyqLf91Rm7/KxT2OEtPXG3PduYJPhVkeQgUb02mg9CRes+vSFEyayx8M+ypTaVso
iqCgER/zzQypTfs8T/SOl3JzQyCa4c5bi8Zo6TB2QBjOgA+BzM2gZeBA3WvNiklhNOHAAimy5xT5
UcVF3QKUEjI6qXjlPiPh/O93ILKfTdvJAIZQYel3sTW1H5qxKNsvlC1bCWPk3cPBjPzJPIW+Oze2
Vo7S/hr42EvQqiUKr+9ZxaR5KCPsOmuKdfTEL/L8QZeep7APpnbYFzgTC+BxWH8PY9J7x0bSs7H4
TUvhZA5dDZqdQg7RXLGd09+pTfbUdR5OA3479Akf6SiDuCQ5CP5PjQcHmmmHQVR7mxRJARs64j9F
mOkSLAcAtLZhDa3gBhtTLYmgANmXDi9pQC/zKTNTUmfRUP7RoLE4uMNz+/ITnJwAjNbiZuJBOFzs
eoSmStZf6gQpevOwHS+eA44FtssX7tB7Rl71yHFLuMvsD1sVcV+m5cRlZIL6+pCBb3DnRbJYwosx
aF5LtziJLmx7UCodgOq+iHltJxVw5Gp7+PUz7fQBy7f7ycDLI5gllJ2/kV1UyIyZ05lys9hBlp00
FMaedogKp9fhU39xTlPMxNgyHzZZic0QiIFOEfFRVW2Fd8YI1ipDKbFTObZS++g+894J4+ETlYnG
Xduy65LL0MFKywtndgU9qXgWRTeboQCFk83UavGYvnnyWMM5ZGU8dXE82XJ5vyRNskUNDAoFgr4d
CyIY+MUb5I2QQS/RaZ8RzgW6YvDKpb5GuKS2a2l+f//tRz0RmHIs0wjaFuKqqJ2sGok8p9h0Gg6B
vLcJHu8BIdvSJgUHsjB3rQbFqMRGCfmU14WqgaPYRZacXYxOqitbjRU5JsaYH48kldpUhY4Vy+Um
i3aSIcTx50+BGP2tuSICbP0mXDfKxjC1773cnBjqaBvqmKyQg61uGXBuSwVyDO4mNroS22dRt2sJ
aw2XtPn+hSY8idHww4JDFsSVsXspwexRtuB4i+VQTXzZpXi+iwtQJZI2O6Cy+Mod/4t58yUp3Nmz
TUgZEgKBbFiKOQ5vbZu/Ip7QiOwT3frdcKcCNTHFGCS797X37Uo2LEAYy6Kr7MSzsDU5BKy3HQxp
rgkUflIl64tEJ3uQpFNeEr9s0NbVbhoQWuG6tFCQdPQqWSdDKphqgMZ773ZX4+1WWZYlqqUdIQIS
TJtjWO15/Ap8pOZpdA3ID7ZL8ooFl6xzEGseEYjsqoAzE0PO4bMdBs1+8uLbd2D92F57l4p3shI0
ATH8+R4mLpAAeKyGkBgFAePp+aHMAp+CsrtjyDSbf8E0VMMdu+1SaIkEFYeg0cib65FjLFlkwJUZ
/b/Uvn2wmAE2xv6EG1sbfZGqVnqU7/EFV0ZU7Z0tiGMHxl7my11toMm4HCxEZFw17BV3S7H4tHfE
IEnzvNi3DzVMXRfRVDHpHOd0Q/fptUC9TW6C06q+XPgpwhtf9scuBzOhSlziJ98/zh/2f/Lk3hpa
OKSOthGcixgmnwIhP+jXifpbMrqyVetaWZ4RdKZdalatwas4Qt9sKzdW05Zh3ymjvnx+nh+AXxp2
3ggHXQw9MQHpXQzpPpJNam6KkuGGN6kmSLHc5xK8jDKHcT1fvJM8nE7iucSg6pXdc9vT/VOOErJr
KiuGDSZlsP77y+EaPPuDiqUXNWjBhiAEkFvrIWWCeZ5GYW520zSx6wI3XmEyRl9lY8p8J/Q4YlUe
wi9ZtKXui3H/iUNJp9Kxv/ndAl7xUgm4JmYt7bHzGVan3DhLwbdlTF0aauDSCOWg3v60wKu4PyLG
m3gBsPvb5SRz04acl0QN2NUdLRlOIaDXIJ7NCe+2ywyZjEE6snBS/x1B2J49lr43HmSXNTRfDS26
qeO1DsGWQufKOQg+ANFPznNj6R+iZnkCHxKDH0B+kU7V2mScHgubrUipnc44cg25JPaEkbaTEh+r
n65ECBxXMG71IDuMmKrTLS/xNkvRX3KD0ikeWs3t/AVw+EL2Dr+njn2wVST51Toc1xfWagf3L0U2
R5LYadRy5vFAimY4dM35vFYjJOLKpLo4sm93+8luRZqS/B+CiTAtcR4TRz+fEl6Y5mFzvRf89uC1
OBTXw1ReIQJHG7TmnpcD2tz8811kjJNUkGBrZF66MiRMnE7Jvc38hx5ca7W1+iFb0EvvPslapBeh
4tVPLAtei3HNtUlN7PS94H354dXStg5SUJG5FBQERRob2UaszccRNcbYrw4i3P32VS2ALm4cWhBw
Vj0/w3K2+suQDOG7+a/gLdRfz97N4HBRTQeygkoqzY87/Iv53OepMUrR8zAPBqdGbGHCt6ZGMbCh
EAaPrBW1RXCMPZzFbjLCUTnYwrt6PQsNWaRuqVmmZC/IduCf4gD9EpGfVAaAdzVz4k4xVloBNJft
hweQr1Bvm/TppJoUxUqpy0O53dLT7+c85L2aO9Dwc7QO6uXKuSzz0jpYCmTElPDa1t7MgsX5qi7N
+7qyCzrJQbDpe9NI9R0GnV0B/kLbVslLAaE1HPkaNUROqzAYw5T+0nWkfiY9yzwm9pzdVyFG5qr3
UBEjAW+RLML5nhbQWZEpl+/hTXamQcZx12O7fjwGsRSvaGH4r5/q8gDoSi9G8Daqk69LvicUNsKY
2W95LCfy/dZybJCfUglr9fqCBHR78oqf+XtBEW1z18wzb23EwkqTvKOIaq3lNaYsfSUklzNWHa9v
ayLMcwxkeOHATbBv3NDBJyIoVg8aIpb6R8DNgtpi+ZpUtVYsfoiJMwOzthD43y+MMMXAyZ9MrM9m
Fz7Sf7nWSW1vkRMyNJV5vqcZkPIPmxP4ab9dmAcA/T1idYtVIYIoXwvTaRRgKaK2m33MY9sjcWb3
YC99+tnaSVRgMHWhpHYVNR1wQWpb0bomk7Hu1s5AZtD9Tgmt65asK0aY4FxnS49GFgL9Pb6a4lyi
fpUiTC7/8zD612zFp3ZgjPPX+x+7g0/81L3+JlYUrysSy1BFRIcy6aLebnCFrzBqhKLHQ0qWauce
VF6eUqitElReDjeuDMaehpQEtkCvjN1Hs7/cxbfNg2BHC8yQK9PzOEV5Nm+5rWwVP/wq3MSqKw2I
lfjKlpiZVC21N4Ip1ioqT4WoC4Qc+QC7yUUdX++gVynwA+nTzOYpNm/mzJb7CQeAaKySVcQdHG0L
NonpSHEWp17r7GpsDjbJpYyID2c2Yr7d5J9hrOQfVqUglo1dlyt//l7DjV5yEVOeBwUMEaJOTIzm
MFGgvCz02Fkeb6oruyq3MTxIBlx75jbeeNomeZTxI1dn71Hphgf1LlqglFb3ooxR27FO3IJG2fQW
RU6HA9DN4SD0Aq9zzBHJvVkYK3FOYIJqGA2oRg3Saz924A0f+Rflx4UDstdsS02r8yOXPxYbA6T2
fW3Syczf9PgZSQKYNCdGiLo0UXSvQQDfZb2Os3L+Bm1c4iEC5AiIv+uwGUBgjyXffJdtB+UZTFdf
2bpQ347Y14C6WZZFAy5y1mGfmVzZUDdp7VJt5quOFAQm/2k92LXCJeib0nkYKUzR+9f9FcOHWL14
cI2fqKrK8uoedZfesgsbebLW9sVfl7yvSLa7b24RdZo8sxKasr17ftYQyzPLJ5Q/l9S6gPdP19XB
dCpqtzYfI91swKTi5mEKM/Nqty23LZSCZKzkYf6Me8RTG/uJjgp6fs6ccdkQ2jEcbx0YVG6aBVHu
LhHKJipT0uVl527Gm1ygWN/lHlbO23q11QGvHIvj/HxUal+eEsc0G77iX4sqcdEQjvx4LvunH51c
xqvurtbUkVorTeltfG4JBSUJzcWBtQcgngL6FoKUXafmlloGTOLIwh1NPsUJ0jvTOwK3kbqGudyA
dngaE07/zoifbrAQOuvMnXW2P2D0LxLvQeYUwsP3FGDv4OWszeqmielliyZpYCmlePMXcDRVn0Qp
OSu3a6xgRkGizEGANYEil0XQ5UJIYoqweooZxLjqbUrtGCuBxi+gd+BKNGLTZ1d2Rq8fZjEpnrwy
p2Vad1i6ROmg2/kR3kF+I2OdmHWkwLUedq2691X0Nf2H2ivntWrpNkAiRmWhwZCGa0R+J/Jo7qpQ
FhqgLSUDuHWuv7kMFkCGcvx7AeaDVyNV9RgBVB0geoPhcCp+Lz8/AtS1NS1/1dURZ0r8ATEQYNNU
qllXpXdeQHL0oa2ez7QC0PYnS/UWaGY1XnhUH6Tf5WHDszEXi3gCESRo9bgGEe5rmv//igurBel/
4J8VtPXjFfV14yKL/clrsvmXVmWHyp8pm+ESU7LuZQAapG1FecE03E7jJmHdXA+4558wjMieeEli
rGaZvGfHXJOX85H6kR4TckcYLV2WEVJUrTOKIJjQ0MlvWKCa8xlngFT2tnyNF95BUVVjF0au+ywX
DGkqlI826SjinMVta9F/3RV92EO5Kq2eP5clyJYLTnhFwv4GoQrTX/KPgVq6oQJjoZZB+mmatrZR
RR1C11T6IE8yBAyvlK4VWs7iWrw2+pJCig8+PU+HVKbDBPvXeB05DY2JAG+PC9J5SoELN7YpiEcF
`protect end_protected
