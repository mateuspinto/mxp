��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���a�`q}�-{7q�s���������H|�?`�G�{s	i�'��]x�r:��ֵq2$�F�����b�Z����%���K��5̛3�X4(�L��ar��!�3>4JR{/�q�1�ud���B9��yw�{R�N@�)���Z[^3T}�{���M�����(x�Çw��/T�� � b�� }�po�������G�$aξ�gw<ר�|�H�&�e{%7su��qE��T��-�{�Zg�H���f�}��$�G�؏�>@n�N&�����J������&�0=��Cq��&��j�^�P��W�U�d3�i���Li�l� ��@�z"�w]O�K�2#
#+k���_���6��<W�b5h}� �\b�$qwrp-�恅�mD�:`҆g�glTP�<t���8��4UՔ���.Uiʥ �2Q'�����h�k�-1�|�*�j!F��5B�� *?/n�>O��K�Øb�W�JpCy�]��]70�c���\j�����Gw�뎛Z�nl�o8L#���]���nۘ�j��~��2{A��섑�� G.
���P?��f.j�2*����˖V��!6���;�{�u����Ht\���m�Qͳɲ]�D��]D��b݁nJ� p���Id�`�tϬ��*����b�jӆ�� -�/c]���i�S �]��]'��=��6Q ು�7�{,�6�DS%�t����(�~k,�+l:l�������B0��['a���t�%f׺�i°UQ��;��S�-��9(�x|��y��QhJ�������sd���@� {e�=3�{Ѫ9�&���ȀRL�� ӆ�C�wo+Q0�Ϝ��顦j<~}j��2|ϡ'F�S���7��D�n�i��5�(�� 1|�+2�4mnܩ�j1
��o��wV�d�A"3Y�ֽ��i�d��Tٙ�n:�3�6/V������ۨU�3H�},��m��#����}`QT�P�G�eo��[4O$1�E��@rL�4�ݸ������֯ ��9�ar�ЗZ�ç��Pz:�9�� KS-�K��0*U�`J����"��\E�Im|��Mԫ^��!��MG�����)����Ԩi�ć̲Z;N25�Z�Œ�H��
��[�j�sݥ3$�Y�m�D:>���Ο̕�:�]&�Gk�\Z޾�!���'��T�d��9b,�ð�c�n'O+�4'��H�����!�j CM�=g1�Bh�[/��͸H`�4���p.Rӥ���܉����ckoK�����O��Y^|Ř���U���f���������'H�Pq*C���?���/�+��d�
JvS��C��m�c,�:��E&��7|��P�����Np�|��;|z��ESU�\4��K�u�r�Fx��l&���	{���.Å�\����v����Z�����j�3��zYV'<G�3���`�Iİ&�3��Jk?m�~�!�[����=�lT��[J���.(_��@1h�\R�j/��������cԦ3�UC�#`/�̼AEp������C����0d�(���*~_p8�c��#��Z$��Jk���ֽo%���9�h�Dd��u��2�Ӌ��=*���,|S/kE���028[8���^���N͖�<���i�ׯ��Hjũ_�? p�Z���X4j��>J�~���>'g�lԤ)+�� vkZ�3���;�;�1�竱:�Gi�����7��"�i�S�� F����!<+���p�D�/Bx��71�l���!�q����JG�J @V���c�~c���C�XĖ
���v?A���2�,�<�6�ID�@z�6���f�N����Guv�m��פ��=A��_[f�4�j�s(��*e�a&�G��ۨ�;Y��Y� ����(��x�P��
] �������y��)#H8�1�<��/K�6���Qe(�HRO�������=^u��<ۻٷ@��g�2� �3K��t�ޫ��σK����G��N�v�_��c���ζ��5��͢��h�>�m��gCa;s�_��8�K����U�ߍ&LN%��ms:��3�% HN�W?cApԨ;�U
�4o?0�W�
�K����7�iW��Ɏdɫ��!��J�%��ɟW#�Gjg��3W	���:���>�M5,́I؅���/���	�m�t���;����l��9���Έ�{�2͕]��+
���/�����9���`@�*�|��}�$I��&4�эh�.8&p����<NP��k��?
sQ�AY�/&P�q.E��ÚT���{l���bnȣ	�.&���Ȗ�wA�X8��:��Q~��̀��>+���4�\���@��o9� BMm.���)����.�\�r��R�pG����3�y��o�(�hb�L���!Lj?p�8!�*d��8K<�h���\|�.�I�\��O�����n��u�6#��c0,b��R�u�۠Ջ���c�*U�CӝOh�qc���~A��* �/�"���'��eq���Fˤ7k�1��~)y��抣�Ѧ���x ��FW�.���F��rZ5�h���{�H�76�`1��:]t*f�=�g�;�F����Bs'7� q��B��,������+��.�����ӝ�(L�3�k=��*a���k��"�v�.�61ĞAPun<����)�`�]aS?�\cP'ߵ#!�	���W�插 �|_��;���כ)Q�[��v�#���_�}{�.ߙIxU��@y��uh6I�X��[jqJ��V��K��r�_����1x�Ǔ���6��}��U��gR�7�]ǈ�y�9��0˪5v
���.o$#��O�"����ˮ-=	K���,�jCZ�NBr��M�ʝ�ūUiB9 �P���ԒMz5�3�b����Bǌw,W��%�o��*3�K��P߱�W�c��$aa<�˓�1���O�_�0������O�ɀ��74�"Tݚ�f��	�oy�Q)�ޯN"��bF.��S@A�`�w/&H��)PL䩏Xr�b�oHg�ϵ��q��"7Cm��r�,jY�bZ_͖h?i6���!�����7��¶�?f��Z�N�#Gi����6����	�����1����F��(h�1 ��Ai}k�%tTy���7vqz�~�.�RƄ���Ȯ�o�>�=����-(z�·'ю{<R��>Y��}<u�qN׌G������2��2��g��O/)�v�3��['��l\%e�3����#��5�Ms��3�$f�2�kF�{�m�Fm��£z���,�܍�_���]�|�t��D2+�%̜[��&�Ҍ�bL�2#i�Ɣ�sdT{?N%x�V���Gї��Xw�έ���	q�珢�,= l�sJ�_�ua�k��@ܽ�9:����,˦�4\��VQuTӎhU��zK��pŵ�398�g�[�y|��xR;�Q�N-Tm5�p���(p����ډ��fu�u]f�M�+����o��Y��iC���õ���x5��Y ��N�@y�T��=�'Y_�4�D��7:�PE�K����`�K�Q
f s�Q�Id�(R��:��|#[| ���̊au�|!dLQ���V
��G���5,i]��%�<"`^�mt�|�����]�*ק�AҺ^j��!���_�+d��U�E���4���%ǂ!�0~���^)�܈ϾD�Ĕ9�?!P��W)a �t��s.1`� ��럘���㬥P8
h���Ȋ��7�ǂ
���J���>��b���T�2�O�u`��Ng�M|����V��Ý`�?>��-��^֌���tj�6�"�O��ʭ���4����U(����l�1��"x���z놰�dȖK�K��K�u�<������Nv��Y�~��m�i$FL]$:�<���`�r*���.�Ѧ��y�$�@ז�7w�6E֠{`�)��y)%P�-9�Qst�uC��>�3�!�����c�9���2.e����x�d0K�O���zy��Mv�<�/5�{���āA*5���?����Ǉ���	�E� �6�0�z�� ����;�ڷ�U5�ԝ'L��Gˑl4���P����3���Ӽ�Ϣ������`�n@;ҋ�Z��G��YN��,���Cc/�n��n��ǅ)ᱨ�Qt���`õ��Uo��+���!�x(����A�{Ӹ��j�3��IMq�Z�k�GA}�<q�:2���b[�j|1?���(6A�PP�?F�!/C��^n����󢂣��v86�4�l n���)�2�XÀ'fwi�W»��}�N��wf�$\�4�Lc��(�vP*R��M�m��s�Y�[mRu��r�tǶn	��򪢷y6��s���TI�u	/��h�7DE����\V���Ɛ�t5R)���]�1�e6�\�Γ������DOK֫eT����L�H��ʼ����·Y^ރRH�R�5<�ѴN�?7��'��I�0*-�%f�=E��c�L<�o�N�ӏM��
3�tT2�C2���]H�������H���B5Tr������N/����>7*�:��2t��a�}28���7XN�3�Am�C���h��QD�!+�@]�����0�߈J�U�������Z݊������y��~�� ^y�k�U�O*�N�=g
�76:Z�o�I���[�
:R���6zE���cĘ_��S@�і<�, Uv��Ʒ�(D��Ω�t �T��mޯ[�6�0��
<v����W���/�ymw�0VErN�(����dJbT�`"H�k5��`[j�A#��� c୳��������&�1�4>���-F�Pz�����-
y���R�����捹ou�TQŔ��x�'�B�<�;�ܖ����W!�֊�_ʝv�X�,�)����,���`ľ҈N��=�-�uʢ@l���V���Ȉ:�q�kظ�%d�؎�Ԇ�X-��ڤ09�$�?�m~��FӌI�q^�<�q_:!"1s@�yi�wHt�2�V)oA���δ`�I�r�Q�ڴ3HJK
_��Ua����-��c����J�@��hƞ�I�r�((g���8�5�q��ѥ����G�%�F��4�e����T�lڙ�& X�����1�5������M���7 �V؃T�.<aU^C�(EL=�df����$Kaz:7�|�����'�y���Y��	�<�"����૩�A%��K������vjvS=.]�
$����-�������`�$�qm�Ih�M��q���I��^�`���7�}��� �����!X�~�&���O�J�q�H-#q��A�0�-�į8���́;��-A�l>4C��i+1��*���c��9;�0-�=�Pi܎�3���p�ݏ�t�@/�^1Ah��{Á��\���F���е.�G�*$�~�C莳��!iŽ�X)�+R�Jۄd��0[�`�v���0���o��}?X{�{Hı�\Y��*��O�~��uV���A� n&�GSN�c&	��Z<�0!�V�$�	A�\�Ch,�M��{VZ�&;�v�n��ha�z�P���&�yv�������1���C̅]���幈U�G���X�a��� �8F<��S��4ޑ������}a&rBWqD�Uœ��X>F��ql�@���q����JVN�ڶ��fH�eq*L�#KO�kI/L��Z���:?6���H-����n�V|�qh���u�ģ����%��S�z��=}M�p,�� _�v:Iob$���,�]xoVT����`�¦����.�Řd�.g�+*�����:1���'1�AΈKE62Ea�/�S��ӾU�����n��z��H�MT͂R�nUQ�`�!/ 
S�.T����P�̛��K��]���7sktr�w�?�������?ĞzOn9�e��&�q	,�	�Z�}��Bw(� �`Wf�$yr��6��Ǚ�H���D!��]��0�����g@Ѷ����A�7�D�d�Qȴ�3��.by���u={e��1PJv��L��a瑤f�2��o�8�N�^��R$K���4����c)p:���,UME`�F�E`�[!����������O�ɭT�'�띊.����@|��tz�$���ũ!��V�ZP��B4�N�+9^lr:i-j���f|���7����m��2�����5�1�c>,W)�M�C.���4�iT'����� bc�m��L��[}��.������(g����4[�̲{��
c'��25�"iײ��imI]2�6J�c�³�3�|8s��=���UC������L��˶F���<��6���^9O�\$���tT���HT�nU���ۖ�n@%���t�Nە<�g!�UF�����eɽr��RMv��Cy�a(�L{���)���	R�O_b$��*�?Z�)�j���ec�Í�ֲ-a��|��ɉ���?��$�Y?z�E�����7�
��:D�r��H1��L�6{��̒s�o��Ź�2�U��+�h�{,:������^z�rX�&������n$v)U_�9�kr=!�]��z��X/�
�7i�ͯ�"X�[B4�铡�{�課�T�[V��9E(8��;����b����dK���{��*$T
P�� �K��0b��dW�Ki÷aOGo�E�ԯ��3^�+u�BV��'��<Q�Ic��b���q�ھ�c�D�;_c��)auN,q�~[}f��L��7(ڍl��RM�%9�1�[2ylN�;f<���j��Æ�K��w��̞3����ۃ�����a�EV@y��CIJ�EV@�{F�Ѱ|$�f��rZ CQw	�6R�EÆ2D��f����^	����E�w@?�À��>����u�P޿�-���`jʯ>}�?
�N�k�mD�sS��Z5V �������qd�3������[:|�f�7d�ӣ �[��s�B��-�aǻ*������<I�Y�F>�[��PbQ��E��;����^���P]�F��?q��w��w6��������l��}��Lf�;�x�����X�k���10��h��H}	CU�s8D�e����L8Q�oq��~�.9Ç+�����FJD$�,�0E%^[Q�b���NC�NI��Ě��1�������݌S�|x1���$.��ŧ]�����X��_{}�ҵ۲�J����S�S#��kږ���bh����*�W��j�8��g�H���5��d�3"=�)�ob+����<��E���l$�6
 ?���\���ELM�E?b���_o����T��}��0�ls-�1U��?�U<1����d`�0�)�	54{�V;�i��Ԓ��>A�����mB�訡Vܥ��^�RZՠ?ֹ�*��4Đ�
��c�YJ����d��-̺�h˔��ßcM���E�|�`����+̪F29���#q��pٍ��#�4Q1F�q�9�MOS�f�_r����r9Oz7�^U��T��������7��C
�O<m��26���p��+P%s5,'|7�i�|��W�q�������b�������I��%�����M�=W�P�C���?-�&,LA�]���7��K���]�CU��7�K�֛<����֥��#E2��'Ɏ]�A!�!{U䙮��?��\1�L$�n�t�h��ȡ�36��8L���7T�\�l ���P�d@$�}����P�e��H�Ђ��yv��R"�Q������"����[�=D�T���b~�4t�4�Fs�z/��إR���Nx2�d�@��6��*Np:K�� c���jT�¿s��T�ՑV�o��o]�6�R�s3-�ߊ5�kI#n,��DQ+�4u��5jU�۬�ɟ�F��� �
k�T	~:�hu}��f�d+�O����`��1i!�/��'��°�S�3���D�m��58;<&M���I�i1�]�sf�H28Kg�ԁ%w���i.u�s!��`�/�z���N�4ʢ�DR��F������}<H�#
pZ�E���UMFS�mȺ��~9:9��-VJ�_]��h��dX�6�̍���ֻ���'�W�}��i��!w�Et\�m~�@���f�N��ւ�]'^��&bw�#���1�1��͵2->��#|��Pį�,Q�����b�q&g��]Y,�h�����Q(�[Kmh�ϨX�����.-�󾎠��[�^"0'���ue����kL�[*�4J����T R���8d<^5�$���"\���f4��1(?\��(%4Yg-Q�SN�����3�>�Yϸ޹5��D#��]��7�G�g�\~?f���ʼl>4 ko���ͬ�߉pܢw���m	z�H�Ƌ:]��1�e�����9������T�^�0��R�/�<��w���30|q�$���e��~�끨:#�����Y���`�&:@��Ć��}��{	^Xj��(A?��\-���Z��¤~����A@|�UNn~u�L���s��z���Vf�3�u�f��m<ȄdWA~�4�]y&������8� Pwz���8+c䊧��ysI�G.�����R�����pK �ʈm7��C?��	��Xւ��52�L����R[.T-7
U�l�U�ݦ�̞regq�h�����$$�~E;�/ːe���v�G�`��hC H����O�}�����N����t/��+�|s�r@���nٰ�S`a���0k~gШS�-L<���g�e���&s���SܲnJr7(��C6mM��_o��Z�N�����j��
�+�pP�Sۃ�T���V���)c��w"�ɶ��}�%8�|�A8�������RN��gI�)��m�?���q�k|���$���;��`�2�,f/ �3Ux=I�����>�>�1,+-0�1��7/�M\�N
�Bm5_��u;�n��cBox1|��M'�[��&�7���!T��߫�4�W�.�1(d����'-���J���zFB>�)��x-3W6�s� ����>��Xd�s����q�Uڬ�n��=7��TU���v.*C� D�����Ւ%ú w�]Pc02W{B���� E�����C�W�'|�R�)撾l+[�b�ؽF��K& /M�6����
?��+3�da���l��<�>\ރ�w�k��)0�
�����dۣ�B�n�NA���Xx=*E�w���ʼgД�?��:#�����G�=|��4=�����KQ��!���[�%�������'L}
a��C�G{���+{����$,���[�\�<��jw	��?�τ鿏��B�(J��tM�&���J���8�� ��"���o٧�<6+գH�:�͙T
�H�7.e��<�t�&fr�.O�9N�-|,�������\�ud�0�s`��[���c�.�4@�A;1��
�nƥ@�4��������!�?{k���
�n�����4��*����I���+Ns���<Y�^\HSq�L�@�ӊ8��K�C�����G��?yR��d-��+�d*����o���ZH]��-<�(%�8=�ʊ��������-e��Qa6Y'����?�tP|���Ɏⱃ3 (0���TZ�t��&r��δo�ϐ�M_�'R��jJ;rh;
A�tM��#�ð"o�hR6o��?���(�棗F�؅�?�s��Z�0
�G�,��u�Amv�Slֆs\)�2��M���i���@�ѐ��$G�7�>Jo�^��܄{~�OݮLgQ/U|m j��.2^-�?����mx,s���]ˬ����E>�'����	�����o$]�� fRԣ���p���M��{/=��IY�z�����-4���7Cj��U{�ɵ��Ndbf�������f�b:0�2Y�!�v�?�SB�Q�U���2�u�K�t���'!�tX�؊^�m�_�s���F�:���#��d�=������n�g����/�&Ĕ��*������P	3�zO λ��W�`�KB$��ߕ��(�l
U������A�����\|�s��C'�ݢ����Ϡ[����`%�TEY��RAf�����c� �q條T}CԴ�U���aj��W,�p����N�� ��*_�<�s���>�G���q=b�-�='7[|Ɇ1ԑzx.�P�9�ګ���v��׆�Rg����o�D��4��u2��Q{�g�_����3(�q��,�4���V���̨;\аmG;@��^��H�1���Z5^���f_�_ϝ��Z�Z-�A=� ���I��߾�}4�ND�c�%/�0����="��e:!�Q�BҚz�����ݧ�Ly���=rhd��+�x�~����M#H�f�;��,�G��r�>��JTw5TM[��*Ӝ�FG�q�(}�S�Ȉ��.�w�V��O��7�q_���tNJ�fm�Y�2*�jW�H���,v��=�����o�$��e��J+�[�Gu��އ#,��IY���\��'13�,���؟&7�� I���O
�9��<� ���E��v�W�l49A����Jܪ���-��� ��%���*L�'��r%c��.4� �Z��a	JI�zI��L�;���u��By�֟����'�/%�^�T'N���#;��g ����Dh�ja�8�*�&�n;~a5�0�b����N�����(��6�O����+1ă�D]��N�D.y��tY���C
|�u#NH~	�3"����>�}��#�M�����ƅo�IX>aI���u8 �:�~<�e���$�IS1�IC�}�ڇqpE4��~����c���yکʼ���e|�]���0c�(��p��Y3n4������a_� $D�q&޷��{�/��:�a�hLpV[�i1S� n*���Sp��P���0��D�R�@�R)^M0۝����(h��vs��u�-�\v�φ�Bb�b�_����n����B+:���U����b
K_3�ﲶ[v���iq�7�oKN�!� ���TYɜ�6�y� ���0���|q+�nބ̭�ԂI	x�#H�~L�3������莞Wd��G�
0�˶]\_B�WW�~G-����ޣ�z2��u��ѭ���]#���.�6�
�-�)�+���en���'�YƴY������.D�S�
���F;�d���,�B	Ø��ԫU":uipT4r�ݣq^��Ҽ�c�b�������ϱD|.�2ߑZ6�\�{fۙ@��u���FN�S206	?u<�ݔK�jd	Gm�U��K������������M�@��Wˠ���5�R��O���j�!@�4ҡq�c����?~n�`8�T턇�K��)��k�m�4�(U-�!!J�Z@�)�����HGuVڇ�#f鵠3=g��k~'��st����o?�q��
��'�֙DC���`��}q
�~Q#��fc�1J�0�Ѷ��a���--�ϻ�y��@�'�B�8u�L��?_Z��q���{�m�W��(�_ ��[��⤆ ���6��m�����?��ϳT��Ý���_��[���5��內�\C�y%��-5������]`+�� �H���Ȝc{���l
Bh�䗿iI��������c�£�#�]�K�}�t���)@U�4����uz��V70:&P�'��_�6,vw=Ԫ;����G����X�xn�b0>b�<��h��_[/vK�������lj����	\	����[�X5�MJ�j͓�2�Ww��x��d�u��K'�A^Z{'�N51�P�\�b��$QKź���?M�_��%���&����n�V'��4���Z�Lɲ[����^����!D���&+~��f�o.�j�IW�r�_��T�5�U��"mǠ���Rm�e#�P}��+H��w'��n�.9��������[w��.x���g_�1K~�^)q<6g�۟,�a��)R]�j���D��x�F+ ~��~z�z��9CG!Ԧ�og`R���D"?iG�4m
�����6�F%�UPe�;�?�.�D�����,��7v�\g��v���,�f�FV����|�a���3��t�$�;��D:s�:~C��u�4
DQ﮼�2�F�ʦ��q��$d�g�͵> 厁�m�K�Ra�km�,G��'���uslO�䜝�X�c\=�JD�g�'��]���bO'�7��6���=��8b'I����wa�IB$���gjx����46u��r��@ZB?=�����#cuS�� ������l35��$d�Tc�k����m���i�yW����[mq�����Ou�|���+�`�����8�"v������8��I�g�/n�@r�I��o704�{�о����[�K���=>�X�����vys5q$��k�sC�Θɶ�ua2��* Y��>�C*3f �)+�G��	 P�}�}݄_~BP�6@�axy0~Å�
QͶ�?�N�A��a���g�O3��Z�h��y���J�wb3���b��IzWZi\tY~�l���{�Ou�}{�T|���o�"w�"��G��Ð�/Zt����sm�o�-y��aJ>Q��/D{T̲ �H��)����!?�J'���U��L�佲�������TsÛ_����$��r$�#�����y[�:(tN?鲖�4�Rq��kE��	H����EZ����`�����bV�_�)t1��Ҽ"k�lH!bE�������ss�hL|3h$�k:x]ZA�R�5 ^0QXq�;`��\[)-
�1Y����5�B�{�&Y˷J�:K��?�u�DbNsE�ֵZVj5KJM1��d0����� |2��#���7�L�U�@@ß�'Ѧ�[���ܸ9��H�	ٜ�x�ޡ���m�Ed��P�k]�Wӧp�𵘇��	W�f;�9ŖA���P��j���L{�-��ۙ�Y^mи1|-�?]��<�ԑ�}���'���3 -
�z��E��%&�|���bm�S�Z���O����y�,mb$�nb=�M 8��%�:&*�1f֍!w�E�OpS[��r��-���Ad�XKmx�c�=�y��6WKB�F+ҩ�3,��(��C��=0P�U����ŃCU�e�¯��x�_�1	b�Z+1;�_��1[��j��ꀓf��-%��~rgJRp����3�/�Їiݡx�-�����a�a��*�a�t�����@��{�4ULA��B$�Fq6z~4�hV�T'�n+����8X� 9��k��PwJ�k�֯1���䡤�\I��E`J���BA��	=G��5�7]�!�s�F��wl�:�O�� �A�"������ApN@������@|�Yj�!ϥ��f�p� ���]a]��ChQzfl�@&��� �
�H�c"��:mye .0��D�1��lzE��^Ƌ�uߋ��K���v�T7����]c<�\Z����Z�s�����N�ѐ�8q5���b�=v��E�Q���5X�s����40;���w����o[��=��%�q�j��%�OZa'U�,>l�g�hQՁ.Q �V��ƫx�h�d^��$өGDC�4*�zq�8�u�"�3�����zǁ=y%����5������&i�=�T� #��۲Z�\6;�U��A߃��Ū��\/P�UVe�.������� ��[�-���}h\���b�ՀL����vc�[��G_ij�;φ�4>O*@*�6k�d6Z<`�������Dw�Q�=��t���4O�� #�����j��|�*�y~~��C7�8)�X�@M��)1�m�R(�U�D�E̗��o�KLy0)���jjF�/^��|��h4��Ǻ�(�H����	�{Y�:�3��,��=Q슦y����S$凌�������Z�B3Pc��L�͵�e\-!��7��$;�C�-u�Ŭ)8劮f�Jt�;n��,e��-� �SS�L��x��eK֢��cO��%%v��I��V�eu�_�Ԍ������"�]�*���ۖ�xwAb�;���|�c��g��%��Q�h���:f f�	�W6+-�(�-)��(��t���������2�,��H��^4?��~qjq�L���*������ \`�L����$�〔!P�E��	����`(̈́']�Lj��9�%�=�hE�e8T�	��n��[���T�\D�	(��?zs7lxJҫ�5;�+�x�:����f'�>O���AH���kK��5+K`��>
� ��\*� �$��H�2�8���Wm���W{l
lo�R��	��UR;�/N
#�|�x��۴ҏp䘟���c)G|��������x^J�rbm�9���I	���<���Oz�t�������z9�`�S&�����K�@[�qz8�|	�6ŞXB��@:[�.�6C���2]�T���1\�T���	�\G���t�oZ��y�b�C�ƾ�\Gy7���0y�:����Z%yk��+?�t��dG:'#������qjՃ���2�(����_�}����S�>p1-��xB相����E��+ɰ.��ͳ���rE�~um��k1�_Y?#ʻGቺ��.**�c4RO�34)ͪK&t���q�p>)�g��K�D��N��BsN�35�HO������7Iyk�Qw���<$Kς	�����7f�����4�
����R��vA�dY�L�����ٌ�݆;��+�x�S`}����X�KK*�KB�����C�vs�˾���Pö=>t]��{�C��웨�/0<D��Pו*�ll4ߗ?P�59�ܜ>���sr}�9��W簇+�}{[��$=7�/!~�3y����T��e�����@Rd�;��k�&���&���'<'��:���0Ff�(&��ԡK�w0��e����1z���_�EV5�Mp�]�	>9-�T��-egs"���F4��^�C(����=`z�	��eG1(�(���Ķ�R���Ho�@��G��ڐ��'P�Աi��p��vHY��T��-�����b���ȕ�%���^�:�K1����$U�m(�ñ)��4+F)<�4�uI��N^!�rITO`2jCM��%�c���Nη�A�����$�_؏�9��$��hmA���u��%�R�*G�7�զ�R ������7q��#�&v�$+�Ko�L23��lgF�9i8@�p��4����lp�
�]�ũ��1ƐǕ�tOg����{�y
m�e��)"���W
��*Q[<y����`f��];�0� ��5�ʘ���j2.�U�f��]o��ńi�<�|ο.�ׇd|���^P0y�xҞ;��%�D������	z�'�q��n���W���������,���*3�5���m��Փo�>���@�,���+�5���S�n!V���~��J��g}�ru
��1���aeͧ�Y�����ҩ��M:��Ĩ_�7)`�s(���Wy��0����{��ݔ6cSv�%�NZ�����.�L�ȝ�SNO���M��J�#w��˱�L��V� c�J�!��BC!"DDpҿf���i�~s�!��p�v���E�L��FCl�����0�d��~�]�i
���C�H�Z����3v9��/G�_P�/v6X��R\;��U]������w�D����O�F�MZD��<Rci��� R�XsS>�Ffo���$43T1W�8>�12����_���5�Ƭ��p�H�I����J�6��~��1G����Q��d�°�`��WaQ<ZO%��!>ގ�KhⰠܽ=~$��c��E����G�t���l3"(��Z��ɑ�
˳���$���G�����4�}�V�i�V�}�u�oC�8���$�XL���������k@�-��U�C^UG76�u�@yJ� �������6���Za�֕��z�C�U���g��#u�~�E��AjG�)�!�~���-�R�x"Ն�e�!5v�
�t��W=|�%�{��c���>�׋�����<�6��*�	M����"��nH���`�A�*l1|=�ӷ�9

�1�'݄,}pt�;r
+G�Fm_��;	������3���j��Ӏ:��hRd�ʉU�����grv�H��vq��`��5P$���`���%��pu�um�?2i]����a��>�I"2m�1��r�� ��dOrn�١Zi����u������Gq�rS�1*��h���iӚ������v녜��x���}�c���8+b�>A�p�7a(���z��I�eP�zp�	�Kq���AGh:�������Ηj��:�B�!1�C{���?,��}IX��cj�L����[w��B�0�,0uj�^Y���:{�g.Up���^��c���k�d�Ҥ˝@�9�m� ��#fͺ�3]�������ϫ�-J��OXr��@��O��	aY�F��(`��!���C��Ћ*	�i��u�b[�^�������3�$2���?%}�!�K7t��
￺;:b������5��� SU�;�]@�H��W����
w�o�ѷ�%�a71�"M�Z����&�rBZ�Da �����|*5@����	��eeW��g^�y!�#�A���a���<J?��/�J#���"�aP*�����b�2`�t�5E�٭A=�e�a'�1j��!�0�ݓ�V�F�r�qX4���gupD;�2�6: dd�5���ӛ���6!���}{IEP���;{c��rDѿݚ�X���_����n���tD��fc�@M�.�鐙]B�ޫdo�R8��aQD�	Pqmrk��<���O��B&����a��x��
��_�'歛��`��Z�]5NF���f�J�`�}X��IO������]���V+�@�?}������Y��	����<	8�~-��,lfI��%�j�i�|q��0ؾ	+:�WU������8��}���8��ҍz��,��T[���t���h��$I����X�qg�b�u�u,?�}T?.�Lܨ-�E �㪓n%��d8dd���FK�;0s�l���W�X�L}��3!��Ҍ���I��@M�t@s@�v�*"�y�\�����D�M戂������U�TŝP�i�a�z�f-Tu�j��e[5j��k4�z ��E�v:U�O��q�ֱr���{��)���*��4\�:�D^)��%dAhc$g�7��� �܉?��>����FטJ�[Օ�$�}T��-�?J(&�D7�]9 &�Y�.k�n����d��g
}yYG��j�Q�>1YN�|�Ǐ]q&����:��
=����ō��}��=��[�R�	|7
��ֶ�IWlOTb|g�U,�Md���
o��}��' A.m��bqM����F��Ͻ#�b,��X��d
�4�!����>؀��'r�^�ć��k�R���-�.��?C�^�-l�8�k�e�Z����;���8/�Sw=~S�A˨ұ�����]{,c�X��
�|�o�I�� o	�<gI9�o�+�؄(��O��i(�(M��� ksB��2�щ�BP�G�`;��da��������t�X2S�sV���m�a�ȹ���eOУ��u龴��О�!}`�6����.%�>i���{�p=*�E����<a���x?����<7����<G<o����C���ϙ���;EpAϛ;�W�?��f`�����/�<�g�FkQ�s�`�ym����V�6ݶ;�����x�'|3\tbG�h&���d�L�A��x�3�ꬣ�1�x�Ư���d��m��7gm8���h'��R^���i��w�&�X���D�����YY�c��iAjo*/2����I�*s=��a��y��z�AJ���~�HWp�����7#?ȗ��#2x�P��4_�G��:�k=�L�t=[�/wE�$�� ����p t�T�O�莦�F�2Fʬ��E��P�f2iucg�:ã��q(w6��C��Y����$�ʖ�Wn�<x�먱�^���4�%-�p��V(�����̑<�PXIt��y�s%�А��qܬ����%�z�5���F�A������Ɵ���kS��r���L�yMC��v�G"�LR�F^�q��u�U�m��gj��#�e�+���������a&��3t�qFss�����:���ǃ,��������W��w�`�2��Ԑ��nW,����@�lX�z#�ut�� ����n�Q�ɢL�Pϳj�p����'��V;��^p����(���ħk1?/��]qP��}�|�Ze`��T	}r�vN)"oc���Y ?�@ff�i7�  &�X�:�H�w�i��3��7C����9S���4�Y`/��1 �>��z��M��_1,���;Z}����BT0C���;�����(����qX"+�������I*�d4�G������F�g�U�G�D�ʚ��B�؞�ʼ\�>�
�1)�2l���2����'�0�"]�ز����ь)��)N��4�7QPX��M뤿C= ot��^������y!*�~!/Iq�}w�Ơ�$}u���#9�����x��|�)|$/`^JS1�c�� Gm��ꪒ�=���ӹ�����d$���
.2_�8�c�oYk�\Cq���)�wU�/L���(i�R�:s�8����AZ�o��#�tU��g祈7�)(޲!!�F/�7\�A��B�����ƹClJ��6T
@� ���f"F��:5-�A=V4m@�C�a�#�hI�WނS�`[X�����}p>���Ԥ/=9�9���� V�ڋ�$�`��4��^�b������2���g�Dvj���NS�0��Ub����,�F`��I��j�:��Yq��-̑�s��_rW��3b������ßF�3��/\q�z���֠	���"�\��rǤ��i�M[�1�% �g-;�E�>�����T�.٧[wؠT^���Ə�spϤ��'v��� +�O���r�l���A����ym��6�C�)���S	f*����X��\$��R׏(ɟV�ò�Ӑż�4���N�ۺ�49��vh�&��0@����~)Y��K1U��|U�K
��7���R0"a�8ׅ�|>�?&����վ(˾�C%����dʙ��u\I��F@"�����y=4�s��h���� @yIy��r2i%�`�]p<�/�����-{.��?��\_�ʃ�}�i2ł>Ÿ�8�k�$D��*��3�]C�!h�愈�1#I��^� �7�K�n��ʗ��!��k��ÅdV���+}�)�Ͷaq�=�"F���L���Y֓B���Ϡ�mG�B��B��Q�w2�z�fϾ*�3���:�}�<�N<.n�>�~"��g����^�U��CM�y)]�yʅy֗�k�lr�t�؃�|k��m�:�U���	�.���$�u���4�c|�V����a��l",�Z�)�$�}�����7��0Z�2�����	��$^?���Y�����3��m�gq^Nb�'2歶����}�%��	=��	��&����!�DF.6�N�dM[Ǜ�w)-�<�I�$b��.^+$�����Օ�;��_У.�-�ݨG�*Uk���_�����BjȠ>-*Fikv+����t����Q5��}<��ޖQ��`/i��P�U�B���3KR<��.QD�J�X��frm'=;�=1F�R�]��@�4��%�+~<ֻ[
���!��$��~PC��;+C�X�ت���DR�F��Y�|v�f���5��ٚWa#��خG���k�gl�X��ғoy���H^ZJXR�2:WjvY��y߂L���\Ĥm��05M��Lܹa�	/!$1��� �ݪ{������I�cj�r����t��p��;�1u�$����jtg�D��1Ɋo6��{Gfz����ou!���{R�Ru��9ij3�b������H�K�m3��. 2�:n(.\�P[p��d���R��RcҒ	-�9��rY�)�Zn�F�zoz+�l_�\Xa^(�']_adj�Y/����>�ؒN��������*K�;�N�0��S�܃�X�C#yU!r��\��h �̏���M�.�B��N2I�ݲ�����T�,;"�%Ҧ>����g�D�׵�\R<��\�Ӱ%m3�KC���!���va;��YM�����LK�C�=�W*�҇ nm�Z�����k�<RT!�F"��q���m�Q�%�A��D_��X�K+�f�M��_RB\�/��q�2�� �H}�T��QA�D��bM&�:�s`���{��L9���3Z:k�$�:P�B�`��v����l�ȇMKm5���|��r}�뽜���]Y?1٦��a�2��#�rO���V ��vA]��y�%ie����3#=p�|�Nw�(Ha��\�`������cϒ�B��o��^&Qy�����D<雳��Hݞh���o�-G�n'`����̊�2>1�
.��VV8Jعl}�w�nlj�vݽ]X��&��*�b�|2�Hn�hc}�1�W*Ǆ�(4��?6�����8��%����$4ǻض�A����7�@n�\<\zq'���ybWc+�g$Hmҟf<(�Ek��]:�v��	���?K9���j:�h;���#�BB;k�S]��l_�`�|=s�7d>Zs��՚v3��-jw)�3�1"�Ji��!"�=��Օ��h�=܇3���t�(J����F#�D�H�utZ���  0�u����>(<��F͝d��������]E���+!�����v��Du�vD$��\�ӊ��|H MO[�:��u̨/�n�na,��XePZ�������t�����	R��e���3��E�`��v�s,���6+d����2�і̟�[&g��]�P�cEE�P8Ӓ����"��/���6��P� �1}��r���~�� ���D��x�6�4c��;���%�o���shv�9�T�G�z��G�<v#���P�a��i�>F޺c��T?�Vqq���l���� ��hAL�Uf���|3���3�wJ�UuV�����\
�Z��l����w�X�C��/;B1�R�F���QMK��z7E�Џ2	s�a�Bf�e�����.I:����?�+"�7=1�63�At�!Hk��L�V�Gv�� ��PR��������8�(�]J#ǯ���C/��}�R�	�$�OU�{��g�3�����VSc6�%�}���l���ATVW<����x �D%:S1ӵ"�k�����`��4�t�gG���m->k.V1�ԙPK�uKt��[ɾHG�`S 2|�s6<����$��C�����l1|f�}!�cX��.��������,�ZG�#c�f�����l�P� �����z�+f'�֩�܍�p3�;��;ɛh5'7��g�*۝���#�x 5����Zt�Sd�!�ٸ�
�l���
�a	��5FK�U����҂,����Y�Q�_��#�7��$�<Q!����ܴ�Rz�oq`���xM4�#%���}��q͂���M�&m��ļ�f�{lb &�����άu���"�_ �Z<.��o����˅x�.�|Al���.���yաYt�БJ m=oA�]�D�+�_M��!m�r�"�A��¶$�S���2�3Z������R�f?�*T��+'�8�R @*	�,�<����[���4jB�*̡���lG�A��2�❼l�~|���5��N�9t�%�B����H�f>����<&(ː�#����FX~����g94G/���J�R d��mNQaX�6��"����G��<Q�-���&.�S�!96�RW��l�<Z�b�Yƹ���ë���rz��>�J?�?
M��*iʲg�-O:+k�('I�a��%��|��Tc���۳�=��Oux�A�ί��� ��NO ��~W�M�`�i�9S�"J���VOj�>�	�Q9��J}�v����
��8=|H]�_2��W��� '�A���巄�.i]�"Q�K#5q��6!��E^f
��ALRM��o�$7��B�"&�b�/���^wC�iP(6ė������B6�.3O�Ѵ��P����H�hO�r�ǔ*B�2�{��I��{|�� O9K-����%1��I|k��w��̪���s��a�����2g�E&���J؄���/���鞲c	J��� �zs����^�DBdet��f2.�`G��;򂼦<%���joA���bk�|j��ے�a��9��᭄�_��K.�XoBK4=~4����>����Q�X�I�wh�>O����Y�u������	��qZ�|�#W��R�������[#6z�g)AF�*��al�l�8:�RH��7k�*�)g�C��<��ds��/e{.pT6�2$��������?���dhƈAH�=�Z-yȱ����d{�)Tw6�?����[ѦԶ_�������u�)�e��(��Z�#���v~�J�9JE�"/�O�{�0��'4����#9y}p_X�>'c��J|� �����tH7�Q�Z���M�%g�+@1=XU��a:�G�;��J1��xa��Ɇ4��	���:/�?.�dx�+�V~*c^)P^d�صr#/c��rzI��A:.������� ��9k@�G̸�4>2�j� �]y���O� �\�����0�Ym�qh�T���/�[\�%�x�nS�K�b���~D�3ޜ4p�,�V,���XN�~R@If
=�E�`ol��?�|�tH�����Б^��I�Xyŕw����&�J*��&qƩ_����#�R�WP�x��V3����x�-)_�d��^�l3��^�`fP�~N���������4E��O~nz�+�-�Ki��\_�D�T	z'��Do�3�uXU4���{��_�Ep��qS��N�c0I��PuM	UC n�� F~cF��Oc�"����	ʇ��=�k{��v\Fch]��ى�o��\
~��r����o���k�/YB֑DB��͛�	�C��Ls�cu�^��{��e�D7 <�`���7O4R��`}L��oSj�O�C�XKt9&�y�guc���8�d�*g����7��v��aH���mYF��1H'�L�0�P�-u�RS�P���2<�#m���\Ss �1�Wv���3G�h��yQ���ik֌u�h?0�7<�	����y�/̫�����gR�����4�(�+��/M����)d�UT�kOf����С���6�<�|��2�u�Z
pC
���p��-�>	t�o�[�����vf����y��u-2��L���!2m���} ���@��T\R�q��tW'�V��@;���e�j\��N��3CK1�������w6��6d)���'6CO�X�G����;x6��G�->��9��ل���<��.�b\*�z��z����gg��g�<�+)����, V��nKNVy���N�cs¶C�|�Y%S�r���tз|z�ͩw�����b��㨱T��g;X+�f�>H����C�5/y+��3oӑ~I�������CfjiQ� m��
vT2H�k�yV��Ò��p0!oo��3�0��t���	>Շ(��g�> 8	M!�L�v�2F�-���E��x{����B�.�	���3����b�Ђ�O&�=����m�ҽFM0 >t��w��*�)#o���>Q�M��(1���{!���,��YO6ic,RB(��Io��/�#�ͮT�0s,&3Q��}�9Ԟ���1aY2-@'�6�����OG��i�󘓌�>�!b��	nݳ��-��yȧ��%���󧿉�ZJ .zM�����X���Z�pD�r�Ǚ!��s(N��oԽ����}kURz��r��]�;�VA�4R�>��`�|-�}U_�W��,�n���D��<�Svr��(�w~�<**��l��}8�I�h������J���׻��;�W"WS��@/�&�o��Da_D,j�Ɨ��-��'K�;e|���{�Z
�1s���ߠ+oW���<C���aW����H��Ktc8��h߮ه:��:Y�=9:���j��U����CC��Q���mn��X����[�jp8�e�/�q�Z���}q�3K��Cx�%�6�LL󊎟ݼ2\B�cSDܑ�7%�q���:R�]Č6��a��2�f�����^ofD>k��5����dj�����/�Smwl���A�қ�5)����R���r�v�)�°�yǸI`�Q)�H��r�U�W*o��Y�����y,[,������7�	͈��/lڗj*��Z@�#7�R�{]����d�� ;6`{ā���_�,�_�Q�y4�Sq�F�����L��K���U�[]:6#�G�Nh�q�
g���p?-���ι�_�L�${t�����d	�3�M{Kq	�孢G9t��i�/}�����ʐI}�k#)�wi6�S�˃�Eq~�.{_d&�$?&>�=0�a�箵B�`�y �b�Y46Ò��gx���[�lOvZ��ڪ�+����:�ZMC{���_|�%�H��#�a�sL)*� \Gg����"�P<v��^�}+�$P/�h0G]0EǍ�%m IW�6�;��M�5�֟2Oq��W����=��\8,���fI��6�6e�c=E�)���^��4f����/9=�K�RE��\�S��Ҭ���2�(L��=6P���l.�m��Ɵi�vF/q'yy��\Sy��L{�ɛR5���!Jُ�)�:��
�WB��l�W�z�@�8�%G/��d����5�����dKxb�аq<k���Q�zk��r�n�r�k#�Ƭ;�c���#X�������L�~2�.æz0�E�µ/��0���������jx��3q(]_�6��bm�rr��B03nΉ,j����A3�uG}f$:
ЖA�C˓ЛkS}�{IJ�
�^\C������BFI�j��L0�p�q�<%��P�q�t+7H�0��bd5���hߟ�@2.�j����e�V�'?�,j���Ɇӽ�O2$�]� ��i�y��RI�u�k��O�Ϧ�F�a�1e���@A���y��g���vo�X�`�	3��󈂖#51��ɀ�"�R됤�-��S����',���'�NWvB���{p�^БX�z����mcbؿ>vC�?G}�̕�+{)f$�a8+���m_�y�#U�t$S�"���*c�j��&Xy<Ֆ�`Y�7I�P	�n��n!`��<�+��]P}����gf<�t^�7u#�vxꂥǶ�'�ô썫�� �J�&8���|�#;�Y��W&T��a|��z-/�k80��w�p9�8������v�՜u��C�YFbXji�c�������[ac ӛ�4"�J�x�)�d$�ݑD�����0sL���h}?Z7 ֭Z�aڏ�ҋ�ה}���A��n��+ճ%h%�˼�ٟ��xI��d�G��#�'a����8W��9�ې׷ճ9��ɍ8��=�C0~t�$q��0���DQ�I�Q���:� OH�[1�?nC��N�L8��g{�����R��#�k�FtӲ��������ܥ�ު}�9�
g\��N��ä��ڠY��]�ࢿu%����$�M�!HCCeN���Ѫ	 j���*�r )w�i
�0 ���J�������#�7G�}
��X>t��`��y"2�Kz`�M^�Ŋ��H���v����$T���W���ަ�$���T-�l�n�X��5�5B�:��W�W����#��-1�Ȕ��'����z
��w�ٹ8{6
��%5�����v2�k +�C�1����[���������e�� ?�P�&/�b�@�#R�1v꧋Vyȴ�nc&*f����l��	<{lx��ģ�Y���j��B��N��"�iz�ǆW�q�B�{��տ�yYW����ʺ�)�Ar|��)i�Y"wPH�w��	��i?�/p7�l�H!����c/c�.��>;��g�~�C�3ش������Ψ#�)�)�����j-4&[��;�c�[� Av0n�6��#n���14�?<oS��]�	F�	ݿT9�˲��т�S�,i��5''����M�9����T�*k�_B{4�vW
H��Z�"��F�� `���2.����w0f�II95]aą"��0Z��hk�5g�K�:',�\��C@Q���}׭CTf֑8�D=/�cZem�0C��\z�ڭ���v�=>+A��7�-%�1�%�{�����Jm�Fɥ叇�Z��l01�i��(i`+�C�l�N�0 ����LĀ@�X�?	�Cԛ+�"�>XQ����}��e���)��#�g]�TŒ5��gw�j�y��x+�.�O��`�5�5�Jvf�4����R��Q���|K�Òt���4R�x7��ç���]\�\�hMN��[�`[f/�#ȅ-Ox�4���uiG*��{��e�`�1J�i�I�&ߛ�D�t�w�^�p��Ga�� �X����|vZ�)l�	�/�k<��0�J�u~k�"2�g�'���2+��nn@U|b�<�Dil}R:V����)'ş��#�a�C�S�����p�ː�q�P�ol��v�~ҹ!���(�,`~RxH}\z��S���J������.�چ���&����+z�������e�a�kƳ8��w:(�T���sJo�(�)�HtW������	qJW�V��!cps;���S��SH<�L՟n,�E;�'j4�5�D� ����9������o��<��������<�
��j�,�22���U�a�5'�eEdI��b�:�Z�h���򏫷�6Ti�c�������R��1��y7�չ���
N8;�~G�ز�ǁ���Mt#5MF����l��c�)�}Sn��x���m���j�r:��I�{E9��y?�@�aC��%�䓩˓�&bv�̀�z��y��O�4���ty����;#�ꎓ���!QE96����?)mt���Zɷ�U�QbD�A(vm/ٶ�U�����=)�%����,b}�^���qe�G��rh!�;aY=!y=�V�~��Z���"Z�Bj�&�SM(J��%h�G�u�I`� �Mv4zT��e�����N^�m����=�4]�F���̓pD���t��S�m����|M��%c~Բ+���^��U(��ş9)6_�<�mI|>R�e��,o0?o*��e>��(
v��3z�@��6���w�-(
6f^v%��_q�y��{e��C��՝P1H�y�l]��,%�_�k#��K�O8���U'3
E�/��	 ~����j9%��ѦF���w���0Z5��!Nڧ����H�Y��	�>lu>�sЁ�Qw��f���t��!�/�R`ZQ�1�?��A	�*��fs�z���\��I��c�Y4�[نq�a&1�-�����>��?��n��?]0*�O�Wګu��q���yhl��8�m��l';�[�!9���sU`�Tr����F(a[m!�U�Ñ�͡�(�2�2�n����E�I�����X���7��k�nuN�B���_T��h�:�����9ffC1^�/��62�8�=�� ٷ�6�����V���\��kĹ�����J|hq��0T�a4�O�f��ܮ���	.�n��'��a�#���qp�˸YS;T7���Fsͼ����n8��F��h$��P{^7��%�6��YhO*�ʈ̴q��;��h����*(��>�}rBDG�/y�_n �V�F|6�h��Â�}|���v��7g��E#��
q�϶8���p�ޥ��벳�����upfG�! �(!�`�c��d�,�D�n6��yWAj�0�?^� �U+4��2a�~k��eZV��އ>�8�G;�+�e6Ȫ)�P���sv]̥�i��~���uJN]��?;<�f�F,�0����q�c��!)R�=E��K�F���7h���r�'Pp)�{L@�1�cԖ�˘�:���UTlRI͚9"��H!0���H9&i:1' �����e���,Ev�B��B�R�~�.Y>q���+D���o�a]��;_�&�+W^���o��t�?�7�������y�ۿ�d�&	��{?�H L�WQx��	��Sj�@�[v��(�tu�RUE�\��U��Rn���NU�Ha>�,�����}�^|��/~Y�:z�4h�]4Eg�qG:��y�/KeL�1�+~�����D��AG���cdT�f9F�vZ�י
	r?>�\�����+���,�KN/�>v|D�*?�[��Z䓖��!����=��`9WO�Q��w������PTSn�S*ƥtb����~Z$T�"-a���g��3�or��^#�h-����ۑ���2��圃�0�BJ�-J�+I�"�v6�I�Ƃl�� � ��4A �����E؝�y]0�}rD��y��m���B$i�,��ۖ��������,$���w�f���]��`r��*5y �Z�ya!�|a�y���N��O�D=�����ŉ�eT)e~N!�$���ѥ�"&]?�L��>�	͔�r�����sґ:�:r��I44-�XC �a|k7qe�z�:�6�+��|��J\��	�	�N�u��9�k+MV}�#	b���	�BB��-�>i�h'���� �_�iK���'$��G�e��J5�)U�X����k*�����@�a1�7�K�eV�
4���}:HP�a����ژ��ΦV
�euS�$C�ҿ_q���k~k�F[s�++���W@��#QD��U�~�&ȕϗ�-
A����[f"`?V
|b�r�O��/�p����]'�y"V�m�,������+˄�q������r�=�g0-q�s���s���l�?�	������k0��A7f"�)�\"��
�ϲ��=����Nm��'��ߴ�H��=�g���d��ɁU�\�#��m�P�7ܽƮ_�JKw����sc�qE#�~)���z�p�z���4��>�uK �\��Z&#�:���5p ZU�cd�ɠ�Y��a4�0�yJ���=�1ݲ����"�S������=4�}�r��'l/<���o�(3`��)�~�
�����5['hem�8$+i� ֘�����XJ�O���`һ��D=p��'�\��x�w� uo���ׅ�V��9�J�/�띃=P�jA
`������h��?�g� d�ϟ5ø�U6`�l0�����E(ld3۽��U�$A�*�ҕ�SuI�ޙ^�6�K�"Ϭn�L��U�r��ꁕ
�;F)��sB�d���4��v,�4ֈGa�.A�X�~xv�Zl��냣�R����R|T�ؾ�IE�,��	
&�3g�4�"A�6��Z|�[=���1���up��1RhPj�v���?E�|���K�������]��B?%�M�M�?ǅ�����%���`�<�(����0����Ψ��%�U���㐴t�r��kT}y&.�a@Z,O>�A˲vxl�oQ8�mY������=N��i�(��C�4��� �a����D���%���$��Ңf�޷�zg@���}��z�ӑ���C��Z{��!,�;�֯�����G�].ȁ��s��c�7^q�L�W����S��+^�����;�\���3E�fG���0���f�W��	9�����+�HML��
�~��8�,�He����w��#��S������q�"JDVbs#�e'*����gG��I��؜�-��t�QI��?���	��mN��~Jn}�'
뢂�i�M��O�˪�=N�oD�u�� ";6�YV�pr�)����옰�����`�S{5��,=��/���M53�F��3%jD&��~�g��p��N�P�1m.!C&��5�|4j�@pfH��m{n�����v�!���o�-`��ܟ�>:��� ��h�����7O�o�G����*O`?FD1�9�v7���/t?8�\�@y���0��	i���6������y�E�O�LeRsc~R��4`#WN�j�N�d׊�S��?���q.�ׄ���$�[��O��������G��<�g(%)����c8��̘��0����8���`�D>��nU1��0h��oSbH<ާ��U�m+�:\j�Lp�z��~�����/u�z��	FY%�n��(���,q �-��r������!%=R��9}� �m|�>���Ҹ�Z�zX1�m�C?���q�B�Ւ��p��##Js�^Q�*V���Z����L�5���+߷����:"��i�d�/�ox���Q?0;�@�}������A��5L�I:Z�+�@�F�o��N�"�h��;�	9��(����
N���4����ۘ��r��s�i_��u�-eUY�6��i�U4�� ?|.�^on�ER�@`.����q$@�p�����LצQ�=e��Q�"V`<8s/j�����-�쾙���o�r�g��r�F�m�A���"!꟠�_&WyE��/s�O~��]=k�r{j����u��{��9�E�3�a��9B�G�6��ZG�{a����Xv�m��8��<�Y�*1���0T���n��m5c�U����:qv2{��:rP��]6cօ�]8��]Db'�\�w���58Q�o
����QB�2��QBơ}FȈԯI$ҋ_�gQ�ۇ����!���C�^�M���6���&���r�$��	����c��Y�J+�O�	6n	t�+2���_L�!-By�Nm=a�w�N�\Q/�E"�Ђ������F�*���RY �k��t���s�${�P�p��U�;�e:���PHBK��>��T��մ�3����L-�r���¨�}}���J)GB�v�+��V���8�񛙎!�Q�g��-���H>�h5�,s>��!���w��3R�{���w(j̡PO��;^/�b]������䨰�j��� ˧��[���T��o�H]���(`�o�G�t;TFO��	���gH���b��w�Z�!�~kd�4UOĠT�W���~%I�5p�Ki��]�j*t>�:�m�d^Tv����_|*����Hj:��Q�g�8��<\��	Of<�<U�$ҨCh*��)��?O�����k;~�z!�9)�) ��	hM��p`����=.����d��S�|&�wcAF�un���.kn��'�j��v�uo�P�Фͤ��Q�h�V;�XQ���3hj{lk*O�g������E��.l���Ln\YT��)-6�	��J{�	�]Cz+*��ٌs �bm��1�ѩ��jl�@rq�mT�	g_-�Q����0��Wb�:ms�����f��'�2:��\���X�رGڷ�>7N����l��J"������i8�G�B�ԬC��)m#�P��D�lQ�U��{>�e�e��O 6��b��n�(�<��cp�b��Dj�uMOoR$G�L�T�#XB?`i�B�k�uɲC��1��i�]� �S��t��1=<p�x�Igh�ʸ����j�����Y>s���qͷPe��|i��j	
|��[��_︋i ��dV v���A����悒�sm���tvf{�\��|ǑSZ�F���sq:QRMq�Ƌ�8Z!��ůG�69v�A�h�xVF;�h��>�x�g�d�7l� qaYְ�ж񱪲`����TBk*��C����~y�!Y������d�J&)L�L���u)d�O�'�j�Sd�WV)�*���(�sV?,�P������K.�<0�æz$��Z�� ����C��pȖl�.�R)��}��u�
`��"�-����T�W���p�F�Z
�!Or�)�w�7�)���LK��D�0u��hC�'�rԝ^��yF^Os�M�`���'�EP2�Z>y} )�a���6�P��`c-Ў^'�yH�s|��G%K��D�sq)�������%���F��)E���bivr%?�hyEk���iiW/H�����]m�V<�@�`{�{�|��X�3E��z�X�"������`��&,0��m����]�H�L�iޓD�4�i��^:B����zU��������'����w�7T�ˡVeˤH?�=����Fg���0T�zWX��j{{�~0��ĺ�_����w�:�.d�e�Z# ��U��M����/��u��v���[��L���P^�������`���T:;ܪ��/W�b	<O�RM�B��Hj�5���V׌7v@=Ï�F�7��8	5�f���5Ҵ�����OS��9g���)k%�R�	蠧\���
^�u��JJ����M�%Y��
ק �H�1L�:@�i��:��3�钠�X8Ru�m���D�5S/�Jx�[p�4��1�P��i�q�&%���2�8r�l:�㼪z�0MZ�/0��#'�^u�Dߡ�CB8$��"�fX��	���A;���Bc��a����B~3����t�B)a���?S�\�#�g�>�E`��J	��MNV��\k3���F�j�7����洫<�m�n�H|�N��	3�ۂ�(�k@�;
�T�ؼ(nxm��4y5L���#�6X\,�
�iT|�_��/�����d���o�/W����-�.`�xXK*$f��d9�3�ޝ^m�)��i��D�-��|����?Ӽ?�{�i9a
T�&+b��.a �Q����� ��kB$@�/����G���_Չa��;@h,ㄱ�}dx�BN��r�5���Jo�� �ӡ���������x��t,��ޝ�J��>n?4��r��(�9��S���>�%�#j���Zxs����ETw�k���?�?j_#�E->m?=bF���hSd�2�ɥr(������}gWӰv:f&�&k� ��N+��"^�WD�k*�.��7���I������z��뉙��߳�������_�M7�Y��cq���I��q<���y����?	�S��/���h霚�C��
r)iI_L�D��ɷ!s���̺Bw�r�ƛW�[|��0��M&��ò��!��8p�A�K�����:��*ƴ%���Kc��`�h����+�U'��G� 륈I�����m/��G��f�=G��,)aHO{��[��]4�����	�b����M����ꗜ����c@��r-C����Q:;��{��ꢗ9�{�	o���'z,�1Vq�i�"�~����#�y[ zgt0
�A�LJ,��a(��;���6څ'���'�88�*��_�0�!�n4�l�T�،�.^DU���W.f�:��|?Y�_�=��u���Iv�9��n�s|�
X^~��M�z�p�P�I�M�K�PJ4���k�S�ũ&o����,mv���>��6N�$�_�����bZ�V<��F�N}A�E�����tO
m0��RI|��A唼�������u�;P�/���2�RdX������#]����;�����ޝ��i黀�)P�+n�w.a�0D��fSљK��YWD��9�T���T�#I�HϓK6O����rL���n����	�(h�az�x/�"O�Ծћ�+dT僶J��RW��������h��(�q����p�ɬm�+
?[���-	���&����[�b��0dbR���>����o`I/_�b�͜�=X��yS�C���俼� ��Fg:)�D�x��:��O<�����1��ʒMgq~��EzW5=��<��1�|U�	��i�k����>�QEc�2����0.�N 3{��dߩI8���z/F2��q��^�[�RN����h����>C29�G�_�k��I&�39�x��z�I������O�n�])�U�R�%�ڊ9jQ�$��C��q73u��-�sG>�`�n������~B;aB5�{��v�U�����ť��T҄�Ɓ�+�w����$3<*��Z�%�~ֵ����)�>H����t��b��}�#K�_i�X�;�z5Ss]���\�e!�;���XX*��+�5��>��mq�UF|C����\R�/�(,-���I�7v�S�p~e�S�O��ѥ�NrD�������FEI�f����ޘ9 f�1C��vD�ܬ�sƯ}|��H��J�1y>1qW�s$��Jh��q����#ϟ�o�Y�ԍ0Ty�K=�	3�ǥ�T�*�Av`�xK(�9�����0�ٳ'�Z�8lF������x�gI2�^�3.�X�2=��-�{����'�rC����f����2"���v6��J���sR����>O�dQ�j��p��_�t������Ӱ�Z8�T��\PY��T��crZ%B�y��=���.�l �TO���x�����xc{p�i�(;��2�/L;�fNiY9��3��^M��#���-6��ԇ��@�{����Bp4��z���X_1�]�%��cf1�aD6?��[�Q�x���;)�?H�%�6YoDa2Ldby��չ�U��/Wck/Jf@���8��/���eVf��; 8���al��oi�~�F�!V��	`���N���;�H��`(�BhQ�q�	$g�������~P����"9�6���� i���A�d�x`i|1q�e��3�ڳ�.S��\�o�����!��Ҷ1z��/)?��.C�zp6�z�JL T�n}Ւ��<�e��?+�
נ�����4E�L���vԁJ�-Ŕ��XLkZ�S~dL�<����h2�t���e���f-��#7�#}h��LϘ���uF���ɮ����H}���Q�<ݑ}�o��V�ኮX� �cͦ��������'���r$g��`K[��(��V	j<�J\��F�$p��3�uP�৏P�1,}29t����|��|H��S�\� ('����[w�7.�ΚҺ��⢗�fàg����?Y�,w��n
��%�8���|*�~��Z�::����D+��]a���'5�M5���ŇW���kWi���'���>T����n^CH��-x?�[���M�����1�P^�ǵ�����a��0E�c�}E��u�Q��QM�x$R��?3\��#{���)ޅؚvѱ���s�5�#:">��%�g�J#r�o��ozX˝v�tw�Hr�Q[���,�嚄��9� ��0_
�&��xAe��5�C^������3eH��Q�>�#R���Q��a���z�ݗ4^�T�W�I����jgA�b�8'�?R�^c�&�#���J�W'u�JL� �7��cײ0j��S6[�1=���|�p��'��;DMO`L+Ĭ��T�?��tz�B }�G ϥ�R�o;�H|A
�}�p��[�3@ע80�$ ���u�$�w8�{��K��^��q�}� at1�ͻ��v%��C���)����Z� J�C�s��J^g�$K��0�� ${	|��Gx�C�:�ـt�6y�(X�m}��R�Ԝо���/-ߛH�O���ʡ��y7!x��,�Z&�J����ǂ������?U��h�Fe���.�����>{��Ԡ�F�[�2E����z�,6/8B��ė�,'Uc D{�^���*1�Ho\:�2b�������V��5���	9-m��3߿�ma�b����&577�Ih�kW	ژ
��n%SaC>_�@���O:�G]x���ƕ��G�����(�0����h�$3� ٚ�7|˼��n�Z��2I$/QUt��Hcb�����b3����l���t�GA��dɌ��DV~�Byݠk��Lb,-�Gۅ=�T;���gu��E$p�k��̏%����ޕ�JgMd!z�[��<��bn�4O�t]pL؄�{���,�X�\I��?��Ǚ"xi�Mu�[�_fUu��A�8:/H����0JX�c�����t��Z�;oђz'�^��TP��^� 9����j������HT�J0/�:�� ��$ym��!�j��R��⢬�M}�3Q,$�� �5I�h�7|�<��T���s��m��sÎ��\6��i���N����(������it߻�M�y;CU��9t�M�d��#�;��-�zD�N@:�u(�O�Ы�D�9R�Ъ�~�&�t�yh��+�#+�^.Юo�R����z���Oe_�$F���(��9�7ߪ�p��QS�TH��Қ�)�v���Q!�Ve��@�~_���l�%-����$�m�f"��uB���/�c�7��)�w��puգ=��a�0�౱�r�p��>m	��b̌��P�m$��H�L����N�3ξ�C�r�wre���K�PR��,
	pյur})r'
��N�y���I+����%Y��RM��5���Z۸�i%߂��"DM�?������Mo�q9��I5�]Ȍ2�$���f5��uF'�`�?�
4��4�܆0]��O��6
��\�Dԟ'I��|����ġ1��H0�!�pb?܊�m��0����y��Z8���JR��m��������gʑ_��R'��4�Z�V���+ 'Ɨ���v��/(<��uc��'h^3����	2����|/6 T�o����d���N5�9Y��3��b[iv�$�M��Fv��Nr�9�~2
[���;]���ͧ��,<���[��j�hQZ{:�j���R�h���}]&�F2_�y���Og����D�^����ɗ��y��<�Y��M	�o��)&�j��?�����uV�޹$ �}�Ͱ��2�Qs&]�p�[�������I�wP ���P�<�,⡔��9�ڴc�2�c�'J�Κ�W�S�WYNJ�3R ?9���-n��d����,�'i�:�^j�y*��_u����g�GD��~Ed�����N�����>�
���˯�DF�X�rxk�(�Sk#��t#�.g��!I&��M����|�m�iNKn���@�]���e�"#��1tX;�x_��% �03��_YU܅	*��˘o�-w2Z��֑6��n8��PdyT�V&s� �;�'0C�6PP^�-�R��`8��]Fq��S.���8#�w�Rׂok��~<�Dw�B���POE4�%ݶߜ|.���T�,J�/�)��|�I����6_,U�P󃩴ԁ@i�e�bQ���՟+�Z	y�j�O�^J��n.Ok����`l�*�'o�+�x%u�<��}���OҔ����Rگ���LB�J��p�\��z+r?�����3�C�=&�^7���UjR���̂)�{*�����a������W�Q�R��yѯ#O�zm��q�d"�@�Sؿ���b��=Z��w��ʨ�8��b^�%��+�K��n�Kf�����!��n_��YD��k�h�ƕ��'�H�����l��9��<<%iq���
6�������M��cm�D�8�~���Ժ�N�H����??"D'Y�$�q���h�h�j���@W(��ݭH�yJM�L��ӉDW�f�F��Tt��ȶ��B�����c�����f�ȯ���ȜJ	G:���3�Y�� ��ѹ����(f�������v,��.��R���_t�&I��(Y��=�ZG�D��@��H5u�h���#�qQ��T0���!eQ�:~s�%H�x���(,ڕ3�@���@9߁�3��8�+�s�"1�<F��hN�<嫈Ԓ@zV��tf��t:�k���ǩ�1�������`nMS�k��L8E��]]A�I)BJ��~n������p�G�s.�����	cK�ڞ=�Q���hԺ�z�x�'��:KAF�Φ�G*�QCz���&%��!¤��O�4�z��@;s���x�m��w��YR�2����Iz<]/CE�.��K�}1�dm<����VQ�Z^�#��m�lcW�M�w��s]�P��A�[�ƭU�q5�j�]��\:������5⭰p2�\3$~1���OO��)��Tm!�AV۞Y=]���!�=��z���;޴s��0?d����Ŏ�+��\/�;�E=~��������?sx,*�;r;$u6��؎]�;��\ܓq�<CFt��/�M�w@��������h�=��
�+vYz�c�Q�z�/P��@�lm�A��j+u��ת8'�$r����� t�P�P%�M>ɛ�@����&�W|��cmi��܌$���lduy!�l��	�Ǥ��͓��4�3�82�ذ_a����C�E���Ȩ���;��k�����M���{��k,Ѥ��w�㛌!�**�|�b>H��#w{��.���e�t��D�LB�~������-�/��#�HE
��,����Bkǥ01Γj�p
tR�`M���>G5��UiaL�J����W�p%
0���_�i7i>V@����P��$[3T�IGx�8L�)�t'P�N������OڲY�M9(�����Sl�n���2l_SL�1RႩv���aH�7`���$����/���T�%�@O�jlw���
f��VM��>�\ט���m�� O����k����5��~�J��� [�F�&��̙=8�*h� ���Ӄ���]�M�����Xj#�/���:^X)�p���+Z�0\��,�_9��9sl�[�}�S����H�<M��v����36�{k�W$H�kW:"a16g:�w(����4�v�=R���m�Pm���Y�-b(/W��Qd|u�ʁ�I�
��<��8�TE�{��VwX�fK��7��@@�����zi<iKx_��F��~�݊Z�иa~ޣ�����,G����z��.e���*c��|�jE>�L��ÖK�I_�aB�х�5��(�	T�"� J��*)p>m&:"Rv��0�pf�&oevB����P	�/\�Y��ug,h���E ���z�r�K_��eW�6G��c?~���W���5$�0���ר� L�u�cI^�
nh�J��� X�d��"aBW+��
�j倖{���X@bMXr�݇'�sj�� �6�r��[�;Ug�j�]p�b���2��e%.k6�P�o�g���7:ק/�MdDD�'8�{u�x	�n�����N�0��q��,�'h�
O���;X:nEC*��f&h^KaL����ܞ�G�����vÉ/^�����ox�R��h-�Á�1�uqf:��Q�ǿ��\�G!א��ac!�Ўݷ�_�����ԑ�@��?\(X�>��:?�&��
�Y�*{O�]�3CX#>�
�Y��l�}j R%��\�E6h-�Jw��J���A�	�/'�5���:���v�H�'��aryْ�뇼���WnpS�gZ1���u�M�L���ұ���k��]�-꩑���b+����Ǿ5~:�;���`a7��n`K|a@����3 (��S]�!�埞�^��(d���a�:��Gey�d�<{�Mr��s �D][	�雔�����x���t�԰�d�ɑ��T����#'0�֠m���(��<F<<{Mv��<ڊ��ߘ�#��lo8lr�V�=VQ"�,�*��'��[*�5ꡟb:��=ۖ���2�t�;��AG�t�|��.![3�m"���ٿ4�3eқ٬c��1�mg5���?2�2Z#A��F��E!���7^߷���^��h.K�P�v 7.�Z������#O���D�(Y�-]�-�{�z)/3̂ {za������������w��P��S����A?�~�(��ڦ��h7�%��p�m����F`>��a���aB3���pJ9A+�Z&6R^�%Ѡ���Ujm��{{�������2ӧZ���/�~�"I�'�T��[0V���R�ٝ*`�L�l�B{Ä��&��$��sP����'w�~�u�e�j�Rĕ�0|�ҳĪ�"���c;I���=�0g��2#Hp�Yۃ�M�ޅ��{E6�q>W1��.}!�8ߴ+Ef�#�`y�����&x^N{�f�@;"\{����A��c@e�p1�Z�~.�BT�*�b'��!�j�n�2�]Q,QM
�.a4�Y\Nx�1�DT������dsRF�
�B�ޚL\��q��� �����Gt8�`!�n�l����(�6�W�$�˓�Z�2[��6uRګ
nď������G��+�(p�U���ﵗo�a��]�t5t��Orށt��}5 ����!��Ɉ

{��ƮY�0ۉҙVm�{;[�B=�� ��+��0�p2���O���i�\��lr<�W:�^m�ڮ��<ި� 6���������M�_�X`����m�]t����S�N��g+;ʪ�l���}��˚�zs��q-$��`�I�����ĵ��KD��4��H�q`-ݸ?� &`�Z	��Kݩ��&(�|N]*2�v.=��M����V�p'ٹ&߀�n�NQk �����K��z.D�B�2�_�4T&���N��J�͢P���``j]�}rA�ũ.���~1�l��C�۷�N�O����ڇ�w�:���ׯ3	�D�Y3s9����yl���b�,�,S.N2�kh�����|r�\�n�nz�Eߥw�R_�L� 
�}��=��j�%�v��G�@�:���I �n-���Iż8���6P+�>CG�䉲�}#���)��SS]Pq2��sP:/N��|q��󸻣cg*پ����FL���s�O;r�Ģ��5�s{"�4Y�L��l��.j�v64cY͜^�(m���@p����o�2�����tt��q�05�21b��tꄹB�؁Ɠ糉:Ǻd'A?d�oiE|X�<%e�
�l���;oЧ,C)�p�$j�����ڸj4�$e}P;��A'��l<P��v��$�qDh��Z�ê�G�&��x��"��|�v�������(6����eq�A�8|��PT`��2�E*i���r<��S���Bt��?'\N��b�	B�V2�W9��,ED��zH�7�:��_l�D��#1.+�Tџ/t�X�_�90W�l�c�ȈL:�ڏ8<u��J.���G�ȩ�YK��eT9��F0��l{�Q�D��)G�qwl��5Kɿ-�����/%4�$��O|?���;�E0�E�6H;v7w�)�J#�,��9EC=�*�f�U���_h���(��Ga�7���o�(Ij�؂�����3��A�� q=�v��L�I�Q���:.����ރ�=�  �.�q����R�:н������C�9bq�i��o���X��E&�Ir�SW�F���;ga�U�3y}��Fބ���R����q��c�w��Č�Mt��=��'���zL�~ɴ"����o����=~���c���e�5���������&��y�s��bX3P�aoB�f�~�~Nivzaү���m�`�އ0����������[cAZ��R>b?���!��7��l,�m	�Y"�o���VF�j�.�a댔�8Zg�s�p�]R��E n ^}�z��@��E�zw@l��xN�'B϶$Rn%Q`��L<7�A�M2?]!�*��e�r���f��1!+��+���?#؋�^)���Y����ш���6�x��;c�R���?�)����{#{8�N�n��N����Z4��%���.���Ղ1�N�`#ꋳO�L�l��{�i�� 4���!��10�����XK�g�tܜ�E����Y�r_0�g��T\ $�a��(���ME�Һ����ک���SV)y����E�fd
^ʶ�c
x5���v�:䠂3_vl�U�h����ez�!9Es�kGxຖ�]jqq!�	�+�s����!ΰ&�H�ה7�=����t��F\�ֳc��<�X�+��=���0<���r��� ����"S�I�c> {�R�%����G��t4�9T���)�'P�6�� H�2P�a5pE��z��võ�(lͺ ¡a�+�W{��4+�a�G �A�^�2Z��1i���s�9,jq���P,��%^=�]����p��X����Styg���P�U
��2$9�:n����.���K�U� Y���2aP.Gv�C��Rù�L��$M�$^���R���X��rd��r��؉c��S��O���t�/dR��v
�Dߍ�0��t�SĆ�VY��T���zes(�zGQ�Ԭ��F��g�S]mxdѤt�
��;b��3@���W�ģ���ꊊ��$�ѯ�1uo��
��a1�-� 	X3˱����t����遢C!T�+���Q����>��u*�+��dl�x'�Њ`rP� s.0Oϧ��������Ff���T9V�&)�(�ƥOH�z+���w��8G�:��>+��wʚt�ۍ
�D�r
��ڤX/aY��^������Ȝ�x���a��;�y�R���_� q����B���B���-��� 6%+	y |(���jU��v.H�����$��W~;�W�?��m:�L��+��,�y�P�}}�[=笽,|!F�x�f�a��@s��C���Y!xh��cB;���Aj�;E��^���G����x�A�)�uR<KVO�c��<�<[��h=)�ן/I%��[��+�ݩ��\�~>�f�"��l�lB�Aܔ(�(�	���s���x������T�u����p0��@��|���BtVit�Z%^Q�{<��㎲�N��}(Ɲ\?~!����״5���:�y�Q��$���^yn���2p�_F)q�l)�s�&�o-�����{sg\����Jk�:����S"F�����.
(v�X�	�0�d�uk�I�����e�M���ץ
��#��3(���Ɇ�C;[���5��1���#C@r������!��FKW�;!�6TT������*���=#�s�q>���������f0�f��@b*(�1�q��݄��z�	N�;P9��p�Γ��[��-���H�.�oR�ڢ=|+��D�R����$3�C^�0�ԇH����]U�f��k���X\C^��TQ�a����ڥ8�ǷK�AJL��3{���I�a��a�/����/����w!���2{���k���x�W����f�Ӆ�^x�S�v���ԆG�/C |1���N*m3�xv �cu�����!e0k:Nn)���e�c�-�:�!��B+.[z~��u(��A7ܟ�o�v���s��[�ϭ�b�7�_�@B����?Α�)�X?󨕳�%���솰����B�D ����i{)9s��{h���6�'�ҸK![�~�d�4�
�����e�9n�5c3c��Ɓ�dZu�u�A�U��f�^5�r�'e7�=g��F't�=������uJl�8$h4d�+��̠H3/�.t��sy; �����4���D��V5c*�(�Ś�Ӌ�C>��
�rP�d�,�� �[�֦%q��|����k�4a��D�y���tKԡ��<���+�უ��g����7��͊O��2bPDO�e��O�g6a���*�π\aSSՒ��m����f2t��X,�n-�_a��k�U-I����VM�;t,B�G�Z��d��L``�%�2ח5k܆=@�}�Uj�ou쾨R�S��h�|	�ru���-H��yi����e9�췞�'F�[���ܓ�]DrM�ZLh��u���bM�7v�l;,$>۝�`����3�� C������"Rڟ	��:����윩��v���iv�yZ8��+�Ϸ�-��������0>�S�r!��FH�D���}+&h���k�iVu�S�Ip*®�����s�'ę�`�T�	P���%お1k�gzx ��.��O�d�5�4�����ˮ����T��,�U�%�?)^�L��ݦ�5��E��&׾�?�T�!��������{Ɖ߿��ՑD������~��Ӊ@�H���=h��Ĕ�9�|��I-WT��u������zv�~��X��f�\)���F�~j������M6��<0Eafw�|v�y�Eܒ���$8�6]tl,I��/N.�ъ�n��V��U�h{����M\��,�% �D6�_��H�2ib�_�T�љ�$	��[S�K1�J��;�����$�Y ��4P��QuÙ��w�Yc)ލL���9���\ ��2Q	��G<��B`�e����*}b�Q*�	�qީ's������b����ˉky��}�3]|��
9;�cc��C6״Y�Q����6~V�o��a���3���������o�>�o)�&��2f��R���%�A$���&��>��]��5�bHv�����Įմ.zYj����/���D|̴nbҹ�)l��>
�NojP�7�y?�2��v"9�L�F݊x�����q	 �{��pxٴ�I ��Z��ڡhU��ܖ�I�y�M�&�����e�fJ�D���MrZӿ|YBgp���o`���?�DQ�Қ����N0�Je�1���ПP{5;;�(R
�^�;�6Ok����}���!#J�h^�����y���O��8�j����^��KUmt�gQ; �fr��PFXM�܂��߾4`�&�ꨑ�n�~�z�9̪��o�U#�#�X�T���F0�FH!bG���-]x����#{��K����A�#׸�O����e�GD���~OX��H^���d�85\^�6�)��qT� �
�1����;6�)�D��^�9��<]r��A��/��|���L�b2.��M�S?��Kǣ�X:���i+��u�m��}���47@��%eC?��y�g�WL��S(������5�I��ʳ�.�}�Ki�����׵���N
��5��l.�C�rśL7D�{
��r���ӥ�O�l�q1��w|�G�6X5�Hª=j���3c����������J\�%Ϝ�.��~^�����3}���BO����$���J �&\����;5��Q�����2̑��&�W�ixD��|�JJ䖌�6�Or��_S��b!Z�����O���y��r�7�*��Jw��GL?�j^\���o��?�(XD=�r���N)��v��
댫yo���k�7��\b�H����y�>GLe[/�I�'Xy��R
cyn�2 ��
�.����ȋ�{ ���Me�_g�b]]�yl��᱕4�A�*�[)	�L����k!���.��^j�}�է([2An·��R'9����c ��^�\�o.�Pܢ�f��g�AQ�DK(��x�\p�A�p�Y����J,i2t/�$�y�ǹ��E��˯9�-�8(ճ�%>�ɝhU.��`�]e�=ߟ��vR�cd�!����t| ����[p�GhO0�.��.c�I�?tO(LjT�óLt��ػ���'�cg:�a����pt�F9�is#�g�=��*��eѫ��K���%�ųc�+t2b�2(��to��GCC��N��Io,BCstB������7R��� �<V��vj�&����<�
�h��PД���)��@�c*pH��&+ǆ�ŷ֜Q����z��v9����A������ɕaVW�Q�z�ٰ;r>"�r���h���_k�A�Fg]5F]���4	����-��V��m��CΡ<�5����DK��^�r�H����}@g�B��T�$���tl����,r������O+XϨ(�_����J&�+�݀���Fs��9֦&�o΋"*l`� aPh#9B2��9��nK�Zm�v����A8��<��ƴ�(S9�:\d!�};�Ar���vb+��Ff�?����Q��(��4\aP��(1bt��q�Z��t�AA��/�i�s��z74	�
�<��nW�]rPۈ���S��kU�~aB)�C���D>���$���V���ֶJ����,�G܋��z���Y�y��k;����"��L��rU�{������H��*�6�y)�5����O�P�4�4~';ȯi@��6����k��`�(s�PŤěk���uʂNwښt4e�b3����>�Q�z���h?w�M�1�Q��Vj$������ �Љe�~��O	[˵211}'�t�+�@,Jx |��0��o�X,[k%{���e߂���gw��w%�4
)���_��(��*�|�t#��e7�T����iS������w�Pp̷Cװ��j��R�����<�yEM��&
�ÚY��u���2�Y����:��^��ۑ���Є�Uc�	�I��\�+�B���<�Y9��kOHN ������tiM�Ieq%x埜,�2( c3���U�ԝ���3�{����(;�9޿YPi��j	�9K:�3c����''bQ��E��;J��k �WAy�u�.	P� ���l[�$f!3p0h,��^�[����z��ѹ=�b��F�b��2��1����mJS����P�6O��ߣ���*���,�-=J?.�w�U��p��EJK�`N��*��q�"��ဍdW��'��ǃ�n�l���dll����F$w���]���"���V{s�vd�P�zf�2�zޑ1Y(9<.�������1|���O3����W�o�Pn��HX�p7^kP6R������o���]��vlCd����[���I8w]9���MeOz39o���'_(�u>���B��`�Ћ;:�M�l)�?cѮ����j���p��ߦd�di���F�V�
3�P� �M�a8���u�����5��'��]x)�7۵tO��ն��A�t:��q8�=��B`-��ǁ��;��3	�4��N�v�}Q�&��Y����a{�J�����l����,a�O�����R��~L��P4T���ϛ<�p��%#S֧��T�L���
X5�^ΘnʖH&֒�r0�#X|��S�n�h��;d�W�%�b�C���)�\�K��U4����Y#��Z|���b��R��>���M'��fF���]+o��4��vYU������%�2�P�dr�}�s��1Z.����#��kB}s���fhN5UY�W���ڦ-O����c�2t������l�"�ﰘ��P5G凪��rl2�Дqԉ��ݗH?��b��]�� \�㦡��-*~��eZ8����\��7W�Ң�P�5L��ܭ��2���9��&[���������>�xTy�`��Z�W�`��Y�_����|Y�dU j�A
�H���*4ǐO�<�s\܄o!9�yՀ�xX��#����
]o��^|>c)���2��VhK5d7���N8�qfjz?�~�=�9�¬aVϪ!�����hOX�zS��2�f6J+_x�>�R��
Rf�B;;ok�$�T�3�:�Q�4�Z�x�q���E�b�3J����>6B���J���O��s ��Y��KB} �cMt��������������0ØP��P�.��!�L����^�3���seP��'g�S$Se��K���ej>�tҠ�nr��/�
P�W��A4�g9��kv1�Ts%_���g�IJ�h���7;��i���z
8J�<�$3^��K+m2�\j��J{�Ԁ��ZS��6
�{c�홑oXCLY`�Q��z3<��]w�E�+��x��i_���D�Y�� �B�&D���'Ǖ��C�?t:\�]d�M����B�&��� ����[����d�Yτ��ݣ�Z�	�}�w <i��6��~��P��2�I�|��y҄�d����X��
�<l���I�k�զ.}�����B"#6V�h��n|�LjI�9u�@p�^�����;I<� '�zw�<��y*k~�ty��-Է,9����oHC����Y��h둂�-��V����qۏ�[4�{�+���b��o#�Q@y�o梛��Bun�=���J��E��qj�#�ĩ'�6WRv4_�HI��\غz{��H%:�[�1E��l�={�o��!����.U��G&��w�un|%K�T"�.�0�&��>O	#v�$6�5;��v�N���q��]h/3��{$�f�U5�����	����u��ܡڴQ��8µ���7�+S���������;E�́h��l�_&�i{�]k�O��1��W,tH��\8{��R�Ϊ����={Ǡ��V�'v�'�T��i7���N�QP�
7&�m�ն��y"c�w�r���ޛX^��_A㱴)V��|k����&�D\�J�'��h���X��۩�e$��R�-E�`\z�Ɣ}�Z��Òl�s��U"����)[	'���WPs�f���So^�ҷ/�ql'�"_s�\q�ӷ���.�	�>Qup�#"t��I���$�D/N�\�T�-x�b(�B�^r�?8�k��bL�Z�5�@΂�,��S�(�����"1+q���nw5$���s����3�uwG�i[��ǫ9/P�5@����u�7��I5Ä)"Y@���p��'��(�8�'u ��P�j��n�C�A�&,�7��T�V�����#�b���2�����!F,g���]���X;
�Q���wGe�ma}'�Q�;+=NnV�f�8G+Y1`2�$Q�������k���*��;~�Q�SJ'u5�
Ѫ駝E����t
ã�C�T5��қ��/UR#_V��5#1u��l�ו��ж=P���#5dD�\:���r���\c�������#��6��֝�~�P|p�(��}��B�˒�$���� ���<�8�����A���t�� �	`&�����#/G c��JiHQ�����R�B=��1r?�1I�����GOۨc';��{��j?�1�4_��Lz�z��
0lԳ6Q,[��p1g
���#9U����%\J�7�J|�B?K��J�"6J��������)�N��o��j�҃س�NG��qvmR��"�=���`�UKt�_�B��6d�?x997N�%lub���]���`m$%#��e!,���P����%s.
��pB7{���x��H2-�uG0��5*^AI�3�k#+~FK֣��T�M�܂�t�Y�Ҡ���]F#a%Y�̔/�T��egk��m8|�?8&G�Q��#���e�)���_��]̏03��L�~�v1_ܣm;��Y�-������2�cg�0J\7��2Z��I��v�U�������@)�����p�5(鑌��Gk�C�$:�jM<����N��ɪ-~ �%�ke	Y�z����ȭ��xu��c9��A��� 5��E�)[%I����=�y��Tܒ��M������'ض�#g>G.�N��_���mY* �h�G1t�6HXGte,L�6�zG�ȓI��{uɪ���g2�E��A�E�$�o�sM�����*e�QD��]���8Mfk�G" wZ�nY�l�q�2

�}*���Y�����E�gR��2]aJ� U��p�@t�KN�ջ�C�
f��T�6�0�:0h��op���SB*v�\�8��xң��:�V҆�:lk�쓓��mk���o��p�)��5ط�"���s�Y1�`#4�ӹ����`ly�_�Z�1�ȍ�;ht����N z��i��ֱ��֏4��`�%H6�
�p�Hμ�u��Y �#�����(	����c�`S G��O�=�(Q��q���(Ǝ��`Eί�� ��5��0+S�n�^	L��/Ӛ?������#ū���p�MS�o���w	����R��P����H�#:2��}��#�X��2�H��@$g5��[�U�����|Ł��
�L���zs���X�qe�ϼn9އ�h�u_��FNL
�d*g�m+<��th����q_��\�-F�+��p�7�D�P�C�>��UI�J���\Y�GBw�^#����|4��o��w���H�DZ���0Gt�3Z���/�" zj�	�~줄h
(�me�l9��L�#3P��d6��$}����UP5��N���e��V��j��\�����qM�C����Oыy`BR��$��ꀭ�kb��=?���Ό\й]�O�f��R���szY�z�+�=�_!�{�ogb�8�n����񟿬q6�5���d<|�H�ʙ�z��F����c�'r@gT�����y?!|��*aB��7�X�x�޲v�<>��a[	���'��)P��6�g�
�-��Y�� u�m~�y��~���	��h"�����h?g�á�H��r�N&�u���4�8/:Q�������|�c1gJ���&��A9�R�}��Qօ��5��Բ�����z'��Ʌ�c�����3M\�lg%�0��p�T=r��Y=��V�Zm;����9�M��Lݭ�ڨ�H�Aւ�&ٚ���e����!F���lh���L�-�����ti:;d��z��2���&$d3�)+�]u�=���HȗAGKtP�c�]5���T�`b��w���Iߦʰ
{68��Qb0"'z`P�M�{����`�w���Y���<<��]3�/�R�3��ס�5��h@K��cx���}y�k��}F��ke��TV(��[ҩ���@��	�G�Ӿ�����08 �o��h�K�b�q��""��4Xx�����T�d�� �w�,k2`�p��lFH����s.m݅E��H����$�G=�1��x~!������'L��M�E��!̔�2�so�  ����Q)���E�Ulu��<�-�E��0��8�|��w�B�g]�z��|�|5�B?���u�O�t*^p%�Y������*�;6F�~yĘ ��_nmf(����R�,|:�]D��`ȧ���%�?z��/����/����ݷSAK|}4���_
,@�W�o��y���Z�L�\9(D�$D�^{q�~_�^ٻ����@�e>)��l���&-�![g�?�^�|��E���XԀ}��֥AD�(�� ���DI$b4	A^���*@P�����P*�.�O���T�{]	�����"�����z?c��bG���׼WeҸ�(�d��bP&A2}W����Ua}?Ũ���/�'����Ә38��Ѕ�.��W�Np�Lv�o:G����)��wKm������oBӪ�o��خ�$=�'�c�?W��{�kH	'��[����
%��X��x�ͷo0
�w ��ttl�~㓊��\-�8	͟���a��,�ې�iOuu�ןx��}Re{m�"���^2;����tc{|�E��K_�� bϋcM�}F��e��k�oZz
WBs��J�"Kz����g�<���L��Y�Z��4^�D�%�f� ?��:�ܚ�\7�D%I�EgjrNk��x�}�!/����S���3���~Tn�('&���q�6�y娹��Q+�
ҫP��~c'F��v�$`�����x+N���y|#���Y{�Ň�G�i�h'�t�y����J����2|�/���#5&��,����?,]@���X����0��_o���F�~���U��_Z���MeU���'��B���5�_��09w� t �F�ا�mg�Iмu�e�V��0խ%�k��ֳ�f����5��)b�m"��n�u����a�C�K�Ado��S���,�=F�۟+�L?~6,��`9�B�*�+�'�;��Y����;����d#��v�Q��|�[w�k�}�x��l@�x%��0����	(�Wt��\ǔ*�{Fˮ���ѻ�ʞ,ͩ������{i�ASE��~�����p����CI���ছ��Ť(@A�Y�}(��n���z���~�5o���<���B�Y,ZYZ��Pd�e�����8����r��?OaG��ȹ4	�Ml��v2�S��^�Y+��Wu�� ���E���}<7���+���{a9_�{��xҰ����K��c���~Ȍ�C�mH���,�������]wV�A_h�:e7��y�P�=K(�1�ئ�0\���v�j�aH)������z���48KƁ�b0�X��p,�<�P�|0XH���P��gL�7��}Ί�������2��Ȫ�:���"Fw A�",
g���!C��6�.7^B�a�.j=$�����Ͽ�,�4o���%��C��pp���0\�=j;OIKz�џ�aO���$*�&��/������ʿ��Vǆ��/Ӛ�*��vp2���R�0vj_�Y
l[���5rc����d{O;��|�s��V����?�l\��BП����u�+�4
W�d2�ٞ	���6�U��ݎg��'W�L��.;�.��qM��h/��,�{a��)�Ǧ&� ͔�@�-��c�<����E���4f�*F<w/�=2K:]�s�9��d{�c^�7�2`��� �G{��J|���h��Lψ�8p̊m��d�%�����W�zZruTͱ���~�?˾?�׎M ��7u(�fg�ݏC�#������J�i�~kv�G�TBy��[���Q��uC�w��Sߠ9d�nU]��PJsBa�U.�
�w�$2պ�fT���o_Y�Ó�0N��S�0�!�>�!���Oy'$��l�$�M�b�2q�I���]=�?���/U��)9��Tl���Q��%��y	r��I��yiw�8}�Ǚ����&'ɘ��I��;x0�,�,4�\v��rƻHWa��/�/:��_�[��y[}W�\LB�) �a�)�/�'Di�e��~���޹�_ٷ���E���ۺh9Y�E2�i�m0n�BN�R���~5��b@2��}����2��aTx�Lﺤ�Y���l�/c���8�`�R���JV��ޣV����Gګd��e�\���1w��d�װg����a#���ĈڑM�[Q��?��a+��}���5�ΒW7o*�/uO�N�X����[#�=��_��kom��� 7���L7H��RE�5/NV}X�o����i���I�����a՜O�s��A�G��v��[�5�ޙ���h���V�c!�{�Ra m�'��H�5|����m��U��9��t<��r���*O��?�$�� �.�֖.�_��˽ S͎f�D��B&����O�	��P;�)�Y
�@�F��K�$<�F��c�*XhT��:KTʹ��	 �?i�{�$����B������E�!/�-N���]
_���g̐��M���J��te�彳�W��`�ԥ�����;Ac��c�A&+y	m��x@�ɟ�WL�l>����WW�����ԮC���gZ2;�tp#}%�h�D�kc~�2/7����W"��侹#ߦ!�3h��a��P�4Xͻ_A�1K^}\&�*�w�O4x�F��paੂ��)��ğ6��P�U�K���{U7.c2@?���M�>VG�� C�%Ҋ�݁�Od�̢���K����Id���eg �N�`-�Ƞ����/?���Dm��r���:6���N�˥Q��2��Y7gLYd�?B=S��U0T��y�)l|T5JÝW�Z��}/��0T��&�x:B,�q�\W11�`�IY��Q�|�/�h;[� >0�ܝH��]��KT�wTC�B� i�I&xݽ=�B�J�f�����g�>2��0�V*p_*g-���oئ$Mw��ۯ�dY�=YFG�~Y����ɪ��q�J������fy*1�t���W�����}�`�_�+f4qf ����d�J�ct�#@�B���ѦfC��l*�����.�r�-X��AP�\$gڏ��Byj�O��{�MTS��\���	��x����p��(
��Z옒�+�ӕ��Hn�XM� 1��f���k�TFY�D=�	O���&'!��`3��.$�bP/m/S�C`�W�r��$[=U^��-k�]E�f������"uq�#%��B~�p�qk��t���Ը���&.�����-S׎�h]�;}�e�ۘ���)�8�z̐4�Ӻc��l��°��G?oͅA����M;u�\�2Lĩ�F��8@+u)��s�	�V�o��Z�&A�����y�ʮ���R4�5���"pIY�t��%q�Ebɫ􈚉�k�����I���r*��K��@����KF����O����P��2��,���^�������ou�6[�%o�f�+���-�W�BkA��l�B��e�:�{�y��gLC�t�G[�P�j?+ �Q������á�nt�i��i:ۤ{z ��A�$�p�Kr�p���
��d�A�X9��+0��gG�=�[�K������H�j�׋���=O٥q��DD��ja�S�p�A�
��̋t��i&���Ȑ�N�r�A��vy'�n��������!���_LE�w	d�㓛���u���a�5��8s
*�I�Ǌ�A�M�N���
~1:ZZ�'/e��w8�i]��q�����j��1���TE��(P���JU��c�~��N����_�$�0�=Q�*��*eҿ��~�-�C\��(`��n�C	�W���8FE �$�N�w5�*�C�$
Q'��`�!�uH\Y�oݢ�E�G ޣ�йH�p��7+Qb���a�RQQo{џ���v��`��������ۺ-6��jc�� �L0�C(ଵ�1i(���"�]k��^�%e޷��%~��A�߭�h32W�d)��D x����u�[d	Ý�)<����+i�����I���Ø���� �F��t� �JQ�Ӻ7���v�C��X�K�������v�Tٴr��Ϻl�y!��?�l��>C�z��B��.c�Dq�,6�� �w|�s�����L�_�u�� ��t|F�����K��|C��\�����X��L�p7��Q֨����D���+Ĝ=|�����|B��16���b�Ĵ�K3�c�a�^`�zN/C�{��/��&�X�"1� 33�A �Փ��� u��F}w�������o8��?�Բf�z�%�� o�����5��kE��&���YD�`��ĳom�f��E��*)�I@�����nVBGA�1�\�2Fuho�����
3���r��coinP�8�!(�v�����@pD�>��8>�O�D��@_ZX�b�ኲ���=�j<xf���a�U�ɴUa��0�Jj=��e'��D��p��c����4"a��Y�,+�{e�?F��b�	I��l����k����͕D3|sy&�k���ZO�]z������Þc��?X7��m�X�!��:|�>�����b���
Z���[f�G_�OM3;���)Jx�y��뀍P��O���6�M��q��b�@��t- ߍ�-���nv�E?i��x�U7�Fͯ���%(J*�g����t����"q6~����?�ő���"r��_�l�~y�u�y�{�nhb$�]�h�5g박	#z�V�p��:À�k�R!�����c����ߋ��]&�^�nR�'��$���� �>���a\��vh��oH�>�X�����#q�B���]����a�e����-Y:�� MJ>�(1J7���k�z�Q%�Txeq��X5ƨ<-@Tɩap�0�C�C �g|��DΙ[��0Wh�ߦ;T|��s�n���|�������P����;#n.q����[��U�㒛�»�c'	qeE}���@ͅ��#�,��V�c�b�u�J#�3��2� �u���+巟�D�,0�a��P{�虁���R�/�a�&[l���8�|-�{�0���z�3C�c�Zh�l��!�}���vB`�J[y�u�5�t�A.U��՚��p��W���8X'���*������j�F���� �N��H�~�=U���A�S%�ORʯ7���,yR�G�-Aq����#�.8XL�cV�����,e>�7���n>�3e�8�9ٱ�Gɓ�i���	Ӧ	f7��b�
;��m����Rٖ��2�i�y|���3�\�z
Dh�*�4]��3W�/�e���nW��$
Q�9�<�].-	i�`�X߬��*���;�B1I�T)�!��6{�q�-�czw��.{$B�8�(@	=�r�����m�> ڕPh����B|(�2�@��07L��5k{n&�hTƕ�5��D����gZ#���-)xօ
��K�,�J5�R�Y5������~�)kV�{���F��3^��|�O{�%>�~1��bV�h1����	*��[������U������gͅ��#D*bb�@Uw��߼��ͺ��ϊ����d�[F��YVt����J.��&�����,*��F�b{/l�l�ʂ�[_��;�k�s��x����JG��,�P�c�F�r!KY���۱��X��+%D7񑫩&=��؂���n$�+�&V�!$��5�1]���J�g�?���`4���~x�,a�����o���N���ti�5�x��?}d�%v�P�V�BED2� W/%��b	��7eF�v� ��Մ\X�|�]K6�}i���Y3 �����yD*�S-���1n����<U2^�E���ɛ��E��Fb�(���<���Pq������Y׶�$8N##����z.G.Ii�N�g�U#�Q,�V�����E���pa*���&��D�T��p^�[��LT�L�Qps�������ɧ���<�b�=J9�q3�m���ȏM����+dk��z�a`Q�Z^��D�x>J�O�#�%�,�|qp`d�T�o�P���!�ڴF^*����l���,�9�����C%�l�j����+���In��eOq?��^�kY�/M��
�j���9������~,E��E�u�X�1��"�G�i���R�4�RǆC�m2���<�U%I�:�X�9���$��ɵ0��9aZw��msx�剩�f�4���_��>?��S�+kŔ���4�5��n>	RJ��vAv�]��f��٣Տ�,�M4��y��1�͟+��#P �zҩt�X0G�6N��.IR�j[���iu��|���'N�"�ѣ�������	���<@~x�[�������Ƚ����~F�v)������� 8m�B�
LK��}X/�2Q_�%��l�KRM�(E>T�r�(�2P�~;k���?�@��%�^��\uV<,�]��e��T��W����T�P}�C�ڌSKR'\2�CX?�3R��Ě�jWF>����x$Maef
Kt԰�*�?"��;�$�ķ�������<�V Ro�o tl��,]�i�v}�K֔�`>�P�����X�Ofu��3e���Pt5F�� #���9V�����ܳ��t|�����m9\�ɵkL��R����~�tK��S]�}�}��D�|�G��@c��H���[3��Ɲ2{�Z��7��]a�C�$.����W�����nԑR����^��fpML?xE�7=��SL��G!�B	��J`�a�!e�2~X�r�=���re�쇩5���BnL�RI�0o��=��D��j���Kj�Q0*l�I��у�7�i�p���$G,�YEоXh5���;�-�o�ng"-�ĥő�'�z�Q�'�a+g�q|V���D�q�&���.���0�r�D��[k v�9B�
�.G�u@�V��ߋ��j�0i@]w�ߩG��-oF�:i��L��ߐK!#����[��u�XF����P5��~����	��a+�<AF�f��CP=��+DZ�&����Щ8�t��V����.��� �C��uc����f���Uq T�JhQ#��X� ,��:���C��<�
eк�_��e}���v�:bkl�����Fc9����ec����d
ը�*k$Bד�+�ID�i*~�����/��#��&~��T��g���A�M�0��`_ۺM<�y'r�B��T.0�
��h�^`K�e�Џ�~+0p�����3}k� �j�����"��rP׈�K�h�y����M���J�;�ԥƚ4x���b��c*�:,�n�r|pKX߇}(�.2�f���Z1�C��P@�Ot!8���<ڂ��\����b�b��j]߻A(�|�-n��m�F�MXs7��z/���<9���Ӷk��"K���f�D�|����[��U�����ιDw0��j�3�kcm������-��A�Ҿ��2'\-���O
� ��o���eJ��H�V뵻�q-�<C���p��l [��o����Ub �)h!�ҥ5K�-��e�ؒ8�y14��o����<�^#���j��N���O��戎�=�a褀�Θ3����N��Ѣn#���:��fr�L�ӓ�k�Ȝ�NȬgnHM
%M�,D2���Y�WwfP=��W}~�^"2i;��V�a�(��ő�
A�?���� ��1G���?����I���'#�d��#�5�Om����jd��wusta��x���U�Ő.�l�l��1a<�a��)����&(4Yɧ�9:=I�<�F��=�
��}�Κ����l=I�m$O�.v���C�����V�ŕ�(£ݿ'��J�2�����޽��z�V:gj���:+�.U2[��@��`$w8�e�kpy#O���3P��MC|�'��&�&���.3va:�e:�z�#�\́Td�0�Y0�UEڟ�.��MB�Ed���  �p�j��m����h?Y[�� ���AmTh"I��d�.���N� j��[b�n��,���m�i�dz�����4��B)�Z�f�e�� &l�NL!�	Z�G���v���m
����4��_���$I��]�)�^�]>i���>J[�sv��4�fF�)�E �,��tO��By�|	>zجɁ,�>��lp]Y�0'y�� :�7���DD�僪�k�o]��8Ω���Q��N��a#�~Ů���9�VF��LC��YF� �~����-EH�2��$����Ei4~ƐM`�ٰYYe*�CG�m8>an.�S4�S����&��;�xj��������W!���^o�-�6l�s���Q�"�|0k}�wQP�DÔ�������ٙvE�|)�'�wܝB'�?#:<	��Џ�1Ǐ�%��ϴ_kRBB�;5R�3���#۴����]t8��|��7��Z�{��/x���6���$�Qڛx�ӛ�l�g11��j�ZYZ׊u��H������҉(ݽ�r?A)�}=��+R @6\(1c��X�e?fA�e����v�IsT�?w;�$��3��|���e��';H^������W�������nb�G��P�WM��jgϘi���n|�͂�F����@��Shǩ��h�ky��_$�v�C�G�w!??k�m6��D��Zе�d�6K��H�1��Z�|�FK%v�$T�C��tp���$[�|�դ�qi%X�63DkQ�",g��O�^�K��X�k�i�S�c%�o>�����Zh%�z� �H
13��_�-RVOTH������ �ܱ&E��Z&C�s ��KD�@YS�������a�"���K�W8�S%��]��36�W�=����I_����:@lx��<�y�rJX�{���x,�q���7�����i?E֌��9[�-K��Ǔ��!fZ﬙�TL��}�3����#���*3���xI$Ӆ�(�g������uo���ôP��P/���e%S5�:-�!檂Wb�/a���\2B?koŃ��+kZG]!�γ�tv,!��DI��F��Hk!s�&,�9��nSl��|�,�>�'���|�=�W�ŦI^d䞎+���S�"��KGX1�(ą4C�'�g������<`�ޚ)�#��s�U$SxqL� ��=�ܥ{�(�U��-��r��rs�����H��.Hz0?pр	 EE$ǽ��F�KCZ��fX��[sݟ��_'�28��@��+�"xD�k�`�Y�nB�%��h]�!�W(�#��5�3�)�ƭ>�-_~�;`���G��4��g�W@Y��Y:��&���i&����7�A`���Pq��-�y����  D�)�N�Oa/!#M��`S��	��9�@�
�~����y�ٮˍe^��k��4�+e`�Ia��l��ʳ<��pA=;µ-���w����zЪF�~�4���(&��^�J8.Or�(s4YR���'~��6#���hjKNÃ�ټ2���1nq #�;[\���R��vr�\Yt���o3p���W��!��Da�x�R=埇�m	���:Gj�����f�`t��&��Z��Yejz�9ʦ5�D� ��7�x9��W����k�{�ξ��F��s����c3�u+���Zf� �F�K�'_�B���
�.
��S4�Y��S���pH�Jhq�4k�R�NQ�����P���77)h3�"�y�
{�q���ȇbD�n�H_��������O V��ǿ���6���B�Y����r��Ia�}!��N�xq#ǄL���Jii�ߥ�G�]X�4ۀ��`��}=3bϣ��V��:[́�]����O�:�z@����Ε #E<���;�@�<t0
F>a�@h/q�)�����k��݁����Xϰ�a�i5�ŤX��8�m�C�k�TNv�U�8�ϐ�XQ*#�#���Bt[a����U�ѐj� o�d<f����M[�����[��>g�q�q���s7�Q������H	���cz�T��9�
謭�@I��]?�n��,]���7h������I4?�d}�V㺗��g뢔�n�l%pH��*NAw>Ysn�l)�E�O9��w�
_B�I���>���k��5���^��5�9��aX�2�c��y�A��G�~н�v�F��;`)^�Y���9�ڧ����)G٧�KB,�gWƤ��U`팀h�U�M�Ѫ��1v�D�l( φ�W��?���%#���.�s6C\�J�/���
i C6e$��!>�1	����M��
['%�������PvT �@����*�&���K*R��n8�����Xж�Z{C��\�%|�9�Ԣ�����`�_�J���V�^A��~�9�f٨y�#����~7�cWC\$�X�'<���N���뛗=UWS�t	j��oOa����u�1n��� �a(�&��%)Q\���Xc�QOs�(Un�M�ey�I]��"�T;�&a0��>���`>&|�K6�t@q��`I>3;c.߽�]i���n�|TA���C	�uU�A�t��T���+�_n矑��i�<���	������2����Ԋ�|���E]���Dy�X����������BCBQi�e�E�"�::�I����Hp �oGc�+������h��S>5�t�XH�(�]�L���p|�"��Hor�y/Y,��4�&`E�[�h@��p�i�N'$�?�D ��H�;�B 2�7���Ԇ�^_7���o���J�T='f�i�8Qj?'���ԺH�̿�|;3��/&|�Q�İd�c��^n-W;�*",�v��@���xޔ�Rp�M�y�qe�����%h��NS,T�A��&��˄�A��f�ˍ�"���i|7��K���Gͱe�B�Tk�,�����z����ݟ̼�?1�DO����$Ao��'��9�{��܊1X,����u��@�r�۔�Z�;8e [�n���I�±���a���sɅaoS�^N6�';�M�8nd���Uu�_HT��)`�bk��>��&^`��v�S>�F�`����Qº��ȷ��G��`�ճe�wu����]J��?ݳ�ɏ皪�^��t;�5]�>`��vn��Ǭ� ���QǕ�{�؅�<V��p<@Zaϝ�$�6��wE��wX1R��h�b�}��<4�:��R1B���B�ȱ񨑄2���:�y��U�G�7�>o�#c��6s�ZS��n���X�IB���6��w�G��EЋ����RҸe���ǡ���@O��Y,����G?ݣ��/_a ��$��#��8!��3��F�q%��X<V����)������,'��f���Ф�!�/���@����@�^6@��G_��hf����i�_z$�ֱk݁�J��,.��p?a����<�E��`6�:���^O&�c�s���YD�����Ъčׅ�[Y6��m�y͕N���5��ttKۉP3�����ް�{����˪e�	}���Ӊ`)cB��)?bc��Q�,z�!�0쵎�E�܂o�m��EЉ��7����f��5V�x������s�֑Y���μ��!}zS
k:�uiq�QaQ�d��ץ�V=�[E?�~!��8�4����k�E�d��s�К� ���ADF�~o����ӄfDu�Ӝf=b
}T�\���c�׳y�>B9�J���s�b<������M�鞿��-�'�oK���nE1&CQ(yݼt��<&���T'6�t.c������D{�>w����=)������֫p�x��?)��S��Z�)2.<��`�/�U3�ZP�ڦ��k��CG�� ����VU�D�w�'?�T����1eX�ҋLV��o����������6ͯv�_��������Q�������(���e�Odn��_ʓX�Y����u׻[�¾��� ڝA�o����$!z���{>Y@��Rgm��=������R�<�w��$a�FE��O�N66�u1u�*�k�.���$��ZGY���&ꮈPP�~ʹp��)!���.�����|p�\"��Y4��9��j&�^c�|w��4ˏĜ��6���='���w6Y� C�R��K/��7�aem!�`���`�i�����+������q
����1i�*޼�v�K*��_���Ra�ٓ8���_,G����g�}�W�atqO$ޯq$�m[(ꅏġ���(���:�/�w��_����>X��U"�Ό���g횾ƅ�vQC�h����EeQ�c�ƼJI�'��E�k�;�R�V���F�0Tӝst��8-��4b.a
����~>�� ��3fe7��VOF90	�)h����AX��B������	!�܄M�����vpo����gk.l�`s�+�6o��5x�a�FE,����n�w�{M�;�u
ǔL�¨�V@�}��w�~������4�Tv�ɹm�N��ŵ���T��}F6r�C�5�E�2J�I�����w��|K��u�mU~1E/������E��d�z̽��	����߻��01Bx���C�]iH1���&�	���;r�\4f�1~�џd�?K�-h1/���
*�����"��.
����Ρh,����0��2�D��֡�w�7�&k��������?�h�p���3�$E���4���'L}�s�1箕1���+�[#)78${����֫0��K��[
�I���-��8�Ol����ح��#��Hq\���M�j���S��Y&���~$<�J�Νr�sK��[?�v�����t@[� ܈Pq]����U��m����ecIV��t�_e�Bi���ŭ�z����P��b_d���|�<v  G���,q+�轾^Eo��yR���S�b�!\Q���%ɫ�u���@�;��������݄�z����4��0S򢱻{�_��?%:g�-ٺ8*RQ66h����S\B�RT�ϪPw�y��w���J���0�bO��0M��_'�� ��C������ L����̖�%��sYZv�(f�ܲ���YKȠ������.�W6M&���ѫ�w��x*�;s9LN�U�t7���x��'v�f[
THh�Y􉮻G�u!��	�Y�"�
,��2��d(h��y���n @:���l�]�zFYa�8O�"�^ �,�[�?X��o��S��C>КE�k�M�Mtп�PeƝL�4V�A��Ɗ~B�r2���r�+*qo�_`,-o��"t��RK]z�g�փ��!���)W��ܾf�L��j��#���Y��>`��>���@�<1թ�󄙿�u���T�0i��E*�'SH��'0wӧ���]lI���
����}�j ��.H����QX����73�w�$�^ԅD�im+��_��]�]޵��uq�W��DV�6R~Ub'z��q���ae����զ���CƢu$J�6�$���*�J��`�}��$��"��X��4ċ/J��Og�>rIz���S��v�,Д@U�p�,�����=�8��hڄ�����VV���qq7J��HZ�����.dkA ��Mо&�����i`�ǐv�dlm���!S͋¸��>F~Q����0\v��$�о�B�b
�X���w�B�Gjt %���-Xb��#��c�訮Fn,e��;H�	�y!晣�cPhq��������P+��$�5���B�ʐ?���^�{I����pT�����y�X"������TI�̘�F��9pLV4ĂREw�~�qs3��`+u]�T����J�:zC"IO����A�9R�����΍Q���]~W)g�۹��a�Jr	������r\������������SB�<��A��Ne�Rg�� �����|N��Ӈ��w3~������e#��
����rS�b�z��>mt!&�;m�H�)^L'l{��CO�����߆lEHնE@es+�ݐ��yg1���C�����9��AUV���|E�h6�Ĕ#T�hY[�K��̐��ȕ��\�(a��O�����I��J(1��d6�-N��Ԉm�^/za��W��=���
kMV�\�\����=d���h�X��
��;ݓ��D�����P]���T�anX��u[�[��m��>��?=�s2�T3���j�jPh����qA�����.T�*���B����`'�I���F�S��<6��L��@[�v��y2)z<ǿ�Xh_��T6ҏ�j"��iL*���@É@f}"�UJ ~~�;��B��X�	5]�����6�[T�ł��7���oA���fq��(wօ*�:l�T>�c����7:£��2[>
c3���0	��I'wrhc�M}_�ڥ�����])|~���*�%����(���U+���Xmja*
��,'���ͱ���~�}F�\"�������0��H3`���{1�I����C}$O��X&�� �mc:��m�����ח����}���4N��M�R��$˄�Ul'~���↦=u칺p�������>DpyI^����v��즻v��P��C���_t��Js.������@�����X���]���:�q0	[B���#�Y;JQ���" �H��[1��KQ�	�gE~(�=wZb̯��Z4~[rb�T|(���r,F��X_�5�y{��f�V��i@�%^�wL(�s,4q�]I��g�ϵF��I$h�ot��G�(�T2�I�drQh��	��r�ÊP�a�=�Ϛ>�cd�:\�D�A�cĴ|�m ���36�����0 ����-P��Йa�� u����.�w�d,�B���D�Z27��?�.�m��y�n'a/Z��O��"���������݆w��9��{�K`j�������#瞊��;�dY{>�����9ئHahT�(���ȁUJ���>��W5��!������?�1f|��.hN,���Z���X$wǟ7��]
�'��X���t	�X�s���¨$"O)+�B���d�s�Q䀎N �C���*5]�c�ǖw� b��=�V� ^3c76�$����1��Ս�uT�tqg����Pbw�@d�u�5��A�/��cO�I�H���'��\��!.���0�V7	õN�~�;A�$ˉ��)�2�9�c�_��>������>�쐕`{M���[(���SL�p�./Q�qK��׻��� O;���\�W�/�A��0�	�Â"ϙbd9`��H{&W�jD1ԬI�is/�,VH����L�{�4�=�%���lVbO��{�ݪ�ֽmS�t���ܨ����U�g&��"��!Ց�3�⦓N*V�8�@����?��:���#͡���	Ȣ$tܹ��*��'�
�Dak��i�uι{.s�,��r�2��d	1���2MSx]��q���'�����ۗ��3ȭ2� B����SÊ5/���c;�י���E��u���jAJj0���d�`��r�?����7M/�#�V���s�T��<��#�\٘.�A���)\<�ȴ�`�^��c���x��U�</��A�?59 ����g�4�!f<9_�7�=�ζփ,�|Ez-��T�	}"��I��@��wj�`���J�i�y.Gu��crI'�i�����r�;�L����˄R�O!/��pTW��	����ڧv�}����M�e;?���FQ�Ә3��qep�1�������ꦠ;�C�W|�멞*.�fހ��^m�b�EW�9��D���N�5�S¿F�8�+�*8 4�����)ğ�u9�f+|y�ػ��b�������*.�t��\�m]3E�\N��BA\�F�~���TrQ!�M��I7Q5�{�>�l]�����k��̀Ӟ�q��c�^3�3�P|0���h?�Qi�x�s/}�۞�T�'wh�!L�C,#���h���5�,b�3�K�f�ZPq���]��X�߱�������8'��z,)C=yoԂ�|��^E�{^B��^���s2'	>���v饴V�D0����WU���c(v�.�dw�~��O4Z��i�Y���� �0Ц-]�1�>;5Q�9�'!��ҥ,��KIH�+.��-��ԽÎk
U�=�� ��	|�G�I@��+O��,��j�+���\�am^`��Iul��_P���4yrX��=Hp�����;�s���6J�b%�\��T�9�b��"닸&��-��)���w�Gşr;�4JU�����"���JXK�D׆�,!q(Qyw^����W���8<»E@�J�Z�8?�9�O!64^3.�HRT8��qսk�~�	�
Bb���#
g�i^-5�_/��6sgM�[F�X�t�)��#�b0o�=l���靶j������s�x�f��7\͑8��=;�fyj�O� �H�l�Nq@$S�h�?��Q�C��H���@�@�m=)��n�}i��
T:�E�H���&{��5�r���I@V��d�œ�"*,(7Aq+�_�j�s$^�T3Y(��٠U��+:��qÖ)1��_DV�7���$�Z�/ﲿ�Y"�a�˳�B|�O��/=M������c�����$��v�l\TCu��gA�p��Ы�+�(2n�ό ��78��ҥ9#��B�qE��;̄�ҍ<�*���@wS���~�_������Y�B6���y���3���+p��l���gxdl�:X�@Ea_q�g��%I���:J>R$y`�G�=��rs+ue�y_U�@4=8~O�8�x�sM4���yb(���Û�ƐFYߵz�D���9Ɔ��DKm�U�f�Ւ�%�<�ϒdi6��w m�c��ܺ��y	g�� -$Pj=u���`���tˣ�t�k�7�����S�����bţ�˻���y���<�'��U�G�%��U���
���	��`Ih�{��s���Tv� %~��A
���ģ-�?f���w�͜�SG�jC �����v�n� �o��RL���^�}��@�}3���
���ܲ||-�g���x�c�c�Զަ;:�Y:�z�u p!����(�D�������5R޻ǘ9K�@�����i�Ү�L�f�r�S�{�wv�dU���Ș�>R҄��ҁr�B���@�F�Mh�`�Ys$/3���wh5�
���f�m��gʁ�i_�-A�O��﷉u�N��ǡx��U@/bս�e�������Z.R�E�����eY����S�@�L�� �f3���9���\zЊ$��E���Kb��7Ut��KKڅ�dV?4P ����5>;�XU��UNR6%RR���N����fBQj/j��e������>���h��Q���1��.���7���(E%e+?5��g|�.;�G�B6�U=�c�\0��2xwT�>�`Aگ����ش���&�h tM��ͻ�{wYf���:$�
�z�U�))i�yR�9�z��T��T�Z��__ڥ�A_I�