XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��QU1�t,v��J����l갺 ��̧�O��h���c�N
�]�3m�T��dh0fz�%�B�4zM�^�?���^V���b;7i�ϡ�`��[���T^�8��J��޷Ȑz �q##��Va�Զ�A±�g�(O�*_����R�~�����pZ���uQMn�,�e*G�q%���Ikd������Rk�؂/כ�oj}�ĩP_����>+	ބ��,C���1�t�dI=�r���F-K��zZ��7GbD����W�R��UP�-_q��L���W�{�$[�K3����3n�}mj�ߵv:dc�H"'e���E��[��\�$.Y/�,��+k���O��2�^�������ʥ$�(�<)��c/�c�<���q��u�豐�l%��vV���3ι�����q���������c�&�D����vw>��8<ҧ�t�AN���BD\у2�`�g ����zu���r�P	�C�'�/2��p@�=Z��Ա1��emϜ:/|�u*�����,u�����QLE�[2�~��]4uT����IL܈����;}C�~91�>�֡P�r����}*��S#��B�1k(�=0~�PaRxW���l5��W�b��~���.͟�<\�ɛΌ�z��?�I�ư��#$ק<��-����<N��p$&`����d��?#պ�q,^�J]�	��8*�ղ��ڪrWX�������
�e?h�2�I��Y���E�{=c��
�5U�`�!���QG�	��Y"��GuXlxVHYEB     400     1b0�_i4Zm>t�6�Q�w�٘�U��� �`	�K���q[���~��6(���?t�r�9�Elq͕l�3Ԃ�M�����x����}f}<��]�q-ARc  *3�B�-�	��ހ?���%��ϊ��D}Z�5�Ql��6��*{�i3�)Չ�/ޓ��N�fY.��Cfg_@C�_'�����06���i��R����.�.��ۯ�XL�g��iW
�t'W�[]���r3�ȹ/է�LT� 2��f�B:u�u=7��漺�ZQ�G�����:&g��{ߺ�B3l ��Bx�!���`�r� 3��Ce����\��)|��ѧv���&����w \�ns��q�Ccԍ,��0�`z«�}�o{D����Ѐ�#H��9M�n|���-]si����R[�ğ�����bu*|�Z��G*7N�M�:�XlxVHYEB     400      c0^qR�I��h1�?��Y��B�>����T's�f
8��Q6�o���9�����j�Ȅ	��|��wJ��S���_�\ئv/wޚ�ү*H����b'h���I�ζ��I��|�T��xh�,G�:7>&5O�o4<���]��cv`�Y=���v],�.Y�|�P�sXd����+w��j���f�(�XlxVHYEB     400      b0��t�ʲ���Y6k�RuuNO!t�ش���A�mZ :��Ue��
h���5��>Y�̸��2�;"|Q�Nv�|e@�!:��^�т���\�׵�V��['��]1�4��@We�$+0HN�⅙�8��	6�0�e���|[�\Q���B�Y��[��������pߢAXlxVHYEB     400     130c'm�Ǡ
_r4��u�2�f��T�;�wN�h��E���~��-$"~�ԛ93<��Ug"h��m�a���4����iQ��n>$Dx
�$Cڹ�z%���[�b��p`M�`ȅ��H�؅d�v�*�m�i$gE
�����o��w��}/��3����+�J	�RDͥ]$ت}��Sr�icP��[�6g�������&�:#!�;�y�E�iQ�}8đ赨|Eň��0���r��K�N�[�^���M[��:����@_Q�c�B�T��v��V�S��\�h��c����s��y�l��^D��1){�XlxVHYEB     400     1a0p�y�m[�	��[��(�i�[1#菨��?��.��O��fD�V�u�𭎭H�Z�8]7����F���T�S���x@�q�e�����#?���jD��#|t�7(��&�(_O5�L�:�����s�Leh���ߗ���YE�ij�Q��ư��A �p�Nb�~sɝ���@�J��fd�������0�L��˧Y����H��  ��2�~S�=~3kq����8�۩�#�_����B��k<���c��k��nl}��T0��K������t�,�1Cg&L���p"᝟�'��>�LM3�al�=V��#^��ʴ�#c�N���:'��p�Z+AX�w�	0��|� rHtH��lP
Pr�&�ԕ慩�"R|�kl1��G��@g�:�+i�,N��������r�G��ݡ8�ȥ��XlxVHYEB     400     140H�#��N�|.�n@�r�\0C��9��?#H�Qw�Hhn�l�u��n�i�ۊ�l���O�����Rl�`�����	2|������x���L����vy��!��ެ&Uw� ��nH�2�sŒ?H�_��Ek�,P�ҐOİ����ɾ�|�� _�Utg���Z��y��^0� F$���l���p4f0y�b�2qh��IIy����]
��ż�g�>ڈ
��P�ȅw0��:HL�$N2s:�c}�,G-�n_�}���Z�J*�l�| �3�\��5m�|V����P�ϑ�Lp3��R&���2WXlxVHYEB     400     120�,@X�k��O��@ݏ	�VR���}ef{��)P:ߣ�Z��.�7��	:�|��:��F�^�L�k��J�A��w�O���׏� =Zs"z�\��ƈ��)Q��zq�]{%z�ؑ�X#<��z?���ۥ
8�e����SF�[�Y�y��Ɂ��tt��Oj����|J�:(΃��&�"����O�!��^�b�1iZ��aԯ��qo���C?���5(�P��ɍע��!M��
�������mZ(����?D������ �q�}��W81�Xܿ!o=
�s3	o�XlxVHYEB     400     110����W�XAp������1�|A��^�j=	��LpS�:N*2`�ƼEpy�B�a�[��$�MG�k'���^��y|!��	�gpѬ����$��T�4_<Z,I������&j�g@�A�iM��p/ ����AU'8K�b������3�ɪ�<���c҂F�ࢁ��A���&���tTr4����q&� �݉���\�W��&ɜ-~��\#�	q�퀶0��	vF@�q0����>Y�=Z����[���'�I�Rw�X�7��!�c8�?XlxVHYEB     400     110a��� ��ԒȳSui�>����}��������]J�,�0��;�8�(��~�eMS
��m'��wp��˻�M3V�;��!ӟ���U<�+L��Ԗ!yr����ln� �½������5<b�1 a���
|?u�l7n7Q���!@�m@P��L^�ckW����S�#�GtS�%��5K?[ta���x��q��Q�mC١w-4�HUӵ�,���ͳf1�V�%F]��ղݽN%��J�*�^+@��ݢ�gҠ�k~aBWt�K��B�	�XlxVHYEB     400     130#�ŚZ�mIu�Y%��5>˃�d,V׎�Vb� b�6��� �ô�@[�3eA���!"��6������	��,�1R��-��uq���;`�LR��6+��lI��}��Mk�ˬP_K�k��W�6	���ro\�Qk����c4�>��D���YT�.��}��_v��oz�0К��X�Gh�lƗ��Ô�=^0M�)T|�Ά�Q�fE��;9�ˋ0���˦����Z��
�kp�K�X�C����F�J�T%���܅T*�~����yj�tq�������x�Q�i�Rn߇ �J�b�7XlxVHYEB     400     110��C;H�"�X1�0S��`H&P��_�A<�$���ϳ'��0�F��p����Y9��#��l�aKή�.�XǱ�)0��ˑ����ptc<z��@}��R})�3c#<Ȁ�D\��
���Ĵ�O�����G��A�C�9![4H ��q�S�-�v<�b���3�F���`�i�ݴ�y}P��q�E�ډ�s�DK��P�*�<�1]�V�<�\�>3�E.d�t2�L���mX��gXm��C�bN^T(�_�1�vXlxVHYEB     400     120�W��查6m�.DK���y��mZ��i����"���I?Ɔ���WKN�[���a>�>���=��A�>��B��6�y��("���x.6��S��0�A��H�;��m�w��I�;=�������̣�;����EÆi�=��2�og܉�B&q���F?PX����u�[,a��S����cE���Zp��U�Gy'͡7��X��Tŧ>�p���Ȍlag�]�D܀��&�-`���=�M� V�߾�{�ݍ�5��5�{y�������*=�b$L���|XlxVHYEB     400     130�2�Ҿ��wM�O�ʟ>5j����Y�s��N2P)�m�w���U���;=V��q�q���>}o L�Ibe(:H�u���v9eh�t�:�I�E���vr�������JvN����/�h���cy���ʻ�h䑓����]O����A2b�h���D!��Ը�	��4�i@���h�%�\�:���^x!�P��8�Erb\p���Lo�'�?j���:�t�&�m�$BA��r��O�p���Hq�"^y�
p-�I��A
#S�����;�ltͩS8�^�j�t��XlxVHYEB     400     100���H�)�����'i.Y�U�8l)3���}P�S^��y�қ�p�1S$[!]�T &8.�h��>��=� c-�c�p���]Gʎ�{���k��HV
��e�;_���lRi;z��j�+�Ѭ� "��{]�k��(!	�0"���t�@�G3��yTe���r��s�Z*�po�G��׃*& �Xo�c�p�� P�客��m�U���������,%;��:R�&�:�,DZ�s޲�HB�>��WXlxVHYEB     400      e0�.~�t�<�Sz���������[B�=U4FE���f*\��gf��@w=�f��e��V��:*nX�B�q{Ԙ�ڇ�]�����i���z{��4��4y,��%����	Y��B��h� 52:A&Oև�|wB ��7%�dJ7������Ws$r+!�6xKAc��8�=�d�Gד��ZF<X���oY.\���ٵ�����jGXlxVHYEB     3fa     160�|1���!7�:J�\C/Ӭ<�+�#���8x�4 ��vU��=�є,�����Y������g���;�X��r��}.�k�v/���L9�՚�!Ƹ�@��F<:�����/%�ʢ��wXh�}��;��k�������ʜ�i1�>[F-l+�%����B�1�C@>$����'aI&a�t3<����?`♩9@�Z�0P~2Z\����'HQI%�\�-3���?�n��]�W��o,'31���4��|���k�B��ٲ�z�#қ0Z|������C	S`l��M� �q�f��qe�IU�_h�=6���1,v���C[��a6�2�Y���/