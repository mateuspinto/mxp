XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����>���rş�u��h7鴉�7'+!LE�̫t�EFl~��=Ů/��C㏳�a�Ѭ����N����hC��ft�.|⅚����*�6I�h���	T%�)-C�͒C�5�[b5�	���CٚCIjc������yQ��D��D��l�-�5S�r�h�Y�}�p'�os�����Ɲ2!��Ezis��[��g��e��w˰�~���RGd��������>d�Q��V�X�@ğ��q���g+\�)��^=A���A�&�΀�3b���Kx{����w�h0X{��vE="���ɦ�g-鳻��u�0=�(|��΋'��?���Zm���:-g�������<Ѡde�8 ����j�;��'L�ȴG��rH6��}��	��{g�p4)3|.���n5^u�� c��!�`"<_��V��6�J���6�����J4���L	k1M���i�b�:N����(rե�'�h�v34�p# �?J��Wt�)�����W����������Ǡ�J4�׉N�q�}/!��ST��4���FLa.z[SN/���t��g���e(�.�����D�����M)��� ���m���h�m�{�k���*ӳ6�/��
[�r��-Q+�f��V��ȟp�S�D7���/�&V��UF��}���Mt$HC��ƛE���.�}�+�P��R�§���R���3+�������/VS�+oڸn2c���:��4�f�@��n�Ʊ�)Nh�{�[@���XlxVHYEB     400     1f0�A.�H��PY��45���E�ҫ�������D9��a���pt+}���bj�:�6mCfH1�ŝ��IH~��V�ψ�*��c =���(͎4AYm�	y�*<���J��	���2�2!9���[�F�m 8@fР`����J�:r�h=E�TȆmQ1w�k��SF.[�%�C����������	����s�c�R� h��e����ɷ&Ș$��;�d��JP��	�x�!�%l�Z�[�%�._E�\~oM��`����o��b톣�'�4�3�8���~m��[#�d��?�����X�Mi+
�Z0�-`W7Li�4����E�).c�#ƙz�2�aJFũ�5�Jg��V����f�q�II]�0
;	�����ˮI�++
�q�ƀ�t)�0�}@�掦��y,Axu1q�����8tɗ�D�ױ��	8�����OnS��c� �'�)�qu
�2�qo��VB�B�?I�nXlxVHYEB     400     130?\9�ǙK����A���ӋO�y�-�&}+#(nrB�m������AB�ʠ�\;JKi(gvBTwA�ў��@����!�eګV!�/:{d��q�5�>߮G!�teI�.o#�Nӌ-�<�SǬD'�T�v�exh۰��zt	�m�Gd�Y�AS�u�J�<55��{����J���_�y$���o��B�I��tjԙ��o�SFg�5n[��`@�����o����H�ڡ󇘻]ލ�ц���N<�`*�0����k���E�7=�L1�;��S9�E�a�߽h�;969O�`m-4���XlxVHYEB     400     120����Jx���'���Jc�񩱊��W)���4,��z}��aGa�A�/��0��{7��*Z�hHV���K4�5����D�@�v6u���
��k�*!^���ç��l��d̀�ː��k�SS���;˚:A��4�@ 7Bf�x��MG��c���i� EL�(%��^k-���*�9�~�èT��0��~��H~�ip���:�{���1;�T�5�Ʌ��Iʭ%�0��.�N^0~�$����x(��Ĥ��H�hB��Fo*Z����"qJ��x�_R&{XlxVHYEB     400     130XH�ɥ�X���2����PG�ivur	��"�Ut�ۄ[:�g�X��Y�)�t�P����4^���������0����=���=��,q��^��o��a�1�@z(�׏�MP͵�˯e{E�h'��{�_BI�� }����u~Ķօ
9����c�J�{ԥH֎��_�d��p��z�g��� ����h���g}��ԡs� ��O��������¢��t{#��e��ђo�!Ugx�b��M^:���b�B�L�&Ջ���taT�v#�O��NR;�	O6��Q�m"�l�t���7Yr���=�P�XlxVHYEB     400     140���hA�)�Ur����9��k�F��%sP��j���|��
i��ٚ�#�H��=i7=��C]��H\�YUZ�ů���78��-���@H�%̻�Zn��ܞ��>���_�	W��X�e�%�4���8#,g�μ�5���uJgd���
[~{��s2����J8w�Έ�vKT9�;}�&�.5�#�+������D��rkRYw��9Ȯ:��rM��E�� ��Q��~�y~��l�8��3�Ƶ<�rLϾ�[���и�$	�Au!�o��lM3)�M��6�na�S��ˆȔ��7xӒ��p���w�XlxVHYEB     400     180��Ε5�I3�{��$�b��n��x�� !+ԗx�����@������S���A��՛��:Ѷ��w#J����B";�/&��N���W��TL,�����'.C;�	=
��1>CnЀm�.��ɲ�$+nJ��yk6p�܁����Ʀ|�H��%ı�i8c9ywY�Vj�T��g��}�Z6���� �;�:]��[P���ͨ���8��N̯���+��f��]&@�<������\�4繥��x�u�yJ��r�"����-�l$=h��
sWN�>��~�m.<tww�/�=\�����FFG;F�{���:������R8�j��c6k̕ÑJ�����x75f)j �9n[ϓy��T���+Q�+H�XlxVHYEB     400      f0��j��`��oEǕ���0N�
�F����0�� ]��\�Sjt�iQV%���J@s����P��ȭCC�b]�yOf:����7z����k�J?T���r��ՕvH��8bk�xO����M�����#[�*��<A�߾�[BS��o�o���\;M4(4�^sZ7U�i�WL_s�����;H�F���r
��ӪkR������'���Ֆ��|���68ƪK� ��f�9�:Z�O��P�XlxVHYEB     400     150X�f?���^�8F�Z}1R�jT�_�`�M�I�S�ʴ��fW�y�GU����b5�����u\��A&���5�{U|� Y���3*$hT@3=��tө �& � �pE��=Ы�U�b܁A�K���7YJ��x5N5f����>M` x�9X�y$���K�W!~��E}p~���V;w�,���
G�FX��ִ���E
2�a�4#d��;O�P�l�㡲rA�b[�ĉ6�Yd��S�-����Ԋ�L=�V�ӽ�D.����N6�~v��Q���g�Ē�ޒ���B�Ǻ�W�e���*�݆���DH�5�AJ��I XlxVHYEB      b5      70����{/<�V#�L�Ro8%*�qڣ�)q��.IHc�Kӑ�y��جF�#��V�N�u��wΚ	뎬O!r"��"�6�R0C N܍Rp�=$f|��]�[��bwf����