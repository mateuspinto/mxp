��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ё����ԩ{�x'�ݪ�PN����wR*��RhV�c-�	M�
���v��TQK�}�xN�>��b��mhg �`Ё@
�α�`�����!6B�r��#elԠ�Y�C�$�w�)�r�!�[����6��ӫwc����L�b+�#���8�b�@�̪�Du�S��K��:&%8&�#��!�	jkʺ�mg���z&�g���3�� ֣���� J�Ĝ�h�;ҳ�%��ٿQ�Z*��i���/h�Y�t��P;y膫:����~��R~T8ӤK��C0�eg_Z>�o�?��;���*!u�ώ @��}�&/N#7n2a�Jkv���,uD��_os��T��(���u�W�3>�f���������8�z�vӟG��?5roqb�_ǅ��@���J/ѯF-\�p����8�6����V���m>�����L����άR�l�hڳ�!=����И�V3��ۯ���v�ڪ��w�c�*=�#�h�����ђ?����}ya�~g���z�	�ˬ�x,0(���s[2����)�?�cF���<��_)tj�vK��m%�b^=l�]�µ������-�J]aq@�������Y���C�)�un�/�a�c������Ur#��Zm�I5��+�����x*=�X��o���h'�n
�'�7�G8u�5/�p>�(�ҟ����gUy��갥�T��i�	9��P��)�=�����'3֙���ˇ���Es��'u���Zt*�����څA`�1�経��<w6�{��hX6���N� ������yI�;��8]��P婱��L��D�cP ȅt�^��n��,���c�w���0v?L�
�:r�YL}�Ҟ�G�a�S���J��G����q�9TPd1�ɥ2�f����ew�hV�����m���m|j�S��虌��A#��4�\e�)Sz�*�o���_�ʱf!31,u�[	Ͷ�k�=��	l�&dV@����8[�(��t�ҏ���xy=q����+��,�1�ȎdFQ���e[��Z�.���7Y�ϓsf��.�l��0���% �ή�.���+�j=��ּ�?�U�*{0�㌫:q����������x��>?�	*K{�ٶ*�m� ߜ� �h��$=��=ɵ�`ӜJ\խ�X�h����u�q��RLKLu����^�����`�˵CG���-Ej��4��B��"���mh���$��i���hɜ�z���{aL��WH 	��)Lj�+��Pzb(Nc>�Lٛ_�a#\
B/��ﲧ~��ܹ���~��{� ��;��>5�6����E��A��������V�,�=B������4���]�c~UB2B�~��7��;�،I�3�%��C�yR��&���"0��?�e8"Ԁ���U�K\x0�v}	?��"E�؍�[\C
���GQW����� wZp*U['\L�n��tMWwr͵J)�qo�}���T)��K�;�*�N��;ơ�U�\�/a(q'��#Sr7�̸�_���1�ȯt�'���(8�v7A0Rr��7a��~7�o��ӓ�e�*���[&Z!�]h�T~�_As�# �D+��x��g�A�d�>-C����	:�Ԃ�T� ��ڑ��H��,���Xw E� T�Ϟ�"z�R+���Q�j�>֚���b��NY�j߆�BtT���bS�y�he���W��
+��0�������w(m��Ӈ�q�Zji"o�o���X��Nűs��l&�	�+��kƹP��7�J�x�_�j�t���c��~k�Y��;u��9���F󰪳FN8���T=�����|��%w�1�Y��j��A����t�$����'���XܹF�}ic�U�
�u*�����H���a,�<g�KA�|a�?ts9�ߊ7���&eDZ��	��>/n���r{���Z�1"h�`����_�k$���K5�\�װ�0b�%(z�:z���3e�d�?DRT���`J*��sKS/mmhy��K˷znéNT������qBr$r_69�a�JP�Ht-�a�����;:�D��B�sZ��jt�ǩ���p�A���ُ~;BYs����°�Y���w�-���Ws;��;N�d�Fۭr�+�o�F\�\f���W������pX�0�������	�d���F��M=h����V5�
>f���&JC�k�u����eo@9͏���K@A��y��	B�S��{6�}r�U�XE�O� BR�9�Y��FJ4���4�A<�-8��'�x1Uy�ܱ�����"O�	@��^��P��� %òu�q�qh�}����2j���U�h�AdG��o])c�;f���Yܾ���z�0��h{��$�`����km�������b�
Pr�D��w�gƔ�*TB�A�_g�Ez#g�A�=��:�>9W4��A��h03�E���#�U��%΋�7;�|*�y�I��'
V�7��5�<�~�B�3�@�|�^�\z�3=�ko�e����ئ�|No!�"���	$�&	�مH"�����W!���O����|E.`����s� ��J;	�.�^nc���<s���EG F(�wg�L^G�[]���HL��ݛ<=m����tٚ������A�g�� �����撟���W��:բ]a`�0�}�T�mY�=�D�I��PH����_�[��־�POc�`���1�� �V�N}���L���oO)�{�Cß�S2��ϙ*#|V�?�e��P�4�A�̆��p����2�P޶i��B�A�uKyT���X�4��g����9�E�JD��6��&kA׺��Gb�m?䶒�B%$~zm��T��`'˲G��>���f�&��������� �N�NT��ο=���&��5�or9��Ʉb��e#��L�ee�?dU���\U��{`��Q96���/�#phm)��X�[�)�o�g�z#QOROK���DN�������i�p����{���\���A�H6�)�>s�eG�k�P����*�|lr�����<>��`|��i1�v�@9��V�]a�����K���r2N��OBw�諴��U�h<K�+���8m�W���u��� ��*�	NcWp���������b��ޞ�6:��*a_x�и*�`��tp�!���h��N�VUE�B�Q��ۅ�L���.��	���Ʊ�޶��
�PG�&�y3q�3�b���z�`��Q����������@�ԅ w��_��k��ò){ f��,�;��V���It1���9eiU�� ��_\���b`4�Q _�����ZB�&�i�-?�Y����Z$G"	"	�=oE�0 ����{�6���iD�Y|
�t4�
,���õl�#������
: �$��>�:#D�V���)8�L���p�6�BD�v�]�pb�*t�0�A��b�x�<��)�NS���Lv�|%PRkӪfi�j��cj���䕈������o�6!	����x�T��ۨ�~�	�m��͈�ʽM����~d����t�l�܅"���,�.3����h����p�)��-G��'˥��g��%� �޾�#N0�h�{���(���������v��I�2Y?O�$-����0lᚿ�t�`?D��_A��>�z��
��� �=^^��:���yS� �Q���mX�ӷ7&Q�#�\bU�Ǆ~X�q����4���o+�q�(�ybD�MZѽ"�/YMj��%bz�1
xJ*x��Osl�}�\e�/P�0���W�#�N�	CY\��f%��H��"��Y���]tJ��v'��q�0 ��NQ�c�湦��#����!͖R�!U\&hRə��WE����31\��+�N\(�D��y�Q�4C�"��dm�{	h\��Kz)��i�b'�`��	]v�r4�3�A�g2[���U6-����ܸ�ph�*~=E�bRF��St,m�2��X��ˣ�ʽl��J�=;�4^5R�r�uo�ܯ15A��i�}�+9M~����J�K�٥�MJZ47����O�W���1�d�D���L��Zj5 Qi��@2	��q��Vvǅs���Е���̻5�,��{�o�l�6e��M\��q�q
?y#�{�[πc��fm���Űp\��ZI�׽��]j�}��BAcM.���>��Å�q'���wg�a�nL���غ���2���N
H���x
/��7-��c9U-)��b3yV�b��G�i�����C8?4� �+-8�X*۲��n���o�b?Fsoi��"���Oi����db�L(V�.1�@�1�!�y�|��;�8�*��6��� Y��ߚWD���DS+&��,ꞡ�6RѕK��`@m��&��ߩ� ��_.�P���Pi2�ᷰ�c�N
u�L��gЛ��~|l�Ņ̶)��ʕ*=���)ߛz�_Ne�M�]� n�ӓ�A^V����ʖ�W@*�v��<��vi�V06�$�EP��^NeC:g�QE��/=����b�����ۍ�쬩��.+m�?c)!$���\2i��5��y���&e��VV��xь��G#ʬf���\W����RX�>AX��v"L����U���/T
lQ5��P� �*i�d9�\�W������a��Ur4� w�h|u�1A�{�<u�@�z�B�g�����X��.>[ٞ�q��{7���XE�D.���t���9ҧ�0ך�c$zPsg]�T'�G�/O8v��v�M�E���������Hpq��l�;AE:�8omY��\��Rz�+d�CH�6}�dJ-NtL������uft����C�S1��sXw݈�¢���i�8�>��N9�� �����������={4���enpW��o�>���ѼKE/!��F��hq��V�hrz��2�JӼ�Vw��H�:Q.��V�趁�ՈZ��չc�6����T��U��� ]�5�M�E�MN` �@�^n��U��- ��c�\�I�3p����/�|�;���hȪ���e�.g�Ɛ�h*G�(��H���9S���`t�O2���J�V!���`�Z��:#6�����-�gN�&!HN�6�e*�Uߕ/I£���^)6�4G��IkEL�;e��:Q���P҅�۟Z>��P���¡@/ܗ�kSiK�����4�����#E�*����쀆�F�خ�U�7ߵ��8�����m��7Y�L)�+K���5���E[���� �h��ZK���3�6q�T#s/��L���ӕ��1pCߩ߲7�?u�"�c�	Q���MN�J�cZ��UijTJ�XK��һ;��������l�s����3�h�'\K�'�{X=L:��T��ޛ���"u��CD�P=��O*ϼ45��w�$�'�9����_��(���ـ�H���ƥ�����L��{�T�|��i��2��������[ԝ(gaVrg���� k��.��+/=�u�C����d�,zi] [j��#� !�rz��!��F�-=�77< j����Y��Y�t���L*t*�R��XHe��;�5$�/�]k�`�h��-b���I�,�w$h���>D�����qC�s�2��ػ���Q���_���W�e8^�=�Ǧ���@oV���v�.�������V�3�K�>�l�AOv��'�D�to�άB��`%�k��%8uG�]Y���6+gn!��ˌ'��" M�,���x{Yy�3���hmR�ɜ��̵ W�?P�?	w0d�r��yC�����󧱉&�~�f�S%���m���GȢ�5Zv�}��V��y\'��!��9ey:�J��*�]t@#�X6.��z6ٝaaH�4�9b]P��ĈtQ ��g��]VJ������:�k�ޒ��F3ܱ�w���Ĺk\�9
Qg�H�H�s	��1�u�蒞}���(85�e�^q�sm�����Ǯ��Ձ��>�N���#u��0/�O,�����O��\�G��>�Ħ�����9�~.|95\�E��|�) >c�uO4�lL���§�2�$�3��H0mר��JM��<		#���rj�O|<K��+�Ed/���}3*F?U�w�Ƞf�	�ylw�}��1ogɤ��3U�-
d*-�U�y�(Ŀʄ�.H׼N��22�.'h{w����i󡀚�C�29t�s�
oũ�<�{-�a��|��"ix��;B�%�"'>*��#�0̜��4�BCW1�ԙo���1t�S+-�=8�wB|wv]���ݏ҇v�[r�VڬS��M6R����U�
�4;ݗU��	��C�d%i�oA��q�B7-ר,����3����]@�ٮ�Ӵ!���;9S?����ԯ�M��?ܔ�lVf�N�=o,Q��N<K������_�h�����ի��3����z�X�C�[v�� 6��.��e�zQ�۔`�R��O��p	!����K@m���� ����x�8&���w�dх$���W��n�Z��Q;��.�e ��c��Ռ�� (PpUT,��<��a��	���Id.�SjJ\P�^@��r�.�	gT �v�4��-�����\r9
g��MC��IG�LU"+*�[�^9��"��8����Ӗ��$ �(<,���:P�|�N�W�%Z��k�0�{	� ����vM[���M�ą�J�R�E����^�@���2\C$�jbgD��-S]!�*j��8�'�B�swHhQ_�'b�\����2w�XA����J����>�v��Pٺ� �a�fsm8��B�9_j#6� A_�u���~���0i����$D���y�}_����6���b��F������s�
(�n�
h���ͷ�~�/6P TQ�˦�S�md��唻�.�2�l����
�4ND�lX^�M	�Q hh]~̓�3��o��5&D4F-E��蛤!���8�h�o�Ƿ=>4��6r��JUQ��U�ja��QnW�����i�
W�rԕwJ�1_!`�~Cױ����0cx�Py�J�t�?=4���r������Z|QR~v��w��m�i�ޘer�}»���Q��#�	4�8�
�s�J�?����� �(E�5n�DY�����5^84uZ�_{;LT(�z���>M�}�Ѯc(ݷ���\��ʃ��u�N=)<$)<p+*�����
����0M�!}+
��j.3�T%�b�z�'7��f�䁡�R���B>�+������a=�	K=@�����Ვ�������gx��"#���f�\����B��~�ë�]�d�#�����c�j/��e�ݯ1�Z __D���X�'/��M��WMOh�s�<�X3�{Z���*�ؿ�r�wV�]K�����|�7��`�Y��Qv����3�Hq|t��D�cu���9��!�[�O6�
 �T�O��v�0���A��8I�*@Z%*:�J �����V�&Sqd?B6ε��ˀ��t���Oꅵj��n��,#>L�:L͠�
���4��#�e��&�tz�iR<ޕv�!�#-/���ck3��F[6s��Ћ*�0��h���|}����6���3��z��9[�!�� �U#�Ι: �,���iЩ �W�&Iʌ/zS���1L�i��؏(�`�K�ei��Cټ2��Tb ��n�Zҟ��.�q"�����q"�NĂ�m� qӊY�����tg��6g����4M$%nʙ��Zg\�zX6������ hK 9�+�?s��5�� �9H\�I�;�̾�^`�kc�E��V���?r�.>o��	���h1�N�c����0�Ż�J�
��6Ï�nT[V�w���������W���	s^�|�TJ�
J�uU��5D��ߏr�N78���o���H�����Qi�J�;%[�G����:.�$p��9_1`�\j͊e|�
y�
���V��C�y��LVi����t��a�(A�f����0j�=ES���Y�V�'g>¥�mI�B	��Y�}DQ�z�Z��W��͒���L~!��u>��s��B`	����j�_8KSN�^B@�Ax��w!��W����ke�\1���0�ȷ�m��=��ͻ����Hǳk���^�
��!r G0r�0�V�q�}d��ł�G�n�J���t$0c�̈�7�+h0š�޽�y���Iǌ	�[�gAR&F���ye�ȫ��&�������"BjK�^��x�5��K'C#��F.��.�Rg�p���/̕�ш���;�f�����j�%NT�U�ax�;�=:@D�,@��Tn�=/�c�,։^�=V�5��T���m�	&� 7Ć���^�j���fL�:�>1ElRpU- �����Y�B2s�[�#�gF�N�`<i�3�#h���#uL��SQp;�'=K��U�@�T����1l�뇨�&@����p�a*����W=�H�ڏ���ÿ�����{��,
�-�E��@��R-���a��u���`�ʊ���f��]L�����ʝMr��]6��<ZnZg��=�n����vY;S�R�f*��d\	Z2L��]�n�NHw�̬��_��쀯N��z��y�<&�45;LnG#�b��id�&�4G~�������I����Y��R'�xQ�s�>_J4�K��o�t�ėݱ�ft�����I�*xG�$0�4�i�33��Hk@�V&�ª�9x�θG��G�G��m���,-���@�Ig�7ك���ߔ�c���M�b�Z7ߨ��Q��N�]�,��� ǣ-9tyMF�c(>Iym)����"����|��p������=�Wu���dG~M,�۶�K�?VGߍ��_z%� ���cv�,K&�%�����}����yVta\���fh8j�7��˳�H�� �ny�D{c�)u���f���Y��˛�]���\<1���s��')ݿ����rϞ���P�|)��q�>����.:/jo��ۦ�W��quX�=��E!s=*������xE����
�J<b
z�wǧ�g#)�~�v��r��f�����eB�����1HK	���������KM	��� �X��k���X2��6-�lW�R�2��$5L�gm;&��:�i��}��3Ut9�;�SR M�����S��+�)Tb�j3���(Չi�� WBM��g�m�X'�h=PǷ������瀗�j��!��:]�N7v��VU���ZhɮU��H>C��l������E�>ߗ�-/@C��U'��r�M�����f��9��('��k�<N���\a��pL�_�J��$�4��"�{���s�^�;���O�Z]�J�4�����ܯ��̪NNq�A��7���6�޷T�%���#�X9Ʃ��g���M�!"���½Ayi�F�|�����Ma�L�'��8>�/`z��uI%����,��he'��ݔ�3�i��c���:u*1>윢��)����U����:��k���'K��Fon�cY��x��?%tR�cN���r�y=�m�� $)�-kxۍsACK��~�U
�bT����⧔"����OB�T����VN?�O_�Ό�p{'rݗ�E����m�H�����םV�F���j�N�En�ݞ��ȕ92�X
����4�R�ɡ�󉲸 ��R��r���u}�:�j]��Wإ�CU3��=L�����]p<�����u��'�;�KZ�Sn��fu�,س����[���]�FxK�)8�ٸi�:)�*V1��()��{W�`�0|0m	�ʬ�ˢuxNju�3�Y�U���;�Ab҃��,M�������x�o.�[��M��w?�COt�5��~��<��7�����%&fO�s#�/L�$�N��P��l����嗈�2� ӎo�
*�Ⱦ��μ��ع�t�qKo{}$��X��O�ݘ��D7�3�S	y�T����wD�̌8t�#��8�nL÷?�{N �tU
hn�e��i3��%U���[��If���;�T>�G2��l8NO���F����x�������|���K�4h����h�d�(��ǅ��+�f���7>�}~�ZG&P��e��@8�m���Ǒ�u3�s�4j������8�3�<㛻6��l�rc�	�-�EK�R��ydon��B4�*q-�he��5�;1���6~ ��!�����,��Փ�#����v[C��7��k�K�� �BVP�w7�t�l����&<��G1�:%�r�'�١	qZ|���ЏJc^4�M�3�M۶џnN�S��<����;	4�Pj��:bI�y&�=����q���\����8��	�1~����i��1�L��+��%�ץy�I����!kmK���b:�?�5�vz�F 0�0�@�����~tʼ��)kz\3��9��9��Ђ�f{�H�Ggo�4�:��^�<5��A�?w~D��
��*���
���G�2�韠Dz<v�&@���+&U� e`�߈����w�M����[��Gj m�[F�Y�S=��~7��\L^i�2� у#@uz#����5�U���W��.�9�T!�Z�]��6X��ۍ��,�� n%�(�����Jܭ�ּ]�S�|���ljg��&�9���B)�%�>1�O.�ܔl���PՌ���_�<RJ��f��xjK��X��f�J�)*�/�3�-�N_1��a�F.�P>��Ug��_�*�β��	*�5	�jUF9�Ċ��A������ʶ��̖K�F#��s�WZ�Y��"j��S��]]�v�
�z�L`N�NU�?^�*�F���A�9����ug�dD����|�h!�K6�>���I t�t���]������D�6(�e�.n\" �}�;��tގ����@��J����%+q�� R+g��xj��X�܆Go\�Ŏ��4P!L�LtД��H��!�G%� g��Q�����G�TO;�Q]���\�%
��_�"����@�pz��:ֽ�5q�L��,����{��ط�e7_�1�W>�����U��*8$�z�7�}�B���l:��h+A����Eߴ��x�$n�`�B(�ڗ�̺Pʎ��95`3��T��a৪��J�����_�SٷCJ���c/e{Ȇ�"qg�7���6�ԭڤ�N�t��+��ֵDQ{9��=7-r�6Y��ˡ�#�q	}��;Ĥ�W� N��^4�Sؼ֋#YF��I*��z�����b��۪gQy�V�	���6y�AVS ��������-ss��yr>Ό����:��X���i?��;�(!�����t�����-i��5��1���K?�N��jF�A����O��^�*'rD^�u��B���K��w�E�034�8�ϴL�DR,t����l�3��^f@p:���h�AA��gbov��\�����N ���U����|���#ꇠ�3��n_~d�X�#NT�&���Z�Q�=x����Q!��ꌳ>���j�*�����߯�o?�Lq@1�Q�F���i5Ҽa�ڜ-F����)8qY�E���ü���y��.��Qc֦���~P�.�b5,Cw"u H2�Ts��� ؀O�Z���i��o���{��x�)R��T�/w8f��Z0��J��<���qC!ؽ;c$.`��¾%Է3�Ȓ���`��8��%��YP���Clp彘Z��(c�.�s�&��
D��_���vS4�ˮS�=��ByM Ӌ�;Y�(�@������':<v�T�Y�E��a�Gx���q�yA����~�1�C<�J�L�PB��YWUe�x�Ƅ�8�׳#����� �Vk3g4�xS��V	�U|�M{��U��,��Mr֑n�U	�f�"��yαkօ1�ʨ���H:Y(��C���^��f*V��^lsf�ǡ�"<��$^Z5�B�!D�Gd��M�G=�(
���}�%b��Z�W]>�hhJU�����գR3|{�-$M3�} Ę;E�	�e9L�d��ࣹ�S�c��yfN_�?��qV�FM,٬\�c�	Z��Ab�_�9�B��f3M��Z���Vw��/Nl��� ����h�x^E���t~zC��Z^}�Ǐ4HU�t"��������]�c�>g/F��E������K:����k~��g��kY�����f��Yχ])8��)�#G0�:�x�`�;�� �E����@H :�����'"f}��,&�x�����vT=��'ؑ�αm;�q�
���@�+�]��l���X��`M/\�&�1p��+��P;�ov��A$k�x�h��ͺ.	J�ҟ��&&�� �,g`0	�^ �3q�f���,���iG�!�
�ds��^W2�A�ϺD�]�D˘�Wu�"(O�6�J h�N���Gb�ZdAM2F��ѧ4`�>��?�L�Yg�da�'J��# p�L�;H){���Z�E�hР��d'�Gx(L�:�S�g��3�������ޢ���(�?qnЦ��*3j�f0Z�JpP��l<ч|r_��d��k���H��W�
5�UD�g�K�����o���u��͓��Ue�B2��D]�a>��d��p���%!B��9��an겿�~[ʾ���`�5��M��X˳ �˷��+����efۭ.ʶ�d'b�Ҋ%�@���5�6.��4o茛Q&������
9鼏�pT}�᳁���~tRF�s������#��_��H��[�vH^5�휄�jf��P��W'h���/8\ڼ���x�i��d�R�D��87w�{�� M�WޅZ�gny�2��w��w D��������
'b1�t�]��y/�fz~����e��ufA��N�G����6A�6��'��a�n�"I��kF̙J �t�%���6�V�W�e
}D������g�78���7���lF��{�*�"��d�t(Q�&�N�A'��}lyC���c��$6�ҩx-�(üJ�(������,�n�y�x��է=Az�ԓ9?3s+5ɣ�NTm���{v��2`DG`9𶯙�5&��ї5��M���n����S��4��k���_m�~����.���=c��K!�b�7��4b:��cd�?�2�f �O4����6S
�/����KHF:�,X�"o�=�M�CI��G@X]���h۵ǂ3\� �F���Ү��k�	�k^l�59JὪ�#��.s�2y,S�ЧտC�$,���L�a���7<hF�amN��[s�.I>�1M������4ļ�$�F	`���:��U��|�$>Q�9�6�@��i��?�N�g FM���5��O���=��l"���o��_!���ɨGTg+۬�"�c
t�i��J�����Hy��d$[-��u���Jv�\X�7p���H=�~1 iB��j�Ĩ�^vQ��i�շ�t�=��z�U�� �עT`X��z�8�X�mm�1�icƝ�\�1�ϵּ�M�蛰G�Q���fS4�B:d�6��w���O0���鮈�JF:;[��E�i�W4��[��mD���A�1�𤥹 j�8��&5�JU>��^Z�-b�q�K+��Lh����Dx��g�Q���<@mƟ��k���8�P�E����F^���}����-���a�&"o�%d䊻$M��/�V�����M��ʦ�GrL�Z'�cG��ݟfC)���E<��cE0�l���M�l�a>�����m��3n�0^��pbL�����	��G��sV�	�=|�Q�$C���qc$�"��w;�vWsr5��z��+sZ����C�4j�Lq�\ܼD�M�x\v ��=}�=���U� �&��i�F<7Eijj`���̽aF�E���f����0S�^��
|������hYUQ�&q(B�7��D��7o�@�_�P��ʹ2䚻n�n��'�響*������_8l��9[��8�{0�k����F�>��Ȕ1�m���h����k�h�G->Q��K� �&ɤ�C_�r)�]�L�ǎc�³e�>;�o,�4�}���^����ɦ4hj�2���9��L����UzK�ϭ[,kz/�MW�دiV���-y'�`խ�B`t+x<��yQ;�ᅅM�+{!�PK��3�o���+.��M�_�m]�"���3G�N�S%G���;�̦3��0�>�iP�%O��g�h�ѥ�N��|1�ա����21ۉԋ�5cL��.CK�ZO�.#ED� ��ۻ"�+<ew�dSg�Y�J6�Yl��xڌ���)Zx�7�Ѐvru���m�~�ɵx߅���Ie���/��n_~�_J=p&T�jF�J�A�D��%kM+(3�SIO*I�gKOwf�ş"n�%M�} ��Y��>�8W4X���B�ȡ��}`�G�ڽ�;�?�����-E'��	�sk�����B�3����~-ߑ��K����O5�d�u	�.�dVL���}�s�?%�P<e�����(+�ل�Οi�E�oT���8J��ݐ�o��y����|����q���;C�Y���'B�`��U���ʚk��.�w�4�6e0�I�|������!n�ϫ#FJ/s�'Zb� ��{ĕ�#�r0	�'���xց��F���[���U��#�~ؖ�J���_�m��uq_^b�Ib�<����jS�I����;z������lt_���k�-�TS�q���D�;���L���I1��-o��BY/���I7H���6��t�{b�t��iZѕKg �lW�C��³��y���	̫��r>`{�v2����q��.��%Ұ�� q��'�_�v�+^��+bW�rp�N�9 !P[�q�z�j�XϿ.��ozX���xW8�[�]�>h��\F�کO��$;��+� \���8�~M���L1�Ior�>ܻr��o\6a�_N��ƘX��u���g͟q�6È���Ԏ�uK����|J��u1Fm�5b�ju�_�f�zw���_34�rx�(��kTܘw���&O��U/��]���Z��N%���M?��y
�נ��2�
�C�q��v��w�o��S��>"����c����ۀ�
F#L�\�Fx`�^�����!��r�2@��]`O���Vyi�e�=�ɥ�$�O� 8\����1�N�˙<��Uv4����i1P<N�BM	h��Z��o�U���O��J��`;��W��r�<�ޜ��D�G^(v�������c�mёg�7:��)��E�G����Gp��pU>��֊dwi��?j���o�?Q���c�W97��7��XOB�_E��7v���n\3�oa왌��^���6n�3�Z���"!�Q+�FV�j�;�=Q��?~]A��c;`���ӳ� <՞ψ��a�,��r�0�w#'�ލ5�3�k[z�~�b6��w±�N�u�l`l�E]��dVU��y��G�\����!��W��\�h�xx�"a5����m�� a�١�b>�NQ�´�P)ȼs��?�p��k��)����͐D��Gku�	��,Q��B�������)2��~ndV��f��kk'��Tnz��΃_:��(���7�>�]����4��r���P~/�!#F�����>�ub���4�Ƶ�|~X����J�AQ=���c�������´w�f�����ۍ����������4��t�+�ߖ����'�?���p4�Bb][��צ~\;�ԣ��\�G�m�E>��6�a�j��w�$�\�K��J�����3@�A�&�1y�=���,�Zk���R���$��.
�a;�S��D]�VS�7��L�q}l���4%�CH+��x��Y�6�<��x/����\�9'�Q
�M��>��}���_yu-�����آ-�[�_\��d�ƯVt�����������TmAX��}A���>���p��X����XY� X,!]��s� R�l0���}���x�r<���v��p!|���J�����:�gKQ> o�����m�@�t#�/��y~�;�KE � !0�B1�x#�R[��������M�<���{���|&{�bD�/~Z5���dk�jl'۾$ن�tC�V��6��:�;#x�Gڒ^�?qaL���Q\)��n���n;ꈺ/��阈8
�Yj��@"_�HB��ܩ��3�B��5 �A�дIv��r/�WS�*��Dҥ �ˡx�4��ś��XB�~�Q����I*=3������H%�&�����:�Z�0�TJ��7�@}`t.RDKe�����T��RM>�c�GuN��.
����l
Wb4��>���^J��9N�Y0����Gʫz�],@���\�j��Ƣ�H�կ�� ���ɯ(�ַx)��~}���rXR;�1�
Q�r}Ag�sKLt��0�UHV��Im&�IZ�R�_�`M!�Du�n�PC�bTc+�>:=����юM՘{Lq��o���'�W~i��񻮅�O�/�	�O���O�#�f�7��/�؊��*n�i�,ꝝ�)H�������`&E$��(���|�ӻ5�T��ho|��U�fj��I���]@=֗
 ��^I�Y�I��IeI�	k����ē�_����VM��M�����:�t�u�?	i���^�D��i��E�#���:fP��}lӌ��C�ŏ�E��^)�z}�f�Gё
9�W��i����1u�#����Y��|f���Y��u�����5N��`j�`�#�S��5ʥ�ݛ+9�_n��6�����J#�^�vQQ�\V��x��i���0�ʬ�zi���P9�˳��&��2L�:��7����e����1���)|]�yn'��'$k���..��9��ζ���H�@����|��0F	 �8V()������C�56�����N�)��̀E����>�ؓߔg0���kr��@3'�k�m%�փ]�6_��u._9�?�SA��j�k|e��,`ˌ�}#4���]��9|�	���b�޷�Ku�M 3+�ڂ�L��.�F��
w�0V.CA��c�޷>q!�����_��f��K����ӿ�2���@|h����Bgo�iZ��R�Z��"m�t��E�-Ѯ�4q$�_6\)<��JީU�������֘�!%�2��rbI%G8/;?o�:HG��O	h��˭��گD��^8�X��h=
��	�)=�U'vC�l�2UT���b!f�yW�T�1a'��~M)��0�