`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
osR6ZA9/JfXc+QhHq/Fq+zhs9n6vgUcyC8BjhbkK7rCik9GbnwJO2oyF0IEG4cc/hj94mfajr/rs
7bYtqZxyMuJ7kDi4hgc4g0W9+Uu975wrnq03Lv4YqZF9fJj3hg8hf7I1gHQezDTPJgAbZ01HmJph
wf2DKeT+K5FNE6nx0XYv6Cm0vsC4ZdUXWypMP4uSmHp3v+Oh/pRcbpRrJe/KGrGM5ZhPKfW+eVyZ
FokC4ZFm7j9EUR/umxf4LgXVHVLZXTMLxSLE2YkHA/elppjH1/xda+7WVpMJ2aXrbeQlFOwntk6b
TRcHc4+VlqcwBjq6ySpqbX8xS8rHyCcVpw9gZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="66RHWmgzQRXTiF7wJZ8ugtVqv8cXorE7Lg01bDScU10="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
sJBiNzUCP/1GPE8r9O3xPzPyGDpTiH525IluE/CL0Z9LoGd6QwJA2oqWx+CAe3xxKSW/B662N9ew
9IAqBx+SfAC0j3YoTjP9Nt6kh3Ibq6VhCQP+z7aTXZBzBrlN6umpE+ikwoq9uH1g4a9dn8vnOqXT
q7LRbb/5VMDC4I1+iuIyRtVwtR0zftFFJymns3m5e4KdCuz9ZhEzYl8lxmzMeQh03kjLfYUBzRjG
Ffdmf4l5vcoY/hFDY+f70qxUotZeVnin8SJx8UCPYcJ73F3i4ih7Zh204DqVaDnnmHdqlB1cW1iP
9XNSAb5BEJyT/gjkkt6siM6jMBNG01C2e5hn6sXqQX6JizwfkzbcScyO+ckZ26wdWH7Ct9aD2ljo
ZOcPdnfgztY1MdyEP+Ct7baxzlFOgrm0Vu5mJj8rFMxP3uQ79oUUAyzKKGQUQzhCB+fQdhi2E0XB
wAvxHcuyVzlz1HRKI5sbtMfwdaCpDX8RiwTHWqLh52Lnqke6u96mPsfe/lz2M+s5HQ4CNLSezvcL
YVEj9UmqXt3q+ZgIp1EGTVrxwliC4qabiIoW7vYP6YhK1AoVkqskGegxAH38/9rlqPzBBbvtH/o1
+o3Whio+EF2OxSICr0NFspQX2a25L2q6pWYc79U9HCZ+Gm6oNMkWcetfimyRUjay+phZi2LQHBJI
jAcmagEH0ze7C5Fh6R3zM+sbJj4hjzdLqyMNEaH/pANFbLvUelx5kGiPgAYGgRAhysjZq5rAHXjE
QvU1Bh+L4IfkWi8YTp0+RCSrQ54H6Ol9LrIDzsCsusX7YvuiZrbtocL+PbsgNCq2PzgWKXcZz1/u
OeUEC41ZmN8msLtblKxav1FX0l0zTqtMac2RicsntYhwPqzxTYnUecdfAvNRxXh3WbpKOx4Rd4rl
IB50Ln/QARgKqhhLUJCCGJKjOT0LPp/gtXU9gXvy018hJ+sExNjPUDhWd9mWoMGp9m2DyyC0ToiX
rCT1ioGRatSXT4M7jvldZ3Yxq97vEq8jCdW+uoMQJbWStGBmzcjiseS077mDVyjTFIRvz1XTK7yQ
QDLgYBkYqrvZg8fEPQ9670l45CCZWmIJzyQMG3i64kfLjXQyhpdkSO+2lK4RyiTKuVNZWu1p5bYR
Rn6490vLyWq1aUTyUJDxMsAdKR4NCoTgnKyKSPSCrgqC2GGb0V0mNr9iwvOXVsOs6vEoECbYjNCZ
IBW0ZBd1Y6gMxodrgzEoeZTRG0xBqNluAboPWqHmXbHFmINegeU1XQLXxipQ4wWRLJ5eyySptxzT
6kQqHmC5Fc1f+IGvf2bGaUju8HQqGHnzb/qTlwc26yASCe+qi4jPGymgu/QJoQ3djjRcxk96hM1p
qtLzl8P8txj4CsYYLf7qSeh6TiiBpMC0oWf6yOOg6+/pH8v4sSfDLSYeRIaC47AC/GcICNEdxt+I
CH21P+UemdXmF0MI58BKDq8eOQY0IeOa+P05sOWWy725Hm7CZphIVhKy7T3ain+POq95ZXfWQGGI
LhULBLgUUlxF0OFFbHOvLAKaoa8+nY/swJUkNP3KDBdkklegC3KKWJ6U5Rp+4JpxqT12St83LPxg
77+K28XOZ0IXivW+tDQ9VzE7moqG5j/ag5RK9GhnAS8ggQFrPsL5RkuhuVyFLu+v0jBZDFGtcVBD
Cmun56RnDH8LRgvdEVFW8FmBq31tBqvifGgGi9x3NqF0Qb4mIem/jWO1PqFf1BSk2YBo6QNFDwuQ
PlzlC94n/z3id3VXwJnNStstLRylp2qyBZu9qyYMAdw4doVook/GvJc0r4qTHvqbtsEOdxW9rvWR
2FiRKjdAntgoXVwJwG+Sq1hvzis1NBSKLwBT3XB/IhSfWgNfk7BBMwLTJovYWM+I0uGCscpnt77m
KWV18hFXWm0Qyg4bH7EoCJPlvNFDXIFW83SNOcKXB/k90a8ZQlM+Yii8eNftNgRNjGxBmMu00z3S
mo6DZcnw6+mw7TEgkI9b7cSy2w2lStt3Hgard/ohdIeUM2Qf9EEgvZPpczTYXFW/9gxe0DKtt1cT
roFQ8A/NjKexTECptyIagsRMO4E5J9LJHOL6cJPZuYwaMasXi46VuEGtm1XnNEmB3jIzkLeiWHJ+
WOCEBajfSb3fcL3OWCQFNe4yx7tQjSZiX1neA1BaXA8UVTqBBlHLCvDYp0XmrOTGaDhtGQhsI5kO
JTvNlp9RRjTTy2IdO0KzqAXQbyjFJrMCTOEmxfopCDt9eY6Wth28GUnPpMtng2VeQb/JdmxFLsTy
SChM2sTD+cXKf5gMLUyVPaU+c/2OYtTwvqdfOHgkHIvjSaCfMXXSsCkEg6421k8ZJzzzTU8oszXl
+Mc9yt0Q/nSjLeIlmtLX/fcPKsHhCXJLYgNjd597+n4cqw/lM78NvMLo+97pFBYWFJ8c1rxdJmn3
JPxnTssyKUZ3EcmvUUBrXXKv0gF9wI5cEM5y+7CAeSNgDg43DnpEZfCXTBVELzsEiSfK8jBPo2cd
aiZkNMTTtiO7LDhZhYKYXCBV1Llw53Z8gAcEO3I3xLLb0xLL++PfoP4LllyAYSydX6MN0yaVC2w6
yv0298Hv0Ev3MexH9sIiegBbniXZfFPL6pxELp25tjdK0iabEOnQhHoBZEHP6HhJc4LrRs7+7kG7
0hgEDg+Gd200ifGDBi3ejOc+WFDj9aukp1smY2/6IEK6BziNOwV47tnTA029fZXdO8YlnZpe8io9
SANJ2vdrNKpA6iqUwIBwCVYOaEgTJ7oyWTlezdnC8JfuuUgHGYgyzDsHwKnnd2TArRIJYyK+/WQL
hNVF09fqpw5BU8uuYhN1UiOBkbYxTiEoOh2oBCu9ZYciTHt1uuu2KimFFi9USXhmslvcblKlnvOM
19ougduNaZFsYQ8KhkbDlliyU3h/puaVAzY552JqYA8ISn9SXGziRqRZHT5uYyfmZT8EZLWsupex
r0z5I3PE5AF/rJGGNHP/ELM9Hy9FfThV8lXdZY68OnwTtBQ6oLbo+Vyg6iRZk6z+VxR5X3irY/8Q
UHoT7TiYPiKoOqZZDklIosRpRMt6BgYYqqrvh92olEuGD1dRnI0G6vtIo27R5r1CVY53ogJGXYc+
SdsPtnkN4wNJYUkBcyGzq5ULEn27+x3cGkbNal6ximdVj4rG8DgFvsKx+cc31Sb1BOXVxRHOI4Ds
df/HuBAT9wB1LffpaAFQtpN9EOm5jelIdFggAOETjhS2f7MiPfDEhmTfbJbuvQrHJzzYHbAWfpRe
rZ5T6Wrjw874QESy+N2KGUVITnl/1Qx6Kbkd3pedsFbVO5TCq/RNgRbl4jdILrJjJaIqEEOunpyG
GwBI6F67EJQcfESpDcJUqfIpcvWDX9id77+NGuzNXeB9zbbOgW8GTrIxU4TQ1ZYmg4LZBNMUFWJ5
v4qy/sgsm03sNSqn02VF2SV9UZQt8ZyluFJ4uJg7evGaIFScbrKxewt5FXzmi11jbS2HIvlZOKan
83iPqKJj5fvQEjvYPBXQ70TRrqcCjzMhpcJjqOIdtxkGa1aCvvOKDxpptZ6nHPiZsyRTgsO7xvNW
el2GAZghu4WR85pWuPBpLWdBek+e/UbUqLrtSoGqpACM25cBzIJdGzT/pmvKfIJcv2RpU7C0EKEg
XaucllhZenmwDTDZnGD2P8b4cVYV7j6Bb53YKB1DmhbaTlRCN0WIDMa7dIoTle+hA3JbwnYrD+yt
oLl4wR4i2L31s6n5BBWEU1VcTTuQyApuwUDNv1qOnjl+ytOMjHNogmrktdA3ouDjbGsGHhf1sXrm
EavJlQxYIni7e8qbEJgMwD5fAQdxuQPhPupgCXdOtGbEe8sYv16feGc/AD3YwQ==
`protect end_protected
