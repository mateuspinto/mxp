`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
sGlIVqnV5mdrdBd2q77X0GmLKnbO+SDIDb+cw/UmfOIN8Ej8vfcWTFq10UQadNDHMCIGxdiawauc
QgHIPwjSQqM2y8bj3V9HCZ+fFQLc3I0/pQdPvww9+kXWP1WKs0vw7v9f8CHLMCFnOpGdFY4/BJQa
GT6UsSa3z7VokAWT6XdMcLDGsfFf4ZQAwZI65IefeKauaEGfFVJddkD8MIq+0LxBFm5PDu8Rytnb
5W6AMwFweVk/30gIlASAkVotCLTi+fudUgsYjloUOVtuxPkW/qfC/HHUdCyL3PIAj3nh90anbv5D
DbC/3yz/zYBsbrxU0rsWNqhYe0A7386yUFVo0q6rnb6vtIy49dDIDSTEVL/NsEWQblGMLH4Mn6ZN
okwospY1JBfapO6PdRXaWC0VG/Lb0TJ9rQo4Q5ZM6re+YbH22/7JStyuQscKgY5gKhgV78KhmiLA
vNcENLsDO2h/J3D3f9nTD0fY0ET6kKAyAUkxrXPku24rW058Mgq8D4GnZ9IY2lI4gBE9stBqpF4a
UekmCl0Ban53sfs0tORP6YxC+1Cw6C8y28G1KgOskFSiQMizRdqUuRJ7HaGRf8xzzREbFJFDAjqJ
TswL02z2iPnY2CV6kVlCKMHHKopp/3CiKAehbYf1SQcylkMmUb0uWIXBPei53I8d07KljCMp3dD4
vlmRIdSRnAxs9uFa8AwD8tzBB3HXfVpq3aoc9Qq6mjEEFYGD4A6mKFpHRz0K8l4yZ/d2hrOcvWhd
YMlbciWBhOrye2kw/gzWmVuekSN1MkdSm7cTLbAn5xg4rAwk5q2TPlsaquSHnI/slsdlhenq5Qdp
kklYh8+f4tvg8UmhXE61pQ39aGUjuYyqAmnzkkl/ogAifDPsJVNd23NfTJqN+ZezQGzyFqhRz+ZZ
SQq1fgbw7faMjQvZD0/i+UgKC9knkMH/iyjn4Qs9YlW9X842psDPs10AxiPa62BLkn5VxlC7OLqs
WNcTAPO4tS07VSZaCgVrHgSJyvDzuJy9zJzX9R79zoHej1qXqNvOpBLXS8AzYfOS6qKIYjp1kJJQ
1ZtI0xMAFXPLzVlv7FO6VwFjf+iQKaWtOgconqzOw3TPf7+wDCf9AUJOI0JlaCLQhZQY7WYTQDGR
gkwCgDJSRVAt6Hccwu/h6mMeL9K5xc/scpdA48QRqjJeqQv9/Wxxzow373vgc9rMGaVi0kqtzn6k
wqao/dGUWwYYGIdd039ekLlYTrgDU1Q1cthYxKUzgJz0cjGXsMc+xGrwm6TN8KItwbVhxuq7A0Eh
X9Hm2r7KPJ8VLvYndU4sB1gMssvpM6JpC7E0PYt75Nm2cYfW6RZ0cpEqyUxCDW+WCuiklbF0R4i/
goLYoXSJh1QzSUzAjVEG6ppFSQxaYOso/C1JWOdppPzNl3crmGIND22PUlXBv4s4S6TfQQ1XhWav
R6aqLArZKU7ARVo+mV9DiGuK/HwgVEbK5yXpubBudkZIp1kZxjA7Lc1ZY1/Ep/iDs6jn2vF3rCff
1ZRfN0+Idq9MuMCn+ApVrepMoXk9q1YFZ7+WuPpbg27R4CajaaH8oQLudQICquKyAhjjNcQjHgxe
0gPOgh99vHX8bCCKWyEFYoAwwgeDnS8i5qfFLnXAGbZ7HUNqnjlLnoCDS8PyFDDLI5ka/KYehAjL
PYmPL5THCf0AIXLjdyM0aJ6L4BtsS1EUd+iViJldny9laKuCEsK0GDI2xCDFj5/Vfhqo7BA72SNO
oV5xMRnUPZXrDZ6Jkvl5Eu2kC+J+n2pCDxhF4YrhPuPf4NyLzh5U2qsmWhSHgW2TZH2XJAdtXMqb
YOR0be/3IGBv6/o2SiSt2C39+Un5R/kAs3vVAlsN1TBcsxrDmZ9SBn1BKLl3Luvgg+nUu7I56/P8
UWor7GwS0cQxpmanKxZb/8aDAaxF6F4Uw07KajN63/9gi6/vhLfkbH+PksweaQGsNmqwEvTt841T
Q2kJKWQnty7gfG+l4WcCXjQed5+I9pNPd6woCc4Td7f+v29Er8yEN0wOfsnHGO0avW3sPhJRrFHx
3WZLh76c5XaTPN90gLbMapBpkWXD4uG1mStvUMC8RkLG+OBG+RCaXsugop21
`protect end_protected
