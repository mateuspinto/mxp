`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
nZ0ElgeZfpf5/fUg+kt69EKeNsMLnmjzKs1TQaitYH/G8wboYaEjTraLuzJsBYs0MJfwJDHQoR3X
CVr/FZGKQK+MW9FzRFpkW0a3OaXbrifA/jc4MoCIhkbFRByJYMZkJQCcXesqyeKlzhk4UdMWhv55
Yiir34HAOiLb+6KPYWFha1F42wyehzU5G3Dz5HZstjxngQMh9Pd7UOJspKAiXlzxrBP0fzFajRDy
FeY6AXlQ9xMnRs46TR89Dv8wqpcpoIwlKyetppAb5/4gGCNqSfvix8pRnYheFC0ERAgupeMnufYx
Yt1mnBkmD67I7R7ZbRHQLVyzm0f2tHzruc/vDQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="spKPz58jIm9gH106Wa3GvsvLIhmHN6d1GKfaD/fz7CI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6512)
`protect data_block
W8EagQsfH0Kj+remBFgq2EBj+lCE2XyshAKc837NbNwCQqMV+iSJebIGk92LnDGiIXs4q4Qf9feC
gCVz8HOe1/Q1ycEqxyh5XlYpACWGpFvSrkkaIJ0IycbFWXBwFHrhWB4HAV/tFycM/DaXySp8wkvb
o8ega3AhO3kG5q0irXJUd6aJ5d523ApJ6+gnm4ok+QwKzvRyWSjhDWK2F7hs8lnYRBdQFSi6asrj
QKSy1Q/9seUDF+QX7CWuwMsuh/HKw8eU6fz1aRwqJSYLYFcfCn6uSu7EFLwCSm7xL/eRv0jLImZs
tq/4SjtTca3ucFf7aFDJABEnfyBzP+3BvM6Rpazyh8RML1gLNwGXEgG8msBpII0zcaJVXq0FoF3U
Xr3lsxl7Va5kVE8dOcVOG2usfU49lgO0TMltxtg1v052HD7QX1ameVYbA634L4lf947rgtw9Qzdr
DHbAt5C3eMtqaq/iZTIOwXayETJX2wTv0uP6InEBSMLPeUnWxLew5zeJfcWCssnaXcnDv0jr/uv5
tm4W12sqHVzfvoMUuPIyyV9NOonDbTiEUMVqh4WY3i/XlHteou5vv4SaESHOQsfqfKHLXWE+H3Uj
lYqN0tGhou+Kqzly0W7iSbHB4wp4okmaqwsPqejC1WZpRiBbgan9Y9H5HmcCmIv2WOtmgRdGcfJO
4utJGrwVsSc48JgswxUNrWt2/TNtoiYzLvoLAOmmGqeNvs/omNdK78TXAd7/4N9rKpIqLj0oLYlD
xX+ayr5s1ZRttS7r3I7W/ByDq+VBEzxn8r9YLAHr061ifCUrO5DAqxYu/PjElJuGlA7qgglzKsYP
KYFQWyT1oHMBaqPyplHRHSDRVsPptfkSl4KaZ3RD0cEJspk8jPK0BWrGOuLl1jDnJf6WhPfmDHEI
fISZeCGCM5ZCjYeWcFPnD0yMFDwAUv+saQ8NEk049wsw5h6p/14o1boVH81GNxU6tmZyync5ZZ6Y
4CCxml5lmfKvynYOZrMONUqMGVrBp35wCzryWzLCBnsEaqmu4SjfvSEgcn9WR4s3Dd9hZfCUbwpL
61yD9/Hx5OjZ7oa9sHHZ05sx5fjntgTt+7W1RHUJUVMgZDBiG0K1vaAf9cPmucoh7qo2qYMK2Vp4
T20tr3w13PNc7usAr3eTmATUQPP9FBWQElIlLbANlh3/iouq1IWrh++5cDM1sS2ybDcNszHUfR1j
CXiPS+eCttZRt/Q/wdRnvMsB/G5hUR3JItVlthZtKsjT35fSQNoIgnT8sj5Yu0YJRluPD3Owi6nl
uFkgcIKlNTn1XSFdPsXiJohuz8RmwqHnCndQ3EsQkGnYVCTK3Os4oS8I6MhqpBBxYLzbo3Yu+/nW
/hPccI9DxLslo05FzdcCeV/0lcPoT0uEdzfEbUQpaoCcWqhdDA1IogJ+8xfJZX+jbRTJzYm5A4xQ
txYrZ6cC9DlOtJBCAfiycTvGyNcqdaDzelTCfbZZiSf+r0KRK/KLWMjqSsYNONdszAM2Dxd/fVJd
0dfNzK+qrLfhIKPNWRgEMt1O6I1nE3sv5j9JtCRdkY33nAYei13waIf2YxzcG04AARmOe6PK2/Vh
XAVxfJ0BOhBViUnAwW9THFHGOwnbkOfcKHUH02cL9Pj1muhbcm1bhoVEop1vtURk4CBFcNwYdmO5
mtjjyvbn9Z33TNH1T8dMne37SHK2r/7lhxUchk7scQNKnh5GyoFgVZX96I7dCCpQNuWPaI1Jr5xG
8uZ9BEBpkAcPVpSugcCiaccfiM3hS+LJVp7UQjXXFdqLzkP61dNhLZHmCWambsK8mNgJ9Z402jSX
p4k1S2oIfQ/Jo9bU/79NVblHJqaWRIeP7K3fxbzKE8fYyTxzuAqwxyoOaZoQ4GP1Vz+D4SscboEE
195bzk+Gz7dOUGZAbBWmQ6+OYGJ1mYHYrLOaJJfaGB5re/3vMwG/33bqTtLzV5N5em5lb+lB+l8N
EyRMboValPSrb0rZb8R4cY4panPNwf2uzcB3UCuKrbqFto6z0LYBr2WTHQj3mZZxvrQdHM042irY
Hr2YKhQ/7UdwkAR3DCJyth4GXJ135MGjUQjueEtYj7XbCfhBtXwXVA6Ck/283qZdL1Np2aywM/so
pXs8bEHMMC3Xl4JTjVUglJvSe8TIRm6eI9F16aTIxB175aVZr8ijlPNvE9WlDTS32OZ+21V/eV7c
+gjdMwYz3ZqkuBC7P99vTNEFgptUfIvo8OhzbPg3+e1R9FiEf5XS9KFWy4goKFUPEXNI+XUOddIo
TiBBy2lMPLUo7lXuldOUwTFZ/5z1HHMeK5JJRxGVZKtSnX/a/ivTYe0BXprM924GmGMxI0pdDxJs
wKBVXkv+5dqeY5Af5X2K++pTE+fISao77x9tiNxDC2tZX85ioapA8qR6zaSgYbB0IpV56b/1seeb
jh5aH+hzmPDsB0DLRokYADR/1xaSBJdYkQmCJz0SR4I60aMl0mEqECp2+M14Ssi9rZGhuLDFmvJw
8DxsARUXX6AkirFVgSgIQx5UWvZy2DI9p2YpGuXkJADSq7XlyW/CO0rHNEI09oRaL0115SArxX07
oUKRx0hm8+pzrgHruLcs5Eyf7tfZ1Hw97dVdIRn9LSIFLL7A4+SzO0vpLP8vGCPddZSUPlcOYq3q
APmDJjuFxFmBgRVMIeRLuRBqzUL4P1ZmeIiqn9jJAeR8ALBxCeAUQ0Q/4g+Yaeby5bWYGzO4UbXH
rjUW8RJWRV3+rkSZsmbVbuPLxux/vT+imj5z5P/6urr1667y0LNx12pnbLDZUlDIxzATgx6X2lU6
0Oi/ZvYugiJZZ3XXvvZY7rbC3c3Ri6osrXdyhq9jhxAGrta5jEweeWqPHG23DameCopJOUARQLSL
ZeOzlbrMEpwHqdvGd52kICuiAVpm9Op0bO8cRLMQYsJ44B7AiTe+GpWp8ISiVSxT/Lxb3NaMAMwg
rrd4VUowRrWnZZqH6aZ7AASoTglnL7kuhQCQOieMZtsIo9jlX3KfouQSkEDkhc1k5USC3Syp/ocV
ppdBofelvpNf2cF7ZtSQp90cdfvO0Hdt4Ck76PM24Rer/eAK4lHs5y0Qzgq1uV4UGjI380OcGI7+
+jAWe1MxUCCcHwhva721IoRa2wnpar3luQxpTepoSQDkg5GeC46fPMl2y7jS8tv7eFUmggORYjzd
q6HKkllz9vel56MtNa5j/9Wi/kh4w3e5M9lBsB+xTUp8gdBoWB2UauX2KDSZie7vgqaeGyd+a8gT
WM2Q44k9r+LGwfOIz+uXQQjEZ+/8IyFlaLK10Oa9b+sc/Qa6qQRmq8BF9PJxSkfCsPHVSb/1JUbn
epGwMuDZ7RStDSElryx8jZ0ieK1mCQiYaL1cZxRRh4YwLH3huTz6eUZk6TWuBq7yQEDHcVfwHqE/
wx506mjSbHSnDlspGYXSIUX6aFztd1OWsvLvnVTKMthQ5Zl4shkqB9qc/j0JQKTJLEfkr7T1yvhF
tQgSEMsL+KD3jF33hJ6aQTiV7NbmbUv900SCxMErVc11YPJjxMTix6gUlasFI8MNaVfhILaNoKaO
7Dif3OtMOPjqnn/wL4xspX0uM2teFJax2KTJFvQLyRxIEYAhRxnN4viTLC+R0y3JiAlA40trfCoR
acxdzaV/G9/MEXE2CylQEJ3IIi0mKl3DZZwJlLDrzlrdzK3gs0Q53yF93iD/uw14DocvJTW6DbzO
yeHA3a9eEzjIePPteGs5UPAvjPBpLdfapiwasJrDn4CKmXTUF8ieoOffNeerGrvOHx9qI4mf8WoE
KZG58vS92NeN4bA2pTHzsFaYGSwJ/zSEg1T3AePhwekU+UlHvBFciJUShdIjxSHTpR+wKUPbbd4p
sEcFD5NvwB1pUdbbGAAEqmHHPXZbKfmJnrFxTPX3IoGSbPuKQAZFDUYMIeBTX7lsP9RaCQMvFSj2
R6IRdQbXO3xBU7DGx5oJDuVaYSHsQCFRHMPUtYypZ7L3acNVRhZh15omIxU43fo7mvTEiw+E/Xpw
D4QA46Cr7x/5vNeqkgc16XR8AM1GjkrUW7nssuhRgWx9rnH1dg1bqHH+DQwZMfCgGCN6awmbO3GK
Cy8Pi1bXsah79A0i9AFcHzwwhwp9I5SmGbp35W0xs+iGWmmvR34X3fPGzoR0L5DVdNcJdJVEtflk
WnOfbBSSmXJP4XcXu57n/v/WC7/GKeJr04sIgiW62w6Wn+iBdggPpwJ/YQ5eiVZ3eMA86Z+slulh
Vnc0GgWc45q6LpA05ahHDWPvaYpqOEyXplPf7+zIM+0/7jrd/cBmNmqL/uRVfiRCxw7ghBZSyz3I
7X76n1y4OkdR+xyjBrfcPDflIiwMtTKRTaH1QNQ72ODhNiPNpdvIlIQlj92xri1KfNklkpwbYNNb
s3ZrHdtYhdBbDGxtjT5g7eYe6HR3r4WqNsH9wdRSUrcOPYF1gO/khrrsJvpJ9APxkjvnfGWDPaZZ
41l/5FDdL5m8CXVGSBcyNT2RyMpYPCp0NK6PfpVkXu0vJdU2WvSIwtv8+kbvRRp0n9N7jJwRlmxr
G79rQ+6wkbMkCyCDmToMGiCjKLlrXrybO0HSMiX07rMCs+kZnMATYoSIxVc1GJMd9cHg7g996emO
bdjVDx4zXwoKO1d4PPajOXMI3Z42XPEY+qNvmskPPgEkJAOs7IPwNHZJtQRqRs/+iA75bV4Yg834
RsyCZs1Ojh9fZvgnMc+VMde02PcVEP+LtnUXm822GGmIBngBRGGrOIcBV7PD1lNcA+t94rY5dLgd
dWLRFqIKEhKTxrNTblKFXwQp2uX59dk5VQ9rtJQycxAfVLO2sVa98J+EoSQLmtR8K1VSs1BO4YHB
pOaqocpD/es9yZJtCZX8pL9OZShV6mZ2xZZbqoCZPTSto+EfpUK78qWnXvYQUrSJ1U11Jndc9Wih
yWXLoUxqq5SHn3w8Ip78A4ZbtF2kM9fNsueAi+4019q3qm5J7X7Co0flJ+q/4+fp6A9Kh6m0kFjN
dHwFj5HVBIxDuCo99ZHvDVhnSpwykf6uKvzgFjp4F441vWAMrEw7sUQ8P5WAXS8I7fujh5l4I4s3
CJMw5PRicOcJT2R1r5jc05qtzAl7xiCghszjMIkaaAlJBkw4IHbnjEn0CkjHuNomdqx4Kzl1A5xj
2x0KD01Mn0TKjtMDGRjMIqGJGWvRiTCsayo3HInt/Wk30kzaC1F/xVoAtdWtDpzjXpCjXc3gWmkk
gX3w++o2WspRuUjLuhcxE+Se2Qqi/bbj1D1Mj7xT8H/B2nTBxQo5P9KHPSG03lb8p0Jk+wcrE5rY
XvrzYZ2PKYMA4VtyapXPPHTwyoxmvyGHb2qN2sU5ATBuCX49Fqau+NODVwUWa9wwZq7fb1DcaUsq
zgZeDbXuKU+k7/ENP3DeFst6kMLyF9Ij7sHzvGbfcOaKQOQz9glL3lzijRxsMtHA2k+6DmUdBjEy
yP1ZEGE0+5iWMyR6AU4bE/Y36ptn74/lvO0S1kd8vbptfNDb9y5bQpdmA7M6kyH4T9Opg8BcTemZ
5n8UVo5dZ9Q0D7K1eAAvK622CV12JqxbljT3ZpZQcATaQFy2ocCFmctqVJSy4qg+1rGvu0lXRC8d
3h/ptGJGKVZqBD6+K+y3b/vz/TkSRUoZxhC7p+IncfwH3AKlBV0oNI9fWeqqY1DiC6eBcAZbn1nL
ZhTX0Q3f0jRLY5b2SpwFmOp3hcW4W96dUBF7Gu0bywhDox+1OjuJv6Zqn2u0Q//JbahnNKxn+YeV
rPsVPZrY85vu2/DX+5qWUocjDD0qKYgTxGgRcoTbS9NRsLiNJ4Q9gz6UlQGN0IJUvShtAp+FI8J9
CutQGTuWzl37DPSRXCbOKtv8FiJpD8HlwhtOaxk2Eg/2clZM0B5S+jOeAlvbQX3RcAuflKxOA/sE
jQQ55nCLco/SWuqXNv3qUrW2BE17UCr7G+q6os9Fl1jEgN7jLQH4eIfUlCt1bvF/Q5YgiP7cprrz
l48iFTdd+kaQ27CueNiVHlLgq4pmlfUdVwsB8vaNXype7wc3CACop9m+C0ZPN/NZj9Aj+2qwd8+z
bJUE0QggGcFS38srSO+xBZlzv/MJl6rqQbcpot1dJTCzBbA1DmzE/zVjAEVgAWju4JSA9ncY1YPa
p2S1iF1QNUtDFpS/GQvr+0m9OSVGQS3bmqAPZzdv1Wn1Nf0Xic39YeB6Flj1FyvVyRdWMfTHdrz1
uNCYaC/VGoSD1uS0nPsynWRwjEqPSKWvOiilCR4KN1oBX/3yu3IHE0zsb6xNgggGWRHD9PWSvE4c
pdlzIrudfqmC/n8ZA5YSdDPpaOi524s5pvb64Imlw0/+IyJeosZQgoEj3HszOsubhPCPRCX13bcD
iQJen/XbqEulhRRDRtgrU6l53Lt2xiAOe0FnC4e1Ftgks/p5I27BwdfPvz7iIRZCYjf8EQwFFJ0Q
/WwE2309Ril7yuervkwXrp/cG2tTPYqkZheFE1v0jWsqa7TNflvEQ2cMrnEpr2qkJ+th6MMy97YV
HvkSZH8gqLZK9xKVB63IGZUetf+npP4mZBPTRzzeJ8JnY9ujg41HCYdC86CSNKPZ7Q0/8fBbCPp4
5EplWJ/S7iI3p89gW0FFn2SmwP4EZVK9yvW7Hpu/U/XetM8qX8oklxoS9N3KuVDHygpW/+lds6Xc
kfbZn/LiEghE6jK62Da7Qhpayz+jujDqd01pCgqqY2SThZSnMew5g5viQTsR1Ciz2txlh6afyFo8
15HxCNtDKUyO+bYewE/QR0USXRUBZxJhYnyqJMeFM/6Dupnu4a+FpqgW1WL+RfVksI6gozyEpGY9
KrLapFropxkCw0PXuNuyzlzjO9GhyYHafv4OjkL2FYmeyVMqoMhDehWYc9Ddd19R7ohTDAjAyu7T
4aWM2SlPkTOp6pL+j3YiuRtOI2oG84xRtedLc4SGfbHISnQ4NA/9qMG7uufb9SwpnIKNuOoFkknh
jIOS+dj4fhZtIdDYhD0IUpg1nnz9OZ4y4tCWNjC/CeOnn2KqkpbjYnZdrIbd+jGAC57lP05u48PA
Lshv8+U8WtpL/bPJeRVV+LogZ+cpXavqNp6oaGzixq7hx3Cca+X5vT35n1cHAVjraPrwbVWMrGGZ
9m19Ga8yDll1YbVEF1+4ZlyPxrymUvBkYGcmpFSdyAFkHD8mq2HhkEIPQQZSdmPWyu5ESxVLFVq6
h4dIMPh+9NPtKoLYsVdfdBB6wNg7QY47Dq5ZWzHErsaZZzKGMXbxkMCEjcvjW6SGzCdVtBtFiVCY
F5kpXTyAprVDc5WOxpY972Aw46nJxsrTngsl8rybo54HTG7DXf0gxipC2AMYYpvYRbuKssh0jCnH
Wxo76/O4ylbvc6OYWTg74my0I3nq71zSJJRF05B8qhG7Iapp0OznKI5Ulk+/xdZKQLR8kE0jgb5s
xFdb9FmZGpQkAvyZ+ndu+ZBbnARM493AAoS5Isy3GKhvzfFZqas0DFA1R58/ljrmUNxU8Ljd2Yfg
JwytpCi77NDVDzK0AJe8nLBgWY3KomIuGp3uO9Iyi1Hjd3uViKk0GcKauZXctKgvFScWaO1Ehz5U
6vlm+UMzBDy8xS7MCHlEDbBLfuKm55LXeVyUB4jVJxvxID6oh4ZrLvw31NZLPjf+wDm1c6UBNYBV
Wul7OpHcfrg/02Q/j44pbSqynEoOOmPMcbNjiUYBH/0U1H1taQbpIJnKZZOAld1b0cB+dedkXF4m
zdIYpVB0FHbqzPTGCfETE+a+dYi+DWG7c/uc38KD+Uq1WtKGK48LnsWNCv7fA/BtbC328MafROXE
XdPYRqUKa9/BJnO6il10BToKLDrqWYTQZGe/jzU1iIiVIDTdUT+F8AfwWWE1EUyV1kszeCY3LneY
qcprJimDUsAVYKl7qAfP5hCrnvspFoZvmwy6NGWoX/aATTYpezNp5T67LSt+UppkiCPikryBzV4t
by0J2E6xa0G1HY7oXX2Qace71ziRZ2HppO2V9PJErOdlYAAnR9ZAYWGTJ1g+VNUd8hSA/okCkYod
3JN47e27siGAObRcWIvRc7VY/J4KNu1NeGyuDWzct73FD6lQT25ivcURF7G8KUf2PcGTkx1ZEwr5
zOut7PYj6LV+VUTgRF6twZE/iJToEXguqZwRvez8xbNhBsR6zGF0uFgmDJvyiGvGFqHTlYImgYWi
NQjcCnIHorCDQUsIppeXZnNq3eBLsQ/g6JuOBURsEFNqNFrHhqWp2xqtxORnUuAtFTE1rgsny9OQ
90w+CrWCsJXDC0GGPMgxCsb73ECOUsvW2BZzBPhdbSWR4Fut1Er2/sRyWjYu/kNAlCSLZ/9tAzbD
P39GGpJADZCH2XPWHV861usfgD9paZPxH46zLM3MtFVkoPwZc4cajGAoMAEaR4upH3SZf3tHxnKY
0YiqOf5iF9lpID4dcQFYo3GRoeX3594e8uG+CHKNKohlZFeBx2QdvZ+pR6pIq+p9RA5E58adIhqq
v/jsJSgkrCl0OUF0RYyYcKE8KfgkmGBuWHdQik5u7nkQZhw1IEgfw9t5KghnK0k0lMDCwOrZxbad
PzBzTrLytMqD5gnm3jmivn2twH7JG2oOvCNyHipUEmUSyTb1sV3klTGOnSs3O6vUyHfPqzfUoENs
+6H9LFj9axIV2R8uWAA=
`protect end_protected
