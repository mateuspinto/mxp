XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[�BAǁ�O5�?�\�O;i۹��z�;��阁r�b���Uy[#���$  ZQ��ݖ�6���	��`퓲#���:A��Z˗��-�[M��lے\�2{Ĉ��Ւ�}Q�9��~��iӄ`���c��ۜw!,��_m�@��Ҹ�~?�S=�}�Rd��w�|�wQ#u�C�`~I���	k��W�gv9Y]��U1�;��5����碋S�y�w�Ox������u���c�(���s�3�쨖��$S|:O�@�ى����	��f�>ꨗK�;`G���"pX%"Z�g��ae�:?-.{,0m�&�'Q��$���Rye�a�Ŭ{��>O�q�/���=p�%�h�%W{���y|�	O���e�U"B�7z�V/��+GxV�t/;��]^���}�]Cޏb2W�l��w|Խٔ�8N�����N����QE8��"���D�1�ʾ1^�QMa�8��RN`�mHn��9'%��q%���-v
O�]Vo��.(�%�0WLӟ���
Z�ghxZf����?p��B�jvO7I�\&F�w�VC�	E��'ݓGC���:}��H^�nwx#�qjn=�V��Z�Q���U Iq,p���J/h`������3>�1����ߨi�=�����؋�"K_q|�,��u��5*{��%@�6��Xק���O0rOA&m1�U���9�֞7}W�.6�}���p'�Ǹ�5Iu�-�C�����s*v���D�%kx<��uT�毁�d D_�Q����V��ԙm�����YX1XlxVHYEB     400     190q\��@ar�gv�v"C�މ{E�H�2���c��;M1z�O�l}��n��w��2&xɶ��H��?���\��$*T��`{����o�ѭ�m���O��{��Нj��2�����t*=��W�N���=���=�ʽ��ta��V�F_V�����a��r�!`A$�&�Di�yg��]�'�.������z��������JC�Ƃms�������֚�L�<��\�t�G�V��]���}�oP��9���� B:pbvGA�J�J尿T�z]�P�r�h�����hSk�m��2ճ
�y�!{��twxpO.�w��}R(H��#;̠k[[�$�1��CXz��X�3ܲ}�!2肒�$rr����T,�s'������XlxVHYEB     400      b0���4Z��˦���_"��=Ja! >��X[�J��TXm���*|@�+��=D��Z=�N����"7�V�ⷿ&bU\��<]���>����d�bLR�v����EF
_8Ko˲����������s�Y�F�#N'��Ӎ��$ ��r�T���8�s2Xp��"M����]�A�C XlxVHYEB     400      f0.з=	 ��ޒ�v�w܄�����	%&Y�~�m��[:s�����C(!��^YN���24߱��mB�e�K�R5�r�V����+�a�`��~��߳���}y�/*���_��^3��p+��'�%�&� �d�(�t?	�x��o�/@a�s�݅VAU��ݝ���G�g=�v�D���;t�#�|�^%.��%��5�O��O~Τ���jV��>��LW=�z�a�^;W�N����XlxVHYEB     400     150oSmX0=� o !C�� 3I� ��8ܴ���9���=%F.L�^߆#�s]�;{Y�>�)۹Ja�������+(��y���nU;��m"ZL��<i�G���f��i�=�0
� ��i�ve ��J_�z������Y���jl���;��<�P3o��a5x;K ɘ�,6��m7�]�@*I��L��W���m�VR.@�H���cZ����b�F�38����O"_� ��pI	��@+tb�dM��oS��r!`$ʲ�_���6�2�KO@]��R;�j�������.�{�z@i���#~�E��[_h������Y�l�+���XlxVHYEB     400     160V̑�9���#@��a)�(q�H-�a~�r��n�iZ��f����V π�ʭ2<��>݁O��.w�2�~��c�6N 7��5PikRʄ�����-�ىÅrY���d?�Jy���''DР�킚Յ��9��snM~����ZX�U�'e״�v$;�ъ~��6*r���̻	 __�u��s��9Ǜ��FW�?%{-��ߥ�A�JE����}1�K�˟ZK�T���k~�&2�e��d}�V�h�5�lO�F_!���wts���ɿ��x,�$Uњ�(�+�F��+�v��6�2�V���"�T;+���C$�K� ʣ-T�C��τ'ݛŗv{��J	�%z�~dV���XlxVHYEB     400     120 x!Lb)OZ�/� v�צ��jbG}H2U��V�T	2�Z���ˎ����_\�}�k��{D��3��jf�bL�P@����∧5k����4<�ɩ�4v�-C3��"w�N[����b�O���o0�}!!���U�̜�"'�7�8�q�0��㔦h�Z{]�m4��7���5�A��Nq�1t��x�%�ئj�~�!J�j�~�^c�!r� vq"�S6Nk�R�g)0���[��bvnH�KrW�C�P)b>�,M8V�G�`L}:��1_��|f�(�dXlxVHYEB     400     110�7�=�_��=���*��@8FuN��fwg˱�h��5 㚡!�iK��b�E�?˅-����.��3��a1f����8�����w|vң��Y��_�N�=1�O(�h��sq�h��o�ž*�@��0TҒ��>�#�* �X���=p��{�v�����o��=h�q�Tʏ_�ɨ�:�7oY���r��;�k�:$�I[�\�S��?F�L�Ҫ���x�wi���X���YC�)d7��v�s��h�]SB��"��&-�o`4�T"�6�XlxVHYEB     400     110����E��I!��=Ai	�Dg$̉8q^�cilB`���|P'N���ib��-�"�|�F�y�E�=���j����D��ߙ�me�ՇRr�����E������V{W�CɑC�ͤ����u/��/�a�#+L��	�ڒȖ�j�s;����-F��Ɠ1��П��g(m�^�6Z��H��6�~��o�f����K6�O�.��jgb�3�0є��gp�C��wmX\���6�5�HDۣW�5N��i���P��n�nRY�R�1	�����XlxVHYEB     400     130�Ng9@��|!������2�k�b;��~������j߮{��]��U�aP�)}�5N��wd@�3���Q���L��i����!eS�%/dǔ�-w��%ks�+����Y�گ���ш���U*�C�@:���1xC̭�(����\�wǟ퇍����P��7�Y@��G����`��)�
��H�U���3H;�����m�v��e�>Mc��/��M9����l�s. � W;��ǖҖ���<����-����4H�+���� �0�Z����6P�Ƣ��·��MXlxVHYEB     400     140��<�CT���@�;>����/��C#��J�fy�|���^4�ɞ�Y�嬟¢�;K)� !RfM����ߤ�R�n�K[|jY}C)�xKy^dG�i�+>y������=(�-f��C�6(��1��=W����E99��m|˳M��RS���.)��^����������@;���e�m�Z	� T���8�)�"x��㥆5��!������|F�<t�p_48Z�{�తwZ��GqO|����~Rd`�H+�û�����Z�%q�Ine��9&�
�	��@gYx,��o�M-���t��퀔eεXlxVHYEB     400     100l�*<�t���M��<��Y�ګ�4���D˲��ģ��IFE�G�ӗl_�~V&�CM�ɸV��=�K֑��:b���s�%T�ׇM�Y�U�j[����-oT��A��f�����e�+^s�B��?�I���,�l�m�z:������fM��ŉo�}�ͺP��+��%5NԻ)�Ga|���e����S�[f9g��,��y*��0cX�-T��*wT�	�T��7��O�e��/[dP��&`�5�	v1��XlxVHYEB     37b     140�0k����x���Y��3̏�/�\=��.����:��%?:��<L�Lӗ�8�#:(gV���B[���s!�Mz�_E���y���x�U�ȇ��@�����؊Z�x
�B����Ļ�+T�s�.�
����@�����_^ �-@$��, ��3b��9>��t+���l|��WE�f�����M�=N�� 
ul�n
t�Z��\*���&~�q��Gc�8������{۩�l�钡ӟ��Ȋ���E�V�!�������S?>.���P���\����t�.�3n�(�{�i�$��1p"s��Ɵĸ<�7ȁR�!�