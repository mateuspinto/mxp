XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� 0�a�a*�����޺�9��	0�o��H�,�\� ��@(�6���Y�<�J?5KB�0N$�"T%`�ѽ1���Vu%���슯}8_W��6���[b���X��f������fu�I�Ahj믯pҼt$#����=E1��Ѧ^��)}�XIk~7u�9���Ê�����{���M}��o��>��x�2S��rD3)��\<�Q���2��9ȰTͽ�+�/ş�Ε��9 � �#�!�$��_�_4(���})K/*�Y,���=���RO��~�!��	�r�U�0j��7���x��q���0X��l��~H��/�Z�Rr�Ų!�G��4gh�-`�Ŀ�T:x"M,���k�U�V�X�j�W8�˝6� /�tJa�фyd�kc.�,���NkF�3�+�������#�K�L����>y@6���u�H���r��"����,g�Qdh��w�
��J��ig*�A��Vz{��\���`d~]�
M���}�4.�}]���Ķĕ�rlF���_��ʧ �5���������4�)�-�P��d����8	��jA��{�+h��v���Xv�����҇ƛq����ǧ8l�$����d���R/�:<@0ɂ��8?n�Вa{�6Hי�I��o���/�<f�D�\)�K��L�t�Q��~sn��?>�fT�?h3\$q�u�Sҁ�RJ%�e������P����������>:~��	 �T��ޮϰYV����j�s@���ىXlxVHYEB     400     1d0�ޖ Dsx�Lӡ́T��=lP��(@��W1�؋�Ƥ�8D_�7�m�I`����~��*�����a`Ț���P���ђk �P���PΗ��1Tw���i�/3z%��6� }"��Y����)�׷��� a_7ma����e[#�zL,�i���ඬ�Fei�>����/Hx��e�ӊ���1S�⻪�I7bD�MX�dG֕�z�&&�8}��HT�o�P��I'���f�/�8/��>�:5ޤ	<!�9�]�n����Nޏ/w�S��v���>.���{ip�"[& ��-n7��k�u��2�g�r�bYM#e��Pk C��ː�01 �v� �M<g��GMG8���uDj��@�ݙ��XmǏ�,7Z}:L�6�������mEqϑ���kZR>_9�Zz:j�����wJ%���>|'��Z�9�J}���W�OoU?�TT�n���B����̏XlxVHYEB     400     1501��2���w��C%@�|���!�X��.�3�
��h��33ܪ�I�e�Ꮲ��P2�*cM#{*U��ǘ���g��|���H��F�U�b��.w
�?���MR�����&L�X��H�-��TP�ŀ�:�B��Rt��Og] Z�ս�Δ~�Bq�<֚����*?}�*�OƖ�S��+2��� L:xY�O�`D�b���T���O���OZs�Vr��$I����d~2�q��ڽ�Ғg	���G2��U�,�9i�H}U8*�~�Y%��.(�9FX(�51���;؞O�}e��.����K��	E���1��MRcXnXR��uk?p؃�G�XlxVHYEB     400     180Ie��"��1>����Ƅ	@���wjE8ec�5��^�^ƥhAw>q�W�H�;�6��ֶW�]ϻ`���&�2��2W�Dqun�׃��#֭����zi�ͳ
n�����AȦ�`�1�_!���@	,��#�<	����nѶ�8~%Ӛ��p�%�Nn�l*�Tt�f��p��3�P�rMj.�y!{z�lZ�ٱ��}%En{!�/B�q�1�A$������"c��h3��`i}*���N�nK^ưԇ|��e���cGa�g@㓲~��K�g�t8J�=@Ċ��]ƅU�5�)K|�֞�$(�f�Z����|���XO�J;�Fȋ�x�-��Lr��s�Q�3����Cv�'+_G��x4�Z8�O�����G'���41�tXlxVHYEB     400     100
\\;�b�{K�"y7{R�[�,X�������nSm���dq0���}�]e}I�u��l�^tB�m�k��=�u��Qgm<I���㿃��X/ɗ�P���]��F��uT�� �ŏg����ԟ��g6um5�\)y�;E�}G3��ڝ�T��E�%�l���g4US�o�'�:*nP{kp?U`�H\W=.W���R��l;�fkK1An��[s��o-+=���{���W]rE
���`�ޚX���Q+%��c"�p��Ѡ�XlxVHYEB     400     170
'a�-������.@6��2���G���G6?�����j,������bd��&��B�m��,I~C�j-t8Zpt�Z�Ʈ�;�%*�ŖRgw�)�5�(��-F�;jM��mf�aR�#y�����M�"��m���L_�y�"�F�@R@k�����'Ę��4@}z��o)(w!�x^�Zo�5��v5�! �oN�~��)������%Γs���������g���;���$t����
����.9�ؙ��6��C�W���6���x�/l 
�����ͬiByj��O�k#�Ϙ_rU{L��0�A�-=V)E��f�P!%o����F��j���b��\bw{E�{�i�����XlxVHYEB     400     160O�������3��=���x2��e���ȳ�۟�M;I�ޫN�E]�[2/��%���1���j�e歚t�u�+�ؚ`�v�g�<�mDFyD\��.�N��Bef���ul]�n�O �^�R X���|�I�L	���V�2�%X��H4\,E�h��q"��7���z[�Q(���L}�uP���,TNtj��f�<s��٬�xA��$�҅���C�O�=|>�LsO~2>��"��5�{͠�+�
�͝q0������s	Y� ������Zsa%��y�1�g�UPr�����K��-�
0\Sχћ���}&�6���d7%'���2B�	�h��'�WXlxVHYEB     400     190:�\M=5N+��",?#O����>���S������6n�j�hj!}�Ǿ
���*"O�6Ւ�{��k"s,�C��a�1�I&�M�lҚm��m�v�{�����qf���]��9A��,�#+m�ٍ7����x*�B����$����`�શ����o{�7~��B�	`9�GY{$������X�9D�A�s�;�F؋J�c$�G�wo4��8��+�*�t-��]^s(�T��I��$.x7�1ݎS:>�ߏ�d����o|��Pqa��{�>��>�dV���3)��z��:n�uW��Y�ʏl��ė]P�����?Ũ��uY�ۑ����r,
����ܘe6�M&ߪW�]�%��R�q�w�.�UD�-�p,A��ηĤQ�o��i���XlxVHYEB     400      f0�y�w&W��Y/K�>�Sjr��[���Ʈ�~/a눤�Tr��H8w�u���	��6l.�rs�wr�H`�`]yS�>0R{�������k����WR�ьXL���eaUP:2�؜��F�3��+�A������4s�j鐉$4Ȇe�bƛ���pM"JՈ����Q�p��mR�������k�v�c%�ϡ��R� �?v=D��'͜���g3Mv�8YpM�0�EEP��XlxVHYEB     400     170Q���C�N?�:����Grb�/������{Yy���/K��a���N�#F��n��먨M����+����*iF`�,�R'J�����i���7oש��/��f�K��+�J[��f��&�ɩ�&bG�xt?��M9��<,#���7�A�4�?�@\��!$v����L]Ey3Xk�r�E���bEțO���Y녩�	�hG`�O�[��&Xm��'F��{\��"���"���3�<ߨ��|/�`����%��[���䬚H�Pf��4,�TRW⭙��wä�����ܰ��jW͔�����\��F���2=�($�6��h�۲)��⤎�a��g�����6k5&�����$G�I����hvXlxVHYEB     400     1c0
,�ޞté��Z��@�ej�}��J��nyn�G�4�ϋ޷^:�����"!����jv��٥�$O�S�B��t��C��R%���JVW���j�,1@��pl�>��,��
+ ��WO��p���{���j.��(M�9B����h���I9��^@{L�V��4��I�<eG��|Jg�Q�"?�ʁ���>���r-�]�S�ak�m����R���O��/O�
7�!�蜉(��C�=��rKz���^�'�)��T����z��6,���a"�``�Ģ�S�`}�?nm��|ԣ4��fv����ؽr�;QZ�(�cVl�^��9JraPC%�[��%ͫ+*�5qN;5�p)��-���A�;�T#�v���!��v�gw�6�����ZNY�WC�M���6G?����?kE
��MSBN^VM!���f}XlxVHYEB     400     1a0h?-�A���q�
��p�*�x!�x>VY�I�S���%�3�S�ɺ�S?\�m�O�W�(S��﨧\��� ,R�ʾ��ɎX�S�]�~�ΰqH:����6Upn��}�������Clǵ��X2���Y�N��"�b
�t�������]=��W�ǧ���y|߁�ɵ�� �Is�w4����;��j&�.[�y�[xb6C8#���7*-"p}(��!�Y��qU�[@*a:*ً�g2��Rh06��$��S�����ja�뇂D�����E�<�)�$܁?�eϓ��\��pP�d������.��̈�f�l�(�Z����k4(�t�\J�O7k�xҺ�]���u,��J��w�M�����ޓ8�����Q�<�+�i���
!Ƿ"�~�L	*n��0�XlxVHYEB     400     180)E{�Ͼ=��}�@�
�"��"�F�L��6nyIZ�>�&�#�-tB��5��������=A$y-����J�M��@���Q�0�<��Xʅ('�e�"w���%1/*��,�ﭒ��A`JB1Ar봐{�M���_�M�4���I���+�M͜S��"��� i	��������%�ˤXi�!ҀN�dm`��}�9aLV@.�&�P�ť���ne�h��Q����Pɲ|�
�� E�M��{�6�=��ҵ	x��.)9�A���Br`��ꡤ�.�<�/ޱ�%��1P�͈�{ir���UY�-Z��aH�Q>��R��:�mF�q�@{�X��$�ƣDi�Uw�R����:� .��h�� 煁7ɐ.'+��~��MXlxVHYEB     400      d0�T�� �Ò�I��!�_W����
�����Y�8���j ��m`׵I�\���B�.��\��*�=[8N�����pⰼ9+��-�7H���7�2ȭ�@����'Q����f�j��R֜����#U�?l�NQ$� ʍXP��K=�����R� 6;� ��e���C�u��զ�u�ǝ#:��g���v^�.���l.E�LYZjN�XlxVHYEB     1d7      c0n3�}K���·���kX��i��v�}T�37V�r�4�V�*��'!���Y+���^/�7���ί�\z���F�Y���l��k!���T���AC��@�?,Ȗ[�L�ѯ��E{e�|3J�������4 T-{sV�Z�ȟ���$�~Ք��!���'�"T�oL�D���0�s�M\-2AX