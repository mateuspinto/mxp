`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
O7UnRw83r4I5hksTfcIXJ3pWGb9RZhBuaIX7cXv0/SErcuaCDyx6twjHBfw9wtKcvccDISaxQI+P
LzcfpFfXnMQkdbpAeZJ7jjRCG2sF7IDKIP45eIRSdWNsJ+anj9WxuOV5TcDhSIjroa570lnV4pgc
sYZjk6sTlCK7MPTJkxCGEaf8BUkLJnGKoQfcB4383Qd6q08BruK245OfcNZR3acCg+8v/OI4dwAx
3pY2U+yh8jIiMszfAgJb8KZUlkvysONdrq3d4TgJDrPi2Qh9UrmHhNivnbiu6r9UGczgb+ypCw/P
F6QoUKM5/Mxty0rirYMHI+0JQ3++0bGzC1/d1Imk6tdqLx/ldq5wCXpERadkY5IN3lZ0Av+sEeNZ
4gHO/rFKpKOWecT63aKrg3nBgowxFwGl9vGtfpIfTj7TrLRQedu61gJ2kliR09hlLkbyZKr8DKBv
ItSSpkSceJVpUf3TnG0vTsBL6c47tB1v/Ru88p+69xnTZfufAFBlo1d3eM0VU1ANKCAzcESlyJQc
vnUmxLbrtla7wo8WTKMl3ttlTyHWn/Zfju6sj9SzTxsYCwSnKDzSxnTQMNsUhI1oF8HAuRqQy2/3
EoIURysJfBnFQEIrux2p5oTrcs4MHHe3r9/xfRUqds4o/WBK/UxFsaR2h7hNeKXg6HHT7BhV+qUe
OHZApSMMM1iYqoANuCBwJ/KxWmONvxlgO6Rk6sUfYEk2t7waTS30oZkPFeVhyCjIK98u4X7btWTr
YdMJfuD8RPQrFoskC6juio1WM2whtx33HU8YnQ1UT7jFjEGxtRGeZQUGZ0QeEm6oXkg0atAkjXKB
Y5unA9/5fPu5bY2nLSuoiRj9Bv/FGbg2fZhzuIwUzocbMfKx2NP1891lH4rPNcR/A2qeKzUmvVYz
Xo5UKl/AfP9lsFC4GTMfR+OGeTRa42lISLqKKmQ6PY0mQudxiUSrD2arbLWEcpC3FfskQds+1IPi
HTa+OKImcT/9QV0Dvv9GqKwe8kyvaR/1dwdvy7QaB0UKe5X97wP/Qpwx5Lc/YItJ2W0tOAzGj9Fu
62kvoIQS2o9m2ChQLCzahcGiZGSREHXYUM6585Ht2Ovc+WGSF1QFV861OhflsxuCBvzzbfKa2wcx
vb1Gqh/ouBz+A4AMjONAwkcxKVuvV47a+R0OutQ+Htd/xP7/FN5rQ89aSFVKwtEAx3sbAWeZzXVj
kGKG4ghHtz0GrPOqrpgiXfPKRyLDTkWVw620Ne1vMgEREPizInAakmiykdxAIl2Np9Ht/ik0y6Dk
rrL1zMOvdE1O9U5VbJLox34p9qgi0WmCDcY4lB5RSLcEKwbpR2rgcP/Gz/p4PEwnTkqQzvbpPqiG
lexA2h8UNsxO2+XKph5EQCfdWQ9ft2WIWbHc4+khB7Br81lo/VZCCCCxGVqboC40wv9BIWDWtgrU
iSdxr/jtcRBFzLg+TUDi5/tVgxb9osUHKoSM8f83g2GWDFf73/lK0pP/Hv/Ae3PZjP72MPW/bf+v
tFaeJdJg/zcW47c3y8n3bjYvozNtNCt0avYCOGEBHo4TT110imkLqA7NN956SNNhflxfYpdAYHNq
1m+80MZ4tHTnu1+yY+Au267KJEYLx9YnZbdOaK1lUCLYHZkB7Pl9l3jovHypJTM13418HBjMKo2w
NqbiynrmaS8MWQgV2U24jjB5zx3enG1Ad1hdacpoOjk47r40jps9Hgf5Z3F/tFD4Bxtteyga1sSX
UHPiV6beivTNPcr/d85E4/dtGSx+B3QIVrHqGGRDjGqGhYHXtIhZ2BX+/GcCB4FqUqSKftZvsW8r
LaA2LsNbsxSXpgpUWqymCqeYrzCdZQeubx78s+MX/wv5i1I9QOS8ubaDpTHE92RwGL7CA8Y+ZCy9
7U3j5VAe8T8NNc6Rv1U2B0GFuNwcvZu30s7H5qlS+8tY/+tpndLLkHa4VSX0/j2yK5zIXvnrrtMp
ioeUNhYA+yMJLwFGmHHDvCPwVInNdY5vqX2tNeIceBSYfp4nFlUOvnMtSmYyZOW5H7bFCpoRH0Dt
8QRazO7MoZDAFNzwn372iIcKlrIUyqO4jrximBliObXLa35fluBMxAUhkjC5Rlri2lC6F2ATufBo
061NZP3G47ISrMyDaBDooxPC92W0iAFl4j/XTV6hZneqI///QIQCw3EPIdLuKiiGTgE7jicYglpj
6BDPc8ltTPYca7TITcaraLP/G9SWaKeNHNlJks60KqOksjv15qOIUOAstw9KODC3fv69xnEdGWAS
LYV8d+5+Sc+GaU2ZY+Q2E/NU5HRy0YGkVGdRqRJw9cXUgawTRXgWMxpD5jyPcZ3APxpFHKRxB9Cc
f8r1tQdj+UjgQyR8JKdSStowxo/OdjuPCxp+uWDtqkZcxapLNIPDX/SFZZWp2Ir0CWeKm4/i+hQi
SUyEcuv4Vom88MJrVfxR9jRaRIL1hW/JsJ37u77yLfJxcHd0pRpzdGWnDVUyhhmXolPKwu0j6qIj
yuedKS4LePnU4TIE2rzGnEbrnf/Q2O+eg+Fodn5qfndkjEQjZ5H4U/utWXuRtRSWkcxUsK68kjfy
P+Pasa7aj7mgHP3M+M0WQZGfXf1eRr8TSJQAFJnPjO68ugnM3fqyOii3izpTRlDh6I3JKhSe/z6/
wCHlzoc2HAti76x7/eayS8nF1Wg7DojnPbOpEIMNf5kfyn7Nnpg7fwfnG1JA0HvoZPD0/Xn22ZOE
9Ur46nl+JWKSwdmr/pIiiiU0mNZ1pufTlHLqEpuSPwWdNIcz/TAIL+jw9EMVk+52Ll11cFNgnfYs
ORVX4kMyAKvJhzjuYnVeyWYOXrBcHJNlY3GlPe9V/cDw1hFJBK/tE3ovUoUWT/OzCaSz
`protect end_protected
