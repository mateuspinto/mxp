��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ДėV�ކ6�>z��3>�\{���Ҕc��z�J�9���
����!3�㌸C
��P��GV9�����0��W��T��=�3}�2��7m�v@�=_�I������\��4='�����E1�b�8�̶���Pn�,`��Q�݃�<�8��>|��K��[+���"3�h����f��Z�2��b��JI�d�m������(N$>��[����ʗ�?���$�.�(fd��j���Ѽ$|f�6�C�:0♗�®̠?�� �4���f^a�'�ԙ�AO-�<�����Ѝg﷧��,m�΀�����NP���x�C��6�]�zkMߺY����t��3�&<=��	j��q�BQ���9�kE��L����KJ����(;��;�����m>Ck�q˴��9X	�y�y�^v�υ�^L���S�}K�~����'Y��I��E�HJ�s�[В�Yp��1NL�lx��F]̃�?<�t'E�f)� D�X!����rX��D3�X[���`7�^�KG�~ �cp����;onOr�Ɔ���e{���:��r-�R����p(��,`���2�K!q��`,;ٖ<rQsӁ0]���e��b'���H�]8K�"�ˍy�@�7��,?un{{�k�}�˰zo�0�����n��V8*N�-��hL1gintA<�o��1�����K�ʷzEQ���c7��V�r�2���3X& +����xk��5S�/�=Oa�;�����
��%C��_�	|2���P���^����
e�ɞUj������C?����$�|H��A�0����o�@�Ra$�Շ�?�ؿ_�"�v8�?%�w(U����ʕ1^˔T�1�s_R��k��+b���H�y���r��p��}�T�Ie�M��H�p[w{�p�C��4O�͑�v�@\�\\��:ָ	����±���I�)�[�<~�O �H�_�&�i�����a��_�#�29���u��[����uW�<o���V�>�����_������S}��g����.L��M�����9��s�k��}��HR�[�a�� 
*��rr�a���tn8��((�D�_pF�J���
��C*��:�:]�N�NS�� ��󢼧ل��<��p�����c�<�t~Z��m�'�y,�+Z�)�f��<�qքS����܅���{	G��-�����`���e��?u��l/�;���Q6��UɊ��Fz�f����v�E�~N���F}���y�1l�L���i�'i2�bP�`i���e��L����%!c�T�I&��--C�&`c�n��s6�%��g�Ó����SB���Z�)�n-}馁�-��pwj���5��h|�a��]�~����Qp��
����^�h3��76PS�awY����;M�ح{�{D��F���CU�U���)0k<33s�"4�Y%�xTfbA��|��Ƒ(���ȖM⤟w#O�W���|�^�lmi��u���p} �m �i��j6Qث��1*� ?��
�:�����1�<5u}���6�6g	ٽq�l��o�-�I�(�`����&���?[�":ȁ(��)����]��5�ȿ��E�y�B,T����,�<L1#���7r�+��J����R�����[����FF�ld�/�;o�{���K�KK#e2����G����4�ެ��	�W�P4?Q����1��Q�j ��t�̎�{K��@u�!!�	,��ﱧ���{���<�p1����B�cV|��[�E�������7�V��y�PZ�k���E�Ӌ܉,e�G�b>�{B�D��*����`k���v�o��8^��Z^�xN4f�Ū���"%ݝU����Qx��\,��(s���B=��U�YO���{퀷����؄��	M؉�����B2����s��}�nt��p'�{�� ���q���?�:�js=4�����
��a�!�EN�1Y�=�d4^ٺˏ&��5�8��cV����^��E'���=�Br�C!���d�ϱ��Y�CR�W�>��,�
H�(���#X��@��Ypk�y�o�d~	FH�\��c���y�|���w~,����ν[��fZBJ�tJ�G��Z*�I��5*1K&�Hz�?��p����B.���mD�Hv���h�@��Q�k3��n"����'}f���q7r�5�y��!�ϗ�S��T0"�;4a���/o���'����׫��}B�V;�
��|��-���˔�n}�j���K��t��t�;�����'�m�|��N$��x��Z0�>��㑅�Y��0�� ՞������z�#3s�~��E ��\c,��:���\�󖯱k���n;:4�T}�o��W��l�t���ʧ ��㿏�2Mɾ���kT�:kɩ|���D��aHZ�]��{��R,��'s���ɣƸ�e��������?��3�T/�3��s;ͯ�M��� k��W*����\{���~F�#�� 
'��/�¨��V݇T7��B0 �;<�m#0w�5�.C��/HX|k�X����C�����"Lb0�`��`}���t�jٚ0�������a�U�x��g�.�|��εLSd���&a�=�3��8�ӏ���9�9s�n���+�>?/�*�>�k�.��B7��w=���b'x�Zݾ�}Z� S���W��h�I|�|��$��@L���ŘD��U��3/��ۜ'T����UB`f�@�
���~$$�No�3�ݘ���YW[��2�ar����u]@�,���F�(��J���^�T�&��S�Z�G�_�*"��q��{���)�L�*rԤL�=����E�|n���o�Ş��6���G<�xl�Ak߿C!&g�d����E��d�%���O�a�S�(F;̅Bnv���S�8U~��Q)�  � /�mI�k�z>����a�l��$���O<��eĿ��������+Biio��ݪmx�7z�7/���N7�&`�5'��	�BT��[�Sd��"��a�8؁��T���:�C�1��:P?N���0�^#�Oe��h��xN���6�C���d2����ڀ]@�#T��o��R�t��l:���"�<c��%�bq�}�5�h���g�r���y�C��?����S4y�\���;Qӗ�W�c8�r�>/-�@�f�f�ā�N��uC�*Y���}6�w��8)�0

݁�UHL��XoL7�ƹ����n�m��_tÈ=�0�,�$�I���Ю�, _���6N���.$Ӄ�j�$����'��cQl�C��@�_t)�rkr��p���#��8b:h��������9��:dRU̐$��K�qQ�	"O/��3�?K���m�A��ʁ�B]ґ����q�������&�`Ef��D0�#N�*�:�#F�-���uܔ����u	>�:[#��������KB�D��
���XbZi}}`�
���1Q��| eJ9.Qr#N1�w�k��◷M pv�ے��p��KӍ:n�3�g��I��=pDIF� �C�Ƀ2:?"ْ�� ^$"���	ㆨ��%�ߠ��32�>>���&ۼ�5��ojc�k���& �W��r��?	����ǒp.u�g��s������ċx���Ϫ���m`�~��uD��ɟ��i�l�$��+A�Rb��O�)s���0X�l�� �G��A�ĩ?�~�e`�V��f��8�|"ދ��@�X&G�q`� �+}�"��#���CS�;�:�a����y�[����5�#��&�L{��Gau��}	��`�Q8ɗV<�H��˗R�tG ����3�.��]	~�6pE'���:6A�[�Y;����-��ܥ�V�g���7�%B��Ԃ�^!N��\������%���]�����"��NF�̢8�3��L��T��fI,Z�Ǳ�)3�������nB��{v�:���y��SYb�M�?C8�D��1�jЙ\�mqB�+#������g���{�T
�/���K�TE����wg�p
+�6���M܎����I�,뢸����{/W���@�C��t�Tź"��(~��q��E�n���Ԙ���������{���Hz���tʓ�7����G��u'�������P�]�i/�`a�@$��I�S���I*��A�+�&��P;)�Z �k�0�%_���:�u �t�x��Z�~w�xK�ƋJ��Jv8�e"+S���f��l�J����fd]�y�=u���=T���&��X��"�n5V�7��n�����I�f�H���h ��oE��VP��㰞�������y����W'�	p3��.
��R���r���"p����@)B�o��]v����Azh�^p�&BثK^8������(�|v�1�8�E*2��B��u�^����/x ǲioN�X�afС�6CIHY�֚�e���O`|F�j�ܒ�)�H�A�����B؈���Dpm_����rc�V��j�L8l�X��x �~VJ�N�n�Y]�|o��(����XT��}��N4��uf��ЁT���UC��XH�m殷A^�k`~�kD�U2��wK̴�돢 �Un���3pz1mLTr�z��5�i��1�׬h��i[0|�X��Ø
�����ͨ�GA�c���ҁA,l�	+\
��wgd�-�5����pj�A6X����&��l���c�	��4�/�#锔;9ˇLm>�}�/6Ѧ-��ig�� ̄�s�^�Ig�y���e�:��y��O팅��.��#���Ml��8g��#�ffM�:M�ѹZmmOF�< J��'O۶���h��m��d����j#6��R�\���ۊu=�F���^iV��L�3Z�Eh�&I��d�À��߀%�|��`T{�T_�HH����㛥Kc���(vb`e��� ���Vܗ�/�'ٝ����C&td%ō���i�����p�,;�-:��������[�q�=�H��#MR8��>t}"d���M��<.\���]���^4�v`%�|ޫ6�	��3��Ox~2[X_�\�V�|I�E�z�b� -jU� F�>/�NzIz����51�a�&�n��	� ��H�V��N5���	D�D�������IZ�K�)���������r.���������ra����'0U�k+ʉ$M�T����\Z�;�Ѩ���i�~_,�DS�K�������IЄD{��k���[�ĘB[�V�IHeAl��q�q�Ĕ�9CI�H`u�Qd[�/L���4�)<��1�U���*+0��jN����ِ_x�f�������g�ڇ
�tI�EB��.���n8֪�eF��U���8�eq��
�XE��8�����B��gT�K�y�b�1��G��^L/��l��z�3�E����]���DH���b�%�TM1ܣYW-Fx.��ھn�`5O�<�[��
��Jom,�*2ky��P:�1��>8'��&����k��㛧�1>�S�)�=W^�n�����o�I`Lv��Du7YGQ�vs]N�;���Ά��d�P��v���B3�BK��|����D�j.�60--ɬ�'_���պt{���i���� &�8A���Y	�����T��RE�O<��z�s��l����m���T+gV�_�J!����R���L���gB�� K��=��������hA:�Mh�;���[���� ���6��?�,-\�A����&�s����	��vA����ȩ3�7f���0���^V>EP���@|>�)�}K�hM�`R�O�3o��9��F�J����@j��t�,�e��͸'��Q�������'�U���n1�z1�;�N~�F��1�>4�S�v�C�"�����z��c8lmL{r3�ߴ��bҥ=�͘ 1Fg
���T�rr�[�O �v����I~� ɱ�?�j^����6�dv"�v�A��Lǟ["����7����,Yx�c��ލ wǘ�/� 9K�����7�7�Q��FD��I��9[!ʛ� �r���'�#`��۲���A�=)J��/��ޱ���v�c{빱\���%$5�a��U�W	9�8�fe�	�$�_�X��I����^�lHV��.J&�׊>��g�@�8���QN65��O�3�4!Lp��C��˟�+{q�4�pIy#�ڛhz}����}f��+�;�h�=�A`m�q��Փ�3tG�|'��\n? ��̸3s�i�* a��Ɂ��{���N�J>�Qŕ�E)���O������T����5�o�=C�^A �G	Q;0|,���ssGm6^np*��a�C��̩�J�_S!���4���H�a�99Q�xE�xo��T �5�Ab����@�������EJ����e�~�H��@hڧ�?��t��w��>�|c���R�E�rXR�o>�YZ�qoi��}�h:"�a���؝g8���[��/�X�����J�e��R�����J;"K^+��о.��pF6����D������sغ���Sw�s	��&G&cb6��O���B;j�������T�vv���N�׊h��!���w�BJ�^jQ( *}����qx����;T�ꁅ���#Eoj �%���Az=��Wx��e��S�`nP�s�X5����,H\5f��'6┙��U\�el�>ML{�gc�#�� :�E��c���	���U�Z4b��:���Er���zbx�*�xT�b�l�Gf����D���V[��E쐹��IR������/�I7e�N֜���*��d7�i�X�
ƈ8?y�h�h�)�g&t4��Dk����NA���%�2����
Z*��A�Ԩ��v�9�?H�h�ϒ`�3*N�b�q�G�$[�2Q8s�Է�gC�%\v����T%�t�E?΍?���S\�Y�d݊
0Q�b�[ӽ�O��Y0����|x-Ay���D�l.ޠJ�0Da��ѫ��.���&/Z� � =����_u�,�~���w�擅U S���]��gf93m�-S�̉N�s͊�p��#m�t�_��w�@�43�w��>��ɺT+�7����*�;Ͻ���u$�VznƐѯ }�v/Z(!�5�%�4��	�W�5�y�wW{���o��-f8����B�+eDg9�w������?�C��6)�փ�w��q�2�Z�ݡ� �Sq��cb�6�2����d�����"m�Sl*?����������}Zw�����9���xS�2�6�9 ������G�_��26�%�s2F��ko�'�um쭰�XX�v�f��n����.�5��p�F�M�5�#���C�d>����G-��)݃��2��V/�A�;i�r���Ҧ����y��s5-UnfU�L��Ч~H.ǒ�4�Fw�OZ]�*��Q��/qT�+7������G
|����<$|/.(��7>:6nz��V��9�4=�Y�w%#���u]��3��}���+�4v�Y�n(�2#n��S!��|���5dM2���G�Z�kٰ�HbRD��v:����y����ؠ�g����J��~��x��`#J�W�1L#f��:m�,��|���s]��ä�k�;$��&rF!n�O��kp|\Nר=�,���P��tc�8��su��yvG{�"�>�j��:<܁���-����T�_�e	2����WS�q��0�N.)�c�,>,�:�̛<�v%�%�v\�"�V萁G���٩��S>���j.��U�yO�[A�pe�y8�Wcg��7�k���y��@�B)���d����tΏ��a+��i�� 2��ˁ���Ms�&���_<Th�8��5�����4�@�B�u�3J�Ҙrd�w!����f�h{�ߎ�	dE�Z�\��?]~_U�w������o�,�@I�^hR�s��-^�e
{7���L�'�W�4�]���Z8���S��n(���(�e� =�l���z���:@8)������؊c�5��\2��+y�)#�6���rˉR}�����J* ����=�_�&���;:=��x��¯ǥ�_������M�{/�׶�=jS�#'��d��3�[�L߲�5s�@��a�#�����P��!$���l
8��� `ݍq7��!x����\���Dʼ㐧��ID,��V;7t�:\6��m~�����,��i�!�ۏ�}�:��v�6��q�h���!��9�+X?@��1�#*n~�`� ������;M���N��/=���ΔYQ���� ~��dh#oR�7
Ŕɋ��ʈ���L��ҡ�m�����? ��24h�	��)�߳��=�9
Y�	�/*UuqeX����f�����'[�5��ժ�P<~�n�Ak~}dq:�&94��>g9�h~,}���:�%�w�g>k�\Y��\e��}�q�Y���Sɑ
���M�[D�l�>�ל=�ڤ$�]v�B�5�i��y�΃�5�k��d��n��p�~̕��C��3,ߌ蓓|m�87_��.�Zc�u�4��U��!�3�4�}[��aK�4c�+
�C���q.��=�>�W��l���@��Р
|]@�Vz��ҏ똄�2E�]KDO��ʝ��C{G���>����)R+�uݶ�	�����",�*�%��B�u%>���4�HD[?�����:k�,����՜����5�7w��E&4�]�v}�q��Kwj���!G(V�M��{��lM�N^~pjBo�H��T
d)��{QL�N�[=^l���⩣�i.6�����v,���@Pc��9�vR;u-��+�yS�AR9�i�Ȃ~�5F:�ÉϿ�C��^E���Eq�}��#:¦�,�*�m��&��H�U���EbڶD�p5s���ˆ�k�-��	��9Nh�\8�f9�E�P������ �g�׌.Q�Ҥ���.�G��'*������3G��sO�F	�<��t��_1�I���>��~Q-/�>���0~@�P���PQ����t~<)n=Y���y�V��u�K�if��/��X���ip���Znu��d�$�z|� �����Kq5����C9ғAU���fK<].�l��ښz�̡�W����}BPW%�Tz���6{С�<(��&����z�)����(�#B���+�/U����='��Ƌ�r���p����C� � �.	z�h�����*�۩���U�O4���ⴧ�Z/"PO�f�>8�j���4��v�*�������]�V��;|(1�>zj� ������5Tq��!S%K��IAlL�dv�遼0��vS�m�|"��.�f���}�bf4�p¤����f���)�V^km�V�MY��PW�G�7x�{��?�Ұ�P���`��u%K��u��g8�]>�х���L�x_1�T��/���}G#��o���� ��E  ���� ���8��#��q�.H����G���'D��y�uX�PYb�L��R���56s�bdϑ��
/�O�Ё�?뎂��ۛD�@��$��=����G�Z�)0ι~�aꗿ���Z�͏��f2����Y���L����E_�A��������	�R�L g�%�@���@D�9�(B�I��6v�c>��@Z�N�[�?����7Z��n����~��(~�yw�f�[��c��+7���((ʚ.���$!e�G��	 �ǜ�, D�<��,�������.��nXco�nB4�kZ���0*h庼�ndm0܋o�2�%F��!y(�
�3��_g���>���<���j�
W�?�������.XM���;, <q�yg����