XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;W�����MN)!������@��,�x6Ws�A�]�a<��7�y)����C�8��'�5��!�9Lq L���d�AYx��3��a��Y�͞G&�U=k��O�\8m��B'ψg�O3�	=������5?ٝߤ��pkNw�,��,[����X�3���sy�� �ep:�;�i�+i��_��:!"!;�'�&T/u�p��>�}/z{J�v}ҝ�.p(�$x�n܉��R�e��>Wx:)���Z]�����v[�
��r�G��N�ר�az�]1р	H�vN
�",
���T�V���;��$ڬ;ٹ�'�k2T�4��[�]a����)�V�7�A)a�/E�"g�b�'����` �M���xi�%�L@"�d�w8��1c�������C��!�Q���.������6�8QjԒuoy�6$��n=6�\�AŇ�46�tK���H��S�iZ�uaQ<h� ���;g�؛��8w��37|�_��Nϴ����#]�Wj�$F��Sk�ܔ瞠<�� D/��� �HRl�:���o@�2��_�MX�e�by����E�c}��n
�!�>���F��"	M��l|6�}�|�E-�@-|L/�^�9���A'��V�Ye,v$�l����MS�6]��������"s7���R��O���T��<ݚ��m�1��I/7rf��a�R��ĕ�f�]���:��U��e�=�``ێo���w�,4��+���w11���L )���[�x�᪾��9NT�XlxVHYEB     400     1c0H�*�άAV*�����)�7��V�V���,֋��� ����5U��,��f�e�'�yx#���ǆ��E��,Q�o���A� ���ݗ��NE���Fh{�Z�T�)kT����[�[MęB��[#�]Q�}Q��?ZGI�&	�(��(A}]X�.�J�Q̕�߰�.�o��5�����h%��V��<�	��NS��-\�Hbɾ�S���a0<h�����f���F�lG�R4#0��^.�p�43�Iv79S�t� �V�p��%��4E���=~U��� �1��3��� � �|d �=�$�kL��.��s>yk�S���;\G�8%6c�5_�Ǐ^j�/�ؗ���%��owj�� q>DK��L�ZFȨ�;!g�ƚ�f����)�TC�}�dr(�=BFK����f!�#f~�-�&k���w�g���]'�`�ۖP���+㡪�XlxVHYEB     400     150��h��%��q����qQ9���g�L�'y���E���5W]Bkj�`��9�����RR��������KԲ?U_X� �˚��ৱ�:.�t���zyZ>N�v�\]�T6��o__�3����jy3^��G��Uiw�)��pv�"���<f����������$	{w�S!w�OVƨK�O�֤���I�>�٫�<$w$�X�D+��&�z��2ʮ7��Z9q��D���7�� #N��4��r��3�	
~�*��<���/��WҶ�k��]��R7yb��H�0@0�dy�_��"F������DpJS+��zޛc0�"y�8�̶XlxVHYEB     400     130�1���\K��N~Jٲ�9]�}̯[��^	��r�����Ϻ�F<<*��~���_��[�ٯ�f�¯��%sì������� ��K��G��V^��A�5?�V\���^Mg �|�U��G���kx^�g�v	.>*�7��<�\2���-���@4������$7G�wDf����V �M\�����8��!�-�y��� Y��5�t���jG��G��{1>�����u'���<	���'�?�:�rD�{Kq^TU� ��d�B]�W�0|�p��CU=�\݅6�T!�p�i i��XlxVHYEB     400     160͓)+�qS�낁��b4��ƚ%KaÒ��z�h���`O��U_ʞ�ci6I|�Ci���M�	�O�,��M.�<�����멍���Ӻ���7��'ȶ-�r���r��,��`�>������O;�f���6��]JVPFƴ�:Ըˮ!6����
Q�H� e��麛��Gwa����n�23����1���˿r��n[����dj*�"�a���-]�(����׹=�4f�}�T�r9��{��Y�c׽�������P�M��4H!�n�t�zy��#��Gv�<N	����|���^"�j�"5ulg&�}���VX��3��c񫸃F�[SDVқ�U�k��XlxVHYEB     400     1e0�N�'�%�l>4����-1+]&��s�wc����;4|?e<g�Y��S��wRt���q�M~�sJ�����m���G|��������(�M����+#*_M�9;L��б5m�$�`�O�����f�4�B@3�aN8��"
d��1	Bt!	�5�����J?Fl���q��rs���T}�~!�!��zиy���I��%�u���ی>}Hl��pDF�t����
ϕĲB�y������h�h[\"��ӵǔz�N�%�jlZm�:P���c��8���3�k&�߰;�-��ٔ5f&a�!�����!+�mL"r��y���"Q���c�&Eo[��dyh�!�9����µ��5(��@Ӟ#x����e=C�7�uS�<⨣v)��JV_��x�C����M�h���^b��O\Y���-5q>n�ZC�ĎVsz�1'�I-"��g��H$��=��Z���fXlxVHYEB     400      f0�k �W!
���4������۔5��iz��3Q� [_���0+4G�ݾr�9��'+�[�NM�d&q��x�(�`�!�|�>���K����)���4x��0��h�����h�0���;���8��R�yչBw�_�I�=���W
:h!�~���M�Hl(4�,e��l�~E�Q�W���y�G��D�'�R Q��2Ń6�v]����{s_,�9��tL��� �Z���XlxVHYEB     400     150��q�,'@3,�n*zr�v��i:��N<�4�z��J��M����7
Ex)b��������(��@+R9��I~$�����1?�iV>��aM����e@�=���*�)\PC/����㳥�'m�Z���w�?�8��e�~�!���TՃ��;�G�Hk������r	b��V���-�)����2�Q<�B-��Ľ�41�QѴ&"��j�~I^�uE��$΀p���U���g�1�XT��(�+IA2��r'��68��!GwP�U���KMqI�k�K�_�����{�O�y`@J�}YD�Pҁ+*���J-I��CG& ����x %r�s;��K1u����xtXlxVHYEB     400     170"����/(���H����S��ęB�
v�':wƼIX�s�z�����q�O\j7�z�>`��0�Ȱ�p$�-<�{i�
��s�u�g5kJH�f�C�ALQX3^mQj�}U{�@���&P��C������Gol)�EU::ؿ���#��l�DR���v�=�.�iN'��V�bU.�m]�<�W��0�_~�X<��������,;���� �&��ݬr��0G΅���8���}�rc���M��Lӝ:&��.��߃�3��95u���#h�M��@��
!��
��>��Lf�����,��S��J�@��"x@��M'z��k��p�A��_u��f���g6f�A�f �XlxVHYEB     400     160d�����y�@(�j!����m��ct��4��΀ �V�说���܋T�q��S8���m'�>��J*E#a��O-�\�"\k}�|Y�s�?^���ݪc�y|���H��޹Z��,�b���u[,�L�A�H�~���E�)'�*hd��ĥY򐴕��n���	!�O���~�{���.�U��f8́&7*��Ⓙ�=�Ze|LIʊ%z��nt)��LɃ6,fN�}|?�G�r�E�QaˊSYZg�Įh�qUi,C��{aѲ�MoS~��0E�� �w��[^^�7��b#ӎ��Bz����F6��&�C-�H������dsy����w+XZ�YC�!- f7S#9��̡?8�XlxVHYEB     400     180�����5^H� H����#g��*.*.}�1iӻ�Xg�2�9H��8�;�p��@��������p�AsH�,�h�2�p�",��������4�H0����1>�o?߼��B
86l�gp�
u&IY�$І���X�
`Jˮf�Z�-� �n��q���^N�]��7/
à_�?5�`	�!Y��ry��L�ɝk:��\��U�w�dum���	a81E�p5��<5��Y`_�y������	��j��N���}nzR��R)���M�l�^���`W&NIi ZQgp�n�Z[�p�_�s$sG��A\3ҳ���(�~0���rDf+���v�pp0x��W Q�$�`
ҵvu��*�i���uv���`����3PXlxVHYEB     369     180#�i���������G�E��2���G߭�Rx1R�  0
⟿�44��*��(��R�9`���P��N/f���#5wV�����r��ݻeTC����i$y.��o͉���-���.]7uʵw<�R�t�t���9�߇��J�����c��T�L��}�ԥ�	�&g�MZ�/��j��S���tw�"`�����[�������a�`�;����$]ĂL���^� �R�6���ʴ8�q{Ü�uL�ssm�0�/,�2�0-#�D�pC]�d|��\B��~vJa��;�΢x�PЁ~Tɷ r#��}+�{�P�-��ğ)�ϼ�������96�l�l�
�8Ǥ�X4���9��lv��s���Ș�#