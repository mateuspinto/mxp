XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}D�Q��}��+FYF:���:�a4�E� X�n6��*��"�O8�7��>\�r��S�v��6��t����2Qf��;��E=Q"�6��#�md�� ����V���s�,T��L)��bV޿�R�%Șm�k<���Dr��fy:1�5R�������o�(fuf4�:�zB�� ����t0���Z�^�����$+�1�hm3��.�w$4hZ�^�t���rۗ�Y�Fh=X����r�3�R^r�^T;Յa�	%�0aSkX��M��Y;��(Zmd���� �m�$�{�,:�t�d�K��;���uز[ڔ�Ҳ.�޸2^W���܆���:0����R����K��
n�؅��Xkq˹�]U{��Ȼ�,#�Y�����m�����`����!_u�X���g(�p�E�{�A�r]�+S�(lvb��� ��vkņJA;>Y�N�$^�IK�:W�JRt�����ٖ͜�B�6���#7M��J���%�ߊP�k��"~�BN���怵ʝ�P&U���`������H1����`>�7pk��K����h��~�;���3��YX;�o��F/� ݘgO����a�Pt<���J��7�tHԅ�l��$��3z�i�&j���Rv�lwul�,���d6ОuO^��T�D3�<Y��\�'�y	DJŹ��}��q�Z��q")���4A<g��M��ÔnBQ[�k�ὅ�j�x��G!3U�
�~�*)�4Zܽ�R1�9��s9XlxVHYEB     400     190�3��U$n{r\���,W��Ğ�L	G؎+�M��@߽��E�|b6%�$t5�
��t�q���m���Լ��hQ�Z�g�		ڋ,�jqw��ֿ@	%~H�Jt�sY25�;VK��m�k��䂆r	b�BwZ�Ԛͽ�o�����e�#p�2Ѵ{�� <x��4�$rH7� 'oHYu[f)��	����	��o�v���X�d��k���?:{_6����]��	�nk�@�NR��	΀�ѬZ�&/���z��1�r!~4�S�W��n�r��*�B�-������mr��~�{���h.�~���� �� !ｓ�@|�������'t��b�\�޾���>y����t������5����1�����:�XlxVHYEB     400     140b�F[���y}�E�\G�Ȓ�d(<:I<S��[|lg�|�]ӣ҈Q���|�_����T������s��������->g���+���&�^����<��k��d�9��eGҠ��q�e�1�Us�#CX`�YM�<6V�͆#�b,.�؛�]O�Ο�3
�z�~�� ����ב���ʳ����.Z׆��N���	PO(ͮ\c�c�P��Ĺ��@8.��}zJ�죗�%9O̭nX�LR( ���utXD6(\�ڊa|�f ��ŭ�ڸ4�w!Ѡe����K�%�S��c �Bv���B���f%�l�ɹxXlxVHYEB     400     130x1����~��R�'��؟?`�Jr:��xJ�nx���ybv<�^�|k@*$H�+�/��@�WIf�4�k������Y�»sv[�m�R�����rۀ�14VR���,��3�1�����l��#j������"��v�B?b�e�K:��eq��,<0(*���@2_��`����=���ң9iZҦv�C��9�2�ت!�ܔ��*�&V/��S�����D����镣nzw��f�]���=����06T�/!��y��5�~����&�2��J��g�t�ۍe��"��C��t�}z�&�?���XlxVHYEB     232     110׉��_ས�>��1s�\F�͘mݩ
���=��$�L~GbR��; :�
�@�L���=���A�Ϯ������v8�a�&�ަ'=���Q�D	��2�$4��T���gCg�@�1 �}���L��J�Z���E�u`L��M<8�Z���X�PQ�'t��M$Ǟ��v�6(�Y�7�L+S}@3Y�k6���BT���v�7��z���cֻNtv��x�M������!u׋��tI�$�)t���A���~�7>�D(���.���2z���