`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
Px7LmfEj4vpQLo9J882BfBgRRRPXo8q5Tr5D9jy+JkkbxYr/KYunpI3FylpcYm4fcn6Rd4w8l5us
Ebeb43EPUZoX5w/MqirXr5EFhPTvtd41f5NTNbIHy0Hk2MaFaNX24MsoF+rVm9hoJuB6tCM4Zdtu
m+PXVci++g8YoZW6uCTAxuVQ/NaHZJ0QtFP4vx09GOEQ2FRLIKhd9FGyiAHg8DkAtBjmOZihqzW+
xeBW+VBw6poq4b0/U/gArJjb28uIfdXWQfY+f/m4WadqLcArD1CnfybtFe4oxTi2fYqss4DLHAgY
OkQuIxYNL++Rw1CGE2YKjq9enFQgcLTHAFSKN0malB7CLIiuMELjPCXXAwa+nRsYZP7PR3QGmMCO
wu0VxKkjg5BtwAOP5ElHIu0Xiph9UYqFkk3aHFJY1H6VesCwgKb0G+WIv7UOTwjBzmjV4cK51mf/
XQo19Imdc32DGlBWMvH0J2nd/99us7HSsG3TAdhGGnGawES6hMIzDFgxIRd/1l0957puAF3/2emd
0x6RiQoUuIJZw7ESm4cfM49b5AW3iDG+xfvCQ4hFBYV8srw2EEfxOx5w4KikUz36wvA1omyr19g+
/m5B+cdvfJvTNN8j+/9QAg+1ubMc+XditcjIuVqXHP2IEZ1NFvtWtVIflXPNGLa9xkqvYHBAsGPj
TL5W4q0XPImtcV+bql1A6LBs+5sjqtxgwFWmc9bx2R2QVMxueGI2gpB/lWJ5nOdsDxnYhWSv9Gda
uoKrrmCT0MaYXbQhG0vo2qPryCzXbOFigK54eXlVFV3sWF9l/gPFoeVL2yt8HAZ84AVmrqjMHbSt
UCwmWSI4MK1S1IBPeULfZyrQVGmOhR1LJ3gki7ME7c4kaAqVugjvwcFWhnw7CsuDky5o2kqYGKK6
TK0xomIVXYs2lASlnfjdVSRvaYCwrXmHhtzE+pZApLWgpI5vRxD93jixLCu3+Fagy5P2jM6cCybE
8YSh65aqARmqIrJLe4W0mKD+IBsutH+o8FYSSo73IuZiT67v0PIeDHJ2MAgegbRKoRu/fLEgBT6y
LCzlID+qbkk1nFSz8FfD8wM+EJLn0qct7zyoJndsSPt9RR1jtq1CeP0WITMrKzb6XM2H0mc9E3X5
D3OkUouWu+vfraWY2CBV4EMKoNheKz+/J/bE3CJ6LaXUxGByfO6U0dGZXNLBsCPZCTN1b7EzrkIp
FmcAQTeMdo5GHqHuK17t27WEEuLxTlrDGhupT3rRghqQh2a/fQd0xLZQmExp/lreLTMqlAt8aNDj
Uj//hljd2cEke8TvG1KYx/S5V+vtFlb9m5BaEuBik1K+DlA3sp3W9Qgfi3/RRc/iAoXe/5FmmhtB
a+tkXksILGmFV+UU9b11G3E2fr0e8A6/+NZgtLzg6SnwA4e9Wha79A0e32+m+UdT6K2nBF0o5IO4
kuKnqkYMvBlIh1zXzODPxXEdFhwwxpUwovgX/Icf0JC1pnGdwlsuSHIQWvzuvuND/0z1kKW3QtE6
WoPrSSzhuC4ef0ltqQaLHomOgT2edDQdB6l3fPrMA0ZRjbr3d6O2gaDLO4mCgcpUJOtuMdiJH5im
8qkHGQOkajmEhDQ1cnu9ZX7+/jlibIAUoec+UPofZmUQmGS0b4eb0C37ntXhvknrLB+yCygvOy0q
/anfbUl9Yv6hSqDyfShpGLxA5ZPoliYwIZ7fCiYmaGz0SXz4mbmuPS97qcYXA3jiFJep1sry6OP8
6Q0w9MyHXMbtVIuvdaiGcezTdmCvo2NmxG2CiigdlhPDTxrmMX46E6BC4LrZMFRsD4Boec10znfR
SiCeQ9SB6CkZM2bXtrhKt6zuObg/syxazDjCRu4MjOfDFimr8vrbiNYUxAEvIRtUCYi5DJCybQiG
2IuJnhehVFh5ZX9oW9XgiXOVk70MdVIyG0kuJQ7IykWux8Xo1LlkOanJP1VvVyIbe0kG7UwVUXyw
Iiz63M3zKZjXxEAochYlyTRdRZacj1ZN/M1Hd8j7P/bZKrdHopxf/b1fx6X0j5YoVWbGKTHvLSmx
hetzdN5XaIY/lIJfjUrKLrLno4OYXjvTzhyfhVPtTCOdO3+niN0VzY7gDWvu9IO41loNvlsRCshE
5kewKuGGuFxfqgkxsDTdIs/8caxk6E5QCJkuBpXx0WUHjD4Z8UI5sGgPGnm9Vb8H+3sI2/cVGyYz
488zjkRQ3td/R+UwNK85byTYQQi9UvkOO/qqghmHx4yUbqiFbqN5YB2AycTnqTiP0U8KgAMKmxo2
DXA3maCfFiDiOcsDewI/Lz4FSR2JRT1m4IiB56AXT2Sg+1vZhg+ESY5offFpQqpB5J1luYWpseYD
G4+sTDOIOQcppo1oTGa923scAA8F2pnAqF8CpL9gyJYakupae/ddsWAFkjAy6Jv4ysoOT69mzg+4
JK94Qc75LwapRi567Uj1Cozt8ncsMnyvUwjNqTJrdcnOHvDJdJjdfNY6x4Koyn536GIYZVCe07DY
yv/VzcpcBKdD/AH9tFIRJ126F4dF57p0CjQNk3RfkuHHP9hh4aiPT3amQDaNcXGrgsXbuRJg8SIR
94z4Kxs9+Bbaf9dqGjNahQhdKKyrqn6sUBzQdyUcpBjmSFV1Eug6kLaZ+/Spke4fVboqJZoYvs61
5lIY/mhycgf3dqN4ia9gmVQH+PfhkLaUxhiRHO+vkhZ2FuhuzF90MRFhDL+ER7uv9/6IIRkD1yLr
TGweaMR/IWbPFJh+uPMXqFJmVWWUEAkAK7rGdmRSBnxN8CH/dugbcu7kH+ebzeggnIe8rfRC+BnD
zPyNE/X6yMdh51QJ8gzmOTxplAR2+V6VJia7+8TVnbEhEr2hgVEvltOJ7ieI04x7C6VPfZkFg9jR
yaidJnWPhDVOxfH8wHlOdv//xKfktLgUohwxj9QWW9Bgmdm/ZVraEQcj+adIJBR5+WLraEnlZ43w
xWJf7caWptyJGkjrg75ORvu9DnwGz7HQt0C9uvrkaHQZYyLFBxz+WsIyqDTqK1SkRQ9SHwL7wO8J
UB39H/ms5SWxgnAeSbWU1VzvjyuyUX1FvzV4YvPPXFD6SkJjGQ36KQ+1ACfxxN7wVzslX5l7DwFE
w+Fs38jcpMy4JvGcLRwmgX4/t6CAKF8Y9DA5RunytKl/Lgb0p0vOkGR3rKMvMGIgINpjHW7X5e1C
tJmyA0Z8i2sH+2FwfaZMbzzcwBxi13MOoNRzadYiZ135qgdU5+6DmSSudkqy0wJel+/l875U
`protect end_protected
