`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
9sLZ08b8SdqFSwRv1zIdZH7uNtfh9m7B1Ci1uusCPX2QVGsSpCwi3gPJ9BTsxmULnmBC85QSCQwh
gVWq4I3Kiny6Ge+j4W2JnXF4vI6o2OF3HVRPvBH3T0fDCCSr6IDeuR3md2HnzymUrXCj5LhCab8n
XR6eAqvzPR2CnW3npHedBEhw1Ct206xuWxwJ52MzkOigSLwqJOPYF8xLKbRpsimYkr6zDxS/0NZO
k91/Vm2Bbz5Xi+TzG+g+GLR8bTbfEp1w33n+XE5dTN9fcP92Flsh/m75Gw6WZyPuU9R81HGOVbK/
hVyhfc4oYzVC+X3V/0pOrfKMTrngcpPJIj+XogAdCJ8UoDQBbwoKNhPO/8ehKUF4li0eKOOFTps7
9pZoZHiNqUGRZy3ZGXePnTMBH96x0CYZNn9l6krhsjgrbx52z8htw77lfpMwPZYYO2l8ulIAIEcy
BAOr6UgsjIvef3KNjLn9HVRq+sJdBEz72xD74E6OndPTRod3gW9cI1xZCR0xRyhAgz4EvwYljSP/
ZLQ9Rw0zj6ddtXKE+vlIdz6WR3iBro7CRdVN+Wt82EUNHva+2fyG+y3Hjadx46OnSwpWjQho5Ll3
NQ5G3BPzmaZ8ZwdgcaCeb0zXB2PNgv1B1FjoIGYH9PmVny3JeGAB0BsxlOiMQ1hi4SqYpcus8uJa
PCSQLW861OYhbXAuqcPul+F28m0OxDPN0MEr6Q43tmknvQIty77gVaSICpeYZ49s34WcFaK9/Mvg
7rR0j6kwfz/PjYlanG/iX9K3uDj2x5iNMWVyHZIG7Vu1d+ZzlkMLN1seEBH1F9kcuJV7aiKRYUR7
WFE+Yr0+hrjMU1oiGeHI+Dklgw/vYBp4C6mcTvqxfrzRpBe+/QObdi01+9cls1MfYorJ9Fds+aba
a7In2Z//ywU/+1Q8MNziFzS915KR4wgXfsNfUJEM5LwxAPFTdrOPS7yddxjiyGm22hFmQQPYeDTb
BiMwyTmbfEIYLW09C2C+ZXM92iYL5oCJWeDuS6ckox5YSFB+qh2TyRZdr/qy1x9juHUOY0d5/ETA
VXjOL+s9CwDUR5isi/joSwTiQ+tW28ETll4Nwrp+zu/jlxeboIsgtF3RDjY/D91Fvt/ka4eTizzS
8SbCVi0TuSjIU/VL+bP0JL3/NHirO93mbzBtvy0qxAS8d1NSLUaLsk7TnQmqQyUOe/z7J/wo5JJb
LdTXule5odQGOMxb1xvowYWybKuBw5chGGATUvmLDPbLaWvTbLIJm0gqByPqYr9CjWW+NfmSWmSi
/zDrRR2EHj8zJDd264g1Q1rVLv+lKq7eDoc/0uDA2Smo7H1SS8gqF4WOCe0PWFdlh6XNYW+zaJ58
CKHE1hFKX9LVMs6Qi/Pu/C+RFfGQxxkJsfOtEpsbYkQITdFe78yO3j9MjPzi5Ul5t823dfNKHhQA
O1qZNkt+Mbhdi1sdzENQ2/EjljGOhPmXMCQcDq2uy2iIZBZpF0zFaP9EiWYQB1wLa7RVbKBTGmjU
JDb/qb2S55ZtW7QTlqfAbyW6znMsWLiV+95KGvQfnGd+vN7TXH6hTNDJIr/0cbKlIY0p+sPewhf5
0foQFtrEU05NgE8Kitnbn7yzwJRhEyTiEyHJa/oG2XZuynwmaHGJAjLLiUifZ3ViLIg+TSldnUxm
yrEgaAVtmDE3h48haCue67cccWDHBvGif4/91WrhFQ8tFua1AhcYfAL1zgrF05qVDpTE+NkPShzf
6n2neXzJiKZFm885QXB8fjfrY7XVG81QdbdHh+SMFTIr+vmpl34XF5UtLMkt/Ao4cFRC8k+l2Jn6
whcoaOKcGDs3PBklaQx+k/MenynoBq8cGh2tD43xDskzEubzC3hXHZpFxFAHLKoQXu2TIzCX6sGr
ypk9BHfrmCE1SDs8dMR8JSvI9FDomQe0wOUGB1bpHZWUGXjyCVXeMTtVPe9OK1W/jzVXjYcha8cm
6VZBHYujfrRaBe2IDLhvWpWmYZklSpP6I3fXiImhUON3n9qbeJ9UMw942/RxSq40RNcAAAGea2xU
MMnern7ry8BPDE+nioHrID6NQJ3hrTx7eRNVsV1/YQmR9ShBCuinc4oTevGUFPDHKttIUKIM5B4H
pcbWMeaAAhVRV7fTOaqxBedEuEvgrsNgSMecxpY8lKXYfKewR9/Vevbdq/nt4jPvx2pbToDySeZn
3RiSx7RL/aJ8s/nkntv2OsrvIOzc+r2Mi+9cgYymhX+1ocr0wq1BOAeKXg3j6eVXQZzJQoNvCTVi
CpmHFBRiwgAM1zTlYvwohkDQcoEydxMF/ORkva4VV/esxqDQec/lwmcRFH0E+bAgO5hzdTj9YReH
WhQZkMxVElREimLf2ybnp1jTdreZhvMiAmp+REaKunzKleV2r30Dl3AOOxxuQgaizcpM2O4AxKJi
mOmHcBXqy4fjzWUemdG6sxDRtHne4jMddmmvAb+Bm8NFTVUH5yU3vUvfkzDTmu5r4tLMopZFMB+w
uoTU3GJeq18qgi0GodygxElDnf+Pj/7CvtcNsz2ZTXJFRPKxeQR1BZ0NIAeHxAkDAB+a5n+b3mRy
gYC/Bgu+OYYFzlnh/iJsjcZvDdmXjQPeGiXmqpYocF1ozUx7WIL4OPA5Pc1bjl2Hn8Zulwtgd1yg
XrOCTxmPewoWPafN+GEUcNIH3HGipLTYjgKSYN3ha1Lr82tFGU31tu0G8OToa54+vDP8Ls5JmqAj
Y+MfWdthC+w9UNXbq4So342QCJCJcSauqkWBYz0HHbQ7TPmpg0ugZx7DtjcPrEoFlemOCaTG8G44
VHz3b2NWzeAGRzDhKr7WIYaF+YjMWZZsSJNDbLjuL+QbwuaPkrHReD2qrJ9WVFwgWXKuf+NAUtz+
qFcRzcR5x9g/k7pVg7erf2jwzdXDYCEG9V9veO7HNRiODBegtONHVciJmH3hpzhDCwIlpknVzpRN
kbSdI0YiHAxct2YyHZmiA/r33D99TcwjQ7mqq2RaNjc34GQa+r0CXFYLmCANySDJ0ZmRWQB9b985
jERmPeHpDnVR681NMdQrQ/fXyRPEpyMhNdzixDRmLAmGr9tBstNSdMRT4PRepklZKm8tmkLaM7Rb
5HsLYQCK8GDrc7Kg4b6il6VXCoLtRmyI5xL2AAK+acTZjmLo5sbuFhVqpypGrxjTE9kkGFXYy04W
96QPRvSX7MGQ385AgCTgtWlt8FUbpeYJJzZrUbEl2U2bsfhqgMa4czHgh5M4LpO6+RrtykhIETJZ
rTPiPbiOFYAm8GEEOnhWqibtTVW5/nAPBUN8FcotR58QvaItV5v9zqkoUA5opEGTLuMjQD1vzsGx
MhM2dbYM/ihhnRKf16fWBgTyV4WWAGjsGrh5pR2VpQKFLuv69F8jEKdmsGwq8fQu8QZEkqGBZdiH
E7ymbvrdfLCMRVzWydZMRtFdiQVZURnrXhd035amc0UiuDAIBfMH3lJV7Zhn0v1C8F7KPJhSy2Zi
2E0FrE0U5AiR5aSLJxNIZCsBDY1MUoYfJ+Qqhnm2Iukdp7VmRHfV2f/vvZaLHN7X4uujQS7F279D
YSZgxHXYcODczscMyiw3qzmR+qf75rwdjs2maY/CiCFWeF85eBUXEFxHF1sxNaIObleSGhPm5Lhd
6s1QDpePvCtT1fk4On4xFuptaq1ZCpRpMKzFqJGg8SMGTF9U3g7+KsQ9TwM9cN2yDF8ZUMxK4on7
loIgrxAxUmDAtj8R3dWXGCGfwY8tfiHK6zAOlsR0VQwSiHlMyOKbSug/Boq+i//K4c4rMlpTHcdR
ZRiwUicndPSB4hmvMi9ZYr6t1Dqmr/e6Z7fBvOszGvS2UUYiwLuGZYYOuanwWPGRBodjAmqkydJI
kfF1Rrnh9rz0mfaTfwCaM5w3gvsa3XLOxUOg507AUo8AKoyx4EqHcgoa/H438lLFD59al2/84r42
7IjnmX47ce45IcjLHvtVaajdW7PdM0R4mI3EnoryY5T0guW1TM7fa19r7sjlJzE4KE974QGedY43
dyI+e2S5pvYVwwUw9Y9bzDb4whpkcpHit9nILVJpoicTd6EYpiHxSoTbKLu+6HwygBB9xdahgpj8
xoQVYmSu4/6Mt7ufxsS1YgnlGwKFWpZ0gSj1W5Fxf00QZr+IdTKQMwqtK58ygaVTd4hv6Mfuzz50
9M9pETli49TKgk3q/ee+4lW9QLh2b0K3vfwg9HbJhS4MqxWN346m6WkO0k9pAgLEDUaUa8hI/FyP
EcNYSNnGNksmge0TFRPZSoU6c63DBYCK/hl9Gf5QyJJq4lMJsyk3NrKmLYcM5iQAwrP86kyTwqH7
k8aRZQj2Coaq54ynbStl94jdffIgLLd0tnIXABDU3Ge5KLzX7wYdQDokrBnFh/jJXIf3v87BkFrb
ZmQboKlAZWo8DTBD99GPKgE0+0IycnlYBYcICyzF5KBBTYpSDYuC+MjQTZuZSgdQSJTFvl9RI/Qs
FvNm10FQ6wIstwA0mTAzvnxGOMSUaC3rRnCGFpw1dYUw7ms97Cw0QJs/r0KwQxoXti9PEVsksqDA
0aDqQ15Ocf6Bb5FxejwybVN3axJDtGzv0IdApJvq9cZGTYMsWogT+S8QVPcn9TYfL2j0pn5k5hOS
FF2i3QCtNTyn8Vgsqj1ghqQXNpQ/ZQ6z81TW9gJEd1+QKL8YBlhw7jCyt7NDbnY1eqcY737lJVSJ
Gf+e+ZjZ9zhE7Nq6K00BzFnBE9ATg7cAsvw7WIuFj5mUrKi6ZZhhl9zAnfp7U87zQdbt5ZfMik79
7XaT4EWP/REQv2v6yJ5HimUKULJvsgzHAHG4XQjpCzRtGeR8GoBdosbPHCDgGxtlFXQaTQvTbmMF
otmEu8Olyw8K71fwDRfg7c9IkMRUft6RyHRY1TWXtru7MVIVKIr4OhIot+GQBQh1Evk4kSDAz4o+
th3lbhyMVcasEG7x6lH5k1Elmq5Vb8w1utu0qm3Bx7PSWsFRd+ph9SsvXgQ9OEdhymlVf+bjU3yN
iJp2yUQTrdST88soX28h8mEq5v2uWiKBXzVM61MFzckVMElNTk5yE4ZfjRgEOm7gvtgENe/fuzXw
iqihh6P1kisZ3ydRlZ7/VkMHyd9sDjwAllwLaduJ08cqiv5UbBfMjIsomdtaf4NRSk56/EhENdau
xqAU7vZrKYFTaKe71dB0hdixaf+nnoMn9il0scBcenQYK824wGng2tCHrPO/v50xEGzc5RaSBtIe
8v4CLMBj6fFIIHWzaWSuoowLpRoIjh6FJSibqVWMzHYD4CAcvMc43Ish/NoeH+sOK2vp4fyUSbfZ
WGPXGv3FU1Z7VAYH91p4v+kJQIl6GUxwqDVrrN44ot26J81Wf6j1bSbpAoUk9udQW4dHjixyTTl4
i02Eh6lsTtECk0G2gjXU/MTlwa6q1CVe2UXrxGRI6zLzeW6LZKRa7tHE5ZH60qNGJ9gnZ2PfXphx
Ot0R92GBy2FxVpr0idW5t/ZgZn3WY2dlmimcd6IH9WOwdAR8gTWEdfOZWfEkqngg2Jpw35JeIhjw
pNdDh6kjcbc3lKHL3NslzfjClVu3e9cD5d5RJ2HJO4FdOhf6r2s9ZomBYmxOr4ZsLZDViMfH/B0K
992ucJOpxDILGKa1bOhDbCH5yUE3Fw9ePVhf3xjBXCYoA6ZGm+AJWtneXT4I4rE2LmXTCQMIZ7g9
GLGMOgiZeT2SyRK94N3xiZQ0GqTx8NcKGL1l4mif0GDMTTZYETqbNkc/BU2zXxoBtLYVHfcRMCew
x3ya2n7PUr5nUI/X5JEoMzOOubsoEqk8DYqcY34wH8SrMgmcbn3b157eNx4KgbyuxIBNXxKG/ZAS
Ju4h1tm0f1T+7ex9cSxdetO7v2kd96l5kZceotEwe4VeAUXvVPrCvSYJ1YXs1g70KwH67cuydvqf
BqoATE2+gppquH5XdM+yCbc+53ksRKcZ1pWT42wUwLEv/wmr//f6FNV86dx64TQQo4x2aqoVKisR
GUTKKzBzH9VgOp8sMeGDB2kErODYB9gUq7eA5fKW5YFjrOeAydW9/IdQKyM/MKYm0VXjdxDeZK9l
FUbZysqyDemPQBdwrVp42H7MamMWULw7vuopGz44bfiLGudT1IFIIJlmQr4GWLSd1MOh5dv1ArxZ
iki0JcANaYJoWUxZvr0xhKZieBIP1K6DD/hHVvlRAajktFBswGQojgUJQRl4WmI3iLSk7zg+R5PW
gKlb4lOs2PFfWvStx2rUEG7bn1WnhFZVAHv3UhpJf+nZpJpkYLuvPGKRVj21mqzRhfkXYJ+4tR7Q
8QdEGRsraKaP/n3AyzXF2XEa0lgWSYaJLkAb/R5kjjIp9TbdrdQ7jg4KvmuCfAg5A5/y769lEuwx
UZhpGKwO+fzFAtpa61jTZiSK4HsCu6L49+Z14wW1Glg+ei5Cj1ehtM1zebaPcK5Etowvd8cL4Hov
syAyrs2ZWgvRlBYQzvMcIrfvnr6qsmK4uZAmbNlpClBol2BI4uzPAcd2n0CNqYQPD3j/xG35xOTc
6vMPtx1eBxnoXsUPmauYXjgNUFFOpxy7ne4zCZEB25EJaM3+c7GHRE2UcufuLNafDaFvHBlqCwEN
+dbiQ3RtB7n/qSfV2L2AXz5zCUD3seJxjONYYVG3IgOvL1xgVVplbYePcWzF/AP7V45X2yS/Ue3I
it1O+fe03b1H+0IShgcYqvTSOvtGp+g0s5UQh5A/WANDaNHni8JLKvkoDMwiYs9SImLIVZUVA1hs
6OvD+m5rsAZy+kAH+MjDGyDgkAQPEbrBo7jedHxLttcUX+X7lSI5rx0ZGNxkTrRDfksL4539j5QK
60JbL2fmi0D00owlKZj9ibdCjihE3O2cjHQdc7cR6pnWH8VctWaX/b7eFFIGzlasKi0ZtA02b2em
lJhBwgAI7tszGY14nH1niFnjXyVoqw2TmTs9oBv1CKqgjO0Tg01KvsnnQxaAUIQ7ykc6wotP83Wv
xT8WqfE+O8I+D6zx5/+FX9aQi4goaBPW1nPHJM9p9EjyydV+oQeccuufT1a0trhRGLujeS4NChd3
gKJ24DxmW4yFVfntb9MdEr4croN20NO8NoJ7alXFKpu3iM2zc6wRAbSORbefZal8axPcKB++amuI
wxVLpkJ8hr9JMa5WK8CHPH1cXBB23a4qlmBidxCzeY1gsrg487S6unNX1WOISGracb+OrPs5j/en
GjkWUM+Gc6jqs+BQYZWkvpoaLvmTNi/xUENon7b2YMlB9bC0X+IRTRnIn794xUzk7pvZSfFZ0eQA
X95XzQC2LRTXF2BUMNpas9+ke+vYiJeK+aKiPq+UhAonhN6+23usjVHYrlLX5TXnx6QXYIZLvX87
9cGKBmxIqws6xwMwG7npFMX5VL6DnycbTQZelioyfUOVX8yarQDaNJyp6MrsrHzioGz2lVou43+I
O4jjGT+gZGLs+NBoZPSZWweds3ZIQmlY6BgC/jDNCmy1ZqJoBMhgKFhz3/V87cmNK81kO7rSRE8V
Nl7ju8FEUuOzYDBpE8UG4Eqvt3sXX2//67WQFE5SF2lhzoGtGCmcfufw5JURIKuZoCe36ehRExRZ
W+urscniVAYq+W9m5OHM842ADlpSPkY+Qv2iBD/KIYyimwOzdCrXqpPMmQ4PyWgqAreXEZk0mQed
AdTujj0vPpah6tCex8Flik6QnwhbrvlPwuwlfAyZzEEuTDqJIiOApxSmdq31sWaJPd0VCZ2OoTt5
LPH4JZEYKlp3K9IrNJWrhYFgzngHFj2ZGShtvPGaowsI+ObgP6mGtar5F8dpMSx4q/WsCH0gVNaR
SEv0UuMKIEfqDXXZ8FAfoxpI9gimzt3OoCz1PAvla6HepxaZBTXP8j8OMJjE8zrVELeD7PoVo6Ge
RbkNzne2K1KK+fawNIsPc7yhWxf08cZ8XulQMHKg12A/Tnn1QOGNNyR4oUXZ1fVhxYH/BjUx0Q1X
8Oc9/5rs7NvdB+ZCXPKQVYgpMiHnvux7IRrQSgYASzGmO0ypqFLBw/NhiOUKMaeIpSNeVsk6/1e4
zDkuh52nRzRnfGPr0JYIQSObRbv73KbJDlonfU0qdoNn6N498SBKQB2gY4OV+zOAsUbIX06SglU4
FZN7een50BgkKUtx41T4CUnZXSP+EJwkMF4E1KPrDq7vdbINYnEV6Kq1RSD4rDBParBd16vjC7V7
1jmbSRESEUM2I+9tvn8nSZqLrMRyiAjFbakuvPcZRasHYMKH8w1AjChnNfWuJX2bEoeDX16GyClG
cO8J/mIQwaBkfUThYZMR9leYF0LRmyBdz0zzyS2ed9NJ97y2R45FD+mKd23VPF4YcYfnzQXrlQjZ
eTJmn+OwgJmO2rZtkBOd7qCjOQChTehf0zZ+F72V0RCxrnA+PQ6046TfwpQpptxkIdbIrCZEGn7d
JmddpjTmV5jliij62k22dtDrGzJ1+r/ctkFxjVm2ZxvahGIfu+mILxwf/SItXgQgJ74hntsibQbb
S8Z2TrX0GoTwV6ZABS95nkEkoMjqiQtpuWuTG7StVHoeayyyGt1O4poHGNzAP2eIN+GvIZ0JY48A
AEwL8/L6LHty+4cbA8x5mbvPzR90YVxsDp3qtvOsJtUBog3Hq4M5c7R9Et5YJ/4G3Ann1tcqC3Z0
sQhv6Ln3KbkP9eUHtOc7BvyRS/LMqgfLmS4E/3Qq3NWe3aGsNNC2Ajife12L4iqExW224YH1mm30
2IStWX27PtjMWHpICfoxRycSBYewgzWcftbGEAoJLjHoWiK5Qvf4OfKYWWa8BN2E8FN2Tbok12Iy
Zox4Mg5zh18I9t4xLEG4aU+W4fU6Ef9kmCHrQiVwcE0b1nx9fDwNKVMl1O7W/VuYfOeWWcA0tUIA
LR2/IgAvkWkqFLZOmiAfw65Kbzpx+pFpejkI8bihNXy+qgkHxmODYnHMttXWWkAfzd+uXBkip//t
J4UQJqPfk2t6t3myMqGUiFyuDtcIrLgSmH5hIRwO1LjeSc6GXnuOCTQ15XF/mSGLd/KtPFB7lTfk
oFUZbPMKcbBy61MlDtNyQlqMZgKOGiajTbVaSt8v04VTO1OXH0mg1YeQvDOsX2KiVl6YF2mqPUd2
t3aoR+5XJ3GGfN5yLmLp6vSxzuNzSVS3hbNRIxQpGugJ3l+qv43xxo+4XRWjYvwKzbtmxDYOce1A
xNPqTa5i91sI84Sf31b1SFqUZfhI2gc6WaVc8xLb4uzy3QbYs2vJHyA+hahOMP3pOlBKF221IMce
qWUFm2i+ySxvgy4ewa7WEatTAR2h2eXsdibT4pOqeQHdNZn8PmPTsF2n1ttff2CIlhUbsVsxQpAB
zAoExxTVSqIeN2H+T/yOzmbzMHslFoVWVb2OgaqJCXSTr9sPxdVMM0eW780flCSDeRnAg8OQK1a2
CnX4/kW1ISlW828K4cnNxsr2UgtDVPglfftEVuPheXn4/Kd1pllfXmpndknw4LTnyyOnW7J7WcLg
OxfKYn/+DG9uozwoYW3P/9tG6DkEYehDSpPAo4n/sKLGF2ZnyLhrd5i7X44O2Oynh0X7Yg7KXPeK
pHCmfgcb9UNfu0OPESAw+QBS6RXJz3Pueb5QH6VEGbwNzTTN1XUtxTSjn8OEMaeS//KSkzUoNq8W
eEC3pVNMRruDrmvsvn710+luKPLfYGQLRJFiRP24orfb8j+mjyI0YrDLojpdjF0liyMcOgLPu5vE
8bL2ZFyi/48RJTJiDK0Mf/NHYO8RRgED9upWf4515DRN1LUMZF+Y05kjJI6Zd3MCTC+OFKQJCdcH
+jspii+mZFz5mXetYwOhNLCh1oobVBb1c8I1wghBl2xbEPQYhgxdcP1+S+TIxLbuRRwDvwDuNFKe
eVrDwlHBFIg/vpABTojKZauV3R1UfRngkeOJm2TjfWyXHdBX1xfmfTEGAVc1oxbX3jnVIZs0bGrW
RglcoVm+VMfJ0jn2W6ZbL87nGsdGpWubAucDaQ4A/9MSsNSTuc5Xj47CMuIyVBwbybIzrBUiT7CA
j3ttnhFs+aw9PU7opahDQdrICuclC0nDxAU0oeULzPD1oKZVK9fnjaMmpNSBemn9FWEBbAQeGJKK
/B3YgLrjRJWJVs4MNNYEZUnfL77ckk6l1PJkilplgB6Eyj95nXTVyFww8ui6PKgugqX+aoFwRe2k
A1XhOaf0dVOW5J/T+Ao/FLmv59x376ZTpluS0kR0VaGdAqMp1PddfjZ5Py0w45kbQ6SwBaByzFM0
zPTsxJl/3f8/+gEVAOly9jDUOOcRqRla2B6qfWdn9MeCRRE/F50Kbp68QSma+75NzGk+KgZ19TAs
X6iPr0nEaBjoNs0a7HdlCzLaaUPvNvQ/FCobMtoxlq5uqcAUQrAwxLcf/NCQ0sQoPkMoPG/1hxd0
nHHfpO/omPGgdnqun9RcVNcvWqbA1IwfMJJAqwTUE2o3dzoWTgFPZ96B6mBy4I3YbNGm8F8IeFB1
5qd8AbBAcPh3FPSNxtH9mZquZaowJZXtPz8PEg97LS+UbWYUe/vJEw5hoENdwjmE0lo3uf+t8lT1
er2wiZEq61DdoY9Ek0+dPbUM01mhqBwlZrdFG3cSTI2TEPwvsgEvvpgtlDSsSUL4VLDaiaD/K66S
gadc7RM9OUJirurWkpv91zad0OIlYhoYy0ukz0edWJ5O0hfcBrmkwgNrHX4wsWt9GspAmLH2Uufw
9bn8Vk20egZwP/MD2ikscdhkuHWsUf31WCPIJFtfqb7kTgl9o+sA9DDRTiYdE8fw+1fmDvdctJCm
jMXJCxJaYYQsvDeSGmYXWTz3/d1v+XrWdhuc7eQDeq/oYKADsBcck9tB70LBM/6q5ufoUIgcc9/u
4AkRwv+XUf0dpND9P6Jzq1xD9zUDQkIX81fP7OGCyJGM+iyq618VHEQfVCCn2oSndU+GNPj/gp6a
WNKd0cNkQPIyB8o/4/WVwFxQL+feJdYF2kADZk6XWQrsuaaYT3z6bNo2wRyo8GvnX1iHQ3NkphjM
WNxyzHwdQMYzohNM6kkIZr/kErxFwY6SZ05Yzy8JhGx5IQyzceAGZSTBBTPpKsOg/BDwuA2iV0da
jPDRaYeEJIOnnV+P+KAFZhOp4iS540Mn3lOJGsUT389DEZ/pkB/UBR3H45MViXRZWgazZDLeDH4X
t78Obc5Qa1IDUJlIBW1OZc4UW+bUWrgPB87+2L38ifMJTYfqA+n8o+bVKFbgBeUo/9HdlG0QsR5J
YYf7GtecNz2zedms7+6tjhts7EGJkp57k0CERLvg7aPJtht/JK1l6yKK5e3pxNZO1nFtNRp1RWtU
SUVExXfbNj9D0c0XaTzv+imLvM1tR3MdZwck+vubJYgYmrO18sWKUXWx/yy8P0Uq1v1ZV0g2M5DG
AIqiJ6Y10pRcvyG49OSF2h4/vXLLrkPteklTxchFff2WpPXmRURfO0j6GuNXvbqZcyOe5tQl6pUD
t03jFjwtOWYq1z8svYDsbqJjdBrpLjJ0+dPbhidnIgcxsd7SiKT7/l0zvMzIM53wkvmW1a4rzPxl
YiPflqku3gYccNYQlbsi49nZTclCVh9yEMgb0iSkZkQRK6MCssYgoNXjf9TjYMF7xGjDtmTfEnvW
NP27ttACtcZUXIW/Y5NfsxieLdcVdgl4Y7SqWvlNuVXU3BHoR0pA/8DEIAiLKaYwU+BUN+f5bInt
8yOetQ2dHHNTi4Hp9Int6pvg9X4CwV4xeziL8Rz7MTfWqHsgvnCPq350/qYNAW9ejAcMKoo0I/rr
dUH2wzBDKWUJUafWGcIsPYNvguaC/wqHSdU6MmnOUrjFqAc6DMXo3OvgGHRF3i8/A3Rl9VgM85Qq
TM8H4CT3LBqpSOP8Pe6yW5/3USRoGGNdSuPjeBp4vEoO9a64FEoMpCT7i8wnFV1PGuucNCuadupG
95bElXAD01/hdCmWC6Uhk21RDqBXkaYqB95jkw5CDrLQGRCvpAiQ0uzGNGNS5PaVODPQAnJfgKD/
vYN3tJ9HiYOD+2SwQB5iTKpT3QqT+k0eEXUSFbmet9RWnYZ6xYL8/4fankpEGTr4+ZY2GovPbbyC
aHyl2/ZT70Esk/W1kxIiupY7ckKlMMU0fPR0jga3B2bg2STJroABM5ymOQX9ncfe4Q4re1Cd7tRL
JrP2xaM35DYkeW46jgvQerSEe8zTSrJ+ln1Ftf2Xlbdwzr+mjcOwUJ+cZpf/NKOlN/i2Qbc43hfJ
cpWkR5ltwjl36WzdzflhXbHUTwA9Qp9jPbIH3d3GouaiNnZ1rtSvr2eu/cJYrOllQXBf/gOV8BMj
KmG9dtQ6S2f8ulixdnB/VRA5f1GcXRD+mj9H5FNbl1b88aGLXTAka5gbs6665QrvoBKp6enphM5d
+/m0ZI2cwUMymN9l8und8mZ7x+Vq43JDtnssVNmFEFmvIO3SXkWFT+xwOniQdodYsRLpg2IW6ZMv
q8+wak54jKqw4Ex2rPRizwrMK+V0lNPwu3z/X+g1ZwudmNzRPztKXTsZUKD7w1mZf7nj9kVSTvfF
CX60ZeMZRneX2GXEDdG317aL1ZV13lMrGRDHD1KQgi4O+7x48JMKGtmNWmiEK9uB8ZTQ8kfQjmrX
3VTa6uzVdQ9TRRjyckLvHHsGuTITP1Sntp2qLSxmFPnuHOrxJmFR9kiZm1xpVjS+QgMPVbRYR5rU
4VygbajaXnc4nhlSZyTfFw4+XIe/r0hIgRlafvbsN3wmgra41nUXf7dXPKBUc1tnB0RaIvnmj2BB
R/0HwOcukKnO+YzrG2i9CcXrmYWU3upIErLvGXBZRAEo4nzR9lUd09aHZXdPHApiQP8nCpJTASc0
c7f0Dig7tK4AVmgEI0YvGUUmwDG55vMRF/jiKCc4MaGWWQ8EA0ka7bVUlGHl+/31BWj3ps3UMUDS
rzLNc95FqVPrHNa2z1dK2Xy5ySFXTtq5n91LGM0TIo7vLTg3sGPy1ouQeH09JGe7g584oqLiKiB4
MTIJGp0W/81PYGfo3clPKc0lcPb7yErZNisIt5veoD+fLcuq/BiCFgz8PFbxIJ+DjKF+sAM1yx1e
uCUK/osDKPILGf6JlswP5DZp0jLz0GKQI5iqOllrdao2xNcsfpCil8Xpdu/XWWz5BRgdVVY20NOf
UA2vddn+2JCt3vsh8HvhcyowimdjRhGQlpYF6l9YSGLSKxGdG9HcFO2PasMEdsiBegj4kavLD3w1
CcZli9fFssozjzLBg3VZNNvMaVV/bybM4mj1ItPW6G3uagUS3BvVrZZsrruh4NMoPZ6KRBFSdkcr
YwPyi6OCyhIgmQMw2C0HX1mmEFni4CkbulX6/tC7BJDlGpx/vZNltSCyIY7ldSjhPIGTYlU7Lm1Z
SRTt7rzuSdyQ7dKN3KxwZkoJvAdHQQYU5cyKHkeHgs4wvxaZ6guXoTylvvqZi1qp+JdKi9GoH1jh
KmNtQhuSeRMhOCETMJD2PCMQsah8Z2huoSUkJeAbnR1kqttuHsgQtzZ5FXHmH5m0FpSTcjNf155G
9j/9xaHMt5wLZEosHkYHtgDED7g2zV3a2QjP8Zrrd702eNGKh1zXxJad2nxBeR7+JeJbA3ykM+I1
Bc7yi+lTIlrfbHgwQEw40DRZu4Zq81dqf8UoObKEYEoGKic37OsPKLapl+Ka0pyUXyTwHguD2dd+
4Aqd01cNtYmkSkOrkRD6cfdXY43MOI/acupfhkUy+GTqud/QAw7G/KHQxbCKuXmKu4erM8rlOcJf
Wesf2+nLNVCaz+nqsasJAxWZSWBc7l+9EI3ZmoSbVebWBrgX1fEGW2ju5gxp7i04c0dodOUPOk+b
Wstuwsj85vlLKovHrpddBgXQ/JqSUkxK4hJ+klvzx8vFa5z9Oi4H+G9jxmW442MsxJCbFGR4tzQv
rY7xseB9Svm+TCbMJWGb8UjDrItVyFZXSaI6PJ+3LlDKz3Ouq4YgQpaICFz9D4/vW2JiZKIxNB8Q
gJMH+RQE+bfVsPocw7JGXiol/iCW4CSeQOw/Cf8Hjn/dAYBsRZbeAtizazwylGOWsb868Syj9GoT
x+EyPJHtHyT+3CRxGLIAdOnkaZIPdj9YTd8g+G06ucVNSBopeEzKSzGBDMPBsVR1OEcE1F86GfY4
ZoYlmFugExhmPtIMs0DICuDGOhvyHyQZdWXg0xe0yTK0JKTuLP94+LuKeTKFbNp/c8ez1DOclWd1
av5FNaF74h8oaHPhJACshmBneKrpFUqZmS8cCXyqE99KCybjinyC8RvRWZy2+WUhN1gKWrW6QFd/
s6cQzkkZdZRcst9mAbXCVDeGxZDmiQTimk11AEMfRj+ay3rKvPQ46vHQpxEuoqyOXXDJctqWzxFU
UXkzcEYEso4i54zymikKw4+2JweuIhP0L24gER5N9eUljatbQfyilyYHCPq9RG//k1z5dW5kXbQF
e8WGOci2tN/mN+oYOscN9FZIjXXHsE30mSnBQKbBDjW6jXV05RSF1a5a9p6tD+Z9wiNN8rU2z9BM
G53Dzk5noT8xh7sB/dMxhmzTG9SwFLVD+CqsjryC22Dw9AYFwsCANsRhPO/tPIQWYDbK4CWoMxOw
Qj5dZ114L1RFjO+gXJcCjvzNZI08Yhw/VOlEKb7KGv9J+TNSrtq/IrZWfc2J69QhA/HwELRtv8Hy
FNACBl3aziRzJ1fdHLAHKk0ygGShI27AelDaW4vQjKgjDuxNvJApCogbQzjaYAHSSZTelAKZy7GG
LXyUqILpUuZewQDRbW9pw5io8Kli9qOSpiC6f1fyl6p15ZsEBso8Fig6ygEh5YmHAtuR3Si5RBqC
9109Wp42ZYeKNJT0Zh8y9/w82Ihv/pD++ExJxFMODath08m0va3mgbl3TJXFBK70Dl7zplwVSxjn
mtgkEN+7zZHIqIYfdZluYVbdMxtrlfJfA6xigcVS46WlF71fTUqFAUIcU8pSPIzOX07AHTbfNhj2
B32xIp7BZ4tHZwFliUGta6lP+l+Zy6KY0UB3cLGB7dc0IxQHId6Mcw3mgvdk6elKAbcbwfRNz5az
t0NNO6oxRM53ZnzPLDJLvDZ/dISj5Dyd6sc9d1HFt7HaTdg31xoY2EDV1FUpSyuOex2YsJXbGXOw
zE+lZRyvp4scAwvjTsyFCrhWR02n+Z7I0ikqsOV3J30cCLMVHbPDnLaIKWlfdA62QA5oXG38gCvw
Ta6/FTAnANFgeiaFdikAqr8K7/H1pDXRzaLgQoWf6n5P+QXdAqgaHL1eb+kdvAbHyN3ixoGppl/b
BsJetsrq0eoX56qBnOjA13mWSq2laZ3aLflfBmE9PqB2kDJtUe3J7uoHqYtiOYhO8Rwct6GkUVPP
ZeLlEjnPK8pgRssM9kJV/L8FTTGBFfPXNatBs8kFC49p/L+IGl6Z3TnsR1xKoe2PBOivfXIbwfq6
dckAHrBLYmV7KIFpKAfx08SFsgH4lg+JN0BZKujn8ENMSkuP/q9JVAqHR2EDCmV5rqYTQdHZIU9z
3Uw2MDzJtAgG9WxGwDsw0uREgwEBOdUbs5neRuH7i7qOmfJYGgEsVpsGOa0sx0a1hgAlqs3VtQca
63bvOAkSD5Qp3C87J815T1WwZVCS6kc3WXb9IXltu3oqYskUzOam4FL7VsVh7LpGxHSdhnIssB9Y
NiOzzER8oUVPKleQJ15y7aYhvv9KLH2CCCwAt/PjEFtlBC74srmE4pACQEhYK79UvK4k3Pay5WTJ
tFeDIAvQwSM0rUaQfZzoNPO0zgLjcB/KZH6JktlRufbGGbMTRJLrK2CoglhAHqJmYZBISDnQr8/x
AEwEYIXLBZjNgbgT5keP9PqJJIIZPhrpV3/o+VI7D5jOW/QWWFhOsZDLccERxbjRGcOJRNLNMDGb
tbz28NjijyqM//akiUTaufeP6YSHleeShh/iDhgb87SBqZoi7c9nqlEpd2vHUNdR54/i+KzcMCcW
WzYowBMidJn0oWlIP75O+4xCtG+CCswiPPDW9uYvyVOXM454OTlzFGGa/rlogkFj/tFhPrQ5u/BB
XkWhCowuxIlDJ4kCJvy4XmahR2JSgPQFZTIcBF3f1PqN8MSdAk/QgJzGbyCUAa2kD9ZUrmgJJ/Gj
M8vyMv2UcYTt7J3Chkc1KxO6PQW492/KUuXJ6i+dGOaWpFkN0gC5sa739J+On9mwXUBXP9cp7l/B
kwPFIfNjg58hpQGH2/wWmMwViTAnzhlcbDLOLMOfUJgXmTQKD4fndlQ2lNN68olQbOOGY34GhMMg
oL2DvuwaXDHOxrsdIrjSZ5hDhugIJ62KJ3aIIQXX+FFp5OUWGbMn8nB5ZRMsyAHPRBRg/8MNI4zL
kFyRRIH4fiwLQuhKWBelWQyVKmSmVl1D6IAqAYwIkrj6AHQV+rEQgPYnjAphCS7h5A+oJ/uXwIA8
ZnnBOqgSKOAe3RcY6UcT+3X5lUZURs2IZm5SuaczjHal7HRmGX9dnea8oVai4sdQwlgl0fyrHnWd
4Dmz5xwNNiKRWf5vFA/JMZwj8qYDb1+IVJcesLWOLO+Wn6nH5FkgLWH5PXvk8K0xrqaIIaFSuojJ
5+OpmD27SM4bRleHjjIiAZZxb2PEzU/g1lbljmOlWwzBAugpkYWQUHmrM7edbOu2Zb1giUrW5N8J
TGKlQswe04xiPKIZAL+xCT+UjbICOzvkWzNWT4qaXP3Q9OtCAesDKSYtzIYwqzSAlelgDGNt8zmB
dq1R0tH6PL6YSm4z+B/CQmuG633/efYyUHhFHOzMXYKEYGxnUfBqfI/qCdKl24TlAEqoAqvoBqsc
jX3fuNYRoomArZp2OTanVmidcTXUO5OG+PX8cF9tv1qqQx8s5sGajfsmMQUqZJ+FQKqx+n+u9lhk
BOrCFrkpoTaZjU4nsnz7Uuap301lbj2vFCyVaBQrtEB5A5hy/WxlKBaJ/7VRTLsj0HBgIs7WEksm
DK8GMe8lZGVkwm04oz0oITkZSw6kr5vOaZgAABqyC8uc6PULAU61HHB62HHYglddZ+hBU5637NpX
vS0M2gxdDYmVbQlS4SEwc9bpvNJ/3lrhmXw/C65ecWP5iMgmnicMErkb4cjAaoTmXAfSgdre9JVX
kZBOinDt8WBJ27aryDFF4AaZVETvw9R4ZnHzapw5SDzvCyOKTUVgtxCQz4HAYu0Lfwhr5jchbnnW
v19GTgcBBpsxp3eT+cWlmWY43/ol010oYkw1uWRxmoyLz5OsJOaM7WkMG3vNlnx671xDVhJKDfmE
kujg9nx0xW4FRKgfrkhW6GSLcjGQBZ9l0ahpwqYJ0SL77kweNWFPq+TUnYDnj4RvBeFBVhKcZ4D7
xLla5DpGHInupMtP1ZOwHJuNpx2gdKM2LwKHNZMks1Y6upZlfcvZYq7YDbYZFZTlOOkI2b1NGDvP
EFJ/lagWLEKW2j9cuUADWAkaIiesm8uULDGe3N5MZnTTEPoc//YSSnMAjlnltEh0weNghQgqvqNh
jcFMJp1C9LdAu3VFmQKVho9I8ugaKK9oHVCzYHdLUh2opq/pYWkWKrj4FMm/31AXMyIAdQ8goyUm
UPgdK2ULYne4cbLVswN6cYcfEIRAFD4ydaSxr2wW8n2Ro7X4qjOdIl7KBtSb5gngwS4/Qp9qGB9V
pUwP9n6n+XqrZDnJdX/Lll08WZVaLZilbrV89BYr/XmKce30k1yzWObmtF8uoDP7NIqyoHoFZ3Rz
DeWQKE17l5axtLdk6th9nODAFUNpDWORMg/NzoMN3PVpoPow5CJ7fNlvVDi41wVmxudp687W/cO3
cmCJrzVVjV2cYZrsVk64oSkqEfsdruTVYsPckqh9lqVLgzx+4NDASRkXdbW2XIo0kOA2EBgru2ju
9X8yytygx+xNK/FFesb3EV1s3FgaHo43zkRvRaY5qRxrv3AeXWA1lbIG+3vjZONv/gKoPQTkndZO
FJfE20NFxHeF+FPNurECOoPuAY5mTk2F2c5QAfxv4kHSpmLP7YZH20MNRuqRPMLBYPINUbKbpe+/
Al96QQUyNW0Enqq3M4HugOc4Q92Fms5g9eit2uY625SDEuZh1dg6ZyiM2jy43G2e1JO+OuQfFBMc
+iAq3fO3h9YvdqWat+tyAEw4BrL2RG2CTo/P1PS36vqEKPBu+tW23kahehkVYBYRdt+nUBpFhrU8
kTrb4Z/34+kGyfgjCuJXUH57uYmRy/6E8JVa+otxNVX0BvFhOHkGKD+HD9JIaNA7tSv4qk+YBrmD
/vSQTEXTdJyeExkzSBy30iUg1LxJ7bNzMIxPqqOGdG2iR0xoPdxyNfvqvbu0P5Mtk5QIS+MILaR1
Bo0I8d/KHDYI1JKCtg+bQMMiAHk9TjsX5y46mz4WYFmhMOqpr+ancEAa3ABK6fbP5dlyR3U97wN+
myVzDiBYstX4p+kE6eBJgm/v5Z28vik46/iSTJvzQ8vT5QFmQyofUL1Fm6AczLNdAmyuagciCbRV
esYCgoM25Zk4kHKIWwok3uz1W7TgsnO8zH91c6we9D4WgjSlmDErjlmVDDVdWzTMZsG6Dm206VYi
pQ5I1r7IOaVCKgCTSVpGjLWZx855J1A1256b4359cbmWWUs2zQeQt+bd9Cla6KyqqYMIjaV6BuG3
72HfEr9L5xljFfLfbFXWlAsVs1VQ+Kpo2BQ5OAojXDud8FbgxS4WFCj0D8a7oqoXea6+i1TB0lCs
5gtw3+OosUqVfe0JbZIRCpaHgErqonGUVwc7vuRL6haIQepIhsNUMiuvIAlzqdINgAC6yAfRmlMz
S0qDC6wKgERH2JFPvlILheMP2ssRQWj8FpdiUUBGYEq1iUDWgceoUWCm4DL+m3KPMrq/eF6ajBCL
pom1m/MkrU61t+z6E5fwHy7e/s6ooMan+StmeLXQqHs9TWVm+m98uWGBBrYKvIVI7ND0NXj4UY9p
TMbCULGNLKm0IjS4UnzgHVjxXxbaxANKggXjqfd/7eIMkMoqIrBDTYVXymf6PstQMC8FohXESYIX
PSqe4f4hPSeWAKtEkLFZifGvoLWTo2NKShlwreiD7n7RaZ80+o/10N/Mc0f5mFFSubagcWQ/8MMR
BIteB8ahVuQMi7NRH57lJLYNg/VDmH+q4Uhbetuhf8akMcvq7HN3aOyJ9TeiwBdZSlEjlapMXTX1
G8hQR4LeU9uvJjJhwEe7dU/MGbl0ziS96xEfUIKFJBwxqmO/O6vFeZ8MSamBNwzfVwGMfbqYVau+
re/h93CPMZIneonnSrqR5vZ848XjyZRJh0Yo4lRgGuhNtQhnXhFj8oIXZYeOYFJW234gPtoWPbNa
K5zYtV1ODh9gKWLxOK7DTzC0guPNbP42+3ddPoPf2uYHLTwE6KVk71XqNQh2LdeCEWK2Xtiv9xz2
GZFzkSZ+0b7YHwUo3KVWBaoAPCoEyjpRWZ/vKdPdm/2rss9odLIav/7VF9QowN4pDkn2yznyF1oc
JekYwhgcJZw/23sMb44Ns1n+wwE7z5UG0kKTTmBQcbVv4tt4yQ6q3szZUUn57V6dHkupCzE4ndLz
Hz3rZnUkO+vaYSrCxBWpscqTwwK9HGDSu7hA1RXTfJbE3ri5D3RYLreZG2CmYlD2YWxYLc4YHpOV
cXvBBYtgiGnV56QdmglVyjqoZBsx0JRCGu9p9JCnC05maECl/OOOeJx2UlZYZ6Zh0IUYo7BuqS/V
iCVmWWP5Bu9ftwRMUf74gxg8pVD75GobsQJhuOvIdfDe8KbqFNXffzV+z0DmnrJbwUgeYrPz8n6p
RuC+YMfO8unmeeT7heEK63VAmfTmzFPm5xAiJesvdAWXns0bq6JeLLrF/kteo/b3r5ZuYyiaWpmo
ZsRW1zcEqDDQynyCLW0MXd/524cSP4SI2d//y9aYKt6UJ625AjG0Joc/597FnB0GbaYvyoLp5Q4f
/EM8cpszbUVsAlF+wMRB3eA8B2mqcZsum50Q/bIjOQNVEh3zIRktOg3FvtTgPVcVGHWQ2Gx0jMlw
m44cXgmYwNqMl739dKodKZs/4ByEb2hBV/PrNkvW4NiDeIwsjb8QCiCSFsHCTaBdYV+T8ZgFIUsm
dTMMfr95hQIotCKRKDR6KThs0px1nx1z/1BuQBo6B6oVU4JkjX3q3bqVQEBjjM+ypYATg1yw/tHJ
5bQRIoyss+EXM54SuOo2rNVkQQAXwily3RMacEEjM1LVILyaLTj7GMmNayUYFlyYFh1nb87Fs3pz
zvIvRmBqPfIpm7zzhR0/2AvN3xMLyJwZW/HJsGbUwOGvLTU4sw/E7qvXLr6+nsXWmqPRreNkSyi1
tuD3r8+v4+oa6konCFS3t1AVhhbR9YF6JyYsgN7koSLur0TMUjy2XrgXmjOCBPMFjmGQTwFrgJ0F
isHj8W6E30mkroRG6FwL+RWaCMdDMIK7edV+GcJ5L0AVFPIp948YlpQsTbNvF6u5IvXX1pU6oG4i
VqTydjG5fhHOBvttfTveejhIj3S5M7+IyPVHSU+xd/QvE4/BBNtJeR8L2ukeO8qWpPnJ37YaScIi
KsWzjT5hzfMrzfnTyTD91VDVPjIPYtxdPP+PXyxJ8J1rv8tUH8g8vmD8Slkl065raBFgJ6f5xDgn
kN1VAyF6dHPmTCqVUhIzjMdgN3pzk7KwinqehK3NGX5MszhdP2Q2QZdHiZJzVVA99O3qvTPGUAw0
NFIQV7UxhYaq5v0Q3DKXZsqCCa63JBWryT24TaZRhQw+AFR/hWD4Qn+PY+vPalCizbs+TUT1yzzi
1YHGAYgpAyGSE9aAXpbDhaJ9fJRHEwBLhIli90w2R0s89r5qAjkW+I/v8fFpSGBV9OfloYdbDVn5
XqlhDYildkuVrttosJjkvju5Z0TeZQyiWK8BNqqNG3ckXmvF/N4V4tfdQzQ7tzDzs/9a3If3Ji+E
zuAh8v2Lb/LP5QOIbA2BtcNUfEhwfFDegOKwx747eikVJtYJZFlTxwphMFkxg+3OaTT6dEyo4tNc
F/Ld/lVMgCMpx25F9gBh8O/CXE/JbKt5d/Rl4trPR2Og8b2WqXabOA4dAa0Y+IAMGQMPW5844nOY
QiEjQXdjMwrOyU7hwZXBpAWc0AW4BkVAz2OJLWnl84uocsWBzs6s09wZEcYsF4+H2q8jfyqF6sze
KWQqN8cih67G/Hq3snJOtT/cuCn48yRm4bnrShrYhWtNSGEJLK0LH7SffonqLXkMrMgEYJ5miM8k
YEgu24+137tY/kHr4vm/FZ2t6rRtC/gtuszQ59GrexLeKmgwMmpyJ0p9k4K6g9fbtyvb3cLums94
61GfS0zszua8QKpZYn31qtzF4l0JtEyQpefa/Nfv1n46ENx67B1+AH+dgtu0++1PB8Ju+AFOFYai
AIQbJBt+C12ZJFy4xrENxoxVTV8KaXN3aR/Sjc7OWS1Z7RoZO/2Pnbg/KNEDaY3NcLgVsaatiZJH
Xvp8DoXhmMyltOszpNXmtX7uipEA9OyYLzoaIviW+U2qyMkj9lLtvqe31gzld0QNY9/lXXdsAGFO
DvILpWy7nJPfusW18qrmlOkL27kvCs5KhlFNJccZdL66DYg0RDv8eDA8+qtU2SJAz2GQ3a0C7WLL
YS+LUfulZ2oot3kuvAnak6K14rkOvee5st/u14vUKP95eVRAGVpB3pbdJnesEqGz+E4XY9ZdTCTT
60sacAHapWdi4HEV/zuR6Yt03ltxXZfp3BAkSoxZ4SIu412uFbYpA4lUyGcAjhNFI9ZmOqnvYq6h
n4NA3kHXnGTDmctnOiDe5oATtU+49QrIOF3jcUVgW+vZtFUjkOLgdkBVeRZihBKn26QpufT/5Ov1
ky6QZmEmxqOMM6kdZXqJAfZllaa0HTf2PrA4CGroNUr4ww6nw1rwy8ZDk3+R/Ad0wLrD8RhnCTz1
E6CIeH1trqrSO8zyB+ttxDCokp6k7y9TXm54uwDllYD/NHixX3gBWTStfurHJDUVDilFtOwFHQfO
M68lmLQqTne/+sSb0CEX558V2+2BFelRZc22MV9yebTaG+n71kJwE17lWA3/6sZSQihmi/YsF1HD
KugrXPTxvLixHNro44M1v2baU7XyZoWhtTJY1svN6xSWo60iSGxr/c2oj0pnhXuxa+f8GlTnpKF7
jIoCo89P4NWSQJ5VnH1aLL0pxNBWhYp8Hb/8x1EPpkZ7WMx6Pn310AURBh/7oYEAzJMkoN+0uhqI
UK8eIMU7V2xRj37eppKB7N0sh1pdg8Fnh1jCYOWBlCVIKyoGBJqgNnVd88Gn1vnF4E2nwW+mpQ44
ENS9l/L7RJo3Ll4x2WrNxcGqRmPJSgzaDRvTRhD0cVcqNSk3i7iAgCnishJhrfw2RD3COYRq2BG2
il7mqQBrYXGDw5l39u1UnsrOUFAmeLFQbzqeA7Fx2obBcz6LlTfu4AooxnVwRCFTpZvtMYaNy8qQ
GqlVRbDYLSWYHLGhvhl8o2FFnrhoa8/PqdQpns3mC6eGRBQ6wbksG5FIqYvFzvfK1G4z5Fn6VpYq
n59Tv2YKJc7ESINVkMVsJDng3IA4MUY6fvXhXvwpIXbtCIpyMM9P9+JuNhYzOYMieFzmce92Fdh2
RRbjkOWdbLkivac9Xd9gLuL0Kc/bqmTX7sGbON7Fo3In2027C89ka6jXYC7Kcxs9JTUq/xbq8Pc9
h4OuqUNUEVxqpoJ64UVciTrXO9RP/jAbWpRwc3qoWZhD+wrxSqJ3dD/+p90HV2hR2cu0tTRcUMyz
DEBx7fnnhOEC9002/5B16J8KUHjaKK0llIRwA2dhczAuE6iN+IBsQWLM2h5n+InridMGKcLRDooV
/LKFluAMAVDS4YA9+cKwUNazlrRzO544Yo1agCszN7AjUccGNDOTMLMPb5EBg2M//xAnT/XddQGF
V5JefJXqolPLfD+GTtjL5Q3qnxVQ0mM/Do3Klju2DNNPuub+wfsXoi77UOtJ3ZUzDNvSX9LtKyQJ
U7PE3fQmzaICMtbxJoPRUH480l/Dloycn8Ag4AdfaqVc6yr8RXnbV/Km7DOyDo8xZq6eQr/XCfNO
2I8F0QDTBrkZVniYmJu3xUHUegxh/k0fdI0rhork9hnQ2MXKuwJZVZ7K2N3En3KtrVSqFF2JU0Xc
uVRVfLEQtlQEiJmUwLAgNVSA7qhVPa/efRuQPtN+ORuVkV5Q1qmbyHGi61tTWa1G7/BZv1ckaC1K
c2Kl5dVdd7vDy+FkPLEDnHtQw70euPdY5H9cTb+A9b4bOCVaZsrV6Nh77NqlIlRP2bQslhZdTQpM
WXkBylnV39RxCxDxnHPvQKXjESjNfOunPacI1BCaCYvqP4BAEQ+orMoJSqcGMKN0pOzkmKouOiB1
jFZ50WNuA6Py/LghNi+afj298nZG/4n7cL28Kj+DS2McE8OYWtwhM8G0Hw0AbuW0YNVTICQNxb1a
D3LnoieazDWhkgjWIIn8AvZ5X4MAfRdDyzxh90uJVZjUYu9fvQLl+84wmsJNR5VznBAC/GFBymE5
LQZ/7JDJfHkRW8m8Cpj8B41UkH2Mx0LylzthPDMrbL0otmthP4fYZCK1FLE8Wpj0ccvhvInGfJLi
8qZ/cqn9nYRRc9Ie6O3kFie+az7gmyMy1p7LY8nBK3VOORQ66m9VKVz4KbOF22rnEHq74SWzmC6A
ZdcfGyW/ecdIlLU0RznfvX7s+QW1k+T7IoghVNbA0w30rtbrCQCea51d4mPn9Ciec03gVVIy8eej
RhKA5AGTnV4pX+4xY4uWfFba7rBfDF32e8gSTRfiKRE9TBGoB1CG9cbg36KxrhOnrbe1UTXLuHpL
VtQ9KHtf3BAQnatzOtPyoFykspkeUVyWN6UJVK23u554jth2ojhtZl/C/F3434WqGI+yqydnEN4Y
QnlxjFGx3dptviMQCgu40uvTnxAg78V5GlXRidlxsFPzXMuFW/qiaL7dBFKaqlh7Ulw1QhxuM/D2
ttSmVwv7twihFVfPS//2wbXRF1Bm0/CfJ9aQ7p7Wb8cD+Z4uKX4sRlGF+7ZCczHilMV5lcUE9Neg
u98SJPE7Tmm3iG6b1r02xmvGgYotPU4MamEHeT+xyK6huRrfXxy7H3etwjER0fIQRf2B4JeVruPZ
kqOxlmZyFPJ8aw3dxFiLn4tlrsXnzromnsd1jfgHyo8B+wDxyBV6qeopWPxsJcMqyM+h8Fo4ZHUC
mdCCw4EL+Gep9YutD2v4sWDe5Aqw0/2DZIh7J4IDutz5TYgLcixnVYGHGTSVdSgXQGA4aluJr0De
8AL+jBbphm7oO5JKfrYASX+3/EbhlxmN5YzfSi0QVUsZb19IRbsPXjpJE+3yzOzEKcRCp3wFR+D+
L11bzkwSkXtfG8535iesso+argfNEr2K9dUvrI9seTWZFpCjd3bMmSihWQ3dyClFxkL1I4Qk+V3J
9Ky9Pzs6vXmIqZte9B2KK6aqFJOKsc6YTvttwo/gAWSqbLCQ4Di7zhq4W7jj9/3/UHHCc1CsJyhV
Wd2LwYsGtR69lMGwHXCYpB6EOsGinVzNXjoAGhGa29Y8XMoKNqvRnVsSpQTPHzV92f2yPg+qiuM6
E8BIXUaLIaJnqavdrFTcLHYuPXkoB3Q6WYHsf40vK6A2ibmyoMMVG6GEqBME8voxDWgmmI7c5fbc
atCbPGDUBPBtPuJBGqTO4fbJRoTfD1kE8hM+dqDp4IgzWcpmL8lucKBa6IVRCo+twFyuGow3bVqe
474SqJ1DpFXFzujLathcr36HucHjGtZ0QniZ8V0UzMsAV+q3PjYsnneE3gMwimfwAkqARXtWNjdh
2w/5J7K02UniNndJP1qJXUxS8U9K/8Bo7yrNBcmOCkW6upXk6xYovwBjA+lh/ESn+LbDtUOyAO3m
SQ9tvGA+zk4JWpI3UK929oAYv7oM+6pPU/tNdoWMd8Gt1TEdsWLTZmwSTBJPG8OKfLwgbrKHQo7u
MhDoYKJiS/vKkXcs2ZHQS6TBDTn0oL4XJYYqGtvoIMmPCpePu7ptV1bzrUqWJX1oOfBIloPXMKgt
N8vO/rGB9uzmpjviEJ/0dMgsHYLxmV5MQ94Q/ZIZbL3YYCHfeDR7kfvsscTBwtB4tqYpT9WbHsoK
+o2VJDEBEZcmxtOq1/Ddm87iN5VoXUio0I7Gka5gqOCW1AYIF3K+sIJtgoPvtuDAomPpG+Pt/0iZ
NU5Ue5IPQ0PucOMnMcGSWpD5Wr96GP4lByyn1fq1xLX42XAZc9+cmTmLQEFfhGgScCRhVo/OKoOP
fLpKix02NkXxz+GuThNoAudYvIxd3m3nTZYpqUfgjwlOoj7Uwngyot0TYqFQ+RIrtKR4fm0ak/Qr
mGobuUy/m4GoBKumKJcQDTWksX1Gg8Gbxs7Pwx0Q6hh09gLg/kAV6qP36+EyhVTGh8fP9DPNTK5C
3yaweAHVlGzlquTFrUY3sDAEDt46BxdESUEQ0skJbH+SOhQt4BJrTVjRxpNRcwBLPNHfZ5B0ud6Q
fz7E0zO1sJ/VK4IJeFmDGyyDLwGpa5VdrIEjsGl0OBoR9sUaPqr3/a/00tWNv7eXY1yJ1Ff0oL7J
gGk1KQIyQLOTRDfkoxISYEe/FCoUWabnm5aKZtjoxDKu/GwFK7D1olqGyXdP9kARaOszTpIF8aSp
71Gvp+ni0hwiRGDz/A/l/meyAQxUgzuN356GpapVm40mPOEuesGuM1a3f5sp7zrLejjKe1hvec18
8O3wLmBnCZiwa2TejbRtUEV3obcpyC5hxddAdf3+tnAiYk8i4klpcI6Vznj/osY/5D2V4WgnjGPJ
pJGhsRLZwaMiRml9Pw4OXMEbkwde02lNDgBVA/YDgBoo++H3OJMe8DDlIWRTJXkSGxCmzqrBrW0Q
wgjsId/z83pKBTi7CP1YfV2kxc4gEDZRqS0+Gr2loqBIoLtnyOlxPGDTk7AdiUfs7oqwQZEY8QLc
sHO9YW3l3yV8VxPlB1LenrZASwy+s1ns93lXub9LKnqcjN9YWE3Grl2Nquo+ZJ75iP5Czg7aKFRH
9DdSn7IckjYrjFx1dWckyKOOjKI8R7xzCO2b+CqqskEvDFjfzFpTrDEv46sslqquBz2T9dKEODyY
1mAhPlK8oFp1urGW6gx1l4JRkwd+5A0n/YUgZd8YUGSmyBC/lHLH/FTowIKLmzPyFj5mYiSItIyk
DRfSfRr+QjPtMzODSsYlc+zygnR2vPUaW3Sj40/+Jq2qYKRaMHAjNQ5S1OhLKObjz8l+s1KAQ+gR
KueZldBMHG6He5jZa7NUbDJJv2du71UOXSTCrvXueBsY74KUVX804jK83DEithPf333rtTEIKMxl
YlFCF9rdWG63IZai7kzOdVc7EyJv+h47SnUbkeOoWGfu69ioaqzUJohpl/3qbZXmgkoTEbOzf1BP
P8Lb5LwOTwfjYeFTt4d72g/6qNDG8RyQmu20ZCGVbOqLVCQaH+j5WtttlB1gtObKe8u62yzQIgeU
BiumWoW/M4KMbq/Uyg4KLBv72b2e7Yf717lIweG7KJn88QqgKqq+mRvX1/l+CNWEsZPYZBbTVMAE
LWQWdzu3GCedbvisU7fw7mhwUqfKWY+P1csErwFCQ1j4u/aEXbFI32KejfwT2oHy6zjvtkGWVbHo
yMmTvGXIIv0RRk8hfLoYJkTuFkuZanaLRJfXHEYH+GAN6X2Sh6AEuo1Nw+dJGKXQlxrEYIzscWVk
yNon7eHR8XMGiuAZQEfbuWNcmT+1iiVPXQ1xoJiVF1I/pqhec9xi7SpX+2AGnQM/I38ZDxmXLksw
UD59Iian5aFrUxEned6AvWstNcYSYkrPTO2RDpiY5CAULypMwZajOiGCmuvKmZ9kqWmWHMqn29iB
DK2XlV61Rq467RBtqKYAB/lxIs3JueIG/BTKOj+6Cvcl4nISU8PHgCqXmw2y3d/7c3CMQPZZRonT
lFeEaBaVp47nrv0vntZq3bQqmT+HEOezvKYyEOpXVWU7gFVC5YnmDDXEJxdBmTc2051sDhFYXrNe
kaFQFKxZtrjuxjGrB5dDPkq0LGqLpr6FV/9VhOHzgG8V8NFsOzb7VuAFIpOgboJO18xNibqadZBp
ddC8Vir3MEfO+qbGCeVXKxmxOHU83OoH9fZXIzAluRiOubPb/aDsFwhrF/jbNoiNJbTmyzZ4LkAM
tSSy/9bqElOqujkl+GJPvEurX7p/yVzU0wm/0cHR0EKXdcgTF9dD29uESaMpaG80ic4dZw61ryfr
4EyOAq5X9BQ9M443XrY+n3hvJCSro4TQcVbz43mOtI7Yf7AmqZAoNuZDavz617kK/ep+8L/OLcEC
+lEsNZm6hSOEyG4chwVuvO2muNn//W5YdoiqXplU6V/l7kqgKofRtdzEVeWQSPOetWwA2LRBFPpe
uQlH0H6/cpQRMzv8xZ7AmPcTPrsdmRBuUfPTbjOvmnMPlLAUlQEEmvMlzGYCAutwj8b12cJdcdNc
JJN29pZtT4O/5sLyNWPqXvHDjXcUdR5q8UmazwoahUe5+eKa1cb1j0Ti9KDet1hGWMOcCC0Z71A7
hyyi1hWF5HambyC7U4eaL/c9ZlpOYAMfY2uxH+xs+zA5vtvAQNBgDEEecDDdQKvqwTmJak+ioTiv
KkhDg7Cu5PuD+uMlJEaF7miLzxk9anAWZ7xl+yilAZdi8n5VkvjSRmOEFd33dvdCVeLLzzZ5EzKz
QWdIHLw55fudt1IWt6Xtiagl6BmpF3mZYpYrwr+Dbbps+Ddhu8br8RRLov2UCxfI5vZf9KF3uFl2
R6LU/6QXVodA++MIMhGnzYjXDERomnyap0nymDRE2P8bFEEPHh6gkixEXxw3rmZ76esZLB7cJzio
Wi39oQZXO0/p9peuUSIaLetnaH7xzovTJEmiTh90+Te+fo8qI2x8LQ+R6KcxXhTC1jzAd2ZvLf2Z
hlNYOBKsHEp+2tekYsVFHvXj2y+Q+gnWMazXP5JjRNAuQiA/59DREE8i37dw1f+Qv3LwrPy+5nYq
kOPNonw5mzvPpbNy8SimiYRcbFgNc/cVjfNgnVKK5ZlvVYPYh1LAtFNNrQBCSEXzsJb2cFHe9m+G
yuChKeYcrHOsjOIJTISyzzr7YgqrdoE5CXu26ImsL3zLNpmohlXOcfWgZd4mU343dtUx1kzqeVAf
S3DeUHj87GDGXahSW4rz0tsEWpcYLSlDlwsntnMRJk24gvtU93u5+zXcrNVedu88ABzQn6DvMPDK
kHoDqewSMZTyzN2HTyOvSbk3ugpJYPB6XctDNd2dEaqYp7DDNBI3bobb0TBo6nyA2GB8VexAf04F
QJq7sxuQfAhFtgG/499fKjvngioMKq7Y1GgDQX8sNLhw5Zg2kO0/q6+lyOaE3aebRO41FDoK4aam
gugiiudjacjWRf0pcjXQ2F4jKpWBJh2AbGrpNutBO2SVe2JSUk0rcDDuAVVHJZne25Mxjnl24quq
aa64N1dZ/Hw5a5Sth54hoUoGwHZHEtuC3Ry/NiNL9cicGdr+3rcEDW+7y78tWdhrOjIXIeWpIpnV
Vaej4EqDSesl8u+P7N8WQbU9zxamTAa1rEtfnqqdv6nAcKiYqJwahJ/euuVeHBhFN0PVF1uttZbx
WJ6GmS9sv4OWUAqMXY/ygWEkYdktzZujMwy37xJxZSAnu1JsvpC8BYfbLjUR3EWbcz6r4du7dtKX
OPirJNzlPf3siI462nLYeF/1dSny+9vw2mANLKft446jLBKga2hvj8odQI1YSsZn0rdgVARz5rdS
2LAp+Zs2toEAZ6pxXBdP0JQjOdGRqgru3AeJgTGaUDHChcNxgGVz5c28prCbZyK69vXAwSwdHEFk
OXfbLIcw2dygqiI6bf0f0gHk6D6gtaDwj+7nAiZgB3k6ztN2WOuwyMEpg/9KJIil7BNdxwVyB2Bu
dLEMqQZpZNiRJfCDpO1RZfBSW3WZgVxVRIfbOnZWAvt061ZJeGFXidnbbEPaW7JM74mpryeLUK4Z
TEtERKEowqFn7lAGTOAKah59ncDF4JUrkYlZRX6m17At53tWFHNg8cLqFgrAbitfxchczxMRrHeB
SNPw25ZHHekIiADe5Y5hGxdzotPCq22rSkHemdhHKXJ+NMx6f/0q0bnAYz4w4oieUP2q5V2/8fdQ
m7idL/ei6nZwYEgaq79nem2Yz0PM4InGQJHnRcw1lWQDS0Lz9qHkTTgu2wKaaChwQa8DBb0btOHM
G+G8Oc9D4WM5oAqgB2yvtyMQ1HZipugIj1NTDx4gJe9h6nQivEq2iL8fuDEb80QwalCKnnwmSEaw
hx35WfsvQNGQrF/bPz53QI9cvx/V0dg21UP1WElDbowqQn3nLODrLjTNOEIAtzNdZcc3bl5Szwe2
Vx89xbbaXx3cl4Z7zHsi50BN44wZDxx6T+gguN7MKxKNa9RwTEqP7ECunNN7P3JkGlxjfeW/b132
atE8JgcGdCyusJtwn4VLGVvDfRDbFhC4IABTJZadE3iaWJ8NH6f8j3WrZuWNxt36D2BiG3ClqZs7
Xh9ORpyL+OutPr9pT08rW8md509IdOydaM56MwV3I74HZC5uoQhwcMcHIbq28dqN9OW8vVpwn1sr
fHj2HRo2BdDk7k2CKlx8w/0FxQvpJeQYlVtQ7eULy8r136uj75Zv/2qmdjL9DvUMsrFkjPyf5vhZ
wmjmY+YowCfrsIO5iFOddiQvdip7aDv9C4RuA/PVF7/1vtJY4ZJsf4nqpRYqSwHVO+pT1pGMcfko
BjzFAp5h+kuT5Ky63s8pM8s4JlgUrzrpnUznZeG+n4414vMhGbsmJWhqo9Ojw+Dac2jKgdwLXfXQ
TNHfG2iZLFghsel8xF/G2K0ycSQzpuEQR/MlMi0yB6/c9bttl7zOJ+AIMy8AtTTJTgMDlMAgcORl
KkQ/ZxZEGyGcFMxll48Tkw6GL8yr8i7T8thbPccN9MQxgC9N1QJzQ6t6kV4al/2LMIopxKrIhX71
95jYqO1Yf+vp0BYLRZE/SIy3ay9GyzmzGQbC8bDCI1h5nRT4DPEHpvi4408R7NcT/g6eOF3Cyjj/
tD1ViEld8mzkJ1BpA54Q/VdUp3JaFyk4topvpbJdWYzSaOjVnUpFMTn77q9ayI6i2WXTC6SN9M+/
BT8rXRriD9Ibe7YTabYb+K6Wcwv7ClJa0rBPEOg4fvGYSgRD3+Qt1sYH0ZTXEx3NyeiG2/H9riBx
d/C5xHvc5oOqo+i8/rcCvXp+wRKWYzIA/woukUvxOLSeywyazjrfXtMYXJMOwMECOdgbV7FJgfvb
HMD6Gz8GgxsAgoy8qgm1hGUGbQTqyhx7taLTnRwuqaAl1K4a1xu6EtUwTYXDK9t31H62hZaWPEUS
knL8PDLfQYoWw4vJC7BJQaR4gJflPscE6HYFwSadW4xTVOcws708fEftqLGeS70K/VI8QFTMhjDI
gl6QziuXgfZZmS9HDClYHvhd2KnpATDqgUM1V+K+VitTY0cG12Oa9Fj8WnbuMFUg0Tq701cfZ0x3
xqffS4NIKcZXC0nAyxa1uvz2ukSo+93UImSb3aXKtojzHL3dcqm3HNwJa69nb4lDL47waABI9VUl
pFoR4Rob1biU+lF0uvYHvStNuzYJY1IV+ZrdJvJtH2UvLn9kyOGDL1YleQVodRQh+zm1Gm53A+58
zMUlnea1IDziMJ48NqlFOzB0/QQMbdsNntImLkzf4qonmh7gTCyU9cMGOEL08VtjO/4XmZuvvRwB
aIG7uvUx6xvhKV+Hb4S7AgGqrGzUYGfpIgJE9iGyleYNCxwNi9wQsF+afalD5TyLOajW4fB6AZgk
JaDB1aSX7zw+LI3h5WAzkPsxt013ZR6L0LIQfbgCg/zBrcWaZKS9/uF+NSUohBWcDDap5FwPG8Oo
zr/qtpLs4n1ZEIncPj5pWYUMBOt/0tTcBT37+WJbzCB0Jl3kXfe1skPK/NfMwmImJNuqzynmU+J/
GYYrm32hUe8YHT0VWI71shZoU9fYZ/UIF13uGNj5QRfAsrFl4lDTgBTjKhxWvWI0pmnRoV0Mh5G+
Ip/Tl7eDjZuId6uR+rl3lG9DrIIGkGH4YNq4Xb8JbjTRqRi6k43+6oL6EGSCp4dpblMpA/6nIL59
hZmH3SpNyfWs+YrXQXOdHvfQJtNoMHBwQC0BiGsm0B9enwFIlzfuNOMKUb5pbS4jY7TsCsasoiHA
YvX4q2DbUI94kHxU7lNGF5Nwiau1XovqQKfmPBy+cd9O2FstXJvjazYac1vQD8kzYKjGzgSL5H3/
0cPpA27J37Vh7Bhht1anhMI3DOOko+YviOVNNxPcxiDPu7G5DaiZyZ/YLuYriuXShUxsPPP+7qBr
vBv+lh0W6Z7KqiPrE1jtQ9b1hAbCd7M/6vxs7x5M22+88jyIv9UUT4Fj8TljNPe3VSNROT/ARoEU
AMPlBCLrR/16eNzVlnEdJX34DGZ//VTAI8VZqTyMofA+HgCcBwk4p82ePaxrMWzzC5qH5wUgUE4R
m9/L4/COR4d3qhUysD8qlBat6IERA9wysfO/wFiZwvo8ZSoCDskNvAjE/uRBDC+qUfBb7vy9uysl
02dwr0uaiG1oWZ11b3sneGj3zPm9+Wgll+NJsXbdo//YuNgjQ7qwDHaB2pLrBJKKuo743T6AKMoQ
fCOtC6mV2oC1vPOwa9tHpsk8mtUXMLOIKhKs2fVjyWstItH0zuv2Jvye5N2zMgzndImizC0W3pES
ywaV3vtV1r3jXx5WtjgVf5NrbEslpZcCN1aT1lcxPNcSAWchVc7fnALwcA8xnewUChTxfGfr+CHD
J5Fi06sA9yMOQSucpkne4sI1Aay/oBR6u6qbiv9r03vBU9aL8ybmSTkc/Wuq1agymKyHvdEzfjOS
GKLwQrd4vQBD15wdIXw/wc8t6Pg1Gh7yj1vIcFMiYtaAzGWL0cA7n4/mVy7jTwdmRGMS/K3XXfjX
dlUNKZhfbyhLw5ngJger+VzfgaR05Cr77ziizI4jmnyPRqsVQHxx+zq8BVgV69wfSniReYI8Ct7t
BC1K4ek4hlGsfcEHJwM5MmdWvoBdiXfa87pTS7VwMDDg1DMYM1X/+zcRUBMTe42hRrzQvow0hyow
kjzTvo+/jj3VPlkJRWNuzdtin+18vsvLRRb1PRB/huIV8IjLYzA7P2qu5AlWp1GbWGcLyJosQgZS
51oGpLQQN3/aue/nily9dlCK2DASnQpiA8cbMxYc7+nJFunQE2WEM7xQsK3IS7ppM9OhOsuzWs0A
4RG7nGN2QPpJhKJft72OZrZ57idXFsqxMy3641IdwbP5r2ac/YbeSOXMIv8Zl5+eoKHbsCg74iHU
bZnaWofVpvinAv92DtFstpFj3Z74sPeifDpOzvgoVVcCftYoicBaaY1eYRTUddcZVbRsRNxUW5Ew
ukmtutHEgb/pY1BUUSGF+nkMnBIGOUTXTea/a8fHiw42WOgmRloIyjmUjjgEUe5i+iVBpUi1n2eb
y+eSCZJpqah4+34CWzPfugrNdYCduWkjGyNsQ2H1wYgbZGkqUL7Ispd3fEcJpNOA/RARsNKMMPNQ
gzFgFdmiflYOpJka5b3VRiM9Swx1DP37suOprJqyz5VO8khXc7Ufx8dc8Azlotds2/VDll8Bf7ld
+5nARcJ6lYwH38Au75IQg0ZqBUU2WRCmiQDHrK/CXGmAx04VU3BvmHXO72em1ZkExgxG5XSUwWLZ
GEjlea40twGVkK/ZHAd/eVa5qizFH9WHEFP9MqzbiEFnAQXTs5WpC06KuMmfc3P9t074YzHJ1E8i
03+qimw+ZPDXMSabz79pi+Mjn3HuJKj8SAsfrSQbQ0gRiHHP2T6Fe8nkzrNKIVksSm+M11ieQxZX
DJBJXvGU+ChLJBpHh/Tl2s87M7VkF4ZdYHQInp+g3Mn0gRnDQEAHTGJNMuTS/o8jp/xmtSKfIpu+
8hCBSlx8cNrRh+9oHS1qb+AwoN1QxS84ylOWFrIbZyGOO/XBFtlgs2G2jDKJflrnq9NxHnTvTHQq
ZGvqOu2MKaK1dPdhnMJPExmGtg2HsnJjXMx5GCn7+GOKooKRE2KDcLQyTqpfKtZyyZ+ucCc1E1N3
qyP46OWSisxYsEZH6CZc7DucUUZRbw/BV8MjzW/7YxJA+b8gJR+/uKYwlOYivhrbO1kjdA0xPjO2
mc+KQbCF2H/JxVSlUdvH17Shj6RWVZcLS+LTr6M6lYALw5y7JFVpFlbOVPTa4Z+2P9g8gaRgh2fU
r7ms0EgwDq7o4lsVr+7ASCyT4VmakbC4fSeVlcmzw2inLvUDhUYOSEvfTlrTUOM/BdiL70PHeTQc
qKhDqM1po5eUKcV9KAiIsS8wBtQN8FlOzQaTDd3R5viyHeoHf6OYahMrdXfcWWaRc/1eLLJ3t7Wp
VRVPsPuXn4Kd6igHXJLTLOgqe87jocxt3okO0Q/pCvIo4xtxluBfPuYe6vDQsIWOorpYiETdKRzM
aTlhul10LzmnPTVNZGObTmWUVEYINnWu0CXHeJbKy7HK8kK4cJ31rQtXTcFO3LjBGP08UhTQ7eXr
GscZOp83C2MtGQC2K/740VaaB3MaDu3rZFNygNEpjmsy/nCQoDFzAk8VJj9MhDx06IdJX1CrhfKf
J4BBQxMr2u7Qp+qRm2d1PTv5oRDWLtSM2CBb2uhZibIIYyu4AFC1JP2cqNClnQPTdjWb4qsVQeVv
xbGmlJVMfwwfS2rHBlBZljXAS7GgdGZhZpmOqBFde5bsGBAx866DJru7wQI08qiamJIl7jql9iKu
grIsZwWSCLT5YAQdjznz6Q/Wf5Ue719RI/aarNFeMd2IiZU1Km+poTjolrvGsNTQs3zH53Aof4H5
LepoZA2mNtllh6ifYFI4qtkRys1e27H9UzvVhhUD2Vuf8U61C3PxqJF/kEiVYqvUdMSy/wRn0W2X
qagfa4RwE7QcBuBfsVG9Q1SvOHIpA2y3ZKr/kq8cev53piancmLHtDMObR2MeeSXGv9eL6M68Nwh
Tbdzqir0K2+KFrBMNcrEvTm4VCOQ44QJM2uuZCbTt710Zbk3KoXpMsT19MrjV9ZwUClZ7g/Ehj9N
hodA9d95OqxbzGnUR+ql48B86H+SEm+NryPryPu6BHDM0O/d/LkCQVxEUNw18vpEDR7hKL+SO9/O
8WjtICVv8nq9ryzuH4yiCvHOps5oobTIHx5LZiWvt1trnZQQwfFQM6+V7oyHIzM42TLd7COnPs9s
eiLJGBasZsscDe/lTphiKENWFQoyeEuRbqxkhen/TZyLGhYMvQMTr39A37GAmeqABAT3+XeKYcNg
f0peR/7CsefMbwFga9F6U0byMTlRnCV1KKQeA722tnf1vQNaE11CRABnH1ofnOUVl5yqAkHD6ble
Zr+Um1GuHnSfaFpR57WKWJKy2P7io8dFbzqrMNVODhSYRgjvozzyWpw6QKSytsLwbrmFVuBV3oVb
6MFe01wLpK6YMa4C8G72047XSq7mLGDTp4qnOKL0cHfM/dgjEbL1l8buwUm4yG84rlL7SE8JV0o3
QyaFXufzvlbmBf86fb2VgAwnetHlif4pnWpDW5idumP65AZv62UWclgigOP9IF+/8iZfya242OGi
alnVIn5AhZ3UujX6CIRZNDpBL0dZGBbVsLBBqJUrsEK2MBhbuuismPYL+Y976zBRYHQ+kO87jX1i
B5hFWjEL8uSI5OBYbaQu5r13mZM2qbhDM6LOAjORADPbL67re36w4landN4gBqyX0Mwz94YSAIso
3detSBPY4hDgOaiSCG9w/FePoo9OvfbrCRqcVidJ59QfYOO1xBqOk1eGBSi133TgWRT4c71H5bu8
SSUgvuNvybKo7uJLrKlymbI0mABlSWYA8uA8sN1Az6IRnGBVXt1G0v1plVMKXGPE1Sf+kfrDd2P2
OiJmAgP4ZM2GBgbA6KTE6P3TzJU4LDVXyPXVkMQkfEtxciuewtj+nwzP+LF7RVUo6lndg7ikent0
XWA/xnxqlycY1S8OM2d5j8AvFUoCMfpDf1bgoz2kmFXw3gyD/+FqNVJtB+F4FJ/dl7O/U5yPZazB
7Q9QB3oHkY80smbTZpWxpeDv7lCzfLVK3eyzLEBhiOwMPgtIKzYBi8pM8VC5nOd1cPpA80oLu/2w
vhWYksdXg+o3nGF/327Ema6OcgnAhJyxyk/jCM7M9zpEjJN+6scFjZKG0/guFfkbnZhJeNUe95cy
kwDZo8ezCKC8mT4VstAvD0uqZYyqTscnmQ5GD1VLBYkqxI5jmNmMs79+yFh2INUNSQG+O4qR8lLj
yjq3VSaNZ2MHro9S1hFJsN/E3oOZ8mG0K92RnME3dhpjt8rQxbkTKnjmI85QX31SBrs/dNkRwBQf
2yNd2tmF3MUvKN+gcdl4/xuBASsSDwZVTedoNiueSS1IqES3cpIR1dVtTYcQb7b3ATQrOicNqqPl
8OZc24mLwvw1SclMjf1bSV7GnOXNyS02ICdBApEbipFVedPNkQ6ezSfrQmK2oziplHV82mgnmPU+
2mc994D/vVcbndbaX8iG3Kx25JqPS11dKeyeU+XmbCAUYvE89gPwh9txSSF/k3f94Xi369MxkPXI
x1dEd64X5mDtwgSmBDlceLAOEhcLmPBpK4O3EE13JQwm6RPGylll0bmGxAm5NDVOaFj8XlyeMQbE
bEbZy92yNI5fSLiV1ePMfuoDjg4TfbK9SWfn7BGxdGJw7VbgjswVWeM258r2twf4Q+kJDzWzW/eU
BumD+Mx5saocLxPTIN0s/T7PMa4v+oLCbVWDzQKRg/zJYia94vgXwWJFQPOX+VYG9vBga6bB2EnD
hChIWxWhHMa3RAjJuiW9rhFpMLEbNYrZM5anqWPDAuD7vQ6OMLyuq8UQ+aHyanQiyvcEPJrOdjzE
rhzuXElyDxht2t3xKC4A+Bc5Sn7fkOlzCDvvflkTlNheGlsXlVYSJ7ng2R7vNT7sIGbQa1opynKD
GUX17WlT5zdTaPdTVFsD3nzSYdcbHBpgifcbDskE+MDNAavSM09TLRuj2GPS2L0dFvCJWaIbttts
5d2HshLg5IC2YwLS1ci8fU5TcuQJAcEzKqWEmQhpE3+gq9o12HxmTb/wwCliesuHd4hcDz2n5BDq
nq+p9JVN+4q8fkC2h93BdtCAK6AWizImR+6bv26j7B/jB4Y8727ym4J4vQNrhgV3PjBjy6E6pFko
ZQ9/SeXKiSmzK+l1i0t2b2RqEo3EQhmIZOEjmkSDYhbvnnYAArXnQgD13Pk9xBYIPPmaANM/mw4S
lEBQVmEaksH5ezza96AMkDjpemrPe2wuQMV32JtYrlsB5+YpdrxdZmtyMl76XaRReQnaHxuNZQR0
l0enZXLOmcm+0CPjX2pmqGsoOgKD1wJiss/oDrywjrlnVLbTwOsbM5/6OpO7YreKR01MCXyyHmoP
2seR834wBUoXzk40MAN8o/u/jHaaU5b0rXzUJdwtjlAYPC4QJjkFLoS6UI/gpLRHd3Htp1NogVgr
pHvpdDn9OLlOJ0Q2kXVBaQ9pM3uLKvbBkjTx2IFcNx2wCv9ymkyx89746sRYy5xsS2yp1acl4O/v
LOEjBWeZSnArWvN5NmQZ+bD0i3O2cR2yJtnVUVEMgAyz6vY5diuMDPcbzHgz/Rpj56tfufaD8hj0
JsK2FgMF7J3OK4poOnoC+7HMqj5m2ffZj2Xf/EF36Ak1+bN9+ocXA+ERk8JCBr6hCQhuMqVMOI1o
VcfNl/No01SLbXibfhKO6fiUhxu5AtcMtNgMc+BoZKONpGEdP5yO93GBZiLEG+ly7tXXyOoBMZme
NgI3Z9e10xCuhmJRm6Sv63O6ToRtapm1RquJHnK45GLQsScv0Wb6enJZ8mMlbk6IM9YO7a8VTuFn
cViLiQolJ/XpngMBUGRd1VOqabAgozh2RvWAaLt6uOxKH5rqBMs/ngqW1SUhH1KvQ2bKZfBFy7o/
p1crCVvRw7lo6DHd9TJrs3oGv3udk1WaY23SK4Tw7q2qhHhriQwHLwmDjZdDMd7oqgBIj2Uz1KO5
FWdDY8CDKM6ObXzftiPddrorbbPzonhwP2hZefTQSFiHbXjRUAGJ8NlEV2vKC2T01JgnAogW21KD
qcHXlB4lc8JoEp4PKl/qH+Bdl3yWk9g1V5XX4wIBRRyDsDHymzs4jFWjx+2FYAh3tu1fs8pfGsqf
u7A46+0wLd8mQj8iGc5ntZ3HEEeN8oSSWeCw+qjPcvSM7T7oRi2ICKSAVJiAcbE1kVmof4va09ga
21RFx1yjw5RKYqtlSNJsuRo/Ul/9ZZ6UdCjtI442OAHlot5zv+XSq1NfcvXY5+kWzl3pysVsPZvF
LaZMZbvnTSPDtMTGoHGBHFhy3858JgukAjD7xnEb5rFNkhlG56vGCSj4ANPFHIEUiBPm77dJz9E+
P8w2drR7OAt2yUpZaV5RT86etuWR0bj1lkUzUEdsM6vfiAxXN5dJy5tzA1pwt4BfUgS1AWE06X1U
fc4HLKbpKJLE8TfJfEKfqCmwVHiBqgnV/gMo7aVNXonObjODiIuD67klhGGF/fF3A1kBqDLC8mwG
K8/nwMZGjWsMW6mKuYWtzsysT210e1rpcMD1n7dG4pTHdzsSBlthdDMO5Bjp+PPHogIofwk3xVTM
c5lUDjzYodwIsaIbBwskxtx/d2rOoKUhAKoWwhFnw/TyWGD43PcTU6nVMWvYaAfRa0HVpSz1OktG
BJEXhGSaDD3L5EP3wvfXnTZy+gZtWFw0E5bL/XF3cEeYcyDgWGv0Cnd6n+4eqOwPJyejgPngy/MV
QWl3C3/J2Fm8IwTUN6kstbnED7gI8mX2PmRjCiZ6kL0mXlql7QQiGTo1/gL9Pn3Atelv5Bjwq+4I
Ea2aXIlKse748s4+eDXUz5EOJnToqmSDql+x1o0BFSC5V5wV53yV4dgLTaYsmMA8oy5Dmu9slWfy
ZP+LnJu6WeyDqERNOZY6aCBohnpRrGLv0aDqKCe7l0qZTHNC/Md4/7JcgRPRcZ4+2kuEqk97l7vo
qsp7glTOkLDOIu5W1OHo+l8z9yg/KvpH9kF896JAobtx2LlJWgLbdo4bYXyAxabhT1MyhHSnrqFu
MkUNEe7G7bXa8kWoaIn+rSRz77R2KtxussRfT0yUujlQCkWKvpoxmncUCD/R1iGXMV/ljrwEp5PN
2K7/A+yWCIrr75Lw8aSH1/nSmRrVg3wO9/i5Qum0brvuq7gkGgM6eUwAb3KJdwGlmsZgHb19r+0/
QBXWlSnKmZq6iaiAB7HUGAbLk9et4V1Tmi6rd9RLQ4e+2w8sagXy3We6Vrs87IHjY3b5RduEt8mT
U3i/ZR0WbTeiL1sKDTH/rYLwTklrY3rKaPxjMvkHZle+qWU187x117SI8QynQ9euvGUEd32P4oZB
Lc8dAWUQNUqSlews1iNY/YZobp2E/HMmMn4to1WR0GAiHNIdka+WuJjWPBJ36jRUw3i73cqZjfUW
+27FfQ86lEUKln9Tv4nvVBBBNxwtSDO/r1iNx2kveJT0A8V4+CW9EgzeA4IXJe/qrkLuHxex1GMr
l1odlH6seYIYBRoqHGL/zmgOtOKd/5bV4SfXTVaPWmMk4QwYoi8QG6rf67tqWwwrAkx1vaeIJYws
gQRtIQrBZGzxM02kRuAE9pa+SUSvAB2Zbs6Qpx4/HtZIh7936lpRYlgXh4bDGxKbAekGwPVOSagl
QB5NW9AwivQzx5/ophQT+Pno8eYYINg0k2O7C+LGcfkLtaB+Jf3wP97ZWiicNG4VPNlkxdRnj3j7
X2pn3klq0BJVDvIi8WllR+QxTkvCzVfaOqScqA8zQr9PnkQ7BPVHbDy4o/216yVJ6OFIb3N9JRHD
qpB4rYKdODDC08fkzoWD0q8pFIKQZL0a+Vl9QPmoMldSRMdtnlExXpTT9ME2QI02xU/TSZPnFAsC
U41PIe5+M2wQBuqWyRHhwFpPlLlfd221ZAXu/GUtQZGXqTAPuBbXXxW4/m0EvHJjd/JI/l+Wh3iy
gTUUe25jG4bAhCV6S2eucCKuKY7zoEAgf0QVUFK7S6EFAHDgjHGBe+7xzQ3J+JIVm4uaz3FYKUGr
Nr1TvH4lFYayFC8TxkcXwv2qGYWAZyDPWmUW9e0E4ARyrTzzs25Nbk04uFAhEJo6bUBx1MVatt8+
ReofwLzBHlljftCAnxYgvoabI9T4h/m8Bk5vKhuyDpbXnKF5e5Z1KpJx7lPveYker7+6mF+00RGV
OBn7BC6zVuCblyLwrXVAHvRRIOpJsu1qB4wDfPZyn+aUFzPptRLMDulmFzWXbvX7if1kgpv72yCP
sUjpguoxB/9Vdu0V5QTj94UZtF08LmZxZYRS2SGWLgA9t8jpwLhn8y0iNJkMMutoRej4HWkJy652
W+WXK1BhnDdUoCP2xMbBYQhirFYHM4suZGzw5Nh2AufPmdnVEav8IVzVKre2F3ltDWvMChWH9SpB
TS5Md1nH0bRaqY/nl7E6OIvnyoKsWpcHWo89vfcAV+aZ3vmwyMqYfevMr1/ujnGXETbh0cqohq89
tGwoSSUEWKWzf6Lzo6s1Qv4yqk9+cv/RAcrn3ZGXTwOexU59KuKh6bzlGjerfeqOTlu0zDz5Gi3Z
5EOWRIWJb5i6Z5/QZftObKP5TqiiNw354VmOrVq3Nwszqm/98CvHYeI7D+0G6XOtFjkznaSPpNEV
4+qvl7mkmOT3eJxPoouBbLbIK7i1DYVSUZ+NfA6N76j7cmYccxceq0QbJoOxp+okUMhXaPnie5ow
IKDOdKmhgmwFdiXf2wdwW5FTNY79Xioef8/xWjJ4KTDsTNVViHmmCaUWUp/p9GW8jtddNXV4ZuL6
IxmYnYVdOCbd5njF57KsTDQb4dHQ6DHID/uXtikZ4ibkF7Y4ZhViyTJl3q5+ZfXi7d3GAN/nCuFb
a1xMXV0cbTSAe3Wmi+q2b6HySLz4Et/yQtzXoDiqYRvZqnYsW7nbP63BXg827vD9h8BenGlq7nl9
WSNpiXUjWtL0JGqZ5jUUMP/+lAS089E+WCYpFt2bHQ2WcMcG63duujsvh1SSKhrNd1YELqwGf9j4
cWtdHyCw34vhde+QPEqLoljlqZ7xAFv24jeZtOSFizTccFW462FPp+dDaKpUFD1OyvyV6WuKA3qJ
a8ENBtlu2dH8LL1nwbCEYMZXTB+JIHmZdOZSoR3RZO9fIvf16NpswpqOyulHwYAiPvU3pVRp0yrs
kwkQhlhD725vdR4lZTVIoi2KDa9xhBIO1L1rEnKDeDZuz9FsgWqhNcPmAPhxCVBXKBkZ5ljbNIv4
gPmKI3OBLUtXDCVX3lP2PKp2qoLV6pBORKTlFQAENNhXp8EWLYiyBpOnPMHL59DBbj4Wzaf7z6Fq
3fhk7j5yaz6SxK126k3IgC1iOG/797/XidMo0F26hcWzupDjgPTSajH8ZJvyrrY4bY8Jby2IXEgE
MJ2cJffHby6kPb76ucYLnNFmzBK1GsshVDuBeuhtxYg/EzRWvPDI3O/lAZFmz6FVrFRcbyc6219W
+xiZ2ldyPM2vycHd7WwV+gvyKkSZT/OvVYpMdq22MK8ArL0yHWdCKha51MyAo/IzkgaxmEXIS1Lz
zynInZ+6vAHj9te85NDnYhk+xyU0BCAOWKKsrA/yKSBJmVS3GF15rgJ/5im6bf85BOKojixK0JGL
iuxBuD4JvdABwFeV/z7e70gXJqbS46FFUudpgNNJXLcjhMTs7hr19SEAS8Z7zngHTk5oKRjG6VCW
hKLkxCRIeH7HhKvLQ991ZpQFbWxqZVQ6yZ92YcIgdn7mkuF/tW+NGRcetmNF3zRnioWIXWdZe8sq
Dq55a78CO0kvSI9lWMP+ok4Bc+lnEKEAdPRBD1Va+mBHJ5IUHosDQ+XbXN+vnRon42VGUFDzsB65
fHnmyI7NAW/1fQu3qiEurKQdm0FKDC/Cj/ZtfRPmm3DkHHZCYV8wykOAnJ8sHBlS6vTKhpPJNm8y
s9uoljBa2cwGbZ0aHJz4Mmj6rGLMMM9z9CFFxs8ZaeHjQUT+RZNjIPhrgpnKJ3qZhW3ohgVYsQsF
7ZGvJGNLunljrZwDVeqvXt3rtzU2g/aMVfdRK1SyyEP6d/Yj38uOM1TOmHbOY52vUpKOCzGYemAv
EpLkXGj6xHUkf6YEFBwQo1vrfDyZvtM3dgUpqOL0IECgSR40k73U9gt5laGif9yiCdMtAnffO1AR
+iXFTLa6+sLCpTBPMGpL0FRz/xazc/nhDfZuYMNxJq+eoO5w2W+EiB7c2OFAGREkSgovucM7VJCu
nXKzrFFEZM2KbiELLUqIMtk2XPFu75Pcabkm2exArfTOCu2n4q+MvC8zoDIH05/+f2kxS+T6gTU5
s0w8Z0By0X/UIRaLzOe4cSrfjYuyX3/1OFGsVfMaTw0/RAoofxbMn3QSXLE+AmzR0iH/qrO5HAt+
DeqGOU27Q4fWXhB5AzOFo5tdyq7RnjmzLibaXPyPqThTTVkDVwCHz5C4XLYGKeTCEPzO241VbGs3
i1fD/ZCtj9utSGEemdg1Agh7lSgR6RkwDH5FGqivWRQ0k6o0kfS5qnDK8sD32yJ0FdRRainEDUYP
jiiW1oO3lWDQFOQVfVnk1IW+0oFYLPl8ldoiW7e7Q3VLfWgePz5pU8HUs3xwiAF8aAk9rdRC19u+
W/pgtnEbeMJcDmgogvKyM5qI04MdycUxOP7VFJBJAuJwJM4wa6mUSkhL0QLWCId3gi/VYTZRmxfb
fjm/ZhkcGMK9QIDhHv+lIgX49FWzBGtEACP780y6VjeU4jh6eJu2ZBasbQGrbvNiR5gs27uGDdY9
esMw/Au4KZUnLmTcY7C/6eromLLCJdEIZUd+BKbxno43jbYImGZ/NIuS5ka3RAl3ZrYgj6F22WXP
EEGBREuP486pfAkRkfM+ut0ER4omHpQht5uSetWt3EkTTxwP4Cuzws10Ge/ay+gPczp85H/TSlgD
l4fVET1kLVA6Vw6bIw9oUOXjQTyvryc9GQdnIHSQEQ8yX/lBPWRi8ULYZpQUYaEFeRkCq9eYjd5X
57KjO5kpBVeaefAPp2BMOmYg9FpIajFM6hrsvipT/ZOJlrrloYvRof4ZmQSvyjFWdvkNLg4Yibat
TPEyhWElrxlK7hxwuC2BVAJaxwiEVI2Aht6cncXUFQQmX364BnKLz6Py2pKLMfjBPVMink5C5K14
mhiFFGpsvNedtYZ8uI4K17mEE/lzeWtUBv0NnhwFnnCzjHsMeG4QsUtzkwRZ8RxQ8x6aLlPYO6o8
4HkCzblQ4lmh1lt5jJ+syumq8vMuDv/3Xxpo39AUsjkEsvGVhOBcLW3e+CcYBWavicUbnG9ftJNB
8baksE9TtKLAQWg+o5alFKcSSN2d8iRKv8WKyBtVutgZa4Qaadk9qhCYWktYS2qkoFSJRh+UIevL
arw6YJeDRlSitGF223WwuOwUnnzoZk1bmP71324B4qthjHzmXl5z4KrkNwuKz+1ot69BfX+7EErW
XKP4tqZ4cPKib+iJdsoSidB3iQ+JqMPkTBiXWkqUmd2bV4SC0m6R4xIzTsb2kqWZHvszOtr+bDBt
fl9/1pbTOyRdAuXIANfBspormmhqs2sPD/B+ndwpIV9LSgEENoi5niU0xpulLfHdU6jhZCWGSJpJ
RjTid9tAhfsWGrtw5tBnKH78FgU1zMf+fRwnyd3xFTQhr1uRI/WgVXPyH0prRtoqOsJ62oQc1Hnt
ZthS5GZxFAHUbNssAFmuq6xTuhiJY6l9JnYMF43b6NGE6z45OrGP1Xg1JfnyWzdAL4MwfL7c3mL5
twE3xPE5UjgSQ0vwcWelo2regoNbk/XaDqrcAjSJd6EQyySg14Xwj4Cnl+Op8sO2MIhL1oCoqb2V
DdjJQkA4Q3xt1y29Sdli2ZA6Si+nN2hckIX6u1EsmcHW3BKD0QccZF5sw2l42XWGGavWcIdXfy+3
fD+6kPWRN2a3HU9vUz7j9PxR44AmKRX/ZZQVvU7fdTfMi/i91mC9fKddAJ4fBxvmcevSxo2/IokD
k5lmB4WUZwIg7TEXD344uJBI+xQIfSC5f7ggCeqjOrYSKfs/krV9Y1zicMGa+hmHCAGj63DJi9NP
H5nuU5cae75twLGuNYOCE1mI9v5jAJpiT0UVVMZej1wAAAX3rd8dJ6zl/coMvo5MDnLbk62Pl52p
QlOJKY0cXdHZeFIsxk0YwaUrv7trS28UdAuXV4MOVg4M36BDhxUergYEI7He335mAOvMnxLfrXJB
ARP66xIzdy9l7VJGN0rtRQvL8fI9ZBEy0Zy7pGjp32qrBs837eVuelTbSRmARcFiG3FTyfbbIVSN
iBo+L+jVSLuSKr+NeEfM4W7ORMYevVLrsTxNVf5WR8gGFLe9J2U6XkgUnUhZbuvUMr/y7iDqsA4l
S9dX1ppzu8syIonED3NqFHLOCjQj/4wvJGFhIGF1qipF2xBOnCMNNaROSnO296TXXb23XEylE/Zh
XtEd2iyYODAPHbe4ft2QiiB1RJBmU8Qq0pb8+HWlJ01TPhH5UF9OiukFwiFfjremMa8KR3qQ7qDl
d9n1YaPumlRaB9fbF9ZO9K2dfCzCXE7WqYE7zpNFhycuzOzX23vy1XU6pKdBB0rErdvc543j9KRq
6YwHjUIdIiFN3Qotm9sohyV6ZseJxz2ZF9fuD9kYx0hLOUJWd0gBfKoufue9g6I/TvxPhdA5+hkk
WfgQNDnbuc13tMtP5oJbGKLfty6tyZtFmUMRfzMuFVF5+JyylzoAtUrqsu6Igeed/1ONVg8MTSca
alvME58Ml88ZWohSF9ohFSXZ74L+5YfZmg0rclvq7iOgCuK4nUkNsPT0pfMjwnInmUqm4xzXAt6p
CTBKdnBBoDfAzzrTFQhXCs5K0I+AIVduT1aKD5RgomEbJ1iSu2k+f9fL7O7qX0eqWC9ppEge3gBS
qt557nT4opnRDICeJp1gcHxp2k7EtsGlrYJeEimJh0Zytf9wdXdQhhWHozbL1YaFH9MuFhr1ge/B
u2ZTYzz+4IKwOLaa1TxGK/bcszmf73eCa+w5KIBu6qIR4l0Luy4P1ZnroN4CpI9KcRQIq4MrcdPf
8uHjLQeJTzCQql9JzEbd7ZfqXp92jt4cthNp/6pc/QMhsJreBnutKhz4ENzaOiF9SR89qBBy8qD2
G2xzTm+O7Kofl0GvcjmxyQXH3gxn+/YgiOM3npVkKJCDGflfD/beaHwI0Yqw4hW5ZaML1z9rs6O8
uOfOU41CATdGuQNOfHSELTWVpVfcesNIH/8RLsR9Tb7zbF0+FuVKngXc0k3ynpV0fDfM0wna6ZAz
/iRCXXbz/8sEocJfDwqguKABEAIVVTnAl9AlK9Ka+4N1wRFENAQ5GJSk3W/Ae/VlEM+pPad4Dusl
NUUVz2/gekow5Yso8dEc4BK3jNXZdZTwLXDw4LdwBUP6rlzinDXka8xWbDREyxkf56TKiiwakzCd
YPxkdTJpkkE9zmQh4wS8sx9CxDOguIIpJlFViGe4xxwSk+UVsDcUqvrErLnSYKKwpSL1+Lg7D3Mp
D8Bq1AmyS/h9QzSI0omT5AlGkL5T4F2aEGEzZ/mno7dHhuoO+3SVBzhrngjsQSv9TGtsYolIrOLP
3b879/Ps5ljmbc8l+3wODJzAFYpivLOxAkn4tYTT/onBIlKVbBnBDwxANNHb56Lq/YCCow4gKpT1
8KCPVXAag0fkdgojxAXwO0Bp+YWGFWCqVdIVD3IUPH+PaqsmyEp7DHvarFFlgIrvTdUgH+d/Ie7F
xfX9SZq5RBZrr/YQgTu2L5W1KMRJfqnezEsS7OBqOfq5M7kuSYPDLmPC/wZTS4ZbfKf1zAww2LO2
qHqUVgewvnpWbLlupjOKFsyJXue/30tfsqfushGa1E/xY09AwHgEXYeXGqvrsEh093Xf3do0AtaD
1PV9jRMuE0l7uFqjhW8Dtt8v56E1wmrz5EmX3m1omWZTpGrhYaNVUuzwaLq60hpMNRR8TcLfzTNB
6tB9ZNwViHlLj8Ayi+Nwen6HN0qPannXLq1v5wHdxO/VfxoKqCb/C04aNbo+YxRhrsK77HjPAOTx
4YwYgDADQS21h6dw9FtrXj+WSVYrHeXakwbE27BoOwq+c0qxWnCYxqLw15iQlql9VsYoN4YMMqDW
YNkfMFNYzRGo0r4U1ImzQl4jOe5evAxWIahKx9lAlwv4KeV2T0rith69Xi52X9digH+DTs4vr8Dv
2m6jTX9TyLmQ8JKEzO15fd6gc8JSJ3iXhxaRBb094v0ojf4d3auSQmDEFGbGRVAy4YsMYQtjkyXF
QIxGCkPNymAWyZr7mcOftgow45i4IcA18/yQzg4SJGpi2ooz4XYTTz4LJ6etXuhx9HENdvmVVwWS
4oMKh8Oah86Vmz/yfLZENA1f7YBd9mlMsCpPiLUjOrSYpiBmWWYzPim1a6intnyqm5ULP13cws6r
pLR7AX604HAtkTRq7czgpE2XXORQO8+/bVdy9yD6gFl7aJPihK6oD7swo6lEst08JJf89V+/X/TE
XVZ/Tc+UJaGb3hHIFIcXL1XxG9dL+itAe01qDXL4hZVKa0Sv/N/3GEOFJL/4vlskUCTUxn0JClYv
GrlIsyKl3SZ9QO8M/j1MIwY2ijAvxYaLvinoT0zsmfmt1+wv+PBxPMDjyQQb7+99P5IDxx6Uv2zL
mJc0K3hErqrNux4b9qwiTBuQMcl2wPwD6+WYKZIkXCFgrsES49yK4mgZrWXqfTw9IVTqCxvLdWCa
1pqLls6aipzx1086TDlHM65fBmRxyPmFhSXWpnFXIGGfsyrBUTfW7mvIeCS+fthMSMYvOOsiXpPn
IQVEXvdVBtshLRM5ELclZ6ErCcQ2RzL0TQoUuzq50csQA2HsJkFMsQDyiQy7JVgswkBnYz0HTCh2
rLv0rjkIe+0I1gO9Mx6AGOXDN3WGvwJZFVdoE5Qbin2tbXMu01jpoZ34Whv3LbnO73zMUJxFap6O
0tAiXki6SZS9hcBzDcEvHAwRaBSChbJ/XQBP8mkMj43qjCrjldSJqLVj4PfSLNlL+IWMdoFFdANr
YCviNATNUvaTo6Yl68UEv48qFmPUllS2Kpku/7hA0JVcOKXHlfoJpa/ts9kSPlrE2JRXqCAh6C+9
yqrKTQ9JU+8BrA4ZZXqlj0F/13Rwg4fnYnxfoibvuK/EoMoc6G3SdOnV7O4YzzOqb9tcEFdUeH3j
/uoKaPQn9z95sGIk4vuJWm6lVVUGXDeEJLrOz4tPyA1c+UbChjjI1xOZr0g34dY8NSR9VrzFIh+g
f5OG7Lsfye0OWpYLmmDd6i6LoGPrZxsuyemPnHmG1iPYJ4gXrNK56Ti2qtRdKQ+eHLNJUC9jCQcL
hnj+Kg8lp4rGlpMqmYBcN48qxS/Mrh6sEyNC0oy5zF0lRnes6HCI/oAWRq2HuEUs5K4YUlZ8Riyz
IKzQYV38VefDObPbUzs4zboGftDcSAo+0PF8eZWpknY9eG2PVM1jdUxO0HYPTfkqaYXBuJlBXhkO
ilMqYG+tUIQv6tTVBdnU1WumOO4oxGzmy9Y8pL6afBYte9c6QuuM9bEMO3PObaZMfXlSg9bukDLG
IYJsJvlHWveMeHhwkJchQmPO9FnZm1hdQWwkSY9Rqbav1DJsxSpByEhw+5/dTB6SozIMRFk2/O1k
JTqNmzCVAsgwJzff9ff6r2ltaYdmGOITSHJZT3//4pZxFJ6dhwrjrWM8KkSOz0O6AJGT3AMg2tKN
IvLp93SjdX4jFdejQ17R/XJzcjZTO272hR6R9VEFMs7YGbbpX9zdnYOgNzUcOWOaE330REFW3/CD
n3vMgqNQkM3Yf0XqID2in2qji5TF/Zm4pIvdHhBXZDbMrCMVpy8oZNe+Ah+ManTOgjYMqTig8Hnr
MG3tmxN3P8ZxXr7PFH/tYMwS7wlcCh5wPHfOxBgUan8BvFZkaAz+c3lm120EEieaf2pinozk+8pG
g+63XSZ91H3M4HIJfhR8MuUQZbfKZIH7zRDOcHHigzotUN1M1dnHNcjR/RihiUNQejaSklMer+8h
hHUF3QlfurbeEgdODFAaSpn50tDT00JY58lLPn/8THgL0xppORWd7/Tqy6wl4Wb/5Q1Jb65NMvLl
MA27uRA3C+r/xbo71wqc3roRNgEbXUAcFl8TQiIYKuuHFm/76/WQbYTKtEFZw/Mj8PDY3KMKSpSQ
CBnod1tAFO8Lx67eDyNcVxjZypwMry4UvAb/uHq/NiREI9a4ZPQSCEGWB99SV4id41RinvqUA+r5
J3e76JAezgkv2AOZCXwaU/KqTldd7U9GtOKU69nkO/L/zlZNhikidWQgG/yPPykjvUpvDdeA582h
91L1tWVGiHl3zE2VWlZxq/4ceLUuPCCtxbUDPJ1YG7MQTohEjGe3LFZeWEXlh0WZ7NyD3whJZYuh
cy+dnAjcpXyTbP70GYZIRi8A8LaoLLZLEwF3SChqMhBgKSHjLHspzm61fHRH/mFW0BcKCx0+o1Uv
L+/z1/7tgWTXyVIq2AmRbkC+DBDUZUUlKISk9pGaHYzAOEEjyO9lWTlJSvLGRQk2Wn14VN4NNobw
QlNa6kkOG5k5KU8LhjfWf8E+/m9Vhc+1Z2o0blcMEaMXzFfsxhuNUHyps4INhZ/d1kQscwxA2XWs
yWuoxUToP1+U/JjDY8X+GjcDb3RWw7CaBllbzpa4UwqVA7a2gIDe3oCqsUjkp531HT48ymSIjWLu
j09nvEFQyHkjeckdWa5kkYv0/5OMt5MEy36rFfg0+rb2Ql/IfzSV+IzT8xImEBPd/nvYzYjnnvtg
mhz+Wt1hv7bsmsUEcVbI3BRlqaEMnkG87tIhDnP/vuXLfj4MtEWgHMwxiJFHSmTJWfL7dunyt4ub
DaePfgX7qVK5bqJ2ZjIGMdZd29riecUTnsSUaKKdgKJNgsEGOs5feRH8BJ1aD/flPZombwE9uY5d
iFI0yNCHaOvCXUyx9wTnLpiKZpErfpzmObVff/EZwUvY1laxJHgDsS9RzlotFI5NDAMGKso5TZ/a
rlq0zP9a4FqK8S0gwxkxbfKGlPy0oXtSxkUg2wlFlqYCTApk2QBX2xQVywKUl6rnBCFab+v0C+Sr
KLy5cpV4sKchE3FVd1UR5AZbSYboDfFIq6IlQ0eBp5b875rM3R9mKs00ho34XDeDtf/tSEPFQDnh
8sDaKpevNAJ0+fHjh7SCx1qJbc94l+tmVrvdWHsh2DsJMykgQwHiZ/XkB1cKlabckL8YZ6wQ5HMR
DnHCEjse9O8c/OcOg/edUjWMyJAOc1o0z//eCMo1/2O6wcroUGvidlQskpqa3OzEPh0feiYFuNKT
e4UR/dxWASl1DCmRsB+K9iF2f96i/hvf72L7UXDxq7QxmXd5JlkrLcwFJ1k9gLoG/qK03BkbXnRM
O4eAOXI8eD1tk+x6JOuhFd6XHunoFen3QzPm+SRHK/qi224NMdswxhNlj9cSyLvIEUbgr3/pgIhp
pwP8YriKEglIL9QC/42j5IlrmdH3l492suBHrwN2C4D9Yy8T1nS793UA5Utc+yNAdYkhXgYs9Lte
CkUuaGu5s+JAYm/OlGc5Euraadv5ICH7ThPVCesdHeL5kN3amuhhYAPpGgoEEBxoMz20kWP+yN9Q
a/oFAGc5ni0YtVLu4Od/mL1VLQWG0Kyt6crWmr/4J57Yiu5UGcL/74kNLyZbn02eobRMp/cHOAAn
aFbZyX5rD//kdSSCTZMZtdp2XYUZlUGl3TgUuIqeQhvmNvgCUE1DoqfyiFOQlJgzOOIJlS0crNOU
RqQ/IDTOpTve3yW0HwywqNrsKUY+oqH7ADFmLwE7Vi5ZGBh52BDf1m8YOC5pOCwQXdktnH9HbiS/
qluwXu7LYQawnHb8Ib7LRid6lFuBjv4ZSaHs+LTAh7J3+H44z71bJ7W05d9oehEEByGYaZyJPf0Y
2PtL3cSuzItvz0AtNNgCi61r0JxmIEhCBnCYJ51164Q5gRwKuGrWrounKZEUv1gZn6wzfkuW30nt
6W03jIAODJolU249q6ZmBTKa2+amKMJ6o1S3Gh5ENHO80X0ueHp63W/ksCnQXJwuWhkSioFtIdEp
WdSiTvgBgSbZ+T+LkzVPkwpmbELltT91Ru9PF/VlPPJa90GH4FcBBMyrTguzChnxSuLCI/ak9Cm3
ucSA5lpyQC/bjvmHJ8gBJ88SZO2CnavjwlMdLDo5mjIoTTHGVsxPCJ6hJiEHDNB2/oAXfEmCEfDJ
UI6meVJ8pfslP2fd2zDCVwlbVtyzvjfreIpcitaPOV4R356pHFFkrfVCYEIGuUEGK+AzE0zBcf9Q
7Gm4w+uT0IVI7I94YwOo1j0F9X8z9mwxIwpNVWZU314Sk+TvCmI/KVkS8JvA+UcalkVQjo1tujcV
uuojs0TcPHzXVoIghCbOPEaXor7ywcfJVGlY/AWKOK16i1vNKOvVutALAmK+9EXMu/O4dCBPN2UU
GfkT0UQ6KdclQF2hLwbfiWt7ViQZKZzQKj1d0x2wKfj4tg8v+n+Tus+iDGA0mcg5RaeQWFlxi39w
1eIC/GjnffbLSRvoqV88gviQW5xUfQhn981qOiHTCm51YjO6NZIozdSA9mZLyczV3HksIXQBF9Wp
/yzToo6wDcA57orhe86Cj/Nekz6kuWhtiZG7hduk49gzBTjVC4DbG+lJoO0CH3cbDrC+Nv4oag5I
Of/wU/HvAhKew3AeS8nkQ5gMKM4jpueUvLRsijEgRLPklm2IZ6WjfIbLMlv7klWB7juSv46uq6jG
IdYIjY/+FDEkrYZvTdOvGsDLNC0J374r5QL6Ll1DdQy6VPaMh23o95YlEYaHVmjbzGBOQH59I/q3
LkZzlRCY1NTh6Nu/pt5fVe25n9hM1bEUExsZ8Thr2wm/Mg/j1w5grGNGw3DtYiWc4JtFu+qOsCq1
lSudDLzkbm3B0m2t2fzSHvwzKPOSPhM4ZInMHvPGpP/Es4Yx+F8YHMiSUiavafjiZfps5460eKhb
JcUa7VCNLptMuPTO3Zi+JXhnjjV9ivpHkyMt7lu6DVcr8e+KWXVmYF0/1XiTrxthsnkgROR1A0MD
dfi0ck1a8J9r8JXadgJzRqFkiK36B5+O/yHQY1fd30bD3Eeb4wY2Nr6hjihWfeDIXFeV8AhPY9a/
x968ob1ZNUrnyFoSbV5xH7rGw+Qw61qBNA5apnSjki9U6HM/s25w+o0bA5aBax40Qr7vSc1wCinA
R8+ZNas/5Dz0SGkLKHHB2yPR2xsvNqmDAEp+bfrNEiV0fz9jpk7COph/MMjAx+OMulSihgfHn6Wo
B13XLelMq344sYTxBThNAq/gVR5Mu78ng4TIc8yMvpKtnmzZOSGU7AiiwQ3B+f4JpCpA6LnSoxUc
/ykXkwWr4yTud8oCuwpTSxH8MlU4KPd/7MEYXUlHTqiDf+TBxPLW+yLPxLwVCCN9yZHFENEpQD9r
xRzs2WPDj1LC8fTKF9YJ4nms8nKVuBd9NVEHhucvuDlgHc07Pr4dN2tcxv7PPl6tpU/E2/GsEA0E
/f4WgoSMDtsQCb+GNMirMEPxGswjXZZdm4bwrNrs7GQjVU6QFj9DTE8ouEMyR5w8wkhJ7LwgUw2K
AvrmVTQHT+sRD9PDsSCSFPdjI6ARV9GHmxFHcJd0kzsnizjpOvKN7En/Cki+PAZoyCd4s8WJTMgh
FO/VYMCEgS3BtyS5G+jZLjXUmT9pfwxf3YBk+R2YP9NwvBFz/lMFOG7rHSzr5Nsr8MOL6MfhxgpV
BRorJJ1oAsIYOS2HVvKHhz4VeGLml+iLzSJb0/tPN6cs2V2+m6fpisc0F30N8xcnc05S21hUr8Op
HDSwtpYWx1VDbgyHNJWC1ALG40jHTpUYs4fPpFY3/qkp8AAOfd52J41eAA5PNxA4JQUXxO79cRQe
pJdHf7Hnecxh5hPS7vz1mvGKI3S3Uye+iryQgYD0Km3ThwuRIf7bZgkTjnDFX5C2mcNit2JIed9D
8TmtAZMLzCIYStIfFS5JGE57KTJuUHXD83UoxjPI2hzhZwWe8DAOhkR1Lh8A+SKoq8PNKjtg4n1N
Napr/3v3e9k/G3BtEpw0muMArEHpRRF/TsIbSXAYViV8vJdQxrvz7OQQ2pd+TM5It0IYIVP/9br7
awTPlqh7B07rp8HjTi1uNJARisxIA0Rjd0T4OMbb7Z65qzUO0HcogCOyUOzW72DYQSAGOvjfqcHY
OmUXf5VZ0KoTHkVYjnwfHMTXRxg+M9tKy8g+7djQXI9lLpAtDKKcs6Xe0JuHzf2xd0zfHEEoAkiF
7kV0TpbM6jdM9uX0ifpmFKtnrW4b7MKcCJ+Hl76QRFJOo2eCrdAXTI07VEE5HrLLmQSSCcZ2vbs/
+Q1v/h1O3a7hl5DdBEPBixquUvh4DgbcasAzjKGvRPcLw2fYsXlAHPzXaRj4puzy4wki40TukmGO
xrqh+abgdmGYhAYG3nShiY57EJjy8xvFY9oAqkEjxpRquj1oP0vffbAet6kQJhD6i+AqwX+rrcKQ
i2l+C9kIL1TJ4QNjXPVHeoV4sj45R24ChMFh49znLUJWpP1/Djo8twG271qPnLbXJz7EzAAnW5xo
dCJj1v3jItcC5yGtgGRmJeCKRGmqwVEmZkRU+2uNDXxfhDPoOoeZBWb98u7V/OacwyLDUe4IA6Jf
xXys+NjSCRHADTcD3k/eg5+1HJ23G1Zpl6gwFWsYTzuptxvZ+GBnnmjpyEQ5ZZab45N+6fAN2cWI
sJQfB/mpW85+Zlb7lYs32bXUbK7Ax/F6RTRot1neVVvY+t4GgJnSAsKTF741UHuDyXKvvFa0xX2+
jCjsNdIAHaioBRRy+bl2yz/R8PWjL0HNs8DUP2xx77Nrun51MuHYpVZ17/r8TkMEJUaxJVkvuebU
SA7e7+vIJPD3dTlMualqYZv16ft2CGZyyx27dzN9JWTrG8tJL4mHyxa8m6lgtzNGll5Xnn6amT9g
44P1qVbFqIYXplLyjq+5bysuN2syK08OBJJnAk/n41pmC54WEKoE25oWMWobg8WjAaPKTp475NAa
LV367CYflsQxHLlTbXOcFUsMPjUNjavn8ap17H0PiSQ4Vhveg4f9p19joq8hLqZmevxeXtQop0zd
IyqZtWEkPjDc2+VGLxmP/d9k1l5IWjRE4OKMUda5e4S9EaJkA1tX7o8Gsw7hzTZ9BDVk8Uh7xGFW
HiAS9UzlAAM0+O1oEEq52OUOZeKrS49cSxrvBS9DCb7Cg5onnkzfWNO0vx2gEEvrZt9oKu64FNAQ
ZFrAN1Sz7SMvSeFMR+EFPrUsggJAJ4AAfzAqCRlXS07ULHULpK4HGU0do0zdUgakqSJcdhyodpiM
JTlA36o9PzQzgzTIJkGOwXXgKIIKz7e7/3PBzkvO/ZAUDKtwp2WTw4Z/zafbmx+rRrssDbzSqCZN
wVHDrIki4175qU33KI2jN6qxqKs2otp8+P9qjo07WDSvI/vYAfoNFsOarOW9spYiUZ6SxzxVcnAE
KTcio2+KHIcXPobCV45upGvyT/QKGeZ6UkWDvWbuTw6nla6WrNLcPfnyYhye8s3+y0rAp2iEFH/R
ZlBZwEG+Q3e3CC9ofy/wyHAvfUXmJM/lRW95k/+0BbcWjsVGFT1owKRdRK5e5k4aVlAMP6BK/DLH
Ux4WLiI+ha1qdNs57Ahy9yBMte0rq+Ek5zCtZ9fealW3cvR3ZppNTzl9iB+GCiopELlqzQVqruEb
BkhxH7s7d7+O2moQM9DHqyNpXh16i4a/wEA7uopiBwdYiwshemN/VyITI8QulEGbKdyo1bHpjlmg
bTX0Qd0+tDaK9NP14TaJob9PhHtQCsxix58Z0dRpwJcGBVrb5IHpiVdGPO3h8njqrwGHqlIuUT8b
X4MI/45Mluv562wHs5wahGWjozTwt8t7I8qUMJ+Vnwgx7Lf5ArEIp8A9OaquR19SjlHJVPYsActH
8Dr29ZYL/z+Y71avqEQiaJeSXJe2xIqbA6Sc2KNmL+Nhax5of+aMA3yQyp3VvlDCx/zLcfsz7T1r
qjwgBoaPswXzpP4qohi+fqJnHHirdmHaWj15LSzmel7oHTZyjjVjmHVyz8YqxAecAoZs5N0W8iLe
VHfO3DN8PrrNtaSJnBUA9zZix1Eg51TxnoQtjKWe/mMciNEA7d0/OAW3qC0/GIbaO0I+WskUeNVF
yisGW5tivdH9E8TMN+7sGI9ITnFxzhMy9TGLfmDEHnbvjPuFnG93+gsYB7PKKwp8WBdsHzoTK/Xn
h5W7rNoPUext7iTrl4z/x9G5cG91Stzx1llfW+j1ellhBQ0HX9wspt/MspifdWgxLrZ84YP7dpaZ
N2at9lYQ6N2g7D8Psux0R0xfFzTITtBnpfepylchqCmKLUsSMbDXCwa/ZzYlYW366sgnXiRY5bNO
IqCiS3A/gnwXVnPURpX1sIQyowCWFqd8jDbQ7bnWtCllga6tliCpf+nxysHjtuHzssiMJWj/y28T
dopWDzG4vmwdt2KT+Wf3wSoF4qVL5Tb2eXvZoe6mUJhX0B8cGQI9criqW86g+Hwz64/FylINTeG4
cIsZLSZ/mOcZeOg13ZlS8SpKr3vMP+NSJ2zRp73ZeGypmRv5bb3nq7P9UtliAvb/pkNB2ytu8Uc4
DvDU8ZcxWfcfaNLRv05HbX72fZXFLyO57x9o1DaNiDxFJwWps1PKlBIzfqH7dpIt9TixhFaP0+/c
zzpNrSJ9Z8+qaQ3rNH3Otf7oULKZ6SMQRIBFDh9yqsHWzGgvSwcO0dWwztDjaqQHSKf898hsL+ec
Jaek01vqe5qjGtnviG/82LHb6AYruoFkKDQ3/esgvUsuX60vpjBj5EBZIIWl17oHC2MQ5C2fLrhg
r7HKA6APfnyI97f3o+oy09Ab9AbOAaX1u/SA0Jt9TkvS3p2Q+kCjxF6109JduJpQuItQ4LWRVM0M
eDsjpe7E2FF2TqNcSnLJdYTNg2BH9tvMxhNehtQjQnk4M+VWmRQiBfaT6msFcBtGC/a0jGhRw0sE
Yf34IWZvVaG5VjeX1/uYQ2hgODjbfw5MvPGN597brYqWgvvUrr2TifGe+ovcJSfy92dSMTjtsL1y
rZWLqrM8K1yVtv529+g+2/nVYUwdOLMPF8nZJB9SmdHlJQs3bB/zZFCYBEJng4Oy7jfNZgkDBMWI
6h57LyZsJZx0mVk0ykl4iDmlK7/yg9awhs/toTJPNHh5l/ry1q2asj2454p+ASpBkE0kiUG2u+l1
ziat5lkgELw1gZgqZuRgkNfdX7Z/Kxy5wsCUGu9MEhCcV+idkNXiNOxeuD2+M6OqsVbhK4WvIjfB
EhlSveiTES/eKbhAIPkHp/IH4IJhSxky8YFp20Ee3r9bzQStVRC4Rvj/7VoF2eTbVSpVqZvn0sFq
v/zZGq8vla/uMjMDLdWu3QXAGSuN8XtFU0T6u6X7NsvEmMzXAb1ByOlKcpZUfTYdTqbNp26EeT6e
UhsL4x6nltH0N6+QL89D02W+DepE8VQyQcvJDO9DHENLF6gUPOvUj5oYM8QazrAUbt7waDs0+QI6
uqR0RuOE1Y2b8d3hXUxjIyp+S15WpagldWx99jRnpwEIY2askoW9qlL75VABybVPslREZfuwDwOV
0sBH6knp3S2F40KLreP41+MAdO6AeYtnj2wZ87KRYJCPKi2HtXzU5D4QnX6Pk7EKtdgOAlJOfi5s
LVJjrk5uVyoxMT+thR0dgSV+Sh346M7lMkS8AXRSpoXMng3/jv583Fgdoau7swonSWyZx4LR5M1W
YyCgpuX8rONOWKKdAj2QXesm7B8PBm45Djxqg76rt8ks0x+EjdBHyEzTVufab1gwnCqg8ivr0orb
opxqYI5/3lwVVzqdGvzaJcm3tg9OCNfEjSDEj/vaE/7PMsxw6nnHtDyzhkkZkIxhjxBm9gb4SFpb
EKKemtHtTQ8Es7KHWo7kZMwdZH5SqUSzqZz6NzeO206/IOf1cH/18Dija7RI9adr+h87GlROc1ey
jMe7wIzkQD5N1ATrBUibTCUTuj8mbKoZqODLVzEh2IvEQBEUUfop3J9shGXn+KiYq82nIBRV1BSo
XVNtuecGim+bhyvMB+B0CMNyJdIVIcrscXZh8ZeUBHSWzCrRihpjlmVZDZaFFXzoTl8kvuxLizsW
9npLVa/5LfYwhdZ3ZwPwnzFzvDh1wY6DJU2A2lu+sOQIYUJUbuITzsEyJwpwiy1hFgjUSkmL4X1U
1GU1MM4dnpe0b/Qpo0Ls0M3Uu2zRQa+g6L6vdiJQQNDWOKpZKCtD8bT6DMBTkzumINqIEdREScc0
iuX9ALUNKVJrZWUXI4GpMNo+lEcqx2El23Q/x55HrV/vzFBLwUlhHa2UwGC8xNjoTi5oQDXLqOVF
/jYE6EmkuSD9zG8YqIsXPwfaYLH33nu8EXD8NZx00DXZewU5d6yoVbxsDOS19fKMfw+dasTTLH//
6vE/n0DNbWTooUL0I9k2b3PhPpYgdN+jrLQ+pgKnvp2TQx5DHDjAhfBtBz1+DKzT6tpjfxZ+MsZj
GEI8cM/fkBabmHGfzvLdJz2CmVtKHe4Fw0Ew0NluwbhkRTC4i3UVBP5Ep/7IulX9C6ZXYpWerZIc
YdIYm5npPVqRK9j0s6J1hdUiqVwcOP8ARrghglNQIfAPbvw6Q43RzYv54yfhrCyC0W59Nb/71Wmm
sxt66U9qqNqS96sfMCyNVEHutUPXEc8bnKZwwJrpA/oA5Z7e+8xxQ7eCRSjSPC7qXvT4myPwNEzV
qadl5v1vz+jXUTD5W5NPsYlTVfQRyB3nndfXCh6fBOmW7LMOEVrwuMunZufGr3e2h8+lB7dIN3gi
NR0lqUQ1QTqh4NQB7GNHbQtB1DygrEZUdqVTJY50lxriHDt6DvGcogiOtRX/ZzFG5kFCGnQsGphr
6+W69ZaE4J+7x0Y9kaOsh0gNmFjr1cEceU1vlL6AGXnfJsCttQ49ul4P2KJzsosQOHUyhadOqT1p
5+IHyRDM1hNsxdDVgh8//hEZ5gYobaQKzlb6o9yE5t75V2TdItYO0X3oI69knkl9AZqzwTdyzqDJ
+Iv91oxQ9HAmiTGl26MwKhfeNLd4A9HD52uN50n7AbQTu7C3haUVhfTwAoaogL4nYI9lwZq0vtNO
rtPTLILEBlVXjmfmYQwjezLYqfxXrcmC5MVM1nwTsozxz75xJd6vt+h7FIQGbUrcISHJu4B6rKoi
gMrrEYJL1KL/eKsdkhVBvgtHkDM51lfwX15XjlXJB7M1wXYNkAToaRGNEePzLB8DBqzHAvv104GK
lKg2ttKYHzrD88vmte4iF31DblU9WQaajb0uOpdqMaYmpSys8kdB950VfwRPYF86lNRuDfwoD9Ym
1ZP3L3UD9BJHBbziH6HHe/Uts73dm3Iltsa+z5yaNehXTLXMGXdQ9zaTGkHPPJVr5kBnvhn4kAl1
uDAfCkVKV1tC1dKOjmMc305iMUlyA/z8hkCiez7yr93CQfi7/PIV9UggvmD8wHbpaVEf5DnZigcA
nVACWAdrWj4TFpLYesw9qT74zAy+X+eY/2GiB48AYNuLBSYpgBgiQfVZvGLAj/vgofYxAVgFiU0Z
L/xcvSXg3wXamfA515cuhvdOgGgE4743sjnSvEeB92LVoPHwk5zcmUeQbXiyd0liL8fr6GIpBVG2
y0ka9XsfQeZDELT/gCTs104Z+BUHXEY4vuBl0hhAnyEDB52rUkFgbjVbOFrC7t6uJishd9OMLYxY
aUMfdBZWy6Nx49e90Kgf1VMZY29VwfpXg+iKZRlvMVv3MWefrsjQZW5RBIt7R0GyxKy00mEAyNoX
Omc9Vr70oSANH70pwpjtWXLBqPOENUGvLw39IdEVcAg2tHDH+JFYZ7IaFm/peXaeShgwxEN7unAt
ePg2tjCAUBq5y7D56384AM1dyFinHRAvCIUp382NiTRjncs1WFU+Wju5bao+mICuMvUevOweIDmb
P7FWV/F/L6hH0SqzpEM9MJ5oZuiXyQ2ChZkrPMyHM21TgmSLqMW0qzvzCJzojZGvNbrKvqMpeTEn
Xw8aUxpgz7siVatWqOy83wkFO6d8CAIYQ3tySJe+gM2U1Rk23hDpTQtHWnEGJSzzW8GKRosoy6M5
bKxEiOM58ERej8ofsBrA2CTM4a6JduhFZ0Jq5yYZGf4oCqKrhxWRV2clLPRoyxrmpde/C9+JxnSL
SHfH4TtDFJVsy7n4Ty5oyel+xrdtLEMKQfg1oPxO94TBOQRnvE+PlslU5JHgLFvUTXnhhOyuyh05
VMw8s3oPN7iR5YXNHqKAlyQRElGLXS28/yvB5/Lt8+SWa/P0JMpNjIENRUPtyy14sGLJBAX5rflb
CZa54I9hCzpI8U7KRz1xtDELFfh2HYVdBnOqgU3xQyzun48GlTzxoiYPyd8u591NNdF/3qS6ts2E
HIYgwoHrBtILpKoQRCnFxDWpEOtNQ7q0w4rX8ZvEDmkiyXF41hww0uAOMwrPr6khTyLTI/x/eJp+
JWYL/nvEYGkeUByJQPOWhIYpVLpC/trNCreh1VhYpnvuqpd6rTnnk8gfhYROKzTxC7ewvE393arC
lRzbwkzMLr9FRTLkPXu91GaaZu1e5h11/2YVAfXd+NpHLY+FPRD5U1cRQ8BKFU50uY/Rn+P7aKVb
gJyhn3jyFTM+hvQ1rv1yWYlOOVhjJzVLJjIxBqlsu1MhJkPmKWxjJxp4sW7MjfGDZUiC3hE98iIm
Pxxu3wWjpAapIPfd92k5+F/gYb5KosebJEu3c0PxQJ7VXtmr/fJ6dg4ZLSgPkw3xIURIspVGqTBV
x87L2GKuMglOV0/wWlK4kgQWcJ9/aiY+cJTelfkmuJARwajxCEHnDJ84WaG+wOHvlTuEF4u/R9N0
yCnx/allRyaF3QSMe1L/Um/uPaIf7N9cACObk6M6Nmkz5O+vEnlVlUEXzHdNPOl8j9xthk+KzFCA
scdR88O0ypD6kXpzy8nfgt+hQ+rHi5XPtBWzQVk/1MKGAf0BSU06HTuJh+FRtWffb8KNWonFJHIT
Xzj8K7pFSOkkeFZQi79zva5araq3cw/BGGS3CmaIChRsK4V83MISo71/ZUEtZk7XbKw7saxVRyqk
FLv8Nm5PYCmB5Raut55O0PZcg6TgewLYVmovFX8mWodOtGtt0hJeu2+cbmbjU5489/AKqUQTNQdM
dyRZNuuxwrPthl2CcoII0dM1JX/tb7BDXjknVtOfLkcV14br0/MdSqfF348+tp3lhrs08HSUm0Mn
kcVcpX1oF4Tx/KuZIY28nTzBkBpJdCMhPI9TlXaA7pkHxxxk6OH5OuND1uSYf4SQ1YuqUQR29Sco
gTC3TryxiuTGcNDwYKu9E+HbnF+eiJhQqol75g3PeZLfu/VCcB9ejflKpZTzXIZil0HCTmFd0qGg
AUouH0VzrVTk0hO6uSrKD0aQUcLzUTfNgBU75fJNHvEFaXAPjX5FaZY0APkMpqIIZxYqwARQ5ZBu
MyeeVdIMRbiKpDoeHvRd5efCnhoyCsI8rpU8h+T9qlPQTSn4p2lgzrk40mgV+Om8kilxNWV3nykj
gdeG2FS83KPo4dd6aEhkWCY7bBoxQ/+7dTtCLXS5nT28gyg/753AeZ9nylSO4KuPyaI8FA+i7FPH
odb5y3UxpBdp/WwQPzYKUC3KbwbBTm4O+vzBNcKT9u8fpKkZKildiRwJXF9E46scpHy+JlFVjeDi
1jEhFkYnhtxE8eCuUGU1lbJKqe+GuIYLo0/KJFuuhMZ57Km0FVJyL8Nv5fWbCTPO7fzIQIWVq77w
JVc0HFaxi34D6X8JrlJb0D15ESE/dVegVEZGRQ3ztiuWvWUE/OrT3vTSyCeA3g21UHMdCYE4GDat
b9DPEx92KNOdYNa4xowSjV1B6u8wXmkKwZ6zFarFrMwuP6IZCorQSOeqjJGaM1TZf2cJZdlQpdl9
AX6P0LV6tmMSAyLZGhacgvYsbP5zH9A0hLN1q0G7pQ/ny42vZmmxtjljShBJJQsHE/49HJ+LI1ZI
uZ0aJLAgGkQscmpQN3T5KCEjxeOwD4a8r/ZNaLGsUbn7SC7Cv7S29oqnQ0uuzH2qN9tmg3A5wEs3
NFZ2DhYpKsE7j51963jbU3z0/BTnyNYbEqHvbh6iPr2Ei3xCblYLZLm0Zt6UQ6mX+F1pS90F9dyv
l/TUJOvMd9231gkDzgtebUqxnhD538FZ0/W1Sz7++XinWG5a6fNcjmy5xi5pN1IFUqskRz7yEwP0
ScPiHWwWSvQ/K40ayAO3o5Ce9fTl4101szKIZnsjAPrHjKnZrpV12PUbgkBoxKzJdtEeLLhMrtie
/0s8EzhmW6GP8afMMBtrjqSARjIRtjIRPY0yb5//Ge3/5AXmzqxbTPXNzIcv64DwbxBcLhxdJGXF
OUriFliE6IOUfElHNUZaa/0DHcIg/tpdVskMeicQXb7tzaYOEyJRBQOJROKqvsZTr6OKApLJnleW
KM6UlC5qILGPYwH7ZG5lBCBmm+q1s1LlinBfehXgR0df+5Ip+FLYyjVXr75f8FSuXXa/ouh2ZpO/
1tefIoGalXNvU3JlVoPezbCta7Q+JP7lD+y5/BhTRzP7ufG516x7Wbl1zqli+j1hbw7e7kFmCU9S
G4gQByf5MAHhJRA7QJH3OIJO9kz7Ay2feenNMBNMXsmIPPvCAfVc2Ln5kXAC5dsH2T943XR1sb9R
crq5M+5laK4u46CQtng8AMMR6Y50HNf6Dd+9rfGu3v1XtPS6tOKv/YEfQT8Qm6eEdc1MECToTnju
IUNdJj3FYKWeKgAcV+i0gHV1a3pEntzeEgF7sV0vSMgT1bMuh6u7Bu4mUuYDuGVma/7Io0kPyzmo
NSLsIWztgTuOW9O77zPH6Rtz8YDjgpm/u3XYt4UCP1TgJj5iBxjWubtPEJ1eOIlAJB/hBGVvUVtH
k3dNvWdCDV7rbVS0vnmFdhM0ST9ygSmULmmOfmTuFQWYWdbTEd7xaaLXhevDM8xTZDLYuoeKPdh0
bWyp9X+41u5xJHF1oa3gAx0q4WjGbObINDDptRMPYUY9llAApJddWs8BmdSRQrBqk1Rl9Fr3PEnl
g+V02O88CRpfUFpXXSPadvIeKHPsB1D8uJghIqWQbqH7V2jJY/gXK7Cz6IYzrIDNrHE5OFOpqoNj
5yITK+Ebe7+JQVlBZdGh56HiQU1VK7Li4rBA9KTiwzjbWaxHlI990i7c48FQjZJQ56OJqAlRKhxX
F+bYKMBqy23119W5hSs0wuOXmhldmWHW0H8fKJ30UChwuWE1Lyvi77e+rXZtJMMaDPHOIuicN35R
b/zZo/4ggUEDQzRia7+BWO1txg0KzM7QAHHoBS+ReLlRLPT+ALXBEMJIrIHi7dkL4qTM+UmbeiKM
chvKWexYv1PngszfNuystjoyRHtV3Jp8JvSrDvlnBVsoBjZ2BJTwSjoDsOP7FBUuyac1uzzEk1Ps
jFeHXtn0V1wo7/ylTN6dY8+IbP1qHX/wjGbdTQQc3fH0YglKzazD/P5t7FPGX8BLt/kLU6BlTOTz
PxaEdooICjZpyKHfv5R0MBpKD15awY7v9U+IOQDvyjx8ZScwlF2xMRzI8sIYciclAtS3dgI+eCTO
XysXc+goSj6o/Euj95kGtHsCCVATDL9EH0Eo37gb0AlNwSJe+w3l7qcLcXr2DVUHvaMGSaLo9jmE
R2FAqbLJxViVeaYrkMC9VLRpqCNgyqTW5k1IozEhxIAaPSzt5GkeI/5PoSh0vnEEDQK2evZ3Ro9J
yaJspVj0SoO7+yOo4DvEGiB6XXOGngL71TJFelCsPNelNFYftxnliS4/524VKPLN7nMNY4flkpvR
rgQE4sy+g16Ge14JwVw/WRTqZtSjo04wK/B+Z6aSPXLR6u6l08Hpj7CXPGhDFUw8wRb1/bbBMQpj
Sz5jrqDW+wuy60H73dTrbkR5PH18uXOu/n1VnjRsXLJI5qtgND+ziIYtx9ZofHpb1GFsMNLNa0OJ
dqQ7XIE4D+b00U5zsYbZSls9+cHBGbLWvt2b4D0zxjXu2gcm07yhsY/NPgy4ni5EdlGLf1rzU6Iy
PZ1ciNF0DeOBPmRp8U4Hz2sqbO0J0FX05/hLq+aZRUM3fGDZqhDZEV/sGrW4drWHo8lCACO5/Atk
atXl6dQnKvt+xIMscYVlu1JY1zt5ZN12NQL2LxWk8KmDn83z+DVEoUFYXLjRz9+v3S/ZIvk/fNtE
pFaqQ4NKsVoocpSCgM2DqY9+Atvwtvw+5NTI4/D8m6rsXfHq1LLqpIeIpVu/6fiw8wYGuP0VGQ4y
N5CJLbY+jhCU44cRPgD9yJJaIpj/UAlLo0zWRLahQYJG+3DvHNKnYT2XW8GpKkggaW5AnQXE8UQI
3B2Ny+nKiYutX28G4Xfk3jbz1Jcu3ia0dl1a8466qUHjkZtJHb6yz+TCzDaSDyQ4lP5nZJPkhwGz
8CGSXlz/ei+c4kbUWHNQ87kATTOH6oKl6rLgfteBdiJBJp3BtIo8oUSwRJQPAjXYgpmXEB9Gl2/0
lPWyJThdoTmntoIN2yDOmUWWyhqi33pZ/HtjdRPzusY2R77MeuL4Is3GPUZMHaGA6RNG+c64DZfj
TUWBR55G02B6M3lWefrMum60cKDKel3qmAMuDwrt/dbTkCesjPmRSV9P4BiWCNQbApMae4jvpPvL
d0hc9dhZIwJdEygbUIy9C5KBlDOD3hrXNzPDJbvG+cW5A4Sp30eqsds0JSIeVBqcYW5Ow1cC5DeR
2r02o2K8IKP+TO8QUd7Qczft0vufOXzdQUkaAZ0PaRbi1ygW2wHr2zrZgo214uPsCTzOPSCK370i
UdX3uaRmRaJ3JItYn98I4RFpL6WlsuIaaAqYaNItqQHkIZgKVOkqU2Zz8e8G0+0Z85bSnaXDjHJm
dLXiVoEceS1TDf+erwEpDK1EyfW4qreC1jisvUcikBzZMHLqZdHNRkxvZ2g6f8UqJb8Smq5JWCLE
EKIK6l1qsNqD6SKLc4IAicNaPIDWPNTWy2w60aLU+DhEfbYogW3q2M1HtHmlj/gfAwUwVvsV+o6b
Uhd2S9PXHy83iTkYEm2rBi/oETXitFrcraqKpzJtt+hh38Tvk3Rkc9g3KvzZVqlqrLIqTUkb0WBx
1jEx9ZxsJBVci8hz2KXWFAoAHCXIkctafB66MNkCypsqWAL7yOeON5c/s15VXyCdH34VvV3FuAmS
iy/Hycl1H6kHHuMfRl5mS+iqNBEJ8ZzTpFleIey0KLzLLalMEZZGca/dxtesXuK42B93a982oTug
PK6pMmZEUdJf67m9qpPD3Id23MvPVcVPMhUlHoknLNAi7J9GCkOE8xOfcaOlCzZlZmiBggpxS5VO
gj02vwI7l6M5mx0E0Jk6i3DJekiuNPrIcE4n5kdNGkVoZ4IHKK00D150C4KyQdvf0dken9f47JQH
e4LBxPsdQfEZdu07FcX4toSSRV7rhRW0KQi3t5qZfeJrS7pr4qCO5JppUf/VAORjdgsrPTkjvxZK
l2Ox6wqOsxAh3MKUesyhK0nXiCZHJbgfnaE8PTK9+TbgML/oX9OIbFw+DiP4EOLrI5eZth0gJUZK
xzxjWCSKrg06AnhYDCpKXCKyiqppo/oiCqSnFt1I0A5P0Nv/yv8bP7EYD674TxVD8vj1RGjlKztm
eGPAt+JYpgUZLjqrjz+AOq1HPAfoP0EiqfRtsBMKJPBfjq3ESFFi7pUrVh65pVF5VIpjnimMA3oM
4QgKX9vOHeeZujstPIt2nuwDsD47DBO431JywHOtIPffTheMmFaBpPsDf7+es03GMec3m604w8wg
X+eMwUdhe5sJNWOB9vNqZGXZB7zNgxPGyI0pYtdi3rcEq1Ap2qWOcBsPNDeKwm7TTRGGEMlylL2d
pYMuI3dFYAwJfvPF4ViAGvVzvhW/v42LOvcoMGM/3LN1Yo0vUfqoSBp6kI52L/TOIiwpjT+TNN/7
ftCSOyzozwoD11+a4+c5tUtGCjehQjAMQVbWddirtXgd0QkPUK6jDys6ei4nMkaY1SWFymx27N/B
/KoiM+XClmgRGLeIobG5EH5Puuv6UTL3iRZL7dakTL4YbIGjbz7X0CgAy5YIkiwhqblZxH+xM3JZ
CSJ29cCs9KOytNMTO/TPnHFkS04mkgERgZJdH5BXkJoNu2M0fOKIdHlggp87WfFo3HgmR3H9+O/c
kcM6sfQVigRvb1jHltwoImdeLkJreR12I+nGt6SuTqcPQDi1JshhA2BKi0UK2jC7HeA9Vrut5da+
XedrtHaF14PRlVuacBfZWj30cmK5GGY2N5/UvE+0Sgv3pxlAAg/T/xwOH2kEVgl1HcXYj3zU/mlS
qFfREjnlGmkABKXhsiFl9ffGW6TKdS8aVtthbTitwo08YBOXudYHdf83ChMdA3EN22O2qhs7gbrG
7KzAwk2BHUWYStjzEei+KSemC8GGgmV5uYrToMJwjSGX1KF1w5qtevfGU6y35ZyBN2fWZZf9dDPo
9D4jQDYJuwyXo2i5z8IRdJE2RRXfPECO5Gyva0xoSgywuNVz+za+zfnaKsoJck4iV4MK8y2LhgBL
zvPu8VPnsbCwoa8EzCyw3yQfqY/rAcrMFdacNDLdXOdnZnB96q2sqaQi33wR5eowwJc+r+NA9b7S
1xom6p96BoHgaK0DO7ISNrwrNqkrkUufAYgAHRoUOmYQqJMK5BovJHNm05yJFlnioJurNXP0im2K
R7VT8jIzcZhdJQ4CxVo6IL2JJkT8jTFStUBmHUK4bZ1dVKwbm2FWcC7h+XEIS+plTY2LXgIeAkIe
ljwUjjNSxprKcdKqpQaM3hfpVqcg/TsUciebTqMXa6bJAGTHJ55C2mn6wfna7vzAk6E26oY620tl
zGKetpXShnZn1uckbLdMWjzrR9VAefooycuspHd6F0JmF8JSRdo9gvjEK70u3n70MjZ8l3yxPniY
M4tyAR64voibYKn1B575fuL00AysFscdRBg90vWVibGpNuHaQoIMwAg8Zk/N0Thgv24d6kI4zypb
ObfZoCw2or4FYzKPC2oFVYhIv1V057dDqk+2z2fONLQjGqoey8MR9raKnp2lQaebKq54hpqyurTf
0jy8x6KkRRjlcIpn50qkkZLFcYTdSlWI5MXrpTXJ0OWn8d91rrCm09OOZXFlxRTxA7nKsGOlrkNj
k8yUE22DianK7Sa6CrdXuOtlsa4V1mvZa33y3Oom4o6lDMINXMCNRqUGrs3IWSXaASw3y7scYXtw
RC8HSTU8D2RxNq2RhiQRJDcxezcFF2oq7uRU/u+OSlX33cHhK3SKyNKEo3TZz3PieZh5Lt3kZ+AC
lXFeCvl0n0dFexiC02VOxAQOtVtmeaqjZ1ir6UJic1xCPdVsPJu341lF3SrST37klqvdefq4SMZx
fPcexNII/uN91bli1EHF+pEG/3s4ipn1zPahLicQDOaCA17hJS5rvqdh9NtnEQdfqAbpM7gQWgdG
Oix/X43ag7zGQcfGUssL7Hjnksz++9Y/YQadP62/0g7nZSkkisnX8JQqHaEhq0gzMjDf6f5YxkiP
98kYrZ0LbKiFngK3LWIyWwcQyldTfu6rGS09lT+vVfQi5eLtKZd+U3kq2lD9YrdoYEtqKTGmAIHY
3DGb8x4fCOpNXeAJm17lTdSsAAIqPAScG44Wqw/dP4zOYhEnSMU0RIA6yx9Ymrk4QuwOrAwJMa0P
S14sxbBs7cKOb2klSiDOB32F5LXD9oeYRhqZjq99dN/FnXLdgVrR2/+Qwp+AUd+wRQoiPjJ+W9XN
XG/D8MNnlF3fI5BqHhcZ6MStEXLuTENdQcyDOWWYsy3v2iuhuB5+tpGGFa6kp8LYSqHJ+hR2lOue
+hkFBROSfRfqMERmhnJIRf1w2qY8jgT8d2WYUnGQfFdopv9UQQv8I2imZ61ydQa2aVxtVYAT/32o
lcnxznG43VPoA6n9OboK3SyPf8unCxsRUxQPLT4MivlhmaqotcQIKQlV7k1m2EnEc4gz2kO4XucT
YXpu0IoZG5XrjrDbMo6U6FZXUVVLM+8gLmSqsyCvD0y3bYg4NlNVuB7MKsYms0DhvC5rT4u/WBK5
sP784WVB2gYgX/Ezco44Og31udpa3yrVAZBUohkLrxJ3nCPOunLiIpno8zOXpV57igqpwlUpX8Z+
M0uz5rZRWQ7SkoSANx/xPO+7nyaPM2eZ7/8QMtQtnpLmpWbawVF4UGwdivRtvFbIB2jRVy522tRA
YddK/YEejtoDcL5B6/4gv1RMQ/0ngC1lmW9QStoenGAj+2OeOUYZrUJdXSgb+agj8eZ4N1kPnGgR
XVi+OXv34ArSlWXwqn3u/dy1NabFK2/b2mYOoKJ0kyVcggIvyM94xCTEIuU53c0vIWKITI9ZTluY
mbrDNWUqv91d6rS55KbMJ5rPLDbF4uWNB4ZwJWgWgUZhJd/bKvoYZl4HhqdRnrAs1YEiB7HJA3uT
Vxc77nykuBy6giYzvkS5RTIkuj6pSWW5zUW6TsU9O0YjduTtNdEqxsWUbaPfofCHp6eoap2WeunB
ms7t8iASqY+Ix8KuJinYLR0RfOKL8HbNhqk4F80zklI18Al6m+kGr3QG4AEOxi0R8MQzlSyKNVIC
YY6JFxUCXQBqKaCslQZX4MYxO1hTrpcNrjsDSPlLm2ahD2MAccB870LNWGcEfGbZAhk2iLHEUMGt
PYvb+g+RQiynsABj963tGuGia0XwjWJo4SgozRmSSFyNTHttcCdsdTdk7TK+8iC1ToRvp3dc3g/L
jxJXhrRCjmj8mA+93kiZP77cXsneWcKq1iYmZY1NHUgrqkCyKRu6+hLdnc4BM7S1ahZMFEREkJ/r
Eh/Stoq+rnyHyC8fOq9cAId8s6T7CE53G4PMiYF3g6pqmygaMuIZxTUVq+Udvc4gfX6gN4DdWjll
4yGG5t+f9EIoWl2Hw6HRg7w61LrQ9/IU1MOyo3npKiblXtrqk1qobhvtHLWUj7dts6ZTBtZaFs9W
QGlR8nHGkHh5zgGQ4SpjS4avJ59yAF96bzDNvogNae3+pjTB6v5tiNDt65MqFZdwNyJMo4J/oR8n
DzOzP/6y5aUfobKHLAEQyQ8CgbOaHkxI059on1pH/XGZmHuNabd/uWbvL/WKScX9akqgglig1MKk
Zu1yYSBnGPWUmdTX7TUesOfmnQHGMlbq/pSMLSvKvyryyPb7kiEjyRwE9POWR8xfOzsGFL6/0QJb
E9owwPLQDhtnLeyfEP8fPzfbdJ8lg/nqwqA5aBfBHZUY+0RPhobPec4QxXySuWbAeX9haHjeIdw2
QBR1XpS04TCLuj5C0rTckX/h7O1I5kXq9uWK1llgX4SrnPR2jDOTCp03kEj8FJyyhW+D2AkEZVcS
GnrXLY/ks4vLoVphnFWnpyrKID90NGz+1FupRYM+OLII4Cs/dphj+3JlVAHViFWw+QJU7GHaZm0G
AABNtV4WqLGhdBP3j7WqbZP4xr87YJVeyndxQE3IPm3zhboWKzjJSJAQVZO8+XrLWc4eUtZFKEz8
n4Tbq8jLOG+a9cb1C7qPZjiTX9PbKJ3aBVtVPlfeIDnCiS1Vw26bhjv7nrdGCY4WGLVYtodJAqsk
ZiVFDaCEjwuEoTrDhogwKCIA7jRjNO1tIiI10ZYpy2B/ujzvr4Gv9PbuOh03lqYTZ27fL2Ul4Sy4
Gdn7a5TxjxBWbO/Y7LamBmiab1jpH66QCf7+ATouZALaIhJBgO/ylpQBzRMjnYLjCMipemUHa9/K
3ZPOAaHfdZ0J1yiZS2jotjcfQxm+q7vEKnCyWrIGDqWBNpDdJZ9u8e6mN9ftvrS6an9f9fE0wTNr
DcRjXSKsonSRnghMvxw4j60yJadce71cr83C/stXjFxEYNZjH6mWwppX9qwtHwGdT/gOpf4506GB
ZRJ7mw6KMrnVfmC4ob+iakjbtddzzp6gUm69WiZYXQ0LEO9yMojyAreN1BtnCBMj2dDm01ccvDx/
zi1Uguzf7l7bLP4bppxlByxQr+BDIlYHI8w/YuC/TJxMyz5ayTaJMwTCaGonQ7CzijN2KEbmFtqb
AVbgRrcsm96xi+k1iRz8sjAoR8q7FycLVhVVuxbM76wK83kiPlWeo8sO7pkAwtOKPYZQSWI3eHRg
zar/C4RYZh8z+xSdlJ77RTlGhq4Y0X0THZqt5jeEtaIMG+LtTIp+kkrnGdju9/PaodoRSo7CDW+v
u3sXQKpcwAooYWkXy0rdHvG6yeUea6Y2rX5sp/MwVIi6ljhAPpdGqS7IQwu49J4gxfgwW+26Xa/G
PVPIX2Ic4TfbIqPv9v18cyVbmuxhiTkKi2ExTCeHA9FmmGNBt76XqYlSa03PTzSED97HCE4g2BMi
2dgQJ93asxgbehHoaSEW4ifiZAeBzwtTB9upZ31BNu1yuooaeebBXF6zqY1JwLQxHyQ+MXaWX4Q0
zgNEnpfnFlBEhFXKmuj2FpYl8F43Mfwkcc+uVUGPr9xbvvrDjKQ4cz9QhPx+pt1ZWJNXd/AUZW7j
n/evqLZUaWXqs532uJlb+Fhk/r194nbHrmQaCPngBskEhI5oGgcOfRqNKqF9yls8iixeW6EPU8kd
7DY8lghQ7ujAsqY808dbnYXlshJTq/fd3yqFVZ9rCHvg93LItsSDyKd+dN61IbwTNqnEIkNuOvRi
72KkVr06DuK+kd2pTQkHh3kqjUAhh+6dB2HuP0CC1LpBBRSCKEs+r4m3tugK0HX1kMi6g8CHSzX2
r8VjsjOoYbd1P9eSf0dzgPIaxMJ433GSy22Y37uiYI7l31KLVMdWqkRUK+9Klz3V9+K2YwWLjuZC
/+Hi+lUu1F9fn47Abo+yJakjnRpaSjLX4PBW7drIPeaWjgPGivW+crtJ926q0Ks9eccX7gcpB88S
ywS1G1Rxtp70NkDfRQn81N96Lq6svxma+BDb2CiKsOC+qKf4C3l9Le20Se3ye8a5u+16hTks8tRg
CvBlJCIHjlpN3F46mkNy0Ignq8RKH8K3jC9zrCIfetZiyseYRg0/hVF9tYA4y41DG+7bAFWAz84d
itaUVBabsmHi4ti4/uPTHxErct93uGkkFInkEnZ9tkQCElJBMCXs4qwKOppt1dj+elW8mkH1IotT
n3b10IDZXP46Hs58yGhyDIx2WDcUekUBu9ZK6OG1ThzoCnST889qT7nxQadv1g9562mBfi+IAjff
RZY3v4DN32C3mxcK27NmxtYkDYzPUmqYa6g0FT+BlO0JvrqePr5Sr6Tc3WPCPIxiFhSztm+Pjm7r
ZmPNVIBr9QswJ8K76tiSkDEkkRltGOJVdv/y1O9Dmk2ZwM11xNyhRgHVGwnSDXoQt1x/7EoyUQsK
K3WHgUB2qy9ZDdeePce2CSZouM1dc2K+bP4P8QHhoKtZkHMqB/mHnMvd75J2ck6hwfNpCw0A5yVZ
baHY5b+ssOBob77nslB87p1nZ15lNOsic5Hik5NMPTdzRHpO8cQPDGBiXt4m4BB/d5i5TohBu9be
wNFM9HFKmo6gvblBlQVFWar4fKI9IIp8yrwhXn/DnNXSUj6E1a52xJvOmIbWlh2RdArxlHcaXn5I
aQTpe8QVPe5PFKvocHDCVZgCM5Adsr8OghKyyrXL8O0UPkS2O1xlz6Y+FvYTaRpkgIIP2aEy1UkX
Gz98Jm9SLGQJ70J6Yj9gM8RBvRESIDA1dYmPktJIhIPjgmcaPBviKgc/v8416tBp+jG66HCuqJym
QPXA+krq1qQc5VLQKIEdDZKKrpxwpL5uQsmojGhb87FO8pkh8xaEC7g/tngVMBCFIXuItHPfWrjV
cq0k3PIyYNFcaw8xrhFRLwYVeLIGHzNZ+MK5Y2+N8RChzKQSWxEKDYAGBz7Qk6/EF2KUl+8tJmDb
hTTS5EkjGT1UrT9Ac+XXDZi1923smHGPk9umY9sA1WEh4ieWKwJFYD/HS0SxStUKu/g6UtbLj2cm
AgXI8v5E7yPbWdZjAQ4i6eEMu1zydckj22UKrpdA7YQ/TUdcbBQpgIv6J5aCcbUklZ1n0y6jS7BN
P/MbdpDfbfHKeQr8ZbPSSgdx7E7DAXmUsAVYqoXQLyEVl1godKzbj0BYMIH69P6OUOdD8m9kC7dz
9Q9PDoWtbRsSwK+H81ucjBlRZzFA/zXmEX3qHu1fQ+nE6KZyKXGF0M2pB2Ki+4YUm/Xj5B+ELKbC
4gZrcx+vnwbHTfQ5/hUZawZlTD7uxd4RhN5stpTTcu7Y4amcAUXUjJon2qpG2QbVblcYGWWWkNIG
xcmXKjUtSxiIlQMsceLksciGQmwkv2Yd7b7+ad8AmpCLF3l5S+Xov2IJb2zm9oNMq7q4v4AZfAxL
GblQRQR85G6r48Z3ernJQ8EwfDwI513DsZ4ltmu9ArSEYXBlh1+LU0Kn5rmIauQOXitMVbE+LwUV
uCPoG+Mnsm+2rTGBRlpRjXrt7bQO6x+5NLrAn4IsuVjrel84Yw8lUiMcVzzeFKGr5TownY762Pev
m7cFdl8dmmT0RkYk2pn4by/F76y/hhHEID9+vcp1GHPe80TsZ21RPvduCJgW/yAt9BWM6RT7r9JQ
+MFt4yKDChAR3dJP5sS7iljdm7Qc2Sw6dww2t1WQiDFGstZ3i0UirARW833mIR+F6OkjgIizhH+x
syB+xGdJRy3vGc4uXrkV+T5vcQwRFGFugAj7lMkgYPnldcJ8VDDc3VjxKFPLO276FzG++nVLxAEI
5xGYAXUeL08DQ1qiGIR3RPXGP1FEFK3jr5g3dRLzlpoaSP8xj2qGpJx5bv0rt45SMJj63C9C/gaE
x3S2z+igNnAe4Nvl2kbGgo1LAeHaIRsPJoBJhOmzwiJUMWq/f/snSyay5cPT5O0L5d9gW9UfF4ma
Duk/nsTujOvVx4hJ8Ckob5EnXK5ZlqIsk0vvyzc+OX6fjKyBQaP+MJB1ODKzETexz0I/MCyWxbnO
0TNGEUL49cUDlQxShV1wE6S1TmLzguToArhkSUaw4fEA4E3C6mhi4kDdFpX1frhJ4HmWrSRn0O+U
2HKyhATDmunOn4j/HRVl1jPVm4Vc3X0P2gbBBxkh48d4OAvmJ6vDMj/ak22EBYJl+i/21rfKpeRY
vv6Yufl5KHIdbpLKc995LP3DXe5NgiMFMONc8bonuRdKUxnohSKFh/A5VzrNviNCignU/EidQOf/
t5NxodxRYhxmMF3Ahr8eyyHqO8mVe4oHs8OJ7gVLTRcBRWFwM+bBsqjz7MzLSF4uWb6DJ1noMjNH
2rpecwZcedXh7M2PLkMmtA0gFnJO/vHeORR9tg5TTWjN7KjT/1vIA41BogwGs8C0YyICqcc/epZm
7KQGO4HtCFSiDj553PJWOhEIuE6IInYSTtJB8akoHyqmnlB1FafLLQGSBWMY44ivRgcGnIDGCdsf
5KxoZYDJb/S28ZQaEfvXXUHJKByAkLH1G6ji1v5dLFwmgYAuumWm78mNm51m+TTYcle15Sw1ON3b
MtSATqzaL7s9arlJqVSnvP5QJl5rL6gLbsZNbGlbdUwMkXfdRTMhqkK44pHSDiXcC/Li2fHpYcFe
FPBZKWWZzsWGeZBLbNPYwDGP7kfaqgIJjbTtodD2BKNhYeMCA1g+vwaF9V/EobsaYmu8i2utBTxi
ms7Hi9aOCPq61jhwVki3CtAYsNfLDIotrWXKDU4BQAvY0ibfKOKx7MhMsgYXk/H7ijl5xFTw3dm+
JnKAC3iNZ0VUTnDeuPLVwia7Z+sHb28KpCwNvPDm50n/nijuzK8R6pSku/iEgeVlOmJSHZ1iTHqM
3xFVneWzWvViz5vOpX/3s7NlZrwZ4yFEUewYJyG5CkMyylovyyYmX11nl17XyvFiSY6wpWQGWUgz
GWBCQ8n6xPR80FJLaO6xW/PubIZ6jZKArqTHw6USBlaYfrlP5uUNGwykS1Vpx5DYESLSGQb72HJr
Qo2qZ7TgfcZRq3gzAZL0+u12mRKSh2XsFnX11W0k/otT4y4jgKxlcv0OjPvap9P18E953dLsg5xy
xkdbqZTV5hzWO33F3x5YbIoZxzVWbwM88OK99g2hdoDDyeIdNo5BcI+RIEfyHFb0HXebykbGf+p/
+c3xof6ebdag2rNsVZ3JdfVQEu66Z1OXiYYXRRKFMG8+mx1teBvNdGHCcurjNFJ3fDUkKeq+bLbI
lRtodesoEHOu3v7eKlN/kLtVoThAm+VfwJ8DHPPh2ZjSkzE6EiRBO5syly4jUcqmBrM6RKl5QXnv
dsRxtdHR8MRuCu13bi4dWRPrSOrjh+ftpBUsasIXDrwjSy/BG4ysLrXjMeynarPfwYWEStkN6wIm
Mgz3SbwFCXWQPPm7wd5hIkFK6KBbKydW+dbpE5BkupdYrC5EgFyc9x9Y6t4IeOL9MEVwxRDrPJVP
d41QKdyhPHuv0OqGroMVl/T/tZDFY9Gs5155wwU95m7zlpKqXpfiISjIV3A1a3sGpXJCH/IxXRz/
uWIK/BT+LgnmNz8HE3vfh/6tNhmUpr+HoNuH3Ha8KjaLaXptrTFaMgh2ub+AfR1KkA47X9K01CU/
xQUAndwRO1zd5D58dPMcByQTa5e/6T2RzIZRpvOH9DWypF0BPUCKsjAoytNIfcr0z9pSXFwBLZVq
YYSvN4Zls2/bk/EcWqFemcEpUmR4fSrCbU07gn5ywRblUsfKc8Dyh1oHRVirijeFbXZjYXRXz0NV
2CVP7vhlFDP9hdKQeXe2ZJa2p0HKTzzcgcaQcqunWEBqth1FwknExg59UF1mbSVI5/u7K9I6J7gX
IE7HEMZUOKS8jhh5jMtCvudZGpiDOZCD1n3alu9dh1b5VLtAXLjsTEcYXCe5vXXPuUSF+i7yyY2P
GAgH4Df+nMvAhtM1TV8zV6V9VqIDwwXRwirjdoxZmKC6BIrAOn/AO55wX3JLX83CEB59kDTpBK+U
tEuCsJGW+MtPMifFjUXMFA9u8w65FMgxb3+Am2pIfhMGNKtrZ4qjWyZg60cRKhiQiyGRp+QjzCVj
wbBIlmr/mKTBRh7SgG4fzun/63aptDDVouGRoQKM4HJzulCDAdXpjY0P59s/dhM1d3kttvqhSIEA
QwtFl6GsFx2RQz4tYRbaX/qkkuKyD68LftI95DbbQgWOF6gLg49EtihWMZbFVnHprEPqQ/NS8ZAS
TWxRnu08OVxnmUGe+aEGnVZc0kgXIbhXgteWhdDf04eSt8/WmOmb+wvtvlY1eIxpWDO9ZwYfPIO/
GEturu40j9iY9cLny+994rcsxZbGrnpI7hjDOPsUTEiDH3Q0/r4MXf94pGpdKoT63zfXKyC/hur9
9nauDW4BC4xiTOYFRDV0oW80UHq9lvCTYApijZ+WahSTystQ8uAve/3H/thNeubQH9cmgDwQ9MT/
1Vj0feYq50tXZ43+zCTHQ22TXwmj10jbQ3u9q2Oawqx4wK0+vj5xJ7yIulALUWQvFDotVRdtvSFO
/UJOKr8+DKvUtAykDimtwsGpSOoUEh4M9SkXEUc2jRMP1hylfZpZpwMT36uNIvK6Piaiqm+EcLrJ
k9DqwuUjAjJqlAr0CyQ8mggkDjA/E6VZ051AsJxfEV6HasL92n2DV7hE0gyg7T/JgIJ+Sg5KVwyR
S3ti8s4vdfhbToABlXfI4kip1jliwRJ9Ikbrd0zs7MYFPtj+AaCtyYl84bcwfWzFQO+BnIWjMgtg
iKIMwqpEofwH3Gwf+IM4ngHsKvKJrCY4h1qUSdRL/TpbVSxB/aTyZbveMBb1RONbskCyx1Rv41C3
WC2B2h/u90+4e9y3fb1hJT7cCz+/TeYM9LO7w7oYobTiaPWpUV/IW5NL7ewvHsJlKnW5s0rb4aaX
6jdq2QB4b+zmY8Dy922asQKiCF5GsUNMFes5jAyHlzUKWk6pRYgaYY8IItsUGQH5qYneDYrUtq8f
+jJG//wrF4E+x80DiZvnGxcHWZRESJJ5675hG4LGS/7SWMksTf7FCy/TpCLspf+R200LKSr0yLo5
a4wsUtjcr3I6jR9UYSwcgZB+nrGpjKgCoRHVHo0dpn6pREjzHmUZ01OJboTc6R4KxtSomZWVl25Q
bH7iKIOGeh0gr+pHMnRZ09Z4Z9mNgf27WXoQhjfq2HOJ2f4UbAa/VHtzCIpETinpI11/kwSTQQ+z
nK2YhOdQValuMAJhe7GvAhwRVGpRz07YRPloT2VNhjeV2IASMqMj5/taEYBqQv+rODpdmoEhU8xV
UxdKY9l9btIrqvOactV87RyOzo3otydZK2m18aImGDcOw7DfLXYFe4Rs0y/T2Xy06JDJ1tdW1BoW
z5tHYMJydaTR6oJZ3ce8syYRHTGhUWXD+tV4+L+bERonhy2+IhiT8NqFbmn3VRXnIOK03LwqpN/u
/FcwGI2UpqvTHwWzuWSmxX25ScwXG9of7Yku9+L3Ke3cCsd671Tdd/ToPcCTRbnEl4EHWiPXEd0p
cM50KmiUnhuehGy3oZSsV9fuaEN8FpjRI8BFr3dxHLw+6zDleuZPdSl2VRsN/VVETkv5fQuXc5Q0
SXmxlyVpvf9X0jpe/eku7eUGxDJMZDQIwHtXFBEmSppbrXlFMh9cez0kJ9g6M/fCRCEGBl1QPJFf
ndN9TOF9zfAkz2AjhnuCTna8PnrcZUhWXs0MZPioVCODDNMm5n5RSINmEGDS4acfDTSoPEQQJpXu
Kzi1x/ZhWknfKm+VSs8OvK6mKewf5L7PSwBveGT6JFjry6+unLgA9yL7XgI42ZjFk/34nnFL4+1c
Q5CPHHoFyL2ZoTQZ/Ic0jz8ewdiEoE2pka62d5t7UgnLCT04C0zaOiUwKteuyuROaPyixVVAosN4
mWt6ZrjQGywpjzIrN2GsNn3DsYC1geUNK3UfcvDdsf4zXgK9zd8dxys3Z/W4evXycBe6cU+V5Z8r
uLSK9TRogz6wkaSis2v22XrtWoXwtARMCa98IQiKCzt2ksivddC8vz5LYpjQkS47jGWGEGDqjvzG
ggOcdRC0uGfuE0qHi05rpeMauUnYe89ijHJpiCkj181wDWkptBSuQIRq1TdG4Vc+NIMgoBqWtbRV
LicEJGLDzebnpc05f6r2WSChcY4gIAEDicNraPiZQCDLKBnh0G8HCypC3QUA91NxoBqy+QaRQOmD
8gNNhnYjJPSgAZ+kqbon+jBhNsTLgSv4k4XVgZh/9mHcuJlP6C8HEpDhlWB6UEkbyuOjy/M+qrh8
YOwJ/mFvqGkhx77to0sKAQMeHwwWVTB8ZiLtrxH5fwIMC2OOZaL1fJoW3QHKQ90fNmxXZFl9gLmy
BDnZjTRTtqk4gHFQ0ieWzokhUXy/er/HX1FVAVMBbx8vm+YHSxErmSksDNfPrsV2TNPAI+0c3rwS
kdqKbrnHyck5SC5mcCNUZbenNrthpUOt3yFzpBJsj5zeadGWSbqjtc2RM60GC49BWpbHvUf09klY
ENXed8ery0ZnB6H2cJEUYzaSNHFIAdqyfgTNmAnB4Ya2tE1JqZ7WI8UKQYAHwW/einzMRBGIop0F
LeMSFdzdcLw+fvYMTLQ9yRnjF1BVOdib4Txb/iKZwnQ8/q6IMsOWGWBBc/iEcYul4vHOTYQiyuVP
WyBUr73CV41n8gxfvyQ6Klx+hqWuZAGt7lxK/l98LKpmsRQoNiBcGs3UpAR7hAGiprk2PMfNRuVU
kVfz6rT8S0kHSeHxg+ewDT7uAYkVSsKWWrGZ3PEmeoqIjWiwWwDlHJV+IRqIMEsQucMtn1/EU1SP
1Q3V/POcYci0NjE2GKZjt2t5JpNhEiyLTmxj9xFycemNlg6CzehssECr635nEaA8qcu3jnzqEyE6
wY72tmhFNQU3xb93HS9CpBQR1Oak+AnUgNp+q4OcYNY2xVwM6dD/l883q0vy4Fg0IBwOlIaM47tk
W5oUo2OqgXrCBhiQGA/3AF2fK8fkm5XUlSj6x/14elRLTXdUFkVJaUCPM+y/Jymm1zd/H+cKh0jU
BovfFVTahLHz01F6ZWETR3UoX8O6MWV27dHPElTm4Cq90zY+xVlbGJS77jQrSBc1rxKDc8xOnnf9
iKuKvH4Tu7q4qSKGZVt6imxk8Wc2KVGi+tuo6ph5ktvT97Vqy/zHhD5NOvdSOX32UEba3yEuMdUb
3pyQdbnBU4adDVHdIXgy3cWqTj37h4+pw0lwVCdc4oDXkCo8sLc7LLK374Z8DYlke1Q6kbGS77Bl
AY2GFYcWeeuSLq+4X0CiqnQ/VR8FZBvIe63MCyUUE3dKw6DmTmWIwNdKXd/kvghRGkpz+UHKOYH0
xowP2JYGTxohV/QmM1G2IotUNUZAH9CvtrWBXf/W1fJPs1fXM4aLbQGJUw5AdJR7S33uDyfECn4k
3l1mcfZwNNOa4rFgMQJ/pXiYynVLizZhnurrgAwH7/fFNMdNKxd9uTIEAPO1Y6n/nVJT8E+WBo/h
3jY9DuDhqyuqPECoyOhmxLgJlP535Rn1419hfGF96Yhd8m7KrKHR659oreBsAinlSfGFGhpQGBft
sN208gQECcOaiEkjkzi2c1oGVdQIvRtPED4/UVNhAlS++4w2m54357hs8wd7UtIK3z3MWrSx5HJM
EWCiRdZcw8ky9QumepQGpDgm9HfAarNdnybAYsgIP3WKlzg0ZtgfrEWdeQr4F+r39LTTjOQQskX3
xR5BrNKenR9JxlJ6CBIYo89xsrNHtnoX1H5AqEyGdCov5BrjBs9F+SF5FwXwVgTHAAqgpfbVTWYs
nuB6elLbTYDhbuZpYDWScP6Lb90GhPRFFI/3rPtzaSMykjznwB4EurQFXojCjP22407BsREPXBYU
aLiWC1Alw8Kdd6mrPsOtpsBL2Tb2UN50MobkSlK64Dbpn6Szw3piai4rDdaqkE2wJaII6gj4jzyn
LmtaG5ZHWii/XOK3rQLe98d4mfvvD/xEFqnLYjo6qSSb2doVL/GX8GzaNDx8VdreNa/m3bQMSnWy
wOu5LLtuB3MMZuEqsKjSQwCiX61mOTgKGUtkmq0k4qsaYAjOXtmUGgA3+y+Fo1UcmqvAp35m3u/6
GyTGCb2x4x8/354lLAoqG3PDcq8+dVPr9h9vzXxA0mr8T0FSZrABTyNhP34xd4S9cFxLATMDPesp
uzySCeQUpARIBmxCZk8DdsKqZiEsS++nALYoMEgDoPXff3rBHCY9C2UFwv2vuKcFv3P0JUpZPLaH
cN+Qw1xpGcnxKBF+mWELmdU+Ew+YuJMZ/mZi+A290Hdcxh5mrSviRSED3dYUC+MBwDQZtBOzg7X5
C8qCZJYwYMT+ubY6/Elk4UWgYcXucrH9aSXKjBue/AksrNMVhpydk23h0qyTHzlR2cniaYwFSnP5
pToaUYH0Rxz2A6c5qFwroMgq5r1fWlM/tqtd4M4Cnr1S4PDT5J1qDnFIYI1AbVdJluluEJMcKu2Q
Lr85urE3v2GM/NkSafS24il5tAR/+at5NyI1alO7gURg0wkkRW31f9l3I8klxYWZWAjFAqxfwZdP
vbd9ipIhTqrnV4tZQ/tf3RaXlgYnuzoZRFE006YryrY6icjETF/16OWqc8te49ge97dND00mAfGi
FVSorl8exL3XQkqWM7bobObTccVYl8q0UKUGrMnlL2dN1JcNlQga9P0ve9Og0uzThMRni8cgaQeC
ta4poQzzZYEml+s58SQt+z7hXFF7D+fUohK86TkrJy9Yo9K7Rxvf2Yh1BQWtseIDDC0TocueMKAD
vMXm+7+1xPqqSLySYnQ2kqgB5Ufeoy+7e44MbPbgtHDOYfq9voco+EPp37Z4R8D58oW4TdSH+t+V
wGsrdP1uAWtHmEZjOp7IHyBX5bSbN7wWgLvdX2nroftRYAfeXLWzo/a1uwxRjZOZiBBQrqbqrb2K
nrMf+qNBHpaATd8KVn0wuu4cuGrBUEaHvJfyA2yllMYc5Mu7dRAvfTe1ogsql5GjCTa87NCqJyBb
po83N3xHcQEl2FQZduFYPRCLNI918ZPO2/VNE+rni0o9+dwdMJRA3LvzUYGlQV4AzFpWgIax6Irx
C15PHEf7E+xEFwG1y74hTzJu1+kJJXiUhIjolnWIOiSNUYFFB0KJnZBECt5R5d5Wa84YcHjTT5bQ
pU4rw73gU4tVeVO/wWmZtN1NBRBWhhfFtIsVdXyrDBQtLQGz+lIhYbgHTWJZKFtnXI/lKg5FUkGG
9XVrgrCGBQ+S1v2E39Q1FW0HB+SFbK3PWkzqJz1mElUGXiUyExOa7KFvR8/gtHSeS3sEzdnLY91k
EsEZXIWsPt8xG3ksTYB/xkxf1Khon/hTr4H5hfYtY1VuVCRj7AkHGfHTJaT4YduDqt6hWvMjdcj8
ibclgvcFqqgk+J24G80ajbF+LHuZgizUx084Z3uR3FOXTIFBU/righcX4i9D2GZXbk8Se4wglXnL
ltJcfL/XV0CZw9RSo5l7Q3/yCLFRcxzf686LfO0IhyYQghKJf9iyAHhGkzaQcf+tOvsb2BDSUMag
CihdsBviaLfsdev4602ZNdZmdzYJUvXdgLb7bgj+UkRzTLvWEqYP1kDCPV/znm2drYnk7qEYIbJ3
eXTq32Wt3jY7IOqz45tkA7SZ7RQPtmb2OcqFFpy/n736wGA1t8P7JfZsqXdufvcoK+zwKiq0RGdu
liDt89MfHMT5F59rs1sdISCY2xgAaiItkDm4ty7soWx3/GaiTHeyqx3DzrlYllID4GkAmKByiN8k
8TmvAsYBfgEjfZHgxR+OigBzks29ye09nA7OtAk67v/p4B22LxwBNaDcx7K5yHCvA9i5/YPeLgzG
o3qQFqomXwUtZtgRC6DU+RkNlk/GePjTqOJKafKhhzt2ydfoaG7222NcNSmcTCoFsIepcYH0SUnP
N/KnqI3Q3gWoN3/9piUNYp+ELy8EYw3u25ira4h5zVaEE13wu0vdi3RGpf38Iyra2zuzQTZQ6vjF
+aqFB+9Hd+KXzSVKztZ6B6GK1agzWbyiZ0KJam1ObgfjOPlb84Upqwz723ldmG9SojDyjcEo7hiK
agUtzUcylJDfhB295/QSyriyMHpUhkvAPucEo0fhTYfnldaLv5sOwB7vKbfsAPlLHRzv5mJoTORs
1gpxCgDt/DwC78k1qoUM45N4HrJM7vqN7OMavxkph8aOeaeLg6bR69D2lSznOvylc5tL33DneBLG
KQYVxHb/BI2JAnOWTi/Z1JNHjKC9AeDL7tRm/Cw4/Co6O+TwAWEPhOCMHz3503wLeq/VV//EriBk
tU4114mXXVDUGL3HNvLGXBEob6KpjLhAsGiV7jHrzcYCGcj5hFBLwQiGap2h1T0Jcb078wLTjeUC
WDqPBQ2dEBRUbVTtNd/VrDjuY7RSmzhXy0/2ymTLgAZSvFPw43/WLd5VGy0pAkFVfvKG+Zadb25P
uZIAKCgWqnHziOg05AnwsS/DWTsCaJ/SC9RJsPqCilTXKEGF5JUIXUYfQ6/UQccqd/CZAcgxXWpb
dvToo3jC3ifK83NCKrKrRMlnsSKCnh+BIUqVlpE2nfKUcrZ3SpSSbzoh68z6RpXSAse/aAZjd7rg
O3NFxbX1TtBJykMm+W6k/GdMKnzZUs9muZ04pQ/MeYPgUJGS78B13HhMAwy1xktjGazM3k25gofo
gDq2B5lC0EoqeyKtFP04vK5GSGjzvxGCeAlBabVLFcD6t63rAp+6lKe9Cr/ASB17LO6QrG5aAPe9
RoZLLetFS15qrA7fyqYY0q4bXJ2jLCpH+tSQYtjaRL0u39oY4q4CanrOMY2zvjyInXzyPPU44JAI
a4O19vLvL5Dr0p0xaDucng0pGcuihbjSpUamjpACOgeogbg7ocQ2sBJCxZ4PIQezSakekulRHhGr
q3M+Qr+M/auzGrGSDDVIAqxTla29E1/EONTjHkssXLNjACjTV6LaTUgn9VK+CrnV2yfK4VpqVzRH
3sfzQw8tPvFkCx3qoAv63/1Jgj570vWhSqVM2fVbVKcv9gwXoIVgu6V7cKLQAIPgJdeB1t9FEa7W
K5lbgSRSpIhdQNxak2ojh+9HtDfltTnA0QQh/uizSqUZ9IA+PSGLHA2/s6Tdw5Lh8cCR23kQvJWX
QdYL/FWIp+A0XfMODXK2362MBlCc8PX7cVObCuUeTljjG/FiPrROWD2dph6cuKsi0hAyTP8S7nyw
Ji35GhVFRFuMQz1zS4rcVUp/ye7CcAfOG4mad0A6QRLdfPX2pdWxReOztMVAZwaqVBQKK2fCawxD
pezS2B3Eti+bWBuaEtyY7b2B4Q0Ph+7//6B0oRnYCK7V7PHcoEY8em9GWKST6IvHpPIdnUXBC9OI
ltzoOGPCmeA1cRqrkcmpBhLcmLsWNJb8HS/NiXT5sHU5arI2e4mr6pRbI3IwCW9IPd4bnAjpywEs
yZGEZqWADCj6Cf8CGnHpKuf05FOQBqEVcQIKNjKbhhv4BHEAV8pAluW+8EbvT1arPJXcX37Fk8X2
GlnSpLBqnlDHfcwH53XCvCdDcQV34fe4IEcSiNDpPMp8+jWxImnH08bTljMPz7GN5r3rD2+JUE42
sWph0BxIMbw1XeScLbzEZdiGfIytwbQjimtIjWx5XhprW23IYmaCY74vDoRHGQbvFP737MKaA3KE
nCFytoRwX20n9Y9M+b6EMhUTYvSFjvhHDyVKOR7jljjQNS1Rty2VwngKTv2vPfHYFcecH1KPYUTf
dw+cNdfZefI1c1MoG1szJFIVIrCVy7BG7I2RhVnsezGkYJE+6Am2f+PJdvET2gpUas4ul/fFtP1L
CvBM7pZw24NSJDFYLyrH3Y0JT6Oxh5xFv80H/b0HEUwO1cdk7832jZxysIWWSfJQpYbqLR6fy/8+
c5LGb0rQ6n1vTIg7fJ2NDOfxPyYvMp6llF7GFT/RHXDgGg6+mHYkwE8V4u5BPK52+DiinEjW8zJL
DJCIIWpP0EZv4mgo6AjUcWYND9LUrc3h9lvZhFIH8MxCqjSN+GCwO85J1IxRYjgfwBtbaaZVWnSo
gsbTVNqzcKUj/f6+i6czVCNDN/d0+0A+9wVwuJ5ZQKyn0z3ObPOWiUJ8Yic4DLLQMTleguggvW+H
37Nk0jTZNkILzE7gVz45RClTRkPT8VcBRMYqSroxI40R1k7Z77QXfABYMCwhM82m11WYXOmoODcR
GkvLhzT2DvWNAS2wkb/cs7YMGzKbRKfs/wO7bynd5SxidcmlB17YlFeUwsDMULS3wvtIVvir5TNp
V52zB8jL0WdxXogOKrFhvyFkmJ5x5BvCv9bDJiYEWQkHJTLE4F/OW9n7y3pw/ZgQBVm/mKVw+3cp
nvo677Zsgoc/mj3rrR4HBvmfGmlnylfmwNMnZiZNOxISINbKaEwxPlXsd+GC8jwC01Jq7Lq6scKc
Qdh3B5xZcnRxFp1xMWLA7C2QXsX6X0DdHfa/sO1bHOqCNBSW2uNvyyzXxZplcJf8pnpIWyXagaY0
bf4yVTBdH7kgx2m3Oj6DY2H0cGd//Y4jHYbeYMiuWAH9HwXaJGb94otFw6u8KrRUE85fmbS7DRQX
pbC/74OU3qMAzPQZB4gMui0pfJIGRO7nDWz/evEIG9JfTKung0wmwISJP82P3O3IqntCfM1Snc53
HSnGnFlX6uvbW4jnuPaAzqNuhCSEVVlu3obGQDvRAd8nrJ/p7uhTdHR6tB5TVIyDo/tpeDkOKFSq
AaPK/zjprBrO7iWcQCJlZ38bVa6tCYfn3MhLWFo75aJ8jv9kqTDRWwdKYkc1xV314jrQTZ49aprL
PtdCeaCZn8n1wleMSnB768aUruq6slAebkd3dTghwuWiN/QhJB/TuJKB2PLjQMYq/sY71jyOameg
SqIIbDQrnlBUWkJdbTu1GT7jYRRaJyljiwfvvpMBQjGSiRa/h9tLul+BlPkgOIwLTTA7qs1Axx4y
IP5+tH2kdPqaTG4c4DXd4dcrDwfMiwS9ASlVSNaM12F0vdCDAnANWbwWuiYz5Jebl2NefGHoLGBh
sM7ScQgO69O0nsX0BGB9eCf7zQbtqCWp2sCl5FG25kIo42ehet7d9bewXo5np3/av02jpB6NRbiO
AlDQaQKnG9BMePaLwnppKKOCBNeX210HWOSyflPRgHOwAXHaKFhS+dv7HeOyn6l8J16wwBNPf9j3
ZrRlFfLpHxP+0y30x8rL6P6ZUtgdyY3VMHWCoQ9rjEVgn/WgTOSVHCZ0mYp3uwSxwaBT7QhOEBn1
/9FJIDnJRI/P4TYRwtsKeEI2T4zwNSUlBNx/2LKViIQ18jTf7f7A3XhvopOldoT+rQQrkQwNB0r5
Ie88dxr1J6leRAiOKxhIpqT2ZRowxbo//Wdu5ZFnsnmQay9KLFeRx82eo1SjTsR0fxFuLgNIpdF2
I8w/ijJ3lARHfeXTzABnsUWnoPyTwtLqyYU9YA8ns1bDp5JLnQzw6qDVhBXCVPVARk8/UTlYGjxO
DDbn8NrXug6tchNJxhXDFo9z2kixE8veik/JwzZtkMIedLqb1bo3Z9FZXKOtO7eXoL1XH7404Tmt
js6pODFXR+vpjZMaF5e0kLJ9phnLkz2WKfQP6ooZ5V+q4l7gUU7oiipD5Zz6qJWzyTyMDkSLvsNq
tY4re2GdHt4ah0qwa1+WWgPXObGc5b4NF+4WV2DbnvKI0KMXt8tRRvIy9ToYZUrAhBwESIMBA/+1
amH5c4skA8Oe0I/hkGMzSAlRfMoceOVvd4py3RiIUGu3n2UWC+30i7Cv0IfJtu8zdqxYEmkryKcO
JEGtaRtybNj/T0cFPCt2dS3mL8pw6EqjeQzxh2S1BrYAFTHWG+bA1DeiokYDeJIW8HSdaoNidJle
quQeN7+oaPaeKFpjVS7TJkcn8fgiAYJgkfQf/EJG8hKRuuJ2sdpa/UmjEuhZ87S+tucdGogNM1DV
GWW9HPW0y8TS5/FMcy/sVQt527WDp6GpZYFLOgzuOVa5FYqDb6MHIETlLZOFe924aGObFIdJ3Pbh
pXD7mOfE4tvk9xeP4H5tJZlV/WT6Z48LOrj8A+C/3PPTAzyUCw0rlGHnwl5W9uu1XqLu/8vgELxZ
fbeULbKYTYbILpfr2isNlMrgOedwP8Vl5puaxmHrT4V9DhN5WjBB3bD/Ht9+5YwzGhF8vv7x1dEm
JEwiAee6USvgTuno8zR5ptLsANv7fiHgXGye8J8XIbDyFuKXiV+4ou3ELXYtK2i3HlXkZVLpaqcr
nKMGe/W6oi5v2gL67JBBq1nCU+LwsHq+uu7o9ccvkY9XCHi/WjNi43vDM5sRYgA2WZeCraLZXrg0
W0h+i8hUvTnz3RTVXZF6Dk5GKcWOVGmYkscpXCNMPJZ/StxEKdbTdhT6UlERB1vVlH1aDYOvQvV4
gam1a2JaFpt7ldU8a+gdEgLdG6orexYD6JNm0yeXYmtg2hp5ou3qX2ABXddhohbJWSVRO7PzKrtW
E1zhZz3XlKxCISMNt87zFt6eIkyE9pDWlR9vE/0ateeDQhULubBifPOvdobGf6XiMeGk5nELks4w
OgnaktgzIT738jmPSIXdNikE3iHInA3mPp4ZluIX8jE0SW0c89cgnXDA3YNa3nYe9vnUDabKCTij
f/0y3955dxdiUlx/tBGET8PgHbLnSOdokGQhf8+oLDGV62N7JnXDR+M9IA0TIm2f6CPmL8KawkS4
5v8Ssbmd1XBbQU+FQ72qf2mSAQFOQnFVI/m07W3+2lRU5TTxqNbkPUy1UTV7HXfjRqzRro/r0Fab
XTCuyA5ozXx9JS0xl2tnfa/7tl3w1up3FtbfAVeU899OY2GzOy/4BsRuRFLU/ZMsj7HEA6LPQ/I4
H4SFHYz/xvVNin1MigftFQLnsuJz5kkI9O7UVfWF2oeXBmkkFMi5ZI1yvJsJ0NBiAEYeB4oXH2on
u4rtkDP8NQ3G3HdpANwzgeBdoNfLZTXfAw0aaNqgYG6wQxCFcIsEYmN+bYsOTJ1HxSFr1b9y99nG
8ohebdXUpSb1vuW6MQ6mJHo51W4vPZZkRnMqeK28pQX3ZvuwXKbs0eCBLwOwKgdtO3FonzQuJXam
NTPO2teMemqmeG6FPc8G7i0QCyr5QOKCCMYrxJ4qhT5xm2XyF5MpXHENI+csYWrU94V3BJpY/GYD
+IlWIY6cr2EKk76t+7qvH/o3HEPdNF3RfatZu5vHT7a+ZC3HeduroakWY7Ntplha1jznS74ZNami
8N4Bp8nZModzbEXLHw3tJYXgphNj4gs3Brm39+Ly5sUVI+fK4/u/8imlpZxJE9VLkftx0G17eNv7
VEWtymrTGDT1rq7iZS1vYc7KRy277yJvPRBVSsGJ6SQrxQc9WFMhJXevsjyl64vS6r+NrJcsgzMg
yp4TkEU6VEq1sKP7xUkTK92xVPPUs2yaZ8oXcQXJ8CKYU2kRpTJnTzmCZ04KpLOFIe7qAiAorbuM
WTQVr3IR/sz/46Y7rhRI1/J+n/S14P4ro859W/CjZwex8VzYBmDq3NygzAsFWMOLolbXuxQdch6X
jojrSxVUx3h0OfUDKO9DK6EvfB9y0QTFPiHasku+PDZP6zDuJf+zCI7QkBlkeQR4RatXP74D65ln
wIxzQSq9LfUzBH21dZApnVMIA8ibSMHg4iCZtGH8yF1xg4allX9sUiN6rXnv7UtiLSRRkoHo92j7
D8JX4U0WRXzt/pviw23Hgz4AmsXjckxj1dLQa+9Y+cd0rFAyE/5dmjqGo9+iFf7c4aurIcGRRPGL
PGcc8zH1nKO0XjB4B0lRc49bnLmIOo3t2XxLQ+OMCH5a67BIjjTJ9mFdfBMJLBoKBEtJCjWWDBrX
SGNnwRNNvTz4lH3QLx3nByAcHGIYMcRdusnbV+iyCqmHj6UQ8YqPX2Qpko4xfohEg9h8Lh3HtUC3
NNcwPLdchfeDmfETcr3HG7uAHxjT64GD9pmvSPGhk2yewacQbp3rAMKBxfcc+rnRBO9zfIyvPrb8
leZ60+vS7pg2qZtedN2lQBIgBpg6J+Tf/2ePR7ZA14EbTMc2I6N1Q3KsaT4tsHpBd79P3ZkLhHYb
uMUe0J1baENpNYudDNyPJgczvzhSaFz+EwjaxhWqUqnCoMNr2YXlkupdpPFeLvvzlVtTxSnUr2u9
LvJGMBlFNvohA9sxwpIywoAPkqWRhpVD0LJVStLEmKsRreMYHx24BgCEL+H136OQEKMIf3vLK/of
7dAC5S4GdFfNtRFHbbpVavjyQIHiIQrNv7xknjxblrdVKY10AVZtETcHhYiNeHOMOUyRWr2p5U1g
uVq0s1zWVufH0IUs3ogSw0/UZ1L/Q8moT1KZAvEATpFfqp0Bl9Rxtq+Rft+9cQGOIHGmSUmNCaPb
rFPuokJHDI3RScK6XD+tCYVobWm+fFAodKGP6CvE9YILbkhMgITnDJDP6M3R9/CDdMqfFL4HfY8U
NHiRRfeFdI1XWUNiDu0YIj+Y+v5V6kVEGnmB1Z6GCORk+eNE7lNoWZ7/Ox5vONeL071L+ujMAHEL
htJY5BpyI7LDaZqoDNW5uxBWzxU27Zoj9PaZ4JHFwsyVUaWy5KxWkhlGDfZXURMkfwI0hzBu/M4A
RXX560a9Pg/72s5aLUTFPuS4R7KmnkoD+/qnwzpylvXgN8dmUPxOFfSK4TcijsmKTgqSE/ZJYICq
wj9aksvxbCF8geOPAZ81WaY9DtFTAHMDchbp6JSyge583iKEJnrwvHYUtnmqTEI+vMvCXxF+1HB+
IMvZ8Ojdp7kasgdotg4oo15igTCmMtmwdAkmfM/dht9Pu5oKWgnoM/akq9rWURp00eJH9P0W/U37
oNDaZNdhdnNd7R0li3pbx8AkXiI616EwAwlbKB9xVihKYSwuYeVjWzprKROtJ3HRsT1B7VwzJUL+
OE9PakRXQKelD7zUb4sYEVI8Bo1estDskB8avnGH3sx9zjWLg0GoEZ7uvKUYHjnW5acNAQaDrQfa
jdt/q2lmMsNXxSEEUVLYrQ8azard+Z6bSjc8VAs1Yf3APSJ8fs5Dem6KiRk84NhS+zQi2PMEnyqE
MOe3GwvuR4ATk9Si8l1rrFH8pADjMgc8usuUjS3kEaS5A0S1wFxbHvME1NWPZgt61FsPLb0/JcGr
H3HkmqLmE60O0UmeMJcdL20weJWEODVCUo3mepMXzxicApx1zd1IpoYgL8hsLeZEFTHBMHqXkK8f
eAfHDpRhbQr/RTi2aa/04GENR0NUiExB7zsXHV9aSbPl+Q9xFfR0KgRGILaxFmnh2WCwJod8jqHn
kZhZBZ49GrNnMbevAFA1uGSFYcQb52m9NWVpjQ9tuyiLG8egI8PnUIPTJskq4OqxTQqZeuhaTW2r
aOfkmXnB2pNBQfui80lj3L4xmkFcjNpNMr5gMD59KfDkPozIoQboUWOHlD2r1LYe3xgno0eqvOgY
7UG+IldInUHuehc7l5SFnxiOPXVY+SQcYapDDKV+MX3cAQTCrJOwhvDrzOzZJMYUaqtZGOmjEk94
HgeW5D5b55Mep5Uio3vImdpkTVH2PkiZS3dQkbshG58UuvHse8Hx9A899V1iTgNNGhyilK+2mpbU
YZANaQbEfdu3r6SpK+XXoJlewB91o5glfrPOjK6x3Va/e3FaT7boOHb8k29fjF+/G7ZanABjZ2/B
Y+QpP388GvYOa7GqOoWWBteT8m+2m3bHXELKYU2f3laaEHeoApIaowkrIW2Lm2UJrCCAs1cv+geh
kQ9obJxX90+tZY0mPA4ciHy0xK7jim/jf9/YXDFPtnuacDUFGTe/tV8qfVx+BiyVzf2ZFumq/lQp
A1kL1UbQgQbQcRA4zFriG4zCg6g1lOYnmleWRmzUCPjoNSBuNwpog8w3Y6TK45Evcnc3ghrT1Q3e
V+zgB+nlok2r3TRNyQif7+XzFc+mTchAe9xDGPEXpNH6/hU0XidqNXJ6qO1pp4IE9ZlBJaToYnN4
H+RCJq93SpIwIEh6WO17GJOx/mTYxNbItrqxaEJnMN3UYfJjJCiRHCkNn2IzqMGQYWjzfRGfLhFL
Mg8WyLx9oXKscyfjA/FC8NSsndHyrzXMCzwiq9fLXb4Iikf/MASWfqCYLUVU2edTh7XvoqvV1hQa
KuMi2AtnjLgXRJtxfdmgPDA4RkHwD2VEidI7w5ry2dqE03Kyto+ngHOkVqchpG5FK2hMTnac/HML
etkTQRc2Zse8BMCNbAmtsTKs5BXM9NPVJpY4TWwUw4dM/NUq1kXzvXKAoVRJboAXnzQrs+WbFH2p
TRsgy0wedOg4WXEIB31s45c2n7muArD40H22qWJ959ybQWLGeDv3TZVQ14ENLQ/sdWYPFb922M5z
lhnBTSkGvyKqZSTP2JqgI+HRLUZ2y4cmsTb+WYWcdV4tON9bf3L3sXpZFkC25n8OcA4wF5oQ67xa
bRzU7czg1egVJ3RpvME2pwlhm7VSP2jrvCmr4w1VLPgm8D3OsmnykJhHnfTFrXCd2NnMKSxzZ3UM
wiop7Lpx0pwVoITIxAmauKUHx5ye8XXc+2TpvDjj9etUD7X3wgxApJ/p+pHuK0kkv447urp4oar3
FXr2Y8YKtFb1tq/mlRE38+daA1cHXMLXLvnPAK7HcTzmE7VLI8Wx38HDjRQohQYFbpNnwPVZS50Z
+7amNjeQ/Fn5RE23mwPdT6AVLPq2tDTVLVF7KtQR0r2JhtO+4pXsgPvclq1BjQ5Vyjl7sOvUthxQ
oCbQQNI1loP4uI32IgdVeiMQ5C8mJPZ2sa1Qn6YiKBKsHvZt8BbnuvPM5lcg1E7In0zHw7FXXD2Z
Yj2gaDxX1Td2k5+kK81MQubXlY7aHeBaBw6afckIeoxEQaBXBbUNFQh5GZTxz7vR3N2fwlCWyQCK
slXXqAabMIwOMrFoDomS2MkHYjnejIIBw+vE1ePLG3luxKM+Gf+JkJg8ndWnwvvhA6KW+BcXQsMp
AgChL9xv7QRjMlr+sr4TrRcS/PYg53bgZHdAPslgeFElmmJnDnlYEIHzqk/kFmzdDN/YKJP9Haix
m0KBaTX+Y/PwAnj1aiuaw7hVXtguU7L2ntDs9U/yJDlEqZnmpPodxoVhmy5JTtpa65G7Ye2XvlRW
U36pvZx0WmlSrOo23BUDj2cIrkP2eLUPiURZYiYAKJprFVusY5ueCoDfTBzbl510HtdQo+RECdJi
PsMSwbVzXo99hYbeSGnUXcG7s55HwiXJ5ITIwjDt4jtR3MtFk7/oC8SpSBrQzR4iw5B7YN2zcmRI
erfPqoay1kxBA2MzUoSMCDY4LDuc1QwC0cysfDIxY6aXpRzSgHXA0QxdRfiN2Bn3ArCxJy49r/Gh
1Y2KronGjsydZDIEX83zgxLUxumPiDqlhS5UC7B+JOgS2Mu6xFzdGMgBmlxgIgHP4JwbCvRkQM6w
Hw6r7pW1ob31yAo4dCQRJ69rXGfwhzcPP0GNCOHBmEjwa+mJI32khJpjksMt9mY8rmSb41opBRYk
60qzW8HENBg4jrnaJ/71y2iZAbDdG4Ya1Q5kW89Pduq9ZVPSiKP9a1Dozt1YRwPHiT4inAZdWJRY
8k7WRe74CFoLi4INBViH57A4qrbY4hWY2trB9bLOAaaK0SAzLIpivnvxB7uQpcn4ks38ruTKpYwu
v5B+uLp6qxIwDAbHB2JT8F0cVcyO7+aEyx53x6Vye9kqIeXni9Wk1K3MsxZbS6qgfnA622AQwh80
HNLBKTILhjyLdBMyr2rM4FExuLktvFUpO2Eaqm8yPo4usAGxB3Rd8HRv+kcDmbvS7r9USbgahQg2
NuN0w2A/pLyD07m/QjP++ETTrHbqqTM7J6KuhEsEY5/vqxsCmGlRZgjfNGI9M9DgRIPHkQZT6jpO
lP9+8AJ3RJq6VomBJSAxyjJpu6hq+x0GXPS52QNdhyZiaTBgoL67aBf8pwqJmyRoNELOack5NIDz
ACq7Hoy72DdSj5rj9M+yK4aowqTri2WQcZEtzkj4mCXdUfZG6G6+LDVYV88ZtPYQYRQyBg0RgVlt
5o0T+qb04f3j8Rsjgp5PuaCF6CaT40GG9hpwNLSo/oSrb/1IH+jzs7i/B6mzyVWSneAaCsHKkVS8
czk6oCUuTPadGlV32WYKPQGOT1QkB8szPK6BJXSs+ckz3BXjxvp7lE1has6y02SvmNejf1iV7jeK
KwKeH/KmYPbHSzg0FI0a7DH94jnOpfXU1QqbfTtEgqV2zYMXBTbMlD3jLaujnieWOrDgQvb/Ql2+
ir0qyIs+ApQiFc50iB9Dj2wWXa3RYFV18z/7/hJYYKJhYIkS3hGqFCLyu2t33JE9A0t4CLyiJh4B
du4Veo6bNqVigcSsKlviZIQ5rr0gtsJ2Q413NqCO7sdhk4PE43STO0VNUO5uskWgboJOiu9ULUhx
LJv/d//HKkXSfEY1g2CsZlhXn98pbpO2RFclvxiriQQBNPhLURGEHsSmXaWosjKYBerkZL2gwxIp
lDyXPVMepSJzMcEFjMFwFoVfUTbZcfsb6C2elP0vwIh5uapTP8nW8CCeU4e0ZlO4j9QZnelsFv7E
lraKU/xjlX9zaSeq738ubKNiSiiDsieO7HzNm3xu02vAMYNyKGcMxUwO59akSVEDQoYMHm5dWDoe
Lo4SMWQaw9QTFO767ZmTps6RBOkSPrwF/9liTVEQQ/9t3gVanQD7/NKVjVapUkiGj2Z96WokZICc
k8b48gFVuwwF00CfR7jMYhrHBsMO1ftJMICJ9AX8ml+F442F9OlK2S8nu0N30p6UNR9jkqxIVl8b
ktVkEOYtfF6fATSMti0R5WaOKOBgZwvevPx5H2eeqh42psrrNptpT/9i0c/7w6ROt47fD1MZkrWN
QKEqPBF4XfBhtxIEJ09nu9Xg21LKXOSY3VKxy6JhNv+ql0EgmWTb9uEcVvVqac7UYYVMMwylCN0O
XsE8wvyEMuWbDVfzaau6m6eoRb1Hf8+XtNg1T+ZO0wJxEVnBvXwwQHyFTZK8NYhud9ofvbgF24NO
SRk7qBIJHouhJ/Wqodzlxx1W0ysZjv9ZXCCaslkceWmY64yl+mmOZg32KGLV5IaEQ1Pmy0RF8Lg2
wii+n6a6zOkZk34mK3V3rthIvSPOIlb6ASFxKR5UUlGqatS7hf5rP+HhhvVvKy3nKHNHmLxFswlD
TdsD5SMPt2uZ2ZPYjwldWBD7lp3RZZrOochGQTHCO0mSdrcsNWuRpRuJWuVCCnbpdzuyWDd6+8V3
uBokvBb3x/9bxLAARcVt+oztiMQZooretrmLhOAd7pcEEH4R4vWxiU6ADHNGo8fvuWkUEf7SddWE
PSp69aF/ojQjXpOj/OelVY7gCcxHYmGjJCN3Mu+25njdRGB8R+VGieTrEl1p/zb+HGoSMOt15mke
MEVl0CJ5hMIWapmU6LAgot9bn5gEMATjbxV7qa7U4/eObTrLfcWdtRlArAXKcxrGIhxilWJPAezr
LZcUWIiYM4EQ3rnh+7ytQIMq4dpQACgb2XLNQo+7AXm5OB/S99DCEVf8mQGzjbBkq8pnKSYSIHw+
Y2IJfRkRerhV0Ep67hjPHqLWeB3ndhxnAwR5Sy2JE+H+kyLsYDyw3HYSsSitR720ffyChHW8FiL2
4QLV9/ox6XO+n9jyPLgrQQmF1kw2c/sUIgz7PJRbz94358jEVNlBo6P9Xoui1D734UoQYaKt06gn
dOYdCYgq1A2TxPL+6Sc+93YK5thBQ0qRSlX+EGHjYaBxDSbf3HRy6psCEam0bwiBTBgyeihf3Jzd
gsJYehqnyjo6DonpMmuckdiidKOdTcMefWMVAsKuchdROBerPdZdfHb/yLT1Yd/0NUEmvIqi+U5k
RfzB30LlZm9RI9OtQ26SUyjSOJNWp+gqLVPwzZExAMx5ahktMV5jIqnJEuxsGIq87q4leHvMzV8V
CBU5mIAGj2k3d6//2y1QUZseFX21n3AsRAHXVM8+WHlvgCWMdzooJ0BrAihTNhIJvPW+MDzhi5EZ
H575JO3Tiil7p+WcNk8RrVlnr9UYynH0wW4teukcSlCYjviI50WdtOsonqHl0954/nOAqrzocKFl
6QLkNXLUTB6h+HVGf6bzdqKRxOPmZ//HoE3/33RJDne63VhLkkcGLOMndKXjNMu2JCRHIwAAKKlT
VYbbwZoGuoJcXVCwYvr7YpoeOZB4M5V7FUPUGc69X4CFf1FyMlfUvFhW28tF4sIqCL8ngY8tWXOz
Au7Je6PE9DOrG6WpMNPkejJacnm3vQMGfmL2y5/+AWreQKBDxIor6IFOti+vutd+L9YzuD6YdRmP
3/mvJkuAdbIMNU3p8PKFP6LiDVkCL6Z5Xa/6jteS8on5h/wcW9JAEK3shAxEJz5TTuai58ojWPxq
lcE1rFdNTeT1T+jC+bPJ1//nbjkhZ5g/LiLyVRE2XCCZZNq7acvoWRz5FCchQwaxxNp2Td5Wedmj
a/OAFZ9wyOAJv/GbWXTPRJJE1bpxS2Rdn5dsylIlWpYJqU8jLo+1rGMYFl2Vq80iR8CdpSPg/4nw
Dr5di1ylj2OGnN9QbNTmbOuhLWThRCyga5CpgUIelR6qGvWBkzJ8Z3+JEoSuD1OxIUsprivnVjHw
NHuOaIheRccNR4gw+WOcda5cd3vHGo3+2UMWE1Q8CNoCX8ysB3Za6Ys/pjrpU1X0NUK4F3LY94HS
XiPUjsa4gLKYZdMOaLuDvOYw9/y0yUt4/RtjDomztpUvXHdDFjUD1fNKaSu8kjL9peW5VnYgiGuI
KMXzaDXl9CWSr9BnGwCjUEs8x4Ka7Zjdp7OayS+pDOnmUAVwPn7pOmonKvnHrs52F18ciFTMg9vf
8Bmfw0OZwb7YbbL3CZeB0KBIMD8Ukb87hO+dSlz9yabx5ZPSuzGhh8qgbUPfUeKDJ+CIIb0GbPO1
c+Jw+GikKdPrJUQhD/h8ZCUJw3N+ms658Ev6AYdNoZkTUsqGoL/i6G/MFoppOFcr6qz+VvaB8t9i
P4sImZ99IxD60xBW7JmEXVHKWYRG78mR9K+0hoX/prs2RRDJSQXnMd/sOMH5Y6qDoAvQeUk/OSrv
qlIIMYgnyI7nOwgZhOJjYP/54Lz7JeLjZcnO8ebbZB/3uRTZij2DfL99A0d3vz+eGKrDaQijSyLx
jKTK6u7sGwTL1qq//5MLKyvelFKzPyJoEpAz/wNlKrgCkgLShg3Lg4k4QXX35dVYs7iI7CDT6l+W
mI9H4kyelzldfSKHw7KFAXwPnCYMla4CSTlD9Bh1oayBSHLqwVGy0dHL/A2nuijZjc1OUrxFzHU8
RVHvgZYMtEt+OvGaSA8/fK9nvDW2CW0gH+aGHSjxGrJRkTddjVntyKDFXy6DNFG0H+qpNPsUo1fF
eENfMkRVQrS9PIHLQcSRO5RJAgen/XFHMpeyhflqNyY6sTG2fv/2+AeWZqmSWGs59DzuQR7gu5Gj
wslmEYmux2xBwwNxEIXBG3jrl0VzkjJDDaLYI/aSktNxGVYxGYX+C4uDmRqunSKfjFdruOETp/Dt
HCH1bYujNqt9FzcSPSaIbywfE8nth096fxEdeu3ikJrAaAE+2TVMam3T6XiWeV2m/A6xu/7bMWZm
9V4+xgEzjQ3To1bCE9EEbuFwf1xRV6wzc/mkSSyOb1Kn36io2cRyF2nDBkgOiaPyK+a79eTZu6vA
PVbqs3jEZmCuRfRb6V/nrGdshKrcsGDsE+7rEswvFIwpgsE33NkWz7Lo/Ncwz/PZLNsuiwYwf02s
IvZVCD3qB2oiQLlzALd4xg6nSL5dETwg25cLAe2vtSWQT0PPZrC0FadhuiWmfUbXt7NfMkcSPKVc
SOQOKNxpYCe99BN2hsf6Pw5Lsk4wduk3zaia+/k+1GiBpMk8cMYkZOHSlCzlvqVr7oqj5XBi2tbQ
OwNUYsxNdYhn3oXfaWdbOj4EodrZQR6BucGgcDIQ5ApspZa2TTds7SKCJEuFI8xHOP8YUZ8ebxsB
BTurE4Icl2yYBEgq5vhplL22YQFFq1sPshL3BQMVrx+zb+ZNMyToxIjieBvt1rCKIv5Xv33DDBLs
mxbcMREmXGTm+oOEIXAAP4VNckHaazIScG1BfDqeaDwsJgjmtgwscBKGhwYiWqvjAw991uFyxh0v
NJ2mmSDFTIm1ZhTs+VX7QqZFWLRfq9fuFlnR8DrG93S6seZtEEQ6uab/7Txdo4uQJEj3tBlGNd07
akz95AqdVkSaUAqrbDP8mLjYo96BuVKEWB68LNiMN+ZGQsrzz856YPdh7aQVO33clnpEc220dryZ
3u7Wj8LbOP5BcXaQ8ty83Zou7fEfIy/qLrAxhW7j80RDkLhnt0iWG4gNnCxEm9r4+3qxiPezoB8M
KC7KXgCLimS3yN3N1vQDY9ZEF9fOWDuYyPcQzsrcgc8JBemhb2THPYFBuQebwyT+kplMDBY0fenL
Apqs6gCyEzU0ouGHEnH4kWPU2Z2wl8id+R1zgq7BxO/6YLNQavGcfsAwEA4eYkJvgAlcrffhQcyi
VshLvez8adU3b/B4+t5C9UNVhEkytixGYdGZk/spLiwyErlSRIoVaQd9Q3m0mVlUc0U1Pqf59T8U
E89ja6CTJgW3V5qWE+8Mnu5cd0jTv9fst/EXW2s1PkjChCgvaKgwvZ+nO7GjDOtqcU300pZoZBKx
mImIHvj+dCihrM+CenRkyY2oGp7n41d46600wbj0brLSXNdgXF+PIiZzAkAEqw/zBwN6wBtGZzfM
lXuaal53+Gug7liErslv9mqM9DepPUgW8wqcsxA3IQ23SdRXVPIUUyPrdmg6nFY6fpD3MzsrB4hM
j5YpsLZM21j/vwupt7cHd3NjEMQdAKB69Ng9urz7tPKlCAoa/iNk8Oq11d5W7z20Sbanne1E9ns9
SMII8mo1Uy+3pynasUXXkoaVo7ZIE1mJUP8rl+1gYtloGRuFz5bc/1NZu755HRzRC6cfgupyLva4
lYjZiPYYHsBlFknbGfGdvTnmnOQC0V/ZhvYtGAbIFgzX+0f23jzaDo3SD6bMCs36xFtrO6WTlOvp
FVL7AVoG4dj/v3WlzrrftuV9rN9VieFzVkGeBHyX68hyJQEujUu6XlLARK9tdrxwwwelqosUspoE
FmmGwGXp7tsvWN7TXJAco6dXbJU/j9CTbiUg5g8pz3XmIfo3VNTY8kAizUB+2NTZrrlU65IDp6+F
IAE/C9frOBSpTjGovgK4oH15OGIoSju0xG45dXnJ6PoQG2LATiR2QNLbxIsucKz5csvmh06+PaiW
zHZPzLeAlG3cK7iWkGrNEewLnLvx9GXVCcVRDEnZcIK0aj65Vjnb1g9oX5nmOrHZ+d3qNZ5MGbuO
zfJNNQYgR+9BYnDuS6/7cqnmKHSdXso0xv7Slb5m3vZ7XJSgS5KK6apgORcj/jR2PLO3+sgJFn1g
DJkxJwSE9BTdznOskOsTEfl+6sxwPTypQ21exKA6buDFWSvdLWb8THKA3fBB3/V4Jfwdxsws35OC
w4RnzGv28wQGJ1shi8TllG5+2nPz7ZmUfHfb4BabeIo7k1UW3zFyOjAC999oMvJ4v25fXk1+B2r7
loiwftwpZmmD4Ep37YCUp7/JdMepwD2cXuaUkb8uemz26N6Op0BdUUggqYoE2coLCRZ3sFhaMbsB
CfN1d/Q8YRHH6SrpzPhzMjqkz5/hW8mfZWydHm+inKfCpfWNun2DEYtKUm7piSEyf/fJ4We9NRSn
sHYcBokD++SFuvsN/Turxd0FYNnKQ6aKY6A3PZZVgaKfbEKGlDz1Ngs/O7fS4Xp+qi4dHHsy4yrJ
SpqvMQTFRkIsJ/kFNYUlYKtMOhpMIk14+W83lLePTp8R8r3I4QfzT5YRaVScnO51O/BdGLYJ7Cs/
sHvArzxxU2KOrx5dTQ4yEwytNyob4oLJAvR4VjD3LU3GYksKIoJHM5ZgaRadBMaTeE7mwyFtOiH+
GNHxs/A/58NhSaGPPs+pENFwYLL+l0XvE3UGs/iwKRXvzMVMGG/SDd4HY3BWmkREj0Fzm7Ow/X+V
XH9uUbH2EpBwptsDh5Nfljq72tkE5biWRdnrU/DNCzczWyLcN+t+/yDaqdV1X59mCaA3T62SJY06
4TIyKAFreXbVqQScXL2Z4ZU9/tdFxzoYXHvvi+3lfnyYkKIbPGemGq36s/cPByFDrmwRT7FUDbRi
7AjCrUZ7eGIlzYbgp/Oxlj9aXBnbxAjj0uXnyyfQXMy3DqffL+Y/J10fgUX8he5I904GajBeMT6Q
OT/7thOBV5h4p8HIzLgTflk4cSNnGBuSS/9tRPkHtwmw3OE5agGuVe/o4vEQtnTH062W5Ecc6z75
bgFeJ14OPVFpHKIqZ0Mvq5TiCGo9QCHcMiuqn849U8eJ0MSu3QfjH3D1u9zjsJVajE/St6wrKYgi
ramjqZBB34WoAPDqbHIl76Q3pQLm2hrrH9vFWQi1BC/I6zfQf9Pgkj1/NmpP6n6x7yz6YYlKSsZv
rkg2DUGdwZF7OF4MjOryRHAlpQdjipFo8PAP2wAx/dYgWjPmwC+SnOtY40rKmlf6+HHv1Zf94Ij3
CLCTvO7/IN5lyCwjCLyP8ujgsQ/PhFiVnAnLNOXBCBn1m0OCUvVpHRnsmFDZw/hUmUbGk2dNxh+8
Jmk6Psmxw/71moxqghfmdNG2UjSZkyJwkOxSn0levusf1Rj2wv5I1qT2ya6Dh9JWtJP2r6c4OBu7
OB5yJlIxDc7p92+HcYpmX4dpFpe36geVgjHeY4FSQLK7qd3gBH2eH67EOU+HqdTHapZXsNnXK3V/
sWBpot+Mztzc8VdGWktu4+tO3P+4/LTdh6r+BJxOvZ1Tu0msjIKMQMQkq7x6N+ADxdzU5WtztY2p
ciwXhxADd1xepxJGYi/ZLHM8lKwckTKB+R1nauCdTAkuWaZ6YTMNMDUQ9Ooa0CVUy4nUmG5dqpIw
tBZj8BLBlUE9G7J7Mtxt7W/0lWp4eNqt8FxQBTBwsDM/cHGXXENrmzBLUfdnUemaw5hFqcIYZ3yz
m2evLtURCRRtOML6BOYQidZ1Q+1JlU2dVVOGVK0XS0PrvQYLpUSvC8r8uP/CL32Y2rHKItc7cqde
NW4d4FprSW6jbZ9G+Z/jmE6DB1wPaDieUfFTtYt2lPalfhPyoSpMZV7T4l9nAfCI3IptmP4GHl8k
HAXtBQEnS9lv79NkGE9KPbL+WNnSQwXkaLVr8gzuBHnCIq5xeF3ZdjTN2kYk8jjjLOjRcsdjkpDt
9U7M7VkeF7H3gLdrGdA8e3xf7MQv4EIuPVnfpkmWNM34LkPH7EUE7U9jnfGw+UQ56MiOI5nMWnhq
e2wIpgvWKbrrxVJn0+PLyf7FPo3yt4Zf4Bz0dH37t3V0VrU93PG49hjGVAEvvtB1E2hDyhui/50x
Hm9KqPIJfTaJcZm7m2VilTt9QUf1mr1X2cwWa6Fzj4IOZAD/Sy7NLuwt90aCuMzv+ucNHs7ch0tT
Ibc3t19KigPr/TCaBgRknjevCm4/8HyiiMosN7RnzHJyuvIwh8AMWsLoOInqiOgffBH0UQShO6zp
t/03ARAsf0Yl4nfIkCpACZlJ4Oz87LQFRCTZUEdlHqE/jEx2pioscChKLxkhYZUw3lB4WXdrcIS4
n1Qb6axw0tfkA+ilUyR4Z5aWWe0aE3rujnOsndyVapi1qTwFacxN8mJsKRQsjpFWh061dlRxo1Pi
ek+VTE7oIc8++2VYhysGihvTKjKXqX1puZvgNfwVFCJV0TBzNp94dPm22jnikkiFjmrF+bWZxuAW
g1zmiTdXFFFbnveFCfRDn2wdcronPJbXh433Sg9w1Ld4b5sgu/KZJGxuniR9Ce6BeCO44xMP1+zn
w6BP4GP0F9BwRaMe54P/cx1YsWA0T+T1DfSHawYXIn5cJ9nJNZRXGaGD4vSDO35oKzFJO/74mDmZ
hIScOXvl8KOzSn/Dn5Phmc2LhDcWLmRdKNmNH+oBV1fUo0s261RA/ZgyrR/QFWmMmwyEVirSO1xU
hFLqKEC3MuP2Fmh2+PvWM71A9g10s2l/KYF1Yus1mRrPgV/FepZm6jcv18iBY++L48JNWbP7DfOo
nkVDCAXdXhbRslGZGbV66CUng8UpAPhL9SDM1mY7/tcJLhPlHZYMeboefsy9+bZzJRLQLPTOLZ15
FM2cXP+T+xhq90EM9WXc1Zdtjss1JD9HyHHmEOW1MRX4Y0rYSWaCjjBo7L0+9hdQIVymIOfnhTy1
TniTcrxJe1cxWIevvGqrIQAAnoKoMV0y/T18kEEYxhIIP4rLlMCoCFY8UKmNmS19AqxSOrAoLQiX
jSMJ5JxJMmLmoM1TqzfIOGg0yeSb7Of9sdxCvZQi3tGbfrDtzsx2AKfnV2AckPxNzIFYZBkqAgai
CMrxva2h9kPpfyD1k0RZ3L9I3M4/L633SZm7sa/do/44BrITYX75tJZfa83udfmtyMXWm1Xh8vUf
bEeoVYMM3MWLdGzBIFPzbNHz6myYkOqwl4+OFbX4JYwHbxBwXe9pkZMNOtuCzSum87e5aSOM/2Fy
ruwDmLqQBhmwcMen0jrIu4BYXK/k1aARo6qhlaoWoGx+5UTYIfhRLKt+Kn/yTHYUxRsDC9ySt5VM
uI4vhAuU/8E5RfjIeBmP3rbzAFDeoeFITCm6gswmQsnUpOc84EhfhN8UYI/Dff8V7zl/X1Ch5TMq
d2Acpgg0yp3LunUSUEFKMc/eRG/2BC7+oAzXATrsG3yT++SAwHPSiJWG9b0AMuVUR79VoMBgZoP3
R1jDDb2iCiZU7jdzJ1joryVFbIMJinGdahh+8OsAcN9dPX6Bdjvi8p44gGpuL5ICaZy35Af/0rqt
KOH1zXfJmAvyHy2DqxpxIugllrV+gilM88E31OhvZtVSX+GA9mbhnFx+InsDQCZhyk8ZYUs+6452
U5Dmp1DivuO/J1p/4DmGrAu25JSHscg+yjNGKCufTi0bZGrXswNZthLsxKTv6D7oHxjmr1DkvLhl
QDn5n8zW3R69JyDR1w/05eeGS+A4EFRIdFZV9u/AN2PQF8eq/emFnTwka04s8m/6FLEDV3R85yRr
BnDIdSStOI+3Icazwscqr0dKIoBpnfYVOeQrs9fSwRvnHL9RpxNS/EG8NENGWUQ5m6lPpceDpot4
2/s+J9FAp3LQJEPMA+/0OUrR4pMwksEctfb2cpOCxzIG7PVvbItFn4ghONQ7lfflDzOKx1e2TLRI
gIQr1QJEUJ/y/OfG8o+AUjWvmnTgLZLG72VEDduIBWaUPSj0UVVEZa7+p/+bNSDfkiXPv0obMlsr
xt77QeDhreQy+QoN5d9/ZyYd+Hskk6j8fC39+qvTTJx7wnykfquX3MU25Rg1AoMtM+FR7TwZBcXL
oBP+YN30sFnAFmMMkLdxmzxJAIiVeWGdcWF5w4QnQU/kxoHxB+Qs1vFOo436+yV0JsCZy74/ychY
Yg9LUT0/29VJrw6pu/25XBqFBeelI3wVW+kddq1TkpEUwhLMMaoIW/J8uhYsgMzU/FIi2RgrOmZ5
ghiZ+sWP9JG1gXtznBRa7AGZZW3JCZgEIZg+mR2ktZY2KZLTOG7yTz9jByyi279/YL4MQeuBOobH
ERPSFMHLV7lVbjyDFWcYbMr5hdgtOVoCeIy0M7sCLEsyKqcD47neSsx7aUP9k/7tkr7KC3SgRbqd
y2B6lIFFn14w6f07oQa6QoLPWJogagBCEdKEFm23Yhmdtd+v6sPWNmNYWnt1FGrU/QYARf0GLDmN
Z4obK0h4mqGf6M0g3R/sdaK0HsXqxoypUJurqhYXgnAWcAwHI4Dr0LTJ9ptNBmJlpx0tKRPFUaNe
zyFrrl2RGpTwgbrIp8Zrg9w26udtpAl0w9vp0M+AjPGwtFLLmOm9BJRkqQPEyb+ukfhaK1+F1GIh
7ONvDbwXiP1XfgBAzTeyY775cZeVCKYtdseIZDSHvXeSo2sJdA1knzNTmRqCiPErj2bqzYRGXsLk
MpHTOO/pwCDOpx7p1VJ9DZEFnIWa+Fhu86YY3DJYCwFMWabM2+JJXKZCAGicTokJcoVL0Eq+Ij8y
S93B133HUrTztAy4yLDZgSxGGIVR/nh6b9Dt+RTxwibjkTfG364QgN1KmVaKEyuQ1vxv90uiF2Kx
woiiSNq9avC8sX+N1LYWlw2qOkLMMuDaYQmXIQY23VeUPVhPzSJMfF7QQgBT0kuIHvb7bcOX0xF+
u4iP2NeuxawWbXntdGfWOhX5tVvqWptRwh72rJNJ8CEf2u/hcYMd/Y40LMj9UkNIqrdgOA5x8Elm
+ieUarIRApvlLomKfIU7MJfNFjS/P3+bJoC2xNN8KYNjrP08a9u2CxVQg8Vl3/d459zkIQqG3UWd
V2zZXal4PoVZZOg477t1FfhlwptTlk9oGnr6S9xVrPLfclnJeE1lTejE4iyOHFtaeMGA/kPXz4+3
5Zj048M7aCmRZSv9VvHT9zuAYOxoguOWvbHZ08+TT7z0j/6NBVRYSrBbdV6ZafqQK1CnzgDStGYY
Hwd/ONA0PUKfH/j3an5kjzBB+NNJQZDLSThNIvpter02Wp0qWeGxncV7Z1nR1bJuUBVVUsDOJcpu
tRdSwj0+7QAGa9PR+fGbac65DeiX6OYhHuOYx/SiGm1DRSQJLvNq72Mc1ecbNxzDslwuDUM0ymbG
GCg7WWskCfOLOfxPWywQmZhdjkD3/McPhAtVks9TpLP4kNpNbseNX3YRksWwDlg29Irs4TL+00BI
XkXYlQt8JXsA3jxMQnvicOlwuAtBA7Jw0s/hnQXz/dPN/CXfu1Ya1Vj9yl9yCu78fIufKoAvj3hW
SR+WNl9fo18p7lsT/XPWf9J0a/y1nEB2iN7ofFGuRUwmvNGzlQT3URx7TJl1DxEdot4m8+azHe3L
Mw1NPslfGlbNV7r1tM859s63/U7YxYfmpXQFhbC4DE5wSVsCruGgxsj2DTZwub1aiGjb/XBxLu8y
PMLuAYJuyEMdr1VTi+9A4MgPwIqp18/cNrBiS0Hy3999C5cuyChSBxXjiwViyBw76H5dC6E5v+Hn
eiO8cHqdEQPZMnFfJMqF3m3SLTYRKBSNGj0yEr90EITk9R8gLRNxgSE2J53X+CY2q0I2rOB7DUj9
kImDMm6kBDFELuVBHkvsv2vA/ETNqqXWdelYq2oP32L3AC955tBfIHRQdpYAyUJ1fYNCaqAjx2lO
Xy2whyNaXahiAMrJ8nZT6VDX6fdI1XnnFfcLhrpZXtwEsQTYOGGLXSIsV73/NCuraP6lhZY9zRx0
GY+o0TvCDjhKE1yNbohsDzQ0gqNw0U5kjittHv1WLn8y2tHJnUVycbC7aE8qVSpiHuP2S7Ugud3w
/aP0//0H4FVoiQ7julI0GC6Tvn8y/6QH+q7HAVVn5bjB+8M4K1U6ydeEF23Si2UVDtlU6Y8BWQpH
zlP0qB+RlRUS6MheHj6vo9NSxsRmA7ZsvPKAmISuQc9HOTYTe5ckBqyGSloHA7/OQCPGvuRt6/Jk
brVSRBnG7S4NeEZAZbQj77hooIEDledGKOimzW2+FKOnYoQ+4zJt3Z4Mza9UIq3It8RRBR6IkYyo
ut3TZQknSYo8e2q0fWojAyj5zknY+6NYO3LXLyy1K3fs9S/eySxVocWKKkF86kVcukGoZS4M927D
dtcPGwbO4aETTY97MRiEdpsIlJBtiK/BsjoUjTxnOnjGJmQFHJU0S4IIpTEJxnNEV07dppzA7Frd
Z/NNpSI4aPOP9Tzsie5C6O9ykNlHDNjw2eOB/P1h1ly/YuVZxe/8CutDnZ8NTQNwQ2ddfF8nhpzZ
PQ/oCWui9jA/GZXKxePTzAZJ1MnrPu9eoN2beEmFs9T0d/XOB4XAgpc4sDc/T6Cmzs0ndOSKMFet
FxLkYkQtcwASxsY6LCmdBApjEk/QNZwNOYDd0rbvOnP8rRjSVB/6IQNbuKpCUwqR8GA2yBVBEFLd
7btl+JpflobzcryLzcXAa3FxYrCLEyV6MefXVY9XwU/6oTJRj/RQO0jMbMr1JS5BJBMpyOLVZJIW
6hI6VYamtB9sVBvyFHtAGck1byfb+rHlszwrAUJzXSunpnNe22S4NSHFUdBnyp+1mh/uDlpy3Kyt
CBFUgtkuz3/inMKmLdkmZcwcLrXuLAcpps3nOwItD7mLl4kexS/8pjE5ayX6ATKItaqFx0bUYq2X
z/JMwfAsIKE6R2Q9prCmUvEEyemaQtWk6P+iOlU3Zi9Ib67UZkYo/UO0158eIV3kX9QZwkYhRv5h
X/zyO5DvsQXA62D6o2OMmRP5r8tEnTU15GE3jXqg2Jd8tABOEVANRCU2wxUTebos7+4WFPnB7Igd
K5N3LUUbu8pYsBqU8++/r+FG+P2a6kd5+nbx7lQmnr+Mp+HHPrxkQkQjsE7/UBZr3dPoK2eEHjYK
FbwW7zG+srK61WxClyBZVc2DLDlpnV62tqH6Grc5xKSiE8sCbA1f6ZfY61oXzETyxGh0CTv5368O
FmKJQ8ffRSK50WrcQPB8v1+bYoqjpdi1TNQinhtUIeF7Vuep8htC2eFcP1s070FEFWmqojgqfD2m
sZskd/gOqR2QvgJIrSb6zw2gGG1UMqTMapPwm/iGxNPohiC6q5K+1R79/kvNIuFdgco7q78SmgCO
qv/T+kkrZzELQgmQNNHEUZgcaPqaCb0/niPW+yfk11VkEgfkWDfP05rCv+JbOjKlyyAO7GSR/+9l
RZrVf28MC2RxGYuBZxJwazBQMeMzcUi6WIyj/e/ybbsnqc4U08XxGuvAovl+sFaCkgXl//HcLz/V
K8tHF8j73oJbTxUWgazRg7VYG2bkFpDAmnP8b3zU5un1VGg7J2nAf94BAAay+8ilWMHXG0T0FgK5
DPykqYJO+9dz6zqr7svHHxWRm8ppAJ15L9rSMjNl5dh8TNINBTky2ucaLmqtlH43G3qX4edepj/t
qTf1h4YetCB+f18QXInGAKjrRokd7zr8QEMCSLIssSquyTwFREmES8Ecf42SnsNi9RfTu6xuu8Wq
3rCARGxZoR7rEI0ezC0h0YuYRjnFfLQ0Vg1GVC+H76p68zKHWkp7zyzb+SW+Pj1lxouvTatA615W
lustdXk28GOkvDJ4hpQ4MpLiqUsgdwRm26d7lYcjpCxHQypHgK6/3uUzLWBRbK2eSmt5qrtQk6IY
FHtLuNmVJ6uAOkm5xa21VwyICakg7lp+rbwpt0BeqAdTAe0EXYOEWo50r/B0vaCA/FSCvDBHKamN
pyEm/vpKfCcyMwutCoVypsTb5BH0nSI5Q8yMMaULKjtpjV7ra5OzbxTuxthDSgKfGwyicgrDqESE
/bbZZ1FNNl8pTXnw/TEifCruMIMDX/J6AJDJUwAIx5ocSDgyt2CqE7lOlyvXUsoa+P09IdAz4Pce
1R4ruvuNb1FxYWlcd8w4s3jnhcnroEqfOXcWL+He2y3W+SAVeWPq45qo5qpnW1bHFMyOSMoP++/I
fGkWwQ81qpZTzMtdo4C7jS3UvjXCsYZkexl+xCGYZBynwBsrL4k37nfeDybG84670unVWVIcQ6Rv
JdPTFewz1JAuS1zsdxlrii1DLdgPmn2hCJs60DVb+FqphAKhcGSVxDInmL2CwokPhiaOvdYTjXuH
D+sVUvQmTSbgtTOD54s2mRRs2Kr8hyv27EWm7SHvarZJ7foLAkiCGcATZUzB/nJ9mNbr+ArfRi6x
rCOtvVj7QgRl4cW2ZWSiLJ27cyvQfNmIgAkXoXeGX1E4GprOlxN/WrLnWxeBA2WZ2m8sNEL/OcPp
Z+d/DyJrLuF1RNfDZrE4loMa3ZjsLnwPTZzSiOtg23s9ZKhj/T4dj0rOJ0xiHpOAqmKNMERg22pX
yhfNMNiZeLkLuy7TGvPElAtbrb0Ha8+Z0j63/K27qoXD4xZtgW6SKusn1NBvEPDbVa9c8pgU20Q+
LVATXVud4Ypf2oh6mzDQFyhw3RSWfVhx+MbQLleh32nr3ZU3Tc4mWCKLZEcF4YnEBR2zZuNs16Sx
ra6vOGeo2sSwcs2jQwjCn0QJw2DwEGklJtRvJy7pplMyKAGpVTmBqVj02lHRZOoxdj5MUuDMDOWw
FzIKVZZZ00vXI67L+55b95Ygv5XqixxwOf7RqIHueg7EeKcpNe89NNA6tkBJ4rg7z6VIj8AGd/1W
y8HPrOL/ftB9TyMz0crkHpeNCLFXw2eRNoI6DbEitYzJCfaPROakvBBSjJmhFh938KtOW9PYNBtW
0a4Wut1cxqUGRAdPwUWJ6rpprx96L7Nn8aBX8y7ZXUwGvrck5gouq40996z+XxI0VBwP9tZGI9s6
HfsSxYOah3OIB8cd/bVIkaIv777A7lEgI640gqtruvW6lH/RP2jwzY8NhbFZDS5VlkBj4o/NkCPU
Icia/gXdxdQllopATeHIuvY/J/RkF5e63Ndib8WcmJGIpcTE3QyXrFnHzKrlrLODSozIwIHl+wR5
OvKiVnGOVX/kS2KPggvql+ylfCahCUYAhbfbLMQT4wjEUnB5NaL4t42RI+SjqDLOvrDI0M1gj/oR
d+ahKnQ5E3p9eSK3JKW+5Bys1zbaK6PTQ84CVnn5nqib7hAv+q0MqW58LnQnnrYI/80mNMN8+IO0
NC5hTIiHXzmrSRJtNBtuKjMkJ8EDjmQgGXgWjFgiIxvCAmgBk32iG/OnsmNSALW+9LYD2ZMvd78Z
QiSy5fHQ+P/acdfZceEbQmMR5TapLvwlpjsD81Wlf4nwZK4fYANRWupzMnk8OnT7gV3MnWQzmO0D
4vTIqqJGOX4r/vRwaPVhDoQXl9RbRqjpOgJ0THugzEnNtiKdKdr4JTaJ3e2nRme8VNuv9CfanJ72
9OlG3M7gr3IvQzIgcb9fFJxH2REXSmBwX1rL3vcdoOJJOGdF0o+4FU0vwl7Qx8sWqEqyFw/RtVd6
GHNc3v6CN5vqRNCY4Nasg1Vlc6ETR5g+cdjnYqZ6vdBObEH+J2FbcYi4FjXvsuHSpaotcOkzcq+8
7ljEZ6LTPCfzSaFQT67Cu/4GLQiraOtqBi10oYbImEijLvo+AXZ1+M32QiUcvKCNxKWqSXGS7M+c
GIjGeNJfLUC4wyru4x9csRJvmEkkWyClNkcoMY5TZRRtX5klc6wy8i4Ib2gcy6gFpN44E+w0ZPJ2
b2xaugclC5ezDIE9XyvBMn35jsYswwC9o4f9P+BLdlCfBOOLFS37/Z1WhxgOdUkkBzXbHXiz3RVZ
hHOZl8aR2qUJBHxSBGv966HU49kXjY2xAcjh4hRLiaSzolY9k2Fic5BW18/nHI6wx/popc8099Bj
/3+/3mU6v1C1piM2g9eG26sdedukkI+ezHdoCPmxGNOi1qIuxXK54Pd/AaUxCi3uIkWBQEt/vXRJ
g1EybDczPmRWSO+FmpVFIFmJHmBVcdBbb9Gio5zlm1je/gvNZfDjYLocXjxdATi6PzybO7+hPYO4
gV1itZY9mLZNFvvyWc0rxkzxIV7LCyCIj79xoIKxJi8bTjp57jyWlVFdMGDH7wF/M28plFOYP4mX
ZQMGQF7bbqI8R8LScY0BLPIUQeZ8V8QdHu7Zg3vtVptMxI+UF/xHjfbT0VoQ47Ao2vHMEo8BGr2C
HAoFC+COatCFa4nOEjzo4WNqMzGOIWA2e9i0MzutiFlRrTEFyLj5i38jcFdavr+D1/WUUBBZ5fLt
VC/UtU+giScgYxUktgE6Gzt4iW/3Cv/SQixIJXFwC7drN8a1eeg46KrzV2kXYZlR2cFaCu16gYrb
3PtQz8ViBAGcRXD+KbJ2Bi2pj8I0e9Bvu7LD0qYmtTzcQvXhlsTcAeEuewwHElQv7YyMTBzeV3L3
HnD1BODwFqZWG/gpQ+HxXpHTySCF/WNtE/eBPl1cbzJc54OJH/kevkaPJDW+ChMgCRJ1vsSCTG5v
a72Irpg0snvdYK2nT0sFfwJP5zwDIN+rbY79VqIzFI2n4uv8twYq7xqOaxxblA8WojobAxK0Q0Zg
6lxHSHf/+kZ7qk3gLrm7faYFiTGET8kpMDizilLGVIA9SMV+t9PZMNGizX8/Uksnee9J+IdLx+E6
b+4YaxOduYR32NfFSPteM1PXzIrYZws4/WrC4KqqqHT1WVzBIhyfpqJpzLoIZd+XPUqZMbtLxcc3
hP0GT5D5someH61Pfbm7peGD909gYMmv6rQ25SZ86YinacpiizVgJ5LnLImlWIRIkLqwrrTx+ueJ
7XMrwzc60r4XW9caXtXI7shHv9jUrjqHwY86Cw2+RJq6Kitz9t1uNxlk6g2rgY6lVG/vKbaYFSMA
ZXgUD4PScrbGtDCOU26uCcOw0Z01yb0OMio929Z3/5aMMnWFzSkLXowd823xUEuyFOXdJplu/J4V
K3GjwbvnsJS5VhIvOBSXCv2AIe43gkmQFE7ENENbx9pnHQbWjDquslne1Ut0RXWpGcxh2cPBbGZq
zheeAzQia7lXJKUhmzDa/pZQvjS4dRIUrpps/1V5Gap18/umNFL4ryVPkB2PvAWvjR+h5azrTpzR
48AT4M0LDBaEPoLqq9qi83qjbgao+3UKWBB6uI7+0Dg48CLVO0CoChjaELzf/8S1HA0DLcsxXjnO
xV43qmc/4j5iFyXDv4bxUXy+uLWpFLYvBV4OUeoJnbJ844vkrvVi+EDiI2zzxeGbzYOlONl1DpWW
oRXYl0+DpUyj4t+o97WgBXh7AmE/kRscQfIeNq0WvQ5ujBV8YydSUQCu9GQ6NLzkabaO5HJqWcKz
Ftk14D3rw7MO0lAodIwZg8/DfaZgCeMWeCNAzBOXxosQgCrnV3Om0DiHrJfWfrNQ+efLY4d+qGKp
8NOHl1cT9inCyDNqBDNuAOMVdrlgwkrXii2+fpVIBJO8G92ltA6y6GxgRWbkpVjLkkZD8hDbXLNd
eH1CQL0Oxx9W0fpG+3SohshjGL49Lhyde0jcm3IK9eLc1HnOjbEj6AB6ZeP7j09JCVahCwy7jt3W
T1sDhcQPRznrkzA/tkTBEJmQBV+6ww6/KhwHweimSh8SFaWZ4p3JE1mw8ym3YD7y4r+VO2VKrzNj
KmoBxAGcxuaKiTc3qpa8Hi5ol6ACEGyc1UPSdb/rTL/tDpzTE7iunNH2bx34zjjPrKC9KMQ900ON
RB+Up1ZXfqD78QOju/LtmT0VvqyR5Ze6yrrJaegtC0MmlFoPpnZZOD6X0jjkbHWon9sxXAHuxrDo
6ymuoCyRuhtozKO6N4i49/MQ7xMrI9XU2n+IVcqCNDYLnJJq7LoRjYlyipsvVGKQKZ+IKlVXJG7v
gks98abzjmBvrwo5X+wD1n3LyrY/TrSJgZDAdWm+XrZjmi9k8/LBqxj2HBa0hJS5YHLjVw7rd57v
LvSXhEMIkTpM0RNnjO5kZ5YtEBQAyl3DYK2gROVuVES9YUcxn1b2nA+ZC33sSrp6eCTvJ84rzlce
t7BI2PubtCRtq/YTbbAocCDHJB0Q41SGt58bi2hOKnLkb7ioZWhsPs2/eWcsoU7y7IqKQCDNMGrp
73IntW85su9PmQG6aG8ZZYhWjSAP5+M0nVP7gPWEzFMD/U3RdQ3SDvAGjlaaf4FzP9sA1oqsRLns
qCofLOE9r+dIMNh5pNLDSqdaVxUW13/4tFWR36APC7WgOvgyJWdIuYoPUXBbCmdpUpQpmdwOFsJT
A9/vhsgCkXRDRVcWGuHrNrtVbH4D65D4pbetIqRaE30IcCl+ld1MPSMuIc+7iYlhtDF+U9PNcE4I
b5zDF/OcfMIPGbWl2khjfg5vqYhfV++inLpH8hYHbE/vu7pUZlWTKHeI6Nhp3zNXDM9G6XMCPwzj
FhQ7qRdxFft6KkQ8B243Y9F0pOD+3TdW2fy6cfZxw+9JPYehWLZMObZyo7DbI3VInd+FA5GUQ8de
/aCTONTpQNRB5Tfjt+C+DICRFmq5xSSrdBZtQjZn34bsRGbfIBjRhMbSmV2BA8Sa3vslT5XOgpnt
WEsMvEj3C/ZoMkX9S5cXAywcKaMXH8/7tk30SoDNCSgUfFDUoJRxbRr5IZ1dY5Ddh/7hPurcV0Q7
cWmLzzwcSeKF7M85107BOYkU7luUwZGbLpaCB1Lmds2f1dvNrN2K1V7Zez3Anrp5ddkSC+VFRs03
p5owWZNkOMMVLFFv/jCP5dMx3BK2seWB7j24JswFkFPvpg8g3AtmZ5inrHUm/g/G2uGBc+uzcWTK
i485o2cE3LDqc6RrI2RbK7sd9e+uE00NbBAkIraqJJx8hpMmHePk5l50dR7RsbWYe/545dedWDde
eWhl0/VupR3r23/zJhBlw/sTsKnF4rMfYbzg/K4Llnw3Vtz+8hhPJqkHg70AvaYCaB3+8+j5cKYL
JGbW5+s1jplOFPuLSvE4WOq9nX2M33HLDw6M/wmAFZRqUE46Ff3yPdF5Xg7litX7htbiG96cBOK8
rryZ2o8I1hKf2XOmYaNW82CEuSElw/UnDE0uK3VOkjI8pmDclORmc353Bhw2laRdhnBjSxBYbnH4
wh8XW4GwFL6AZKgTTzylpfVhbiRyMIBp6aYo5Cn9JzGC75CnYxEaoFTm4HZvNNp1HhPTnYpXVw5f
wXLcwQqFBT+ciYb9i8Au0rq35FVvVbhhpTk3OzuAnAHqDqpEPdrpN/MfCDXHijg8uaO5A+2o8VAQ
jESGg9nzIanRbib6Ur5zDtnR/4VMOGZRfXcgwbpr99EGjmGO47d80f85Z2wpfOeW2avDFLe8Hxx4
UXkzA74bpmYh1+FmtoUWdVfcz9GpDG+JCrqy251yKwRYHRcdsoGEkO7vKkfzut+uII+1yzWQT8N+
9iO1B8zMSKu3gIHEMzHal41cwgN/PJHPc/rKMt6J0Tcbz9ysHO3GWLZXaegFAsoNJUTVcFq8QmrD
ZxYO78i0Y+bCOyhWDXzFN6MjHOwCliJ+AbKJDE2ZUkcAnvepdUBexaYlGpfJwbG/cn+GvjZIH2L7
W3IApZpwHsUZqjQzocg32vmX+uHpfHa3WAan7cOHdwH8oYqFhbfD41P4sU1qTRbWEUficSoNL4C7
E8NAPx+07xJN+yPBrOdXx0AxNO2EBHTfVdUh/qJb+3YCOzsiKaS31kVi0qJkHeQQ/tLvJCNK463g
FZZ1UA0/cIzBHm9n8KxXaX+Z1i1ugbqIpY3Q/AD1AQdhTx9qBdG+dhawnKafw/ds6nrMbuk7wSYy
84jOQp/Ue/1quE/kSl5p1JP1+q1yF1ejH7v2yNN0tVdmewN6N+vevbF1B7OtlS7NIAC4TY7mvxn0
di3wb48ss3yrjirBjxgALdweWW0tP0STLA+53pE1QDsfssOXGdNXwX/Witx0jTLRXRTewPBc1ceZ
33JMkbfH0/8+mSSutPR+rR+ROaJvVFTQ9ruLly+RNbUgThu8KjZ4utoZa5COS09zcvKKY072zook
dysvvB93GMLgHErwEMIri6jFSFb0vc07GRHMPYfyov3tOTZ1+vTrTMFwO1I+aGzC77IZYewhkQWS
I5P9njfVEfLswDLo715qwoC43WRyweHw3p/k4rOha5TnkoAjAiaaWT30GBvHxwvIv66O9ipy31O2
lSzsZYA//18mUOlJRflg9+26CXZQQp/FNez5xvqLyhtK4evzIsO5gPRlG6fLh3Ka+LFaF568qgXf
PLnNqnnpopRAHrpSGEQpI/kVxhak/TtJVplUS7NpTYm8z0L5mJb3FluOU6bVe9O5Ux0t06VKTFfV
4VtaK4bOcfcrHWOXZipGAZg4g8I+6AK8Wrr0WU38TmOVXUAis1NYOxY1Zd8whmsNf+6UjTFVfinx
al4ynsoSlR8z1XEEaEKFVXuAbQydhCeCGjhuyuCLGrPmQrtOI9oTSmpQAtLd/EGzhyLtenmRKG93
KgG2Q8t0VYJ4KWdPZRPjdr2lGK+1JrZEs0KrAQUceRvP0AMtdMiReimXdJWBAy8p2Ze3hHjCWFdR
CrD6aW5sQIDMuKe4eYW8BGMoSGNfTA8iTY4pYcV8mVILmpeyR5c29XAWO4IyJZpRAz8VsqKZv+vZ
G86DJ0iZ2hm8vFDC5hCWsLUmYt3BCazUiXDXyLGy7qvTYRvjyc3h+mzOXCm/vfQs+wDF0Ggfz9OT
O7RvKHBfn4Ienl299EKtq5CIYtSzVHMQxv7AjqHTpF/IX6oERDy6BeBAyKtUVp3jSb7OjP+T/EfT
vEhP3qqhBFVQWQbjnsqwVqKktpS8T+XIcmRbB5KXD9aW1RD9BIaEaKXMzm6X1f4NPt6cs5Z2cJHp
Gh3FJHfp0X/AwV17fRj9TzCjwttn0WVtumQYDBT8OYqcg8qsND6my1nDG8sd0CkKAzEahNU5xPwV
YBcjATNamNvPGFPIG3AMMbAEb2ryRQl402mIetGCH9HpxuBtbOu8i0nQ1eNlXOLtY20YZtvSqzvX
h3nkWFHEhifr1RReY4wPn5umhSfdnk6BE1QDobkxNOB37lphRNER2YymV8z3WnQSDWURaY9j9UKH
OreGYHzcLwKbN/3dBXlNle7w9x69osU2Mc6r8xTfDpyJEEyvbtIZfQBNq6a/h2u1FKGi7SVBgtyD
Fc0EASZgGrz/2CVpIEZBk2zHugw8cV6YClC89zC3DNPyKuuRmsJdebfvRNjUEFmbbqWw+g+pLAa2
dgq4kI+bmbMARO+kKhJL34/PpMc7mYXqJs8zm1tWh6aFM9JIErV8CN6oLvvXpceed5XdusiFKZbL
MGb/DvBz5q0eaZQ6Frswve1EMtfYdi1DrVwwKptzOuMF6o3NClHnmAq/Qsx6eTRDhyBt+WahxPSV
fFD+znOZSn6UzrTGvTQsJ7DjGzf5/ClhngAawSzIrM4xLaGnrRNG64A3pQCu62s1NKHP45SGFBi4
mGzpJhvhVhe7GHfYPx+ivkdCUGLcWmjlwaGzHc6UGSoIvP2aLHMlsXXjBlyTT02M1TQcO9cr7I4/
Mv00YBFvmkd15WHtHGxNtxoR8LHYIxB1/JObgK7EE7SjXv2hBVFMdnaGq6TARjMOgidV7P9xFGcr
a38erwnSN1qGGDCpIw6ameiqXIYGRrS5vp3km4iv9eiPf11da9MquX2hFo0/EPviiy0Ks4TvAiHT
zjgImpP2PQjYRE2Hh88eJaOBBsiPJqj+hYH7PwZpurQo/dGZEFvd36jfcl0PeKyGfsUzEtwxohgM
0nUoPTU9nEYiBF46cHmZGJq9F4dlhAjtXh2/kjr7esTaRj15JipKQv6HE68cfmP94V00Uj6CxHVX
3fcRWQrlFx67KbbzOUYCFsAJvDMwK/x0Dzq783+XagxjB23P14sxIV2XtS2iuZpK4anayL2FFtBl
RYvPWpsfLWDM8s8D/LNToI9bVUWcG9BVKO7XPyHFDMu+Ewmi8mw1snSlj+3zQTxbQIFpVUOP20fO
sU+fqzPO47z18ewFNYo+QPyTHCA8AzJL+OVPXQuojkbuOEKUsCJtRmU6G1AX/UuJA1kEzRE/wO7L
9uOENbyaj9ge/nvzjzDozmSi2w/yJjdKon76tpXMwf/bUDMUk5/VLnsv9ndSrA20bJy0SdUG6Pr6
+0yDXaDkF1jaDHrJbm/Wv4gsNa2AF+o7JdfAUGWnyOP1tBZyFw1ft8nvGP1g/JQzJjg4Y8/zGv+X
tsmhO1pSg54D+6J7aYzLgY9JaGzUrNKAiqAmdtDDTQFha52IQJxzKbd0yAIoYX5huON7tbjTTHbP
gHZ4HSb+wAYOi9f5xRyIf7MihW+wNs0LcFgIjeDQ1ELV6484Fui0+D/T6F6FCr8Zy5QNGkfBi9F8
Gj2Xw4F42P1K03X1dbTnTF3Nt8d2AN02PPUl6yGwft5uPA7k5Mw+GTALvpiBr8AOdxauZn/RSU+7
a8r9QFCgSm7pQTsVZ5dirpp3UloB/cCF0Gsd+nAEq9FxpjmAmec6c14Wa76nsRMGIw70Qzxd7bqY
0Z+gkIF6/b1Am2cGuLQPn0xlVkHDmzi2rMEzoYOWVWU/0GkIXiD16WsLXnBzZ3jknC6rrlrwrk0j
FpctAFMC1pDbnEpz1q5HpQzkt4s7Jl0I9Wl15z5te7sIrQc2EWliNoGvc2da/J2iOkNe948ElLdL
Mok5yP+3MvLHPnsjaa8sRDMGcvG2Kf3RIH+LpbaeLPsEoUUVpqZuTUTFB092frz5/S6ZaXN54oAp
Jw6GzGULMYpKf1ABmwpV4/ydR9+d2zeGQUqIXG6S1A+2fmmBIsOEGySZjIqSNDo1cKeRrhxZ0aX6
+yihXxyUQF+La7cu81e6/xqvNceT3UTxKIjH84APLTDEAqfxsF3xZcqrh5EZQoWFB7RTV6oXryxj
2kIAiMgVnfCA2DJHso06QSpVl3p5vkhtOTtWfVwqfj4Kxg2LeqD4ru7AD7TQmaOscHBjyfpneKLY
pHFmEZAO3bNBND2phX9++IUREL5zOLWWLcov+9RX8O5jjw6Mz62Cx/EHJlzVSZEleuBwRy6cbMoG
B9bMw5zVh6kVvKzSHcn5HJGiztygNdemv0qMkFAveOcMgk7688fLY+SlbBDIW1V5a++IqSmFoiZj
1qm6fmXuRuVQmKVv8NAOPuz1l25p1oAMDhX0JDmRCMAyAE63Ti6eOcyOgGi5hQhpkB0Qz2XozRfM
8O1010X7QCPTmeoIOWlYKydpGWPhAPTLUt7DVdPziWy6lwgjUDXaAd/LND28WHswdSohpK2G4Sqn
kmJXYTcsCjRjmusrUQdx9oKPzS4hn2sRZOC6foz5z2ntX1N8wJfqX2d/8bNxdENp9VFDc8o3DMin
DgtrkNBD1uEUOr+8TazL2L2PGAI07R0lne3Iwl3BjbW40cSRkib7u29kltkQreGKj1tESYAdgQIu
/S5BI08HLKrps/mdL4jhVbo5TPUeQFNOd3sbM0mz3CcIjCS+/7ytoY/x6r6Gl4aoTL5TWcSn3xy6
H8VslvnN/UhZtsc2zqcqXIXIaOXHbAsldWA37ClS/PJ+phReg6OiLSJLLQiu5VtPEl/CEluuzxJT
ixuIalVpP1rDlYThk9xb4pKjJhAyWyMk1CZNuSrTFMDgF0OjDgk3C0Gi0giGcJkLF5Uw9kZAmZCF
M2hzNHnHeIZBmfUMZ/OUhoznU4nqs6GUBOFegG6WBY9jvK278KhUp6rpYglycG6fI4gwCT5SyX4v
C2siGo/Z7aZDnGpNuu0KK44TiOrKdyhkCX5qpcsyafU7hIecfpwey/5hOQF5qDcTotl1J+sYWK9h
QO6H/wiMl71oNPTYqrAWFub3LywqYVlSsCf9vMwRVifit13C0UMadaCH0VhGIp8/277x1XzAZ3M+
q31pce1GAfpGIFFUgkz2VWMQmU86y49vGtK4IV1fHRCftXi8NRNVaGFfkfGhIagNQ+iOiTi9pQmY
+DmMowIsOoVcMvaZz+Y8fwXngykkJdhji/FnTHMzguYWZh9mB76e3BZJslmggl1r+pJr8HWOHQB4
IdYYPOAmh1mE1g7av2wyWbmzUXnhMkuFAUkp+83WAFMzEbF7rskOwrbhNdHwW0vXmODpqt0CNb78
YFzyBvHguTr7BJfmrUv7GohxuUvUsbLXuCKnuQ7om+If8u8EXjxUhDnn2fCiDzleuGEf9I7jq0VP
n/GPA2vZNidetbVnMv+c1jK8SzCgd8ri3wuO9Gpjm+8JAP558jqAq8lQ3SHWE+Eoicsq9w9mrDXU
G/wpd2+jOM8BVUAFiq4xMNSpe2B0XM5CIRvssIfPUe6bUAxCtbQMoW2O19NRY8fr1Mkc0hPJu78a
iQDRbB2OV2VZgSgFXeEzP1i3+IJ7o2JdgbDxXON0pzVM1rcY10Tq1eHX2S6BFNunbzTF6yrg5Z7/
oEe0Wu42kBdbh4fJnYXh09an3KTP3lunxOnrIDu0XOQI4q2xq0zsBq5KKJdVB778L/wa/iGBsGeH
LmF7H9UVV9dGVuyNT/Nc4yvr5y2gy6DP77heGB88en97rqOzKBO+CebTtfwUiBLDLzMQXTFABxjN
LaZg6nuuwH4A7hYwMlumFYfp5W24RFINpyed0W+lCDHfsUGXu2bv8bTkN5tvuIlp37Oh0ZWGr/f5
ZQz2gdyVdoDcojAjZk2mqwjCi20GoF7sFYVTSMsU6HP7y0rVHe8TMiCh1L/vuQgAQSCtKAD9d4Wa
Ex+ToKtKcTxavsnRNDFy45uI8wXVqfqqoVn2ivxmLni5TwGqLOdx+G2tUDX2amJnX6HODg2SE8xj
qWOs8C8hlHGf2UOFFy4uA7Zkbe/El4btV8ptnrFK4LWweAtWS/JfmQAHtODHaJuYCaflPr/ipRg8
f4fj/02I8yONvpDFNZWrr/mG1C7RgCtzo2lUwEeXQ0vxIsdD0ClPZ7lT7DqONSusxSthrZl4Npku
srBpGIE8MwgHOPad97ib22pzJDgNXU7F61eL0md2ZqAQUI1eHyaVENczVNIC66F+IqvHPLWUaeS8
hyqBNqPg8BoKvt8uamphdzUcqLfrVTfyDyHrVKGJatjF/wN7fMlwOiaC4TN6cAeJ2YonOSDklCu3
bmXxcuEVciGT4dRhRlaw1WxSD8JkZY2WgVLZriUyT/IaWgG+oMnKvQndxy2Zs2kMIVye2dF/yjHp
kl708T0zEYOgiULjF/ZIHQL7cPACC4o1Jh2fKscM04WPs9njoGlVDsxQebkfP1r1S1fqYJXqInG4
pWReUGsD1b6EEWTlEhXNN2Fpy4cLt4ktVKXLmBTvMKCuuZpc4bgTHeJtIMNDmC9JpgjIUEyIBo85
nAkOoAzEzuHn1HTUwguaT2lFAMUbCV4OqjpNQtk4SnC/9bDuryNuVmCaD9DCmN+PgflDNr221c3c
0vvFy2q841uHSXFw6aNChfEBOMEMxOJ0NaztN5iS59KFJnYHO1IZoSI2YT6NDon824uWDveSO3g2
o4/JIirLuaMXN52MyaiTsS1Jpk2Lz90yQQg5Poyu9eVZxZ6Lww4U2x4VOTAMLHIFVz8vn/8AbWAp
bYLMmk7z4hx6TcLo73mSQDMQp+kRifLp/12sCgNstHqf2VXpv58xj2m1Bp3xP9Dt+oityydnMoko
hVOcqVhqNmsaPCp2thspDM/57QuV87on7yhoRfvm21xg0czUY9nibfNvXBjKtciNv+c9rnx+818X
tiQ6cujOE+pCpxa4B3iflQso2JIX8BUM8LHnxSkB3gVfmWVdB878hP0D/h7yzlDXhk3uRN5lAHm+
5sS7j0YNeiNHcFCORMRSVt8wqyokskpmzB0GOBjqHx88kn5MLm1UUGk/lGK8Fu6icJuc9e2TCI9B
v+uA94wq71WLsl6nukeWobc1oiWO1i4Ie0yat1IcIf5F/VqoXJpJg6n/KgPIG584yANgdiqcE5Pq
FjBsIa9K3gls0fMEObCTfHiaSmXuHEc4H0M/G5E5AMfGjDqbsWpKd6KUT3gFY/LHTJx2KueVCqUm
rjPvwxNLKbkGfC+4nRWpsX0kBEUeqA2ZLFKwh8D3EO26GPs00R2tAmbNwi/AkGa77sK8t4n9TChV
Ds0qIQneqsQCAfYn6I6H+iw0X1MEQkzMl+QjKx/CuhlneAI1IfE6AdU2xobt9QsyJeLek2iszazy
11ogK49aeqWixGs/bW6CvYODK/bkZOv4R0EFO+dvIfLhGHUmyFo81brGZPUTTkR7CkGsHRabq5vv
ZEaaXKfcT1Gqh5ul/tDp3yRbjW8pl/UrrAyQrEvTImakTUgfGSMToddEyuRCPALKCk4PmFpnUylX
49rMMSV7isPELX8QgZzhOjpM8KiUAUi8sC20iZluYuseBHAbjOYWr6pLv1tFUTiurqyb6GU9wqHb
bX28IBEiu63Yt2bYwx1cITNQFLas+vT25hbRAKI2DVHl8qgB3MthThAddfaGjYOt3N08Anu0GF3m
qlmkvBpJHRpQmLj/TOVtdUsQaFhMdIHrYNZT6b3Il/Y/cN52cKcVqwgirVCOpBNpUL5r3+qStPJl
ubybuOHnWCZGwQtA8ugy54P0pKqytPLqo05+9E23DQhY4xCfQJ1CVh9x8b6NYmHyHLYnYw3+ZpLg
H5ttINz9/He5KKYWrGe4/D9cBtHU0n13q0p4DtHp8eWo3alXHTxnPDs9m81XWEJ4qvyEhjs4yXOe
TLfji3Yzj1ZOkfCS6NHTS8SmhUMs8GobeeCBHva+qZ6gdYZwDRtZ2icr6+IBIF4C4gpQkfaZAFgs
ADKOv2UzrxXMMGWlChcjNPatCQenjgtIiujKUsmafAWOYAfY95ku5VzJ8UPdYSm/t4P4WucOgALq
v4+DgIiMY3Xlm+1z+fpQKSIXo25ICRB7lR9Gy08N1acZaR/ojNlzyfEqvYs2/WGW8JeLrsGH9jEA
mpB9bwrxYxI3jVy4xcp+GYQAUL89A2fI6TS3zriERCzUj+s74P4cW7PmjCD7lXpg/K7TKZWZskFf
0az/kyKyHkPkQo40wwqY0ctbbNIV771N5ZSmz3rsydNwENCrwFj2szP1cKScmKKwCDhCB4Q41cDY
fIofhtjXqpuTg2pas6JZoAgyfO1qqcK2r9qgJkyyYx24EDi06g5iBOWlGBxuu+nfNvLspYvCWNWn
T4M7UrpyEBf8jr8331rqTGdR+YuKCSHeuIwNCXafu+j/lYWLkWLe3JpbP0rVTzGP2WiKuvX0hclL
h0Cxqou47Hfu4UEHqkDupJC67eJpO6YxTRIqVWE2Z5VlQunhN/kBq7Q95jJTeJU7SWnnmMV9+mDx
ZLLQ3K04CThlWx4LeoPe8GPvbtI33K20I3VTEkTiA5aTsPUrdc3Xavlcut2FkjUyGdyd8NJPVIgr
t3lSQn5WKFh4vuEZsLjukAxj6wqpUCvPNtL5FVo29ki9W3y0znm82tYmrC9vuz680xhHREDxHVcv
mAEKLhgTXybtn6wBaCho/kVGB0dD6JiZz8qbgO9AmziLj1j29qZG9oQ5xg/ebDB3SprkzDfTAztq
6PYGgqskytvwqyeMxVQoG9E25hWF6I5CtwDLIiwX5rsez2bXTVCRX9ik2955o5YJFUAMmZjW5cei
75OB7dAEgr+x3GOjGYvB/wHWlZYu+MMI6A4ldw2oxNsQJzkVGCUPImwjg0Qh0WjOcjciz0wST638
aD0w1q1VHGns3QlUelDYIMwpXB50WJ241pwX0A5DmUXOcldhtmC/p/RCOKP+Z5hskofI0gwUmhg/
3VLBHasCEGNl2RQrHcldw256chvwpUJlAZI/YXClQEOW9ttuvXg8TGe+ROVQmM2wpM/GmxRJqNMh
xU6eIApGHAaud/IRv5fwR6sAan1G9/bRRO2Ihsk2w3erOiWvfA6mofY3nlvFRltQaJItTy96DbXv
KuxHcbc11ihgUNerckIT2euJnNmJh3ZV2I0uwlRsHBqFIE9ZyFBIzp5t3gEuOGMGSS+ka4DP2cnr
v4bVl7QjfQTtNt5UgJSJhyhozcBBPwNQhttghtvWywWyjiTXv0MLPs2WtFq7jIHvX/gfnGcSPvrf
OqO+zPVFHGlY0N4Az5vvUaVF/2drx77wzsmy+1ND4WGQlO+wy7WA27MaGE/BsylhLF9y1pHvwPNb
MWDC9ONbBF6BkhFean82MlKvu31S9LQtantxgfwjOq5Un6yLlrj9UXEMcnrqIwHzDihnBYKpfTML
SbBwboMJ0gy3OambQ2MCAKVnNHeymrxcTw+1nfTd9kiqyDLDACpP6dK3LLqlH1bgLHkPudFflbNp
TiTuF0X1VjymOfp/Rze595Ik0q6UUKWKraek5PkWjCn9tDDDQkZGL5QJHIFISQ2hEk9HKyWxN9f9
YX2wjO5ffPW0fzXSJwvZgjoqpmEM0fkeOq9OPVL5IWopwGKu/p8SVE8t9S84aY+4n82iBtHY0t70
NRC2HPNQ5LzyooAOzx18ucRcCoKeNRjNK98bFi7n1LS4ZBvXYFzJk4PYvS92yx6N069bJWMqSYKI
24uGz134VmKMz8+Ce1G02dTESV8W3aZaDaS9TdeMVMKYCKw5DqWOIg+RR8Ja29SPMguKCuZ2iVCG
RxsUT2H+J62jpwJsk8GoJ5sETi9Ks9ulMqeMzPa9xiyaH84YfgsFJZ5ggHbVt/dhgg+EcdsY/Pic
dS5Pd/n83Q5hgZxjJ2SF4ByJXH39GY4UAyCiUtJsLES9xNXiekKnl75a6OXRUTmMdLLcOeHUE25i
bB1OVMc0oC31fta6+tjxmFJc6jaDhuXopiIkezsnyurKweI+I97pjqSxUcQIFCrChV9Jc4LlrxFi
yxa71jksrfx0a2knzze4DCZmoyAvj3xex9gVmNtlbi3jWGp1ime2M47RXEkyDlF/3ABuiUfFNbCs
sneolTNq22UPx2bkJr8t1Qm0AtrAonw/NGEFNQZh0+NZ+XPVr4LjgQXT9Z85Jjopp4UB6cboo7JT
3Vp6Zr0468UYyNmI3LUaKzPQ8cqxCaeW+HmAVz1gBIY6h8KWVEdADqWxAOdB/Nn9dXWF2MaV5Mr3
41aj1tcLIbQKF7jjPiBcP0frni1R7Qz9kgGA3CDtQxnphpb4Qd9FXYs/MshX0PydT8dAg0aIZtMa
XL9uUkgSk1ArR0qDQZS5Ml1x3h6n429N2QKZ4Vpk0IuyqSKa9mgW/64rAWbwHRU70dIABBwRE8A1
adCv/TBff7vxUhW8IBTpJvw0rsFJpaaGC2NTIiMVEUoHgJ9FqwFFnvRFLbJCdsyENvL1bbVJEOHI
tpsI/yDjW+r8vkcaCrXc3whV8Pj4mZK65t5pX51onkERHxcvrsD2YVeUgGPmel5YgSwa+/zU3Ozn
fefl6WJJZhJZmi9POc9OHSSLB5RupC7cSC5yhPO+KQskdeHefOUBYlruOUTMLkbZFg3ghjLlNDHH
bLnGoYUckLo7wF+UsjeV/bCRgEgJbN16HtWusiVx/IKFE06BQlrM69qd80/Iy3DIbgKTCTaW/PAy
Q4VrdbnJjHEzTbLSVeR/f862BvW4sMIvo74+vj0hzl7iOwAaYX/+ehWOTuDOHP3GNy+KXzt6tekT
ChPmIRGmsWIdZ5NyUao2ydkcLlqAUMO3T1ZKMotdMm1/oQAuPdaZR7UZAQgSPo72LpS4XY8vIBb4
K2n58mAoIHh7PEpAXxB8wyOy5eEKu7Yuk7owXmlSMR2GSwFSLiSC0VPIfh7D+nUQEXLDbpQSFrEm
sweAActuNz6moMT824ZrSQIDLxZlEt15wWl1ThNJgCPhr2j1JieRMRwbyKhpAaDk6tUAydA6O/HH
1Vf5PmpA/IWhbLwCkVV92KfN0RsCd+SHLqTItoozvp73aA3m5MPgVLojYIY4dKFjPYp4wJJN6l0b
y9HXc9X8AEPLLGYmzP9T0LT1/JF3cYjbdY8K96DDohbtr4V8PF/hvQgrOncYY3WIkZl6pH4VcifP
8KJphhW0M8Q2uRg7rfoB/HdDGdYNFwsJvZkPBNr+/D5CPRk0Ex7XKHxgGiQKn/64zXHe6lJyrZIS
TOlnbcY0hN3DAJBRkXxpqhRucnNc5yjrP84Nu+Dzi887JptPUWUO7WmNCowpgbZASxqmmtRdZicc
PuXAp3tb7bGMb7pvKUS6b6a/+ckmnBS7Lc3kcsVupWEXKdlVx2iXugKzW+rI6s0nFfQEdVjohAj2
wIeGoNr0giU90jf7OeqBL8lFtCkbZTNAUkArgFtZBQZ8dWJAj3Cisu8LP0g7k97q+rwy62rD+gof
ftRdgfiCjVT13wFjBZ6gk7B8nwXtlJ73sYz3QZrdYE6K+xz/a5zhfJcBxqZ31j9O7YiLZZXsbSl0
F0Cl2vLvFl0JcpcFQHUbaozlg0HIGP8ziQsuC7ilU5I8GFaSHcvGGZIXj/AwRkwaDNxr51NJhzem
IRzwF5S9u73SVlbTsQPTzuAiD/umO+J815/BLWmY479Ye072DV2+NBCY+tAF98qGfrg1cB9AJMmg
xM33uPQsxBZNIcApJPMPBSGsONHOuk2XSEUef8rpryDVeLnkls2pSbkp0FQ9RL+z3ZnOPn9NGQ0f
OJiY4Y3YZbhgL+rQs1vOmqWSDubRRaI6Hxn3Ib4ZdlZHTzb6MO1Vl1CKHtB6S2QkvspZly6k0SOq
USVbcUHF27TwAgqf8qCOVybSuBHoz+FrzlNz7bimUsZvbWigHpaoB8Le0vrmHtdR69F5j8Fm868a
Py8KsZgDAs5BddwiugZoqzeZE31oa63jLJypwNlP2gRaN5xjD34qU+E8EJ1W37vNs/NBzoVA+vpi
hgNjgo+7xzMlU1StR/HVUkgsULmpGx2fspF3KtfV/3h5YCkrK8pi6FezW6O8lRhqT/f//wJnwJAk
SfobLsTbITmxScCyP495rn/BOoFHLKudMZBl7PjmRi/90VN9WulL67rtKP6/BI+7CXEBkuvZ/BaV
ev23erbiX41cxEZlDYxBQ2tvVk++p30FDMokDCsxmS6X9vOk4vv06co5fTXnag8mSidnP/jsdTzy
OLLX3/D5xukSoXNxDP/t3jlZV4O1Tp2JasOEsDhRgkqoAny8o1DWphJz5ghWvhzhVhtRBPJaSz22
O5v44iZ/EZshaiwlZX/LP/CHnlnaqD7tPq5Nm/YKHLMK49dGQ/JatAOy7e43w8PBiZWDEoBjM3+E
p5kmdbMfXcQ8PrUxXckcKofxxaBKrLX8q2d4mcI5jzcsRWg+z+taBSiEXTkdiqzMPLFx8xWNnY0q
sjO0MCXYyAJ2WOc6iThH4oFb1C8tUk4gyUUT2pIbrkGrVemWFxWZZBlwwowfeP+p+SpcgMNihReP
z/so+xGVVt4Mane7oM5OlMLoHkRa3m9fDC6SM0UgQlC8SNP4LKxGz9erWBN8cE/TrMwtkK7xqgGZ
bo9iEdTjvPE31m6bdWVQe8pALXLKQTns5Akw8oUYvCbWRYNDJ7X7lS06YKJo0nr6+i5M3jrN4E5z
Z9ggh8cp41Jc6PR/t7B92uUAxdklsnJd0mpgjUNDvrrUvl5xPEFtBNY/z+KoPwdun07JuX7JDC3E
fLpS66Ma1pYbXNUyyWUPqusejl4xb490a4fhUKUZujVrmUTtLuRqlByh4+tpqKi7iDQwg8eOUqej
KFn3FSRBJ6OTsbLd9uZJfcRCV00PhhAuzeME0Xluj9Tgbk72l7TGzD8CpjHr8NxhwZ5pBlDVJj0b
pmkv/aeW/WWcyz/TZQbB98ydUaZz1Pg8NXqXoum94uwVBDTuo3n1sZpeChRH4zu1gvIiYSR3lcCU
8VD49ZT4o+2MPwIhmTDhrd52wc2Sc9boMNopCvfwTatMbmoHirhofo5Z6LqgSzHAsk3GZQDbN/PT
SGStzycBrkjYJnEAKZNTSF/Hl4di69VwRbAlvoD0u11Jroyu1L/hjPNVWr5volNHWFzvayrkZqgQ
mNA1zdj/UGwuptQNTTQhI4pgMrMxXVfV2DveRMq4ooRf5naLRDAxbE9teM3uOWO7FM2Ex7VyhS60
WUWLpuWWKUKp83Juh7TMYZ3Mr1D0XLBJjLwDZMqg1sw5+vocpzwTfQSaDrIDuUf0phxXIYxrQX9L
q721xJ4GS7bpWMGdBHKKBkLanYTbJ1es4tlRNgGoWMVXbWvxBB1fFxRAkxO9z+cV/nJbHVg0J8Lq
MYEAibsRAjhoauKCVFb0CcbumEAKP6Bp/X8tyHgBtyD8tqjyKEvQBmpTd0Q2xRgKKYAv+UpozrRB
+1OiNxyfzPxEG6zDBtDKfp3zEg+Uo/SetVZ0Tcy412iZYwFNQ2NvuD9AN/FOBvYqq673598JbfAS
z/nq30tFF+fwSaVm+OcdSPC/Mbgf81Sd5j7NkQCZAhvVUB2gE/huxMjoZ5veJ8zkramRmg5RLuMr
kC6m8nX7g2fe9AiE693OhDeF9L7UJMhkpnanGdUfQxicj3f1jYjwKggsddNsXDXB1wcMkMEyH5Ad
OG93IuUneurjxlP3+9mmw+dHwZkI69U7w1Pj5zpk3x9/EiT7qWWzQ+tSIDF+kAygEmJD4HfhliDB
uPtVSNcnlfM5ao1RThtFcHFTmYnRhAZop7oU86oWFnW24N7Ekx7cCl5iWbP45pQ6lgvXX7bT5r2t
j2v/FEhoimw+GrGlngz44MMZ4RiVIYAE0/AQeKqeEnwyhA0Njr6D7q0ifj1SZE8xlA5u/CO9Ru+7
cxq2fp3W9IQX4Clq5JkxsTw75T/MxrOI5x9zIPMfO86iuom94XkT+YttafbIetCliH94Qu7ZSCC2
mWWwZbxB7ERqMc/wENwnrJYGvBoCkT5L6Iv8GDnbReZmyrEKylJQo5L1Ip0dp4ZEtMnYhHeoq214
Y2uWqaDQ3Pq2dMCfzZsXPCl/ko80I3Kqgs9ZseO4RhDZPdwUx2B+XB0a010uiZnQcxDtzUx43CFe
YlK7eC6QkDPnQGr2siIFFYxYLKAGK6/oQaCDtgwf8BMLWMrW6+8we93SveLTMeHxbyHbprw11n7g
1RIymFGEzyhfoS1bKSzdSCb8fB8m1WZ/maGuTzY7sUGe/3CsMlXCcxkhE8EaEDYWR+qm7HJ5SsGY
nAMqK/Up0pIZL0nHWnvjuggzJfr57pdnovk16pRPuawG7OBhqwkj/e6bAEC+nk6LDs9HacjhcaUX
DBj4/CE/gjcvFDm6JR6pj6QtYEX3+2xLi7gg4C9CbuAg/bnHm/iar6MPJO7WiNp1A9P/cWux18I2
8TC5NFQE+Xbt8qQx+jIDtU4jVIqljueg6Z4+KhM4VhejScozDTi2WYJzVWm+3aRkpn7vG5k4sSXE
QBfrH1mPTO2Z85sza0MPSUg8vawLa4M+1iLVo3rRTmUj59FqfBBZ3KyoCeFwM8uNVy/oWOLO6xZI
W0C8Oy0Sv7QEJMqAsKOlSRizC7DaPZCj5mQe8RVYHS0udXNDVuQ8HzVbt7CxERRODTGWbmrjKJJC
lnSUp3ddBR6fC0AAnlF/p9DcGwch9v1W5cam35/pk/K/Uy5DFeH/kEq3QeA1LkyTBi6meNYSPF9X
E2GlBFLsDc+XCjhG+bOCEC96u4g/FYeiS9ZVGxZ0FFuthvE8O1MTaU2Hw2DFazwJc93GEEO7MDnK
COpQfhzVsP4luC1gAvXjcSGjPxC7Xr77IFLqwQLzKX9F87kXNWilTM5VUHQ5hgw2nX+29rvW9r5S
StlKtvO1ZUNqZCC/fZQE7kK/qcp1FGTIhi+0UZdkFLwU0ylstZzmOsglBJ/xg3aZgeNpxVtJ/CeC
imidIETT8HPBC1BOsfAOb6N7p1RPBLDwRvcxocpaIJFrngIq1MEuocy+WOhb88rB3d3Oy767+aW6
R2/e2t/5oEJQWBj/6F7c0x1RfndNt1aoa+hmobhtnCEF/oN7mHIsS6rGVJFk7AB5jzzruDuruEh8
269SlwBxw8JSiPwRneN7wUNyfdddUguE4yxutVmFevy3WGXdRkDWeAm1r4Yu9w1j0+dD1w6R4kjy
W+zLq7QGhU3D101+kE9ATY/x4XrtE3UYN5tS7UaJFWUOJsn8DAQ783634W27Fl8836Lrbzr4ECO1
ZeRJEgMxU0ItyLmSn/w7S1PRSozD3ioDH/uEZ8x/ZMI1RaYmUAFWwWmAx0XUtKzsn9btRw19ek3T
hYR/+twtN7CxbT20SlxYrN+Qch7k2mwn0KsJ9ifPLNku9MBxl6zYUaGluvI+OElTKF0kVVdwY8R4
uyn5aLeqFN+QFooJf5bAlQd1EpXcZHlJOcxcRRB3ZTz2nwWsk1dXMJyDfXm5XUGjWzAlkz4MYpQR
jw73vrc+FR7ppvSGytQDDYI6tGC1LFUgMjloJ879mGfCHk7lMJ1kimAA19lm5icjhw6VVOCTh4uU
t2WDVQXRRz9qUuy/SIir7eLHAIG1sjYR/SGQaIVVarjXH95PXxGgDUTrnbRWkGn/l21JVWzczs/7
fOuqlmEUtNv05Zov1mm6xZlWkJJSkpKWsmShNnWqRLouPZRP1gkYO2SUPAehtpMB7unsl5PL9ApP
+p2IycvYUp0fUU29nmYEcIUQOO+W1NxEY3nx2XBGH02g37gDqughCSsS5VpxGNQl9HQaua+4eIqa
BZ/0Ae08n54IPFRxPUoL2oRx/awVqMl2ix+/iqzXolk7MQ53FYFlxTQZBJvkeROX8MnuwA0gYHJD
soRrGUw6Nvrag440Mn/MQ2alWHOXo+0ZA537Ri80DC02IcH6HcS9hZEebXWnJGDYLSpTQ65bS8bn
F1zUoavvZb+AfQ4DBTSWZi+sd8JsEXa3P+AS3wCGz/XFq2DSHvjTc5a/aW89hSKtCXHffoe8ZFUn
hOWUrZB3hxZEEd46AH3vBqaERfkV4Gf1ZmGHj8cGj88/PW84/u/+SQ52vNgLFXQMiM5nphVlGbhp
oAE5jPbWqc41QhjBNqDJUwox94FpxE6VySLgRtZ0M5IufRBTpy/g/NR2maEoPMb7B45rT7YQqAFe
fvFfcoMo2q2aAlBX/nrWkPt46bA7WFfLWn6GTg3/tTJ2JMzaQd1tzhq1sn+WSJsdbrX5Y0xSCSLw
R/qjABqsx57XXPKwvLP1uCQgHSOniELsUSDCJvvwdguggEm0h3p03aMxjZPPYpxEffGrW3yIRgly
+tRy39dcP/F6vRPFewEbRWExVRxkkq8J95JGgltRcIDIpq8PtREsMA9HvsZy2dZ4CZ/NLrKhjcLO
av59y6IbbyFBTcAxuOSsOgB6kfRaxW01IsIobIGRtn/blKBCvggf53wSWtm7oAgPDTIMOBXwND2u
yyqAsWr/PY3DxmyoYzXkYkr7AAChJJHX/PRcWVMksNeupcFe0kN00xgEBK9nPWi/HbGnNkRerZjj
n6S2BH0xQ6GRb4JTz9v7iBVmhE4iPPcpuDTq0RRvf83WOZyxBfr3s9vhiWmIA2l9mBuj1M8EBQd5
6suYP8itMfY6VzEObnB98vJRUTWWxhB7/V1tDKbhayEFmLvAmpMAJmxz4ay8UhVLms8GwaI3HcAj
aaq38JtQyG2FVIlghgwKvONzFQTCEhqrJdyxXkQ6vZdL8qVoTjLpAGaJ0iSDv3qV/mliBNJJRtpf
Ao5EM84Atr8BqZ4T12uA41jQv+J2pKf3pM0wGZ7UxHaLENM7nqQmkqZR6mYJoF7K6bl6LI69pEsb
pPHq9q2GkOCcGPIemy8jPGI//n85s7rrkMa8uszroD3lLzxnKT20bX2K5MVvsM8+aJFrE9vZBMul
R+lVAR6IC5Xu1bTkUvduEJqhD2OQp9EAQmjp46AU6npcGFVUrNFO4FJzAMx2utcm7ni3TKlOXZJe
jP/nM8Zybk3PheQgi9FI7uXDKBuxL3XAR0sFiFWQGKvfjn2MZpUTB4RzYkKYvlCaBdzyFS1X3/mc
ry6B3NJ/pdXUQ7FtCm+0idd2L9tLuOLQMfYffTS1l9EFfK5O17WCMPEmMhtjHJDUVLQdoUk+Yl50
pk8vcv2ecKl4npPqY40KMBuZlg9w8dVtiI2RQBzwAakAuIJPsljYG9eGBDiJHcL1qD2Vr0MrmVXe
C0gQULN7CV+aW8RRf0Hi+1dLj7yAws+85ESR5mMUEEKu5RgyvtXYFlDoBN/sTqkoQsgnHCr7C6eS
C0FVFW24uvtlh0TRny7502LqnddT6BYif/tXtNOjak0PfK/KRDNAy5o+OgoBgTiFHQ71MZuwVXkb
JldT85hIVcnIvqA8U0n8RjsIFXrYgM5k11uP0IZ950/2lgCYGC8Z+4WcUQlxQKYwv5Xz1b4N5zet
HN5CV+9+MJuda+Yg/6ej2506XzVzExU5CjgJAZgB0ebNqmbpiT7iicJn7L+yxgFGu97BB343zFNs
6GEDPQ9gNED+ZdtBkAEfkBQtQVlXbL8NIcNlAvD/VpbkqoCQP/j31+sHp2oSPH2mWo/ITTH65090
84BvDMb7++tO587MqzQew9SVLQ5tU2ZWUpgnZ+ZtSKGx6kOpwwn/PlHVGRFeANkvbln4N7D7lR5a
M9uJNG931F/KNKVhpPgqBNcKEOdrsJ/XiMpJmGa0I+sqali7AkEj+hva2FShz6J6QfpptXJgEA0Y
xlG5uzbgfgELTKIoB11knPhTSaA1Tu41RfdRITD+ZeR2YarkbHWNGyleXN3dQcO+H5waBzvcvaRz
Izg+CEvI6Lswby8dhGtw8fe7Q3fdSM1bgv9rV2Bv+szgo/FdkPXtjeQ2rS12TI+9PU0gXWmb8NRK
bIXym+nS+0jcuGucTwbt1XJgLwqFm+jgWRpBsvF2r2zdbZgO3nEU+9AaFnru6LYnmNy7uI5asvyj
1BAiTJkkX+9Yc5vHZUmINhFyb0zAVeB9cE0x+nPW7fjAZJj+xEUUT8fIt4C88lPpKPUruGLU6SPA
K4bj5SitCbXczJdsFzyVrUQesi8/vTHOdu23wa+9WGmeH9AyKbk8o76SUHjOXpfkRY/g468mCe70
Ug96R1Ph2WMYLtJX3UaWozoVenQ1bY6meIH15S5n+w+bSKJSFfUfUNCSmYqGwpWH/L/hhsurI3e4
5HYVgOWmDncrXwWvU/FX11DZ7t0eR0j3qg70U0ukLNbCrSn8Jdc18imgqT4SpNsiRS3nOnJ0sXag
VZfU97BQICZQtexSLAqaOJl2IZ0337JZ5HDHSqEkoLSCJ29Ucip3w6JwtgND73NJ3wnn9CMm1/x4
0vaqTwuUFJCY4wZdzfirUnwKNhFmEi8X6AHJup+A5ylrjQKRs09VC0QSpYt+s6NeeczdvMUUDhFb
Kfp0oESN78fBvn3U1YkR4aLNMmHhw8ZUzSmpBc4j5rcWe2K2m4PYrFENrny/GK2vt2LRBRNy2QjJ
DrF5tHSf2e2988NV7LnIJS2gof1Tj2FVPAPxLCpkxidsb2VEGCFsZ3xCNMcy7yi1jd0OgG//CXEd
HDGBspBImf/WMnyElW86B1/NQg0oq6HcxNT/RWIfW18pPcKuXjAv5shEh4Fct4HEXXLCD5rV+rZc
ClBPyg8dqOzh7TZw08WD8Q1JVJEwozQFrR46H3hEXYc7visKHv/yHdo/3vEoPlMdl83FLXn0sbA8
VKqRT7VnP8d2X84PwqtfK5uYMo8DxCeUklUbw1VGZhxSmJRsIj528MWf6h+TCyP32xrK7Qpmhb03
ipynCvtUSzXBZ3gwC2fHSIyql+8zKUFhedjvslogdotWXcRD8w6CSRAxgiAq4sGf6uGBnu/zvJMl
JF2RPfWysREA/Aagm1tdIBU1fH+MZN7mGABXdYrQt7ySbRJcl3zDvCHbOz7uxhZMoJbO4hZRdH6c
htYl81gjQYpZLbJyE4/eEXQs7oA0WMHiF15eKvb/8XHz6r+Xsp4R4maTczgnFHczckcTejWdDZED
oQ3+lKH20CVgpztqdAAusBImzqq7UZLmUfg9CHuWgbpOB8JdmsyurnhFzNph5uGgfGAKTiOF+Y4g
HDYJj/GEzQDesPbOUEbYrAcpSd1YKUv+UfdZf8yKfReLJvE2BCqEDQQ+A+yOg8kON2PVBz0m9yTl
OQ7PhvErBN2Ay3LzQ+mgml2LHfjbcmkca8+9j1VumYcvv4TAykQVl+MZqEXpKnzt9MKoPfWlUcUT
JeoQsJZv7MaJGOS59EyAWqBW7TyYkZgXQ5qK69eJym8rF38oImoU3UWl8DryR846rJYkapjeGdsv
HMtFOHm77bdbvJWc3Y2o8/vRmMNsd8WYgJZ5AV7zU4gX+Q9mEYcFmMI9BYMn0K0T2hZ3E2YYm6WS
CxcUgrURg0AqVI20SS43BXleHyR99CerCfdzGvfe/oRd+Yg4cX9TKDWdtmcQt8HqD67QtW2PNQzz
nwd29HXGxouK91jjr5OwW3heYWDgJ7tVA1dozqrv6aJL7u+tnaOL67sitoafqdibyMEhQln2bmwX
yRMFS97R9zNCHr5iuLcwHpmIw2MMghw4clz7+k9goiCeWIkrwZRbJn6f/DE7z8bxTUXNYOqSviqr
X7VxD93TC5vXfaExh8Cz6iOPb5TQRzyv3QFnp0NVIjdy12FM7SGijZZSs3jfxE50tbA8NSEUDIrG
3rTXf8wzKRboOA3CIpFAwOQjFQnPANJoEfEGiuR0AdzViyKf5QgWSCNyDZUwkOnqa5QSY+CeKnIQ
4XsNNs4GyUgakrpypb1MjjLxobGZIkXBE1pbAXvaynn+tNOaie+xvB49rhfImvDoN+Keoqtl+gw6
ZJh/Mq3EAoFl58WaWgDIOY1Go0qAdrtleSOO1ooKGKiZB6lbIWrLCRo0WAv65SSHG/O+dyMh6Icb
gqU6hQxkz50B8ajoQaS1lcdwz6+oupRPXZkjj1B0Ef7l9MRdZjFHyCvmlisU+9HI00egW2ueXm1/
5heQCgoly0CsffH438SISpwIJ6d4CldI+lC6AzawjgBJB4Gd3QfOt2+MnHzuJBKfAHOuX1AnSafZ
NZgm5W0v6VHIgkNpIlFPN7EgFlYbxitzS0B+CzrNudbtEMb+ipo8ma850x+FNuEzhOfW+Lmd/sCo
jlml4qgBS52GASL6PjVRKx8EBuTY3l3A7P6lMafGrKOsIporLNyA6b9nCyd6YFSAfr0L1yxSOqrJ
01Rdk0pRU8uYMGBgjACZgJHW5butXrFYMgIFYy9zIaokbswEO6b3AzxoqAABFLHOHk0euu4zurGL
8taSsvQfq9r1X+70oFAzOAZC2isSbIVMGYdqxIxfeCbu9riWk2lqd5WsjVD1FwkV5x7zaWpRAPy5
I0HpXp1D4Fo3AuHhuR5SfzyPhj2uSadauh6T59rSuk3DGYHmz4V03xzZ/YQtcMIxFRcvS9VgqPts
ah1HPyLIPX59tlrvdx6fZSf65A5UWzgCHdEISa7X6PVDv0etrk4fUFpKcanEsdrwsGPkml3/phdT
NlFnlx7epd/Mr4Xw90D7BXxprUYaozon82N+20ki5LQWbnNQHjyXOKlexBuzJtG+t73lUkg2dYbl
KBukR2AoSacYGQGghxT4xAmV2BkMgQf5844Ta/mkAQhqm507MrNaqekoxRC5fbwq76yuUgqeAE6b
wwPOZkNWoYSdJct80WSIdm66ft2RSvXHmoMk6GCO2ysBvVGkVLGVZmh9+fH0YIh+Nw/bFN8kJU+p
z3lRRBUYOnjE5nkrhu5G8ZjplDKwGIrE/l74YMTQNEt1ZA2MvfpJ8BF5A4iYD6IHdoMBXgtOIjr7
B5LIQC+mRXnSjH/S8eUm3p5P88iXTPB4ZSYCNUEV2kU1xOwdAUBek2nLIj9T/I9NI2bRSxDohwCd
3/4bVddyJvRb1HsjWyVESOyvX24i7CDaxWZmjNQnI0ksErcuizpPiAOMVt+SZWRP8LEjsq3M7zOb
soTWRl7KQQodfz8b5UH2UDt3lXgoezH4+oaTsWQMgulhE0JoViUScWbdAb+NZDFUmlSKqILFCTX0
iG7ZC3WdsPgVKM43W9TQb0S/Oh/in4Y3mmU+zclRhu8DNS2oW/PyDGariFIXK5LfCmocseoWZkTj
b+H+MC10tFle6sY5UNaQQPnxv4BxfvGXAyv40AqIu3O36zxo8yr+swgELK5Km1k5B+OGS1SDph6k
69kJmTG5EjxWOI1pQOXiF8geQgntP6iEOhQDopoz6pr8NSvvbapGDNUwbe0Fp9vPaEEjlCh9a69s
o/Vm7KSHiyPJ/TEtqVwZK2kb2ELuWOA8DPeklV7YN8g6FU40aw07MzZwKy5aWSO5eQLleDtQd8ED
P0c5GqIs+aBFXHj45c9N9VlI/tcWbOTd8XEuTNQfSug+crOev1AM//O/kmOM+QoU8Ror/dGvZx5x
8nHQEjjp3DXpH3qX4L6QKcRQddY0ph2Ii1Lu6wK9+zcrTSlhU8UU7XAtO8o6kC27brId/Hl7f9WN
LMXdkZZVmWYT66WBoel5MfrmjtUEHeaQ3l2b6X4D9As9pjQKPsRAcGzUFEkxqah9sA9ouSTiKgiU
aBz4OMhlRjKw8K7+4b5T6aPD7Ng1Ai0wllnrgnliw7RHmzmtSu3xs4MAAL6KiLS0vvtQqNWNJtfN
DC8zx2wn/tKupOj1LRE7aPkMw5sBfw4QTuimwMnSaxFiU8NhNa6HZPcrWdk23/4/4NTs44lQLvPc
WOu0cmA05+vQ+0Diq7EkJf/xu5pTuJbUCwAuSxAZp3mPTkUwZzR6y8tHvytzfYY2kGuZNGkWFEsw
KOGSbnWriSXamthkLvcBCMjkl6QWeH534tu5z6loUyt2qL6FCen/6ekrHBLhXVwn8VRPcPDp1gek
IHP6qbZ+R0s1gdcCKAt33Jw3+KyAUCsgzO0dzRBqnVAUz+dNGNOHVgSOI+WIuOc405CImolp4qdA
+lIoy8IJimik6M+PuqydTkVRsH/7Wxs/2m/mCQcSQsXtzXHDn96j62qak1VUrtXhw44dI37rlnzj
V6NRgmBBg5lCLtraDGeRmdUQP8ycxOz9l0ButV43ZpQI2/sEHEuJh3HlpRuj45Vfdp09uk0gBeSm
38IoscA3e/nk5WqrJgN7t19JdYqKXEBx8HMYySkvRvQVQymQ02wvELKX31lPfG55LazFosQchjex
wWM0A6iePYnvDIN3346oPqJL7hLr7g/ZqQIo2zSVBuix325j/7nuxesGsw/poAS5fpDvhTGEIWN0
62W7/lhmPZZCK1nvqIGo76zWlZIvj3y+5o8Zy3aQDZBfv4qZ/MeshLWSGNfupSlVUl0xnN6A12Qg
9eQTylpiysz9lsB/TMC0nRzZ9/6N6n4Ks9TNu0OOnYQyXbsBJCDvj3wkz0/ODA+z5PDyDGw8zJ1/
9+Dft9FqCCV4WQKPkc440zSthsTov+aMF54QqSFQSYDcMUqSkzkU9Omfn4+kOd30bWE3uTBWrOx4
DkA/dCG3qRhyWC1wBlpIrRqsEEhSpFYMwO5LvwHEKqBUAPAgDL52SofiBPm8f4Uqv3bUmtwO5soX
dBaEWGuJ9d1Zl178upIo7AY+KaGFVJ/7AI+OjyJKPCvfAwbYF5BAsazv+gybRWIUflmKCCkldFUa
eBiEs3VOmyZbARkdPzYCetmtUyIHfb02TjWzYyHNo+3Oo0xEnUU3YM3t72BazYqv/D72dmI2Z8pR
pFZJV7sC3e7nPaU7be+wtCo8/SeF5np534NwU6AYVwSDXJ8NM38KX7aOkJC26whMwkZXZj4+ODhZ
iO3UWCo/V1BarS8+q2auTTh8bcv0nGdCKMc5e/tn72w0vC4OveD91VFHb41d2Z+Ewz26ywLI1O6I
h4/XFd0UXIaJRoohuNi4PHYzuqAjl52wkGJNMLuc+4CLP2RSWYr17Crq9LGzJkzkEkQKDANPwYK9
PCqCxT4V57cMxvtBKcGtMssaDfg6FZX8glC3eILqXZ0+R2TyXzCsypsaAgDyoaBiBQAeyuvEXT3w
Shvayhk05v2PIbmWF0RhXXzu2iFyTWrS6La1jPYV9W3sl0Q5/ftYQZXzVWG38Wte7ZNV2QVAoVs0
aDe+4HukE21zPViQBwZrG48LmvYh/ufgKAUNgv9CxQZCRqHtF+QOGnZNpl0yKLsXxImL5hy+0yP+
xqGVxIwUIdgIuB5YNGgAAZbmR3eK+949HVv91bqHfyPPnUFHf1KtpQxdG5gxSPymn5LQOD2oYmMZ
FZVHI7VF3AhTHQjO3Y1omcyNdcTxPceuKJJYwbHeu52LCMtsvGDJtoIMxrf2iqqPE2+ttJ3zbeYg
jPtRRNs52/426f4NxGzyJdXRPoCed2Ww3XobbdR1HTsW+Uao02VvswpdEuEUqhisS6lux54RcvAu
sd4/AxLFdDyldWwYXPB8kRhs+NubTGu/nfTc+A+o8DtUybmqXyClYiAxmP1iC5bC9r4RDu0lq+WO
Xocm6O2+3K5SFbs9yz9Jm2yG4agnFMP3natke4fo1gFJXm+8YgfwqagUopyetZWbFAMyK8uDLn7X
GXMr5oVBQ6YFIx0Nd/ljD8/L1vEYSzxgTCc6yJnnurxzIQgXdvGfimmFAINSyqgJbaQVMxJf63P0
FtZqja7lQVALnChaX7FFCO4cvVFBlWodAbBm1KEV7DzN1iCEcr+WL0kxhDPPnUXkzJuV7n3yIlZL
3bI2lVV4agerMWRdrtunRhPFe2ZUWZHTrlPclJ7EhpoPvm55SrciTXbRrBn0LRJlxzSqkQJL3Bnh
htUpLuOknwr6c4euWihRali9atiQ8lZzpy81CASA9NNFrqx0HVj6F6H1eyptSZh3AQJBx5XFEzGn
KbV+PbsIM9Y1syFuOr78PlLtXgilqSCwaAJxXKVv1R4eYdhCGkRwbqbnrtu/s0awPdxML6nC34SL
SS28Xn4nE+6dl5A/0KbpidcxAwkW3FIzSIfhUpGkOkkKZ5nWn+9uPnziUWF7jV21uV6tkubmE7Eq
kWk+M3iTfYA3KEAQ7zIfhi93nyxcgbJ8tPtnxToPhEp8t1ImIrUgXCGPBJ7ZRuaSQPO13l4IohG6
5JKh5s0r37WMqR0AtONhON3ELLwVpeINUZ1o3ZBpJZ/8a9jvAxun5hnygyzNj3NW4O3MBZgKAY9k
1L9FaSnAVIdq3F4UJwWfEa0BxdaNupOr+zqUgfkL9ZYadsogFOpR4ZFC5+f5aNh91N+qcdMNWLQJ
z3hL38anym3+d1aJEy/vETzAni7pUV1DL2he0N37l6UgCtdXoPin5r1f/BKrGRodQVmVpySD/KIv
3krSHqFbSZLUXTHpqBiXMuArJoqIOtpTSD7gp4+CF2wKzcDsQqpg417L0SDUF13O20fxOVfuwHLW
suCbV4aJk2D2itWO9HcaV0zrT5zEMXQuzKoyt8wK+JQPm9TJTo/5QOz6sHZhQ0OXn2VtCaCmZ0FO
LvERUWtLkBcHYaKwOvNhQdz6dLtMrRxzw+NWk0wvTGUYrsTAZTyeZTUu7WrGM2GtYlefYb3aB2MN
U+3XPPytvW27/Hruwpu7+XgfHX0MJc3tzyVtzpUSoqSk/0fHTxT3MbfY5kgfbcthNQMC2DcwAcql
kJALDGgX+FdMpRMNncAnKJr8/UfTP8kRKrG5Ffjxgq6csWh9YDWrVh+ITZ1LJ8l6qActX/z6doWf
zIwlIxs8/g2ZWymdsZltWre/3azjnx4rJ4NZ7VrblDbWp6udDp/dSi6hcacAejGUO9Qpk+Ww1NNr
MU0Kg0FZxo/dv5inMcWTSezfLvgYeNp9BejF+bDwQkt9kPesxu2nefSIpKlTwVLHXDFXUVtvLpar
dvdq03eMVUVL23pWST1e58w75QK2MEd2/yf8/i3CZBr9hZCRpd7oteaWc8y0wL79KDmc0RvmtrgG
HnIdvwhdDJTZ+nQLQzh1uzoePURgUUfmWS2b8+jH18eJpZgi+7qt8EslON/JCFEqWk5CjD3M8Kwc
JqRsTr1ie8C+cbqgMKmYCqHW+DCaBChesjiHLS2GjwaMdSfgEwoKsVq6KFSDROKTNyXl6aI9/mks
s/957lCvIstcppSasV0pR7+Rek6BGHlqlfXVGL+fAHtEgshZSptUammvXQdN04JgI+qsX4MTZZwH
sWxSNFZQOGmFgwE3H3r6mngU0ARmoV00tLETI+sDe8P4TzLShM42H/lc1nqcwFZOaOSk1KOHCdNX
+GI5bQGuee13DePBGWoOwy+QYOe6YwZREYlladjVdDF3QkUV6uUnUkbUknBWX28gSIc/RlDxA+5D
ghDe0pZX+Y7og84pKWu1joTe3wEp+c+xcxx9A8ZibL9hHPmn1KqKRfo1cnvg+y72C73ZFzuuSHd9
1KSbZkhiq5xw9xs9QRFCz4L9EG3HJgF8ddCPY2j9jNQLyF5TwuIELG5y8tzRP1BaXHqiX0LtZA/3
H23vlK8MgDqrGhuBFuRRoXxPGkT9V4tW3omnoq2za302pQPBGcllcB471YeDhN6RV8pIdI3aDuht
g2jyLhX/TdW4EXHH+nomrzreWmko0yS/9N4kObD+QPeNsfqaAPnTeLV8T50Tkk3XN6au6945Mwqe
WxsQ94KS+MGWgyGCd+WFBu22593OaR9jG+7M0pcazbhKSP+HIaI3mT8sVZnP0YytVm05/2cqse6f
15efHfmk5qz1TV8I5lpIbXHvER+Hd4eFjm5rTho7OYdO5q6079spdbxfdShVV46OsrfhpWjMQtTR
A6Uwh/ZFeGrl6A1nJ5ozrBZyBI7NT4/96kkCtXDvvCv6jImN+i8HEaivMg0UASSRM1SqGiuwI97M
hJVI+TQ/OxZ3AT5qFXt7bI7iyENdZcMy0coRQKi0lkYH5lNdGpuQocr7bsWzB57h2kDdccsz0Iiv
vulhx4s78PUNqnvLA5Z/wRpLlCyrcffTk5fBoo1ETKF/WH5RYUq+scVRfVQwnpUph/dUBqI3ROfv
UqHfOsJABG2YzNrp2Ydu1GFR8jIKuAiV/InD0xlOtQn1NTIYJx+RxbgKEHcKIKvOCUs/egbuk5ar
pBfvuldHGSrrEVpv8Eg/DlzoKmoQ7IuZXCQ3rTxxrN2FWxjtiSovUwvfGuhMQJd2xJ+QO6NbFb2R
xu4TvwISVbtxGPjmqAh4OxQSLL1oZvwztbgivwIcxIFdpLGfImscHuxz82o1Dnta2yC41os1QIyb
46F4HXD7YJnXMm2wMEs9RNijuXw/2PDQ1CP8zUvSgdw/MZWA/T6WhuTROYHKGDkqiGvVbxnN7I3C
QUZD3atzxlustCswoadMEnN7oznfb9fDryEUziuu4E29NQAq6DhFvhBYWsRU1nPm+s3p1t/DDszu
82RyHCjwwXOAItmtqUlYrChGWbrnMR8TS0891ZKpL7q/hB5pt2UbmTBxqET38vy0w+iINV3ChYzt
TcUup4AqBL3qgEQyb3pTD9zS9W0AMWCxV6NXUbmIV/5FzhlSRMBLiwrU0J4mDaXGn6h+N69R0GGB
pHd/2oYPYHb/Sa6lwv6jTlvCtvUYBhHOCJvJzpSsAakIKytJgRdBMJkzoSXjek6sw5h7q/XISRNf
kbOv1+OAOo+qSJbKI4Op2WhVZfjpnbWi5Pd50KCE3puX2KB3yf84mjVQJ7j8j57UW97bKzta7wyO
SwMAy602fovoYT6Ph9xOgtEqdvTApQ7fZ9R+513vhStE+w/QNwqn7ECoUbGEae9LtY2DBr4ggJRD
pHJsClSSrngrLkG7qrrDa/iHX5DByXEJa+BLIF6YgRp2e4J9lAbBiQS59VG0DzcigfOkXMWWzvQE
Ln8FxuK+8hNojRXJNgr4OG5OOmIsiOmfUMoDfdU+JWeyqSPU76FZgoXUEhMaCrdiJWB705P51AOG
YytyTe1maetVpoORl5iinrK5655zjCdvV41Z3ijyLXVZUIRCaIdDjur6Wd/pCgQOFKBjDEf7CATY
rkEz6rIqMnbKzDy2NI8TLGYDiIgMWvVE3jUaBazxyAqecbvPbJoWjDF83fUsPAGxqfaT+fT36n8L
dngq/BBQczcvOWJeIsFjC9JR6+MkayX2XQq4olRw+zLkhgK4pD8fdyloH9V6znQ78MVX0k/1lMeo
CVcPIUChQIjbzv2hPoDIvj9VYcsVfsYr2+NU1K3UhRkvxsxuy0SC9URmRiVOjIIWryun0xa6Yurd
fuZ6BoeWIQkaETEWiegO69zAnyDcP1bzBtP8/tgGAhRQYmOmh2fJEaKL07KvnU57x5I+/WrHcA5V
IpANC/yZpZWd05Vmn+uATcTGvdIDxNNvlVCQ
`protect end_protected
