`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
UzOGIrPVWQL+hr/QS3vAGBIt4/yE1zJwjhu6mQdYCDXGYnMkOmfLXzOyZgZ026lhU2fO+dBVQru6
tkX7G+DRWCChSAZmVzX3mmG3yWWV37+pmbxY0wipKe6Lw+Ft2dVnGPnkHW+G98pvZVp7qoBP0d2l
1pp+lQfpqtCwMv+pylqpquNHPuq6pkfcprlpof+lN85Csg3ncdVAstIX6VJQHofvniL/Ahqa4PGL
RyAZJXFNdQBOEvjc/VhbLDPJoH3nGvk3wIXWsQeFUFnXctYWGU5a3vnxqaTTWnmwfgIMkR8HcQ0H
TVM1fmbkYlzsQ6jTANNEcKg1xfG1karCGZdkQg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="sKOZF8vgPvAgbaCID0L1vTI41gAo5H2/kDisjJDi1Cs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17216)
`protect data_block
ZoZXWvRhQBYQWQ9ogfDwxv7/7ARhm3VvwVWq8lOHEVED6/qMr0rqG4E6RB3gbtLoDe5+NSGx4VKi
wyAMrHe1r4LJnzEwMZM88gnoc245Wv9qeQejFuESbuEtkY+jkyxPLEBHC5tcp20O9wHNUM0RJmgD
vgFNGOqgEXnThyelWcVykcxO4wwsNvPjPx6RQrN3/KK5ibI0pQDVtCdw3b7IoM45NlWWz0lAxay5
lq0+TsggyXqIsT31HUNX5rsfVnB6elVa6AB1zsA9OuTavWsEOZ+DtbnaeP0dziYGZeOYr7YgURZN
nSWdQybeIF7lYn1wMJz9bMhupLTq18oQxgofF9p+wRlOh5aQh75yJ94pLAt/VMAvHI0jij5Qd4Qi
/GEuKvwuAUnF/cJY/XudzrzLMohkK+AXdRcjR47df+MSg01n5Rw9oxgC+uZMe3hLWaGHAA10iDKQ
EN1GQOK6T7wnlIyIB/Ta88sINouNlbtn3aneHj2pUiG4VXmPWGTOVkCJ9EACnKkiWi59/Xq9M56V
HZt+RPn97yF6rqNWWmq53+lqDZWBygn3IJPxFetrYcerdlOCraDZi7H1D79M2FTIgx5NmOB9LSD7
ESPh+Vd1mO22o4wbMhmt2b8SEo3YsScjufc6fQopRYQlLRtvcn5uCh2pxAAXbmg8M8a4ddLxRiP5
+pn4bSqyXdGae712jye2DhkEI8H54ER+VGo7e4NCWBAaZTiqbpMuQOrsYjN1x6qp0ESghZFHOLyV
j4PNuHLd2I4h3yf/GeuB2etMQ7e20yHnn0gB3NvVO9NjcwC9/A074CFhJCh1BY0SMgJTo9tV4sau
sNSsqKL1Z1MhYTiCOsCagI8IYL9DzvuPQ6NtzRbbCwkYoxd+b0VVNiOqqS3KO6sMy8JN71RgjbKI
bjHO4OCvNa5Bt7lK5IAqkEPt+RWy3hG3j0BnaIWqTX7nscYbMW17aOMsFLs7dF56fPvO3tclijMz
x1QjZQFpipovlmUP8c5U/MCrSI/5PKOqiHCzVkzR7NeW9TWb3f47bVPOf9TsGMwkvfzC3l6laq6g
N5c7j0NX6i4msWVd1PPl2iIujxJ1tFfXQ6rR/TEqFpFZtmQmg6nLdc2QdyqNdCgf1ImXJmT/XbTm
+T7qqRoTwVQJXGvlGSiuA0+xLwK64PZB+FyVQ3waeQuRBV/Hg4l4W7S44wG0mPEZj3zdoN1wkl7l
vEdvbu2m1NyhBO7PmIrubjYsvLCmWKCgvy2hfbhzF+QEztw+pbpW7E/GTqawzgMiPOkRfV6DnZDV
SiYX6VblVtetvIwtdxrnjR2cXArn4DwFGw7YoKjE1JXlUzprQBCt4yhawCIfdObqCLWjL9If6JPk
bq0rKqggctP+gIKcco8/vNb/XHAZtcktWxkVbQv8KBIvTdrV7Tz/CSIBMGLO5skdzH+0/0NSMNSr
6wXfFwD2yHAwA8fwVmdR9xIsCsGy49MI1C5ATqk7H/g3gdDi81jEvbjSiDbG4CxVwpKD6aFHBOop
JzoY09bPO+vxmdqPosaSgeVes+6l9H9tcnfNvoxY1CA2BmpV3VtDUCPMHzQP9k3OslCgtYnEQJWu
qnA828zIfU8/yrjv4Shd0olj5zA4KLltL06slCl5fz7P+Q6dWONDcU8x0vr3+7336W9ntvPa8G1z
gCOke8YL5NSGQNgq+hKrkHwRBhG87HNpK2KB3X76uispQay1GHMjXzDNj4ynvRtrh6l6VO4iBfH6
YFxByTFz/yhxKBYHW0fMvz/96yMAXNaSmuWbM9W42YHOCQsZsE4CpK3g+hQ1WxftTIn8PRcnCw0O
sBVw7e3Xh7qmvnHp+mHeRerL1b7y5YpergkSrjUtj/RXsliqCOikePihPT0plzhfpnfE0hHE0x86
KPtaMfjXvE42xTm65hwFkLXZu31oMbqdnmCDiBQusaZPsmGoXnJK1LKNIAsiHuHPDSDOPFYhyeGB
X5TyZ72JDKvhqqOoavZz92xPqkbmX6og9/xJWjc4MMP1AAS81zSA8pPK3QJK27vrLhl/jfpDpoEb
AR6rP1lequxwQ4jLHXJbE82DpLO5FeNm4VKXbz6U2rbjXL0IMBrFlqOiCjqHzG+CGIj+Iwx8znoh
ulIqnZ67zBb20U00njxE2fCVi5UyRdni57UX24sw7spvibvCRVxyhiSXLZKXhYVxKgluRKJn1QGY
Fa/fCmfZE8Y9gTdb5Dt+o/s8w9qPl4OURpsx7J3jdIWjT6Nsmmj0zmcIJzeezsGZ8P5fnC9Ej0v+
8qgcO5Sce4YqhVEB5ob4CFysrY6BKtiDbwmlXL5EJg9amq61UYHVF51jtyMH8wUKydbL5vYsVpQL
soFeXZXcgDFmukAnNdit7emzAeZ+bfk7VQXphOj7uzQpbjMcU23CMGv1t63FUVq/jAtwKdfRm1RF
KFhKp7MeizjpQhYaWDUBl26aK8trZWYu9tIfC/fvLZrxnJdPMQ26dgm/2jhXfh7vYbGD7JKA8DAM
tOi2ZZ0Q1HreYbbN7YTKLCgPBQO/bPJ4r7FWfnpZixiJ5sXMqT9JAIjUVFr1zk/H61unaFiAEU2I
tsc70CB9pREIIoBcrpsaNZukK5decqFM1apnW/fO6q7dvYEv2bYT3GhyPlES75eM2BcC4kRKlcs4
KWkFPjpfojlRscVDzZqScSEEy2N2uW93NjBWFMRrCy8xXtJYHSwDd1EMithEE0hOgT5pcxwHw/FQ
l06Bz01N8uxbo4Dl44Zov+mPUg3aWS3WmS59ic6JbezSs2VU3u2Ph4nnKq8utyXe09GnC8mvNKfh
LioPJPXK2rzS6E4ocJcEjQTB/SMlTelHspD5yY9WUBdwwqwmypByS9yDpqG0YFpeCxjC5gPmMzOm
E2IJi7qNesyUNRYeP8N6zOTdTtTzR9+fTSJmD1sr4f/teiYqzZjQgYjkR6a6ZwPeDJen1T2o+TgP
vFrKAZZtF/SDxKK5VikRWSJhGXHh3urPZMr8v6c7bdNVlDNl0KVujckQH04hG7tXIDRL6gGtKEJV
mAZqfVN82PJrvys8T9sbuZXdPM3Y31bM1bvAPL9lLa4O7Brh8gwJnswURVG9dKXTbSEhBm5mNLTw
an1mATB6jUOvCScQWj0v8iiVSLjxSCMkeTRtOlMN9uoQu43WmJTZ4goX8nLGSHhrx36RZZsXF6BB
SwrPa9MPdjC2lX21DKFc+EzJuTvdgPFhryR1PUMKMeSW4Ypws+r5xVw7CcXLkXw1xF9a07iJgVs5
M8oeyRqNGvQzcKk8O4BeP+SIwrQPpM4+sP3yBiiaMqe2mBQNpgD0MAUxep5qBy7RHfsQF7P8VFya
8Ucgd8TbrEAzLp+1UwuvmAfsLoBcgRt2sdu+dOL+OdkgxZlZVXO5mxX5xrV3LadeG+bMdYiuJv1k
ZiGTbksAKyjU1iyaTrkkQRzPi0stjFJhUq+QXmvVRE3OKTToQANTRu9Cf/uVRcRu49QWejpTErb/
MJX/pLfrdM0wf7eRFDGz49c5koSMWG8P0UO+ImqOECDJBie35bHaoIoT/adgvrpiW4VAcBlG8H6w
hFaCLfc23YN5PQPZzsjYJUEV9sGkkhQLAEKY5ZZOuaZPsgUlj2FthnUfAaLjEdnu7/gf9wziN5UQ
EciB/1zvCWnmf2uRmT0my+Ej7lYjHEmmkuOvHZhvY3FD7RAhHQ/QQIWYBQ8V7fuXeMq7ewwVr/bU
89OSuYgyjEiM6iAbqLOp7KT9GhYPyJbqe5+CGwMXr6aEDx0Vl018puCov4bEqCT6240YymzcQumw
ktFlgyVIKQZSzG75prdL9x2DlxuY7tPhvDzJjncPitKUn28xiaoeGydI0GaMasNLRwQkO+UuhdZd
VXT9IIRUUsBPTDBwAL1GGKRk7LTq0fNDAnYGiUQG4nGWpqQFa6UdOfOM1fR7lWh3KoLD63H23oPb
u6aZOkHX5tv+jTesK42bcRdCEnWpSOpbEg8RTdGq06WWDddsNBpNiQS1ZR7FUmIENA0kF8fpgiat
Fo13924lXvHhWlxuKXrWLj46dXujc8CqxeW7zrtSmoP3+VAKfupcS+AlDrDDnvUpZkxt+evDDcef
rcV4Lzf2KzS3dmKx4olw4LdNRpE/Vog0v6FUkitLNSVsBFD3BYaWlRNsSSSAgni4jgVigv2z9xS3
Zu41t63EPE3WdnA5m2wcGCHyltrZjGcPotdm2+j1pv0ff2goSZM7YH6CajDOVlD5CjnWzeVsWa75
F5RO/hfuhoeteqMY5YEfb7fuIBqSktMx0eyNB7vZvULqVcNYxuRP6DLEKD47WEoBsJaPnkmSaSAY
ryCvXdSh5AUgBkzKf2WY44v2dQiICfHVbGuwt/RcbIsfW4d9kzVaWnMx7DbOk7yAPWYO4cilo17s
TEVa91K8lCdZhiABI906ViytGohOFe0KU4mrsi5KaVJ/pJTBAVMJleFp+crmd6aNqZqGqxINd+wt
dp5JgTBPJCoXxmn2m3tw+CdDvIx9AbLOIle8rtaCnteCFo59y/C18db1T3Gi0t7TqgbFhAZ0W9a/
kqHJ80JtVEywri7teWYtgbfmV04Ltt7TYARjFnx4PwFv8cU8NpfbrTBCKtb8mSrwY/LXXJ77obbh
Hj/tHjN3Xa2bHY4Ysd2rJEOnZLxdbKHfEhO3QyWpuNucMFDIcXXO2Gf6Pt8PK/lvdqga13opm/Mn
V4jeTWsWoxjSf6Z0BSU09KrM/8pvNS8h9KJohMa1907swqlusrXhtjKR+q3K3EglmQOAfhNLqPwe
B0Bu/OdWqBGZpYCu3cWZhiZFjROqt3AdE5sqWhfnqa1gOIQMNkO9yfE/9i+JnuZhxEqhIZDcChXA
px+jnlfejPLn6OdUtAQZqupuM1UrK+qqNmVOM/kGuohWxkrwT12i+P6dbHDI33nyVOpOzSwXNaMm
WXIFGkp+puigY/YNFU7Ro8VuArHv3EpUmGW8Y0YIG8JaZtLCfXMgbrDBEUmAMMlf38xDx0AOLavT
HNjLNw8d2EPI3AU6IWMZiywr+7XRs8UtyLcXOL7n4+bo4nlzzK4HxHoQxa8+TvpFZWr28uQnB4Hj
z3g9errvHk4GT0+9psQPFBTntbVN5RFwvnwnMpD7PewnxLjmKFx0bDvpqRcC69KTdseI/jTlvGQf
lnYfHugKyNFjlUm8LeJ0nSEH2lEGnFC5DH6BUuEFcYkg+OEj/C7xF/YoEo/e4vwjvw7Dx7ThppBH
CPNP/BHk0M6+CSmEgk8OhKcxa2A/oRa2H/cVA4RoE77LJ0/qZS+V/oIhY4bzfgy/BNpq4wwQ9mff
BCNu7gZYMdMPW4r7UM9BTZT5FT7z1BxvQ67LDtsUG0njIziU+w36apav7Xt836F73UhiR5GtFm4c
t8giVQlNEfNp0g3urPE5orwSH3kzEasvRGyChF19QTnPV+6cfHcPJCcrst0eTBv+SV1fuSwL9qQy
YYOJjB5g9B7r3rGe9oTJ30lMFJhulCvHrZSZDERYV+qCMmcLbOa+5CJWrmqz/MVSL2Y1mei4myCA
F95AqLCHBBhJEVzmlORMNdcoRj6/LuYfJNdLtLKrwo71XRjnqcocVxKPq8b3zp6Y+ZdBT5GgjZHb
bxvnYNAOVJCE/JxVPPrfD9dTmWZN15MLYqYQFw8lU/3Ta95VOGKi0WMdFXGMGB52x0P6/5B+Kko9
4HqIXXsNLwx1VYRk25/0v+wrEBQDSvTv5ncxAKY2d8bsxCOKapxnvsHfcrRTzPJ8d6AbGLPu6ZpU
d9ieW1YhoNoFsil0CSfrbl5caBpoRabD7SWhTXMFFt+Ct+5Re72S5Y8Tx/gOs5zWKQU8K1OAEcKk
BOzhaUJRcn8H8ZRCbBqp/dC/kIj8sBt5YcIwXKm1vp+5+aKuiSDUMM9cee54FGkDR+Z+t6fQI0Wm
avxte7WWI0WujVbp0SSOcWEobGWQ+GWzGqV8urFln7l3RB3K+e3WK8VKcnxXjglrwSCAFQLN/1NB
IRw7cVErDXtgz58HyQNvx8G6i+9Jpr4vzDxmMPxYr57gGs+oL3L4wZuQmWNqq10hV7/kw8xgdgER
DJAhIgrHgC3yzHsMBGp+skCtC/wfRGLorf2AMr1p3+8MJX/s/i9OqTTMFt4W6t9auIR+VUBHSt7X
9pkAX3c5D/9nEuPYjMYwo14bDKi8zqiXv2ZF/bw2W6MIPohGSL3hXRpCD8r1n2VMt0cqTnYax2se
CffiEYun7Mn9JjQIjXNB0Z/6yZOErbFOCGRnX8j/iEwZyv3tchTnY1QHOC6HQfutGtNt6/gTWBqg
jU+FY3SXyG9fSrVIUHfnyPgnJ9tbKEFCt/LKo30IaTAiWE7uWHqdgi9KHcsbape9m7J4PMt5gCoS
eGvBJPqduOwIYfNwg7wBe3/+eM//Mq9ezVaHRfOBO1OOz3s0zHeMfCXZ6TCm52NdnDgM/dliPQm0
S/x3JEtA9QRkmPD1I7tymDkHXAH0aXbWaHBLhOsFLqpqjesW7spJKLcq3ue5vI7sDpJtehFDKU+z
DvDv9+Gzj01IsweIG+TlqlOR63cPdvp1sFSZ6+PbD1cGhhij/bEGKpVpzEUsGAIL0IUxoAMlqHtc
v5G6KG9AtSBGcqZVFtsKnYowuB2irf6SaHKLuN8de+nPGqc4mDm/AROA+n1FcYgdlWLLPpYb5Her
fsXVKftntQiEwbQ01tnUfo+OHYcMkeKyfNS8bw65G5VAbbeRIoAKZaIidUz2wWZJZJNCxUy+9qFt
E5ejia+H4oELHjCNBv8XYEq40u5O/Oyj2SpnqJIEcDHKBhJpPEqYXH/wLKBeRvZNvHpTMYyjOJGq
SIjCVjblpaSeZnSwWkr7cH9sM0AKDPDKuGxBJBuei3tIYXiDM9VfYqwLHPmIBsVRVYSg+Yqegf8C
dbUoCC5hii0KzIsrOjAqylmcwzzlR0MDGBvb2VgTDHrpweA/CLsDGz88LTymCeEmXzHZEDRLMGLC
KFPjzzvdoyvl7YaELu9Yg8qzgEus5/uiUrR6UcYrGW2qVUgTAM8s2kRA8OfRktkc9T9nwCs5y6UW
LuD9DQeEjE+oJsSyF+OvUIaRK9hTca3coYPWeTnEjEouJ66UAM319zr3Vgu6JGUZXEaG37B+bm/R
q1BitOAVg1t+yQ6aznX37uo2G1R806DzmPrqnfKNKTfcv8ezPuh3t2Qj4FiC0x01tDFhs8voFxXV
BRKrYY3rFjHpqH7TNH+SFwdlxtEw+JIiIgxjCT8L+rrQChBRpmd8AcytT9NqssMWR6rxQQz5EhIp
1fSH+xCrODFSStciETGXOV+zpHxmQS/PuxoEvk39inbypciY1mHiCnbxJzZkQHx/CPmdHvp+3Zxj
oh1ZcOE49F1VU4CLXd0wFcB91/Tk9Eumldw/vhIVfZwlL1OdXCnAIL+gwLmTn3UhpCdbkEZfMFJz
keWSMwB6WqDITMJCHVXmMqlpw7+VR8++5scD3nUgk+cA20kTBa8QSJRlND9c1S6SjdZ4SZORReZB
3cSDJpVW/0XEt6tFUVjc+3jwnfl9cMnkq3RCiVA0qmALBXgl3c/j8LVCZX2sM+MWdRSDCUn+w5GG
eUko1RshvdarQk+9KIsrKQkWJGgVAiVlbU5zj53onxuPdlOC3QCclcbc/mQp2OZwcHR8/ELUgtC2
qD8UzW9bLG8PBIED2qyJbcHv7VILxHG4KZxoPsdeyvJuuxdEwqOUgkHAW+GYLCOVW+LuajU1ebPw
Yy1WtkWroY8EJzTPEEQImb4IynkNsstCphVXA/y/ZZuVu/GCzHMldI3q1w4Teu98RE9ppp9xVQ4e
FdNUeECBLwBt5kwHq5ukjMoWt5PR9Up0x2Ak7+y+9hYaQ17g3Lvx8703MJqq4JspUR4mSB1xUGay
YjGG2MH8fEx0jJ3y7xFbtNFEqP1SfEcpzJssrxKZ3MjfijtRRr0hxmBY5jCW64NGXqRhttF3H/oH
xsccnQW1+OfmDfejwvqSb7f9bJTNQIxBPWtnFHK7qVCWxVjonjLQEo+xKJuxsX6qSuGwA0C81eBE
9M/cEyl9uJbqPpSeAncX3p55bn84L9hqSQvmEOvsSGqF4SnCkVdrDY9Lx7bhckVZj4npgngFN5tx
18YlVy1TLIpNWmFBAHr34hnh4aZpQs9ItnTFlEGzXVGGssvMcbTYZqEcgWQkmyCLIfkDZEZpMdHG
ZisYrNZHFGbYHeDxTygIp7fbb9epHgMpNKvUo+v77AlHHo0fxkYtNmjsI6YaQTlBE1fZKa4UNDsU
KSltY1MP8vw/LbbdL/YEIXWUlP6vg0I24WpBdCVUUu4Qqt3A96Y1TljHfbIbgD5Xih5n/4fbFgaT
uw8QN2MBsiLBYs4vdQLV9aqQz8qZWlEEB8B/Fw0hbkoOxfdxWGiobSV6J7XCIaFfmyuiukLi+uRw
bfKoEUATz5g0w90tdmmpQoqT2O9Tz+506vr4+t8n8WlewWwu1LoBzYo2h/PTAD/XkeAfmMVNMKoz
fLtpZwPY3adAuVe0FDwK2i8hzxdC5P74eZ5M6NyaSBegYp5lQhLyzBfwiG5wQsrLS8s4LGKEhZ6+
tSRVl8dHPAX/M7hxqVYauB+QCFZA4/aQRMLYgspvTBhBj38mHGTxFk9aGnIDjPZ6NFEAsEr1gUh9
1TZUufPsnXwpJ7/CnJGfZS7DZPE7ctSOZWQ0oyTFsXlY8d9jEl66tIr4JgNxRhaXwC3Hz3cPDDUP
H+HA2Mpq85bRlG9hNk0dH2eRDHvlA+111F4aAE9iw1RM7KOk/F/5j3JMCicL9WPhoLfEtajt9sYw
2vrCupr55UNraWocVy+mbV9b3mKmQds361icQq4xw96zcNEKWXIoVdzOai1q2vu9GzonfYjmUIN1
2QaOcC+5kQdq4h28qEFKvgF+PvCKKU9QnVsZto4lPzmcRnviwycDr5DOOaeIs774iw4Y6Xcxrtug
tGB94yHG11K5f6fxgv6XF294nUilem3JcXNdRoZMxrbTJJ7pEfT4PBZfvru4y6wfKBcvn0s+0TJr
+dWsSthBeB5bj61ZmDVHJHtMBFr2nMO/YIvaAtW/WcLiuxwGpKfAUsaesw7qmnT4YCcKg/n/51Bt
x4HmIGN+wMZI1gx2JWf6/idMFasay0cu2YMYYk6AQnPE+rP3WG8bftIZqhxLxVSMt8tpuERhbqzu
GlJGbmQIEcNWkdPqVRZTbVAA16UmLusVAxhiytuUdCO/EzTHKEY6riGs0gxX8avoZkACpMWeqeVC
wNsasZbLlFZ3cFKV4W5eHw7iA5kyVrj/a3xLcemMdQEyPG/kiCF/1PP3e6ukDdWuhBltp2iOYVTc
HCoatBxi7XU6Op8g73kgaM8ifj0LgeqRGWi+c5oTOMkHQ2OWK2Lau3YXr+yuKL4/KaBaLdEAVCMw
e9DcuN/YGHDpfsHsrDxmOIPe+M4BCV4cnmx7dmnadcI8C4U8G1sCmoAs5HHSgOe7N9dDNjUjyQv+
RXx1TRMdH4SAllLBb0rE9hy0LJn7pk8oo1NfcjPjVaQm4eNRrcckej24PjdXJCkbyVC+OTuUCRFP
fmWtsrHnTlYCgxLmnrVsrlAxGXVgkD1iO3T9y/af1sa0VC97cyCpqdIVPF4CKRfvAis012rU267g
dyHwx5L+JZPAhjofvXv8KXcPjtOkR+hEQ09evzcb8w/f7ZuxQbTEa3VYdtvMPmeg3Sy7nt2wRfH9
v49eaEMaf5i3eIg0mcrNYR9LAzyxT20bVPk69TLFau2PS0umOgr/+ttl81xDPBGrlq8ZxsxOvE0v
AFPAhRY024cpKeMpktl+libgpqwbKFtSCbM9yXFvwTlKcJUAKp2QggHYwNuzryLCwCm33+4bVh86
7YhJwGW+uhQDS2ZtPlvcb/idfVFTS4Py3xEQ+RdYOeRZo/SWSxYgtkkXea22PY4956pl4m5zgiLK
xInk/37YMBqyaEu8Y694A8UtOLuupxtWXT5dZLbyoLI/bHyhiUVxqihrz3eLYCv9hkQIXtitDoKB
0xE+L4MQqFqj0NN4mUI19gZb1xaQo4e9riIN3D5dSqL6Uoh8jah7dE0fAoeTZynrKt20Pvv2mKXt
oRIjDjTCjWL2xZjyufos7TsS5c6BA5PlXTr+YpIqSReoNlCQ/efQuRy7uuaAMgCWrmHXS9mhjS0F
yZZ2u0RtbY9J6cScYM5LOhMdM4DJUB/W6JQQ3/SFsZ1VYCmgbh51ziEC+1YFWIUgeH+V9l66qvtD
gRvGCdzOctBo3If7uY1NkTuGDpyMKWknhC5/0bPbwgvocJSy8Lk9KNLlroIdqozKgS2TG7/osb6d
CsC/02IE+V3osuumW+zpzxR65y/zi0A10IKFAf9y6RAsbX/mwNhVxsKkM7sB8/E/pI6pithcCd5G
bhukgQXQ59pORcD1AgbGS0yDA4s5Gh7CbN7Ss7e+C27oG+NNTSKE+2+NSwfMBs0XITW1vIFOrgKg
oVbuYJ24x820kvgI4Da3TRnA3PGMzk/XFcATznVZPoqM4JBT/SsJgpN/qww3Bn0ByWjfvE48VET0
2HYsG8v5w1jnjE2TKqw6sbvz6sVHqKZbq92ZBAosep52mWM254Sgp8bZU77oWfaMO2K05nP+rPTG
AW+MdZrXelVkSuiUChUIg/fla6NZB/9OTMk7iPsbHzTDpp4LHYMECEs7VV6Fv9/1Nmk1L36cY0J2
mIMB6h9XiK3GRzezxzLsBuAUouvAlKzTPQcFLzjXU97CyUEA2hBA+x8WjJWsa7rxP11jqi9gAhUv
iEju5H3a/Ib9e2jRa+gjaO4CAqelnW/vjAaklaFBkFB90WmuSWGwGsqTvxZQmoEyU41vzcP5OMxC
jMWeaiL8aoG5CyHt6mBtdWufbjRxBRGHIIvmqwKkFSTPDkKtd3AEbmm52WeAKcN8LUE6IapyUQBk
cAQFjKoIhJ+3qJeB8gzw9SSoCsem44b8Mer4AUTxz6/6F+DDg6iowa+IzX8RDE4sKsnVWjWwrfGq
scgCDH3nXNUo2HIi9PRFSwdsiP9DWLQfWCrEuWPYIRphKBKwWDt5HcBz2Fx1FjA/8XKd/Oflp+MN
pheju39RgQWoEaRarpmbaUeZ9tPTrCaESvy1ATw3Wpd3/Y6vPrIW2R3SHxBSmKX3CLfs8CTNsn4p
j+CsDI4Nrad+Q0XPpRDvHnJbb8LgCQ6nrGyOaXPC9yt1cYGNmvI3tbcGHRkW2brjRqbh5Di7x9Ph
fn7UpYivWas5zOMgfKa4d4dTIfO53Il1EwPbE747utqoGtamtN3ZHMHwTkloWMcbn/SrJdRVpKKd
GzohV7SUAxyTPUI+jauY5JQw3OQzSwhiLKVLN6TDQbFOiSgxryqJRNBVbULlOjjmvS1gJiOaq5qs
iwm7YiP3mvPUJmm1yrzFcHAQ08x/ekdk1aoUoy+YgeZdGZKbdlY0LokUHkkAtj+UjRQYEoIzI+vN
16SRAzCCU8NtcUO9/KM2B1HEYc66XjG6J24B4Ks9oFntx6acqhltyqt26I+oqm09FjQA18A+zS+o
TFRSUj9OBUw8MDx9mwbce3eTThNnYxRe6nkf1oFsAKM0J0I5EJe31+MM5MpZVxoqBe0ClOU1ufby
sO05Qhppsc03EnTLheCcgo1bUnylo/6jNIVhlImBuw6xn3RINx2k8qtCzZCSUlpOQWO+ZiIfdCFa
oUCqRTtxmKMargIGxQ/cbEHH5e3HmSpaJf9Na0UoikzqrWufc3WR4A28Z+umR7XAVqjN7DaLwqL/
MQpaRi+3RihvubqM3cPyrhr6e1Bvk9iYGrpTkqMZT0dtlznW4iKFVwQ6G9EybLaIieZHu0esnBsm
YOvB1JmjHiyShnG/GqS8VmWe3kVyEdRe79aC/BHsAA//8dI3nHg7oBMqepxL0k70pA+b/CUFLc/g
8GbETAqTlompoQO/wZHs1HUY+UOmHue43DSaSMeho2iRliI8KnuJkIELPR7bBON2GSL4qtUZbcay
xIt6yAjBwdgNwkkzRT72oawaf04SEfEHmbkpKL7Gg0MmB9af+CFHRykIfodJ4j/2n3IwJus+0aGV
Q1h0wwWRTTsQcocngDqty2U5HsaybjSgBlyYFd4hjlSvNiLqZy8pgJ+W7BCtZw0IRru1iAzW5Beq
vyF2SAJSVJx274dR5j3xVeIm7elFp/K8vLXJZvDYzn2a+ze4wdczdTg1OOFO0+lo8/dcJQg19LPw
EUBBlD3wqFvhyKNl2SlwM3s89qsnY7tfB1vnv9Tl7H/PltdWRLE86vaH9uoI4X46vSI7tCRCeqIi
Fv57hzAvEuzuZEWD/gS+AmlH4ybYd4r3nufQyN4jbHGnMcLKN3cyhlglEX/pQCZQmucz8i5uH3XF
QrYQHAVHl1Phn8p4aaaj8gJZI58L/+zntr92I2/wJ5WQpZpjSRBCC30Wvi825hViKNxMz1p1q1AA
4o+EYcoFN1PrKwA8+7MV65b/4gU3rmvg86Nba/0zw/wEh7dt+Wm6EjHGAZCycFiOqUwCoMJ7H5D1
pbQZoFJZFzxrhIiyXAT3AOyDvopLybHgVyfX2ZJF5rgzhjcJAMSqSuu16Uy9/6XOnlEd2GAVPwOm
DY2fbiOUA4f/3d0ixOK1ntfXcMQafG6ak1yEaVKQv8U0NNZAJGmiZeMBJlvKztTYP/IYi+x0fto5
G8zcOpPgwP4fh5vyW3Zm1bQJqAX6+Ph4h9MwEfxrERV8/fS8EH62GhQuFBG3jiUuoMk/XBWeQprw
aNC1U0Rh+l8mT09rMQXY4dzr1/C1O+oxIjAsg6C0Z83GJ/rRmbuJpO7gMMlGiwMOemno1JU7UkUY
clgzSBuuHWwgZGKz3C7nH2rftvyejRg9C0o6bXeK7H3RY8Q19aCpfsEL0uuNyyGPzEWY9HIRXfPW
XiXPzNB5YF9xdzqWUy7F4opr8789XncJo9q2hJF2blTc41i0pGx0iblPFxQnAVPYRLUoMRgnPtCi
n3eIxBqSkylHRO0E4U7dIC6Q2KAjw0sn8w9TM1Jrf5jbBrK1tY8NNU/6qWtB6+XLHKar4GsdkYVe
90fz4slNqzSwsABt+mgwvtCD2BSjllDG+StH7sbNjiM3gUnsFURAYABeVD2nIknF7lj+5QwqeTzl
PpR+2liX0PulXUANXFdJydbH8dd6LfW57/X94niMhf+8CdPA5wr1KvaQw7eM7vn/j9ss+rG+4ghR
M4qDEeiAFkhH9GMrt1WEihxvNXQ9ctE5NlrD6frWSkudeNNoiETJoHeM3cP3/PMKtr3sKu1rPqsY
3ElUSmYAUvwxvEzOLIpZGI5ytyw9Twm0LLGoGy8Qi8Jh2T3XMrHMmbrmvD+qdgERsMfG2dXvELzQ
iVL1iqzW+a2Tkx/iv8HQh33cG9z1CfUtKeKIx+nsHieqqMXsFIwsZdJ/2FAa1/QBIFxJ/qYSvVQs
vjPdsE9sokagAx1LiqYnmSJHUJU+NZCajYIqthPgbeW1r/UruLBOoT2pyY/FFGatedNz3ud98JSF
Puj6EUfcwlLdq/Yef6h9dlLV4uaaCz+ZUwVG3bQ/PKunaBQkiYEFWvc2gjs807u8qBCs4RzDVBeq
s4bPyzC19mk03vMgzTp0DlVNa3zfgFRN8q0GgFOODm/gdNjUgf40nWyGG7m/IBH4aRO1+xkfj4Gu
PWjJTGJbegTJpXn6F+6pjsOER2x1udsydKAUlm35JpN0kZ/KBMTAaHmrnjQ/o/L/W9rX7k9s6T9V
HJTEfipJLNMylERClWeeK1EBmwDnPAdrD4QSbj1xchfanQWx3/88ak9wi/QRGnfkndQT/6mV5oXM
DcXjxmiB5yMmNNnRhUzBXDi37D5YCK5G0v48FxyA+5xWKrfsGA5V/LxhJUu6WoD9ZQa/PZdozxZU
FzcUhKA5u9zoggHixxgqqabc8slnj5E1j2NWLoCM4nq+yzqZvo9U61Vhu5D09/DPG2cE2W/dIov6
LebCu3NvvQBr6C3NMZqn3g9HSgHj6maOdgGa+A2bXQlF9s7htwI0gBA+x0kczGQsD2gJhArZhbvJ
DIUje+VzV1m+UPze1K16aY0dUQRauVkA0dZOFrRHtQL5dDpCmuI0JgMGTn1x8aXXw75t0yX3agm+
9aDSd94li0JUTMG04LC9x5o/kNE1vgKx6DpErwga/h3yFnCy7TBK4IaJEoLJDsQNR/E4dePhTFA8
sdqvrIJ0Rf42K0dqceOzlKTskEodCV2JPz596wL77U9DKR+08bT7Yvq6838Ob1lZPrl8tF+/VNOZ
ael1hBpa7ok6/udVSkEdWFFKW224hTquuqaErTDKuV9IBOdC6WrQL9U6BZd7eTAuCBuXTnjSOTmw
9pbYrUQ9cJnoZeQ2UUb7QqnJbqCgD8pUKUZn4m93kvsdZgtjdNbCpGwyBKMmCJtUGuBLDPouoyQJ
XHtuKjU25GbtgdDWt8tC4uHRlrLGq33w/2qb0K/YwpIZdqBwhHcRSm8RCxJZnjffxNP4HdwQjpAN
NH9AUWaI24v/7F5XBFJK8A2Ft+HIJSPzEwRMKja0zUkNEwCnM7J/Riak9J3Z69Ve/HrNMTgcRUHY
by4JQWSPuRHKaYXodXfsJztpyVkf/ZAtEy2k3FveMlsFxxC91uaFQW5JlJV6SE1BtjrxMAlF0O7R
QrStZ9PkugWYBmvnym9GyoIkUoUITXITNl/vWCBQADJQDLzFW6A8PebvpfNm6TAU2HypXKAHfmuL
eAuQMl2JjaBsHvDFAkvjbkCHrjSoBb2EXhK8VRDSS0gAcKrAaqezrL1setzXoRwfedOARrB8WJ5W
oaX3yVfzXAO5kx6XdqwSQdtA5v1wU4uBFHD1aUQ0XWgsI01tCBQVP+H2G9uMynhDipRdJG/mRJYy
PnMBNvomDbmvjUDhcj6uWVJgsaoWmvnl2/cD17c+oUzGk/hi4Zwo80Hy8pwYelxQGzqgRHBya8GD
dvHjW4nT+Utn7Zgwz2DJLUbPHDLl6Tdrz6QC+rtuPlvXmlS6LquBLJUkuzoXD7oSizc9t65o298C
6GaGHfmRcjMzbh/DCnCFiEgX/XzfPnTr28VNr7OubRCWiG2nz6fNVkLB9az1EZoSBoqq/zSIC7ac
9P99QVo1wWlKPrhjyhw8j1qiJBZlUEaaLzrMubEqUEGirMzY76d1zi0ru2rmeV+/4KF2E4svGKoK
8uppUc4YesG+aDq5oti6wjAIIBm8GDvA/xVXJxGD2r+t4ZjQDaQ91qCpY2U1E08v6JSTz02m2+s+
BW9/gh5ECEpNoHQhujiEp9QyPTFrKSrtXzoY9+CdBYGXiz4wJxm+l2TRACKWt8pEPZ4j6lvl4RF2
J3igWJuNvJd6Y9TzolbwEAlVcs34CbM6Ac9hoplN7jc0q/MY5zn/k/vfsAHciZK3TsAN97p1sFqr
nb7Oh7wHILirTeyoG70vDXkIGxIYkznq6gcnqJWrZFNhfCmPOGx7oJUXeAo02qs7Xs/jMLDbE8WX
ChthIYj3HXkqCDxmtDIb++a7RFH97juF7E4zje6yoQopWl/4AsMhoczStSXAKSSqIiFfdZ/9UlYq
cwbf+PtlptD5RgRYjggvBd9GwYzpYPYcky0OX8x5cK8AumUpf1O7OPe7GZihJpQ9/kpNXz/KMfan
u7d0R0bCZ0GuNmUf9+gm0we5Gc5HxfnzwEdBiWeAPHPKxLBxzHn6ZPJYWUE0O2Xr21bWi1Uv07hz
e/18Plwzqox4jgnlaNpkZHgfziQiz+b/6MpB+UDjDc9KHTrp4+p6J1Yj7p9dUBxaA+XvtFtlBPDN
c+T3/awQ/8fz56Hg/yD8J84awxH+7PUy6tra9CA4oJ+xxhXwD/d0pEK7RnUmpqhS+FgBSDpE5VtH
/WBSvy4ydn6GPqo0RyPYkGE/hu8pE7f47Dkw8m9yBMyskN/j1o3mVuXU0frsKf0HIKys6k5CeJ1G
lff2RIyiJqFLOKx1ffuEVlZTNLuoKbihr2itu/jVQB/fiflabn7lgZBYdWDjcgaMG0+6U5ZedaXQ
e7vth/ljLT+2LF5mRSi5aRITyNzUiiuJksvBI23dKM1Er9zRg0XFI9ElwxjHgtrjPo5CMP+UrQCP
m62hBq0FWtvc8bdykRUrLhEsScdzX8XAyJLOwSaFqp4sDiydpCeEmh/7FURUiZt7CpiCAKUpJ5Ol
Dv5UUle8VMYwxCCCM0+l4dmjRTjV9sAQi32Y3x2aSTxJgyDvrIcmYampBnXlS4COvPs7d/4rQoHA
9kJ9SJVSs8qn48bxod5InFUbxSlNsJ/X21zEU0NaUHkAo0Yz9B7FWt9WxBmzUsQJxpv5ZLp4mEA/
9RGN05fx0DQ2zht98PZeKbidaZJtuxX3jQ7jJSjzvStN5D2VdJrVCpQvfTKARXz9f7xMy8n0VNHI
AVNbRwcX48ICrnSOXsyCIvjZZQCCcBLhjfWXfG3UDNGn35ZqUB0La0pk+V4mVJObHkp4Ejo5fCLn
11BAg+X/eLsRwbaAs0aTPPpyq70O+Nnied7q53unAhqtIJGbRlqxkvtJtDE3iE8wEawVECZYa5R8
xgBMRf0HbGZTe8t44oviLEiYRZ3jQDvdlUz3YMmSNKJWePH5dk2+pUBHEE5fYOM+dLbP8dKrr4FA
+5Wd+CUles70PRANDOYTH/hgF0EdjgVecHswcqDW4/4GBr8g37RSpETtXl7RX/rGJMX9v4NXF4Jx
ZdcB34F4waFpTZF3tRtb6PC5MULYtB4356KTXrtve/j+Q3Grk0whyEuieve5JrWOxRlbdwJmM0x1
8jdzhhL2JNjstlew7pAP9PCBouD4iFqG4W6b95PIVyecsapJ6eLCYganmbBFqtfPV0AN+wIFILwX
JbdHBqumGAeqkvSMvUrC5jX05QzTvNj402IkZMxdIRITJ5AFAGyBBX8Zz/3Z6Af8TzAvtmHj/kkl
MDmlJYRA1F3j55iZSFuiPCLE/2WIHWO+n7aSKd9IH2V9P8NHOCZHaUVqF/yq0nzNS3/Q6ldCIG6a
CLkSSjwPFgMHsN0zPAS+jV/ww9Qi3rHt7UMyYgoYtblp4CqWF/C9tXCDqu2OS3Sgpu6cc6++qWtB
L2yOz8YMmt23kPeyspU6hrFu8Uo7gh/BW08Yj5iAcZxE9w2lPXdZNDqAPTAFlN2MCJ19jQkg1d+Z
T5cCEWgKDCjljMoFJoDGKeq7xQ5XrfUEPOdYs/6P4quRkdcmR+cyX//R7HXDUO0gJXzEZrR/5NsF
v7hjHb9VaPsMB+HQNxnpBCoVTc4BerRY+sc6uGYurZa5/yODzc7aE98EJZ2oihXodLwNWd7LTjP6
C7OvPE7TPeM8BZBYBZAJGsnU/xAdFGtGixFQpM92Zg0LOm2Bc8Do4x1IQlp2jzWS61vM5SEd8QCr
b+ekVwd5fF0sDnn2T+mNeY4tE3fR+AoKg9nafK3OIThyaDRpK3MiJWlIHt6bKr3XBQzCLMuNVqKE
liJ4g1w6e057FV39QPdueN2G1xOpqksnj6entMHx0Q16qKLD30HeXBYg2/DIXVtGVm+3TCS6YtE+
mwVL3LzcFOyOJEqdmP25lGK/pkZ6UU3TOvpFU51itVK87czc35YFCg1NoIvjz/thshZh4f22XNlM
0VD6FNCFzwmrCE7UBB0bF8GVJByewE9xP1+Vq4eAlQXUqaAyCN49RPtAFq2MCczXj66DJT0SbKvv
uZU6C3m43Vv/6eJ/m96tfYUeHO1zWhmmxG5tJHHZbIl7UTbNNq5+Gy8NO5MIBA7uyIAgntEpjd7O
X/mfmdU0AnwOxSoHPL4c62UL1x0ISJN0hL7ocAVrJ2Pvpa9HBDNda0TwBn0QOjmnyi1KdqDplQHI
n8T1J9DCPI9qpCu2ckXdqOI/tEOGdxR0v34qweeN+bb8MgY5UnhKQTZVggLCePOoxnKMge99zSRG
7JcTdXcUvsf5cl+5+/cBpZSXUNBSz0jL85su2fT16DgC2z4hkeZnubLy8JNIwrvCVbTb4BY6A2/T
qDBlrMFhegMEQlaoDq00RB+0STrrD3IbYO1zHjh6xzuLXoVHVGj8FHkMwQ03ctszet7gDJBdFtOd
3U8AR4b2DeZkWJ7QNbKp2jltYPsxtGvaMTE9uOeMyjTrH1+8N/bcqcDvVL4WnE7fgSP0+bU3LqDs
1zpM+koPmbPodhti3nhUk7hipJLOs23eU0GIdojcIrMuayE0ZFgAFrXzp6kdPccrhWug1+22I9ST
SaZsu7Aqhhlm8YJ1w4bodSfD4fQumbVT4h7W719x9PQGIfogBpnEIOuXow3v4XcpKikAyb0CzG9L
VE2mDIO4EQZW2DY/eQs9y2k7YDq3NTEN/QmZIaf/3Xvn2a0GT13I4esYB3TwbUum2z1RXuKkvrma
05XNLFJZGjVb7SjQLBYKzDY0Er6s0yXJt7J9wJGIryeeaFB0CSjzyPeDE8/jhj96nvV6S8PVxHcH
3GFjhH3HvTaPmT0j/iRwvQOvSCnYG+YOtuFLZuoORvqWFqMwPh/C4Z8f2fDoLZJvHH4IzQeEdHK8
3em/8oDGvSJIaO4nINAzm5O6M48Hl5o8OPKl0nAeJZYJZHVGj2NIO9Z7WxvNATyQvmjuEvbk/eIu
1H4MU63UNoY52h8FQ7Nn9gBnn+nH0KINO3W4rbr13abDvJMHfG/7zOgRnXorgFAWd7tE6n80ZLuW
SdRqOW4TuQ+LXKzFiKAtIaaEywgKxZPM3D4y/sejmjaj/6FTfbIQWfGi97rS5nO+fg0jVlLsH8qu
E0tXnB9W/PgMnkA5RTfQSTkTaUOiSk7sT+zGiQxTkNI2gi72mmdt/aPDs5+iw5GmxQSHXXA2OHaY
AA1D/uuIt+gV51JuN660Sag8D9FaiRwzzvAaON+JxGgW8kfBMuRJEfqKUmOgRug7MFUOlgn2Yzcm
YjtP93vagUyCTfB77BxaAc/Z8AI8dE+gAnPOzPhkX087KowZWEJOWXffWzrrXXN8YUOO7mHsgxNS
shFtvmMyDCSVpoW+0tEZ7Z2sMZv73q8ZSR2rru3foqpamNVIZ2OJ7pk+XgyZlgQyas+KlTsecePX
AY4NdhulTeZTedVWHUReKoOvu8XaXa02HtUGsLd48bIWsPw/Qady1B/6XYS8aQtPCB0plgX60Xp/
4NLTdSrXgZsCWHAVhzqqGvZu/XBfTMZNkmmzISX/nrv0JE5AsZQJPqxQpJAsH3ZsMh8T8cq4BnkQ
4/HzwZ6Wt6IaBxLvUlcyoTBSmuX47SiV0hN2ER7ulxCi2dFocybIanpU5GhtYAtF7H2AauNZAiX/
ZHliBz3eUpfCq0KK0x9oMQTULqSyUQVw0PrrYJorCutxwaUzWvDtkHENdIvjEiv20u589C/bvCnA
0LHlY5R5/uR8TzL0sa6O0PIT1//U0S6xpiptItsYq1mn6DBU1hb0O3ADlow6+Nrzbnn8/fPpCqbj
EdIBlwVPljBS6A23dbZTRQATd09RfRHl0z2oQ5HjUywYwqm6lllnyiOY6vSlWaOnrK8WmVFRubT/
z2lrnBn2Czya2878sg4c3d+GUJThTNYsOAynUMl8GhgCEkw6TRLWGrT34SHeTXgQvE9HhFA+M0Ht
hABjM9/47q8ULca+louwa/dLDGxJ6LiYZM0hvdhWE3OBxUdp661zkzoRMJfXtQ/TUDzA1OygAnFe
3iRMIDGgIvG9IDxL8Y2fyS0OKeXYvwt+LhVqWHT+W6SLw/sJbRzJuZmw1zodfB3ohX7MeykMK5zK
8e9PmkipncG2pDnlS1oy8NHvYMoWYaIOfs7wseALNyhHdSrGXWWQbCVLSP3gFC+JUTufML9sUrJT
rMN8yRKdqiv1klO47w6+4UhBXhJQblyODIarmI/WXNF4Yr25CkA+GlY7mPzVHyIwOsqjI+WdSxoE
85fR8G0LNv/hw2vJ2twj9Po2Cm359/o9wm1kDjKcweH92mxM0qNBc3fAP31gSwyL0zzg5qwqAlzt
omd8A+8NTH9nHY3eV6H8prZ7bam+OYaaOBMLMPFs+t/uDGdaEDocuXzaJcgPtBeje/VOPpnchWc/
2G/E6Kbne+kisSrDH0/LDCuMfMo2k/d+iQxvaHiEk7d0WTFS93gpyPDr7LHoGXUl++1i2D5hZzvE
BMKlEK2C9DM8bXECBqeBtVcTWHi74RlJDusXHduwAQIPP8V0OBReWd2w3oL+nEDm8u24Z2PnAHoz
zmt5nXTtt6tR/i71jxCjXRArYh4o8QcExUw6vES1F7hC3DjrJU7BT4Zgna3HpyqYbf5wpGCWv1Jr
ZE0aBwfAf3rIlWTxGn+GhLtS2d6u2h6SJMT1GgO2OYFPQyhC3xvCYaL4eVOxn1p1AsyxEB884jWr
O1ZxIKT4LgbCTBMPw0SA3I9/LioGSq4tnL4+8Pmbdl4Imvf8TzVdnCwHauJhCXX1WJlIKx2mdKPC
sRgcVXioLQbG9fGN6VjDeoypr4etatRBuuTCtMYpHLb+Jx9ak7Mr3627XBFrp4PPM5t0thzMA75z
+ThQ4Maa02od8a25Yr0bUdpEHovpEc6Mu3OmBHhtaO6VEl6muk36M1EJ8eDnd0DrCDoA8wNEBkrY
jJ47W7TKSmT/OB+Pv0RQk07Sxb6eRfBAVu4k77V9g8ErnL4hYXRQvkoJnenf6JNdYQKhhOyXRQzQ
xRrKXt64YAckX3heS2h57pieLmivFErk2pE2aRJu4DSWoEFtbcmQx8/ADszfHU5154t/A8KsfZke
IXf1RRNemxEfDktLD6tqTUPEhcBLGljTRUNtTSyRrByKWsYn8LUGYANQvBnPwn1aYBuRfYk6ZlPZ
k5DaXxIZU24y4qwIiZwnpEEjYhunHQOdDTaCrrCeGvEp5DczyCJb8bhSAi+Lz0wSBOWk1gWFZZtx
j9ttGqYhjC1LWe91D9HB0FJB4A+CPc57k/zbLqMfaz9jIMskP29fEAXrUUUIWs7ShkOGpnyAF5Ph
/WFysaWf++YXhxdZgzN7zKJReK2Ntm3FumaDBPfaLPAZa3fWHIfnE4StDRQcY3Zq+kveBzp8bsjg
X+LiQElA08PNVgfSG0dZHAeO2AJLbmsa5kpcu/Td/BAB9+PcywqGo+hlCWkCjTZnlWYo4iCAiIIL
I86K6eK+qSTtNJs6TvWW+rLw9o/GkHk4w7b8n/nHTil/NtYl8PLtJbhEqCX6nC7wPx314PO5TLvr
YabwnC1cb5ceHaveRYZu/2Ls59ZAvBLYCVg/oINx6pWZC+oLV3BMrZoHVduMbII0OCEx4aOI9svj
1xfX3nVu4B1Ag4o4/muI5JB1smTjkhAQ5ZzVWCbGco2dsGbevNjOyo2qiUiYuxG/MhNaNq62oWEt
hTD/oMtWlRNNXeHJd/8D5lPCbnvkFqAM+diJKU8sbcpZ02yVVkTRmalUrKwQbTisprf3aaYp2nIz
4AYYPu4tGzlpaOLq6xCnITDMFoGeVKKn8RHpi/n6GeCiunB8WPMtLXYq2PkpVrFVPVAig04m9Tl1
ncmZ0PQajoR6yiaG5PtTBSCSKKnfSW2hbcPysozOh8/kIpGklqsTIYP5DkeY7JZBQj2U3Rj+v6f1
JITiumR0PIoCJ5YJnvaPvzFt44ezBSf/Dv2MAIZWpxcRVmi7XxTlohbMDr/gse5JCU8tzCEVl0Ye
cBufs2sm4s83Q2lCZWuxU72Ut5ajQZfp5qYSt+QOjBPAbbAseym1V7Kwish6ppLRvxOkvdpTwuhF
VNbDqCx+WRG0PxTZgpDEjiOs/HLH3QHHsQ1np04NZYZXGrW3xGBA9BXGe/Z1JcMxNDOIsYbweO1u
h3ud/L0HR6p9gAxtDQ2EAYntHmL2KkcFEeARu6qf4fsLY4z4SBhZcgiNyhAGOPs/Qyb2MU14sIVS
qGoHm8dFKxQZMQJMt3ERRl98gFbG6iNfuDUaKYfnvyiQisF422C91tMcJPP/18gzHcDXmrB1hmgI
+vocf19p0O/IjB/2SsDhCWPrTlt91p4N56/u2XyRd4eTS2BbXcaOtpJmYLRz3ZwHpdrrFxPi8tQY
A9uqVCm2leUBuNHKH8MR+MORSAbvK7wxDSpXIss2gJpViVSIVZlajNVxAwrNBpoKOOIbI/0HDMlF
LEQ/IJgj2fLAwDUyg0xxm+lwMn3K3k3lKtrst8rp4a2a+vV/7RbI6Q85zedcR/Hk5w2YpLJdrut0
FJ97fpXAaMlq07XIy41gbvWkAajibrSdu7NPffYlIxeBwwOxOOmD4GqxYA2Urk7Dv1uJJ/Q5dsMR
3otHqC24LMYDOQodokAOZfi1b1NhDwrm6OU7ik5outdsF79byJykxMTgpr9+UsCoWr+PQ6Z0BdpR
PWTt+RcgEKM0BfxL9+0SYSnuUnWZ2zkahV+znSgXw/ZTm7UcOG65/nw9irYNUuW7Il5PbuNVQ4Tw
vCuzAP8zjGt1+/+uM9QfDR1yqRZbCJvxlKAnFyKjnvtf770VzSo4fStOdhi0lyz+JT51pKdRU98m
j4mUSNCRUi4KncIZg5YJasPfqCFqaOM79wudjp8RrphPeXBrvCUS/QbrxFuc2UirogEGZBRcQrKz
d/UQ1vFuCbsWfcCPErZvKDk8cBcukrg45idtp2t8JJdeqecxc/nuqYdP/lfcF4InFXcvZ/0VIDRP
DRyJ92yDs6rnDeeKJfcM3dltwoXKJ9uF34FEs0UiVHqADJqbo71MTkdyKlREoGE2nPQICrrLHvMy
Tc6yJ18kp/oYo9E1Lse8K9SZ34krmrVjWg8azxGKLUmdEC8XpNBTrEb/jq6To6RwvxYjemASkqKK
2aKODw5YQDBOxaM4/2THmyMYoCDF8elIc8yHGtxmBt/pWzB+loUMsaWMmY3BuxBlyOtpy40ycNq+
NdO3B2gw9HKqvQ9DsXP8pSaLhSR8PYMiiiQhHo2KkZaH3BRN7eSw7br7HlPVUMfxYOwz2cxClfUn
yOA=
`protect end_protected
