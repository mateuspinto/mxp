XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��׷м�]�`�K�Y@�S95R���3W�8�z�QŨ��z���ȡB&��_X8��C�rݮwT�.l�m��>?��}�6�'1��1�P��"���R���g�C*���-��{���+�9������I�k���_�(��s�ԔS�n_d��|]��9�����ABz�t������sA��u	���%�3X��Î�-��p����������(� ���h3.;4�h�c��L��p��oh.�YI�z.d�J�_U�?i�j.P܊x3V�(���3t��OJb���0|�s������1�?<]��=tz	&��|�,h"!��3���{�Gl��b����5�fDF:q�������e�B�$�rA#�%���jv���,�0@@���>
�"�����_��̹��[�]X9�N�]6���֚ɦiV�-��
݃u�<���k%���.r���@���Ã��&"Ɣd١KZ=��H*���f�)��x=�%��ڹ���^���P�vT�v;�Β
�\1 �=׬��+�p��qh*�.��������Z"A��t��\_r����K�@�H�	�L����d�6f�!�ֱ�}�]�M��r_G8��,JE�� �wbH�tU4�}g��r�S��^$�=�c�Ԙ���*���J!�Z�C/h��I�l-���6_>�a7�K�AVu4�Md�pp�4��G�;C�ԋ��نU�}�l~��R��<e=9���f�V��V�(�.�W9��\G�(3lXlxVHYEB     400     180�*BĦ�;�܁�D�M���81���7/������z�I���Q����ZeȮsuš���s>j~1x�)ݚ��ޜ��LfQ�e×�{u:�t6�!:Q&t�&�Eȭ�0Q[v��QHi���R)�g7+�����)�J��Y���P0�6:��'�p�A,�u ��~c�^�p��V������S[�dj�yc)����TH�D혱��XN�H�	�ó�"�-{�P�%u���}^�7z���X��V^Ǣ�5��BVf��Sҗɋ�
ǃ5�t�*�>qEV=��,.��G�)���"�ŇV��2(�e�����h3���~Y�lwvS�$�o�iY��6���s���
'Nƌ��OWץ<����Z)��4��w����-���XlxVHYEB     400     180rk��C] M�O9^~�W���p_��^7e�ٕ��&�\����L �����0Զp���a=o$�����K8�ka���`u�% �&��nOS���?�&D�����F�p�瑠��
��E�:��9��pƈ�oR>Y�E��0|�,�zke�Fe��/=�yC�#mj�R���rF��4ѤM4��2�$x���g�R�%Rc/�g����Km�{�Z>%���'�F>����mAx�	T?��ǵ�K6��JW��y�o�6�k�h��W�I�D�5�A���b��f�}��I.CTc?)��:4�q�#�=��&M�=��gWt�خ޿w^��;A�_�����*��$^Դ�bұã�n�e	��,[U�J�:`�L��G[���XlxVHYEB     400     170�h��9Ӑ ��E��Xg@�ӆ6��,3��@f�в�kSY�wGEz�h�u�D���d�yK\ɨ~kRW�-R�DJ�� /6�"�jgӈ������х�A*~%��"Uc��t�K1�Y�D"-Yc��G>A��]���1�V�,=D�X���3���n������l�a�"�~�B���פ��h��I��^���q~�����Xn�s3t�[�~]��ᘞF�kHm�N�8}��u)Z�p�9�Ab�;�O�G
�I|�� ���=�G��2}�o^j]!K 2xh�>�1P�c�׬��ش�����id9A?9+�r�QG���TN߃�-Wm/�-S���	L.w9i�g��Mr������[XlxVHYEB     2e8     120��N��ǈ�&SU��� 5;2���Q8w`@�*� ��@� �*���(�<6��"�Ӌa�
�n�JK�8�E���Ωꑦ���@�F�=e@㌬ێ9��FV�B�{DdZ$�����e��J_�W��k�_#����.Ug� f��z�e���,Ug��bև�󥈱�ӰYy_ӑ��[�U�[Z7D�N�ٿ����`��>߀�ͤн�v��a�'��ɺ`�'z "k�`�͆����`V&�iE��V*< ̈́��(��
�����U�����Xz�8�