XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~T�g�1�Kq/o��Av�+�ʅd��\0|��)��o3@.��"��VC��e{G�%5�r���Y)�E�+Q$Y��n���i����YrQ�,���o?V|�/�Q���0t��w�v��)�7i6�x�S\v�o{��ñx��K�&g���^����(n� �j�ml,���'Ǵ� ^"�ܘ�<9��>N����S�e����xS��{K�$j�B��@_D����HT|�x�����S�H�G�$/��j�gsd�}�'�<����/{��.h��O(����
��7��e���O7OӠgF�l�����l��"x:Jv���f��n)�!G�9�˥f�|QS^��+�fdm�]E�NCT�>��q�Xڋ	�"_#��ր��͙�È�h���(T9�U�Oǀ��f��w�AK�y�u֟�����9�O+�����^�_~�|0�ŷ���)�����o�&�T�H�E�_����%��vaqM���e$#|��^{x+�&�q��f^��T�BUk��,R�j5<U����Gc��P;i�5�|�?�K�ZZ y����	$E����K�1[p���(-F������}�-&�Us����N��6�ҝ�(<b>��%�P�^�{�1�9N���Q� #a�ϳoTU3?��v&@'�h�ޯ�A4�Q�iD�5�Ɵ[�[?ֺ���X��(�3T��7gZ�)8�h��75���W� ����@r5Læ���h�Ft�'2����M��ԡ^��)XlxVHYEB     389     180��.��)�����[ȡwk�xV��h��:�Qb� .�Rh����
�`�1?n��
��wx��^i�?FK��q@,/E(��&��+��
���	ER�<*t��������Y�b������M �f�f���#Y"�7�K��:�zP��C}J�oo���6*�k�3Ksݍ3���YQ�(��L������C9HU
;� G����=&
���;у�K���o'MO"^"�X�%�x�v�TD�X�TB��|g�a��L[꿨;��s6`�:l��ERֹ2�C��f!�������D�[8�f����K�z���lN�;Rrt�ż��}�`����M��.�n��gt�eWVЩ'`�蘊Od�)W<�2��_�-�%
��