`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
n4VkW17rK/wr2HiHvLVWqy16Ywtzkta4E6cBhv2NP1rfnsNhoPNRVyrwxRRz0ZvKoO8lNxPeMMed
EjQyMFYNtFP646fnWxl20lGf+d2aXpAKHltT/47Ad9VxaEOCxc/CDoRuOqKyZdBlFbxNwSTsDoJT
n3gM5KTAUlgDuE0mwtRhvI9P7/E7XgM5Cl+YFXIkedamjl70RY6D9qjpV3NfV1nuOvPUttYQHwG/
xdWu8oHvzYXda+PWvrEt2fNgJR6j9cBdTimXBOt2G9DYVXVIUJQMR2CFdI/h6b4lhIzTfdYz3XpK
81lZHAGMuTj0qLcvzuDIah58RCbKmoXIh2phvg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="iqkkHuCJ5LRM45QeftQOrDXGmpUA4oGUia5QoJRab+M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48352)
`protect data_block
KNgUx0zYfZrpSFuWvKHDiY8VGUTjRQ124IZUjjiJQ8Cc00udml6CmSFy0EFeefihfutLK1IABKQS
5WGwytFL8XfhhmBd0ZHpu6RJjAgTfz0SFxaYMIaLLAeDsc7dbBuoO+48gPJ+JQ+OkNVLE0CAQML7
87vf5HkF+r4OLVARoB8eXLAcmqi+DTLKDlx7qIFwCfN8fwgHOIOB88mG9Sr5HlT42Y8cE93RwhFY
kX0SfbxGQ0JWnjpqgHHha4boLJcFx6cdyyv5FiGw2+t5WxUD94d11MgMQnWHFnVpNgppNoJxBVWx
0DbR6skrBMZbcBsFYn3XkdIgj9Zzu93XsIaT2kfLXY3hO49YAJ1+HM69ur7bAdMT34N2aa0RqQ75
yzZWY126C0eydN5r6YVwau6d5ZKX9YAHyQ3D7PBeDC5vZtAE6WjmqJbYgOk1XC3jyYgaGSxisMdn
1lpgfQhJEpgo9F8wayTfKMv2Yjf/psYYHj8yN8Nf6fZH2ESJ+jHp0YrUQFeuaiebVOZzSmZo3wAH
mU/LaGfC4HUwXPNE9nZo+ck+ezEMt/bjeVS4/Mg//+hepJDGeWvmDPC1WT1vuukGjqZRBpQ2vx0l
RUHK1TME/RowToXn5nYhZ/hk1L/G+DsU50ee4Hsz6Pesb4upqUeSTgtJ2pJM/u/Zc8ERQahrVBNp
6h40svMh088VaoWiIvOJPcfcQA9pUZcSb0Y8hJD+d1WABNP4Inj8kZ43mRxxmAAceUM0ffvE2gF2
Cc4iJmVwldESdyZURM0t+V1Lziw0dd1WHcblnbXJC5Y9Eu5eBNHHjVGNuj7UGQ9UfWWI8n2381yL
IbNPSIszsuhx9nf++POnXVL+SpwLwaQeyIiZMaUFZJ6j1BjkJWuRwEBa+Fj3PJm7pd6YU3PtRclq
Le0l+tYkJXYXsTaon8Ga/rBukof6O7ZlRFfozIX4fKOw5AGO0ot6zP161jJSHg3spZWGJixnqmoI
6pBbWO76zVMLJSjEdcDdym0+RgpTkXKnPOG5rVZDXk38a6Uw962SPQmjZhA5wSJW3dpZIjGuZdrc
1BWNOPOutjb5Y4OHmRnVhSByTLCTGOHF7hoNA0bnPwEesrpuevHsOy8c0uUPCTTw7zChtVy+De6Z
K2yfcvRuiu8NakAs1sR4Pe1laW0pLp4Iu3MP3t0v6ThpW1UIkWnkQB55uG5qDgxIaiEAj39G90Bs
OpnPZkcP8YE2OfaF0swu33fRlB1XhQS1fcldRGIIs/CH9Prq/HpD40i+Ti7Wmywm7X/05KGpbjGv
83JtMn54UFlGB2UfxYbB4Ljrtxucmn3YVwVtJUj+mVjz/bZUKdzPLMEH5+Yq9lnwRsVtZE6wo0/3
1ttiBbsALAcEWt2jN0CQiNudCHFggVWyjmPxKOpMKspZz95RG8fsyLM2dUa5l59LfVV/KaYyTaoP
iEXVybZ29IdeIaroaL62ETHpEH6VNpg/0QiTY8n2fgDdGsR4g3CbbNs6pCDc02LEbRWkRQBJ04nQ
YdIMRlaofPUs3CmVkHEUHTTit4YI5tvwV1fX0qJnrVSVIMimYRxzhtcKkvBiNeQw41tPdE8HvxlE
c19C7bVyLWMeU6jPmdAntVKLmeNOGd729xqJqf7ZTP2jyv0BCDXTRQiWH07FiIzx5OV9/h1ZCSz/
WDU+7OaL9coI8XJvFvuyQ294MNYcZrywPZxWeKM9Iqs3vmsmZEiao7AeCBFrDdeeP6PF8s2+rYR5
RDlboF2ZHrLq1BmDW81IVpSMjkkgyY5v+4VLTFqmPVwlxc1o9mXgtxtlUXY9dK0vquRGAOWHJJ7o
8dbOK8huYXRSgLZao+Ji5DKzG90h/6LocrDGQmcGWd+/yF5clHIgiWkNh0HQLfc5ejGgPRf4TV0U
t1nQ+epUmMCTaOxvkFogD9ijSwPVGXhfTX5w1IZthofdPJp9I1PpxWkw4sIffTyIWHHIbQakJW+v
lE+0aw7gyY+ClUzMzUZjucOBJhLHh57LpSHCVxlwfoXEPjW9dOVw/mJVS5NBkdzmAILH8+Ekd5QO
okeRjmCtgQtWYSWvofPvhzE7RMRGq7gtzACJBs0mBsNrFDV6R5SIjvCl2eTNkaccMH5jy/7tbj2z
IJz03ulVwZpsS0s4VRQZMUbkeyF7xFrtOaI5vOjq9hIiooROV0n8ATQ3BPG02fr5jLcTlwpwX8Vy
SreGlv2krgpjVGfpJyqMO3qfdLWP8nlENRxG+Z3kU6yhtzjKCz4c1AuuFbhooyK0M/z3h/llhyvO
4dY7hWowvdi/oWMlgwExOQh1joSfHEaxjUVdvghA51SgkI1laKltETDtotWv3jp2WFwFT32aHBsJ
7WGyN1KUyM3QsAm+cbnHXNKgm+a65BAU12XrWSMcO8nR4YYeC5b7/8YzevuwYc4FU8BzxExktWeG
SPEFuyqWBnxAfwxzb9wzWxhU0+iyABVbDXqCfRLd7u/kh9w65kb033OozuwCkxzgjMdGhDzGhMz5
jJ4ioiMTel4QxlQ1gSc3+16cDWvJoNOZ7Lu95YgTYHZ4HYZudgtDX8aiLBbkB20lpA+pciTDGTMR
xLzj7n7CjbAYa92CNaxaCJvX1B6H9y6P/Clht8clV+Xdp8yu/Ear7wqOxk/qqCoX3xEfk2f4bkuJ
Qc1cQ3uTgfKupYZGyiKnTzbV1obUWLS99IJRIlcBF2uVa9gpM11UdyIR1+N4JfZIOClSsAzjIXcJ
aEs6DPiUXtsKcbXXzv9gXRuUYYosUCGB2Udghlka56greR66whtEAOd55lRAyZCU05/Zi8+D7/j2
8jsIE0xRCceRde60ipeCGtoPRpD2hZa4JCYM6qfQwO1gaEAOLhrJze9rL24mf3wH8mrrs5l4X+2j
vFQuczpZZLKMnQ5AGmPgsXjNxTr/mc/iqrnKlOv/n43/SoYapbVfP+2eMd/Kqyr15kC2oN9wOwpY
/1mIbmo0V9mcpyd7cDvPl8vOk4G8UBE8rs21h1++d/+TUIV4x6pj/HYgDrS+j+RzlnxK9JfF3V5x
v0NPmL142kWdyAYlfnK25dYRqh6HyboiKRqg5/l2G9L/gSbyN5o4+m7OavWQlaYi7hrI65Ui17sT
dxL5PkPMSN75EDus8x/sOjYnCAA/Fgl+odfuMCn9LqlE9/6Otx/E44u8c2nhyvfXox8wncyWOT6I
vsAVl+Sev99BhpQpYtRnzyLxU7ijEDqr12Ds+lWVMFytV/1z8PPN5HJGAYfH6n4WTFQzJH6QFCf7
hTuu8S4KNh9Qq4uQB60d8xJ8o45lL6kFSUFkTsZug4pqlkHVrsV3abxSqZBa8zygNursi+lbuKDZ
DkBLuPv6T9Ih8L6S9tJYLz1hDMyobySqXwykZ3CUQdaPgiJXjmVpRxuzLIiWlmhLln59/7Bxzm7S
Jd4/f8Az6fAOWxgmr1TCaHVrjaQ1tA0xTO5fDQKpu9OPx02lCq3aOlcg32rf13JZ6wLvY9vPZX/V
2tTy6nMK25YNGWGaHl+QtJRe+HT0vo3ICnDoKMxcGvqC2aQZBrUaGa2VHniSHpszyUj9P3cco4rU
bENNIO78kgGbyq6d+zw5TdftGNkqoOVAjpHzxdbWZio3WCNLmlDP8YcIeKb5h2mykRLRqrznFdsG
hGxTWNEZk0reajglRSCwiPKbp1NJVl9lsuRfOYogZowF54qkXme95E/tiEMXL8BpRY2cY6j3AKF/
x5bBhbUpt4Iqr8ZOm64YiHx8UH8rVYmHe2VTPnRE9QxhswvLIeH65j/EgSyvvOAJurDlO/suZ8NM
Z07S/UvohR4h0Wx6mX7defK6VfmBY8NuLuHbS+ed2YlDuyIvz8aGMQQaGEll9UPfxYKlksgr4LMj
OCzpDnqyH42cu6cvE/9ifTNd0ndIS55gO7vvW+WmWzqvJJi6M4hdXAWoleE43F6bYSWZJI1GLl0G
4rqoCG3rt8lx2YyD1+ootaE8d1sFgKDpwxz4kPLqAbDIn3MpP9dLAdjmQEKtee5wyZXq9EDzdoST
mNNcZPPBxJxF9neJXXukqIU67pDV1CBTmKuNn6i24KB4X+j4hUTSUEtTvD0mcpfY2yPOJ3BmoUKf
YNjpcfh78vJsXpZFtShA03t7fxQQpc3epfWOTwAhYiA4e2IAkTdLWvT8DRZQf/zjbf0hweXfw7Su
UnzwCePThuwvz6wlBsAN/252Qut0w5seCzrPLjG/uELIyDpSBBJTnhHzNPJJUXmneDA1+9CkCTgH
ajB87WhHuzuzzVLHyN1ltkLLSsI5zuZgzAUglu1uwfkENthEoDs3YvKGXe5t9cefg4kVEuwjLzd3
CxjJrkC7t6BbxrfoHw2M2s5kMfxRzuRKT51gTK08SO2EdENC09clO3y2CG+mw0nNQGhuNoeNLNfC
fA4+/ZyzR1QEUqYgnpdwwM+JQ8umrqnpDya5p8OD4T4bDXtB+9CQ4uoj0c0S3NF8eFyrfmVQ8LT1
g4kH5YYt7Hgmhu0TnZCdehJxNANZRQSF9uuQk9VJ0Fe0KOyzMftHGFKU9RwgqTWEbXQ5jKuTr/N+
tT+HbIGONMCHMHL2i2V2kU1W3dxxc9yDdve2IG0baaHg9JsyTrrPyh0LDkvCGlT7zLzucmklzgIH
AsA25RHknPwP46Bwwq43iKyMqTiNft7rXdA3WFqmwWxQoEmPsXLHkurUxGQHtAp6Ay1Tju55hkSf
2Zkiutwv/gYYb6UIq2y8x5OQC6Lh29zxOAGWjj4KjaBw2AVM7hILkY7/gGQKHrZ4Re+yaDl5YvS5
Ys6Hpnag7EcCXixbzSK2SsuQWQ8HzM0y0CZM9O74Yc87EyAaEe0P5kgb3UysEmFTegV9oCN8XA33
CyaiMH5jj2/MMhx80UyDSSv6p7QnSR7jLofAuLe9hWQdU2TwcUbTvgvdkNF5+HAbaEuw0CeB+3pp
ty53aIguLPbJ/yaqLfNqFnEaL4VgPSSaxcSKlgRow0j/jzao1oMPIP6SVsH7pqhEGt2ABpBURHo9
I4wIJGqIhiyzx/EEXrY2rCMpdjLGq1RsnMDZaxetXQ1ou48dWJj6x8jTqYo86jfMSnwW3bYbsm7q
XuzyxGtI1HmbpaahW3958jx8/4mo0k5tYa8gmE8aNfCZCK9E9y564pw2lllJ40RVx2+zC48Cks7M
83sgT2q0TtdGjdhejmTykzOv5ksIKZsgEsOccY5tPfuMAp/rO0pvgGuesqdbU73afx86eueOg1hE
imtidfc3w6uuPWsKQoRHM1xPHGULJ4v8NBH/HuEJkOffca79asTF7wW1pNW6Hpk3IdT99RHEIRhb
Uh0x3fpvXBTglEzG9HKshupH0N0UUAWQngkvaIJy1uKN6LbbH1PiUCADMf+HRzTGkDtVXpW2mD6l
FtXZDoTwDwhqLtUm06x42NEizCe+RMxl89OUNuHj+NJmiBw6CjmfMmldFVC3WhwK/au3si1gWtnl
IbNLV6Dlp9G0nixmC0otYN/6CdbwRfJod2C++cOBhWdG2TvPro5zS6xCWBxoeRSs/lHdiXQdj+a2
xdNxusZJmiVDxWNwxrMaq2/EnIBufTk9t0EAbFcLal9jULlfIFr7qcw1DUdidFFzC/0PhfKvB+g5
qxKOPChYoYCpERSIH2QifxR15234YyEsxuKzyJyMBBxTxeXCmEtAM4S/ydlYgizNDLgy1Rqha7hs
hhQLgU2O1eMBCO2gr3Oh1NwyUV4VfUbbHqj1U2YAE3rP59pkuKHFG5zYM1DaDZ6HvNzLsfEyRyxW
HwX8cpW8t4arBfaKNKhoc3M5wbZZKWsxJM8MtfW1X9raWQlu6uDo8+GBIZOOseKDURlw9Nijeamy
RqsCwSY8r7ZL8X+ZHSpKawxGErxY4Zfc/t1RdO9ZMS4VhW0R5f8ix6TuQYzshqYTfYwjL4luUMD/
FMZziYEkA6vAVygCBSqhPNVrOuKHs45AGtAUgzU7wrd5RE98PwLhpfZcTK+rNPhCWy+YS5wPGwBr
ajy1S3SRdKoIT5Jrw1bGXnSJroveGKDIGO39OQLuyhRSiynyfBFoUc92QAu8Mk5tvdMc/P0U6Ex1
AvqoNimXO5sTNyRo5r4BHU1uGUGF6SnFT8GK4GWdG4ASc1mNlInGUcqSaPilbfF0OHu4amGoHEGp
i+X4bwVzDt4VAlnQOwe9bURMYpnmDW2Cjh5Sexnh3TlcT4henG1GN/ocTccXnKG4ip6CRyMI4hWb
rAAYjJrP4mPoHYgAMegQZdQMyBoPuQn/9a8vVEiw5LuptE/9B5C2gTEFLmS7Q2ApLwBW0iq/WHNj
MsO6i/GOutZu+MHO2MPDhEYTF1FGjcCw7quN3KQGsuIztYRUDQWvPTfw7mtRzfHPsgaz0I0a6BJn
iLb3MDdaZJwkGJigcKnfg+zrLjNbc6B8rxcAkjSfPPlbtaPMY+PCcqGHz5iRT3svkyuLRqaTTOW9
e7mBDVS0klUeGd+uqea8JXyC59czKzHlqZ8ZJWczUyAJ7UDZZVYVBDO9mvXXvNMG6e/YI4kVwx+H
TmCOGgwGeQRcQnUqsPGlDZWuNqJSFrQnddY86cnNb2aO6aIL9IHhZrS0yTt1dFb8NZwkCGTmanhc
FluBG5udQcOUUxzBPlpen9ndYdERwEwQIlwQuRVREuCOfDXoIxM95SbmfEHl6mAKR0K+dXTT1VFX
Pm4W6QRHuX4+dyQkzr5bBAoiHF9V1pc31NQ4OlSTZ9kYXLPZ/6yqPNwAMntJVNvMkd0BCa2s6xI3
Yd7byS8WzDRAa0p3+2M4pGapyMlzYE+c0POtqP+rjEHnzXhqdlsJsy9LUAdS75FEfXpnbKGwYDX4
1R+v0k5GpED9GsD8DQRWh+eZ580muaRFAeZqUli8oXQIYsr4tYsRZLk3tT+CRH6i7yGjigOzNibA
sWOSkipvMFvMoG5G1NPBqTdLDhy/y7aw3FL561cX39S/FH+rLiGmIKTQombVErWnGZ1AnFTd5/nY
1/jdXf1GBIExuX9kOLwYtMQawONG5ygUtoPbCwacIC0edpivX5kXNsI8l19+a6Psawl6W4L2iQ3i
BrNQ68qapy3iMBIv4CiCBPRKxX0N3mDoSRVTiet2pcfbzBxfspTH9Uk4pLRYTEqOv2c4bP7zd9O2
/6rg3PGHM/Mm/x7Xyw6CqVAf5nS81guBXmAgoBCFjTMlC8JUVilTtofK6YgzJxyRjlraCJFiSD1T
eeoIs7tUhdqlsrzLKvXbodDE9y1+2EpzQB6zpm3GjjC36+gIicldiwrOD9vHK8Y3n+/t3DGMh24V
jc9DHUKPLWZX0EtaYLyM842j9KhTQK9gKTutsoE85iWixYpk4Q93PlGN31HFWosEQs3jlQmoniyu
c1vAk+RzwV8uMtP7dSHzXsdbf6xcj5leaewHKLC7EUGEcjGPoATSwHZaguxYAumvMdTDotz2M4cZ
1L/CC/HBx/51HCIZPaiPmJhObwWaXflBHsihfPh3X8zEHUItHYBOaY5KDJ91pu9gkT6MuNQgi9gt
0FyqBgV6PGVL2alOp1ZVNMn1N1HJyVnvtkwO3VRPXc1xJeTZiEEXOvU+Kj+QJDgm6F5ZxUO5+eAP
A8ZJw9nvUUWlzNASzcZF1WNIBmT+Q0GBYw8skRdYBADwKlCQ2kGnxYWjl41DHo4bhfPlpYTqzTVW
vNGTdepNQIpYumbkyqSwL0ZGiuvtcXz7DgmIJoRx/S7QMK4lwznquywlxVJ7YPskQTtwM5Q2q4cA
9yQLlcC3O8sB/sBRU9WrxzEzIEjJb1pQzcR3yf0Qbn8S/Knu5cOYloBtG/Guk1v71GwPiILHz7t8
MiHC449aO7Bw2rgPyaPRgNAU8g4HH1EZu2CP8dtlHeBkrU1J4OutdCgLSIKiGoankS4ESuvnurzX
xx1S9XXy/sg/k9VGUgw8KK12dUa/lEvgBbSsZ5eqNuxkfHW43LQs02snHtjj3Tpnaq7on+KOn+nI
qUEzT6XQf9RONR9CEtId5/MEnMbZ//ta+D6R0e+s/4Kj2/JMd4y1YEQpAPUTzVFskxPTjf6v1JXW
tXxHBwNZ6ESqkwI3W9Tnv3jTsnf0UprQ1/H93FCEJpxRXYqP0L3QHcGwu5Yzwlu3dcMTKyp7F1Hr
O1j4ZDhEwRMifzUvTWuAwAagLgPz1B/433R6Om/N0GlvOkmNNJyY3EPyow1tDXQIkSGMeZFYnPHW
8Cy8Pfd1V6M6Gqype4C/PAqj82jDHGn+mU28zxjXlgdj6U0/xc4foAeiUmUR/4bmixt4OVWXxHPz
DGzz+BI66EgW+CswNxNh1/G+HKMk6pyZt6XSCoQur+J9fI7InmFcSzl5ipIxujsxcrJOQO8U/HLg
jhBow6B1+dBF+amJXSse/rpIfgQnnDcINAEdOgcS0W6s9A40N/kni/0GbjcXeQ1goItMQvZjtm2u
0X9uT47YzGAKAAjOMJeddt6EP/HrD6xoEVxlHf8T31Bn9XjlrEQ0cuVpjQa282YFrcfgTfc1aQ9L
GUdl1yaRtHxjRL0XHrpg2DmY0R8EPUeAfm7sRqwZ9vP5UDofiB0UVF6gSJRhbQ8Z73/i5S+AQPTv
V0npyQ/tYOwtCrxfaeLGnbqPXlQ1tuu1LUCWRz/GyhritgwKbrEIUUDXciZApQ2abFXstCo4zM4i
Q/Do6ygVRwwK1vISdIARgKffjE87XISqiCnUkhOvmIw0wdrl2XGEKO/hu/nKrz69YeHWzJ949kt/
5CunhIgcqm+YRQbULNPzaSVOTMKRT80m5Y+aZ+lFD1ypziHGiJ9/RSycCUVyAunBK6KqfkTy/Sle
KvR4D7N2RKhoj+z2KOvC9CLbGkrtLUVr7YHd8Bk+/oYlENlVZvBrAGGCvhVuVbABJ91UCOuazC4F
/0Hmi4L1sGITsRDeSHJCbEPp1AvPLAhmLlJ6Ij9zYr4bZJnls7LI1LEO0acYUoQpsEZLtndYgYIE
gH4UyIMVkC374uAuiiLwZAaRh7556OqHavHb4vgWLakQhyORFfUal2jKPazWz/7mz2nmIRnK+lfw
pz/GmVDQC7yG8SnRRsztnUzZm/bz7wDEef3nX+rxM2k6KCa1OXs6DAZorVwPD7hbL/Y34jSXGdLy
N9ahUncKABVIHC0IdASnpBfghX7WHXnoWaxsy7LIFvqGvlkwAPDgoFXtjJ5uEode86h80V1AGqdW
BzSfiU9LB8sRDSwZITnef8iJstkAOuEgQyIcrsoyksxQxpE2sA83NN7oKQ8LXat6PTPxymeWEMfU
4LHROBBxxX+PDa4ZKQao5gWFGkCmKBvr7y2DoigcayR5I/cmESGxlB54KuA6Hzf9HDrZsgha0h7U
CQUSTwx9UbtewHy3oG7E260atORnWs+PXfckr7GY7DpuQmXbjcOQZjRCqz12YP/bB0TM9zerVwT/
fvMyvqNDnP4glxyjtTNsGUVWCmvDgdVLvhdk+6zX7rlsY0ap8a6CX0UzAayScN0RehpdE6671nyb
5DPvKGzOfSKMwla3EnKI/NaQnP/32rSKmVcZVm0GqqKYX7QrA1myBWaKsNSnmPdGdIfBI9/+q6/T
IpFsvqmudAMTzYi8qJW3MD2ZcPGvhFA2I7uko66hrfBrNI/R9SN0vx4sRKe+JTv5zvakmKjYFCtK
Laf++L4oFehlRh7aFAG9AM4ZSaWzs7z9IxnoDLm2cqlzJQcEsw8AXC5Au0SvkbStIZqI3AeyPjuP
K/D67TDDzuVurr1P922TWgqiVUxy4PkvAERAayGM0+QCk/krDazlFcCqzACfcsyxdt72PYa1MdcE
U8AHjuLu6Ru5f+i2dInTMjZNhIcSVr1o05H/WzPuI4MUrEWib2zl0iXteo5KnZ+5w4/wtAjHjV9+
2PuKJZrhFKSi2v1i1d5KTco14x5wdfIo9OU1ElSwDyIJ40vuKuPKT7EX7uLMkPL2oyLBX5LhEk3b
2RjH3G/xZsUj41jY3EFrLPr3/mwyg+WPg1Qe9BjN+SMUcgvZlYo/+Ra8pp1p9FKEV4LHP36vi5Su
IUI30POOxq85VrUGVzcTHZIgYiySlIMHdET2/rTOqAUSkFOMZL82A3Qm7myHDu1PYmMp7+PLevLO
T5oE+xU9WE91CUbibrwIZoC+kw5tsTVU0hbCQdi8lpH3Ypf3FN0pNiEZU22v2oguKkYm7s1s/ri7
rFXTQMPcebUP9qJbxOSxdbyOO+vPVqlHoH6MUCv5l9bAMvSZjU9ipCx6Y87v2pRMr6CYXkq7BjWd
NssbWzFRT4hvcWDOqqMJjm+FEk21NVz2MIhWssKjlaaDlkXCqf1bqM8iMvTF/VWYTu/bu3ggz3/U
pZK95kMFZRPD8994VLPK9EW/6YMdA6TiicelCoBtvphprJHklWawtLxtYWjVRJ/O77GJ585bByNR
V7kpw2gSEU6bYIZ6YPL2lzloF0c7T0f9AQ3HgBAo+ZwSuOLQLuKD5WmSBKuON0DBOp+kyPYQXH0x
j2sbRK6a1FjZngMpyuqQH6BvNqxDPXBz2RJOBMgAv4GU44XE0ztzfsH2CYXNBbMeL9Y9mGj+Xdnw
Z2GxremaFRnA6MrGo5SixPaXVAkJJv/572GV+9BI++QgFOtHvKpEArd9W7Q1c10gG7mSlc7+gnKa
7mo6Pmav1zruVDH7mYLj0uoBWZXDDs1ZPAhj7FbBcju+SqCBTGOIIh1dbXeye12QOCBMH5RcSRb6
hpuGz9W2l1BUw0A4Vn1gmi9K878qGzMgUx7B857bpVrf2g1eJhuHut+wGTtus696MpGHO1ls8xxu
wfFJEk30GnUC04w5NumZQgjHcv1ZlG/Vd5eiw/j7mc96LQ1OryBxehhlaU+tGPpIWsqCeqpG1Pw5
SLnVU2E8d7/127bdBu0YkG2T1VCVo94pfMcHe5Lqg5srGecxP9pWpJxm0nS+gAQXNNR9qD4ddAKK
wBuJx5nmQiVPkmQJV9f/e0Ztud1yp4QNewpt+/l7CNuWgWv6t7VWwa1jFoY0UGOcKVzj7fsjWIb8
cTub/oOiWao+VyHdZPs40uFgRXMnR2g1aTPS5pe1+8zTUOxmehldB6hOjIYDSmeYQ6Eyih1vSshp
Leym2Rb32mlL7NPx9RVve2kU42GdAAsUdPzRDOW8kzhtrZVbD1dIMICYJwQl1UNdREzVicGpYOXS
alBRxjeyr3LHSIhKeBGrzjl0f6TJByxLWPlANGRMbZryXG9obdIn1q7hwT8HHeXajySfmFytRtoE
On8+my/YD1IuWp9PZApWsgUbVO1c1irCzfdZAVAWQ15yYrNL+8NCh4dlaurSy/iv+loWLYo7KFcG
PoRxXiG4DSv8CnVQYEWTwiJ2/vYFgxyTHAH8A8IJlRRMpB25bo0mK4yJtBx/Wu/U93MLbJ2nlfLo
CsGTo78L/yPwm0KrT5lQ5AcclJCwSL6K5XaYgs58hkR8AaA63945YLRtwd36r3gjwpFPvwhqFfSk
53u7MUQ21t09nITzL/2vZKcjWC3YFakUYQIpAOQbFrTrSaw9h5CtSS2uDSwdnhTKtLkGTx3PywL3
mk3rFu9JByT2m7Rhy81CpgHo78eipbbInya9cQ8CKQQYOOjeUcw8H2iJ3NqYL0LEZpfZCOU8ZvRr
hM0DgcL0FEp7TSIcQw646/FB+hhEEFD+lUUS2rdoQoNMLoQyS1yIasUfBczuWn0HQp1M0R7BrgXB
rSlAmgZv7lPbC4x0nRO0KkwwxtgabiHoLqFNoHQptNZUTWZh18n/tGpPJK419r+jfKB0MvKc9eSt
wbrzW8UKp+jXlPVlMIyeSDj4ltv0gjzTtoRtfwWsuXN2quPwlYFY6F8z6pFNfjCygkiowFNUNOdR
ovzbti391nHuRQlusOjjfkMRhE7HHxy1LnVBoynSCTPnSvytoFuZFciaqS9p0DmkjW7YeqVexsXH
b8jBtBZfvxyXY+ACvG/grTgE/Ay/2V4dW6E672WPXVotrYHoverF7v7Pxp7YDMk/ttMsO8IhfeYv
nk+knLFKG/1ctG/3oY5lp6MiNiIumcl5lmLC+umZGzoJ2vNx9pFf+4AkdQCUjywrpn90WDUP9wo6
IgWv6K30ekMH8+nsSctmi2fUiGSZ9d+66uYuCVMytzANLFEYl7aeCvIICaw6JPo7IJ3GgQCKIBx1
3w5I1hgJPoaWCb+iuwKaJh67+FmV6YZrdcfWz14roRXeI8w+nyEQ0QOtByLXPbZtppR9GQulHmlv
WQxfdqqR7LZfPfqyUSDQfVNFiagba/duB2bjJSm4QkDbAvdI7krchlnViXwGCVOVhZjo2zlIkOr0
QZyJPniRP8SAlPyVrX/lbUuLNkXviSFHhRGfHzkeABGvxCn7+8nvpo62RFOB9x67v/gAjwQdAouT
5XmAQ7nWTxnhC5G/0Jjk0PTBXo4DgY1QdJikl7yF8YOsXsQK0Ao6IFTCnR+WzqC8H0ZktGtQmfZ+
2tKZfNnHyMHC00tLPUKQDgRbyLF0tqhuJu8IXbuweoKQBCDJRqHnzKYtZiZyz2ib3UtNt135mANX
tt17qYo63Pkx0Pr3y1/utF7ULniyO3oT6DAIjL55vyt0QxrcXGnNKXW6W7atU+2wuj39rSDMiJxM
GLWcxiTPzBeeA4sIcosmnrpd6KVThFJXlVwRUb2F9Uod9i7BIcqtcnemjPr/xXDOfxIEblEQ6a8O
/BLpfOhpi9Bp2V4j3LSXXqSprxIQc+2PgN8MtqfWE7Oz5jQq9hhy8UNMk4t0K/xmDRwi+zE5iMgo
GOtOzfE+MLvUTzrnfNZU2NYz2+7iUaHV999+DB8wGV3dTQ7oppNOgqIHwRnjkxc9NnmAjcvJxwo9
UNGnHCDdwCDa4iscCXfYa2DhhfIkAt/7FRySF2d+1kVlDBtcWufLxcSvby566vfSyoh0Sg7OzUdy
g0cr4g/U0awh0qhyg9Oaf52by8lj+tNlsScs37ATIUU9GhBSTtXplUUoXRK+6mcXT3vsAOgpeR9B
8GsN0JJpxg/Q0/fM7nhBri0kTisFZb8lPWDZ/hPO+5eeLKiHp/V85eUHnMeStC3sVouqae/YZ4vC
tntiuJ8UJwC5b5dviWApup6qHPhK52iAO47s+u1NTNz7u9EPIgHNkhR7porxRS3KnFtTp5V76jo2
XP/S+RLJ3q1qO+1yh9SWysqE9A7CaxepM3OJAk9ObslL59K8K1I9zXk/y6EC+he9Mkn/qYAYO4wT
/zRvvSZhd4J5PcQstP3iaLrlHD0tiQ3IdG/khho1x82K4JoWTXO+nNlS6h2cjQu8ShfaEXyJhQN/
dDZBabC48qZ+cIh+CXyvyKGyazdWcwVYP4nY4qdf4PFRb9euYfNvI2nhznF3U14DlQP7FrqEB+MZ
/y19kJNJAlo48LrEDvcIwxhp9RSwprhR9lbYy02vt79dznVL+h54ICIWDWgfsn6mt4Wr0naluFk5
TToL4uz0BKtI/VSEwcMpfwu3zn9aKnWmPbOA4dYanDe8P6H8rffELK8ko61LxMyaNYMjSpIvQKRi
iJWJTpwI8dHaYvr3+tOGU5xbVVAXqx6rhyCRgqVZyh0tWI/Kk5tTbLFJq2COn29J85InonhYg37Z
GkMtl5bbmdkSGmCh6g7pwAqELu1O3/GoSYtQLFFe9BlzuEV36t4Hhwggm5O3vUKUyQUaTHTejVms
tEk6PjlE9xZWhi/61U8SUFaY0041F+Hcmpj9o5144IxvJBvVM+cR25+bEo1DzIDlZA5HVpdrNJYh
KaVDfZpNlqtDaDtihxfQsafR0/KhLURAmUKunXCr17kxUO+kKWxo02EHOQY8r+zUgM5AFXmbFKvO
SM1ggZh9iWEie9Qt5U7xBdamcoJEAbqZZ32NIMuhgCb9k2KYGQ5FDjfEY1UTup0JGrkpBf9WuXYZ
pgnFN003QpProcfU5kGfx4DW7Umb/w0RcXhNiL7bE7aQZ/sP5os9g542NkQOOypjF+7Zaf0C/4xy
VY3qc5OxflNsJ4EbUfOu9f0pkTDRnQ1C6VuBUPzN1f8nliANgxqS/d8u64srfJrZ6fw/KvmFNOs3
NJugJQ8fWcvRAI0PS/xcFJgLLEKSbaryvNmuHIVE9HaQluTRKZ8wDmhxlDBJkr0dEljUcTZsLG60
qB0CFB7ttzAt0aZNxqZj5IDHRu/S+PN7Nea076g9eYFuhbGjl/LrDrJ1bAcP+sPYckyIB+NU+DOE
FvDH3MRb6hVuDphicachzSGxTGS4kvQtuUlNF8QELvVTaAa/e64qlGnlzZql/fP/9dY3dEOAJ4wM
xO8RgfoWrqbdDTUfc5Lj/ek29FU0dLJ/mAMB3FDXo9K6dPGe9BqUBK5FHChtIu2QJ7EjMB6/wuqA
n7htZRMpXDe646RQkYeyoVoD4KjIL4ocNeElpRg3B263gl/gOsmdEL6cdMMnFBRvQLmbjuQ13xNw
f9eq6h+saXIpyca5pEQL4U7wKvZQmhxhnldcDZ3DbzUuzzppkYV1nG0GA5C2Qr4bH7v298ZEsLzJ
bMF9MSoBoJMI87B2VQ/UCLPcpGoFDjTvI3TqrCkK/qdIgbBw3YpRQvD+asqc5YHWXfGLX+cbDGkV
aYDJyzdZdefPcD76ttKPeS+0DMigVklzJlm1sYlBK7zH2690cvtGL9SzG/OHS+i4WHL9/VPayAiE
yeB6TLlLWEMT7DFkoAA0/JNxs+eAS+1lsLNZNXFi84mziD3io7PiAMDGCQuT+cXh4OnxqFOUut8P
9WMp2v3gOX7tZFR39bgJgfg8rSGT2bY5RO+/saBsYMVP2hH/k2Oyl0FlU6HRpd934kB7QrTWiFyN
f2EoEx4WKtP1Lp8kPFW6g71HmOjiBZMSJrEe640l+R+RD/+YbyrmjAtT2U6HfPt123c8R8ea17wo
VejqwHizU90GTFcSnYTDryWKrLUhPmbmDVUXxcrESFhaqgV2EYkT/0z0i4wOz5mlOd4Pt8fwXI8i
jyybRLEBGHcbUBUL3q6q62IAgY8lxV5i7wca4oOQJQkKJ+GC6DTuJ5ii0OLAozz6zFySZ7BcG7Q8
X5XfwLC0Io1Ho3AOSxN9s2J/mojry9RZyb4n7keIUyAWAFsoUW3kD2BnslPpn26LTg+S30Ra0E8r
gXQoQvMqABcF+e8ZsU2qA7xe5PYQYk4Sh/gxwm07MMONBeer/M60OLHz06Kh7qVbW2KyulklgVuz
YjIUJkV7smHYEzUwb55lG/igEjQJfzYY4wCB7Topv+WXzxtco3jJSH12tqKwOAVfOILX9Zj9+bmi
CV8jASM1pF9nu1R+6J5Yeh5aDfE7f4IUrTgSL52LtahsTHxR72xZPMLiUt4notp1x1OLhmlEWQZF
PvyS9A7trnjtZEInX23C9haUDvEJFpq/x/0Pdw1qmC7tV5hLbjbtxh1hJAo1Pnrs07RGp+9alyLD
hrtBz+xZmg2G/mz57UVX+Rhh1g+NsnQNfRD6XOW5YwP86u85V32ldPC5A9ewuEi6qTr7DIkxW7Ab
4wAdyhEgknvS2e/pndAuhkkHNIY8tISQfEOK30GU1gVe06iMZHz7BuE4cgEwM0nzJkaKpFe+mTPW
rmZIQN4O3rHPGuYMmAKagrdRE1wQ1PmnSRQrdaGVYwCHkYAeZ5z1EG3QIN2e9PIjTjbEdGxzhAwh
7w6dGXG3X1tz4mJwq2z/Iv6Iu8Li+i7C1G6KzonnjzDhQpgXN43qtdMPtGyS1vzBWe302OYQooyf
RvQxTs2hMlK/vrlHwwHXEWS21fvlqG+W1lzRx4mEzeLARuOmOsamdx3keHukVLcP4lCxwW6TMpus
vgcCzKsdGpeH5l/22bAXfwpw5tW3VOcicx6GgoBgLk45bxBZM9vYzeJH8YGxA/mIvsrlYZtL8iLD
58fkSNxFBoMWmb8ZSa11H/xY7bJ9nqbHC1F4xqJX1MDfOia3HpyP9lo9DYtIiMzbBnQk2qwSxZkb
GPmECNLwsKhx5k7YeOhwVOG5k5WTm+Eo1aMMK40DeshhFAXa0P86dZTJu5OHtj1ye2NTjEFdNn+X
U7dY1V0pMrD435vYCz//5arVUgasUma6VFH63K33W8Spku0hgdIsMvM+ryuIzbWqdBR3T1Rm+wpB
VRwI0krsIIdAL+3DwqRIfVL8OP6+0Hpu7lJAIKADHj6MFO4grWPuxvLEbGa/wlQCGV5bd4UgZtc+
Kd8DdU1LSr8Ttj+DgPCz1eLs/8KV7vEGS7j4Zh7Daq4DQtVo/T6/V0jNjCypaxpp4o2qoyQZBiLv
W/Lnjcz6ArX36UVYXb30wVQCuR7NeDErFnVrlNd4hqyzcZcnkYgpNmUiOK+DnZQJkAURhShH2l1Q
MiFtwkA+Iek0wstW4t+U1EB3XPxP66CvvJp7Hs0NduJOMyq8U8nYVfW+o6WZfcktBKPp0lgOpneA
SHhviinmv+xVFKty1uh+HFaw0AaSuHjZIUtV9ujLR5ygFmveh2nJlomI5uLKEqRFJnQWnCGbYPhh
hiTBU7WNYea92sApCwB37kXw1aRIlq92xANsStLUSZ/7zD70oFJN2ZBAHbGYBtFDyMNykzvdDf5Z
b91LXcRwU1fx4ewkF9TTYsq6xR9z4NIfzRNyRAyFnfEesDVQAzadJvLZyV3D5TSaB/d1oq2dlJc9
IS3+10IDQg5TgKw8IcW7ZoZ6JgOPSxycCmj+QNs9I7T0G0Rc8HKj4vcTRGl6KKliMA/0Bd3oUWQm
58kTZR4ZOJlWR2xw1j/F4n846Ty0TP/RYV30wGhQTfrSVczgdBLXe7jnZ91WTz+jpYwlZg0VJw6A
P46dATzf1jIQDSxo6MzNANcl9rcTFw5UCupJP3PELkQtdKK+f+oaU/C0virq5XPSpmpU/4n3+CFD
hD1/0bxtX7siR1efT6F/S4inDpl1d96w4HemUN1nCfqI/JG3Ig32EyUQT5GFcYpCQt9p2r7/Sb7p
nN71jDc5IxJPhPWTsu8MGe/RIFFHo46J7Wu3s8LLae6ZVsbx/yKA950G8zNxsaGrMunaPV+O74bN
fd+96xhwS/W81rsB1tpH99yqXZ3x6Qp3c/iqEzcqXtAax+77VGPtEJSC8GaboSRVsPQTAKupzugq
Me3aeYsSbgucXkuq61zkfv+wWpKsCJ09UqqR6+FbiLu8khJ/89P6eCYLjfLSx8PB9SF5/dfnnjOj
3b5we+sGofuinHiyRW+ReP51btWsdRvEjIolPfiXDJ390X7B+xTFz7fBpC73PtMYZWuSdtdnsDZt
DMMg1J58SUCwPqVk7GoJbFc8idqDDdqvYZJF1mGqQ/Ysx5koeyVzQWaa4DW+QDkq67KfipcqfJAT
cZ4iZ3zEpGJ08msMw/M/7Ws4YNXVFeWs/rpDG0yVmgAZfjYB1fdwyvFU6ubEnvO5zL5HMzUyujGU
6Z1HkwxFmFM9e6IYd29mgk5trj/fZSDf17wrMtAI+dF4k8DMfSsCfPbO0sIT/5+rKwbNI+AtR1lH
wf0gBYV4FVS+qh1vCsFhLy3X36fddpV+Sq+GATOH2Uv632uv32mTp2gbsQbBMLUzbvjj2VkBU0Hu
x/OKfcyZDRX7ub8pVEYB2E836MudTPgX7DCOBwyhW1fC1bhtMLQWIzr1TNgArSS7el5RUUeDqlOA
T57PRhgK0rqsLQ2alqO0nzPhTPFhrnmhpQwyzfDXpWT9nxP1Y+UDmhLNmPsb6GNaBKhviEjf3nUG
27KlyUmNz19ZuF55kovU7XyrJexwGT0CGQo3t04pbmQi1XalZrV8kcF/fkc4hL9mHlaEdjyAmjSK
p0oTefGKG5t6LSWMXYUARwFzWJ3RaHmlmC5Ot3GYS1/WFQeAzIQPX/P4Kq/exE8aiUjtizvpY3NZ
l35P62A1ECesmvFiRufiUBb1W6fh9XXW4HmEesCrhl9eSwXKX/T07pWmIgGJsQMgDflTfngTBcUu
wgBdUIzaF8a0sQsclIKHoHXTUt4tfWvJbTXGpzyuGheWV/Drq8eJdUuzvI70UO8ykVL8V4jg1OAC
Xb3HhxvH66p1kSpzC/DyKCmQ8t4BksjlIh5uL6kM70HYM6gtP0XabohtYBdKd9CqIepDUpMPFeR1
gJl0RywFOvOCPLsROGnZ2vK6byWjn1BFIMy1EsTh67WpFQfizxgsGtlGJOZKQKL81FoCTd4OXPVn
X0WEfppuBrENggIGYC6/AnGXn8O+TbHoy5HVSZc0ZAQC6AIz8t1M29WQdmD+KhKbKN/yDOKQHEPx
WzytC8RlBQ256Xdr/kzWGNCeytFgf7bbBHvykjBeOZagEc1kAXSJ2pBRaeuGbcAuH8wok9YU1rr5
+40stOqUK31kECHjmS9frXNWbAKCgYSQWJI9vDnmL0/qSeLjvpwV6VwGVxn41ZbJF7Yxon8lrNk8
66dIY2EzUMk4zGa5LCtcx9UD0P239eaZuDFmBNMtv6li7AnZSSmnLgqIXo/Nfo/LHxUti66SDUWp
mXl0ZDpFs9PhBPoGN0V2pWkxvAQBlafMIWT5yAvGalJzCrSxNDBKgI9Jk8/twLS/HwfoFE9kTVGe
mtb5eNUG7REY6qkNaAfCSxSbIbdbwNttSD300Y9X7i8d+yhyp3Bq5jpJFPOizSUrjOp5/5Fu3SVI
P0Ekg0+AdabclRPNLgjnAEUlxpNkVGBVULGiGLm19QjscSSyg71yHigttdrAUSB+gAYDdsiOMQIi
Um2UWoLhsoyN16Y9dJMzstb116CQeNQzyRAiG/gLYw6sq9lzb1MX9I0WpC9yht0OzlWPQtrPWLY5
/OsybX8smHmvaQN9O3GyL2y7sCXjvZba9VpjSkhcsr2Roa/vvMDjSa5XXo2a2XjRVrmC6QugU6Pw
ZIDWRVYkvad3hgYdx8ontsSoAGUSV8Ak50iE48hjMc7OQmtqXe+1vHzdDgCoILB2C4hY7QU86azu
HG1nZzsXWvrNp3bedYi7oF1JABInfq5yBeeiMsnm7zkIoUMtnfxhoETBKdKvhv/AMvdgwidASuoU
SPc6PGf+FujZJyg9CkyeAHYEAUjoFdktzmT4KmIbF/7i48Rt+3LkFxFtpjU/B2DWtFLCoD73KDLd
apI/LfRCtxdCrDzuECl2D/dfYvOBAtVm3RDWq7C9wbCMkOT0IYhQZBp1YuqKggBeGUleFyhQI7bR
YIuHQi7hhjKdTe/udflhuud00Car5kzQIyndWjcMlaxPB5lpVC8P8MrEr4FJq88R1iNexjBs7S8G
s/T0m/F6oLgQI+YfRjgQeQxn0gl1afz8n9B/u+im6YFb+UqPBG0D4II4soPpB1QfbRZXetlu2Fdf
OA4XAnTxXg3kf9j98xpErbLvF3pcxWDtcH1MCVY1umOPf27zmISaDXUrqREmjs854DPJtVPDyr6c
4VBZV9e3HntcW+KqR+cmmrp4BzVqwpiEywnuHZ55LRc4GKdo06o6C211vulLRpy88GTp2lAevBVI
TkudM3RYtQqDJF1CVwuMnI/R2VRvBjJCtphiFjPKw9+B1QO6vNcSiiEXrUQK9DFd1bKIH+GnG2tL
Jbt6I70nS4JtOsPEhEvSj8rb/0K2sHYcSDxQF1FvnhdMgcfiAPJKaUeFyTM3Cr4n0gzxmMi9jLd6
atk3OYn66AoQV66mSuAVooIasLm8+C1sBOIYakt9m7jBCG78HBuofrsqCsXH+KcmUSMw/VGfPNM1
tffPZjOkMV3o6WnoxwAASIWdP7xJP0fvL8LZubjq8DBvzZk+kmlohBPAqxzogyCzg5sol0v4GMtL
OSXLTykeEI+p7DKfaalTzVBXOf7OoW2M9FQXdzP80SeELX0Z+eLTgRRDJ9FCb0PC/au0lqAYHxKJ
VKFCyra5rWUrhqDUsv+Np8xbyqdheJtQbjY3krEtUrPxts97HnJKp5bOC7UVrGXCpI7tVpM7tpwW
60d3LP3vsVizMrNprYxXXE2zeHPvlqNYzmVLhXJM5xnBd46dNplo7vL9V+0nTZrg4Eh3yroZJeeB
XULz7TFKPso6Npyn7361uMxZMLTcI8X8RIlWMptGusTG5g2QwqR4+rWtLA7hvXgtGko+SfQF6ea4
MyLN36v+F/IqzbJMfnWpPro+3AoR5sRlUerfoMGoXU5+KdyK3/vfoNv3L9U4F7ydXdXAwMN4tGjA
2LaBDPv1AevuZZI0Zw/LLoripveBnXE1Q5BVS0s+kXzUdFhb1PrvgxLPBSndFveJ2OWMOOKOFZRy
bVjs7Ix4zusliNTjMHkwbh+BqKt4Fm01JnM1DMJBoW/wm/4Hy3994P6LCJsA1V/TjHKeTDACOTVp
6FPnVXP7VAXcS+UOWojEj0NieYMNwgcDrv8wAiWGhuywwffScAmgjkqpf7rPqVeuk3ccyGLGEMjP
OzjcWv4Ty0uivv92LOGSEv2X/HxaGnxZ3UIL1+dX75HhEMiYdGHBmTLPcC+S7lRU8CKQgZPxQPuz
tpfrdox6MErwo/BsXEg23E+/16y5kKscsT+zJBXiKmrHG9CSsm3dCF4aJ1ezf2l9q+yiLFKEUbOS
OM1yYfjsNUB7TRVfXc7H0Xz/6qrEAzRivGrPMA9YPCUoVc2LLXizqW88P1yElB6WB1KyE+LTIZWx
foCnEGNzb/dQ0+nc5JHEZj21U+ugxnYRPg9D2BL1SLjNVGKU6j8PQEnes5YrKaWcWUV0Dew7I4jy
mWy67jy0Bn0tCYcPy6jYxCdnpKwWSLjfNXXhcciJDWG+XQgeQq6R4VJNgOhva6uMS4C5G1/I+DLy
sqFkdVsinu4pI1gDwqGxSgQYW54Vqtj5WDS4B3ED7D3qlGJ77C4XPMDxJsi37wVGOSE7y5G/9qDF
y874FjRq/Elrfgn8+naIsGvn5bL/F5nngKlCGK9l3DSCYnjYyztu2OfvWiZbhBis6B+s/ACOyVa5
j7RWlRjeqrAok8GUHail8wneZp+Q6yeMVWWDWcJUSaXbnr73L//QJi9QR4hQL/Z3JVGRfIx+8g2k
2HECoks3thjhMeEgDt0In0MgyTrZkCBrLEq8gBw624podaqVANzU4r3c+51wqW+waO8tUSFpFkL6
3xKVb5vu9TyUJQUNm0VAQgI21QyPO4zbBVqPtyXrTeYJ+4s9fVojvxeWDHjXbLUK7OB6no7scCsR
4QrQeAmWWaxu8Re+gxATxoDMW0UZUSfZlSZyqoopZtgX//fNu4eeC9MYHK+3JH7UBusDgmWwbHUH
uYr5fmmgmAtnrfSFnTHoY3xbJDlpYNYXtUboc1IFhWKZ651e1bmKlghqNlcyrgTDtUq3iv9witok
tWhwinToe7FcestE77BATJ0s0BX4iZoeYNntMrxby3E5+NsIM8i+N4MoTo2ktUKZiVDR2ltQS03p
n7LVmAlRnUCo5it7fAk9pchJKa/Z/tTQtlJTFxzSBveQWao7guTynmlgLg0CznTrUeW7hfb+ni8N
KIY0dGF+EhS2U0aECRcrQaM6GPEroCjXEE2/o4epjyHxK2y+DVMLdagUZreMil5/l62P+7jCL5w5
ozP9QYqFRnyBGochoJZF0BIYTpsErca4I7/lfV2t9eOM1xWz+fhs3uj7HRC9ItlkBG+I14Hk0K1D
SXYGgfMC78LV+pYnulhLYklxpXuh/PSDPSYki5fr/5tGzXM0jqeRc/aldU9gHyNg++1fIJ2TBlVW
z4h9oBsgJxdvcNobS5k1Olw/ez5ronOHjddkQVS703R/ju0bJvxEake5sUbJwZ5DBOuFng3LQiIX
pqQViHaSS96OaiEAYspbrqJyEuheRECWjlotigpoPpq2Px511qFVxMONm38cRM37nWW+6KaMK0Ma
XPXv1LvA1hC+tMULpmtad4jZUADBLIJaTLy6piBFd8RXa7/2zmHXsVNdf560CAU3+M3LUlqLgntn
jLPL/RP9ur6w2hSG8UAiEoT5rq4wj16kSaIQvXXhJcT183TQfIK9XLQFlqw8jEqcYYO7r0wjDIt+
hvult9ESsE+Z2NkaVTGFBIoIs64OKa6GoeggE85X0he5xlmkqkzKLqX2B9p5+nJu30ZxqNMDj5K9
YUr0rNgRR5Ib7Rw1c6jXIFWa9NM73lkctpmd+v0iwgj6FTchHvZPSngMW4eVZaa5GrkGEYbyonwa
WcMqNYf93SrX205orxvncntwGyeVWv8nyfMtdqeSl3ApcL1CAjQXiEpYS8GnhpD2DifW0s7Iol+c
1zH4coqy1UfIuQSwues3FVDkw9jHhUT68bs/g3AJ3i1Rpur1LYqrRoTVClDUqru9aWuKR7r2mJJA
oKrXieAEZrjMvH2jHLTO4r85kk8M2b8ul4qDuwotViqs972gHBMSQF1Zy3ObbQKVgkW2ZweCFL1w
Wikb3xKkMS+7QWhlbVcfiDuQTJ4dB0RMwpq8KOW2KC7OlkHwpYrfp/fbMjxxzYdFK42XBaCAl63d
+nahAjzzXzSQauWtbfSdf5t7CdApDXy+dNdi4C4wfp9mh4ldlgxnfvvy2DIUqLfnd/TkROHkPGzo
86M+6EXzU1cC6yREPeuTdp2lAOMApQwjXC2FOagBRee2qbyl5IUV/QdmiGG3x9Pdg+6XC7WN5/Kx
EZzdnJjI1EIaVCvOcXeHYvPaQQAhFl4mm+9jtuz8cpYEBq+eNd/x5dWcbYJe7bF5ePtOdhmivd6t
8tNC6M1q6MPSXWhJ6Ljc0JeDSdcxc8uCXRRxIZZTdq+Kh8ffCkZsDv02hbVJLc33mn/ey/53oye0
ToVYsiAXmBgnVqvxp5bzxr01PnRyqGwsn0SKdVylcl5Ce+ln//yYjJg4DPu1fQwKrH58sCwLtJd9
/f8ZfCDs1WFOJj1wGu+ZftbnrnzSDQBmD0e6A0Q3uvnzh22665pHX/kQwaeR+dDgG30tVYIACBIR
ODc+l69djVHWqbt9KdSvI+7sVFoef66cVAQqqzjdcqctLcy6rEK0sINQhH1+4Y/dVHvvdJHhtZJZ
5XUsMOZ7JzvvPlBDXONOabzsJ7TdUdnLchAQURflrXbmi4ewdtQGwHvL+0gYE/2YlevU71jzbxcc
dcYDBuiPg1T+/fXkxhGnzwIWXtN+sVDkycbEsHgG/KgrH7PLC2ncWCjFNvqgI8ppdDdPjsD2f10s
61fD+8PGhHY+AwrGdYKR7o35ro/EjWLZLm5AaQcPyKBFUuVVdZNiQAMIwlno5PZbqT6aY2VA923o
hf0IjgXufoeqsZlf+lbmz68rJ4rlWTtAjLjBDpHNhB7vbefAsQdTSqJXuT5rZe/J5oMZfXZag62i
S/Ep40iwBb8pa9DJZ/k5OT3YJJ3n7fpOAzLDJBKwHpxotXfnoyofL2jA73SV1ym8jKZ4c9Syi+Dx
32A04M9LqUFwcyo3fEY9+6mgAVrchP9AgFyBLLn7eAf7/pmRPmuFgAI3tPABf/+nzq8y38iwvZ39
V96BnCgZyJr2m2vah+cNaZ9RuoTAbEOdw1cJOIpLlaQ7JBnzvjDEGmxWlDRZczkcvEX/D51asrbN
vXUBK9kHXpFjVB+HKc+6jtIkb/hsPx1KKlQSo1nN+0GAeqQNeRf5Vn9HcDR4JTpa6XUNnW0drcNi
HipSi2Mqh+Qrcnop16UzEDMnuo+fg5Ee0EU62JI/wdWjhyulAdsGznBrQwQkr5Eb3hr7/REW7jzh
587I06FsOrV81pAR7NTt38KLyo/U7rKVQWaqooAEmo3LYUHCO/h3mcR1JsEEh9tLC39MbOyoIMTR
gznwPQuotutmy/K3o4uQtBHo3/V2/vQqF/lh0U9Z03QrKSA+wgcYBMhOwfUVCPrY6ATA1v8RpbyM
YIGbLGbG8LDEXwpzrcCYq4eSxFbV6tUxLZvc/j0bRAI8Ym9j6lJh95Fa7gYIVYwFQjD4im5gSxtt
704LIztlEjtf7uq9h52nxin2hBmkz8FZe60KzkFO1rtQ567A8jbGIQzVAhyfC2jTH8f+N3Hjvxbo
7f9O+jgFU+PEUJYfQBMeDpvvg5WwBAOA9RSEPphYnRlTEP0omAa3o91RM5ifcThs0B3f7VugNygW
/qrRmaJM0f8sTsPVuGCzsap1SXoSuLfKoOLHDbfLNhmQhml5W08fcHtuc4drMW/j8Y+u+X21247o
I/E1wznY18el5iGskxZdCb6FK8xV+/vvTvZrKfBvRxXp3Gz8zOw4d5qKAfIZ9o+2hNGOqHwyTqsA
N3CCeZqANgSzDkIuoeauZBfUgRQSM5PL1vMei/KaYyEgxPzwPinUfcDg7Ic/I4Aj/fLSxSUkCbEt
mF7fDX/JvvM/uSBQlZk6BAyBAQVI8gYdUXcnUrCV3bxeIIbhpHfwjg9MiQYL1c3bwdiiQFqXlJ2+
c3xXll6+P3RFQfVBvb4nVDz/SNySVtrxzo/OR5gCJuDFoV5Lzy3Ju9HTQHjzuVuYA+J5RzX8uyJL
5vY5NFHPdN+Gbm4i3Ana69/zEVRzz7S4GO6Ryp/P+i3fpeq4q6eqN6Nd8qaRMvb2T09vYWALiXFt
ut/jIXSBrPXoTlHQUPGqlo63Nfu1J3T+mQ+HD8yPjT+s6BNikYeyh7KBtxxUrkA1E3mMhGXWZak7
/jg20QDqw8Hcf6gKbgTg1koe0MWQnNnEtFK18JalgRznaPAKuadZO7VwjqgLjd7yXLOyXlpOEeGc
i6ZZohRL3DUy+qlpogrxrKH4W2ALk5rwG0ay5CPSYC5ts3sAmyFDjx2vP1m9G8JNSeaz5BdY418J
2JDsyROE70oTLlqkOFE+JjWJ5K1pjKv0HRXCc4Iv8HVMnppVU5zg8Se4hVmu2fB5XyNwhKQGBYbN
NvMXWCwV5fDMRNjsETLl12zEViOE0aog8X75kZ6SRJ3lUiagDN0+SioZ55qg0EyXOkHzUqcclEfE
n2f35NW9IMI2w6zbp7rlhT0aTMuC30qnqkKS7z3u8u3PgATI288F747DJG/9ksId+7cBwCIuU2uQ
v9vtsLoggQChtxpNQ+xWDtCD3ty0DXuz/LsYy2g8Nfrkge8NdvCt4ctH67aSzfGnEedV40PixLh/
wwpXfJzsQiTYP36YuB2lsHLeVk8lUgVSSGYO+uff6XkNTGOWk9Y3tImQhRELdv50AnlIMk5UbDCZ
A1hi3NwDAAUZrsF3G0pQxrzcejhpJob+rhdSbqBsKETzeTccPFVcaMEJRYNkmd7wWm5NcvLs2v8Z
D5303yGcVdojdVjjYRjgWtbew8YOpA7htqV1uGaWNkwpP3xXTJhZLMoIPz4pzkQHChrUP9vLCL98
II1bxLDLtO25/HD2MzHAyBzq3WOtHok6d7oCxE5/37Om0dud0as4siCBtsOzcz9HBURp64iVPrrL
MtnLfqaaFLeP64XimzD5Sw8c1I13O8IgNU/F+P4fOfhZBI1hABMRoOPfy2/uuB/qslv4aSLgwV+o
CcR7ps7ubAXSNuWjZgQeCbCjZcc6HuC8te7Q4IKd2aqDFWMee8oXAcVkF+zFQxecjUNMb+5yTjk5
H7rhBlZlnAAWe7BznNrrksO1Gd99DnWLUcstGGqT744sai8NVNiE2GO8voUEiuc95t1FPbr6pZzW
XNdNpf3y9sDdD5DxzsdlewCjgm8fe07/I/5hdOkluUZlz2/e6SUl3bfVzIkPf2A8EjoVpU8tq9Tf
9k7+4Lx+7eGXjqEWEo+A8QwFC3y0I1fQ/gF5fKMnGeK1ylgjLf2R7bGQqqt4ML+H27WLvWV86Xb4
3a+jdKJbUJy0JfvIayjMNuJijf51zV9SLXJ2ZdId/UOQjhOLDiUszbq30pXEcZkIiiqB0qkxpjcQ
Go/d6o7fqJ3v4JPJ9AKTW7iuHjva3xbcUcYcC29SKIJG/ewH9mtWB+aad06Q6cB2NUS0A6oXTb4n
mMaUabAV/oJzKXLEB27G/QjODognKFh/V58VWqggtOT3lU/4BkyPo0wfCKVA777Fb8MAuPVfDzcl
Idxory5xYL8wgdmtmK9xqaxQn6ezefPa+SnBGZw2EyKjCXkJAPTpLt+1KGYm9gvlfSBXOo7W/ggV
ovxJsFiQDYhUMSaF6fN1u2qaMo6Hd9Vu81aRYhE9h7eMsVlz+QAEuiMQ6+pNK+GjPQlowFTWnrkQ
71nUe2u4lr56LB16H+nV4Oug/e3ohJDJUIx4mrJoNuDnMJFl6QLRa/7CqdGZgIOY9uy6pSzurlTk
5i0ejuijJZj1aUSzy2ktI+5J1sAyNPFI/iEY9S9xh10dsc+ds8AAobviPmiM0nVSjjhV5ir0IzIf
vOBj9Mow79SJrrG4CEFbs5mc3MW3ct5DKHt6wakVbNnuVMmp73bGRgX+NWL2mNzHfyf5IpbQVr2D
JUcL0M51rRXKsU3y3k9UyZvwZXHoN9ko8A68g7hHLkD1LPCOsryiQE9KPQr+59Jh4rL3vQRq/hVy
mo9AN3dS1g54zxBGVaK2yJ++aAFqO4BubAoxI0ds4HNOK1hSTKwJV2nqfVsONmExLHf1Hi0TFIk/
G5tIQVPMLnU3KYknOHp2mVvFXB7UkFSG86wvZb0GH5SepgHNERPP/8KOmlsn/b38DWr4u974xoaN
35JEhwz3TF8d9uCqXavRP65mKqU9UK5rIDVfWYpEq57oWJmFOb9ObX5iCA11uk/GuZNfMlk/Do5k
1UqxHfw0S2uufGUpwv5yzTCWHdrqIa3LuO4sZuzDOTRrFdkU+gGQhv0D7GekTEcL+GO4b9B6VDs8
ETB8i8f5hUvwIzfylVM7VKnVGw+h1qzeXMpNXGsp/Za2ezNDNkO8tG047Bvp4mjTVqFkb5fgiZrJ
h75c1CHv3B91r8yCESNtqykWqThJaCyfU+Q+cZUDHqAw1sapEktPIewZWY6QvkKn/L9xPiwKZaVi
gRzVZUNsM2HURDiGF+Jhkj/bHMme+XedPJ6stAulQ/vucGtLXBMA5HrZLGD6keCFTdjb7p5DZo4m
pKssSTetMtU7ZUtfmFDQKyrW4QIT+W8e9Q04D33FUCYsXg7vlo6hfBUwHTtzqgg1ub/D8UaSsw1/
mupD+QgKSJ0BEJOYg0DVvC17vzMv4eYTOpjr3hUN6EqOFZ2s6YlkkTH9eeqTnufjuAO2LNQV7IQa
XKAIpZlxNikU2es7hgsq67DD18X4NRYjpFGO4dkm+LLlZl2JDSqM3XCrJeMcGtD+xLHSizdNvpbC
tvo7Z7/XAuZmiNn/mVSvJIjPDLG6foHQQ7qgQQR92i0T7Z8w73TuysUJwKIXC79hJwRfOeXadZiq
OZrIT7rozpc/pOwhVsHt99y/Chr4e2yhCCfNMNK7mVDJYL38KWnYwkFf9TxlTIm2G66fjFsx1jlo
xsuISaglsJC1yQksiZJPvO7RYPRhf0BK+h5YbcZ3nAFPRNZQWknOkhfAkMsCLmvGh74Wpwu5QzfB
AeqKKRRyGDgI/731oJ4xSS2F36RUGbHRDPnHzm8ul3rXbeHxQxmABCwS0famAvJn0nkxoloHbBih
k1F+AzYpwFuLC3Fy67Bt+72fNJMQD9EOjER1DAtd8JmZzUs50aIaP/UpT/OytejKH5Ka3SHTqHpA
OISCCjifuWWa2kqGHwH6ziv7lPZvzPEhYV5ztO/KGMPXRtg1a4R2SfpuAEa4WDw4scsWpEjWlBD8
jTEhGhcLoelNrdOdcmQPXS7de7T9F4Squ0/srr9KWhWGJRr8GSsgRHyJj5Dz+oVsV+0gI18FPe1Y
UK+dTLsYkcYNzkaNHMzFQ9FhQ6GNdkhkgHN+W9TNm8AZYMmBIqQaQsKkWm5zS0RbDSoqHrmf+BHb
YWkYbq995/bp/VCOKhvbNVgiKuvXkRkUKAOyJwcC2nJPnayiUBJ+DECFkizffPe8pUIR37AOe3I8
E+SuGLBslNqsrKuGinUmEAbXmU2ejbNaRAtCU5G1r8RlZCQlJgCVxwHYfM/tyWqWfhRfgKmMPb0I
yL7NUB2n0rFEB+PW7gweP4cWt0f1j8lrG1NNUHFnIM9t4usU5DBzwoO8fIJuySxlvWdQnG/YwO3f
scZEQ3irXCOGxp6IofSQV2uguJ9/S3rGWQEcGY6rcyt3GAyBTl4B8bZtr+UXEO1+k0EHNFCZeb4g
UjpwivPpWf53tnAkJxpiJkueFbquQ4Aoxlgsf2SVBAgicaFCN9u8HxQpUrwEMTB+5l1yOur0J/yX
w3WhRTBAgde39Nzvpw8xYOx5XcnnU0HNFIgAV6ySj+19Gcyd9PgF0qwQTz6MCBOe8ftqpZsDxX9q
xGOYqpbVoCLFH3HEc7KY6a9tPWlC54rG7nQxLotbxiGfkbttSoevwzugNBbe5P2TUrjbZRjtPCzy
R/0nYfDJ6R0ktvFljn4CXDS0kCwt6BYeGtjjqE7aeGDMvkTmpVG04mV5ae2Xl7sV3b1XeyuEyTiK
4N9THk+e7P+8HlEqOufY9mXPPbqZAQREFm1SQr+bPp/VJhVrTKT0D0KXxVjC7ZDI7UCchF92UlHO
fQFcrbhsMyo/WMw8y7DbGQxJNr+BN+9uOe8xZXD7OBOHulkpX72q3SgJZwkD60wwvz2t4dyEIUpI
kt3Jp/ZhXhVX10qA9PmnPSjrboUmmRAXiHoYIQE45kjegHhMD839CwTjfASlTVWAUq9P6gjIkKyf
ujjRMw3hFeFFsO3SiWKkRsyTaKcNiHRvJmDBhGwQMwC7vmNzjfiCVrJQ7Dqh3LV8HQIjfnbI5Yyj
PXysUxaUURsWAjPWEuu3wgWSwAzfMoL1Ox+ZoEw10KU4QzyT+zxT25WAsKGM93GzXUeThQHMIZNr
V8YeNrJIAnAQqtutvq7TkqSrbElQPr/F/WN0jpU4nIONSOziir7k78CvjzCJTBqNPQY5Do3cgPpH
vtdTYcbI2wylLuFXiifiuaM4dQ5k8tOm7AbyVt+0ROjwUtI9MbUF1UJ4vkc0HCFA05QsUpRXUDtX
EYICwIjIwlmhUiQjWT7h5EEbOfnJBrhJjhDfSJGzEaYTHNUFnmau/XXaCBR7M3cSTB/qYGc2SFs6
xTXzl/QoLro1SYqtn6yrvSr6P7FG4FtUWcvbPswnCPC2r0Az0VgoCYkZNuFr3Eclkh/TUY0E4GMd
LDGcr8hgX3k8p5Uc/T02RZOVy6vgRpuJSa9GceWAYWNYNJlpsV2vp5c+dnXsUC/DnIzH92criQuR
0Ka74snhjBKfrxST01FAxC6Vgc+ARa4UySic5c7dr3snduAXrA+sc3o6ZBpDwAv7k1geb9UqFgpl
mUX808dIi6zbwcmd3ZKC/CpyPCTSb+J0DE+qqA70dKHU4PEeR93sB7WRgQKQM9bDi0MpPJohYxuV
9y3jN1T0V+5AiK8j+TkSO+p/wbXKlXQAypd7ON+JR+3mH7x6gmSGpuv+IM7CupVMmnfpVgDjD338
9gdtN70gWOnNDVxCIaL3OHUW25P/YkkX+N9i/VMj7z4pN2wwJwf2F67JHas8wyw3fvD0PN0iqlYx
H0ld4LmD9TVBAPjP0z8v0VSR9Kl0QaNbZ5agJLVMEujM2xofDI6i79/6nKBGN5bnBq7SuJJoWzOp
fdy7TMhoroPotUTvCCcCwfhvrTeFlD3iWuuA4cC1RT244xD3+2qvMjeGO9cAiasTE0Dg/xz719go
4CywewB/Hwicuhfk40ONO8Nm381Z/Oyqu2dgRX9C/+c1SaCa4Nu5RGtO5Fn9cQPB4vKzq+DIogAK
E4jjpN/kC9G/AKhVFDjFOoNgUq/gd5gAdJnAIYEjjQN4TYbCYHziWttZR93TvfuT2fqeWn24IfFU
ZZy/PCENlB2uDuhdex3QhSZ4H5UXdON6LcUm00z6ajSm3Pp0NyTcg7cte7GCIex5wWAZEOKZNIX9
vJjXzQYEaNQTRArhSQij7J34FrdzSq6L0goYcXYaPBkvqr9o3g41gl1DTJDWagpveiQaQ5WUISuj
3D6YabJvmNYD/qL40WtV7DXqLD4DuuStsNHQkPK+oKqcq5wrNg6wN7e80FpT8fr9VPzZmFgQVU2W
Ks3oFfYHo63+UwG0WNguy07Mg2JQL95JbgJz5FAPxUAOx56mrPJUAJvn3fukk8NIIoNkByfmCpmh
vHRAuu+EfolTdezcjzgA71mbonFfzUYADAtKRR8Sau9A6rwf5psnK4Ji1X40QItoczNvXUbn2nBG
iuWWMOgICCOvsGQ1C1xt/CJGmS/Rz1ae4w1OEUrtJHnWnhj89vtX1IfrgTKgyokGPC5HJQdUuOIz
h3JUA1z/xARFEI0FED03kxR3okgCAcBP/Qfswotr1aAWLhYAA6/icYmLiZZW3g4fvS71eZIhn2zc
KmKe3TjoJoKcN+jrBiwV11Mdo3MCaKbzdIBsRBjI0vCbh4MPUkLuIzg+ncw2ayWj9evcsd8PkYuI
N0/JaIuF7KmkV+cBQtnal0Z9RGZB2GpVU1JPOpeqxjeBSW3etTqoIdkpKgPiGf2nAJYZBIbZDu8c
fab8mLwvb/UYh0wEhpzuozzM0GaFy0ZUlxFbvefhuxZkq6dFkZfEZMkeE7Gj+EnTMywzGHqxg9by
JoEx9ZB02at0kPD+9VGORY9c1H0jx7x1N1vGIws/jnTVNdYDwqNSkrZsVHz1fh2SCyuCXHtJvkCS
iUMaPs0tQK3XiaJUZvkQW/1QhnePJ92vRPlhX5hpiSn/hWoamPFYoSR2A5/jHdd/v8Jd/2/8za6C
yBnL3pBE1T7fei8ehaKYHvTawWLZQ2VXUhG2MBKrzQsPEVv+RMiZvJ5l+TPqgDNhau+x3+pfQJWv
HwNPOnLQ7jmgkPNbGlI9lP/vpN1G52V4b9mehdfTeMWWZQReYbRpU//vE9WBPA2Nb28q1KBigvSC
5iVFRKxq7LDrlUA11euNn96OuTWD55SFdbPLmqMhatz8D2DN+vL7aAaBpNHguLctCXIZV70dDR8p
JLQv2VKKOJ8iIaTBQv+heLGXRMslQshTIHtZauyWrqazprylkm+l/rdxChZbhiX+GoNxzAF2+vW3
e5seS1BX0HI5FV27uhOo37lmo5Cz5iGnjO+quwowenyRFraIWF7WqrD4RPKs8xEpYw4fQUYkGjbQ
QCYKJ2vU5hSM7ulDvvfEb8OEoVEy9eSKE4ebvvFn/zfprwG8lToaqGXDZlxX9m17XJ77mpImkg1c
UmXNMyoxtpvHWrI0hSrdifGvu1+4NAlS/RSh+tDSRp0hynG3ceQJaQ7mHVfQDjljQjvIlOjWUFNE
fXmFRKiPYCKKqQ1/QXO2MCgbM4KERjs/PrcRHoQPee3E01WxukFuqamG7w4G0rLzoYLcvVr+mxVB
VzU4LTeddmIKznr0LTXSJ6HA4RhMACl5PTesxe3w2TTEoITKwz2DhPRGGqBBmocjbZTLUNnYIuNZ
LjvS56edHreLJBHXrBix327P9P7SryAojTVNB4SPby5v46xtBVzmVUGdOv8+bCWvhyt1ZVQniUyY
Vujr39VdfVtEK3Ec0UgwTDdTfKXPliFqEpJiSYN9TayNcb7MmM1ahg43+5p/MPbb7CCF6lXV3pMc
kCE0EvE5qegJz/dCmYCLfzn7y/oRC8En2Yi51MVjC0glccnZi9A59x2v6oO2Z5t2ZlXsDEV8360E
cpuQN/2ZzNQs+KoUck34fM9ixGFklFbLmZJr2mJ/hholcz+ucDSvrn6OzpkqPoflNp2L1t1KDiId
54Ihnfay2aRAz5TTw164TGuNkDZri8RjCTSxbGpjsAy64iI8DPGtlQ38AGdeUR0xR5yU92jFUJ2b
AHKSMYOK4iUpV/pljFDM2WVaiLI/DWDREJ8id3N+Ak8eGeBETs29AYBg5nnRKa/sz/okiB9/26LP
YvtbQ76LcTaMwl2QfRkskO6dNTxN9SKEWiVGTOAuiCI8BpNwkU/jiflfSppi77uB2BQ5pr9aW7je
XW4NzAZA/SCLEZsx0BD/0e/CNgbgGI7mkHpZoKR2Plzc+ZgIWSgkyeFDP2BfRbtdWXX3oyYOQhIy
J6WNbXSv+8b5GQzF+Id+M/g0qauKPfEIgAuTQow6vAQ2Z9++tarGkHEosssvs5qK7arttCiGm4uC
ohtp4S0P2WsJPWrkIRUi47Nd6Qlynh9S9qW7L1vsKNfQ0ni9oR9xF0AIZOXwXUr25ntjbb+F8xH8
d+57dHdPTTnQ/jKBWXpEr/Oys5QTj+Rp/1stC1+2X4o/juwq7aI66EOKt4bMBDUACyqwcsT5C2WD
oKXe34f/Nm+Rg4VRFqMViiV7f06xDookZdeJKB66BeMAaKJ+MXt4vR1ePqlab28GBsMJ1e7qoY/n
zM9lbsUiL7DNljwJcwd/Mvte8QHG+dRvzrFHfFSBiOjQuA3gZBFHvkYbP0VHMm4lzTrAnTV6QpMs
Qsyz1AAWgodD6gzuOm9+U8NFEXQmT/fPlxJF5AQlHyRBAlguYWEP0/d3k1UjD4nbTizY2ybENbMv
SRUXb+eX70cb0r04zqrFQRmCZ6Od38dLOl1B6xdMj/KqJ51fv96C2QUPdqFYdxQW6huUiV1/ODxd
d8Hu4RMgnUeoSBRxHmrx3OKrcSWrxgIVHZ5/C4Fj+iQXJsgxE8ZbfiubUrDvcH6NkngVcCZabNd+
2p24udk5nXbu/CkQLGpOVGR5zIEU6nYBZR0pZ2iiLDoa5aHBygnu5iaGELroYEAqsCvZopHbMkKV
Fd/1GxcCprqq/8d999NMH1nr+9UiUB8EdJ4xCvGfHd97cgmwZ8+17eB0Fpo/eyab68uT9KGtAT9Z
8QLGCtY0MQSl3KfkHuLST089+xVpuRhU26mLzNo3AGJvbvGb4QlRrAJhtHnMhEwWvsvD/gGAC6cc
GvHvqTfQi5vMj7sSOAKUAO+CsEn1WsMkMnqZklKisogECSSQ0oD2LWQivCNXXhHCPKkeEcr0GGBc
BPHv6lcj2vXPicAPy1bnqg3dhuJOgXEJw798YChuCWSg8BRZG+T0xnPKuB/s6rZ/b5scCMvUIZkH
9p+VZ4NkYkiB3UQ8E+mWUlBKepmv3WvJQCdJsAQyqUVBfMaZlf1a/1Evb7Ko6QhNEsWq242/kskt
Gr4K90aqM+LJg4Dx4cKz4OWD/9iTuq4ordZrptTqa/VgnAoX3yLW4s2VgGphQ49ZYOdGNRBJLpDU
qZZfc1wFoANzMj7JOh9TPEWxFNhN2ga7dAE2dZhAlMuW/8jVKe4JWNdkI02Xfjiz3sRmNPa4Xb6/
xu6vbxYUGqAxMghl9qvnTPg9HFFkQoGxuGfnFXdhyOM8shKl1e03wnMupDXzS7D9qcVyRrGwIQv7
KnVESW3JKwPTz/O9Blo/42l7LmIU3jlZZKmbrx5lsuogKS5ShEI8HNGc8w1mYpLTaNcmeQ+wXHTm
eNaMYjFol+2424tkgHbQ7sD5ZAyIIIhL/Po5/qSGWJL28Sh5M5cnP6g6iy7QDGezE//Fe5P++4am
G9dkU1KIWEoWfqzYheb8UTh/uGcycXGH07/ffZZVXIpfUVDhO6Qbf2MXblWeGewq50ljdskN31Co
3TyffTEZEMV1zEy0tdlJQmUCpebwq66Fdd1G2O9qXV445WkRFqLGkMTfbbyArEZ3INmNVZcu5yNl
qBmLlzk0Bi/BLKAMcOPgk+AxTmQE8cuVUL756a84aaG1N0HNcD0me3C3BJLtlwBIP4gAvE92uXvA
ccgn2eir9tUJwv6OjBQTecJKOygeajEeHdaYa6Lq6b59rjl0xHo6A3ztcMC86XlQ6rXHxt8SdxDR
EWmJUB50/FBCjU2ShFQuQpH8m8UbwglZmi+Nr9tsXbmt3OL7jP5cvjImzamaGB6pbMQ8U7GE5E0L
V77vU9HCdiVW5HX3dwjcj5Ud7/mp9A38Znr2BI8DZ/eWMDtfWJWAoZakn4054oL5+1IOjq0yFUj3
NBFruGcFr2ZFNOq965bqeotNzrf/s1HG8PX82+KA39/qWJQFNHcg3KpBJILMRa2ZUd2y58PYBATn
LW5I/5lzq29jliH2VVUhxtob9+bZ8hYB6pDm4/z6f+aiXuLZonpqn34Zpf2j7uE+ZJtxNTd+5lKn
AY7s6Z1TitnEbYf4ZFQm2lr8S7cqEMiJruTvhISdLIJx5Nls7FTidyZ6fSvONJDoRuOPa/lAYK91
ZM8Vjh5F8fQRH4w4xyTyfG3KVsNQ9ESB9l8JfEKta2aoM7Q0fYJg0/SARtvWnWTnMD9vwPOU+vCz
nY9nCto2jhd17qDQPreGrTZLRjYvvqJYcKEQ++N4VwacdbhqBp4a0W21me3qikY8urMTrQjivV65
gJhr8dwFLVViW8TXPeG48Ij6ZxZJRgy/zL7rYurblLJEy2ebw0gm51IKChjRuOaXQbSDVUjcOLdi
44d7S5NxOiE/y/CvPz4lOvs99SnIfeR3eqtRIViXJxTt3H6JVTgNFqb7yFTar2VMhwPN5VZ3QEVd
9gLRDpi9ZjjwZCa2Q/Ixcq1xw6esBPQVIezdoKQBrEVdJ2mEljpVRppVz4R7cAQV5oSzTcfgInyz
5Y6THg70mRd6G3tA/8jjVABWdRncuOuaFsIm5a213KIw+w/oKNQCDyXcGxAcCc1SPM7QtldEKwZE
frXs3pU8IDyJDnGvqUy7J1cViA7EhxA4GTnZpeMto/eweRWGvDctXF4mYOWbDYNgFMPX/CUIhxVZ
E7/HwzVVuPYpKMNzgtdUiArpU2a0AX7pWlaAGWCL393X0ib1ZpuD/3M7zDJOnf/rxCLVZ5BixVoZ
yzqr8CePwiD6jw2qEWNSt7J6fuT5nBN9u6uVxcRps1CyICvXyevwp255aaZMM71hitUJWuJ7O3xn
g9N671ZVW8doNoX53e4ZGbuOutKTaLYOjRX49vA0xDIf1T5ozhmTRedVDDm7UYWnUwwHGMQDUu4F
tm9Lwu6U64vohd9U1gYPXYmbNbI8vaZmErtMscEJr4Yx/TIfwt1UlfOOPdk5TG6BLQXd43drlVl9
T9xzNTg02UTIJCt4kCcJNsKH6oe0ovqvYzqpH3koC6sHkAL9iTI8izBjVluOgN2QE4+huw0j1fun
fjewrLtaZSarGFIO5y0bRyQ+QnwSAgjrTXWAqLNFawQSKl7dgXMHB52AZtqukOK7oxt7GibaPSGN
f9Uk85V5oPWM9BYH0/rdMdWgHCQtg6Am/UROHh6YZ8eywp/jv1YkNn4VGi6ysQVASoYHFc8GAGbH
AW+OtjTkORlkC/jzMpoJPEfoi5PV6p3m6dYGApY0psmGNGpBWCuKhLJW9LOPoTVUkBxayhi4PopW
6ne74nfYgHsdapy7OnOiF9eL4XtQsbIPMg0/vZ5BuKjVoiobw/buHTUKr31QP67ILEnQ4H5WvUYQ
PeCS7AQ42MWjey7lRloQLJvIAjijXphq9b5g6Mqu83SIz4rRRuCGhU4To4zgXq1FWDg4L39PQhy3
fJcjMAwY8SGCvTF8rmNkbXfCDhH6wB8tMXInbqy3PxML4DcNWyfLj9HmdIuxpPY8Z5sE3QM9BJLy
rL7JioVztsjmvQ5YVmjxC04OSFGgZgm8On8Q4hDEt5icOOeEl6pADygmDg4yiQfkGt6d3F3O61CQ
o0rR91ekbEeafoVUdSD3Hu+LIbAqvRcjyhmt6Jh63LhH2IAOKPEXc4sqi8M015FC6jdcaLRl0VtS
F0mQozgpXiic3H+GBe23frl5Ffq9FXEyM0ukCtfenWVarEaJPPJtrkee4y3AbW6Kz1ZEZ8ptKLC4
hvBemfx481DBZwti8K4EchmAchXWt6nY5kG/aV9sZE6yS1dY4F7qKHErqt6pt66AYpIhtuwyiXGc
4PKJ74GxvM2s1n+pEVmtTapezWGP+3zfjbNomw7QrtwQ2br8mWzw/lXpLdqgiyaH9uiCnq21npGB
f0WebHtB+o1QtFC4ZlQMNTpyKMhmiHaT3wK0QJmWuaBXNF71kHtIGWhw520IRJkjrzy36qKJKQUm
FxZcwGNPmBVMw5Q5mJLfGSkYkLhA/BS0DtQoRJlnNdEzaqw2z6+CohS5eYjj/v6VlGAPYvQ04LFz
UNtL7bxBD4Ag8SdHB6xTT7BC1HuOZjutvVvGLgDayTEyCW+4o29mf7hgLB82qy3Fk9kDXBCtDHeO
+/IPdXHUwzaoUSiTQ1EAAe6yY6adkRJeorfEEmMEnfhmJ+nxdgEAWHQf3Z3fALVbdwgnrsAtoF4t
gQSN3JHWG1s5KQxOVZNjxq7EBYrXVlTILJ00Q2dK0WqAKj968sEgoR8oiY6DZciApg4ncknxFUuu
ydbuhZFVljAcTbfIqrAKTHhKo8yuPV7rLB0ZHEqcqcpbqY6tJL3+CrH5kV9nBwqgm7scDX2zzp92
OSv1KDqi+bHNwa1jCXLRENc/4jPDwLhpkz2xox/SycOa+tz243tHKsmAO3EYy+g+HmOR3GXYb7rl
/ylQKzpjIXJUGvjBD5qpqNf3u/hLAzAJQFuR43r81ixOassVdJKKhP49FblJl+u/Np7bfG3yRBo5
mT/RIk4OFDz7yXcpwd3k+B4F66tLUMC7nSDjbr16L9kOko0z8YF0uVAyoES6a83tCqj+FJkI2AMD
oIjVAMxz83b9iFgmsP02yDRrfGMOV6M29Q0qW/ymcMYVMSRIKBhqhUnxvc22HlmeLGObyzc6aKFq
pitdOyhldCEQemEFlTWgJFyILy6/s7XiXlKaCzVbicsKiJAKO4+h+pb5AEcO1M1J/nrU2cDZ94Ld
DbdkebJgToSpfmOHxppAgm4TJq7ZRxxBAQzfbDzh98IRj8Pax96gUqoT+dQpUwBuf/PHFbBdJBQL
vf542Dp4zfdoErLb/uYSLb68u6Uf/Oyf54nOWm1Nggdmk585mffJFwjfS/kY+ZtoBEhF/VRM/ybh
3Ob3beZTYJbaSPknsrhDgE0WGrGqrfwH4UO4yN5nFt3KaNDqQEoVyZxsCJln6/PIND62fnYBsq8J
Qryo4czoOEatfLFuuSzqGjmgLgP3wzXR/j+k9E1W7iVOwmWLDfHJg7Zx6/yhXJh/DplSZSKJk92D
iGCQPTUPHBCxWs7cDS1hdT3Nlozjle1mImTqtVhO5MkOgp7dS1dRJnqnViwdwpTeQizxQ/hpshkF
3Z1x8UTaVXqvKJqYY/UsXo7W2ExHXYw9qwoXkkf1fyLJD+s7CxWBn/uopZt8whHUYQJLXz80N4Nc
hlo7UWdhR02pYCxyURBTEYGtn/6DN/kdJEGHL+GHMmHMkSyBdRVU5ZV45YnV93cBrJxa9VVLWouG
WpmvzYk5qd5nWUxzAlNtkVzQU60eEZOHv/v7vls6tXzOfbuSfBz5Gm0LfoXSmLqKFK0A87CZpzEu
MVi2gNt73152jvZhi5CucuYuBBkYHu6TjrzQGnaEmAJhKng/Fld4o16Z/NuVHIzVE+5PbzCXOcAB
s3NkfF8AFG4mOT9IcUYb+7Zp2eJ793XNCbuPqBjKNXgcm9NHtWUcwwZuOArpMXRM0/cfxH7+YjVE
XodI3FzrrIqRZQNs3Kl9wnUe0/KfeAVo76nbwrvNHFtRWgQqgjoYqcTLx6MV1a5o4m7/LrE/QGH5
hMB6k7WjXIElMejV/cs77qvpovwzLPwchMyMtT78PsX1cu6cAMilPdkqbx2LF2hoUnqSf5Dx0Fi6
EMl53s1pF+rdipjBLOnnbOBzSdxrL8hW005YwYqw97iqIOhOaQpZe+PWauubuJswjkOt1icWWj8K
ifrwYNzgyvk+Z+2bwDFheehb7T4elZ9Peyh8UuSbfCBLGUytX57usZUmkfFDQJ10l8nAondNIutU
8hHLDCMOT7k6Ks/m08vE31QHvf6M70BOLnBdXXclxp+u8vV7Js4HgEKQ+XBCg7hCzgGJZu+OFHKo
cKraRFmUgP2/jnD0ycKrakPPzixvdDMSFprryvUp6D/dOhLlX1hQDUEOaegDonTIcWHaBUKil8FQ
wLRdpDtwF11mWR5nBkVNxiVcEKoKP2SUDfLYwamHUu0RHSfQbqiIZfJVIrwpHGubD0Rx0J9cr6Qw
GSSloKMhSNmePw1sV5SjLnMRURxg/54hSo+f+w15GgtqJd4gF18K9Ci6VrOIAzVJSX5aCf8SdOdE
lN3kcnhYK43Ish0f1P/l9tqROoyEbz1Jv/ZAO7QFw2iDst2aPc1i5qlND7iTCpSpej2eh5vlxYzS
ORDa2WSeKnX7KLGi9p8cIHEFMQbfMDIov9bly+5gLvy8XXOlYGLvPiVn6ieHRDWzTgplenGNIfXy
gmvSiH/hyfl2T9UNOJxPHrK5JpMUqgr+cC7+XHc+lNuFmQif/Ov9sQmtIv9WGA39xcmMo7ubXRlO
4XlkqAwe+XeGTkyK6ockDF5tjJURo2TrAiOCFTt61YmEAd0E7phOHxE1CA/OXdlnItdjPgCvPHzr
m+cFv3fs5Q4GvSfn5Y1bWyq7prcynDg1hDwQi1AnvhCwVkuQFCcLW34vwk4jfE8XVvuYqyj4YxA4
PzSIEW91KyVo9Py4famQIGM9iqw16Sqx4kXYb8hbn9xNfHjB2GYWz4qthyhGuJPjXgBw0DNMVWNX
eNcpTmRNW6ZUSCeHBG69Y9wvKjki8epUh44giUc8uLmSGNuv17Tt6B3bBwv+8V5tlvHOwHkbqdES
i/AqnHgxG0oaLsA3s6xHQduHGo1f/TfEBVSZ1FtMTpr1rQHeZgVVHmmQiHPAlpuZa+348HZMuB7h
lJBO0lnOLthzqbtcBtYWMY66a09V0dyG42KcPDpyDgl4ZZtJeR7iVQJNeLEEds4fH/tn12syQ9Gq
N3VRIvxrnAlyVhsQ+iiRKxr5zFfIwUKaq6HYweMwgLNUzYyizcj3HBm9YBhT99M2QNU1egJMyfOF
VkuT59uLMgQgErnJ4uH4n+ybEcEaGqlVb3urh+5Se9hntPOoKL9Qd4pUeWRNo1H6g0hSVZOaZltD
eLbi5gUSynuw1JyHO0kzdEAGU6zEbb+ugz+T/OmSbGc0wXOGpCcJDmsccH/stnN7iQ6r2+tQCQsK
t1wXlp20iIhpbj715RoMPR42yVzHrVo83iV57exjAl788J3c5KsSDyL2Ce2B3RWIbErIHY+QPtz5
HsoZhnHWhuAs7qOzsI86nYgnL94bEQqJzP0SE6G61W3ypTPzZCK5oLdFTLccMAaYRMR0U2TPYvrR
MpWi0cy80qkup26izP2e804HO9anVjVJUuB1PB9G1Bia7nHWtY14KvG9dcBPSIwlXje/3bWej42i
dCFbOYjLn++u2MBUwbSnrIVdtmfYkkdsXbHT56++5w/ULW38wV0p/8s/uiRRDPnyUufRmZsYKZW9
L0jvLp8FWxfwVo7su/hb1Qzd1O8k+Wa4WWtZ8iRPc6cwotUbDv9OjW5CfQ3R3bwCvEzrJKLAICkO
+AHYS6EqKJSfvHE2Hnf2IRIjnH0jvStqanf8pSC1G87i7HyoIBRUjVQ1bXJ9sBJhTw58KNNVWR4w
k5i5mMxlwZqQjDKOvv9vVJpSEhmza9WMvliGL8sLdFlrMkXyb4QtShz2JDKW1uu8SMfVksIrCgJx
zog2Q5aRM+2gcqvhW2krs5ZZINFtNl9M2NAiCghrkW0YbnsrQ75xqAoS4FSS5rJivjWWLxo33apV
kNhbS0RCFnoYcqb6FEzN1OAvJjJFSlhOFvW9nhtHOzJP1c1y1qJOYI56Nv1JTxeV5KNXW5JPg/eE
6SVagsHmuZk3MyjjlFJkncf+R6A3JpuuiRrGaLn7A8Szjx1yI5t3jTpK4HwN/zRTV16o+P4PPsXw
56cGvKsHMkZY1Cq1iKshpJKDfEZaExobwtPhcJO9JPl4EaL6Q+jQaITrT33c/Nbxb8qeTdRLhn/h
CLRk+BXtChvcH7K+3OH528NJxrMYodYHWJn9g5ijM/r7D9ix7PesrfIm1vxj7g+0BOLQ0Ad29cXL
y9KpIjI5TBb+CgrYwmwbeIJqIKBwF1sGrm6gEzqCLOmGilu08cktCIhW1MRWBWwHZUlVgyIvPprF
abLx19+B7V+KxYG5kXwP0/PImjiQmHbTwjm0Us09xbCZOtDpmCs9OsUubzj0Ya+u0ghwI8J0dFSQ
RZJ/n+KAyVpfch4T51Q+/hU0s7M/mFYbWLRXjhm2uQW/1/aQerpXHaD7h77xcCuFuLaFNtirMtlb
/+uu6dQkqNX2h9cyp+pi2zHSdrqYxafeLQNVNWbpJYhDGLF+UP6CI2KO+BNmGh+gA60267bmrM2u
5y86FjI4oSzsSdVxFb3VgXab/aIdjbsvYfTyzQTfgs5rhaE8qi3Fqh2mxMtTiS9W65uUiYSYvis3
S6w8FI4mxv1tRf1DnREW9MDUxC29y9AZBnJPOWbAZ2MUjToMqgw6IaniSqVA7T1U3YI9h9cDhDVg
0cwiWo4ICERlTddpFo5+tZBAUmhY06Ey0J5xsd0/QFZhhDgUm+xCChm1gRrwWiWSCkcvPvbF6F1g
Ljl5sMkkQ3ihvRz8k7ci6Jz/3IbK8pdsrFfQMw5IiYKknp3cPhp4LCDnwQdy/M4rLYgfI+t9C+pG
qWx3xFratz2gQEjWbnMkcRYKAZPWxNFRiTs03GnafbJNNjjLA+OMGFbxPsN5Zvsqg9MMWYJRKDry
VWHPYtYtk8O2Wclud2SWxKIuKUIbT8CG2idfxTvJex2ycuFZ19djaeg3hVDWTas7gvhIKV/OmM+y
v0vJ1ahc//ZYQdNCISxnwf/5WR9Q6OcUFCkKSMKcDYVaw0Nr3MfDE6oU2/h4RVTmqJ27OtwHEx/f
U922CV60HsD5G0mEgPXa7R5Qc/Sl91438Sbyl9d7zWVmfbgZ3hCOFd91OCyYeAstPyZ63mCG5pC3
yEUkPyzjxRUgGKszpt85JCCq+jLDFOj9/NPrWgOqe62ZlBnZJI8pIhOIlB482l4Lj55rEHG8vesC
3hh7qO9HIYoWenj2mmIqZiohki/k2zpniSr2sLXlmf+nXgQ9RiIsNyasCx8Ig2sr57cYpI2+OzMY
awsS7uwomEJuPMfHx7JM8CmxijSPo4fcTf5sd2+hgb/ysn8qZVMJtU7t7Qd4z7bp9MaKYWzO0Gfl
NXcQ2uFspf9hWAIwQAqRNW4Kj7rVjWClAdiwkYay+QNqYZE6t7oU5+49eB17zqXATUqfcqWuGaZy
lY6oUmdUjMlKDV0fF4RClhkuI0l32OskahVsdHLCrCJ3APmvFalQtZXzDdnS5h/mBD1XroSUXsxU
KB9HPcouC60I6yb3D2foASJvZgplAhSf4CI1i8sgaFsqTtDKQ09LIsiMHizAkG5w0TTw5+c9pALr
IHCDIpHfonz0Rm1j3fsej0p+610S4tbXg86EgjuHidy+8gVvjF9tyD67HxXRBn6Vjtq2rv7scJoo
zejYoz4Mbwq6JYExHe4o8lyrvOZJcZzujcdGcKuoJwq9WsyFcDYRSGjqLlAG7b6K0boKqDCl/4t8
MtO9Nv7qQttow8xC633ahId/GI70ec0ATYoch+1mfpgb6iPS2PcYhaB/NhOa5YyDUbPDkDRDRU3t
kt+Ri1s5zwdVeHL45e/FcUvLU/39fDfzJX02f6+sAbf5k8JwylWl8wBFyB/lgNbGi6C5sQK/6MgO
8pXrfmsOpiQTjtOmRKQnObd2X4i7Et+Gu4xjNPMk0mMIm/wZuhTEyL73RLTxULxAI05caIBKjjPS
+VN8dl8wxKPqn2RB2Z/uJiXdG/jCrO0FvC0uicmQzp7ZTRPxv8v4gcfYOypUZalg9TpJoTSQaaQi
2ww1GDpBDeKU/LndC5mg0DpgqZbugNoIVhgdoyp335bRqQhv6VaF/SRBVNTP+SqzuPxvL5Xp6KdV
Ge3x+qEKVSiHxLW6k+FxhI3/ThEb154OS5SFxTAHNWKdwnFGE5AgWNS/+czaNMrK0ow8PWqScy2M
zUzRgA0V2/5cBbmqgWaHD+tfwMExvdLqxlA5T2GMXI1NtZ4GDW4ffyIKU4k1EGyAwfkxt2/eJNc3
DgqxSNaTuqYOuDzUemEXErl64AM3bhAzZD9ybS/dD7KjMlNJyaWp/kKxIa5v3BA1IFqePDDlfyZZ
kLTE0kkwE/OKeyCrkOxzYxO8QNP4YeXlaDEKW5pwT8L9/nm0yki2wmuGyc+hAdDSEOOOrKaALZPZ
FjI2nAPQcqERVFYw21LpZCxwuaFlBgEhzFO2UNSGIaZjkF8dS7vt5T6IcLemJSwbzdOqrydxvOzK
UtirM+YPzydCjX6W4t1Vvu7+y3HYhHCNkOOJp/N5AVCI3xegGevJOpZfrgUJIY9mTegplYE4m9rd
+9iAhtFbfPcPcCbwhPGePnLnim0E6EXGPjOMCFyPdDR/5qehIJVGdzupfbVo1sf6XsyEVTw6G4So
L9jEcHk6qZpzWsxs5Eymd23UoSHATJeFEyTMvZyUoo4qzVLqGgIms5t+Igv7E084U0gmNxVao1nd
yp8vmSo/j7RZOBg0wSkvjcrru9b/+8FwxBF0T45K73aKoT2mgDrWqCy4c3zThM8V+z1Y0FT+H/LT
CiruAhQVEq/sVMnH0R9SMzrN4J67xLlXt7X+aacgCw34mJz4SZY89dCI/ps5CDEEzwA4L436oNzL
nM8uEtmHffXQkUBe551XH3dAdGiIEq2+ulv4J4HUvWeN6mDZ2fav7rH0NvlEhihTdPe5G/QAhrHo
mMfGVsfXw3DJW2LxC3Hn2/Z/qvckFqWM52Mw4fFkqvUlLGG+leY/oQc1JsV6XgiRL9f8aEvUGB7Q
1rdMXSCHvF00GLUDLAFyLKmsnWSygONeNb2ox/wAgzLHIOLvkVGwhz2BwQM/+XoseuEgdiAbJW79
t/PuvExgvlmSAxOTq/mH6baMcOwDmYW/YpKByJjBYE/k3JYbUFON4yOStRpPAIcV+Brx28wyVcXj
fx3MVsW8CfXf6NqabtdbfbF+FTufbEZv5aS2SHkqPzSS47B6EKFn4Xle1H4F6TxX0c7u7aPH8/7m
aYuGXJQ0/8WTeGo8z8bTrT0kXXbzjzac+HkuIxCPpHr6Z8qmGtl7GFAK2WRqVmt6Pkyqb9VkhrI6
N6vI1YK8bQOqjCNJ+zJ1NBrYXxHcyzHU/0CCL/EN3vXQNZIaaJKIvo4EzSVRVuBIApxmzeShc/sR
5wN35Z26rqRpF/wjNDb3q9apn4BtPP8hS5Oux+mqPEVFS2hbaa3AhXKkpHCuKUTEgMVFpPDDjYoL
jtnmdsGnuyxO0KUE9JmvBJuVtnnOSdRhEBmLa5TZ5+09tPDqPkZMS7/qeI88HILXQdmUntDaRziV
uGZtwfPhbJeUJYVl+xrQHWMzV4pSTJj0QH9IfzOQquYcXNpaYxHg+gRi+QgMVfeUaCJStt7jRgLZ
iHdX1h6fKLh16Sa6+vbOXmtIOJkhrthDXeq22Ef3bwILFPd4XG0Ieg6zWyV9uYWTJPQceNzo8dYP
r0MdpjZ2Ji0At2KCUK0O3JClV/6eNNdt1cu1C2O7Qc1g7GX4bpWiwTHjVyiqSNfgBu34R0pEzhxN
LpElZVVgLjJbp0lkEf0RfN4qW8YF3ij4oAZNCc0SHqWDC5kQknOskrHhBuWHZPfpqaTYYeI1qL4a
hq7l1bycSxC496fmHX2xx7E0DfJrdM1U3yMZjprXt+L3Bq3x7axpkPW+tsoU0G31Z2A8IbiDAdK5
qWUgs2S6TITBtoBr2t8qf0RwsCplwLJiTOOVxDsInERzUVrTU1QePRVQpYnhE6UQnReS6ijlFe1E
Ce3PZd7vNo3kn23xajMcheO1qvbUq1SJQWheHqCZZwq1JLZuBL+6BbUteBT1Ir3VI/A6sKZSyJzg
AxO/FPc4IUbDOEzMQ6HyZ7DjrG+iiWbOKoiIqGuP40EZyfzm+heotePGZPuqv44ft1LWVRP4+7WJ
AQBkikmjl/hfY2HVIb0BQIFWSbsVak7lMIms7w3nl2dwVzJZckrOP50a884sqpM+7ydrbMc2hRKg
iGPYVtLv80gsBJDTzCGXUMDmb065p00UQM6VzbZu5YVh1q4HMwKVz5IQJjjNFc5G1yxPDie8H5Qh
bA5xP627do1K0oA1xdWVB58Hk3mZgRkd+qczrXhlYowrg0zDblegFRTFzi/J85EElcpYlptp+IY/
hVJc6DdKVqF4/1AvGQb8j3k7Qm8qClF2vdgjvQSuhRUpFojCwiqEE4wW6BsyF+AF18GpK9/BrHHe
7ZPFAeEJUxuXzmNGWJCc69rBVjQkWHi8V23SLD2OMc+SCaXKs9hhzpVI4dtGiVJ5r1+aMQXTnBSb
zbES3uiKFLZo6KWYSRbvr6H1BPnAPvGo1EdR3KiFHR61COHc55ElD+mCWMDZPh3u4MDnIma+wyjK
dRlFPV22si/jJWbinYc3bKM+Q3YhUo6iGUKAX3eTRULeEWju1h0vZVb8gJ88Rjv+kl0SWVMJ1Fa9
f9G1ZxPUYcUt8NqR6Jd8q8agqQOA4POrHg6WM60qhSiTdSJvCJotGsugY9LnprK0wbBCBqlCVaW0
wTaWioOFoNKdHHXfD5DfayNt3TwgMXzrGp91+1yzPIQJ0p4aFVonQiRC5MPB9lvIeYIS42PKfiky
UcP+m2MPEE+rf+DQUdQS0V0eYHCEeWNrF88IfyZY8oVYj6Zxgsf3DsYG2J68hWYu1Ns3lrVg7nME
B+s0ZJAaZ4oZpgmnHvlPDW0SUYcTFcfKNxrXX65ne4n+BPWaFZyqA32qglBH26sUVYZN5ipP9bel
MJvfRf+71Fft2x0VR8eYCUZMSn0fkgnKKjmpWO3ztkdtLe54v0b59NZbGtMDnZeZt4Bb+gXzR97Z
273FV0raJRMp49kKQGj5EcRoF2X1OwdJVVEDN0DF5Gfzf6lSqQsIt+PevMbVD7fasPhhLk1nqYvF
BQdImBYcg2Zr3UV+et5rlMu6Toubxp0EPrVc3iDqdMEYrDi6XDZY+eHCtCElnnaS7jk8vSpdeWNE
VrbGd6XAtfLm1XOzBy2zdSfTVTMCDHOzOrbSbvH3Jsrkxw30N3bPyuOLYKR7sQdRTttQ37FNLap4
e+gmbQk5FvJuMuO/MKVyZYAE3/fjRyaR/yKE+XOjwUCIUlwtIRw4Lr6kAJAVr0ADIXKX/rO3sjkY
tPX/jkHx7nIHSUiic5Dj7UsQUOYWbpuhxyQmdi3125W7xIpPwAlrXZDgzipnzUzabO/V6tEf9bKi
ZT8D38ng83pvcv8pEbIQhT0LweU/zDEFFb6V+7MK4kMOcd+1PxTLupBJzmNZJl7mjC0K1HwGDh4m
Ejt9rosZecw0wa1xLcEjjXY+6S+aj999p8dTM252wd8Niy9fzO/MWXnisWgHksrP1r9fvQjwX1zb
XC36NdqeWrXg8W+S+p/+oYFbvIf44fMMP1m7YIU7Bjso1GLk+F3ZMak4wN9gGQhKFzfP/tLeg9KH
UFKUGhaLKC+xpctvdIj6GV65AYDB9T0DmVqbIRaODD36LMt4J5f0vnn//DzIT4Yh8K8ieAPGihON
2CGNn7EQJLwsgnTL3gAoQSlqnde3ezX6lbJlg5b7yKOuxUBEI0QZ6dqjPHgIimcyb4xYONbrJYB+
GC8iFw6A4HVfZ2atTKxPLLEEs+N/+NvwwPiB0ShwRJ3WyjwtqbbiHWgH5xkM5gZPdi6tgpCJko0s
qAgOqDzi3Aa1/DfSog3FQRVy8L/VRbVLFCf4mC+8Y1qGG7tTeR2j2+ymr1wnGlPSoa94z0WTMd/x
KrNYH7JPFNn4GYNMaB4vJVrSw0Eud6v6uRlrMWW7YOyXYoqWsnwitUtObGQj/J25K+GeDqeVG3iy
U+Xj5oVxitKNEHXcmu9BjmtQ2qdJsJvc/AL1LDawH4uu5gz4jMdPakk90Wc7CLzyxzWn3THyCJq+
C+n2AjSXebVlGBLwUykP3kRW8JBtY95dSFWXQRB/0YlBlLgd+uikqbLSUx1zz57WFtZlEOCoBMGt
wF761ixj7LFNzbEx8g0xH6TqqAl5b/XDI1s4CSttJinuRVT9doXWfBp+oCNFCBIjc1ZoWoiP2eK/
LYi6tgwHJAKYMdaI7o+gdJxrc3gBvVcoPg/JpQ6frn71MeGwP+H/1XymVGFK+G9IzEPdBrwYHa1N
v+Zxb/Cesee2q7DwYpUqYNZl1zne3jT1K0IllIYAKJV+nC7dqjQvDycb43q9v2GFVIuQAQ+askQS
ufpm+tyiNt8/ymb0DFu5535JqIpRC9dg8R3wdSjDLRODI4ICXkQxQtz8+ZV7gSYATJHa9WCYHzVM
etr9PMV4ZIic8JBRSpkTBlGaJT7oZyLyaoG5eAxUOvltHcxZHWRu8g9+PALPhZBD8gl6hNY0GcEV
UGVgsC9FlkCMHQv/Io9PRgABOQ+xb2UGOZotP861CAituuRR6p1zazkRIApHwXogvypcjx92D4tR
e3uQckYEDbRAZlkUrdeRvazdh/V1TnutVfaUug7dVc3cm7e3YimHAWKJcNQQxYIFRqH62u/sRC8y
4jc6ueP8PM9xilTYJqb4pDPJvI56LKBd8O8w5Ue/Li6QgybaaWXeEPb+SE8iR/ENxhy4ODms8VW2
MHiFFuZLD9lIYHUrSfyWEP+4rXWNzXwGDqT2CXm87akymvk+M7+5AQlnbYmuwFd3nOMxj9zzfFt/
XwwGzlwyb7ZMSrlHqDRyyXPH+SzfKUCAFeYHQaIvnLEew/8z7AOAecMT7tbCyqkCNawDJhcD5A3E
GoWht2gHCGWVtsgQHYhQNZ0RfHreaB4Mk3reNEDtd8yjdC7GavlrmQkdIHQZrOV1DTC3icY886yV
drX0g+d7BjwcF9lxDbFq2wXpx1/5TPn7tjd02LvnC7GvHgF09PXpqLs0MGHNKFHcCLpK/j4i+eBM
lUpzsAZHKl15ejt+kJon5M9Be13bf4+1ev9EV2b9mEUWp8tHIr2WLlouE9mQW7awwS/qkviL6gLH
bOIDBsQmXvzNxKSxHoJ5TJPS9Fmbzr4GWuPphdETRoFg6IWLeE6V6eKvy0nnr3j0fMNrF59SZpAw
AyzPTrD2EZo6X/s3X3FDqJUS8mbldlnZLTf4iBgFs3rVJfTzI/wTQPVupcN6e4FGAg/0tKeB80LQ
jLQHEXEW6NgZJj8FJXhPBRTE4PfHvWUfRk1owCdn+rSc4Oo0cBTDKagoicPGsKG848/+WL5cbj94
ZDFFg0+WImO/28qWvwTamaokbxTRmphviB5UuhHoSj7mns5YTA1VaozwxaZQBqq73Ds7k+Fej++8
7GS5j2pf6qUDZeNAmtAw1TFjIZHpf3PJcfZcVeO5BBIwgxsICW88snL6qt43I3eMxI6S513Nxydn
QsB6pXtg9o9v1rGMuvj7vybV+Rl1ZQFdmOAWdP1jjjFjRIuuyvsqAQ7dWk3bj56zGD/YNVc5BVKx
hFcPCTTg8NV2wA8slPJhEducVtoCOahPyJS6ydFo4CzuXe14A7QpvhP9viqsu8jlpuiW3XqtDAKG
2NI3yC+wRFqVTE8brykjxJgQFIgiw8g1hIjS+W8NllPtg62GqvU2iChBJ/bDtAP/oba9W/n7GcnG
NGaPYMeXkBX8AA/LKdI0CqgKBw7N8ewgxG566cnOMY6CjS+AdwJ1+CyBEHDqkpPxkCNbnthpenQh
jwb5gQjOGO68052MKJOp3YyxMzqFZ3tfXvCkhDVF4DObRLPBGzT6ZIqfzzbIupeNh/Aq1cJ80ez9
phl0Qm7Ysb0xqHcfMzAAn8oHT7HLAu0IKt+Xetquo4rpkF8iv6DL0B3P/56EkUl/2R3jPO/XXF6R
5EdP+3m/F9Dz3ElSEtUgtrne+K95sU4fUYwWobhwVf9sp7JE1kdC9V1SMfDUN/sHixZb3nDPhQj1
gOSZBgZE1Y/cmmS7LuoqfdVcOvpzKrU4YnlGiofaqRi2+r3u8mxWfdhUmDIdD51koByu5h9xCF7L
ndT6LVJUTAnkvr9fKuUPtJANhagkgeZdR7PPxdbj3zU2sFEEjJz/MPH70Os0fv9DqoRszo+Nm6nb
3u21oDeLYO4PW7tUWovr7YuiNb2ZrYeoDSLkWvkvNS9u+52yPWVQJ+PG+e7I7Fod523E3Zu3FbUB
AppOKLwlw0GPyabjTYb3uPc6BUqhb0OZkTls+rYD/Umcn08saNN7nIykboUimINH1bE+Djh+74/y
0hSErGsBbHQfxehTvFVnrC79q+ZErlzHuqXlHbpNK54lL4A3btwLIslYPJK0Qh7nN5kCqha6OmeD
Y8s39CJk0BJa8R8yTLo1Z4V1O8yG7fzVlbvQ5xCfbdSFnGpZefBhqz4ciO48CJPPD0MF861myl9e
YWq1FzoKdB7I7hSkVZoI2yIAEEKi8F7Mf8b8FtSVvbTmaKCEMIS/8tFMuYii212nOrnUqm/nD8rq
14I1N/JpsuxH1MMJ6Qg1OLJPENm0UDCQTHoLKsW9RkPiv4C2Uh8bMLm+izItxLFXTjdMazp8r1jY
rP48q0Mfeosg0Pi63gjfmULmZOiII1zDWIuMB+FdCGQ/z68lD+vANm8gXuMSUl+I++nAHdD0FERN
Vlvbpb+ybvQBuS+nS91L1AUGv4W8Wq/9ByGBNr/Aned5CITn7TPwEWCmi3A1JvGjoRWG0F6Pzifz
o20mOWmayK1fsDXiEIntppOHxQvQlL6HGx2NKL6arA4oewCgpc/HAAJEfinQQTGncArziN1YBeg3
hzRmo0xVya2er22nmL2xIzz6XOD+bbmJlAArUYJmaLSoddi2f5zZDoVYMVZN5cgYhD36bputsXUY
wHhZxxVZhF8uhx0w7IP/j7KL2k+7+iPsQR0x2lsREai3zd5BBNq11sb7btGUYm5W7qTqF83Ig3qy
9INysuv4EpWf8CJIWM58Qb52/XOjdUmG/8Ch4kbV6cXaOZwYUmjbwv2RGyMXcspVRhSHlRx5vUXq
WoEV4akiUAqogqZz8IqLM/E1UXOf0NwgMi1uO/l3S0TkoRO262iOg/jRsY+SqV4YqsAWhn+LBBMe
/JKvCcEPQBsysmpk8OtaqCY9MGGcrwQUxwRkd6qzdW/O98k83dZd19v5tDwj84zmrhTPBmEAddHt
sssc18kgvr5sz3eaiQl4eiEIUSMOE8pdUurcfViTFR7PbiQrKUNqXYg6nMH43+bByOsBCLH8h/vM
9jDHxE5x475NQm5f3yyKar1nOl7MHKgxN506EGu1+mlaOGN4zdUtgjStC+XKFA/OFJ/c2SiNPy1w
M1j3uscUsRnUXqT5UHXHLrcmv5azf73uzsZWd89BFS1JnR601sXiBKNUbUmAAtWsb0DpBTuONtt6
yAI6Yz8J1xC1qdxgwZDh8ZnBinJJVG2CW92zw2p8jGLn6f/RM6wNdjCp1mHe3qwpkyXf/I+fuX+s
r0lmWvhfLcHATTQqc7HbeXY0uuLe/kDNNC6IAn/Kx9uyizUAD4/PmtHJU+AtBr2nJxZ4mqk2/vHg
/tlp44jaeR23/+0yBrCxisxKN6y+5qkuAlVxFCrYWKwyQgBLLAs4GjJnoPVOTlboTLsFQsTXUnAj
FxrAo4LQjlHPQBAn0d9b4W7Gg41E5UllkjIAIVbIVIHLKQsczohdpPFQxLcwwZdhLXR0wpu2GGu6
UuQYMUgbKEbPsTf+ifUFl+QGXff47LGv0My2xZUVlzafCMC51V4p8JK8vg2WkITeHNkv4EnyOQaU
iBa86Xw15xaYueHkhLZuPcmvJnY4teuuBm/YFxgdoRkYZn4tfaKAAYjDPEDY0VZQbiiDcfhUUmb5
ed9hAuBde/Q2QdSnHpMmMuJ4H3pgEq7DxoN+dxgS9UeXh9wzo4BfHNcd8trCrzRygNQcMhggvN8R
Hnn7HIm6zfl/1h4jkYftH1YMdqiQ4Au0I4XAlDZY1SzBejs6VAD97hqNsNHpo01O9WC4LEAVMkij
rathmUL0kPBOpbTRIYOdk1rKW4XB1ifoaH9Oo0/rbVYjX+A78tcoaAOIvTpNZs6YpxLtf4DQAmW3
7fZOFIQ9S/wr6jy+FFF44BhwM7+60RYqtCx6YrAJ1BpBNl9aNt0kcchpNdZlgSvFPlzZx6a+yR91
c5gmrppklD/u+3UlOBtQcWo+f2qDQTbWt3EYZ92XyGaAC54BnrynZdGaPpGFbEsT9Q2eF8ITNNjh
2PuHROZipIy1MNUAv8Ah/Ag29+AnPwclnW4AQSB6rCFtF3mcP7d330Wuvm5+NQzfr43WhvkEs9I+
AKZwxkn1+quu3YeI7liQQNP9milG6ViNMqb3y91f7FbgPbfvwuMcFcY2piGAEIhzyW+2ZhxNuJru
aD8yF7Xn3bGfTdee8bsibIEjWv/mwsoCHHxs3GmKLUZehwDPtcMYB96obncNRPmQd6eQ9hZrsjQn
r8J4s6JERmK+kwnCqRbUdpUIexUX5M710n3YmdXc1va3oFgK57TaikI59aGKbljA3lhqXgv+nkir
FDeyM2vsbWB/Nh8FtaOdFQmshVg18i4fZrPTUa3Ybg1vFOUx0cvhGHuYtWvDB/H52ClNYUTOht5I
rXgIYrxmmoQrSpnBq5XZ2iEkv4oXZn13kVPgjosSfqK/vqK6h8jN8M2H06VBryRpm0eN5EY9wnZp
/EZ0ZQEP6kX6Cw/YUJxiB3Bb9iUV2iagr8gf036G75DQElQQUtzaHoSrEWnTByBUhY7lNV/djF0e
k5ySQsutuK9okWTq9eCFRkLeep9QplCEgd7o1skCo8QdAoFLU7+jUJ3/l0OfgqahHm47Zhu7J+KB
89SXkNt/pgA/0/t8bFxrvvLv3HhNICyKQS7o9FhAcbdsL0sl15wHrO6vsGjHPyD1+IGTkG3NVhPm
5jvVdizBzmazaClUaVXHg0A3EbaTZQK5cx2/tdCA3ENm13u0pbu4fNzUbggpQFujmz3Q069zjPsc
/TKT9BQQBvbHbhOPwv+PdnRrZbJCIR7LIw7M0i1wyEmmZA5sLd44JToQP1XcbM2sden4067X4gXr
aaRc3iZcEzVt0/Bm1Ndhm3fdoqN63rdEcwgLJzmuOEuCvUdEdkyn8RA4ptIH3WveBogN2uMHXCeV
aEWmxTZOBzDq7RKNv2eKD1hiQ6HfGn8866Xy2CYvJ2T8snhrZ454vLEDhgk52OMYCHpUWsWksj0n
1N2OsPi2MblnQKZT/7xXgrwAto8kZuxPNdyWFZvFrNugEwMDnuIgn/cTvbeItfeCHKZjdI4x1Pli
ud9CuZuu87WtRB+P1all2+75Fd365VBXxY5aqyjtGfbN1CeFvq5mkRE+jLDQPTAGMPAMVkKvftuV
crx7olTxucd7zBue2y8J10C/2Ta9VA+PKyhJjtq2YtKmEEoSVgEnUpKXdUBt1cs5SfNSpOiUJfw6
yc7/Vd1MS27cynAITg/wHTv1pB65aL32kaN3uOc7QhnDf95VhOYciLCJvo4mdBz6JsEtdZljD0XH
erSxIaBUUfEFQe6ACMegq60JaVezJl/+YRSYFJDomOHNvhhimENmSjmXd4fWDUJaVdS2Uew+Mtug
lwxMFF4bnCNcdCdsoEX0T1c4V5T2xR7lxoHdVUYLjW5H6mX28n9cbkhXPSOqvXUHFBGC9tRImhwh
7az4odPYwE/ngC4/fBeV7faLUhm/BgErT715Cx/XiakVVvVXyrq0lpQBrcIqeHHs3SzAgHvEaqya
eagAMEg8bAMFafuwx/sg7tBt2v2sb5c5rPVwCjENV/rVeWEvhVYRigexm6TRLALJBQhKZH8xvWWY
UmF7uNJnb3OVqtazAam0bm+Svu1dlMjsRXmvXuk+z5zi470QjtB8JeujvPDIZu8Njnm/CojuYbkE
cqm7uUhjXzvU+Or32qv9li5cepIXX2AMI9mhSyi2X/WH81k/umNq/gILLAEeUlrbaJ8BqecOq6Cz
X7FZ1z37FzW1uLh3uyGeRzr3F0kHO4q5ag0/NBmHVslhJ/reEyMVdCTCiWHajXgbUtI+XqqzB/kp
q+SE19Ix3nDJR+Aio1t8YZ3/WYxiGRpsIQA9btR2F8VDy6CGSNCpo9Qgj2S3LWk3B8W5RCyDp3cL
/SIz9WP5jMqQTxSsKzQ0dNxktC++5xq/ZL0xf76L+0wldfzwyHiD6bSA3Ed/m/TYdsifQVGYNrpB
/mRTGqFXSkv5aeodMg0i9pfk6T6oLm5lPrLwCZ8RW+EvjItsy6CBPqwE58Q4cpKQRBFo5BWhiiR7
jTJFhS6izNsdqzwiGxE9xKWIPvaot7xXFatSZYsPeGda2jqX8e6XSd+/hGkwhJWVi1bymfEODYuB
iavK+jzCIFDnCDcaFKiSuleNA1GYJt6lVVJzGXMs6+CEMQ/djh0pMdCFDE810szWfsve1SfPcqG1
o64yIHnpvwjfQ3cvwbPQHg83885z4xKyTLQAkJbi9aKYBFnNqkulDP2oUdeys7g2/ZUMe6E7KFuy
2GaKD5BdXmDN/ABiL8gbjwDKO0sMNG3SDUUyDCRWrGB4RjQFxYT75onh0L1bt6S9+jDYDymumXTM
CNumhMTeUwV470HyM+/4sLftUZG0mSFvdHAG4Wtce3hX1xCmBHUTJZG0yhha5ghm+U0TIym0fXmR
ppirg+eljII2Pl1Ti00mPlgAT4N1cAKNiQkDCclCO7gCjV0aT6JuN2bXlWnSKt+ApG5bSKKwpPkS
BjvqNX4rM4yjJNXQ3rzM98HTjlvtuNlccfE83oHB9qa1JaCU7ahR2LOj64MeP2WclyP9UNNZHr9J
dQ8Moz8XfdOVc/1IwOt2zaa7ygMbaPFycZ0zbtgymnoZJDx3NnlOaqwyRs+n2GvMN6RsSzIjRyTJ
bgK4Tddp6mhg+YHLbI7UDnBLUJ3ejpmOb3yF450hgUoupAYpLKl3o9UvkkqMdv5Iy2d451cNPNL0
nT/tpbUJMQY4LfIXzbiclUB6qWiDnt1KN+93NvT/hu835P1gokF6qj0S4xtjGz/OR+OF8rzRuZ4N
ppQpanZmy+GQrGlPpVa4AqgLIEyZTUtrWLPMZ/qnONjKe5H3il6DsGmDHI4uH7Z2HuL1h5aQOw6f
2SWPM5aINHqMynKWZenbC/nfTNyHbE5smmputsEMfzHphNmW/IlBoaKefCzLBeuyE3YGTWp2B8oT
RPnV98k9KAfNsxwYc52hF9s/CLRmtlaMNS8Mu3gNyU9SGip5b1uKU0MqD0KmOBvfXVMLijftqpwn
DvLb6GFM7aOKx/u/0d8KrkNR7SReYBK7vgyeLDdMTwjX4IHVBoBDMOkHQ970y24YcLRuEjht/1j5
wei/B8cM77nrnoOmZxvjm5jL7+sNMrjVvJRMw9tO6d912FUBdi3A65ZcIFs6g65qvntLJkhWaI86
NDl0XO5lRiOabNIBIfmaeLHEe9+HlAMOZFgTW/K8YDtKVyylcHkMraqd85LL+rVwwwq+chJ+1F1v
4TMFtqLMpFcKUkJaIwamyXNbIj5T7tQqDWA9zDXhmALeYJRxPxV1WA4Pvb7JXpbT4wmHEnBj708d
Z9C6iQuf/fUjQ9OMRgub1RddbZDMci3pbquD9foiV5ommQa1qGjohL7/Qmq3Oz6gxirPpkOuYjPH
/SEmEPPwwqqAxpXcZ2qjuL7UsvSjfh4jD4DtpfcEeGgqEaQOZ1ny+oDjGGqE3TFUHFYYOxjb9bDg
ckReHWvLHPqtDe5sZHC7ND/3uK0oSe815XsWiVpCUIurToPbmv3VYsO6yVOTT5Z2kIaI7parMfab
BiVKMyWTaYaYPAVVnUXBuAlEB1wt0Nzfw40JN4PTK/YOfkBBMIDksCVfy/6eJPPYaDW3CL1StP8D
8uan7/Md/HGY2jVSuIKocUd/qpS8djQQK7sjQW/P8TXVOJ6WFFROcwee8Z1RXaiHMejuZjlm4f1e
hjTvDmJDd3E5vwXNGj5HQoqfLkuelhi/UmuxzJQLOZAp8IkFKtdyHHCPIULfWmB33HxSmxF8E7ix
oGHvVViIp9vlrn2lklN2bL/YYTP/oboEypCFziryXO7fqAS1F92RBGBCQqDLZk9JyQvXLOSsLkDL
xE2EvIZGQHuF6XlWI1d1E3T9N0iBtyIWgVLgyjjLTmibVG105dmymr97j3nI70+xD+aQKv9mc2bg
krJjw4rtvuY5WXjql3thGbirkUxZWLhGGgKb8aHXqMn2hAipmtnYP2JjwhBqaRCnEeGuoxm5clhC
eJFi2DCs8fkhC0+XLXHif0aVfvTwg1TFGh2rfUkzLvem01zBLTfgk90vhNBtW6iG/m7oiOwQJkYa
OZUCkwWfJXKGx4iRfpG1cJ8FDme5xZSeVYEXx5x9HM8ViqW/6F7a7nxf0aVd+jaeSICI5IJmISai
29GG5LhnrPmrgTNRdNAZHQu0qvSAxBhrRetpz678zJf1QAnSt2+zXFzo06daQXawqLsQ8FQZYuI3
0jDnjo35or9h68f4bDXxD+SzvbU0RGgItHJt4wOsVskZAYOsQk9eq28UU1SyPnB9bPSWqpuE+IZC
H1RNmsUEeV59tfFad7MgGa1DjiEktEfBNME3+X8ivYdSTttSXixE9Y2Gd5Acj2105RYHZZziSCAY
+GoGsJyBe1vC4M25OiOnOFJjcqrfV8exewZJEvSf6FQb3YB6jVAmMfYgMuo9IaxUAxwc73WTIfce
mEBEisfYSPLCyGFtNKK0SsR18W8j0jVJHpvwXf3h7OqUWkhqt15cO4ChIHO2078fXZLCOux8CKEs
jk4IqeFpzBOH7PchnICLgxqrp0a+yJTzLzlZIIdCiaGvtGOTsU9nrC++ntIiNMRPtgAFprHtK1XG
n0pkxNJnzwQxi2raZLWUk/1/WB0ZLjeOeb2m7rWcvyja2rqvlzMNRSPIY19yuMpLuLNyNP64PHIa
+YnZsNCaBXWM+AOqZ6DXzqIRuIv4grXWpbsY3GqHSDLKQXgeZN4sZggQfCg5HEavRicK6vT95CPs
zlTFuMKyDHDblGAfza64/hH3nYtmi/KeLt96h2BkCbif7qzy7VendLCX8FIDRY+1pGJsTT8INWaM
mqPjCc1xWwWkfg7+xz9MzRapE0iW1t+YBmqU0f+zDXu+NAUcW8FwOeSOMvPFTB/6cyYwcbNL9MUq
XzT/Rzbz4izlGFbjx1wQKtITNM+rcD26JBrIG8kCVN2PG3eg/PaVl2FAVTXSwRvErXOBr/DL+te/
tYCj3ddecaPeM6xGveOTw1Tj7NN6GRsf5lynGfa62WVG6DH+zwt+7sOp/Ssf+zB+/Bkzb81Tuom3
2EXYBJGUOI+ck8gQxgu93EoQTFKCgZk3G3x0fmMsMj+K2Oj9O7xIfhIeRCOs4xQCGEANRwHov6Fa
42xzEDU20ARGceVklWjJf1CHBwj3Dm6tZK5YemdDGhFGNiP8uTEiB9Dg4D/CIxSjerEgtd0gcr/H
qL87Lw0UbxRcHbQmzOhErmfssaqSwdkKcbQii7Lvp19onuOHO7IWMC9kZHuWkeimGs+rlIMRGdWJ
xedVU3mSh06K8zx8tETE6lPGCUI0205TK0UjgA3SmYNQKYX937jGJuTqBzoX505e/08P1Z6ukp3A
HCLzgdvVWPer0xNlmBUgH7cBbG9zx1EpRSDG+4t70tj+0jFxGfEaEU/CLSflenqP6NBzhDMk8yFD
idqZbtLQzxL7f1n5X4Mycz6fPbNccZX8xXyFAXl4YWC5W0+8j7YNpfndjz66ZFQ3fXETagv3pWxJ
i3pSPzKsuMs4lwciFIGF4gin1RkWcndVGFuqyR5WJBxW5AhqiM1MF1XZtci2uFTXBZ0Qu1SkiH4D
LcINMLVey/hfPGlHwPoKKFQcaIa1cH/eu4SmLImex+XtqvlYyJxEDygugGFxLCyQUwUSr5XqJVyK
usHquEXWwcvrRxsIKSctGJhtVHmmNXk4A8jkRSZ4g33c8cpWMeJHhcfPWI5+nULkYmPV6eC60WDw
BloEqHAea9kxAmSaIYN0rxymoH8RLGaJyF9o9IzuPAihjbCgc87kqez4wdPXmzdd5Qwxv8/PInTc
dcpnOjEDYvpjRFyp9xb6jZbUmUuDCfRgWPI+gV8AOGuNm+5Ei4oUl/ZJd3zMEKfdkgjlZU8m4T9V
88wHe8QroZobBqpnNrUpYxHAkjyoP7q+ULTn2XmLfx1aiRs1CZqEknM1JAQ7QNLZKgjgryick4E+
GHbsJkdJVOYASpgF6MXVjWbe5XJ5etxotgMd4TzO4b3yvDEOm/kN2s4bYrPEwXfJhe8Z7kE46ne8
wBnDnfbKP1Rft0uptF90lxMVrtHPIbzlHRHssKkpMEBI+pyoGqRl3Ts5K/Dupiy0Hq83sLT0Xvi3
yiJo9HQFgVYmkRvjgMS+hS3cF6teVpqNE3zK1JNPgk5FrbswxNnO9KB4Ygj6Hk3/CV2lQw/+1ZjT
ukHtS8GDiszVDKKgWX+QkqFrKW2QpnYMa7aEjVlsZ4RRnW+U64l+XADxez5WO6uZQ6j0KpNz2Xtr
DUNGyY6gMWeRnKmJaaBrZ5kcHi4QZyTniQT2UBF5g8tWIBH4GAyF1kt+YtUGDiws68p8rYCx2NUT
kLA0hGgbzYCNPQRhLnTwYsyL36t8xI8E9RNOsSrCq+wGXALry4ifjuD8f22i3MysjMi+8JmWQ5mc
4H6kTnY6xSlNHjUHHr/av+QVtyapB5kVjrheAreoZLVotdxI0BR4pVnkVtQWLeu9cJjOdXvBvUjr
kMn4eA/8g9xNWAHkt3N1BQpb/Ou+upxhY+FoNBLetHHcrGuKIbxbkIRJqh3TTK3X6MbLUUStI1ns
C3aGF88yiVDu09E0YTihk/zUHPFCnYkfS7bZLLPaJv85CGobLhxslbXVaYTW5REn5dYictSCb2+c
eToJKnvr7XO6DWeaLbYhCMfHGweWp0/me1KH//b4dW7wyiGvLVkT1XIy6Alp1JGhFICZwoWhfoCe
EXitCvDx8DKe6n69uqDPCke/Z30lOScq+c51+r5c3l6Yj+TeWgnqUWuahWIBk1djfds3qSJJb474
WkTCGfllL06p/AjCnxEFEghfiPBX/mDMdcWXoBzC+npoNlEaLqbVDaVwLprKdPjY2vp75qmiMJaj
F3kWXaw9yYAWCV5+sRDIBWXJUvQgllR210n+ipfxXxiqvu+AWEB8PRBMcbgnrLAcA+ZS0Rm8aAez
CyMNundGmNbwv1vzfEpqHUXhFO1MJy4YI5e7aSPjwP0xOw3kftxKHXz9EbUajxK+VjttXs8L1Gq7
J92kF90jH6Lm6hNhG9J83jPScpjBzA3LZjj8UawApaW7Fy2dtrN/47gMqEMxawJwIw0imxYbcfxl
yma6KMiDdl+7n36B0JYMvlj/Ke7+jg3Ypw6VHUCvpoHFs3kK3OaaS+jhZYcQzL86dvwco7d+zl4S
Pqv7ZIC+6t3jJ5xSrzaTTwVFg+CMM4e+Cmthi7Y6JZd+ohA31e1QQsiGhQ+3uTlyJuASNyj7nKZ3
uVMP3DExIuOegZu+Br+sOvc0lM94s+oY/zeFcVmbD6CFJG950WM1knrHr4gGizktrgTUaquuKbZL
avHHR6lBsWP+Xe0i/IHeGhrMWKqnYnvp5NkvacZUZHM1ZgX9BvtsG1TmP9AtaztwxKVnuAEiwb3m
mO3o/DrxwKJnpD+SjFp1r3/K8jBhawoxt4FtyLuBiKfUhmG7eHtHsDduImGS/Dnin5zagsbWIXfn
oIpVCKmj9m7BsELJlsCxYKdWn/uVykNWoXTyKvb22xo8yN4xP6MeVx19cBE3msdD4Sl5FSRDOaEh
NhMjnTZ1Vg82dVgP6yJxtvO7o6gCe91YPHJts2SRdlEvSv4JbKTi/filKPViVbxANJoSmBEv0xpm
cVyEi5FTm6S74wzd4jZ7q+949liGwPn0vDkE5wQZT6OA8X4sPoLdru2NkD1zDfUXRDatuk5QaNDx
qX1d1G6+iHauV9I6rxY0KJIr0oBE5ou8/Z758zH5fH2ITrOKm1npeaimDuQzXyuHvlU4Cogxhm1c
CKUN3DjdaWfqf8T56gkgUdDef1lGpUThkaXyHyD8gsb1Txr9ojqaXxczx8KH2OOVrNEzICeh7FSX
iRc+cIvPqd4Iz91sYgntpYrA4AFPnnMhyhZE5GSKtWppMd9JhbtIasUh//ARi0SggcNqVZ4cHDyM
K+nyud/UNikLwpIwydJsHVsbyY5AN6OSdjhzi12mnLYpINhjl5jtfSGBbIi0FKWl4Bd+kRYtMMBK
BJA5vwD2brx3jKquKe9T1/HICaYcXBwnUOml1VEJ1VtnEElrD7H8UUVuL90GxvMylQquYi/COhD3
8qf2Es8CShKD5O6BEjzouES97O0fS/WGT6eU8tk4mjJKrlTlCmtSVywxlkNJ+uaZiw2610z2YTEf
vOiSg89NW+zyPa9FqdaM5dkZ05DvqD3SIXUQzehFszWhvQPmhng23xeJoOwnzAmS9OKV1rsCYDtM
VoJUhxkuBxkue3bLj7nOfsqI2qVN16qhJr6ajoax8GX2lDpImAUp5B9evOV3PhA5KUhwFwNQaufc
s20iM+pvBIHjYqBiK6Hw+A2eowboZq6DrXww/zapEcT2ZoA+BX06mOkFegtJP2wMnCJUiO9rdtEm
xGJY64JktkCIpq3Y8z7qgfmO9RX6KerwMRkYri89pam/6VASZb80M0j9k7hl86ophX+zKchnGmFF
92xZm/m9pA01ggUczMLQ/Vf/HAyAomIwbcLxiihr5xnnorJ3WiMkdJiGgrXn6EhHLchuAoLkJM1Q
Ec7KS9QoqgR8ApIRSAccyyXVJD6XmlRpEfZrRntsR8gu97QCcheS7zZcqS1etKqxnQN+wO88RHyb
Kli+4aVZrXKn4Zqea3ki0hDSQWgp/fOVuXSwP14Sy3yh52c0EEB9edAhROmO9E9a73KYlMXigXuL
7JPNffGl0MT7jbx3HcORcfvt0fjUHEjlS1+mZXQM9gl5xMNitIFnVlFBPi9NNZ/scHznX3QpK8hF
mtiRTsf3RbQWT9kF3RBfA/mfoMM1ggrhgz3pFTbnjtYxJxXM6fFhoH3q6IC1mhBvc4ygxrgXASUp
gMgZms7ph68RNsstayLkIvnU1VS+2tavCvqO1Ad4TsjjfwQvj+WizscNQya6ZRMs/a6p4dmvRRtd
XAfp4KhcAfcNPHk1MkElEVvFz448Eyyoa16durcp9Gtapo+ozVfnNMxOMv1OaSLF6HngtGLcGOMp
eKczb/Dw9oHUql0u2ICQVQ64XjYDufdiT7rWw/aZbyv6CUlTOTy1d3bDY/Jy55YrtvwDAlRMPORh
gqrhN7luyqQL7CddibaI/pZNtuuVi3qFZFnO0sY0MiStakd7aB7XepS83J1opugtTBHjp0p500X2
eG6ReAj9/lKig7DCBZ3+shjlY4drtrUIv8hEMvTgQUX7qnv4lwiwq/deDZ1Eux1V1T1Ih6PYX+iu
bILFnOfqzJTidGu2jdyMhalC2f3nx+fRWhjDzjHk6q7YwtDOjI6S5X6vI5iO1xk4Oaiiuf/ZZR6Z
qi8czaDYVBL0OhbbaRLRTQkikM+ZOnfrIllmP5HmAfXXKwJzXOT5qN5d17RyXlVQTeEz+ji/1gsI
JAZFKVjaR4+sCYZrWXJEuaPnVHrB4h/Cprh6bsGY1+w5fG/+pnvlYMv7PjB8Htn9z7XdILHcCl78
yzfLZw7u8DyQDn6HzxFRN83SH8WiPt9s3WC/vG027J/0xNidcjK+MvteG6EwEdz6iUbcebT3VTJe
2QEsg0LSKgTzcaV9JON1yD1layVxBHMa6OsY3eu27fBkW4llOUu/HBq/izzdMASaaIyzz3GZZSvy
pbAfd90l1O9m5LClsatuLXCXCK3GfNZA16f3YI9GTvB1iR3BRnOCrJ5lFXiL5oynl/lUV26Wb4e5
ztOTHiGyo+2XMGF1ibECWbcl/grESS1VWKa7Xi4DgQ85n9cPWc84p9bYxXwKKJgojXVg0SOUphPA
7KDrnzumR1T1sibGIHI5sGXwHfj0FJ3J2U6rWnv3xsiSKaQHzUV/Le51mmg2bMGbCvPFkp4YYCws
Q5JLUhgmY7b0/kN4J/5RR9KOCD1blGOecIf+RL7ED2+n/oLXE2jkGcsaaHYo9ufXFtNK8vA4AbBC
gpSyI6hzChF1+b4O0yvT1Aig8Jtr2TIVTLlaE/NqAlfnltkze+z8yISt0AcFGV0lCMZ57zUtcpzd
KnVvc7ahzl9dNPNF0GzJ3quZz0TjCVWst77B6OAqOpSU0IyOzSEIramydWheRj3OBcMsyPl5IssI
N4QEjuZ4FmIZRkB0rf+nuZFLwgOouSCB3PjDUCWj1nGUrl/MgUxwS4C+GxDgBzNnZPL+x83AqFLM
LkU8pQE70CMo8vbxzTnrt/z1iGTyNtHPm3doyqX5tZHbKuy+l2vBAx7DP66CuvW+E827osiMcnD2
9G/i6+h/cdfiKnZeHpvQ1P/SH9hAUGKnC8/YIJ2tCNIBOeowfSYXXGqp7wTkyqRaeaGnmT5o2Nlt
YPKjcpDQsNmnigiovCP2y7CHY4PXQdKlsQ6hbVFXytbbVqyDEHNKs+XWFMeHB/Pi6X53i932sN9y
nTbVbDChNYnQ9BMLg7xl4nCVAXo0IDfxeaHU6/DqYxtgReKirYUjQ5tmIXls+QH+g9MNBseYj2+P
FkA7juEbc2gTydVBvVfM+OrnmD3HKtppe2u3Ibov7HbmLUtenZGbBpsyU65SiZTqQ508t+oZ5e8f
4dLCDI8k8HNRCFmJm8UqftRaYoFEv99Yx3ZjZmhISbRJq/OKiwQxXFPxWQqap3YXWzp9qwie1sC0
szFf0u74pXC9FOol4UJtu0gGsNnNTnTgUaegfVEmEmWCkmypzPR1BgidW971QqgzCaE0GNluGBvJ
BRy3WqjfMoEdXrS+6NBl28/hL4MIE6FhDCgeI/uOzJ1Eshr+UutsC5ZW43fQuD1qi/CF8vtWKc4d
TcOvV3KWGLRJ/eHnHUS/VV2ms9QqXReB/zOU3z56dSusg0K8HNRHhBh1FSeMrMmKVdfnEnS5nlCt
HrQ698LebrMlGxtYdr24OwBnWBr4lq1enqfwhv7jXasWnwBmZWozihxLV23UCICEE9/IkcRvqDqE
F/BvvdF+aGsldqk2UaxM9FCwq3TAV7Vse7jtkZjzaO12jq7Pad0n5itB4QY2p2fY3hIyjgKkuav9
gPvIryAcGnLtRGCNNQehma7k9aEwnskQOsq0uk71uqqm9j8uaE9B7NE/dWwbe3dfnFGQeIvYAlQR
VDtNgyt+tTN/xFQowxwx51un2+6GLLo5+ZbMLI304ugZQ7rMJu/+mZFzi7HFNPsPSY6CYETlRDux
+joTcFIRXihE/PQ04PessabHvmurQMpAfg1kwK9gEbTuM7A750I1P3eyS4WwbPQ7NgYJ1LiMZfi8
ZdztLdygeI8wWi/JcT4GElG2ROi955I3BrgfdJqTz30RlP+5ZU0CHhkB/t8NQZct4MadvOsssOv2
ePdebvHi4/FPl+zVBQsjOxSg7Zj7IAinZbnyETxEm7i9u786Jir/SAnTbLzqgditHsaDz4qYs+eX
5CUNIgX81GSJ5qX/CboEdv/e/y4Ib2s8Jvwqhn/AVhRi7+j38Xev+X1KbbQOBznZrCvZsbh62wIY
/JF9A3EcghkeUi2gM+NFSQtlhgjBXjZP/Vl3yYa13qb9TqpnvuSIuEP/pB87bQXXUyZUfWnkKqq0
a+yVWA/GrPvRoLrCsnxZJQbr4FxKTsfZ5/MEjNoXmVIPk3vnv1YQAsQifOUnQX+nFnLkEG/c92T2
4vxK72Mn3GkELE43abEp04uhu9kq7IuWksRwGVKcWuBW1z8UxaD4xhwc3nHTCVh5fYjC9bflsG5/
CWtLuJgC+pQL2S8iMwwpqkyXHnYk4F4SzFD0MJjUlVR+klyfg/eNHoYoX6d5MAJz+Qg3fxz2T6/8
/kLnDwZDIn9JIBEYUJ5mJuJY8rYxm4Wn10PL2ruu0oKSIiIOcOsV1RIYREVGRG1J+iIsNA0syUME
rp0FVqEGyvZY+RXUd+vBv8QXmm7BWj2ybfwPP5i5nmXB9fTMG01YvGN3hYiXJbKGI4mib+FP/hs9
22ytroZSWoev5QlShknPasDNFlKlOqSJFW2oAOc5pKoK/hiMvZNckFQcv5qzW5eC/NG5IYjBfMR8
eAbEWUYtGPfcN4ICabtdsM4EYHT533I5rq62Cj9UZwjUaNeTzdosZx7OYzqfkAFvjNEIeAleW586
mI2d3bNTDe2WFjm6FpOJ2tglTBkSesXtG7YDrOg/qvhOqRTYMAAr8PIgO5IGdZnwiFCK7SjYJ5nH
VNsy05ZS7YzRglE39WmFY4CzMJ30UhGW1x+QlsjLtugm3XdlmuWZ+iFDdSeE7oD2/9vuww3fDN54
uat7hn3rAmbtfuKqZLFumDFrUW/ERwXDaGDqtMjhUvtklB+PG52HiLmZLBUtQ5Ztj0xRs4dARZa5
yO/fpu4Lxm1AEIJtj4jf4lD2K6eIkVh5JBYHKvRRVrO72pqIXzKomvzB7tQQka39rTGqrOkS99zM
nsuju92tlsLB+IRl37OG8WHLzkQgMlRHGq0aPqAIwafXRWT4ofPcw04unqcp2Uzg6UyGa+00qvs1
PtizXdoB5vTA7Bc6ZlPfCT+1sQac6Jwv+W0RhW4Ieo9rej+W9pTmaZCFUrHA5Mr1Q7UlvEM2nbp3
7oGkftep9QzbSPNdXzUyiw125wLNa83AoY+Q1pStl6hyrfZcMS3vB8JQHbtPTG29XZma8zsaqSVZ
JWxp0TfqsPikNddAxcFIiHVdm6ISPE5myD8nm2iRps9EDr4wN8FURQay3GI4sngNve9IuD0U4HMz
ZGZSkaT1IhoV/rMFjaDOoQFuDgGMKaadG+qY7YO+QiwwwCEhS5ndc2gfw6zQKO28+46u+zQdsJYU
6UbytJeDfqmbc9zwvEW8e26aorAdEM88824YuaptHR9CdEpIiX8J0udw694Go5VNg8Mj2ag7Cj1O
QNNSmpgeDuF5NLgxmDVblBtGwar3K/4wCEO+VeN9nheWPb/rQMDYFwRpQHtEzzXC232H7bhO5YKt
bJVxqktmHH7NHFLH/Q3KlYzuzB4xZXdomX80+ZSqynFO3sfx4qOof+HmnMImc3DRhSuv8HyDMBkD
ojHQlurRuB1hjAYcT55B5EsRmOMDYeg752qG7SWKH9wAmrqLlG0Yinofd7KSiBXeLmi7CUg5KdqE
1lMhmWvPChXiBpzkibzhMVP7RbKfLXtSWjdOLDKSZSYpK9uTiVlYFKUMd7W/OaLNfEtDivFoZVP+
xhVsF2gjbDR2NOQah/wHqAH9lNwNiT10u0WV57XmybkUJRXL8rzVdiWwRhYFYpIfeyMFEfXb3CU7
rl78RNf+oUuPopK0qpztbZNDrwPI5PcVLztELDymhPb5Wgk3DteFAipjh9Jh8qPAT24OPgdwlQRe
Bbuo2ryTTnSIRWNAEwiEOMAcu5K0ByedszGST8JIAJHRWU0cVsrauvGgzPgvGxEvfGliwHyqOJdM
tX2NWxEkDGrQ3KLuq0x+EDw2ws+Pl4Um6ugzNVGp3idZMLcSebA6B5ujUeOibDpp/1TH7payhpA+
F15a/ypA6lu1CEtpy+d75OjN6wc2kjmkR6wbXQUDkjSzVV5XnIpt+qzBkWt1LEVh8s5YTqJZV7qk
6hgKIl3WfeonFL0GiylsBSddjjf49edUdc2Wf+cku3f1bUpaz0/ZFhxBlbE17MdAg4djOR4icOsh
2GVNv1uX9u7CfWWZd4fhwSzudeooYxvNdK4naQ1AQpykuqskXaLTjLdpYe67rQ7Ay/ZxrjdPZ1gc
a7HsNfO5gtYMhonDHnwo/87Nukm+b1sCJUnEz4BA63X8JteHiEz3SOcvt1+QWEkRNvVEiXqtQ2W4
fdW55LfRga3HtnCS/RaTgts7Yz/W1MzW4JnC+XFAam1WyugdUWj3C7R2jZeK0rcDUCox7pkq83LH
qW7aQvjVL+qiiaNZIoblT1RVvzgDnb3NOHG5e+Qgh0F+eHlJa3bhQcp629mlRlX++vEgQUuKwYj2
WKr8n+0ZnX9AhMW93Ujoz0yUVXcVVjBE7MBmFU64Upd/geG0iKYovzJmINLMjkeXAIgvEdDcqKtT
KIv8kmJsaFeydh10Oie1jivuHBUlDT7fS3iNBGKzefq6rKld89bdU+lbHhrAYbJM7gvQkMlg9eN2
UyvVF3Cxwthi+HFof9Pm+f+6pWWUzOHTdR29bRmEBNKijCOWw852SXwueX+za1UStXlZWVoob/7l
iXYHKbU6qagCRrl+HDN4ee9axxNEL0k+KEVMQv0HmKFxuSWkrpGtBHci8HqX8fClxDuzoQL9QRH6
uqEDlB4Pd3csvLlMtJe1FjSHcPqR9Q+MUrkrLmVzRcomSQ7U5E9jomxq2heGB2WILm3jwSliskRQ
7u1xHfwDXcgrQ8hJfHDq2ia8saPQJ+220GBXXit8GYE+VD+zw9Lbihh2j7uddlXSpR4Dlz3O94KU
P8NRI3pwKatK2nCrcuXVVpME5MVumIaR3bWRTvKbGfn0sD2HK1+RLmNwSVGBjbb576wqrXiQLaFc
vANBX/h7uW1AoRtPLapMTQ==
`protect end_protected
