XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}SΣC�U��0�H絢h�lεP1�M�fH\�X����'>^r��l�w�Qׯ�S�2��r�_A�����X$��L:s�rc��f�i�˦W�iڦ<4ˣB��F��}w'e�'B��f���Dh~B��z����e`��D,I�c�d9�[N)�-��k:o���Y��O_=X��U^K��M�x�M����TV��]�Tfi�u9|�-��m�|P2+ԃi��'�&�|Hχ��ġC�ڗ���3Ң'��z�C�0��5�������pD>ם`�5MOfJ��faZ�<2o�7Oj ��i���������X#�U��f��Q�C;p���l�QB������U�d��� �K�d�7���S"!G��y訷	7���o��uW��߈��"n���09ǀĳ�pZ��.g�Aj%!�xWC�9�>�<-?N�D��\"�4Ź��MS6�c��kҷ� L���-�b],]�nw�3����H#�9�褓@�5-���+$5�>����p+�en���fa䏦�l�yqB�}���"�v��Вws���"*��h��Z����RȮ�gTC��{)���Y-�:�߼r˩ǭ��?6���TH��/�޲yS��Nh�Q�w�� Q+p�Ь�'�h�KX�c��r��w\L�S�D�-��4nd���7�ЖoD.�ˋNh�l�A�%P .��n��>��an���Vpa�X�mҾ5��/�V�2��b����Ĳ9Sõ���C�ʬس�`H'8E?�XlxVHYEB     400     210jkV�,�sS��������9
�p��cJ-U=�K�$7$-����W;�;`�Pxy˳��h1 -�+�q�7��e��J�1����vs��ϣ�у�*J���F"��}�eJ֏����r@6?�6��,���2L�(��!���%q��N��hc��Yq�w���k�yۢAv8�c���0V�{�KS�6T/J+��~���'�7�x����ؚ�ڸƈE��gbMgYP8c��1W��z���,N>����,�K��Qj���r	������IE)��V�W:ex.�{�.CıD�D��B$
'T���>�a9��"��r{�A^��$���m�q�J6"ֆbK13����*�o�
xJ�=����;�I���(��*WwCJM
hE:���C�ܹ�r�*����d���2��R�
��kί��NV�;h�(s�h�� �� ��B�p�3Hߥ�M�����HĮM��8�X bV�,�۟H]�<g��jsʢH��=�S�Q�y�F:"���XlxVHYEB     400     100�+���~�>ύ�؃�xG&��?G埕IR�����u
@v@;�s�QC�e�2ݞ�&ˆO;��,�Ƚ��T�ދ�r�z%�Gt�g� /q�Ԗ?�ka����K��CH���
�?"�*B^�e'������K�h�@�
��f�^�[���eE
(�-��#� �渧���~e�Y���<�%-X�i�Cg�˘;�r%�E� ��gO��>���+)����!v�/���3�Ъ�Zͦ}O�[�,�`i�7���t�	XlxVHYEB     400     1f0�QP�-��*�::��l��P��
v�İ����?�{�p�z��Iƿ���;H�&�2�QJ�y��,ӛV�6K]�M,ԃ3�|�����ZO#M3-�V,}��Ϭ���0�B�k���ߩi�ٴH��?� �1�GSGj�qho�Տ����y��~�q�V���g�+PQKA���`���3���ө�C%���;�}n[���9�Ү���9񪞫����_sM>��$$��W�!� o�����f��ozt�f�;�
'N�D̵�.Z���j�F�CJ1k��T����h_09$��N١6��y��,�(��9����z�=7՟SI/� �y�rb�ϻ��Ȟ�%�-W��kY[����&���x �!�$䅕��,�����!I�d��.�G�][? E���<��th�h���t�����Sd�̅^[R���(&i���^��eaA����A}�b����!7�)�퍪�]��� �h@]mq\]ʁ�XlxVHYEB     400     230չ�1�f�9�&�_O)l�`իK��N�%��#��?ȟ�5d_��A�R���:J��*���G��]y���	Mu����1���T��^���|)a[��i���6?�玴^�'5�L�"{ a��O�Ɍ����iP}[���	�Z-��$X��-���C��A�n����*�ۿ�|'����� QS�%��d�P3R�Xԋf�:$d�F�{b���r�E^�bH�wAWf�h�Q�p���QZ�*����_V��"�.�Z�	e~�̮%$'��ou��2��vÞ�c�BS8��^�4�a�1k��z�	i��z�k�?�3�QL�:�o� �YQ�]1WjږmwX�M��^Քj�*ҭ0\��h4��		�~|�c�h��u����t��[���ںF��K�1��F�\I�����Ap� ��Z>)n�/H��˝�Ӱ1o1*�S%>�aSn��~7��B���z�ճM��N_��X��{z���5��z����K!�"
�;^jM�>���l����p���>Þ�W���͍WI�ruhK\KXlxVHYEB     400     1a0,�@[�џz�/f�:��m �vX��L�2_K���Q-�A��Pw�+��@ukiyA���ߟ�иo�+OY>L�&\��^Xh�uK������~��3�;8k�9���F��4b�_�~	����Q�>��h������9��2a�}4��p"\��%K\���v���bc͙Y��E�u8NS[�׳���p��}��,[<D1k�`�CInV�)T��́��E��$-^��E�%����>��IA�Tkj���� u� �n���7p����\-<,�+A�t�����9ż��=qa*0���OCxU#�T��NZ�Q\��Z�!�a��L2�
\X�8��GG(fsB��E�h��hBN��:�Ӛ(Z^3�8	���ehQN�u�v�'��bL��Y�I�d��ZC`���������XlxVHYEB     400     1a0�1`d|I~����Zz���jv�#�,�f��Z�4w��hE_�p���y���( ~qݐ���:/�s��m��j)D�*����=j��=/�� o�����#`%nZ�R���Ò�Q�G6���{>5ط�"6s�r�K����6���C�f�X���˜�dNaL�����Y-o1��S�0�T�^^��s<�_���0�4�AN tB߁۲�y�<�̃<�D�@�)�wנK%4�@&C�95�Y^k{Ƅ�<�By�|$�-Z�:W�4D�ᢷ�tE"'�]A�5ґ�Z�J�����B$�5P����������6��d�G��隵c�o�kj�cڰ������b+�
���f#=r��]�cٝa���j�[���{�8��Z�]�:��#�#J���A_h� cp_�
�u�
��bbjXlxVHYEB     400     1d0��8�@j]o�	1�P����h�7݉~�u�X����	�\�#���wya �V�I��Vi׿�Á�L�LXB�@���֤8A��b[�5(b�3���h�a�Nmo�Gظ=W�b�Ȃs9:l�wޏ`��Q�b2�R������3g�>��9vd=��!�^��د��i�����o~����H[����dJSw.�5 2�ч�{�� �A�=y�zj}P������Ц������$�s ,�g��U���Ew�:ppI_�6��Vg��Cb<4	[3@PY-�3���#��-ygBP�k�o'��9�9;f|�.+�f���J��L��L�c(���wlE)�ܴ�B��v����Vr�t'���6��g@�4:�޷A=a�d�Oҳ�wWHiZc��` ��e�1V3Ԍ�.�?��5w��r�A��� ^���~�f�zM����q�����K�c��q1�L~�@XlxVHYEB     400     170�W~,߇�F=d7=IʯȒٰצ���#;���C�2�2:4{ng�7�u$�.9L�@(Ԥ��*~�o�}���p���2��ͬ��oi�*i�^��z ��`��Cp��SwξT[p��R!0��(bM��s�sL�^�	�O�1Zj�T Ru���TC�7�A)�pΆ	�3ϒ��*�8�H�]>��vO۩A{T�y��\����U�8]� ��!J���;~�~�x"`�,�o$����&��-^Gby�c���yB}��j��E��#��F �m�p��'�������X��_� y.�-�VTԯ��D0���W;�i��6�y�7�R�N�4T>L�`ǅ��&Ĩ�~�BY�m�Y��P92$}XlxVHYEB     400     1c0~��^��2�F�.�>p�S�hC��쒅̴��R�U���-8v�2�'��Io��76ʍs[F��t��+'���:�A��Z��� 1�-����V��3�ߦ�P�b�J�N�F���WeA�"���B?���2@��Y����l��uΡ��(�#�I1��M�NE�K�����*k�{��[Ȼ�TJ��'�
�5X�6����+(8\+��$��R��*k�q��$��U=a����n�w�9�l�M�	xN�9W�w�d��1�I>�$nnmP��	kȆ_��}@��+J�d=�,R��G�Y"����5�QFLK�O�M�C4����%�5�!b��bHER�\��$�4���/�5�.F�aדr�U��O��Pl������H�&��+�oP$�:-`4�����aH�ef�*/@q����mKバ�nf������I�0;P���}�߇t�XlxVHYEB     400     1a0��c8��z�^o�Ѷ=�v��alE]	`�w�Vl�.-��TL�ڀ�%m㩷�k��W��A!+�_e�2��/2M�YԾ�#���ǧ�a�T�'��)qr���ۙߦ*q!�t,	cօaYL:4�p�>�6�f��������H��@-�y!��]_8��D��2;φ�َ!R���U?��� �����2t�d�H��^�@V��օ]��+�*!.EV�u��]7ly3�}kf0�E	�O��#�ۚM��(��,�B{�3LA0SB_M���N��2�~�nީ�O����`-JN59������8����.���V�?	U�"��#q34�խ��2�6A��X'�C�*KQ)�����x���#j�F��A��.)�F�*���;�3�~�����f
z�Nˬ�Ȕ?�a[��M�R�XlxVHYEB     400     140���i�)�أF!��A��	�?k$^`��`Ê���c��H3<펧"��,=�c��l��y��U�n=䘥�s�o���YC��ӁwǬ�56dU��"��V1�2iF�Q)����W~�h�}c�,������F�)��K%v��zǜ//��q@��̜03e�6C������~�+�,L��Ƞ��v	ԯ��Ѐ�78{;vj�;\�S<�|�h���[p���R��a�VA�	eW���y��(;q�|Zl}��y���f^���vSk�v����AU9�RxY`�b0�P���R@��1���jnT(�M]�I�s�o��i�XlxVHYEB     38a     180�ʱ�+M�0Ё��܅���(1����$؜��7 �!�R������~��	E#���5�~0k���Tڵ;�z���"�2K<Ȝ�|�Lb����*�{a�$���+��o���ɇ����^gd�>�v����e��GꮣWe��nn�m��' ��VծKQCI��E�U�����Ɖ�h������#�/�#(٧������k2s~ E!��a}߼O·����u��|/�Zf0M���^chf�T��:-�\���oEJS����^�[�&��[/��j��&dO��i������ny�����ϻ�qʛ����� �l��OLk�
��ABR�3�A�C 䔄�0��f���y� S�vGƔu��0�N�MՅ��