`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
jJ3BUdnVVfGIN4GgwGpmIb1xbQSTglypuGZoKt4Azj8pMQJMIxIAkKCoQ/2jeJiIec376dN8F7BP
Z9tAx85Z756Byrq4XRD8vfbj/HlW3XdwD+CK3FC5SqeIyVIlh5lP5jpt6dqtPlz052fm0KoOBg4h
8zM87Po4tUZhW+VFyw2MU8GSzfwLewBGSzCKYctF6KIfEorwn/RFY+DWtkqQfoRGqOjyf9OWQetx
0dsG2N+yhQ7sbey/Cb1lIaTjhvNi/oHURLlHn7FvrxSW71g0mm7W6f7k+JLPug8gUSwmKhzI72V8
3Fo26gOynAznBsFrVUN/DFvoqNjeEWibhIO3dw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="p7SrWziqPrJxd2K4/cHm0TN7earhq/aC8UiHeGAI1Ks="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17872)
`protect data_block
WPyF0yxN+QFRLudGzLvPHHzi2MEM3fQconZeBIljOsVv/8IMbMbvPMfL+P+pVQY9YV3L047x0om2
m6SAqTfAS4L5pIX19ChCvUnu4rfso+yd2xFP0z9DwpzwwtkcSZVed5MXmOcHiUIeNETyNstnF+MQ
qK6W1m6XKRVJKRfIhS+r0PKt2fGzkONMI+B2XBKtUCZWaZQZW2p2xvIUMQLFvRQkf26nVT06ZtNB
KqHknRoLivm8butxShFTUeAEInf4TWfqHYUSXK/S/5onQwujJQ9sN9h2nLQQVxB0rMhG44cDPqiC
yPOoIXvqYXaphZukB+OS4Rb5ZIASkzoNvrcr/spMHDE/Xvjy9ZG93DvLEY2hJ9CsJGRWDQyTuPTw
qBaR8YcnT67b9sHut/mezEm/NRPkviXH42hBnlmVBbNbsY3OWwRTEKI9t8xJBrWz5Bu0rboA8zNX
EyDMiASorfJfL0FSSI8KII7ON5Lc1ahFXrb97HT+SYv5expZ/U3gb1C144tTHin9QTHWRjIQPAGt
kJRvwH262BDyroI528MTgw0pYAlr0/ZIhA0XG0sNS46X8K0ajJ78EUD8NmN+66plzWcYN7p8eLyo
lLNLzhQcxzg5Nma3V998+BXmKVD/6QiONgK9dCmGQN/igg0nMM/Inc26+0DBi9H2vtl8G2spHKfX
6V0aY5nOTbx2/YdN8vlG801L0tHPcERCdGFU8+VK/gX2kGqkNXxo9dOLx6ix+5cm1IY3X7+peocx
Puq8V8YPKs15/MDpuSc4+ar7mQLF8HTzk1HCd3xq7l9dPMExQeiacNN8srsGVgpPMwtJjIonLOhL
RBFvwd6Y86txpw4O9pLBf/rMr8YtwVw2W0omiqP97GsAGXHODQSvSp4it0bGxT/K+c6/xA51e179
ijon75NkPbUOmi0GdkXGNy/UeW5q6L5UaxromjL5IVHk7d/+aZGc7HbTq8c3sgDeN4pexfwxAyke
qUcShF4Xhfr+HQJoTxUClxYgD/dKaUXuimJbU6a8xG4yFBucyMoMJMzfgxg+EylFZeIyc2QJ89eQ
fGpbq5c5sh+Vb/fXknZoKUD1fgoZB0nTdX2wRf0B/esA3UgpqQf2WGn0UXxvDg5oPvhl00BmX9h0
G+9VAOi4qIP3XgDdqIgWCL7/yEATB2PQ3oiQPD0D8yKPpOr2uMzSzH9v4fmKO8C2fhOQy6ts1o5I
ofaoiVsMRsLJmZvCRIVJMuyIh0SvrWRby00SMhu/PxNaJRcr6t4aUOpF344ic/ud7FSpmDuSmLL3
UBsbJdm1cjelp/r093rJ28ZZGNUh4nzj0+hPPaOebi/dT5jtGi+2hjvR6hsFhrSoqPAXaWr7/cWO
2qYCl2sCPF7JxT81Osnu0ab6m0Z1b2vTkILLukau1D7KMv3fIm6giMMN3POA8IbVJcoZ7C6Isf7z
seZO3slhCalow6pdjxwU9vpw2b3dKy8QmES8alJaIZd8kWCp8Mifl1iOrtI9F9KHGIO+YL6MvBgj
X7jpHNEkQW7C7uKs2EmXNuTqGq41FqOfZzpntot17hlRLf9sVyPSAjpEOYI5IPrzSefzgGAW3XFR
3mXdFkLTTKBkhJ0+o1Pa1B+sotQwKIcCa7Hcvwf2a0fJdpgq7TCecj/aEHVbmMrNhAfEKnqCNC4w
H+0KffyQ551Iuj/A4nU9wp17j8AebiWqVaXzgKril6kPddFMfhXcFRrhRJ0IYrBr8LZfuBRQDubf
/nJasYFvhOkARMa7L4LYuJDE1KlD16+9FtNRvHN9F6ndu3cMgmE9o66y8F72UiMM+iV5LPbFoA2v
i9le+f9QOz7x929uOYlcDAOY6Ne0s6X0zAy3JbeJukMbPY3bpwgldKd4kvPJZHVvwWyLo3wSWuHj
7Zq/7c9vQkF2zX1tVndCHCNGgmVUhEW87pJToxpY4l4KJLvgrhPLciN++hpMJqCRVpCKRKOU14iA
zJzb2xtfYAqwUZJspm+F82xL8NC3ZDvzTjZTlMCyIXuDU6KFu9d/nA61a04dvUCVr+3Bj/Jqaj+O
efxIl3HGBA1FYLxF9cWeQcNum5vrLde2ZRwO9wRXYkdzQzbQ3UC4BhwCYEGeGYYdTZYxV5+/QOUV
0KAoEwhLHvwzfhvxNhxPPylg4SFXRDgcgCedWpiWcexfooNpKZFlpBtPSxonchlPxITN2EKYapwd
lkHsPz7lhpxVgdl/Tc5Ib09YuM2Pct52hYPN2juMqxSVWBuZ9U9V7oEeNKocPGUgdYR55v0ouNDd
9ac7PWnqTwU+cS5sv6bc+Rc09D5yJXJPsMpcLmj86JV/LvQLV5K/QOhpGkxiBpRXLNMnvxT2u2+Y
n0m64MecMrqHf4OyOZhD6LCi7ECMr6sNmq95E+xwqvuJTQyIP/3vKyAP1WFsXbgQMZ9i0ZK3F2Xs
MoA47y4E8l2oQ7XZGZJjXBsB4efzUaltKNvRJ+p/LyrYkCXKpZtWE/0AgkStpbN/TLmTt7Ges6bX
3IBXvsEEo599DyBIjOMIKLvA23ZnGr2tz1vnZJ+sajwbUC9+g8fwb85UwwHGcTCTnEkEOmXWlx64
mvuTIN1XWZ++In3Z5AtG4oQHjWLjISIj+oeeOeZjUDCimA91vAGk4NurOe62TZH/Vb+czEP82gWa
bYlcjL1ZmgXNk43M2e82Pljrtxm9D7xji1kTs/V7j/b84ZnnpUjx2mKr+U9/52Kavhl1pAt+3l1E
KwBqjtot8A5+RK3k/Ovj9qoRdq+QSztPuDFaVXG//ycFsbX2fcEMNBbqQgnHBYVLnvmLVy9s3zP4
rYjA6oTGeMjkyR/35VdmE0+zZVALdMYKuohY9kxkiCx2JUXFLzjRjcl/oCklUpinaNxOrBuOCBoI
t//YaEHu4Gxb/WWdqynqoQXE3TMhvwnoGhip82GAH9auNtQO3vMmO29s275r7q5iWgj4v09UTua0
MPvsCQPe6lYG9MZyxV/TDYd6OK33W/VrnsggLQfASjrDVHV1/HiFicYM5pD7vzQ/yDV0Fh2Ou2sA
fO8eib7P2vb9LI1TAK62an5D7ZSYgXkJEZuL0NutOfaE0nh7M/CEY3r6tZbDu5fcy3HmR3hN57Q1
15UNhLAbT/EgDynwtFpeRUUi6u5eTy3VS2+wPsz8L3nzdNoSvB0kpoQkCBjBo6/xwdFMz3uUQ0gK
QJCVvvD/pcf2b+zDqdm8nA3nyzy9ilDCjQ+dAZC0SYw0d9HEsAxl1OloLMylqikKahI9qjmFPxbD
DF1Msejkb8EhQhszBJ46Tj9ko8ji2DF7AVPJcVMLuZpjEmbnDzWFMw9hdpJ2Fbclrf1hwH7BNDkL
LRWF+yjw8EXIurk0xOPknWSvK4w4TgKGKzFdohS8vK1cYqReDIifLvOSnyBVmftHo0GF+FmmKzrX
Hi6shGJbFEO2NXSgyCISru7TgQVpik+o0WnzbfS+bBb4VImuoIq9Pdr9YFdQAoMtPaCOfpRp00IY
qv5GC7wW7h44exog0vLehFaht4LYupVTkYqDwh1vJW8LtomSwAPHNl72ku4mtuQnEdr6Cww19mnh
6d4CUWNe2abpoxTf+XvyltZQeY/MZUhEBL39dLS9+N+jJgnWGfdS9wu5H3TC9AkTToglO9Cpo47K
nqt5PchH6R+PtNbo324Jcek8i9nPQTrF0mfzs2n+5DOW8SQTNep7EnxpqfeK7b8/1fnm2h0QXuzD
5Mi2QeEewCi3kP4WkyehL3iFT7uKEVfU/wTi0wR+RX9+bU7fTmzX7yZIo2mjBVsRnteDB/HZ7StG
x65+hplFNrn5Ui9Txa6vlTVYxy0oJXfu44bdYq5LQdVEdUy5Es5Br/OcTTC6akMEI9ctR1YNfUl0
LoKnMOSApppmdBpDFufolL7SdcdncB3QX0c4UbusMjAfIrh9c67e9/M+KiwmRCC/h9BPNa6fc2A9
VtauH2U7POyvX8uapfCwfNIf1nHr+5bpBCZapHTwo98hFXobIz6aAtm9z9SMntiU9aeI4VGqLuBW
8ENv/rSFTckVggmkAqQ4O3MuakAXFJw1N+2W+hdg/+pHDNjUYfwCL+nFsFywMhyXNlyymAJjB9Bp
TDhugUtzfrVSKPSvbMiL3XwicBhO9q0HBSBMTSiIkhMBqCcN0RWoE3t2iAtXbSWfXRMcFR1njbWd
OoRPf9ONSEYbG0lSh7XTcrOVbDsEGeDZE9qYrlvAsQVBy0wYlzqEXaL0byT5KwEgpBSmVF8yzLs6
hhV4Yf7aFPRuIHIP+D0HuxH7IwyC77fzxT3UGl3IdG1R2u3kcc499u/ME2B/PiU/cxN8REup+P0U
xAu6MDvkPa9YtRnSQHTaORc+MOVzKVmNxq2qzdOawOagWg+KmfsGLGxJGF/HrG2EepKGa8oyQNTt
cLTSKyZ4l1YKZwLfawN0StSSh9IyJPYf1SM1uuh/GEkoFHG/c2zaiyExuvfp+5TTO882iwqBs97J
bh6f1bMz5ZPLGQ07PR8JmonenSJ+FfZmeROkrzf2AzsTeCEXTf+NyEgr3sqtWilf4zt9+OUV+gPA
IOm7PHwwk9JY6hVUriZ1qNgRlSgqMQSa08v+wVIAVUxCFFoGgMo36ZlmTJA38EmaqvMdl+x6f5/q
loohOe0iwz0j9NDwibXw7Sm/MM6CKUshbhsKkTlLTryxbBFotoJL0Az2XgyAK4M3yn7OVZ6rUKva
t4INtKRIl8IdIE8zJHYOzvjtkLGnO4AtmdFm3t2th/iP3fWjGd9uCpulLHjST+V4KKj1OrxTojKI
yCFEn0mib8h//U+PvOvhMXwNQe6cUwGcWKB+T7PRmwqJGmDRR4SM9VAcsR17eUqQmkmJ3i5yI5F+
yWhaqJuABcHYcTEwlZSxKgG1Ko4ECuBNbjtbKndzwjzOr3Z09sdplIxI1OgslTt78uc3Yc8UErKY
Zphxb0FIAQw4Dk+Gjpz2PXyI0vsuR7i9teqWiUItGeRMK3G10qoOBPNwdMLzT/H25wCyC4/7fupB
deB0vPfvjQOAUBNObYAmgAEbdO8mPL887ia9pnHfYESMTDWq4uqyT3F1McFXy6CvfhRJQLIbLYi6
FE74pAJ4H844ZgdEJkJ/zrllLk9xecVKGuTukVZLsOlBTUpRBwWKBwm0iklqBbJE8Ih8ZbW9sSu7
F3NP3RksuD8LFYpXlrMF3W7qx8rtHhJs1TUgxz00s5Gyx1v24xvi58ZeLeS+wM4B1uk38zNjqyyN
cbeFutxZ/ajy5J5Mf+mxjTG60exrI/cmz+blRaoyuLkNuyO5JDu+sIDbbJo1jzuFev7rGjQfOaLI
RM6PnVX+s8hjl0+dcj08OZAJclHg+w1Z469mXkmXmbW49CI+sEQtFKKrx86hCZIVAmCmRktCP/cg
S6AzA05Xl88zZUbpA4hOHW8BsiozDI7EvzzWLkT/ZEG2m+T2Nnfo+M3EWAuxkmRjpw8pImQYifFe
3jvR5VpKTLaiUiDfBo6LvCyBa6MnQriuBNRf1RXI8cVAZADH5QpiyFH3kW42DPB89GF8R6NEjBCW
SjVNcEiqMLB9jVS5bhjK+kgcvWaQq8xD80SqJqwPnE/sHiKoA1cdqrnW2PIcBlcjfRpoj8xXVZTo
MXwfXyUUEII6U8g7wh5nu4mfy3+O88F6brEiJL8P5Swl1MKQS3NL4l7XuDTFpcFIl+aQ61HX3DKr
7OPq/oTQvkyzhf7hHxQcyShQBTSDufQCDBjuaxczCjtvfAe7r6DTTTr1higDBIehw2Nc2t60WEpr
EuGks+/72l3X2TSOBWVS+wF4c7A9sKGrM3YNuJ+4r1KMKgy90Kvsxq5ApQwSNssFZrvOToG8mxgZ
4Qg8mnXhk9rzxKrSda23fRL+8xKCOF+/9uumRJ8PA65p1dM209CcvA9G+p8TNfGcI0nAE8tzSRpV
NJiLybXlQjfzYcwY2Hqz/72pjmFs1yxnkbipiDEIIYcJf4OF/xCQhw/nU5qTO+krcQ7BNrnaZr9J
Qa3HMOSf1/ozbMwFlFujNZe1NZT2diIn0BclExhTDHXPj40+T68SK/LLTun5MJqsNm0StE98FZ4E
ysFNQuoa4PrbI9C0/b12qoqwOXbJwAjeLUGQHXLDlqyimYh1vD1fpRyuFMMUv4yHlegubw1WiLsA
gtj3jjBDytwSR5tz2cdT7sW0+WdPPFjcdNhnoMDd5e4eHur6wwIyx5v/1YbaqXncswYZCDR+go6N
uB1G6tWyAnn9idwGDZjchzKHuJ6Hn3UPV1saFCmXA9DLn1lqSoBuFXaYO/cNrQii4rvBoABoW5cX
EF/6TxasUlSmCX7UB8pi6cBeVjEepoCIoCKArVfcbxoJGgwR3UiDxl0OSkfAd9N0mY1CSmhmPyrK
zhU5kMMTL+2thJP9RA4eCQJV4q0u09YUUeLhvuoJUDLB3oR3mfZuwBHaeWQMBWMSd3q8wPkKbo6P
PX4RcRXoY9V3rv2e6GrCpP7zBA8NZUmHT4ap8yijIC7cyN6f73sajiCe7qmvjKtRL6f2VV7io0GI
MnODuYK83c+eNila81s9KL/NcGZ7apQt7XcV7NteZ+8+Rju8tgHFJJ47yIzlYG2GKRbJlFGVmowX
j+itJIE/Mk+a5WEWWeCeitt3ZtP7Bcg7P4K1KPySsFnh23Jpm9d9KpSO0ebHNujkv8EfRWyQmXYd
D76Z555vv6X52kV3PSoEM2UGBUblqI9mYA/9xpgVfS8shaaLb2S3O59isAJRCOcnmE4nCeF859qO
DcmrXcAbLBGY9evWB1wMpCObVj4x8swOn+7Is0l9DiHQhQBtcMrREycrl9twlm6+C3SsajPlIwIH
YVcRGTTQYbmpN82ff7ROpwezTgxLoczLfq5chSHaUfNUOcQ7xkniRYQrY+r/fcK6OeHgEhvToMb1
CBykYeu0nudT2yQZBq80qNWjuYkJxhN0otCCHpYu0EsuKT6eaLQ2mS8xESf5oXv5bXro2gVDMUc8
TD5OtHAD40omM/IU62oEPB1DGHeke3qLBXEyXcb9Nr3HYK7LPUj0KronMtmiJTSJCRqmn5Nxg272
EmIDz8K1Rqo7FdI5i9F9hTR0KJbzY1jXZKBfeQYEjCtTf4U1/ba/wLqVb48MA7NlytvgOpgMF68G
UFou2iGYE79CpgiKzB6csGfWZveZN7wS7grkdKD8LlApqHW5LnrhlKd/svKtueBLhXKwP+VIQ3CP
J6j/JHv9AuxfkgFYO9QoXAKJlABQj1mr2WG8wkPFaDTs9svnharPnWGMRYDcJGge3/CT+46TWQlt
/AV2ldwKQRrqpMdFkGN6Hx44sWuf60S1Yu1yF1a7N69Fz5NPAQfPjmDXwUfwNcC5eyt/RFa0YTPB
nyI0WlW72K41udtVOP2/mLNTVIytzf8LxhzfUs0+Dj4cD/Wwd7IyRNYJa0RxJisUD5OEvOnDN75q
qm60Wvt+Uj03BBCRuAGAVSbUJJ6xAFQ4j8FIVD4fl0hmQpZBJEO+Lv5LdXrlEMx2ew4HXmOE9GBQ
LBlBJoUOY4UtEDUcYPbLSqIkaIdj8wJguspJ67MC550FQ+NaznfRdVrFaVqqJq6v7e+LXnOueKn+
c/IgwcrB1dnYUPoqhfFmIByXxBnqhJITOMY34TTJTObndpq8r1uOw8MWfckb2p1CoHGfgTBEcKUr
xel3WjB4sas+TD7UQbV8R7q42zaa2x2898AwLcBWkr20GnPtELna8LcXpr7OptwsF0SK/oBxmq6Z
+Yhma0KHe20DPFGbHo4Ip3B41Q6pLHWD4sRcw/l+Ds1zl3souiMsujPeyMWQwK6d0ZF8r/7S+x+E
m1cQmLxO+sIoKQ5CPL0GBcDgckM4mvBmxe0Ewx8F1MfWnIjrp08nKcCid7emrQNcR//m2rMOswrx
/lUqM1iNRAEWdBEUzcF5kwRYkwWJQcXlssOuD7fMatOGVOze7NPPNRAFTN20oiZiFQYRMvhRYvkM
g6HjbJieDSGK7fj11i6Ngat0v011QAfXYTBKZxf6IpL+nro3dwDx86wzZB/AJag6kYkGTKV2VY9t
66QhzGhTyv8kT3inulK9DM0MFMblMH7K3WrANXWJiUz3+MpxK1mRGa5MzQWUjZtgxrQAWPxP4saJ
MguX77e0MDTWywcnYEvB4AfHWWvVjTZxIbCwYVsLM8PGKSdW90ilHTViKkczyjsIQfn/OCKTfeOJ
pod6DdymtjI2qp5OscRyDZoPQofBqBMFjk2A6nLHkmABIRMC7Dvp1+2M6BTpT7L2GMIbcptormjq
miZKF2hrPpwOh8A281M345AVXigshyWkcmAJwzUQJEo7LrKRiOEP9ce7/0L4xHzlBzcdSXMzJYrO
Zsk2og9lak/FPSQ1SJE+eck9ZqoUFL+lL1FCy0f3DmsTs2IDGUAc9qU7VXm1YRWGZQqMWbBa7goH
jujHMdPMJG303k0Esuw4eOz8WhsAdvKv1FgHrB/Ldli8NiMRBpmaxzFeYGd1WpWuEOejxFYvRKqh
7Xpn+EKklwWtTdMzKwfh+ZI0GqJipdIj0PRiyRt9jzSeZp7hbw6v77E8gzYEbKfVQFeAjjlhGDrI
SRA/lacS2cCTqWtryF74ssUkgOBqK2vFlOImtOVlvr4fF+vHZ9MRblSdVpucBs6puwjs8k00eCAm
mqFUmHb8O++kizo3lef1i/oE/UV2zIqhpVgsSjfEmrlp5xVRq532qEI5EqH4TcMgPjEYOtkV4u3j
KHZVu1Y13cLqkGiQi2/mJ5/QoFAeEhZse5Mn/lef+M96+NiLYzExonZeBhreq7BQKGJ57h8Vvb3w
1PbFjSSkC5gfMdDIoy0dDJ9uNTmg4UUrtUsx/wt5dc746bJ+09zKrhy0TJ0LMse5+0OY+E9Wx7gT
KTBzo90feK7YfHHvNN/HsxECZBL9qWiODr9In42zzu/xoOmo1EXcXWTECWKxC8LHTsvSVAj7qMBE
f67PZo0mInsxpqc1qPP2leJqnCfHgM2I50zD7434xgPkcgMLILmsOJH6ieEXRoClvphGP4A4r7WT
7xuTDXnqklCRiVdCrKcyyUvwcoS9hrr6OTe55v7Q9//3xn+xULrOXhvAtBXPErd6bJvmgVY1Y3th
oc3Z7U24TMbp0UGvBq/q86DSF97GXShlUtf22MBp03U19yXlYPQarEVBGEp+1OjXfGQkk1aR4GAT
ylDUiqt7CEBJ4biJ7rlYwphCMPLSAMNRKyt+Auln50Cm9HBgZrOMDU1aa9SIZsYLTofnT4aAG+Yp
cwozxzuKLi1OMdhV4Hnr9ZEFKDJPsdFWj6qf0wrJQ+XnftXaXhogR8TQJ7qBBKpwpdwTOQQzys2L
583ocpt9TUkjL6Bp9Ojh82YowzGVDdLraA6apliZcUGBtMupc2JSVjUgirjMamyNCiyO3zjAejpl
2i7MRJqAatA838H9ZJzmECTRrOatMoVPlQsExhLJ1FJtnDUJd1FRkvAnivQ4pudr5Um+IrOcGa8P
ckUzxUH/ZJ+r6gQ8lrPGgspC9dc6sVnuXhkPa3GBfleo6ZOi4kMt5Fb6DmO4eGuWc8X8xjZRqthx
zC8NXdnHMYwWWfDImFI0hWCzKfhzIHJI/aaQ63jOmaORLVr2y65IfLYTJ5+4gPoyAAz8JqGYKEHg
PIr4EvE6BLHzeaRCpJR5EXhpIRi7gaXeDDobTBY7g+nJb2nYwPYQ1NKtkx0tZ3vtdEqiDq2DZ2/0
j1V9/XFJoYRRc6xfF/sIFwW5XKg6dKaKYbC7DDMGU2FbPtuPI5h3RuHEZ9vHwKpZ0b6n+IYVgQ/b
xUcDyc5fEzx4OhFLfBPVPUF97r4Y3KlezlhRdI7kYJyV8oqf9O86tf3QuC+kChRJthOYgjsXLEWl
BHUXop6QaWEMuepuosgP6wFGw3MS8FsgINGuqW6x2EXukjSvuUuOIXbMPq6mffAHi3O4nMkf/Ftn
wCQkH1j71ZZ3E8RJICQasX6EpJ0c4KS5yPmIf+ry3ayuXpDOxA0OurgMIfZccFLkmOIrYqkJWeI8
WhP6ndN+ClSEd2jkcQwXBejSooY+RwSOmExge3EUOgtDvVQjWvLhGzajYcMIuNB3V7tkmWXCzRuD
L2wWza3Z4KFY9pWdvP0sFMrVd3fYeFsxRtvwDcdr+zj1LyhmZcYyEYOcDlvgaPJkBfawbPoT+3Ui
bvU3NGfn2B5DnOQAFIQD9IpqnOEYFGIVYmggzwPsO4P58rtJUy5A0wwSPuFX+Wit94uEYxnza34h
Di0GQMtA5EozRHGm21j+Tao0etZveZMEWwitHkkJzJuHvNblUpUYGWieegdccDaC9mzM4Z0jrW2Q
0/z6QvycfvGoHY6sdUvj1ys23GXMOLpwvROIEunfnQLe0oqsmk8DZgRWhXG8AIzVxq0LPZGmmXsf
KA39rHg6PknUeIJ9zFfYNklj0+R5idCNCWonA5GLqaONc0UU12Cyt3JcafPpYIk7tL+2idzk1Dml
nz61dGYDLSQ+OtIB9X43XwDR3g1CgL/enB/w+GdHGHPw21LCuFCVMldkWYgkvEi2a3ohhigZhz7N
aFCySw94Gl5+cRj2NlcIbhzsw27Eam6O4P/aHU30F0j+Ayq8NgMkIibVgF8SvvwF/2ihGSofcuVY
tVH+zOcB+1Bxu2JixmVdVzhmzffWPRTA6tJCO4NMNuv2ujajjOzx33pBbhaAUODZ9viCkcjefR+B
+ui+svDSQmZUyi7rE2Pf4IP3PJjQPedcdlDM/yDUfAvrLDyJNC1zXJ/3R8kqUNYL+82Ox15orP1V
d7QluIDPTqTaFcZ0sMdYUAT+NOpuAsGLgciY2jkBIcudRQwNkq3VNEXNlCBi5Iq7wMh60iJWsVLG
T1fOtAbirN5Z/e2iQUs/65Wd9BgwBFlA67thxHsrCsoN41Y9uotZLRKgPGv6p1uhQ1rMPPsWS8Zk
biYqw/N5kdsu8wYCRaRYlaheCU4Q004gk24gi6iqXsGA6HK6bQYcVGo/XLH3XQI/jypnF80/PxBA
c54DBJCfMJQ/TuhbE87jkzKQU+5YPCbxbRuaWwtJuyDFt6IoM1TkD5fKz1op9FZkVf4vPfda47GJ
iF5n9h8PYLNxpcLw80c66cANpjjqd5zmo8cgMbJHM12pZLQvHSMe81sgoyJpMHNcYuKFe5sKELCs
OKgUjeFKDIA65gUAA544OTIrEgG4gl97J0FYKZ/pcyROq+w9Txkb+vYS55otNdj95krjtAFjQ90W
tMaZcL6Jvks1UgQFKDnpwz09rpimQAajyITvolIkQUOrSK/TaTXQ8dboWf7qn/ra7O86w+0V1s7t
kqiBkynPCaJ1KSxg4s0x54uu6f4N3rTvEHAXIREivPSAgU2qY8ndYi+yw1ZTSAzYB9WPQvz4r/UW
W/1e9FTqfuga1aK5gxJtuDOBw89T2WU2EWkxD7zTxK4YHE+Xqqxj6lvAT9VOeiZPcLerWnErUbzC
Jj04CKP6AHa/4LlHyM114QF5ILiqT8NFw5tBBGlp7VWwZV6VxlyAh1lJOGp/m+W8QQb5kGMgVzp6
WVoTX0smnMy7ZXEsV7Veg2FveLmyhNGqWQVrLLVqkIGORXY/GXzgH5w3VATyryhgSF5y6mQS1hHL
M2fzGBdaXTalBPM/mu3E8Dl2pATPxgkySbeBEbt4cTewg6P7y6smV6kXo1KxsggBoDj0ZlicB4wn
ag7arEkQ+NpZNHTUzgXJ2WHJ7uOzUcbvlyPqZeDkrefm2ZZ3ZUS/AeK90YuA6FnIBjVeoMrwt7Yd
GC7qzbCBM9k3fJfDPTzDvTLGHr4/9F9Vq87Y6fsxAV1XIhBmVMD7twhV3gDKUVCAb6kf6msHgHmN
2djRDi5+4C7vVZOkzv8a2OVm5EI1Tt7BwO34HLhgWpfLJPIrr4UDe9kXnere1BwL5NceqsC4eHW6
sxKhNyuXR1LDVFGJr5XeCSn41ctznrsb2R18EBkBfGng84c2Ur2P8Qbo8dGYIqiSmdksgJarcbd0
GaZWsWeaK7BCW6HQH+4HVf2+RvAL8jOuWjSsjiN8og0PpXarDnp6X6Zja8OiniIo4kN5qsjkQUzt
fgDEIwQnZJSSik8hrS18AG8bwBCAu6YUwCvSN1a08yDZd5PxWq82kFGnyThx7h5Ntnfemwz62GdZ
K6BIwD6ATrM0YRDpFaEEOhvzfr2w1ei0vR1+qw2j1Dm17VBKm8WfU0yZ3AM09rjUOSxRibgArmyI
IvBsDT6Vk+VbkiZ8RPxwPDAz2m5MSs3t4UZILv/pGkwJG375MfxgnW3lRSgJWxUYEjuQYBTCKm9W
YUDSof09PuNu7lntGgUCTHi9kvxiXuu8+TNnGv5xiej/3OHaJWOD1HFMZA6co1b42/bd7EbN7ALu
fGrn76cu7mvejCR+d1Tgx4Tdq8M7s0llfqB2B9Ahy+9tn6tpzWr0rCNti4/GTvNk5qo/nI+vPi03
7sECcIe781G9Of68Ma6CknFa4BsYhhIVFhCUJ8IBSIlOqlh/jiIXkQ0vee4O1cIgslFxjLhL3dy3
l/8AcJQhPACA40v9Akq7tHcqmtKxdd3o05xYfAsoX749EcG8NLNOtVFFm8Af4dNSy7p1UCkl4/Qi
jmbuTxtsqQWVdbS0ufnnYgW8l0m5i4iLoEVhHY9RcS5+rQkyCEb0u32f/8yTW7dyulBN/ThucM8g
6kagsnBUr3/EbvmWlZNwh6IDmka5ylHY4WUfVBhOTR4mWrcmhOYHHKmTKjlphh6sFgDDpvfvR9xt
5uJzvYL69d4iG7xFt3Sze0czMZ67zaDIIgOA4oiX5O0+SzNO2igZZbsVgdMkpDzAOvvNG2y07VND
mEwuogi4FKyfjnd0KUQSfGrwlst8z/JpMFFNONk6cJyxzSzGVJX61VtjbKKb55kWlI6ETNIz7LZd
Ze8f+K0PfDm5HBljhU5UTJJnU+ZahaJmhsfZBvLWr+z2SikwY35F5xeFU6iElrtBJV2mHYgNK01W
UfoZhPsm3EqMU3cimS+6XQwZE7dJetZrLlmZZedW0M+KLX2sOYAp4I4gEjda73tAf/PZq1FG+Ocs
DJqcxfgPKHCbKNLrl/+e53OTtd+TssaLMg5GdbRVqVMpNfTOR0ApX3ICu1nUShTkX78RS1Svdy8K
2jf5m/UQWXbEXI/0qGB434aPy5Vt9d51bBHYxu22CRL4tfAw+gw3Piv0aD955X6DgCCg+AGJP9Uv
6bChMZPUoeR02u3RKprRTv9CISOLfDwdnLXTJzYPmWzkFj5Xw4O7LA41whspx/4WIWG6bKsJrCv2
IoWZibU2I8GN7RcKAp7F5yUJsyQqx1PF4EUi522ZEmkcTXOLCIfDn5Cz9avp345t9jOtOP17PgZh
499Syv8L6cGN78XKf2aCnVm3UeLHCWGENgaf8Q1d+vBrLOVtkxBur0AsydS+MO3o8zIgmPdeTFcG
oH5hryTXRvze9JVX+NPUeFU6KRwp5g3+g2qdFxV3S0415ga/aI9gq4A7TMmue+Tv+TazoZ0yL+bv
I/1GrxqFbQ/mxxUB03UmZGS8bEuvfNJhoO6RETHnIVkOrwn7iE7Us9qf9MxBK8PRDV/kODtPP8YJ
qgtggu20R6pGAQv8od/PfAO6ViS4Dt0NmqdZXNUrN2jF0ExbZkaFiJ+Zv0j8OGLl75G2JuvcWCP9
OZ1aXCW+eM/SUIZ45Ux6S98bDjTYcdZ1vycfcbYxmrhiI836VJBcgfNvhJT7m3GqexM8lPlLCZ31
MKa16NEbvttQaPfv1psPot7AuNG0VQlidJCUm62vxAXDFzjIMvng/3ZpyXR0UXna61FOSDAm+mIl
oEVoRBPiKTDazT0y77c+VtR4Ucaf+qOxItRjpjZ9d+g8KODZMKjSHAq3iCk1VYT/aem3406cYwhb
+cb5vXmzM4WVjHfgA9uA2LNwvvjMnuIDgsYolWuojf9CmJxJBCGCoMk7+tB4ai1qerznmYB0iaok
a8wDmvl1AMdN1swtgZ6Wlby7STtTkOT4vejNCdDaxyS7QlJc9CcmiHbmWvIeCCMCcl4wHl7kznGU
brGsDH23LFv60oaTN1M3mKD2WlOgYmCUP596xpsZz3hohHv0l6F++4V9Zv18z8LTMn6Ct9whL7cU
gqHtrUJD1GRwD1hiD1TtbJEwrf+uffM3+dhcOLGOdeZ4m7xFTHfMfauTDHFCpaME578Q9yalkSLF
3/sQxZyrVnW8Wx56enuaNF955OY6072DwMWP2k1oWW25Us+ey8U8J8E0YrbJs6+U/GtZHGkMVLPi
WUCFtzUXgStIFjKzkrHgVjtytkzA2yxEIw9MbicJYz0BJuh9KUtAEU6gYEHqBbCwrpNz1NnQdeMF
nTtghvAWkxzRPyZnwDedvwowgQ/fEtwkqMTduWCb1aKGGvRpopBmdE5MPoS1T5VKR9c8sfbG5ZAz
bsFI6OFCkxuofseDawesVp57xn5HUEKVYfvRZrpd+rdZnJ7paM6XgnKvNNdw4Do3AsgGAMZZKW3p
qZEKqtb4QLLvcNX+mNLyKBWye1B94u/wrFhUoWaXRLYURJlxtoMTogXt+5Gb/fSCahw9CRA2xk/e
83LPp3yrXakY/rxkbylgvkzdcgdbVceOnXVZ6bv7M2Vub+UXE+lgcsQCTX4wQdzI7FCuQy5pqtgt
jLty15iwJ3OoRf+O3lolWKpDZatL5zPnBsx+0sJU4zsBDBwAnuQnxaHZLUVhijt72mQXEs0mTSaO
4e5ehX+6tbiKLG7vF6KEpRHNHDEnRocTEsOcq5i+NOpMo0Uru24CkJJI4dAbTtZqmxfcVOt94/qd
zqWaHBycUlTLI6NgLLWTwh9GgYCVoDXVhTqyUSgDjBo8OzV+4//dA8RmuMa3Ai5YN+rVqc9nPHfn
M9PQqFoj935c/b69bRXlytEwdRK+RKBE64rrlOkS3LdfGiYCgnLpa+YL9M7ugtqH+Z6yGl7WrFCa
CuM6+iOCxCbZVVgCirkjEtKVQchG1yjo7aiVTEB4mhh+JtleoirTckvtt2bgcavO3ylDVaeDCRMZ
P8EzUR60u5OuUdWrEtaGOEv1yoew3lisWu4JCSHCiXDn4H3NY7G+cgPC67Cwg35FKyZTMMPoBB4r
HgZ8y1GcOxau8xG3GumrKMIcavTwBeYaKU/7BLnf3j4UN5irVkS5tPrGP1J+vZ8ssZ3WOJixQdgT
Qx8sGLkudunpVhjISHpSBMB06GNo79LdmtYMqvJ9QIoeWNbjPivsPJSAteCa2sDcRc0ScKZYECYp
snKbCsOIytm3FyoFPnc/fONJpX0pW3axBVBbO8XayuvIvSEAmCfhTKIM811S5h4BkB6r3F4IiRis
ffQ0Uss3EeJdY4e4bjhs6ti7GmY0zuwT7iJE9/D4sh7YfnXLLAm7nqbrpLg/YNsHlRyjb6XgvZyd
rTuH9xgDFpUmk+wFxGTONCvFLMXLFJnJ87McqxFexr1+br05U5IXNPLYu83Adp+D6ZGntC686en8
k+1pFblzc0NPsMwY+gn2JC94K2UY4e3ebj2VC2IxnVg7jtdHxxrJHIPY99eOF5flcRNifG7Xw3IN
SL3dCkAQ+sl73RLZpBG1jC+UKbrjcvqVesa+EJT1erAmh6+IVSVJPPXDMc4BCUERv3VkPulok4yd
MCiUXqk6IKKaVm4D4rKzndhYrS5BgWa67BATE78LVhr6xGnBydMKxk8muFQAlRz/42TERmjad4Ji
7naRQr+9zNxt0aS+eqnnJpRNhO9jE2s6uR8/OWnfTV0WzWDrKW5BzHrbpx2p6hwu8LIDQKoOemQ9
l9biIov7u1MReYba4TDZ+J2CmkPveYXaIP5/+0ubnyJmFhQuzUY5Vl36YY9ijtcTgPB00SqOAvQB
0ff+D/GhvVGBbyc6iWiQsc9AkzMszzYggJOj9hqhFIUz87CQCwMk0e2nEAbZUQwYvpAE2rtOImuO
MEVUd9X8911a0eQFZUkwNAjgFNiQ6c/2xvCYpufRufsfICvfwU1HTWWU+xKEFVYBrCwnErOkLvqz
zD184DnmFHUB9NjHFhY0AgKC13Rclp+01d8Dw9GUIoMoUpOHy3rMHwpo6eUiUk6fO6j8cXD9HH8s
5s5SfUkCjkYG5LhcqMe+WWpWK1Lcw4egXbp+w6/z89clTR5AxdRIqntdcYFyPBBOivbVz8RI3d4U
bS4UO3bSMqxBkjYX1YslbDgDx2jTtGKSI8jSB8MYE67M9fGLpx/Wykg6L+cW71lNoevUlh4li5Zo
URfbkBXK7H+XA0MPekVkdkDRtNSkWLaDHqMF9GrBZ2KyrMdRKpO+tx+aC1MMoGSuGrghDbp6+u7o
5+9XodqdV6EXgQFuDaSSCIxrA0be1KeBwddrg65VwDWdDN5tutk8b302ARsN08P8PZEf+8kgwW6U
lL+2am6qe/bTzH1OGgS7ABRG3vE3M06xLGC+M6X3si8NJGw0+gA5CGh1S2fwA5rtmASA7KGcxvui
dQzw8cEPdWxpu3QTQQqOAtV2M1eazXYOtHAHqXXc5Rm1/kdMIC6tBbtPthv61gYsaH78zKCiU0rl
M8hUNgv9nxyIxUIOpDVmYvfTfG+fI88QEenRtQuOj6Rfgs9HbL4TATBm3P81mkXd5J150DcQn8Ka
6Cm8/svY5uO9xSmhow0mBeXqhcDWCAtsdDxizVMreZiP7z0qHdeHq0av5kVn4l3KCiOf1oGq6A6y
A3GShgRpv+gHgp9GCZQJbS8p8BQcYuFuUJON2Dbpga0tNCFWDYZr8uwSZg5g6f1eY2+VupRN1MBp
FJf/DrsVJKyetToZcYvS+256zqvoQmvB2y/bokPuv4ISwJ0pgx1CWuucO/GLwfQVRnbdhcHSl9rR
yHyJ7LA+aFaq1lRLDNf0gT9zY/mp0aMyAym4oRZkNnVs0p7axq5oUVQqGX6sYuqhvGqT/+zgCCOp
gGvV9K55j3QJaKS5bg+oZOuQvAuET02/YreBghkoHP8s5Vwxlx2lDADuOT00N7AT7DYIzpWJjucQ
V/Ask0hEIND3yNzN6L8Lb3pRMEsIkNK0iUQtq+Vzco9TLQ5gqGXo3nxLmdT+dqHyogqxKi3dXGcC
eL8sKJDjHz5Oi5GIZ1xAqTH5ul/PSzmLDgyjKYTHIGwOBN2jIsWeGiCzMSinCIdIqw2EV2ykvFrx
+YTrfrSeau21BZoUQT1TBicsaJgpIX86xgkzZfDX7iKiPcRE9hAl3GNn/2D7/kHGZoVvF/TUmiq4
Eu+U3ZIUft4211na8eHMjYXivdKf6QP5n7y/yJCgkpplb9bwAG8KqoFOymRPFBvJJ3ChQ7HyObzW
Y7qaL3X61GVMphj72sn3zbNlPQjSwfbZSPGonbC/e3suAKCEkeCZ2IQbUELGjNaDxc0MSzDUOj6J
DobT7mZsN3qcKi+S2efULZK3dFcanrScPj2MOhe+0fSYhwYdx+TMomblCNnR5EPQzc0VgRn6C27N
6if7W2mQxCc3Qcoe1HUHVWfRItBpNepSH+uSB9TAs4f0aUHLQOpENvUix0qRgJNVYNbvAA2evFO8
4BsdJioZsWxFG9bqgXEGqGmDQtScsueZFojKZtLX5ey2jTQmO/qs08O+S85Vi2NiTsaHWwnxETIA
MBeCjUYWdCHugee37H5ZqnDuIqIQ5wVLNtieSYAYqM/qF05WSqQvWj3OymjER5iW8XDanhhZ6QBf
UrClqh3meieLy9HeXKaxty8K/1MIIJRYZ0colcFXB3zgFaBdTTo6O0KH2fROlde2ZUFgUdyCzkVE
Ib5O4daXM/VmzzBCsRXhzgGBZ457M8uPpZzScoYIswaoBEJNKBMELgP7oSudaS/vEFIZHxgTu91j
LuAejRIXkuSiU8g4GDuA6nbpuUmlFr9XwkKJmVhYF1jnSItg5acAvnzf1ufowtRgJ9HQIwaU9qEC
N2kQnlysIliI1DRLNzMvxAtld/1uu/V0hQoSCVHrRSjw/fgjhNDQcWEINocJCoRo9/NeifHL8Jxt
+byjfB5ZcpbeA/2+inCBjKvB5CRhFvfbpgV62QPM5z6HtqdjkLgWDrr4jM+qxSVQnOb6G8Ut3m8f
Ts4Qj1m7Uh8r3F8ioQAECJU+RzlhEBURMofo78wUjh/ykbVOYIPR81JhWEs8KaiKOqPHdHh0Nybl
WUKpvrjrXZhsYLS+R50ymx/GWADbNMHwhTnla62hD/Zc6jeTqNfKbcwxv8JAcZFaeU9TKeQPNiUk
OrAz6zc9VEnkM1FrhMKEq7nDhZB6zv5GBAeyx/bcy71jLPjNvz2wSqM/mUOma1OkPtODh73MNK0V
ajVkxPkhLDDuJKghKIoiuFyJcJg1LPWelDT6jwdLo/Pj7g8w4FvgqmSMoqHmA2tQGIlI/0Ya9AKh
fRtvuU9piWa8RpWDPfUapu7JTiwE9rhZAaXOh6/4aDTf9GBrCATXNBkyotax5eJUH9e/9eyVXW5A
VkkBWkwG16LD8m79ZQTBEHAPt0ovZsBc74BucvnSaXC5o4rXIpbWULjWAkp55D0/DmaqSQ6vq78p
g++5OD5a1Qc2GNvcsACS1sf+yBUYtC9YpYDovMux5LpjAmniyU4lfYnLXW4sR0ohKRCSYWcICXP7
bgsMwib8SSt217cJRCpH6qCPWN61qXlNxUHxg/MuMM6x89ByO3Hfah4Hvd2PxTrkTL0omQ6ZI196
Ow4kMVwo6R+qAcJznFqHR8GcU4exqO88VxqaRZ8UjraklFuGlKxyNEGL0lem9XMh1DF1nvy02Peq
Pis5cWWvt98RJJFXHF++q9gMfsgCCOcwPGLRIRL0w30rcnLS0V/oDVZ8nDiuYzCUQPJrIMaFdsYU
cG36g0HFSoXj0jgGN6eJrkMJk3HjEfhBQHv4+GvzlwvgbAeJOfCgVUocEnMZ2j7sWLZLBUm7VbRB
9c2sVqOk3g53cmtBg9tc+4u+KhGewluD/HK4JxDDAFANSygNQhMEN3QuFj11bResN3gZ+qS7Yil7
ptdTlTIlHIfTs6ALNeBpFOo+eb7SWPLlbBWf/ZOXSAUndi2bXSeeh+ulU5isHNwwrTff3awtZbCj
jHkrlIjpVpJSCq5GQjaEv8D0wWPX0H4fjnC8FAlKDYQh2Pd/CYOjhWx9J2pe60ftVBx//0V7yl0A
mcsk6ZoAMjZCo//pDQSrR77SvzJGpJHtXjIQKyrRceieeueqBgYQ3ECaKtXtjomH7Ea0s7rTHu6I
bwItsFJ1FScs0XnWCKs+HVJLHomz6o1v2MrUfm0Dg/ARLL0O3NQ2ZVDguspqR3U5BK0NkMZyJv6d
OWSRvSWkONNbNSk3S3OuDZVOB1TKZSiS0CFCcL3EllE98ZguZtHm2KML2lQhqHYy8EkcyHG3Yri2
lKyIk6m9/7IFU1pQO27zdUFT2Ngu/wd5RtMiDvBJ8PsD/9euiJu0fVn9WxpUmjEHAEj/cd/hy62A
kIcBXANrD3srgv3Jy91HFNmaTSmeP6Zxf9jkZayZGIS200Vc/L45BKLVaCmfJ4ILFu3SWneA/1jj
Ac79wlg4YUSGz4koBGdF2rj3brvWA5T124BUDbRscx3GqJqBe6bCN/hE3MEjhxtCNK8YL80cMzeW
V0bpUJFBC4K6gcNiemZheLJN8HhRUoBg4v6BLdtSw9+UNkWfWFV5PJAYLPDUqbZoBDQhPla8fYBi
GYsI6LKp0/AQ4QInJ+JyY5FULvkB59ALbq9WJh29vYBkIxijCyTkUseuCOzoIhOwDJMxYdrYA7Fu
U/VjtxRyTAMD1FmFKVuZFiuvZHbiA+y8/5/vcYvtCYxStcyxezNkxUt21rD2WunHP2zfEfJnNJsX
HfRz34g1KY6utfCqnWagOTNF/83/IcRL7dCeFR0FMJi4qE2qX9kAqf84djfJLQPmUX4EI1WfmdQm
2Vxsq6Z0RyZCf2wXBWe6qQlf8ZP5sqC5qvNPVaSKytf0tLI/tXJ8TBaPEvQPjdO99KikPsdr2++p
2ZmAIiD3bFPfbYbMgTQD1a7kgNOYAkP5ULy3ck1RXhcT54oZf9Lc9c79SPNqKdp4fwqXy99l/x6G
7wfkyI14vu6aGIcj1ZeRmZaMrUiHB8rhAKosE0lfuqfVcBRH9xL5hycKDPxEQ6neeWu46mavODal
o+tWMRPih021Z18HZPRsboXiFWccUDp25lOImqqgqeVZOJw/kMMQE7Cg/SzdXsoWAsW7mPi2HVm5
4dKv01iJeaeHxSQgwb719qy7RJiIKMUu/q3+ejVYMRcwe8VwFGkbsAK8hJlIdjKnnpwHcTGpA9U2
sO0+xip6DuiDLz8wTE9QCStaU0jxlLNR1Dk1BAtVDmp76EMP0bUnF4iC8tda6xzyAYZLUR562F0K
ovKk2P/4G+hpdSO+hkbm/fHL77mjWL3vCUp0cG8qQXCyfx6rrzD8Nn92mbZrwjIQ9ZuRuh05k6I2
sdCk79iwspbGkFEWKuMBUNZC1mfv7CP/bKLldf3ndoMl8cYpDiqXEvNveIPti4hlhP3LCbSHm2iD
Ka5cvKHx2vN9CzvQhjxk/bcqj2392vOjsvOwjQH2fLIY0dtnawsqxw1DidU+NdzTiCDALPH5R6U6
IknshVRTWgOz6B974jVjPSHyi4tzf8qnHOJdQWNysrHe1efOVlo+HpXQLbFj0DTkMYQa5HcimDS2
o+O/3N81Z3FRWhUHY9FWKFkUsVTCh3pewOt6uOCmBwKVhN47yd3Io9tz0JMouTkgtuX3x9tKdp/T
GdDj8jf+Pcowp0cBLhxs3qEPlK9Wpdabld+jCJUEnlweLP8a+e8XAUMPHF3lifEb4kCTwqt/F0tu
qGXWPy07akBhcNgbO4scms+JwSaVJsaoVeA4xva906/fTRMiv3LnguNv3aBW6hLEsU7UMSrI4kYg
juKfj2GIiKtDs4HF2AG7Pe2gyvphzyjE6CaE2p/CTNsD4vfszJs3GFjzir//3ltdiOoRReRSC4oE
ed9R3EipNBCZdBTTUBGvA6+cMrooGz0HYzJP5SpXzodeveAR24xOMX52ZKQAnqK2s9Ujz5JbAlVz
jSLCWIO+pqtGSWHotbsDrO+HRT24bY7nwRiykT5Br7/ACR7wr/aUBbVhMLVoaqz5oC6ckibgazwO
VP2oM2G1F1bTOdii8fjDzw6cOqA24tpCwYnEeRkIwUarnClPi9Ya6UfqQAykLgZSwryfYOzKZMV8
PsKCH2YojwmhlUH4sXihYmhMlpEw0/hblGARp2k+xDA/7OWJOw1AxxUGKEeRKM+DMSGx/0hCwosG
L50HZAGKBT/l62UOP5xqilxt3KBNEQeIW61836tOc8n7knEvZ8qKdWY74Og+7kE9gMxPY/2SXV8s
oLzVmvuBWvDVOxyBwji5P5n+2RxL5u+xB8jypaGT9RqTNIMDMyEq5mNFAIKyVo0MPQsgB6mAfI7n
Z7TNoajh1AFu+wLgukokoNi3VztPH6oAWHMQPfZiCgp++aGD5dgO6KRML4FGmy5aRNNQDmu25phy
NG5mOGsqYz3soHfABRftr5Cd4h7OdF8HjrUELKNXfbh0Bn3XZN9O30CnHBkQfVDXIDY6Ts1MjlWc
SekBzm8Q2JbTEc+WConZXmST4SeWEVvK4FKnm7K0R1pcDumod8PC/Kyp+xWfKLw337imfjnh0KQ4
ESpHv2epOd6bqFE1fZpCJNxTuqIpXr8tJz4GiBG3PK7z1VIM67eGmhm4k/2RYEl7XHdP+D86ChfM
Aro1Qs0ZP3d7CCgtBKmH8xayzOoN03CEZUXaDxAnbNaR1Q31Xb4/OUSfcGPkRaqf+Xd19ul6rPix
lOs+iB4Ch8PMod6MpTfEB9cR2erQIk/GmyJxo9u8hl3mS3okpvM4oxPPwK3w/x4U5n7FZqSBk9fo
KFmBSX3YwugGjyeQZiJUTI5oBUYYNadQT1TI+6jRYu3OxXPo2fAEhD/xgb2MulfR+O06Taw1EVLU
FuqGaeKKnsFBMyVaGotB7nVscUITpXBOyD/Nn64lTOvlYPLZWGMWDaacsLHF1Af63zt0NkMcMRdZ
QoBM8VfDp2UXQI5IaotgSB95sAmhHGQrg3ENdrH0cOEWQ3Irg4YaoaXWplr9dupmP9mz1MvRFxBg
hS3oGJkDE0hjsb9vqmokYoExF7esXHHE8l7h+aARG3t5hgi2VT8PkPhJSir5m0C3qrq04Hs6ll3g
iOyvvhTYrm6kpsapzCvClSejRXKOB7xwzNn1v2pNg2knwDqT4O7cV7BNUpjKFfEuSzyotXTrBkLB
EmzQ7d1vEOxpE0Cz2K8+HF5pPvv4Opvh6ZLY8YRmV0RA9f9FlCqUnmdd5BhCM8tfPm4OaH84Jh1V
TFXOveuHTZZ0b1d95H5O4dXpylGN9iTyR4kTHLTAt1v7x9fWkAQNf8NKubz9W2rl2OiA4+phVsig
yRWDVXKu/33e9yzDsd0/hYTPAWvVNtklHGAs5yX0AHtQRUsS2S8jxbsr0QVEL0vVW80MjyZ37tUz
ALedyL0Shxhpri9AjgF/2ECr1NYO5pxCJpui4q/LMOpprtiYcxEkI0Uz4pA8w8sPDcOSLXK8FOiq
A/7+CFW5CA+nNpBZrrZCF8MdR2odTk8bVYBk8jKeWPZP03lf2JtPTKtS6BzennHFPFEB20GzC9gv
x+5B//bq8aXz4Lqj5XpjMW/0vzPv7wXIpfDK41G6cc1E6qRbrZCAWEHZvJwWbkHAxkG5GScZ8re+
IuN0I/xi5UQhhKXnU9XIVJXIzQTb6CpcGmAza4JiXcmOt2zVFga3FMZEvDcczNH0nYs8tKLeIb4n
F+RIeR+vFC1bcDaKzUeYwiC6N6wXf0HutJIra5B4vs0CHTg27XuVIe2YFc5jqF87mHOS3Gje7U/j
ykp9g+GK6p/ULpwgsSTTAMgyjprpyn6Sxk1o/xxiQ0oxLaSCA13YMvLX+yUu/bvGJHSuQFfJqD/H
zyohwItxvZvplfKU9ropF0RHXD6Sl11MMd6Ra1LZBLKoIb7F9DeI8UkllB0XhNc5WseY1pEmb2sQ
9NjQOzyKZiPOzXC9Kw1FDR6e5Jkda6UpbPF361sl3E2SztN/tOpry/ohwMMHDvdCq8DBWuWTxwgT
p/woyTbY7v3IGHSjCu/8vND6Z4whQA784ud1NMwE9hvR0HMIcIuLC1XZgEqHP/iazs6VPUt8P1UQ
EkRcXTqnt+nO/5+6ilEGsO1SLwFsgr5iFFm8U/76mxeP3VNm2qFJAA1dh8PPUV7U6AT4Cf3ACtu5
S+iJerDxpV8yYIgXv8z4SGfhsjXd0c0ZQJJmRwjSC9PSwMEOlon70E5fuJO2B/36YAkwuctumS/5
Nu+g+/RDAiPutIOykL+oDrNUrTAz8kWqKHY7e7b+NJ12FcWM/zGZM8hI3z0obWDAh1/eP/BJM6ka
mTuUdgOiAh9YNefkjt1Y0cT24E66ilQ1J9NyJ46pRAYzE54ZvIlnDquZZNeZq/ohuf+v509XLGs2
GZ9Xs3qApNj7c9BrtsaFqSwowwI3+/cp7QNGtjdqFU4TeO+5tWGDhdMoJ8YkjU8wlttLSBmZnGYj
ynYqq7EXwXE5eAEaJL01rNecVj8a/WYn17U0Z649UX34nMosMRa7pyvCqo4TVrjepDlm9JDJkdAd
qKnbZK5KiX7BhGfDTbs8gJCZub4KFXCc1K1Q/QtLcB9B6jv3jbTFk/qQk12HvTQiGT3P4f+ja7Nc
dEojyAsE4KeaovGqbpFWR6RFsa2clXZYxxi1WTZYv//v7xEA/TuGckudcxjWCWG7qyfJH6YGHfcK
QDoRUGYqcy5aaG/0yX0oEcLOaQCgOaTP31hDqdeXiA==
`protect end_protected
