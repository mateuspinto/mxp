��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����<VF��B�k��o�*D������b
/�G�d�}fW:GW�h6��$6^W���z�`W��Y0d#�G'8�y����	��{~�W�C�������^��z����O�:*4�$3��vƧ9=���Vù���n����atu���V,Mr���Ͼ���ӡ�[ȁ.d�0�JV}$�����MS���I4��9w1� ��U��ՌMԤ�Z�F��øǼ�bЬ� ~J񮅴�ў��v�z�o����G����)W�SOw��\���,u��W���'w�+i`��:�)������|<��cZ�=<{b��N� !��~@��]?�R!��Y��l9���.|-�6Ng��`е_����.o@�axA46Ӧ�Ҏy,�um:�>�m<e�h��ʎ���g����Toy\!J����f�."	8�
���wd�13A�+��.��$gd��5�����0v�Y�n�y�Iw���B.m�WcTJY�h	��5Q)+��?79��Ⱥ��s Ė���0k��7�":
�6%�.T���F��"6�G���ÚN	&Ԁ�b��Pۋ2Y23))��e�Z��.	�?ʗ���,��=A�=0�jlfF�!	�,U��������JE���}�d�+:~�%���? �[�g�SB�D2�t
(��,�HG�`�Nh�2va�h�"y��5_x��P]|�D	�FS�-C��4cԟ0�}ߒ�`�X��k����+we��{P�O\i|*L~(�Jz��@�2��S(�b������l�����|"�}R��l��I��H�/�\���ኋ������!�W�y�J�kx���Lz"�S���)_��zye����7?�c��7=�W>mNy�(S�W�}d�X>S�q�����3�����#��ς!�|^��@��L�;PHH�x�����=�����	���-D����aRn��b��G �\ͪt5���A�y�|�^��
H\�G�o�*
Z��Q�3����5�˰�E{��9擿m�whd<h�{x@%���:n��q�Tj��!Қ�Q�{O{�X���kd-E��kq�n��rxqF�R�DH�(Ei����>W�@X����ea��˥������r�e�lS�Nς?�/�Q֩��K������DKOv�ԧ�%��󐙬@�E)Ι,;ZL�r�晛d�6B:� ��j�g�z���Yt�w��l䖂���R�,R���`j�XV`x�Oi;K��X�IŻ�=��C5��N#f 6{@����!��~ ����b7��FX�Υ��|�iu������gH�6���*�Lh!k�dS��pqs��d �X�A3����ct�^R����s'�0�dZ3��LQ�3���i��%�>˚��F�9q�Ҁ<t��W+����$a�����W����_�yNz�|��}̎]���j�d�?�7g6���w�?�ɂIy��/:#;̡���[D��fx��qd�W�ӡ��jXS!�m��0E�5�g��dg_kz���I��|^<���²��??����������P�:0��7�P�t�p������Fٳ��&a�-/cy��1.�1�wu�E�DL��B�Sa����n�8+nթ���� �Ӭ����b��V�b$W�n0<j��6ݙ�Fut�*���v��si����x<gY�a�:hI5�3�z�p�Y�^��?�j��LdJ���(��NTn(�s�Q�q@���O{����ل��!��e/^�6(8@Y�t�.ADK��Ñ��1�L��y�'4�����^={�R�{h ��o���Z�_,���
~Y�l�xy��i�/��V�a��	Œ���x��K3wW��:PC��4��x�b�.�8H�A͎{��6�4Ɏ��$�%/��G#.#:N�s٬�|C5�B&�YZ�u3����׉||]}����6�%x?#�^s=�����tYv�^��$�M�\Y��~�{� D�����$�����}�`�,⨴_bJP`��@�l`��������zΠ�~�Ҩ4p5v���p�z%��=�W�i��s�I�H+{�gv}{�"�KA������9�Q�`��t��N}#рfu��xnu�'h���`Bb���W, A\XjId�b�;����J@}�$ۦ��/�T��\�ťYpBs�Ã+�P���y,�<u�$y�v�2D?}� 
�RY��D^O���D�PH%ۖ�Z�q�L�7>�O��c�Q��e:^�,�a�����w�3Ν����|��l�NZI�6��z�W��܊��5����A�[�*n����f� �A(�̃��M�VF{)5���.�4��?�a�/D�� p��;��ZR����d��&�k�W<]:>u�����U濌���{6wl�% QOQ�B��T�Hf᡻K��4agt�'����䧌 @�ՖԿ��~�k�y�tx&�Ͷ��]\
ՠE��2ùNw�vbԂM�^%�m����}VH4�2C6(�zߩ���!���X�98��������n(xH�P���B����J!:�<��Ի'/��vr6!���h�w�f���{������f��,N�>tD����	��ASQ,�?6n�)؅KY=<�[���ݣ� �p�$MXC��r���!?8���������D�>�Z�>�����r;,z������_� vt�Z6�Ȩ{|Fq�p�S���Ĵ�X�f��]|ud�R!l�ttM9�/�O�V*M8�毨�����gZm�l�kHz�b�%�l�F�l��X��廵6�΋�^Th���$&"��4�1����^{6b�i�>�A�����8m�g�tC���K���jP"?S�x9e���%��������A���z·H&U���_DGţ��v7V�a��r��y���1��N�9 � O�����'�2Xl��vt6 ��;$���9�G��\�k�{�@��>�{�U���7�am7E	�����?Ȃ@�x���]�>�$�E Ik��-%�!�����,1�]�����`��*}�ށ�%��a܄�~Q/�[���ۅ��⢡�2q��b����?�<n�����AJ1<�Ppa,��OiA D�J�hѥ�mdj���IN���rqT�#�K�aj5�K������g�k8�e��C��)��N�������� ��$FMo,�"��;���x��Xފ����/څJ:(�Lv��9�-�SQ�A��Fb�p�3ʹ2:L�o��A�8�˻����WGLί��.��hJT�ӫ��Ok^,:�Pq�f�I�э���F��K�<{^�50A<Ny�1FS���,ST Т�ف���P_����p=͐��	��~�mH�Z�Fr��-g���<�m��_H�}���V_���p)��9���p�=	k��S�aI�!�il�Sbj��u ���#�r 'T*`���5<Ěe��w��3�e�!d���zI|��-dI�$+^;!�� ���HF��$��1�y��b��9L�iP�*���}vbԩBA���Ї]��8i�GF(�(/��4t��O��@��a�&mX�'轣��
� �̂�\�B�]f��� ��aq�*�r����mzO����NDܜ�C�� �W��<�M>v��G�ϗ��r��-,.6	8�9�-��+i'\m�e����P�go��jB�q�mD�Hj�\���C�3Ͷg�x&6f���'���-�����rz�H�u z-��Ŋp/��X%�I�sޓ��\yG= LC7�\F�U]��u/�������_6ԈU�~��*q�)(Z:�k�({�����%"�{,�3.�D�B���E���0۾y"?/.�ղ!�B�ט� +�$nr>�u�X�T�#c�HO��h����~���f��(��8�3Ոuw�7�(KV��Ť����`��}f� 6���s�
g[��Ip�D��~���U�c�p�P��@�ZJF�uj���B9+fG�	+ϊ�� Jtod�Q=�T����G�ONή��~�J?���\�x�����7m�(]���^�)��)�2D�]���q��P�zh|�k ��إڸ��>������c�8Q�a��h����T�:$�r$�݀��e���0#mxE�����eVE-�wp-��#U�T��XK���2Ǎ)�����_��]T�RW��I4R��a�����8�>P���=0�9�}��rkvz~��U�X\\R���1x������4���D�ν��s_���tI� ��v�?Ƥ��qY1�b�|��#&5V���k|5��D�;�|��1���e�K��%���W���뺆�E��1�i�u0��w�n��aU��Ҏ��OpbF_�� 0�D��l}�t�M}��V'+Ŋp����JW֏FA$B����h����!^�p����Y�F�
J�͹�ʦ}�pO��Gf����`��'[��9����a�3�pN�J)o�!�pqe=ߘ5^�V�	�Ԫk/l�]��gq�]Q��tt���}��כ�M�����x��Hڳ��f�vз?F�iM�b�����禿��OUݛb?���n�&��M�T��d�ꇗe�´tX#��� �_2&�n�(n��U�"��"�~X�d�-��"�5�FI#s����U����T���jB`ڦ�./��(��t�g����(m�:�9��(���)���c�~F�� �#n�V���:؃�W����TN��h�,Ttݬ5%���k�m��`�oi�35J�
;�,��_F�1Q�ٱ��RF���:�):9��h�vSH_%Y���S˔բ�����H�|[]���U���mΌU1=�U-Bx�Ljק6�C~�\�w�'po�b���F�����J�@�r��}%��`Ӿ]Cŝԑ���AI��3�;�F�0�P<�E��)I?$�N�h9�w��lwj�l���[���k�L����-ZͅZ�A�a��A�����}/ؓ$ѱm\زۯ��U���9h�rî$�}��8hV����7#1vň�>����}�z�vTcx����т���s��}Hn83g�#�L�I	�/�����v;�+��B���J@�]�@$��K&�������w��SX��f]�d��F�n�y*�A#ă�$��Q���9@�%����> ���&�0^Y,�Ԑo܂��V>��Y�v���êgt������&�z̢�Z;�T���W�R����0��E��X�7�*-���l� ���>E��3Lf���҂~_�U֥�W'���e�7�1�D��ޱ]�)3�&�f���8|Hou�i��+$p��!Ӂ�2fz�۫��2G�^xtk�TP+߃֓�	���VK:�uB�[-��ȋ22."F:ՍY�
��-H�d���i��lӋ�l�(53NaJ�.P���wZ�r��+�>*$]E� "���z�mҏ ��q�2�(j�$��k3��S�扵n�~���[˩f�6�Г=>
TT�� $��w@�l���cT��qa���|�\��7�'Ve#�֣���(AH��~�?�TY�G �=e,^g���d�.HP�����AJ��5�2�����p��H�[�@[�3�'�)o|����J1�jܤ
PB {��c)Ȁ�.X+ ��W�žx���/�u���fx���V��S�0�N-��z���f�w�x;g�ec��8>�H+<%w��%s�·ҁ|�腨� ������9$�K����te9N���o��RvWG �#�O��Y+��˙¿�Tm��yˢ�"O�^	���+��Sk�2��:��tZ����$=�|��tqijT&�l����=6(���R���nX�/"��f�{�OH���M�?�h�u�1�h��⏠ҍ&�w)��9S������?����|�b�.��7X��[��� �w�{f�X��	�D�J��ع#����0륑|%�f�l���ρ%iÊ+֙��Y4�u���H�늢vvӬ��[؟��I= ;�`�urt*]��4!3��~�����E�@�4��_�̢�c�{��Q_ݓ�y蚹Xo��"�3���\���@"��{�,�p���5m�8�����O�u훃�{�\��*Hr6�^�Э�YP�Vf�q�{�YQ �k�|�c�8�V�7��8>�����C[�m�2{밑�k��"��J+%Sc�p$?����B����a̜Bq��JJ��b�L���u�F�G�L�� 5+��B��1�|j����T����h̔B,e#v��gyD�Z�_����r��YQ3ɱ-8��9�b�D�	F��l�>��8]��AD�����u�I�$������`	Ή�e@��x��h[�f��}����WZ���&���Z��}��R|��?ث*����:G��U4Fİ[f=*y8�Y'Rg��_�r���'��xX���]ҥ����$�d���%�wr�/���*_��{r�!L8�}G1���@r�����ۅ�#��(o��]yƏ�A��X�Py�R�Wz �=��]ycJK�_4��[;��p��u������Ǿ��˘ՈJ	����'�Oy��}e�w��ˬ�W|�ԃ��v�ڪt�w�e2�L�D�ᵸS������Qq�tr� L)��^k�䓩��dfX�A�T���ڙi`�	�]4nx+�����\}�|N�����ϥc���������]Z����?}�b`�cB�o�6�'��3;�&���q��Ջ��@x�|0�o',%G����f�<Q��Ӟ%��h���>GTB�h�+�z���v1�����N�)q��I�sCuX�Uv���f�#*!�  �k�&f.��
q����Lhƭ��4���������F͐
1�'T9u�+>�b�|�#6�l�Z�F���">�����hsl<k$�6R���?e���Y�=��O��8�~n�:��J�0ۚ�M�����#�IpϖP��G6ӝ'+S<)��G��.�����\���z+�����/��i.�Ҳz�`J�2ƪ�lᣐ�!�y/���h^���Ѱ�+��E�d����x�UR�ygP�
'�7��Y��w�7�dv%��%u���z5x�1r�����ClX���.nhEs�R���'�1j����w5;���Y�
k,lh/ Ձo�UЧ��|�����*}�E�+K9�N�v3,��%Uo����/���`ŐK�F�%��~�I3����ǒ�����wS���ƘB�pA!_�7$0G/��fs�p�ǋ�3�b����vt�Z�C��2t	k`��o�fږ��Q�B6pt޸��'���<��k�g
������J�����@�ś#��Q܋����'[�K�SQh��E6\)�8���MN�4(���N)~�����xUb��lk��SF�񔓕���_o8�9���Eۍj����+(�f�s �;��׃E���qC�=�J��-�bD�HG�����҅[-*db�������'���@�����zt�#c����E.cgN������>"��5H�0���'Y�H�g�*Z�Te�tMN��K�~6�����{u�(���γ�vd%x_O��r&� �w�X���|���١���sكS�U|���0Jq�
nD�EӶ�lA��朘i5�^���"��\��eot�땾k���+>�C�mn}I]p;r����}���\��PV4%^��8!�x���܀�w8uz;x�zjC��9�vY�hq��I���-��ܟ:�Y-���~
�nd$Y��"o�rd� ��8�]*����g�T@q�o���������G���y��x_c��ٞ�E��#_(�Ƞ{l�b ͼ,�����m
^`��a�v�![��m�K�eɃ����B�x�q>�s��:`EA�~���=�cK`�#�ҡ@��#]�A���w _�2ώ�!>�_�����-�.�>j�c���K�d%��*I N�����4��~v�t�z|�,���]���~ޯuS��5k��L���ӌ���T�]�Q¦���}|���gF��`�Q�m<�6V�υ�_�I�|�*S�FURM[�:O�O�naμ�]��W���x�6��"wY� צ]����S0V�������d�޴ز��.5/&��tӇ�!Ԛ�% ��\������d��]Z���3�~Q���j]���:�`�=`Vq�4�	�.���k:Ʌ�bn�Y�?t�3w��+�Yy�5�N��iiF⾢VIƢw����ONm��$�";���FN����B�Z��Y[?�Nؗ|�1�noˍ��*�X�e6��SM�9���=�< ���~xtǪ�u��z@#� P��������c{�������MҸ`��&7�)G���w�+q8F�D�$<,��`���=��
8:�ģ+H>8��L�q�M�Y�Z��v���gv��MP�@��L[�O�f�1՛��$��-�}u�3g���p�*4J(�) ���Y#K�{D�M�"̯O?,�'g֪4��3����%0�O]�d/�ZY�hQlDA�%� Zs$xo�v����%A ��9Ոm��$�Ҡ��AtB��lK����S)��ρ~3Å����ѿ�t�DϪ���e|P�>Ss��{� �\�F��Z��\�^:l�i;��E���� ��L�wvd7��}y�tY�Eqv:�� T��m,����[����۵��{"��:��t�#�*I�ds��V�Hʰ��n%��mG�����Rҝ���-a�k��*�ANX��pw����u�H��+��S�	G�M8���� �P�y��I���$E�_X�( \�n�bv}��0'hGl�f��d|���O�o� l�.��hR�2��?O7(%�#�W�	<��B��އ����<�(.u;���.,�Sv�|���h��"��U�]j XbC�B't*[�b˧꛴�::�(���d	Н�n�F?�e�0WpG�b3B �T���HE?^a6�j��5�ܗ���(�c�
����YkV��k	�D�E�����r�!�����o��U��e��4��k_\-}F�u%�ú�?�&I�n�-��`QZ/s�.H, Nc�;�����gTE�-���B�CI��X�p�6?��!����wHs%8�xCI%�k��;{~㌏ G�[3�C�O>���'�iO3�G���?�v*���F�z�H�N�x�5'��g�]�M�5��͒�~�������/��d����9tJ>�q��1��dn��k"���A�C�	�ȍ���0��4��vWl�
FK�y� �0��/�=n�^b���zЎ9-�\�Of���ɺ��97ew5�X�S�l\h,.G	�T��E](L�S�T����7P��\��s��(2~�l��?~�-ĥ��C��V<�Y�qu��û���J,��e�{X%o�j~�s�
�[K*��頔2�����������T��)�ZS����P���2�j���pe�񞞷쐟:�cw*��65����ݨ]���Fl�G�C-��x�LG�Y1��OH�d~�Ӳ(�@���z�w����lH�Ⴀ��W��g����"�I��B�5ag�;v$�^l��۱|\y�?_V��N�(��o����4F��"!��Z���6��� �{z�E��X�p�4ڶ��TJH��� �<�I�nz�H����%�	Íaõ��'��;8>^�~c�T�б/�ԧ�HnY�s�8���g��iu�9i;��©���ع�M�%Y�K<�{�@�"�l��PfQ��6��b3��O��E  ���T�,��Ҫ�
����aƆ|"�����8	k�4k�\Ѿ3�2�*�!�Mx^�rA��<]2^�S��e�����Dm�]g�2]+:0_�������¨kQ�ί+1�� 0�g ���AX���p���&�h�8a��~a�#�� Ϫo`Y4�P��N�^Y룩�[������{q
�Ւ��1�/��ތd���31��B�-�֕1U!�5�WO)<���- �4m�ؚ��e�7�a}:д��AE�^
�QmA��,��	��|7QV��*��&�/0�F`j��{�Q�R�*J
_<�Xe��g��
��u:���;��{��+ܱ)Xӡ�����X����}Y���Œ�=
��F.� qW���1	��y��^]=C9r���+�H��?+PE��y`�ۯ�Y]�cS��5|��#@>m�g���g��&�[�b���ú0>�/?�bvV֯�����
��5���A�]"]:�2
��\|2NR;K�cj�1OiI�u���l��6Tq{u�h��3�b)��荗��S,�`���&MA��H)YGa�����(�X��IL�nMv�,��
eHT��u�~;�qr��:9�NvpQ{2�^�M��@��+"N3/��uXG}�`'�n�|�i9�9�g�G�`'����ʓR:Ը��Kv�2�|�@rVK���V*yP8���_Hx�E�%Ԉ\���(�U��v��O��ءqm���?����x��ڟ&��8���%�x;�^C0g�@(?���>��;�r���@�
��U	A�vn�{�%3�۾K��^?%D���^��E�EN0_��9�̈�$��k?�����[9�����pǒ��=P��X�?�zrW�n�O`���-��N�[�,G�"�Vi����˜r���g���=���wNZ�&�&nd�(��Qo�wY:�����r�1�Ŏ�t���;J��Kqw�(�h����:-R����>n�.U*����u{���5k
k{�s��\|V��E��`u�&;�z���[��z~���Qף�~�ݚ�z���a���pA�{�M��A-NJ��9��5����h[v'<nC�[pjqy'����@���鉄"��W۬wZ�Kꊙwr䲄���]]Gs��~Tw���e�?��
%�d�)M�z����լ֯�E�:� tC�p`�fs�fl�K�e�HU�J.��_���H���޶��\m`O饭0R|V���cJo��a�L�$�'�/���eq��/fq�����>�S�A��oR�ሡ~����ቍa%r�~Z�ze<5v�Y�d$�~�n5�z�u\���6��A|fR��p���'�˥.i)�?������JQ��Y���X"f@Q$�%�/�My/	�ͩ�E�"��_�4�3� +d�]�~>]�gR�sb�����II�TE���3�Yl?И�Sp�IH�f:5�8��aXy1���(��hitJ�(�'y�p�,��l��&8�n��>��&�C�lK��z$�$��0t(էZ[�Øɠ���ud��͈��ap��\�*��)��@�zXg+݄��.X
m�@���-iz
���h�c��z�� �
}b
/?�2��4�i��'�)��ہq�S�6��o�8���T?	��D1���9Lp�3�{
v�Ƅpo��x�<�F�+|��Rʑ�GVd�ݻ�֒��\K����`�Tf66��|�#�����<�#~K�[j��󰅽���O<�䶮��.j����[�<�������4���~-A[��	���L1����L��S��`��}����xj�8�>u"~~���]�4�����z�Y�vi�<��`T�X
���� �'p��`�b�Y����t�E��Zk�q���}�zro�e�kN8�����-�d���s�����7��G�&������2ӆ��^��6w=@i�_b�jS/�6
�G{������+���G~$z����B �%UeI{����x:���%��W��L��wLl�T�?����`���_w}Ro�v��N�0j!)���a����ZK	��⣑]� �}M�z1p�����)t;Md��#��ĩ������ �Ox)�fg�z��ܚ�ՠ��B
?�u&.��z�]%�SH��bb����k�����~��,�����U�Y�9���>�p��h�U2^��/�C��E1�gK�-bϭWI�����t*���o�g�/?l���b�h�ǳU�r"1�Z�T�`V`�Ҩ�Dv��H����+��2�2��.����H�X>D���RMF~杆,y��u�˱܉��nm�09�-���A���č|о��-�k�;eL��{&| �p��ŧL�}��� b��d7n�]x��C~�}���*�~/S�|��[�*T��*����orl�>���u��`VH�\*�H��;6V�P[H�S��Fmb�T�Ţ��6�^�,[̯V@��<%o� X�$���c�!��,�6�dB��[� ��$�[�����/>`n��eǊ|��ϩfy�Ӯ��{#�o�g��a�BH~�����~O�6�^�N�XNɌ��c��6� !��IM��������3n���nH�=d&@)N�P%֌�>�t���K�,V�G�]����'v[h Uf��"���ț�Q�
���a �I���E��T~y8( N���n��ˆ�G"l#�o�ǽm��yX]�<-�ʐ��
�����x�9�m��TvkD�!�B[�d����A��&�g�\���X�����h��j��Ӵn��ĿCQ��=o��HĘ�T��&:�JX� �9���?�]-0�i�1J��Cm��4�A�)]��nGl(���rx�;=nN&������|`��L �?%�Neu���m�!m���;�S��@��6�C��"����Zds	^8H!��$p�G�0���X�9��8!����{Vp�G"#l�\"X��n�t��&&��3OCΌ@Us�V �d���exW��@���$
�"�w�G�Z�`�.�t �[$5?X�g��$���{����f��8���� dO�M8�W�\�j����J�o���@�7B��i�~��qT�r4�o��H%�чc��G�&��T�nI�g��r�&�;�Өh��q��\ɗz�\I5��7�~T�U���O�-+x|M�/Hm.�.I�LT
w��%�MK�|�7������]��"?J1�׼f�!��W�g��\? sk]�S���C����6�t&5��H��*	3
3=YX?��D�3���1`Fq��b��FI�9+	�j����~<͇^�lpl����@��f�%rV��E���"y������
�0o���w��sHu�sM��c�j��̶r8��>�5���eWp��`��훖��{r�sZZž�S���Qok7Ѷ�d�}���	�mw]���U:�j7=[ӂ �q�|�������2��#�H&R_,b�~���bp�1G~�Xȱ��C[��*��lgcY�f6�>���|�lYc�j���b��RJZ.�ke�̕�>�&�+�B3:e����1dۢ�~5��h��:)�㥛y��jk������܌߁Z>���_�$:� Me(���x
��1�3�5��E}8 n��fX�hN;��D���LX|��  ��?��[��qo����Λ�ډ����:@`M.[�f��P������j��T��$�-��+�+�Lq�<<هg�x+*Bb�.�ku�0�'l��B�L-o�g�JF��2^kۿ7��>�d5�Ǹ���W��XVt#������԰�<'�� ��Nr@7;;��WǤRh��G���QB�H|EK�Ƭ��Æ�K�wK�.�����.��l�frp���KB�v��F�̈́G��gA�����\�o$@��%~e|	�H�UR&F �tA	q���P˓��F�;�՜�Q�{�γHl�5%�Q������xi5�0��֑����k��i��E2~*Ef�&����c5�z�C�V.W��������i��]��ɂn��o�91^���U���5ߺAy���b��q��e�b��F/��\�1��lb��Yۯ��o��r�s�`����#-�``>��� 9�T��#ܼi�q�#=�s.����! �%%�����d���KW����$>�Ȅ��C3�Y�I`��bB�l��!����fd�g�6����x�_ռ2V;P����Ir��|X|in(g�hOēC��u:�7�׼� �rү 4'$~ARt�GF��> _Ћw�B�7�Du��y9�(h}���O镞\s������Nӝ��9RR��c�ɬA�|y?7�W���;�.ǬnWH�VA���st{GH�{��q��*���,���ۑ�X�h;�\�-fUby?�h[��b����g��H��&�g����Qn�H�����cB6��#��3:��RE�|ݿY%�,SB{π��L�u)\�=I�]�2K�~���U�׊g��P� �J~��W���.?���je΍<�i�;]�[�f���k���(���-E'W��B)� ���	[�q#ow�El$��6��|���e��ݤع��P�_��gQ S�)�Է:�dw�|j����$��ӷ˸Җ�E�X�Я�HS�'Fi�"�`J,�/��Vǧj<��C�����ׂ��kY�"P��U�O�É��e���o�E��5'�ƅ��1ߞ�`���\Ǆ����k��i���tP�*S���Y�(�'sJI��Y-�)	Sh�'$Jc����˾2g;N�����r 6::���]=2e�@�N�W��uI���O%��r�%BB.`�����gt�k&��U8O�[O��p��hf<96���y��e陏�b�E��7�$B�`�mȺւ�;䗽�N�t��l~F�B���������j	Q-P\ ��2�ɍ2 ����s�]��īS�&�d/�F]܍z�xR%����RԡgK��ӃF���< 6����q|{~}l�&���ǐ&q��5o�!�,����H�l�av�C{#i�L��8��p�(l�����c����L �Tˉ��9�
�����ru�	%��bû��}��d�o��!���`�¸�8�rN�����;�Z!/��+F���5+����)����[�8���	���r�����%�Gq����J��I��w̯\��;$����H��y���䶾�G�:k�0���\�?k��>�N�{(�����!��x��^���k��<�rϚW��D���^W?�����"('��sKdԇ�/�SQ��N���c���z���f���$��Ě���d42Q4�A���R��W�m\����� �:����mLw�\��%���d�k>�s��_;c��%@��ڈ���0��(՟�f�y7Q��f�f��E��?�h�ڱJ�������%Ǐ�u����!L*�W��s��H�Bw��n�~�2��ots��ݜ�XY��V2�_�����$��'�QRFv��)v����k�v�;��	��|��h�7�������q�7�O2S����-�۔9!y*�Tz�i�qho��AE+��P$o���d�PC�%�R-_��I�{((aoM��b_0����vW��L-fX��[=i���K12�L��������x<���#��{��A����F �[��r�����%��qz�q�4�.�][�<��a�����q)զ�������4�1-�8�e�#�N۴e[ ���O�!Y>�dR��^[dx�\�@�W�=-���`D��0u>)�u<��
fc荭��7������������{}�0��_��(o�6u��ed/�H1��+�E��X�F3I,���"ޜƽ�.�h!�q7�o�f�3���O��9���1"sP���s\���/y��3�y�҈�4�չ��K����"��>m�k�.w��y��jD�Ê&�,G�_2���X�p������� �!hE˃b{�?��;�;#�S�@Æ��í�������r���1�|��f�g���uU-���:�c/I������[y�O㾶 81 <b?G/?ԝXHB�,�����:�Ti%�U�`: �Te������u'Mk���bՈ���F	�\߲�2gnG�G�� b������>�+�6�qi	ZvR���VH�g}`Z{�"����W�bL��w?�n�D����@��%A���ENje���vP��������Y��^qX��f��г�M���Ʋ�ܿ~�XUŘ������G$�q���(�e0��}���ƃ��-�s�S�Oĩ̀Ie�h�实t$l詾��ŭ�����r&������4+ut���4�����,(�*k���0З\�ʓx�UXٲ�]�:Nj��b������Χ�Tʘ� 7�����Tl�s�J����߈�i*J9̒|mH!o`b(P�$e˱�.�a�>r�h�2�����/����
�?��z���)mR�ɧ�E�и5���:��,`�L/rMI4T���Ҭ��5�*c���8S�W�%�<��K9uq�k8��I�*
4tw�s�DaHq1�bz����3���VRk!�DXl����}�
��S,)�i�mҰ�;	���j��":«q�{d�@����@G�}�r��.�U^��Uq�>�bʑ�ZF��F]AN�dN�iO�߸� |R�"���}��.���]��KI[3֙(�	�:%�H_y�Ⱥ�H�3�p�2�ٳ��SS{� >WWu����Wh7��n�~i��JKy��fR�R�;ϕ�	y߂�`;���"����B�C;� r�c�
ѱ��Nr�O}��A�!�F5�B�H�Լ��Y���&�R�����|�~�/ �U��.�Qc�1L{�֨���Qz)IUV�A����si��5fB��q�� |���������v���lMޘ��Ё�/;O�ܸ@p���$�LJ[Es7w8����O�9��7��L��y�R9لwo��eS¶�_�B�;�bѻD[$�����[����x����D\M���ϪDV�w��7���[�LL�x.�A��]pP?���[�6�^`{uҎ���<eaq�(4���5�գ�����A�Q�ҳ���w��������}T�SX��+�t;e���O����ȣ�H�ˇh�`��z�����_Jv캂3��m��t����.:�G�>��,��#�)	Bd
��`jM'Z��X���Gk�κw1U֢��4/�x�u0�<v�Zi��h
�i�r��)���iJ�P��/�>U_a{;8_�Z��}�Q�+AT�QqŊg ��֊����1�Œͻ���5�f;7��a�y{foGM������i]�]U 6,��m�/�4rn �ӥʩ�~J������|�\$f`�7�/��i< )ms5�.]2B�?�'��\��څ_�+|���\p���4ɯ��@�H2���
�
�6��8W��7A�tJT�� �e�H#�CD�W�qp�jѕ:a�v_5	"|l�n���WW���S����>�s��u���Q�Ų8<�;0��D��iPiRR��FO�X=���XI
W3�z&����A�����.�)���J�d'(�Dbh+pr��*7�r�Chy��8c!iI�i��.�o�S�<NH�>�Oz���%$�#��ڝ���/�'9&��Ї5��Q�8-qԕ8XQ@F�����c ��������j�W��]`c�N_�2���Rg�@���Z���,a!�)c2��`�GF�3+ith�EI/i�`X�6�I!|$������@ԉW��?���^e��=�&"K҇�NS��y�j)ܬ�%ퟪ�ŘS��M6Q3���d�k��/�?���Oϑ��D�zJ���1�I �r���Y1�"��|��r�fh+�wP����BD��������^��>l[2:%HF� P�j�#g��c	_��߽�j�1�EnF�j���*�ɹ�����w��R���\fE�E��ͻf2hXY���աC�1L��h�j�ezW���� ��q`4�!�%o��r��1�{��YÂt�y^U<3(�nZo�˦)�|�H�)u��� (�=��p^/�pF����ǋޝ�E f�ʲ�Gs�CC sd�Ӷ|Ǎ�����.$�똩�#t�����ן}���G~Y�tA�~A�>�L�8�7ͣL�{��Tuz}�r�e�`"���"��3���C ��t�<2z`n�e�?��%_�Y���.m5�k���o�%��/#<V+�{;5�p���ڭ7i�T�v!����n�^�.]���9���y=>�����p�5��H��i,��]`XH��8���2��[�Ϸ�Ol���Қq�:�H?���R���߯<'f�>��p1�_F[H��G��E�ڌ���Ȁ$������*�3��Nt�y�B���҅d��H�Vb�PWFg�S���}kΥƂ����^��^դDZ�۩'݋�\Q�-�G�.'y3hӀ��/�d�ޮ�����!n�C�*+���N���T�u��wZ�
��O����*:�)�ṋ�C�K��
�߸�����1f������*�NE�o�:�E��8k]��R��+w�(�R[[�%�����4	��ҥ��k{�܅ŧ����Ӊ5	]�*����o�nY�68kT�!�uZ�בg�kӹ�'�
��~�li!��=Q��R��x�*���h�=����=
�(.'"��)z�[:�X���$�M7E��)DMБl0��~�ƍ�{�B���<u��?��_�{t[���xb��ȅ:_�%;ʁ�W���-�1j�+c�<cT�e��lF!���h�3I=���|�»K*k�T����,�ȗT�=<o%7�_�	B�m��v{p����e��� Y�?���\h e_s�D: g�"��	��f�"*��~���4������`ȵi�]T��"A㥃p���h���'m���S6,gz���������;T`l:|�ZA.1��|/�K��Tx����D���;����˞.�l2+v��I�J� ,t]O�C��� GR&Sj���W�9�B��Xđ!�c�{��ߵ��ߺ��1�W;�r&<��=��,h5�;I��j6����Ab�`����H!��EI&�e��3ǺE������6���f��ꐙzj�yCqV� �@ėp�$N�6�4�r<"[��A8�X]�I5�e�NAe�Fc02��#���/T�y缷�to��;�Gk ˺1��@��e-��}�@�{B�là3O˵93K��*��1���n-�J�h:���m���N�b=���?)�<OoMe��z�+㿳k��=D��D"u(���ߒpM��!_1oo-�i9Ec]�3������0�����lbF�" �V��-��|�3*���}�+��`�DO��n�[\7��� �m '�<�~j�ӈ��\���>㽝&� ���f4>��Mdޥ$���'�xX�AU�$T��̄�N�b�B�ϬHT�������`��lc-��[��)S3M���]�ο�W�K�".'ˎ]-��ap�?��_ K
[w˙ꯉ$�s���_����#g�n9��'[�#���������M��ro��Q@�5X��6��Vr1Nᷧ[��RS�It��F[���E�ܻDֲ9	�)lr�?
/<����_�Z�S�2��"��z�{˶*ag��q�c�Tm`����J��\�n��*�g��$E6��$�h7��z�?��H�"G0 F��i��o�2�i��j���sz'�6�javh����Z��3���t���>���9��p��>�?�ǔd�� �5��8 J1�\���v��A�>��c���=i��j����o��V*�C�3���N1��uoPc>Jt'�����!�x4\Q��m����	"� ��k-���k��I�`ިd2�Dt�7.����[�?��q�,r�!�W�R\`��8xs�Ƈ�Y\rۢ�iiW�s89䖒<��_-�6�U(6<A��iUMN��ʱ6 QV��H(�8V����a{8iʜ��.��v>H�΀DV���÷�4�T���*T�*6lsY�קav�-�e���==��A�?�sG�&E{j	�������E��+��鍮�H?cq�$��$hZ����ж2�J0����+h��+y�`c��7��u�9�U�02	Fuj�����6��Z;bn&&����JH��F�UB~�$��ĩZDw�W��X&����V��}Vw>c����1��L5�V�Ayv"#Ж�k�B){bBݹ���"Z��"b��ZQIQ�B��~�<!���$���e[4������u��O�Lv�W�qӮ&� u�m��ez^P�z�a�r���X��p� .��&SJ���C#22k��@��rK��e 4ZPW0�E�����`��:�x���Q���o��@��a�Ӈ|Vu��w@�#�-<4���xCrb�y�2$���(*�^��V�j��$ p�8a,���oT��J�L15��-ǎV�Y�m��\��Hm±Ԝ��p�4�z`b����g����!�'!���S�E([�n1�4�z��{�ũ�*ab�^1J��h�1P[D�f�:Ba)���\f�4�h�C�x��`��b�X;w�Z�"��%A��<��[;ֶ9ً�՝
D��평�`�Իb��th.0���$�׀k�P�u�%`�F�lP���e�9�10y�K1��R�?
�\�Ԗ�Rq����q��|j���d��ޤ����K~���}u![���P�W�� �4c��'�0�"�����71_�(Ǖ
���QX[�+P	l,[;�b���y`�����u�sN8����s���F�!�L|;ƣ�$��u���W">��t��Ԑ���=���[�
VE)��bc�0��|�:�dnGi�DcDE�`k�j�6(�q:��3�:��P�����M�9�
 �Qƞ�\y�����Msk����g�^��[��E���*P��;-�`��T;#�$%�x=n�:U��W��N�[mL���%$ oР�p�3.�~z�S��m�'�棘c3���r�FEk'��P�uN��z^��d{��vl=:m����kɮ7�*a�`�ak32��]Nm7�i�{W
��� ��H(�a����&s�C�;WP��!^��kpa4yy��
z���ią�T���Z�Jo��9�ϯ,�m-C�r��Wyl�Y�Hn+S"�#�3]��
�5�o!n�7�/��T��oFh�#wn�������><M�u/�!�C�"htY5s�*��n%�9kz8��rvm��B.jnm@}˔4��Y|5��r�Dv3Fn^�Lϳ�|��a���HU��)�G�Q��{	�꟮y��0��+0�*�؇��?��E,n�
P��k�B�]�?S1�U��As���%Bķ�CS$鰶K��@U����1�:Ⱥ���M+/Ҹ��5�.�v��΁���6j�U���4����A<-��M~(j���l�>��94ʤ;�Ӭ����W�y$TZ.V�(��{T��Fvq����&�.F�fE�d�h�Pm�\�_Z�lN��7��X{�aE-=�'����@3��{2Y�
�&q�le�* Q��w�#\'-�xc���6kܾj���#ߙ����'~�;��6|�6���U��ϵ�J�7�����c�e�A���H��|TU�s��X�� ������g���P�Ş��F��V�q��ൿ����罂�^OY ���gA)mi����s�j�l��,���O~�L��9�Y���va�je�7ۊd=@r�f,���'��\���Tx�e����H��ޣ�54���_u!��<w*ݒ��ӧ��g��:#d"�h	ȃ�����*��2��n%/,~dm=~H�t�5AMNZfR	kn@�P	���~�|�^�Pl�X��c�ic�_�I�q���6�0�͑�~#P���7��u�fYģ%ow��V8ԗ9�r�>, Q�Y����)Yb������>���3���Z�]��͎��_��F<sbaP� ���K*P��#���:�5��:]T�&o&���=dc%��;�Q��H�2:�vN���ր�F����p��>"�ʊ���1�������(���E��D��C�v�~<��_ѵ�D�S%?��T����IC ��m�/�>�@QD�D:C��]G�j��£g l�Z'2�Th����|�JzO��%4�?��j���WZ�BC�1Kp����L��W��ǝ�9-�'4��)P�&����zˊ�:e��YO��5��3��i�OyĢ�<c]=��d��������NY�wS�z���� ���6���5��z�V`�=�
K1 i�������ȍ�vBl{�#^��}��P	�;c�erۦ'�"R@��l���~�w-�+���5� ����(th�H%��ڰ�)Q\И.񎯍�x�69'�$x�T�٘R�_�,"�����u��/&�f
���i��������c�5�_s��yo��Y��KI��
��1V�sQ	7�^���yab�{��}�<����{"{ޫc0(�g�j���o6��d��p%����U��oN�i�E&�l��<j��&�g�4�ղ�雨0 _�qo3w)!(��͠��*��!/�鈏��g�?�t$�#7A`q�v�Z�*u]�'�l��t��6�bK���%_P��*�:"��FdjXB�5�Ay\�q���
8�lE0�!���h]XR�B���� _��>y��P���4<T��xM y����o��{R�j��E+��w+���ޛ�# �f#�|C�Z�f��j7$hYY�Hևg�D�?���8�������^��)������E9~��"s��<u�)�@b�3Cn������vjxʎ#�[�M�t䭉��6Y����`ܠ^/4�3�c��x�5��XZf��n���O��4���hj�k��<�U��uj�+Z�P}���s�үWk�,�|��3�t�i���Nr����o��\s$�^C��2?��*�Ё�O��)����i�+�u��t��ǋ}6��Y+�Wy���x���'�L�s4tȧ�Е4�]��-�����7R�+<#�1�{�x"3{�&������6�8  ��.�����߃d�%�!Z�׋��w��K1���^|3҆9���!�*j�+�>X�@�r�����]&�����4�������ˆ�R����(�Hn�¬��|�3 J_���Z���/�V�9�[UU�ে)�s@
d,�e� e�߅˽�=(�Z����;��>�ޝA"�k���1� }�����h�>xy�z:��B�e�'U�Z}�]����2�O�������U����?��ռE����9��*?��{�A�ꆖ�̞؀�8��^|���Ӛ5=k���I��9a�L-!��i��mO٥"�W������L?����Vۡ��"�/� Qt�\hi�ݒ���<)�+��(u��k4ڷj˪약����U؇��~�yю[�6nW�"$L�Z+bj冗�&I����W��]_i��@C�&ٯY����a�cj���Nd$P��l�#�[]��(P��o�f`FP�����'�p�A����eW�`V�M��x���J}j��ic��������=TkXF�!d���R�66ɛ��&?�6�r0�GL�l�٢��c�o����tt��:�d�������pBt��{�1��v�F��=�� ����~��V�g��w�����d�Ϲ��qO"	 �U�ؚb�K"�ޭێy/�����f�J{�{I����!�N��)�D�wO@�>�o��������CP���˫�w�f��]��ε���lƎ`*Y�J�g��ݙ8�ƫ3d����W�应��"�Te���M�Ӵ G��Ǣdd?��ɡ�!�q�G9�Q�|�E1;��-���:��d�/��oןw�,^��%�N��X<|��X�^5�#��R=�D�6��5^T��~��^yy�G�<�O�oGt�ր�Xb�5�w@œ*��Ԛt������MK[�g��!<y�]��=�u�*�P�
��t���˃�<�֏W��o�h����v̟�z�p9iRNj0��ETI�8٪H��aLFw���d��M5@0Uo������[�wP �x߁�X��� 3��$�딶$:��)̑������@���M$b��H�,�V�[0��5��$��>�Oj]C�-R�v��ͿY`I��{E�Ŗ�A�]����P]R�(�ZO�\Nl����L('���s�d����/ɫ���c�Zn9��l��H�w�5r�9���g����2��_)��F�m��w�����L8�(fx�~RG�=ȟ���5ӿRت0Rk��|��|-2���mD�"��Gr��٤�[~+5��s��RsVc���8���z���p�3hGT���wVY�*?��2�F#-_[�"�7�}��@����<i?�{"֛�wul�K���~S!����رzا�/��T\:�N��ip��*�~��U��'�Sߏg����Թ�����JS}����|Υ#���{ߨ��֋��I�d� W����(Ro��H���cRѺ��Dp�"��&aU7����V��j��@U�v��.x���!j��}a��3�0��e㵵|bl=��&�@H8-CGp6ׄ�k۔>C�fhn|(Q�s�����.X��1n�Vi��.��0pm�����tE2�Ђt`ހ%��9����>�͢��5�9��c������@z�7{�R��
ǀ�r����J�o�k�D�u<��,���G2�u>�1����5!���� 0�v}��-�����H+��������7]h �}	�@��ZF�Dr���<�A	(�2W�oFG�nJ�:<����1���<�j8�-Q15�*_~j(M�߃ڗ*q@��K��_M��(� ���E���~�<%�Gg�����ewo�t�Y�� �B��>���$�X���2#����T��{V��>tk�nWo�=�#��� ȩ��.Bd�)c3p�t:�����l�M��懩n�$�
�/���\����@9�.� &��ś���Q�=�γ��2��q�0c1F�Z��G��հ��Ն(+i��!f��3�SԲ3ΰ�,(�������"r��Я���ԗ-����4qʀɫ�Lbr���&F����>E����r!i<���ŏ׏J�\�T���6G��@�./��hX�]p����������t��"n�0¶-Pp���l\S�>C����3գg�Z��v� ��BmRc�#��{�'!v���<�(K;�BD�v�"$�q�0C��ޥ�7[��X��Lͷ~�/�W������3�� !
Re�o�����)��;��(@�ڱ��6���g�)�Mm�-�Ƀ9B��y��.�ck��V딐� ��"mQ콴�qm$�����N�rr�a��vXƿ�����2~�46Q9M��n_����6F����,�,�Ȉ�)�8Zߌ{"֩V�i ������чl2�U�A\7�k�$~��x8\����r�$zv�ʠ��n�AC0��U�	�h�Z���z$~�I��4;���'���\0�ǭnH�/����o*�Q�C��,B3�B�xa�_�f�d�'<�?��ݑT�����p�}���SK��@�X��ןO�,�EH�|-a���Bk����g��x��[�~uS���\���nN�Q;Na�s� ��T@%�G���e��ѱ|r��%k���S2�\���H��($Ѥ��[�"��C2��<����G@ ��
���o��U̗����D���5r!?I��<]h����`E��%�wZp��yw?0��mpK��=�Y�7<(���&)G�]������}L-IEt��mC<�9v���Y�ww
Ϋ��q_�O�V�`΁'�	�o��h+�l��0�D~�m�c7�ʜ}V�c�[p�;�=�߳��*��%���2F�����JRa���m�A[DV����1��ae�7[��-����E���v�]���QKd��J��9�P��h��ǁ�4��P�N}���{C����������'Y�q���|t��SH`���=�>O)�f欠���XaR���Eu��9=5���C�U��"CE�ʍ����Y���W�c�@
��TSw`�@���62�nU� !���v;�/����O��̼���S�/rj	aޒ��Fҹ�l���h;d���\�(X:�6|?E�r����y����2+4Vg�Xx��bekc��`H�����vIʩ�q�O��Cb�T��/�L+u�k�^�8��|Qzq}Zq�2��ǾF:ފ�����=�����IaqU��,�"Q<A�BL���y$R�ԇ2,Br�As1^<�T�(D�C���M�6��@�������K�:;:�A��6�L'	q�и}�&�ތ;j�Em�I��?��Ӹf��h�+�ޥ�y�yͅ�9AO�Ȟ�B��3�������e���G=��8�@1��h��]YZjO�:�0w�2v(	�r>0��}�� �|�?�R(������{6�/au������a:E��ka�94�awwf���?�.�4�N����u�a2�E7����z�N/�c ��nl*Sӫ�a��9��	R@ӇV�ݣ�8mr7����%��ڵ#Ѧ���Q@Åa�U�����װ������_��[|����M���Ta���n�/Udy��~'���Z��v�����pw�� u6���cHAp�B̕\|��XcG�/-�x��<S���_�~�7�9�I�k<�͝)�(�CD��Pol�Õ��
��,vLX��!� ��I��RwXD��hj54C��= 6M�P��sJy�ܩȊu�E���At1n@i��]�������xf�Ǳ�v�[7����^: J&_�D	̎�6IE�#�l:8](	����I:�>�T���B-�t����u�N��~q�}���O�QR>#V3��5ƍ_�)��p�Qҩ���e.�L�����:-�ؾ�"��3�l���,�`�T�
�����GB vF�S�m�#�(Xڀ^-ʛ��Y�B�g������.Վ�C�wC�KpMc����x����[�':�=��(11�7t�W��L��o��E�@<9Vn����x�o�;;f�!�_Q|+��ɹ��)����q����;� �ۃJ�y�Dl�@
�1a�
��֘	��xw:0Z��Ak���
a�uo�����i�(����OCt7 ��{ދ5znqc���H��xE!��W�� ��׿{uK��pbܵ64�]�{�» ����|�����a��
�����HXy4ض�x��~�Ѧ��_5C�����Ͼ�ڀ�}���F�����N��)>�$X8���k��	�Rb�&�(��3��W{޻<�kL(�)�ԇ��Ñ�b4����-����"1V���kP�q����Ǎ�Y'���6�?��b)�n�Y�N!��I�%�Ncg���[(D�!r�����sʧ���g��/�Z��R'�-|�V4��4�r@�\0,?����K�MV���K�]t�~k�O���V�����UN���z�o���r��"<�0p�x�jO(�tH^{=�Iͦ1�Uy�!�&� �|)�u��9j� �[���5����M�ZF�O�^�plk��^(d·?`"����h�k;z,4�6�;���t�.�����	\�?�Y�����A�y~"�����F�:����)��f �wp����f.]��Y����5��̵XXB�u�^*ܘ���]V�h��r���2]Q��7�N��z��@�fz�U����ґ�a�ʠЊ�2~�}��#��=�)I]d6�lZ�7i�$U�+�R���*[M5Ī>1��f"�{Ⱥ�DX Rs,�ɹY����L�b�s�$i�Z.���n�e:�ĺgCέᴾ}�(���%b8����-�TuMr�>�d�lV��]�}?O}�~>np'T�#"�������H�o��,���c�d�s����lY�����z"���1Đ	���Z}pp~�W���W[s-�i!�S#�7ʓ�/E��.�W����h9�f�p$���Ӥس�Yד�r�c_�K$^�������tA!�)����i�t��jp1�V�
[�`��[�z穧��[.��
�A���������H�qot�_=4eb} 03(:'}�N/����C��W��VE��m��K"�*hWԻW��@�!)����8��W�#p!ܞ��J�	�M5�J�ܶ�1�ἊX�
�~�"�O!$��+�!�^�
[���W��ȺT ��M@ �b�i�I!��R���?Ǫ|���tR���T+�$�#�:ĕ���..�����7;�e�8��a�_`�fDEu� �>9y��]��*����:��#N^�ӡ�N�ΪY�ǯ1��A�#�3I�3�����X&�F��e��l��P��K��K�;�M-V2�:�^�ֽKE(<������,D�P�a��8�M��p�S�������~\u]^�\/'str�i���\�n���<�ґ�� 5��P'ccm8e����ݦ%x����P�B��?���wU�O�����v�U5I�;����vsM˂r����t�:���s��y�=mL�0ǆ��Ѯ�'Թ��}.�>�%fO�mx�L��	�T1=�+6J���1�k�����|��@>��4�lS -�tKf��2Dd!EewY�� ����4�|/0I�nr��6���u��O��Hq��N.���x��9&~><��-�"��>:�H� ������/�UW��o4+�Z"blH�������,_�	�.���e���C]�p7�kڈa%�r/�Y�q�Y��
�YB ��kKP��K����/�L^CWD�l˅��>"-�C ��=�Ad��򉹀+��{a
�&��dDR����?VG<��Wvs�!�QOu
��݀����
�</Ҭ��pg�����ߊ�D�W�u@{��j2_�_/M4��[��Ԟ3:�Mvx���(�c��������#+�P\�Yb���ˑ�� }�1���"��SGr<���!e��| ��F�b���"J�Ʈ�G����d�% �#c@z�����Ҵ�P	Zu����E-���M��G��n3���1I%m��? +�C�/��^֪�!�����6wK��w]��V]�H?�4?��E!�9C�^'P��G���_��G��o˜~�'59U>�Q�����(�m�U�\�#�8��i� �~���<�E�%�Y�	�61͘��"EbS+�١�~���Z��m'����O���)_�U�0jWݣ%Y�v#M�RYC=dY��� %�i>��~;Qb���t/���wY"��t�
�+����w ��=���S����X�$*�ˣx������W�``v}<��L��k&��.���Ҩ��[�>��������i3ׂ�毈�W�^�3��h�q<�DI*5�.I���L7͜φ�K�?-��O��oݓ���}ka4DE�';����p��V('6���� ?��ĵ�'��	+O �_e�y��?�l�Dk<��c�v�}!���DqF�G�f#���^���Ȥ��n���s�3���T��TL��G㩕���J��Un ����V�|�0� (��V]�ʄ�ҁuGϵ��n��>�b�����@ ���7/��)��F��/��:tZ�S��W���W�QYE������kTh=6]2
�WP2��z,���$�k�ҳ2L��ܲ���
�U�t��?���G�����1+�j����#H��t�7̈�=�ŴŐ7E��ӌG�Ye$GI�*���u*&,EA/:�Z��R����f�/�3ג:��vݳ�5i:i�;�p�I�d�f>����{� *�̡�M�|=jϞ����<y}��	���k���!r-����|����Ӻ��e���D��R`����=�5K��:�Z~W��&���w˾�-mR�l.�ZP��^N��䊍4Rƣ\۰�c�5��LApŷ,8*����2�j�0�m4�
���*|�^;�8���ȵ�O���p���9�U%Ye�E��B��`y���J��څ{M�Z��H��Lu!���}J�4ֲ��֗����+��W��9�����L��c�Y��m��/x)�T��7׼sf�Zn�SD��~=���=����0�l��g�>�i��x��G��:<�i��vO��o�-�X��U��W:8�h���FG��z��%嶗�mS���� ?�|iK��4�gY��7)��S���1�	g�(²��Wk��� ul�4N^>��<�#d��)Xe`�ď���C� ������#X�/�~�=�:h؟�^�(i<bV��z�,(!������W�����.ɓ��S�/k���b�pgw�?WC�7爐�JJO)4�ԇX�=���~��v���f�$�N�b��y� F�𙂜��=�Q���vnL�	=T���渔�E���\�B��E�>|#��Z�٨���m�L��_pjP�������0 U*C".�2�FJAX:Ud�I�b��j/�l��ݯ�[���6�I�?�)>`���@������6-�4я��%�g�19ً��c������|&�G/��s��M,L�3��3UF�Z�9E�1D�~Vk���"���F�*%��G��(J����Yh��~�>�1����((�v~q��*��q���������x\+Vs�s��~ge�o0d��-�aƱm�N4��6���O}��Cz:c����c��K�u_ �����X�S]��*��P˾�ۥ�1\�)|w�*�H`�W[I�>�r�^zHH�,&��&zË���FxϪ���P	�����gZ�ѫ�?�
A�XJ�����6�_���� :��)��C����{�q�yM�4�RU���7T�oE�d�"�@��K��Y(��zN�{@U/�����I����U@W�����ـ'J8F���J�I��x�5 0�����Un�xr�N�EL��d��u�\�(0�YȎ���1ʍl��Z���;h*ީ}�_��b�G�MN^g�S�p�R�U��G]@D��dғX~k?ۜV�<+
��[�����g�DgWM?��s͞�����r/�g�s��$3�2=u�I���<�������j�O�O���M�1�E
 &�B���*)J�I;Z�Dp3��<�N,v��VMV	J�4�(K��!�2��&H��9�̯-b���L��%�&��Ѻj�Uy���z�,z��[>�~���U��l�\�,W`���J5�|%��jA��G�&CZʴ�A�� �59��m'�6
����x��CS>�`��\φ�=���tڇ���L��5�K���G��!uYPEiT���vڨ���I��Tc�;��es��6d����?����������[�D�w�q=�R��U��_L��=q�C/A��J�f���B2;�p���0��)������J��~?�zS��*���� ��J��
hw�.o��D�(����bD�	ijӯr"i�j��3}���yjV�1y_��k�����Ռ�!�~K1�(���E�j� �;Z�Gp�aɉ�E���49�a)a�+!�~�
�9n�$+%d� ���X(���rf�@�]�����/��;�81��CZ�^�ݪ��x#`�*/�+��G�~��)���h�������ʽ%�t�T91����v��Z���<힤�e�PVH��A�!{�?1�)S2��<*y)��M&�~�m쏭��?��Pk��ZL^FD�=!*������C�}&�c���f���ǿ0UET�  o��r������ ���  N��d�(h��ۍ3�km������ނ�k r��i(2��rP���B�Qd�+N��d��ٯV;�<�W٠UA$�19�@*�ԅ��?��**YI�3��S��D�
��Qை�7��GZ!9Q�-��.�6�k�V����0�{$�!��~pl��;�V�������#��IM>�X����1�L=",�YP���Ԋͽ�h��'W��@�����}7C/~�p�Y2�����򭿽�m=�N���D�;D��*�:Z� 8
����Ri��4 ���l(j�(���,O�+�D&����5�ٟn�\�	��ʪ�Ѓq�|��Y��4J��?J�_
�1�+���*A'}�GO�ﶕdjV�(�_�-N����q�����[���=���`��W�<A���a6N]6�3�d��>ࢴ���@��hD�b'zm��n���	I��g2Gx4�L�*�/%�G�{�|����ƹ��	6\�M"�UUc�X�E<KB����3X,��"Q�%���V���!;^��kV[RA �$ܽ:���b�\st{D��B�Gz��c<�F��\=�@�]��	����2a�I�tbf��,���cB 1M�{���c�eX桵�}�O���f`=���L��4�]wd�M��u	������ ޲��pB����/��s�����������l�X=D�D�ؓϟ��7�Pط6e8�<��f϶�"�n�zl�>���̩��).�4:�5c��J�;�	�6N@�|o}�]�:��~�+��0k$F�Z� �s�rs)��gmд���=�{�L�~�!n�t^)��Z�y���u�p[{��	��/��?�pyI~�����[�	f�[�[҈��	d:���I�*�Q��sRs�7W��-���{�w�8��nd�N��;]�'ˁq�
</J���!�dOاR�-�cdQ�Bhj45��XC���"K�`U���fAa�����lP"�*k��C4����� �?�B��Q��.O�M@��<��O�H��Ja���.Q�g�s�0�Y�i���#�����3�����-�N�D��lU�����0P4H��4:�O#sD��r���x�"����#���V�(ۼ�&�����n�c�}�+V������S���Xg�ڛ-�����3Ъ$�L�,�-#�����dV����T��o�yũ�:��/��MJ�9�\l��L ��X�X �g�d,ͭ��'J�X%���l����s:;(T9�p�0��� M�������i`�S��c �-Z
X8��s�Dp���=%��J�IڇYn.���6�s�|�ǡ+��-g۞L����DxC�p�$c�X�3LOl�{(�	�/N���}V�0ƚT�#�:��j���f��`��S`����X��޾%d'~϶o0��fN���k�(�8�:\�+�k�P"��8��ʄ�t��i"��:\
���C�Ґ�_38�����@5ͩI-���c��P1����T�w�8�m�����?�F*�V�kA����X9�{���(E6?�F���zz-����i /u�w�L�%����Hp�0�Ztk��;�	���zd�r��E�?R�r_����j�N�g��;��3oF� ��Z	�����9һFI���q���_�^�p��sº.�ܯo�?��B��Y+X���"N[�.����z#S�S2���`	�i�f.F;��1Ҝ�I��K�ně���/�Ǚ�fW�/e���74��XN��]`�f����e ��'%�6�����UT�]YYQ��{@ o*}ƴ�fPT������.Zt��<�B�X���9Fy��?�ʃ��ß��� �՜F���m�`��rJW
���iY79���Wg���/y
�Ot��`$zo)���q����ϔc'�C����ªW��@�giդ�VB�=��r��ؘ�ȫ"ʕ]��kS��s�y<�D��)R�����9o�#J�,G]!7�o:ٹ�S�!�8�;�k�H.�|�E�u�J�Lf+�]] �-P�Q���&K�w�y��CA�W����F���y�O�!�{���a�~�P���B�z��cS)�0~��s�(9�M����ʏƻ
b�k�~����1�&����!�YyW;���P�����r�_�r��Kn���j�`��� �I�|�Hac'u~3h�!�f�437���Ot�&��ٓ�<(\@VuQ�����~N���˘���e����HG)��W/	�,�H=��J� O�v�.}��c�P �V��{�-�I�����*/�N���Ľ���$�f�
�	#-����21Z}r!�MO�(u�q��c�w�Ʒ����S���WN3��=jt���tA�(h!���z�<���w0��hͯ{�xW�݉���U���J�:J�7:��g2���C��8݈���}W�<���,"�.�������~^l���̀s����ư��~���Xb��",)���C��228���g۶��W�c�[���_EEl���xRyf��O\�߂F��a�����Q����<� ��T��@u��� P��M}��t������rZja+�����@CT��y7�oX��$��[��l	=�h��)z��FX��S�i�ӈ&
��!p�HnVUr�Zª3���O+�䠓��$�%
W�2�[�������Z}a�pܰi�u�Gx���7�0�(B�hI�^����2�Jb�K����z���v�����M�TTr��)�q������2��^��-1}��#"I<t�d�,��<���t�m����+���� ] ��s���šN<�2>^z�c�v��b�����P��~<��i����l���ϭ��nLo�<6bu	܎3�$��(^������Y�|�R�$m$�?��{+G�Jx������r�3�r�{�j���Ќ�5.����h��=�iiCU� ���O�������C�h�f�G��O�/�Qf�U6eۤ}'p+���o�f�w�Q�DLvb�K�!5i����iW-�l�ɣh��o� �Кq/��!��gzv*'��?�����b����{u���cW���v!y꘏8s�[�����$/D�?2��٫���$n�ڒA�/X���\�*,�Y��t��`s�ύ6S�;F^���3K�^ԕ�Y��Ԭ�TtvWv3U^��Z�Ƙq�[/~�)�E;�/H(3���41�ٌ�̣HG!�!'��]�fO�n�����������Ko@ yu[��M�{��1�Ұ��1��O�[e�Oâυ�_��-6���-���Z/i��Å+���U#q���
��0D����O;~D,#�LK ڹN3ԑ����Oy�k��Q�v(������n�7]n���a������e�\�N�vs���c���Vm���.��R��`6�!�������CK���t���"�Y {�y��26�Skb"A��#�+C._*�ԋ(�.���$O�c	����z�7b�.�r���,�^Q��V���{I�t���q��u��c-�'�I�p�j�����+۬�S"����`�ꯠ.}�7�����FDI����vRKN�pA�
r���Z��9� `�-�x�L1=pǞ�8Vm���HF��?��X�S꾋nH0H@����b���9J�?� �!>���@w��#9�^��E�F3:���R�8}�G-���b��Wh��zp�>Sf�/toA�JO�C<���h����DoiƟ��ˢ�����G���/e/Ӌkԧ����3F��6�6�FS�{\�/&�1"��etB��|����n̺���2c
:)ByJi�M,��L��7/��8�H�H5-d��7F+~ѷع�9�ǧO�W�v|Ļ��)(Q��ם�2�P���;�(���e��0J��������Uoť�dh�p[���n�?�e�B��4{��D35O!V��5S���3�n�&��J:�h�1�	�6�g;-��
�eA9Q]�+Ge��Q�g�p��r�#˫P#?^��B��UCJ`�r	n�'ѻ��ӴV�h� 9�TF	"]Ԓhe����a�k"'VhA�v�8'6J9��]�:����{�S�Z�9��"�yw򳲀���}�)U�7ݬ�P�j��'_����j�W�}˔�n�M>�p���%����;;�П%��mv��+�x���c"�K�5a��kB�>��|G�$�B9��\/Nl6��"���QA F��X�*����qYQ��w(ׇ�Xq�;q@鱒?^�/�ړ�"oq؈�i��|ɹ���6n^�LG�(���$��L3)*��JY���b�5ػX�<h�S�w�v5<�	h_Dl���o���G�_d�H{��V>,� ��q̰����/hV/]p]q[ÃQ^�˝g��11>�h�H��v��T��>(�d�
U���i�� BV/)�t��Dmٲ�x�7���^[�3�Fv�c��Qӓ����]y���B�s�����@8�)���G:���?�pTb�u����D.�Ft�9^-�CBwr�Hm�*�V����BS!���U �^J�ʩ�}c=���X��Ly������zt�N�#�dU#��b�f���[�~������۞X�4�L��*Fn��٫�
D�=(�Vl� �i�J�p����7�:S�r�~6��0��(f>�J�#;rI8�E��1y�d:��5���ұ�>|��#�iՆ��e����ϯ����4�1g�l��TK��ei#���H �x��
a�)8��i���	k�'AJ�!NW��bL��XG78bH�	'�jxbE�uNk���6�@��)�eA���,S��/���J��L�1%@�q�t��!>���f�y��5��)JV̹�F���	�)�3��(�H0���Ŕ�[\?}��&�Lߙb��?֘���j`�_',ȮG������jO�i��I7�9=:�����F7kҝ�I�Nd�3�<ɲ`b��ѤF�$>�n���R��i�H=�3-6�w�r�F�A��,�T���LQ�T�S>���T^�8�X����D�r�<�_d|�J��V,�O-�f�c���W;N�{j錜i�&+�}T�ᔞf���>-J�c���#��u���ڴ���~ 8r��[%�6S�;�7&�l�&D��i�.��;&pc.�D[��d=�.������V�( zN���ߢ�e+��ݐ5�D�zsl�{8�o�3o�ק�7ޥdJV�h�>��p�!��@�������I#S�\~�v��?b�����;�8	�.<�Gm!=�}Re�A�v#��Ŝ��d�� �u����UHrl4�q��,�MG$�C��<&���gJ���|�(�*>E'F�~����9���&����c��Z]0ىV��Z�>`�b�^���=
�����LGD~
^�|��k��ȝ�|���K�)Le�Fqn�,����f[ �1>m���¿��N��ƌ1ׂ�^�̄`�r�J�HnNm����?�B��F����qYB3szr?:���G�{��A�-��ke���L�ڦ�-�xJ�`�)�T�ҩ��nç+�������B*d�Z}��v7�ȽV��|t"�l`���e��q�D�jY;2o?�O�����6�2�2<�V��n��͋Q�0ܤ���u����D}Q��6Z-�� ��\�z�U�,�f(2�h�UE|{7��"��ig�{�N�@��&囯4��+���!x���}��.��z5��1�?��̾���,U���~��
Ȩ���X���mX �݅o�g���+Ā�����SP��+	�ݑR���т�������"1����䟥ZA��.p
���I:�W�P�D�3a����RMO}�>	�ρf�H�6R���X�������1		�Z"9̴���=��0��c/Vޝ!Ve����3�&7/�T�W�W҈Q�v���އ�?m�sz�R�� � >^��0~b�<�Q8H�\��0΁���>��lЇ	��C�9�N?%Vô4V*b)D�0~��P썗����[�G�v�wr�y���Mtc?��Q˘޼D��?&.�\K����8.�y'��&B'��MK�jH�TH&�[��"2Y�:+ǫ'�m�XH9�6 �����bؐ��fg����P�:�<(�NQ�~�ˡ�2m�	x+G��x�%�����2����2!@cA��CO��cebj���>��Q��
c�+���۟�ujE�M1�Zd��y}e\(�16�qw��7=C�%NS�o6Qm���[ߘ���V6�%z�Y!�IA����c2ߗ��+��y�M�@9wt��B.XL8�ϥN�Wҵ�<�W�P
ٸ�LҚ)�ſ)��̪i�)
��ZF2��xf~~���ZQ����O�T"��r
<�_'��� Dۥ��5o<�{yg���Oe2gr��%#*n9��a��X;�8�·��H�u����!	���U�]y���:4� ���*R��x��G�{Ȥ���0�y7�6��&H�A���A,��$K:�����eq�w����j�	�K���}�<�=yA��Ģ=�DxS;���#;�T�?��Lh��Jf��a�nHH��vh�����cG��ɛ��9�J��Pp�԰�Ik�U`wK���X'��q�c�hJ��}��0�	h�4��q������&V<��F��ɢ��Jy���>$w��}�Ux�O�q����dhi�W�	\%�FZ����
Kuկ�<H��@���S_cWs	W�j�d���s�p�`����2�.�G���V�YۮVH�׈�������|�����=ߌ����9"���R����xQqRrś?��(��W���>ad�\W�U�h��z��Fk�]���[Ȑ��-��Xs������XR��-�	�]�L�d�4��Y�Eﰋ���_bN��Z,`��?�
�k�?�̴I��(�
�ڎ��UӜމp��"������l����ߢ�
��u�
$+`a��~;-K�+�t���r[�*��f%8��8�r�#^e(`�z��,!T�S�ąD�	x��m��c�;ʱW�C�,9t�-��+L��A�H'��2�M�V����EnLp�F��I����ܼ������<{�২B���_��#Ju`�%I,�)�J{�-K.��ѫ�D�&R�M;�FxӴt	
۴���}��Bm�~�@�����G*Ff�Sj�x�$��A�c�O��d��b+��,x�z��퀂V"Hl>��1~���IpQ6AW���m&�?Io�#�F�k�Y��Cwq�Ȁ��i�����˲���?@�KE0x,�{~��R�U���p���`n�q&�|Ln9�Ƕ��5Qm^eW �[H�N=��E�?bk�lO��.@�ٷ#K�7HU���n�^ʼ���y�ͤ�'�)[Y'�fTPkEJ�:mI�HH�*�	�&BQ;YΊ���g���H�f�U:�_bnt¬cy���t�a7���3��z�
�%�{��}g0Kxru3���T�
�t���F1�_H�n�s��S1(� �i��Znϻ�2�:U<��l�ghdw}� ��ML�pp��fC�a��n��n C%��I2�67}L��MN~��V<	�i|9��)�Ƴ���о�N'����/�t�g�"P���-Wɍ6y6H�^Z�{dy��s��fz��V�2q���'l��s�5�v�9z�������٦�#�ؠ.�� ; ��7k�?�8bp�T�B5ʨ{�6�"�(+;�����P��P�Áx��>^��5�����Τ���Pπ�'�!�z����'bY����B�+��\!,�e��˔��Z� ���YN �Bb��0��fZJX��Ҽ5,pU��4�����y��{�;�f��E(�9�8E$	�Zhu�U��VކO�����|��t�盺-_��`�gH���O��j���z+KH�O�,6�#5��>�.�u�BKT��`���}�:o�^M�h,2��_.����D���224I5+ad�k������y@0�j����\e���nX�=&D:ŧW��XO�hŐ�蜍J��L(*����i�R\��k&w�myLݜ�c����w�nu"�8O�1��u�g��n��N=^w�z)����-K�,qu�BH�q@e��Ro����m�R�RД��ص��9����ݔ<�:j�� ����8L�Tl�`x��,Ut8a�1~��r[!+�u���������|�OxDr���7R_k���{�8͏�e�I�&g"��Xl�.�s�ֆv����f��cS����a�<X�Ǒ�D<=��������x�I_�)f,-c�4і�w��D�L?�ER�ʿ�u�G���ɴ�p8GO�e���H�_���_TZv�6ڍHo��,h�A}]	�j��"��"r�y]��|@B��m��gw�(����2th���+\	k��9l��)j5��0��>���)@��DE��@��l�]�_�"|��5��r0@�\�>�0]�f/F�o������
���e��~$���s�������t���I���n3ų���S6�S�A�c�^��n�Ϋ�3��SS��Ś�C� ��bd��T�6���q֕S#���o ��"�i�����h�����dO_�:0���U㦺2͐p����BI�����y�R�������iM�����M���(Cm¶�ݣ�ӭ�#��5 +F;ה�Ur����bQc��x�{����\l��dJ�kq1���U���{�r��_������։w��p���8y���b�c_?��uɏ&�o�*�E�~��:qQ/}����m�	��Xo	Q�{_+82�/���9�t���1�tI*Ϭ�id���_�.�e�0���VDH0��̥�n�:-�s<|��8Uwܬ�RLbԻ������ ԋ���O��5�MQ �2� p��8���˖U�\\�T���22}�4����9�3�bB��}�������[�g>Wg�A}�4����^���J��񔔒lߍ\ &��&-�N\���{g�q�:�1�<�ߙ�W/�;?�B\5�M�/�#�mimUY���a�p�wT�y��"bK��wu'�68��Vگɂh��	P��;#��a���Ow��r�k�.���wѥf�[��Ҫ��82RZ*S�+�d�u�v�v�-+�;dV�p�ch� ��ނ�.
rm�b,?�U l�RlP��P��v.��4�O?�1��=�!eo
�Ѫ���,�k{}�Ւ�7K,�rFx� �Q�,H�B_���x�*��e=�̌���A��i"�4���d�%������
���ӃX��QM#z
0ņ۩k� ��a΀e���@���t<���=d\���-��u��%��w�W!��4��]�<��-W�2E��>I�[��?�Mj�w��7�`K:�"�U�6�__%�۠�cL�BI6�� H�:���ME�i8�_s�Tr[i��Rlu�u�y����	ŀC����ئ=u�A�#�����9Օ�Ż��lBANpNisM�'��
w�*6���j��tnjP2����{j:zG��k�Hؐl�MiA�J��6��ǡ��LK���"��TA�$�p���0�f��%�fn�zK�>P�Wxі�w�� ��	6d���ek��eV���w	 ��.��{��0^��`6�g�JEwwe�܏h�l��ڂ`�2]��E��{UC�������f�e!�N���FM�އ�Y��{~)"uH�W�n�fˉ�u�U�r��j�|D��f�Ɲ���}�0ط�ŁY?�e�s�aީ�qЏKw.�~��r_�1y=���Y�ˡ|�z ����,�c��2�0�m���M�X]oq{��+���K��	� mUi�Ɔ�vL�(�a*}j��R���l��_��Ē�}��'��)CA4�/!��H0��!���m���V^��p4�~D�,B@U6f�0t����if����ʤkIw�
��y���U1\�ȗ9h2��$6�l#.��Z�Ue6)a������=E�j����`&�j�w��"��z��8qpt/[�8����[U�l�w<7�I=�Ȋ��0^�M>��]*�za��<��0��M��
���u�Ht��0���y:@��A�!_��5:a���>��J�����gt���E���4$</�~/��]�T���
�� ����=y
��[�T�͢GX*O�6jLJ�.��V+`�`lb!W���W+O�����,D+A���p�+���9q�sJ;����ŧ��*������Q)գ��hp�� �֍��g>Hȃ1؋{�QЉ�/��.�<(o�2�+�۞c�h.W<3��}�<��H�DH�֋��s��u8	)V#�F
V���=΋���� �����c�:ν�lE��>NNӚÄ@�z���:�&Ԝ�?���	��3��Z��c���`q�|	��崟Q�@&�8�f&�O�/�O�İy��VfM�um?���cͦ���������~���<��=�T���p�a�2����IĞ��!p@|�=�p�u�if�X�UqВn|����b��>�!eh+�H:����L����V����{��s .Ӽ�4ơ��HV���Y�5H�-��ST�l�_ w��;O,�ձ��fh�g%�������Ѡ����o�Β��	�GiLx�����H�N|B+��\Z�?<��h��pǏ��}�3�WF�n�>y�	����+*]�H�N�6�)�D wZt E��|Tm¯���z��B��:�������'I�'7t��j7a�~)��	����~}�T������>��Y����B�������G<�W���Ȝ���]6��EK��з:.�����ݟ�t�� ļ�v��o"f�|���DK�ub��+G�d���|A�t:�%�����]�j��>;�֎d����^���5�x2 �*K�4l�Z_�����}���s`�4���dPz����&�G�Ip[ G53M���=nx%u�E����J2�7��	�$���:i�Y��FJx#Zi����@�$7ۼ1c,��z9��`�����t����4ц���.�7U}A���l)9�s�j��&u�{�@)u'�r�5=��N�9,.Emmz�ѡ�G�8(�	��D�>9��U�uܾ�8�FU����?IWn0���F�
��3k��_0o��@T�Qu݉�&�{y�Rܭ��	������ƙ�:�(�,2��s)�)�kK�%�}�������k�R��|��(*�#��N��f��'[=|�?e]���'��ʂ!�70�s&��:�v�c�����ݪY��3�1!���|����v�REGE����!�?�����}&�Ŕ !=[�"��+�M/f	!�CZ���z<W(����Y�������GnDz3���9��7m"��͝�����)��I�_�T�+��~���ގ�wXۿ�)A�a������k�:�[�j"䤾�v��7�唬jY��-�;n���[�wD�5�)�!KB���i_&��oP|n����88qQ���?ʞ�Im��;2��*p�G$���+"˱�tGF�(�Z}��=|��u|�eyG��x���]�w_�`4��YBQ
{s�͠k�!�5�7�t�BA՛��y��!�����+p�i�ak�NSEI7�"��xcq�;P԰�I1�a�NZ��<m'3|;ΝEы�����>n��f�-ߐ�R~�����&�f2�H�pѰ������4�{��'�K�i���;���P�e�Da�>*Z���>a�AX�Z� �*[эM�g�΁����ġ�hvq?�U�=�:�i��$��o���y��@�Q���/���WŠ���ϖ�9�V�dn�ޞ�<a��o���E�� ��hP�j��z\$K驾6�3�b�x�� �,�����JJޞ�g!�#%">[�Z�W��Z������CoW�Wqp٭�\}�?_��w	ݿg7�7�� �?i�VJi�e�
6��5�h�C�ӓhgDֶy|�H���YR�m+'1�S�`L��a���f@ڧ�ߴ��v�:��[�w�胴��������Z�6 �Kj��Ʈ�ڡ�@��C�Y�\j�C����T|I�`	�^�ܖ ��E�G��K�\^��A�"��l{r�l��g�7��5�ҝ-ԭ�b�ux�$�r�m�C�@Fpߟ��#�K��G�4��Y�7ξO�rƆ[�F�=V��$�R�p�\�qR ��y*��{����/��Z�U�-�/��0�+h�_�����!(���c����qv囡q�*����e�iǈ������2�2
�x�V��4��5{'�_�����Lk�Wlx�ZbG��I�$��j8�VP`��7xd�<2!\�µ�'��,���9�֓�`k��0�C��<����R���'��wEƒ��ad��n=��b����M8���S��Ob�)�X��q�6ێ�ܞ��-B�r�p�8ߐ5ވK�Cr2Lnhڏ�\��Ȅ���W��Ca��3ww2��k)���|����[�k�����fR�U>�)r -K�l�J
m
�-���Z&,B��:XLq"^�E��Y� �0�\�/-��s�ԁ�ݢ'����56(�bm4��M�)��	�����
�~_ф���-^c ���F��?��u��}'���LޒFa�j+��H�I-���V��{^��9�Ã6��X�^r�P��终N���i]L��u������*��_�B ?�#4݉�i�R�5�%d<z�Vy�k�������0�"�\M�GvI�(�y���Q�����]���K��z��F1{T*��:Ѭqs���[����h��b�Y�'�^�]UMA�}�6L��֋)�g�۩��5��%�{k�5hT6i�:�ڹu��Kf��{�]9� n�s��ݧ���| �ge����Vx��?��.ңQD��|��a2��O/^���M��������֜�L���V�;AQ�'O}vc���j����)'�釓C��*�5oM�sܾE�z�G����EH�m�������9u?�h�"���Vb�c\�	��r�i�\}���t�ր�[]pt���o8��2�̳�=)3�T���.#3��R���
m>\i~��T<�]-t�)�`�ں0�S����5�
l8�PM�5�l,�DL�~�4w{��l�?ʡ��oLgj���j{i�t��>?�+a�ژX)�8�uwig^��r���:5�^4���G�^d�Ď��F�p��;����3��ŝ�)i4SV`mg;X�̽Ǽ먇�%e�I��2�T��	���aO��7F�e���I��脷�%�R��T�W�D)���05*?�T�Yk���͐E�I��μ���)�S��m�ҒKU&?�ɋiϝ ��|T�:���X�{���l.mkF��|t��0aP�hֽZ�#����蟅����m�h'<b��i~y�C��4�{���$E=�ۺ(�4�̀$y��*Z��p��I�J��y [�:$K[Q��]�S�0���B%5����1�tR�N9����GD��@^��u�d��l8�cqħ�N����?صg�����C�����}�����*Bdh�`e;	�pH	4�f�:�m�=P�Cɖ���'�+h;�&@���i�h��;Sm�SM�?�	8:h��BWFׇ;;Q�d���6\��)�Njw��s�^\p�; �����߳���[ᷓ����ڔ(�
�]�o��	�,�����4�I��\���E�9=>�շbxF�e1�ޮ^=��������?�=�,����F?�3�'|����/_.��d������;�'&;2*�}^{�;7��1 6�d��D�WH�����U��ۚ��yK�E�p���v����)5HP���IA�[�K0{����zŏ���"�3%�B?��{]���������4�Sܤm̖r��E>��E9�.�5� � W��-�Z-~�DP�o]���+�����&q�4�&�m�1�:���KX�`=Um�5
����p=@=&[YN�cqU_�uF�H�&M��.v銈��A�	$��V[��D#Ν2���Լ{M
m
�_���v+,��RQB���y�pR�}O�sA�D�ف
��u��:	�n�in�0�:l	5|�S��fo���|�#$&e�Ğ/�+�_�9�W`�==7��|:�Sj�,�Պb�!�쥘��δe���VB��z���1#�I��!bAg��-5�eV��TA�`��Ԟa��&h��D�(��ͯV�S���4��P�uy3`��R�d����W"�I;f��Ь��F#x�q�1 �EF�_��Z���@Is�
W�C�-�R�h�[�)c�yQ3%��	fgk��]��%g,F�qcT��l4��z#��W�v5�w�|�ǫ�Y��Bl	s|���*nu�/ջoL �iT �x4�ʅמ�Hz9�@�P��6Ϲ����&�ڋ��]���I+����"ϭt� 0Z(�[	1��U�f�S���
ױB卜����b�u��l~�� ����f��~ΐ��ԕ(��z=�`?��"���y�	��?�L����wۆ�0���>G�_ig�l&:�ǡ���I:��Tt�|�Y�q��A�/y��"�Y����q���seh�	ˌH�Qr�P_�85 �f�C��xΉݙ�OK�P:6��b�3�L��P׸Ed�4��p��rv�F+�y��g�o�̂4	�Z&��`Κ���+K��sV�4'DL�� ��>`��HN5���]ҵ�Ҋ?5��19̤��pO�m��U5�P���۳�hԠ�?*7�=���?jּU�ئ���u`Z�c�����E����c��`�b ��0�
n����}�q)�"ErH���-�+����(��H�c����W���a0�x���i! 5���]���д�X㑪F�(�h���� �m�y�L�3]�/IG�7"�w<z��S[&�t���n�H�͢�b&���/r����N }���0���=�<"�G�W�I�N��z�����[�W�Ǉ�O�Ɇ���=��6Qc���{D�x&���ML�v���O�TQ�J�}؅���~�k��Em�2
�'?܏{��-4�=*��b����5�_G�,��(�O ��L[%�0��Y�>�oљ�ѩ[�2��X?��/�E7nn��¶���3Or������EO��[�Q@�Xϗ�la։� ��R�}g6Y:��t)"��0L����{n�������ZE�6	BĶ}�)�vb����<�A�x����ˁ'���ѵm&�^�C�� �0�Y�_���p��@�����c���E��6��B� ��[�.���x�CN�lR_w_�2��b�gVW�_�/(���fֹ=�q�<��Ȇ|y�'qW��xu�G���9z>�,FjL��N�K��� ^���5�T�oQ���g��c��A(�:УOm��񈧋+�H�e-qs�f\'��!��5itJ����qm��Xu�v*�\w���~֞�����Nl�cKO���h�;��k�]wȍ Tj溅�k����h���W ';�����|�����]�Y��!. ׅy��g�ٛJ�U%�jB��������ro{nXH�z��#�[@58�&�ɰ��?h-�?��f��{�8�xC#�/C�3��@0�ٱ�?����&c+z
�Bm�$�1a2f����W��������T>{
�w}Q�v���Z�f���DT!P�2 ��Q��⟷���"�5�::����d��P�wQ]�a���G�$ym�qSX7�f� '�c���'�g���b�r�	�[�\�!�}(��]�:���xy�Ի�B1M棡��Bw��� �0H�{hnFǟt��_�d�'�.��,}ٔ*I)�D(��5�w�[ȭ����z��95k�5��,f�k�H�.�@w)��vz�*s�Q����<T>����sM+"�Pt�aO���%�i��}Ҍ�Ԇ�SȆ�+�;�?�'z�'㈛F¬u���A}�z���`��*r
�?hR8�61�l��9��c���o���ٿS���H���<�Y�Ӆ}��c�,L��3�\���na=��ޢ�&b_�B�K�)�Ce���lx|����^��(��c�?%�7�~}A|�6�H�k��4C1������t��R:�5��~ha�/��I��.�"��������v��Y���}6FV,���=Xa��.�H�X��Q�-f����$�����W	ʍE<��r��տ��X0KV�����F��Qzs���]F�c���.��~�$6Sx�]|�=&����zv�����ܛ:y��q\DZIȇ�M��6���|p��{��|��,�Th���>�.y�X��Fe�O��E�d, �Tq�޼	Z7���G��-������ډu���c4���hD����c�݉�TF�����6)2>���p��:�܁��Jn�݋!�vD�R^)�}1���(�&䋜oBտc�۞�De_����Lf��x�Pု�W}ض0�M���3�G��N�~-����,�W#�W>�l��3
��Ga'������x7�Q�_j��ᚙ��7��W���F�|F�PɚW�E ����5T؂������%����v�ۓ�{)��m^|:�Y��[J�O�0��+�Q�����m>��"(�nZ�m�bP�ҨȜ��`��z	헡Y��9勐<�l4d_eд��0?'x��M�֢�������FPi�օ��#�i ��asbY�S���=q�l�] ��uM�o�=æ�Z��Y�v��6��|F���������� .�(�ȾD�����$~�,���v����m&�-�2�"-��qNaz�g��
	�П7�=⮌7V�x��ͺ6߅N0��q�Bh�<#��n|3 ���Z�v��#�9Mk���	4�8���{��/��>Ֆ��ztwpf������Y�)',L�ff�i���y�[w)�+��:G;q��o�!�A��ƣ3�X11l�X5�Kf��B,D!���!��&�~dO����q��l6�D�I����uo��%BL��2�LgA�x�������8�Ԝ	�s�s����~^_�U=���˃���ߝ��.� 
ч��F�ň�6qE	^����S"-�v*���I<no.�֌�#ӝ����d�E�:�ښW��Q�q�$$9��n�d+���@���R��j3��f7�҅y�z�6,���x$3J����0_����y@�0�Y�<YA��}��f` ��J~���|m��YH�S3^6��BX�߫��3C����M07�Y2hXnT�'���s4W�1%�Q�,�?J�����z��i�o��?~-�y5�N�iޅ��Ec�KT�Y��Mn<�o��G}����I2�WL�!<���$or�agJό=���H�l@1D�9��͙�j�S���E>�g
�# B�M��\DK�3���CQ\�\�3bg!��l4�ی��Kn�!�7?JٝA����❊;����Bdc��}��Y��[Aǁ�n�/�!樞���$u��a� ��6�P����\�|7��	��1^P�z����\�/�C󜋼LQ��ySz?kMkAn]۴H�(
�T�2�:�uݾR,G-gmR�#��`Z��ef�$SX�L������Cq�b�C.�����w4�V\�����*Vq�8�+��>��I�~t����k��u��):@kVB�\����`3p̼:��4�Q₵r���`H�:������陏�9j����]p�X��aT��c1�x.G�����O��PQ�měP��o��K�%��wlH��Eī�"&Q�]�� �3U�v�3y�5�N__g�W~H'��C�>sR����3���0~1��V?���Ȟ'?;�� b#U1���R]�D�;��=�<�3
�R��\�CE �	ߤKԘ|�
��H�>�k������b9�A	�O�i���4(L9����Z2�|K1PNa�FG��xu7E�Yqɘ��*]��R�w�a�@.�`�_a5"(��9��D�%'e��e�ն������Y���y<���b���z�Dh��e�>-�o1)g�
�� W�Ӊ&�]�f�P�J��7&��LȞ���a�Z({�j{נiE���9~���\?2�>��>w4�+<k���k��H�oA��IH�d�h�!�08�8�b����OX��~F�`X4�XP¨g��J�c(�e�0=n�?���;��ZSZ#M�.2��"OCº��7Or�,w��s.x`�7�D�x�%3����[3�/���P���v��5�Bf!�aF2��mZo�.��H�G|���%���6�Ɯ�c�e����
ͯ3�d�OkCL<H��)���̡Y�gK���']U!�-s>po3~��"@���/I�z�����)���K%��v���[ɋ}�S@3!�W4�	R�n���\�/�:����:�����@.Q��sQ�e���v/:I��X���-��a�L��,�PE���R�u�1G�U9���wV�-p6q�1qQ�9�d@0�����5�W�r���j��<�[��t<)�Y�9�[��8Y�׿JK&�O�5Ҙ=Aw7Ԇc��T���'��~��=���ک���e��h���вy2xzd�:�^X�e��ݻ���P�������[1��A!DF�:��I�_j�z1٧��@����r���d�W�m\��~��̻�������[�݉���a��p&n�i��7�\{fT����VO �v��x��MC��?��	G�:�pn�(Fa(1�h\t���-U��j��+��I&1��J�JBs�k��BJEP�sq8��G��ԟ��u/=��X"�Y�6r�^}�,��vX��}e_E@L��]��u՞����w<W���L�R%�C"7N�H��r��_J����Qy���1Kk��Tf��J �ƃI���I�yM��ky^ %M��-~n{	�����m�n�ր;�7mx�E6}����0��SB�'���fn9�V�	"��hP���� ҳ=�����s gu��i���W�W�O(t��Xv���2��;�0O��ݿ3��o�6�>r��Q��Q&��_C��<x �������v�|hثyk��D����1/�����w�sQjԔ�z�J�A"IuYʮ�Q��xZ�T�����U���N�tāJ�t9H,ϻ{!u����R,^,����!�$D�g�}�C��`��B�R��
J�����#WB�g=
	��"CC��zq��zi3GD��\{+�γe�/Y�E$�N|6��і�U<T�}�d�R!,�Zf�C`:p���s� �RIh&�փ�2o�L$�A4� M�p>׷9�.��2������7!>�D���������2���&��$�N���������nb��~ȍ��Q�%U���N'_%�yUA��Ca��q_1�{	���+��B�����5a�֦y�]#}�c�'M��p�Ǜ��K+���ejw����Ut�����a�@�� 7�j~�Q�G���L��)T����7~��"�q x���t�+�֯�Htl;W�}A���ǔǹਃ���=ٷ��Ȯ��k�1Il�=�u`I_a[�֋��	=����	�EL���[��ڏ6p����Q�l�t�F�߰B��-���}n�WA�+TG�g��`��Mr-��?׮�����"���2L�K�[�:B�B���V�PW%.@��;;�@�ޥ�W �<�UBL�a����߶��O��6+�mW�mmt���*�T�v�A
m�#_���޾)��c�%X�~��| �fY�|{�l(+&��:�u�[T*�\�.�a��r����<���K�m0���j�{��!a�o0o���%,�<��#6R�P('�e�fg!�7P����nȹ�z���N�.� ���|�Js�ߜ�h��h��7U?|7��2���u[@{}�!��}�u-� S�Z"/��F��o�|lqfJ��Q�uF�C����&�R��e��CQ���V5|�By��3a�j'���K�J�n%F�A�V~�O����&1�o�{G����ḭ9 �&�Ja=�k3	o��y���p%ٻ����ev�s�)���h��jE��
��9���5k�wf�]�j��\��MR��	l�A��;'5��%Sk��7�8������}j[���+=�H�ߏn�0W��ܒ��h����+��Р.Y,XQ%ң��U���)}��;��7�ˬ�hx���t��2����Ҋ�`�.�`�O��~&�.�S���)�&�L/��Ilއ��>3��0X ��,����y��� �K���r��=���(��9Je+�0o�mμ�j�	#i���������L����;���pf.6�X�n#K�Xq��n���ޖ%�:�NzK�'��5Ǹ󅌌헕5��m��m���1���u��]t3��۲���򑇄df���pTa���1���H2����T<u�{�$d�z�l`<�p�&y�6t��I�N{���V��N�3N�SU/�ب�9U)s�QAK�՗6~��?��!�G�j�k]5��{�"��G�}k��(��r�E��K/l�پ�9Г�y�9�������D�[&�����f�CR46��.����i-�)����p����Uq��897eU�6�0gq��}ږRJbA_��$>	"����EG
��ۻ����< <HW:�^M~,�{]޹kH0���]�Q�K0�m��3o��p��[�ݧ�@��0K�ξ�]���٫�ͩ�Vl�Ke����-pվ����k+R�4�z�����
�+����cO�� BB�qh)o7�G2o��}��)�is�EK��%3�w~QI?�ce��L�����y����T�M?���mH8�߮-x����H
��=L-��6�S�_�H��=�f(4z�|�}G�-7�^���\2 �Р�vA�C'c���W�Cƺ�!���������K���-p��(F���['� t��nD��k����f��%WP�82����u�ɪ�cO�Iz˶�c=����
bB�R��k��Py�Wv��Һ#�D��c�Iz�ȳ�(��c,�����"q�~�tЩ��e�˖�H#B�]a����FGC"B:��Z���o�2Q�k�M?C~!~�,lG��~<��e���Q6z�/�jJ��M�����+�A@�B9p<P�@П���M5r�x��H�9��S=������X%�Ͷ-���`��w���K�(��Zĭ�+]�O�ar������졍�4��`uǚ���.4�v�J�K��+/۫-0n3$�N?�yi�H�lF��cxˤ���: ��MV�Ay_�q8@�1�VQ�7�=Q�,Q�~��x�����Vj����ʛ\�-�7%�%��2�Ί�'�"ݬ����Y��*\��l|a���<��O��C?�;�e"�`4��'1L���_�V�.��Lh� ��#jO(�|�HГCp=�f���`�я����6�Y�C�� � ��ީ�?�Q�'���>ٳ�����ľ7��Zv$J^��.�٩�������9�e��# �}(�Y�%��*M�^<O5�ǯ��I�BO���MS;9���k�nO���M����%p�ڬ:[�f�Z�i-���^����v�iC{r��Ÿqf�	u���t����q��ò��9o#	���[=���z�4�e�RͰ�$=��S�*[����� ^����=b�/�ѐu�j8@ͽ�'Ff}�=��, b����?2֒@�"Tp�K䐹s�H�ϩ��5	9�[���$�g0E�k�y�u'R�ww�bq�����l���̕� �iZb���ޕ��0�A��ထ�SN�M"w>�qA�T_N�
�f�3����\��iB�^�l�����y����E$);�Pf�U��}KV�Ň:;1����TZ���AIn��ǁ��������Ia�)N�D�r���>����4�q��U��M���ֈ�홮�}�4!EK�h��(�;��u�y�\��#��n{������)�Q��P�m&|�����|D�p�И�}��� ck�4I��J���Np��Rlڂ:@@���� �].�[��;�X��^	B�ޏ�4�����np���fg�M���Y�,x���r�ۥq��m>������d�تg���l�e�"�����k�*���S��Q�|7��FK�Av��evN��ϯ�Z�sc�<�g�9GL��Οo�}��=�Xd��I�rG�8�1K_-g A��b����|�Ċ��<�� O�t}�?!tv. ���kH��W(��u�%�_?[AcҢU��`{~Ɔng���Tt1�<��8�6����,xږ���`��K�R�@|�9�'�T���)��i��w~`�L;]ᕍO���ŝd�j���D���Pɱ'�p���������iO7>}��� ��>�i�m�i��k��F�
:�����u�քe�q|tF �-�C�R�)$mg��X���%��L�#�plW9�]���+0	��Q3��N#�}�^†��q�������ܞ(�R;�.#n׏��O��0H���#�]|~#7����+��Ul7�&a�ʌ���7��ҧ� �o0�L�a6?c�����W>�W.�3��_�g�]G k�o,K圥W�������=D� ]N6�1�W"!#_���[�x�eA�0,C��Ȉ��y��Zb���y�\����7�Y]� N�s�5<�����4.��N�uR�$}�����4v轸���º�5c��d农�9��ھ�n	�c��Q�$�O���p�ŋ���[:۽;�K7�?5Y+��j~�wM�,��Z���k�87�?"m,{��bI�3�
�6�M��$G%�2��C=+�!{�S����JR�
�c���h`w3������ 	z��V<����Y�-����/��a� )_����\���	fD�����4�s�֧R����r�;�hy��^�yv"}�x�9����X)F���U�̷��~ɱ|yQ9�9~���e�������#9w5�K������M�0�qT=�*$PP��@���:	���a]�|�X���h��H}�����Xz��31�e3���u�ͬ��2� ��.��V�v^�!�c�6�2���u@�T�!�Q0���aq.���u=C~�Ux����^*�ѓ�9�����1����R�������lP��cb?�`�����,U��9� ������=�}SQ��m�E"�5�4� �2������$���rr-�:��t���3�e�vn�L*Y���b�^�I*O��HT�c�m'0��:�G��q>Kg���������;_L�e�)B����C#m�)�D�[ɴ={ֻa,��w�HsA�&)�tRI��^gF��V��Z4�1K5?ob<�`�b�.��Nc$�$-���&����"�1�<�_�^��^�n�?��EyQ�8��@J�&G6�[�1ڣA� :H�4/�[K��ѡ�4Yhe�&.���;,�G���N��K�-�,wp��ߑ�(t��N���w\��ޔ�}���iaG�ڦ�����C�[��<��m�@�X��'F �t��e��ћ�Ѹ��a{�Я���J^���̕�3n���}X��gi��
���h_X�%5s^�n��<�|,�R�F�ڋL�**���4O��yw�aA39�x�W#�"���r-��ӚM��=%�6	;��)� άI�q@�;�/sMj�`��trѡ����m ��
M���ޟ;GW�S�9H��oi%d��oUʸ!�¸9u�J�V	C/H)�R�H0�*_��	��U�9M�{U;7�!7� �o�3pѐQm���a�L#R:���Vd���A*|X�p�M�+�!�0/4�z�ͫP�t;��}TA��#V���ۜ2C�T.  ��h_7��u=����Ԫ��	��c�ټL-�f�4�-��%���u��y��v7��L�����G5�D)��|O�����=���P�_��d��腭���״��@lG5�~���-5���XEs������E�H�����m���5>��"��PgH4 �8��,vR�wb��坺v*ih��>8L�!>1��n�-��]�X��:���yt�f�)���ϬjX�rsD9SP��-�OPr+r�~����a/0�������m��b�}UZɼo�������Ne*|s��֘E0~�����#P�Of8>>A�5�#�q}y����?��+/�L�����8�C��2M��W���󙘷_��}2���.Td�eٞ�̇�e�֕\-��ɩǆ�+%�n�tJ�� ⮣G��W?�C_/�4"p�7�JV�|�������L%�RE�Y夒�4� ���/�7N@��Ԟ���e�����F�?4�&�-�z��h�@"P�WT��K��P��	>��»�	1�4���cV��g	J"���C�oI�`ށ�pBxu�_�<�`=w:�^� ���M$Z洯�I8}^��}�L�M����A��F<D��x�W���=��$_ r	��~C4�|=ȭ���4�<H�E��׼�p��kY-ikkGG��-�˛��΢����9���+fH�a��4�Λ�_5���ꠥW�h�P&�	g�]�^�rP��6t^�n�舣�VA���&3�y2J)�I掉{�8Bb��]����vj�>�GfX	�����\ݾ�&Y�C�xWV�p���Vo��P.]�`�>���VW�8k ��2�W��)������-�a��U��#y������_B��5�t�|2��F�)��"ü_<� K';�����q�/֯W
y���}>�T��2��&�H�]�1V�!p���2�*�9�c^� CR�צm���k�t�ƨ}���&9
�	3.j��o򀉌��;�X/���΢iX��]���`vބ��R椦;3����Z��I<v������گ�(JY �a2�븈���i�#Ha�#N$S'cGyCz���Ur=��y`m���Z�	��*i]5�gڻV��Cd¡�皘����^d<a=�J��"eZ�vIm:�8��fw�����I(��7(?�7�9d�m��$��4�J9-��DCRc�g��Ζ��!D%�G�K�w��m	o;fzk�q��~��~U�Kk֝?�9�e�4 ٺs���]�R�t>��o��@3\�ine�^L�|]��̏�,U��o�o����S�tRv�z�r�Y�?x��_�s��M���4>��o�
�&�1ܾ�׾��K�9ڰ�%��Q����aW�SP @�8~/�B���<[@��b,�<���&���xc+��\�(�c�pW�3C�p�k��%�r:+(]٠2?z��cD-�vb�Q�����j��P �^3�'���7䱲ءz�͢Y S��՚�����[�A���d�2�\b4	��&u>�'����H5j,T���� ��`B��
	vt�)�����HtRpX�$6�����"�%�D	��ި�L�B��vK��ti�w,���y^����xa�SF��;Гye� c��wLP�ux
��~�d;�[�֏�:/H���}� |w�F5#�z�֍��|��O6ٞz���?{~o+[�*��Xx>ŕ�� ?W_��m�#K��/g�{�v�Vzh���f�W8ҕ{`~i6B/'��u�D&�9	a\���v7e�[XQ��=�kK�IBM�����͛��m_K��Eq����H7f��9"�*��y�2�-�IDL�,���5� �����V�p�5�W�X�ky�/n�aQ+O ���rQ�'	(���u�6��~Dq��@�F��;��J�@�O������p�{=�y�����nZ�)�ی�Xb=ӧw�����}&3u���+%�	>|l
�[�w��Qg��>���0�{#��jN���C�g�̔�*[���,j��q��i�V<�A�!|	����{4�
q�ȳ�kI��t�1�)�E��=�^{4S��|φ:��X�n�9-�����e_��Jﮋ	@���"ȁ����PĲ,U�Ɵ������v6aKŐ��Ѹp������6PI��I!�Zp�+Fީ��Q��,�a�k��$W�Ŏ����0��D���+�f�?����:s�)��8{�������>��T�3��y7~��j�����;�ƐW�>�*���w ���Tk/�������hhT�(�S��a��$� b<|z"�d21�+���1�&����^�1-P��g4uׇ�xK[��Z����Ǐz�������W��y����˅�N]嬑�s\T08�b����*��>��_	�Ɔ:�X���s�b�[,%�? ���.,��yކ'���[m��˽�)�'ː�TGV9�'���>���L�C��kS^I�n������j�Uao�sqp1?Hۍ毖��0���Luң.d�&��xJ��|�zuTV����|�V�r�(����"/�.��a0�{�q��֗��'�`NN�m���z(��v��+pQ+/����h�3��_�oR�.�c��
:Q@!�6���� p������+�>�x���=�I���M��9k��P�E7���]��&��e�a\��\��q8�@h�3y \�o�T����s�ǋx�G��˅F}MY�<{�-�*�EU�-�r�Mg'��G
�yx�ڒ�dn�<^~�WșQfI��t<K�tF���4�qy������B�7��p�s9���w��
��Xr�%�chv��y�W����iY���e]@_�Y����s�D;��N�}A���C�]���*|붖:㉛]�����c����{���5��r��Y�N�B���R���m���tڭ��no7,��� Q9||�w�Z�e�I�4	�1�V��n�3+N;�a�i�]Ρίw�9�r�Q^���]�NF�.OS7.��I-�`������G�䭒��_�<3��Q<3jIRA�aqܾ�7k6>\q'$�U��#���獃�"}8��L�Uވ�*;����-��oWK����y���dT�`jcܾg��9��g����&j_�c��`x��vPP�rwm>hU_a���b6|٧zѮ�$b����N+�?K��SuKN
���NA\�$�H%(��M*	��n6���G��aJ���mh��j�q���L�M�Ȓ�{��O�Q_�T6G�n�*�{�����f.���K,���P/%�z����Ґ��]m��MVg��8�(��k)u��v�ӏ�?d'����{`I�R��T��V�5���<j^cnV�E�՘��Q��"���v��z`�Z!�󃧫=�܎�(A�5+0�+�����Y���3�k\��V�o��Ł3/!,
~ܲ�P��n�L���j�QF�cG{�,ӺK�t:':���UF��(ZH�X*�m��	m&̀�Z�.���~�F�k-<�v����v�\�YGԫ6�.�1�����$�9�׊�#&]`�0O��ТT�*a��C�.��ݲ�B�&dR +B�������;�Q>	�|r9Y޻1G[���FR!�M�g?8x#w�i�Ѹߨ�X�(��B*�؄X���cׁ	H����2������?KQ?�0}Gy5�P>���Z�WĀ�M^5�krG��
����|&0D$d�^��Ta�3:�����t�)�&>�W���5�J^3*�B7ྛ<�\���t�j��ѣ?Io�k�쿣��Zz����Jֵ �� �ڟ��/��\ko$%�Ai�a��#�կ�!c��)x �mh�V�BG���d܌�:�ڒ8<�{d}�HT^���u����I���JEe{Y���R��!�)�!'��p�J�*�!�V��%��_���1
�[#ؼ�fƇc�NQ��fK0�'z���Ti�7iC�� �����@eCD<��"f*Ǎ�Gc.Ah��7[�rT9�9f7���tS�an.�#l��4�v����[W��U�Xvit�����@)��8zu�>����O��i��Q���T� A$h����Xn��K��`��jO?���*w�Slm)a�~�����;�d����Аr��J��MT��z`\��9�R2��B���>��=��޽�K�V4W�~Ρ��:� )r�`<���`�s%��Awݞ����� �����I%��9r���<`љc�9���k�2�^�L �I��|�* ��4��i�Rg�F6��d�`��$�Yjd@�_�P�M�I�Y��S5z��> ��r�Z:3��~�C�
��˿��ƞd���a	qd�Ы�\�coe+ ��E�O���`�h;��SZ���0�.�Qv���� r��h���ٔdڴp�6rj�O�=%�7��փM��w�Ԫ���`RI�(Ro���Ǝ��툩Iק
��XA˂P�����<�8I�i���i혊�:!�iA������f�.���B��JҶ� 'j]t0��p�8��U�z�wRC����6^�tTy|�����}R&=.�.�9Ϻy�9��z	*��|�̯G_}�!�]�h�,�2��&�3�#$��v(`˽T���D}��<@����-y[t�x\�)EH�֏[�-Au]9N��6�ԇ:y �(S
J�f+�8X�3�.�
��1X���/��{,���z!��@?_2��6� �e�S�q��m��\�^r����XK��q?�l�Ah�[����w����ʆ��X��q�sܙ&�ːg�wB�B�$J���~��f����ͻx^���?��h�͖AW����c�VmK�AJi�F�'|�؞/�(�0�LU�,�X՛`iڵ���A��"FqQ��W͇ ���y����
h��$�����By����&��O�Cd[��g%�����O�4�. %�O��������������������~���P�
ք���K�Ӣ9]�m!��'%�@��3� j��|L�`y��L1��L�w�\� �\�B<��C[��XG}s!ͮT&�*Rvsj�;T�̚N�v^�d?x�nb�� ~���7'�8*��, ����<'ܽ�[k��󍲙��^��
5*�x��R��s�V�B��s�{BZE�Q�311vޠ�[���C�֚��d�V����O����K��!L�zM�B~�vm�S������[vh��n|�)��w>G����p�gq��}ݦ�RH�Z����ꪚ�QN*|Y��e�X��A<E&��/��_�'�a��w�it�����y�{���1�k�6SJ��sf$�j������$�d%��U&���"��
}��_8���l�KN{b﷫ ��D��x��~��#��~��R1U�ƠI��9������G�|!Q��:_l�5���������x������p����J7�.�HZy�����N���}�9'̟`Q��u\h[�sEBǧ���,���!��}��b����c�(����1f��?�x�\��A�Ϊ�P��1')�zx ?�����H{|��]�(��-�]Kԩ�g�8g:t�	j�`g�Ϋ������c��n�������<X�մA7#@j��+����Wڀ'��O����Ԏ)+��*8:�1��g�D=��G���a��\��a}Im-%�F�B]��\�TեU��7����3,�	z�`���n���i"�]�� h\���|j��3��E@�g@ϽNAð7�%p��*�h�e���s�x'�ΚLz��c]��1�v���9R2�2ď�{�r�L�$;!F7!��3V��(�n�0A���<����Ssp��jOO�%�͖�ℜ5���6fhq����=�Ntu1�����88�;�_ z�6���i��J�{�͵r>�°�N�1ǌ��k�#���V^��R�#���x*e����CD�����Tt��N�}����z~�#�ν�=��8�	��M�{b/ϴ�͢d�~���_��%͂�� �-�z�dvGRF	:�Q����ᔟ�y��d����@~2U��+�����^(���sB�K��"1  �I�6�qG���7gF�p�Δ?�a�?�m�x�;N({��w���Ű�Ę
�nV�4T�TG��c������Y�3 �j���
j�ǂ�������GW�v��ey���1@5l����6L��
��+���@���͹i	�[s�Yc9�fgbR��rs��~�4N64��7P�w�k�3j�������#�y����o�|A�W�p��O�J�Yy�AQ�t��q$R�lЎf*0���H˸�݋�&TfL�~J�$7А�9��DrgҖ���ti#pg��BS�|%���~aYg7��Law+����O��G� -�9W�C��/Cs�c�'���Y���t��8��Lq|�}C���S8ӱsصIL�v[X%�	�,PRІc?u��Z��G�,a��7���jk�}#e=!���yB���ҁ-���<`���,(��eX���Je��J7U3��[��YJ��f"M��iaԆZI�:��[��%5�5�����o6���0�'�-y/lk�ڳ�÷���.�A����iC�r	4
�G�2� V ���[R�*k�̢Y��请_]>o,��P������a鑇w���X��c�Y8�p͒GNf��uB����/�H�R^��x8=6�rHP�Ydɑ�C��5B&�i�0�5���=E�)��S��AZ�_��]\g�tPܻ�]�ҹ�s��`��a.Ad�\??PiM��@+!�Z<�=�)ȳ�\�CRڞG���\���tv���[Y5	ё������X́M~L�E�$D	n�Q���WJQ|��	
O�$K���b1��39�Kv�zR�ΡX	\z'M"&��3̗紾Ѝ�!N\�ͮ����ۯpԭWf�2`�}M����($�#?^ �7n�@>N�xm_�e�&�����qQyݒ<��!v���J����HAƅ(���テ_��yD؎���89sKPX_��Y�c��,��`<��}$�x���U����8�Bd$0��TQ��ٹ�F+��m���g��O�=X��Q��발8�5w���󆸋��5 +��Ta)�!7�φ_V� �c{�X�}}8���F:��xLB��x�4��wӒ�hfv�O�M��B��at�$��L�y�0L�kZ�B`���H��2*-/�J�g����V獍�{��z}��|7�pE�]�!��"GLM�V�����Q����Gڿ��y��~ (z�Wm.���R���(V���~&��K��(f#�n��j|UAB�DL?W�N��9��џ6��	�
�U:#�:��dj@Ѫ�����ac�C,��u�2�iE�j�f.�h�w"�x=T0Fŕ_<M��3{o���k��i~�nyn�qF�G$���qߑg���p�u#D��;T�ZEܡ���O��+���D(�����*%��)�"vA�sN���[��KIR�ݗ�M�߯�B�զ&1:��0w���p�g����xRfx�q���Fg@.��`-���X�o	��'޽<8���H&��Q��?�,B�O��?��	��U�*0A�6�%A��3�'x������z�ٕxGy(?U������E�������L������t���T�E�9�l+X������Ȓ�@�/��w�`?����؛�V�ܷuT�Wy��˫d�Da~q�*E��+�U�d�6��?�P�p����L.�N����p�I�'�o�v1��_�"�Y���_1��{.�����=}� �h&�}Ȝ�OQ�����O�9`�ui}v�5t+H�}���x���B���~	� ��Of�l��y)��1KF�o� *���6d�ĎJ�h�F��G�hu�&\���i�����a���;� ;�6P�}�� ��>_�������;�����p�t��3C�<7���ʃ�ܤ�H�6MV��	��}�2^�!�@/��#4����W���8��QI����
�6���'�Lş��T��0��[naj	o�ဇ�~2嵨U(lƎ�bqGQ���k���1�	��<�j!�a�7��m�6�e^p��sU�fa�ϒ����;u3+қ��p�� �\��.�<ҭ~3Rf�.5±T$�+�~1v���ټ,�0��
����>����ոrv�g��id>N����)vJ��~z�w�뒷��߅�'P�(�i1.�2U��Va��e��G�"���Vn�����S����3x���cƞPRߐ�l(����e��!�KP5s�k�ڬnF��������ȕ�jX�C�80fz��f鿾q��nf&-��p��׻�yO�Aw�d�3	��$L��S/Z��nl��������O� 4pq$%��dIW�èS�*5���&�-�4T��� @��U���,z]�g��������{��+8]�+eQ�����z�UðM�K��svHe�w���`�Ō��Ǥl�$���C�Ǒg����@�v~W�*w�7�-�� @��J-b��h� 3�v�u �a+n܊�_�JU�5���/�I�H�S�Z�F�\`G�v�!Zm���*��?T��
5�����o2�3lo���\�B����|r�* 8�	Nv�Țglyk #��9�H���Y1��ձ�_�j'B��_��d|�WĢlFMfQ�32Ȯ�-r�Ib5�Q��ټ�C��'i�8���	"-�����O�zv"�;��1�Y�+��I�Z�ó=�3{
 j$��=�A��I�e�	��ѡ����L{�XIrO���"wC���#{���aL��C�M�l{�]�˂���mVB� �	����Y&����P���1�8����.Mn)�w�I7���������a�2�CΪ�Vb�6�w��EC�>s�t��f#d �}�ߛ�h\Q"2=� �M�[��$T�b_O2W��+�<�O�A���� �N���@P'7U�Zp5�g�/z)+׬38B�]�+������F����vV6$-��F�NI��NpWڀP�t�i��xp!��'�yytz�%�4���:M��'� ���G�kM�J �����R�������j�:�����#�ܡy8�a&���x�F?o�悑��L=�0e��/��rl��-@�S+y�!>��ʓ�f�?5Ɂ�9�����U�w��*I#��r1�H�O���=����;��-��O�C�$M�����P��8�D��� �I
.��z�Z��,�~"�2��M��N��>�a��E@K�poϋ8��������ё�V�Ŧ$d�C%[K�q�ia��f�II.v�i�$%�e�&\�{�2��ڊ:@:�S3�U�&��Q��]$��&��	�+J�ې]&���/�p@X*�MJa��Ӂ��9|m��Kol^�y|ݰq �_�G,^�vP��j���;8��5�+���s&Ή�V6���B�}�ɘ�<�|���t�{+�j8=�LcL���$?Tt2�����_c�̝�ߒr��P��e�%R�~^�l�e�j�Ba���V�|(�j���^)�|ZTNo���!�mn3�.��`�շWN-���a�*l�`�������H�4�#�pw哱k6���.���[��|�_}���[�m�;}�'�����4dt˴�O��3F>���؅��G��x��H[����C�CW��{Mcѕ�gb��3GhZ��F�DeÅj��E��:��d���b��\0�ʣJ�'�;���S�2����D�8^Y+�"�Ή��q�s�gh���L�jw�X��V5�GC7�,˘�|N˩�"���/(Ԛ����lF�=�zY���1.��:MF���T)��7	X�4���ڧ� 5=����a��s��7��!��Ԕ�@��t�/��s��`Y�^��s�����2�»�k$��!�>�p�p�1+����Bə�=��*�]P����f�� t��"��Ds�1Z�8���&Y�2��qɗ��J��9 ��1Dx�T�+u�� �?�y���H�[�Ǜ�������_���z�������䛛�b�e$z�?��t��j��$g��}�Wȉ�o�����.<��X��_��(�l�]Q��5��~����?g�<�$-�al�M�����M�M�$p�m&[ ���w�T?R��Rԅc�1ߢ��R�Q���b.���H~'8h�X�]�����i�r?az�{�
���S� ����
g8Ȩ�X��ǂ��\`�T�)��5#;��}H��u�X(��+L��e�ts�Mj��ơ�Zb�ގ�K�}W	[(�m����֘�,V�Y6OXA�<^?ʒ����|�T����x7��W%CXa1u�D�������>B�h������>=�t�fd�������9�+�x	��&��j��>��̺ޔg���S���;�5��a��(W��w@�x ��YE|S�4 �V�#|�u�0��_��;�z�,�¨0,䱘s��A��t����(Y���)�6�&��w�3�>n��ǝ.	�ƈJy�mU�i�'�	�s���u�@��q�=���}���ޚ\i�/��r{���N�~#؁�1��A��󒗪S�9"����0�h��ce�~4dǊ����Ԝ�h^�{T�0��~�E�������ƽ!x?�pd(����:�s�̮z����ȳ]ǹ��y��VST�<�Vo�?a��Y%_[(`��;�����o��5�����reo}c}�n��� �
Xʕ(D;���X��0��[x�¬�۩
qA�N8�I�=Ɍ1��`��G�Tcm�'+E^wo���=���bc-��G%O*�q��ZO��$����.�7���tZ���	���u!!��(��	��l���k�������g�"��d�'`b53#ا����8�D�=38Z	$d-S������������i�T����>��'o1�� M�}�E(����Ϣ��F��o�+��R/9�[o�̔h8���BK9�V��'=A�