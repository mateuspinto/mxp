`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51552)
`protect data_block
0USWSUGxovGsyBJteYpEoRnANFXLl2YaLKb1HPHqYwsXDM7as45UJAwwWR5WUKZWguzYAx4ZRLo/
JZAtykE4JsLJtwByte237Pga7/xz4eeYZhS8Y3bmdCemz86w06GRD15lMir+tSpMtrViZT6bWD99
Of2VvthM3Fp/HTlzmWeAK4wV5JQB+1sy5jUaDTadE7cgrTrCuX8M3H2wjkXx3vnMavgMw4azz+bt
yFidg1Tm3Rz1WrXwwKgKIpYo8/+SMDE5TcMjAhG5JZwGFw8wds4OWN7jRYb7SllgPLA+IhCidzp6
m8Ao1uD5EsbziwvwDmzdaXvkT/jFfH455QDd0QYgzhLGjISiwvvgz9qMRfY6NeAnH9qJILqdD1n+
wl/NcZYvZE183D7E9bneeF6z6T1Zcfi0OsVGZSHeE2iDWpccxXXqt6r5N/b7PddrCD60Ds/UlIE3
RS5unfpAk7mdquE8pjkj3AU+r5CIiRk9MqPcy58+MZKWxinkrrcokzhtrYP3D3sXR5dl4kR1l7IH
w7udy80fDw+dlu0TvCtaPSZVemRcaSZ1HjnXfnpsnnteVlSO1VhpBghLfe22uwkrV33KqD88o7Xt
ZtSEj306JeeXB1UJ8HZewP7L1++YXLeqAkEsSduEzaegokEbUtUSXWHtIefIHDiaMId/ldkTnGev
SANJh5xIv0YfpP2xa9WzQomXO1oFwLI1fxwS15kQbgILq395vYUOM8SwyyOl4oWhMs/iyBzG1W2+
KRNFpndrTr9dkO3IAdD9DQtoDaqbNqvI5V10YU7wMRS6hSp9PSBtOC+W4tFnr/a6NNotMmfDA7eA
W5qPCKLylnCO9S/mcfzt1Ib0pffBYfGDO362NiOeOWRNXynFMqPDKv+4qi4HVmazRd23sgDwCxpM
6YI2wZyadL3L+GSXrOhQIHLEER3i5D21DkGaMDbMzXfy9dZAtxmSaKMi6Of2WBELbbEIia2pIoaY
dgOJ8DvlYv/pYraBkFiSb0ZZfrPbfXxCwQLlNheL7DqioE8h+MHTQbQJYj2Rj3Z4aeATLhTVEXTc
zFsGkeqmFfwPyf7rI/Ptr3o0VqNCnv52wWehfEY4WNjaNP6sZnDZarS9tKd7LZW4Xt7Pl1W+L9U9
LcOWLShk7/onUQlYoahy2X6XMlZz9RpXauBeuU173zkPSGCgW2rI7TNqZ9h+FLYTuLkGDtnsL30a
lYZgYO6/2N11mZAXfRwZDa/aQyMlb6WyVSoU8H3M/FfyoVL7M8l2Wb0DfPVTXtrEiStN57zH+PAk
5GYEMjKnCxrsWIAfvU3W2RUAno2ODsgnQ/fJCtFAMBPU80XbUohmiUN+vYYTk8NYSmvmH989muDI
PGcb2WAR5FKuePHTfuVNUnhCIVVqeC9iwklfiOdbaM+1Y/7utV2AzHgqwhuM/70M8ZCDZVZImnaQ
M7ApD/uUdbeOdbMESR7zHPClwOjqLr16mRK5RwmyZxgTbQKqO24rqDZeTFr1yf95KxVb/swulnUy
ipNsHP3WcbGS/JpXIWD0JLPy2ltJgbfq6NiZ574AG2w765A5kT1C5FkfeN0va3Prl9kCpGae91eJ
pDWFxfPu0FJdzgorlYNHIJkFMDQXIQEasqhz0fXJDMcNF0khxjQ5Z5IbI7hzjITPks0mDYSpKPoH
Nr/oUcvj0px3NmIpDkDvhO8hS4X6pwo1vuhEvuth1XuM+9J3abuF8fIE3QlH+3yYIZrUXdinfDq0
CMd4sr8N94XikSb9P8uIx8PrFWfK+TonqD1zHTa9sl0bLw0Vd5VOpHer1ueHfRxUxm5jJVvItcPs
VyIbZIhNCdmcnu+Hxmthk8YxDooCn9A6mi4XXLkEjiC5XEqqAXGrfHttQTzIxKHrsoDBHa7D8Gdg
S3pWBOXCnGlEqe2QG7KMPOpYE63BDfePFasLAmw5A7HQJH2dFsMlhRz5P752ikXxN/omJVvMYmjl
I4xq6SafVdj6kBWqI5q/KKZevAOAPUcF6pHkxsu27Mr8QUFl0bQH7s1YLqeBAxuEPrjmZfinvHnN
uQpl1h3UCfwnBcTNnChNb8t/LYJmkkLSjtAxzi7+GiyeSaIkvWU+5Ug+u+2nd6iAmfpASFSP2HzM
dqVn0JfziCRkutuY1MND3ClYAa47ZRQUmZx+q6qSYVuYo75/HAqjljRUT9wzZeFSyIWfaYFLMxTq
qHz9ENO+QZdaiE0XgJW9H5olizWcaDyx3iaOBF908IMvYdnmT5out6BLFk42SVmg7hQBk5XL0uhj
YxF2SpDjr/PgWU/reXAoz/JxpTALzRjWnzEbb9yec6wegjJdtof5F4hTAkNaoj2uPe6h360xLo5o
J8JYGPBHirP0ZwKbtWLRmj+YlyFDrlSCY/2CnYlbd4IHVra0Cn5Kqh3BLmYGioSWGj01qz30YYu4
JrbX5aYTQIV+ZdqhltlBYuMAUY7RfDIRlA9BlpPyb2jdNEVnIbHjTUNDTVijopWzk5oN2p/VmAZ2
MVd+AmwLJBNwWrZ+tb7yRxI2/bRuh5Ioivav1Z0T8MbC2YKYaasGRV7fnZ8ev/HF14S3eX4W5y9s
lPmDv5KiSLUBaB6huXqjIJYY8xi6aK8OGySgafg2rbpvq19Y2kU3KVblFAYNKdxS/TNBwyKfrKp3
2phjznyrkb/+Csomyfd86OKoHxrZFPyasSwUPw9yYDvYBUA9BOgUGvN3ex/1tgkKZe7x2FzGHZVH
9Rvbii8ISUeuazxHj+Ddo3MdWZW5qxK7YZ8/fRG9nrcX3QCsDymqGy4LjjKySlvAAXy3IqEdM5iV
kEBUPvRLLQ4q37TNHi4ETCu8gCF9eA4jc7ofYwsnN5VQXM2pZhGXusqK+uZwz+82/T96sBBHI0zR
OtlB1v7JX21Kbqn5z2UShBnBW37z/qu0HCkyjIKZAgCfH+F74nrx9t7XoWP4ZFBDxiIZSHxkfLC8
C22mnmeSZ+Yomdq9+2oTRZSDnc/v/bOMgS2LeQSmjOHJvUB9hRQkieFkY3FajP67fc/doL+eOrxQ
7O/ViuXj6hRtbR7jDX6cdzYFpYGrewU3htkFer5bIZwsGHS9TwyinQaTVcwtGdO+xyjPv53JIzlv
AUCW6htU7XVoZC329vWysmrJesv/SaVzjRSsWY8Q/I7sKW8/gsaJRAKmEW3o3HeINZuMFZ9xFG44
N0rsKwJCi+ODldEo6mXXiQhQul5a3WI0ADFjt/Cd5/KFFhFGb6P4bJyycLNVIHX38HXj3GyY++et
MmEXJIUx9nmChdHSBVxBRSzotIXSEwpj/hz/KwRZNT/8i4CtififddOj1sHAqxU1yYjhLeOlp+dG
5lzBWrRdlE2+88MpgpijLi3DcHQzn2w03FLGgvQymBn/SiRbWypjC7jDZzii5NvOxrv1LTnzpGBh
ooA+2DyhtH2PBcS9ArjSU0TQd1SSlitFoQeqw7lLgeFTTzi47QkMJ2oKdnf9VuWmSw3+Joxf7/kr
BRf92LMCSFkqKhJoWqihUXzI808dUK3727ZetacQj0PSinRYj2xfGpUQB++I1F7mKYRfAZOM3LR1
lG003i0vmdfBVtUni5wEOMvp1a0kk6+C3jOCFfCfpu6UphK9DxUwA4gUyR17gVLIiyrkxo1EtdTy
Glju4fURaxD4oAu6AmLNDiji/KHACs/Dqpm2p4VAsMVulOVH3RbYyO1yK3u9OBPofIlIGJMhnI92
Ixo6xR0zQAVo65YRPQuLYpbYEl4gddcBdPxsN3MZvm8eF7Aq+15xk/K8jRkaK6Xg072Z5v0B3PFr
F9zq5n8B/dan9TaXCMsTCvu6XLu6XsAxnTUuCSKo4nxzLJPMOY8rqzb9bIK6DyX0IwY4cU2gh6ur
9NokljE5JwR6WIGgfdIklTaiwxDET1RHHjMxZ41PUsOHnswXCuyfblf+ZyMGIzsPwDwpB7wtTmh0
I7vccQNmp8HWnmePX5JuAqBmW2CGoInvVrxVRefYGwnjfaBoCDRLXyCuCKQ77YqYJMF7Zr+W5Q22
BTifK4oFtP0QqsRPVsPVGkUjSBIkNW1GymMqBbY0WWKOK0RMicaB74lvkqpXgDvDp5rGLosyK1t2
khnajY/Zp/rufD8G8fzt2B4GfLoywHAhvK4Iv+pv4d+i6stu8EUrE/EFy0Q+pUIZAr8hTIAeLJW+
McatlNi0HHQaZqnbPryY1MbR2LqBqHU7OpBtlsaGVaYPBk7smArELlxP612PINxyYQ2wabFlJj1k
HQZOAlIaAQ+6jb50qIvQtYLK+Vvj1HB8Ru8oCq/55eyoAyrKrJpfEC7g+328el1cGsVknDo3xtOn
AyZ2cmCgJ7/I4SXsU7V4Lagp0p0QOHlRbjVEm+LrtMCT/xrL1iK321DwoUpKacawkCdiyEyFBbNh
dEnV1g6YvIzZ+glNzJb16OdcRJAVSTuEpS4xltCufyG4NPk8Q0U5lTQvPsF2M8i/xDltKWRnMUvY
wqn+NQHyRfX2pW4lOhZf5KCHqDtJ9tInAddhqtJXvR2Jss6sdQbHyHXVVhUa9C5vPhUWHPwmMl1I
U8DlVZNkFxf2z/VClOibDfczCSa5m0tGcjeJ4B37o6t6PiFwHcwjPGUqnRFogkXvG2BUYVHufyf9
ugRunF5nuTnvNhYsDErKwmHNKD2yKQS9WbDuHoUQXFfKgIM/WOiKzOE5eVMJsLVI49SGj1vFQY9v
BAZtg6XqtVhvDGHrA48Eb+E5HglTto2m7cLueUzePQLBKnF+uISVaAzFcaEsAqJO5xXYNPi1mkEW
ps4cV+FcsFElT77sbK8JAGlhTdIAHAYlKNBA/idOYAGoqxkPqO1iMvqV2/LXfVoVGW1xKDmK28B0
J+xGraOHDes4QtQikLBtEfk+lyzhuZT+anvYR3Eyh/wjgWji0wCXWipW1g1vQOaQmJtnonTjK1pr
QzPJBwwGqLR3R17xo3Nijp6BbVD5ZFBFuBt/J0af9SVQ/0+C8HsuLkPwKdDFs/wocUJecq43lCSk
2+Fp9wH2b3e9JqdK4VVkpaYrfTXI5kQbqEd+If4Y7IiwKZwvuwiA0byCLVNx/NslW8aZSYH2/8UI
6X3jtrbDxu3Vh6ws7Ae/QwEP2nmFtEWML8+QxqF86CLEyn7EC5LO9EeffYL+LEtmtBuzfnH6pG6T
bd8eOtdJwM71MyV+EHmU+pZeKn9VIYsCZAo0Zs+Y6wA3yVOEhWZ6Ih7VB/wUHkucMTHYJF0KK/EN
jI33W74zPnu99iQKPdqbkDlAtvMGfi71wV8xdz7Es5rmQ9pq0CouVVCNo5UheXljbsWK71nxDYv1
bI0x7a+gk3lhtHCDaraQEWxwbUNqMN2Z3RC9tUwGVlGgCDBPN36oUPbzqsQgKN65oB13CnLtSBe9
9vupXChJJAeC/i+0oNdDMT+8M/qc5+ZAc7fAQWvMvJ6rDtAjM7DhTEVYpjUKzEKyoa83bwWw9qLr
1lN+OzFHt3QMJkAk8oyzUk2E9VTq+PH4jn6xODbWWAG6TwYiS6ctNgCTlNapkXXK0TkUATsk3h6M
R9peT6nXHcTtrkYZAi6tlb3SMJoUHvQ/EXQBLG0PX90VYflVK2UlqeUsSegsAlSYJfV4m5c1YQHe
ehzPElMJ0g0cL0+qXh1zVmRc4fzE30AMj25S9F0jwDlsLtV2a8ZfftSYU/pY/3/PqnRZdrRSX/Zi
r0q/0V808TZADSFHem49ZnGy5pms2lgq6ibNGyvgy9FzI7Zyozj2WVpr6bP7nVr0byiWvHr4taue
fGTrZwEM3MGOzUor6QXYZWJTSEmicM00p4hgvZFJyBLWVzrOj2jBJA6N080hQ7gq5gaMO9eAjmSt
1Nv6YEdsMKq2kPvsJsVWHWbvKRq53kC/+YUdsCmFWJqnrFcPaM3b2zTXP9finLfwvUUAMAx4ivlZ
ij/eLE8GZqa/6QSzEQbRyYkwC34/nG2PZFFFepC1WFrEnvej9h1aqq0ggYhBbkf5+A6r2ufOq/B0
7/xp3BGUSEI+tYMeJpTza6B1Hk9DNqBuMpSmqDB1idvwmjWaDrcYNISkFUI0Cfuo95hSeZ5+WqBO
JlE70Y7DGAfjacwKnp9r3pva0ehgvtsMoMaysYon/QvAQ10jEhwKGr19/yhaJzGwudmGFVixSyY7
9r/e4nPwhDU0HEQNXFB5y1BUxr/MvtrCeTqleLUzOJt/ECJuCU2mxjy/koJKZsDiwyF+JJhuWib5
o70A1Q8qif1ejvr/v/m5kvUU2AbDZR8jB+Xm4sTDx/n4t3gXXOxtSqE7/zAbHNxwySC9GALQEDSZ
ue101Uxk4utK5f/UrIH3WFDSA9Gw7Qrwu1vgytYVaxSDLzb1T4rEMx0AVpSTOicqmmRLzNTCpnuf
uQRjEC6jHVVjroqDoyinXtQmXbnveCRT+V+x/rv6GzzXkFqK47YgSy2EyqKw2cQ37NBv/DcMZbmN
rf4IzSFX+beERZotecf3mYAxE1lk8LF8Ne6g/gaQ8gatug/esqNgU9aDyeEn1vixeoWA/H+U3Qbg
ikeCyN0dalvddBS8XRoRGQ4qafsLlIxAY8mABdp4mvUmnRZyBxSH9F06ST7tdNZOyn9Y/lBy0vCE
JOxKOJPvuYbgxwje3feXBdNxAGLVyaP4RXwtcs5LDy28/lslXPemnSPO4pw6MP4eIbrXx5veAiRt
txdMGtBM7fuMpmeOx/LAkwyolmoBfqXgWV9ZQZtVNtgVdCTkfUpTzkzuA5YFjvzxA33ebWSmYwen
MNK31bAlVbOoDwVHM7bVg6JPtZYvV7teBX/08h6c3DrqclK+jya4TvuhCWPqa9Hav7O+T/ZzvZ58
iOMm/5hbH7bhX95UKQjJJqodRrdlK2HwV8Lr2B9SlMCmE4YjwgZviEGflRv2kzhKCkwu8LALcb+f
k3H5StYNCulYRqIl2UqgrzECAaWSvfJOpzZTNCzXJPN8iwTaCelrEfoHyOwbAGP6Fr22dMy0ekbG
uAGw+RaZkoqhOtuJ5W0EBR0nZ1T2o4VTyJzq/SAwFmSgkfdp37Uha8lQagcM9Ulja+hT15G0AU2g
DojxJKZeznbAjCo6NQXg9SCSuD8Y2uTaYhxZmHGgoTL/AFP3KEWZqKv/wZYtSfY6Xc+PxIJ+uoyv
plAyDyFGUDZh7H6X+0PREUSujtsLRL726zn9O8MO+ytcCidolVr/jKRAPoNijvr5JB6kLuF8vcTa
fYmDHclZ3RTFS7iCRYBiverVFFCfQ1sAbMLNX4r6YcXjGIk4fJqxYRpxxZ01wrT0CFoxaJNkkfA6
/BcGjChRvo4v29KaubGWy8dg8LyL5G3XkOhZvD+PJyjfFUWYEYmUIu8GCXshT6jfN0ZjmgmdNML3
Bo294B6kxHulWOvQ/h51LyZAVhn6JFFOzoRKcbJ2xSmFkAv7Ckb2mlGIA40xIYicHeWoXnYS8IZC
0EVrbqa/nTiKZa7/wkFPLLiESqWKPV7bJdEMSrRaU6VUU5ssh3f9RStNEO1lWOFfaxRKeONPyl9E
bgSIPFfriOa/ot6iEQ0fpSEHvINC1yKcyI7+6UPTtDMJqsXrBReQtdvxM78aKvt6pwnv+/xlRF+7
+faFX3LJKlieM7Zo2tXA3U1CACpSQDBYQFRmNvJBlUNEuUCKbMf40FRrt4q5/cP7cj6M/SeXOLbj
Zj2giXYfgSyNOh/XYpCRoIty+p2dMqqxGaGmADRh19pbLNaRBWsdrXoMZOpRuIjbW83uwj4j5hr/
2smMFeEbwbf/hZKTHkInDYmKcxSDCoQMeg6yi63+WHKsmDiPw6+/qOT5quQFRtBHL0E+k+KNCzwC
JoLcX/7Pf7GRFSA6rSsmoRa5B0A+QSuR+9FzThS/WuK4BR423EY1yGHRP3uV2dfdbGcEXqJLBLHD
zzdFRukrcq+Z0SEUhnFB8S3ziRpOsPVG6y9IUcUGUuWknKG5OqBK2kc8XP/x85GCd00z8HZn/pM5
wEUsOV8egzVuQuVTqJlrMn4ROA7tAu9HD2blsC1MAk5wPOyOMkZp0vSoqeTmSNY81B1l/I1NMEYA
s2iihvD1SGYz+BBO4baXDlX4T8qTC2wuz4pnTIFUD04Q599kECZznNnlkVw0W2h3GRauH/pC3g+Y
UmBxpjgjfw75UMydgbxiZdPTx2k5ZgFIQu7DlTItvXsWZ6xhAQAAfcpryYVK6ClJ/7ObqPi8XC6d
Ov01tf6Y1VPoV8ustygHHPSpUnNQsX++W5mICcKYz1ct4V5ZDnxlthGTOcUf9CW/s1ypzT9MKVBx
lAK43va6hbzePMmKnx/9sEsU0zfNyY0NiPJG5XHCviuqs+Gr8AU/+phUeJljxiYvxISJRtLVcDXa
QF7DnE73TDZDs9CAZlNvFJVoANbOLzl0iYM5TAOpj/nwrwHtNRgA3fv7eumqvymH2zi7d1e4DuYk
pFUCRKidnOslYH7IwZOXJbmYfXaaDkYE5+XphHh2BxB5/qHvTQFTT1lbgc582jnd0pkQILmpkH+3
DCJZ6eq9UdCEy9vPX6IT7VmD/FnCtwa5WgSZxWsvjILv7NXSOA+czZivIAJpbj+GhnpPbSH1UAYF
+Zv78gqWrGOtrZnYrwxt8j7WBmy8b1O6E8VJgXFM1IJniThGsO6cXTDj6i8AJlp8shEHTLiodsOx
+SNq/DQVqaQcLW/ta5fcc5eXnxztOb6VgIbcGCliEVl3wPOXV6Wge6o9LCGY1OkYoHy87gqpN3tC
ct8WyPKclXffL2PixiT8lPlb1SWnj9gen0zt5+IFyR69DFsYyfcW0oiXw/rAEjqfPpt2ryTZrqOy
9Rr2PAF9pPofSmRhgTW2jLPQPRJxKY73mnuf/UZvedikHB0/wQapOKzhwgrPQi8UhdkcpaPA+pap
AGjA9KdXTRDmwrCVsmEYJg4c09z+ev0q8vwi7JHEqY/dWfSJsobMSEHt7vkUm0O9jMTGZZXErdMy
z+hYwdQcE6fk/+eBVV4SO9a76WgOHRBXKbOvnMv6Nu6d6h0gtA19dh81X6sYUy1pldmk4ndBXPyd
l+KM98aretx/QqQVtkmVvBZS2UD04FZCeIzV8COqcYh2KZEgcqqmM7IWW3FQSvgIRYX+Odtn/RGU
HPkQNE+wrBlmX49L+bAG6ubOGZ608nnhr44fygLhfLbFr3nXdcNA1YO7YGMW5FzZrbISRiHtr1ri
d0IcyH2NVPPjzZ/yUnq6Q8knUs4woaUvtN+AxZHFOGcKMEJbbOuZ2Fl2YfJmmyC0epnpeFvpQmGQ
fPvsbNrqJlgB2x60pNgEyoKNsuxKhS9dCyMSeZntdzMf/MWRu7BYmAzxhRV3qzZjOcp8Zui5it5G
MVgeBjdEkbykpp0u2/QYqmZxel8QPFzK+8JvOPjvBShgdsu7aaTY/CGtR5IZIjrSRWvVWBIU3lW4
kJ2cw7RKJrsz/4NjVwJqYjQlx5mywzFJsPiwCy2tvRWj2xpS2SBrgZGWzFTE+bmR1UIcfH8HKzUs
MX92m57jdcpmgZtR60bVzBqcFdLCYatKrL8JIv50Lto6St68/FOyPHz5lXSMhtKTqJehPpwS8NXm
TA4K4rT4NQ9jvqM57xZyiJSSkITRKlxLfy+72r4Wuw7IQYkbdNc5U+ZrrhLTA/RHsHfe0ElPd7pH
4s3iL9Ji89HkW5awi0881IM7EvtpGDIy16ZZnggx2lWJ8V2iIejDubHqJv7I9HZkgXy7zPDqCx13
lxwG5gTmiqKeb+52vUBhGOyVlHyFOo9iirjqGoz5NDFO0ag7WEgH2HUiNupeDHPYdVpdxCAUhncm
cLHVbm9gASYuculG1ga2p8JxbL7AzwFwN8jVx98zBIpbFaABzvDkb2iPEPop+KYHX46jlAIW4rPG
17bu/NQK8iVpwDJse9bkWONfsMhZ2D1xcjN4xTvbwtBCOsZ+dJAmntJUp2WV3H2MiGCEhwyp6J/3
sJsVWU07/3y7WMgQNYan19pSmO0A9iU7WMGXGRB54AfmVf9r/AyMxKfxxVp9oaIoDAyymyxsjHYi
S2Dpc2wNlT1E/EnDrztbtDZDfn5E1InQPYh4WHLlAoxB3hn0rEyhSSILfoVTu4EL2YpiLnqLMP8t
gcw3bMZi2kat4t2FLRQ1QpoJ/syt3I5DgXVWVJ4sCUqowVy2qmlq692jBO/uY0VmL6eaAD1efjiI
n/bd/vBrg4w+cYf1bwT2bA/S3Nf57Jq0veEniHQT+Ez1HVUIJoPqAawAgI7nrXYof4LSaC/8Sh76
6dSX4issUUXF+V1I7HM31yJ6abAZqPOrJdmIJ6BMtOS4QyNy7wcbyaa+ZoTlljnw5ngjGUfjgki6
GpNItGORDea6IIfBXQ/nZKHT9t3SM6EwxeiDeHv5+mjKpw4CzZNFRfJeqCRlv5w/GDF50GI6Vmqa
uimzqgjZhStKBDmQp/0Agp60T8kRgBwWDqR+HGOTcL8+l/MBYG6cuf08grMsWmRMhjjbY3X6zdxZ
hQEM1aKF5pz+GdTfra4ZSQfbQboSbcdQLKiPoj1wTQ4IocmKwYrhHuvBeWKbXgekjmntfGpTpmaq
viKpixUHWil1OaYE0+9EV3jUMAQLHlBso+K2rSClvHJ+vN7bo+IonR/6SyAiJtXAAHFVVSleCFPj
3BHziMMpt6rk0W6tQKCGNFoszIHuzoxmJ40RDnc7R35lxu9vHMVZbFMErVKzzlnHE1egKFPjtDvf
ppIXzXH8M9SKpjz+ebGEXUVNB7oqSiuEqv4mbY93uQXRE6reOTpbX8LQZRLbKGAsz7bnMj9aJXS8
dlvMSEKTHUq6Y2uX4kkd6Jkr0+OxIcsTwkOaIR5eWQggUpDpq0St0zYKa0eGa6fHVwQ/lDThj1H9
Rnk62mqvwV9SpXrpoTrnkBXF4XcNAUXYLfeQHfEixfHPaiMtMGxmVu8pkWZw0YrejQBBr0GZpNRZ
OxKZXkQM3+9dhUVpfnQ1AkN5pM1pbHHvEHD09xspFdWWW92ghyvs6vlyzfW943M2JOg76lzRO1kU
1K32OEQXYGrI2Ji6ThXNMGuvzIuINpWcP/d9rtW8V9WZ5ISaY8RGY8qkVGvbX97mRZ0s2Owy3UKM
00rCy6aBwA1vYyCZ8XLT1bcfDR3COs2fNSkZWegkhvgW2rpmJiKu6+AtwB08GZirC3pCMsrb01sp
cYX//90oMOZ3AIfsrBH87zlN0yJeQQQUW8gHjWAWdtVNaqOXtuOq1bX2ril3blqIM6OHoDykkGZR
VM0UQWFaTCIAx59NHnwdwrhQujrKSZMEJv7WVC1YzZDcaAT8Rqu8NS2b1oaM/gMZyW0Yrv7ZLxME
mV/g+CJ1n+8vIzGYDAxIk5VHEMjqXy1VKc6Rr73Q9HykOQO5acljIsRHan6N45cUamdegr+MJa3k
LN5i/T8IaFOEeGjnu10x1KNhpWZt1t+T1H/bfQBx2IcDG2ADDCm8Kwk8CpcSszleLYlk7Vt0QuKw
xMSyLMoR86n2E+Bks1KjKvodMQDtrWDqm0abv7tslzy76UW8ij5CelR5L6WKeoducssA5BM/IDLP
wcxlfFd4WcSgTq3w+mnDTIs+XhkXA/S89fzPQBIy+2azmW4rk3JaE5XbC6k7lnJ6fATb0HSEwrGt
3HHhB1SF8gXcNtDEcNhenblK9VmEnRWQubkBw2uKDCUTWCfOPy5rVNFg9TojqizduJAahnGQxiMC
NNUh0yPfjbUhzLF8ltB9+ZZSM1mitCU7pY426E86kvV9AB1q2TqdzByDqpUfrpOTmi5U+3LVkUCM
cZqHAP5nHliyr7ABr3j2WVvj2z9nfOO/5ktKXzuWFyyhn9fWXtTioCh33abm2wpAqPzHpmFvUdOV
t1v4Wk0INNUcSY78W7P3Ck/baZGsr7MtBxv/HltBP3xY11PDyRLeRHnKENzdBSZkP0SqY9WI2fMg
UBKE+AyPsy98ZU4UhjGSQPtpFyzxm4Zba9xJHfGGWTlYFwUZCqhVjT/oZhpqBPEgBcAI22hN6sPX
hR3VE8AN86m3QK/HyocscgFQSPgbWHXf9fqks++dZZOCkOwliUirUc+JlCQniTRYPNHHOF2dhd3V
tNzmQfyds54KULBG1vOSfBJM2qFL8O3ePPM2ynD8d4dBrMbIl2QzQB3G3Ms9TjDgLyP+48pYgqH5
STLVkFlOil2SaZJCr/RgCsqPv8HY3YfyM43w8hphN8Gl0f+lViHpT9HkBLOpEKcormkMihq2eLpZ
BWtb+Yc5CYeD9cOz+dL8RIR5mGBSXvl9orZ1NdKmhrMBQitPy3ydMjoeu91vCZ4eTrGZ3Xta/Ksd
7ktr2YF+mlP9pk7dAyU21z5YJt1pkW9hubCR3gxkeWKW+K4+IuOYPD/SzTUIGPrJND+nY3WOMHQn
7FVQqyXfOJbTgmYUkCBIABoT+bYv/lYDpaJ0a4FoPvCsywDzUpmGSSq8SE/MIUSQZxQteNZLN5T4
Mk1/Di6fuks1RjktZfJa2r7Sq/tqP70mrhAV8KgRZlVv19m2AuY/mABNFkdRdD6rHWiWeNTqRPaZ
sIWwhU7mL/i+D+U74R47+Tp6DYuw3kAAauuS0LTKXcg6dhuN6ODJseB+Fad01nfM5t05kAtpVigp
k/2wqlcM5oyN8Dah/Fs1VIhkWRkyHFc30dpdExtxmzymnybX/MhwXC0LujlPYUU2DdzFw+QZoInQ
4XmJ+pfcLYvsWZTzvHvfW9rWu2+Xd04sCfMGl0ZvUs2xuxrEJgzAjpW/Un3yl/RqtvhRW/OAEX3g
ljYhTh9Ty9385WTfnrLJBAqrHayOPg24V19qkh9hL2DeOjogyMUCDFHOgd0VmKhCzetHSOAaU802
riQbYur7u1eeZEsZiYqfLZAfV9W7PUaO8Y9RwHtCAQvlDDL2VlV1FGjbn9+v3f3E/k8eilymL9Y+
XrqZGkeyIFDPX2e0Lmb5RxZTYkmR5rYSQs931P0lQ/bvmdylpgbVkh+Obvg02Q/Udx0EIMMD2TBA
LQv5OpTDbxY2NlnylDHS1EufdPh9XEk6mvlU8SfVQjpiKBEJGK3dIF0Se5VqIXScCz5PPdRsPWeb
tc+lJs+JkP7c9Nnpi2SBoIXBvItO2sW3+D6lLAwasm4sCAhoqohyaFcJSg+i4dZ+QfQWSwjiOI2H
SupwuEXpTO9IQyNRGy40SaiNS4nOEg+GMXORr8gnPtCZ6IcKEZd6IWpFYrvTANh5duWNlis1NIGc
mC79odm9twWj+CrlR7FAr7ATgR8jCrVTOoCIzpf9f1JlWuuBzJLMaQ9CbZL1WSJEAh10vigO2J+6
d1Rj2Kov7Q69A5JJB880uUlxYnOnWnsYtv7fP2MpmmDOGWVz8E2fTXLO0VOW1PCtXjb1kTLEF4S7
4x/boJsiGcovwKnBqa9ytr17igkqmAzIOsAfzRgS9w9fPyEgFKfgUtxNxD9sf71kHYmC8ETpodxM
P/XoywDU0+1NSRfpt0K1qPTHStLny1/0SCHrBQg+RtfSRHVmd11w/EJU1CujIlv8aaKZzvaDdWmD
sndvidgtrUjzqARbVa2+4pCVb2Ob4bI3LF3dPp5xSriEuKsR0YwAin4YTvR8dogenGW15hISLCZK
70bWA4IxnSBzJA4B8c1KOzn7Qf3IP2rVkaMogTDeKQ+bKB3WZH2WpkIG5+lo0xngWPwwiCmJtqlt
FXKpKyidGCduaEoMR7X/3/IZNXHCjxzUnqWVvMd5rG4PtiMvSBWfJSn0dAL/9R6F1NniyncZGsoo
MAabjIqnhP91Nkl6o5axnecJhhA3SrtqX8Ob6D69olKE1ND4QaaB/aWqWxwJOd/MmnS5pQPk/Ws+
cIgwu8dqY3VWoWcbf2EhHBD8aEsUwIoGSWlD0usykP9narSvErGo7wxrPrb/WIzjM+lzGJF1Suah
tAKbSf4aIXwoT1K72ru1SWvbMFOxPl+/7aPf4DJ65qJ16vNJXPWXn3CD0PibzabnOV94uZmemn9+
6qopLzvFMGvNUT8ubU1/G7yxVbkH3NjzuNBH8PE0aart8qg9USGClggfD9UIfRZ62gseLImiRSlm
GI+b3lD3dzZEx5/KhgmUnWCAd4sAdveHQe0T67G8pqnDFi5cOszKMMjoT9K4GR8+GWvXgqZs1XPE
hI+WhyGHepO535gExuMa0SbZTp0WFUiulg9FWPsxiG2x7R1kt413a6aFfQRRlETgEXR92seGmEPz
+OFOPeWScAQp832A6Zw6QGTxKHpWJZtu1EmBCRvUIDnTa6KYmUIJYzzdTTiVVfh/4GFmbI+H8Efs
wEBQ5O5C/m2nlnOkAZENyYkiwCM5RPKab5enfKVQjWEUlls3ILd60HsrKTiCCexANLQJgORINUv3
TlwVA21HHG8Z9/vIawllWEFcNghI6K44/SlVqYoc2+rAwfMvXfwKI9SIbzeoRk2/cYiA9RCnMYAh
PLvQlSUXTS40O37p+RhXeBxjT8RGATuJxgpqTisujk1UMq3dxJbMTQeqXsxTXdWAWQ6YiJb7FF6L
fcwmVQvuF3bqTMP0R2f2EeyuaQZSX801M80KW7yzidwt3TP+dnVcNHmvMvuZ53B/pp7xNq2XLeq9
ofDQwp15NU3tfUSwz3eVVSKrXisKJHaD9J8LUCJgqFbNUWKbOF6dfDKbJxqEVX/vFQuqtFRGppZu
KAoAO9fOtpUPct7peLwb2qYHsSjstMEo+ofq/lAcybRJv+y01R8BpKo/RqvwdO26xFRUiW3ro4bN
OYrmXpbmplRPDa20gx9AVbw4TDL2aDpOMxyivMo3nMghqy5BeaMf3rjCONHYD44R3sP+pk2PyY55
w8JwV5k4Fz4WtncYMhg7AHNwS8JTzLBYwht5E2lvLodB6spJdu1VBIEEUur6Qt4ZJXC+J1YEzZ1f
E/oC5ZWFg1fFxsMKK0iNt15Ct8NAu4hhINCrKirnbG6FrLAXnbw2D88mr9SbANDU+/IgTOjSDIty
7ErSTi6xifkrPvNbtt1K/gQhwBykqu26c3mDL0rC8H10MY0NUjX85SNlPDa2ZQy9iIEh05w442wc
h2FPbKGMy/dclC3QUL0+OTfZuv6yBtr7kd0/THQCVKxJgg56rqWRgMAFWhiv7q2d1w3M8IMOjfXe
w1UWb6sodQN3O1OShrlZH7VSYP6Bl0fCtJd4XUnOr43Tagq4DIwMmm+GgbjlOAO9p+fr1Pn59pah
FAhLNLgTaN0MR6+MVFl5Kzc6XnF4F49T9vJ/Tx5SQWiXwY0EfaxG0End9pxcdwFI5QtOJ7TeCs1U
qA9/gtuLpjXAz0BsMZMqAOpxJyAw/JZvhR5qdr3lvkDC2is4GLYDmUhZrpVyVG1PKpzSngrxItUf
wy07kxkmiuuTujUXNaXwG/WWgJmx3SHyHMt9bQMXDdbEERzLWs1KvW80lTcAAaGDqijWdt8DQ+UT
cgpsxGrlnGlhV/O3Eb3a+EQnT9lotMxzOWWFsdPsmzowW8+w+QngmxJNiArazDaoYR0Nn/8zOWyy
3cAwPQ/0D1MOe8P4MfnNLCq19A9qzvwNgHON651C8rlOiPTZVhL2pnE7ftisXZ3PKDvlk0SGVBvn
MEife7pfJ/sTYbLifsd7QSMcvdmAdVRBC73406lcl2nRB/EmPB426RGG6tiAFo0zId0mX7OY7ejw
TEdH0kIKWBVGiXAu/ivhXvzZVq3WUJ/4hAprzgrcEWQykEWBi5fEWejWdwmBWLzgAF7svd+ki3NI
HxVJFwMnjVxWAIL3R5aGFVBZeCzKqG/nYeDCHBXxynMTuCSze3adwxz1YFW7me6QS/zWiPNx37xG
H63ce9MGgNNr4GMg5hBlYLZbkhYzRwPyDVVsJt1LcvIQ5c8Dvdrut2g6k5PeopeOOJ+x0UaartKC
/x2FiHHq5YH5UKaR08H4U8DTz7NXg1rG1gLLKB769KqhpnD+fSPr3NNFsHnYj+r/B0isRsZ5Qotj
Mw/wAT1Pxe4N8es410OFgTAKTkayaElP7vaBNaB/0ByHbTjXF92BTV6w+O8DH0PJFt8qaUhOM8zD
ke+gDbER1hIWiNuhXbBDcro3niJwkOhTpexjKRd0UJgmbQQ68F8xpWjdJHIWfwn0DoofJSg3Pkry
grDjYfmdUhUCpfE8eZRAYA34E5GgM3Sm/qwQzzIs86jR2c1I3kS4x1LLSTZU+YBNCFpJqMp7sYlh
QMzg/yPZuHhnquAXmtzA7PieJtoZ71inQkZwCB+wr41zmU37qUtiI/4ETbCOqWvCwxx1HKoVZDgP
6Zx+n+pdYQ/8LvDLlgLVlnnnM+m3BJVelm8J2KTkiXCeSkcgdcJBOVPII2WQgUcOQyiAPDoSAL6o
CEYQJS/Hjmf5ccaWVStFAsM1PBtxKUw3w6ivG7DtPZnSdbfUReKrMI54PjdD+8y56Dk+KPSOEEvf
7M45f924DmUfLR/EGXEubecRUVVwcRhjQOphniPZayAdl0D98s0eTNiOL+w7l7AxFWRnk5Ea3dLq
2klaEQ0ryDeMR3di1vK41RIfso4LX4kr6ZvS20Ajhqc3DqKf3LrkgsTBIoKn1pHoqZ29wZWn4gdr
SDfqK2dMlK0eyVDzrp9d+TbEWFf6su7zyKYyD8EejBDzZ8kNb4IT1iuo7ZNGOEq4e0+zHjVaUQSq
sx0/T3YWyMXm+0UmQiX6wgoO52If0kYaU7YRuAE1yWKOog1P/nGtZXAivx9zay8hmTwnw+89/XxC
c86wFQJcYh8cDZCr6A11B0wt4CM8SL8sVvHOi+pwkfCePEunXXlK2/IQS0z3Lj6q8p48Wlg1exEb
kbme0r9UY/Uuzm/nHkWv/g2Xy9qa5vMU9XpbDsaLiruBCYeHshr35v82MiqLgm/7YLUSXfF6zOOO
+SvjOWKLanHJgab/JdkNlPH6ZsrRcz9TxLlMccCPviqsdyS04NGsxZoy2IkV7H+TEyUzn3Y4TOmM
oFoj/gokFTGBj69OhfT1MQ77uAtaJMo3fGENEC2pDvsHi68npLpS7QBNwvmvzTwSwO6VQ+RkbTPV
0yTDPfuaeBfL2HwxTKE5cqubnLtNQ17pCaKit8EXYBDeV0iv5CKINzZhFBcWmn0ndVfOk0lXCrV0
o3nOv4qDq/JJOleree0Yr9W3BwWinUE7KDyRm5jhW3gVKMMeAL2y0SZM9I+kfLw+l43P1v2iiZFY
6mLI6vMvSTendwR1K+Va6PKsNsoAZl5itP1bYagyvnN1plm/hYZ4mKHAAQj/Hi9+FkagE+DUfM6q
so6CDYSlWoQfUB3eintKW1ejlVp0A+8SKSc7hH0JRlVL9Kp0KB9D3UeQHPAPn5xvNh5T27koP0sr
XKrbhU8a4GodBikj6uYFwVPaoXdblqs0YITHiJ3XflA6nRK4WoqEDlc2kGZ1RpZz7dd913wkC/gG
7t7tmMhubWR2jtpy9+aw7haFBbte0ejXskioQL0QyMfuCoGty7M0KPNG1H9u1nABHNS5XXY8x3MD
0vX2UjkhDImpk1VxgiIQBqzPJgmkTBrPFpOXM8B2/yK1RTOfyMv1nfmpOfFI0OQiYIVSwxI2X/Z0
+kUg5rYyKs1MZY6ehb/hZ4MCUfwTBMl99SSr4F5Wd4gdqgJF3H7N6FFXM/hY3dtBJrQi4IFaVKmq
y7VudhNcssXKGhrhXBwTbDytQX7qlKyb9rKFkPq155fjW8DVAE4VNsbE1pFW3bQcFz/zeQBTPDE2
EOdgZpElZ7nlMcO37BSxn9tCqDEvCq3uZc7anntibt1rQXUiBE2a1EMvuTCNWjesQgut1PvXnjGU
dMQjuJxkgh3dDPQIXlJyLVnNk145ZGwNgf7YWfyIDkgnmkNyzh3D4VdyHNC6pCMTNzC/zJtyyR6g
5yZkpv5HhmPxrbeAIVSls8soatULvT0JOZWHzbkkAJudG53h8oM3wTXlTYmhvyj2hJ6i2wxtthqP
x94j3adTrrJJlHdt3AWfzY5Rc95dg2eeqkozRrnf7ADMwqmt8LhScJSAawa9SrSSgbsH7lYtlnq2
v8DEwp0y+UcSlTp12rssR/oyx3raHFnzZJON0wxeykfVCr4TRh/9vJKbNdCd0omXP07hU8qgzzZ9
k0/x5XuDc5LVZzyKXCECXEKX4bkObz1OuBO7YHbtD4TXyWlPrXi8QH823rjfkiJVlqHsfGmMPsMz
oDHJHXHzj4iRuTn/Z+l55WwyUwZ5cAKxhLJTfvzcIG52OWsn0u0H8/Ez9vWbrXcmnfQ8IFBDYpJk
zS4EqUCxwuNw0MI9Nv/g+8KCW5lVjMu0xgRoh1eOamvY5StHTh8GHIJkR/D/ftr7na8gxUZoK1K3
x0X2rWtCplZGtjE1wlhfu8+wGK0zSUUyDRtBrCzMY0Tv3M2w/GUcWcu7G+cPqeTSdCbwUrArziFk
pq7WtSdBl6nlsuqtLnVG7k04hjjPt8VE4SOiIeQI2kTmlN7Hvdkx4dkAj/21+FJ+6cWYrA0yYYP5
/4/u7p5NejkrZ/YJ5DIj97xNdQqt2ZXUSH2dke2LqUQY/e432YzD1CZewHBiyFsGH4XlH+42GFav
4edpZ3oBfc2Ga4uiYmUIAUqMnmx7ESs451xMcAMljmyTr5+WAN8jjckYCLPT5CcJLcGA2U4xjBFe
iWRREGbWQmzUr9xS4hkWSm7JG3mhMgoEhS2p+KEY982DBi8fqUMQqbNs1pQgqvCFEkxv/Vlin9dI
wHrKoRP9ou67fAkeME/ya53df5b3O7WHD9RxNUxAzjV73d1P79ua0CszWOWRhpOuPEKs637U++Xn
d+fg/OVeGBID1Y47iVc3PNPqccO8L+dTZI7MwRaytIEF/FC7BNQ1gDvb2nGtVnsOHX+Ok+aNaVKu
3MMX+yr0968DQWVTGge1xBu88B8qDmvyb/ytOrm2v1IFu7bh3rsP/LJCJn+qEDMD6tstPwkDXp+3
Kd/XsdRh1VhIQO8iDbyX72bpDnwtjoVhlP2HesOAN4Qy8d4J5YHIItgDtcmgBAYMZjAoK5Whd+Th
zDddKMOX74vf3q4Pyf6/HPnzl8z//LK4v1uzAS066qbOe0rK6anghvYFkB2WY3aiQty71vpy1VZS
rXQEMuaH9Xn5rz0fltjI+roYdYM3X61Oz8XHfRrQQoeBpkltaVk0TCeheELBsg8/9fvjVuUr/luy
XYEIKM8TXrT3hG3OrVtGuCjhf2BuzWDGk+zQgYxD5bPUzjeflXxoHKKthn4xICG4im9xYg5wYH2L
6AYC7Tzhv5Zh0v+7bTGj+ERyUDSKL/iyrgl5J9BfnEk+mXf6i64Ko3Xy/mF0ovY/UYsRbGK0nOEU
7OgUJcqtkmbllXZGrvva60Rgj5ZVrGyXKubU3/IVIZuppYfMgG6mhsZjo/vF2lk9ngBUsOaLIIsB
o4Rq4etaQD7NebiIkj/FDix5ebRc0jhXb1ZyuUx4Q3pHEOaWGb/AdoJbAOD51xevBWC2V8i3WV+H
q14xmVXGOYighpf8l8kE5tPQQkAij4A2YL/u2oPCOph7kPl3+uMpSO95iXoouRTdg1JaJM/YKt3n
BJ9iAatNoMdzGt9DMFrFzRkPpggV4xgiGQGBQp0mhbpbStmIn9Ywaodc/IFZ5klcBjRwghbFv52P
mvbRadbCYdWgnMP8gAkmDpsBcrz+mFuho49yCZYpHcPXWgKrjMWOp5bB8tNp2/VwHPmW7X6Y0jGy
as8tSdcAMG3opcTxuJ55UIxgcAjSKHllefMaJB8znMG2aSvYaOwJBDDgVFgGwowid8SnnJKXrWCR
pgvwX6DfTV7xbEYAXhPWHdiimjOUiB6YjuIhicU4QENPxwIBgKq3lMaEkmFz589u3pDOO9N05GZw
InSjhwcWav3wZXA1AjRTOBbzwjDARiSVcPF6QkxjGQJbf1uqHu2zfdPJMAmJYnpBSimZt2Q+9wUM
eHzNT5NrVeZZg5fv3xAAF/b6vItq6NEyGqM9UrMx5cNZR8Wk+9MaXrDgZ/vj3EQsaEWzwiLEkbOq
gMNrHNSwCeVscbnN3+vY9pCuUGJjfv44viZzOQ4gK/SVBH9Ox2En8GYmzBACKV6c08bai2FgAPf7
gewtIxQa752mEM8KFS6y6DwBY7Uk+s/6/1L4JTkj/ZUW5YtSBU/cHRG8jlwMuV1GLmU1yx3TcmoO
SQeT+/uHjDHk5Ij0jeg0WvQFyeNewqxNTRLyb9E7PlQJ1ytb66woMx3MXSc2cLKzsh1ES0Bfk7bL
GRwm9MwMpgkHZ1ZGBGl3yXf6DsD8GDal9FwglCH1T/Twmmd7r06TFmPyk/jd4UtBF13cQivsgdMA
ivyNn9AR4/rGqVBiGOtL2gHXzbyuoVtqga/SuX0oFDT7DJdC305FXkJA5x1r5B4iwAFNgQp1+5Ku
tSAZOEwDmEsA3n4A5OgyijZ7LbUaYQPXm6cMcARkXlSc+OCsyLGoMG8MWTZNOzrwX7S3TL71evb9
YZ6FbMsDTQ2v55QRJxI584dsJqFlq4L/pLkQzdfEw6tr2YamVm4duk+jUUkumjX75fqzoI8htQn/
39tn7lXG9SeeZbNwdgSfL3yXJiXL2KxliXbHb1dC1xHqpqdfY+Sbgc5DrkQqYPx3iB6j0oVbqGMY
C7KZLgCvFDsqpUwC1M2wEfS+rVdbuVNIlu8+r89R6NJgFKU0tZ9JPYxMPgI6k+QahM912yrWwDd/
f1hbwQ4jqeDWYLlk+8XZ5Yohd8teBTIsNkD9T2FmGmdTaXizCEdEIHjiaYaVQGgZ4xIlUK+XfQT6
PUDF9wXCBGJqCG9/rGAlDBGe+Ii659IYW39jqBAItrxrHOsArSjI9t6EywqLdefcvCyswmSAMWek
ktFdh5S7DR/VkZhhUTDtm9nRKeSKSMioh0rsD3XJg5C1zQhnuqC/QNqVNF3EEBa9PMN5XPiK495G
n+aHfLMi1F2xUGLv1s2S6NiFonWvj4jN9FGPR/+se+ReZwFHp818rmfZ5671jIMVcR0pax1/StVe
Wha6US3ytvOg7nzzrsrbqnxCHekl8PWvpt6Apeb67EF5culdajv4SHGk1Efg3cZlhx/3n7TNcPra
XCemhzhMQp16oGyfVn7C2cQs0Ajy5Y4giRMFXaxfnuMjEUSloEwQF77J6Zb/RZUYj8dJGPmydd1a
ntONHuax7K2pkHtgsYuK9Q+Epp5ooV4mhL01gTVLno5ZysDrL+Ml51BxiU3JH2g8MxDQue0jbrsZ
7zmbyG0ps+q8Z+J4UK1A1dYCeZVHmtn4He0mFIxGC25C5nKkeFyQvGpl9iK+Sq22Nea/c5G+6ONT
QhZyNbAkJs4JsFNex3jaCyLctpIp7k/kjV6TuXK5jJkpNvZLO0K52olf8tDxKqP7HL3MRCU9/oOA
TRTEA1QvdWdum2LQbM7ELE73sTO920XWymmAOIeGI1JI3gNJ3+Oi3JNEe3BEc/e0EAvGTAFvajg9
qWrwnrjSomr29GFrz0oSI1lwKz5iQCGhXg8K9FK3G/uUogagHJHHt5y3rrQoHTaLtbUeK6slX0nE
Rg05KQwgNK6/2Wh5rHmurZJyZKy1/1iMWB7cfeLgnF+8LZGqkA/yU6kEylryTHGir19TLDXn3anS
3GRf1unLLrtRcMwZMPDH3WBgdhSX5TgAE0MUuphk51vLE1orKNy6RoIawciSHIVQhgr3s9bNjOkV
BdVuh3NgbRGUFx5Ps/FmUKZ+NPhHw0+6R8o4DDEHIrjR0NK+xcHwV8ydQuNGlAI5Er+8/QZpZQP3
43E/4VHnmucc+L0XoXUIe2QjRV7sZct1a0gFh90JjQdJnkWWhizLXSxuNSDgFXHxqZiCtsGYSd97
EnOu/Dad6HWt00IUacO3tSJBPHM4Y/hE0LS75fs8cgrsggsoktoggFCyLSAkb690BW+V1iw5FF0u
HG6BlKB1ujIQ1NVSmlxKUmE7q5Yz55fCPU/G1pAugWxBTi/1kAOHJMDB/YlVDPN1JfKLdIiIvQ52
7neYZaGLjta/QcF0mZE9kkpvbhrEAB8HUYgBGRP3ZWhtURIaAWMBcftoRard3XPM6Hgw4sCrZzC1
OQ2VaEmjqMbziwCKtglHqY4T6wlMxgFiLeplWFL+sIFOyHnrmELVg4zTSnUqWZRugAn11+BhfOF2
fbKb40OHE8u4QYmBAEKW+e/6ltm9MA1cdjhUFctgdMtbdfCTGT37JIKHFO6RwyU+VylyT1DnHtBD
wzWwVylq+Zu5NglY77qbX32SyTCaR8blS/si956BscRE/RjYUG/fZyDmGEvVneXFsC+4b8qv3KEj
pb/z6J7opOuKN9UeTo+7nNStV0IxhkzQKsrwaI7O5GcRk+wJCGpmOn/rmR68V++IFfyKHL7GXGCi
AtfUSQcEK8PGq6xUZY4YsiqYGBoky+ivw7ZOZvy+hm4Avv5PAa/FX6yzO+jJum7HQGk1GDwZV19I
RE69g91GThTzoNLM+wN3jFvwn+bd29NPebU8DFb7mrAziHv/G+mPwVfd9HXZ1zjaff3EZDSJLSv0
eyS1BIWITUN/fZoZUXBFiJPFVdWEKOQsN3uAFugFgyFDkFrKIXWHgRD+iWM/LKzzimMZ5s/PJI6c
l5v5lgw1zRgCvfk639DldVuBT2gas1VDSikNNjWsQhpknjKawSrJq4jlVuOEV2Vw/r+2xciXu2Ss
bTAqdmR/GJZtmBhP4s8vr8CCGJs4nvRAq/c9P9ezzmnH6++UdJ/PTEk27MyHknIB9NoM2zPyRL3w
RNyzSoasuVw1RaMKkX0C+iEq9qEgQ+tjznItSsRDpAbgUPFA7+s8mkNQWRxie5rA/kJxDBJhxc5J
iswvJiGfRFe130mohJcAT50n8V9gSl+kh1b7hXGCzePc2ALY383SIX9JP2aFvhHE6G0VaQzaJWWh
oHc04VvZXDLcEKtnYKOGOm2jDPsOXUJQbg4h42Ebk0oHAi0WEcAIC7GlfojcfhTeEZvZaXPvj1kV
kAJTeQ8CHgbV33r5RRFVF/zbXKNKkoBQQf1QSN9vFH25j3+7K2n0VweeD2qIQH5qLo1akT0rLt6M
9wQbKXXGXdSWViY4cdWaYfTQMJrAIzBAdmiKDiPkfKUbv0dz9y0MJPqMwgKmemUu4doG+SmXsMwm
O3SKA9bu4X0SoqCY+yq5M/6ZEha4nmgJT4N3E4MP0TvxEcxTiIBtVTAC+1x7q9PEw39DxAkS4OIr
cWb9XT/dSAkZ/j/CmjCoWSc/zBLyraPy2esXP+nY0ST8WP2LqtSQHLrbCHtsbxmz6YaazebnvoUn
gSFINdv6AJjtrdsWw/5DuXPUdLleGQxPuBJN2vsSVUTFed2u8MpkHEMzp6lNJbpJ3f0XnYRA/TZ7
MvjlRlgxDBe+QBm/Q6JeDLt4PLpCAnC2jpxmAVkVz7fC6V0ITEGwW8K0zBGuRkrwfhW2Oe635lb5
sEUHj3S7P+knFEYDp7iWfv5U7dBEE18vBw7n9Yh0FqFkO4n0ILn68xaduWMHyON48ncIErTR3vDn
5f+2yW3nKt5VmgrBbCYVnflDF1IeUgzmMZ5+TRLtoZIeCVXKhAC4CT4ymlqyuEAfVX2u/2HR6VI0
8+h7S1L/mAJzBoUR1qr3Ki4xrEq9vfrqc/saJ0fpC6IRmtyGRvqn33fzgtzmWdXB9YTivzXjlNq8
klfuS7TDkAjMx6LAF1J3ByvO4r1zn1Lbfqeqd3GvBhj0NU2t82N5E0MBsA7LvR8lyBqwXG6yPe2Q
Z6wBGKP9nwFUsT5/FEfhD9OEk3lmZ6Adnq++r1+tbgYAv8bVuZExbjYql38YxaVpz2DRGv+RyFMK
BEFLVz2wxBGn54vtrIxqnaz5At8HCC/kwiQdrPgkcY3ttPfBONfu4goKiUM26U6VpJIpvMcpjXTC
exsvsqmr5PpMi1AnjcNwHWJew5vI7RquQ9H7EKDRYLiMUbXrBJyaeskgiPxOURfv7MxN1sL9nb12
ZWTqCEGIG+q9hvACuScAkW0s35QEDzeltWQTh3DVph3WsUpLo7RHgoq1ZDhcavbIup59MLxSo+EI
o+wVrkquD2JG3nGlxMhEtV5/HQ49rI8Z4I2HGXh6W3Gja/LYTsSZHsX4RdSHjHS28hnEXbXmkkl8
9DrtsfFxUi6PK/3tACG/qgem0fMS4m819F0uPGTD+PuRXBxEl39HUsZ8BpkZARTiQjF5X2VZwlIU
wDX3PFNGTGcJIKWdHp0N6UyMWd7sa4M2g2XhYaLKsmRM3I6RgCPKcVW2KVXiVZ96y4o7MrLuCb+S
bzWthxw85vpGS4bKPSAJOdPlzG6nseNaHakpqMcSKDglN3ymc0vpFPPjLSjMwMHZxgcprTM6DUG/
8E1Xx0D3DFPL/RZmGcnajBKMXRvn4Ud4gdAYGzGO+TRL/35yzS31l3vXJ9MvkclNHVhUafKqEJ7A
iWqyO/3LvD1qCOn27GWVzInO6GFGekCIZfcx74PwmwKtIPRftbJjIjqz1LfIXU455fQytohWd6RG
kW0zJAYEP3WaxsQEdHPK+4SEbqaLaYS7uuIe1A/sOTBd6mgEUmLdadqE4qvts8+vkUvcb5wBhab9
HxGWJvgWgPe5OLGAI+I5HTajhwcEyoiXsCpVZB/CpHrKMZYT/1l4XRiIRRcZ+nH/1nX21cqtOwPr
Ee4xOklC6wUz6j0nFVcgF6IbKBKckxE2Nyfg1J55+eRXyTQjaOYysXE+gz9NSwn73Ak1lz4hHWMc
8AhNB9JCJplRQ5XOrPubu6x2M9HZAPpXdeduJHnvifOMHGmISzZLUIu4/LRIHFedPO6y4mhlTgwH
KVzz2e3siSmrx84cmjpBFZlxtrDzqA8VkLY0ctrKYefDyK209/M1nxHqRZD1fsKkfZXjhkx3Jzed
TyDvoHGtLpDK32QFSJoYNWP/4T0lION/DynrLgo5727q6vMemHCHTeTWATsKwr7I47ONgYkPxkjO
/Em3pkC/+y1Aympg3GLBBrUstc7qj+AEwgqIUWddHbEdv3RTpQMP+OPWULt4cFDhp1EE0d+tCWaw
+M9g9v3RXEh6GdRb7ZDxbzlUk92AEQZjoPF4Sq1mg0CZHufTux2h/E/stXjkMEoiVNW2GKSNbdcQ
q6RUX+nCwVKMIOT5h1vZap0A4xxYdvyMp6LTrQY2Be1aGPLV4HtdaNiHPDyxMGUiBanckQn5CobT
nIJ4+hnVAVO1GyGbgGAZsxkv3Y/Ht/cepQDcykiSdN3FnyBGZUlodWkF/6zQ10UNdwsDNqd5lKPV
FE5+vBktSUq5js7Pnt+9EB3FEPo9T1o8ZyHPyLQrdHTwcitkgsSS6UZkPSx1XzgyWsBzJ/CmkhCd
EiGXShuzUYD5Xpv8cUKr/mQMO2XVlXj1IJ07zHgnJygJ0TF2fVqwHrZ0AuLRO+JSa9qCIZbX31Gu
ScW2ZXvL8L1p9Rufvk9igPR7YAwRAqOxne/DPS7XQV9hzbLfeH1nPx3kT2k6YgjBPGvSCD8takY7
LY0SuKppE0WCHO/NZ83+4zidSE2FBOaUKS/2ivJw/cBZH/EoetaELAfnvNBqWloVtZBjW7DWnh5v
WbnNjwea+q5uFcquxYIAkZvSuif31NhMhe9LkC9TKvH5qViqqGLsJf+zoSpHikdskZ23CLd/4yrx
EOCkL0J2KWum2yf4eL8vv9Y3reT1kCFDHiGKHKu0DKRooWj+o9Jvk4PKz4hPHnQOTIe2EOsvDKxt
qt1F/s9p1xoQZt8aRUp5EOzw1OMAQB4972jsiZNykvnBFiedGuPTNPyKmPTX2Ug1wiL8iw96bkev
sc+T+LFzRxS0/tJhQ1SrWn5GdUgBAxfVzO96zxeOoTCsl4Eoe8GeI0mGyznyZtGtqBsTyKrQZQyV
ylJ44BNr5T2mAyKkc93ulTL5srHHsrIc/9zX2NKCkSNOhm7MxPSUEw7iCKD5FEK0u8xXh4mv3lEz
9sfRQYMPX+PY7BeX9IKDPjl1F1bAfcJIPdjwVkMv3DaP4O12KZw87GngURLOsbj5nLwPkSfgSh7e
gDwq1oETw7hRdgqSwHyOvnToS4j+YSUU02lWsS6Gy822+wlYjaTvaHbAgldnKHOQw7/0zI+6Y6zR
vs/dtUuZg8I8o448VJU49LGiBsr6S90oinNg0x/hU+aszPYyXkmX/eexA9Uo0CD02N7i7HkT8A8p
Yoizd57RKq4R2XwsxykD9KUcOq2Ja5T4rAyCL3S2wttkmknA+xK4Jjs02u7vgunFOYkUOTBCjKDH
cr66//yA5J6M4ISS9fyjAJRqs6XT2IaZxw9aGGlCL9Ylv3vuJpDnSgB0vcFFyDXua6GPfn6G1nUZ
RK9hFaTnLEa/O6G0xZJYOHwr5dsggHZaADy5nbq26zHl+2NUklZiAViEqFh6XfWlI6R7dRMXmJUt
g4wHuPk4PKJNbMsNyx1Jt4yoVuZeya2uN+0MlMsa+vPAbrHCW6SGoz0f8LOjZrPCu5Z5Jn3zjxA+
SuODnt6bLQF8xUAnP1xepeqmUCOdPcY0HNK3etHqvfDtTZpvMfos6HrSlZ7fhnE9OyQNc5RO6iXs
R+Nle9ykwcCSNPTX65zRmG8HsLPMDmvGpfNVRulnh9+VuVQFU3qantgf0EeRWIg2+s1jOR1jhBRX
kKojfBwyurR1bhlPAgjB4R9RzBcmKiGq+9rk6GnAEbJxygqSJp/TVeQxBkh26te2P4DROZ1W89Mi
E4z+ryLrF2PfDt3irmPy66JM16cHxz8cLA9Jq9wRo4Ay9yO9/ovhBqhVQzRbKhPIa/teFpKphuGu
n1XR/KeUHE4N6Q667XGFQgzla6phR6Zo5ZiokuhT7lZruLfNcnADeEpAOL7sKrt5R77iX50tdTLN
BefsIUZjaTYULbOXh7mlHaLep3HfVPk6hEYC5tm4FVGj7N9ZtwwhsTxr82HB2ZBh+1uwHiSkGTU3
EDNVKgWY+A5ajCS38F0r5LiuepwSsoaW7hZbQ8V+ov4rQ3IxAk4DDA6hGi4xzxHL1eBtiFNmRqL2
qGc7HXsaU6q7GhL/A8EM/scli2D+auvqkApFNU5cws07tf8hNuVBBSroLLRn16ATDQO2v2viwNwy
ArkMw8aRRALcb0xwa+n+gdV1MM8KQ7ZHRgPgoGEWpcYdMyFMMmy0wFLJ5obJw2n0ezfWOAIVWY8t
zYzJfg5EqGuor6vZ8XsukO65+TLOT0fmJZOOfYeOI7SJw2OcwG5G37kmql5i4PzYu3SK+kaAb8N2
xJXM2exM100NhMuOrOxvNHM0Et6TgCTtAwPJKoNScKG77wQjoDT3QRrJnoKY7WQOy4Qy+JgwMkfw
c7H4tAjwOZKOjeNqeLA+1qKIKG64C4C2f2Rw9WAWfQHSskZvB25LWGU3v4lkg5vHZtS2ctGc1iLY
ACZvKvZqMWbPPcTlzhdtewsGNbDADycv5JzTdjCpMgO8fy8Cmo7ISnp/fTaF2n3NmcsEdQI3iS1f
iweS6rbBC6VIwJnd9i0HsTQTrIwjWp8cRxrwjgB9JZFgr2ulPc+HNj68CoZXJyq7IJGUk+1NUBaU
dCavL3mVrzkNPfYdlocXpKSIvW9PT4GDKJbhPpogE+/S0iPVN7hID9Jh4yrI3cmWio+MKuYsN+xd
6gFC4U9UqyPQb9EvzjeHUPXY5XLF+FWtj6JXLZIInZN+faAoF5US2TywKN7AYFFj6OMcUrQ0I7xS
cS3jUbzrvOWSQIsxMrzEK9uxFgTo+XE1oB6txVZzFG3MeK9RLXiGlONzQvV5heRsmq6bU+bT9cyJ
QpMBAEcu8z25IfmLeJLJnk9qDAKKP+J5cJQWe534MzSpu77X3Xa5+1mRb/dgRv79YzNpHkVT7cyP
A1hmpqpj+h4HBcY/MvmSWpS6m3DMV4yr7pCthoaiy122WzJsPKvpFKTiGomxx4PH3c6ZZRjdE30H
HtGzK4jXqLgyrNGaGDr5Em5pb/9V7luXKRODv6pFnvOOuz9N2oXk84Qq3/zwuOI4TSpyfMzNMdzX
oFmaZjBQXTg8w5y9b/cogAL/qJMtaipjziOtYXsgWxljPzERXFKuWck3SI4nregxtT6kOoAC+9Bp
OBm96ofeKa3MWQ/uUPXF5ZxBoMEn4b6ccnvBdyF0mgaI/VebPyREj6ilI8jOncHqZNBNvUoTqqoE
1mwniYzxVpta/qoSEATZX9HhiJLSyq9rSwnkXNn4u0l1r6EzlCoLmjviG5zIT7kZ6EPJwB+hdkQU
afaXX5kOjIb6yOJtVW2+BMd9+G3briYMdwIYeYQFlHoKwXAq3vMwNxmmyJ17SXLTot7rwvFtNabU
CyHosMdAuAvrdnIV9/TAVDX43mPntwQWiYDXvsehdO0RZhSKDICYArD0YmISsdWIEv5oQLoEo221
k7fV2pWb4Hu5+wRr7OCyhHxf5cG6D+CxLIba35ayd2wB2gLwBEKR4bobjAFetcUP+ohmZ8RbVi93
Pqbt42vyUGLjhFYc3yos5jAECySxc41aVU+Vuc/5KSy8Jo+tZL4hiyEwzr4L+PI+ETyBs+nat2+v
AkcutN3TtiEjoDH0FSoeLXTAjeFN/2FFDqWEln4PVpWVAVBd32Bi3IIYyF8xGsfHuJbVNhK+6eo1
75D3MV9U123or3vYb+abu6QzxDTNgp25pz8UZjvHDj+1cfndX++CejgZ4dTqtwcfk6jbV4oamN0a
4cJtVKFRUInoZDFJ4/Iby1WoStgOOqT2WoJ2xI2HhqreYYiV9BowQepln+rCkdnZZh5b2izM0/HO
YU/L2xDf5FwFnpw45TTr1IemQl6bcpY1WzWOQvFxVl2JQlzlHsXoXLYOhfAwTipInf2Kl+uxaqWy
O27LnRZWMQe5OcvtGWdt+E9epEfMRnPI+rNYGOXGsECb3hofRj2jGALZkVKG6IDV3+RoSGxS0J+2
isHomguuQviABP2Snxn57YQQ5QrT5nluhHYcgappf6q1yO6OFH6NPfgOddZaLYRdRjPUiR26AyI7
Df4GmOjmeYIpVxPwQq9lM0eFKDkzhLx8dbKZ5weQkCde3I6VkBeF1DBeK4nFrEGzyRF4WAtOeBOV
A71X/tsH+b5TXcaDJR+zUwJMSpCisSe1d7975qLtXl/aIIVePSRZxFNWexwTvg7Yg2ftdU+JVT+W
GqnZZEjB3qlWplb+EpgTba80cks78zCC+lU3gxLSWD4D5i/9UL0OpPbob8i7gucP5pWgsrXd8Lq8
KQY5bCkeHbc5X5bTE0O7kde15Dq249i7SGJAFYOM/IrlZS/p4XN43FeRU7ivQUvekiIInxv41vxK
IV6kUYLm0JteRhf8thJhU3+c99m+UCxTM2hxpMjs+MBHWO93VMr71GNQ7iiQ41BkY1vm1I2tknh7
WGzlibivK5zKugbvUiGZ4XTf8goPP7Norw8CH3F4epKBwY/3CyYtp4JPuuYPL691ShIW3vJz+4LW
oOdCU7pvExzLmMXAGT7oEjBfqZaehc7vImZcG/KOgL/W/nyyx0FYOWfKkIsjnDfFndr+LT7PZwFQ
FyU2jadiClqDaWuzRYANvf5183Jef+4eWxxosJCcpVsK7V2rJ7/zxUnzves0qx3u/6xEjrEjAW8V
TUVaLsAFRLkwfr5CkeTp2yHcuHTB5xXumAmCBU2h+DW4q3l/bbbONlamEjNdCqxza6vwevNRoQqk
Vi4seEdx38EuaPL15JRBM4kk6kdVc6vuJdk64oV8/QsqcfO9nJkuaQYOPhmHHlUnHygB9993jWRz
Os9E5v1ZjkHUmAqj8NJ0Qgj8huWZejHeQUSczPfRk7REKoIB9tV755SbLuibnYsDc6GcRdFJTPL/
nj+d5EppdTq/0llrvLFPft1d9iqM807Oa3zT7PNGofOQRRfq03x+DNjANXi4uxePR3P4aa7rFQhK
3u5reyqRdLSAWqWA9ULGgEQuHM2c65ZhLgoRfdlFyK+Z5gGqJh8p18viycXYLUqa8+sYQMhUm+gR
A8z/SlHg9YPbVp+wl9fWEum5OILjqeGmGgkDMP0RTI/QUZ93ToysoxIxeXvUBc+H/EGCIZyPv5eh
Nr4ppslWFw0rDKBn4FKIJDGRH6dYDQYSjTnOCFx2/6K9ehoaD7luGbGDpdxEw7Db/tDVySbcr0DH
sSPvyVSW0qwTioD4LYgf2mzKh5+DWHANeiemxRXPGWMs++uD2mgxf4PYKjk8WicgawQ3uRtIbTHA
/SIH9Q4ttfik+kCQUXm1bPcLLxmpwTlT+rVojPO4RSyFkwHkQC2DJdlx+1M/uNOu4FKpaagWPa0w
9nJK2n95hxT0HX6LvhC0owC8QHjtJc2GRTiN/sr8/UcHqqL6zOqAISG76xOSSDCckWt2eM2i/fs5
V1XMeIKqSRdZ2mm+S/KDovwdWmWU0PSnzqv+jv+wlBOva7JkTE5BZr8TShgq4x2OwQHQUPwFjVDG
Cf+aTnHH61EbIQJxdKBgyduMJj+g/7kgWImhGyQnLVH3UdAFnFFcMUAS8D0imPxSn9dnIeoqeM+y
JXD7X/FnLAjH4MKcOLq4kW7Eok0sM0dwNKSpy6+fBFWJ6gg59m6Jo0qurwpsk2IHR8NXDjN4gXus
dVusyMm+8/w7voWaxKmVXcBxImFY/IO2sNGTDWg7kWzsBDgbhm+230FoNUrUaxAjzDNQIiP0CDTm
FJpKKFT6QjENv7lX/H9YiMGqwQDJ+iyo9EdeHE1yqT1JLjid6DMoBITdSmIIxPveduN4GxcNZdGL
KoZ5iNHWHCVLFOJNrugrXADeq1ApTCWQWl4EhP+JltO7Gg02Wm9XOTLglAZSaQTw/LEiuMSPWObt
Way2kZxddu8IAaOBK4khZgfZ4g+Jq3GRbUdYs7ttfiOgloFillYOK/3aQZbVWP3DVKm60zGpkvZc
liqIzirhCct5V7pr4BcYYFoLC6jtE0+536cDm8518/uSJCZKR+5pJOOo9mOq+41UbetxM/XKmm/N
KZCNqzXjVM2gEzLuAvbDcWjm6OX3LVqJlYBHMn65X396sADofHJQuii2r/CZSJbdNPpa0dpdHZKj
1EyI2juWMXwfApEltXcExqcIuXIxlbtK/tevnX2BS6Q7DwRCYIa0gcdL7W8DuFmnBpWUtz8D1IaH
FXjWGYR5OG6o1lbGTC72v63vTMu3eWVqXGvonavC/WS/T+PzgIBz5VAhd+qPatGQo1DM8HgE/WwJ
TGS6LBOckSUbpVZVGjkKMulPH7/IuWAnBC5ine7O5Gx88rab8fQrt9Gcr55y4moQXHv8RRmPR1hb
0BmMflwFLAu57ob0vQU8jH4MbmvWfo9lI0HtpZ7mFzXRZ6WZllT2Iu+SoK2Sa+qJojTxR8VuRIZN
5qrD7QecfTEwVu9l8LouzBHcyAoASCDZZuK2i0XimayCQN4pnGOerhNpcLZss4umKSVlUcD+aIld
gt+JR+OEXrTy8BX3ONziAFBk3DIgiCcDpSFhfO0J6SXCvfxDI8w0bIrkqBQpkQGRfv6GHQ/l0Ij+
kvylb8RNLgOTElmG0vmj9JIVIsduRjFCXV0gyptGt/WdiLvSUJ7CLqDnJCc0EX18Nejd7XYzAMqZ
J7JNtPw+rQBJL9zZpCfWWS5A/hAT2tE2zen/26Zoe+F6ixFm6LOylOHGUnJboq0ma4mO/5mUNJPq
3U1sbiD2rLjfpY9Lrow7mOQhJrUCWm3NZXSgLlPcZX7/PJ5SEXYyLRrrCC8/bUxo8hD7e0QCtQib
TnA1OZ2ImNBvT3AHPRM1MmlIfwvBW/fsAweQ44X/hPpOjKKX1PlFsm0ArbMUr0r78dNPP5/WR9nm
SwHwTgca76tMRXdeUeZaH1H24eDc5fBApOn7+KafmBogXfdG5Lg4+6W7Rhl4qmAtlQ7iParFg11H
kEpschyBX4uzYSCD5C+OH3BGEzS60zyVkaVobcsCggZLa1Y00ZqKiC9tlIx5f0oMdqkmbOxtU2lX
SXUgnZv5F5DwnYjTwYUBuQpWLnPK9xlcJ51W/p7rAAYN5xoSg1QQ9tDR/53GVx4MOE+Q2c/pGpV0
qpAWARIj1+PHRj8+fiLR3R81wpSHW2qFn0ZoSWJBjuDgGhYNoydL4hGKvMTgysD7ZPDHZ7n1BwoE
M9zLsnWJya5ZXIS1EIA+bBbVSE7ZbAXtNIVunh8sxeg0Uuw3G5VmqsP+8+Y3vy8Wdh0A5LYMI65x
lot12dZ6VtXnFl4UBzzA65rOKha31+U9Agz7kkjIykYxnoesLroCZb1DEr2Rj6J6BrQ7pwuad7Ji
pM00rXpSnFtrQOrBqQopDZl3q5bpmxt/dgTnKO+TOPqYBoN3vJaAaNP4rFiwI8YDYLTMgTyqKG7H
XpCmFoqE8wXtNZaUxmPFCIow+aZc8Fhr3X3nHonR1wo6Xz+nKCNhFi+/ywqJggkSkQM4137JQQou
TdlaWxqaGdq+U59i/ql6xCN6Bw5FauxwwbXOp4OmenDKZUkqkIb9aW5c1UoYy49oDL4XboI1MSdc
Sw3LGUibc9EK/wLJNMAHGIKcFd3SK79welbv2XLSXD3k6xJ4kJwOWdcNDKPROlkj6pUqUg8NKkSl
kgW0WMVwHgGUQ1ZdEFm3kbc1cUbqJOYdNpmvv4+znfShIOU3becEvN7SwVtvaZkKeBIc8t2G5Yrk
/JjanctWtVukCGZUTvYiOsN6jF3R/rp/V2d37BA+wMThoiduop7fK4f2YyFhLalX/5UpJlUwDJ+h
yW4j+EncpfP+kO6+QYuLKvi0kE8itpYLTU7whT9SgE9GWobsqmNwCWCCMiQ5a2GQfq6GBzilLjBm
iUzI2ruvEkbOXE4x/IyzFv9ePHzlPivITKvAH+Lw26xmxya+9nbiTN7sBSn+OPDT93DO8BBhU0/q
RiszH5BigSoPbERHmlnvfei1UEm2Z3q0Vshg5CreKB8d52pcUce6rFMnT43D+3EJh5i6Erjs0+Yh
wj0A7vLMuQSXcFVBmPc1Iw8NG6+abP9n1tZMe587O6F6oql9d/594KI65v/mYmxctWstO/nM2Bzw
tKm/Tg592PGnDniBNdaXCQQEltFQQNWOrzuMp5XRmEiCks1YVOcW+tpEQtPdzphpgFkp/iCHCBqI
oBqD55CU5hfZcKSFcsKjWFOWEGrt8EQD+0Wb07+iwpWPizBIgpvP6nKz44aKrX/e3YzBTMEpJhE+
h+h6onZ20sefJRjaN+QgaeAxqRZPDBtOq6OY/8keHbNaasEPFm83bTkD6zRyPuswPTZpLFkr5tax
fLQMlJH105jP/UuOqXCHEIzrXoCZxlDAeI0gkAgYaVcJFdOeG/gfz+JtTdLW7LostURx9xxqFOXp
xF8FTqClvgEypwd6Lmke7ne4SjnNzh9RQz53ATXbtowbEeCTL8DQY7QnemmlGGqIV/qxIMFkX7tG
C7eiLhOZQPvzNPdpxgQ6TIjOXcWFOKQHzFM9k44AwzmBEn/TQCacEgSSdrA8svWmaWhOEWS11tJ0
BE12qAIm7lH1mq0aYtzllk07QEKaooWJ1koINW93nLSAUlrJcg2ifmz2NGGF8DU8U4aYQJgXSKT9
y53czc3KACeOG4KwcRJwUY+KO1/b0wOGYeZJLTsBU/thDpzQzc8iCG4j7xtXfiv7upX0Hrzag92t
QFNneAGOailjp2Gr9fduwknfQc05oDJjaDsgNoqRWMJu8Od+RRau1QA5syE98X0KWvAeNyGPaDrm
H1x/3jbR+msP425AffWS7zRH8acKCHKwCRRkd2Wqw5nCKQ8C7dVW7mVdstuo0UQHBa8u3oOcZt+X
wKO3uqSDXqja71PHXg+fmeK13HauUxcI4OH9OF7/u6D1Hd85PXuN+cYz2UCWqVn3sbjjJnyURHsE
y6BKAUdDMDDF8NyzHrm5lUjlzWse5sYtAphvy4NHVZ0qHGM16XklHCSdIN4Z2GC/tqG5XtQsQOZ0
A4n1d6ivk/kAyorOoar14ss73AQezQRBvdZOiYWMKurqAJKFIuPNI6rNs66TsybERd4S2uQyXPiO
MAGzvCjVyuH3Zxxvn9O2Ckh3nD/8qVsvq3KUhnGWiESlPMxneYvxERLu48XyQ/EKSJytJUewU1q/
beSrEJWAYJs1iaPcnY5IwtnBa65YGFQhuYurQf4hPL3i74mKp2X+vRvXYC7GRdg1YXFELTel11s2
SGP0Q41X2MaYP3ctWahTzWcs1IxtSHqjNpHiZ0dhtNKrCXrTljpEEDRZZJsjb91yZYyWP0uHSQpu
IjMpW7lHH+aE84Y198QH2gF60bgNhkSDj/oolEhajTz/7IA0kHJ14vQTLTQxB6GdYycWfrxuUzVi
SQhoKJxmqtKv6r4T0E4hEFMm8ldm3IAon9ol80ykp9zdPZFp2DGJ8Gx+38VMslIXy+alzV3y8XN6
f3l3KFPWup925F1Y0/Y2oxFH8RQpJQBmDJDT23ANbnbbHeoaQv/Yz47rPsLvkeJrncHfZHh7T38y
24kcHYY1+fUTv7AAXO1MNps2fM0O6kSIT8H0M7DewdHncJbYBv0kvYBTisO2cA86DV2+s7ZDaEHk
i6bnN3JkggbOzdH6FX2Q+z2M9H3jz+apiZdQqVX4HbiaCTo5kkDoxXkgX8sTkaNTmc+q+wbJbeJr
uPqxi5Fm4Cq4lS7BH2gvZbxygFnbaS5of1wawK+0lkHG2L19F66bbiuwe27YmVaQJOXPuCjK7oVh
HNQ3GG87kSOSNXTUL9FMLdNbzD6WjMjEmCchssmY9tH+HkEeXY9AdWJKoc3JVJJfySOk+SY+Lm3g
MmdZ8HeRNtUYxMM9JmAyLZ7QMvWUT0jMLypoIQpMStGFTwZkP+oIvHNTiv+TcQjBfF1EzuLmlc7m
jS77m3kVlQs9UPKeqUqxhYvs6uwhn+aFehARaB7D0SoOJD5yfkqYvhWuhKdyJba5ySPFu6o9lS+j
zeWfO+zv9wmnVMtDr4g0i2zqRK4dI4OR9vb8uIVWM4VQ0dH2bl2UbbrLCYA/FpvBS4+EY/TMxoim
gnjCpdS7WoiNmspISHMePgH+0dEko1XML5CJXeg0R9DZygK2DqOiMIRRuQcMtOr4ODb8M550WXbM
FICBEvAHTtTmVRzstoe0bx9Hz15og0Peb1nFi97HgvaZ4pLGi+NIywys3tS0qLFGyTljfkxRRhY6
liUX8hTEsYY87pXIj6u9fkfzA68H1yQ8c3sREcKy3aPv2G5ZlrbRHYoX91zjq7zT3QAb4syuG2Tr
GjDVB/J8lHqUO1Df7Rq1jF/Yg0UYzwRJFqSV4caD5gClUrVsLIXEhj7R+czU+cuAUrjDrWjQF4i/
GojXB13yME5oxvmy0L4amjhjezTYefr/BDinRY84cE10i0i3uqYzLUHWN0g1GR+PAmiGyBSJKx5k
43Ll5GEho5RzJNiotp7bmvEZzvUd/22GDeS6KMnUGv8qw9MddQiY7dk2I37x1nR2ObFWy8KWwmnc
DkIc1WdkBze4cZqIpPcfviug1FoZPoU9UjGYaHu2piw8oEpC3P76PnSOFAzyjqyaXO6mmJJTkAF9
GGRDvMZYiX3BBkXXrjy7loMA2bThNUwZ3i2ORbx276wxrHYiqRCZpk+NK9loVSy3HySE0rGKxvjP
6vIHIpf9rccKNIsca85018ZwPgJRraLTdZ1P9kJLyiP1E1pvZhopcjclTbZ+Sn2wt/DkupQHjbt1
rLMy57T7iEr+ISA0+QcKm7U0GppEsMiToqDMyd6kte39vgENdCFpW9TjcUGIs+kjgMpk8rpqzuFz
WXS1y8+Iu1m/YTvyfQvyD0nc/QiKhja7uUwZ8lt6PEYQprlAsEffoZMxrLieskg7tRFH2++niwoD
tGjMSuKfab/4OzXCzamdY/MzHhTTQnFZ0gpmoDoeG3eYOtGoCeF2OZAxXkcfZCFFy0vQdGng9OjS
z6LjQSwaXxw0RY823Bhf0P5x9d2b+8sidImiEBWUGm9fLv8IwUWAXL7N5/ZIiTKRFe9QSWjksJoB
RNSvJFDMhvzzZILXIjJuIly9/AMPr6IABx2OG571myNfk+H2QzW+RBIuWXam01+kO/3Y7P7bAN8Z
Msv0UbfxyOIxSsT2PDUQu36GAVQke2m3UzZdhtkj8J8XqB1Q6fb3sE32pJKegAJN7kIFa4zVoagG
nb9wM/XF0v2DEJeBC35tjDoFkuKGoNNaI6bUz/pi/Sg7Z3BN5ibDsRjl5HWhtfCv5vsW88IU1WCz
xusY52tGJiNsYMFqKTfyVPnIDRwWCbSlQCglfBksRIh81BLvSlP+EELfsBOGZGNhvzKoEh29A26Q
U650fzmMxy98XcJDqAFx0TzgR67nD4dCo8rBVFwyi6NPTTHzGPNawouHaUJEIdtfpDYzbo3OPcBQ
gk/8x0Fmq9+62b3IPPOuV3aek4NGtMISqdqAYF4P8hVe7gZ7PMqld5xrTpvz8hYZX75wf7MW+4CQ
gKzpMMAZ1VzHh7/YmE4w12Vx2VTNoe2IIcmPq3pcqZ/Ujj8HO+K/XA4Re+t4UN4sKukNADCct3nR
VujRxl+TcVar2oJnNDHT/Aa50gytehi0ozG/J7TlHnBx9bD3CN+OJzU2gXEX4ZdksGw/n+FiRlIc
b857oBxAM18vPmQFAODIFhgcRYesbKS+4LVHMhARR5U7Y4dtFqcn0392u+XZnueMN91jZB+L0Ru5
sDQn9o5vgg5EA73EhgEabhXQZvREt6f/qilnG7MHeHb3cp0g8YILjKOxfU4EVHRI7nxcdGBrjyQO
2Qjwy3FpCRvRTEhDYFGeRSfpCfbKe+HR/1IZD0D2Vz3U7miUCQ2DW5FMRZaJ6sPqYtmocCcxZkdt
QjvC27eTNqkFxoj7AnOiOtpFqUddc3JWU2ckwUEHaA57nRmrbMn/r8yMVRod/m8JGRVFadrAYtmT
wy0tJEEAakknxHP+C9sn1XD49cX7lOfqwt8TuFeVbxfT6FSg6TVkr0gt28yYboApG1kZjxkiW1Le
D9ob3hL8HxM03Q4RrV8gTgcLytxs3L2nFAo34mGHuJJmyAMt/7xMZE7wcvZP8OKDZdaMF/RJHuvG
fLgL9JXUXi41nX35IqRKHTYnsaZj5JRNgJLrQHgIvgYXqxCj0Wm5+DFwQmj37fMzZwh7z99LEbGG
616TvoWrJOefQAi+qxn+wWbCXFOiref26dh7Mt792uRLIaLqm2CPncCtXJegI+DtTFYSJdIbFABw
frLcCFphhJcr++SsEOnicsBKLTz60/M/HU8VlqiEgRcGBZmlCqn9ahj5NVrl99WoVgC+zu3TLvCc
swMGppOghGizfTDhmquea1NrJ4dLt+xlQ/Qw4fKzMHEEmEJy/tPZS3NbJ4dhpRlmkxpGA+l8xS5k
Hf11tPvTRnoYME2IkD28iLJX7dkeEnR/OVQP8gekkBxzaOJ74uJwWNcCNwrEPBunsug2B5g5kv1N
dtxAetroEBc4bde2cxFxJCCQkaNUW8kxOfpJsf1vA9MUosbtI0m97hyXzZCzMFwN9tGB21wHaY+w
Miv2W6tE1TIGwWSiQ/lbCv6IIvpXHo40Jrc7fHmYWd/Mzn6GI9O8U0xAoSDylZYcA9GV+FCwxtuc
b5XoqSFm+N/TGWWVuGaw9np3nnQH3KK8oqeRuqcAZFZ/SWO5o9+RtZLwcnMkXy3LmI+YfqiqEhBA
Ybg6o4QiiPfNRU78cwkxAdDcxj7BCGysjkPXwTR4n89kYkc13RVuvSoiDlDssS1lz9ji4Qoae52e
erTAcGbD7lHZTIBFn3mNGz6LZ511HBBCjonF6T/s9UCBdTW6YSDCD+jWF4T7ZGcZrV/ilLJKemyZ
KvsXhThlW+KWVUls0aQt9fGpfT+hWbri3AfqQIqT8pdssS4rbD1AXcFicD7BGai3F1TBftZ7Ri+y
k3USUdD2G/UdRMD4tGlJGfpztVdBjaONDS0ndYZX3VXMtc6VBMnIoEtNZaE3gtGP8OZQ4mZ0R2Nf
iXcBFL5ndMb07iW27XcR3YnEZuAWrDXSGRwHt0vy+XqtSE6XtMKZRlTumse5I7Oe+rhMqnykCk5n
iXTkQxyndKKM4uzXQbJDb5I3pD59C4IvrFMQgCeaWt9lI08K5Y5AEDfEa47Lw4PtkQDL+7BwgsZT
A5OxTAHA2ERHg3NzDBZRhVHfYrsQU+97OSUZM9+YBZpDPp1tH4+xYvstv5OaMM+uWnS7d04qENf+
uFRj/swrY39jU+u755EgJV8Tw4CVBlDm+oBEfAYLDz17EOdnXkh+dPqPxfl0wBWEc51CjpKghDiO
EB3Y9PcRMcRjwqwweYDcu3/G2QOpmVhvi7EiCWB7SphtmYgNNW1CQfIcRITzQOls7FO9F2bMd1fH
7g+Ehr6QKgbEgY8pWnlef3Ui3EISHcNoWW1XJdaQX8ZPx7OQ4v2iUNctw3k39mlhZ0t2vyW3i/Y4
WEpLg854adayF9rdjyMeIblIgSCsUCqrvDc49/+AZJuvXtGDEGDxNawdWmvs7HDGMCy9hq3YNvGM
frf0SfidedenyJrZE9Z/ATLZxs5gW/S3MctS/t7VwpxkQD2n8ETrPpbdMALy1SuLkCRwLCVQEdhO
BZH3fOsA7fC4v3eNw1T2DUs9bQEx/LdSMvIFDfqdLQh38GPFwkk+87+SOrNRT+3yL29evVfbCzsG
AOvvsIBz/cOYpdtqDKjLIRnlB4tGvYwGmSDdx5eaSoqY8qzBdvaLzNdL5/YaaH/Z3BYKwRCalowG
16vwgXqEON+QMEUEhRsMiQYBB/PyOeO57nuyDj2KzzuEkzSUcavGH8zG+A0ylnOoDUZRqLkoT0fy
RwNfVZSTw6Q0Zr3i8k3OifAMwp6ujlAZe1qYO4xc1g/x9fdf/b3nprELqpB3p+W/qLiT1Butzd5e
jMhxx04rOh8Wu5SQK7e4/Xe6UgVQl4uBh8VyqY0waGNXDmBK4rl3mMDupBN0KWnMeJMDHaKbcVMG
ucqZ4Axs+dPczA+c1LKB9OxvxU7QyXQ1JA6bQdGPcfQqmfhWsnehEt/MVS3bvvRAOVyR19ZbZayQ
Ee8UMLJrutuZybMrlc8KN+SyhKTQmh/w0gMHmwuyYQNwGjkqSnOUVszJp/cGG+bq8XdhasDrKy4d
PQnxzRilObZEGt56/iA6nioFqwkfpYzrVzoO6K71o8oHm1J3xgJDFEE8IsP/5gqY5sIPJnjKEcbR
CNrTZ9ozIkmJBCVjOAJEzNfAp8P4cqiL+ecPHzM0znyPTk+n5qPYbU3+c3My2Q/w9BkOVBsHm2Ds
O9r4KJUcVNJUeEQ+0FP6FSEzgVH/45o+6hgpNS5FA2KIqtPDJtLl7vcSY6cqt92IReQcN4Ln5AJW
KnloBmjznb95jy5ADWT5V1PvNzn/duUp0XhRhi6NTg+zh6iEBbDQ7FUTBNyezMD3DlYvFu2FtORa
FW2EPCunPyrNgnz6hgX/HufgPSBIZmLc2NlNv6BzZxWXyU16H0z2FZ4Z7oZYYQ1XKsItH3dzV0MQ
zdH/8YHM/bfNSP2gRkg+sJzZyQSMevrwbei0aebStUwuYQqd5KEK/pqAcPWVyRfp9weOA0vwNtkz
As001xSItrrELPxEujuAbZEJFmKgyInFEf4c6i5N87YrWNeJ0pIa0mEkblHW7mfpd37SInGXTUoH
ILxDEOZKcXK0fhiraSUa6YQkmxEgJ2acqR+Xx41TR+PpNUPes2bfIT50OXK7CmkmHXlYfYmCpxL4
Es2uowMWf1Judx8oPmswbRCx2RbOWNfZW59m53UfV7g26eX/SD0sOfRzkfS/3qfJD20LPq7VWQct
0EXMWF9TWXYvVIo8r6RFN2xyAjTcLGehSb398mr0JepPLMQLB+0Z0pmbVKjASsQphssoDS/SyfIJ
QueB7zZ91Ua5H8p27UhBZOclglPTsMxpqcIieEyAAk4XM/0MGL7Zodz37YCJTx9qbNSFr02yBypG
qBAG6zpHHNeVxSQ0/+8JOHuh+4POkfWDbqFk8Gd2+74EjGSOqHWi2fJ8Da5vFBVuafQirDNfigHS
LWGV/Jfv/wF2j+Q0FyEKOeGwW4KnClqlnjbomLvxLV6IPGzj4qa+ESC3AE8TKx2reI3udTIORu5H
XJQt9VygQk11Ox3NyK11hg5rFOECL5+Z3RtkZNMZlIj2BGwl3WUNM10qc2UFSzfjefPGCHkF6nZ+
8b5r5dBHbqKRvMBZm7uRxLVU2tBd2ejgM2VXmzxRclThkU3NtrJb/OEGacTan9bsBbTIPdHLzKC1
HV9mxmUbR1A4ffzJh3LTOrBawquwCjS5vJMQTLexaqgxoTfs8mjTm7wpMIr8oSzvCl30qvag7DM0
RZDU4AvjhpXp4sOldtjs8v+CQcUDeJVo7fa/Qc8ol/+kRBwYdyqEvhCgUeAEu7HZNwRzHsdmtPzo
ymP7tbEdfjI/WhNf3lPX2bQBE5zuh1jW6tmfg1u7gKCLZU2fwWcz17vLaezg7beGrK6ou2/EKl41
FlYNqbZkg/8432t4H+X5yL96h7NSmomXiIipWwIXIEi2KoQVw0hm2Qj26/FliVRLhWYrNrIDndxG
FwiaqGcelWkJudot+SgTlwaMED+Skf+5NqGl0SXHzLzHl2M6EgnPsGo/WUAP7sylL5tJ5OGi4NNI
7An4mXbLOMqBk3USiAYVVMI6H516GqfZ9uI00iYBSLCQMFRip1uTEg3BcpL4Xk0AMVzK2dHrJe+W
ZfDWYn/Qfr0tEDH9/ED2DB3reRbWdeeW1hq4ooXDZwWha+c/i0F2EmdjsxEs6BCA3zMtgYbyS0aU
ZpYXH2hzgPq1VWGdwbZ3SNTlgn9c25JguPGu/OVB1OYz3JX1OzscsscU/ra/g+b1e/EMgrQRtlXI
N4eRzAZCUD18DIoRR8BnHXPL4seSF8tLx4a8U4XRGpHhNIoZ2RJCGnqd0G1w36+6fg4h6WHySKTt
Snh1WF15uRiM9RY7bt0yMT+giZQHbud39RSSdcdcHVid34sc2vnvzyztagsbu3zfkjl8DISGgl/x
JPUMBs8X3f5s8gCeJSxPweh+9Fb9uN6y88rgIdzA+RmH1KkHy6qAb0KbATSZwSpOCgkyM9kdtWUn
26kZsPCxVD9TH+pYi1caf5uw/s8H0JWMjnB0B/V0HXD0XUdjww3I0AYcr9MLqzEtGdxG1xHEG9G4
3jgQkQk6aZRt3t62hTrX6Lof7soDDVn8vujVeyhxGtXF+yX0SMq3Mrt8ga4bTBoMEan6XjUCKGR8
jKOVypwVuKaDuTCxDMoHI6Nh47gSeJQmWnzndfxKQtIMAfrEFIzV7cBtgxcd21xCGe+qNFoBp6ro
h03acP5oQ0wR71mr+Jn9/7xqE2wGClkqxbrREJ3QId+rmI5MtvKYvL1EX98Den7ANyrFV60U08v2
kcYKuXt8FgkFCFlq+3BEwwjgdDZXyIebiEZWxv5oc4JV9aqZzaMjcdnSsgjOxziqFiQ9zae+tzfV
/rW523A2W8GYt0HvRlQ2MNmyh9za9gbJFagsUwmsgCnI3RiLI1kM5qY5sKtUXgME4lt5VjUv3wnR
EM9ITB4ZxnZxofg/eiJ7Q0ELw/eqr3AB99oAYtQ1j9p5mb9Wac6hH81RMJTrcP9PDU+U/UbsPtk4
L12zkeT6KBP5subd5HcNY5D6+IroNLKbFQ7pVi9AG0hkCk78KpN+T7Ss8uE4Xna6bdIaDfopVkFC
A0XLHkAEEue8+Dz3b+oIdAAx72KJdwMAjrX/8dgQLjRCq+eUTvKH632N5RIQRQyiB6MFoQRsalO9
K0DEUd+vUqZQkw89IWVHFAsddX8o49rfadyXRCrBNAjdj54lKt1tHr2sPJJazZ1fPhesuMky73HJ
LG93cPA/9V0TcEKwuChOe9/A2rk2JSpKawdSm2kzoQg73yv8o1rixb7RbtK1OJW3xizA4VrVUDJw
NOlQsj49bb0ED4I/FWzqFz8L9vJJJrO0F3uRfAXITH3fWmoNvdPpbfKTCdjP0J7QTIbFlYZ8Rgnl
u+yZEkwQ5YzPn3loLb0GGlbUybl4ZgD84aHlB7mRMw8F/r7GJHdbeInS0QrxuvW+ggHBYE17wcBm
nfYVSU/q2ZRkh130pooSiRxiNvBZen7Dpv1yhhpyOU7OcHJcXcS6vCh4hnB80TIZsMbPDjkSWpE5
enb0KSkBueh4b0RjktMNXUSaNRqscyLmQHDBblxtN18lfmcKbuaPlCGwlCDjUKkA+KG46grNYz2s
pX8CSjpfrspTdMEAUriCLVf/dpB8eADTmX9Tzyt2GRYlJBJ9XkVmdjm3kPbjI2Kp7ugkfgucwqaV
NAEokjQDLqR0cy75DFXJBoco6LJv44zTMsPW+/rjYwerVaJWT6rAshg8eDW+aMypewH4LRck1YPR
E7t9vMi3stz6u9RsvVKZOVlCaGSo2r6OlpjwzjnUiE7JWJHjrmXT8Ns0Std5/mHWpEtVq/B6rrgc
3XBZMVsUttOmglY8gse7FRMtPy3JKiwAahxDhImlZmpHmwIcE2Cb5DFlf6Db5hBAPx2CEC1UG+G6
hiGbiNLc/HII2JCUvM6blGpZW3gNLLE83FwJ75xlxvXnSJlpLwi9xTqxMRD20Nqj4vDLUDmv7rvo
xeMlM2p6uCEKRWZvqyipiodi08DTaM5OY7Hz5f0zqmmw7PwAVa7Ogdyxj/otnOnpsalSxnBkir97
Lqd3umQww2BvCLPecrx9VX5Qiohl/ule6ynHqHeHUD1vO9hk+mRmsTVcwzHZUE4fU43z4ZWpoGQs
MVzQ3NXgoU/ty7+kWqQp5LocORwC9JM2rBxEIyzaTYJEJb8woAQENms8+/JHzni8GGoEU/HgWYph
XzLUQclD2H1qH5o+v1zhIG1Qr/8hSkHJ/w/m8Var6kfvsR0vbszWfdTTOdzWFCZnYtqhcadGS+43
A1RSbISuKCvMd1C8z64XTdByqR3aflWGAgUCmelg2t/hSPbflgHsWq0gXg//JsSrGBxm8VGxYKS7
TXXaEvxqd3k+ntHFFGSq/b+yuORTU9137QVsYkKD9x9eWRWtNkaxMUKIL1Y9pQrkWmZmgJNH/17p
Ty4G2Jgp9mdXm8ANSyUVMNXx0INju5qNA4yBx0xQRgJChMZRdxrb3Cnn7O/ZAM/dtsbFCqC/z53L
4rGklQH0Pwuf6wpa62GD8lSHzJs4W5tbfP/LdUwsGRAElw9vITwJpV+nDLlTUC/Y/J1KilM8O+Ek
D+JXer8bPpnpEatqCEG+6DllPXp8PKOKwMZHRFTa9awS8bb7AbAyFqKtRCr4xnQLIomM/oT31xcR
1rqV9Wdll6IF7qoH3I4/5SeNtGnHAIsBNiQNweAug9GvfKNQPkISE5czoG8bHCvSeTgLZuNN5+5x
/qYXPCCJY8LMcoFlBt5RQF6n+gPymlhCjQ3o6DFP2d4KSnwA4Pwbfejz0Jb/3kGmPrvLBI4XJSIy
I3mxaEeSeNhjrOjgprVWv4ql37E0SNkHXzZzmX+6siXdTVjzRMDQ8zP9/QdqL6t7s2wd/mNvm+gj
CzfQIsSetoT2wKfTwSaeU3xmgbEehy82+XY3aa6zIIlVDLCNqGy8LdsqUCQJKMul8wZdOLeCwNyQ
eWBRmW+1chPDv1fR+5ZcqLmVTI/08HL8GE2+mB80W80uWPG7yfZQp50dBgwAILyRUONXTuYtQogB
HIYeQ1nEKxOsDhlQgSoRUDMd+GsgkSddQ3OPjHkpvwXzvR6FjxZ8T8m1yrnh4ApWa8Wa7ba8YD/Q
bRCHEGFIXoEQROHMMY/NgF35osQwHWbsVDTBNTw+aMPu1JibYhXg5jx4AxoZyOj3YkoPJOzBg8Sy
NKnE49BYvbAGw9i5FgQMUxJWKgqoRbiMBOi1d/bZq4/S9TjAy9FUIv7nxyEAa8/Iwlxqo7XXLcY2
XOM/PGTM9eFCwz5ch2GL607Am3Lf0PjkE8d3O9nAp0sZiF5bzNPhkt0wHnr/ZlyzfEx/xg+o1Wgo
3l34oSlYbdobc0I7HxipL3pYrHGOmwMtdUlrpnziwwYLUmOzNrtGaQEFubxKVi4vg2gb+AFG5SwI
bU2wluC6tXPY+bacjVa+/1p/Sg+BupUbjMBZDCvzzQf1ZmEHr9R7dajOupcwJFDusKXQYuJvDYAn
scHqmC+Q6QtaNaBadbDT3+w9lhDyZ7iNki0sogxTJ75TS5nOvCcq7aSP8neZqpkb+Xyi3YDn3leG
R7TbXBaXttnY3/ZEMHPSphLfLVYhHVoXDrm25TrxGTZyXzfaGA48AoFERwnCrf8XC4enagxLxLk5
PymUIK49pielNOnhtJzscXreYQMulLf9XJunjxPEaqguHSxQRpsT7ASsoch9sd1uSGgRgOSJq7MW
Q19cW69FanLXBiFKdcsSMqRhtXRdpQqway0apAzULnPaZg90oah4Dpubl8iHO0JsVCdyjp671tTg
e6NCl+zBm4XRnfq4u2hyP2hd4A2/Yoih0oKhw3pUOp6E21hoTZ/+5zn0HXNuGGREXe8cc1WBBu0+
wweSbFunp5BUmEbLJVHFykPdJCW+Ta1qOG+YW7+5qa2Eo7OSlC45AZ9lqyHlWh6KYAhG8PEgOMCJ
CCllFqiQM2yIjl6z6qOqBO49SvRbMtjALaI7Zv8G+zYAMgb7GNLvjUeVVzBEZkz0llgciISVDNpq
Y98gUi9n/kqbFDenhDnQCxte5a3Z6a7u63FyDyCznRkuaYRSLOVL6/irucGIOw34JVqY43odzo5q
bd7jCSwvTdjKVaBZUS+pU5L21Mz2HJFFcmGsxSwsJomPkDh6LTeYBfSn9fqRLs+MZkrd65RM6CU9
F8+VdwtE/tOyZSoLzBBPTx4DJ80O4pC6MgHLfKPALoOH8eiKsZF+43uL1gTe7JQAsa4QE37WFdVJ
/MPGzMxLluv5DZdYF6RjlTeUP9eQa4UOD70QYciqt+0EKxarvDTJb61WQ0REmDOP+tMag/d7E7dc
0h//tq0gCEolNUtVLDaBOzyhb4xqdQMX/+8KqaAINz1BzvjBHUQ3yrla/WzzqY6tyOAZXQcCnfRC
RWKrv+jQlzuKZuK/hKT+jm5RvDKalWUn+vfQOQt9gDnHMcQVXA5w+KGhYTeNk7ia3DMhM4ZqzHM3
Tp9vsqpKswQfmoxLBkBw/rTiV84hgBLrHpR3kaRV8ICcHo07yEwM8nPmP7VRSzrQlI+gmwyIVSBB
Znd33ZdbOfYu0ExSUJT4XLODmog0p/xfHvPjyOEjkGUpFqswCtj0gW98aDi3nGIa34VFwPKbRJ14
/R8eifW1RSYtYffXasRk5yfoIWFqz4cD5JQ+wCysjUcWbdlc4yfHY72s4YqSwzHpmevLi/iy8mDG
i+Gtzxlliox+WCSLPG1pne6rYOnQk32ryGmZKuBbMR4EPwLhV62cuvUAYAEpN7qvlFhlqHUsPoxg
RuA5Nkd4b+TvG4wrafzzSqmkIf9uafHnCyJaaQwKgahaUxSzv2L/c9InlzndfnP9LVUBVtLIJ93i
5K2zYNkQ1bYXSc98xNndu/60GgItC2NDX9v7evlC/NmRUJKpNmG6mzEnb1WmxE1iPOy2adFMlSF8
43xw0XQAXQ+dLdEqXvm3PNdVXHWFm5b1lIlvw7e7fKIPTeT2a+ZPhRG1RpNsEpdjxe1Ub/K8wrhS
G5qLgPBCBBaL0cq3YQ9wWPiI9JDYz55HV/GFS9fERu2DSK8+CFUV7Tdw8xgtIzMZXl+bozCEmUUE
xZrjrQU8GwOgLJkcALS0TPYS/EuXssjE9QpTE/cWDZGVWOqMJ+RfreiD7IJXdVyO6QzK0w2y0hzz
LHbZPtj4wpH1+h34sfj/2k5XmxKIhPPSbPNCEHWMsNS0gyLlYEzgsaiR8nqtqpnku0MsRORdxtQT
gPKYD7Nnj6AawkVBwjwM98GhDk6Z+lhd5sqEMCDIOOOnEBuq0PQE6gW1Va/p/6T1wQs8exOyk0wR
+CRcX4QlYADFByLJmUggDRP/u/k+QeKfYHdz54om/N6uHyAbQ0IUBxGpPtHsDz2bOpUCuJ7HENSg
IbfV5CnyxfzWQ3R+e6WWrBk7YWCKw+Ip4u244TMm0xq3SiTolB6x52a54jKH3n3tMNg9q0DHNpB8
ZiiV/3FVzu2mkvI90foO5Tw/Y8smqMcVh913TFTbWifth6wAcCdhtsa/WR5uvNpJxuy1tyjx0nDh
Qst78I1ddA/0w4Aj+V9rBBS/ofAN9AZkAyYIUunmWrK9e+NE97wB6RtJx7aM0FTAuhY2z6Z1X5EO
MK8Vj+nMwrYI6FT9bQMg0pfgZJdhUPhOtzLyF7pDYATZ+aTHBOPlyZPFEC/OuZXOpxBGR7Ws0qw4
Ne02Bi4+2sdTo32c7FVO+yKKokY+kjsJMNX3A5PotOFM+nIeP+iGJWndYTMVJHgXTsKSQQVT1hLl
Wv9hDgEEid5kvNRPgMoAonurphGCNvRtRcqGP8WfyxYVbFW9rlvPJH4Df7UEuhB5wNuwJlE6fly6
IhvNoIhVKv6cAF3gWGONj1dtVx/jvA4PyVsBOkxMDzkQTQ9qAyJaO+r9Gwn7gl2BVAe+O/yLyu/q
Otz4kNfK8X+j5Dm2No8/Zh0sbMsTYoLk5fG5Eed2h80JO0Pf05pLknXeAPAHBK4DclCEwydZIuIc
L+dBV72oYSjy8JtXkEGPQfG+lbbOPXM71cE107jZpezf0NpCTO4mDqBJu4LpsQVX3WW6Fjr1FGW9
vnHtRbVoJSc6r60qYIHqgopWZeK1IaKCG+BftUnkKfcyDMl7BO0xrnHj2e/T04uvb+iTs5R+4fsZ
9fQoiwZprAgqBN5WQgyjVkQcgT2Gtw2nzMvLOvQaQ+q8zevPI13hxDhNy3WpZOqjR4no3lpMLHb5
YKlpKewpirOBvbcJXyZHp+MtxhxQPN/XzszkQjl7YZNwO+RbO3doJfjrvq3xgSlCAuDKHecnRCpu
alRuko7yn4b0GtQCytzNO8O5lq4/GirF6coJvHjbJ6SH9QXMEImma0oQbDrBMDWbDzbcDyUntRi4
YlhcXtCfCGaCgsV3Wj95qoRW15e8PCTa+mPEeJlzRYHBrmbwZ74xkiK1WQmd6X2h+QeWhGUWIrEZ
l7a2QeYRAyi2LgWtT5Tx21nDz/5Q0xfSAot1QOodZzZm6qxwN3LTObgxG1YL2l/o0wDqvLfJEEfk
n09RzmAhSjvk309j4cKDp9FpEyTxpmHrXUMQjI+b72I3n+STsHzutf6JHkuchHsARjlcKTNzRhAF
dddlLy9QHA6icRj9i9FadYTlcSuAgrJEdfv0de4oSzB9iYIwcilfQ+99La8L/b88s0tIwIVAYS1b
2wVMBfYOnPU7iYuCULSdX8oAfKuMt24DNIOKDMO33P3k/LHhJL4gk2rfOtkkvqGGMpkmTb59pnnK
+ZAaFFzdBhiF8devV0Q28S2HObYRZGb0ZPW/Cy7Na6C+xpoM45XPZX407/1lJPW0PFh6EqXF/o3/
38p/D4moMdAA4+/lfKVEVpzJhY9Rl6AbIOsj1SfmYe2sH+o74WU+I2+dTnyM62hQDTsW1u4N2qvw
Hb1FJicaqYe48ZPY8NaKv1QEI7JFCS4dNCFbUfk6DgXFl6JjE/1kr4ehM80WAUqCiWINf9vjQ76K
3V9bSH/IKiCkTfrlBWTZUin2HHMxPxv3SJjazYKDIUXqyxF0sWWoxuzhFRmkGSieVMTsU/7aRsAq
jZZmJqe041v0UwiRF5dwAC4UOkpHlydM3q7MlB9DaQ+w7yEc8TP0FYp8z7f4xhkP7XG6bME/nLDX
0rVDbS685yUU4C1+H9V0zn3UN8paAhrjvve7MQKm37dUEgfCY3ZP5cwbb3C7TN28fbIxKAjKnPOY
KfGPOl5w+ShlLFIcwV92QSuusUEO1j6aeVDXliGbJp2CduZX0EUDO4iS/ahUmZAoO70iNAqDABxY
gfv0VGW6t03mBRl3Zh+7ugbDG5ONOOUkTndlaAlDGlwBKBCOJUaJVbkR3NCnWLYA4UHNEYwe+M14
oYUpK/8ZCiWcmnHvtdrCxJ4BL78onmW9rhoZLPIVwnNwuNVhBIlZG2Gl/S3X1fbjpRNnRitIH8s3
wQCwb2wKtaDSYOVipeCyD+HBa/ooZ1ikK9JVfDe6/i3smK21In63R9kXCmHYFJ/CuiDk4o5xCn1R
1xVEltcoYz/rwSBAp3qKhuUDow14vy3lsT0/6fdM3iP15E/F4bX8w22v/Dr7A3LArEtzKtri0vpP
ljOktqmwf05ImH/3O5m7TrZF10QyHB24bMMNQGOe+KanEBclex6d1E5N+nAYi2F3nEVq+6seJi8G
hndDV4QOJl4g5/u+IHgmTdbKQ7PXOzzVU+EqZrrX7hQ70cOSMGhCrBcFv0b2tQJL1qYMrP/rsviE
EujNW1JA+1ha+rv25+/0gl4+7dfmJuaFSOv1qtyCzwAhIEhIz1Tv6UhkSRkXmySzRu0uHb3KGWFc
Ib8sZMqhwVdoE3SOZOq6WqMkQAoLHb1LB71b5+/t4GJwNE+20HOoZcO3iahoKw0/aH6oeD7baRqr
OGnJ2Ts7b+XU+ut3TEDs3tjHD6/xG8OgC5fh1ydSs8o+TKONXouegon4YCYY13PeUh7FQed9SJSn
BAZGq+AK11wV+aXtCHoniYKOsMIiTFL1AEkO4HK8g1VywBEDQxClL6ZRS0j2CGUA/ClWiucpUZK3
5ZM1Jdf76MzQBRAqSGnOQB7OBll+/Q2ImMz6AalKGEV5pVSucvNjs9msvvbhq+hOP7w6Dj5nsPXe
txUoLPDxi2582TsF0CPLqOB6GMf+sa3sp12FmQFY3ovGZOO3P5FQ2GFTFgGbt5afuKoiD7gotaon
jYLmulathaZKYIyDWcNn/DQEXsrA/ApKpa+wFsIl1v7GsOXzE7wFj+kcE/MqYJPv6F21S7VYqgsj
FbF8qPFwXYmjW8vP4EKGdKJluDp6IS2/zmHlgXK5OsMLJo5pkkM0TkMf9+4ARPHlFirzSY/j2+ER
bGuAQ1/fr9TmNJJusi+N64rIMon+0exNNC2vzy0kLxkhUK7IGp9/MQvra4jcIN8ZcIBj2TfN0vz2
JzTcarVurcJ3PgKVTwXSDKTNbntL9kzRBQzD4iTxgbg0DydbtPPNmz9zAdyjjU6nmBOLmAT36na7
8Y4zU1XpY0lr/jMibOBXNwLMncMjZxM0LofVvyvWcOzYCn1E5gf0PnueUByYIvDUGJrHpHlCXa9N
ZMDW5NBonpPBOegGHnJpJKEJ/e3G+brczH6LYX9lwVCP21TdyMEj4J1pFLUq0MSlRPf+l8mUOtc/
xuJFwdnoh+gYyKT+96HkNLT4+SnaANsRs8MJi6U7TRC5E1dMULlPU1FWmYhZ5qQ6m3wt4Ntk4M5+
8JsaY6bi5pSaJB5jFqtIFT3bY0SRVPwEQ6r37/K5Sx00RYbMxrvpOY8cLEJVUSeQLsBHFgzS3Qvk
PV6qnqYFpxMqh379IPSlD+liqpGs++iHKlCuggI3UYje6Ed5mzKDvEvq6ocJRe6QCEk0RZQ8qBWf
wZYafmtjHTagOICBPt8vDOPJF4FX1SE016fsMQIuQ5kAOCwb4sarWFzXmyOQyWqQzmwF+xMMqftQ
Wb6ndTgKXH2H1fJjMvKY2xIUMBu3pZ2SuwRf6OlDDZnn4+Ouq0TSRcZ1NSVyEb1Wmy9LshbzBioe
nlUFjLtaXCYC4qGtj5eF5LfQx60z/qodmzJbYP8obEHcWQGzVZMS8ShVVf4uMrySquenYroT9+TV
f0ANuv1SIisajenM2u77lyoAVhn+vfKRQGlpf3qeB2tqZmWeySEfYxOYzEOlC4DH5Pg8hFsRALwQ
hVkrQe+roa2XjodzH7Q4BATYSh5DSLNTNL0OJQDpyT+l2tYiKLpuoWW2VAM+e3eUtXY00mkC1yKd
5xRSA9XkUVd/WXmcZ0y6HLTXe5N91ZF6VK6cuPBE1ny93lf8GvlnEVRBqnm85C1mBoJSIWpr+8R7
80QR+4XGDI59vpVx+a+1wk0ldQw8m6WCM3rBOwv0AKJ1HYiOq2J/7ml2M1t6ddYEjrDie048ufov
qXl7MM50fKg3+JSS9qtHHpPxWsF9RFq72RcFCkRUKgMVRomnGL87z3aE8wAEs63cMVoeLDvTc5Da
bobDeVOI5VnQJsCja8HyV8L2ZemGWDByrhhbokmyV7+zANSTnfLAoy7u00KsqJyPSUVo5OqZcDzm
D0SZ8U3Ohjdw22HrKQuLizg1dUNfMr6YVUHwOhFXSCU7QvdHllOL9asxGRVkdXcIgzxuXr93jg23
i8t48PucskCKuI3YaQptougbq7f2L9kFyrh9fsvDukqSpm1eCRnYgnxHMyBJFkKm4+UeVXyayAVZ
MWoAtmOCinOWLLIlxluEePGJcchphI37jCBmYmXTowQ3/ldHaaTfVmEw0IGscPj5EWeQ0X0MpgaJ
71qxL20U/GIuBkcOWezeBdjQ2cFBAZqI2jX0eVBRtmz46ACGZr5pc9oLnSDiTSVNnCFw+sS1XRVn
tv9zWyC5VIdaIQfbvgWH7q+hOk+ZZ61uNWqoO44yCjtFsq3uyzwY15s5fHT4wu4AG3tUo27tj84e
m53xkGeKfBQr2tm3mQJ/5SWuqPt/vJ5vdCDu7VDMfeIOuV8gmQ35LmAe/4fQ3DYXW1xkzGtJDH+F
1SITYJNv3lpSBE10lCX4JGsC4lCBJ9zywJqaOhOH7ybyrTV9nej8KpQk0YVwB2BCL10+C0cm80Se
kU2H721EPUFiiW+NBmDakCl20Achi5oPDVQWj5fSF0gNRIdvtNlRCpZa/MtmkH8rVjbg4XDWfUVj
dBEoW4xA7j1yb8owlI7qodo5oea58SUylYWnu3AMZO60nyEtp1k+U/yDyk+kl20ztnwNpT4D+q3N
ed2AA7MW0QMmKsojLhcLfcSmJDcFwHJq3n3kUZ6K5ZOt59eQS8H9LJu2+hYsFNBgQBZkUbbDtE0z
DQzNWjrlmcC4sZrDZgQj0Rxb8u6/6M91uWf67qC4Qlzr6Ya8iLvfWj4oYZFUdxZ2Truy1wpjIfnV
nI8hkVFFf/0eeBOEZeVzJyWJu/rko+7gjr/kbTFrY2CnGnYtpNi1DHQlvhgM6TQ+sgBpHSu7ggYH
TmP83WIZVLLkaNntdcLb9hMKVEAvSXhdYjdYmcVFlO18vRrY5xZv71BYKvTerPJ//11dKuN/nveZ
X77iKKql9qy8Tp+lEF2Vmv9MWi9GqzLOwME9gCB+oOBRtx4BhdXYg1nsf5M6vLJj/aUFGqhTn8I6
vttFSEU1MjRSjuguoodqHOsTO1u6dLMAhM1kLc1iI54r3xVUZVboucTXDJr5YDokO8HlFnwLHylB
YdIi3idK35mnQmwG//N2UbVNJqwyIv34wjRjGBu+TQWKJzxY80F0UkoFb6FCBCoe+x2btNOqDXaN
CeDmKvqBoy6ry66B+LgLhSsOL815JyGynRMLzcAUG0pT5HYLt6cWzMIzZ11Pff4xcfH1tjBZr3V9
qxu/ly7FKtbx+ia9JTTUpCS+AcIrbkf+XWCFKpljguDafL1uYd/kpaiE8WjOs69uZofb8hEStS3X
mDHVgQW9S66xDsmBJYtjVnXoI9ANHVbUrq5JUxXqTfuRhC2InVDUkB61ORxeqfaSn4NUGd5yls3c
92I4SnntJ6Mp+yzs2lP+9UasatRnLpfJY8kRNbjN9XB71DpPEy9zJKHvjSAniM+dwV0ZLRGcY3dt
yGRSoy+x1/7G8NmaLzIqfSq+rh48Bv/Ju9+5FzmOe+WorZPVkt7jZPAEU6XQgXqo1oGkTjZ2vSkp
7UnQ1DuaTGHYJv/C3XIrjRIasxyQSIPJ1yjuweg4CMc/R/PLnPcloKjGJJvA5NJooDAedgDj874y
+5otl/fPjsZtdnYrZV8xkaA+U07MO8OWK7cSvbfTv3Ovw2PIWn7MP0sekB8AHRDcerYhkEJfdUlx
5jLaYS9Y2IOe3IDB3LsBRSGNt8Go+7o7jZwD18+VIjgzvk+xHYPROnDWl4CMkpbcfhi6qBqVsmcI
KIdD9HlCQgImGVZbF0GgtzPozWrcha8gVmuPlZFpl0PMdEx5nQmFu0u4wyIr5txBs67LdWmRl4Va
s0U5KhH5wggUOSyiDNzRIMUj9TCKXUx/OUixCfBp9SmM/bIVQ9D9JtzMcMtUti3EkTbEFlK7tkb8
diIEygxnzVT/VeamMk0m8eGAeTih0iT7ZGB+o/S2X9lQA2RqDA2RMZvXp2bLRWp7V5JDuwLw/uax
QLESAGduEA/LnYxfak1jMJ7JEPnRozze8N35LVL0OshXC85dFuOGo6Bv8BHipR/PQK7QhnZyoyHx
sNO4WgTpa4UarWp8Y/RPbwMxP9PCAToUWGPtX0MhFGv6keEzuoJzHXnsLxQqMED40yMjRU1YqYOS
obvXLZp0m2a1+TZYqafw3wdMRK7W96uOzNpDHSiI7AZ1MJ10uMKngjIEeE9jtGYwmTlFF3rppXue
yhSCDWOlVJJGoxRE1MZyHxtXLq8FH0ye3UCO/Okj187meRuTEYpgVTQfqmJQZ26UIAKj4v+27sg2
KSk/Fj2//5VStbzz39uIR/768by3E/m1tXeOaUzWmIHs/8b3SYpBsFAir5p4Gzn+QSDafc/5BA88
kMh1GiuWpd+5OtjD4MQjZb1TEo2OyiqSZi74njDjiGFhcae7nmkPhcKzo1/HNxbVuEiyL+vyKZPI
oifc40R6/IQIG3nFk6uSYvkKxOpUwpySRxnIldKciuIR+1kPAYvBjkOBZE/VHg4Qr92VqxZwpIgi
BZUAtRxfpPAhnUJLLJMUUcOzRES0ruaB3UECDUp8NNK1WYaCeUO04suFYYElXp3/3NfYgYoe9MKK
jNgpNpw6HXSrZzkk/i5aqd+Bz4F45sQuzvGGGLeFutLNtsaTBX+fEvqm/QmlCIiZAKMMnNT9eYtH
redjsFgwksQQcnimO28w/+olds9T0R3+8EaSk/7wK1ZCXH89x1cjPTY9eVb3TrUBSueFLuuzdEpi
eTAyG4f+/2mNtnZXVPNzacOcJXXabSZxcEaG/VJJH0Pz1yzcxYGdGOgjcXpKzvvddKdBTu4ZYiOT
GlO9yHLT4NIb6mmk00oUQRZp2wN9iYw7mJ0WFwnDW5PP8a/sf+X5dqEx6401kaXcUXf4vEigGlaX
6rALznVq5cAhikdbVhgU+uznaE73gxxAIZ3j/l1JE+XFdyQCBOECJN6VHDrhV6EP/3ixpd8Ax0wP
wMUWLyZTHyKyoiNQfnXou+qAEG30Y2NQ1akt/eOHk6gdTRY27gSq6zKAFRiHfFGqF4bUOfDkl/UD
ahjzgToZnEEw4+/b90H3or6mC+is+d2LsVJtWyvdZpdl/HbRN5SNbqOJDAwbzcWXlZKWwW+pYRBw
1IT1SH+gio/D+qB8p/mBg+uP6XHgPKJF9qfDqltE+r/a7TPxthulQ3G7RwR+FekesY4seRJiF6Tc
iANihts3D/B2QiG3uXCOfBjsQHJLw6jTUQwLAnMSBAjL+2zcF3PUQFfLUGrw/bSc4Fj1BjSBzAFT
yk8OqZzYm5q2Z0JZoBE1jpwYqu92YJ7mdEzmaP/H21RooPdutPysz7c2oLX3nWxFNULEhhmMVpnH
7iJN5/FYJ5Rb7Z65yB5OOxKHDsCfAe1UeNbapnA2YGT5WWbX38FMHUvIda+xaGYB2udVHoPTfbxQ
V0Dy68nhaEXjCALTYz7Rc97bHsXID+oJQRRA96IsT5fSrtqBKpaE7NA31BOz13ZF/ECyEr941kxz
1A8yWjXDQh3KHSr7XurWVVrWmYLZqRhqX4fCN4raKg8P5SWyTtTjsOhVnDBFLxKjk0SmwzdUVEuX
L5MIfnRpeGoxYEDi8eXCq5MSnHAb4gmiQcjUZqeKgkWb0VOoMenC0n5lmt55XwSKjxSkcETMv7My
1Q3a1AJPANqhiofJAmKdKfFwihFI0JAxzM4ETHcfJuTxeK2DPu0D6rnP374lQR7jw0WsmOs1K3h7
0v2hFq93xbgNao3r1euzDIJ4dabzgD1uZQI8KskbC5XtzqUSzTFC6q9ka3P+QidFtf8LxtQKX9CA
CHUFkomeaHWgr7oGSskXHsmOt769UoWelZMXRe+1Grz0q0qeIXlqd7vz3ocZajrVm6lVFWrfaCvT
Eh72RO9le92GL7qjsrViuW6oyJTRLOKgtek64kX5VsdRsXiMSPok57FKBfcqb8O9mUu4nc7ohk79
DytK6zJNJDvwcxABOTrxDo0xN1MYq78yozKtiyWaRRXcv1cH/0658Otoocb6tTTpJN2eU1siacMe
Mn7ong3YSG63+uENGvYmJ4aNAtMfAcApOO05PfNUGNL4yRfShoQfT5+ZQ/sbymhRzUkBaKgxyu06
2SzPSOw5SCjVHffSchgLJJNro/JeHq1G7Zv2O3d/S5YEahJBN6WHbuBHw/V3PgmpHI3TA4wAH0OX
uv3BpVZzJutALF23jKP69uV1MIo0OZzQwlpbyq/ZiKqSfcgRbU2a/IbXFppUJ5WwPotO+gLM2Ja3
AC/rPhKdgN4I4sStp4Zz6QDPDLzPNVRFiRPD9SRySPB4FXplWbUdcLL48D+K2v3AKfmhFSVfCgft
4AGFOFJRWNi/HHsmmQTkSUYqpkMlMlcOjQ4VUiQfez1yqy2N1Glm6xWm0jwbQn4svaHMmd9mrRrT
3bqeQLClaYuW9xOXqQZHFyop8SN9zFstTu978jE4KOG4VG+Z2YgH2Zg1fc7imn6RjUmK3yw7pENU
pGWIAZPN8+yJxaOlYqsv0ZLYMdOPuGM355I/SHXR+9XfVQzArXPgry1ig7s/bSrVgD0VLQNwJi7g
HmCyOrJRinKt6lf+gOqepP7vXzwROed4kUwaCTObchf/nP/XZC0Jta0oGkSYKVS1+anWk61im4Xh
jYEa722IwRZGXiF4DOJXODRFOnXPj7j1CD1wZiv2Z/qqSNnvKBSPajD6MEGSw8VuZoP3xiK8Nt/K
UDK4Ix67VqH4fzUn9Un89QPADT+DIPbuZWpH/U9vTkOX2JPobAULMOpqYTC2LbINkBJOcuo5cnHj
FIvuPsw6vEpsxO7WIAB2RgK8alwr6eJW99UoBZU/ATmTNh/7fyC3/WcbQiDNrDzAokLFjvkFuCJf
wZb15pmmduXWFyPxebN0d2VgJKMlpzTglD7Ubch8gmVyU28rW6ifO8NaEHDcgkxTkX9J3+ikLdeq
KdQGDV6SZ5AKfcaob8GTNE3yC+XLvwLHuzzCZDWH6ahB1d9zgb3jSn6KslDp98mtZhUz653BAsdE
EEyvRtwHEIwHaXbzpab6cYRRelus0wpj+kvUkDgpZobWrDAY6QvTO5iG0tupIaAa/ZlXL8c7ERco
c7z1tQSVGmU1gqv/hKW+NnxMutfn0sWIgPOlXqx0YVdej707nox6IDiIL/1Jp3Sq6RfdrdZeejYM
mXdLQBT5mD03XiMQ67dPFF2Ejrqo6fBu+OTokxVEtgLKORfAPxMYxSpxWQomP//GGCnxJ+rE+5gB
ElyyDdw8rD8rAUTqc542Q1JJrQDszvJjyrwvYWd4BAJ+AC4ztFiADSTBckM3m4xzjY84f7iro5Xx
AvarAUxxJSEazd4SzNjhl2BNumXpEIlBevo8wPTDVj2blY4ZqbWFsxav+W68PM1VkwD2dIjOum+r
WSDAzGN9jTe4BihZcRLUuzNzO8WsZyM8jaxce8UTC6cNeQvk2CcppnsuWGSgqTKBtfJiOi13VWRI
xSEF2MYWRrai7OIIK25T+JBNtBYYpEJ7KCKwZ6uALWcw2WDKCiWYht4ObLZqM1c3BEg08cjiVMzO
cvPMQALkPjfWXua8GxCEk4OC6awsJIhfY5Lewn168kCS+H+I0OS+HQQZDLFnQUyoeqtcpPu5rTMr
1EQ83LS5WLJk9U315szZ/NOaILgrKgBIdujrfBqa5vHDOgQSkuNwcPWudOoO3qI/TmYTJ90E5wCp
RwwQ4/CFJTRs8FNh/8SozGVDJuzvNFmUsLi2QCo4kbAyIHtwq0qhwLnMKlbIjNPei1keUF5afG80
ipW0B1TH4Ez/4Mkn9swZSfGoQgGSiGonDYAPjbzwtGns1IEH45EYpuaJTgJj94teZHeu3fZ4QjzQ
TDmlH1TrjTzsFQGxtqN2pdlboDir3do+qYxZ9wLYNPuFovsdIP8OG2TmjArfSVrxyGV54NJM1qFa
GvGETO9VPlz6omNN8aRww5A3PVK4r1ziGlpiM+gLFdSA7n9kEHD+tYt5RiEjqKs7GuMvuVLJH8Ka
SkYfjdW/7/H1X5cofpP0KI78EC9RKhRDv8evhciSPkUFIBv+zlBgSLMaoRTK1glD+PlLaXlHcKR9
Vv34HKU8LXt7fchwYZr7YTK0rfcq1PyNTrhhp432X1j3F6EQL4ucHd0y7mGuOWONnbJZFkF/5KJe
lSLd44vSlhupYI/Phvk30tsWEYfA+wtKp6ssk+fk8vHUDFb5t45o5AHO7s7z79snXT7RBcW1PKkf
gqSgcwhYFrgcDd7cVxfs347ElrWy6nVHlqdMQXlOBj11oaOKQFav0VJ+KHcT4TZojAG4jL5atzCO
qjcXEiiVhkM0BvuvHfKWRe2fXhzT5/QrJYcKJKfIo2Yj57tn39AMIG42m8GaGpED/f4TzqaS8ZGH
+qTMvXZJnH+N5d5c1ZIVemeH5OGhMSSxv0Ep13h5SSuv36iAn7A+DjXxeb0qUITcu1+/8qllA9wB
BrnjyGV9H2ZOyWJDGMx9+jcRUx4yMaCfrNbbo2s+DiURnmsqgs+YHILqClaJt+xgibMZORzFriTy
WnpHlYDVkz2C+XaNyQPUeRHbAdroz7JhR+P+Aoe4x1e0IeNZTH1niK41HSbAa4W48X9cZqyNkWcb
WnC0fN2OizS/G8obISGU1v5KuBAq9WMTlJiur7let2k+Ck2lDtuun2x59VZeiM3vXhE+nf36JMea
6AfHCoG0P05NuyR63PhhSBhiCw1d/PVM/PHHu9uCzWBLbbeXdKzVr/6yRtfFSYVrFHLI3tSpRaGA
98IcRTSFtK+UoKvdirrAJjqpTcLi8VxsBPA9au1VhBxWiy5lOLoaWm577dD1s8MZ2AxJ0Ycb5fUv
vIwYn6P9tRpgXJRS/riD5tWOb2zsDB1Cv5Dq1yuKv9xXGN8cIlWaMc6dQAVAcB/WXTc0PzllyWdQ
xT8xAAXHaZiEjUa//RUNfEr0PU6F8OXZBAa+dZGwQhntS04swc3R4u9JfubkVcdbik9D5ZErM1Ux
dg5YYtE9U3wZhQNP53au6iQ8I0L0C9/PKEmVyVZEoOBD5hQ9dGzFFbZrOkUFgJFd4BnmQ91olmVO
dqU/6vxPSilTeO38La25Ia4gNhIobMqP2mwvW4UwkxnnBFp4IcqMOAJSct+CQoxAoWBnPabp8IT1
mOIYJ6w9GJRjFpzGT0qMzXHzYI/biOeDOBetPEW13/4+3dNVKbsfgqwIUiXWxkVfki+HDt+mS0x1
yNsEHSLOscxu9QTH+3nhTgadlrG2WImxSknBEnVng4El11Af4cTv7LTO4BfPKPnjyaQye8ZJwQ5X
R8O8fcNtnWyIkdN8hLfA07MTJAEyMh8ihXJTpboWkDJNpNUkyBOpcA1tMMoc6HnYACh5HbwxSshy
vvm61nwQupCq1cA/al85uRYquryzJ86J1QLVVILDcPLdx53WpqR6LSyWWtIZF+8598ZecSDORkrK
LgWKunSgRv2qiIx/RilmiAj2w9jr30ZZTAvF5Xes3xZOtF3GuW9fyBlA7GDd4QeRiCGvkeHi8Juq
sbOq49CusiswFsAb4UCLaN/RhyZjf/0GasteXtpXry4jJIpJfnBZ9M4/BekPFvi6pbIziebRKEIg
wljNW6/cmSEJ8Fw7TkV02Rv3u/poi6xm58HdxPPgT+vyugwAJjxs9jNBwGNV98VB45ZVzVj79mb7
xJKZ2ctjrWm7PzSz3z9U8STvqhxHwNOkR1bJ6wsJY51B8pl6V9XvX3HOiNKGQ81C364mOeRtKwGg
PYsflczBLrv/zIXwIsKeFmkQqUReEqAAMjcDUQEgdrXzptwN44Srlc6y6G8mAaoynyLEHLLd3BG8
0CvzmQIiWj8uhJi/rsrQ5nNzNhb1hyuIFa9YlHJwSMVqp4fGQlwwUZCCGTt5r4me7GetlDTms0C6
ik9VALvIYhhp1mkOuTQ9vRV4YshGtVDzc0GgwbZzFOkhFoLBSAFXeCcAU5/WjlLJIn+fAJBPPkRK
cj16U/vdgCnfQlbvNoJF88wM4CUM0VI5J6xdDPrhX5/dth8C9GRtJ8Sq6RD1kBkqj/xpIG66dYIy
AFHgEr8ebOOj82vDYIyN6JvQuFLUsO7p23KCqeh57RXAC7PBINwemiLRm8C9uxKvw0Nu0VGIcZAw
mSduf4Dma4R6uzG7tDJsPg8gsPLpDMLydcjkGs/FONknEGkm2iGdTuze005Jor0Y1dQrtmchX38X
vxJdy2SFLemQptPipzM5mFZuZjel6NNsD3j5sOVyG6Eizogzm0zUBCwVGU6EbHoQBI6A04qBCE8l
FNY9obYHh2HowpQ0WLwOcu3fkCEr0uzMGIuEw960IzqWqDxKfnmgOSt24oWWzSGk63WjdZOA9YL8
juy0MoN4kN3NC+uSG8c3Bvger9CRhgsUDQVcnCVa+fUaYWQ3cc8hOvRKJxXwkx3tASAEuwfTfo3p
gqDn+lCR6SkCCcOWNzriKS06nTzY6guS3yLf3OSObIcVQE08uFABfh65I+nfOpcYU0bVIAHiSH35
psRC21/hjxj8+3bO8ZeZhDKvTV2uPfjaITvz9RUIlBRmKuSoG5MdHeUm0TBoNLNZeGgia+d/Mssu
mYtm6zVPBTP+XOXTiFdgXpVqc3ntNBdyGHByJkmvAjYoJKfCt5KWfEo6KokszEVcNO4wAkjho4mc
L72eI7h7fkXmxxt136kurggEVa2jYW3+z8qPMEPiB2HZ8Oj7KSNlrds1vmDnb0UIx/0KbAEmiDCV
gBJIax4rMK6DAFm81kfLiJXKlILmo9zBWgOe3qRmlvg+ZjNMy9S5FxJT+514ul4Gq/GHszoFldMh
CHs21KwJC0BE2Mutiycn61O+0VYGyNXGH2yYnckeyszn+v+J2tWB0OkqnuQ3/vUa+XrunbTNv+lo
sn3vqpCSUYQmYUQPVHZR/tUYgc1y9Hczqwq2Qmb0uM4Dypw+BI8kmHNDQESMS1QXigKbsNbE0yMh
xLn9RHCrOsmYnzIBGuaJB1sChvTGE97n4aDwhHkzkZh7vQUmKF9YPmbnvgZVke7dK7IVwN+lUY7y
+S0CoyH/ZkjWoUlOAQeziSa+FXNJYSXU1YydawD5WSO8k/9AswRbv8/oYIM4G/zj2YNxm/uYKcRX
RRrLSdG94bfFZxceZiupagpypg1rEZKKcjivMLN5WYKBZ2I8LhLj3YLcUysty8iYga0o5pyW48ek
ULtD4c4mcsiVoNFWPuZ7XqHubLqDvv9qS08FZPXVHsLkPeRgOssGa5Ms6Ac3rQkqdRnlOSNJr9ad
Gy9QWBI3v6+hvyM0DUZKZm0j2PUjh5UH/ou6+JBOKMf4oSOtMSYkxU9m9vhid7MQ4FxnXjPJIEq5
GD4o1XfyScfWyoZ5vDXJmvBdbTYhw3jSoQidTF3bc/BDnl0ShYFLEv1fHCet9CvzUKTjxLypsi2a
rtxv6f/TkFI/sx7iNqqNtnGpIbI0IOv5cI6F8UEnssvROXf86y5J1KEWVdeqDs8O+57TBHBus1pq
9hXD5adDyc2O4HTpfV0cuwK2mhozPafjQJOQcUNZ6Vu8SwSmaSUvcWSlQFiIcf4yY/nQfcZPrmYK
5UBMDMbEsu6xgEjaAwovC/BSDquSODLHh9mp8cpJhIkCmxbOx7VLWMF8SfmQtR4WCNMzM1MdOps5
CmS4OPlomD4KAA12CY6L+LhfSduptomLri9svx+NdPpKUkdPXHFqX4kHsf6CxXRS2ztJ/LWLLU4U
oDidJn4y6KCGPU7guHopenZm5UL2V56Iww16ZSlJfjIDrNih7iok6z7vd2tADFwwjwkqDSL752Ef
I4u+IrQ3Xys0uL9J2C1i7vbVNbz+aBolhBaeSovEWskJAS7zj8yuaggi7hPsus3UjVkAipZBbHq5
VyAZ2JDAc0vOg/2VHvta7+8rJXfK2ZHM5fy4OXaz6ga0W88QG1S9i/D1ji2cLzg9Gi90Znsn4dXo
tBb5fcA1SaPy1FHkBk+vJafqwfLGNWzd5ow5xX3Mr5vc9ocVgtONUUcQz65fCUkFBYB1W0ZvVST9
psPnOKkR/CEQomjpv5CxNVYIjfiLJ6CsxRuM53GbXKjqmRxLpII+abquO0fzZ4U7FP7gNw+kgxv2
9WZDanO6IhFSQiU+iKFS9RMvh7m7PYOlpP7O6nM62aiUOt/9L1HE7QYnTtvW0s9GR4DJE5gdEHHI
MCxUpFGzPOUhBLigBHMkPB6J3Sq7MomxHDUWLLvFnFoIksZcS34Jip1PuAOCXUToYUPUMMmImwFd
k62J6+RXhrpG1J6AcEU+kQ5DGTYBhSyiV8LhPFNNcJTBF6+lG/2p5FHX+FVtb+AAN+5Z9483QeS+
Zbe+pGwpf//n1Bn4iJpUqV7LrzC5aBkpHJmYBnbtGvN1RMPnUj1VUydNO87BUtrcQ+V09KXCVWCZ
b14qmaz8N1ej4p5I9RLLqGkx+utyuklz6cbO+do77MSzP++IYWvGp313RLrnG09Q2FKL/fhDs/eV
ycchzTUUCpkU6HbIpjRH460GHasGPofuklDuGVUAkYxQvLWaFGXKY2RkbChxJ7hidJkaIg4d6sOK
KbGn7ICiA51Tc5fUT/YnhbNJ9LzsYyWXsDvJxPx7BTJvOswmJjnx5wVOJw2rhTe527STBMxY37b7
T9ElfhZ5skamrQkbAp6csLNxYns3N5OJNijmPWAmRL9eQxyj8+qHdu6FgHuhXhGbpmDeskeCoDO0
spf+OkaOGLeNai5Bq6uLPPZDZuGsEvY5zV7ft+gjUAqkd7CYUCJCU7tgneKp3/QNOvfNLr3atI7f
L1YTpsvFRcSlsH8pmYc1pbjfM7gBU8ZWjMvtduVK8sKlUkYUkeXY3eiJiqhoefdybtBiAa5A+rJY
obWh5F7F8UUF2M3Aq5qrtHd/zR1TPSXUEeYA8ZWB41hNXQEpMyL1/9+WpP+B/FDeaAtEdNV0WB1v
Ur8s7lVNVymYObLR9iEHj6f+cbzWmLCreul4ixNrNJvmylIp9vVCM/TzPsTc7OKsZh+qibfOHnLo
xZ0ZhogVU4q9CnZWQftKwUHILApNzp+utlcD1Ss7u0QxKNcxYP5CQ6jOkgfZpuMSIPG6EdmaaFZE
s4nhB5I3oC+7PmG3qG4rY9lBcbaklsMbtxJMUhO0Mwvt0ijMdbMRxsoMNhHe9m35nBZXPl8ctw4T
AqnRyGHgEuJMU60XZvyxKgtbXmOT5Nj7P8DVBmF1JsZqwKKvsTY6Lo0TChUVOy5RQ9zz2TeIxvQd
1Q06d1mQxoojNDn0om97EJRlY93vxoklQVrkz2+3DzlDd/uN9WDiDwnDxVXgesEPfhOAFkNdIMOS
i0HK0PK6/55jxmUpFUpXvStNQMbesIf5bpmPog3EI6VIbc2stpBxktca7YgnUc1W/eIqCMtoPnXS
qsl+xKGevf4TnHJP7ayaE1/MmznKsP0tsc2YP4A92Nu5fAdTMRfOSvd6jMMfdD7B6RrpXemdlOLE
3sSPlJW5/Dzh8KX6RJP1aA4g2IgTOz/4BFFNLf26pvX94+ViQzWxyy14cmNZSxG+1wQEWFsUanU/
ZaaLxIkIKrBVqFqwBsFZz0C9/2RO6Db1RcdZDUe7zfimbFOlwrBrUmxAa56x7tn61P9ebsLO4yBp
nBVbNCiDRISzaOjnxZgHqkIlfFoFNKgGrgAZifI14CXVSE8AcRkhGyen0PLG95GUdtMxBC1A8uOm
nj/+HANa+UK3Wv90nVxPls6Gm8PY61i2NvW7qFt7DeKujqJc/5fRhkicI9nyMvQ07AuTBb7oJNZW
IFhlvICuQbvjd6f3Goy5A2E4T7GppRtUP6pHAx1MboO2v9xawIqXhX0FrJxyUzgrdUBiCjFnQT0P
Xf9FQb8x2EzTmhPGkpYfTy8Q8rgo9n5gj9sNWgpy7wqwUIGY2D52EMQIducp5CoQWzUIzaSdOYaQ
l4YwqoOztY8VQ0jzN2/WO/n6nQcWxFB/ea5rNZdrc4aUeYEDZEHAeOnUfx4PlBDrTPfr3D4qVLVl
2kdE399t3e9qaZrA/ASTkez+UPK8NdTdeBuCibNFYndO3hYwVPWEv4vShdFntkw0faPr84fsgKwm
jGAPZkkDTVf20tCMah5O0jTIRqE+4iifjwD8UuC80bXCFnRitmfCmOveDB24Bl8thhS6sJbEtyZY
QqceyYwzhOOKADkG9MDCVLdlSejiTdrcezsm3lCAnoUvTod4j69s0lfdwA2MQt8y/wmudH9l86Tf
ptlr6y18fnDYSg6qCkSMfRojtCfMn0u+vHRP/fb0XPUnPpAYPUoonaEv6sBj4td0TIr0hWorq8Pc
tZDilmyTZwZ9tdCAndXjFjuxVk2OgIka0hdUZAr0mwda0sze6mHtPUBnaP1kLYtCWPcBMf2VmU6O
1O/7xVCQxd3aVk9dPwngbVDckvY/eGks6jq8rGxMUqNJYEJjoSXc6vF9117rIShIUoCXOLAoyhrQ
4kXoftKawuQ/YYR6Nb8GA2jJWaEMqX48I57c1IVHMI64H8Cb1bpIov/maD9dtlrsDr58J7/vTNqG
IqMdhuyXohZZgdrL2i9rKx7DlHfycSZuCVhqNuuWauxsxKtrj5+DGlMyWydN7OuY7GoHpNqkOmjK
uw2CmdT3drkZfk2SmiZyy2nK6ENNqwuTp7IXkIO/45rnB7snJiR6FI7q6Kr8Mn7qkwheHIpl+QAQ
hDdqffjXdZGgd45zsZ8jFbrmGYNNvezpR9ZpHoyBtNxmjgzgfaQLu2ny83aqV1pj7GBy0ZXNsddj
i48WJH1k9dRG8bkI6i6nn3Ex1tgDD7HH1+WRtUWLf/ImavIQirqKx6bunnvoOYLvVvkcYZikiYTz
HR4huGPMnwbGwwEj6FuexCqPP1X6BSj1QNZbUCQw7r3RTHe7GLcxBisYQgyfXD/C2o5a1YrLtzAQ
XRVnYbbaDhlHVF1P5LyX0pOiRF1Qhvg0TAWfqCO6kE5GPwlj3ARC2PqJR5/v4pFrQ907BSbcixbK
v8BNOVdFgWazRpAcpu7bjmqJCuoU8TUFygMJjdHLM60eIDP07qZXKT1udjIYldoGsag9Gv1XvKNd
aUwM/zI8MoR7GDdJHFf6tO/Zk6WbgoDCal5MVBgzzo1kjX8I5JA1d7mVIOUM6+CkIM2dZO9C2zb3
OqZPpI+x1V+RanhHPHbBhauB1omGq2SEfkx5bJ2PbEUQht7P7pU/pQKDPn9IWm3pCDeQw7ci4388
eBVhznL0kvDnuRKjBsHtcSNwH+/1SMtO11fLdn3DWpv5PrkkDqseEV81C01wLoSPjI9/pP/oQhO5
Nwi7Y9b5VLD0YlxZUaprUPsTnM+tRSu+bKD/ZbHh8Exh//8sfM8oVHxnivT/VXgXPzMesLxK6nsM
NcX5oIh2RyjoEWxm4F6geA13WGvnlrH66dSGHDvpYzNHnBCfrF6if5ADUxyaPjNHlLKg5hZrke52
3hXkJLSRIty6bS2MqdIDlr5Nz3N5TpgFhzF38sY2+agREnHLH6dkg+PEwPZ6DuNXeAqHUZk04szx
iGGlhKXjeENmFNHc6Z6xA+aECuMQj0+SMM8LPY3hisq7fi360EyAI5YjCFypY2BT6A/saWMjonu9
Kq6ti4pXiU2V7Wg3+x6+WBAxkbueB4FVklrPeIYAM4gDEmmPz1YkC5EtImVQlU4uZyODH3fhA1EE
qCz9eKWGN62317elGgHCEr53CvI8uSdOFc4lC2OVfgV4u7XjIeiqhS1+HtdJxOaNL22KkCPv8g/t
nTGcCF7sOJGb+0ZEkzHJjJiPhGVMUMrFnmh4LldYlHg9TIGySoYd1h1oFNNtmxKfHdBGjnbEiJDb
8guLRmD+HVO+CfFP0ighwJWNUf413wYZtDetqrylUlD6B5AxGHtgFBvCEdxr5uOaBoS9Zl9IM+RG
uaGkyfJ+mku3Ayft2/uOAqTxN32vfsawIj8zIpdCn6UFsjktx3srJ8uzk2kGwn7ESTV9BZQ/CL7R
7wFtZIGVd7Pc7x7fN7gpYacJfyYFhpunXkRzbHYaLxYqnuQUANoZuPvdP0RMtgcwtIZAa8jr2/Sj
2bT/4NlWHH8om4Bmttx24Dm5/gom81x74L/BalxWoz1haKtYC7zVhLvTshFY3bxL8qy82zmX2Zb7
lKiUucBSwJvbMzkIWQuOBAY35Sgp+6lIg1V20YApLol2KROGEM1aGuMQjOqkFzNRncYnkVKDNukO
maY1va/3EpFdDo1fg6PPCT4Cq5+r1vaQ86E667XH/yeAAJ/mt9LCW0TVxO59+Gte0YLvCQTrQWsR
F4byH4brQH/1MTe96p1eLpMYM7yGdlSD4wThRQ8IfuIw7uhHzdBGnvQef93hR3dEX/Pmp0WjQY94
s6tz6Ri+Jf+4eHF64/fHDNnElrW7BEqi5mUXywYJV2iwxSfOmqjk/pkjISCarpv3CBMczt96S3v2
jjM9ZrPfc9OrhVoUC1E7WoseMC+Gr0lCfvbYgs8x/TDjVWcC6gsC5NALO4TJ7M+CCF1LEe2J+tCX
F+0d/AYmvoTbsfKa+CDNLRxFKjTl6e84tnygP0XI+9GmIa8cNCPTdCgfHQkvud0S1nA+paRqntyp
r2a0mad5V/jdWMuRzInSUiwC3Bho1hCJ55CjOGdheAHxurE0t5Ap3Y0hkE2lO/WMrtrnfrR9iNIj
r2wC3LRR5oXpsP9+1I6snd85YfOJtSGo45v4KixgwPd71jV5pEBF38rT0qcyh7oOFy4mJhbvzAlZ
DdDd/8/u4koTO9Anq2TSZzPtm3197qwjqCaO3tf8ejoh77JGv35tIGDmWbBEOTlAqNyvzY/u5IE5
Fm4H3SCfT7E7zRX0VetpzHq5Snu2kpBhr0rysQ+HNQKmgtfP+9L500H3I1SvhhuKZWR323IeMxPO
mK5NhIoVWrL1wQJqj+OG6p8lO4uLWVQQoWXn7owHzH7s5U4PYjehb7XowdsJkHQU1vYr3kXLyvqa
2D8BeIiZok9z0cbsg6zvAHq1ODADXkGgFMyb9dOmBth0mlOcODw9GZjPuTyQqrOHeI2hEBJmOL2q
AYKXZSb491uTXB7K9EvdDCxbqVMgJIXp0yS47qar4RCbigExezjn9UhToum1qlRPLV3mMigLKcji
hZXE9hF6pV7KsZ6NrXbQkkEpqF9UYAAItO+uPRJW9C+GyQYTE/zLaDq/HUJqL4VLBnCDvat6RMWm
aPxCqqZG6bGKClWg2ai7fJLHECLsbC94lL6qCRnjMhBxwU42E2vK0DceGDnNgg1bNjaxRsvMWsog
hdDYN0TQclTXSsYPw9nu8fCIlOQaJGE5AYoJtjoccbBUK1NqSb2vBZFM+64NeoZ4wbF56zjCHRCW
TN/b8RykS1HOuJ3nmU8XvbHczNQzeSnH/gkvbi+WI4TeZT0MAwfPYlm/HMrT2VgYr4cGEh5i7P57
pKfKPmtBb1vSnA3+9pNusTNCTAdTZ76u9MZ2+mmbvguT7MBQPwJnP0UoDQHy3hFhX0Eok0unMbFU
sRkIJ663bEK+r2UsNncLEzEWMP6StxDy+FLmFeD3S4IZ1d7oDnB/Dqhzr79Ay0xWWqmPUcsAVs2I
zF1rk9iLxDyYYdRaJP+AKlYII2C+vQzF4JaZWf4GVXk3vK3MoxcOIJiuEYuOjNudFxSEmOllyTCq
DD5eTPdTfWRdSoIo9ryxld8w4HbohtwJKZM8rhpK22x1hwERZoDkKXvkZ1Dbq8p0taEKKUF3WTc1
5ZepoDKnwxKFD4dVEiB2E6bbBzCeSXyy1kI488e6RDSteA5D7CohJVobj1ovk2ZrrgSgyfakxXYE
tvJfJ9CyH9TQh4aSGdU6IXGZtQvG8zKp6r9CMgOXuNxho8MJEyVqzC/LcthhUclE5NcEteAOyY6l
Nvc6Yp26ry0nMor5DRhIsICLAjL85zmwMF4UaDsRIhODMZr4XWSL53FZWJxaJ44RI25491gWuZVX
ei6iy92Kq0k5vWHKBno+vXa+RW2CS5Ougb0xlpsJ8HA9N9A6CiZAYLqnUBg9fcXljhAOhDHN8h2H
c+5rdyzzEpFHKFMwHHcNqwYZG/3+2+XamY5zP6hLx2Ph1nyE/bpyIj7y0C2l1g0CyYxuDpJ0eUdX
xcqzTY/9B5kUiCeU62iqFT5SXmbzhh2mItEkTZyn7aEL6xGemLkv4FEiS3UWEOeGHieQDmgIUPj4
vMkamZLhF3OOw8rtff68ZFbfPkujmSmaXllrWeJisCv9Pb2Tslp7pFfA5hZ3q3Pwb9fjq1nGSzaa
D03ILDiXmRZW2oAPqoIjxAf0i3jkVD5NouHdEZ0CN+M4u+D/gvYxGqRa725l/d0i2KLLRmJm9Fdb
72gAwbAJTfkkAvGPw0QDQim3Z3d0J+/8bvaclbDxs1tHve49p6RTIm/brJWwgvYPdu+XPCKDYzQV
OUsVdfSWSepGy5tSuq753uWDh9MpjzNpP0CwT6U9pw5pcFKf6K7YMvee8XC78+RFnORq1cNuj2st
7VaICdeKFaPNqfQVmSClohK3/gxPjMHrEZHpas5iudZtk+opG484YS7IyUmSZM3g68mG0Up+oY8S
niVT01KzuzPy7SmA2qdlLA5CkAXn12sEMf89VQMUCJXmrHc5ikddwgX4Leff3GU69HOPmXCgIigi
vGdegesLbGAKllq9R3wj3ShY3fblTQwc/hCfDj+ZbDp9nDdBqagnYNpwY+lhrRzrMPttsLf4xxn+
VSsCopMKoLoiNsc9uZmxZNwgGnOBa8/qegGmp7b4lf6J/wB/WThfeTdBUPJ3giAgf6WjiY8aRP4+
kAHxqHr+EBge+PrXF2nJB8zXFT2kUpg3KIF05X2/m5H15arnlxOYwxqMRaYMxMEauFpiLEP0xqAd
x+/1q2/Bby6EAvQAUUzyf2p4Gz0SUQLb8ORWqRVKzXLhKZYiDwpKRgl+s0eacEjItQQ/sroF3czJ
sprZe7NWmSWVyvMYKlgFcGBybHOAV9/qR4g6SR7tpIfFGXj99aC1ZIRLb9MGJ1kZG7Y1l07FF0+5
1YaZwa05w16Uv7ia38bjTbJvOLlQxI/SpnXv8ntWwDtiW7+QQ0PvR9h0EdtMz6lhfk2syVch4u8B
v3DgMd+4Y6ped3UP2z2l+D314mNYiG9nX+LydUAIfN+2Tq5cHLBtjOAIXVf3EfMq0+QNYEg/K3wH
ewLm8OZW0uq8KfnZ+SGRQcRfeQXfHnsolqfDgo7pnoN1zdeENywSZOmosXB4oxMz6iAY6XMwkyW5
v44liucYCBeKLbQGh6mMzd6jIxGy17//IPnUAApmJt6jh0G2PXCx2NY3IBbskFlTFD7+4bmMkFCS
iJpf5qmo4Qma5yEhU9j7wgB1gETVxZ0SYDr+7Cekk79/t5sR4IK0yhD0D3aE4USaoaCdZ4Qw6IOH
qaMfuDTLSAK6iem2XA6GWQRl1rgdPDOMoKskNlaVgtFt/fvdK8gzGG3MgQmIsmUN8uEEEAGMJ5AF
+XrsNrO2idQRNu6lF2nJnxYF/DStjebwmYeHDhIv5XZQMBkD4EOX/POFtwVwVAjm5YEojd2Kn6cx
9/ZBDy6/iFTGH4lZlJYsAK4sM5i4BWXg5haGxLIWJNQ59DkphxndkWZIDX6QoYrAKDv0l4pvA51M
ZOAg0sqOV4MXqqejO4MaLO7ijR+zrwO7LPnye8GKDRrPdD33MLclpt7EIhyg7/PP4gg4pWADBzJB
bhxqChD+XUXhFh0c9E6UOahCo7LClqLtHklgWKzQw6MzTvKcC+QTey1DRnCvdgXv/cLBj2PsIQ+R
PlIGwtvxditgan/ZDbnaRSnelWispt20kD4OzLbgB4ETQ8/pflQoLjauzgz9SlSpWwDGiW/gFOxE
E4lkCJflAFhrMR/NpFLstlaKD5aH4m3wHKOoW2UXegkVFdf2seME+yvBNTF/BywrLrTfY8cR36Fg
P1SDXAU8sqEHIsdBKQ0VXL6uZp8x5qV9TK1Ni+f5Qv2cc8p4sQDhgZBG+Ts7HoLfWPxeydzlisel
qpl1mAnHMLOh+jocq8Zw89GqIIMy3AaA3cyKcf/WuDkxWt7QB/4BBnl9xd6pZ3q5FWnQvZPQjb9G
7icCG7Dhnb+1blGlSaYBMpCGpgr9PQNx4MonzTZJUT0aOfRvUsbVE2r6A+VOZMcvT0Np7bplol2w
EkS+Aqf0slHqpJGU/kcbQj5heqocFgfcbPJU+6Yy7fsm0Qo1+nmrug6gZKL646V224JobFZ9SmwJ
Iwrq7O+D9jIOHfordrDp1eJmrt0B/50glaTJDdwNAPmv8QyG3MLjoeY+xEMLpnV0ChBrRJago+UC
FIPPw1YvDoXRQ9UutOXsfYF1ovRqiplF1Ryi2r9OhVuRbXxqnIdHueh8593kWlj5fPTTw21xT0Bn
1vgS+YV90Pp0H1S+EWDOD69L59GYdQo0Qzt2CfbYsSbgy42TSJEUHeNFxhLWmiHxe7Z6z+KU0mF6
FV+Qc2nVUaXKAFPTNA0Qf4qq6FHRsjPq
`protect end_protected
