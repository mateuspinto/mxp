XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"���>��I�������+XE��e�ý_�]#�4���a�J�>|f�#��L�C�?�|�v��7���OV�lF��
|c.Kn$d����l�+�j���E򍳴ݦ8f������*z�tL{��f�{�����&
�b��:�%&_ ��e���;�o�Y���*�Ӿ�7����eV4�˅������{ڷǽ�0�i��.���Fg�A���ߒ�y�I�L?���%#�f&ƹ�v���=W�|������ć_����/G�=w���Va�����c�������rJ��`9�a<���l��u��IGw4ۂ��"�/>U��2,�I��L���M�U߱���i��a/�9D��Kw]�41�� y�1�<�4���l$^�#/� ��mPx���_nr�#�����ė�HZ/����� \,��q&�B�c_�z�;���'���H6�c�� ���2��<*�ʡ|���b^(��g���_�H	l�#�I�_d$!�DfDm��gld�?&�@|�3�S�����$��8�S��������K� ƶuiH���L͗��."N���I�f7���q�$�y�n�[�²����k������_���,�<+A/u#��׻/y�%ä�i�g[���rǰ�2h���0U{<�Ϲn��!�7��5���pb]�jq��<Vs�4>8���<4\zЗ�=�6UP+Όyi�|�gN��`5����
�}�蕵�W�{&�Mɖ*,+-V�2L|XlxVHYEB     400     1b0D!�����6�80i��>w�l��eo9�
�1c�r���V�[��῅e�}���˃%:��6�3~6y�s�q���+�����P±
�
���E�N���Jb��j�<�iz�(��gI��''�{/Ӆk[�ӖL2-��'��X�N���X�Z�*����(��X��KR�Ht�(Q<Gע���]��^S6����Xi!�y<NV�(_7�����mu���&�46Da@��Ch�a��TFj::E�L�������ߗ>w?=#$e���ߡ����i�J%��ߝ��)��Q�:��=-蕠���O$��M�o�'��{�����$���v�������L~�`��hg@T��`��DfA�%ٲ_A.A���n�jPÚ��p�7��o�u����NU�63E���Uv�lvG�>,���������qXlxVHYEB     400     130��/�SpD�PRP�,�ȍܶ8�>J���Pz �m��V��f|��t=S6�G���ݣ��c!位��Xi��oO���=��E�yoJ��\���
,�A�?,�wf&�����k���u�*u�A�ҷ2��MM؉��lsE<D�M�1�@���� ݕ������n�t�}L� M�_��Ԟ�U��/\��s��ly�ә4v���kJ�\����t��훞���ݾ��l�Pr��o�UD�)�`r�����+ҮSےdE��#�=$�9�/*(�F���#���X����7Aa�Bn� �@�PM��XlxVHYEB     400     120:�Pϙn���2������e'�d�CL�L&�6��I��}n\����ށ\�������ۘ��u�����1FH@�X'��ۑfųk�n.蝵Jy9&1�Z�RȪ�M�ˋq9��_��/@Fޔ��h�gO�fTV�r�x�� �r)��Y�A�=뱔윶�n5��Nq�iہ�@�׳\��lU�~�6YɢF�l�fhe��8�n��upc	U���o��l��P��Vý�b��/�o0p�--����M�a{5�-���Rݴ�XJ���0[��`��S�ZzV#��D�XlxVHYEB     400     170�R��Uc�2���5����br/[�i�����xR��N�7��+R�c���2�=4�G��,(�r����7�8�dw��.����&�dj(N�-vG7��5HCeI�E�8+C�����Z8�xQ/���`�2	j�����E�_���pN� hm�ƊX,gR���wTK+�j~N�Z���Hd6��V6xWOzT��'0���S)b��*r�y��G�gO��F>w��"�6���;!�� �W�^=���rZ#��a?�he��Ϯ ,�X,�{���]�7a	JF���ʚ�J��m�|��WrMfOI���N�k���I�5Kw���n���baz}'�*��)�٠F�ÚT���]��K��XlxVHYEB     400     1c0B�� .*B�N�������c8l��3�L�k��G--
̥��
ISޔ�v�(��$_x�،����{���g�`Fo�t����z3@��_8w��!�����YN��y��}�%�V���7�]7V����_�X ��-{45�\��F%�,z	+���VpOHԆ���t�}��E�{��$ c�E���F��׳�U��� ��Ȼ�WZuNA����Pb(�ܰ�R���ǭ� "�������I�U� kn��K Jun��$���{7RU�N��j��*̐�g=�BR��oeԶ�P�ߑB�*#1���Ck۞��a��U�lgB�;��W���ݲ��d����U"�em�)j�m��ۏ$����%�g���x8���f�t�L�#�u�����T�Q�����m�n�ū:�j�y,�E��3G���VϧS���qQ�����4XlxVHYEB     400     170aZ;����Yf*�ț�u<Һ���䴚��D�*����@�,e�Ϭox1&s�N����H7i���_Gdb	�#��Oa��-�tg�qY/�{.�?+�͖B��:I���Ժ���Ӽ��ąSU�]#�K"'a��ё�p'ʻv�G�<�M3�.Q��	�
0\N)EĚ�d��17�^����V�W;�_�Z�<���|*�+M0������c%Z�'��ʗ����>�V�bf��t���/�W��JO_��X�����4x�8��=�3���!� ��T�����ӳ4@b��3c��x�"���9b:I�3=�\�=qg�
�<6.�7��@V�߅W毪�����y w`�}]���*l�񱬭XlxVHYEB      5a      500�n@����I!/��:�+k�l��d?oi�6ˠ��	�~�њ�����V��S�v8zmVàbAXz�u���o�Z\;