`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
puFGolSwSoWBCpkLvcuiF8NCdbZuY6hZ6XglmYWNuWOJdMmC+cXBYgFdiTQhLNpxUMiqKM7NNEuO
r83EWUZNd8tG2kj9FZeSnWLBlX6PJivadEE+UDkark6EU49hhGoeOVJoFc8feVmGvgankFpOaQo8
tt8CXbCnsmCX3LMDsCw3nKpVRhqjVtWTJ6WaIqxcypNprav7SRXhhlYfg3uqJgkncbez2cGaWdWM
cfWyErgaDOYUiuu2rzfDx5xmsSJ7CXccGq7KmM9Z4BUqPFRfzASEWDOjY9QdgjAHNifWeBH+d5WJ
Uj26WLglCoWLBYFD70/m5qTw0PVseJLbd8aomzQtEo9UwhLqF1DjGXfcad5C76qRbpc0q1dzfVNC
cGF9sfBzgx0HZi/ZiC5A9uF+hzlvJEhCl/XZqS5Anem2uhwcd6F7y67cIlj/2FaTNZ5v4xCIdFBW
F3MFJrAw/azJyG2Sa/5yFGSDdOd7WUstLKLZDK68dppuC7lYi2Wx/dfcuHQpIZ3oyZSZY9vY1OLC
BIU1BYHofSX6VPv5kkoi41pXW/vdOUATepit25ucNSJ+d2EeWedtCV6IS24YuzVb8m67xIqw7gEI
Ev2e7P0iMHRTtc5yCmgtdtOOVaEoRmqr5ZpxfLLbHOZFMFUCV+LEGKcC1JEdwg8J0R3nZsLFHDKN
aUfhJJMmuTpXLDbKyPaxiCZIB4mcYS8HctiUXYZ4dsKSlt5t38fPNSE2FyLrMewIj1xZO+D/EjUL
6T12IXJxec/50I7aEgcmQ3NFU48Bm2qBlIb4TJVXkO12kGN8smRGLhD3xYzvjHPDj4lNyJQhVJAY
UTDSBTXQLjmfp3/l4bRhjLMxHGN8BynF030hdIlBfWNXdSNqlKc7xOu7dL7/o6T65R2nU24Jqmw2
O5hj5w52pWtB0fXOGeqtkUYA429hRJAhkawTTsMP7Cu3YxPxWS/2cmKAP+2gMShxh0DPBuYyh5Pt
VkARD4PYwCDgjG1WxbUEWt9naoJ/9vRarjp15HuVrv7H4uysVYamAkXF2sweSwQ/WIlhv03mn4DI
Jq8hchBSOOAo7Ir30IBjAI+wjlvibuOLQUQnJaifGoHTIdZdRDLQf6dKF2uKcLpgD+dutMUVOnfN
cgkj+un3DgMnpHncaEuqyHItnaCTWRHiRQv2XfCbkU/mKM4L2ja9gntCcgJdR98KVn0H53TgMCtF
6wSKWT1bPKcEZVrsvSOfiXuo99qSdJLPMLlduQm+4N3sn2dvrhORpHJ4n+048DC9W8XIHrW7ci0U
/n+G6ckB/lnAq5YP6Ac01UOmA/bxhAiU20Jp7mUvMkmUBHMTaxI3AM55B3oUKgJbEeoO0GW9xjbe
U/W87Rl4Z/LfRVXFcx8M1VwNbEEVk32CGBTo61i3GozIqXH84Oo3DD+/dS3DzrHDGDgMF1JdNG47
fJJ6Vw0iD/7DvKmTllOI81w2woWzP7C2oJ1r88OZN3gAhw8yKkB0pGhfEHM5vu0lHvFLTTOynBBf
4eo3QK3CtcBwUIWageOuE0WL5iMQ3y7fchplj1aZARZLSoKjF06RGF4vuoEne2FfwQom++iJj8Mb
+P3hVSTrDShnDqDCbCVd+vZewmYSzwh2U8I+owtKXmMDBjRA8LbmZ1aGju3nzt6mQuOlo5UiuvMM
2cXx9uZEx14gzylx5X20RyZSAAp+9qCn1nhepg1hZtfFJsrUwP8LR1URuNYWvmWXw22ho/mH21vq
26WIcHOU564w5qxCilJzGxmxT0EgCh1VNAJvu+H0zFHYMQOakcozQu+tzhhTlI8Bvg1U8PtpsQq9
ZRGCAHD2svmbcGaM+2SwaNw17r+48iB4Ipt7T1ctnpQsfXaMWH13kskf/hr0phvZ3MGtDr6lGKH9
Glw28ePtPtXXM3l1NwY3RKny0OjvHcejCofDPN8yccnEWl6pN4NiuH8sV+sQFLsh1IcJnCpgen0f
VGVyw5wcw2+E+qmxMmVF+w1jOp/lvKCckqbVF3qyFmni/2thC4+PgpFFz5Sz3fZ04GEByFOVkTSt
P+nrevDlS5XIcSQnE91ZjDnDeySdURKrytC6sncPNeS7nOWvwh0OHQviaF9YSlO8oeFMh0+8jpWG
B2YalEyPybB36Ch01iKvghtWQ490ILdEQDAvLfOvdgvGOQ5UlJBVorKWLnmNvED8bCnvC6pDBFHz
cZ5RAGgA/C+POGCkU2FJA5uQaVNxagcO1l3eh/HN+hHxMhuxi3jMgCQvsieWUM2r/k4uSammmMxA
Tz3G6vefLj9FizqTzGHRMDPGXvIuidT2yFvDZ3xQrg2j+6qjoHxv4uWXB+w5SUkol42krRnI1qGB
Bz7RM+sFv+1lr6ZwIS2fr/G1sNPn2BjEfu+HDNRZlWXTq6xkHTv/a2C203QfEP1TG6ejY+lKIA29
hoQzxjaIETGNftS8R1O2ul9MQfCJE5rGxkMkH8UMogorowkAP9/4MqbPMAbqDlM4J/luwiQ9rajW
5eDNCPV+iISBnkWnFueYpvdhDmU2j3n65MkOYJtdOoMPvenOwo1q6nRVCV265V9yIXbmuMlvhRaw
NTU++KkQq0UesOAlww8DRj0lpZFsSa6BzPqxR/B63JWW3unVx/9GGuepeB2h7INRjT/U10Ckk3S1
RLTcIpug9hx8xbsefJEAK6z9F93CQLwOXTcK4Lg6yOcw8j86eHoWzXNL3xk5biBMvDTc5CH+f2uT
nPjY4bEGl/BAP64rhID7Pl/GtBEPWqiYYumEybTrixy+4q2QBcelP9lVA5/4eRqN1s2UZTYf+qmS
mYc0W1RM7+AqMO54ANiuF6kUdd2cs/XPUWbslQQ/6CtvBXh+I6HNryny++6lcbu5wezdxYwI6vTD
3Lny9boOm2o0GJ32QCVnX2U0JvqNvZPurFdn1MJAuqksC60oN8g/T7kBlXsRzoCc0xqGkjIZDWkJ
UD9n0sh2h8ePMuzUwFCrAbzPqeNEfJlI4i80yQox1zV1OswkbF7AZbuV/dyUN+d8qq8i/xLCIUY+
h0Ucqdkbuo8+edoy/Vj5cO/R9xD7hGkoUodWIffGcOeprYCASNsZfdd4BNOvAuzTjO6Eo+ygi0hJ
6AX7SVU3WKoN2LfV/dcgDxPPhImg5XmEwBw42+hsCHTmaN8nt/4qmTNzxpp6I7mlU9JWtNvjo7r7
YyiREZFHFmYhkztclCVXTYmKHtxUxzRiiA6muOWE3WZsIymUdYLA2bIrikIq6sS6PGAYEVQ/O6hz
BmJA8oeKjCo+7IpAL3ufigzGK51jglwlNT8CpCDaS4dcTIbheSje0MSSernsyV1e4ELCo6+U2yTi
QVTgIdrefiyz+UbWO3oHxu4MBSmdOOy6muYPR9GwcnwklB098ZHlTqitYq/c6yA+CIrGO+A+Ex9S
YV/VFHBLRiL4ntZ7nzZOK/AwmqiRF3svyszZbdUy/OxUgfaBbv39N/65/MQsyzyQ5qbPxRaiOkHT
9X/R3T9N1xVzRrfl82bo7pDQOyvxGwIaFteZKMFSqYYl7gBIHPpD+fcCjTRNlu7XF7OwiRaxJgIH
4CPm0ldWcvFMxQTj8AENDdOjMF6PN7NO/EAZJbDXTIV2UGu7ItX7/3mnLwckS/YbZpOHGuV8xUFw
3ow1Q6nvzo9TL7O4Tt6jWdVOp+Tz+VXvO1uO6E2iAfJggACDFUKIVjMwPRP1CcAoRq8W0Opy57A0
5BF0Ivcl4t5IIgicmYo+xd9RjzFN1d4Wm0aZVlp+PxGjhrF3vEtarDRXmyaDMK2UQ3KS+3M3NpYV
+WFWG8mw5tKggv44OaMS12wcPjxZEvEbGyIJGFxnk6dPl+EstUVmB6p/n+TVCPL30N/dPBZo0KNb
N1h+1FO2F1wLkahieHGnt5E7NZ2ltMP9S2aG3mGtawq3cV9SOV+inblgBH3ITneTAeBG4ZnF5UMt
8ZG9KUnnd2aT1MiCFwQccdPSvhPw1V2CE8YHJJrw+byUSCLud3p6NgXLNYWXR6zispmj+NVnPTZQ
5p+Zgvlpr29Xrw5UPvQ73608crk4Hco92pa6d57GUBwpTp1obvImSRboOLSJqRoRDnhwtiBEyIGm
ZIc4tT5x1Qt0xj7NY9WYZzhbCYDoUDGO1Uk6QtUEtSQ7BDAJnYB3RyoWnANDL4wgfqF+6P3qgRJn
fsOBsaj7mKE+PTn3NU+t1uOz1xP6KxkV7SxVOCzasAhRrpbRR7ag78o7dJFI8Es4+ZcBLnGry/Pp
MNGZWUedq3OKkHfzwmmxlBmJT1oEFwAIpcJOdk+wOgYdUjn82QIXbL4fV0it5HzIjpSPUgqcxSrq
OZbkuRVzvRXsKAZ65TPvIgNu01EZryq5j7IEXsBeeVegn9m79ZG+4LfGH+2TwwouZHSeW1ncSFB5
fdgImtWhe2qaLFQKrrDDWqpBOd9/jQKGbrGNUdXL6B0TQ6/c8tI4mineNnIektZqxrSzkG3UAhrH
5oRoD4m2WbTs8gRE5dgcHZKb2doJH8uu6XQpuBVG9Ama5qYOcbM+Q9pf6HxWUhsCyXQSrN46ic95
WDRG0DZ2+VnzOm+bR33p/g+YUVqTgJ/7iby367Df1I9jK/6bHYxobsgECKTZoxsi1l145Dj65VXc
m+EJAGA+iHiWTFBm3LGW+XsUTliQuFCdZdFVtPOa1DgJ8TsIswGMrv4/mF/m36QzyGJAVJXsMFt+
+kaizp/6RJLW/enXcdLKY6MWAhOMNtTPqz3LtiVPrWFO/5S7mbNaH+LVmQ67h85mtanTPfutuGE4
mqDxBcOl3wO8Z5NiTBNcLgbfFmHq/HrZgO9r7FdO26FAbgWElc6/IIo+fqPVILZPKkNGxm1LRWn1
2U+DiHyVpm82cGs5aYnhOs9UE9CXCgJsCgdvOqyOanYM64nH4YblNDZo2cxFvI5yEwOej6QzJoms
B1FLmpNSRyvNe4ARVA05zQM86c54zKn/vWVeLv2llOk3dwe/tgRm4PtocR2lIAugVsJKYGd5XjnP
E0Y/+R20ePpLhhE/BMlizGjCaU+hha87DWQUcFl+tA3HUUVq4oUB9rj+MG8lOBCqCGGlzLD5ralG
1opnTAZsfz0cWhN4txED5EPBMQJl2AaFdrYmNB+85q8ZmNiTlO6QFfq6FkGspQqShVYoJjY+29eN
BeCYglaeQveDd9FuuejiGZvqUMxC6TPJvP9yjVVJlxdzfMXJp6UmxZ+FzWEYwJYZCkd5m6Jhcyj6
ZJ8SvTC8wOURr+ZCeafbbTgN9Opinvsrx0lkYrEWUsiBPHNt9Rmq6kGmriPZAKZB8FLgwDwEWGSf
/KCcavMb2xId9jFdOmoZZ07Hlj75j6ewPXA1yv0mOm3Fo3M5Px58p39xPRP8sgO18ne/Aw1lYmfH
AosrQ3NedfAaMu2eEAaJT6ZE8vw16QXRL3b6LhYayPAaFtuCIK6xGON25NdsVQI1pKCVbx5GHu48
wIBGBCWJkhBK9RGZmFE8rUhkUS/Z50HSqXs49o6qAbqhpoGECsPf3p0DADzzSIDFIrDkREv+H4WD
mJAgVABIJHwfC05f++tV/d0G4RokCF6sMqc+WqXqRqPzLNsx9s69pw+BcPrTjhzvZLZy7Q08NvRM
bg6Kgm+SkZM6Y3BJtKmNdI9ADHRszXyWMc46niRkiM6lXvL650LtrPulj1Jdss3fPsleMX/Wzolf
58N423scV1Rd4uQncBdFJpbT91bHUZyZjtUnsXTfiBRvoZ4DnlLxaXFHwMgiYz3MkhXFR1oCK3fg
/X/ombAo/fVBdGhHK0nNJRNMaxT/sgH1VTNbAUA/4v9YQthmXGZ1SkLQloNk5a7GYISIK8oesM2u
euAf0wCWdFDcG1+TpkRCRqGWLJh+G9t7WZ13yEV0dYLJfWgYCnlFoUBNTk0ExYrNFXtizlmTOhWt
KZeMS74qvVKUL6i3igeZTxM+YNDCEucDPfxwJhcKFyYO3wBPjKmgJjWew+7gA+FMfdKqRMNy6uVD
hCXcaSYzE3ob6dFCKr6HURh9Nxv+MX4DDfHYpMpHl7j+ayXlKEX1nK3lBCPJBgKH2+Y4ebcrBDww
pv7Dw+bgT41HSuKBnr8A0ROunWjYsZEHH3c0OLbUox01YfxccEeFydAISBjNPTMFNcR9ePeij+QA
t4Wg1rR/jDO/N8yGVHLqRzYkvbQB2gYriCE9QLqKsfcyVqOKK/UXzJA+BatbxFhYdaGt6IHpkV6y
woT0bgXV83p+IwF3XJSIWJ2oJ+zOnjeu9Rmmqk3eIacAW07+R5qM9DTl+kEx3mWwz5mijT8L4dsz
p65cbErWNIceIapGxGfRZqYzreHWeMYgBOTh9mQJDio4uOTjBplRwsutXuqZC+7Z+bqgLdjOCFSR
virwqSMjQtpYHd7h1QPgJC655FaTfIFauiHjySfC0XAsk0/vKwB8VYUucJc5AhgG7TALHnH/nDYx
1NiE8jf0YlfW8puq1Lo3R8CNC4o/Byra4WryhuBDhfljBGiAllny/2ZjGYSiEmnI6sHmeSW4RocE
Un5xcrBSHNaVlzyHbpahThGMo+QtupdbYYwMB7LVLxDL4+e9dc98LQapt+jKm5M0emC0jmqZ+EV6
Ra4ft/YaTugfT+UH3FUWbVj3GWcJQYs7DJ8Z+ZOUSqc/yRqgx5VZ8A6aSOdD4ZHQ8JwfGlmDbyT+
etwUcdT3MeVCZkREClGi1VEs0lRiia7kJHm4uGAD+P17IXHeHds93iRZbuOrhgEHtYzjZ9EcKgI0
Gch/vIy8vd9ot6nqgnTkCpCiKj17VE9na9iJrpIjCi/Hqxn6byqTkZJENd7SbOaAlPCBB1NDPYB4
LHzpBH6up4D/IipPUi5Te7stkbOo22bcMvh0crYwd1yCi3lyxbK4j6IWcAsSaUIgbs+urQLFLftk
xW8SXjA/TpdfMk3xAa5k3zZ5qgpj3mPfDzHhoKn2KPSZIkHB/vrM9LpClqtA620HJbcjwzqXfUJT
FeJMUNYxbx/XUdqnt82OxjQQHmkG7dDqyY1EeOpzOTLtpNUHPeIuhEXbAx1qqpM5uuZciQs3SFtI
/hfS4S8BUBoyhbYXO/iTQOd3rta1+7gdtWSVPqTyR/ZUUOvbF423AoivCuq6KtDjp96DUyqI8fmK
jn10TGjjSkijmz0y9w4uMtu/L5EFGr37+/ciTATbNaXeYWQ+AfNBNkwyWKCW8k+w1YpnVozN6grp
F3SAFHT4E7a+tA65oHwnDHuX/nzfgCDRHTrYhY1BhL/UkWxlQPkqOojqcntFELQnQTO+X8tpVxMi
YkyXVebgYr4X5kxmIwKteeJhnZL/YyBWd8lar+kYYMO5z1aixTWJIW+YFIMnWHUurf9mIvmhQURY
GCVqAy8fPQ8mJbYhuM8YHK8AqNnlbMzsOqavHb1MRQd14J8LkSQn9tKIRxoy7JD3ff1I++oE7urE
UxS29S5BdBgu+8Bxa1otI0mlPj8mEdvUJeV+qZeWKyA9+txnCViE7V+ZUpcqTbJ3rw226FoUOFwm
SMBiO+gDiD55VYH8mjO9CWBLK/kOcrK85wvg8Hhh3jwU5wJVHXxx4l/QttiQJ+RW5RHuUFCQ0Fup
YZ8Xbk9WCcs/REI0fKqQ3k9uJu/ypwmDcmkJAfbOTk0A7IdhQCz/T8zzNcWaq72Xmk0zjy3SrK5P
YesIXuBPDCzCEygcp4EeYfw3jTSw1qanvbgNzEcWF0JiIhz5/ZLk+paH8Bn3VF5m8GGif3dRft2A
Mqm4/zxMMUWwlGSE3vfgzTouT5zx4xgJNNpF8x9ITfDhqI24FxOy/sbwpdxurQRy9o8WiNL5H2ZY
B1VyRvw6B9DH2pzACqqybw+uO6afjzf9DHZt4+ZuAMVDAC9vo/9777sAoeHKUEA53A5hz8ZYcM4t
n5xhhydf8P3iyElYEfCq977agrCkgRz1iBVm5H/mVU4jFEp5obfqBb4f1Hp4qReFEI3NtNnGAZT/
eZR+viBdaD70AwdQ9aA7C4WeNUZwKmmzqFgRWoR/YqZxpWEtuUhABQ5szKZBc0scx6GpkGLCxRZJ
xGR2Dlu/M5G9x6NYryN4dRXaHQKWkF05AvUcXVb1i9YMqOlThMPCwYLQIx+2s+pQkJ73tEOBpZLd
o7rN4xw80r8FL+kISfoNgbIABvX+WoAd62eBoPpziSJhsi5ZjkOi7wKc4knDKPZ/E0XY+FKvt5ct
HZvPRu85YTKPBK4W88/6vezRqSf+nDJArcrl7ugJlIxGn7Fxwx/5Bh4K49y/91Qhvu40rTzyVvyQ
t2NgOkdTAFuvPOI/x+3W3b2UW5NPN5GnQxL0wq0zn8U/ZTKsRJN2AZm+jtxQvxrudGeVG7VnCHOu
FS4CcarjhTio6BVlS3PCdJmBwefrcEx95fZir57qrUQC0SJImJi+EVQpb4XGsuHHiwKPjASdjhrx
hP4WnwRqUh77UN9Ft7xZ8/QZo94vxDiJXXpl3nYV/ul2WaUP3ohoym1jEqHNslPuJIm7aHTHDS0h
hfNUBynqq2bfPsfxQextPITdyxlnlIyR7SNbuh+WpSBXgUXlEdM5c1T7jQcEp3x9NqmqEoGsG5OK
QZlAxPfrT3PWpB1HpknwaNTL1/e4XvQ8novdYP/JkdEwhYaw+YBAPVnnyuPYLUYIqRZbMM+QucLp
b7iTofGp7/rotXVkBroJefXnxd3THhlV5VDrFrGfgCIii1oiPUSX6SS+ZORtX5u73l7/WcNHTKC4
IgS1kE+U1fLjoCY7cDNUb2I9R22sd1N/LW28GPIYgTxGI6u+3MH/vicUuN+XjjNVrFLVduSYcheM
K7WZ6m8god0fpsSHmBoMuWxb9CxE2gOIotz2TvbjaYXdrWiadHgsl0h6RDiG0hkk/rlmAKJXoJUO
EOHDUcA4RL5G2Jzt2c6RXdE1kiwikZKxctOf4T0s9t3XPXWY1JZ5D7geffPeT0+LKfu2lWN+XqlR
0a8LYD1r0qE/A43jj1k0lgn2/Uu4uArYOXflpG0bG4g8WhkrBubste1HODGqKL2bPjMvxzBEBrIr
zL6zZMWOkUgdt2wm44WalrdbVG7MG8xKYPhMhVNtyASGfSxzg2hm6TiXBcSaWj4haGo/lyDf443F
Vs23+9yuST33/IrHoiriVoOW4nbrAeaMkUCtsd3KDFZnfuChS1f68WWxYMw+YZZDFdLx6lI6DtZI
yOeR4pB+TDBtlynMGV69g83bO/pCYsKoAPLRCxeUlRkKiytt5JaMK1rmVj7WQm+OSC5RWLfbKchw
TDCCgSRqw6z8phuWFhW1MsGiGWLmmXyjqleQxZphM7XiOPbu85+aOuLveRbOW4O8WsR1xChDBRP+
jGhrwEiodIns7+UYxbOnsAfeH4jyjEz0bFYXeeLUrSQ0v7F4oNQNWbuqXd9k1pQD0LweQUTgmnEV
B0kpvPiGNiqkcxN6ffh2ZidCJ1w6NNE3lXZ2dl0SdMzB/s3LwiFKZ7MvrNFn1aOm+IKD6AGsMxHr
enCWcCSzdMjRkbA8+ZgD4OQzuuMfBgW9B94Hr4rMgZGfTaHM+xthMKHeOMiq/FXolYxFCYQbIx9J
9naxE1agNJf8sY+Ckqw0aLn0cwcOFuVi+/ZLc/asBeSYTWsHul9qtCy2kVfA5/0i1x8dzIAHiiJ+
xTiTd4OinUSU6F9Uvncyj1uAkDFsUvjca9wyGhYQ4xLCwuh8XIsl9DVqKcxoskEIFSH9435HR9Vq
O3EBE6jfzYsDv7Xe3qsVpQhxXSFY9cnLznWJ6CfvVel+A2lvbkRuTp20he1+lCNKaKizQNYwBSwi
Bm68wWOkW+XPSDhycCrpuVMpgJ5yTqMFxAd6R+zpE7Z+hHy+1Kh+UGa/QdCZjspaCa/YPcTU10EB
hN8Pwtmo54uhlZuRrQb1ZZpq6eBIz5lrhLfLjmb0fiTNX9oorOuyWoyynuCNPczUE5JIlkIcctii
7ogtjLKi7XsruOyQMtNOQfV6VWrr9LCDEh3r+4daBLTflhTfVLnddGIZzDaqittUKfHOmHZ1thcv
MXtwnUZI+0jqNm01R15OrOg+LVmLV8XDXA/Yfj+1+vBf7dtPa3Q4eZ5PWhU1vbWATBfjKB4cbqvy
HUCCWddT4lkDTEhT2EwEhZZNlZpwOh5G38apdtNp4EZn+GORVyELZacl0tyv1z+oE3Vne7Jy7FLM
RoYOFYkCRLu5VSs5dorgBj3U8yGSqXrZ9HIHjLbkzbhm+aqsBNyPx4vi9UimwQp1qw4bChIv7TfW
YzpI1Dn6DHO629pyTmaqg70uGaAWYQuZ9zMm8QjxAzz7A4k0vMIz4Qwcs+u73ZhkOcz186XL8OMW
+GB3c6H2EU5dO8Xl4fs7/JZ8KnkoKxulvBvaUbwMlH4LT3xuJET22Eo/PB7nD01mFUOh8ug3MNz0
ySJ8WzkUsd3wQIMMDKjL5xeIdZCr1ownGeAaaCI2fZEjEvyrAocdICYAPWQ4RdRRTG2UUL1eLORj
y6iiX/WYiv0qKLnbA65ecu+GsEFvyDP/Lcazuc5Ey85s1rEHslxD8NLRO3L41uxqWEu+y8lWR0xY
E5+y+LikS/8ZvHYVPZYSXzBI0LKvZJRLfhL1bVuWmkZ7m6CcoXWiqiAE1qu4+1Vj4vPzNbcAdJGe
YLPlI94x82LyVPac5NhCTQ21xHt/gV7l0+OHCgp++CKfWzE6dd6cy5WvkSM1aM/TgAzeqVD9ARBO
ZoUIgHOTpTCjGAV0C1G16EwsODOV5RO6RxcJw7fkJ3iWLMDI36kVG5DlehCAt+/lP5YmrUhLzlMt
p/yHIvpQ5p3qcJ7DTHhxSnxxFrgXrn/Fnqrl3twVHzVWEoITFkn9HRTXpUQ6rTOicV6aXKx4qFG4
ESQsiK+HcbXDCQbiYro0VjmG3F9FQOK5lVHT5t58z9B6sOvQJ6QTxRt8HmpuZgTSuAdiYxrq8d/B
KLJvGJCiiBE+byJpLDv1pky06yVv2AXFIDkOWuikuAcgihgrj3j4Ad1XXdPHUQqqvNuvCs/auahL
tuAbOITQ3MQYCgXx//uJ/D1smUWFalXiI5RQAwu5F8osl3X00oWfkMvQFVH9nWttGosgeoND6wKi
DCk/SjLcCHBXiBg/VgQbrmVXmoF6x460tcZh9tO9UkD4ro8WT/LgTZuQPNIS0KpDevXD9SSI+yUM
+8tkPE+2JbK5bF5bU34WeNXJG3Yw8Ts4/b4GKD1O1VsiGllwesUxZ9FNhDVoDeLqRiQTrVUoYiuQ
N1UiyfGlcW8x35jNFmGUCgtPDPXLmJoNHgKq66zdXN7va3mQ8bJ5wZTrFBHT6lQ+Aa3YSpQhFonl
StNo7TAZfBo+zZs/ErWapTj8EpAiCQPCiY27/Bt4m4ecYCWVdxvSSdcuBlZ4N7SSrnQMgGV35kJZ
hTvIDxGe3I9QVHQ2ttNLyHVOgN3oy6qRvpAfijaolGrQ+vU3/lpTuVVha3uouJYeyDjMMxNqUcKS
1N+hovFrLRMTBOT5+wem8dc/m2TgSYv5amTIdovK8uV0ZVXyeJoesxiMs8eBC60/AN0J7b74FILB
eYIByvVKK5yr9K4Q+iKq6D07lY0oUlcNzFytjVfDwVFv66s/DOJ/u5rNNFhtc1ILa5RA9/+vvgrJ
TQHsSfoZytEASsH3xwf7IljjLWFXhikR8D4fqMttiqdnfVnbbl7ecNeLY+VgZDKLYCR4wZNQ2K+R
ky2FW10oA/pyqhz3Uw2EAR3RtYR2puAOQZvF9/LM6fN/DbBnUWVJN1yhUJPdCdsCvuQu8reFdrtZ
JOUfG+zp9h6uz5i1PdZu8r2WJUrtVGAb/w3VcZaZBsPLlw1fvh/7DRhfU1+ZHYrDO9XMrkFklB9V
TRtHdHc99b/csEWVaM8iEFnpFy8F8gAMAneCFZ5z+zu9Dr/4JjF2oa2H87CNzwx5SU8cAl5gaJo9
p+PzUvpn8Wv6ce6pNJg4jOmp0Fmjvgu3dzwa3jIhkYb2EzV1m5EXz8ZNQrGxQ9PHnokn3Xea8ziW
uvAZWQ7x8wB+i1y8928Lp2ltSsDRzR5R/d0EwQCLQnThxsNcYIkGKrlabtR1kaNZ00PGl3FkRbXa
5ZoAavuyoOdxUnRRoLgZBzMojuxb9MqCHAA8lFFp7g+Jnu0uRqRhQf6vPLRtXYjrlypUucuClvHl
w23Ny6WLI79Xez0pf7v6WznSdcENzCLgozwot4bjoJcuSBciEaYJf/WeU4X2Mal+SDbyZrAo7BMl
j4nMCAY/elWW6hIzNMPJXz3srL2aB/Pi+pEz01GeQQfAvmJwIZ/baWq77ehElTwq7zoPja6g3czK
wTDz1nh5IxCBT1fTRGmMT5w0FsdsWIXHRvyyMC43MLVy6v1n02xksS+BuOXUKnHl4IdCdzHjmy5k
AQXclrV2gqF3OKti4ajDzE8R5zQe8d37bxAbgHvRl5S4n2cQsF1pN5vs3ljkJ/l9bNbPpn25iMzX
NPlv8Uu3CqGiCzb4uOshKr9vFA7mWuGyAudux0sQRcoFW1VX/OxsFSYcNjNnV1tQj0wIQZPm59hS
ZmlDd70QbFQisGHlTJfmXhykUnHidMUxvtiGRToHhpNcTj5cLVIqGddkWfGn6HlUviipbZQCFFc+
uGVvBBdNU/4N0nAXPP9zaM1WVztlSVqrSFz27GrPNRILfi/ed1lr584dz5kwkSXIEeiFdy0dVmCv
BOYVPauve0oIxQfq+9PmmZF0LDi5tqmEL62pd1Nqg/UvIJTaNaQYd+dczJP/6qmT9mcbiPPoEaxN
Ibly9PJpInGs+sMZkF6Uyu3NATTkfVqHYOqUnz9v6Hg34QyvAZ1XBYjfC+Gjds6nwt5OMPk6EwLp
/TnVHVlDFAVdOAcJA6AuxZ9lXj3Dpw26B39Xp04gmvrxDKYtnVsvkXGa7bld8ibXhQISXVRUmEOg
qqDRH5XRptkNRcp0u5KhrT4Hde02rLA5zw3uId1Vezemuu6MBfGfZxfjJHDgrW/gp2MMGdq1WJ1T
yG9280fpDtPh9uEe0ObRzlHuJGB5LP1l2Tyb0aP4BmT2JMGSOpHV8zSfWgUD6aIGyEcWLSAHsoXo
EbrSn1Gw+s5XWDay+ySgzXGTX70vOAepXfQz4Hq7fEBL8zgBmmFTrmRgWD7irpaeCIVzW19yjAGO
iLkBSpVctLyJ1CbHgKxotyWoo8Nd4d4H3ViqcuFr1CIL0TcWjyXsX63Ejy5y+KPdxY+aweMkv9pH
Kyeybd+fBq3NZY5admdhfJxo9keXGnLIjP8VCKMIU1wHZzzNvb62Ma9OQAY/5UtleFlXHlda0O2B
YQpdHFHBF+dOqp2n+A5smI/dyrsK87iiwBytu0ZvkiQZ24O2ogpyUsuV3keczYtfvbkn/0aZw9oG
KUKIPNBFYBftd1All3PRQZoqHfrY6V9PSYORiroSvDqsW5mXtxkp9Ubi/MEZzKB8sLrmyRJ/0vJN
VkbKVirjQSrIZlu6yeUKyX2mY/5Y4AbXfun3aKYbGcvthhgX0C6xH/+y2FCrzYjnYSNfGoXJKns1
z+ovzpasIx8p8wiQpAOKq9B80XpZ+Mj3dkYDX45X5M+tqRPEDyD9MBmwBhbdBtzLxq5kE9p+4xGB
ax8YmOxjUNbJtpFLotbqHHhtPsq3iXNWuho36ww9r8nKPNc1BYmhkI1s9JYLEGebaIg9KTty3a3e
6DUx8kIR88PZ+h7o9kZGCEW8zmQMdx/cj0YQxco8USvXj0I3Lag4rK/jeFS/iR4b7M8+8qGRSVFO
U6UGPkrEE4Vb7Io3aEAV0D20YV6fRL+FBOkTUHc1OnGhNzUj2rToxfX2+WXYVeo9v8wzt6tPKyMY
3Mc1zFhE8AteO8Wq2NLkR8NWaxEjqZQurAUT5pWKKXeXCPhhb91j9+GHibeg1ICO1sXiFufPIN4D
m/kPO4ByAl0muCqUaSImbzKnVsvSHpvRoaKOb8x3w32N0y5ttvL0Q11PR48vZl4RSrjWYnUhxKCS
bAT0Yd9j2ZzrOnvxZ41XNv+dwGiT+CnxfNtK6Ijajbm4crEQ18UMaZdngnKFTYEYo+skoiUXy1Jx
yH3W/jZX3keYP6Vq9ai+A2eC8hvZK5rJ70IV8xmMVavVgVBxA2J2XZExOJjXiO+UmL2KHrxJ/x21
srNwO0AZLz+LEnEYlBox/valpAhQp7hS+Id+WIMQvzWG8JLq5pmA8wbtaoZpAln8HoCK4XBm6WlA
GfTqQ5Ev40y76YL9jz9PcXWL+4QgcBmBzCONN66QRVwGh+W2vZg9TNHMLm6uzFOTtGIYV7JZTZsM
ji6XNCdfOFDWgVYf5ZRbFLoStAcBkTa+NXauzj4A2aOBPqfNi13RKJpnRiIIdI+zrIQrAh4TbV7a
BcyXCfD6x0G2StBbF5Ufa3nPoqmHYT3+RGS5QJwEelNCW5MbVCCg5bagwjEMk0BB8nR44zgu1yAf
kttJtH0KRaFc5YBTXYZAVbTYY0rLfTSBFKgZxCByCuL0V9npkFDCZPRw82P3hGrNREBy9tUVfuJg
kWRohtNu/DxySicLIptqIE7LYavI9Cg7fI2bEk4i9t8qxVSsPTh/KA/xdpYd+xERrW+DX1KnDpJ4
8l+8JSI3+scBhUmvqyh4qwrqyd27kEAapoPNpdAjufE/CwLwEKDZ4sJXM5yTlx0kkRO5p0orrUFe
kEq1bHH9y/eB6wWc3YK2vbWUho/soLDEf2C6xBUJS6KVrOfRRrwO106JetMAHKBWWCALvXaANe9t
JfDGJ4L7DM3YqgH7szIMT0cN9FTM2zU9+ow8ksjNjBIaff7WNz6K/TqeD8MA02wOwWm/L42CEQvQ
heQU6itmoFWsUuWUI/pDXUxrnDk+pII6/Y0+ILxLR53/lA0tYZWGB1KalDZF74h58MWJji2DK//y
1wLqvZr8NwkbfR77q+yQ4T+C/L4q3a/Ofst6YNhbSrCKEf1baCEyJ5Ni/nzCEchttqBeire5rNUD
aLi1ReHTycj+notwoD/pbALN6iA/iOn26Uog5gPdozbdiMe7gXU7KlPXBWzTv3yxS9gwsPHXv5Wl
dwnDdjX5ftox3c9Av1YKnRnlsBN3b/naVCnRyhbjrAcDJMxT18zMbSedHHODoxumfN8Kvi+grh5d
Q4TjRD99ZXf3a3kPYiBYh24PBHiXn56dyxQ6AOdBPLnAxqOqQNK4s+YIytOh5hO4RtkN5gzFfbJp
pY1tzXwig9txhY55DOMapxeIs8JktLduubBFxn9wrxZn0RzfmIMmqw0+hTfFIIWrfIsS2EvJgDyp
CGaP2AMSaxZLDaeXdNnuP69TBKkfp/NKofHehAYGYsC2rkvOFQ2Upwgx3rXs8YhLc4VetT55MJ4q
+HENyBiisKF0BFUTM1DIWjhf4obgA8Y8vn4BF5OOFdIRRyN5MoyELvAll+mUFMe/B9i+WkbVn/hS
SJwjs/ywaCazmUMvo2XC+/GOEt79mwfhYVUmUzhz5IE4uDzaKgPi2oHE1lQY8d56rcw7/0lfNdyG
K/+RzOXAyOP4XpJKV0AcjzV4JWwi6QGUpEyfw0yaGuGDGnB7kMwxtxbbrthpjHWHlFQa7acatZgX
B6ENGQnKWsOQwC4ScFUBwHc8bHYxM0a9vALknUaMxGlmntiW4/Q8/0SD5GP6lH83Wu0tzxQAoeBa
gphqGa0sojldOWGOaNUxHDefZadcJqWJIJesGEqs112ygOIHbb0sotZo//HtLQaZ9yYp0RvbG6HT
+6IZRq7TbaTJo/JTKrlyfaJm5yjIO8/OYtRKigbR0UkQCzsBD5cFttJcOloJuaDN4gdSRcV5K0NV
wYu7+l5nj8li+Y6wooZcfeOQiqqQ2P0C+cMrvaayOySYDt7mc//FeYEHuq0hNwl6wkAS3ucRSuJF
2TBrBJmY9Q4J/GfCR883psVF1vA4UYB3ehjS9wxw5iUP4G8R2xuzoosJiOvSZ8RYaM4p+Wdp6RV/
xX5HWCcyCJUgDnuoAIbhIWRLvOG0DcuiS5ygievaDesDP8QWCvqowMZcVwfVgsrjEqHPFsfc8nHV
ncqEJuaAnKq439XPy68/JdzvL3nSgrcWjLK2j8H/wLYS256RJznG3DbY/EjUljV2+77p8GC3iv3l
LchBoHC7B3qh5NI8XABolwNzqljNjSHql26i1f4e8bijxj6h8aMXFA199XRlqo51N3hyMcOZW/06
0SVmEScLYFDHk3dA10Ol+LZaVfUXNEL3XGMHYaxVuxZgcB5NMLHhn4Xbq33SrX1psHTo
`protect end_protected
