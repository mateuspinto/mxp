XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���GU�l�gK�ͻ��8���e��(v^k4qb'7�z����-�;�98��Ҡ���P�˞���3����b�)��g�EUid�����������2�$�&N.6�;�+���#d��1e.U���sZ��$ ���'�s����=�+#`�'{?f	I�m)�I	�F�?	��x:XSӔwLf̊ %N}�b��{B-}l�)]D�g1��˙�� ۭ��7+sR�C4�za�T"�}�I��/������%��0x'�ߞ�-l9{������'�ǹ���L�-��*��y,w!D��%3K��Y����JT&�\�0D~P�w��׀B����`>]rz@���~9/?�(����[�١�nwyɀK����y6Db�<n�)��o��w��S�*#_��}J]�?�����ӥ�j��7��4��t�o��n��a��Z5A�o{N�h���+>@�i]��ƶ4'���i-��<�p�(�cg���K���9-�a�.��d�TFK�H�#��>0�uv߈ބD��G���/x����*��>�6�`������(��j�_���uS�:����d�1��3AS���`!��c�2d
F���.O���'g	�R��u�0�R!�D¼o��[��%�p:�C���+h}ϟ��vȑi�q�/L���K�#�+1���u��,����'Նm$매�+���k��	a�P1�&1���Ŕ
ih�s����	U�H;�^XlxVHYEB     400     150�|����
%�'�І�P2�HL�Z5�=ӣ|Z[�����!�'���]"Q�KdcX���aV�/\��ىh(I�>�%֪_�� ݐ��|�!����"�v���Y�}}�y��@V<h��,��T,�$<GN�:�#>�peЖ^���nI}�F$�9�Af��2X����F��`bX�<'K��԰��C�į�PF��t�qψ�qb>�B'i�M̪��U��k�M�9�]|[�=�Y���1MKs�I�Ύ��ouQm�����&P&�Fe�+?ր�ohg��fB}M������u��L�֭�&}|���rS����G3�� 9̼M�JfU��/���-N�93XlxVHYEB     400     170?�<��# ��'ᴊ�K�cm����/�<��3󣔠7J�3�ò!���8��?�f��b}�v�VM�����;�i���L>����	6��h�M�F��7�X��C���{^vKǔ�؂i�F��9p���H��L�D��,�À|��|��˔w��(kh��]A��S�Mԁ<7��Y�`�����U *�[eCa�r���s�({�<�ňv�f��)k
MC6i\60&h9�l,4��Yp�5Q�q�}�_��	ʿ�Cc!.P�<��U�W1��z�2�Aj/$����ʻ��>^�$�rYV!X�H�>��Z���V�� ��6��	L
N<�GC�w�9R?�;	�9�˅2���<G�sѻ��RpXlxVHYEB     400     130�a��Q_���nb�nM�u�8č��T�P�5f�w&/:r|��6���[?���殷5dZ��:I2����>�C�^t�֮Y�|�o䠣�6�83÷�X�P�l`���{�.��l���$��@��<^W����V�V͔�&[/�^⠄Iv��e�Mi?;��$�KYKo�0[l���>q��E$��s�x�5��ѫ����y�WÔ��D���.w%7%5�H�Ua���U�9�Q�X�Pe�7����E��u����AP���Q¢��:\�gG���oȼI��J(w��c�%��y�3"7��LXlxVHYEB     400     100��ދ9̙*��~C���uo��V6'0t���JVe�P5Yy�o>� I^��εpWm�xm�Q ��@k�[F%��S��՚�f.�� ڠ)�P�bWp	-�Fy�s��M�)�83���1Sug�`�.� �ͮ�L�, �I���{�E&��僘lA*����nr���;��=�P��1;�ۗuL2<S���:�.�~,5^5�@��Yے7nm$u���$)c��\��2����6��˾�|���5!ȱXlxVHYEB     400      e0k>M��4�����?�Ba����n�][����/�b�Fy�u�@E�q,<v:�.�[_w)��p���
ΫhB�1%N�������(e�v������b�H���`���VM�na��ݙHa�yCR9�$i8���:���~>ɻΨ[ں�d���t����j�����te6�\���XE
QR�ú�D�|��ҨM��@�g��7�`\a���i)�XlxVHYEB     400      d0&FV-Ӷ�7rai)Qp���/ �кvl�9:Hmb�ok�&��uQ�A�$�TN<���3{��N�}��?o�\��V���Jo���F�JR�s�l����\�r���ܘà�����Rg�q&x�,~p���U�@,�R�f�O~��
�
[�FYCp��[tD���!���Gߓ����*���F�@�{��5�~Zmx; �Ɋ�(!�b�]�0�0XlxVHYEB     400     120H���E궳� ��o��ܷz�r9���֎=�����m`ZE�z�TN�*9~�v����z�
NAy���+���R�hh��+���R7��*c�Y^��*��}��*ʚ��%�j�kQ��WvG�.r����V�o�d�?�w�v@|�W��2�6�mY��@K#��J��.;���zE~�C��sXl�l6�a$^�n<7[嘎-4@�wA�f��B�������N9@��Cib���`\��d*�)��Ïςr,n�LAJ����� ,��cv��>���%�+�.'`XlxVHYEB     400     180�2�1.ry�:8*@�c�=��λ���\X�D	��vm�bv�i�������9Pvi����Q���7&�{q8������,*:<�0uG=�%��:��F��cv�--�����)�C��c��D���p�?`�<l�	�e(�f�[HN�� �˞� Z4%@D\�8n	�DP�c��|��T��Xz���Y�'E:�:p�����i�nj-i����NzQ��X]���'����\���*늳al�C�������*n)0���:\vK8�ꟀrI���q��J�[X����OUOh{� ����G��[ߑU���ēoyz览S(�F�S��f7�N����=$��EL�ʜ`N,��hB�ÿ���"�T�B��mR{ ^흺^�K��_*XlxVHYEB     400     140�N�yPϵ��+���%�q�,}E@�7K���-p7�D�9�<�"�iN����N�2�/��R��d���]h#�����K�㾱N�Kx_qWI�#d�m��
!T��I�W� Ak ���}�$��0nc���K�K�<��!%�WA�b�	��"���q��؃�=�]닀2���8�¶.������jA_C����x�UXaޅ1�(�I���0�`cƤ�����4��i�� �TOq�A��G&���h�3k,L��hN&��._�'�(��5�ʪ�P����D6����Y�<.WL��W��t 2���_���El�XlxVHYEB     400     170�r���}��-�����L9�]Fy<��W0(e݊@c��ZС(��.��"��a���Ȗ?��b,]� ��h�_Nk�
�IOȮt:M>av;�p�>�P%�ep�+EA����ƫ.�~��`�C��.dc�x�Oa��6O�+��^��"2c�V�>���U�����s]��ߦ�Z�����ef���my�-q�.B�Da�l�:¯-��,\�.+�*9���V��Y�f�G�Kb�W��)�ީց��u��#�ϝq&��e�(�;��ש Ky[F �s=�Լ�@�����C?��1A�?Lĺ�j˘v\x�I���|�U���kCO?|�3�v�=^�(�'l�����:��f)���Q�0��3XlxVHYEB     170      d0��6\X���W��J"�Å�2�����>O�y��NH?a#X�)������c�"��^S���A6�ԽE�h������A���U�4�聻�}��H\�\]+��-K�z����ؔc��A����ۖ�8)�X�!<�7������PJI��J�~~
������� 2s��UP[����.���=��w���B���y����a��