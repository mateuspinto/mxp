��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���đƼ?F?7�
�=�Q)�Zi�#��R`P���^��W;�, N�{�(�CU*i	N��"�3�PR�ZX�i�������$�rXM^���3�W ��!Y��E�ٜlژ1�<AJx��ՓI��p`��;�4���̉�wI��o���m�FH`|�D�=�O���'����D�jL��A8�$��D:�An��"��Ok篬�<D9uY��.M�J��F�|���~�X~ef'&��c8�M�7����.���k�Է�N��͂H�HQ�Gu�mS発�a�d!�?ђ��:��(��U�	'<J[)����Fb�@�  ��1 >o.;�NpJ
��;qE,��C�k9�.��bn��,��������=/Ŷq2`�e���+��b{7��}�yp��wܥF5ɌA��T��6����߼��ۜv��LIW��z.RfծS���n�t������H���e�ĉ3�.�ZU�J�W�_�r�zLxRJ���9����	�����To�����*�m��t8�C�uA�4l�����&8�{&�	D��D�B"_
�Ғv�+���E\�1(�������A��������@x�O�Q�}�+���G<�⵵�F��:2Sk���!zf�|����RWڕCo�|�dQ��j���T��v��_'�D��Y���%^�#���bܛ+�"��h
���eZ��Q	��!��2��2}�p�Q0�ч��Jn��B��!�EQ�ϻKz�rᄾ���W��0dIH�n�)ݒv���ͨx\GZ�N����m
)v�{^���e�;�9?|S�)O�"C��N��5F��(��6oH-*�_|��<`�xq�x.��X�`�\�u�EIפ{��|0F��ߟ`B�ޙ��[q�U��׎)�~�	���h-`��u�;O.>�_@�s�@9rX�ҸA�K�+8�b�� i$�ǜW-GD�n�$�-E�����ڐܱVx�Є/�r��c�g����4,v���%n�2�������LM�[�ru�~��q�0�ڵ�4h�49��g�*�ʴ���q$�ȋ�2���c�*�v�H3��TLn��E�/���+Oc���{ |�Wq�P㟗�g,����]� F�B�6S����f��� ����i���L�+l������m�%B�_0����b!D�t���+E+I������M�8n�y^�p*}U�	�h�H�	C<J5/�ͤ��]!�U �c3�K8�U�S=�vG��סiD_��s�VɌJ ������o��x������]}MB/+��&�����g�P��9� 9��%�'�M���	�~�(�����P����`ϓ4���7������]��-��M�`�,��e�e)�g�V�j�<�W�W��Drm�'��~�u��*3�w3E�������x܊�/�@J�u�Y���n���N&߳d��4�=�P�a��� ��[�k˨,%{C0mj�醠�`H������5���S��i��l���M~���j�Bd�'��{���O�4���Y`8�Md1���f^���ܣɾ ��d��)z9ԓC�r L'�Z��!oCy�Ќ�����_�AB��7ܩyX��C�����k�KY���9��WP&�CF��X��G�cClzE�"��PE��ޔ+��`f6�%��x�O��|�~�vJ!���À{�I���bP�U��}���9w�@�� k��?K�m,&���*��s`��"�
r��0��Z�H���?A^7Ҟ�\��"�Z���v��F����	��Dڅ���h���	�YG�#=>d6ǐ�@w���l;е�	��~R>{@V܂�u���#.��4��ǟ�����O�[���f���^�BDB5��*}�ȼ����N��:�7}�@����H`YX���yQ]¶�H��_ᥔ,�*Ӥ���I�������Vt ���2<�%��8�$äX�Ֆ�ě|�F6<��VgY?�H�Y
H�~���n��B�L�"P�L���Tha.$�&ND�J�	풆�&�Q"%W+��{�K��qݑ���WL#���Ꮟ� ��J�m0�d�?n2�y�5�2-�4BT�*���ǂ8<*"$ZUfX��Xj�M_3�ϳ�[X�VX��~yE�&�d�^V��غb9��x����ִҐ>�,c��5�n8�L�A����wxZT7���/�-P}��Γ<��_p���8�?L>z��V�j��o�,�}�*�����@��
=d���nhKk�Y��**	bM������M���*t�R]��dk$�^s&������=[wX$�`�R1�j6�OiLX����$��4�4 <�C,j��>y� �����e�B��s�Q�w'*b�����t���5�~�I����F�D3��n�R2$��-�A�:�i�!�V=yi�Q�/��coh�l^g|V-�u�SR;M�J�aָy�ŗp�����Xyc�F���F���V��	��cE��%n;A|E��y
!k��+�m�{�Aښ�2�Y�+�ߩr�
�x8��P{�����3V�Q�$�W��V)���+�z2C+���'��&�����k���(/X��0�%2��G��:�u[�*�F5���뜸 [j� ���!n�`�g�Z2�>H/�1�{��xC�E#v��^2��� �~��y ��Iێ1�mB�8�e6����3�דc�~qƛ�1" �d�aU�X�aӈ��b�]G~��b���%�|oZ23�kG���i����tV���?�<��9)��Asn}O>g��v�#�g�S��H0.�fi��g��Հa_�N��>�18�!��P�E���L���-O��ɺ�Z��� ��:7�$��M;��)!�M��l!@D�^�m�D�>�Y'��EM)b`#pF?_�'_wb�|BΙ����vk����=0��$��Fq�c<��b>^sj�L!��TƩB��jU�XG%�����֟P�ӽ���_�~U��b��<���D�@o��<� ���c?e�V��������0D��rhe3�{2q~y_|80OI-״���]6�=��O��m%)܇�ϱ�N�v�0M8)�~RVN��q�X߭�	��ϫV�Q�3�W\P�ϣ l%M��萏}VSÔ�sL�n����Z��#�rDjj��b�܋��;���r��F�F~�����T��h/�����qV�f�vw�DBG!q���C��U��lZ7��=$&n(�[q��L[4ݓ����g�5�lS�����{z XnYh،ژ�;�a-����9��`���򆠑G֍�u��,
��9�#�Ш�(���_j�$Cm��5`��;�=�e�@�A{�� M���U������֢�K�����xx�;����u7]]ʒ|�Ѡ���LD���>S�_��⚈1.n\��lB��5����n���]�(������p<^)B�� �ޘ��lW#X��BcT֍�r}�0jZ�)2����r��j�.��|t�_���y���7���n>����=����hG�9#H�Ґ�"D�C�3���#���o���:�t�Bdi���K�@���a0i:f��TDW��۵����չ=��,��6���\���iP��*��_�i�8@qUx�¬��Y�1�ŵ�+��Z-���q%i�br �Y_ZK��̱-
��'a(s|H��;:j�%" �����5] �}�&ɸ���l/�N��z��A��R.�å�����3٫�Y�5��XϏY�5�&+$���y��=R���,��'tRa��j�Rx�7���ow��������4s�%N<��
�G���ů 5p�j���~�W�����9W��"�p}�t]JC`�]�� ?N��nP���Th�Y i�`�%�ʹ�+HM�i צ����F�
�'pϴ.}���<�}�A��@�.�L���2yjqE�>ّY{t�*T0\�l]��Y�(Xܿ������R�K�.��:4�L�X3�͐"^�ߖH2!1w���x����e7Sn���fs�D�"��۔�t�gm ��F�̴�ȱIL��2���_�����?Ih�"�2oN.�B��	#²�>G�L��@���ￔEy\1%�܄�X4��i.��D�9V���s��Eױ��پ~�!G��������M����eVص(��b� P��7�H\���T�k�!_�ED�i���YW3����7nH��Y�>�>�%Q�j��԰ H��7w�T�m|�t*����u��N�.�(!�Ϲ�Q{��Z3�K
eG��^�^��ȫ3�H�3w�U���r�2��4*2K�z"ԍ���S�ax���$���k�����r�@ls����U�a��#~�<r.�@$҈����*�\��)�zh�a)zXྏ��a��������B'	�-�Mz�s���}�y}�NO��a�J������(�����* K��a�@��6��x;�<MCO�P�v�n]�8����ʂ�����MF��5�0��љ��@7���,!�wE<1"�� ��z%X��h����^Pk�tw���'G�A/~�g��b`�4�@K��cY��/�7��^���B�R���G�l=퓳��3��H�N�,`�Ѣ���E+ؖ	�ß�c�bP)^���5n�߼�fy�
�c���Za,���1�����&��"F��ݾ�6k�2Ǌ�"o�0}1��p��E��j�{]O<�Y�|[�%��N�j5����vhNfu�b�,�;ŷ�΀�S|�9�*3�m*�7�C�ȫ�|����m̯�@�<Y�����w������t�K3K�	c��j�Ջl��R���	�]�Iu.5����Ք��^�N9h�-A�(�����.�1��i1r*%*6�g����ׄ�f�5��
S\in�e�z�})� ��\��t�D���sۍ�Jm��.?K�v�ڥL��L4�ȹ����'�o�i�����#I�����>"��b+_ �gA#�q�l������R8��T ���Z�����R�%�7���֏�����8L�џk�Q���.=�K�M��f��Ɯ�䁧��������_"����I�Osw닰
�+2���g3�$���=7���-D�Z�X�_�L��A����qzN�u,9G��za2�LUį��_Z��
�c��w��C���'�p����l���b���F��� �{���?���pP[�q����P=�T�$>:
sU���an���t�>{�&�����g�\t�p)��?<���ɘ���6��8���eQ숛ߝ�F�P �P�!	�����k6�OyKhe��E'@뎵X��:390���@���A�+�%�w��j��$9�NI`������]_!���"��H�qb#���<��[S����
^,l�׫-A����e�Z8�ꐏ�dd�(V���K��G��Q�L� �Q�|( �.����Y,uf�Y�y�ˈ?��l/�N(%�/�f�`"�1NW�T��k�Ѱl����*Yf�5gi��3��v�-l&����Sm�#��%*�f�B��:�Ѥ�@^c�c����,���̀������u���2h�?�Fz�����Æ�R���l�&'�>otg�H�YY#>=��2�o�E�7!��!_��oo��X~_���~Cy�ط��g����J�S?�r�x(���K� (Y_�{O��?����)�yv�<�\ ��)�8�}@�	"�q;�2��.�Ͷ���O�	�R�NC��-~���t��[�7o�u�L˫����e�^@Ŵ� lwJ���MbP^d�yr�H
�;�d���&w:��>KV��ñ��x�d�qh�"��s�y�T��:�a�"����<���s���쉝.곇5#�Gi��X4��
�_��\�?�JBF�O����%&-�qy� >~h�V��5A8~�xӇ�T���%!�ޛnp(�u�5�c��w� �q����{�Q�C��M�X��~�.6��1!EA�M<�}�kU�2�~a��K I����uDKT_6B�C�7��^����;��}�=k�����zK��r�Ĉ�os��/��'�y�6CS:�K��f�a}��k�S��Y1<�2uF�+��������׭C���س��|��U.�׿� �n&�@��y،o�Q�뫽�+u�Y���F����XY!*t<˺�C`�#:�Y��e{E���=��F��]F
�'E9Obߎ�o�<��=M�;MW�Ѭ(��M�E$8e���6�`VC,��8i@� `�3oDܓ$���&@M5xW����-���W�n�ri��RM���G��Z���e���.��&��1��1Kq[�������,%���a���e���"�_M�<�с��nάGlx���p�� zP�_�eh��*<�C�p����!�c3��keis��W-����������+J�O�ȷUP_A4����Fa�A\�D\ENq1�8���T��1���Li����8�a��,J��C+T��Cq�vM0�qɶ`#�(�_���pf��#\�8��ۉ�h������Ɇ�ƙ#�U�3g�ݶ�7a��V i˱x��� ��N��)Z�Ñ�֘`"�0W���xV͕{�_�� �_�1Y�2�΅�&�|���9��G���rmr���go��ee�]�?�h�V�8�txпdo��N�?Ɉ��%u	�6�B��,��Xx_Sx�z��&�{�Ɠ^1���m��o�3Z��-���7�I�\p�jE���J��^�����*+��̱�,��

�Zk�3:-�^�jȥ�IYح-sl{蓎��kO��we��N��7�>F�������g_����1�?��P=�]�� "���j�dy�ҦF�@������~�7��J �2��
�nq���}�l��m@L�v��C��.���6v����3��A%8ke��w�����YNhbP���+Ȃ�2L����nR��¼[	ȳ��'DMga�@d��i0&x%�u�b��@
 �5i��%�7�[+hZ �g�!ң{�M��QT*W��=4��i1�t��/�-�J�Y���#
t�! 4�t�ލt��7G��Z� �E�:��e���t�+�7�Ղ�����V���x�v྇(L�;I(/9'Y*sst����W?��������k��0 �z_r�����l3�z��{Z	�;��[�j�v1@I��J���.�eP�ϣ��`��cu)�������bW�����I�����*;�.�1/(a�Y�;��{��%��d-���%��>��d��7փ&[���f�f��q3��#���h�q܄Av?D>��J�	��]&���"�Fu�ǵ+=|�ׂS�{oC&�El��.�`�+�j����с�Y~�)L	SRE�1<�N,Ў�q
k���_��p��sS�p�5�w����;GC�Dqu�|��H]��<ZA����]:hB�)��r^�xDP�9��,���ӿ-uc70}�ق��5�j����M�_,:�C^��SӨH@�p4�q���~t��b� ����3�FzV/��M��w��fp�f#$6uK5#숩5
��R<ܯ��h�>��X��>�:�*�� s���1F�p��)���/Ѳ�A)�/�d�"v('#�<��Mg��Ύd�����W}z��QG��ዉQ�6�z����L�o��0؉�8.��<J}�}��iZ|�d��Ņ������yeGƸ�Ñ��Z:�t�<+x��֤�v��<�!�E¬��q�f��I7�6r0_t���T`�Mz(���FEr`]�m�4���+��GP���O��Mu�I���>����E�g����7�<������>��56��ݦ�qJj�b9�Ai�h��p��r<�Fp*;��p� R�{��t����dm(0E��{��ݩ�]�>]���/�f6�����Y����]o4¶uArT��Qe���3�C~U�A5m��%��lD�/6�,�`��!��ᶽ�Ȕp��ݟ�#S�D��r�jͦX�	�$��ݾ
��e�[>Q�%����R��m�-���d��o5ѤA�2a"���$n؃�u���_䚭�<j|l'�@4g��eA��"%Ŵ�V[�D��y��&_R��`��J��e���U�ʽћ�dkb$Ef���:���/��bB���_֧����WIb\�N�Y�7����2��Kj�3�3�QI��[���)�K��RL,'SZ�y��R������Z�l;	�dg��?�c�3�Y��Z�!(j�c-�ے�|;[5!�N��9�h/��'x�!�N�Kѥ�l����2��/�my7kj���6^C���ƠD�ȞɌ��Xz��Q����J>x"�}�0_�<J�cLG�_�lqb���PlT9?/�iO.����ɂ������� ���E�y��%.��e�)�q��r{;T����x�?�K*���@��v�EN5�b����0�Fz����R�V�b1Q��K�Y�n�D��������g��1{MN���x�F�S1��SSo�	��j�T�O�ÔȨ��91��e	�x^
\
���@����8��b��G�(^���]���L�ÿg���Y-��k��˫�z`*�Fb�F�ټ2��mY�*2��[�(.�K��Gǯ������m}���Ņ���O���Q6� �o�[���5y���q�˒O�{�k������a�h�ׁS��A�D)�r��.�W�R���5�n���/+��r���Y�+�.�y����C?��
��l�Ǣ��]>�����7�8tL��(=M������֋��F4Q3��4W��wh�!'{�L��4�?�)~�Z������s0�l�q��͘���uPY�I�':?U��ޜ��  ��v��+��ꋦ:Hd���E���3�:�e���ei8@�%���@c'*�)���"����*��_���I [:t�C]��F�#���X|ь��B'՚ �{X�h�Y8�bFKɥ�S4wN�"͐9c���n�~�?LV�95LSv��KR`��u��`rw�A��=��~6�D�"�q��pɥP�-�NL�0�{<sN�iZg�0��6ʌ�|�w�F��p��V�%��g#ĵ	��_�.��t(y�o����U�m�#̉�D��u�u����n�Mg�h��ny�M����~J_h�;�#��d�1;�VWww��y���Ƚ4��F����."is>�ݧ]6'���.�$�O��~��j_PގvU���4?� ��51��#�6�L�t>�\:/Ѥ/�������׭XUi�$�+8�/�2�T=�FK�Yv�|�OF���[h�՛rV�ۀ/$o�Qd��;ISm�ھ\Z��ƴu}��T�<�4�Ȯ$�)�d�d�]t�LP�(�i?K
���26M�5�^��#�i4�Ÿ)��K�[6}.D̀\mͨ6Z3�,�����*F�5`��[�S�z����B�����m�O��G����+�%X-	U�&S���Y쁂��~ǣYǓe�
�6��h.Y�J��]L|u!$���F�S�N�V�۬k�z��%rZ�:L2
�oc,�8z��ێQ���>�~��`�Q�D�HF��"�Z��
��ŝ�q�_-z.�v�?<�-RGi��Llyu��Ѳ]�~�g��jA��1��ۦMR?��zd̓z�ć���"�F ����w�:J�J�w& w��
��S��[�ʚ�au|c��꘾kS����D���5�,����h7�<L��?:������^̩� !�Wh�TլZ*��,��I}��!HWg�^$`��{
�Z��k���.��cjb�� cl���=�j��%/�D�-}8��:c����f�7˲�/v��9�tH��{����dQiܭ��j��T.�� 4M(F��#�Fƣ�5)��I�Y��p�ؕŅ���g�e�:��	҃����	��5j]g:��KO���Rv���JGC,�msO�ĝ7�)����ΤM@2u�ä�c,ǉ5P����IH���e�i*�lG����h(��g6u�5=��HC-���1Y*Q�),�Ri�֐�5�w@iB��)-�,q3ڣ�>�A�������-�sL�� �5�آ�:�����	����"���@w<��Av�pR� �%�{S����y<A>E��5z�줶�pͥa�MlY0����f�� d։_d�K�<��~�7����T�=���P�Z���Mw����.�¹;��R�Qc�U$�67�?��pr�f���ŒZ��� Ǥ=g\�X��9ǳF��L���H�|�f8u�c~I�0���O�+�D�(m�h0�Ƚ�!nmn����}A.%

����+1����NE�(�������F9����u�����O?|&Ɂp�+do���>����Btd�B�_:���̣GJ,� ��`�)�+��g��f�Ԁ�!�%�hMQ ^ �~T��Qm.����	��_]h:�2=R���ic$ j-��y�A��U@��f(��~ۑ��$���<���?�����Y���/���X��$a��d	5&�-\+�Ҁ���#L⧹6y���{S[�Fq���`���Fh�} h zY��.JgUw @�\p,p�Vm�2c�(	5��Fg�v�e��<�8�Q�
B<����%���5���gN��cDBq=( D������z�@�<={�#��`�}^˺ܑ�B�=X��+�UD�k;N%�<z�kERZ�&�8�����`�"Bl�5��O�����ЯA@oG`wW|5��Ġ��
սuvBd�F��xr>zg%z2]��sAe�HKC2�L�ȧ���F6['��~���	vzӽ�k��3ֆ'U�"��}��|?���&�1U����9ލS�;�d�_yDIa*
����e��9C�8�#  �K�Ą!��?s���!���z��|^���5��ΰUQ�������.n��rUh�5VßK�d��oܪ��s¬�2����曊��(b?����� 4����%�[�V��8���-��d�Ng
�!%�,�}�U�L���0���t๶H_zo��/d���%:�RB3|��I�,8�9x������Jm���Na��W��h��fȘ�y�Y�ٹH&��r�OM���r,��ʀ�a��!��:"���lT�zP����)ɻ����_ �$�˒6f�����-�o��g/�	|c��$�4"���S���lߖxY�k�qћ��N�2爠��J!8O� ������U��L+A���t�DQܬȸڞgҍ�Ґ����+J�-��������eML�2k��8�}4N��������#�>ܤ�﻽4�X���[$�@%�v"V�:2��%c'F�&�)�-;Y��`6�U�5��@|FGO�|��HT�S�\�:�Ho ΃���!)v`��]���q����f��+i=v�Oe�]^�X��A���w�U�:�7��鎗�����7b:�-n���Ѩb�XM�P��M�(����|$��ծ�j�^nv��bC�aR�@��Gv����*�̓�8_:)�6�I?q\_�9>>��|�yDs�\A�v�صy�m�05r[g3	ʊ'���"ge��8������r��[x� :�l���Q� ��7�(�2�(���}�u��Ŝ�Vo[9��ޤ������W��q��j$�+Ό�z>�1���� �Z������[�r�D��'�)�6����=�V�C��q���i^�E?7�.���d�_],.�]�A1����TcOO���)ȗ²��E9�ʀ����<x���y(,_�'P%4��+�B�!v�d�U���Y7�����R7CF�1�"��W� P���u�bz�z�s HK��u�ܩ�g����Mn���S�r��ī�x\㬣l	*V��?_L�(��AuMgؑ�#)�	9����lⅻ���柛8ƽm{̦,*�P�4���n�@�d-�D��~7��\�����}m�Vz�6a��|k��8_ݞ;���:HTq!�m���K�"��Ox�xz��
W&�WU%DS>��A6�~%�`�m�H,�'��G?��!�o�r<���æS[�(��FZ4��폋*u�``������Lb�s�C�{������5�d��%��|Ԕ����Ru��͎�؆}�/�\�0��rݟ��X�l��	��,�=���Pk(j��'D����ԱΊ�uQ沓�7f0�̽6ۓ� ��H�{�$Y �]��?���C#��a�ߒ9��yY�i�q�9 ����U5FH�����ܭ*�1�ޒ�m0����t)�Ҷ��rR�A'|8;:�b�
H�H���sk�A�3�{a�f3?�Χ1QXO���iþ`i�줜��_Z��Gǔe�П�&�����\�.�i�,0IL&�a����b��r�W��"�����EC��pX��s%�⤗��t�Ҙ>��Ԅ!�4�>ds�TD3��]����/5|*L�:yI�;�����[h�p
��I��\��;e�둁-d��[�46z Ήb���{�_Lo�a�D��|�լ