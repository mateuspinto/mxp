`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
laYJEQzVApU1I1BbvoIR/Ee8Avm009TtAlkCm+lquPXlIprm+X+A9v9Un6R/umGTHLjUkvloZZ+u
jYZVgeEaqwtnSXO39m2+ScYB4VCrD061o+aMZ91RrEylKoxih29kPUtBDE7gJZLxODgUoHYQvscm
umN8DCEM9d6mwIh2TURkosIO+q4JAjQehiuDGTfGwETytP2HipjcHdYRLc7ge+EK6QSPsV97iKGl
AwC4x700PHi4jtOt8MK+9NuIXAk0Mdmuz5gnn3qh1AV2E0IlnJOwQOxjlfVY53e3hVmrLsOnUPY0
GJPi88FTTH+XnEXQ1stopVYrKiPAD4Fila+KcGVjGIw8rmkfIm9moWtbRNfckr6LLHHgc9Cpl9zc
09ZUBpL5Q16AqEF76adg/ocqd9anSG2385yzCTeQvC18bPuSRb9PHPkFB7ZXYEdljRmz7bPwpyUU
Bl03S5NrdNfUplW9+CQTGmZJCn2YQWc0T00JjvhoGM6dvq1nKwARmI0arDoIqi+H4zRr3ktX4RI/
HY+rcyxOVR6wMcAEEpkxQ/ie4luQ5IQ7KvPbUX6KMdX1rmw0PAHAjycLrrLP76yCIQCkQVghnd2C
jFsVWXf9FuSCRSGLU57LvtxwrnkDnVXN6RbKlvHJ/oU478gphxmbK3rTq+ICTJKHPUX97KiVEsRh
5p7Q1FczCootUb1Nx0kuV200rozM8iuH+5WlyuJ3exlrnpQv1lT8MK4k8rJwcxESGp5sfooeWYYh
5mAhsoNs7YhOc63gkOAc6BM7gv84ZQKAmvNfAFkID7R+LigQQE/0P0mo2ixiT1yKaPRLj3MVhqR4
OmtxdDDzMwdv7mEkJexwAyKyBB6Bqv6ww0xRVdFvXHPiZAWIA2b/FUwXBPVFpG6RYLMgIpy4rphw
lEqv/08uwgc+QMb3Wjrad7eez7zGl1cWs4JqrTsW/RbvyzP8EiUmSQnSbU0t4uvsYstvSeNYjhJA
VqF0mPV5Fy8QWjl4Bi+zVhhyjse95RkbCGxDNGwliu3V/42eTNkEYFf6YmjoTxnWQ8v+lfQsAbDV
9d+QOJcbngXdTsaZyfe7camt135I9o/CpjLR5Wj5KTbetv4Dsj6u00N3KUOml0vNdJmbYi7NsAqh
taXtC+PHv6K4KrGHJHd2dw2O19rcypkSgCGtPy2zcOtFElI+d0V+1kcIYBr25tajLoSBenSB9k+K
uxg/SKFnoRl7OKtcLThucLKLsSIDysqT50GvyydgLhdL+uCyhF2IykIZVJMlzHLudMVjHAOOxFAn
WFJYSsqP22bIHG7KvCRoHMiMH3WPSJPp8CfYOjLMz5GaGcYFlVLq5MPu5c0JEENZ1ddkIcFuN2+v
yIvjYhACBU1zl93iMqMFBQqSl+NywTGs3c1oM39Wf8aI0Dmj44m64o2NHgyg6LhHIxBjUB+aXvlp
HG8pFQ2FS8ql9iUPo1EedNGS19uv5sPaOH8iejniWabs0CkfmNgKUoA41DVtq20p1hxz7bTChiZc
mgXvh+N81iv6pgpjcQ/2oHgpn1F+n9oOLzahBC5QAFHQX8cibAPWtap8fi1zvwkj4V6/GlE6JswA
EkOr4Runmhm0/YKByjeWDM/9CyXni4zpD0Cc3Ek87qaaK5/kkrTCzmUteThrKxiLDsoOKFmWEf4n
tJ6z85OkUqrL3n9XrHRjrhVUw6r4zFPOCdDiZAcmG2aZl5TsybQInItzEgnpWPpKMWn2Kc/GPZ5n
CXboXRhHCB/XyFlWJw4O+NTrI6XQmlkMlm1vyot1YVxit8Ls7KW2DYFxE5RLMZyL130icpwCeWr+
TXi8ZJ6dDVYyptah8JSL11UpwLi2wsu0tJA2ntR4uj7oMpPz4ZaO47SRdvzf7av6ll9eyWujsTFN
tdB3O3APTr/S26Or9yZOW+KD1hFQoeu15aNmpsvwhHXd7SP5AqZXFS6zF65sP6aqJXNlGhwD8iaL
DryQwFyockWgk2wLKarZOZ2Uy+SzSkeqyRfZHuJW93EqEYeRYJq/3pygKy9mx89+h9DeCUKIKJHq
vstYrAUu27Akiw9BXGw+P/2MpARNhx1sr9gaOVGUz6evotaDfY+AuFixHdTfsYdTw6v1HYKx/A8M
ZqoViFiba3jZGn/3SulSZcaIpEWZe2LNc6QB+Jh+2m6C5oo7nKasb5tgpJY3a4RkjB8oe6zysOrt
6fydF9+ilOW6iTDW2SskJUtSl7vvKBKhIkUAQY/PGlT1jcSfZt30tGoKP87oJz+qy4Z2s7KIQ67b
nOBXiNjJtL1fYf0IvVrD00B0jAw8YoAky8KppQet5H5UDOTSHm4lea1jL+O0atyBNmaSqgiwin4s
GCTi0qp1clHijK/8ybwGemRUVYI9U0GBjejwbiU+FNPveQYKYWiZNf3rvdRKY6gEb4PLdFskyGnQ
t3zO2cENKR0uYNjy+aSiaK+zIHzF0eFqUj2btad1zrYln+5YXhxRV8YC7qukxAWOtLZuXBE2Ob95
1wc4O/gHXGmJv8UsNeyhUhYzTJyyqaPtR308i62HYWt9G6Y/Y/IpJwMZCQjNYO6Mb/R9WUdrgn8v
o6f4mmv9O2ygonVadu/BtS6gpNVuOs1Nxct/9103evCuj5QGVV82gxxDEo+8a2ktaufq4VpdjY6q
DTJYaZ8cmhIg206kqODLM9fQXFcinFOWm59O3yM1aho9jkreyVw9ZoFYib5SrGTxj4Z6rHqyJJ32
fYv1o2llT/tAFH+yU3aR8RDYXC5V7Ko7e2f3Y5tLr625Wt+H9G/ikLVjR23Moo2cQz89xHZcUowe
YEtsSbvnHQEXv2ZVp0ioZtWpN8OPyU8oXwL2LsmRnI/C/30ub3k6EI1sDGR3hmFxIQurEKXonIxJ
CiQxExXEy2w6/sfJCa+MeYBpWSt6ZdGgpAKeWMbPz6T+0TmQhuHmFSvHsONhV0VaVg9GKkbI/M7v
QdThQ2W9wtH1cSjfOqw3jxmWc0W8JnxU25QqyeH3kvsnILRsXbK9MLYXMSQNE/C2I5wMZCJvdysz
vfRVCZrj/8Jk5pOlCrEqwsNiSGh04ZppltRbrr27hZixs8HJ8US6ashUtn3hcp8AHywI3fTn0CAy
nxkh09d8OD4tFBiRnfnBvmIqyBBPzf6x7aI+GBJsUgasa5XyWihVRiqqGHi6ZPy4XGuI2EDaS8cm
iY0EQTdI112U6vyYWshysB6g2NcoVPp4FbGk1LAtH2JRkVSJZ8KhsAXjLyyU8F7HXAkXG5Zm0UMa
Nx9Sc/Xg1c3PGS4NwxDNWf3eiio7PrM9lVRcbr/6iaHk4D3aIzZ3ESEubtuqeFhV/jqVODGFDJim
uoiPPqkV4bwgaT4RBjCfjVUId8Is/v4/eLKQXcl4Rp4m7ONkdJqZlik7BP3IBPwS/zPnTUTu6T14
K7NZeDTNP7D1oF5YcYn+Qn096zZ9uPRYoAalFJ/OP+o0cbD8UH2VkwQm88tYY/sRvJ9ix2G+Qfny
XBgWX52lkVdzfWxUt5/VaT4OgOAEYRKZv1CvlVsOG5iZUNEKIjloXCh6w0aenSwpftavcjwhbPAo
A3EryMQK0GTtv5wVjwRTqXzzP+T2y1aAFABW/XLeD2jHQSyO5WtfDKAycLU0RJV5ZE50wv5gYtOX
7Hh0TSKyFZw1LkResBtJTJgZXYa+o1u6dKpLOr6wspm/1ybqnisE6ffJV6skDnEpEGqG0qNB2YRX
k1S72dISx9a5d931iD8WxWmKqzXGtxaBzAdDftwgwk2nVOGbCHln0Aulg+wXZbysmW2Di4o6clmX
99zkPU8SgyHfDUUo5orOzlMMvWEsgULZjZ/lWxmfLfhUbT+mCqAqRhE1e4+aCD4hM+IvPMWOTqOg
UqG/PBfetpLu07Gn9uvSrf9PigO2wQzAMLZt8U6siI/qFxtbdSz6m5xxVVkJFIjpT74cxGbN9T7U
MuQ2qKrGQPkk8lwtopfkKDAc6IB51AEPyOxkLmMHiDp4r0nIhIUyzp5mqyEXfKfZGyAEi0GtRuUl
5KTUjeo28pgQD7dwQaWJH5I/UXA9cizpqLfR63y0OVn8JV9p3r+pKv6mzllR6OFIv8VW7pTWd2bi
yOhXMk+HNqYcfNsHN8ObJBytAIiBcsm3qYYYBRu3E/vkff2gydRnhTJUUAKO0/+ahEl14fdPeTGX
8lMU4tllQRpDFX4+5/YYyVNBK5GSc8hq8Sm+HBpgfkPiHQWCzfyO0+GDfVAuclq/vtBi2h0loLyZ
o3my7j136oB2meyvLmzoBAs6fyGv4eBNhLjbU1/5G+BwkBanAbX2SwuRTIHimG9tp9/TP9gtoXjY
FPiL+HtYaeQA4chmKaT7nUD+n5mclaTZUHlgVhmq1dQ8KmiSXvdca5YvTZ2Kh5gQIJYXztbdlXqi
ipJjMduXwx3zJCEEDudUTb6z8YT6pgpc9akFZ3AQyiSYH4vynQk1k+hkTTPKHoi74uC/jeEqbTDd
djiscTHzHsUXYpSXMl6rs6p4BQvhjyrBFq60+3pvEj1GV85Aiqjt3733p7qv593o2PZJkXU4iQDi
hhhiXXANmB+aScuZG/yKsyITgaq8khAIIU3KSbxBKcXxwYTyvJc02I1T+A94w5IbUa+EcdV59qe/
VC5GLMwMwv2UjvE=
`protect end_protected
