`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
onV3bF7qKhy57atXsUew1DqWd8awvqS7uSv1egpZtWt3anXEXhzS/1H/RV+9X5xJ/aGmSWVlYmpi
ivwjk9F2x8ldbwyFr0Y8I3tA01KVZE70oS14yNNdHMVRYWKSkdXNQdP3ZuwYtHa4Cm9lgTLYwpxx
THfUuL9ISXwp74vSxM8ViQNJzgsRvbiOFK6y1FKhwyQ3y3ch+tJXnnOj5jHilICfOG6xb83mZzs7
G3fsf2KonKiLl7e4ccKXXkQJsokXcgKnmPUIukshGd0177NDewqaNM9znXva+zFGnGFnROfUrGnC
CgArASGmGaWUgECvA9hv7LXbEZ+3+9Hml82FI/1XeDf/mT/Djq8WfzD/DGJSGGamj32FoABW7byf
ihu/HkVUbLktKufgk1pjH089Ph5bHFD+BtVOk3UhtJMaQeZk7fnjDzO+mGWFPXgtsarD3EmR57W1
90K3nX4pIu/hphu3su1+gDdI0tTyWyxsMH6DYWqWqK4sTWBvcseCwez0AiTvwHULzIwbiFpp/xZT
EN3x4PhsU+aDX0o9ivozf3sS7gZEOffmE2v3u5Y41uADXHXhLh92BLrAxjGZFGCMbtxZ8XlTgbV4
1DmCwi4xxsiOZaUEF1ckFFz7S/HvUuxpbQhLxi9yKLBB0KzwW7n7ENVq67PpIEV7pHK1Kr3wfkgv
qJZieJYYteuSTPnIDGOjzOvRANmXGkIHOrq8B6BD5ksiRMtCzoTcVdIzRnJZbLBZJvNeEza+d1os
50fHxRRXxxrz5yM5Wc65HPz8NDsPlRI6ikolBjwEDZWhpGEX13yNXUg6CbFir7U0AO705DPtafhT
fnKzZI+ZxTRWYn+sFIgTniohLJ5KUB9kudVNFBqvyHQ3HwNeVMIVwYT1JBAeNEIN5lWcZS76s83h
fjPnDrhzEWPl6sWrhlCdyGkuDjvrF0HMh/rOeY1EmJbT0oHeNdwAERI5nfXv9Y+cPZX+xxq4bf1c
aL+GH+FwV1bLKAYT+xBt6j88ci5zJDHhaZjK7kUD/Ai4etIG4BQM2DIkLAVyKoqXhPp0N94LQado
EME5blTheKRF7jUhjqN/F05X24jDswhpJ1sg80qKcsAGMhLsjrdRLE82xErQMUSg38OPD7GkgmOI
kMlLTft3+qlG0ftElxWNkKk+sdRebpP8ejTofq7cvwtTyxO5b9Kjk9xNyVZyIL/cE4hFOLnbKIM5
2+ejd+cHL68mQYER01f29KlvfVXkhgAZUL0KzZ8wck8WkvS+E+v1KUYbVlD6YjU0em+xG4/SmLQP
750it8RTk+yHvATsCbCkTOyUIoBO+Fa03iaU+NHEJ2j8QTKCX5b+8uRI9IqIyFVI8zbcshRiGjq+
XNGjbXeXJ56yXyXERhIuO4BiQ7XyjGE0UJy9T/nknv4ovUKyU7jdjg8GYdmGmwiXt0B0mG1bGGeh
6zG9Zrg7qQHPoYRE66lClR7SOFg9cx8UFXLg+N/tDxNuvw17vk4wC7ec2SBqSFO1Cqex3WEO6OmL
YwLSplIjCVpQeLD5tc1Zbv6cRDaxJWEm086zwJ0wxPzdFGzLGdkeeE6cIz+C6dPrnPK69ViH9QHO
IZ3LqOziEk+YO1PjIYeJ5ymBUkbslVHYiAuj5hRyhVmOtvO8T08pBsqL+Kj+UGvWceyh73nB3G1v
b3wZi8hGhLwAsPHLDg9DmNKitfALhzLf6mnYA/sZce14TVywp4z3piFs+/yuM+ckd18WYEZgF+3+
imjB/62ZVfSP5TjFaDzG0+7FeRVjlyuQhRffBa7BzKkg+akUtWnRiKX/q2+XPQs1iXIjv2vY1jmi
RZKHaRyt0gnwIY75IzPLsW7FndawA2cCW6LFBRkWQL1tTbTV8mSyWfG4M8ENqubztpsf4RpaCke4
tAVbCcXteYD7DzRy9HRRg6XCk7qBZYAyKibjfD2Vhs575yYIVMPmcJ1m86v6XEFVDQTjYU+whC3W
5/2BsmNdXwCRiEbn0zpCOJ0eQ36bhvYGvlYvF/ak9wL6Utb93Zq1TvdDoEdYFnMDh+pTNbMfmrrR
Uh9Oq2CBVpbG1NcOlZcxKq6s8LjqPpvG4vtSeH+CsYjy1JhnMOX9bgcTcBLV2g0AdmmKN21h8esj
cn0w+VZ9bw4LoK5dXxw8RluqKRVE65apJqFshRncF5ApOVwiI997DK6518ZvlmZNNicgn6M+bKSl
px/xBHRYiCdhxJt8JRvYpEz7GIiT08LSHuagB+V2JVeN4fgxL0sXxRVv+64v9dHGS7UTrp02Acfh
6/IVH056MIvVMZWhiTBf41Kk0sUyBJpPgmjT1TWVhvVuLPPL0Fc4bauhiMPCyLzwrT4lSsBtJ8/A
EyJXKU2YzmK37+TbDQZw7uemaiBz2/dE1Kqi8rYuvF02Rg0YrgOMxH1CizhHqS0SQCWVYdenimkz
Jaspv2yxlYwvoqvGHWKUJOV2IPr6FtKMWHJ6gjHgpcXsDGL79oW49tcnTRlxW3nlNd07GUgEeSLW
BnOwT04PC9Nv1oof/56DzBRNdCYo4wujnTwLhsb0mADRiMVwQ6TyMr8NJXvtkVlNF6JIlx2+CPEY
SbQv2MkqjYdaKJ0d7s+EkYj/fBkkJM5usQrWtyWukxhCN1b0CrWBPxl6S2fCL8nFGlIyVUEOJi4a
ZV+rWfaRjuqRQbFHifzJ+07mM0u+owEdAarUZmxXGTEZIq1DtW/TEvLfYdQS3FS/JjfcsRGjU8lY
aC6DptypOcZzcTR0xCEC9a5sLPC9mcejGQPdkHbtzkWypFBSsuyTGMFeIcGLs/GPh+iw+UTXKql2
lK2LHDGxifgNXs0NAyPzVbIusu0EylO5ZUmG3UlMLANFD7tjpM+rt9iCBiukIfjE1Md45DnQKgrC
unPI8vHxKIc2vhZeDRSpzx4+LIb8la+vn/gn4zZaju1uCo2Y931klQ0Ke2B2NGH1vFaW6VdNUYF0
YyP7J/Qk6ENhh8AQihUnO+Z7LquYA2bskfvvSs+2dqCUG5JwVFnjWxcvD17MEUJN/01r8Lx7P74p
ahRv6wT4s/+wtrnH8Mr2QJR5+wTFr1s2R8GDZoQ1whsYoYEOU4ieSH+V0o8dyZfbkL5WZh22dbQV
xQIa/nc/t9aGh6xNJOC6QU4MX2kz04RH8DL9wRB/kw==
`protect end_protected
