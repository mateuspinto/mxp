`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
XYOBtYIdOulzvLOtDjjJ+r9q3EjDgUNttydAqaq8UH/iDxyHd7SCLl51/4fou7ecnFHRBKnrACVP
smI+rcdJy3greNDLI+dNqHximDv2UHR6u2f2Mb9uedZ5QYKPYc+b3R3h35gaQlpSgVMiru4wg8VF
eHnjPva9xTJfPx75O8pWi2jGSMl1yERFzFcBsLCYVplZFS9Ih8opFCU8BrZsRjNsC+8oj2lceMAl
R7b68Z3u4WyW15qPA+A0FD5HbwRHE7WQCo47+RoSeh/QIknFovwarIgONzjyxJHUyjZMpqSN0XaL
6ezvla5SbsoZbkf/NFphPP6n6ypZJhwhvwrkrwueATT1c6JS9VRaM8KPbubIVyAXvfBh3rKcoU12
YibttqpZK8eKMdn1ir/uboJQNqkRC8MaDxvQbpavti3b6MjmKIMmAiRT86F0KNsRLO0xhuQa68de
J75Nfd/04Pu4Z96KSVoPWWf/PBfoaoNAxeyOCk/DmXOe6zfE2x8q9AH+ncTqiXQN53NmMQU+srC0
2DjjQE2xwyZbaj5wJ73kTklsRjzEeVaZdhUPEztZADaeZu63dvJSSRY+afd6Pna3Y+mLUbR2gy2v
rz5K3aSHJ7ZHtfyzS+LsMeYJ0S0466egV2bZZrX5swxtS+fr0EWwA2Az0U/tFnVYUYYlIuAphWjE
ufkc7gQxo/i6Vh1wfnk6+zFrj1i18B4q7n2dnpSLAuxxeuW5QPJunaBxQRWS07701EE+o6rqv0cL
dTF2GYAIOkyf5v6NlpXfY8l+xUxvALh7Dd6pJiHzPRcsfdrHE7PQ3OvJHMLYVNITd4g6NfhFgjMn
bWWPQrHqr3SZlzF2p9Ugh648TXssmPKj+23qHyJosFeNtIIJxjwoL6+pudQV+rVvquRzsL8vJaSL
6+3Irg+WGs6n50Wre0cHt5VprH48rnoP0bzykKuhkjFgtmfE7C41t10qKDCsFjyLdMa9mKXEMaRE
iY6fBk4TrRAWw9zGldqDFxwWLiDbrJmR3p+TcI488U/QWj+6pvLl402Z64isP1/PbLnrWyXRVJBd
MyrbKL6D/RP+xgMa2nYnqGICOc5SmyaoDqrkWWKPGi5coELpfIuly0OgBLmxV+6yqOk8iplnlFLc
Rf25dyLom4FkEGEEVGhzgFnloWTD7dRLEfQt/9Wt/dZbE2S28w/iJMNNZR5qq/RBiMWLBz19arQV
JWW7WHIsj1Y5pDHLp2GmsK4sxvaioG6RYhGF54OLrmGOs05CD9jwXKRmmm19PR7jaqK5h0kbgZ2c
qe1xwio2z8ig3li4HPJjQM8E1cK0TJoGu+WMg3tD2KwH7qQRPurV8Gyb6VXWg+i10bl2HDHuwFt2
zR6OQucTxl0xikW8hbpOMZ0oJc9f+Ap1ndEEMasfdP1SNzGtGI6MABTIh8aSMs7LahaX1Otw3j9U
xg99XJh3l5MCZUcAVOjDJXcuRLq270jq8MSFg6itfZX3tSczOlhVOI6rDPs1v29RYszMwheg8KgM
Oaurz5uzW35Lsnp3kwZSQ3+54CQh5QiGjuFASCa/FbvADOiZI5wPdC77fcSVwKX3LBwlgdHWY4OE
jfMW2eFKseiQH0Dw61ap5R3Iv/fkbiofSns3D+F2l26dlXCOBT+w5efx4VpWwEgiTuXyROPgicPB
Bxd3qfgnAVIKEt4eK2moOwXcu8QKprt8S/xQ9VL9ECSoTYmwIJfQNn2aDO6u4PFJCm+JETNwr8yW
Jk7rocQvVDadmQaH4jqPqeTYjdms//JiGRw1bKdqxMPgJyQTkIC36eDqpmIUjSoPpwBk2HDuQ5ny
CfkF3d1f8JdG4rOHBWa1y/a7lZRJixDi1Ybno7dlFfZsR2GNwsMPcPSZFVmPdgqEca6aZtPOrM2g
GtXx0VgYJkqflSPXBhkQ0O7jXuJIPhQko9vB2Ourg6nZlbE9Txm9zGd5wq6pLYKB0QMXtVZEw6hS
B5amwHQV0t/jlzjCz5XA5A4jskBRYgL3WjlJodZbREKbHLvfrWrZmHI+opHENH9xqS+/z3V2kDgK
fotuPL9JBm6fuYbp+PWM0Kr+6OHny6oqnNiFrjuDQ0l1cjLmi5CvAa34DWwj
`protect end_protected
