XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Au�	V����K�V?#�c�� �C"�̏�,�d�:���YH�2��VV8*~�:��)�) ��pH������}ᣁ4��v�$����dX���Eh�ٻ���)	
(7�������A�1��G��@�xG�U����|��s^�ȸ���Y+�':/�Y��՞���W{Ѷ�$X� d��X�Nsk+�C�K,�9W�(DнZqO?u��O��Z�P�?c9�f5��F{˕���5�L�aU��{>��r�[&��	k�G���7�C��N�����	�;<�9��'Ϙ��X18(M���nHe:E�Hk �j��I�	t��u$+�K��_�F`vaP��6��(UOؘS�#I$W Ǖ��2&Qb�P[�z^���}�C�5y��`���v*;�ޅ�����ffS����p���{.�f7I^�Gߖ�@HMeWvv���J�`�����L`^%4�s�dy��G(��?l&�By���mn��
��U�T���]ag�x�3���|N�][>1����fka���ϟ���L��q���\X�?S�'������<��[��N~@)�Z�Io�ɘ�9L������=�ovD�r�M4E0�q��\nA�K���o�� �o���j�N"���Z7X�q�zl3���T0+�~CT�m��j��> �dV��~�_>�HL���lf�m�~VXb/a}A�`(�j��0Ǖ�]a���~+��+��[�)���1o��eΤ&�t�,�=E�n���� ��jXlxVHYEB     400     190Ś�k%xe����p�~?C�c�=*OY�x�jK�����<�&��U�y�&VԔa�*؏1�iH�R	�/��v���8gbKfk\w�'��6|f@��	���1\/�6h���b�� ��5�Ό}�Md�B��W
1�y�{����#��ʂϟ�HR2Ş���`}?��#V��#Q A��:����h	�'�t��p��.�f�J54�xP.]P�2իv��3�/kXlᲔ�E�6Z�k
��������!y�؆&��;Q$Λ���U�c{�)�S���?ߟ���#{�$�yrN1a���)�i�?.�"4�^��8�vxd�J4�#�JH��f3�.���) ����j��1BH�uhZoנ@�}�Vޠ?��M���XlxVHYEB     400     1f0�%5�?�G�ɫC;?u�<:Ur���'0���0�K?V(�b���8`G6m-�B�a^'ޏ��s������Rٖ���Vs�T�hw>�.�~��s�X�$,��e�q?��Dw,V���|���¥�F�	���(@�r-�;�������vH��̿-HS)a �=����M@g~v��@� feX�+ֵvd��.ڼ�y6թy��e���YKXn�w�p�i�R��]���x����CU�VHF:�^��O��v �]�밿�h�x�·��18�Yҷ0��H0'?�*5�7�E�pv�(���ַD��kc� .M�h�6Inf˪'��u�.���w*�4g����+��C)=�inr��CJg�?`EI~{]�x:�B���y�{
�����v0�[��V��sG3bqX��� ���͟�u<�+:� �y�WR/~�^\]�{��fX�yrwt��w��N�"�ݟ:�U�qr�!XlxVHYEB     400     200��;�K!*ܷ�I���W��s3K�.V��zk�%���Ҳ*�%�LJ+�[������m��C��L~�y]�O�/%�}+���'羺�=���bP�OMJ��&�P��,87O���tI����%�,�e!�;Kd�4� �1��Ǽ���+��l����5o�G��uWoH�iO��Z���c@ش�α^��)�G�����H]�����w�i���PXG|_A�ς�g�)��Ou��ѻ��ֱ�c�ԝ�O��4�-͋�L�*��hdb%����)t�ER$�N�s� ��������$��#���l��n��0�S)�_�� ���=�NSQ>V�G��m�?�ybt����*^P�:����7��$�!��V�q���z��%lni�Vp�*�<�tL�	���I{�'��@ ~pWN>�5!5��Q����ak��qҭ�)z3wk)SS�Ue�߱rCZ	���}iJ��nòܞ�xm���7�%ҝ"弭̒ޚ��%v��>����XlxVHYEB     197      f0�aB\���.~�^��"=����_޷1��\�T_yີQ���S��rH���[��է� �0��E�ϐ��-VO}W����DY��U��_�Q�q�">Ow�ތ��껛yf�0�(�ؙ=�Ӡy��KO��D<W�%i�V��L�;��XK Y��g^�)_*Ј	�)b���D�~C~�$��8v̤���d�TdD7����l��X�CC_��\s{Z5��g����