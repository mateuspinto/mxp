XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"O����zOC��N�eps��G����y�/Յ�fA˼�Sߡ���F^y5U���]�*���)N���V��^�Nb|Q�d[H�e�:�(�$	.����,7��uT��`l��&�'���O��M��ߓ�6����t��ر�DxQ���=ShMB��=咵���j�s��z}�1H	�DC�d$R���7��V��Nf���w?��W�
x˞�J�܄` ��E�GG�|M*��ճ#_#�j�Շ��4����"�C��A�^2��"�nd\u�%Eq�����/�����Y�+ٟ�4� $L�ym"�5c���dD=UI2��}�a%.�d[�H�N�������q���2U;��f'8�ҏ�����?pLx8���%���.�.|80�G�����ǚao���Ϳ��fz�J����2 ���|Q/Y�v�q$Ef1�?�}Y����a4�eCY}�?u5@�m;P�_���
T�H�!�6��Pi$�HW[<��_rٸ�{Vث�a���'��9�MK�3۫�8P�je������s��=g��-��\��_�lWzA¥0z#wSZК���P���|��P̙nY�J�*���T��� .�̄�jJKg��_aJ[�1M}1���B%�tZ�s�����l�_K�c���}�6`�x�Q�ok�T��p��y�D��}P�'W���2R���v[�Uh�X埴V�^�eN�
#l��[�j�'�����.b�nƴ �f�=B-����� u� U���;69>�XlxVHYEB     400     1c0��RX�j��X�]�u-���j�+�q����ٰ��A"9?Y�F�{�+���.'�O�`��hl>em���"0��	�oZf����y��U��i��eY��'ގ��a.��C�iRzl�ג��!��	�'<\9�RB<آN�1~q���mA������;�Й��:e��K�Ԅ�$V�mP4;$%�,^6�KbLcs9��V�A!���a�̦i�DјUI��b���!�W(�ޯ%HW�G����n��9���]���Ҽ�,��b�*���h�889���Ȝ�%{�y_��Qϒ�`͐�<�}�Qm�jw�Р��WE];�ŗ���%?߲�hR�lb�T4�NY�	�;s�o�5�ϡYWf`��	�["D�
�vX���uK�c�І!��PZ�.X��"��BqZ�5C+B�q�/G�JAI|-��Ʃ2�\n�jXlxVHYEB     212      d0�z��X���TJQs��bV�L)��\1�͙��Uv.aoS�ހ���� -�`a����C��U�Z�0�3-�xw1�x�&]ʌ�^H��z��WD<��*u��)���,C�qX�2QQ�L��{L�o�ϝ�����[�oap��'^FrR)�+h���#�g>�j�����j�85�"��{��#I&i����)�
������ M\4