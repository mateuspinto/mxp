��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���챲-Ȱ?Z�_���N�^�J��6�Wgǅu�9�Ճ.y�����)xi���楊>�����H҈!y��b�G���c��sP��@���g(�Pܹ�o1���5ЦS��(�d4�'��톎ydfƜ�/Ϋt�pӦ�之��������1���*�K�Q ����P��d%@��m�dV��or�B*l�Q����duht��X���WI�[���+��sz��;��2	n�]����>�^��`)�IM��X�=�b-F������U��혅<���S�p@h������.��� �h1�?#LC����x�[��{�~�;<lx�2��FFy�����i}-+Ux��NԽu|3����3���� ���%����C)�x%W�ǩ?��>/��,p@f���&�j�[�f>��_�r�����	�F��6FCҲ�c[-GF�P�T�.�lLt�<Q#��-8?UR7EU�J��A����Zn;��x'�G����F�>��5N���Vm���*6���-���{ToA�m#�m�(?�1�Xx�uM��{���$q�J�ʭP�	��J���*n��G��Q�n׾� *��8\
����㞲f�d�v��0��C&È�B�	�ʈ6P=�_��P����]�I:197���:�A����Vɽ�~v�jNU��X��o����a��c���y�ey�΀����|�0�X� �+C�OU��ْΧ�CTs4��^�%Z�sc7�>��+vϜ�K}�l�lQk툖d�#�F���ɵ'�E]<0h{�2�O�(�mh�G�7.�����U؇��y��
D�H��IY�3����p���a�����}��=��ie��Æ���g��m�Ʒ3���"H�S�p��z�[@��i�_*�7=
�|<�b�O!�^��_��"o;«Pҡ���c2���\"A��Gl�=�S�l�eR烲E5�;�����a[/���m��,Nb�Tw�(? =Y�	\���9Pt\ub,g�I]���%��-�q�4�q[�e��i��3U<�:=p��CI��� ����u|��e�y@%�=˘b�0���˥�VSIؠ��ɴÎ�45_�%�P*9�Q�l֫ޡ{���/�'�7�t�KKw]�s޽^�U��.]^��0�3�x�
��j����Hq!Z��Kh���}r�����QE'��.SAq��
(�E:E�[i.tV����W0�#��a�ά_gYy��P���qh���n����O�FM~:�O�3�U���v<}翎24~�y��ٍ^%�q�m���5�xG�t�^�-񝘣�LT�[NjsW��E@��	��5�b5@��hP2��f����V���ե���t5��WƮA��=�z���㢚۬>���Gvp��9��y���Fn�6MIw�x�5i�{���UK���5j�FN=��6P���慘�#���q�=bq�54m�[G�&�H��;�h��yoF��!=����#ޜjD�|.���('�r����f���
�4��9r�A�%�E��'ms% mW܎�Ӷk�mof̂�[���L�q\8��lW����!`��>�?7��@�m�������nl��Ԡ�iVP���^%��Rr��LE P��ؗK-6��j��*H[��:�e"#�˽0�M�E��g���Whd{��K#�VfK�A��p>���,#�F���p6ޱ/l9���e��F���>͎;	�Gj�f�'g&���v֯�Կ�V�ǂ�*&D=��E].����b��AF�Ӥ�a���^�]�I�[lI)~�.����&��A.����3u�3϶yү�P�Ya�9ل�&Z=�L��mN8?X�3��Ģ��/,��qS�چ�^_97b<i���x�	��	�����{��a�@�up?��Wwib����.C��� ˯��#�31xԺ=��f�V
![��4���KA��Z?��6�X��A�8z�y���R<�_�ɮЃ�v����FP'���[�!��Q�K�sD�[�xQ[������A[��|l�9-əv�ei����ـɺ��7�F����O�ڸN���1�D#kK�qk��F�,�V)�Ɣ\S�3�:�P(+*=ߔI�L�an� �$���镦C?�?�l�DѦ/2I/��5��YT��l�d!���2w�_3�0�]��h��u��Ck�fO�˷�?���Y��@�H�ۍ�{E��	m�#p��M��s���æT�ba�n�I�9��K�����v4�>�y��X�"��SL!���2���'����(әR�K�{>�C^��+�wLX��{2�;�'�xA�`G����<�� �:-�X�6"W'�8��!St$������X���.�������wF�T�q�/���'[�&�=�c(F��+�6��q�Cjd\BZ�ev�z���ԍs��9��.�b���#}9�1*���7�S�22�ے�C�1M$��R��%�e���ƞ�N�Hi�.��e�G�Z#hM*~tcf�Ay}�bf^]R�,l��V��;}�0e���$?�ؖ���Qd��f����f��
��ʂ��#v��e���$�*q��������.H5{�?f�|��sD�	������+B���'$L��;Zyw�h�8�x�^�ŉ�'�-�\2�jI�,,uQ�E|C����uc�x�C@E��捉��u�Q!i�
28�ʔ):��b ���qY@���4:���������x�R}�G,���� ����0�r����'\O�$��d�o���I��#��d��'�F����M�7�C�P�6.M�jK`�+���Z���q����\f��Jv�3�xV*�:���'���{V�F�F��n�j�W��G����b����<{��'-E�zw�w-#��kkq��Z.��K�+6�N/��]T}n���Ʊ<V_���Qy �G��1�)݈W���$J�u����4W�Co�q�$�%��)�ܛ��p��9���9�xL������y�3އ.*z��ն��H�8�G�v�YyT@�s_R��>�؛�3�U�o�����e�G�@j����6@Z������'j�:��/�͌=�9�Zܥz\��n �N�k�ɖȕ�Z6 w�
����\/��V�+���,3�9W�[�29|]����W��N~��v�j '�ʫ��惊,��M�sӻVf�D߱t�����p�e҄ig%9��}5���.�o�_��TB:�9[��Vʮ�C1a*w�eN� t� kY�1�}��d�gd���GL3��:��Dv���a���	��Ѥ�o���4��@EԔ��B�/%���2�F�W=ڢ	�Ӏ- z60Y^��͎��dKq���0j�e1	V�*�-����Z����K�����}��IMݹ�n�is�]�L�?���u&�B��:��?M͂ J��?�U�
�B�8M��[ػ f	)F*�?6��w:=�E�4�#������/�:<�HWjP�g�Q(�92ɿ�wB*�����?䆼�j�,qQ#�av�&ЁaT{`VX�0��g���9���2E/��3��X��FœZ.�Ξǥyr���c�N��n\��Lw�%���ڎ���2��@E�|�1�z��ϼ�{X������ՄC���	���l����PW��{-x���`]�6���9?�&NSFO���qXt��x������j�e��5���I�/\�����W� 9��aA�Ė�d1�"���l8��ʘ���.d £���� ��a �=�z�ӧ��/�+P��)���p#����7r���m�_�ģl�?�f���I��E̜]s�Woea���ky�*�V�C���Z��F�X�,����ԎS��_�<�ݤe�ILx�T�v�g,�Nb����0��w��!��K�v��[��x��߷Jd�!�����$�1Dړ�eӉ;��ᙆ�����89�z��zrp��j&J��v(�P��|��2��kV�/$ل��s���w�����+ڡw����9K���8<̿�8W�Sc%&�E^v��Ǜ���Y���F�9�D�����++�/y�M�ղ
w�������tߩ���oy��+~�c������r�B�F�9&�k�iWDyW�c��:��M��q�Ͳzj�i�����9d1�ϖ�,f��wCQ ����@�1�d 	���[-��gs�ګ2[���R*��:J�,���h�$���	�Y!�4!��������*!�m�6�L��.��Y�p���fY����~��|���νn�ӦÍ[�1Qۣb�bC.Q{��4�b��+�C���j߲�����g�n��Ax>X�
t�*�ǘr2��J�4���4'$���"�OW{��P�m�6�kJ�a�}�JMewl�X��#����gWa��R��1)~�`�l⧪1����{�J���`�� ��ϲ�2$f�n/p7��}�/ο=��G_g&���nօ�g:�.3�
`��ki���;��?�#��YB����k������Y�����`˫�\�n>��onvl'��v22gݷ����~�r��9&M�@^]w�6�cY��f21.lz���z�� ��T啱&���']����O��j7�cT��un�����Y3���v^�K!\h�����荒M��4`�Hƍ�t��G�p)O��A7l�>�+�2������^N~
�5��ږ�51����0��eY�L�@�k+�'�~m����1�Ͱ`A�&��ɮ�1h����+-��n�/���� ���U���0V1��5I��B�#$�q?0l�<��e��+�A_����F�G�5p���;�wXG;�Ǝ{�me{-��U�{~���	�<�t& ����� �m	
�x���#Ɨ��e�BI�����`��Ɣ��W�p�>�R�4��j��P1d��n�Sh�J��TVjm��=�s��@�����R��og��/��a0�p��s��$:�L���	�4$�C�%�ݐ�-p_� �>��[�ɜ�ٲ����; :����u@�R�ʣ��#	Խz�Q�>χ"&Jqi�l�l�#h�dg�%���b��z��ŭ���Ʃ2� iM����T�n?3e�?~���F���QP���T�Z�*�@�����&�rs�3����?�qi��X �����aFY��<�N�"f�4�%ԽR5�af[�j0�p��A��X�\k#�Ð�=zc })2��O�.�Ea���2�Ig�OU�w�`������L�$�(�X*��	>>�ȶ�;#d Fe�-?��A����.x�_��WBk��7��x����m�Y�^���c��u�ۓW.h�����}�4��37L\H&��nC�-xCT�)�n4ӌ�������,�~��:N�BH�X���N�9t�i�xv�6��1c�d�Z,'��z@�'B����i���L���uF�,ton���oB�V�,��'�=�z+����GE�"{�Y�T���u�K�P �
3%��S>,i�]�/6{!M3�-��d���;��Ϭ_��p, �s�T�%�xK�)����+y�N��Z
���0�e�O���A�l*�+\��z�g��N�H���9ݖh?���tk8�;��B��OK��^M�XA����;�Pf�_�aO��������`����ʪ�o�G�>$������:��u�8sEϖ%�A��dt���;n<��	R*#Q�:��Z�`��(��uj@>ˀ�L]ܻ�<̌�����މ0(�R�#��$�� ���c�8�**,�9C�3��;E7b0Sn~\�bB��p�!�@A�:F��~1��[�J&�*�3o��G���T[d�b휓Zf-���V�!��ɽHO"���g z&H��,6�ҡ	��/�h�[+a0�B"��n���}i��HS�er�3��1Q��J<|
�2��۵��J������~��Ւ�N�#t"�Nsx���ys��g�)cd�5����)}��.f��c�6뤰\�Z�11>��~�(�W�Ɏ��pr��83���G�V�'k �������AG�/,�@'{��9��߶�a����N�7�C��$$쯉�l
��3q��u���b+;E"`��kk󹫓��T�HP��c>�����9`Vy�M�t�@�
N^"R��!��{o5��28���h�ҮPe���I��8�c>i��)J^�0�z�7��w�8�����tJ���B$6ﮏ��X�~:E�[v0����x��D�����qM�\��t�fM<���~{<OClj�fX���Wm~��|_6c�ߣ|�PՂ8dCH��t������fk���g8���U4�$y�/���g$љ3��9�T����h��?�mnX��{�.���+c�~�e^�͗xsN���N�-
��������5v4�,I�hBc =)t$���Lŝ[g���[����GB�U+@�Qf�x�-v$ҧ+s�|$�iBG����~��(\*�Y�M�?(˚U��2��{X� �!E�N
����\�'?v�)�����uU`�}_B��<D�s{�c���o�9?����&���HBŖ�&[7��-I�[J0%�6���Zl�6g���7_Sv�(_
'�(*���`󰴘ݴ#łm2�j~u���&�C)��OR�A*r��&fB�&$�"��8��Ч��}/���%�3����t�@�)^G���>{@���#RR����~n6�D�`|����@r|�R[\�7Ƶ��c}b���T�g��:7o|���ː�ê�Ϋ#�KZ���
�К�l��(�:Y�f�Q�� �l-Z{��2���9t�K��a�	�ҵ�~��H��6��H�;
�ao���
���$� &{D����O�|$���U�wS�2@��@���1Ҥ�cd}���b�J�(�(�S��������-�~�/t̛�C�K!�C��5�"��y�coFd�wj\�C6�����3*B`�ųPn7-&��ʈ5�.���p���dM��|c��6��]��P	w��wtK?���O ���XD���R�)�q|�Q\�nGe$����f�<�a��}$�ʺ���	��+{��tK���������";!�N��[
����� ��^%`�sڍ�9��-�Vg�o:v+����!H��j0):�O٩�V��aGc7 ��d��\+��r#M{B�
��� C}����!(��(0?�Ayӄs����Ezd��"���=�u��f������&H3���JOmW�Ӟ��G��Q1=�3:�,cSIj�>0�S�<�m��v�#�(5�}�E	w�#���i�������ǚ�B�<�D\o��.m�r<��-N���������Ծ�� X�t�&1T�r�i)
d�I�4׆���{����*�]L�����(>��P_�C��ť�d]�%���-��w8ޱ�S#q����Sllr���e����^���=)ļ8���Y%H�8�q.3TC<�TX-�`���ۨ��ROv.�G�b0E��T,�Q_�c)���Ll�#i�x���i1r)���cB5��!{��Uǀ�L���=ZHXI����t)앓?(�⿲cB����}r�5���NZR+IC��PWD�&���
��yD����v��3�V��T�f��$�&���#gQZ����W���T��4}B�Wb�`E!n{�͸m��D{4^ �Y:�8�AJ��ag�����vi���!���r� z�0k"�v9���i�������b2��x��$�����W�^�"U�@H���0�����bP��KX��x���Ұ�|�������5�fcu*Dc�a�ɚ8K��Q��|Mc"Z��7�9,�
O��!=v~��;T�i몺j�J�7Gir]pu	;��3��R�?rm�A��Q&>���<�'�>`�x\]ag�M*Zb�r�J�z�h��]{Atn#����7O��%|C�JG�Lm���1�5��f@[{b$33�3a*�Xy�'C�l#�� 6ۆ�B�2�����9�^��̔]�ͻYVF!�:����p��оA���6}A&OW^Fm����t�Ӊ�ԯ��0�
uȼ�X�)eih�m:;�y��Ƅ��/����a�[���%L��v@+�n����ی9/O�㥣h�ء�:�6�u	�<ˀ�P�(�L#L͞\]�=��P�q,`c�	�PDDaꫨ�̚$�d`�5���Q�A���,�l�ScgP��VTIч�S�.ơ� ��g��b��V�~�\޸)���G���u���ds�K�xz��d�\xZ�����̠V-���0Ҟ�o���4N��@A�]������0��������J�˪2�:>�}PL0��Qq�4�����fLST������d�̅���|VHԑ r��O2����B��}�'hBSӗ���3� ֠0.ȸ[I�`�̜ʟ-���ޣEY$�ah5�Q+'�u%3�
��K/7y��&����B�ł �'�v����Wb���:N�'c�(�(��.������t��35�	Ӗ�Ӭ��|ٜ���^��3}W�ŸQ�������7H��#nj'䣴^����wv	«+���𧤝��[XG<������L��Cs������kc�e%9^�A,����R�L2��_�����l#�zgUo��P�i�!���3�uhA]`��`p/� �YCh�6�ܳgI�u�)�y@�%�����B� ���m*�:�Z4SN;u���^�����5Շ����=�YiP1bD�+m�h�yM�9��P3<��l�H��"H�mgG�
4$=��R��Tb`��n%�mz��Њў�y��ѶU��c4�a�3�x���+�6���b�,�U����CMJѬ��Dm�H�@x����#�@V7��1:e{����9U��#��($z�e���G�׵�4p2�-��!|6iD��λ3�Ъ/����Nn�;K���g���������j[�y������>�5=?t��,��n��Xr�Ǘ�eF���*mDa~����3��g��PP넒Uôk�2i`{Nl0�E����=s��(w��+�����#4�@��N�ɏ���F��ɾ	�$�װ�}��`Z0{�aH����}.���~����EAS���"�Z1�"^�аH������-Y�v4�o���-4|E��
�l^� �F�?��И�ܥ�~�A�J�/3,&�H�uO�
TE����oS��o��x%��2>���Q�\��ӓ�7nu���-F��T�B^u�r�ZR3�'#q�f�L����<Z�!�������\