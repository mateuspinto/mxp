XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����w�̔=��։�脘��i7��C��E�T�M�G�f�g+c��U��6�w�Ҭ� �i'ie�,�9z9�Ak�:5���w�HO`2�Eŭ(!��,�������'?�M2�l�&>:gS��uI�g��ZV��B��f/6�K�I���4�;U�K!NˎA�cB:S��g��	�i�p������c[7�h&1�̍�7W�����va�9��,|�)Q�Ŧ�9�c�5�oRf���"H���c��Wv�i�`!�T�R-�S��L���C4��Q��a(coI���	�p������}��շW[�<g�����1�%l��������=�	�AC�\"��ƶ(�~��h�����nKBKc��Ry�=1��HQ�-1`���⎶{����>�%�b�G�*f������aM�$ g��Ͽ��(Mvt���+K������O{ֿ�Oz��æ���O�k��o���lJ�[������#���8�w^F�%(�)�|�M'kHf�Y�g���Z"f�����mV�O�֦.�k�.���#%E$�?ع��0�MK\|q8�;�w ñ��4�Z=R		$�1�L�DA+:�G�e䧜�8�l��V�5�Vƻ���а�4�<��荷���⁵#njF�B��4Mx���v�ǟY��V��4p��m�]0y��EvCj(n��Ϝ�uE�(T�e]�xw���bV�.�9&v����G�N�J��f	Z�nɒcj��x�6ٕ��D��Y�@:����K�5hkXlxVHYEB     400     1a06D}Ó-Ԋp0�N��d�m�b8uz�E�����.+��|;_-K-�V�<��lG>�%V�Kc���9Ӻ'��w(�+}���k�B��fRR��O.�[ȣџ���������&�䋊%xIf��g_���&�.�܂xs�����^�T�7Wq� ��]-�1Y�|��R��~���:�l}朩� @Am�ޙ�E*�&�q��/��53��6�r��rk��m�ղ��&�t��t����B�O��>	 :���6Jo� !�����A��h�@�$�vil���p�{5g&Oɐ���f�ט���A�u.>Q��h��yIK�#!Ԋ���Ȱ�Y��V�BF��'����q��[K���1��'7P}X)|g&m,�euգ'a�(���a��Ѕ�=yGP��ϥM(�xT�չXlxVHYEB     400     1b0�ш���'7V;�J�1b�hvf�=_v�&���L��Z6'��M�����`����|=�z�0-ﱝS\�'/_�W�h%ֲ5�mA��n�V���@QB���Jx�j�����m�]�Ϛ(��n�Ĭ��Q�������Y]3���</,TT$v��/�֪�yu�-������o[D9�ߣ��!�Ex�!V�T{1f��ŗ$Q_���Q�p�+�N����E9�<�-&�:ש��+\���1k~�D�e,v��"��gՉ�v��`�<2�y�O◒�

�����`�����Q�x�}^�ߢ�m����lm c�3l�Cxſu��x�c�I�SCΊ�Z�q3�D�qmG�/�M�5�<���U�Y#+HE�-�܇&~g =,��Z;�a���<t۷1����rN��l�7�p��kKRqkj�쏨XlxVHYEB     3f5     130�
^ꓬ�%�=���U���g�����,��U���,ޞ�*��}c�ᢣ~*�	:Ys�OU噤'#�6��R�paD���-s��n��0&EB�u^���'�eˉ��/ܭ��=*������t��ӨR,خC���Z���D/�։�!YIĲU~|���(�Yg=�I7���	��a3{l�{�0<'�B��+�"���X���ۯb6P�����KU�.F�\,Ȯ���y��w��ٿ�;��԰6�e�9��_g�C�Dt�Y�7C.N"6�};֣>a9/�@