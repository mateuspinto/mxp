XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?,��b�b�\R��1�ݿ�'����� ��c1�O��j"�#u�I��ZP#�?
b�����Fm��R"�7��u�p��u�\1k�͏���Ui������C�����)VͷT��6���Ш���Iq��|��۱)t�|=�*��n�ʌƵ�
�|��uE�]iX��X���2��c"���%>϶T����,�H@`�O�>ɓB9��ó:��=�V���M̓8�J/2pZZWV������=������MHJmꝽ%ΡC���Z_�"�����H{<�ҭ~\L �|9�:�������1->�cu
)9��SDE8f�I��b���^˱}����fg�&�9�Ȳ�*8��[��p��x��焮�J%=�"q����$��1����#�::�Nvf�+�3��]D`Ui��.8�3`�my�K���z�'��v

8e8�-�b��:����}�q�Զ}���
�e)��k�g%n��k�PG=����`���� �F�3	���{M4�c����e.F�v�NuI��v]���2�}ډV�UՂ��U;�Q��0�'�`��.-ƹ�!r�԰���vM�@�8�p���sФ�1ެS�6��O��Y2>ScUx��B[�u��.�U,LU
��/�g�$�c�F�X�FK�w�h�%4���ޚ�k���S�mtl]5��)�Ԝ�1d������:=�	7x�R~�^Z���g@��j�*V����]c�
:6j(���	��E3�m�F�l���Ͷ߬,��#XlxVHYEB     400     190�ᴊ`L�e���n虽ٚ���c����UIS�әB�|�Qr��Q0��yJ~2�!{4�Ss�U;�����_���<2�R��ٮ���� ��?uĝ�G!'X�0|���Ҡ��i����pG$>G.Z���/�$�0��	1������xP�/��� ��D�F&��r��x$�b%/�A2��� ��$�����?:o�������n�-۳�y���Oڽ����R���9i�v��ꇤšTo�����bP�L�oM�<	���;SQ�
��Q��h�K�&��Y�n'~���h�[O�Ɇ��u�
�fu�����-w~�="�(�R�dA"��?�u1O`���(=�$W�k1��$F����Y�1�3���n�E�`�/��G��>aXlxVHYEB     400     140���=k��,�O��OX'n��f�X�!��Va�]�n�.N�K}�9B&������XcT`<=��EV:��o��W�������R#ypB��o����q��6!�}�!6T�k�dE�?逰��q�^��ΐ ��(NwD;<8y0"@e��U��y��d�,��R�،8��+S��>��g*p>^���,��Y����{�| ��c������='�>z��NA��&i*sx�X_�&Ae����nO���@cxpP��$�h�0x��f6�:c}PzJ�怜AQP��)k���	��
���u���uc�F��}�/�az%�ZXlxVHYEB     400     130
�,���v&��8��LW�"���������87�J���D?F��1X$����-\��z��=F1镵�'�N1�Js��/(�8�B�	@�Z���"P��"�;�4yU�'�@�|��3WF@���x:8���w����}>6�k��v~7
���y5�j�@����t	�&��|n`��b����M
���:������)�7�q�:�������H�|�.Tƺ���T��ƥ����]?:AO�Tkq0O�P���{�q58^e��q~��0�� �L���Ow�I���f�lqn�R�f��$��XlxVHYEB     232     110���p��Smuԫg��Src�M�U�Z�;�aZ7����|���V�ĵ�w�(�\��9��;���7��$퍏�?qn7 ȱu�-�b���_u"S���� m9�!�a�$Ӂ��%�V}m�8):H�Z2k䜻��yE,狻���2�Q��rd���b�D�
�CJ0�(]!�Dt�����`����Y�؋#�\�9�pQG��dx�y_�$��y�`�d%�-�(�%ܵ1�U�����wÚ1��Kv>���