XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��CϠ���Wn��M�I7��q\s�q[�'��U�k���O��5�B`�����h�y:�pqU����|�@�h���f�T�R�.V��p��4<Ҭ�b�i�ؘ:Vϔ-��!E۱D��D������H4�S������Y��z��@�Q�k��'�p(��vp^���Wi��x<o8��^���4�����8�l�U���K�.���1]�iK��.���r�!�����)3@��-�m4J�Eܴ0���l�Y�FW�88%�07����N]�R���g������F�7[�e��dq�7ס�'��5�YP}6��G�]�H@���/hym2��D�S�0��S�ؖ%[3����e�I(�Qu�I��C�����g�ϸPؕ���O$9E���f�J�9���;��j����Χ�d�]�"�$T2�}S2�\�[�2�L"׵,O��{�����֟�p�d����!h�d�u%7���XS1]`t�@�N��׷ʄ����+��"�b�Ku� ٮ�2J
�Xi�(�Si_WĜrw'�!-�,猪�;m}�]��V�`Ū�������8�T�^߁mF��)��b*4�|�os};%q���8�UI�cx)�A�z\>�X6ץO�)�5����d�[��5���UPqRf����&��qU?A9��l����i(`�GD�4�L���)��m6s"g�Qݩ%��) �]��D�p����0��t����s����br���!0b��ED�䲿�!yXz�
����=d�;�k�cWXlxVHYEB     400     1d0A�s����H�FQ���R��)g�� 53	xD��S��8o����8��Bʝ��eNi*��Y�U��ʹ�����e����������x=5d	^Ю���i?��7��ħ��rb�qr�J
) 0�C�~�3��?[�W���%_���8)?��߱[��vٰ�q����r���`ٮ���A���ސ��1D�ƏD��׏�y�iB�.�B-�u�s�*��o�����|���.�@3W��9F��h�����uJ�j�$=��{��263���|xc��fz��}����-�}1G5O����q��{)�Y��,̴��t��e�����c� )�M�*BQ�����Q�4<8�O�j��;�DE&�q�g�Cݙ
=���%k�Y��<�.�o�ͧ�q��=
@� )���]��i�R�,�����'�Q��̀A2�z���t&) ���QĬ�ȧx+�Dh04XlxVHYEB     400     180��q-1C��-AC:c>r�|��S܅,-l���~TîvzaF�?K�����+l�R�ټKmX�[����$�R��s�Y@J�R$qZ{qw=��E��E��ԳK;��@i��k�������pqP��M�Fz���y&�s��[�Ʊ훚��C!�N\����ȍ�U�wb>��ZUtr��M~L�S[N f}"��OTC� ���[f�ǥ�$a/}O�O�P�$�UW��_�W�����jp���	�%�'(�kS3r7&r4鿺���uԤ'��*��}���jq�����QH����#�5Y�����y�^,ӏ-����7%�up�E6�<"Ű����l��"���a�;Մ��V�|�$XlxVHYEB     400     140��J˴�fN#����_0p����z	=�7�1�������{��L�4�2�8F��-c%/�w��5�ߨI��*����"�$b�hYR��>�������YpbH�U��X�t{�3��8��Ӧƍ��J4v[���g��F9i���'�o"RӨ���8W��`����<��|#�l&�x�C�J��B���ǒ����6�9W��Rֹ�]��g��ԩ�����T*���SJ����'������.ճ.}B�yr$/�i������*�ˑ�s�X�^������7���<o��}���[N�I�çx\Z;XlxVHYEB     400     110��}���AdC�9z9J�����!" ��e6x�sT��Xl݉��{�$5�U5�d~%�7�H�U#;�x���Į7״�em������>|����+��t�f�C��"�q��Ӿ�Nk
��n\�7��\�B���iA�L$w��&����ql�+=1 �J�q�QҐ4��=��XV^���4u�+˷R���/�_A
��"�\�y<&�� Q�GdnR��	��}�_р�+;ݮ�Sr?g���"�r4[�5d8�th�0zX}̦!J��TXlxVHYEB     400     130�����4<#���s]��c�b#0~ph��+�m�kX��k�x\㢶'~�;���Y�-����h!s`C�f�(=l#� ��P�,��/+��X�f���YX�3�&vdD2ɐt0�M�R+�gV�;�0��=�fjN:r�8~�`��Rą�@e�m!�og��_>�5[�ş���(O���mV�JG�֛}��=��k���K��9��T�.������;D�BY??��@GQ�_�7@�_�������B�v�W4�ɯ`i��Q�|������"Sf@���lzxwP�d��۸䌀�XlxVHYEB     400     150���/R�����&�*��Z�%>[B�e��E��w"\�G��RR�3����D�_}��9	a��?L?qy���1=鴁�I���i*����S{��P��9�9Ƈm���rAQ��ԟ�ۣ�� }`	�T��I���3ra�Kn�u�)Л"k1�/p�J�<t��2���W!���LD��-����>��6�4�0�8���`b�ü��U؜c�d�V|Y,�{Yʶ�`��|>�ĠP��F���j0}����4]�@���Y��1��rI�Y���c�|s��=܎<��#&��lU�H0b�mm�n�ܙ�KBja��(?�[.wX3ϼS������LXlxVHYEB     400     100�%x�M�s&ry	�E,�~�͢h)=fe�"��%�%/�o�2ߴ��i����5c*Q��ߐE��ᾭXZ���i\�{���@�м�ᶵ�8�W�vA��[�²T�#2�6��;W�o�3�)��w�u�B�2E�b<`��ȍ�jͥ�GG\�g]��޼G��}���D�R]�Q�\	V�<=�)�Lb1��Ҽ��$���{������a-�x��+;�����<M�rU�;G]�G�+x΋��ao��UXlxVHYEB     400     1c0�w��-�7��u@��y����O�"�֪A�qej	7���&��0%G`��P�JG�O!��ǹ�L+p�=)]c8����2yL�ת����g��D���g�Fs��A�x,��Y�.6�+i��8��3�U?F����I��4�p��|� �={Ym#���b��+X�D|"�NeW��Y	W�x&6l�yG�{,�6Y:�� )dh)�ګ�ߡ���ֈ�&߃�6�`P��`�E��Vv��\8p�(����PfՄ��]�Y`wW\�&do�f��3�k�����^���!6W��PZ�8k�ò�������#c,=3ġͮ��B�5�VJ#�c9����I���2�@؂�<������G3=F@���0�āU���s�e�Ft(���p�*B�(���|�X��ۚ&���+������2p�|�@o`�+۱XlxVHYEB     400     140m>��+հ�X�k��z�lԸ���?#E��D�=^�؊�H�
���#|�wrOj�.��1j^���Iy頣耽���Yi����3���k�@�l/�MJ��pr�k��*�<Vd�&%�%�6�s������wﮞ;z�<6t�LT�v��kk��Y	o��@sR����.��~T��e1���o��)�_]�G�I�_i��N4��ЕT�ǣikaĶE��(j�kK/)��͹�#M��&������{�I�����)�<�$m������f���*	2k��#QH�}~VG�V�����M�/H쀓5Ca20[c
��� ĭU	XlxVHYEB     400     1a0LG .�V{��\�����m�Bo/�)�+-aT:i&Q�o�43�c��m>�)�1��sk ��(�g������_�cv.<\�`��yg*m��3����UlU���ѽc/�=�?���5PYt����_y�����l^A-�3�A�H4ڔ���Qa<��=�]W�T4��cp�g�[��*�m_��Ⱦ}�,�-��"�:h��g�9g�oV^;6��t�󈹸����y#��d�[Յ�ӏ�_��<}bl�����7qmz�P9]�"��="�sڶg��B���W(�%��U�G��z�ZI��N��wa��_�@�e�*>�W4mt�t8*q����7��c+�u�OC?���'��Vk3(�c?��[hMd)5 )�n��RY���SYw<T��,�v��>�|W"{�T���Z�XlxVHYEB     400     190��@"�>L4�]!N��X�|��4P�]�E�p�G�� f�]�!^�c	�ca&�8��]�	N�|�%vMk�>[���}�>����?�R���تFH�L��^�x����ՙ�h�U��9s+�qp����#]b¼yk8_��5ǰ���W�R��1��-�U1�(��!G��Y�_ �GD�1ʙ��A5Gf9����c������V=��N�3)�6�\�'&9f]�w!�6��Y��������a䝢��R�5h�A��0��;|��.������έ��w�q��S�Z�hm)�0�x�
��	�њVܒ*	�H쎧������LhD�|_���[n�^���%�K�@I;l���h��K#p37��z���p���"ݥ(^���tm��Hf��o�49�KXlxVHYEB     400     1f0��i�6 �p�C��:�]]��qfǒ�[<���>��iD0C���yQ�D7���A�bY���N��5ܥY,C��))��p9}��Y��^4d~/�՝Ǵ�"������9t2�H�����W`�q���<��څg��Ͱ�t�U����t�]�r��,�:5��g���$~ʐ�!��	�96ݡ�e�Pn}'� �������y� JN8p�����CR��?!��.��1���B��1' {�j� B��'s�5$2k�y��P
5I�&�F��7�a�1|�n�f��e�c�I�*|
wu[�#�3ɾ=�ɋ�X��k��օ�[�e�W�Οex��b�� �]�Fƥ�	G퇐��A�J>i+�o D��� 	u!'�j��ݧr�Z�)V���{���v!ì�S'(��z��vKG���r�xV-=��� W��+�:��Q��i�����6��6�)�HY8����H3�R	�fZ�y-2�9�i�i幁l�XlxVHYEB     400     170š�U�����S�M��0<X�{4�WYN�W���_�iI���ʘcș�MH�{�è �!��{���5m�O�����
(�7�A��B�p@u� �dL:fϤ����Nv�C�f�d|���U�-�bǘK��jx�׮�������m�F��
>�W�s@���nN.c-�ci���(�X2[\�b��w���h�M��Gԅ�52L[��Lի�z���:�` ����R
٥�)f#�x�4��x\�J��u(�]�4�e��S�������0ݪD��`�����R�\��*f�8`�z���@g�,��ǒ�ؓ~������2_&L�/���!�C��ʴ�D�d "J0$���s��D��1��Z�XlxVHYEB     400     190;���ǩh:�jV�Չ �QȉĒ�cCۼ�$��﹐f�4S
�@�λL@8�*�ŕ�Г�iA*8�j���+�zdꠓ��=���z2��@t�	Yvi�h�;�D��9]ֽ��!7�#ޝ�Y��n��	�Z�e��C�
��Ҽ�֗�)Da�#Oֲ�(7B���o1_a�#R�y�� ^�%�W@��"���WCi���̿(�P��W��_75���Q�oaW�C�yI@z���a��t���6fx��i'������1C8�����k�5z��L��ce���k;:������-���~�;�TƸl�	l��A�Gї���oq��,.&�Pٺb��QО���,�@8��o��r�Vԍ`��@�G^�M�':u!f6K3�T@X��v�~��UXlxVHYEB     1fc      d0���o��0K�qR�t<�1�8�� .�f�ks>�[}C�G-_����=�-��iZ�.N7 ��P$t��џ�ZD��{�b!Kc����E hA57	�������H�w7�1r�kd��M�@���#����v	t<���ri�F���0.�,G�=��D��P/ ��2��D�A�:����}wd%�s���I?m D�53��C�Tь��1���C