`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
fIuyD5LqTKJwWu/0kfEx8HOVNxFzJS2nDcwsMo5Xy8y1RXOHYD2gkLGJrpX9+KMsS6MokxC7illg
avhd0FZ5EEAQvYg3GYInDqkC2mMFkmykIHXsWzrzmCA4q2qzWPLgbLM1tPkVlkenQma22Ge/MlY5
5OQdxkuAfNoZRoLiXU3XzEPF3gBmIduKYsuDgdspu5UwP6NTa4brn7aYgpiDcbwD87OvMI4Xb5e3
3lby3BfrHoZkfMzqTPwIwru8auMSiMnQOz8DWyzVOajk/S4qTV9o5FKRVHue7WZQlYbS/j2K46MS
A+gIc77JS2HOM5UpVmtC63sRJFUdoQCkU2Q7gA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="bejlSWKAcuXve1g05GmSQ4OIDGBnmcK+IYa5Zsu0lLQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
wpQZDe0C+uWCu1PcFM801EggZgrFTc+037TfBzvkK70Aobww661GuBmzPf4QxePULPWSRsWAMDUW
NCuhLFDqnCtvizMfbf6Hvhx82VBGhzDt2TVsO2C+Bj+TWeGrPSq1F0ZB0xoWvCtZHtk2Jkm0z8C2
QREL3QiNjYMW+cIrvxlU/l+T99STektfB8N2RmYBtzwIb87ZSDhVxAEVF1PDkxuulDm619T1CsM5
adEZ6Hc42UzxYNOs9lx4YnG3VJtWB/Ns96X2lff2KbGWbrhmblmsN9oSs+G8MrkqFrALaTmVS0Y2
+5QjRRe5bOdKeIH2tIesHfC5/Lq98lyWJT/8ODjr8QKIFJYsJX4cbDURC47NfQHO7p7+vzUV8U/t
90S0fIptAlYvotKNg0v25QhPcliVvFPK5jeW7N3upCoSKr2IvnpbqCaZbCA4SG6cUrm4p+UDZ/yV
JsrezqEA4xaEWGNCVeX7+0oHXrxj1E+q6TjgaWBlzn4L0VLjNzbSDoTkkmoOXDfwtmEg0CsBR/Zj
CErzFUfMgbMHT7kDxI61xkjkcwA54A7iEyeWA6weWygdaDFd+xBMyA6d0iiapDn4EQm70suBZB+f
3iRF9mInxGLFPRxD9IBNzfar0R8rSjnrZDh4S8xOSEYRnYPnT9BNzEwKJBcBkjq12fLWUXyDS7Ta
sNyqbEoahnrWLYpsl2CywDth2uD+tR9xLUugJEYDZL3nNoV1zEvi9MqRe9qioesOAl8Y+b/CZL09
Q3YKxXQZIYMarK2i2q7jkeEQpehbjiCOqjDFEBsOzKTe0uIWuck2ecnebVmbK0Q30/OxxKLVsjSh
xE9b3hZzHzs7sNLip5T5mSo9fGeB1lx+kQUpWGdSKaZsZQWH0fjbKL0euxxK8CRkb2260GiVSltq
i5Ils2t5DK0lK5SOLflekZZerzAfCNq4o5Y6ap9LOiqdvElfvDZSW8GMEh4hvG88cLkXltvvky6L
ZDalFyelN/yJFbdTg7MmPFGQTLJI+PSetaler82PCeAMoZrOt5Q2+DeKkC+BG85c6MciocAbnDhW
qE+LRS39MxnN74otq6dTyFNZHSS85twERen32nQdCKIEcBkPlFr74Iuo69zbih0sh7luTWMjde3u
JkVLST81SFAQYjgSLUwYgsHQTqle3tIumeSN4fPqV/n7KXUWRWJ1+BlCY8Jf4IGFi1ojoQhIT39o
bvWIAiBn358juxYBnjNjNSPkQNvU/AlGfG1Wrh3tz560XX6+wTm6d/HgZKAzXv4dj1bOd8nwJ3hz
BOY65dlU8qP8XJbBwtDTdAolzpuBmPHGAABYljNFsKhKjKHDxmF8FyR0uSYCuiHx0Iy3RB12jolj
w5JP2Omdmie4rbn1dFzSpr2+nrI60PfXqWL4445gERVymtxxEHpWF5mIBkj0RxNq5gCEs4CyvvhB
bHnG9MsnR9ha433Y+Zvo0QUv6ZaZ2US/3pbn76R8ajpvETfZ13aHqNEzV5iZLg/9WxGawkr+UXLl
MJMeLOHAj+yYDYa6CZOKl+tPNs/DC2kbWfdpFW2cqi4eTV5r63t8E++Pl9Hw7sdlko5w7lAcF7JY
FVxB1dXzPEbBsamS7fqMEcNuVNP6sQJpUma19GR04pHPjWmj7w6z2urDCDfsgGKXBmSklfoY7z9S
3SANDbThFfcRx8OR0hf5hleiny+0gCRnfTupI2+y0XQVO1BeeqAaamkc3/a+4/A9B2DaPFG3P+pr
RfhwQGhkKfondnnfAoS6FeRBxcX4yzvSivxaJmpw1hnitdfjM81om+rNpWeIXMkAEVkUO2t2LMdM
/gWgyRhO1a9nVO8IseVoxsPhaGGpQgXfbNF+1mxjcR8DXzJYAf8Ps1aLzwRn8BWnFPqAyIgLop1C
0Gb3xUMoHhiQ9XgHm1QwTw29upQqqvv6V2szlvnvBSgQNlGyTTqpN1CApnAVm/yun4IrkzLkOCG0
HHMCDWuChfpxav3Pps7qYDU6ne/lPLQUfNWV91C2QKmoDvT3al3RE5G5ZwFMJz/Wojzghh1r2dom
nMcsY2RKFOJwJ3OBEKdhFlds2JxKEz4w8AvS93ABvsCY8tTTfZOMORJBaK2N6vHicrAehFgQQuPO
r+d8FgvH2WKJ+5NZMO2jkrJIHaMZCyKNGsu220o12tJIGtvpwy0WbgWifW/kIWLluvAKuaiHz0dS
TZjNLmdBBNrvt1tUBKu5gT2bPpKDpPOuLfsT8VE096LscpHAfdMEEyWmrpVrkeOOR2j9YxtAaQqr
/mfKxEySZAlTj7Jexv2G8o5a+v9aPc2kUsOQ5vbX2s83mruF5hhj6uMD9jxCwXJ+JabuGhKAScVz
/6GJQ4KqN8eocuwMGi7wirRG7UfzySCPIthG97qF4coD+jM90F6sUtx3DbLUOqIadVz8VBb6LggR
LJAck/sKd9MytbaBQB5mkYnAkudoY/IkuYd5GO3mwjNeyAGCcKaKHV5F2vA6AevjfYX36n75HIt4
p92zCJ/N8Tb3qZHXxOJN6zHpfagPwTc460WeP8OfgHkHBurDDAjmdgFz5pmmWM4cPrsV4wRTCZ+w
sLK3gGuHd6N8HDP8p3b9CwFvFYSqhs+JXWahiPDi803aHUiT0AQBE9b7ADmQ1GsA0yEcuNxbJk6x
nQM5fs1387HAZYjEpnOI1YPaPxLHbBhDDQ3fzaVpmY7EntNzP9QgxSRrdY1Kq2/NJVjcxVzxxI6c
nxC5XHycSqz79U0DJStuLOFJ0+T4coyL9pGv14a40+QHcigfyNuRJRFDDasZQB8Rk2XUAZLn943d
YJqw9+0+wG9IoA0apFkCP6N6uhaAm4z3Ioh+btJFJ8PmVr9n6/g8oxnXm24AQFbuhj3SJG00OfGz
6Ttxyvndzvm0RGZQvCSB0iHn9cMzk2AJQo64U7a8eYRxk9e/pCwrpyEd0UNfWdo9BI3/pl7eLjwo
c2eBvl8Dir6b+DjbJ/m1FfSKd93omwXeo674MlfXpdTV9X0ma9P8gN892vnbdtNVyeOEFWejFQSU
a0JFpqwCmxJbXlIzb4AB2y3cY/Zab/a4pM9RESo81DwobJOGqsdimhN8GGlSk++pJja/+ubIL5za
KE8S+RjCWTgeRn6tue5QNVKu6ZGwBj6hh7OAHV0owQ==
`protect end_protected
