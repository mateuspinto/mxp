XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����#���j��$�xu UW�X�B�3u�(����6~g�T��t�����4@��f7��]��)�NM��
�.��lD	qɔu�e����T$J��Ƭ+�l�F���`M�w����ƼC0��nOa����xv��,YS�{d� ��׋�Y7��H�MB�*]��@x&" �JIJ�]^oHs��v�ʷ=�\a0D�>a����
�R%ǲ�o*���օn�H�~ *˂�85-�ź3U$���?r�6�Ɲ�?uS҈((z߮�y.vM�p$��\`܍�����=�a�(��!&`��l�����2�~���[ތH�h�܁� h]�c�٣��U���l�q]���.o�ji4cȅ�mPU<$O�M��F�괟���H�y�5���t�^�@��
f�����hO 3��s�x�gD�jy��k1ͤhEF��i03h�+u��A�sw�r}�G��8K͟W=p-�=u���?�)A��&��4�EQ��}5��w��G�!)TY�-d�t�h�O[J$���P�� (��,��!�MSY"�$Z���S�ze�mZK8�<��7����d����m��>�5;V��zl���%ǀ"[�[Ҷu���(fT�VݴF��);`���\+��"��^z�hv�H3�*��8:E�kQ����>bB:Q/�L�?�w"|)7\D�ۂ�m��җ�°��
W�ɛ�
s'����&�Yc	�^!P�d��u��Bf�u.g�W�,5��XlxVHYEB     400     1d0d���S�#�?��� x�ij�������J6��<�񧈍�������*'gbǆtZ�����aab�$�	6�Īn��F��bj��5��4HE�L60?t���"��X�e<�"c���ĞAh}ġ���R���t��0�x�n̽�h*#�a��p0�\�`MYTI��� r�V`݋��ׁ�cB���<��s�=o6�AJ��x���q�p�bgT������_�BE?<����1-^q���|C�㵊Q|*�r��:{Jf�<�\]��]{z��Z����4��>�WZ0G����g�YL�}�7�]�=ť�ڵ���ػEx�}���K��c^�ԣ��"S�׌��2W�9��B^;��If?9�?N����
 �W"��$g��zI�91�a����=l���=*���j3!^�,��M\�����H�N�ר��0>�s��C�,XlxVHYEB     400     160�2^@�<�Ң�������ӼRj�ՑZ��6'���U/��9������M�/oR��Q�`�.)���&()�Y{�(M�3�j���m���&���m~�f�W<�v����u�c������;���+���m�]����J91���m򾴓�dk6�f��Or;D>`O���o_�A��`m�OPKs�2Ӝ�� 5(z��H;am����~O$��Ԏ�}j��x���Oј��CO�Ukf�}&�.u�4�����}���5�{aؗ�����T��a����yb�egB>P��ဟ�5����a./vrC����٥�T[�Cz,P����Zv�G���BXlxVHYEB     400     110���ת��t����G�^��:�a���Ɂ�C)a�3v�j}*x��0-E�`�Q���C?bx3�8J��b�J���Ug�܋F����-���:�H3�q�yhM���Zb�+���?}83�&O���3��y�>3< �n�]eA�e�Jp�G������t(-ڼbf�L)�è���{�X�IW���>�/�zڵ���M�}�Ƃ�]�3��q�V�n��`Az?����KŞW!b.����Qb��U�K�q�I�XlxVHYEB     400     110�����,,���5�D&_���~��ɞ,��`ΔH��}I��m8�jk���f�$�?Z��t|�qyT�:�?��%l�Ɨ����}b1�y�i�Tm��:8�t��_wH!���
���R����>#5ʉY�c�0�e��c����k�w�}���l�V�r� �r6�XO����j��oU���]�F��Ğ��X�dq��u.�0@̱}�_]e��iQ�|�*u���=���/���%�i:�P�ě�@F �6S�����<<sXlxVHYEB     400     150RC����+p��w�tI�R����Ƽ�*�����o3�z>���p:���['�������%z���ϰ���S�Q&���ׯ8�o�W��y2�@U�+v��U� ����%�;Y_����i�ηEt%��.�wn<b�������VZ^�[�«���28��@�E���]VQ����J�W��zJ�]l��^��",j�#��jDa�j�EP0:�G^u(��}��V�݀;_�����n �O�Ѭ��lˈБ�{��q2c%%�͘3�
xE:,�)9�5*���{����Dԅ���g���ӄ�Ej״��_Ø�;�jOXlxVHYEB     400     190N�%0 W)�k�jpI��UPƝ��b�� .*Ɨ?s���]u3���P�Pi�HY���\�ٗoº���(,���q:G��Ӆ"�z��EX�8���\@��o?1N���=K�8SW� Q�բ�J����9�&G܉A�!r��4`A�/E}��<��49�͊a=0L�ҟ��s��X}3\�@���b1��3�O�-�C�ѿ�t��l��`�ۗ�a�ж��y���s>����=dK�q�+�X}������1/��S�_�_����*X�^�|�ՖX@����o��Mc%�F��l!o{^:X�9�W9҄�h��o��O,�E�y}>fR��3�C{��k;��wp�t1� r{�tG���2������׍��um&v����{�,짶T֛\K^��XlxVHYEB     400     150$c�p��)�� ܏lgN�s�9v��>ۡ[n{�y�>!w�ze� eEÌ�P,�/(��3�ĥ��B�3 f7�-Ef�^̖�1V�~~��Q�ӧ�1e�q�&�?t 5�TQu����dRL�s�-�|p(��@����)�88�7����Plp��]%��vf�O�wpы����f�ek8{P���C�v����t���?�*Cǘ-\bJP�B���އy�׋�~��:e�#%J����#�>����6? 'yg�-�+���X��;�](��+Ɇib�З(K�+��'!פr4�	���y�)U`t�TWP�ooԉ�܋���=UQ	G��BSBXlxVHYEB     400     160ɓtU֊��s(�Gl?�[�H ���Tr��צD�w�~�y�ܝpO��#i"P��ؕ~��|�N����d�b�L�hΗ������	��z��qW�\w�f�ѢȆ�d�����,�rA�wl�J�U4X���������h�����tӕ�֘�m�o���F��r��t�����^�I�I�~nlg�ئ/�jay�7wWTm�AD^�>��><ɶ�O��4LeyD�.GYw�uӶ�c�Jn�|�	+åO�\��`0Vv0A�j�`�1]aTo�)l�y��rе{fC<?5�x�3M��Y �H�����m�#d�i1?���=x`��Y�����V]�8Pj�l��XlxVHYEB     400     120g笑[1)���w;c�C������@먮���50���	G�$��I�֥����o3gF������(���q���X�8�X�����d Y~�(7��="�6m%t�
R�K�.MI���$����)�3+DBcD=�&'w_ح����ۀ�#\-����5��(�M��|��'��f��Ž����H��DagzόSBG5E�7�~�G��0P;�NM��km��Eͯ'A߮�{}�~�k��s�‟��W�H�ze��S������yI�	}�� �Bq���XXlxVHYEB     400     1b0G�v�rK�����ھN� ��|iqF�И�X�4�����դ0�"��d��T�4*�B�b)�u>r�v���;�`tZ�ͪR�,��"	TJ��,%�~t8CJ�O�6f㡐�
(-��ק7"Hm��=M�"�)��F(#�]�OW]����;�E�f1���jGc(���Y�<�j��
,�o>��E������H$�u ����ԫ��W�}i2f,ZS=ha�4).��;���pR�A[{f�W��3
���&����r|-l�B�2*;C:����?�ڱ�9��%��s2Tq�^�Le،)�d#�?p>=7%4�=Q�kZ��A��$�3˘�=��̔qA$��EˬQB(����4��'m�v\�[źjL�wJ�f�W훹G`X,��Y��@��9���\"n-��}���R���+{����sx<��򹞥�xZ� c.@=�c��XlxVHYEB     400     1b0�=��)O�V���� ��^�U�Й�ɛ�ؔ|"����+��I��"���dO���	�,��o[{�zu�h8E>�*�Ex<�o<�R����q�H3n�O�ߴ�Z�2�>Z ���l�\��Yt�5�S0��r��@e�]����HƼ#�^I:T�k���f�L�!���-f�J��M{夹V ����E{q��?��oi�Δi��殮x�i�A�p��f?������W���,a�˭�HU������"��G�&W���&Αlٓ�ϸMg��˗�k�l��kC0`��9�DE,i�����Ė7��9%`y������4y�}�C^&q�8���D��_�|O	(�3\��w����s}���Z�����P�9���Pe�J�6�]80�!��m:a�荑�8'��,pj�:�XlxVHYEB     400     180�MU#�i��nJ�~��;�ۛP� Ոs�5m!lQ�a��̸9O��V�O�D���jL]�Iq�(?l� ��v.,p����W��Ə7�G/Gٴ^����\-[grBU���f�,�Z�% ��cL6��Ѝ)O}�>�:{�6rמNZ�mR͖+�\O�]d��� ��[O�L��ē���A;��#OY��zmU�g���H��kM�4��S������u�Л�;�E�z���^Ȑ�qO�l5�wʞ"�L�����l3j��ak���u��4��ߪ��?�cB`��f_�$�O�/��,�4�>y�4~�>�	�����@�W�8��$���+��`F��@��U�j\���t�I�ƾ.[�X3*GI�R��eQG����N3XlxVHYEB     400     170��cR'��F�Êk	J�5�����ȧo�\��$
l$�\�鼧���
~�����m:"�͏��G��/��MPBk��Ƒ�/��sR�y1ܾ/ؑ��d�<�#\�%�A%�n�s�Ƚ�#M��7�<��6��Ϲ���J��u!J�A��};�4��μe�mϝ�F�7���4�א��䅻%K�)�h/9�����7�|�jU��D�݊�Ӷw2�9���Xa0؄�V�$���Ǜ��.*��I� Yk�Ѯ��'�Dzfrq�y�3S�F�
����;>�\����0�O��`5� ��؃��F�
�fm�I#�	Ħa��J���=�m�� j�ۖ?���˟~e"J*�?���lY� t�XlxVHYEB     243     100?T����t����ȴz�dc$Y5���q��BX��\��E��,�!���u��X��=r�O�Ը��x&�����|�1��uVL�kA�D�@a�y����46���ic��M�S���l߇+B���kZ�� n�_زJ5�d�g����c e��a��.؈,��5F[%S�R�����[�;�%�-����2�QH��VT�:���0�Ϊ�/uKP��`7��פ�)꿨X�@[�W#]]��'��٣0�|��