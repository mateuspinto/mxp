`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
ejmy5WJSG8/SA+KcWL5Q+uVqrvl8NRgz2VqS6YSn9PCWfAQPBwDL3Z5YbjU9WG/oOqoW2QEHQUzC
kiOizFtI0DA6a4Hv2S3ECyrLUQf8CHxSxBBl1BUkdp9DVWLtXI3k0Dl1gymO1UHHF59QLhJKC6XK
nX4OA/oeeSsI7kKuhUb/4he1QNZn/gY06DyQszCr0JsLv/QMtEpuKACSbBbkfhH3UzSrUBMhw3yn
hG5n47oF6ShAGuGujfSke1yLKe34VozGGJiPQIkgLhCV7VXyoaLGAMECtLrXTFe3wJlL5/UU+TIB
pGGoYU9k/1XWMeUwtYwC/IjDZZ8H0KEAtwKfJBnq6yTqdR/TVmoM8kZR/4LS0Y5TKv9ws/CBsF5d
t2216DrEUUvUIGaYjSa8AzCka8KG54SZyAug/MakGdvuzt+0KAhootpHJV5MfI69NngC0zO9sUjJ
voEnYO/4IcQGapALiFgEibU+ZfylWy/yHTUCTYMo5QT1HrTM8YUpTP9ypMfMzr9wyPqjVdg0FenW
M4I762D1lDu8ekF3h5jAav7ZTKtHQPOKKAf/7YdNS3J+Qo5nqN3CnriHDAagbyzxONNTHYsAzdCF
c1MxvIBugDVnnvuzMgXwpoCDAYiDZt4LgOrIvBfU2LhnLxMfWEvicAq52uKTzF1yOe3pf9zeuPEw
rj1MYBHVAFRemij0KCwM1fH1RW9Lt8mu2l/FuLWENPjAF78/nThA1VtFZuNaiNdXYrdgZHzteucc
aGV6BlhdfhHqEKhINCAmPLBSPhdO0prDmSkjaYnOQ6iusAEBpr+8RQdrRmnmFSD69V1KYxw69QUu
tFuk+EvB9xXL2TF4fTYMEAb3RqvsmVilmzAe6BMsYyY7m39lBGza8aUjUhWT7z4qxeRvTMB2ZSzL
GuZUAO9KoM8U4bT9UAlEMCMGWwM5H8lB9SFozs5YEqidregH1PzmppbgWw42/QFMdh/X3broOPk7
7jXNB2YI0XYTeChZW++y21cChuUtDk1MvhQNKMx27Qppkuxju/PCbZcwV74YatcjdJ2Vi23b4mjM
AHRYT6ZH11xfv0VJSD+divUgj74t6uR5CVsu2aVivlsPtdVhN4kvaq/jZa1bRTUYO5vIFsCgIAIC
4aHRVwhjsgIlJSI76HX/2HMG8X5Avxo4bDL7khcmGqszIs6BjYu/MZMIZQJzxFKIqoaBQLP3ssop
84NbhI3pb2UP+hN9m8BTI8R6h7wSlfMpIa8A5ic754cotHlSUp9+ZZteD1qPCsTj68QniPk8yIEf
iqv3/1ddraVYN9AgbCs/bdphRAIflK2mMxL2ERDTCqlzedY1fG0w3e2jphwRMfx3qoge4te7eRmf
adHyvtY5QHjPk5BE6ewIbJWUuK4Z9CCU0H75q0J47YvyRCQc/NP0w2TW7lK7XkY6BdhgDsYnjQbf
4lvRkDpV9COt9QuUtTO9EHnZPpeuvGz3HY4UDJSuO8uLR2GCAjG8DtbLOEpIfxtBrIiLLIm7SVTY
irgTl3FxkgGVFfkHSXY4WaNXTEmG0jPASvW4pOgAMwY5gKZqmMpQv1ce1ITEopaKRmNOoqtSChwc
oakgatgGhhDVnNATEK6OfPc5X1fihfRk1YyDtoDa4qaGQodLdDJyNf4GiWNexMKGHUCH3aNeNe7u
6EGfj1ORlgv+IczSUKi6Yvcu2S+uQSlN+PGgeBwknA0bPqKptjHd+WsdmWtRXGFHUh81ttJ1b8Yi
XBr8A0G9nLz3sXX3o92IrFzPEOAyDJKJdTSWx03Dp321NIjxWRFo72iNpCDUE3Ziqeyziosjyn1n
GZl1jM+Krg+saw7UdahzmwkzHWVOSXOo+vsrPu6C9R4EVZ7769C03vTGz4XiWKzhByT+5qDbn2yg
k8AcjtrqQ0ogU7nvVFyrkpcKohv/u9ukgP22/oaHVe4kXyhEGQLgCow05CQ4Se+5wpggiMr8vwE/
S6jDSFogXhC04BBGUDWQXFUmxf7/EMVMq/QzPwiD1E6R+Ho84MFf95vAP+9CyQgibNAAZqtF7V9F
0VZBbGHcvLwOPOuCnSLaN0IB4iAxUWfklyYG7tfO/FpnELY6Wdls8kZk0G8VQC82mQUrwqaH1fto
qzBhcm9WL+eC3xP/e+2dRkEHCfJEf70M5/IgNdnUZ1rj0CeL+clmBCAMCNICuT7lyIyyLpAsRGrg
O+wPCNbFJhgpS97JglpgnDkEJ2TsdT+y5jm2XrU6R/0M8UWigsyLgZM6cmqp5pG40iCWX8ruWD/I
IHST3IUypoGK/ubnYgQj/WV9URYf0wypldysdpwmBYhtS6oyRSdpj4vXqL40/dTn71oi2sxUQkVw
9p2JPRj1Ipp+Q5ENFfpm+mju5aZJcp7cLIW7W+6CzN+PFcpQU0+78TGHRn0R7WzCH/hsA1bg2F/i
AU8Xsery40xYcij1g8lbXzaSVMWGVD0orE5C8MmItaElEcj4wGLr9Xai56q+FLJbGNK64k0l1xRo
vMPIeOxhY0nVRzgrKw0ITFWeDwWedLDT+uOfvU0STNIFfrGkvf3btUnVOZc2Y/irDbZJHh5q5x85
pzksManOxh2PJWrZEJtwEqGhD08tQjHbCzcjkLgn56MpuBAjisSpzp5pUoJnlmNiwv2/0QwkvZc/
OIo6Vzx8P+NZH21RzPgcVn/QbZGxTIXPMTuBw62kKHIhZpssODxgN7n6zZVJLhp/LwH1jH0omauK
RCUw5jGdbtTEhkJH4AUeJznxiui/cHHmmUSPgyCZI3RxMl0teRFMJPUPOB6N49eizMN/W8IyRYFv
qs+tbXDQ1P6YCdSmQfv+9/b/B4cDzdNWg5muuTI2XHjUoIOkC3VupyZ1hNCQcofFSlNrB8XEWsdv
g7SdIT86hFX67+ts0zYwv71nZ6gTzyD34OxGM/hfMCTiG40AhsXMZEdXPmODc849DQFHU5NivLoA
aTUPfPevDEWqdObthAgUdNWY2lBtOpKw0KAiKmpxb5aE39TmfO6uR2K7WX85cDvPUDvRen+tcbfN
h8mBYpZZr63IiNskbXtiCwdZ2Mh+3TArmVLXHdnVEmveyiZdvxEx2g+LBfhKOziuNTEh+FklGPCq
ZflYMBlJZbYWSQ6uDhArkTvRkIMB8W3w2yJ2hezLVPiirerUW6x5vClk3nbhq6B0wyJ41Onu93xx
zDbEf5E80+EBJ9enfMv7oXgHPGc1cg0ZUvujB0tKy+InXvjkA0L0hEc7TkD5gaDNvf/lpw8MnAyp
JRlteLg92Po5rKcO81EalKEv8vrMI/7XVl76EHW6wxCT7GofIWVbsa36ke5yqyBTYcHirdu9yq4T
qbWnJtqkqD9Xq7qpYrtntUkTaIqBu+LJ3MQlBix+2VhHYC+Tno93NDVeL1dFLMQt7dO7m8Bf62Cc
0PHCiC3joW9e3qDd36kDuzSaz7oPoDEsSbtsaCxbz39wrcVrrNQg0QKF7DpBQVZThfibd4N3h7qo
W195t7qQ5+0Qv6fk+1l0E/13HGS9qOG1djwhAR0zm6qXZPdl9T5hVf5J23PvppN9rIU504foZRbz
cKcFW8JJ11YMK35Aocs2A0MpJseR0xWXRlMOn8d7Q/1uA4AjZogTAX2FgkKsUp3tNaC7cG4Lz5jp
SXHQV89UmtBPWg4I+tgMpN/3+8D8gvBeYtKPI2dJjlqHQPWdsdx0QjDML1mUQtpPTWLkv45AfMWA
y9zUr0XkyPJXN5BXctzKhMIyN+Z/ukPGgfh8iPNKLXNz6ObjjBhT/GulK8tVKZM+NQcdrAHsymFm
FHe3IbDm3ElVP3T1/1nMh4wPQ7Z2z2VAZzdGmryrPnDGEcaz4EbjqRT1e0lZQm/iiOp9CfJo92ov
UZRH+n60WTDLNlZBbVxyGa16+UUixzIj6+5dlc0UNjafpB2fVVdhjiw/II0EA1ukAWuA4LD79I5W
3fcE1Mjnq/QmPXLZbF/7/jONPwbKMDeK5Wk/gBG21jjMFpwV2OcKk2BgxTHhPNyRMahiBBJgCvf/
EWrEuDTxrpF68aqqECDGrROhLF2LbnlmfAmnfwfINQ9If1Oa0/yTB08hN4RxFwS0Pf8K1/AZd6vy
M0uPbb/qCvMtSxiqaCCTK2ue5wURcotWl19kd/PfAtzKb6MoP8gaTfw4XAWh7rpw8Sk0PyrrLX7r
3B61jsDSzUYkm0BMdb2VJWCGZWK6vk0MN8+DxedHcOev0Q8eX5ycg8OcY6zhsSufZXqNOQM39v3L
skV/1SjNxCGchXxrTxVpQdp2gZkbWUzHErnCAg4pJ8G1VMPYclpDxRpzCqp+lyEMMSpZp+plrloe
3tGohw+naH7hqtL3vpFRbiYN/1li0vgXnjcLxtXQY7pWBcZ6a9lQFrHJCdnScy5Nlmil11lysqV+
x0gFUdpLdnuGtoKMwTnZcT7AjZFewAAu+iW13XSHEKt5BxII4dSw8gfbemrggd9OKqkErJk/BQrr
OQqmbo9uDMaQOJiX+ytX13SmUrmoHjYf80FNVpmFFy0Ohv0uJRBuMjkBdbTTYNNVyWheQ8S4Rwje
wUUJ7gwFvL8zZKpBys0PkjuBQbM1ixW9sqtEnlFy4B17ndcnb+PdvPsdvyTqXcfRKKpy8Pd9HUBz
Gv6ZpLI31vR4gYHHG5bAWiEhiwdk57cDByCNwmkh2KEK/3d88An1XGs9t7rK3+lq78aaiiAjIJq/
xKk+7ROYk+AVFzbifiX2j5l3gSmPucvkOUEs93eVvfDpTuZvJpFQ1wW8i61VGBTimuyY1sHo8NK2
24b24m/f6UCvxrqMGuRS/kXz6ORIuDdtOibAgHDeXoIsCQzjAZcojSho6aoMKF50CiMftMl6/Gx5
oRUauyHTO/7bnLAAsT/BWd5RBYkhN1Uq/SahLso+Q2DoN56eMPEj1IhhHCv/OGJ+jKmQ6exczckL
bPoA7Slscy1r48LkusX5noy4RYlT34ObiduSh7oxptovj8lGAfuL1ASHpVBkvXsfrMlQY3Qf6oE5
pUlwMTVBS/BmWHsLOFezS7Cc2O0Ym1Bet38+9bZx/+rvh8uz2KvUspRT2SG6nI0mKJ9d53bIBHx1
OXP2bRXU8Ic7Pr04ooLoOpChLFhkTLQOQkXh0VssoZrup5PHG5prku+P/sM6zNklyT+6IYAuliKP
OdXnMsRYoxMO4Z0cPF2cvSmFzCp41yf/AJFAsGACZPUFsldYaXhZogjb5FcAMknfrZ8O12hxHkwz
52bG3w1GVV3TOUBu7RZUC16dzJq4U6ynnCg+GIQinZ3Ifr4cH9x2jyF2+D/vHyLY3zXb2wiCUUoF
3c5N9GZyKuWlZW7yETpAzMRTv3JpJfFrUDGAuamaz3bz3ibk8QDuW8mVV9IYF1I5N0ZGrU+dggoN
S12sXthRPKqqnCNjgNVjIFES27skbfBh6uq1CeXtDYaMAwZYT820svjtW3ZCdf2iBygnzjsES6YO
BEfsaxx1v+SVStroTKJJAcyN5Ut/rMhuMcjAF7FmMiSZ5tz195DsOwWvGSGHm2zlmrCmIaJKfdrB
OK/h7eBGmWNU6Yg3/+fo2+Y8jrwIVJhBaY3qxQ+KqUSGmW1kNV8inohwTBwjo4lEZ7AdAKf0OBxE
Eg6l6G/+rzKEsd4i7dWy9wMpVo0KkijIqGuGGy+2gJ2xa1yeVPPsylpz/kExQLiN8NZxH9bOye8B
pMCB9OaHIZWHLJprSCrQ2/7BycJz2H4+Tbl0/+nnSx2RGwpfLCd53f4pCeRdy/7JS+VsAq0e0ZTB
Z4bqHK2c4kxCnERSdyQei7Gihgsn+Uc1u3LdkqcjGk2K0YDd97xwrc8SfMdp6/nJO1QgSqgR7TAP
1rdrRoDsQZV6+Y+IMBstFnIamYP/ZeDljgQk7n2YsKJVRjqDTCtaoIyqxE3Pd0FlgE9kt5o3T4Kl
4rtYmReS/oIZ/h3BBrtqPqCSYR9bAx2swelMsVFODklOt7jFwOWWqgycWUCZd4rbq15QaE4RuMvG
QI8x+zdUpjuzSqn5nohhdYG5Mg/s/AeChvz6LvPv7aLi9JJODEJjOLHsUn5fggO24mVZfk2CMBO+
limYzjhMl3T/OY3KWN2bZKW1etbVfhQ7BG9jU6yn6hy81hSM0tjpQQUZNnB+jp5d2HOJoIcTA1Ti
LpotofgTRhHrkUmM39JsPBvthIXwcxCcbGnUX7nfyjnZKZoCwr7T4ovBxC/620n2CIcqUeUE74mv
ZPoYRypqQB33iu8yfhbJYPvNpzvz35Kry4/05kXIRikb4ztE77b4vxHH+03oh/loTJbqwkMGNSyw
X7Xg29rvMdbckAfYmm/A5IUm6P1HPjAeTyPGcHhKT1pW8jTmzQyUJz6g8XCKaOo5gqTPx/BkAMlV
c1/1BmPkqFHkx8JFYr6H+e9EpyyYUQkdB3gxixg5LjBzUfBp5tyZ2BWoD1bXKBX5/r80iGWOywNN
OD+YuX6okNFN4i/8s+/0kIt/FXbo0hKFPJRNXW9BGOP2IH5FFsYyePIwRQ+S+kY3j8A0omQGouw7
uHnZ9aUO0Q/HeQAJ61v05esuiUTaoGIHVqVL0L9/h12cCDOLYqgcTprxfwmPNZ4ovTj/7ik8pm8x
wmRgIjaYS2EX4C5qbiSFBXfTKtR5rfSdBgFLBmdsd5kh9XBx02A1ZaqPx0UNSX1N0r+O+HZqIW2/
oe1PSqc9zR9lgUcPdWf2d6OIBqCkjRJmeGNJkEpNFH9Lf8Q0gksG3krH4Rgk0Fp1T3VeWbsh76Cx
+Pr7ou5WG7B1Xw+PzPGNOpqRPVMPbGIWCD25l8nSYrP2pEqkxgk7/7aHu3eviD7H+lVMypDprI+A
B1PYpP6It4IEOrwiSc4btVNcBqN36+D2/7xJPU+YS2bFubMEMU1llNNbvu13HvjkGuo/OIXCPf+l
4dk3sPd+5GJelNU6mFa3vhvNNBPV5jLZ+rPRfan36kRTDr+9HlbB1vYA5/YPOUIN1NFvqZdhjUQG
Qe+DJu88a6voBFBvcXpAB2OK7EDankR7ASl60zgD7daT6qzUlvaROgBcIwHBHVZztwJKNx+tV4bv
g7Ehp/Ut4Rto025M9vAwL9Gl2n/w+UYsL1sdUdtlyEN2WA19AEii7xxCYewz6hPVXZ1CEp/CnpsH
gTi/BIDLxUE44AB1p3VyIitgVgR7nBuprrYeZAGgxqtqMrIB+34fim43cRQLMIIpDwbVbMxlnnGv
gXFy8qbvUC/psHHPzMHWeKtV3OZIgOtZhdxV/4DOCPHh8RSQ6sHBVJbIrLWU87ThZrK3iZjwKri+
o/D4aXAJfhHHGg28PNN8XLtfKhfyYpchMtkT2SzSb+LIGP4vvh7BRtn6v1APJyDgpxjpAVdrQCT7
Z9bIm4LCdeRb9hGKBRcCcgyuRiExAtRug0bl2pDOOv1jFUDgBMixd6zynrNTX0PvedlzoP0Qpb07
BqVrlQXTWgmW2QJi4TL+yzv4FKch8R8K7qvuKh/4rSGQ2k3rQmGIqydTyHH7K12nDwHjq7nEhnTQ
2VMVEs0fK1G1TmCWZg/yjPzztZBsiTouOZiJCxlnZtN32gtnSDIDcjlU9XQwtPjbH6tgdAgPwb48
Qc3f5inNLDBJWsQsMQsKIZqH6YQnlE6t0hO1avxhGd0lgSCP3L/0OH6AVXOAGmLbn7CJaQDwDN2F
yk3fPeD80sSoF6b75BPNsqU0Z+pQextIr6ZZZz4kH1MFcun44NzxEjd3fCkuCJGZMm8umW5AwGy0
5lkB6nxb0lPpUb1SoOUIkgl4QmD+LmwqDOPih+1q5xFHx2MWW7Q4Xl+1z8c8ZuBDO8jJqOHBxVPF
TKzq2qtMaFcsMG+sGWZc7xVkjFqVNv17KAduifi20ca9iLh7KgK8exRTtGhsYbexD+aO8ZO5IZnP
cImOSBOHnRfiFXgpALZCVeevK05patbQOjyRbfayIdBxrHRDHRZOLfJOR58UeUqOMLCLvNkUi2Bv
1+venEuDOLENBiIm3+5Qivmw0OF4XUT6F0qekNC9qmSPdMVJa+2Fy1wntADB5hmMwee55wMJ3M/S
i/DDYEyj+qEnuU8JiUMtDXjK3djXy71Bgpl56rJ+CAbK/TajJ0mIYoyAhE75gSb8aFRCKlnEMAIh
vlUfaPjxi4juYb9c6OPHPX7++582Qq96UULxEO1NdenNkPHcMkNZ8w/zcKIDR9gcimg1yuCYcrlw
ZQv5/prFK2wbQEE+NrbqBcphorXZ1KJugVBsWs6Y47HgzP+O6qp6rm7Y+KegKDTY3YmC5IfTDuXA
HA1zPC5UZg8jueyZgnl2J76+YgEb7sg2eYT2K0UO01Jke2jlmt0NI8Sbu6X2jubuxRRuDdLJaUnI
IuQAiEg5EuYsXOeFKvz9U1jeTushVlXLPYPAlXEzMovJJr4iQOqeuUgDSC2CcYu/G+df7L/yhKsE
fGPMzfccNREtrA0Tuwys54+PVM1+vpW01BmCy1YgtVfv5Xo7RJAtVxqy55LmL8nHHXbsylTV4c+f
vnyEBotUyoqMl5QU5RsvISRj6L/r1GAO+oAmK7DAvv3xTyuXWzgMt7asUl8zFKf4bxiexYuMIjUx
bNHx60QinZEHKsdxNDroArQxrWAIxyW56C79naluttXV13+fgVl7VD+ARt/rpsW7RAIu2UwO0aqc
RHq1lmoDo0AXYNRH6z6pbXE4hus76D4vSyAH4luFfKt7FItoA7vhBbPEyB1t0LGD5Q/FHY8pBs2f
dZiiK7qGUt4ieyQb4qfHmQiiHQzS7UENPnI0LQBS9+7DdDzpEpeEnEkk+hAtrOCu2SqMLcYnjnXx
VVlG5Wgu/aezP6pG3KB/p8xvQKfkhFOlddvszJ9CECWRMejHqmaIhCmzGPSgmkelw5zwCFoRxQI/
KzXTkzMlDS1vJx+ZUluEN9XA5YkBijq/kLnn2Z08jnYiFohHnxiaEi0dbC+JPRwwARIUHIlsTOPY
beJFCRmaDhWtXV7WNFPo2kM39JKOBsTnOC4f4P/zlE+CQ5trz1+hFgxoDT710GVQ/IiPcL4E24Bs
cxqiLKPYxtOflzBe9H32vZQheP1OKdxoN4Q5IJWFBc7naG1eE5RUTpLS7rtz9W5yScH3uLcs+zl+
ebR6BHO1PyLHKLETmDKIdgz512bnC3JNFkMDtw5gbG/6xN2/Z5PVf0feu3kO/OvgmcxW/7emqj/S
YNDF5+a+ERELG4aNiHlOiLRqttY/7UUlw4agLt4+59XTY79+N2ZxnEwkVodcj94i9HyPbEa1k9jg
tEH5vh4oNqDV6ddcEonk28MxYkFd0tD5eeKzZ0hjTlC0Y8P4/lQ4vIu5jM0zhMGTNxKSiqz/19zV
iQE4NIRgjp5NF+AJK0xnm6DL7evJhKWgvLh6ElqCRvWbka/GrzTw8TYDYvY+2glThe1Akag4lUch
S1JNOsgckl5yTjMrUn2FDmpg4m1UzI9i+RGImeP49Pc5U4Nslws2SdnSKJwTGhHZwq4/IqHDBLsA
QnWeiSDolqiT2tOUa/7fMK4ayb/ivog8zeUW8my1Ixw/ERTgF0Y7QnIbtDF3UHgxaQDIf+zMmEnJ
x8aoFWLN1h5vUpnyNhcvcaxrXiLU5bhfBrX6fKhrqUkR8ycW6HCVvHqrJoa92JciE02+r7e/V2cf
OjjKws+IyMHGvE0da0mRvOOrCODG8SLyQZDuBiDbzpARMIgPd8GNBox91cHwFxSi3fBK1wQg5Job
YU62NfzEO2KqfpkauXp/TySe35ULgSwKvXljEaqWdeic3Gcsy8e2VbldmmyKZUya1uJSuH9sT6LE
LOA/2EmnBYpnHGQoZch3HGAkMBAPGctHY6Jd/5Mq4zbPK+lin+Yef6b39f+lnKrpzV7XO655Yv3x
E9DJiqUjtbYHMUMm3FKHD3KPS69IJ/cezB3oK65SFY9gMqpBz+uFIqr3Ng2oSzDwVdq9V9kPB1v5
FrIT+KGuy9LXFe8t0fq3eM0rh6CMnQv5qAZlthCuHDAmRqVxBmNycUgAe1lopQvfsURcMU3Dm8AL
blUtu4ugGaE3FTfrU1F19FHqTWfUfLNVR70NXvZNcQVRhZFw2ofaCvl9YGNPXdi9i/KuDHpE+BxF
3c4gFEIYDFYiGWWrd2fjcV2v2oGa1+OV1HTGm3nhvtBHKcs4IPfDuKg9aJxR2GAiLynlMXPyt0si
31Jy4kBG8QLEnl6Snsyp2i8HuD+QQmEeGCvcdLnOgAVFH/Et5vEBD+PPYMM0tDRddXO2IhYSk0O6
IeFpfTaqjvFyoP9UQeGi+a6OHFUIEY+YqpfTUOqMzbNoyAfm+Ysnj+MuZfj1tLJ+fu+BSX1H+coR
XPcAIaCQtQEM8HU6O0LZOutkW8LHx00p0bEuaM6VUDb44D/YQLBrRrqMuvSYpgWYGECJFvyE3AZa
5i3m+w2Y8xyRtZi5z5ZRpf5Oc9FZ3iyzwNjp2e0I5fEzwPlNtwDqTZr+x4Nd34c/yT16kkkg3kVR
c3o+6gxo3qt7nB52dPyIRkn+eM2VAT4lOkpOUqk1mechDNLHBSyxoZ6XxfKw/1lOMiwoW9J1t8Ky
FmORGEHhNPB4TH4EMDBdNuC0ut/xij84zGH92rjs+IV6JnDVoyWWEbze1QQ1ApawgoXggPV+mDWA
IMIp+HiWYQ4Nmxss3gL8h4/elpWnQ9XG2/56YrAyGj513/qxM+0RRrLC2HIXuYKvZvfiqvZ/ZFX5
UvZSY0odFlsilEeJPQnumfptTokQ2ptJpfYE098tGtaP5BSEzc8a4NMsNPkBDQqN9Et1gYXf1UHN
O+w3FVU2GycWs1B/arS/OoLEXH3vE9I1eyxDCnfvFig2dnkVue2MU7ehmwvJZt/agtMD1awF0cEY
TUKWPys/2qnh/vRxatr02EqWT49RxgrhokIWMBZXaKJxpRWMkNbL1Ug7r3Krxq5gIUVM5Zh7uJJh
qNtZDeCOogQM9aqvh7fSxb7W2ivIsJkU6Y1XV4oFXpCMp3JWyiuG/WintiDAmbr67N+pM7EwEWQj
sapBW2Wx6bKK9k4HdkyzFHyOpr2n8HbAwUkgfrETN9nucV9Ck2GFdevVMSj2pM/itjbvLSH+UAN+
EPT8eLX3AZMTiWYN+/6zDpoxJvKH+0sY8/vlgwIHoSSDuFxwDkgfMHomWRA1wQjLgCFjgX42ddOg
0luAFUas8d+7BzAIb8Qbl+R44sAp4Y5zB7duADRbpdDVvGRrJc/v5Ybx2Wz6IanN3ApNeM00VqRo
hHa6HXk1MnUlK0Of8rEsI9UDeo/MvwgJDffRzIaeoujTsKrDqphN9t+lZfa4oezIMto5L5kPNKyC
GecniZpF/pky7x4faageHd1XdIJp+47Nriw9HHLDvuD89+AW4nBFuroN8FXE0CLmLAKPQnQ9eioP
QFlaDRg9IhDygQbshMkZMVCaaz/0vbxQ4sEins/kk4V/8GaViHZzFLkcRl70WRfiDzC7RZ8YlKZr
t2AEfCW52dV1UJjy8fvgCyVj1Zc/7XClp7LcwUNniXOa4k+DZ8Czt6l2PuzXyNh32qHyZQXMM+Gy
lJ3leoIWfpbmKqNgbpAUL86zp/nFulI9VaRi5u5fTOpUVjTcMPA5C70DI37V8Bxanw7llgJv9F67
C4zNO9if2wewvl7DG6axmY1qVfDL9VF+HUbwcal8QCYL6k0Esc7eNTzPPcH5CXhPwTVx2UaOqMhw
5uiZKjyjj1C/fkMXkQXJ3Xhe9W5aMzZux9g7hag1jsVvFtCTMbQxTAJ8lWTlIrT89RTYmS2DO6mP
zSpHxUdqPEa9gFwuPbZMHbiEOXyr33eIwBoXioVIq9gKzi7P4zELaJSyK/0+HHmrgrAZrJHR43if
pyvL9+Twn4p3q2Bqv+8u020eZn8YOdXwIHosgMuwDhVe60n1Uf8zWTnIUWCLXOO0wizFNND3CSk2
5Dn9YO1aNuVVwoRHF4NeTfNpGHbWvyUgSz1uSX6o4yRH3hq8M9QzsOaAK56mgsdc/9edaE2u0iKa
EzpM6AKPG02tm40dIeWIgenELNLFtKUjWvloJqVmqxju5AOx9VH5J0fBs+SfBh2G1yj6GhU2U8XX
e5uUo7+SI4NiQURWxGmDjgF2BSdecMElSOFipeRsADBYU1FtiY5wZ7Men7p2nfYcotKjtn7zWIxX
Io2pdtzDL/lSiqWqN9+392hDOeKwFzF7QTND6HMoicuQ7H6zJNlYBJs5+IpwyU+MCmQfPi3VVSmN
E9eh4NnxPAQCRuWcQS6674fKa8unZKDKqkCPDZWfhjj8BsRggoRE3YgCGPXUIwMbS+Y/aty8wzqi
qswGXJhjJOpukAwctYrWNFhQ/aPnWHBmjvn7Qq6nk4+0MQm/fPeQnWiirxxrMPnE9zF6lcE93OuE
wglty/jXq7D3u0I8AM8hfQVPvSNjMXifbgS4AcnAWC8UHA7xvf80rIHxVhI+kwv76PaDVEYI8Oj3
01M9Ob47E5iIgkX1qHNAzqxsiTk1hEkYIR5UoM0PobRIxzbjDqDX8dEGKOIvAaqeGSn4MHge9a4q
06OsNONs2iR3VScw5qdPrMi6gqaTBR68LlYYsdSxN0j56giZkh69lQVpSHQCfu54jejJCr0HuGl9
Kf8JD/6775928LHy438LrdfWltFCv4Ih5TfaRw/vE0BRbdvx4LW0ggl7PTUNG+8+tO8sJbkT/L9n
0/P/I2vY7TEpyJ6eHShKrEUE7WtepSbXnwBu2BDxGyGd6eroQRuzVtn1Xs0+7VIs9y1T6ZrXsVXh
W3nysTOLwyYLUW2AOaifEINJGDQBnYcwpbePw7e+EDmK4y2LM15DXzoiJqUHWfkode/JeYgPHegQ
ii0Yk6MmjdiZyOkhEtO2Qmn0+UlJ7JEd1bglJyKyRApiiQKpP4WkxkUonZ/dBvHXDk7DnokVkWGh
0sEXTxOFMON2JYAAPqeR4tRv4fJVkzj7SauMbAs0XVi23bWV6ouZBR+03yN+d7cQKI9JaqM21nWG
h3YC8kevcgvM2lUN0dyvqULxTkPoAWASkLQzrb6M1uPvASdKRVA+1DMWT3uheJfnq8fNxsl4QjPp
Cw/9rA8KWFZT6ysGSqYNRq4gtghNyAK2LySh6SAjslax4qRsY0E/PveQw17LLByXWcL/syMO12g9
5rrvsqvlKO3O/SKUV05lc1UIFzLNa/oWwSnVkXPDv8HuY1zNVI147P1EkecFWpWbxVcJiLOOsQPN
axN6Vmf5IO+pQftsZzUrhluLRJmw0J2VXJgnLIMdQuMqrfHIo7wKZ0TuCrTBh5iinXnVP6cnQJMX
y7DI06ft1Hkks88j2kwJB4rnQtHGC84Og6Wa13QW3oaWAwIJZE1h8H9jLc6X7VJFoX1H4TQqfQCm
NcnHes5h1THbPFOAygbYsGcsHmjzEBM1gcg5bqH0PkCK5Q7xBLbopt51nOUDBx2bS1U8yXQF6YIU
amMtbm18sGoZisCC+x94HM2mtbRVe5R8sPh1pPFV6zy38CmA5ITbc+kldJk3+x6PXzHqBIa6ciJP
QbaWRCJltkkHtKt7bLjuEewR54QtUmNBNc2g9grlC9bS9T3Zjo7f7ayz2RtfmqUdO7w2qo4FN/ft
xAyrq7PnfblnxHzlj32TR/GGlOrvRBP6w2IgjXck3zJVUzLY+fjEl1Mma3ZfeDJ6jZvASss7xBo+
686WpBDBDzIcuPVrx/9NzrfZ7HNXcTjxAou3V5kSTQv6j8p8kEWmRfKjUUrCsZ7r26jD9AC3rbBs
kVWbsF6Z4vLw0GighHusDPUn7+QfbBTj3jjvUaDnizKoqK3uCU+5qXmLaZ2PGUMAMqw30P54yiUQ
fgiOfXR3O48y25zEwIo7SnMfZF/kbj7nsRFwyFnqG2zo+gosbEwzv44LAwGydMAqkRIwIUBq0Q1P
QbkAMC3HQuNHQvW63gLPi2BRlw1/deGz9bjrhiRaoVZDHeH+UaP7AZqieh0IXdYLGOZHBGY8xJvS
ssWmGqFvqij9kWAeBA2Muuvpjzv9t+krG8+i0Re50ss54QM7xd++/frmZGZtWuEnjpvHZSa03JhD
SmURDoKuZeunocgoD+p3tzAQlkDjRIyzfNfe1id6OGCkoHnROQ4oAhLDxo5PfwWg+niltVzPMMcz
U5pXlHkSNsM0XYi1Z0Y5KKFm4qpfde/rV76mW3x+0qfpLlMgsxvv6P3yhNjamsuTtl0FZuNb6fa1
QzBCdgIyiLycUy0PNrLCCU1wnrZmlT1kO94ah//KM/1/HFUZq93V/CY1uhSmQoM5lA5emcAI53Sa
yOBSCJ9NePcUmTji3cS8mJy1qzHfTgZBAa9p36lm7AwOrqwt7q1FidamvKpwtF0XFvwixKYw6Ltb
YA5hxh9+tGyCPxM+fYFzDaY81b3KzutxGTTo9a20lR76Y/Gba2roCUSPpUvCOHXl7gtJEsgqcrb6
/nOqRsw01jgbNtzPXcrqq5dnvafwXxasyWR5HcT2Pl4X0M5QlL1/49K0t8cGB1p9fuCFi4WKYxGN
Mtgzm9a5mSiVMoa31dyrgJtjEETCyuTRIzlklODoLZmJ2yau+tLiu+UfArPfbGYAT82VvcJUXvF1
sHr8VPSspJ8AgDAZC3MuEWNR0D0GytqwthBri5p1Qk1pDKpfq0x8fk5N1a71R98Y3H/HHeqRqn+g
Fze9BkqpeN0pj2Wao2QdcfHNmCV1zdq+aI7ulvx2LL2RGROo9JY2tGr23VYGA1hsQ5Ay+xOs6TfX
JwAWg9kKwTHSIqGx4Ycw/5FErdPeauBVKuWhTQC99+P48hGIXp3HqouRlIsPf3sucy9RpUx5HhOa
VLshZxFus3ARnSQdDUMXJSe2sfpylLNeq1POHbGwNAQj5tXUtk2EUNmq2VA/tmnlMAIH4X8iokJW
fLvNA4CiVkkCTq9CMqyLsBv6LYMgem/1SMKOyqVuLL3hIQrYmDQCBsL/G+gzG9dGPsqs8LlyZEgO
dmBQRnD5XV3rtOE/0JNeoNkNJsdm6dN/0xVEaj41EPE2q7Zhw0DMdoimlZ7HxBx9CYaAeM541xLr
DW1tCtrDmHvTBgQsiDso2ah4tlxQh02mTiC06/9dTAjtxH2YTYT/oTLLtVxKglIiDOKxEfNiUrTq
2x79vcrqugo/mJsgeCvns1gLyJiGgLC8RgI2S79IzD79/opysOgRb16yHKpfFtmV0Ev4MjU5q70C
bIsBKzHiImJ1pbSXQylyOU3gyI4sCjVi+mi9qmDqNAJaqL/5CZKTaz6cd3+EsnXjZUs1/RVeVjr1
3MivR9UoXNSM90EWJCi4QhNhFkxzd0NvIeI6sYpqT6fQ1gCUywyn+e5Gf3vHup2wy0p6AO11BjXL
2l1HBrmMpyaszocEe5sFxn8R/4lA2wauIAnQuT9zx1fFMDczAzKaEvsftVRZNBjsV990yqN5WTlo
OHcf0MW7qSn5z+oOdRZTn1Yn2yPF0RAykhVjLV9o1Bw7SAJ/tfGTjNJIyNE7WHjQhQ7UWd00cBna
Cb7MfzWW9reRkR3QQJ2G/Ibz0Kj7rXUYj0OYsBVmYTPu+hmRnfLpwhGsDUVGuNRCkLGHK7axVK+o
vYHWgW0e8Eoz907tXkiLTdZnGKyGpAovOaAy6jRNTHfuefQhcHAyYUyWPJPcDTVDy7yha/oxsctt
KOi8GbnaKW26APwYyDS+NTMWasINDW66n3CLnNsD2YEtZOtT0WlY812QWxe+R9MM8Ybmt4kVV77b
cRDfw9U4U8deBlz7G041mKm3jovrxPf89+/iqP5vsLWCqEA7H/clh/qBfG4QLZd56wP29KRj7LDB
S0cMHZHxI8iZjVoW5WebiHnF31JVNRk5PO92lMqm4otNQsgT+qaYuR5SPm4EZn+PhhgOhl2wyvDX
n07qXxCrBkXS3A8UgmHryo/cdZvC1TWANopm9uonYRDZGFlq95J44NrJLb4QCGuL2gF/LCOQrrTN
BRb2M5XxQboqb6Ah0K+sJu6R816a06NZTpQFCnGIpAI6WnKoOWypt7fuwqMIhUCKx9VAOh/qvTZC
tUiD4OIX65wXQa9qtJgtgEWLDjl6Aih2awHHRJZ6NIUUG9GMIlushSMl3uB5AIcFbifEtHjfjJlL
PDm0i+k8BLUkKOkyeCwVpdtHF2zq8wrlEn6kdA8tzjL7YpgtJ73m4jZuHRKtA9i8woSnjXhzNFRo
Gp5oNbnr5rAa0YijV3LApEMpkzs3fe3S6Hkt/i0/NqNrwnf9tKfPy/OAs68e2lVeB9VXk92udrNu
UD+Oby/OJImLwXhImd4M8oOTCoFREsSgXHMcfqogGzXSFPsjReCf+fk81Ca44BBN2Xosuk0qF4ZF
v/KO0fsxKwAJuWQ0BiLIOIHToNFvyFoVJtfCsNond5fRhB8RjSPJJJbKZWmgni/YOuUyB5ojbheW
pEQ4GF8evovKHd3sHgRK3vNBySmy0JpHdvUItJebwqzj7rQd8kxc9Eu8aqijUYb14Kcl6xqJTBIr
eOMmf+n/9ZFjPVtMV9gheEtOEmDaBYx5axI+oNJOhK+Wv9U/O3z/Zlqeb8epdepoLJVImLGHlQbR
z6VgDtStKva4t4BaqeAUlFWc2hmg2T0bQr73YkCiuKPIKXAVLh9cuU6x4oSQvrH+20j2n0+tg9ST
GwzMabp53ZKwsIYH11casAyalmybF6z0J5JbbkAurbR2Hkvq+UznFuUXjkUS/MGzCx/UTDms7XiE
fV/RpFBjSQ5wbMP/cIhLB7+sA2rdeq4+fHrs+rQq7vxIBBVla+d1wIL8p2/WWRad/WM7kk8hBv6F
JE0cdYcKbf2SKqVe6964LM/KP/Ine31jtueKa4ECauQONkYFZWOeaDnlnlSYE76OHLkpIiHmPQkx
O6OmaO7NbsgmbWJ6pmIp9rbLfQof+FckqieHdpMTC7sxd5oDSMER5u6UFO9t0wRaORw4sN86lNTK
CjPtmu1XePpKJdAAKcyPnLdguwyElsHS54sLCl89YPcTdeP+gkMyp1KG+XNhnMmOPEn13bDJ7mlp
eo3XLwdq2ieRHgzhcM+L+gfTvfiZAteAZN6y2afs2nrwmu+V2tV1s/ImtT3re6ouknRxHFmNLaM3
Gdlpi8yni7+B/95PO6MGmtd1TRhvK5hzUC33GDvI1ruyjrBrlOmWZAeJOak+vAkVVIZuadS02pRL
R0U7P5ASRDaFcaPYYQtn/X17hy9MkKOf0MU2t3fX7cR8ILKdQthOHVU+fF7sFcMT/sWsmj0IwMx1
eHQIDRxdd/jZJcF/jwpuse0VwkfLTGosciHPlr7Wj8cg5Z+wiHvpKg4sdfyHMLnvUu/VznLqK1Tt
zwgjzq4jEqJ4z99o1Q0HkaezqkK/miywEtEZdXp8PjcS4GUFjTg2GwhBFUcpssBX2xm8KIECOdtn
R9n0of6EO3iRQW+RM7iv8MZYwl13tsBKvUzLN1FFEJrOTbwcv6Q+cwrTpDbDiYYUYOPClddUTzmv
tpafdavq3g+h7waANZxMAQQ5nP6kuCatnQ9oPzmv3uqvjQCHCnclCoVABcDPsOOpXr/Mz/gu9EYP
YSoSxAf7ZBboMg6yVZYkrM9P9qajvrS2c7/Ef/WD9FZHYguF8SVVY4VN0IF01KrqeCDTsAw6V0jW
3QUDvQbZkmlL0Gq1MhrpMr23TUsIObUjF/d2BfRWNn8e5wrOLAIHE45M0oe2L0cJp6yaElsRW45F
mHM3Er1RmMCMSk/ud3s4SjYl9Vq5IG6MxGf6KP/atviPqj/U9VwKWnWj6FXh+GHJeUpGyOZGYGuV
5RdTy1GiXFyX/l02ssmTdWBm74nSGoOtBTphJJZ+0QYEUMch8y8QU7mreqnihq4PnakwMHD5383a
oYQFRm5jmlghlfYxuYpxp8zEgNkcSKrnb9QkDB2yF62pfcIX560STsy54zzl3VILy4Ct37CFP3c5
LDPnpxNJU7dd2yUWlf26Q51ttIyj68JeSXnsxpoNl77tMzbMs21YvXnLV3XcriE5g0JyMs4IUeEj
3AGuu0PjFLWi5eCkUF2symIUDQLUbFUKMKfktMbEzvj3bFXY10Yd+2/EjoWakKv4jU4Xcy2Ho2AR
YTUAXqOiOujBPjxPTqmGzRWTCOCODqYqryKqkwcD3NKzZZGGKUXSscC29s31zXJSkKFijoInQnZZ
+Ms5NgctKVkdmxwWheNqhk2bbYE3u1mGR1p1zVyKXm+c88jUEoknxZLLxYV+Yq5XWlQLWajlyYuY
5nVwHNmoSAXLESvqlLF7aJqkkYVD/FNbSQJZNLhR9FOtjHfO9sEQSfQ9bPhvTcPIw37vsvT34+Hh
Ay/qEU+39fkELolEfgBkLk+VEAD3qbn02dKjnR7JpVhyqdn95iKs2p4X3ZgSDkjJ6CI1sd5nfibV
9TeI5pwvEFtsb7EOSMToRJlmhOxItushvHWLhXd/T3xQbpj9wOOzPFQ2IWQIkXjm/aX+Ef2ueSA7
zJl+kONrW+mhZ5UJyTsapLPQ7+V6fb5fpI3vYTq6S8vRIyqsKNvqbI6UmW6lMWbV4VromPIwQMn7
W7MCBW7Zg2X0dvTLTSBrLDcoV7gKej1ZkElRr8R8Bl6m7t5ldGgoYXixejDYWYQA7zxkkcuwsjW3
hrDS8MwjfJt889lC+KrLC/LqQkJlrOuzezOQGUyZFQ5nAXv3GmWWhtEwhyfncqeX2jj+t7qD3j9M
bNTg5Hvbyi6nw0p7UWs0YtGZ+Pq/XzF6h6qYLo9pWrvLntXci1e7EvlSi44lthciJ8FKlgeITFxe
MBhlVRHgJYlAJBrsBwO40VFZ5PquiymifVq99+tu/eGXHVGY3faH6aSOpH3ayStM0bRqZLmEsL21
zFQZfHL3TfweVEDNXu1t3You6p/0DNoo8qHI/45XGpctEQ8/duVn0jNReZH4hPSXSJ/UaTXPx5+t
qBz5mtFZAPG9WkGRj8mNKnDgUea2wIy9sYuO+VZRiogMIbc0zOR5JW7ATQRfK/KmtHM8LZqJjOG7
seGkM9tj5SC2XdL1Vx2p9jD/AffcJKJ8zKX7XR9PCZsWcsKj6Uent9+0BOWLBiOJoUAKzTdW2YSb
YINxpzOoKodVKtyVX29kpboUYT4x7unJMjEAgdblPcqX0eNe3lFIRvyW9R6XyXTd8vqL0tBDz9Cw
YfV2v7Sbv7UwwWi9U7vMuNOqok7mlVolqBX5PwGZFf4lstxTzHRXNSATpk63JHFmBWYsuCXiSjkR
dfA4Az1bqZvI3lbY2wiGCI99oPoYdNSBLQHq5EpFl0WE0vz7eDKQWNgsXe2UCz5HB8buZHqoyuZx
kK4qq4/z4k/YWtFH+4+2SC2ApRqr84u2hythccg5cbVUBROQ5oQBbTSaBdZfXp02E/E2Ugv5G9Xu
1j5lhE8Ep2wXQFl6H0aGGySg6OlUD6WzIugxA7VC0cX6pWY88bBMuUgzbAZ+8lFDPDGc/8BgpHjJ
UY/RDD91nE1meTsLBJ3BU5ekvgrZG9i7fFpJIxoQj8RbNJahjkbfPx0ohoBRcKIRUsSU6+4LdsZi
HLTcIaEc8t0uFCU4G7v8imBIlfq0Gyvcfa60xh9ijqmBKhWt2jLd3khAVwp7XF2TPukNtlBo/ejT
XEakYSXJdNtFxlOoj2d0U4P/dxh25sH26vq/B4QwWGIYddyxMCbJyfoo9b9CjyXjQON5jmzp1w6b
4+p8pE4C2kY+NixxdOzCDQDWZGT9d/oYoMldNJcLh2n1b8skcdPiIAUJ5FBcumUF98e6lQzsAbA7
pLqPbb8M/Bnr2ZiyYvz7cEmENa5J+X5RcfqmVQz5hIqiykHl7KbbMw24Bg/lsw43YcqaRu+c1t2G
NKI64yZUk1Xp2CkRZ15Zb8vBJJvVhKdI5ft7mMQuOmic4T0AHNy/LH8W+RxVslUgZ9Pwx2C+n9OO
ZenYfFNwA/WVNLW6RsxIIl3J9sDwjsPV6CPvrf71z0bM6hxxiMStMDRIWywAwMwhX21euQsdKBea
crr+vgYshtuSV5UiQ060kvWNx8KjCS3HczD0S+hbT8K/q+PKpOF+6Bw6IDL5LAfVh501J+TDQmzN
KvOhn4OEMWTm9m2wiYCcooCMzMa55aWtJsONG8LnWRLx+4QlLxXTtWAAdsvd0yBrSBLDSZ7qRq9W
qN1Cs23oy6aYZ4Gzl3QCsJYS3XSnTqrCCf1vUM8ELXXWm4utaxVxi69hKVBd03OXivS4s3OpKmDn
eoeMTa8Ic617WPDMmin+B+Epok2mph4VJxmYJZBW36hh82z+GeSl3/8qIvRstw1ZIF7TF97lIQ1R
E2gV9GAp/qpt//+ULBzv4585YPM+dnbrk8iSp9wfI8jkLwUcoTu/kmMwikaSZhmQfQUz1TSfkJ0M
zYdQCQUqav73hrxOEsZBqi2G+EZwVQ9ee/5GBCV2UZGn1iFud89XkNQ0iqv5eprAMPru2QfL2cXA
SlLrVnrGEvv0BQdqStKrK34Yoxj8FSKA9AEXVqAE2RCPrIMpBJ5fNWJE1mk2AoNDc+e9M2veRVb8
xMFDBEYqyujiPMiLMQQkS+mJiZnpw1bZUKszIm5YfDTJ1ryRE1XphOKylWhocpF+qE6We5sVwjSu
qodub2B1LCkkaQZSFS0UTHCSS0GjBFZFxiic9q/jTFWD82vNK5mTG+duc4Jcl8MxIyIsc0Zm1qeH
zFf2qLDeXxHo+FcCJxTRRKZS4NW5aNTXRRDcSYP2eBvjKbFUv78pGzIyCuQ8XXVyrtdCmuH13NM2
Oki77hEOy6xD1ylUS5nTB5oQ4pRU78lbA8f9BsK7cI+Yu+K3cyemysjs/Hpmr+jk8Pqb0P48Ljqw
AMuaZbDsMGbEay/KyXSCgao/YcVlydA/8UptPvPQ1vzLaGMCWX9D3G2Qdn1NLnfnBgefhHnijLpg
DmehJ2x/BxNzAtgjKRXkYpYqzFweXVf9IeVuZGcMaUSH5OGFOBwmj0wgIzDzrEdAF57WKcCy96o1
NTRe1FJWOvac1t2JM/uA6m/YNgeh+3SGqxJvpmFOMPpwW4ccnwcpBiFIpLsIU/dIfsdgKhZbhMM4
VwVPP6r4teobOlh4zU2ZjZjmoLhG9wwlhFuJ5tSa0PRNagU6ADhVmDKFQO24PDlTQZhh66UC15kg
lqtHMw0xVffhAOLsLZ3ihoeEH8KNkg4mPqztOqBKTUUXyyHPzOmjfhpm4kIBWfos/lRcz+OKnI7w
7G2TsIzG3TRA8p2bQbcoxfoEj0qNx3zzwMUPhjtBjeDbvuJn0NamOLMzrJexvQimqwa0T7KNADoU
AE4FDAzy8s5tnqbs6E+PDgsXEEPPVNd2ayzXtPbr3tZb5aH3ZvbPaDhhc27rW0Ja/VeKEfC8NlCu
3Ku96yKSF/JwSZJVTwBGGlZoTD/I4CyvkfWQETshr8QxqmhQaNs+qZAWwPjTRE4wmgMReBBFcAmX
fx0EnsxeNDQNzTDJf1eI6BJenkm565oShsI1X8TuY12hgNakoUwm3kr1/p19+xcDrZxuAbcFsw3r
Pvgtka+dr4fVdBRB2AkRqBMFLz2O8VRLsSpxkecRzBRJih3xkPttdC5A35d4Y4KS8UmyNwuM3/4S
5rMflji/fGDkvCmMb4J8jA5HsoyaKwKdLaCxVeDCiHwLlpH5fuZCDHGJq9aaYncfbsBAz0GDzxlm
T+3dKmMg9G0vOpW4tveJFqrlH5x+LlC4c904bdi+dGHSJnXHx+DiotjLLZ4edC2FVOgEid01+pYM
5Rqyjjq2KK5fwxC2TQpU3o+ew2ra5XpdRw8XhBpMJPHxmG3k/f7/PhbyvRBnQrJZ8MsQZKhix/sd
puSJgBIx1590oHLdgSNEQQJ6beOEPBSnKvOk3jMa9reGsoyBbAUN0Z8+xhRvWe+pjIwrCCxtunDv
TtzN4y1SR61JVa6X+GzpNb4BtDLPfoDdbLby9skQIrmPw5TAp5MPgC5KNiqFF3SOBvTDCaKt+E4p
bJFT4lbTsidXL/7gQCu/wtK5AmgSi3Ci8XzMVnhKf+2foiGzmUTdgeMwrc39AFLJh/PvOVEdca0+
ygEcsRALsjShnsXqsSz73kiyqF2VQd/lwgd7EcvagOVlr6ZQ3ZcrXZYZeGLz3svFAOvJ2T9sddHB
+tvGlHyDOn7zZhA2bYUUYEvaQJT/X8rmiFJ3Bszz46y8WG9MysRg/hm6+kwHWrBCga7aD0N8TtWA
5BA1lXGeZkn13q1PZSoABcu4LJYSlSU2roMDJVn4cKJ8rA1+tf6RTcAxp+7xxxmEW6uRiXoIF1dH
z+i6DtTsOjaCgoYBV8oFY7y0hnHLV2Z/b+qnuOtRgNJUpOHaT5cBBdwtDtg+kt2fttTPY9HfFQry
Mqh+mA03pqREY5c5INlz2jq5n5QVZqwjJPxxp11nvi+PKL8g1lRKZFEzWQNWNNKhloI/sP3pHnIg
5HWmDHffvU91/K6kCYbqq/ZQNWuYa4zRETGkS+IaV+zbe+W66gTgs2KTUB5Lea++93Bx/4kR63fs
4qmCuWDBpMlr4oFiky9PJL008MvxU9Z8+mxlxlZjRSEk1Wi8Pyiu0Oxv+SXWvEhmMEWwRrIblvti
AAy9SPly+cStVMSKYPUCaXbZDd24nq1gxC+Pf3kdvCJcYG5kG6z+uXtUcQWM67Rh9bnFVceToeXW
xBxVoBb7pqeEF+kwQCvv6/LjFcvFgLL+Vn0Nm11wFyUHpXMQP9iv3+/86O8tFDEYZoO+Z//0bClE
M7/XhmRRibjv8/9IAxl1pQ1tdH0bX+7B7rhXaYJBL/LpUlFIzKQefvTUdqC7M/osJ75Bi+1sRI2m
VCeGSr1tCRUFKMcFX/N7u5w8qVqnjU2GOM4ClaymtLgdZ9tzsWqVV9dJwisOwpC0dRVn+vwW71Pt
Dse3j/3jCtBzGjecmCjCBRTKUOMoK/jlf7MbseuOjo1EH1r0j2vedsRaI9Dpqbb2DphTO9kp02AQ
DaRoluxPLKFmPkodausNYeuoWL9d14D0YyuY1RFe/RpIWtbjBKNeC5Xici/olj7Dc7znEOI2TaQi
ofFc5d6d2/lmyhnglbZmI0kCBRk4rRuAbp/y6hnVS27LTBzXdUD3YoQItq+nsaziYmTv2WY3nT9q
okZHhcayDO5wt9X+5+biQoRDx2b411Fxyuzr1Xff/G6j+rAPTk/cyeTgNKAuEx2aqOD/K2i6fJJj
EI3Ksba9+puGxXsvKNXD1h22KmpSGubGFXexIehdheOl2v3LTyGQHsgiexvVeYfV8/K2OGaOOd4d
NjsEXKjyGsARne+9OuXXmm915nrYlWpbbOtNuG/WhtvBDW6OCA2NH9vhnDixc0E2T00cCubrQL1q
L47O1wdf4NsWCvsP//7PKXE7PAITtjZaNB/S4DaGZc4TI+fV3Jad5j7bhkM50gwHalD/49qDmL8G
dXIfxcYFFbCzVzJJIqyW26d/QcxF6CMCK3XXPuwqJY2K36TLlI6GH4MeBZPBUC66Rz2Bx4cTXAWm
haQQlSAzF++5kioeT5hjx9gnvnBGMB+EM6BOX1N5qlltOxz4wMn1WpOlG35RiNmesi5TFz6+GRGq
r4kHU9sDXABQ/HGmDiPtkR2BIgHyBCGjtiFkBb3auDkTggqd49KFozd3e2udl5tXGISipnNlNPJx
Z1kcsr0yL6bnTdfjaTDcGIIqXsMvU+U2tQrlrK/Yr3FjJyA6p5P956rpp/4s30OJpCvE1YkxkXCB
Ztb23EPxMvA4JaHm8DXyY9qXvkPIGLzwWLiCbJshFvPVVUDMA6XyU4AIIaPNy/6em2VvEOVzAoMz
eUB15Z+D+GLKVRUHAskrotjEGwX6IAgZVY1TtmEReA+QPdTU9lLjr1kx79uYvQfIQncTeWFTO83z
UVRaXwcdsJCN3e/p5eJmZYmmuwZ8mct1v46r6gWNhMfBXftSZ4lZNhkDb7sn+drs3dbWEnPH+kci
b29qhD8rD34UiRv7zS57Miab4ZFuxlErZoIWbcxw7kPY9iXJ5knJS9e3DZyusyMuNNrhBe7Zsv8f
u97RHztxrO7Mgy5Gv4KnISfvDSvAHk7qPYOWKwH66RXCkeKjb73QJESfC3z7m+ArL5D4yAPtwoZm
cmiYyUeMIPXo2TubBKxanasgqPdyXXCAS+yYXflqKZpfzfNl2WBi6+BUCBg3+fJ9Xf2yhwUcWbdA
///dA7IJ4G3HIj20ib7o4QCYiJtENRXVVJ/nPmOMAWa6h/izZIZIMz1zx/aPe0A3ygN02p6+4t3r
fjDxX+BiXx7MmmYfRyQhiafozpa2vZUIdBzQmXstS3KxNfv5AE/kIJ5Ai7Bn4xuar8PIlTk6kAwe
GEq20ed+dunQDS8e9mGn+bKnOOtGDzgddpYXDBoW76J3svqWrpCLnhqfqvDFzvi/9+JK+mI4dgOM
teSPHMY75pNZ0MfgTvJqhwU7VA2tpa9S4mkKFBuK+RUQ7S/tmee5By3mMSqD4vwhwTguArQ4LJEu
0hvV0jIMkvmTLZMVhPsC0Mj/xjxDgvAHjXOvxemegHWjTudXP18f3mi1jYM5k6yFmOx+8zG6sTnI
zRDx4M4zBorImuhifAjvNPhMGDul035KGLXYoeTrDp9jU3EM4yIzeyFPGPJdk+IHIZY0L3rkWpUY
2NcuXhKdF6mm99kV1PfKXde0AA92BRhyfbFbsABaFD0qkPKPEa8O4DxZI6svyMhGlk+aYhu5Hksz
03cn0E3d2oJWa67QXHuSzigm+e0Kwm67VKWyxe0fqSCRyv1381RFlOXsRXVA5b75d/PskQZlFKj2
aRh0Dc5Ag7V6HET99D5IG+MLhuMO/jW9GD3WLU/SAfd9beu2IL1Mnyjlmw5iRybVEdnVsqg3xs6h
To5iZUbkuvmSHx2OCQphGIZ+UnWCpw6Br289WLLssX+Rh88A7AJ+qvuxR4C5yIqOHOw7ZVF2r5FB
p/OeqsWLjQ5isyKpRYZ5fE2kDUVtZYMdUSCJM38xwXt4BRwIoBfSf1CDwpB1sKYU0gn1HtGK/THy
z4rgTaB6ytfCxZsDRVsUrEKKGebE5GSshsQWLT/keBHfTkY5EuNpIvyOO8AFdkVJ694U70qZ6eBe
pgRgE8Xl1zlr+vRxFK6doUr9ylc0z+UsaEpCB8VWdVlz0U0hyiUldUOOksLOrjXJ/OEeRjPH+AW9
9M5F0EM7yq0rhPoF5NkrjO1T1n4ggr+CkHkFAxfNIIl8lZ9BGzSJ2BoPBwYSxDKa/7nQfvYy7wxQ
mgduciKDt6myo0E1GNiHoW/siEUoTho9MNoQQ1EiGysD/8780CwVZWfZtszHcV4mcJqnUxxYi1Mw
isDici4JNWZFAyVbQaQ6yRnB/HCQqVt0jx8/BkLTDI0dlj4MIXdbMmnF7mbNarfxDHDl7/h2Nbi6
tbgHIEyvTd4TfMFgBdEBMfgCr1IEsdYtO6GZzbQJ4LWFmrTy/s1uAcLJ5ZN0WkYebIzDyTKe3iF4
tWWXKOc0HQ/KVc561+tuYLL9YN/2B2RV4LWg/YyxHo3idOo2S5E2gXF2ZaYfLwlJvq/r77jAEO3L
vinPAQxKU61m2FzMm9vvCND6Go/9o0OJXtTmu1EQznu0nkzIwWYy0t6v+qPRL8iKLnQW6KMNQR0r
Y5dJ92yuRrFJsV7hpc3tkmh9XjqrigWpCQis5+rPpcQF9iYPsfGom/zn8EIjwKKJ8aJ6/4TOI7bT
j1LTfCAjah6SfQPhmvKlvS6HtHmSHp08YyiNNyhN5/hg6ZbS69h1L1Q+aS6O6yaw8o+xZf79vurk
D5NcarkG2K5ZOTK6fxNdnAaHWW5ZOTH7/K03qlr7a4h4SYPKn8vqEsFccd+XKrXBD+EAtQncFv0v
JCrYuFRGgMW8vrn7DYFRq5To37Ebj7YEMWETLf1EAOGWGR0uefSGf0EEmTlkCJefzCslGDZbInQX
oaKl+c8sIKMbdng12G3aca3yDq2BFwl489z0vy7rEGJ1GavU+/9vFPZQqvad0g3qe/y/+/mkg9AP
tf5g+vnOLjBfdojgsiODuIyZYdjkm1U9oelctAgOKvF7EGSiex4/hUqYeORQl3Ethtf0OJT3f/7U
VoMtdJuHefrwbbhyJG8dqY9wY5BAl/qBgt8HsV/9w5J4kHNsrCBOqpAoAuiyaDoUHyW1Bd2t1tsn
OavLYS5ZmXsajxVNtxXDAQxfQ9t+thiEx0ywKdvzo1k/jrbwTH5xpHNHEQ5V9LNHs/JYGjO8zZWf
yq/cW2ZpzVdfOQbtAxC4SRF8gGPpOTQNOOh+lAIOmlYUqUVNDFsS7QzbMcXUqzHVPV9KRGBPbmK1
PrULS8Pel9NDbEJCvGeiXmbeELxRa74beYzXVgrH3m3GERBUSj3dHVp0PkL3hwKGYD83rerD5bt6
QdQjWHNodSVn6dfmhOyqd6iotCEocsWvguWJ5cUh589UPU4P5IqtV9ctLY59ecRB0Iar+qpOpCp4
sLJ6IPO7od4b5bHmuvZ1vbJJbtg5LDDxKb9hfrehNonHqD0oehOdBm3ow9d2zE6ufz/YzyCV3KQJ
PZVV50S992ruxalOyYH7uSoWhxHyhUd4e9LymWkd5ghC9og8Giei1n1izLuQ20Owz8B5HkcQ4esK
SJprJAONbQRdRlWwm+8vcTzMyPqFwnc8RP6mK+M5NAIuFfP2hBtXQFWj3kshO2bjR0Mz1guE5oNA
nzAJPO0wGMnsigwb/xGpBWWuLEiXicjvHwVVBz01lTGuUQTrUrX3BdTbi0Ic3ZyUJ/6Nhjb6odSM
lsmHyRb/6EJv21RuhaBbutoASac6e+lX1m01CwcY4Fye0CMeiOko86jz3Ix2cSy8BMUMqGHHibVP
ZrsQ4T94rtG+p9o0l26WrjsoCZ5srGfqknsGaT3uyDKCKiIrhs25luliPo4Z/uFCtLqmlA56BSo7
ImhGFpYx/0xwpW2g/YA0sBhIPYZbx/9QLRvVp8q2dCE3InNU9dRmQzU7mQ2xQkV8izxaBfzcYyAl
mU1xNNTS8bjiS1V9HVnXQlAuzVfptCCsePwC2Yt5oUeHmG6PbCjmAnAAolJxqf+pCrFpuOFijzYL
il0UihbYoIUgSmOoQFHz+XesgBwOA6NHSWIbt/QPwtJa6R/z8AkYO6+DaOwA2+KpOmkQjq/0MeHQ
5XppELwt/Q/Ej/kGkNfJPwDao7SLWK0WFVKeRUB6U6WmY+M5msmJ9ZbqcmfRzx9STmouYmzGGsL+
QB736Az5KmzxDfcYNqwT8DweefeEgdnXQ/CPWZfMbvwQBgAyAyj0K0filxhG4IKjdSiKomgZ5c8s
Ds4hDDxRQLuEYXTCc7KnDMuxQPBFKioFUDFFMugebr7KdTwIycm7gnMnm72uAjpueyxdeJgLELV3
ExnRsC8LgVVGo1vZgZbaBTljDLl2KXvPjli2RVUebl71V9LlrUJXCVCHedcJnAodKjW+urO487Oj
Y9b/a/1SmO+bXEXJ5ZtI1sZfg275hWUGBOt80HTXLiqwkUvIW07lbaLARJ2SEOrRBzwBNkCvZ1JT
OI1m+y69dthktIhstxFVdY8ISv4ptgr+D6y2MGrigT85aArcRmFVSfaYZ1n4tlsjwSRY+RFQG+Nl
iDk62jryR5/HUZykh1h23Q4ge9qLfmuEn8EUn9yeJPrFIXlZXf/kn4PCowayT2e44UBjUEi/OzeH
gt3tkOVvaSyfMGRLzXWlpWxS8K9vR4zAYA+9EU+dBX35BWBLHNpkPVXZHG9tM8oBqdPStQsrVOYs
u0qFzYuEd3QvSqvEOegJxdu3YnAmiTqtxRfuGNTiQ0mGQEVKtejgsuYpIG4yeMMK1I8W8eHblIWa
7zC/O3EtCGF36oWrfgsxRein+pMd6c+rSrn6axdZ+pA3zI1M6dbl0ReguATsvt0J87UOKhP+88U4
vJICEvDKV5F4TJR0yTaGPW6FQ83xVxV0I4OIRzjG5NwwdVkW1GEEfupQojsPqX010o4b1tw7VxHH
YMzCURDtMiuJuystqt/55SG3iwLg9OEmfQI/eYdGWIV8Ytw/9bKKe+PhYqEf1IYKhR3LkyT7iN47
EbSo+Zh9jp/TArcadBCz6yG1bIxiEjKOmRdT6CGb0NpyP6lxZuvofjAGOxnU0vjp2NHJXKUgbChC
kTbppZncl+kxW5MzCPR/53FVweldQlPi2omPkYz/PHZtyRSNlbtinc0EW+NnPIYyHI2zTdsA3UGd
yzdu9WU9SEoABkui04pzVhDV8GDUfGNtEC7JRp/4FJa73hqOUeyb2HW9Hee1mtLrkCwz5b7mtmN8
HnMwCvJbN0cPlSJJu1ONkgY5gdLQS6K13ZCHYudtk7tRFPI2+QDqVBmsPILxK16ypONa6Q9GOfBY
hD057L0UBCnpaCXd2GUUhvbWEfzedH4uQnA+n+TQFybYMdE5XF6FItLvmU+1YRE5p4V/F6uyAZ8x
kWsaz4fpIUr3Q1yyHMHXlKA1RIEai+FHzn+RKJYohwWgeAgtJqkAJ0iRrFq2ikPRv2J8ydtFdWcu
Hn4Iv1aKps+dHnToYTrCZfGj7hV3CHwpDYg3ausDTmN05SgL35DKx3LpogwKeRD4A1U1bWN+jaDP
4tujSg9txHSP51XR+VRHZLtdZe1MNUI0FU/E6jcu4DBHUWpWPYe3I9FBwUOYMAthgTvSBcN9WrmQ
iNWtybbAnv++b3weRb7bhwnKmecHAgQVDPu/xM/1CYpvxw8P/vggoZ802BIQA7jOoZFJByKqpMZx
PMSGyz3rSvPKUp6sjqZjBVxzdv6urJMPFT+7NMOI9XJdM0F0mQn+opWyY1uqOEkzO48VhMDaIpoT
pVoEpys8GzUCMPFJjP16FmFsSt54eGxlN2QkVf8cbIIiu3zMSkTrCQco/a6s9TxYBC1q7GnkR9KZ
pcJQQ8PGUc/BCgatEOfhxiWWBYNf6jQ1ZN9qA/DwTyW6KFj1TKv2Ah1y3TqyGTzGNn3colzXXiQ8
5g4/sKlpWkpQrrz1j46TJik+7brnCL1p9cLfDcfl2pfx8po2hCm7kSjbqRib5WmbfBjjIA+SG2lX
+J73O6ngLuKkvCTCjk1M7xKUvPWhV4l35zE35wJ/YU3md8kwN0wClq3+IiReW7rZvAy9Oag4JpMQ
XV9p2NTApj6Ck26fo4Gdv4DtAhBcscpQ3Nc0Wqrt046yzziYxc4A/Hn8Y9wek6P8NbpacYpaQDGH
GW+5N52Wo7h2mS8/oWB4Aa5ZZ2xvWLvTSurbV+Kwt5Tk0RDpQBCPShI1pjlvDqNMjruVTlyErcNe
x4HRHNX3MIdResC+hpXLbTYv319v1fqilRbHkjLJ3buNpn4G8xe9AhXuQ99l8HxSPRo0f+yZFsx8
hhCPZBrxLhFZwb/GzY4glkEr/FDwJ8+hbIQIe7SdmYhBAL1ysUSlj890FXFJdqMsFeKWVhWThm56
uAmAd/ApTJqzfz9s23ld3TGOc+wPYnnDMbAY4GaRHgh5bvnal4bM9TZRvmQnVQ3vid5hBJc0MhZT
I5cRbedjzubAmdLJADb+HTdTPiJ3hzxug49g4+dYKrqarLtN0junhrIO/adotgIagJAhheQ6SGsg
KlDZCLaAh8hsBZowyyQextWy6ocv4RLcoMvN14L9YZ3IjB+aq/zOsztf7VYovRRbcLgfeRdt6WQ+
bXd7+b+w90ttofgcnTxQ2Mlub/mPKWfij4QSFsfCqlnX1jXMX9NWA0gm/7KlubbVualVAneLHcoB
Kk1acKqeYamHf3F4yhI9S1htLWG7n9p8aSHNEw4WwbkFjju6d7YKHzIMU8p8MG0wV0MaYz5LUw07
qCY4Fh70bfvmZK78i50YlGl2ZQpSCeeNZNdDlfp4OCTytg2nKk4pNmfzN+7WSHPp/2lqZRbqMps/
/BxMreP4Q2EJCNyRyy3cerQsZ6iRFroF30fknwOYsnHo3HWyvzYkCXw1so5ZIT/YNhmLKsHbz9YL
1JrPCPzjzPHwa30SBQato9DWPxX8lHdic6cFno4y2Dq4ucLPjr2oAQ8OH8cB8gtKnpsaUlm3gp1F
HYRje5v6enWVzFRaouJWb94aChspC0VBcHHARW9beI1Y7LWJDiBoEqy3l3S/O0yMUC/Lxs8R0eMk
aaTK7KwZa0MECw6dobYmA+cGBSjQ5+icr/ulll6P5DFbT3FIIX5KTrPZMGalE5N67FZ5HnRAo6m+
8E+/hTTbsyEoWr1oQ+X7XX/9Rs/L2rBiqwDSVpOlynLNgwLOcls288sSVcGEf5gNXpPAy5cPx9t7
MoXm1ODzcQVr18EqX2SSluuyMh+bo7Skf7zeReQ0WU1Kch1vyeVm7tQwhcC2dOpNqkHHd4mlDXV2
oFsGslUHr4wGbrVMzmPPhklHE31GgF5RfG/lwIc8WFGWM7UEgpL3Hl1gGdHVTMkFPGCrSFZo6+95
JiGi/qAVb6pGjlOWcTWR/wzTWYZu3j+rooLCnTFFd9Klbr2leR0/m7owBzeboDn5CAnZraRhS2Un
3AfCOQ8mEdaV91FVxukrgVXlJbKpjSeEo8apw4qZO/RMCMQNC6F5zjQxLEsTHco5ae1mor/TWi3B
8uu6ZZjyOboC/EsWjYMfg0YVE1bODwTb/x4arlsJGqB2R3GhYJJhBP1G64zEopY4o41QN0JcvWt2
bvm9fF0mFhFBJFUN3RSc6v6Ibxv08lzSsG/BWQjJoQFk7DVEVoPmC1hDMUDJcdK8ltaJMuZr/oUz
Q6ZuhqnB2pSy2jySyI9YjfMfSAEkTpAbJNPKQrulnB9cPzoRNbXSFWDyH3Vl3GEOoBeB83fwLLAD
SaA0Q5ZTxqJivZdPOCiLRMDuhs3QaKDW+UlmSo7Rq8S2URFXNLXQ8I4zL2PZVgQR8//LUb85202y
12dhfvsgPEfxpAUAUYEo2muf+jeEwkv/uvtdrZlvEWCtJpdHzqgNzRVjsxvhJDBTO8jY2xWS/bIU
WVxl3UYZzzRQ7OazJopsvD9CfvVr8seCv7E6WNrvhYY+mZmdx6Fxbt1uX77UbYDab7zy/4Cr9Ule
aG4KW2vTDLoVZaLX4p9JuigcC0nXKHUZWhS25XlECS68MuCea14uDgfQed1aDgbPcB4Wk8Shv7WG
GfPNLlXbFFbSjfhApwS8LsycO+EK4ev6BmQSmMoDOEQMGvslTZT5gBJCyMsa8Y25q08F6wGx0dc5
1eNhoiNTguWcRbxKf0lfXPYmJPRGRxE0bJ/y7dzFw8ewHecLC+OdlX28LX5DhS0+ezuuBBUKAXiR
EO+VVxgstJ+z02LGQ6dOyjiT9OIx/Iqh3hMHGem5DSFNjJjArVok+lUEVysYMecneSw6H25oHHV0
exlU20RcYQ1OWujBMh7UpauQTzFMcOfxI48qGqT6dX89ZCFTD/X9tA8GtJgI9pNFiiqka98PI4d0
iw8KNsw+5W+B8vSrVuFrNKtWWdQhTAU3MbrQLVYXRWoaEjbJxCHD5s5x8BJehRmW+rM7zi3Vevxb
IZclK9AaEsNB8KcHGaoLkA8F/ewGtHwQJWy740pkLsCwoa5PoGhtmavOdRJN3K9IImRbG45T/7lN
QdR29nhB/rNGqU1NTih3+E1kAUVNzfjem8N+y0gdVbCQNxYB/Yl3nhNOGzumHW1agSuM76HiwzzP
mj9I9hqKe2U4tvweiZFyCvkNWGTaK7A+OwwLb1v52XZtbW8cnhqyWl6u6QlXn+fq0ySchTZlY/4R
W+/LoHRsyQ6N7AURNv2dCCBbGQcGlNroPYbEFEYT4AHj78W3gjCyGeuiwiyNkHqV4CNiD3R1pKg9
Am+si4MRA4OfkWq7bBtZNlH0ouFUmseKrGWfW0pUpRSWodMITtVdUx+cz5YFZnSpqn3hn83AHjYZ
3SS8QKxBLf5RgzT6DSyxYryK4sKZpr47gSo7gFMc0vyEYtg5syFDg1uDK/UvOEt+x5rN9v8irdCe
YNNEuw5zgTpfl9GuT4WVVBiSqpyA0ixWc/QNU9bh8ZM/0OPZGQUI1mMFC264L9T+5+WJtgi2psGl
t4Um+m76wS17Fu5q137locoyilCk2FNARgns0/ESWC8gKPT+1tjh5/QAoWQzDo9/7Lun6r/A1MEA
8FRQ12Z9NV00KFvSJkBdJ9j5RD9MeI5ELUl3rogo+RKaJGwZIXAv2wiGopbgbDHGwdHlZh/6t6tJ
ORP4dKxhxdMY0j97TmOURmQCOP7aofFNJ7D05JfIf0TGZqoXLRU3HvTJ0gdBYLy86CeOuNW4w65T
Sb1KCpYJvMhmUMR4d4LUgcbXaPeByN41tTXPuvSSMZ4aoyCeD9YVdIa5bzqcbrqxNLXjlrGroz9m
TzwEyP3B4WCEmMkoAOWwA8BSva0N1szxFAGQoo584xTMh2YeW927Q66Lj9hh1vBo+UhU2vF1qY3z
SJ0YccIrm6xIwllLm0UpcxPqEKtzDWOwmwzNsmeBqOLla3WdVu1QyrQvCB0EigVFcdv1e7YdvxmU
THFQn0e7e9ITvcdH94+0jHE4Uo2sRu7mikFKM+zdTjyQvQU7uC4yQCwimg+hn8XoaZgZ3hBBHR2K
B+FrRRrrjAEBUfPj5NR2iKLxGFR40NlpkQ4kjmR7XFO5z77htOPA8/ahBPRTtc76cvNDS2mdlpI5
2+uyDTISQuqtGQz1do6z0zkFPPcrGUpWfVbK+X3XXXK1Wx5yVae7IxkUU2uhtAXd7OUAFNu4ovbm
j40EE2GQwW9qR1TzmIanL2JW+s1Z9VEli0mjSjLeDyUIH5gJeA6E9RaN1xbpb8zULIBPts9+Pdb2
Zof52eOjbAc7n5MwRz43PLIqTB+xQz61rzESqrDD11EyMWXqGa/IKWh3WNPFPpRCzaJsWj3mt2wr
tafsy9BgUqqqizAeeIJepGSFW3DSJm1NiMjIhoAO2W7MVAGj5YGT5Ovv0xpKnSPpHZ1LIhwjxr+k
n3ee32ENUx5wigBwndJuC0IOLkjQbXGG9A15jiHqRGeUW0MZPdYAe6qY6bQ1M0Ew38BdwqlDMckD
0h+SeVvOCv+wfMotSrP7nLoiAQJkPpu4KjU7US2RDeQaj0VIBpTRMjhYuHLEgs99SmoImrKdbB5e
0wan2OFXBXn49Q7SZA4p3sd0zvNluKKzgCQZzQRtYSHlYHgUZIN4/vdyE65UMwzCibk5bFS2nAC6
T5FNr328tEWNMDmAbhr3KXhIyo+FwkWYK3LNwRRWKudwwnRvbqI09fqPIeqtdl51MpOpTcDD7t29
lryzv6FC4a4klS9uaEiMC6o2YyfY8cOmYAZPBksMdKA6RKIne9geFZSQmMiif57mEFsR29F284jv
hJ7jax6c0ubqU8sSvrfS+4xg51JfOAU0kIlp7pn+wJx8UAzDM/NbmSVnynRV6sSE6o38wEH3j/SG
gktz+iii9R6OFQEU5enkHP5MhSte4POHCvmJvzb1PVtatTRjcRm2Rfn0wwQqwpI3DFU3D5QRPrbp
vEEA0DI9J3R6zLJrDzLlFI6sIAfCki/9Fl4ySFmy7x+xnUuwj39WSTP4USloDgNKS2DSTOb64ohH
wgMg90+ptmrYX66US3y/2NFi+IRDETtupku07riC0ik34HiSNxnd3ezO2pwO+a4Si4gjHfqAypSd
bEss5VQKU4w2rZPPi0+p3Itj7HrRrK803VUQus9oMZ//omva8sghYmphn65gkr7HcZWqXNfqM+YC
Y5JK2Kd0939xIrNs9HK8uoVEn6B/Ky/W1LudskRvQ1wk2wRcPUyurJP6Afvu1F+8OGdOO1cFPkBE
9A9dkkkfNh/geTH6fnvGnAoYBwTMbJGDqgB1lS/4tfrUyETEKWq9ADYk6tu6FbBGX9TnMg3wQSDr
ibkWw0DKGhpjeYoCwsba5w639rBiNUAKzmN20dKooD+YPP8WFlpivshVfUpZgJCASK/3TLfUyiEQ
tks/EJZiMxRcJNSffCUnH/7HToCgopchR5goDdS1KiIhkV4RUF5mpjDxEkp8ng8pgvI8kNZFCPO2
GOXkZIedwqPpWEdN0S8eLo5ISRj8immGHJciNNhu2fvbFd+OOfvzSrbLaw0ZaZhQPQlS7QOEjEGz
zjKtc9z8FJ8i2CZF1+ad+vqSInW2g4HkMvxqCNCYHJdQAhz922BV/n+AitUtodsiyN4TD06DWfUa
Pjy+VCHSQkoQQ7o3rsI/YnL6MytRUbghSM5GsMBs2zNnS6t5+qO5NCdqAWKnHXSU/ZUYGTh1DiuE
ZWXbJZMVPsgHx/BEs8Yc8t/3o8a60OftO73SOPfMRkDgznvyjhuBFJswifQBoFv/dJM5YQPjc1aB
XlEQFhMM+QzJGzpVRKw1eWXRnob3gj5Rfq6QnDkV1fMvE3bAmeagV1f+Mg/t8xySgJS4hlDYWI7y
MpgiunuRCFrQn7EjTLFs1QUi0eryxZarZd45gDTQMxE3OBAaPTHA33VdDbp30iZXSVrY5Oi3AQkc
2CjbaZy+NlD6kz+p34f2MIVLnTi5py904AKVJ2qNY5i271t6fH9hSMOgJLdE0YttbYju02Kbwr9f
cZzZXzfuFvkw5eMSRljg5zVcKthF2q5c6658hGMm/6UHqaCe9mFLuW6R0BI0+NH7qgIdSoDmmKuv
LjHVKODAGVkl992wU7eMWf7x8Mw5HKHKSrNiBHWhk5Ab2Sb0HbACsZkigWyKilWGdeRe/gDLE90K
4/MkJaxfXKlLAKISY3HIpOjhE5UKq4KYUdGfVUoJb+lk6PaSJC2jYzxRxWnEs4d0yn3zM/C6dR1K
3ZjrxqmJ4miQxvDz0EPUcTivyFKTZoGuwtOHsRJz1bzD416hUiwES1e8WQjFmelQqGSIVQ6pwEbk
rNQBioa9Cdir4F1wfzTcLfe5a6cYIawGzmV6nOj5evTUBKbZHnMJlYnBUsdcqyg9tVpOUHB7v9NY
9Z/+T2fDvaixb8odKxWa5aDFjAT6YLCzmJNbWswcdtD3AIqeY0pLMWX8dw7SFSkYu/qo4dKNfiZp
bQYsuwrIJPGKcBdr2Ir1COBALPO2vFQ1pYC30RjQKJjlydkB8bequqnanUbq7RzyWTfJm/ib2Uor
Z6oRXwetqMB5yQOVghD0gXuH2+WnfJJyCO/wh3DyGGlMIwfJX6kE/W4iOW6xz77+HYtDZEosnaHW
QW6NPFrMHa3RE5f5OQ9XIL7wZKwHOPzTe7QwCU10DL9lK+P1EX38DqDSr0PtJRxxh9HmALKjyMNc
xjpbmAOQNu/xrSgJ8crLokNG0Kx+ovGdXwcTs+ir5JH9u6kSIOJQCmCqGXzAXjf+7lSXZi19R+6o
XIYK87Sr+EDxNTG4jqP+aPzgrjjwovH3myDIQ8wUkh9P5IUyP5LapISKeblkujOlWPSLgpcdyEQ+
1fAwFLuj9Qo/Qdaiw+908gvdwBmbxyTr2mY/ayZJo5MmbH/RiWwUm4Cw3Th8BUeMJ6ocFlWDZHFz
f19lrlrTtCKr5rHEE/1q8mFX7cFBpaqWgWOcNQsvDj1SnUk0PpKS6WgL93tmeZaif76YaygJMs1I
iJ/VLvcvhTpn8c+SXGAkrG7FIJJjFQYsfIybBgtG+wy04hV6RYpDIv2jGo0+YxN2+0lN8L1L0kuH
qySuTKrr7wMYbSQSCxpz5lCz5CwK/jElFyGkVoh91LZaHRxlH7YNxsZN0NQptUf7KFo17DpUUZoJ
EJO4u2z6AOFbCfOlfneyA9Nfr7ZzxHRrRhbPp818A0rqwH6hrd1yDrZQX0vrhJ+rN4BpIagrXR6j
1S++2+LfO1hbE4wvxVUzXKbDKAdpTFtAqTa8Uc7/H8vq7Gd/2QkboghIMqWarKylv2Nt02NvcNpf
7lXz2w6IGOwxMlyXyxyNXANzDG+QEz3KwucO/FVjOFqhL2eWcQEGMASsK9DSzr+P4/lnVQYdWkvS
QxlFA70FMzld45XeJusxqoK16pcXCenbywf+tWOmwYrwHFXF8N4lOVrUUSsfYJ5ujt26pkHiRguT
oxPNq4DuIIMCMURFmlaT4E91nmOaxqooo6ISLyKz8PIUfSz0BMbZV0fbfSxQByL+NvzkePWF9ZLq
Q/+jcDPChLRWxiy+QxXNYMCbzPIeOWLNJ2cTkntvWSAjDdvXATyKLxjJ0gNcZurxHz1ObMF1/w5w
YSQhpmylQURl7GMV5JxFZglS0AJjhzO3eijbYlZAVi73BuwWTeavM6HPwzm2AxhV3E1nRjhP7YeI
SC3laP7yxZWnIT3StXO1Jqt+2X45H+Spui8EL6Y2QweBPtkEz7Xl5uyEGoayYCM48TYIc8aHWVC+
U2qXJi0pEALmEdet9ZLUg3l4dGfCUBocpIOpk6rGzH80AzJt/N3WjfajwwzGeT+tfirD0BurrFfM
PqpKmTXRLoM8UmZDuxu87qk5F2VN5Oto3KbratOs7zAP03kPAZ64VukpOkrWEYyf2cTzFnYt+2fZ
GA95LqVcggm8CQwahO3yE9Cztqr+Yica0Z2q/0KdVpPIS3RJqrLxj4rkeDzr6xikh+IISwPBGbyz
Ef3/GsLRYcr6G3e/VLx1IeggL83qptvWN143pyGgznXlkvQEW4O8KWzM5LjY0w5l8EHffhvt1vFN
BVYGwjRLyV70otG7fKIuX7/RXjP++6hlhmTzX0T/XnV4Nl09WrJ5zNY1/6BiN+zPWHExu7TiyuMd
FNUccxpEiDaJITuBlvFkiB3Vguo66LJ8yR4mB7MFB632z/eg8MzafEgqLzgmDqo5NCxeHQni9hMT
xNxa8dveqasCLNJojCVO5pq6ftukCAXeyIMTAQafEkLccWUKdNE6Sam/EDUAlesdcSiNx6cjd6Vr
17Xz01zIMjMySH1DkY2uG1X1hEjnBuLJq7btvrzvdF+lbeuJtCjukcVi3Sx4gV1rXwqqG81jy3MU
Nzd5jar7dAxrhAl17ultvBX6EDzexYxE0p0ZdqJcpy3L+1TMoBiofb2m9j/4EUBjAPUjD2sMYahu
jtd5u7gYSkk+2WyVL58rOtrjuBqOvCZFNDrOwfU6MQzVcGcu2te2FNEZiGAB/nlH8sFw9nyIaP2H
S1F2sGn0A1EAjHA5vxEwf9qoE/6f6ypyhxdOQTJRSwlx7Wkzrl2T1vP7tML+xeo+t6k/O7bpOn5y
aXpUYZMacLrYVe+jpQZ59/wGdC82kbaswC9kvE77SjonKBiRgOowaBaChr4JvxdRBlMxeo7TQmCo
C36PHIUATTgoglXnEIUaTIpeBtyoL+jf/3mxcVBBGgPclHazjspUbudTOl6e2/mcs8FNPDxoQXzg
2g4CuHcPUrcAr040+m0lTqZ2uY7hGGsTUCd87BihWusao5h/iMUS8rgAsttMvLKs6loq/ruyzZ7S
FIa2vTTNhV6jXM4thw7WDKpXvL/7abWsPf0YKkGlGp0fLu5AhSsqKH8L7J86v2NzrwOW0zQirhfT
B01TeeJe3UaNiomiPJaJlWn/qht5RDbk+OtppF98dsA/PahG7aRSAXUn9NAl0oG8BPiItElC4XjV
6357OzTsgFA7iPyIajle8Z7hH0tw7kq3wdnSk5U7/8EJiuAEjsibPBQ3RBo11hbY9kKREFgG8QTx
qfwvmY8YSImd+MLtO9mTtOV4DSnLITreDtYJngVSJ1h7uPG72v66J5F5ONuY1l3mnPKFdRYX0kZS
lzZUCgMbv7vi2uFIhx8w090dF/QGexEdegFCHSExoTlI+5Ngp8cMcFgl8LQBPHDI74brV2ZmrxA4
7zdxrqHgKXU17R6CND9tb0yjHbHoUn4j3FKll4yxvRn4sKnvR85+BtyhrDl3yGtF8wqQ+nUK2JIz
+kpP6JYLUue781n6KdyeEMyacqXj6GLQoj8H9FnauScsPbrwQO3yfTC60jw2+zDqrH6QuDE9W2XS
IImUrNMLTn71C98632zYg66hNsqxol5VYRNYi5ar06NsicBGnCv2jiUacs5c95a+i6rFtmSY8OwE
6ZwYTPlxepz/COr7x2xZiDVdasmaAaFg0xKnU5MjEZKIrAy/FtVyHsRozWByqBzMIEHlV5uZrXuR
Qv04KmRV9zZ/QSihSVHIP/6PhS/YpSHELB75lQWQGuBf6yeOWxzd1hEVGVJH+rLpWBowGN6gSDVb
MeXxc+jXdmUjH0B89j1XiAa//pc/j1ZwEW3Noc09u9Mtt2Inhv9WI9/3jRt2qFjiojsCHyK3eHki
gmk0m9u/S1vsKXhvuCMJk8KoWmtHXu6xJvN8VGfVsgIvk/rzXIK8+j2Q+eGsaNrebinadJWHrxrV
qegBKJde7HzjDb3qLx31dEDZJKzhwCl6s2tB80U9W63m5DRe2PYA/dWBUVFMWPshCu4vskMy46qh
6cyHsoiSdU4fSBx9Akvy6VKMqKXCGtbxgYbV96cbW7YjHOcogsnjc8SWw2sLQCEReLeinIuepWOy
BWVNOBaC3exRZdMdczCiaaX6LHUVnQCA20BsjjowuWC68jte3hQYfAyhqgH5rKHT64ofs6F5kHrA
9Q8qPYdQesZEwiJ07rMc9hiDCuX036RpXRTtHaWJHuj/twLZXJqMaEur2GHxfcwdnGJ29SC8wq/y
9BjH2sadD+vgYs4+goY41V2yZLRToV95DcQOEkjuZo1c3wzyhRlScUacaxFKYMpsa0eIZbn/3c5t
emUffJqT7C4j2ybpEXcCUAZvf1+D4QHcxU1nO/PLZw4qmZX2qgdH5hLiPFNsZaXGScMdaYpyP0vb
ROxwo6hemiRULPLks3IdvIMpSvHjdSPmg5QisfGUBkh0XxrBcrwxQ4QfwKTxT0IVGs/i7POsY2F4
qQah7Sksr9NxHZSfx59p5MG1wzzxBwXoyHH7jiBh2cruXgNMp+M7utGVInIyKN40r+kIMahNgZ22
MCYBh790mURZVhXSFonbez256z5LXYEc4sOuIuZ54jpSANKzPB/bcx72zJ0vVzls6pd/v+xofARq
+1OOLlAYrkLw8+hiDvxyw0l0IvHP1f2AMiaeVy8iPZAiqMfDbWfRtaS6sRchRcR+Eu+duUIoJ23O
Q8Jd87nlDCHNMTrdMzq2r0fAJfu0YplWZXWzVICp++ofZ8vnHw7KnAp4j4D2fCPmaG8EBJg5CGWG
tT65lJhuyk4JzJSdHENEF7P66xZKcrh05HDb5VklYC4HlXHqMYsF4oQ0H+VjObe7lerXU6Bltgly
ozGL6OVmBan+KiBjPP4CAcVXw3VanNd1Ow+qODJf4fkJ+4wJiXJHT+c7VvKInXmVB//XZ7X12iye
T9RXOrJJjRoPUx3+mWzpBf00Y65F1XlaMev59Xp1PP7/NGBFn+PfKQigNivwWeSFMmSagjNGMtqK
eZyoenKhb3tubi3Crgd/rfAnitRrDOHnnLLxlRu3wNBXI4aHRj0xA5tOy4XHooc5IoAZNu7xmpih
xFncP6UA8y8AlSXJIgcrJZwTUoTpwMgKsvlp78qQabFtiJFrt9A2pWyg5d5o6X3KEn9bpZU89Sw9
WqwM52Y06XbBttGU5hcthPeJK1mO4q6lhXcTy+iry/PUC4d1cf3bUImtvFExB3HvliqoRQxpqF8g
OD4g//70ORD9sa8AZZ2T/TZV79qigU5+T2JmqnGgj2sjr93gydOQCNXjJbWhBe7kOiPdvQAzeuBh
TwQ2hxLHLflYtvlJzYlzAnpAufZ2qKC8P4qdkyDCYasWaZdf8TL/OfTnXui2teG2qbMBhnFjq1Fj
wJapqEEd+b8sXVNBTlPPYUo4meEQOx4sZUhqrGBadDlEZEFcJ/WfEdwzD/1BARIi01IG5Jfp89Rt
N3X4GD8vnhmXtB9PJ0Cuj4GQ4wZmw455uFB7GHVh62kevdhof65yNfBC127+YUb/VdHINAZWU1Ca
wtC4E8cyNbNVVUNx7B/cEbljzndaJR0SVNDqN0d62A63QWJoOHSuj2vzZayFTTx5kbcfBf0Cqhjl
N0RB2cBtkJoj81uWitBHLiDooNKHimT0dZE1He5NikqUMxBnMKpl82+8Utrn28E++iTnivp8n55K
TXkXWB7OD9aEuArPKTAnziAjVGwGpqVFc5k7ZfkKYw9wt3M0v8egGFmN+ssYeC8VLVHMX+Gjttxj
XNAjOg2lunKlOAyhs8XYk01MtMT1YsNhHtIott8oXtuZd0MkeIL3xCfD2ddieDpP74VMUjYifnhq
Lmjx7jY1QuQF52YNN8WQDkTvJIFyK3j8mey/sRLxBL2mhIA56rB4KzI+IrLofuMhizwesG78FR9t
7u5P5NoH7n2u/mBB2a4g7xVn+BEvF4XR4iaZYjOd5Ozf6bl1Fw78j4b9qv6kitahAlhEzqAyehJk
PxWEVq2bEgUOSqaeaqnxWq4mL9kZP2gBPGrIOM4ynGZRYNfg/F/8CS1qGAe8NjROrTxsBVwxk1s6
lluzWB36vN8I7+B80kYs9e4OnZ2XwQtoeBi42ez5uXmGHUgpfNGeHGX0yKA4erp6qy3kzi7r9Esh
CFGSBbHOMvSrN+EET28h2YZSwqzOYC3pmnf+J1r7Gildo0hKX3uVhICdFihPe2g3aWCf24uiMtrG
6pbpoxXpDSo3rG8hEkKNowsNG4Gp9HWXdh1zI11niO4fUAZU0eFd+16/lxVDBoCAj5plTAq6SSOI
8kdmA8KeCdKUlW/hSG9Wk/sHe9Uw1ZwEX1TM8Ev7aiGFdy1c8WgNoSMLTuWfBoEJz6fegU4qHTWZ
wW9EAwzjop3XX2jKql4gbeeM1768BxN/h6StqX2DS7asin+8s0il+6uG/QvnrrTg4w6bKfWsaOUs
tqBzMHMQmhqsC0Zjn0dpaiYLIMhGdzd8dp36Whgc7jfZoBYUXYPtvSDZElDFAtUkUsQijzBWA8wH
OOzw9ui1M1kZOc42JUVW7kg+/UxRf+KJMJtcuJkJ/rl3ikmIiRu17DciQCk+wziToS7X/dA/GiI0
YMLQTZaK/8QxHjG421PmbwB7/ElZgeNgT5lhdUod1wwk+O5dAXiu4+D8fWV7BUqCYfWiCt8hyG5b
aEL3wtf3K/Y1MVNln15uob9u5NBucqChL9XYIm3HuAIxM7un8yPo8LZnqvVu8bW9rbOwGkpH6oxJ
4Oeke7yHuact4tNsEaar9RagUNB2LPDFVlVYR/S3TibXSoVOiJkzP+dkJCW9Opp61z1CpeuJa6e2
iigfvfX/QoePxqNrMMXE2L+otWRMymMCcLrlzybQnos0wKEt96UOE7vS7rrgk5bHJXiuNfXr0Xka
MqRINvmXKd9u/MxcfjIsY/1fQOPlFKt7qFhH/UYdXmiuiqezDpZJMKV10+D5B1rQS9UqJvDR1gsg
i7i99XQGlTR+tkgFHZ34+RFEGqVIgnJY6BvSpaSkyxWxBULAtOAxcFJpFEHdaT80judsUZJABHyj
NgN3WstjrhVYSGuIhX6mwHUcCajmlLGpML7NoGxivWsnZoA981YQnjX41P/EyUZ3Y73284Bv8wzH
dCXgx0EmRdPOKThx8I+byuV5yVOJFZedBn+cdoeYFLd73nNEyRb249o5w9IreFoYVvjnIoibI7dO
mRDaGB+AdclGjMvhfKzDT0u/WwT8L5YwQq+ULaZ/I436MO+sAAnkT0gSrx2abKGZSE3jXY7WT7zO
tw5JnyobxpMWYVO5b14KV+IotB61kAbRfDlx2iQL7FwsuIa7+fZvm5gx8z70aS5DXpFU3iyjegpp
plt4mV+L90eYZiPiGYW8/CerHSlFhBS2jthmDQ6rWMqlwYVYcqCWUXd/bEns8oaYTPbFFVmCeG9R
AqZIIBVLcICzYYg+66tYHOkdj+mbE/k0MCaMhm5i4ufsEzaQURxDx+RhY3EH3dM/s8PGahXFxEV/
KE/H+awgNwYKwZHoTJmrgWplV04wKLEp8Y0LXB7JBSfVDfTbKso+PK781jez+C4NtDqHoHyndCST
rDaERylh0TnwGez7VADPxs9nLmK8XW3JCTzfpMBtVKUfjBQXR7/dLPoGqSRjEwFuMXIJr5aq8OEY
pbORhYoVj8erCga+uf6H3N4kTPjz48QMUrmV19MKO3qaadNXPNsFmRTRtkpRuEuS2QsHTJavuPrW
XgwZh1y+DwMjxfLRCNUKtLEQjfv55Kw/NxZHHD491FqYJyxSrYKIhJ4r72T00upm9jaNmy5B+sRC
INUGTqaRId8DQJ0z+EtkBG46OtCr8Ed3aokfhCeXoFmL4Eb/iZ7EB0lJ4QaJVjY3da2eJgBYY9oc
KqjrRY2YUhmxmt5RXnjoRH19IB/YZMpxdXVU0lgOssXOjtHjELvqNjeqxwE9rq7buLDqPlFQtfZI
XDzbYQL8dDgAGs3Sk9tXIwR7YCs6Hshz0hEeF1CikL6uBXpKtl6Icez7MKQ/u6tjBz7S14g88Lki
SpsHVyFUhYjXyElVlD5y92X4ceir3fspLmQZ+tJXM+sp6bubcAOtVUXydUyc+rvFu2CbCgfDJYwa
xJ/wbs4mDfF4PhEJxG0wb53XAobK3MjC34DBpWrv7P9rtKcmx4BTyHpIZ6XGkKJj0Htd/Kv/vClK
160ks+TPinp5RnAPTScZUYqJTVlTbxQTZ3mZ0/LoL7v4IQ3lQKY2LgZKjBAlS/CZ+1emTxDd96Sk
v1EStleZ+lJeVhb/Srchue/JP9mPnkZmyrSaluUGhsszhLZrof3tM5g3JHdQMWEsesDcYRRcRNbk
xhi5RkTevcZD5urDE8/+0vw6E6IRrL4bzPd0gSzrQaiJ7Q6afDYRMdUe5S2MxZRL42+v5PvSFt0b
EysdapfxsaZfRMPOiCYiHpmJIDTOPRi4x5IlUYVDmInDjrNtHdorBhFe/la+nn8n4IeGMzD1ZeRV
nk3mcwDpd4lsy+e9Ubkqh1GyvqdcjxyGu9QQywaw3zmgLpIdY6VuoA7lQAa3u3ujRDVT6u14wfQx
84S6vokQq4GUez5UKiEHLmMDmHKKNAeqWCq1nx9fR7FFqgXZh0Qcmo54abPXQwOTFSHXqgAh60vo
P9io+/ErpAwo06Pmp0oqDoYGWhjF0+dspBUGF0mGI1uHX3mVRe6QRQbdD5i7XRl3/eY0GE5GqzNp
7Dj10xwVmAWw5y/a3DdC5lofikmMeIQMMU/VoYQTW7F2uTo5/xfBi6HCfQ8N/tpSwj7fV6E1IY/2
8IMZtMCz0sbTrf1JSDny/5BPkHUGUAoTvMmimSzJizLh3nk7eV00TmjRHY1u9vockCeU37FB4tQg
FZVkit/NjONdmCfjIggcNeThBTuYDDcaBDikpIGf5OkoXVk3RnHR4Ta+wQGDKuleG0/Q73VYZB6m
2Nm84VkA8SBxBDC7geXnuIfc4n3m2RMfHCMZoi9zIykMl7u2BMcuDY3+6D7WVERJ++JrX0S00pFK
bdYwD4+DDyOJd9sXN0x1VAcmKlsvky3gyKjT6NgpA5GBBYt8UAUaiEzsIbJ7W28fHbNI1EMgBbN1
OF8rpFjf+cq5w4JGwIzhZrQv16bFaNeBOOYxebMDah52zgIA31m242SDTmXLIoMlh9FoPH46G8wg
yIj+y6TJ28Gm4qLByjju+IOCC9U7sdFm627nXQKWyB9//8tMeDIwmv6OWlAqTFZWXjT4LMfs424S
xoaRDzjdTN9PWwtJeNs5VXchWaOg3fJayJBWrKiTvW08hRaqNSIz/mvYCeax7CMe9dK5fTsM5oCN
c2UV2YSHZQK17ja6/fEMuFZ4DSP9UOhernth2sZ9awJo434q5/FbziWmy52mA5w0Sl62+yVzeHen
DA7XWFTyKJZJHOEDrlVy572XVXC6FlZ9e8pMuviEiJCVZINqaxlYAk+3ZB7B01ZXpIJqng2Hv1XR
3xpxudnOpc09CEeCmOXLZR5uKCqfUYffb+WPLZbxIj2j4v8P93Bn+TZKF5p76GGK6EMGC6N++HrP
0FQAwpNchrm+KhV3ZyLRk+Vn2M6+uNVavA7TBOHdCJbKm/GfkSVyfgCip3ROJMJ0NMh1Hsy+PrM9
f2pj0ulMmv4c61MFW9hAm6y4HHvVjs8qSp7RE5saDjIKDtYYDf1XY+nW7pi18TtUovlwrAs+t3X7
rsVDk6UhJEn62PXEaWVvDRdJsQPankoZ1XAhE8uacX5ONb/bwg2psoDAHmX6Hqtc6pvf69gR++fg
5QVlop7waiKPDFp+7q1aB/d6LnXqvYzPFBjmQmG3olcRgO6tWIQsRF5ZOJ2UnJxnJNHzJmND+rAi
QPjv+V5GpKHUM18Uu87Ei3Hy76Bsm/tyNoKOyLPuV+0EXnku86CUra9YH2fDxNI9YNdxg3PIojEl
yI0ljSnY2UuCKmntwUnOZmqhq4jq7bC/NwoX87oOYJR10+62csb+wr3dHFm6hhj84WuYgf7fkvZo
AoeqOoaY1X+h0CMO5N46CPfjJsVp4XcZ9WSRGrBibfQDTDbuyxJvFzRC4HcntCm+2HMpVSn4nItU
cPx1hEEhFZe2oSz95h14EAkIovPZsDS9IAJy6Y3SOcU+fKCIEvEu4QzFS7AQr4l9QcihVVasttw5
gamW8+ptMQhSPMbvlMWphmN9IDFHHoHZaIyZkBjl1AxrnjQ2wr25X+ki/3egVDcQ2okL7gc4bLQM
I+ZOUK9oATVtbH7zUyHPkHQacttuCvf+9tXflENVoTR+gjhJE9PoeHLkCAJ3PNYp92wF64zsCiV1
lps0RaqfX+G0lL4fzR2xdbekPqZfOqAaApKI3ZIGnGB7+prsqO5vTiRDR1PuXk4h/Dhl3c9+ADmJ
SEwAx/Z/Z6J0vn1yXuTep67eF/0AqkQCGkvTeN3zQykw1hRQ0f1iqmfkktffYcZ3GWDuMLVhBE6y
P0IFCoVeXsd5fc/drNm6vdXkLQv885qMXI38gD1p7ryYngFWxW1iEha7h5LWSmv0sUmngp/L5Jxj
deEnjy9A5cw8R7J8aDsACmjUKG7+ISJusof//7VlDNLIKFr+hUn9B9BFwRsZ8PRe4lwrHobAI3lp
UPGucHWv2fY6tBhXWM9KTZSfygGEx0apSHYLABX7eJqBYEe66VsKtHPkoNTlV7A86Xz2eWQ5JFRl
2SkpZZZQr14DsQ5uWV4ogDd3GmG/YFePu2PqwNHrTmr0ypBTS+K3qZheJRBbcZ2te1muBvroHTLy
s+QlMeKKqvyjDb4/MFc01sLS/mpEFOHz0T0Iee4eieUl/QLFM6oRbblg1wgfY06UkyTI1G0zhkkv
/3mI4CdeR8SFnHhAhGUJaL406GgJ2uaPg2tr1XaoJrTsLbds1WAj7g9d2upSmgd+dSlU3QTMP9wH
0tCg/XL+dd1WfBrRfmsGjAs3ywsg1b9si/ZQVAj+eFhYuRxRuNEzrYxAngD3WdqcrmhnxLDEmG4s
+njKaoqQ2cB3Eax2drju4R9NkQ/udSCezYZIBjfEmX80ybPZjUGBpYe7zcBoiZi2qYBJOqLkpxuB
Q724PryCynj4Zf3Tf/kRfGOk41jIJfuNZ9egIalkNvHxU6AWzcO8urCByDhbGrDzEHTfo3CgbqA7
ZVXFErf7l2QJAF+Kd/5PhQ5slXqOFpOzj1StDOT8eDz//tDbMC2GcvuuLaMovRdxGem0BmIGJYKq
GImJT29CK8yJPDgjODcvHIZoMjtv7ZE+mdTX/wpU1p+f8VRDaLS4Gr7QbrmxhKJF/DpX+s+3sAJD
oBdrIGlXpANMRXwL15NmOI4CC9V/6iE0/tpBtuBb2iYN1YFbOHuu6xrRA6FP9Pq3M853xHfKodZg
YUMy45VNycpJo4zZUK9XRqe9a2ZKC3euDK9HgsTPnNsS+qoxkEn7AQZHj/0DBacHJRv7pIA/y0K6
8Ydfx0iiC/LWHhoyS5XD4SxllROjMsMfP7+r3JdcCBac/9HGieMmgtO3NW+P3OhLOImFkrHUTaAc
1pH91eI1r5KVp4IXrArWEUwKUPtQKHroSw0OSUOF4vRMr0NZ0m7aVuzHrePIUCKmr+TucJvNtAJP
GTj2WwXe0KAYY84gNgijnNCJbhEH/FuGi2lAht3vRvueueIcQygMRCRDzqpk7wCtG+nyW/Ui2wxW
K9ItVAy71/3dSomHzr8jCASvbyCtEYrEWbR8paOzCKQjZESMZFFlZm1Tu9TmW1znubs7odJomFr3
pK41Yyeuy5Ym5NfASwzx0nPjNBeropnWG17nDptCmy40OJ50Q/B2B/kftHFTN2BbTHpawhg2hNrC
2O3ChI/TNbmQgnlPYIh52qjjzzN916RrAfyYqnnJe/sC03d2FglGEEbF3QLldk9zgo5VNAC+VVqn
1fMm/Wobr+FGXll+Mn/cmhkCrAO5EUSxpQKGCPlHISujaxDByIOua5YMgvL95RD7K3iPYpxGSuR4
5jCqKfBOkofGoE4WqZjnbnRU8H1V41sYHEYghMS5STi9S5P7nioT7m3es6aYJmNHkOJGLM1IlVwA
xZ3eWY5QnQT3TVf4oKXbV9XBOhRVCX+j3YSWRZEO9npc3YVcFsrY/Zf4udqRQleSb/tElXFSt9Y1
5yWmiZTXyv8VYyMDhx0P+ixvwXkcHy/nIn1wI2x8Vvsv1NfRD+mZOFhVhPPBd0G68MrS9bWVxTjI
Rm2z8UhBM5pooofdNrohNTKUxFr8vDdJiaeWzSey8t3e69pBh75H4mV0iFgkQT0BzdY4AA91VsSb
opEGKT3itakQwLXt5rKoRAxGPDuSiLehYxM7mfj/21glfHgq8KZ3fuescNeeH5HBkmDlttb9GklI
f48juwPwVHS8K2TEOh9LP0T7cGJSdLvwkOQlFd7xwcmrFWyxf44pOOTTAyease7lHhZbf5WtyA2g
pW3Bw1RGO6VLVmWnfy564zUV2+F7jmQW3qetzjyzUQmQFhNiKM9wKoj59Fw5dSSPE919xeiGzW5y
JJnolrhVIuDTmzZkUj9rid8GkEf2n3HHg6qlbM1N9Kl0rnF7/F8/ZNWIIe6ihevpHsd6MLOVYWFp
J/Gi8MfIRyCOHRM7WjSPhcjzOz5BFoeYup/uK3d4eKBX33nNu9iRpSAMt1lig4tht7xNJADhcXhd
Q/wKaz+BPj6zBePjLla2dLAHz8RRnbsKm4/v9MJk6bquPmR0wHhrEnAO8MoPOQ80GOxxIscgPI4C
2/PofyIzNiHHX+1V23ohrMIUy0+tY3Qv4PtSv+A8TtOTd5kB9zOMCHIpkIkTbinmlh9JKVix0/Pw
RlfG8DYzcMyiaTjTHKR9eH4ccdAcRQM77vG6TxUvDzExK85MrD8oXOa7/5xsNfcnniFxMZHWuasH
oickagzWK//LfFk2Pp5S6YWvzBM8PJCKRohg1mbV/V43/DXeRimsmCJRNaj4awgqdW27RsUjLfBS
OkgePMmFhp9u2QKHn+5jfWpay5QxqMyEYdmslj3/S77d6HL5VG/a32zZOdybIyxmmMB5Hx+kGd8/
e41wdhWIbhWEfFGivHcwGSBAkCw9gGuPzxRIxpeduwaGj4cIG4jrsBImgmvvr8hpkccTcsl/+y7g
PRFG+hGu7vT6cf1XdIaYkwbza88id6bYNDyWYZYDx5397qsJ+0DNtvbPB+ezZ/sKDg9RAWYqeezo
UeohofqT7wnA3Znidl5YrAzu3QEai2CwZBrjbLg88mW36lNK/jbpyaMzPKNF7++VgdzFCNvAIIkw
EHR5wEkCE4+KeWuwTt4rtrr9x5LXs6O6BmPt7vaDfLucMiASkYTqvQHZoLPt8c7q6a37vws50fYx
I4MbD/Savv/W1mZCog/E14w3NpfCLUHNG4qNhVb4mo8vzdxdagMYP6GRmqAqfPl0M75YV/LSjdNC
AlMquCTqJOdX9btFQSpsQuiWH3SCirM9o4bataxA0yCrCBE1ya2vy1ki2MnveMeZvn+CaWF+SDWJ
/sokuJUhf27b+S7/aJ1+JpTxkknipbyZMwAkH1xI3401NDQhpZwhiYUbLm10hBi2gE2PxVIVmG6j
8HaXCEqJFbNFDOW08LULHn03XDEnqc4xyHVAc8cxzK2Qn9yIY9YXnTaZtKO8IwaXdPRE7zabEKb1
zRTLsP03tNWQ3hwsBvJJGW4VA3pqsYOMw3Enu+sol90YhRk5FmphFSM4bS17pYr0JgiW7OXksShc
OOxublzPmBT59M60mXHgiXL9F3sSGNTKTlW6cNhJCImGVvuNXKr82ad58a+qmoHELW5AlCxYI0Mk
xCFsodCzgfdvQ57kSjPRcy3yEHR2Flkv++yPGsLnBenN7zCzGGrCBJFfph65gGy6XaLzpBDdaP6P
3Gf4OGvJ+gQ9tByD9f3NC45obCvLV66RDF9Okm6U/JkaQtcH7vkfBeFAjI4eY99yAZz5iJqi0bqb
91dVDddW/KVzHCUowkACtaA4orPIYeoPHUZWmWay1L1IAbfPJtIffT0GLezZPEjlS+AcfnTbAjlG
4QOgJdB3Z+C0ioJgVYf6qSmiYPzCbwxMiys/KRQXeRrM9FnXsizC5MHwu8XAJeYQjRvqGq9IfgOx
kavt3JCIddx5mlGHvgcouqb+fKCcs0Vd4pHkVlrBDH1j90gPnQoIX8oiVg1/lGyAWE16tR/o8w0u
gh1e3P1jnEnPL/uRZZpYgqkx40hHJPcQCZ0A06SwGzdUWtdM/i+BMbkDvvJhYkQWxtEQf5IoWmcb
UnyAg6E9VCM2jOy4lcKFD0LYwo3RdWuSqEXzibcFimlFM/Vw+aRkZyBXkFNYxFN0wyl9hCW4QXXi
yuSbL1fGwSSSUiewHTSUQ/EHtpETAB2DpvE+xYS+SEdtYHkTJnOjO1CQbLtJRXhRl3AaMWJlgF7P
b0Wk2vNPdrUg1xCqSYGS+gOpAtfppntmi36apSIouxKVJyOeKqy2lmrpmfM4mAr/LKsrc+UuCpQD
sNt8NqvaFKbxOrMr9XPoD3xzbMszwFdXyEJ4QHwb4vSJlWGx0gNfWte4JBzuKf1/Frd+i/iSOYic
7rwJNx6A2WPSVXlm3azp1dxe3jgQjqEu8GTclQvmbVJOX+Vgd3gWuaNugfkzeTb8cCZgtU/BPypt
klnEFro5AOJ5RESvqbb9D72/vqieUnJSq5oo0KPxVpT3ebA+iCt2ffg27XRylF0z6xNjs9f0iNQg
wOARguBG8kjC79U8no8nlihM4yFhU5e/oqEpu7LahZvXNAAvSFg0NH0dfwWBcAfinfCdTRJCofCP
J+LdmfF46+LeiPgwRCJZn6eLIRigT1M8pbZ7mr3B1FpcNP+Eha85Yi/geveobYLeDg+KmS21zusU
SfYULewSdIeiH5mCzqUuzA7kknXTBIsVsErfGQh/vWdp0b3Tul+yMVo6QmGmUeUAUvlYGIrtUwbi
poTyMugMpripMv1vbZPt2pAVhU0Q4UJTZf89MGBM60f7i+Uf7JM1IicvHz6X8Ex1quSH8A+osJ1O
cl6umdrgE3Jv+w9hZRMa+vexCdOykYShR8g4T4OJy6h5Zu7oSjw1f+yWA/muttMs9kM4ux6xaOro
oUsXA659AkSy2pALqvJnZWnLapbDa5veNcnYmzBmp/pBFNVjzVv9srhOpOw77bJ+G9WT1iYVnm1W
2xkWY3G74Mu8RmYgGTsK/+Z/iohv9/c1caEJw6rjPTzrfIRozZVKjcm+GoA+UoTATsW5V4iuZ61d
VJSJZRaP8WZVOqclbezBVBybLEeU4uJEW1HBE4CT5vEooa1aZgQ8XsdY2IYi5Wt9hBnQLQKoUJR5
jXmAq40rVQyliqvHnovbIGzH0mDKqqQdyaYrwj5Tbm4u5l7A5vGxI1MCbcc0GLGrYpjNWvXmv7ry
K9wom9Trfx9xhl2rWu0Q727USonZGPbqySaRTfFjEMe50VIfiRSKZIRxBZxrnkukbJnobzT19WNa
xokSm7tZJIzCEn3wfbPEwrpmLLeFSX5Unh4zIp/j0bnYrJcfaA6wIu5AEkOi/4TOyF4dQi2/ZfLV
xRs8vfJmS45kLfOvVZJO48j9jLFdPYlBi1p1jjzZQ+x22dSS50VgqVH6UECVsmToF40trU2koenj
6AvFaA8eBLFb2cAtjNuNoHh+JNYTRSTxR7monrDWA+id3XyzPr4RizcK0L1HGa1cvBFaLNzcCWE0
DSBTPbGTa5N/vP6I2b+s0917pHX5QALTJMT1NgKfqjV12hRZWVd4d6Ze4ZOs9RhXMf7JSb1KiQyQ
qPI/TocEZb98+DMX15OXpOqnXrtzP+uxrwJgcvYeE7xaNpYZxMDx/VtVOplzo1VQjgT3kz7s2cox
5qm8GdGf1bjVnLTh5WV66iUEB5K1ckByeL4MPpPxqyBNi7CWW1tA13MwWpzcejQ63OIi0NfrmOZR
FURYsZUr6b6Gi2Q+CWm4BZ2PkIRxyo58R2ig5g7uZZQUqHX/g1MQibiacay9xvMZfzjYSqzOrs5R
HC3t3NNdioWwqBaDXxKs+JrIpdbmxAvU8YdfBZ5tAlgC5eZlfAdIWb/q+k/I1HHikkGILG2Fsj6Y
b1WhekqCYsIVC4IEHxL1Yi/TN6F8gRQWLGBg9/btirQVrqvR5nWtnaUInqPtkzqGl4SV/OevdBvg
/jHT1XItogdigDec/ZFH+300nglsIUGFPzfVCE9vQegBS1HwqYTw6TxWeesbAKSCk7VM9KZfwSKp
1o9VmZsWYifhpws4lD32JDfXWhcXbCCAe2cuhQJOo0IcTA1a/q+MGAiMaUJMQhpH2H+HZyNwBWh2
juh68ohWVr+SWMyCVWKPgq544nV34WQe3P4Vpu+BP0X36EGXYuU4/eXpSOvUjlZXHkJg2qO3h1E7
IWiCiwnKkBAUufJNkRRUkW7gI1gh0y3+V1t4bozq7ePbG612MjNp4KvB6Mjult7kLZA+xDnbBVyn
bkR5E2HPAeEMKdxrzjgO8pbC116LvrbDjwprmrkTdWPHQFzYfZLhJTqFXy3IJqdwbse8q5OaW8J8
UZsi+X8DfF4BjH0AaiNKSLIYrV65Cmg3RgRKYiuyjHAIYzi6/HNRsmj377G/JnEpj78ZYX5WA9CZ
8f+J/gFe53jR9v7rjiSFVTDy+WKghs5OkWNdMTO0GTfV+liixlg5iqvwSmEMhaP1nXxGp6QpdXGr
4XpFW0qGl6amtcauNiN9hEIJuF8ulAkyWcNE1DkD8SwVvXWIaD8kc+npQn8UUhs+erp1dNQ81HQl
LFEuL8xYUzn/3O570hMeZS7LbETO8nmQqsSmuzL9kb2Vnk7jloPDmvVI0gslefnu2JqEoPFJkRPz
77yFpFSfMtlz/SPTuAkNFOE5YaP5aMeTzNZWeoQVUJm4lEylHRl8vC9+H3cK70VoKhjLOpMHMpsz
pWgoj9ot2mALhqMz5Qa1dJ0GsUciz946dso2WB4WuQKHOJ5ezzWopfV2ncU8Re155dJ60ip7qJ8D
pKHZ7nEqGkWA5Jh8A+6YnI1U+VFzxpsj0s6dUaGVMpSlqq6+fVWt5PGitMBd6DW2Kmunu2yCj8Vq
R73SfRE/XLhw/Sj3mFtCdYvcLTIXyJemPD3gzj+zEXFbO3FLyvN/hgP9WxvdsURw322qdrgDgExs
U1PRFzcHuPZxNokT4Gx8//21te7Ir+uXBpY3Ut3RFugSBKAIPkzXKFsbCnOc1a/74+vmqBrdcdug
SmxQeRhVqivDXYkUnLx7Sj8MKUO7TV1pkfBu/kEoekn/qrIbk2F40z3BH8qwjqJ4EJGP4yYAC2A5
pHYQFnT5YQqhK5uJXhMbqex189yT3N0yA7KnOiZ19u4XZ7tv+DNykq5HScuauKyokHG3lWsbvjYt
jFLDbyUbnQ5vpjgz5TSqzqvda4H2ihBn7wHrIjeI2bW1V+2qTRSswlNQKYMfpV2WzIWixaLIJ+oK
P1AiShU2aM4fkqgOg+ShB7No0B+ETdXfzqLccyHTP5LEbtUkZcienWY6c/zlUyBa+x5+ibNlImqB
8x138dNg77nTCSuMN4BIiJtCTQSzCjxi6XPzjPayqM/oAb/fzeFGuIW4sS/vB7AoMK7JFOoJo9D7
dKhHN0xMzwmJ1n6LqaYysXJKw1Rrps+UcSPn2NI182rq7sSCzyxQwhnDQB85UOwFdsL4yDTthWXH
N0nk32UDHxCd65IZqk70efMbr7CnGmS2w3C4DN3C26rOLQeuHQGKJ6fWEBRSfZQ+gsy5W4FjsJYU
As2m5er92WqtoenV8SiXb59UVb2xhbpjobK0F+GoJdjE337+c3U9f68mDS2j1Fx4ivaI42VviPy5
mV9D4Fj+oTFG2NG8Ww7qmOwQO+AyG7MCtg5kDTEBOzfzu3X2WLHCR0BVYaJrI4YJ18vUTXMK/9Qi
VQfUjThqRVDM8JHkKPiwrwDo5mD5698W05Bpwb4xAwramhW36iNmRI4g4x01JPG17JvVO1DQstkY
uFkxw/CsfV+2mdBpPgJD9l9Rsyn/LhA7ujR7viJJblXnC+sMA1sx+hGkwJ7IcFoUPl3aWeFUMbCv
hRw0NBsEozqUV0HW/NHgYs4JAaYw0Ud3p6ISPCMbMvbWBU8b4DXtHPYXpmnk0rRxfr/HlCj0XT30
UOQA5kA8uWNdF5wDXeb1FKBUJu1pfrh76CMZYmPgmTV6eFHCp9ueboGxb4h4sJg3hKkTk1MdqZR0
0Vq4CzZY3L7SXj/DL1Mk3GLVpbiKb+d0U6+gC0IuaNecrupjmkHxrSRAaS6H0jhoFHBjK4ARCxpF
OZFSbFMjNzMQAqdoB6WiiUj4nesquypYw6D1bO7rQ2BKJRy2SaTTFQvu3THLyEtswc3j3Cujixgo
IwYhUqETXRwaa1vv0LbukPWWprXUxpRpWR2jvQ4G8z++wFZPpkD9HZsHuaxJXJ2Vu6bJ5jHFleoa
gRGdzRbCAe/TcHYdXw7ZQZQ3+lHgRFRdwrsa26Gxw2eRoQftp6jHm1mQOBUszpT6/Yc49SBklDiD
isekybzMLQSUEfqG23W3q1C8HfdoJSGVujUPoe2jrkFf5zU+EQIIKBXKluDvhc5g9GxWlYGOg8Kf
RiFk/sRCIDqFKqVyXaYwXx7QjZZPxwT1WJokrS5NxHAWmc7IX65+7tLDFEwCCJ5y+zPpCNO/zfan
2964DUgVjDQGhFY+F7yFE6rpHgxylxrY/YSvPtbzp5M0q6PF6sZBNnQIbMbrYCigkN3o6C1k8ERQ
9eTmlhWi3ouFLWqgTM7NfLqHv6ksDvPvMvawCY39jLPMMCnLsEe/jAOMlK+R6IJTfWu1dAhEU/Qm
lNBkTV6I5dQwulRes8/DonaeAJ+IrALe0kNX1/VleLcg8Fle+wUU2wrDRLiHA/lktwHQVAaSm141
PlTGkAN6l/9ifUfkJIAlaMoi2ai+LYrFe8KC6Bejv/iaAtkP08oOIZZ5GcKrTa3Ci5KvVk4RTuC2
My2Ak/n59PT3+FePopsbGbI262PIUWo3OZQbdW1fdTdTGyzMsMhxc4NckaNVVky0i7W7FPOrBXX3
7aLu2hoPSqlyy+wIrb3F8LderjhfF4f6ASr7XuaJBqijEguZQVVoAwfzMVbUJCvIKgIpLfjobMcr
0fsnVrJkndfT+UQAWplosugygX/IyP1n0+0DLz16QlAKL6azmm5we4Do5sgnzZqLYoEUgdlwb9s7
gbo+D4tSIBF7fV5WhdURlbLUXmI2owwJ4eg+Zb0lG30yyzff6FxuXJhy+BZmTvV6+7W12Qsy2WSm
12kfOajHKcnn2RJHQ93NfC3V1SIWDqLJJhYzl5jgNapvcSAFa6FBWPrUh2JK3smNEhjZ2NJWD/v2
IK9b4mLviCza/QsYF6rs9v6L54KTbxaE6hImMOsGMPWMBWekC28QKem/V0X4XJVZd1O2DqfIJbdR
Xc3C0ZEO86oU68Rxce14y8M5agBd8taeq+2glTy6/W673a9Wn/NHEkZdIw7cTHwiI6O466bC4Y08
UPtyW+vN9TZbt35iMPbkm/zOnjwEzNRYsEmroxAJXEVsAKN3/i5rBGPrpjh9NdFtcvC/zo2iDR2v
aU76ggSyHI3qYPMhgPC5g2IvA2jHGPuPRNKqBbJOKNH/tdDx+WUuVZzOlAh9y9BoBxQilgXOTGE4
NK6z0n2wyFaISjFoyDfUYPudtLEJLkY5Jy5+Q2XBsqRd10TZ4ptymdahwcjv9F2og7x4FT+0uyhX
WuTx4/+SHRxmXTKuheQio2uYyEF0EPKNu4edEAZkt9SG07Y2fZRbfs0rzdBiDJlQB/VRLVNdzPEm
T90pjM1YZzOqotALdgRHkOg/Oh6uynO0wFYdLXqN8tap+3Ie+wD0Bi/kkdP+12bE4cLL4ZaKC8Ex
paIJNpTCQLgY+skN+hSaLQdoWyd8+id1DEgu1j6tycF0IB6JY50anFBQeeEsW1o/aCr4iMvgkQln
iqvfVZkKtlQobkR+okjstZUXHXSxGTF6tW2FnsTV3CjSfXODE5Y5ttky9yH1oP3oFwC0NJs/o/bq
wQM0CgPOvGYT75jBXUsibEtkxzBJ30usF36X416abZnWfPGH4LjOlD6kdEfQPIauJQINZCHEmVJ6
Xpe3On+WUZlDpVK8LLpYHveMtIOqC3Qq43v+NxO2qq+Qgunet5gdcMtp5JwONvXspnbh7acy6tCY
dY+EOHPIVkQ6AV1mwgPHBBDjSPOuc2Jddq5VCOkSmG/6QqS0AXiRDhnARrqOXr4b4C5acybLSDqk
7y5lfsmUw7wqsyhJUf9UVmtU6d5a91BPXjgZMN4aDl7tNTyWBSAwVDPx5RLf3WG+ivTq9cd3F3sn
LyuCKYVcCxdsLKSpCnsD9Pb22gf6AOVcNOO42tlh8qvvGE8PoUpHyqBvs/Kz3udct9tPo5fdWgy8
xS9GyFk91NKaRdHYvPWRcnCx1hmQ69GerirFzEPgDnuz5/6kLTAivn/NQN3b8FXWRpkAfk6pfK/P
5PDIIAIUizJVkf0Oe1B3PnKVF3EqzXhHoTvHTFeZKTi+IWkG3cJmiIY/BwKDoU9kCCXn69Mvaqbu
mqjq1oWmcLf2tH+fUT51pJhO7P2GSoVxgpLJb5+UsNDq3oh3p+FSNX58uPk4vn/j3GK5RCJnQWjM
9imhd0US0HAQ+dsbz+q6gvvooH93Lot5HOSwlBWRC4dkDTw6P45t+/4fSc28+Xg3MjDHpGWzA4LZ
ihaid9CIgCrSu1LBV/uLbL60/61EkFBbzsJBHPYdzFZtMqx5dJAhi3FQGKLSqhbIskrbqrKIDlGc
0tU4cbITPU+sAVvpuDzdhXYUWz7Lrkc0wyEBIroL3qzrPl6IKCVpfPv+3p2qCNoBQAhwOkDlVern
K4ZJJ+2p2bWhXKu4XKmVtjUHBXanYDPHZuo3o6CMFCH7ZnzXk0WBRclTdrbHzWeR18LjqjiCGGws
XJOd8QHpPZxvY4l/T1UwGD8fE0dZa+zRXoBJerwvCBt0RHw7dsYEEBtYL5IJ2zpcci+S7+NmIS9Z
4WKvH3YezRSbtNrQ1nZiB/2B3ueVRNQqCdNcxFXFloT0Zj5a7h5rbXleMiQdMDqiXlKiZEvq1vZs
510qiXUrDoKi96j2DOc8ZDuMUjoE5hQQj3/FFZSFXcjtDML9HO0g4sO6mp8Uw48a8hxmRntehm+N
TQV0TAd6zrqCcZ6y8DgSMJ4jyRKnHQ2teYQhrBS6TQjbfqBRm39l+OrYKdJHKkIvwYoLSz6+qgiq
pFLwHV//1oQ2TITAD3fqDGpiC4Ux8jZ8/jLF2FaPTYsWSe/4kXfrFahfanGKfPURire1Pl3AiaDX
7LDhwhhAfsP6P0e1aNuiH58H4eZid1v/M2oI+AB19LZqcGSngPP05PJVAWla7lg0UMmXhFjx2Asy
UHq8HjsjwlUu0nGY2QNQVRJkD2gnTeQYpbZmTjt34k2XAwckZuU90mkHpTLQ1yFX9QI5O+aO2iUm
l9gSHj3urUv6SJJ2xjHlCZJLUq1PYDL3mVG7S5/TeveT2AX7Y77W32PCuOHi4hzc1U52dYAi7udN
dl+u47mzmDwBf7iU7wwj7yUi4tajqpCQlhnL5b58y0Eo2feE9ko6BGbS4dKjLU6pOeof53AyG6cL
yYatajvkFX4CTuuAXHh5d4YliVqTildUtrDcnBzNj7R9nIoirM377CgH32q4EcaKUSMEY22kKDHY
ST3fsz+TJpQ2anvZsNwcdm4sMB0UQwzml0jV1qioFbExHf8TF00J74uROU6Q5ZIA6RctYFUrLzdK
6RZOdqSMyJyjh8oUC2Ly0RDHtr7d1nH+bH8h28NLXj46d7Moly4KPS9bXX/MkclK3XE2Mt955zqj
7vLWeTgHaopdBG8DsislsLVbJjbtHEaTHF/4BPuHyexwRqJxg7ixkrd6ISYi2cZXPMkUzRQMPm7C
EP2XWPrVxzKP+JEqkHUqPlP70b1ryHVvhFGRPs+fHE3VqAplMKhLfkj7H7dksJJDAKpNxr3oknE5
kbHGFQSvQeUYQXXGh1SBlKoCOl/AaizZw9mQZAQd/NOn5tp0N4DcGwJAUgF4Rk3t/94QlyasFpQe
4SQySqdX76oaHZ1r5yb+hVrnY31SpAu1HdVgPdajfXDpXwlwmh0U0K6W2cSGNlpum0NpIKkPEFO1
QKog1mv7BGSpIMkxE5t1BfIaRZpi8ZgnVbTSI22PHLQRjbsDfpLXX5FoK8SS+S8MRRjZ6AGXMwdi
OxuA2Umy3xntNt/LZ29n1bMo+xuMQqiTKU8rdj5X+3mjqLKu2WLWBXdRp23cd1lHEDUfPiKcqsit
zstI6WKa+L5d8KhyNHTUOnD6igaF6kThElAn8uwwAlDs8YHXVZqZgquL8ly+Q2wxEmEVva8SAh0z
msYehjsDI+knN8nHeHedPNbnUWW0rM3bsYi/aVKtQP7XF5YS85YWUehsoOi0kh3ei6QdU5Wk67cw
OVmL6CU4oPfWmnHGojtPE4DiwjNktdhJNUCt43DbYn3vaTP0erH+pS09pWiB6EH2gkrY56GAH7QD
L7pj7jzQ0FinESEaahgyyCeAoIDPqVCVo27XOtpJx+VnTSfoxo84kfD1xZnu14aDfpFWzu3jqWzv
+T0WRiNHp6PfD11KFeUjr5Oou8jLI9egE0bdKSl8dqCvuS0O4no1uefvpMc0MkHVxgJAQ1Jafjmn
QKrl3EYYH3jJi2MEeMNB+Wuks+ZCFiQNWGUG5LCDYl8Db0yN/JK0Teo41is3h/xWP65lY1oXy0bn
3IK3i2Ud2VpZfybRvZCbnYow2Yb3lm/N4/D3dZJ3Ln/u1qlu9OXOFkZ79PabprIHira2aY7HDSH4
oRgMxCfyd81NUWoTTI7cUEyfzvmexKEn9i23kTRwyIBsFLt6BwM4D3wwFyNqM584UfjNqjLvPo21
8hLdubZIuCTW3gzZQe/8SFoZpJDAZ49msQ+2XtiCX8FU1rJXaEcEOFP9spVWW+JEE7llF7EIk9if
iy69PenXIkBTYo1refj8ZfxPpNrOh27NTkTjQwPcPTMahP03G3lBs18bjeuE0aTsF+2GvdiZzSnE
QamYLFzEr6IzcSwKRecxpUfjExk0ojZ3KnKNQmpa+SAr9BmrZvpJwI6vtTIONvEdaBFQilzB6mW3
tq3Dei7YeZlgZ2HMaRgOwvwBecZ6NPajSTHz249NpKffUQsRa/gp/nbU3MN5VOMNmsADMofdSgG+
LHxsHoEBZuHj1gFKs9UVNaWWhUcucaErATLGe9NIJb4igsEL91MTLxXJ+2ujTUrKDfoZAhZSMnYb
FPGQA+1Bn5kPkcyyrjdBWk2RewkOI+4tkfLCxFdnH0iDL27pNULNZ/5+92J9J/2WbgXigsJ+nyj7
UxR4y16lsVYXqFSx6fVhR4m7otqKENiOQwVT8b5yxRJ+KCyE2a8HKtiGQ1c2dCLkHv1WjRGUshyJ
deJiftHpLCv1JhuntCCaKRyMSz4EpRr7VkA3QfH05JN4IX/QWKEOl7eGQTbI16EXOa7jQiaa+KBU
+yUpxIo6wuYEKtryOjBv1Ub3707+7/FoVxXJS6X8tr/A01IvJzXs8/EcZdymjjGOqAXDpiiFTAfT
0OTRp2RGQWJvieHO+BO3aSx+jGP4YUnzTiK8BpmkjrOF3nVURZtl0kHEWYdRq4hf8dinCUCqBqmS
F008MFf3guNYEVBwf77h32j2STMxV19RXIlsCk3asAvtw3u1ZC+K0N35vuDGqLSe+Catrqb9dB/k
YRB66WriqcQZz0O1A6UuWdjcRV7DQompnEnD3WzXveOQ1lkUMv1in8KLtNJuq102e6Ji/ewzUY3d
3kP+2H8nexQfUjZJ6pnKxL6iwyl8/udnTlUvza2LQyxEvKeW6bh7ayJqI627BsWvqlbFptRU6qEo
ogflSv2OCvwp5ycb4cb1rwDCCi0dsNxvJzVfiwjem6eD/wXH+WPazZhdrqLgqWGOWrDdCnyapIAd
+tjpimE8tD85VrfpNBFH8RM1U9roF7/Me21G0FE0S50qVuCWMXIURBgM7QJnoEQigK8rOFy8UtQi
ONlajaoFFRWKeGf2HQtL6zdgtrH/mt/kChuM+RWY/yo/tkXxiz8cy8TX2uIWk9/SeCAsqDOxVZ6O
yVF01zLuETkgbEqcUEU594ps/4nR/O1O6KfAq15cicc5iHbNG6XcyCiT//spbwq94+aLLWUt0Pg2
ON/Yp7N4ArHdFhPQYr3Xrsz7HJ+Ox5kop3otOtt1lR2QEkGVT5Pf45ch43OWMHEVRGLerwGB8Q2x
jrMqGx1yERw++kc/oIf429XbwzX3DBSaoPsXXAAk/LGBZ+C2O7mVy2B0DKI4w2KOv1F94wHWgz10
Lv4Hyj6ElAv59gO/lofzrqAgo2CVygFN/0NCEOVgLM0bwHHi17TWgF0XhetL8lGmTeo2GAFC266z
bPfZ3JVWdFKPO/9Jdq+lvMu58eBM4app6jKsHXfMdH59N1TjReodo2lHCZFlf+EyM7SzHRyUweEI
RE1d40XaNSMuM98a19g963t5Me0mCvt0M/uZ5zcj5nG+7o8cP7B+bdSbFbj1fiFO8MkLsDSApXP3
+H8Gsdr3jlXlXiUpCwcKTR6nSolEiAP4o+CzuW9q9NSzrgsSKVnRKpseAsDkWjXTJadgMBJVKNLG
gGcPOMqs63+ou0heQge1A5w9caP9buqtBCeN7Nnhv31wNuM2PZWlrnkDCcoP4F80SmxNqwD5No6o
AhqhxbxqYP1mI1nHDtFOEDwJmamjLMZuh8pi7Re7CFt8FWs1PtScW6wDGpVkX1JKccil8F+MBiFH
SwkXAsh3wv9Pex8nTw64bq4kN9VBKPfPZODaDI36d2EEgDE4bqFx4wvO+k4j0vutkQBUAFU9MlQe
iju7E5eodCCxhrTXUbxyQ57oUnS7RPSKj0VA62KWnLHPQeWEeYD4fPi83gSfNWvLBdR7eWZ1IAOn
wORH1D0d1fUbnqlCtF0bWPYYxS74mkmqg68elcdUeguGUW8Cc4lhdm/0LSWLFQ9HaeEg+lZLuTMO
nlGpoqkKMAeeSfNEwegbWyfEYvQDKhe1vEFxfBdYeipjnMxXrcozZ5bbFXMYbCqn2WcgErxyoeRU
JMaJUfYFUKt+IJig0btI4F+1354VmPONixUWD8ZASZwr7Qo6iwln/kE9+7LVeDeZMsPl7q8RDa/5
udDrKXfYIuHIwn3cye7IcVneJh2P9HvohPsRQkpNI/eYXDAAwjIY5Z4r7nJLdpoRsvk4RakZx6S6
wTcKawpszW3DrfU1kXTL5fSaz0PTYr0sHd7XFpVeoSEp/071UQsApm0TsoBAJln/7d+RGIjWosbe
OdOEv1ijhJBVbJo45Y3lTqAokfDfB5L0lx+Dut8tYoWGchJ0glz+w2/xBPIAsHZzXqS9lyla64am
SBZmkILJKNAkn3VV1JXt9xDceRKWGyYY52nRFoi615LwDR5IAFS5mFGKMHlzcl/RlLo7Gg5I0GJ/
Uo7uUSDzCZKcek3OJ6+ZN4rqevbRnulhf/l/eqfEA7TaORUcoH4b90tgI0XSAL0/8wHEqaaC6xkw
VSSWTRrF9KqzpRW9GRRVf9ZXmfYUnF+dSund0aM0mncVghQW66HnkgOLJSDg4tfWS19f6qE0kSIh
B/H7b469/swNDDJ8LbxyyEzXy5ME0B70pgE/D1oVxqoOUlzfcVMImKPOCNIricacyfOijPooz4km
pJxFzGXr6h2bOuj4LMKSHIeALUw+iDt+dJuPJUuWFjek374vgVjiunb7XLvx4NMl58wt7ZyjT0fB
0MQNE3OzfU9+gYn6dVrfoQTvtlWzeOhIOgq8GxnU49dGZyYqX8NTAH+Guj5buEh+qgo9/dkRUPww
daHaec/bm+UK2e3djb59QW6TwQo8p87Lcp8oyS5g9maLnbojsbuT2w1yzleJ82kZWMRRTD87lMka
Y8lckg041iIqV2QPB6LvczNAYA2GVtpElrZojrQoCBE2UrnugbRz3AH0OZvFRFptkXkRWPgTQwm6
faGgOwnZYRN4UwGYP94DqRNCkyy0dDW/YbhtNiD8PUOkc3YIXs9EXUqMT1b6V9yBzWTvri3wDW+/
BB8qPpD+p7CYYNHGx02lUoM9HAZ2yhzLG2/47EKMZbDAnnOxGh9SfcKwH1obgbXO1H/SCYP6ax0S
N93tCwMH5Cf6hDNhQ5wYhG2z+gm05dBKjHYqBKUHh79WABS63qdRTU9bmRROWbnnXOjk1O3SzT5R
3314fkEvghIZ+9Z/1Usx78cXp+QLddiJYSHnf5GfrqvjTsGaMLCeCQwjEWghxvcFXkD8Fyb+V4V3
BPbVZ1I7Kjmi3BIomFYm95dSoLTeeS1piKjQ3S756UV8tIrSctqa7Xbhns04A6TcdQvxc0PYiFrV
W5p/MejI3G5v+EjLo5IrFQhQfY6+4KRfXpWgqBLxj8ZAMh+gMJfwizA5nJNbPij23ZtYgj3n88GT
Eu+181qrzaKjePZK0WQHEPY593XPKPS6XlM111QYQ0hUxsCAbMkbD9BMOTRqyOo8dfDhNXHdafOJ
qjPano+n9fUdqXLZMj6lsyv2bB9NBjwPjI4FzPTPh0EynLZe/g/bSLVDt1FQtLVdX5YAfQSf1HpH
oJQ3qw1irp5lZW+tCtcz0kZM8m4hNs60qihGzyZV6L6l5yQcxaFC70nuWRZvFzkDjybSw7LXD2tX
Z1SRdxqJ8P3ZUrYL7WdcUPUaNvAIYq5GgLD/yerE9aELxYb7/k/ZjJHCo+PgjW/E2u7R54WYDj0p
BGnl6GtqzAO+zVVtjNVxR0rV5PYcIkNcK9CzJPVsxXniufOgLaw40OpV5rAlHoFZD+gNS3S01emY
xWXZyks0Bsn5fCgJ/xGTLEFQcb4BbOLWIKTMyBnyASeVdyerVU7ucJTiVx/JuXwcD+wcGswQmWE0
uEDK/A3rrhogtB1wJmpt/q6sGkGqtAJjV93mxGsj5QdBxhJmB4wmMkAJrJUuliim9r1Uci2mcxqn
ZFoG8dG+5zab2b9oxX97pTQxbTRhOaOP0AuolqWrO4mvChvc3YTeAn5cIDpn0A3bUz+7uw9As2R7
2Nc74zwhrvMxnvjNI9lk0ISCJ67a0EIaselsA71TIi83A9B6jV8A4/VauJqE/JYMsY2IGaRtkPwu
WI68EJbA4GMtiYoCkWDjTg+Vbnf0t7aCxvznWr16GNQU3k8ATeid/5BAxmS+9p7aLi7lcAmKDhNq
qRB2lnl9N+l9A6gafRobjHAaFm2BuHlCl4eoUK3ntVfaI8Z/WeNAx26aH2HDzuFP3Gt/T7g+kLax
tYf1kq8NaR3ALPVh58CNNGPhGvjxYtJVD2cak1ENmZbfzHQtDeaEn+17HOIJtVrkDWmXROwaa8Gi
yg8NTv/CjDzqJ9mDwZZ58QbRO+727cUE7JxDNx5Kng4WatbvoX92Nddv5wb68DQ8FABhxnzd4Yls
Qv8dVuoWhAVlo0heb3GOlW9nLOalXGNBzLNO0i8R8FXz0R5DEThzvroj+KkwdcaVaVQ/3BXeSX+I
n3gO/5ILtUZgZAAvYKcnxMpRJ6m9bMfyzwQYfkm5Cs6Q6ywm8lDYK5+SHqP1D5OG5wp7y0vOxigX
tcy/HcnBEo0l63ji59JhQ/Jjoyy5CcR7VEcT6bhua2JaCbqrmhBr7N/VAzxjfq0bnZ39In32qJh5
YFZBsvAekuMGGmgTqISG4lkZTiTwwy5/m64Xlqw+On9czYLLDwUzBf8y0FOqu1E8IUMyT5L8eo4o
ZCcReFoZCqB7iY1YvyF373A/oQ3iaQOqisX3DfNZlIArHJH2+WiZNnAUpL/cl4Ps8o+XoKIjnTN5
365MHCuxaaOzfbenQ2tOQ7WvybZGoBVzCSibJSUUnDOn2+fjfJTVcMlufqAVOel1D9er9S4h37wr
myo37OBjURIJCDrfhl6Q8sArj4atttFwYRSXQlK0jxsVOzzJuWAENLgr3RpOJvPEWJxwiUmv8L96
VYgh3DNm0s8LZo9/QoOQfrFVe2/E36r9aQHrqsQncFsApT3eK7nUkcqExEEAIiMRMKBuWpUkbzow
oymP1xRcYcxazuJoQB1XxXJPlet+EV+u6WCpmXVqSgIXuAi2ToA3oPOlR4dwn0p10hyE4IEiDRtw
s6aRgM2ZO3TZm8jbvLyRIghBvlPkBYAKTZQeHQfQDD44V+Tc4AiTGB/Y6wqRoLSUIqycVILgUxwp
9ZmhQQmCyEzHHCxDcFK+UQEB38+cN32xeI7uNZQX+W9z76jkBvQ9jh9Coc1yGUjubtgj+HMZZmTA
51rtMyRHx8rXYI9tyY0bX99YbFyyzvw/aq+ZkN+csLuMRP6JKp5EwMNzrlI2vkGPQYb6xNm25+4k
M+Ms7sBbdImBb2mM4rJBaJp07728Cdd1vGbKFBnWcu7yfdsQymNPxm82Yq5D7dScm5NL+QDXYx/w
HDa/pslomuanms1JSFv1eJsLV6gzmTbLph2ZcRqhoHPoqVSG6Uv+ieTof7ARVmBgB3iW8MJzIyOM
VLMxxevyfMGedqa1Z0cFhbRqMbz5QsglKxX3lLlhinUMmgNP1M0l3rMAL68jpXVQn8SFJWHSrp9R
8TtYLeoCaDxuhh8UaDrDgNM2zhGveEIlOCHaPpW8dB7EECXhwwZn4Fvy8QpKw3FMxj7BaMkfnYZy
38qYow8CX6tLQ/zMlb5bVsyztLWbSeu8hyM2BP0Qf4HbeaeqFi37CmK6AHpxBmPbj16NUYyK9iDn
vsxbWqMiQNIfVllot0HZZB+8Ep4i5UZiKBR8cGWqif81Vxgf3KJhzS26PedUYElG43mQgwCZmV9g
FDI0VP/cUDkWTEe4x+hbNO3OfAbH2w2u+WojOE+VlukYHYUfszKscSBgIFfH8TrnqnDc9gmXnNQM
vJVqZB+2Tk+t/CgO6+LOae3WwQNf9iRWzg4gt6RpE+MQEdO/lQxdudf+FA2dVGXxSwMx5vW6ekv2
QlQVCTv5mcrP9VyjCi9K0BdbdD3nx//WygeU/CDenx6wHWNB/dtWbfXpHJbrrY+E3CTdaQooS5+g
DAl97SKxYBCaoXbJrgB77LN5Gk+Qlv7AyK4YVsJJh4xvcdZCAKFViiziVYQyAEnUr8iOqRoxpY1/
YM9yuKN+o6Es3S+WT6E2r1KZCtMR/iDHal0OX98Fn7QYhFsKVsWLyYPxjYHFqwZBCTM6U/N7RChX
Ojel9iSeQIvHwEufdceRFpxOY7AHTksMYQgm8jL9V9mwdSeTJHw46RUC1EKH8v6GUlqXxT7IQGfs
ZiQhmIn6C5RLyFcsAtU72hj9ZUer4Lq4U2Qtb6751nHrVldhjIeHSmJlzLjRh4l6OI6LUZRLc4Gm
pwvOFNT6pRBKfMe+DTPUhw+tgr2f0kf0z9gkCPFUGZGhFMVVhEdWT7t26QDu9iCGZMtvC/G33M3W
rKQRVlR3UEd8SyeLKl0MZ+EEVcZFOP4h9QAhiowUdslmAjE6eS1pBZD0T55TrvPYa0KCLP/SQn2A
ygd2olP08xX51g5df0LmNow9aclRCcZ9J5xrmkxdDby2MCSc70BHT4vyfScdDTVXAmPZFWiKZe7w
hRbrNZKW+1bL/7GzECQlSSUud6oQszdhHwla2BDqdcyFuo4K+Y6p+jVMHTp7g1jHQhNFoYz+IYOk
CTL7mOXatTS/lltEhhhWq3Cs6nlAkQ60Gn70audE6jy+9bmXgYeH7GmPy05iOX0aiyhD2tNFWw23
yDGlfGzii5YhrKcmfD8Oj5c4VMKrBBFBK9EDnVkJU4AC7LySmnYHhIejLT0IN9uZUhW4+lxg0v5S
PHY+msxeCa451LcBNXEpEPj4nb0Vwr9iS8702VxVd2UxPpL9mY3OUsjLYIV87wpFmxjePOChX97/
cSKDOMrtkJVrsGP9czw+4v81kcCCFyvPOisF+M6e+sOiRFIBq7DH+BQ8MDehNXTfG9kVqt+vj7o2
E5ibLO83wYyuYogx0aBNb5aPARo9UrNY6MDexKpC+UtuYPMURxKxQwQjgpr0Ps2I0h51KKcdiIeW
583VdWqfVs43We/HZBiEk6ukM69IsN21Kpz1GihdVLjgn5ibPponlW9C9lHHV/W6aYwXi6vtrzn2
KI8vXGOK12cwQJxFGGFdZYpqr14uZhxOBrOCgNUzq7AbLDFJ/DjgH2M80pFUa74BL/8NBN+Ms+FG
w2INz7UllWq4oLbIDlIjEShuRpRuH0g2JiNj4wnfdPrcGHtXsUFweck71K2HbW1wl46/eeH3RJO2
8xdUMAhhPGenUpWwTnLsx+8hMu/oqhqKvxY/SVsxxHp2uQvizDPOSRTDduFTJaPNeNpgbf72Cjn9
ZJHVg+E1NJahhEpNdLqworXqxMrOUExvkVcgr1/DIJSNTWHoUhKEWGsiKubBBYQORbcAPGMKn7BB
ZWx9jaDbZ//5qUVhoUQdvOpxGCekJ1etoSFZPNPvaKa9xYAG3Wq6z8dJouFinFZLds19ayXZEEkc
bX7aEtNWwZLgHBqCYyG0vpGVMVXQwTSZ1rEkgbdllD2q1g+1a/wn9k/H4mVR5x6Nwl4435tYHpII
/Xl/plbmeoyS9yJJyM/1TPgzIK7FWNmhSHsBmayF0FhNHEb2/cVDtrIXTa+7CzJPraRaN6+zuai0
hUiO8nWxvQ1tv1m/mGbSfBg6ZKS7bbEtX1z9AyQzPXWhn8YFXHsMi1Z55n/KgJMienO/ITquIPZG
qEcrWZ2Xxl6qEmOqgAKBCQCXY+gSeCItFjH/yNurYZLMs2vK3CSGmqNog17Nvjv+BCjn2Op2Xleh
PShcQ70w95j0NuOxJGNehuZju52wt23n2NZy4+eRqutN0vlLoFyb8SQHwevpDDZYTUs6M/E8tLrz
WlYk/ElDwLdEFPkYshqTXHCddUiq0uvQnnLTu+BLfiNSwo8q3k11vD7ANiRQFRefi7w3nS9PqwR2
dGvHRCXVzSF7EIv6y1aRoBzdmwwDpmhQk4f1J4DhT/ilmuKTVPKz78asbbxl7U79gc3pk7dM/wmU
WnMT76ryLr6hxsvI6PufdVtPNI4hex8Pl2JompzFURFRW7ohQW8uOGCsKCyXP7iArwSRhl2xc5MI
AJJAQ+7imTNJANasnPD4dh+PWmxcSJqhUN5ukdYCDM9e4IwGnGxL3yA98c7OPzSmgM3cvpfuAZHk
8DXZbjoYnVoUuNVho1V/2FWzyvO2YHGrNmqPcMNhlUP36drWT+uwJuMrfezGmEZ8RVF9EitUvLtD
T2gry25mMbzJSA106uNJt3896s8/ba8IhlGItrqoZH3Id1nu9DA+vy2mrpodIuocMrRqaDVEaEM9
ZrvnJBZdLFBihWGU0+5XW4aU7+JCxEw41S7pR23GeduGxUYVXYrpxGjm4S5R2vzzBm5G+8QP4dz0
yAvHrMWitG5FioscY4ND15y1WWH+1DrS1SmUf7nDEXkJTffCthdXv+eWmyI58KDtDCKJRmM3Fe/j
n0VpFvKkdmZtYQduoFO8Q3Sr3lOIaGXbYPZM9w5itbX3F5DJw6IPNBDkQU6Iyze6UC6OtUysWFCf
LBGGrCwmniKA5qeiPXm1b8lLWJX96q5s2ie9iQO56rdelmpFb8nq5ZP7KUtN+xUKZVbTMA+mZmNg
lKkVvwTNNSIbt/wnERpqw6kVkHxQjQZrWNlPNUQwii0E1YwK7agJBIRiA2BsrwfyLfZTqRxqZvoU
9ZtFWg7hBd6L3OoS8U/SZoii3JOgbRxa4KPTfnemDLE0kNs64tJ/mmYrjeggJdSMDDMv3pCxTukX
0uJ6SVe+maRJD0SmRxoMj66khEyHvZykgDU1NpdA8AVnE1JJX10ju9l9Z90EytLxguGDaB3e1GHj
lKplzDkrPWddksfgzjDhFFa9SeMXfZfO42R9IJtlLYZNB9PxX21VKKPYSqYnOaSdOC6SjgJmHDiJ
51SD4b/pK2Kfr+XEF9cVD0tLW0dnv0MLZO9xtAvBEmy6BTyeSTq8FML6qORq0SOZuU6+72l61iXX
cDOVRZVQYy97yOXNX7cKM+7WIIJ1HN6p7/l+i2B2nyQc5u/n63nCl2UoQU/R2c/168kDoRi6G1BV
DtQv3j5rFqLENiI7dG01XAaC04HPrr+VYmAL9cyOFOV1e52Jdgh99HpCsk6/nYvuuQPGrNvAAEq6
kNtBlHAkeU0zlHQ5Ul7RONbqqfxAG86z4WiHYqe0q7dw4CNPJc+8qTC9MjcmQnZyNXoi7tDbJQa9
NJNDIWMA1qFvm4RBKIaIQwWbsRpiDM8wY0h86BJwyK21g/nxZFsKrL3pys23sPgwfZmHUVPuQcZV
AMzuFrmiaeAJCn0UEZdyu6ZKHvfyJPrXZWiJcYmeJNRD19tuAaM2qnExZcgu4sbwLjP/4F/UUuur
J3L4tqxQPDkMdwRjGSWzZasdR7bPjk1h2Vby+ujGFUSAO6W8xOS+EednDkV46b4cpnkQcsd5P0DU
c/zpPyqrTJsoLJ7wuisNv9Go5S6AexPGuuZNSMYxvHmjZSoBR+aZjJMP1E4oqo6bcQYVS/RDgKKw
SauOtsjeXVlfIyOqJJldnkD5JMDOQzC8MXjzM2okfSkbfJ0qqhZaEGDfHv+I5IC620TOonElYh0U
UIgCOPaPgrAvauXbv1FWP5rbzDrovFpbEkH4c4WmzLyFYDJyTKdByp4gDFAbfCja4E043j5Q/ndQ
UM2p8ey6lUnsFJMeYBtB56Xo5us7QweXkwC0dG3TST2zfilxl7/uGBLc0xsCwM5ek6HM37aTob5M
+lshHY33KknmBFfILbnIhwDB5b5IVnf6Xt9tH4boAh70QEqC4Dnq657vgGVTVnBg/Gs6YC8lriGe
KBJ8YqmWjnvSckjgN2F1meYOcTlL1ljO/+UaTBuILMx5FP6MKRdjRH5ssznzvY9k2HyoVVRo3gQk
47slqVc3LoO0Iy3y39J/a043EfCzA+/pmv3a64zr2ZhURserOOYf6cYTBUHOwKY40AGYlBUpG7cj
/dgmQb2r7iPO2M6dtgfaUXP3+P4SqyqMBag95hppNRBVm9B95Pa/UgveepOPH/iHjRRbU6/7Kzpg
q1fqQIRJ809UbOl7tN0+tGXEysHE6Cgbqmw4QLswKtg6WyO7w07+Mut466utQXxZl/AeyXCr90VD
YrqWo2iBih9QjTDPbDqlSwjdcC+Hd5JUUFR00UmKa2VBb5a0K+G9snSYrXmVMI0qOaIKf+kE/IeH
rBp095k70i32p130146JVoHZmr8b1kTaae//0rUPQej7wdxbVNszHjVKzdeahTdr/mHgnaKHh1fO
RxUPEG09Kid/swD/9VTatTGnsCPxyAytm2tEmNMLa8xFKSCfJ7XExWO2DW1f1ugD3ST12qPkUpUn
lPPyPo5kzu4vxmRfzOAUWkEfpVS3DlguD5EWil880HMAgH3fBTY3Ow5MGtQU+YPSu1W8lGEi7c2z
sQKDX8KRi4aIgCqdzyF4jMlmp8jcRfpxmjed/AWorVuqp/R3Ih03vqd8/ts9DXvTgm3J4k+2UO7p
/C2uhuBfWwravLLaFdk5PQJTkkGNnaZrA6rrli33yveI1uBtSh8wWPUxdFy+URl83eRPFBzUl/Jl
A4gb1z6CDILLIZVKC7Jz2QgkSPxuqJSodqH830eRX+2UydjtDMGmqirPmATYdMiGOVkK1+7c7IIj
SwVeDgCX3f6cxW94HIIU5xTGAs2KCWzIbDZxGkfE8334f3o3tIZGIAXm+4jXpdY9l7HD0M/PZ0vM
c78U3yOmLKkEi3ZAwxwk19jgvXIHUDNPzu+/50KIuNxxrWCza7xnsmY9IcmDwGw48xLorMmNTq7P
D8UQqpynh/a53R5Vn3ZF/cxrYbjCZwTvawKNz8xBRXZncxgCnn2hYaocodTLjqcTpgJcDhCn0PkA
Qj4Njk9NirTJf/Iu5oOzXXsE0HcKBfZYhDvMJlJOFtoX7RXH54DQwf8BIv4wwixwZVNMPuAgSmJ0
JKPbSZDNosGv+R3s6ch7FFUbTsqXJp1rLI+9z1MD0MhDQrYf3afF9oi8lp3o45CduFzy/o/Cs/6i
Llt8I7oNFN8a4XEV5YFlLlQKeL4MxP5cGg5QHzLfaDg0w+/yRcextdUk4t4WHfUm97QUJganyyeH
Ny43Ttoos38u0Ykcj8lTUCcKDgkSOQM0oobdlqA5izof8wgKdrJPKIuoHaKtRKkSnnUQc3gdC556
qZZvfhsGKm+dTgPGnZvulSBpyK2JwUe3EUrGJDPXbrJxkB3itk9jURCkcdsqC4Bc2S1BmnZfGKhG
qJO5KNTsTVEoQAdjeNP3YN08RT3zoBMj+LPmf/Tj8jDYMuWEWiPlLyd0BqD7NKgVDr8lDtuuJriC
66bMv3I8ecHlGVmYtbRcPVjOV+R91aVR3DWuEbvJ23h/GmAuvz9j19CTScie/j1H+EjY3Mpimhv0
BMNAWmv80r70iOexmDph/ugiDq+yp1woqJ8vROhpZzuz6MQe5uZ5KkOdOyeprPLcNhq7tTKPFRTZ
yNWXu85izh3naAU6oaXKPUxLA01kzBmyFZgNkwTFVQPKzTOYbtyNeEcmk1gzgD6+jRW2w15NexJ/
ch4B6GHTv9mpm8rAKtDzd1cBWZae/2kTzNVGJj0pTf/QDaOIpq9vAA4nSflTYEl8pPYk76GS9tKz
tMj0QiRHp9NvHVAFynPHW3Nz0TcudaeMY0eB/4ftUR1MrTdAuZU+DGqpnbDgoj8spMhFivkXGrcb
nzj6oBIVYiK6kIysyoMabG3ALPleaVapleY9IHTbEpgTAOAbsg0H9lxLZ5r9fcuCT8zwu/vaJ+Bf
Y2prOK//m7D4Gde+4I6XbCpqb9amLTrz0v73SUxE/eJGmD9wGUEaB0jH83HgbaPu9Qsp36qUDx3P
s8uYpCoDY/lMDCTwQEZBFj/KCFB3C84Dp7ny8CRAjakDV9OuJOxNvhxbWZaKSjvX0nXBIoyi9h1y
yux/TGFu67yk51q7YzpX3y5kCsZQsIcR78tQXlU2eHOBvCoiPmlngByKrthEkR3OuA0JvopzWfld
kZQw1uVWui91n5P4tp2azMHemDQz+bbO2arNt4i+YvsObvkTnEXTpxKGSdBLJxVOeXYi2xy67XMF
MtSNynYG2ikNCHAkar1pnk7mNU2qD52Hz8RBizz7a7sOS2HLjqWLnr2DDTufxpXvNd29oSD1APas
5Y49DzwDOu5yEmpitNk2+v3xY+RL6XvkaHNWhCtMgsJ9Hct3ay7nh/WCpFyJtTe48WdI79LzHCjv
bFF4Sfd7WwE4je/DRNTa7A+wlAHiqd6JmAc7ALSWUQDyJI8liIEzkke/ctmlkvlTdBhVz2SUcTO1
9tkOIpGc+D77cdrCMQRFLl1ZRArRcZc0JxECOV59tL/fr2LlTFafFpcBlGxbd2Er0dZqKDY8NA/S
5XcL81e8nzcp/DcJNP7+zoDpg/duwYUOi6RuGGD+V18EubXOY2x2QHLvjL/aAXKsnoM/jG+KJF+d
odaZ1eI9b4saBylSx2f7c/sFrzZ/ubxmf9J8kSfKfMjde9UVDt5HlOrk4ZfhYp1M8u48/E17XwYw
yXVFA4uabmk/JNmqRSPDo+S1VqjBea4kHK27I4HizgUH8RU+HXuIBv8/1U36znhZK9MaprZeUv1B
X7y1LiZGhO/IjUTUXoS2wZ71qDTE/psjJ0AZcsUFI6v8N+ZLGo1GV6PtOYo+TUEbnSq48DuZ54cI
OLet8qDyWXZkUPeIcy9jbdP1TTgmlyoUU7HNhQ09nuCWpxbThMfBVn/r5bEWBGRJi0kQPunry2Px
Wyg0JJjr/5fofAulXSkdgbL+YGnP/cOZHftSZNVn77l5q7W97C5oo59nb9UNWEdh1pVp87WXm396
C621lwdm5P6KEBxlvCcTNQ0iPBueJcuDJWdDV7bHb7p3kEJcydBuchUsjye/E0Gc/SSrLVe3MCp7
T+hmdPH9cbPYQcyJyobGX8Lucv1+flTXu8Np+wtbp7kV5p5/c3Av2Pbl96pCUom7iYjD6Y9wloE5
sU+TTakZNNnJScD2+dh4k9cTnx+8FJGoNrfwrnlyYpjLK89xU1ELJjA/o1qajDllaHJr3p/9qtWP
lY2l0OikcHxCTI+mXGcjaKdWFBH34Cn/AqCfnVXQbtE+3PGIf51Kn17BRoaZM7aOl3srhvu8l0dv
8Medmrn8NHllxO9cU+scmUEJ+aGgSeIR+Wf/0wwjgUOa3c8TNxUqD+v5JttHL0sbNnwxz5ZmTMhY
D1McIZ/a/u3gegWq7vzgxDTVPxoVICYCDSCRc6MWFZjIEkmt5CmEmyJcNCWtYhyWG2yeGvqMiWeZ
ORLSRgvAGBtGxxaOCz+1cQY7FMtrX4ZMas47XmwiG410Sb2MLOJ1fYYxOizBh564f6eJ651j7wna
gBZHEejKxwncxJ7VlGDOUdxNl/pUvbEQONo5yk2DUlhFzePMPIleQoORrKGAasQwtqS0M7tIAqf6
stBEt5X9ZcCmQqsMlFv1sY3slK4Vc7hfIVTgViTv2t5juog7/82MwcUT5fudXId9MEnWFGQA6pgr
Tq7Pv4ug1V1mHOEoQYt8qBIqZsOqy2/RQnwpJYbLvX0JrXrM/i7yyFhzhjT4y7zzWx1AQjf23zzX
C8wYuEftLzr6G7tCm55gfV2OkNrUB2eDytfXF4y70qF4QPKMD/oebdSfUzWpSJQrB9MrYlZihAPV
5mYy4fkUSB2zqfyv1yKYTr6glX/canF+SsMid+rIdQXw3nc0JtMUlVAOmaS9aodfZpRxCB5Fw5fl
FKrTUR37vYCg7So3kHcInx25UN+EozdXG4yn+DzLkppLeeJjtO6lhwfnJ+CxtcUV71hJDxFc8wOM
bJmevBpLgeBKeTjsoVFe/FRzy0Pq87sfnjKHdbs2dcIe78XwUKJ02FDt9CRc2z/GvpA5zdqjyNVm
Y4X3tmIZTDdAIGeBeKSTDQ6Ql9lk2cfNUa858qKVpTHW0zNzJWZfE6VhSpO1Bvvc2Pnt7DUwaoOx
m2bOZMrxbHrcRxkbsTGRiIPCNcKSWE6p8eYwxn6pIxTuq90AegCKgGJj2/7oROnm1+7U4b9NVHwq
U6yLecGhc0svKKTkw/QOpgdROoh46sxcZ93wEBZ4F12tP6bVKNHFT9kO5S1wCxG58Zc9JWZ+430u
4iCZk/oiQIsvPbXU56gzXYSue1y8kgSKGQkSseWjTxNlVg36FyJK4J6C3PM8sWHSEYPpuxHxsUpX
9IC11xk5npOjUrZd0rPONa4f11ziWZsxi+iOIGxs1SMsmLeECSc786dhpNHBQ1LbPQA+U1Zmdph3
CMvqtYpNYvLG6ksaTnvJTN+bupRgv8yy8Z+cTUljMDMBUaG4SJ9DFMZV4k7ingLMPdlAD+5CtALo
jd5XUhfNNrcbwPkWlVDfcRZd13fInr7BJvdY1PGmEW93/EyYzF5W0H6qvbHGy6wI/jsOtijdhz8j
xBYhWX2YEO+J95EYLsVdCQEWvBpPRHIvjYRXoUyNNHmlzuPJCJYaXQt/ih9VICexLger8VdjIJmN
+wO7I8OlLnmPMTYamWTWchBSPECYN/AI71tqC5fWCY4TrGydY2/DYzqMexZlH/ZKKQb46k2Pjebj
bpuI1NCNs+HQXfs8Gyjfj7HCZnoHyO6ERFKg8lrq8dvVRA2Z4VIBKy8PqleJ5XeVojoo3CYqdXcz
Z9Q6fg3RZV10qRu9ngg59vtZEsmbXAr9dKSBfwMxJKEDkEyB4zFdbgNUqjSJRP0X781b0/s6RInN
hhUTtLyGpVHcHg/aALUT9E5aaOqtL9S0VIawAKK6T1o0XgHrP/026Y3O+EhPZzO2S1y+hLhr1CEB
VcMqXemzRuUmHrPcM4kRxnONcCt2Goy6wt5VBlPQxW8dIYWHO6jjkhy1o/lSbwF9ga5O6BA/udbg
Bl2BculbheHsh6s1navFA8OSzaVsaY2mN/21DtyvKDSVuAPfEHSeOw9hk/GB8Z+Zd+nt0ySgkRE9
G5hRel/7da4oD33U33mgY1vXVjc9BHMDoz2lFP7ieRMnTAD5kMIneshzQqAPPdeHjh1pzYNHJK3M
Q1FyYwJ40D72fjun6IPag/aKohbkKHgmGzQ8fpUcWxi5RHKZ1uCC9eFDwAoI4IAxLAYl34mPtBje
g1/qBRHr1S5flJa0G3DVvwg5rBHN+oFvAVBJIw0mAuC4vYMSjFmQL0rXONP1f6bEzWf0j9vhD6+f
uumkAhf0dcib4Bk73Z947H4sxABXdg81OdbIvlQ2j9c/eCkcwfju96qBOV6Jq3/eww0bSZnw8Ng8
U68Lrqy9oNkMfDHE7BomQpuIqDDgFQxnUPyXUVhFkgNoYSvn6U8lN62+VbDiokaLg18UAMXMooPu
BSlpocyxuJ84meG/h4dNKocYQg5DCOCEjiozLSk3+/6U8YfKr1RzGOMpbJNOfqfXnRGTwv9t13lM
CIRDVfmAgutICoVJZJwfvfiVf8TJZU9nu5ejq++7hQ9hhJ+aKSqnvqOW4vDaOENYA3u423sDN6ay
rUvg2AiFeECDNPGaxPQPCuYlH+lYUE+HxFVTV+ipiaxKqa/DT+GesdoQU3MciCcSGUti+GD6i1jN
MEFpvM3+KoTzBg57a8kJ391BQpci8zCtKlmr9ikpmKMvYvIRV9PnL0joeY+6m5tGFSwTP8fB8hx5
3eQgY3EeBaCDEldzrfqrVe6bat+KsJiGdqnpFpfUIhZcgD0bAdsD5xgYbXRmEqgZzBzy71zW5Lph
eIvmBMrOVnNZ6DCF/+DNrjP7r0ZLDgQRowqFiLnEzvXfm6qWOs7aGfmnFbyr+VhB39O4SytvkkAQ
5D50LEHMirOGaDwXxs6ebkPg2Q8V0/iv4PGwoJeVHRWSJpLZXIPPgyb3Fl81IrjnvYdhZOTQi4+c
va8sJ7OEsANSujgNspDF9fJ0kcC1L7vfYs0S31gB5K4VYbIzu95UWmcxhf9mTY8bQEDNpQEE2s2+
kav/zPsEYsQtKnyHdNkJpu6P7MPAha+H5aAN5piN1DLpzciv9IADYW50IcFUcbmWQS1bmYdpso1L
OniD7fZ+HJpddqFYp0yGqqxoBUa/Yg65GLukvXztgqAzUX6GgotpSGPeRZAxgpj9qetCK2l34+Ey
Jyg15yMzNcNLZUzVVoOJc4xDfNMJ8ydT7b3KO0O2nofmUFZbjQmrQcT5C3xLy/+a3ob5CsxgcW1E
fLnGVCAu1nLkhbgNJF6hf/5yBeuIINwc+x+jfFlKfue45Wahhp9+BjDzdBZBReooxl9VwVm6rq02
vEncRFRFwUIH/VjJg0TS/DGqCP+BneeKeYgLQPu/tnVz3fbF1bwSYuSsXjzMqdY6dHTfN5UCv0K+
tLcJh2bTki3M2c8UYdtxAtMcP041ZBG9p0n2kIAfvtaDOegzi357LwPD8onulsoS0wsw7gkPT6n4
OignMqgHBQupiHDnPcJF1cSZT/ulhjIg/+/xpI9F56Loun1R6f/3d+V4LNJCpsOV89xjVWrkJkxo
RuYIHBHtP/g0gTEhgRnN0IvRMnbXzI4U3kGG7QoTKVk885us9/VBGNotY5/8YH1DRegM4DYTFONF
Egy2/4s1UaSDA2bqqV/KNCyILvTNS4Z0C4gtNZS+4jdzm1K6gXqJqNOgOrbBYKQsh/Gohf2AH8PI
TAPgAE6NaUQGOePsdYRR4cyGxvVm8Y6T7YD5jN5WvJdQzPps7g0FpYBOUnU4/DYdjG4UDFlV8sRO
+WKxKj7bgwCWHx51bEz7r7b60hs0qmn8Yg+MGAY/v2gExveKQgZWEWqN8U9kqLmQUUARf6yQtXVp
IOc5FFI1fwDKjHo0/Z+7Z9znIekhhI4mjTA3HTOHVLzNCPgbSIyNc4vkxwIjMQeUnk8qGbDsz0+Z
EmyUjkZJ/XGuql6UWycacJbGRfYBy6c6xn7NiOZA8REg6yly0jsPRHWDcfxv1ZSRMs+gIx1s61KJ
o1eifJIbTYBJh86yYpz5aqxXpWQwqmQZE1xupgDgZG8jxwGbmzaHEt3BBGhzQt1NeqhXZB5hfm2N
m4+zs432KjYC2dWvvHbsJfWjADfXiucgoT4XyJfltZlakXiysohpyZH8Q0MKBkkF671ctXaVDpT3
aPQ28tC6Uq9rpIbSwbOO4Zne+ydWbGNpCXkhZN6kjlHrU+CcXAD7HLv5ZEO6YROT/BeIINpSjQwY
VIX6RT3WDlwwsvI4J0nyQ3XWn0xYHabakR+XGCdMUON4bufZGxDaamj+5GuxUFI16CqnqXgZrufI
tFHRyhnM9uyH/t8e+uiL6QkjXy1u2LGeOroz8xN5KJRqEW1nirXuXlMMONZVj9yvYMrElJt8e93y
ehsHQibb5jtky4Ai9OCeaasjR8QbQ61KnVfNloLNHB+Vq/hikON+HNMc3z/5LI00pDSVRNSRW7ww
+NG/EsCzAZdm0NT1olRi2RtPTtmSoixcwHWsplUT8JYeiBL7e4sylYh/UCNuKSUEfxWoxKoN41rI
rNnQh7Owb6nI7bBVeiwkBG4uYzY8M9fy3o9c7Kz80dNccO0DVciOKCFyJyLSLms0I5f8zkXb8w3C
ZZEt62kr1UgAtvUisTa6VY3gK0IcHcKAHkwLmTm6UhlBaFidGS+5hh+oBqPzH9vEuUkDeRXjfh42
NIDGg8EeBF6RNYxg6Dsd+JQcI3F/Mlz5Xp78Z0Bl8yBrhM88wCUB42EhqOAhup8Tm4LzsrgUJrq0
gS6DL+NO0bruFoNEYREt8n3Gs/P+64rfceRXidsFLI28UubE1v3ZYaX1wNMn0/MIgyUDRxHxneEe
ajnoyI1vttsKrmxO6YSBKd0Uy4g0zgenv1uPdzESMxm1MXFZOlDf2ZwBtEqbbRc26/YUjnSdpBpv
3DuSi+D9nRAV4fDKo85d0ibwRXsAT+SGt4xQsAAf/JwOF5oH3ySZAOOz4yPcpN3OUOKFw/eYPuRv
9ODcQSsurj9zrL46I1AG/hQvNDkOy4FYHa5FyGPHGSeW5Bq0Mq+QJGe9aLfugFMXaySC3n5FvC6R
c37JlLi5eP9OLJ9KUeHCPzJa3AVgJwBqjX3WULSdt748HOt+9yyQbBZGZVEv1fBV9sb0vEVla1rR
CqujG0JGakJBKdKz4HWlqeRCOqE0ILf8GAY2295bATK/ZL8TOadvTR+tWUPVWOaHPfhaep43Izza
DAPpsX78B+uu37LuOSRZokiu8K/pWLTkJgnHiy1MomZjftI/2s/hlHm7PeDABjIGbUw/odXBsTAm
TF9V+gijby2sVq/VdrFqGvV8hvlf3ne5wWXdvgrgsbc2xdZPiFXUq91AwWSvrwSyTV674ItPw9Xn
RgUzBFNaAytHvaGV4f7jcJPARvRNsP3Ulpw4QmZ3PcVS5rad833ut3DU339bTjDXwlpre7Kqp6bq
gzfyXGkSoJ/pmCHeaLeo2t7+sFxIfybknjEoe/AlMpF6C80e0/NE0yEogg+6Ck0zH1+A+ySS/9lB
ULAsNUgPZU/h7iZ1xuxGGm6oja3xnr5ylLQbvEuYOa/XrX0iiOCoAxXLRrH1lePveW5Tb+XJeC8P
DHBd/tppStj2lo1Wncs0BBDpj8+FQ8u7JDVV5h7bzRb2KjefCXcjIWeycyY++aoKVqgBSio84ZYI
aYqGKK9Zu5i9ocr6cpqMcWkiehJ77vSJ6tAJ/WTQE/IbMCNRTpyX9UY0VLdgExj/aFCTX/YKVZOY
cjTYaMNcRnNjIW0ewVqCcS5mJHP06R5ymdYTheZv0vGJi7okCp7UZnK3PgOSln7Xr681XPc7Y7lo
/wkIJgKwwrmwR18qMk8m3Ex1PGcAa3Au0ACBeJXJySxRraaKfV5pJdkMGl9uD3RrU8HwuSC7rQy8
7/SfWvSUCkplj8V5fgGmrUm1b3XMkmSCs8QL3op3P/3xGocZ7+bvjPEX3yMQH9HE6kOvexVLNAS8
OECxvUts3Iq/acLn89jXbFvvk/K1vYo0YLDv4A4KMQ6XVCm+xO3TcDoD51zWTPRBhRaiE8IaUCH8
4iPSETZ9f38UrXaCqpXelsdLUkjfmn5mULh3a3Wlv3Dj8pQvS7hingPPefI3RJ2skxq7p6ty3gfl
G0pMV7Y9SbToTiPp6H1Mu2794KgG829TkZfCITN2IsJVLztuTBCmahWVvM9LmhILx9/2Jid6ETNO
cuC6/LV07wJE1B5qCIAUTp0sPQOT6WK0ynbPL1qK1Og1wp1it7iKL4o9AJYkidxwqoPVh8beKelo
BAxnejGokwANj0tP6ZoM4WuK68eeG9b+T3ted/OSjPPXXXjRWWktmrgAUM0pn9Gub1YifwMh7T71
XiY7E/MRnAwQxyJykUYmq8SZr/z8+GFZQf3OCaTl/L0iEik7Qht9nrVxoQ4y0f8kcK9niu9BoEi7
BYvkqzj7FpGQvR+ZzKuXucxCa8sK94rMf5HMrJmvrq+/8WZnzu8ZgzguXehE1HCAkI5gJojqvgIZ
X+yoBmfoanTgt9xi79xO+oItFfK9G70BXqEqrflEcN7Rc9VocXMCkF79lbK3pldM/pDHgOA+iYPM
Gyv+5fv2gjo/2ejBW47X5aVoiT0wPe8wVPrWWcdxfd/DyUL9RYIgkL8jGvF5QrCi78B5h1nrSELo
comA8fAqf1LsRVKTQhwJaNAySeeJBjeMkk7g44X9eh5+GjOdEnJd0ELm2spBeq48lf82jH/0oeKT
dTUJHp3Oc9yU4VBnwS9xGaGhDMC3ktZt1HvlQRtqRZjdE7pK9XGsHxMOPAYDBAkM3VmYpx+cZHlI
uNLW0ZfL3H6TCfK++wcicuBrxHbeX3DtXD73FRf7/3CHoJro4FyIy5kZyTAo8tp8ng3T+s0Pbhfs
zBa2VtFXLnBqt8syfUGOqMAhmK+56QpI0yjSCnh4XM0C6xjfAMwide8aw9QytUVjDEK0E0onODlT
Oi/KeYsErrc7bYZzQEjUrotTZk1fxy20dSERm3258EhyjuVctofh94JOKQAZO57vGzHnfIAeZXai
tzPmmHqtDiGEhI2hcFMHZsfeij9w7y5D5C1rOWKIXfv1hnDR67Ovabk/OzDGopaAHkKl9GvtN2xP
XPxXII3zFxTyUb9Oc90fDzBeQ2yZS8YGs/nITn/oQACcKs2C3qEohKfLPy2wG/t6pPtzp+Vpj14z
HMPgwOirclF27PgeyMy52CGHUL6iBHfIXDAfcPnniCzWMHl/nHZeq33rL9pjGYWU8T7fibClc+2U
2TuBlFLKGgeafILrXFqCMuLwaLQcAHEJVmos5/dUNnxQo8vONqoDh44HL926ZAkcKDG10qw6b9ep
ZqL1l4phOvXlgP685wrUdpc7sStw4ehpiFh/XpItHFJJZV9/V6wTs73qOjNMUI4RaDFwYwyup9no
foapHjePUwX+oIVfG+5cy1wurFXTuBDtRSCN5WT95Eu7uVSMuEEDguwtJxCcqAq5dNag7KC/H1Ud
PomHBhpzAiKop3WFxlIvSsasW1RisLPbG2zpIUuAFtNZA/I4az+3ZYW6qVLfRnzozUzUfAuNat8w
8PfLYKOHNhJn9z+4+SK494RFC6NNx3XIzuHa5BU5R91ZMNh7BtN2JBA71xQk91lGFsKjH9sorUCG
lo9yzgXP9+kyWr6OOnA6BVjDxL58g85MM+uoP+p8i/dsn5U1GHxEHBzJei9pppTxbJArGHz+5nlp
dp44MR7K7l6xSuMl7I15EBw3LKRHq0/o2ppqc8gWJimMBnIlkgg3u3TZlY/DaU1cr6n9kttmsxdh
KjWR1ODpRtA9Tt6ErN0ZbjvX/B0tAz1/p5wDiMzB96gLpMh69ZjoH1CA0yUbIqhXH/ppr/iALUiU
EamdM5gEnWjJir0C9VSjDJIn0AOJbr/xn0x1wPHCum5ipsjKckuAOQ8KX96e5US2Dok0KcDTrMYE
6TrgJS93odOQ2qSZzYkg08bEGd2eotuiaPzDS6Y83BRpgwCwORPCF2RHVCvd29EQd6muiT/lBZaC
ga94/TDom8vm1JGYxq1oRNKKWT48qeINpYaLmzLCkLGAUimBa8Cqy07n8iWRgoc+l2r8y/D4ejVw
MoD4J+pdTGyAdWJaIv2xEKGXgSHADSxzZr6kscI7y3wHDUpDDWxWDDC7XrbonCGF/kPDrSsyP8W7
7tR09dACapESSA9XqUsFF6SRxhheBX8lFYcBQRHFIRKoy2+AR8HDfQGDhOAQfhJs+xGjmF/opE93
vylpaBKKRf6Pibw0ZXNi5WD+fOAPDoSamBQnojw9ecs0FgEz5OZrQy4LTasXHWhUSrADft9dYRfg
NsH7ncln7Eyy4lBKhc62FEL9CTqs3xD5IsYv+I7VdF+fNetm/5useksT84DeE1TEDg2TXDlj5JZU
4bX+43NP5WfaPp45DNm+NIaTqy6r1Jn4VnTrtX8yqDkYt5WTSaSqQ6hW0qeDN3wR4LwcXq2O41tf
MikrpGAhNWYakPF3ybmHPKsE8GhK8zJTIr4Ux5rh3qVllFheZXyDh6C57qlpW8/kUEzOckyHz9aP
cV0tuwUwwNas5pJUQv9hsPWflCHFK1LaAT3N7gsAZsqy8jcmNYs5JV3IZ57c28BzdwU61cXJSfzH
ekqV7tZqyurQByg8jQOJa+gGwJ4/HWZia3VDVW762moo3RHcVLpkEgq1VrUFIYNZmJIbWHcXWzVV
gMlpUfiZLBFC5t4QWjkhdOwQvBsljSbwjhOHw8o559VJvU4dcPEcYPeD0M1cuXVKwbigv3xgMVXi
whuLJBOKD2BdLDGyB0RZlCILOTqYuSihftOKSBNfoyJx/RMeyR4I80PH/WO3jL6iEqHM7PYTzkC+
MpjBlbUIPgCm0YyrIrlr5ELGP9SfByVoaleuKIZ2CJOXF43A/gK2QNGPKTB5AdbpVzZ0oiv8ZlL2
5ke8KAJOeVkRrC/y8tsakGKTpnnLs5jinW+ZE7Ju9j20ohm7yFCdE0XCLhuB56mN8hJ2G10of9Hy
8Y9f5Tg4xvNu22BfrSHdowVRXO6655dAvZV+GwvBXQTur+EvlRNj5gJQZWGo8C+Z/XU+aLX/QCGG
X9ULlcPhH7DsfPhSUYDMqyjSzMa2qlrcxb0dDlIFd73Q8csgef5Vobnta6aF7VKrFTCBzMKKjX2n
wzfwJt26CSOHJcpthlnVb6h8UM662hfIJZnCQ7Bz+eYlvK1NDnMZVApdc9IIdz73LxTIa7xQ53Wu
8aOyqqQYZWsDNlf8HBneGAo2lSiAGN8m1oLsz/FELrfMIJ1F3KDwKQB7rYRexuvM60oPR/1vgJjV
cn83jAxrtmEQt4/xAa0a28ErJE56Csp4KKV8jEi4T/MhFdaVW8XHoy+W2XRCV5Pdg79q+doylA22
373RcckpRXCFFGY+77cN2I6BMGZr2C4rKt7OdcXDqrdxcjDSrCSwGSD0jqpaKZU4dOCKyjG0LVgJ
FKocH9I7IYaX1eKqdfaviwnByl51LLHbGNuHF0d4ZZmaDqK3jVAbuGVH9PSCkrb85WuhE1/1y05/
4k/uLd7ikfHLzA0JKv/Nc7kflyiNy+np1JAcZWdXYoyc8FCbGwHCMA5f5QOO5/IE4gkwi7RR2wYv
KdR3y2SfGQLX/uouAej2KaFbCv+ltLxcFLHmMUIJ9Xy6wtOqqSUUKLh/1qnBluPdiGVVD20WewMy
TjvbvQBJ5LjETRp9V0FgI7cqdHgQZt5VX8M3+CWgrxAZcnHlFPzSVnOpFhP6usa1v9Gxv48sPFxt
YkoCziKSuUCUBxCvwp6Kdzo/24Sytnd4GGbGPuMBBnqm1GNQPr2m14NdA7RLMn5iqu+yGkaVjcey
6VdUIm+2XI5S4sPZkcfgA1W3z6Wr5CvA7XAhXXjYSprvBsg/foxtSv9XT6LXmdapEvegpk96cYFS
9DYSqE+q5p83lXPohInvyqh+QsiMSolz/n04VLWKXe41Z7I0r19YTeMSIXUd1rlEk+ftlwSjwqlp
APB0/hlU1zf6gX36ElfQ6a+08Wba9KC4xPhX5ZlXDUTQAlGR9DQzAlEYyna/K9tqO45EuZ37MR40
S75A9vH5Opx7CVt6HQx32/4Kl+VbmvTedFtK46U3iKFJndQTSZ1E3IPmp8GbI4y1hOGuE8fdi8A5
6bodnWPcNHBA9Za1ezZ+aoPPBUVTaNtZpxtAOQ3y6Ey0+emUIpjOWQpEUYNUP219p7mVqVP3TDgv
p2087HfPpRHxZt0Qhd7YAZ7W1mmLgzMu2CZ3GHyBE/Ms9OT9uyWL1INjTd1YH6Y0C2edsNdyqXtZ
EY7AGFFr2sM4xLuO+NJMHMCwq7Vc++ozqu/jsZd76f/rnnhMw10YR4h4E5o0a33bP1wFa0boogqY
MSqbnJCix7P9BEavAKJ2fj54CUKHQ9efxYiw/VzDqake+cNiy2RGj3DW6RzXBBc4aW+2WWuSapXz
yUPLmT7tNp2HFEn17EG1SCwcYyVFM9UgJn9WroDHdLTZU/grtI1M6MvpgwVTXmmSCi5ed2dLl/xD
ure9SjjMp8BYdJEf1Y2CPbiSCTfW9dptBrixpBwMmix5ra+hSznOLMZZhzCl0hHNW95UOD2ZCUke
ocbcG5gKYwUVniDY486prsafBBJeR+OSF4KC1f29VXI2R6/AR1yeFpg1h3sQbj7pfPkqHAMd/Nd7
n22Hev1IxNx1oWCnrTRcEWu4AoV+hfosBy+lEYjp6YGTkRXNIHjYDyID+oBtQHif1stM8OX6mO6Z
gvOVcwUwIyFjx7dvHOeLR5jbP3fFnAcsvduBMu0mces6K4DAEI5C/pKGKIaR6/W836TfpYTx8g8+
G8YszMdsQ2FJ4uIR1zasH4QIohXK0lmQqTci9MJY9301Y0CfTA/LUZVknkowGFw11lpRui4W9QJY
Skky9OX7F3KvM2SJkQqZivmojvmV+7bNseLtNJffTzxhRu/T4wLDLXqTjAZx8UkPj+HijsbR9vDj
mo1m8VY+XIUf+RedPUoDQEFn+PMKs+IbvB/07nsys5N4IScrNH4dgYS2Ay4x5fSsRxnhXGvajuVl
4nHoalItaGubnDb8cK4vfZuXXOMbqtejPOieKJdMZTV04kRQw8lSh2S4XB6DjAxZ+3f9Usa6R+CL
2FqL7X6ddIPeI7T1+h7qowM4VEQoKI29LtV9M4kWW11mQPo0d/K9CzhAuu8emqfUQcM1tF4l2rR/
icHgW2uhPYJjBMxPGTL0Xz78EXlSk3Aio9ws+BDuAbkJQsHV4Veh8dtlM+ZhnXMj1TyIOcIEa2n1
GpiSiXSZE0hyrHLtmJW1wKMDCX2jqdF9jKDDbVbpGeZAgrcH7ttuUS3EkMl1qy+2RjfTD7GV2Kfp
cvZyF9qPbhym9igDh1ITEH8DGhvzND81L81w2sCcTNv7Zm8PNhg7FUUg7OxD6loJ/RGpD/JZMZyX
ZA/qlkfNiccbTikyd5oRAVzyrSzg+XQD8Lf2HHFcs6M7XAfXaXrQZjmxshQQaAbtYYFzCMMJVgMY
wCFTFPQ0vKlJzPzYln+anFjuoFOI6bJ7Gx5JZjLUaqbgKTB+OtApF+DbvrnrgiM7VG9Yvco3bhQE
SZdS3/xaGO6PmXLNC51liD1H2V7q2MVh88W7ETP3L4NxBPX6pTaQRBVvI+xPvqKGLY5nJLxdnQLX
/0g35fNPo5LvyJnjsr4g/o/PtPIUyppbUjcKpvavNdeN+jun52PRYsTbNmPEcZcBe0l4BGHCBO80
0LPBJlG/8WZjYe9jR/vkvAWu92DdpNOcJvMWotF1RiDhd7VywDr4HX+R0BAnGuSm1ewoMtvpqtiV
a1Q+yPdtdw4P9dJbo22DWUgtg0WKdcU+9HPvarTuh7+0MgCH1uJsOsZXF/6KdHcVbsyLIOEXrhC8
cPuR8M3UsYfckG6q+Pumnr0xv3KnmpHa7XhLdyG7Gdroq+f2ZbpUNuusFIikJaOI07TSuOGUAX0y
GzCaF6nPdjGLNC3TthpgBFa6jyFyTaEHZLxgcg1zIkZbSpYUQd48j7BoHtHSQc/jeIUxJgMmPuyY
pLDSntnBs5oJumu9lJUhXqEJt+YQFN+orcKXjMIzFGkMq3LXA+FTp3nHOR1jpuYgn1CKewlXdShP
6A036vcaneqimgJdkEA4HANVTR4/ha9nNrF9pYgoU/GgOlydHBidgmsxAc7xWegzJAPVB7mmo+OV
JeyuQB9LNITBxOCutxgUtXoGwDehy1S+QUxdpxOjt+VIjxrwPlJnYG2aKFlMPnXui6JHTpeK9DHl
Ho0UAj6VVPltm9V+Pyh8qUK7kZuHMhu+5YHQt2g0u6A7oXOnbYA4xReE6UCg1ZWjKBEYURKSiW5Y
rP41OE1cllr6bzd5r1Srj/1QxDs/cYcst+3a8tyMlHLLHb4q1U6cumc21JvhW6QfBNvl2nkd7Qe3
oPHAaP75hcjg6J07Rcs0FmxVtLSiDHX0xIWa08KCGrhmTWxryBitzRMIlb46UIvAtq3AzOp4M0ub
M5zrX0fnQ2cRztGGwGqod7hkaIW+7OTvHTYMwsIgsiy3VHxtksaDt2CXsLqdYhO3WroDOyuDrS6a
PQcETxVVZTLBasrZeywmDios3HmNxSvpvkAAYWnMDDgFCsLF8wfHBAC7HXIpJVhqwRgj9XdVpiRA
BF8c9aL+r5k4SAyJcZnOFEf/zkAwqSEfNzVZ5+iQVUJozuw8u5tzXaNSEi8/PStutOeZjnLs5cl/
XWqP74XCQ+UUWw4sowsoH2hY1ay08TuzP4tTVqwuBxpYftl7mENC/qDoEUdGilEkkd846JRmce8i
o0IISR3hQKjZhvTU5Z3nwG6n92EQyxICHEj7vgKwD70bPybOVYS/+/CHjHq9O/vVTsR5TxN8hhdw
SjJGeChXccgMWSRIZ1k0BZ3BKsy57ftp9IDdTx63jxkoVViHid3c9h4IBiqEqD0GWVyoRd4EYOJT
8nCQIy5ODfsDYipIlxaybBO8xW1V1Uy0eITVWq0oFEHEcwWr0rgFd8XFJ1WURYrTcEvZeOOkfJH8
wi9qgq8VCvYl/ioeaQZxKU2J710E3hp0O1JgvlC1U5fOerrvLIMkhFWWfPQz94XYNmlB1WcY8FBi
TtOyfkBS0rJMKRKMl7ab0DrebZHSy3BmUt2si4nBLVAj9gaDI0aZTLtX5rEAObMAj9w3UmwvsSYQ
23iPhvdQgOK69JVZPB3Pt+PP/Sb8VRLxzfvLXolYbbSGr5IELwMrcNqecj2Hurt8qfZ239kkoII8
WUIO+ZkO5hvgXNsj+GjkZ7TGwYKRohzaWunNpIes4c1TZq09f2F3s18/Y3AmlhR3cAqxzpVT3ed2
o0xlc3RahM/lP80C81UGWwMs2JRHIDQyUl3NYpybnYEViHnebQ9YfT/1r2L/aDbMMz0XN6aWUG3C
WzsRN+qhM+OcZQjR9MLNkSFsKZZ+ka1L75pAhYBJKOym4+yjS8w2a7LRwDQJiRY/No0VFFTAugRX
49fNAKzxUNpcuUMkaYRVlR5Bxrrph0Fc8XWgYPSf1cylfNT5Xz+MZdb8vSImENNK+N56xSYw2k1X
6I7i6lrTKcvgFJB6MTkg2vihktBbLkechhj/32dclDfbJtjgPwvgIWjYV3ZjOAQE/0R1rVOWenpW
38/H6QPQ7t+lkfrLXWKGHTl897et28K50QHVuW4tTIImldV2iBH7VNtnAjP9NYwcyfoD5euhuKYa
sI7KJKE0ZRUjcxSQImVOlsEs1rFgvNrbImLX0cc2k1DbC4oa0hnCL3Ba17P8eRivlB0VM5wcB3f+
V2fkXsXstMV16KlM74Ab0gKFpsuNVhBUEr72S5gntERyi2X+mqoQ/KYpWC6iv++tLRRrFzi6g9E+
uHNPffzlusfQxXI5mg9Rppj5YLa/9Pw363QZNvtQHL5Ar4REDmPc2NqK6GSDoTSy+TGyIKMuGogF
9zgumRzMEbLRJsDlUkA/nU+uYIYSxBv5KFOyr6acbImxDKaR/FAgFhnn9BeHICpRhmBKXbslNNyY
9DzIWLyvFF2Mzvqf564hhdS/q/57qW4T0zElw/Moix4oqi93mAkN6k7JDEo3iSlXh9SWuJWCO/k+
s53uYi0x3Xuma7QUuW102ElOIKvor/q+DIkyMGjManOwcBkQT/y3y2BeyH9+nSWQLLoNw1yryH6F
pExv9S0JSfxZkTS3aLQGkNiPDz9Ga/HSwgpTqMgjdiwxn1EobpMVCqm/sHtDIfL5cxxGpUtkirAJ
M4Vu5O+spAOmMba+EUgeA/4yvAck3gNg8lJOwgUN410XAdpstOzUXKrRi2fIdc3QAE1Ujl0L4Zjw
qwb6SmQFuuiO9unhnh9eAmlp5ctzJ0HcACs5eSr2R2ySTikNJ9Szar5GvzLns9+7vch3MsaErhpA
tIXjrBnFzgvCWlW0vzu3wzMoUnHcL31ZmyP8NbYhG4aUYthOTGi/7MZDaD06D6t9pgI4ziVUJf1K
7wzDOAf1VQibHD5JBsyc2CrswYiLVNlNR8jfSpCcD+buIpvZm2gslOIptu05BOoY4+vYxSn/QbJm
gbfDUTt4GVONzjE/i6V57bOPwykOb/scQirrfdSldZ5vAg5/Idfuxwc2nJ5EwDO/3MSDlzqW/NSE
ZShipPQ2/Dh9gk74//WXBFtpvTD1vcY1SY2psRAzXrIHWWDMLKfcDWKsS+/IuJ9MkmoJpVPzKWDT
hun0Rk38hbpvnc4II0OXlnkGhgWePZyheYNl5eEpa/pz4RlKb8bRnovVeCIPslnhIuiojs7sqOWU
w440PlYd3xVTtrq/YFHJhfwD0W/Tupp7QQguRxdG3YFTU2F67WZsWvupgadXOo3RZu43q4NQd0gk
NgXyrlFhSSs62g70JOvrSxmRnHuBeVcLIl+TJYu4zi9cobH2N7i1ocIOHSs6NYRcz5OXkmHX3ek4
LuayvY6XXgWLry3OIfWmQPJEaS1LDGWGxZ11VxEHmgPWq7zf6FA0WqTdkFSvMVQ/7yW8Z/p7WsmT
72+GRGRTRhFMLJO2NBZ5R+89pxjcy8jgmNg/z+F2MQng05U0xJmYXyO5FJx0S5mjuGv/zmgJABB/
JkFy3009dOB214KVC1iBOxp2JmRDbG4e41+iCwCltftP1YfzwZai9culwzUndtAetU4k/sN9q5Yq
qRJNTySKugvUEa10nEVclSxlJLTDMmFMt5/ISrDriwj2ciyduUUY/OzRY/Cear7VSmlWewiKlZHQ
VXrobIyBm7ZCzEAR5YnaC58XvsepT/2fBEBgWaUL/qwkufP90WzXW3TJOLLb7KUtsWM/mk3p5fNh
y4sj25JG3ZoivujLMQ6VTUgZ7gVH0jOfLu8lkCmF06BQKY4TfLqVgvSPZx9wrVTRWGOfTwoGC6JT
cXM752pcxFc5RPBpX7YggKTHuBoYDzZmj1SORzU+bkeH6KHd/2Eo9wj5K4rqigGOIEtd8I9bz8b8
61KxfGIlzPN38ADrjJFsPYVvQtL5FgXpY8FIyPf1Ji7QRYMBot4KPdmRfTz3ArXcQ/7azq5GgKY2
QHwe54Z/bCH39Ji2+sWDJWQFS7ouKBXko6odK8pfVWpZMdgae8SIROOG6A+sCF5fMGcgmnEgYfxa
LG1YpDndjc2LYH1tBsHAQqZolW7hH8+wuZiiNRP44qKwdCLHJJoAqd6KYy41GOwZD+9tgLs/Xz+7
xSkxOswz5qR6BKk1aulleo9pYC8T+ewrNc844dfciOzQ2fp5fnkAgWvon5P8xx1bwhB9VpZxWBUu
2IOIDard6XGIMNDA1G7U37bv2pOQDKYgiLf0FgB65YKzqxMRUC0HgXLn/rX5ShLkLKiCVlzj0aD5
KhuUkgl4u06xsgKitw1TR47AlzS/F3imDHpB7C1SmCaAHiIvdZl9xmcwK7c7xh4eFYOHiVmFYGRM
tzXc5r+YCT6W/QpidGw5CfXQoONVKxikJ96nq8eD5/6zdfBBYak6gK/X3Id2c/KtvFH9408c3IHM
qxTl9vhy7cS/s3ZRd8QlL8sRNnTN8UA1zvTjN+dZNIT12suGfTP63OIUgnphBnosGzMjpqWNuAGN
ts+hBSazDvmf1GhMzzg1ECxvumRWScx+AuP9ffZjchvHIeHSJefHBay2uqTmjCv0VlgW8Ker83PX
fjgl0LQ43yXJf3cANyUkkyxjK17T0rSbtMf+SP9vk5uy5c1ZDCy2WQkQwPYI4aykZGhhDfqvgjyr
+1J6qm5jFpoDlOxXXjE8LY1ajOguEtL3750Id90JgjgB+eVJfcqGqE26UEKyjHZ4VWG53d8cziOs
1z3I1a2NDbn5PmqJsQHGKNO61aGfgUavkDPS+T5nE0qao23VouK5JRcRrABWV+S+s/iO11bU6nOR
Rd2+QxYxwpDEMmqP2X0E8YQ0Dkuedu1Is3KM0Z4BtpJd1cWfcmIo2Z3jkCJ51guGsJLocnrXBnKL
2RmMkKKSuFt4hUu/XWHaAnPV8kbIAjQWy9EsiemHwXWSS7oGV87IjuucolqyiWgg4F/EMpZfiY+g
MAUdR5A8202ju0kuyCSB2HEgrm1Kk0NRXUSWBBC4nt1YcslckURWsFOMORmc56i+WxGwVjBEHFJQ
Cr0QhKuE2v0qJL9EudLhFAgDiFLsmpGMjXqbqRw4VSnS2uE6j4nAdfPi4GCHBsSebKMu392wrPRE
2ipsBMaOGzk425xyXMbn39WYSElx/dN1una46qQrXBEg2My+tKaTd+RMMU1baRc4HSBV3A/2Oun0
/wTmXoWQGObtUXGS67xVs3sRTh9FIgiqzuw+RvAGG4f31Cm+1z4+uXKEnaXXMFvtWHoGH86YIaKD
3Ahjdq4mc3jGJc4tEonlSDeof1c6l9w+/xQCoJ65hzwQ8eB6OtMYsk4/9yvsRhG65LqnhVEzFB0i
9gpQt5ylpEVFW7EwzU02ngU6HKUAQVxf9uRFtY9uePO6xm1rPefplQyvIORhLSuUjS8mq2NRUnq8
4mWJMSjNDQKXmfMrCCOtAQZPEFD29SSc4pfS8xe+l9d/CMpQnnXw+N1e3LvzQgfTSqZaz+ZeHAAb
/yXSjJ3U0487hltFrHoK6HCgfWZZ1biToWa+v+MdDNroXInBxG/9v/JKWHoCZ402hlGgm9JZ2/kV
cfNLS7Y47bzD0CaQ7krOrQzabsCqi/XHc7UteND0xgeu71LZC+4r5h+QmmofoojLVR9EXIQaMQjl
hNzhdMOYJDrhUeSA3Qv36NgsUr9XSu+8U7RRlJn2A+knnb2GfA/GGb6nE89wCL2kLSOOEmx8SQfw
8eBTs+lWZM0tmYMYg2iLF/2dhSawbLbSL7vaX5g5yToohNbao0Id3sSpLurV47q/Cz75nyQBH+CE
xBCrQn9v1kLMtgTeYL0eNfe9/62G0qwBvGScdLZKekyH/ytn0ZMzDONnDXkPobuieoM3FvfDNSx/
ES8+W9BJmQHmp6tz91JTD9bHk9I2XdGYgwGRnUP1/97heUD7uX2tjw8ls/hVAcu1dIkWH0KT+tVy
RgSkeueawkK33kFzgvvcRdR2Uw3GkLd+3TK4OJbRcO6qIPC87AL+gpjvwWlI3fWtBj162Z5dQyPz
04/7HL8QI4fTgRjbWFgrMozG+XnxbhhEbqBb7HRxho7HcHFf6NyHDCiTvlw9kyoJ2g/T3CI7Niy9
txQyFAS2T/MeMTk2AB1r7DgrQHesUMdFCffS50j11Y28oTkNrpxYjvMQHDdnFSAIUI7vHyYAHpr7
pPBTX7PoWJAZ7Vtik9Rc2Jre6bj3065nIazifJzxC5MNM8Z7snM8dBDZFxWZGizcxJxO5q5R6Lnz
TnkouQYfouVBULBhX7SuA25gphRuhIhrpbtJml01NuN2Y69xsI1FI13tLZHl0xAQqtbEekvyiCE/
xaEBzqoieSv6BQgn5QRi49QWDfktl9t29ENIoMsESycIfHbqGgSV1G/mRij9Wy0NTPLAbolTaS9Y
Kt++x5FNcVFkJDo6bMzB1AkGYCysd9Fi2hlm5P3UVyrGCmOe1XsfbzByKv/2+feFMU30CoO/J9WG
zgYIO71V8MA4tvX29FsvJjP8HEXX0BrcT6TojOe30I8jxtfVx9KTPhDQeol14RegJmtAoSVm25PF
or4bP2wJOX8D99c3IpWRz3GpjkNY572jUrV/qNRWn18199gcNLPSDBYkE9DIqdgLeFy65Avke79j
TB5EkSw9oGkfdayB8HBfPrG6XKwIDl6RcHLCUeUxvFcBF7RRygLq6nxBmW0+pJukSDcOGnXpoKVu
NAA7aj99AtKsSOJeFpgWCsnXYZ3LQX0PsrKGoa+8PtNIT5k5tVW0gYe3oWn6XycXMkl9LhBpWv0T
AW3PlPpLY5Odfu1Fkh44le+oVRL2VBJH7Kk7Q6EYXxE2MmMQvCa0IRhzEd8sh7LUEqrmCmY78F8C
sGYqYHTrQHyU61SQXh+sgaTzfisGlvt4e1c7mxyCui7girqVtAJw/J1QsD31vVt/fUX4vn0wMjsU
CrfyDzlxcrtxpDy6gx/nbQF9u8CpWHiQ86+NfeAtrUTXNuy8fo8Xx80BFvxBe49JOt1oQUOB78v0
rsOXQ1Yx7IvLdD4D7TgctgaTRZnWv6OMSWtJnrCXROhW4drwrpHGCWEw4/N1gjeoEb3XorrmrjI9
68dH8HK67iD2hIaQBAYzfal6/ujKzAsXWWg9GEFxdWlUhXEz7aQUp7FaWXmloNfB51rN7bJn3ePU
oG8cYEdQuCqoU4sTqnjrgBWI/Si9ogWZlbjVXeOgr8v+T+K15UtI7eUKiyydRUhgNWdSETfrav/F
ph+vTE6n5rkbwy6RT1QnkS2vXG4iaEf8BLDHdwf5PNS013VhHey6yt/gOxMmPYdjQdakx+Ibph9b
XPwZauW1svE3giVxvJiT/kv3/2XsvIxbpRg7+y7fJZwHIU22Kco/5i5hFpcAg0S+8+2Vpc67N8oy
G+Z9PhmJ+pyOUMar1XXMZPKtoA9/RMhnmg1JYP0VEPIYOeBloAd1R7Qz775I0iTtJ9Mb/pkofTOB
5EtjaBtyJL7qB3AO0UuxcejopbyuxZno6K1StQjxHsyBMk/l+J5A4bH0NaASuinIRWRaDhwQwF28
9SRQqjvC0ogQXhbiPPEpYN+4qimboZ49r4eBgH5v7EuKrKSrowf9MODT24LjKxlVy5Wmd/aiyN+B
lkEki2cn7n8bltK03bRnTwbsMRee+k9PaGbzvq6ACr/EGjqr0dcsSLYJ8xcn4QgUsrkVpgZlfHCu
NyfjLIfS2jegtLBwHAsMn9Um5dpgIXf7E1Jg3UK+Ef0LTB6f8lv76dyaX6D3RedaOEJL1nO38o2s
MMqx5aMFpFKgdMCZZjIJrhlmjc8/3svVauZP5N8j+SHUvEs9kobdJ7L0ye9vhDkjIciDYec+6UHP
49wN9bJxpJYbYB2B6t9KuXW3kxVPup2uoNxK8FR6bQ4de9bhteJvexvEHmeegpgVVdh/WaH/CBt2
V8Y6uRxWDUfxU3UWcAsy8QqvEV3pWhD98lvG69B/vD6ONsuEQdXvquAqY9Gk5hM4Ed9BkzM7z908
QW4wMn5WNDLR46fMD+qe4wszP3aB0ftBbvHr46NXph1c1oOEVZeuTqByrjxtytSmcwRNIYJsQ8OR
8cwW5PYaZIR4mP60YevL3/wJr4f1KIsPZmRKOc0uwNroRCIn2xlHLBqhjR+kkjGrN5BHnVOkO1vj
ZKlIX1ym2oR1MXiEUfjC2z08U42B4ynAGo3967QRTnfdGjFC/7HCloB7kfcWvIMjv/7qnfgYHqt+
rNExWY0aVW6Ka3chs3At+2lSOmmv0rT1nJoyxQez4Wt12le+9xrK7lRWj/OnMApSQU4JvZ7Am/w3
Y4qoBJFHbA4MryUF+PPBcy7gfMqNzsYeVsscUnWGwosVQ5SGQ2PavoCZD6STUEyko8IxZyZ6PI6b
c4SD1dYFCmNAB64I5930TFgIHmjnqThpGjFq/QLCWJ4XmMjKih8zVs1zOv/1Pxq1hT/Ul2b4z5jG
izyQFxgH912YEuHKe5uDQDtOuzeK6heaJ/aYGn0di4XhT16DxaxTj78YswBI25Q72bx1sS2Cw9Bf
Sm7K1jAV6X0yXOhRf4QJj05KPoSgalLDl9blIVzH4cZsUcnlCgOa7R8gMt3DQRy/x6ukeBDszroi
Q8EDLKEplYXNxSJ4TDez3DHnYYSowatvKdWL1eaIsTuM0gNsS+JcKMq9nQrz8Bf2cdYR5fdI021j
Qs6u9ArHB8BQdgShBUOWNP7syO+fXMVsrOfK8ZaOoid/7NyiMSI9vvWE0MXYSvg95e6PbrSdg9F6
3MsPuTLzyAlzXT8AHfClUHuNMDezXjlK+EkK89wUciGiaANAyiqQe+Z41LAhas1ct+PDRBLXWeTg
N2CaE+EjUtmtJxWu6Wg4oRGP3auHk55VNwqN0n5K9vwz7RzHSibWLb8OQfT/OjNmWNmajLJ6l7WC
qzyUK5E8Z2PlXv5R1fpXqyRzsNz/lKDZ012X4D1LYuIB2ane45iYpWZEoGu6ZytsiExjP+m+8bDY
0mIGO+Ohdi/JTUpZp97fzMnBgrMt7K8lUQpmitDPTzcFi8MUv6I99pqMUTSKo3MdcYZcWiuq8DNe
AknW8vTESwKTsbMbzHUTTZ/8uZpeambHUGuIBfuFfVKs8jfINcQZgSa4I8a33qKVVoyCDsM0Q9eE
9O0ovzB5vaYeZIaKBtU96auzlZCbon53XG64d/jGnyqQLWXNLB8aXO9zWKAOjol2kHx7kvv3+mZV
IRwob74QGUEzwUKS0ERikaJF96rmQ1TOJzqRTi1O9+DRt7gr5QuT62JJZykVnBF4cbPbBGQi7eoo
9OEBdvK8W3nAf6E9G2Xx1zVllojrZ5qbCQ3BOmDOHuksRzOdA226txFsp6lOjYBaajkpHvWr6Be3
1H8OiM0fBCztMiU9r9hWhoXDD83NWKmy/TfGnxfLgVDtoJ3xqT9nsMBf/SzkDipN136Vq8EAayxB
IHPBefkiBob87F9b6xcdU3JNEsamfjGjT99rYqFTNYVUEqvfB4FVHO9UOsvGQSsTxRE/EQk62jE4
R4LYrLmYIVMC3ICv8NvG6koF0XTyiBkFPncBnqg1J7DeGnUuUzMYb6EmVCDp4oJNbpu9mHw5WA65
LJp3Vam2GY2q1P7fHRoHeMt07OFz4huq6uFfnPh5B1+a7Kq3bamIXCojHS2kCGcM/B1BLd/ALQZA
i+Vf/Mq1MUuPS8Fa+xlMlsZ/mSGcGiKZltIqYy0II19iAb0lTVquNOl1lrcoQGz3RCf9dLBD5Lz9
e5QwqxACtny+CxnU/go9cPovVvsroauyNK1GjpOkoW8bBU5sWO8lvMb0ek20yZmmiPDcfw33z6De
SO0YmJKNGRp1UCLwFaLz0quTzfUsrEf6ODChK/GLkvT+jnhAkWM+4Qa+BR3uVleL9Szt7osq5qYp
ofTkiMffD2jUtmSFR9NJUJzlHLH5jlaMUDpL0HhAu9HgwhyYgZErmQCoE3tUpn8RMkSH/jGi0i+l
cTxqfF730Ix9BB59+V7U/3My1dnQHvL67uzptNVrXkXBQ4vxjDRNrCMFcLzkW9lgld3JQTJTqiWl
GKL8+6pQPEf/asbEe9h9tZl3XYXlBLlf3aYvtMermJRc41/KY95vBdp6QpXcAA/gRmXWOYHxtKfe
Maouhc9WY447v/+GaX8rtZM9uv9IFqvC7uT1oSeRrrwR4GDcyKxvn8Tl/+wzc5qhgPtfkdGbcQmX
bYcCuY4sIsA+UfnUFtIBv0KEnyTMrskd03YFyTU9T5UU75egGpdfdLPlOuWBzDhmYU30IHe7aqDt
HjCv9vpfWbmKD73KNUxm4sCDXOrWmxD7M3ixhHsquxs0A059bYDC/4DYJWAKNnNzdMZLA5Jg8RDg
feamywmDDq/0PuvwYDC7ZUu71IO/ON9FGV+OVwDDE8yVmOz/pMGXyLcVnpLB+tlA7lYW3htt9lGw
VUqWVxPn9Z4yUYUAsxJGTh9ytILupAiuQdiDxicmulNXuK3Th7LSJHFlBA4E6fFkZ4L2C8gDDCk1
wI0v6FBpxZ9u6wn5AJ+VdMinsXDLR2RZrB/iw3VhUPIiXB0TaecuzffasTAn/5Pa9CT9sKfnzbF4
BFLTV3E74lupkFZCb5xNfzcuChD3NMYsiWiaWExUu4o4Fuqf432tAsw7zIRdJywmXGBxFam4rWc4
Vd5Dw0tNH4e9N/e0YuPSfRo2f4If/kcG8GUStX9cVBcvTDe+e4U+YkNuFMDjNHL/bN2v3zZKukkw
2znNmhnqIp77uh+84vhL00ePLn0RXijPrP3laA7bo9dNEbGdZ+1JGyVTm7MGGHlcUU5eJ5gxbziq
Axr1RCMyS5g6wE5Lg9It9ZffOlWZ6kqkvMCttEmn7RDlVwoVtWjBk45/T+WHRYZeNOgxEeTSE9lE
u0Dow6+1tnp1ov1PY9lG849p0MxseuNhSVvsrVYrxSDeumN6U5k7oS1+y5SDr9YgqUF5w1Sb+z7d
VsbgPqDunu+5oIgyoKOn58zDNdXo9d+XVxPkjmvi5CMwxL9M7vCdtrAExd2qVpnCFLT/uvjUc6+w
fPKcCpxpyluSeoBMucdbQuE/0bPpKMZnW2mGuvBOx42QbrfGWiaQJ/wee8Tl6NUYW4DbLvEF2TCJ
M0Sy50VWzZb9oCK5IIB0qSxA9xoRrq/Wbn2v2aXC3373ZBYkgpUpjl1ow6sVYqncmmAbmyREh/Eb
ABQPnbmQmpDe2PnzSJcclfHF9T1s9kimcq2Rop9EdmTEfJasASGHcQYJ/UgovjXIViIqBUStI0+1
y5pEgeVGaQ3m6zm/SR3zwss5xGIweSIdrpa+xxvL3etdiJT3hjLcy88nai6ucuD7kKqLQSaWtW3b
FvPpFLNjEStHp19nVOvHMqmzOaLs5VSWCOF9a5KJ2I2WKAu/9sNV7zm1Zm42KzHsIpJoNtSYYyiU
Gee7BBn2BiJwaA8ZL6vNJXpiZu12gVcO3asCg+jgqkrduIw+cMhcdcA++q6k27tPxDxapDPz9kAt
I/ufvW9jhKZMO8ClgV+lGHIYgn7+BEdAGdyxJPeI1BDgduGdTU5X1n2pO7BRRAIYfBYu4hvYhEx0
XF20t/MTplSHJ6g+3jL/ZPTrZ1UjaoVLypVIio3yLTzNQi9Ssr6B8Z+GsYnkJ2NXBvkCEKGK8Zci
52MNSZv4OItQmpf23kyzkoTg8PC0K0H4nQRicfGDKfgtWBdOtF2+EXgCoT3zgyZz5rzsmmMOfrpZ
vtcWUEiapDogoF/wWLIl3dh9ixgbD+yJy8E6rQWjN8APBD6c6AOm3HTkfj7/RjzVN21Yi7bG0dfm
FSUCwuEz8wJkjH4pE8j1IYnX2iuWOO7mTQhsRqD3WZhfmlGOc2wSfdyEEpXToIpMpZXz7iPSUJHI
wGtaX1YqKwj6ti4P1zzLjRHCbFZaGCWs32FQINgE1rk1rt4pyUWzLAMv9A49ZXXP9uIdW2QxvtXU
XYcBLKEXDyHC8DdaAugapNKphlIOMGW6cMuDF/t4vArBJPReJLb4yDKHmsbnaTBZx67SJ1uVCGxM
QWpMXsEGI2Kwff/DKjzDBbCUWah3T7yNend885wgRGcDMfsaPCBbuYp3IEnZ1qqCyE+U4Wfitgj2
lOr3AxzWsyBydG/qF8rTdp2+5row9zu5O8l43fvPSjsObtFfnuB3yOF/aQYVwUg5uJwRztKd85N3
Odhul7QIAx5JOOhrKgMoX5Mpj0lyeAHY1Ar7M08dxOrrChmsSToSG2J3ciLr9xcF64AMbjUsi7kA
ZAB2u2Zxy3YxcGDiYGdpatJiZQsK3QB26LsLmLFB7CPiMnzBuZBNg1ainv4yyQWA1biKciUB9CPt
p2PVuRxo2LvSlMuhjwexZ5UrZvANXEzl8+giKGC4jW1yCv0C3INLUfckNHaIfzq9/KFhLOaq4sVf
Ks6Nd0Zyar14hMS+8GI0/X1LnhzNZK/SKzQPLiMv7CUbH/Z/neRuvtQFyp6zoCshNcAyhYWuCUAU
ejr2gG8VFxYJyyGCpJOmZDXLsOhXSvqBc8dMtnA6qc8/97TyADQEHN210WiDwEbV7AeIfpnKVA3q
2nLasVDQ+58tr9+7qmIrwafVawnlrxXWxsd2SVMac0Edu33kgd+6708DC5Ilm4/WDnKsuiz7GTAO
8YgJRt9HQKJlPefK7QAK1Uf3lhbZmrudo1ae77ZQe9rR1YBDL1SRH6dR0IfTwNoN3hlaUYuPX3rp
34qPQ4uGeLnZVDUpzwwv/sztPDA1/1/VSMNjasuG2PplbPPPrloHFWlRLP2XKx8P8pWhcEkyJN3j
H2Uj+DmLLiCAi8LLXw+oYM7Rnlh6dGTfJaJmMX2bY/2vCPtY4ZVemAPK/k00UbT1qxZ6vVsfrNQ+
s/c6bWmP9jZDcMzZ2dGUCiULjDJJ6UiP4Y26tbMI2dPeh/rDduP5qLn0EV/uPp1p+bOC0UYGezVI
Ra+REp9b9Q2I786o0zheMsWwQPRbQIXgktKVp+pvnz+zVDiH28zGniswx1JfA1R3bCvDhNrB72gr
j/mJ58kdz1vOGOZeER4oGKwNM5cxgOccfJuN5F7F6lCYmSHg1lsCMo9zfuc1sztFu/odtkPSLzS8
H9miFZ9o3HVHyB9rX+JTzEVxB5hdZ57QBLEVerxuucXneVIhDtJOHpnO4lz5YXYLkA2W78Inm1wy
X9jUmH97yxRWw2DJNykJEhdpprAtV0CLZ53Mmd4Z5CFYg3aNgjAnA2zs9TCACQgOoFzrTg8u6i1+
HiWt0WY8Cm21v4TJOtyopVzXvhkQaFL3D0LQ9qd4neObT2hOQSnU9O0GHzMMvUA0FbtEM3OG1Zar
QEsyVy/WJI3L0Vp3AaHP3w1Byv4nGtNTWLVKiopxOzwv1hf2M406ehy3Dq/mVsEKIjhwEASbpNX0
wv37U5Q5b1zIEeSnbcaV6A/bLfJD7NX1fncmaKcfbtpBFd8JrPSHmu38ozetCtB9uM+cL/+7hLob
9lz0xnYeSQOS9a00jdIqfXuKNxPk3LGzKVtHh5cwSSL//Xg83AsCH1rap00Mz9iN1zGKdKnQHeje
LgS5MLTnWeIyaw4CMN4RFrwPhXgql/tR+I9nv+Mb9TK5hjBWv6/xY7neC92h9eFCb67+zV4xMUBp
rM2eKbXrM18zG9PI7JzSpS+3ZxbzSphGrIr+Z9RG7e+W3u/nUS63ccon7gcoIYIxwf+S6wMWdhKj
bR6UbH9/JFz+UpSEvC2i5EceDp+gd1NJ+YncsmMghZe1Ia9gWbUUFlsSVoBOoThJTNCv43V20sik
hqtnGk2lERMeXhOrSMbsQFI5nQtWRgknur0D7NUq7xOxKAI8F66fB7NbsDxuRh0NeDkLba6sBT6g
ehlVa3ZPplX1pWplYyqdzkZ+1DYR2YTsv0TpRVelOHQCYVfrvvb6imULT7c9lSr7QVqyPWWDXV6H
A0YmJ79wyDQCPZjVP9gpm5NrlLL2EuFOxJ48Uh4RZKcBoOgo5x1d2i6andyhzDY2Ylh9BAO8nBHT
FlsSndzv3dTnvrub5WjAxlQG3bpD50yCBvNsPLYa1zwEnUqm+HZ1d0d1RsqpazOa6YL82xBq9Omf
TpTuP91MNlcKOH61zoiOeSu/bpOwCXLAliZ/ZDj9KXSnuLmCkopI9XrKSLUsO+7UwQdAqG/mciFD
IEECtm0uBIRY2LXKvKwqRAm82TrMgeDHcKNmERCqXgOz9JnT0KUmVRDd6thGJ+6Uf/3YA9ubPqGW
wGlMoboLeUsS+o+zp5bv3s+MwaMoIckwPXvycPfBtMlOkmBd8w41GRnlQmH4vLdwA+SczeGhAd92
9XC9xUspEdwybSqtUKYbluGsMvNDTI7kvIQcT5OYaspYI8kmK9v0QkVoUXmYR3VShTGW+5KCoS50
cZ/v8ZZjRoC6DbvIMYuZbl8nEZ0QRHgQ3XdrDpxeUWRykW56A4vJ9J6fZLoLQ4lWxUJm1/+403Oo
hSyTlrS3icC/ABF55u5zXOuEwQ0BTnGBeuz1jmpxLT9XQfs8H5FCvKQyP86Zcd6zIXU8xpVTSS2r
zBvs71HvLN3uryD9daQgYTdLvEUxA94UoQhm4NNEDKLTmys3UQJlXKHfGC7hUZCPf5nLQZ8toqT2
Ea3eq9flwxbZ7VoaSk8SH1n2fFzFcSivP5Dj+OQg0d91fEEt0ZBdTfVLAiz5cDbCdZISyblo43qz
+XsC21+XTK5NUhQnwbIG10BNSudTGETmOvsXVyfHxVNLTM0ow4Rr6R80E0/YjcG3+9rXnUeatbjt
oy/LXcjWVyDtzMSI/lf1dz8rmt6dCx7TjWw8J5oKt1iwJlbMOSDNefSx+y7k7JwtoQufFtiqU2dl
mdkjUxqdkFeMWIUSLil1fyi5xQoSM6aZh88I/uq/MOmxCKa+1SzMHpJC51Aq6Qc1AHxy5jEy7KPI
WYdHIq1Lv5U+/G9ucwHdYG7ea46G/dzynIr5TZS4lmjcvT+m0979YhUnEaVpwVwNKyq0Rq008Zp6
CRRW67pqHyWz3OiQCSV45fs1S7LcDOD8eO9MXuCB9swSPIy/R0xRORrkl5MH4QSLgveeUYpc+yvA
0E1IYVLHBnunRut9R5CjlF+n+JsxGLeCiLnHoLuE7Ez7dcPDtBxsIysWfmy6BbjeTV6BGkshRsLj
3qiN4DW7fIBac5SXR/Nm2x/DThDXOkZSW50flMVqHvJ/QCo9HLus9DynX2hed7t6PfDiZqv2SsIz
RdsIdV7DZr4BK3jgPPJSaEXBtJ1pJPsp8eEZMk91KhGFHPUMmkSLqC32Bzm18pfWbModvf4Ph5dj
7gGju46a5EckksAmKvFLXWUj9+Qotp3ycEoEM1PWJ+2PI7K8T/CArZW77fnybOvsjOoIFTurLwDm
QjmfxrYEM9mPy9Ya5gF4OwyPi+/y2EZcIlWiwrdyWZGlud4P7yaK16fA/u95VOFBjS1O5qn8mTN2
gr7LFNGMHHfTB+anJzmo8hvefcoyhqIsTxnDQeacY5y1TRZI6Kgfyiv9h3AVuNDw+3W4bnmQwpGu
H3THsPxoH8WNWHOPTMRmJ/GbGcNFL0QYI0EgUQqmTM6pgmYGuS51XyIT8Ekpt2Cund4O3kooxvOi
+rPa86k5fflAG7TqVKImy7vMAuEPCcZJ+lLvpRD5z54Dsp//gSs6gaNoQRDJ2/cYn9jB4Pn+5Ggq
nC1F3ZIj2bcCqMZOx+vpembD9H4HYJMhIhByTWPb8kRpVeX9t4YLZy4tNuYI2v3xcJW8xkdM3qKt
s9KYuGCuBMPTMcZuytFSyUwVLme7BTfbCr1njEYOWvDGljfqpAq8lifkEZSgE0/EPggaL3BciUdz
ZMKDMQu9S1XCtUWBLaJXk+rYfeCLC7IhkO7S4iWhmaO8rQYb1RfWCR6gJ3/O1fdzNt7iKa92YorA
BHy6590IIyGcNYv+yAKPtxarc/NQzjotK6F/Tc0/eilFA5JXzqKHLQnIoMCoyrZ+ae1/eViU0XRb
Hev4Kl0RY+g2xjSTTS5Hj6yB+QHyNX4jH+9T055bljv/rQ1rC534verF0x8NOAQ0KkabNfOULp6w
mVN5m7jMT2y4nIlm/BRcxXjFJx32J4sL5lDVoEREJnI97UFvzjb1S7QOIweEf2IW0Szufgmncs0v
HiW5ovpEz0SuHOeL5QeUbF80d1FAnW1mIlWtW8lbePSr5qk7EMbWtxyESiCweXNYmLMDcUmaHCZ9
hBCsx6yBrvSf7ndZzsIVFeW1TdsuXZNH9RiC6sCbwTLbtUQ2U91YjXMKB6+YuPetMirGIl8eLNOX
/qcKXNRJ6uShIbzulsMD83uU7+YPW1hj9wW3IVL8gtGhPh2yi5BKH++3Xx2x0surGAyfuH2TsIt9
ROsY+1hLj+QE9XJe9kPjjRfvbkuyESoNJehYvF5B7INEqxW/Mk/g1BD+nzqOqYCfL6D6z0c/RI7s
OWeKR0W8pcCz3ilfNakzl0OZZkOXyRofrp/w6te5VAEuESt9BOVaMwoeprTUbO97gHlQnwxktaBG
OSBly/ur0lNJkr8TMxDMI/3Tx2EZEaZAlwlpZS3xP/Y1ZaI2VRiehNxGI2cutJBCfsC46OTdTlvq
o2Pe5xx0R/cncnljxTKoGgKppJM+fHV7DmSvxW7GAfJ4TuysPfa9uqP/8evkjHqnLaOYvaiY0j26
mtdbhI7pcKOs5BqZeeUSZIem+nfYmhj0YC4fc53vhu0UjGUixm6ZOTZCE3Wu2IMr1gVi2XB/e/0t
WDoGNfWd0ne0QwxlTGY99CWyCmvGDAPzojGkN+87L9UlLz4cEveEDlEr2fN3qU9jKadH8+bUc60E
cRX8pkjS5zsOH0OK72bIAbqkbblot8JVA1Vv1Yf3Xc+0fkuQFrINJmzgMCwHTCh5eCYXFiIOAeIy
bxgJfoQdtRcJm0dhGjjgLgHjW2xO5SQdHNZ7ibzYtu3JlJG8vntnxRaMi2KCPshUKPAonABbiu4x
Wincj7sTh34X9qXkLyVEwCoEcR8iw7vPHenx45jjBbHn3onBGPO4NfbpphONeLUT3gwGFlD0s6Lb
Srpvn/5heq3khCyOj78xkiT9fc3TkPfNBGTknzvbhQmJqD5RZ7dHDVAj+oeSvHSlGn135nWQQq4A
EYf281Iy39GW9iZTin5s1rtuipyz4CJUCFrs3eqfqnM1
`protect end_protected
