XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
� ˟X�{*�J1�u��V�Y;�!�/����(��csGcbgJ��/c9�9T����?���&� �\���P�[.Cy��ޢ��,�O��W���|��x��a�.)¤�b�b��PeH-�J<�<�A��q��`�	N?��P��m1}�Qa㯳J�s���*l7:�w�̑;`�/����aݠ`��uȎ\Q��B��p(d3yA��a1	���ʜ��j=�� )�)T�L�邑8<�+^kCl�� �
�~��B�4���;k��Ui�g��D�<L(����ܕ���$���6�y$%��g=�|F���8&5����o�b��Z2[�Dv��uw�ա��\��1�o:�V��+���I��H��b!�=�i�T�݀<���4�1e�i��؏8�g�p�˺���=�XI _<=h����h�"�5����B�0�,Ȁ[�񁘉V�!q�Au ����~��v]Ƙɹ������q5�{5�P�6��$Lsz\`V��5����
��ʼ<2����[��b�f�c]+<4[�PPy,����c`���U<]|1��СfG��Y���?.);���R|�(��x2 �)��V�fE�>�J-�2Q�c�a':#K�E��ć7��]���f���_�ttqEH�>ܚzy�)cG��{�Uq�����H�]�>�A�3�E.~����X�c �)ɷ��y�x�U�D���u���/��Z�,]K{j��G��%l���yqm_H	��j2�#�}n:�]V�a�q!������c:�BeXlxVHYEB     400     1e0ʡ����K�u�d1έ3:S�	���K�t{}PqЕ�j��z8� �0�}\�WE6�5t�ʛ.@! V�R�������(��a���?�:E/�N� ���[堨O�H�ͧ.B�)�]���^`PA+}��0���P�]���Q�ZT��~����
X�ZP��	�ݛ s�Nۋt�u����z������M���P�ŏ�8�?m�!�4��h�<��Z�-lD�*�c����"O�o�=���%y��f*#)��X�+`���(���}�롊J����.G���C�1�<�����7�0C�P��E�#ܠst��;f���Mk�!�;�_�I�)�{�tuk����Wg%� ��N|x"[a��-�6V�qN�7
w=+����(�~�c��2���nZ�XR�n��\
2�Dۘ��VW3����3o�w�ߨ;���>v>���GrP9��W(�ѣ�S���S�|(mP�T�ePj�XlxVHYEB     400     1a0��JgǴ�@��YX��)e�����3Z.[���4Έ�n�����J�ܐ��G�z�f�N���?~�F��zn@�{	x� ���N�g�*��#�4�R�E���9�Bg��Ӣ>I�B���U��|S
/��gw��|n�h���jB*��._Ƶ�J߆0`~�O�xD�#��˥ދJ��̄��>8���<2�'e_9��:�r4
v@h(���A�c�~ɍ�	��a���'DX�+������>$�.&�{h�б�Ckeq�M�䫰>�uF[NO����sr��̃�C.�'����Ǵ�z+��O��)�<Y3n�"v���N��Ѕ9e�$�ǲ����enH<2}Ī�����l�
�	�k�W��!8`q���P��q���Z{�V��a�Ζ� ވ�R���{'��jȰT?��*�P����XlxVHYEB     400     130�Z�P��鞴'`I���\#f�^[�u�k��v�ym��<^���.�jn��m�b
���@n�	�^ڻ�%��HV",#=%I�ɜ3�H��������i��];VxCm�z)~ڈ����O��甤G�	~	EY�n�[�+`�#�	ګ��0��F
N�)�� �<�񾶅���a4딥iF��'�Ax�]�	�x����l�9Y�R,�&3���G�s��;�:w���4� ckf�N���K��7�i���p?� �D_7�fC|-zo?1K�G�aT�1o�Ŀf2�}��iWx�s���K	M@L�XlxVHYEB     400     150����(:�XF=A[f��y�����zv���udmj�6Ұ����m�#ԧܖ|��:���ǒ�l��K��{4��R��91���g�Hx@񃅠�`ߨx*���/���]]��D���XG�\��7QJ�-q[�`�eBoQ�R�����	H,h�۠�Z�N>,4���o����fh.z���D� C9���V}���{�P�}����c�r���V�Q��W�9��/?��G�:,ol]Ǣ�V�.��W�|?�"�CJa�2�M30���O�lj[�~c�7	�s/�Sc.~^�h�M��F:���L������ȡ�"�#��-y���ZO?)XlxVHYEB     400     1a0���W����tʵ =���u+o{�u]���(xct�¤���ʲS�Iҹ_��
b����3Mi�i�T�l�ٶ�1k�p����j7��U��{�/���?����,c6���%����B�hr|�)tC�rPɟ�̀�����JP�%�e�O�K�����X_V䶖,+2xԻ	a}�Ͻ4�I���O���1}�0��mO�t
�K)�C���p�?MꞐ*��S�LC�3��L�������`�'��dDP���s��`���B�<���c�g��8{��pƗо��/���@��l���O'�T���s�!��7�TB8Q��kb.�#�]$�/Z1�B����xW�ZA.�=g����w�j}�&�{�M��&��o=�p�n=���6Ӛ�m�%�>�4t���ku8��XlxVHYEB     400     180%��L!h�ϫY�>0пϲ�� �ۡs�W�=J��<�][FR�҇y�.�݊z�г`�����5���T�UZl�� E�42i���U�>Ji�1bg.T�WԤ����S���L4Bqq�\l��F=��%@��d�C�-�9ʦW�e3��#��`6��Q��[ט^��ο埉�w�V����ce��m�jT����P�e�f��n���[;\%x�UOU��]/�ꮌM�ɓ�M������OD�+HWE$m�,� &.ްj��g�1"n>OUE���~����ޖl0���ʈMmbgx8�y-���q������Q�kD�陑p�v�J^��n؈�=�"Z��N:l����?%M��� ՝�&9&���;�
���XlxVHYEB     3a0     170�\���D��Vw���GL�e�V���|�
f�?k��WԶ�����v�.ۉ��AR0�N����+Ă���n��_�q�G�&1�w�䄖�9~N�T���������$Ox|���%v5A("#)!0z�^���ej<�*yO����+�[�e=�bJ���y^|�4 ��/�|�W��e��zd�D��$	ǭF���'��׹7[��K08� �R����u>�(���}.T��'I�셞*4�O �Q�г���X�e��ŗx��yg!���	���L�����v#r�"�t�%b�2>h%�=x��f����C��L��z+Ң�n�����?(�/�8Z�&�+��:pn�t�5c�e�ҳ`�[