XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R$��@
���B0��Ŧ��x3hIv2���!1�p�B�`�,ő���g\��E�.���*���>s�7\�����~�ٞ���tB����N�����Ej{��?����9�F�Ma,���<��k��-�\�ˬ%cn� ڠjL*n�uJ�*޲p�-���f�T��C"�vD�\sU�{�ߵK�#çMc��$03���y��"���::ڛ&�=�L�ZY��S�a�����$�3|h�����$*+����p��g]�',��}�;�5q豊��M@��FۮZ��v�i��s���S�ЬT�iX���8�:l��ސ8��[���
�^����<e���(�iV�� ]�KX�n?���>��
w�"�h۸��aE������R�-�R}��G�;�Lf/��%^Yb߱ñ��mGG�ҾwH׫�x��[d�j���!Rΰ�,��s�UC��Z����j����M)]���$'�+�՛�Q��A��k�5��u�G6���|{�2fd����������g���w|��ۗ���b�D�MR�R̃��I�U�N���]��̖Ś,T�Y�q�Pt����33��|1w��Q��6�s������t.Am{Q���#����_ę/[!�B�����B�`�Ka�0�}:��n�+A�sʃ9qc�6�z����P�#��2�QC2zx�D����<��kq��Q+�'�U0��'0�M9[v�>*��f�f$R���4���a���u�t�ʺĺD��p&�V�\��ųXlxVHYEB     400     210�H���.Y����~%��#�sZ�A�{T�	t���Jb��-d�$�Jt�j�������L���R�&k��&de2Ar�6
	�9�΅ޒ��V,��!�S��;�,s������`>��_��-O�*m��t�0�=�Ld���?FB邁_�&^��[��+��gw:�n%D�5I͵5�Ջ�*�� �
c#m��3�����׹��yc���V�fĜiQ� ���̫��~�#�"�zp3�T�|B8O-લj��X��I�����q��[���Q�����cR��>TƿF���)�u��H4c��&r,XD*�Ϛhӏfz��i��y�l��:{�g�uY���"hY�] he��h5����
w��}�����p�A��H��~������{kҞ����f������Phw�nUB�:]�������g�3�Vi7��.����9.=fE�#��z�IJ���w�)�F�L�)!�����L��F|��	�O�*�� �/���D���p���N�-��XlxVHYEB     400     100꪿��3�[�V�U3�)B�4�D�o1Xá��I�"����ZSq��5���v%�V�M2��8�cׁ# �� 3.�;E'u+����ͤ���?��s�xU��k"Q"��HI,E�?������(��F�_Vgᕇ�AR����:a%���L��D���`}�0�zF�G&��61�,@�י����a��k.w��S�e�##� �ٚ¬��j�4�۾�Y
�	�� ��E����r�;��s}�l��G��XlxVHYEB     400     1f0b�;v�-4a+��y�����m��Kt�8��t���֬��;�iO�i�p�Կ@DIN��0@;��[��z���r<�0Ϩ�r|�t���/�1V�K_A�믛���T�J��_o;��u��� � 9��E��JE�L��P��&;5ROF*���1`3�����]2g�R�$��E���ԭ��B�D�J8o��D�1q��p�巻�.I�[�I��=C�,l懝����V#�S�xi���1��Iq#�M;��JȆr����D�����d���"?p3S�`�Oxi*K��k�db�ct�?8-fM�7}T�Org�m�Z|KH��1�����0��䂠��e�i�J������3f�М���6��W��^�$z����.�D�$0>jt�������^O��ҕ#!���sO_2���Yl5~��\֗��Z�ґ��w�$Cd/yn�#P߼��I� �+8�c���*�n�ͰʞՌbK��`�iJ��?XlxVHYEB     400     230��0l��k�&`��xjuַ�%��u\mh��O�EO1)"@�PO��;a��v��Y�5�\��� ɓ8��H}0��{%���`V,�k�x��a �Sk�mAO��
Mb�=^�8�DZ�e!S~O�]�-�ϸ���O��N�1���JR^���J4����G4��CWc�/���	y4"� E8a�N�|����_��m��=$ާa�$��]h+�d�C�z�������r������8s(�l��Z�<{��^'�� W� 
.�o��J�Ѵ�����4C��G�ItLasؤN�*NUANƼկRJ�^Djy~)wǙ9߫,n?���7Q��y�cl�$U�[���C�F[�ljߥ7ǣ3���.�K��#y��X�F���<��w���0B���	���Qۥ�T�&i7��iuY�ʮM��1#iH�d��E����@�#���:��!d(s�`|Ql�G���MFK���eT&:�Bgܮ���:��_C�y��(��5{@�j�e���o�X��VAprg�(�w֬�u�O�ݿe�J�V�`���Bfo��[XlxVHYEB     400     1a0����gnx��R�PŦ�Z���uI���wMH"!��߼����C{C���r �b^@k�F�*Q�I:v��B#6��'�ز�W�S�J'��4�*/�n�)I�8�tQ��<-�Z��|����:6e�c6x�Z��'����.�M4N���͔��~�@�'F�a�V�\[w����"�4���]B�+����ϼ�z�zb�r��|�~��QP���<�}C�'�m����(8ң�H�)z�*��߾�Y�.dj�&#[6R�GfB陳C@�ɝ�[Y�w���o�Ɲl�f�hB�u�$q~�H��)��=��\;�G��
���,��w���
�ZA<Ҝj6I^���̧�pa1Th�6|m���.����V[�1�c�� l���3��U�wo� �>c��XlxVHYEB     400     1a0 ��N�$�QD�����#��x�֎TU>"t���QTv�튋�f)�ȅJ�a.�Mg$V�!T�/�94��ǃ[�\��,�9�b�P'�o��	��E�H>%��I��׋"qH[��n��~��P!3�Dݮ��CR�Ϛ��'d���j��U�'��ܺv�q�:X�r-��F���[�V��G�]���>���L��aċ��>�̷�D�ӳf�e`�������͚rr�T���b�D�� ����R'��`�D7L!M^�Fȧ+U%��)E�,+� 4VAł��̦꾗�x�M�K��������P)��7�J��:��0xH����̒*����t� ^J�zg2dS5�3��V�K��#��-x��#�5B�d���m�n���48��!����-Z<�M[XlxVHYEB     400     1d0�3n���o���]�V�)�gB�|�C�&�1@+���.mS%c�	F��~��̮'���/��~t�M��=�	)p:H
��*|z1��Ŷ��+���Q5^�n}.K{8 ���4�(�b6�����*���R�Iވ��zq����T6Ԋ�\"A��Ē�I���f�y~ǅZSNff�`T���l#��&*f$���7,/��،ѡ�a�V]�
,u��Њ6�?�'��8�9�i\�"5��`�x!���o��m��O��, ����Q}��i��t�dU,�aUK�%���kOg�Iܐu�ؖ���ݩ�����_��j��U���p�Id�G���i«�`L,	LE�ZF���r��|-s�g�� �V�d1~�YT�����Fc�C3�;��� ��C�n���1�׷�"��Km�����wK��￈���=��3aRD���qn6�XlxVHYEB     400     170�g�\������v^Q0�<��D�l���`=���D)Vޣ�愚��:f������RO:��)���>0��>��^�!7�1��8�:��:\O�,��Z@�T�M1q�dS�+fj���1�Z��)�H��sC۪��0~��iY�Ř��=PK Ε���Go�_�'߭� 9��\5����9ୁy�����R��gM�P�UA�B/���S���[6��*H�&s�f����l����0T��
��'���g��[��~'MQ3̓X�-�N��-��_׾�[�KjP>O����8�jX�?�����������MKNQ%�oWaR�!Ax���Ҽ���nX�_z���X/XlxVHYEB     400     1c0W��G�����8�[L�Ӆ	'�+��b���d=y��1>ͺꠁ��o�N��6�{\�mɿ�!"M��}u�i�%g!���K�ey�ʷr ����t�8VI�5Γ��Es�]�0]z�`�:�Bl��0:cMpC�f�y��z�ȝ�����LS��n�3�FYGƾK!�]ҿ�,*xq����K�hc���x-��-���W�u��X��F�To�m��pz�fv�̓0*@�Ed���?�(:��N����l7���+!�G�F�j�3upg3j������ �.-T�q+�c���3+���r%��΀�v���l���F=V�i\��!��ԩ�H+��,��	�X�*ۦ ���w�v�Pp�����W{9�A�� 1����96�:u��?x�\��'�OE� 9�>U��㛙i��0�5+�%�_���dc`��/[
qz"�)rXlxVHYEB     400     1a0G�,g9�E��Ueyy�iGߟ`� ��Ӱ|�0 �A��%VP��ױ!��V��zF�  �ʾ�߫���P�z<�K��A��z>���}�,��@�l�1�T��}�,,-(������Ԉ���w��%h�P��,������p3��3���5[��J9Obo�䵲�j��p�!�>c�wr���$��"�%�NX���,#)�赑�e��z���>6���l�0��=��e(�J$E9��')s HH��jj�*�d��R�Y؉�����8�m�@�(|E�soDn�$�r#��!�8�?"�	B��"裭�쇱��)V�3`�)"��<�^UFܘ�5h��6�ޜ���*�_
��x�#o��a��=�^F3��
/u�I�\ v1K&D��<R&�O�d/>��o�\XlxVHYEB     400     140�w+�{!�c�=~s���s9S��`���b �C0w���gjM8�2�3�G5/�s@ׁ�M���@�V�#�.��\�A��x`���U�i�%dj�߼��ʘ��ݝaK����:X� ��lM��&.��u�©]e	&���*u�7��,����G�W�oǳ�U�ymr�)�p���:C��"+o+�G��D���:��^�;^�ك�i��A�g�90 �nR�u�_���E~^Uլ42� 4c9ia1$1�B��t=6���:sg.�)*%����w�SHm��ح5��Þ��8�Y��� >7�x3}>n�+�l��XlxVHYEB     38a     180���&m�2�C�]7o�6=�L,�}�ʊ��
o!6$�Yc@�ߓ�1�R�G�N|�!�(U�=3�'��^�)xa��^ֆP����N;�@}c	����:,;�E� �((`mݳ�[�⟡=u�{�������yv��}�]����"s#���ι�:q �G�'=������$�̯J ��F@�K4=�[����Ì���Jpљ��b	�� ��1�4�"G����ۖ�"��)ۺ�n����c;���T'TY��jI͝1l嚇��BH�`d��Y��Hv3vJd�D	��=Rϭ,v�?�Y�i���^�r	�u�˸���E�V4��gH����r�?�D�f����w;�;c �?�Kь�Cеɜ}�A��+�)>��~