`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
MPvb9h+b/PRyCkq2D+pdqJqDFUvxarrTtpNofn99HdItv8zHl1RA0iEsTJ780TPo9obcT/XMZHph
vqjuQfuJyn/MLaEF1EjAnXTDLUOpVrTajUw6mk7WhTNgffMuXXkVNUAjvpp6q/dcwQaqu2qTsFSO
SHzgtIZnQ7bKBOBUqtnixDdtuAIUc+Uo68mERJPzE8WO/I5oLuooHAQ3j9Yz/cYM7JQzgKXWh/v5
5y3gb8EFjkIGKyUNZXCIs6mRJsi7w3GjR8GKZg0Jh8fgskCHeL8XPJSVov34a8M7TZSJbtmPOAM2
+XDI7CXqSPAZDTu6PO1orVRIRX/AokisQtoC/HZznzlMUVhp9MlNRdxYgRY+votuYugkAeGr8mOJ
aQaEfzGQSFuHLZccTxSOe87btKRw2D5eR4BlwUgYAwiqWdIx0DOXC59t1eDTMIj2gVgSTbCTJrH7
a6IsWlIXW/kgtDTGHXiMAE8gWszeeRp4jHN3NdrMq1BWmSlINonrfUoUAKHw8c4Aq7pXqTyW9F5J
zufWOmmnGNhcOZdxqvBHWhNxg7binOkI6/Z2mebnpJW+PI4+ZtXyFcZNdzOkwM8KEbz1fEflLf1j
Dyvte8g6Sw0MUVRMTg4GxxbM08g4iSzn2WKhbW1bZAXfG8BV3IzJ3xCPGaF9VqCB1QYGLEMyEe2O
uXz2/oUHN5gVjKf34XkpcHLs37ZGYivQX/LDvhA0+u0QDLERbLrEwSoFe/1Sm9UWDwqPf2FQsC8q
IUpEC4lqKt98KVurj4wUmMROXb76jwlYNU4bDqK+FSQtboYWacwkZPY/P2X2LA5MablEd4BHfGSH
hC8lGbKep6xV5qBxKfJ7g37VOgYCKDuljyy1xiyW0FNS0dpQEUC0RXJ5u0wtlbj1ivVD7ft4UXlV
eP1d9mSIexoOdpFHxuAx9oSqv1g8psMeO9aiUCkMSMpNQTSgW/l2wSHOeWiipESGSl3xRKvmy+6I
fIxZXEvuIv4oVflk9JyLUbWFdiIDuJAp0gmoikOmBgTPy/P92QyyRaa2WI8vto/xvFoUNKe0vkvY
B1X8bX6oo1lDWjESYdZnDH9lm1buRXnjjJ5Sx/s1/gLb3sJG8hYziGRyoR/qDw0n356FmIX2rbms
WE7JDSC7R7Ni7nzPyeyUIA4fGal8dMhlaD2El2L8dQh9Ew9URNU6clcN+p6Dn7OS0Hs6nzXTWEHl
a6UJnAJ4u9//J4mqefTjaYXE1yiFD3XVqfxh/7zkrEdf6WqMlbs7gEVRO3lASQ9GatehrKbXs7Ik
O4+yF/ySrKyxRQrdHBvwLNI9180C7Idbn5N5ysmdtgTBkBc+kqnpoduNbtFg3Bd79ZaKHZPiwRAU
khtKOvNwaxNY9uBHW3/ssnyf4QiDFiF//2IFdAwYZf8ibt3tgRMNS7z3K0LdLD4ML+fCDYVXOnNf
q5z6DUBO/U035uQ/nAuCQI59uS3mauIRGa0LInUx9ssQH6iuj/kbPZmR38ChPX6TTsQ5SPbWnrrI
TqkOpQE8lUytWR+6YoE5vU3533ywORzl8jDwLCtyFQVs7iTtRM+H3fHlVzIQ564KHMzvc6ZxHwGg
jtVt+BgO06YbMgUaazkvyMamQ/PeKA8URLMedRWjG8iKQsaWYaBUSbQgOAGwMBK0xTb+83R9ZXRc
J9HgcvQxpekpK0uFQxBLeL0CpWng1NtHOjFSqRhAeAD+WI74blrY28A4lBTnNlNL5D36raHbqqoe
aQIeuXh5Wsp4zPDPhxsklvot76HuI4xkxHNayppRUloghPIoh6ABvVXvEbk6mR0hd7oK1tNEsBOD
GBd+yo6Mnx0UL5N1hBNF3ETCNRRImgZYdy05PG46RHWD0XFuSZ45YM8L6vPUj6XQSb2sjMzvPUqE
aA7zJs6ksNahKU1Elv5QSUnsEUjwJnjXvgNHvT5LtGGDNdcZzvY6mBRM3xGnJIGRqTlVOY38BoXI
z2ab0P+smkUtSWY5gi8VceEzpXJVs3ToQdEbg3xb/lVQdlR48aq5U67YpSNFGA5t2QPQUWXEVzqb
ZaJSODmo0b4+/pUTwrJ7Vfd0u5mzZs5KGDCF6TG9/IcwZm85MPzOuFxbb244fn5VxBLXabCLdCFX
2dWXfGJcmyDx65uyh++o7JeTyLFJq9aQrIuYDGT89Exf502sNWqpOjgwazdHymCTky8MeLtYs60b
Daex1m/GFkqtNz7o2GeNE6T58kXRIjwKt8bYTUdxAuWoHov96wXVjR7Qf06wA6yGZUmIrP61Jgzm
mh9vSjGd22A7O4WHo6p5tEgd6vyTJLIrowLzSxDR0wQ/iFJCDsZhKXHsQpo/uah7YU+c0jsGgZXK
5aTn5M3PTkIUL9+erAe23uyPvrHYa0ErQmF8Eas+uJMp7zlQAi9RcxpIV+mxHvi6+21oJortS0MF
Z5VPDzBaPcbF+Euyf62O57OIhXlexrm786cMLyEuaRtQdAlZg8dFzBcWfwXyRP5SuMSWvvhkJI+q
vlFmyssh1qhHMdenKfrVZ3x/i9qc2otvNiJH9S1U8jZMhPMJE5FZhw6oiq6mWbaP4hlIauZp+t6o
YgdknGspp2H6Idh5O1iqj0Be/5ulHxwBCuSxr9wWoTd0lQlqqIXzrCMLdbQEj+7mS0kFjuc8T2nW
ZD1k0TuHoK0bhleLRWS5uSuE5EziL5IXld5e1jS9UxkVl9J2vMfZKHv2dpajFho/BHdko82ljVDY
V+TBGVb5jWMfucEwKAcASPilGxcJdsGYmQ4Rh/Ou4a1y2WQ21jgfPhnkKIF08tcTvmxHk9uzkPgk
1rvzvElbM2pp8tq7z1lOx5WRuc1Uhstroxfm+TRJY+/ZwE0lpjqHjdEuB2vxXR+nOMR3kwtU86sc
CGG6jK8o2KPDHYNPKAIeu/fTqq/6udRkaffFExc7EMzDDEb+jaDNJdUNItdF5RpSTvgBOdvw+NYH
07acysSh4HDClcRrKtL8jyxq4sOZEoTkTwJ3F7EyuRQr82TukfSGtdX0k3hH1W02t4dHrQxNIw1l
4puSn2Vak+VBWTL2600/R5RW9merSMRr6v8o3G+9GWGF9mRAZKzWN4Oaofkczz7A5AHHTHbpwjNj
rcEBEtB+zn/543Lejgpzt6V93QTAQasyH0xEb0P+rX4trBURZx8ZhjAO5odrOkLHHzDxZgkbYwIM
HBvO1J0XGadRIClBm3z0gIu4Wrk+Aha8T4qKeZLMcFTCFKqiqL7fwDkV7lQq9Q3geKy7Znb++TGR
ypzRbje2SiQwXjJn6IYcF43rUF9vCXKzmUFTfkMDB8M1uC49x9II3B/qze71Tg/+SDkQJzydQvNt
sWcagfZ4lcWc/59dV2yZFEc8ULGp1P01sUokBTUEjrkrK65gxJ+JyaB33nkjmvgvrUnZ34ocHgIh
F0pmVpsBFWh9oJvP24fy5S1wDrJwY5DK6h5BABaaFn/XzXoT96tjthOTsylKjFXF5egPiHMTlHAP
RUpChTMf9M8weV00eXfy4HiP66Nu9FQLzXVWvggv8G4++NIXSrr/esndpLk75rdn5UBFAVLx0RV2
Oayt2jd6K3IXDON6E64bCxJLr7TUa0bvqS9ZLiOQOhO7BKO1RmvugcjV7qLXcJRYAjPFDNCEH3xx
2J/kU1Ss3LTUCPJqt+cs44oSk5LRnOIOI5mTDvLM7hx/7K5mCVvX692bZi5TX4SGsK4nIvs2pTL+
ycI9NcwH8nElyu2s0mwowUH/sTw4lueGJ+g/Flq+fro8xDX/EUa3Qsk05QjRCN7KXBVFf7WNIDDN
vb1bu3+ZThQkey/waats2lsa22owZpcY+Nyr6EjHLa1rTq7uUpiq5VoyNRt+vTSjHZqcI7mTYaPd
ZcBWrP1Pd5ahFp8W4qR/7NtldpLkRA2CaMm+Q9GBkPgL2J/EQQpHsufyLdzV/yt1R/ZHo8HcmcNE
tjWImOQN0k4v39r4+u0w8q8XW7sG2bZOAoc9jk0TfrHSgl1howkOolJ8fJuVRqkpMNrkYHY2lset
ULQi2Q6yvyk8WBqcBzByj44OZJvYrI8opA0RrlSdhcNYTUi1s2g0r8XqQGxQ2BsPZA7ptEZQWdGD
bBJ2cGLCEMCacRqBpd1lIB+f409j9EvnXCeRCMP/sYFMjUeEETf1CZAKqkD9CAP0JC53G7FsqpkB
+5D/OyMd62lQRJQ1bXlQ/3OEgvx61+VcUoVPiHB+Y4BeCGC6LL+GxpUFXKlvv6ZmyHO5svYPx4td
EnkrmtgM87XVLVHivN6lDHnY2uzbTh7Xc+3VGdDtCR/lytIouWiZk7lh0+EtjLc8xRZQGCH0FfMh
m9U4uE22wMYYGVQz8YZsi+vtGnWNBPSkbSQz20ecwCZKAbcUmNVicGV0K8+uLdcDI/UqRd+5VsMS
ZEV4xEj/lmDO+Ay7boFpHG0SHqz5N8dzoV+VoW9QEeaKRp7zwbNqcjg691WkdR5ANUi8ioEctzT+
zoYxQJlZcLgqhOmMQTnzTq6WLYlWH7hcMPxVN0+6OYlfn56OyJmg3lv2WgaOkuzbIzhOH4su3X4w
r+bTkeCEyusfOQGQgMThFV9fRnN3CW0Dgs84hnmmFaRvIg3tkP5AT3dD5jR4z77ZlDDb4zalsfHl
lLzdyaDhIB9AzbVUo4Q9wadFBIIap91Ow5ajUpZqdqA5u4c6l4Z3wt5QEjT2re5QyaJGwnAjTjHD
cogVauHEi9kMot5tRkbePHyrP7CCuCdAqRfHz2Mo4jUS5xQ8GE1QL37//VlDWJJynHUCfzDz18ot
0RgVWCNfObDB6obYTtZ1OrNbLeenFk/KH7PCvlUfaXhwGfRSnz3lgLx8QUmPjmd57SO8MHSuWchJ
ZBb12eZOZz+VX9TNCTASv8qdQZvKcqvHQ4cjMe4/JqPq46X8jssx+z+ZwEPRZQqlbCPTksTCyD94
EiA7zJo6+SLtIKONKULjBxEcQshM8/LTwLkVQUmMTAGzWoVCz9BK94uZOCTfDIf68yTwjvgexx8R
6rULS41eyNjwaswrGYrfmCctYEMBiCYAs7Ou1wNTkcMl1lo9VC2hAcMzlBFgl+oeFw1L4id6rboz
C7FmWPBi1OXzUHZzy583JsucpM8cnOhtjqxEu3r8oAUiFdkB92QUU0mYWAZw29ZgczX+bu23KUKa
OJNoUI+je4OV3wtdCHppDtjxPNdKgh+yl2ab0DFDU+ga0PBVKb1EZ23LdgP5riVv8JCKLu3aBqy6
VZuI8WXjYc1pbja6D/LoPS6tC85OusgaZ6CTAP0F25u3nAAYUR5OakKHEuuVOu7/8G2EdQsfdoSi
0uuJv2N6G0P9wyxyyfiSOV/c9A76PaieQ7O/196G8DPiFLNFp2EZTskXZBb/Xtf2XXD1LPj5aiUv
PQMAEZk/7izHx4vqKoq/PySwIGURQ4T5MDMnx9eMJAz+k2KlnDEzev8skI7lsXGBLuAlUWVU116E
86wFLTDYWPRqgar+OOr360kKqHdo/wxkZoWWmRPXNKYWYHsf4VyT2VSSxnD8N0zmYWJUiAIHXzpC
4XAmV02YshWcI4NVGmabbbloGpdrvfmdfuUHJhtJMzBqQmihIixKVCh+lhI+NpPREGwu04lA82Ag
vtcqPiMGkL0QYrXLsHhzQMW7XADY+ucEDZrBE4sb9Y6z/q1ZqPPeuirZ6GxjUdLIGXYc3dg5+aAc
9d7irsZYRDMzi/JORx5514CLA8YwmPho5nuR7F2nQpAyM/nwlGa6E7N6z0nwi0BR8X42EFUZzbyy
RQvxYks+NKUXTKJwJPSIyW/xgePGDis3EJhB6d9+An0phdn4FDhpZfomWCZ4+Tk1Cst7m382Fgk/
XVTDyEUtNZLqgYpqtbMgOWhlqb+GInr08j4L+YjSRVt8rnP3pWRx4h4kRsi071J87pV3rakVoPmH
yz8Tfg6i4IeE2LRZBDnA475ZwSpD/2Q/zJhY0YFsk5yI05mz3DSDYg6YP1q6ukSc7hU8+/6DLAIq
RQ6dpICSIXVBUG9VP81pdBUIOSwi21PVeIcetI7PGOuCS1tAPO4IwFbqaTk2v+hASpSQLi6JBVjr
7S0TWLuyhPqgmGdiVAlNXrfw3ZduCZqcOZVaiMw9ja1vrj2v6Or/xPKv8L7+pGiudRVSSfDWPJcW
pABe6VuzxpEOJybvTNVAICoSxIRbbMXXXH5DoUUfjeF9kupAv4LWpAmGlF6gzDSkO5J3BEBti8bP
4mewXE98yqywAi140BvD+xoHwPeztCzxmlVd2wHJ+00AXDKSQoT8UZHaozTTCJjyPaGP2PZCgsyU
rvOox1MwB7RF9HmOTzP/kZZPu358zHGG4iOEWeNPUBdYkq57AKAO6n4dlo3i6Lj4yAPTE3rPy9KI
FhiPVeuYiV3gjJW1ldHUT487qZXcWzuvwO5ETFw3gkAZU8F9B+Ki15bJzgMj8aA8UACR5OuX4okM
dF5M5pzeZsRznCtUNc4iehNHD0hLw729M5/Wnx84Geq/TCLFurjhvYtLc3ZkIOic5H8n+vmvyJ7l
Ml9um0aZ5lDC01P442TOY6+UMvHhTHyaDASOUIucRqXhc/PwsaFQlHJSmNXlHr0hDrDfnbh1Q7yT
doWKGyKROHuwlHEr1TTcNPNQsIzUemfhbdmIVDe0OWYrTEmA9G7JaK9mbrsWQNM5r6iPmfNe6i2Y
qxI6vjP5SCr2w6rOkjMFRdyS2d678IradGVmgSWnMNglVH3uf/PtHuaJXSdpAuJoelwrdsE2IXyc
oY+aZFFrDVwmSsFZdpTCtBe7gF2Mwi4lAA++VVdri2UsWP6jX6rVhXGyLpojcWMrEDLkJqMU3q1T
zQtiZ/XeJRtgG8blyg7Qgv25RpRnFCH753hIjZXECAd+k2tfBG/EBn+n0/ZjrqZCrUHq91mLgv09
xAWR3kG48Yk0I9T8V4A5wCsLJUYlvccM+feJ+gHlUllxvSMO5fgK374m2fz1YZKdkW708ukpjWoV
yf1uk3KVCG1iYALvMIjtB/+wGcf5fD/xTjXRneABNuG1ZtTS1NesirmrJTgXTvrJjlLR2MUziq0T
DZLIs/IRmZ08FqF4Wba82z3vyYXy+/UnCmDyVN7Ktsx7cFzQjN/atTByL/pdEh83ZQ573qEWTF1t
5vga454lMBm7DS3FftI/yJVifWvZROzCEjrQu10jgnkD3bDYGBvTp5+ocgWFHDrG9J2SZHmN/Fgq
HM067uHKk+hbi/+ZqymuJua4TrdaGAPK4QhOxWu8QvfIHMZDP+qMrgDMzqTIBKfjKB2xt31mgfiX
pvJzQLvl8/M401cQNa55XbOrNi3cBiLE5OlDUcruXkYlHuAKrX9zlAU64KZ+dCxJwlYQS2M8aWxZ
UsTAIVeTv+oiWeBJsUvbzYOeHASblGte/lQh+CpePz4N2HPn2xVT1qWvkJ+1W+UO4Ri6c+O2Miuz
V6+GFzhzbLEFvmlBK149Hi/+pVFHHd3q9YF6w+Mb6s8aL0xb6BzoAVj9RB+ufaUv1CgyA2rO1Ufo
h9jbugPBCx5bihW3kvVDSqmHCh+h5LiTB9uhuncw/Wdo7lP9uxLuaXgzXaNhFE2BJxibu3od3hJM
6+ZtAx02D2VZCuNok+z39hmpBsZFuiTYT6SmjvuaiftGiUXQZdKANWRx6pP2xFR7b7HmI/vYsRTG
N80Qfm32IuHpCg5RUO6QCxoCFz4KXG6AK5JXYzp1VjoTbgMAqonpgmjY4Pa723Kh7Uq0PPDt27lI
fGx/IIIbrydXsASmo1jqgouxy8Sbv3QNasv5vQLMe0YT349JUqTkOQO5AIMR417UGScH1g/hDH/X
Nwz7tAgI6Wbosltsdyy38uYlyExz33gQf5yuiE0DnnR2GTCKTSqRgnvXmoubr6WZibkuaMRAjM2h
yJgaYBrnuJeMxNbC9zC2ZNtjXNjjx3QlelCPmY7rge/Ql/Zw51h7CYPkZjHwd8Yvew4zml169/x7
yqs9ynbEX/8lM2ah/TuIPOIcCjmQ5TS+HmvgoQGSMzyGncrMJ2WHea9dnjVgg9GAvhLMaH31Ukj7
damEV0PEtDEbOTu1sUUQK+HFctrQKlzkb4jWgEFASZcGcT8htXFrhSXEIL3fBUaIL7uk0SAFlvU3
hdkhRfq77FcNXvE596IUBdZwyPy6D2J8aykok9W4l0i5V56DJgVAYpxTsamoCaTqPpqKPZ554IdY
n2lIfVtkybQfqGn/cUtYpuYWw593FdcgMle2Yx9tJbmMO3OQlHqDDUunZfBuZVxcK7HR7J8y/la4
i9T+vVWr6Fdb2UGSG+FQbhEHk65v+kExDbHmTICBECIHbBbqMCcwRaC4sWFobwMpWPGyEIUxknLo
B+IH9QZRcfXDVYjuahISD1z7mXsGCO98cfTy0wbzZWkXdlk4YIEz8lpQELfGGKNGn1D1i+x3tzCe
y3sVDI6x36Rhnx3XrxoLykaMikko59CtfV7Mxml38EZ8rGZeuE8qctSssUafZTrURoBmIH/0HSFs
kCFD7zyPd6QEnikrkoRpiF6+2dDqbc8sNx8rWAc2jnr1sOz5XLUJvFF27LTMg+KQ0DlZeUKXymxJ
BrSBKP7Mn/x8wcVkFEq/YXrd1mMvkZzJjHfUsIsImlPmfDysl96jxzfedlP2NIvx1TEkzjtVOgeM
hBic+BeY3pujEYeSmrRwri4l9rfngwTUNipFslngaqLAJPwMBbdkoeXz8TYUTXRxzUZH8Hq1zuea
3H3WtysPCFhtl9W+hVBiPfaJpE6+BqNBc4+r8e/IvOOUuw5d6yXAHt18fZaRU3tJHsmX/4vtM+zH
6tCA/WDC05enGAxIKk7CjHG7ifL9An5xN5fjE1jRolow+y6c+yh2IXCtnRRmoGoRIWLcV5os/YIC
f1ewyYi3EpxvreX1C9NFBFrfA9hCAqmzqiOrFmlC9FA2LAiXGdBdEqeInTdOcPEMFulhD5zWAbNU
zi3C1cZXUP5/pUseYpxMIzT7ShUflUsLGNc9PR3VWfda734ag+fMfQG3hlGYduePmTuU5Sz4Jebg
UhbLZQeHGFb1E34wppk4QZRojjizwO9jFUeJvy/FMB/0tMytWjOT9adsX/QVH3fdaOrTI5AM9hir
roBayummzRr0EZddI3lYnZFRHJXi/ZCJKIB+UnaY3wXZN8fLt3i3JBk7iTcserPmdecV5RvbOCSF
kpy8+mmFe41XEca9kdMYxskW2zwgYtVWWd+IjJ/pDD1zJmuYCVoERDDoy+GlxnlyA0TLscodmdpH
+KGT577YGUSQBle5qeOZqq91gn9dbZVxwkwguB0Lq3vA7WcpHpXhDH25pxQpa3ifxjWLOLJN7rU3
sooSJFgK+FCmnx5Ec4jp8hvPs6EyxBKU4eC1TxLwiGs0qA+BeWw8rPwq1akYrIsDKzgJnzDWeixy
SjNFrUSJ5LwniP4LBOIerTeQmP+/Fq1rZvvg0mcHg2tT6msXF/RtY4B4dp2zPyHX0GyHjLTqJ2Ue
b+MlL9BQRNGQOTVVTrLqXtM9utPV2YbRh2oDTEtxtybgeWWtIvtAphB6vYGQmgkZ6gBLRyXGz9i3
GUwIbuJqZh0d98LoHb9zlwFghvYjhYKoVhPKVeMUoPKh42WLD+KZOBSZAanZTk2ceRA1kSsDxDQw
ewbGvCvfVpsqz+5R69JH5nLqSyB9Mkdr+rCw82YtgHwyGvERH05jc3V3zAxRP3sGv35VXZcNvJqt
oJVPMcVt2XnC5VM3G5pDkWGEGjeWlDFNcOJCMS2XIIyaHGsdYe7ulxVtn9u14nsEXCBsoNwQuPRz
3okXInNKqEzLzdR1XnMC2gNp3fGJVNzd73sgcCTupOeX4UQOGvXaq94CS/J7hk04RjVqXmcPMQMd
CE68LOO+9kBV67xvwB2BYkSBqLlzjXorF7Ame6OM3EMtZ1WVjZgt4zZ+8/AZVWzZrhto7oJBSsF4
ysCMBcrxXSrbfjZSBSHIViqVoKgi/DPjfuO5N3AZEMIWmp9+FKttQEWxFEo/sMZTCmYqPeuFvYkA
Fk7Mc6Azd3KIpJ9T2mw4DYrfwyFDPqj2fFAUmQ+xzASAcfzmqHG/tqxi2WsozU9fH7qPaF7G5Jsm
hulY5f1osk+ynkAROBIaJNqc8aGFpBW/JLT1SFWSOoGPmCxUUl7bYLd2VvA4cxlkrB3p4B+2mvLj
0UEVOZHeJRxbHPCuUKW8gL5+HiK8V3RQKlB5zyVblpSxYzAesNOT4KYMqtjJI0usNnZk3cVnxCzz
Dg2LTb3KI48UjA4QOQln5Mfm5dtDQN6vqZ0S1t9/mktEW6pFMwquyQmGZSXuV83//l3/hNJRxLZh
Na1uRQRdD8wsNQJz05Nwhfv0I1i92hYY16zL2VG2gpJJYa8GlWOG0X6m1e4YqfdsBFKaXcQa6fqj
6EvLwZk/drBbnxlH0XExRezRPD8qJ3R/ERvtwurvR8NjQYbf8fT7ze/iGc609BvaW/DVui+RE+9v
BsVj7rQOObks0bIviVoT/0Lro/u6uk8pcOZmLaXTXBABQy7DIF30az9oSyxXbTXGt8uBtlr9GRe1
cXu2NXXeyr0paLTdm2aZ064SlggCKPKj8eR6MUXZa4qRUlbj9eCU3KhQMomlBoy51hIy5ApfK2nn
l098eTUwA+TwNNviH7kuwgn1aqcEXFlzbY58dcKty0Q+yvNlLHcSRe8rWJgDsG0SHIKujtBOtCaX
SE4oDA4/49pKbS+hRzfp5rvXOkkOmLKyaAuoQzURGCQ14gsH5X5CFEVbaX3teHw0P923waIva0M8
KHaV5AI78rT5aXXLSKJ2mAH8PQjPRaFwLAHd2nZ6AFSldZ68boqzl0U+szPXsRZ60nVpPHerfz2v
K6pGu1N/U/8mjPniz05M4OT6rDiLl/ZroCU9Yatfxs/ej9nZhNWj/HCXGdU47mrg/Wa437/EmPSt
lNvb/zLofEQfxtZTlafaOHviE+V2mF4VZfuczkNZ70dT5FEAZQ4mYzQnjl2Cz+MvCa4ZIU72goR4
mVXclkNxGlKXnfjWl6/sdQ3X6/jQLJqOw8C7K2RBho0/O1OjO5nDqkzTGzbNtfMKCj1KXiJz01Nj
CQPWa6WKjMRttZFXke3zUf6XaE8W7fWYCR6/UZ6EWPl5ky8BdxEre4A7hi5jiSFfwTbc3BScnoSA
z+wnyT55XBJweLOioYtesQ8ex5dZxGcClc8HeQFWJZ/LJ19t0doe7gBb/UqRWZlMlMeKZycPwuS7
dPXaMWZke5jFuPJvLQpY3nIK8Oc13gN9qnkby9L6XlshEVQ8ULiVFFrzntI2lbjvDy1KFpWDM4S5
jViB0s0Wlq9nhcrI07gBD4eahOGAH/0ZHB+1TG8HoT7oVjLoRpXbYwGS1xF6aW9dl0Ny8CKW7KNz
i7i/GaS5JzEDpBA9/ZtcR+dvhYb2ScL6UsMvglG3wp5oJWzsFEwsomcNRHKo8sXDG6npuz3ANMQo
XFDHNYtfT7lDrNQ5oWaFFhI80iiSAKQ9mUDpmk3r7WyKubXnjqVDNL7XUTu0IoZp1+JKe2SCs1pX
Mwvq//GWoKIUhuZLtQh3jJtNMwD3P+g+QXcNgXrbbLWugs+Os0VlyafXU5xm+5R3nxWkbyQoixgw
kDcLc8AYXfBFkC1Fa7+FJ6De0X2uL8Thq7WqkwtwWRP2DDsCRbzLakxJqsL7f4Dcnj7sfIJq+0Lo
ohM+KxszhXSi4XxwUbbQqzNiciVgz3awNKS2yLfAmWGLdeVYpfe6rD1FEjckMIS2vM6Z8Zyg3tsz
FyyCayajaZiNrJ2iS4DkgpnqQXyi2KELIrqMDBe80ZqrFlDRTlmXeKVFA3icoD0a4w5BlE+37xuM
3tlm199QKig/KLezW1kHao+BT933HHCKpr1U5cE6bUCkyNIoH8lu6wSb4GE5dl/ekCIQkB8KFSTj
OR1xzrmZORpjTi46NEtWBOP3Dsokma5Y9IbFLpUrh7+bNphWtwXKifBkjuoUAc5uSeIallf/YcKc
ZHBLT1sDsxORdDZnyrdSnla4hVxbxMP4eM/KhvV41yV2In2OB26V57AGEfTUtvfZqa5imEPm0SyB
hTj+7MdgI21G+aaRZGf0vcb4KMKo4VbEwe3kmJ4dG9tq8djGYBEywTKl0NBDJyzQNoveuRASccyI
lIJkRkdmOzGb8pHMsldF00VY145V1FM9YnB+ywTk6O4sDMUptPI6U0FdVd0XnF/Z93jJ/T8yFZUs
pz7tv6KRbSZJNZGxFJkwIN4erf8pKQ+Exu2/o/i00g3ghqWe/0efJPL3Obw1pu3ZHJHoLgq0FZ8P
jXypuWm+Aj1ZsrUTuxID7bmAA+zjtlaLF7zQSb3XGqG/sfSxiIqldbknLiPpj4TKoDaojx1yVGfR
T1SxHF2Ir2qn/wN7MNazflQLWvgF1Jw1C+tjwCwAoz3Z19fN5lJ+qDJxJvIOVTvsEGQnU6vgSez8
qsB8Q9kJPmzxfl4kySW8lrM65GOPi5kOt1/ZNda9G9mC3pL/RNcjs2B5bxYa/NouoMrw6dYWMtqF
mILIXM/h065+YDoBQs2RSJlV1BR4fvmUy5Ik9V03UZRo/mKzZSmhlHotDE1+1UtTVIVQ9HdrvFZC
sARPKQDzWTJv7ZceUyz1YwP063CfZLnYURsm3HJZa2EvldYto49lG1Qd8QCdunxG5EPjdGDYFz4P
3UeuN+hLUob4L0l66FYXt6Pui87bcIx6/iJU5Ykn+zpEa3sNftfp8QDLjX+4MWyLh3b7Sfn+VkQU
c/P6OSk9PXrgU4BQlI9Ai/Zh2rj9CvvOabaeYqA/uV+b+qY7yQ2GU55lhvxU1MCO4dAal0Hlln4Q
OfedCww5YRFijL1hm9VZADELdzDVYo/tdB5GPXHhOjr8dT8tUOU6QL4/4XxCP7bb9IIL2T8aRKyu
ODWjV0ZtdKfNkQG8hPAgv036z2xlkd/VxuaZqP6smHfASOXuIuoPNvy5RntcOTU6edXpfkG5hn71
eNupHjdymuA4cO8xMrck0JU9yqo5eChxJ7IPF0xWUtCmVmLG18LFooyV/bP76tGGN8dfMQkrr3uw
BbiVupIjIDMNFIPREMM79hHaYXg9wEAoeBoySRVzahYDNv3/vFWFZhe9MTaFobdn3///kJiMCeUr
NkCk++fEqWjPysvTEtfcekdDyqvw4zK/yS7gz8yFqIp9iAbaS9AYTsZXhOY55l8WkSHhAWurz0k8
/kk/fssLRFVBMCOfJbtFj1W0tWi4wgTP78FcjbFvo6eXZo/e5HVzBFOTk+d03UdHO/LZAg/C6etn
jDqnXrJJzBPyt20jFmOiPdieplDb9icLmyoRpq6DLtBuUblQqmBj84S8x01JgM8ViLAUXWwJ8KXy
BwpbW5NGwBRGzx1Ealta0MYXtWN6PFpV8rIGtPA/1wDs+cAKMcW+v/UL8g9MsdkkNO79wTmGyimH
sOn0ndbQikj0QdtiD1D2qJ1KpNk3oa/e8RyeOe2ENHKGbtWheH+V/ClTysCD6uVKXyQCizia/AwC
gt3M0Z2yt/3CoAEts1xZmwrN44PnNfM2bdd620Rr7SDeN28ZtLSRbz365jibPt4Bym/MHa814rbi
rZOicQ0a76Toymx0jcviYlp3vdBElEJD1r3CBsHbiZ+bHcTni3h2NN4Ua55zXfi6ju9Xm0W7mkl+
XeLxJed2AQDWKoqNp5p+jLdw2e55QOveEDJRYD5lAf7fTTs1Bp2UjF+nBLwY4HLh9OydgaLaSkGv
+GCiEs3buJ7UgSNJev8gIDfU7qaKLoY/X9p/vZNCYRcdYZDglTcU16CFVqSrN9gQOmn/oydAiGPv
tkadnslqqSQsnBEdK9X0gXUkyfDdnFzeBvtuHLoeMHVl4GuEd4Hdl7vOzZUnEAHpd9ZAAD5Tjk5L
twEj9oN+JNanGwfOfuAy9fmhqcNjLRteaDYou8EzpI9boqgCZXP+wJPv2CFVn7huTSlaT89zUQDa
W3D0SR6NYg8G+A110rCQQ7RcViN4MMXUPIztP6gCc/sHVCEPWe1x/XU4g3GxISpPZLLfDtLCPQHj
L6p3WcSrBZSzv4rBjZ394Uojp63/SjN9T99E+3gYIw3mQnKTyWOPFwV0XUfLASCN7jskom8XNUG6
L7xDk8ACNwPGu3FgZeX10CnwSKvChH1XQcME27jYNav4zEsJR6AkxxhMDEIqbI84PVgtnu+wko/a
VNQn/vLwGepI19BH/qJ6v5Lpy78EIRLamLlavUINXPStMKMEREXBRO88yaNCygR50VJahXxfGZLp
tGupi/eBxmav8/AoAdxg14fyEKu/eCNEZ3App9zgeUjPlA1xR2dcfVRJ5ZhdmKZn6lPNqygUjic3
RPIs3jyoTybeU7bDfJbZR1cBGssDQYmryhfhXMb0APfPX8mN5bXoqOQ2vyFt/aaERZODucz+uBf6
ugESIbusInkJgYMhAaWng8WVqM3RSa0CIkzhlBvLhFmXCi3JEdJ8oU9q5VtJg1YtGnqiP2SPHRWV
hc/k/5TPgmG9r0ti7mcy421eFv/9dXImwg9I4zim4hHQdw4aSdBiFzIzY7Nt97d0q/6ic9thy8kv
91RMNBNnYLJHXqooEb8VQwF8NcxWZ9BIjju1KsP17/AN+ugGpGr+3E8+szlt4snAC1jJpSEETpUY
mFiIC7LoVheVV/RRBLJ4eumzCwRwDuq9kPEFGfpQJE6OAlyTqkn+QzLW3BbITp1C8PwYWPcoEfNZ
swXeDxwjKboAk/B5xgDSbAP4yCLnbAiVA7tq+Aptibw3/pWkvG5Yz6vc1VDhbqBRhuhtoiVIhJ6A
73XBsJ5d4J1xX1jH50hOGTnYMkzVJbXGPZPq0xZxSfC6IIde+o3WGAQwge/v0tUk8kt3u7n5XZb0
SRPsLp2OJoPMPwG8aYU5BvEWFzwBxlDya7EClD17M/9ic3nJ5TnztAbrRcrjmVcN3gZABgqjeOYe
4kiPPRW4mjsKHiRYXmqfuy8c6/oDqWEn4sJPFtXF7iXcUJbiG8SBrh73uferm9dp0PHozCOv4qkq
Y81UfM23Alm2fDY0PS6aJdJpVyTXbjnbYSrk71Ufhv3urUal2RAr80ow7yDK0KWShu7Or9t4xpP3
SueENuN12CavMRZp8OaeNqV99y1VKKcNmHmpMtRFXZ6spshAsamQfC9TlkfvZnlwQ58/68TBgRsO
IDrgLcC4nSGxa65Ptno/tjxnIO2l6EPafmK7EKK67WVXvU9eISRGTNwevUt9Ot7uih/+zhBlRqun
NvHB8d2/KI0brfhTQMsLuCzeNly4w/ywFkk/lxfVcrGIyfjq9H+YK/6JZf+mATR2EVH2x+qelHdJ
guT3bPcjXjwHVqpEysSpgoITtYp8rh9gE26n4H7Jif3CGndXoFCU6lsVpR1RRKWk8ncGcFQrhSP/
6Pdl/53aVFalPooweYj+FYAXyCeGTpqXSBmnOLnlH1aiRvI/YB/hZxKjdFEiPGM44BF6VsG+5/l2
GHJ4viY3cH46JrPMggFpaDdxhHRs//IIzIDGCaSBXXBD5hB65h4j5q4xy9zFGWdKuBGiz5DncCp6
5xH/vm/Kpw9b0O78TME0KBFdlWQ78nmL7FuKrvS1vTUB5dNB9k6Izt4hw/EDTO8mGOxzOlyrChrX
AuqrcwuIn7NYI2F504gN2ZyGk89+q6bc2s4gRh/mpC687DZhxCx9qogWPIxCqti0GJhsN1aLuxgb
paJoXdsKb/ab1fzUjHPrlD3HM224VnBeiKdZl4KoPeqpPYD35c6YyMa9IuqllCY59o1q0kBJkEh5
UIZF0LXyEwdrJV5P+27hCsdkaYC/85rDD3ofXUwHr99B+d5+I//CpMf97lDXjeG0Rih/bXumxtdk
1IF3F6ILlG5a6rJLmbA2HL/iYBL7J6cu3kyqTcxLR8YZ8r8MxvrQ3zZdONNyiel3eoOm+71KPCLh
T2eBzgSTwNEAkSooabFfVAt+ESHaCDt5VPV49O7b2iR1B0CMD4wMsg2UNxJ9EnMMQ+gERrjcwv+O
F/uWqi/LZ5YrbmHPq6Bj4CtwgI02kYP3UDm03z69Qn9gdD+iag/Y7fFgKeHWPhc0mtmp6Mn73RIP
Fyiqh8wcFm6mX4OJ8W/V1qKGFNpO+Xv2/bjopsAHF4NSHINLzxaOHTmpy0UMzGj3sGFB1lrOxuwE
LJobzmuFI06VaZuEEMbQo3WSDgxeFyV9AJnPnxAdRyJj8jpfpD+2b7TyAOyCGZAJ5st8f0G2B3X+
P5EfZ2k6lIYOP40Af0ONQXJIljy62lNKMlZIwlvNeWbiJ2xY72SbRHHURva4gMqbc9prQn1LjDO2
stGkX5dwrGn3Fcm1EC/VMMRZJ1urlJu3kuzg+WXGAv/9uAH4kViSgT9KKvcTewzcUu4VG4qbti+V
UNOpSK7SnHphvnxJQ2oW5fy5aUpbYLlqENiCzQi5zlbmXJRVmFDza3rpVzzxPOsuXN7eTm7Cslqr
k3JZMosXsQvXElZB0xdfy1M81vYQ72wJJYFgkTpOtWt+Tkw4mrxy2S1VmPBzJmHQAaacvr09c0qe
vhQSJqtnT5wDDxU7xka+zuYAYs4Wv6EMaky+5yj8+h3PSpPwRfCAnvgW9AI9OZWnKWB0ifgO+1OA
yVAlgpn95PFCl34X1gwY1PIBuI9OkDqd04pJfY+ZdeD6drzJNb9Cxgj/9hvNV52Nzl2LH63jnuTm
XCy7xzCsjYgIz+63m8hrGSAr7vMCnuztC4/EYeiQl7vC0B2E7vgeZXkr6V6iLinL2fFxcgTUHQH1
OwexyLMrCzn4hK2v6hx8MhXP1FbWfcMwRWqfBHJy9ZzPwCBA91+3sllQtbYaoRGd/GYR6EwQQTGt
NdIzl5cjjuJyv3NmARbI/pQwoCzwJg8PCYL1nIjHdl5KcF97Lv5HA4xd21dGxfhTNkhONWV3Jk9A
pRDO5U2xj9pxcsTh4KRc4EBjmUarnAKvTArWUOUI2ouYeo1TzpT+WjhnvAF0W4IvxIA1spo+TVty
dokiB4qnGk/m4KB2qwsRB0QOWr/UZFlivBsLPBG6pnE+PB6MAQuFGtsQuQWjJigoqfqgYnSgTXTt
eP97SOkxGh4uNqKNyBnapo4TJCnsjIzwqG1FFUidF/hjLM48THs2F+Z0nwkTcquNv/X5k7Evm7fE
AuoHLysVImov0MR6y9rZx32WDgPm67Q6X8TbWWLtZxAb+Wof18ZEPNeAXqRiz59H2jx0fhHaLU9U
s5KeaoZPpwvkxNlRG56bwchdivP3Qbb2Ek5RB07lVqHZUdIHgEXwSY9HW3ZU0RzA1Efa7EIIU+EP
bNFq6Z0hegfUOEFJG9pLID4zR7EIBLM0njuB7sj/MNHxUGasy8CA167oBsCjW09iTIwLKZJB+71H
+A3to6eGhZWu/3fB+LZYn6tUYGw5er5YKHOWewpmgRiqR+vQIBMGUokLJqpv8WEn9cOZCAT4rnpz
NhbQmbyA/+C+zMugHZYSwyZTe3zK9OSnARv2N0SQvdOOZ9sbqoVh/tvgBfovPp70HF5iMwMf2TwN
x+7Zhi+Eeuk1uIbHjIcmHTGE56i/hfPr356w8x+NnzjAEblMFjUF3FfKYL0ePHZZQJjfJ1Uz8lHA
tAHxlVcaTIRTFPQrFbNeK8A3bFr+c9rMey9kUINkmBPHKWFIsZjr3oXRSEik7zi9MSQbM/LLZPOr
qTWsawxKRzXD4wfu5C/z+hw3Vf4cj6iDhyHaHr60p3q7cRnPR+LX0CvKFdpSrKhrRgFtP5gX3Fu8
7nRtXPO3TAIt7Nk1aedgS/JJ9dFISvQlBgk7vEqOcKnmW7jPhiN01QuDQaPYRomkGu4qVOoSwQAN
BELy2RngZFXfGCaCSfBa//9qoO2dRfpKsb0DrC8BRTzAswwGorWDoB+NZMqExjl8/cTSWudcv3pA
DRdmNHumrhoXTZLXknjYqg6qhJA121DKefB8sx9twzCbQ0H5DAcwfPi0zUMsKwI9sm4U8EtBWo/4
/nHt/8wWcs7IqZauvrqplQuNZnmFGSRyflmp4FaSrc+D95Vflh1j+sJsKv5ffWypFlXzyEwXxREg
V2O4G1CUBniBkGhE4Lc8IVsvwEXmYvQWqaq6H6N3i0K9N01bSqdxGE0nV/edjIV8F4asyivm+aap
mtcQ0mp9fHF7P8QSoIDU+pRDm4g4sKjUKcidyXf27gCh7EWnuvgKBTzlXwK7BJXjcDQ7TB3azhre
RqOx09mk4yTgjqlUDs+V99Iw6DO2k3fXaW0GCO8ks67akId/a4Ku9Yqap5X6C3EOzaki4TMkndpU
8MrgYKd8epQRtFXbpBeSBV7wHqVJG96ExrQlPFbRvxxEZzD7iV/ZYwTjtn2GTOwwfZEOdhB1w62l
5+Z39ZNQqfDOxMjMtDnXV3GeZz1Xbm3igquxcKcrl6cm6SBQ13e068RFjnTiFaYvbILCEymiXo/+
UXTzbm2RMZWeTP4Kuo+L2nHxoepfodfAGowiAEtmaJNetL2gBJs++hnWKdhE6Iz8bDLZnV25qw2T
pABO6VFQ53QIBM24T8qLKuCwjbuO5F8qsh1ybKoszDR4QnHon89TGLsYJXD3OLKHB/X0nRBuIAfE
IcCmeZiRKwxJLr6ufoV99iHfOSM+ZtWLbWOURdliTp9UT5S4bpH729MhxS1k47rARh/xYLWc6hl6
Fxyif+bnRAOvt0lQ6VKlGiP6OIbHhIDusFeJDxX5UVWg9Y0YhnCuPr88RGAOD+56MKKiPeL5nTNX
2Mt4+LKOMIUNJrIzileMBTbo7RmHnvkJm7/6oMP2cDC0eqjqUq/SiPOOES4/QCNobz5W3F9rREcV
/qQCRSyrVrqbtPMiSUsXwxKqpElM1JOqCFPguLJ5mlIxb3FD7KS7LFx8swhN5IcXgo7WzooElFvV
FT2Pvr4BbOEVeaCA4VftLOR1sIA5WOAt1uAIQlQErNZviW2HlZPTszFiT8veA1i9SbK8QXK2/DYi
OON3xz2137e7QiBse9O6ocJ/yNWxG//gW7eHhnApWGTJAkspYRlN09H2FJp03AsytI0UyDZPopRz
s4zwr3JbMYu8Bxk3bpD3UM9s+LyZZucQH3qyPUquwII5gEaUqZQwSDjp6jV8LRBoV36hLpWB6y1u
uefsonBggffNU8L/2NUtUgguKw8Hv+vhY3w09heRS7qP4jTIzd7gnX0hNZM+LnFuYgQjcDIi2hqM
vR1uYZOINrF1+LL4ssWxh5m3SYgW7K8L1P0U+KOmIUhSqYjAnioYUE6oy2LuPFdBJok8TiJQ1p94
4Jsqxh0WQrraoMXKz9+dsJ5GgR3P9PcgTdJ6gPkAVeAn7CqtsKbAEiSXq6j6JO2UHwsBHJei1gj/
eu7bELUsL/knSM4LesUbQi8is5AJaDyhujxMfFeuYOKo2IGXmwYjpFuPaYqO+VDOiLTtTE8YJE5Q
QmSqD2QgT59cwsQRonl3u+2e1KiMatG1RoARp/CcfbggKZGWL3GCHVx/6NRyneOM23YWJ3Gal0FL
LBXJea2ltd9DvM/WPOwlc3LGXoT/beIwLLKR/S9Agfw0nn+P5Ko9sXbML1VO4IBI7zDiiHdR4edg
LGylRwwkbaNxlYMF1BYKnNdedp6JQWrhTFqPiI4svb6Ng9zlsO8rUwcS2yriXC09K/dadeXb/Vfl
0VrTWe/+H8MlxEXoKx2WVNMQSUfDCfKHEK9WZifRqD/8NsPDzZuT+pmDAYEwDTIGLdfEiaWo2NTB
Xo+sLRn9AT4Z+BCpTCEwm06WXk2lVW5JErSJAltAk1ZhUAra0Lxw6WgMHk9Dtk25U4riUc9qU37D
RyH4c+XolGuM/7HGDqhm5826mKNocjaen38E5aeHaCR+72FOQOborXGCgJVS4lzf6ue8z5OacGYQ
pN3STya+RBwafG0Zzw4k7q/NWkOZLDh24xRG3NV63xUQcQwkVBzBc8O5o1C1zidXir6fsDD0bRsd
wbCqKpJcAi8TK/jdqzN6me7v/vhVRxDjJ2uxgYvm3tuabDhDzaXpUDRnvAWM6n52VgDC5drA2YCi
FuOr67zZc9iOIhq9qFPxC6njuw3/sod/45nfhhjljlhEIqfsdy3CMWN2ED4zx/srw9iRGew0hXXT
i6KSAhr3lA9cSzULK8FgmlXeBuRbhGq4KouHkE7rfI0xGUcPN1jpQmqo1n8UVPdxCS69FkOefqtP
KwmCnY/exqYDyRZhOAB+17+OcxDFDuf0tCgb2TdIFsS37S0N/jI1+EtDrYuYlavUf+UeTMv01a5q
t/9C+GgJB8m0WyNTfW8lrjlsK+Ju2dPI3FOZs8mdwtKiAyCU0ZvxrdvNUyyUAIdwPZErQ7Y1N9dy
nEqdLTosuokmvB0nY1//Rl87vCQ2hpipXCFR5CwhmWlPYWYxuHiqBMegGRUlQQ0s4pPSqFfJfl/6
SBN95HQZOlahFqRmWkTioux9W36586r2ANHYQuhQMH3RY+H0jV6yUJihvJx6v4frmRZu8nG2pWXa
+nFu72AGZ3iNWbqBmB6Vg60edRcfTpk73wJS34Wk2kd8v21ZzLHlcazMlWAZmHKTT1RWTJj/3RKe
hkFfBjwkvxRz8n/X1IJnXHr9e7HrZjhEXGDPSegVHyzLLcTZ6ZoXPi3mmr8UfD2bPNS4C9Or0vzL
czteR3tdOCZk1E/rp0l8iONlgW7Qo8XLKlZFN7RKeMlltqZ91Di63NDsJzo7GOY890BytLyfmsB1
HlYarbkgJY7Y+30FBlweqyOiRz6IzUyhOlPkc+DUrg+Eeo6RW1rFGcWICRY5+Uh9+nwRw3BCsKCi
13GZ0n2AqZXYus41R1aUMdpGqkLeUrQDm+xzZzMAAKKb3WrTU8xtLseinGOmY0SDdGS0pNvis1S+
3BTM7Xz2z2pkaiS5zdyx/TUh6FAW3mC9SHBo3HKT1LZTknUq2E/5EZfcyWQei3Dziw2z8BZ22w9q
HoSX6I56woLZq15adhrrOaEh93axpk495TJBg6eQ6YWQQfHDmM3wzth0Var+NeSl4j14ajyCJ7Mo
jaGnQAg/swvMtKtfry0eeV66MOfZgKf2EO/6itcdT0XKVtAogtXY936133yhF8dLPWujfppJJkgE
jFlmAWBn5/e+A7oATVeWG6CWlTbBLJaKRv4pUrWE/NyZ/AJ0jwVlP9oQ82WegTSHUjkz8hpHR1Ml
pXxAFnmf4kcVKbe7mCJ+Pc+tciB5bO2CNf9miIKEEeSDlxJOp+KM3+uUMhz5f69QJJRG6bGbrJ1i
/oFHqOFsn/Is0qGYkPoSnxg0j/PATg6RQJNaojGlFgkgvC8+WU2InWSegXwRunOqVFX8v1MORrC/
QtA4T5l+n8hTzw9YqLRjmAydyxFF5pmYt4PIlIYGMaIY7l/GXP1nMMeDaxGtImkb1Lvat4jezDrr
hxFP8joDes/ecTn9s+RPmOALskTr0Gy7uVDG4TNNB6A2EMabvRuWs5wfnBnnLtCL3/KII4gPb4VS
OuIt/9PxjD1WNA3Gv3DGp+OpZsPbdc3Xro88PHm6rC64e6gIz3VSYhuBErKmsznSIS1FSvunYMUX
4zz0KBnA2dvqC5derirsTb0F2L7fPtrGObZRLfBxoLiHcTKBOajmEd59Actd48EoFFej76ASjwn+
PBDTF7o9xREKuKhwPKi6MGTFzSjm8GyslpGuVABI9cBy2irzAaISTI5E4VncS39diHcuXN4sC4A9
kB7X7sA1NHVkkzp8brueu9qnpqJsof5nFbF1SjWC37eYjXaPJoM0lJImf0qEeOW4pjYWwCCQ/Q4R
79CE2cMYgJRgXF3gPaPSmp1kngNnEZQqXuQuaQ/TOpDdYIC/6QTTnaRNIE3fCtV8Pj8ZyvjTEmbY
ETnO06F6ikvCMQMGOOoStDpvAcQo8zWtTllxqMcaPp2ybMMXzLBaOwKLTiZfoq1e/2Yo4ag+Rw9b
noPepW1peRpRn8LKpfPdnD+yHWwNcssaM8hI4BhXSiRInNcz0zX58nID9jI+hYn70EvFJsXUDKZU
NoUN4UD5tN7mdB92Y5WvxQ/ESRE2K9j/M33x9qe+K7h1QAEK8E8f9B2l0+x56QKGYrL2Jhz2Qruy
voXSBzg2UKST/Q8CQ0gGt9Ivt1nT/HRU0woklx/HChoYBd11ZrTF113wOYwBLJPQoFm3+8HFXthS
3Q2G+/yBv0pdReZXaTqXUHE7Ouo1HNXu62ewXWWllDEr7dnRyXvntGDbtlcCP3J0RQjaFoFSVWmM
gQwXn4ruZPjJs4vZVvl5OBcVPS9FY7f3bEXWuZD+evMZdCm463ZcDuXXdGUff25p4yd/q7EIVFOy
mLhg2qygI/uKMv/DK60+8rUNEDdcGicXUV9pCAqcpQ6jP8ejsrhi4ya7LeVQ57UpsU/uJd79c5Va
qq1nPzIcTkMOgxphMG25k2Vzh0bcZhViVcdxDKAYEibVzB5juMv5fOQy75f8nGGi67Manh16T9QY
5vp9pzJhtH6wNnqI/MLoRIZ9pPDk8iXrmd/ggymsbKxRXtot2v7CoIt6EU6PX4SkkTtAVvl3KaGQ
S+gtDeoPu2bBvrBnma7bAtIwWdQpgykzpg0gh1Tzi8sr8bZyNo0muHs59eE6cObA35Ib5bu/rtcR
jJV8DdVHsEntz6M9t7Y8QUmuxhMwG7bRv4yNXoVw/cWr/NJJRPArpYt+uh5h/HgQ5HCgCGNMMvWt
jcwJL+X3b16kV/mUe73aUJpildPPTANcSCBn5Ey2xgL27SwcWPiCG8Q7O8aVywul8+pO4jwGLcz+
ybzQ8+x5bA7exhB+7NdH8bd/BbiMbZb09/tSymQp3tZxsrI4uZJ0myCXxUY1qyMmh+S6Q4BOXSCT
VgMyGo5wkCCiIg2bkk/QLfmr1HzFtaZ4I0bupG0ki5oqreN/YX96mI903h+PXCoqvpnknebqNvug
PdGzz4zsGQtVrcjYlcZ6iUjUaWCe2KHSeCjl6tLpCv1UugRBc3MbjwiZ9x6TQDwg4is+LsOcfz9d
tkoS5RwdJomM4k0JKIPB359FzPhmOEEeNHtp5KDqa5tJTqvwUAqf5Y30dhZAerh1sW0y5DflTgXm
cUAwYWFIcHhTX0g5UW9YsUW5CsApMigpPInbwiVOd9GCpScuxAvkZTLeIEa5LzaDEFnu1oNcXSDV
ELk6YGUrHgllkE3jQzA9U+gP2juQfAGYL2FEsaiIWL0tHraxHZ3u1i3YzX6ehzz6obTOvh6Q6NbG
iwD/I5HdLGdzN0EAZ0ghwyYJogY0/0RLX7SV288OPEU8XRb99jANBZgdQFsEIlcsVe9gAc6dDRdb
x2lqZ5nmdvOfyWTsZtmDad4boLmnELFJnGyoeeY9+xqmiU57fIRqzO5KDuOsS6qhHU42liR1rN0E
cmj6rGm8syTOIXUu2zH/YZRisSqMlXiw5SIuLKFzuKjVhYRNvP2eW6dIroqmpjvOW7QN+AYE0Yhy
a4kFCnysPJMIyWVjd84PGeMZ7AauTmn2XL/hQZjNyx/r8vxh1GNEeQzBJHeg9hzeL1lCG60f53N+
yWUt4Wsf1bYxlolspJpyGvRmhjRqvu4M2JsmvjzwcisZD6kgbbH6tbWWgzQ/ztbFq8eNFplIX8FQ
K7wjdFL4NXWLiM/FqS3quyAK1rHw3TvVDhd/Mdiy8qXjEfFNO+ApmujEghlmw+NY+cpAFOb2NAV3
4Tndcm7tcOzZ0qSAfMeAuUiVn5IdYdIOz/UbBypvwUg/66PVrUlqOudBaVyX1RTfrAQc354XNPeR
liTwnVqaGoC654i12+j614p0iXX3fdPbJVI43rMtok7Af+qfq4JLJxzaWWEsxcR096g7Y3n4/x0L
ebc8W3/RzwYt714CHoYfH8eYe4fjZgjuOsS9CAvtCgRM5cV7SmFlkoEasEwSbxPcQBMKsSIkkYEc
dH6z/WyrNE8OWRiM6MnyFx4EHbkFU+85e692+Ffmmnfp1e7LPCspROIyBCUEGOvl5XiL+csv3Bgd
1kEc2jFvH5GKjqgl76akfvIfqzLlUktOWvk35JDDxqgzLorRZ4tHiW5jFXtXoqEsEmYudyUquK1r
N7I4WsWacgG91UWq3zPyFj3kcHRYdX0Mwpss/oh4ke34WoVY+pdfNzh46NoFPnRLigGZwrqPHpfJ
FRxLnnz4vS01hcOnvyXjpoNox9ye+PW/GADB9afAKxyqVd5K57F7q8rPeTLBaIzzrIg6b8uwg4cJ
01jDrZznaFbcijKWGTwOJy+rBFMSu0sMi8qI/9WWxPwyRNEajXasCXTBYEgae3LHSWlEVZPhX8lk
eIoluMCQ4xxvYcmC8Kybt585nffgvHQqthyYtJUaKfaJUtDFZzvmOY/fe3zwrZU68VbPnapuTSfX
rj2GVA4NIwg3KG/7xhv8gllUF6m4zQ/p7eM+UaPn52r/qx3QP57tzxOI4osqIRwi1D/LXY76TIae
i/S4LLC6kt+1sCjAHshndiS9+B5MG9W1+1Lt2l8oceqFk0ktole48bfXsC8/RZXcVoBCnl5EkkeE
edad4sCQuh2y5CXCnnikHOA7aKUf1pPUecpvLOpue8W/XBBXidO1AZ2GV/CA5IuP2yVeVOEaNs9e
gYOZX4HUBWPE7JEmghIJjkCJoKoYN8IkuO9lhyxzZSouCyhHJXH1XVdT0Hhu1U5E6Rh8sjqak+ZZ
9+rp4MXm1CavDyGw9xCoZEdajUgnxhh1GyyMLMpIK+/rWWdMxOHPTXE4hfHl7FjgFPh92/QxLeNg
z/NDfYW/9cNRX0e8t2U2MfyRs/rIHur1lXHcA9akKmb3sFBw/1m0HywPiY0JLxY5tq0BPnO+w+va
tqQCYpat8Rv7KffISbyTJFCbrM4gnNzYvW5uSztGtFTeJUnmhk5ky+IqnPrrpsIif1O9dIX67940
pxQ7rXBz4/ng/XtEkCa29ZwjXPwLbmbBDxxyyYMzmxKwEeuqL8CV+I9vkdabA4YCABpjAkVwhhyW
BXa3rfgxc0LcQtJIQFgRubqVWwX+H6wxG3e9V46tUOpR1BtARN4gU+x+PJmJpKZQSxowzDXspV7H
4eH9Q4/86JKDqzgJQz9CLMD6s2XUUMPsC/iAvClZY2KfiFB8I8zPyFhWhR7CNogGzwHwPKab4gJj
3ALl0bflUTyW+cCOUrh6SO9KO10PqEVqteVR9oWc+3tTjCjGkvJmIW0pdgDuA10D8Ly7kC72vruM
mBRg149JyKKFxs1S9JxrJeAaoAbkYvbEQNSM91gyqOOCa8/TpGAxuwYVGLdqEi4tus2w0TPJZAnI
5nup4tGdYT91rjBEAOgUHriiPne7wY8PUr7e2voaTs8PgTqoksJhyMHL7uDH6qmm5vzSi+pZvdht
H5W42DyjaYlVGbFLFBNPq101+D5GWTvlC9Wck40B21RfUbgt3XLFxcaDxGpqzM8y+5QKnyOiBT1D
hP+v353bPnVLC+MF8xDrFzk/bQmxQNUlLh2z6SDBDMwTfYJIRbgBA4fQn5wh8zd1Kkd4I4HbhCt8
RxoSHL6PzktWWjvWydRYkbAjM4cUF8DIgqkRnqylGQOvmwIF+rzqVADVvkjgqRs81YCrTff2YYbf
524MT6ult+A0qoxcd3JcfcVB+pwjJM6rgJVorJY6OYsCbd0ZgyfwrfGMQ31ulYfdhsd2lmDiQXTO
+SpxBhsApfH8hIQiRgF5qSNW6X8VkujCsq82TApJIfl1ZVanPA67XOvLn3E1c7rOhXwGrbzwfx0g
Bxjw8DOp9cilpMsqyzYoTBQU1cDwkgPKwbfb97YPsehNKrApNRQXUxDE7e4M3dUbBBoFNfF0j3is
7ytAuWfaJz398y31Pf77GablqYNWbIo4t3Kf6F8zaWzekUvGroqIlq2wdNnJnM5pvZCWhInGtJVl
JdV+5LU3n8mYOCOIfEiFDjqIFX+dDBvsS3ik4yMww5OwwA3i0NFCnl7ikCX5dzrmGuPgFmczcqF6
ii7ZThnpRSQAmeB/DAY3+WXb/vpibpLKgAEEcQ6YvS0YU9sB4LqzmUE/U/znisQbSM1sON5Vwgaa
+X57+qF5T9aQvMby1CtN4nBVPiDW5WOB8YiP9dyTDaOCfVZnLacw1R95rwmkz+bvcBd/VQcGKyA5
/fdUDO90u1pAmOp//5IwkISNWpXdjUf3ATopcq/pQCKMmABwd+Ig368u6+rC+ShVDykHzkws9lN3
vjisOQPuDnt6nLP/Wae+9MIDCxZm0ogFqSwgkU09e/BMjQ17WsJV+/5gLeO2KWi++nDYVNFKqEUU
pYxc2vVUe6gyOvOPD34ZjVwYZ757xPxsJ/ecCcCYuGGLctQYUdwg4pSCoJpGXcHNPUBwMRiiIyqO
fLnwWNazZ2WcMUJUhzytNl6vJGzlAduvI+uGfn4AL6JBhC+H0906PHAOTjUYgKQCK3iQ4g5nlQpg
ac5cGj7jRw7NjaXULzlfaASx4EMHyv7u8doHaJTzFuoeCXqR/K4YurPDibKrduqXe691rTbMRMcH
w5DhAtGTEEaT4JFOGofi/l5oCsrvMSeosfQhcz65QeGqTYKXgxIALZPF7YUaJ29ZbdWP24voV2Gt
Spmdb6JfNOMHv7qpG3nt+r+gZJnFjWO9INwbe159GBJ7TfiWVBCbIyk8FT10D4nX1njIbgDCJFDR
806lVaR9u+ARR0DnODh85VawOrwI1kt9DK1s/Na7aKE9lJk1vhJAMP9Us04aGJyNmtJ6yo+jCBc7
RGrnhsgY3flcfIrhCRkHWbq4VvZ2SQcWAXKR6bDkF3Sbg7vUpSB3+aL5WD0JZBOFGhQiAoeSer3V
QeoM1VvLlmS5Pd394d1AMVttoAETuw4XvFS++Y/b5QanMNlorihQxSLY7uCMwzg3TYzknm/CbHdS
0yyzxQJ5CuCR8b77zqU0lTVfvX+CMZvoXbJ0dHcfbCrXHvzYtgobs+EHO5tg0umETDdnezGsUnid
aaJI0Dn+yipkMjq3VPqtM4Pku0Itns6EuTRDXyo++DKDfTRlKR6Wm+QSgkLwoAEMHUqAKcHs0IBV
ENs7C4aZHm4Y5eOXkBP7qVm1xd8PyZs+a+ihZaW0axu5N/3nylYE4uzp0Y+2L6N8vPXP+fRKGZ6X
5jpTnYn+qHZ6uy2m0o7fl4N2eSpUkgrXhxADau7zDq1WIIFBsXqXx5aIErDb+pMwB4t0F4WYCkym
uBX4W7RMVG9ykYoXJy15AverqKQPVLpcRR1CF8Ogcmd077IvTmrHkNeqB94fb4PAcmen9H+OYMIc
NN6F40lthqMEKY9caP2OpkgPb97CCDSosP1/c6W9QZ/DtRwro/KYLT2Xoq8fU5evzRZYgZgUq8ZY
Gw5AYSbfSnyWFiQ7izAZQOqd1VpWyghMTUfrklEzL0Oh6wXjo5v3A4EybCwVzWVORxRUgzIkQTcU
I6t3yDd5q01t9fmNmgmMjrttGKUuAlMgyipKDOM5MczKd4C+on5FURYnWYD1h+y/9fXETeO9ieBg
h5OJRfFq1IrC2GlG/IY1NU2JuggDSBRtk+kcueFK+OoJ1wnIWBJ9PcPLIIHLG5R5nUKImmx06Z16
ojYvTNI9VHTltgnniFOdxXvZhnO3Y9rjpYQozmkVt3dY7xMpLdxTO+g1JyD0FHxod0iDuubRnlms
LQNgmEtPaH1Law/ghZUagR5x8e3aVyJg3Doo7TvAcWPmOWQ/xUsXWogCT8vhH/T9gyOSpJZFzZt4
qMlegBZ4U1/ov+0tkfn04tLnzpStJZNktGvaAE0zuQCXxs4gfGmIE5qmj9bJdfMCZmQZLPY+oN3w
J+Zc1q6kMHc4BpyLTD9SoASOriDrVDMQinxtn+ZZudt71SvDegcVf3+hd6PamiLX21TExN+EHXD8
QtgDrj0TPyYbjMtcfGDdKIAHYof1xkz3uuWCbMM/d1aM5S3Z/G6pVL7ybPWNue0+G1iGxXhIiGIq
734bKd65t+i1OLCm6qTb0Lje/z79OceW9wdVA0XEx6qC3610NblrTQofWOXxQvw0NwlnTJrmGFgd
0PySdUf5AvruMql9ADFBK2WxdAB50Oq63fup9lRqFnQ6rwlVAAdvdMjumCnNIM+wEkQ6+o+URLKn
1wK4FR+g6gwOEvsKqHLwTs4TAcpZ/tAPbCQX8hxa6cwtR+gLiDGJ9NAkKCJaPC0Js1K5rfYctp5c
kg5KEpdLGLPYVMOhq2PvJytQ32a0Caf6fWUKHCR78wimYTe/dcUPh2GTKyRwzuaneqZAuO0rYzDv
9IV89XqsJ2Gz3TIG/awXfvPFJZcSRYOloumsd9kXMUS6jvs+n+Zp24CjH164GnxPNGprQLio/82G
Qa2v8DIICz3aJeZP6JEo1fk8DvuLVg1NM2e7vCIi3MjFDffEu2ahhbVyDfIy204oRYyc6ZqHGmFs
1EZHjE0svktNRAIjER2xzkG3S8ATMTWIcP9toCYraNi82RujYyE4DE8m67Wt7bAzOSKx6a41GiZ/
PF4O/ZB8nv9coQmPmp5PyQ7DE5a2ONryLGOLzk0gR7ymyP7s8FWS5VMIjNFnnD4cYWRyCjvDCB4A
F1wlpZ2Ca7xXQ/84Qjnu52/2m7xB7UhDzGSrnJfV9XqIfiUTwNqBjVhfyNLsy5IdlSEI1JlBaD6b
gFKlW1qBzuG2jHSO0gIgEA6bKXOFB6zNkPKtIanuJMIzao+RJOdKxmsi0tDZGJjykJpOmiL44CTh
2QNVN+ifZVDeZJHpmXDmJFpgxh2vU+GrHMvPA0YAesEbs2S6VEbosVq2oacKv0asmsiqFVrvRDCq
3anf9SOduasgU8vFRJqMEF8S3tbdPegiTOvprzLsP34q4pE1ZVb8ipb1cRhNJfXq6hp6jbBawTVp
Lydp4omLP4UqkFKpP3csbKpKiGR8SeQB7P75GC/z0e23Lc/1fiMRLtPmYM/Vf0LDFTA2J/hn/jZ9
kROXlzX9y2YtX/U2P96ElECldh3iRQ8raPkQCXWvtnmZS7pViNkxt6fgCN2ncEXa1ZozibFit/z3
C5CaVjbuXcBI+bDTBFHmdqKx7wKQuoqVTNBRanPdKYHS1FWc3jyeoAuex3FlRg6THSgqZVG8CrIX
EuBAVWxjbjSzlUWs4RruFkReANozto/AdaG2x8pVtzPA4+qXZhEgv4I1Rf23IzoXs04WXFrnT2b/
ukZkd/tZ15wDqowx8L0R1d3Dvy3enKQBpp4GKvQ1gwcGxhT2zAGRQ8jj8Htkf2jCPJ49V56yam0w
YNIgtLguJ2mXwDCLToya2Kmbwe7IF8/a3pczn1FFVOOEzzCRYLtw0FkC01wIzGS88DI+4KiAm8OY
W88hFzlyTMuFjz/9cidnPq6MV/pGbL7KakPxvn/yMcf0GJqoduVNsjykvvFAHzZ2vdLPjD9P/UnP
JAGjONYCWQeNwJHCRCWLGqg309QlpHwwXddI0QC4iLXazjGv4+QQpAi87gQLxDXio7uZVsF5qINX
WM3GWl+RE3vKmzNYr4h9HzbHU5TWNJ3g0+lZholFsK7ZPHMBYbQUf+Laykt/g+cvg+STuDl1yVpq
sPnhQ+kJdRSN6I8cGOur/srVNEjJ+1k85GpPQNp5vRt/pCvqcy8o1Bjohby9OJV6ookXTNJUAYwV
IBWwBQc/Wt4q9lWBwi2Y23IfPnhK0K23aehHZGuI5LafyX4eQpGU9Qm6sRZ5bcpng3rMRdoeWocC
6Pa7uU/PjC5WTT5kTpQuBltCh1hFdrpOjTL38PaHdihMovg4aQxMiHbCC62fPpfzFZZhaxwTY6sr
FbWaAkHTqX7XCZg2yLLpzQqFkk1Anyo2DpRldjYtZpmA0DUcskLOvJ7SbJqVuJyeUfGpEnQ8RZok
RreYd5vVMdB63FBvlP28JcQGkn4gTqX5Gvga9yXXRBLsrPcY3q4Ne6IZph1sOdyKEGkAJxuirxIJ
IuXFfRpOZScq8tr1NudjoZYVquzTIRoRchZFctZfBReQz6AOwbVR3RxbJ+igVuqO3m3yX+LbzvD1
UCY59mMEwO812p4tn7EsxlQG+PtQeCtE13GBncaqlUZnTx5zAq3aBs1u27ng8RNMUb//XPcdf2W1
k57uq5uvV9AbC8so88X87bcPoxalpqZs74viMnz6BIjdWatdmtt8A66UgeoHzJCgISv48s9APrdS
AcYRv2pFrwzx+twyKVvEu0dkHgmv5xk/zW17JWoUxSl89Ee4/1PrRGiTB8NR+sbKS3gmP7jPXL/6
wH0q37zxTjrC9AkrwH3koPMLexHY0Sekl/qRUjrNCo39Zq8Yv2BpOnXFcUOf9VFsnivS/YlwR0lT
zdfY7bNtwJFskgUIhTbTPB+jECeM4FQdaNwEwqtCxPV/J6zYnrZ5XY35WQHykMFFrZY7GUbTqEGn
PHrvF6SqpxUhNQuYPE3iK5HboG2U3B4eN0ZngwJzo1N97eMOOgcfF9Zrt9fc++5lB9vDDnnAoDa2
exy8oyRrpR1F0/9l0bvXrXitX7bzrzSUJMFsEma5Uk6yUe7vY83+hNEwOtQ9LRmdWdR4LXKF9VMd
X4WmsSUpz9HjV+aGSnb/XsmPlBv18QEiSii3VKU+KJNtv1XI5/aNkarkvfbk86ZsW+Ng8b9dZ3VO
6yudfKsydp1k5IJRB+swsE/EqScXDep/RjJk6f8gKrg4y4UbmHUjv/ZkfDq8cbA+g8heNvZ95kfj
WC7mO4dEMvhgCjenh9KhHYK5lbT9j74xzUtBYwX2bRzoTkv7tNEz5C9gMvzuL04Ml3DKeYKiAL1n
VbMMNvrzUl8t6r4aFqRp3Q0wy+0D4wFWOaQy58s0P6HH8K5YY+6QrxhPpJlmB9swxKNeiBzgVfh+
yR/LDDjBzM/hpUpfIKh5n/t0HSmydBnnvPKA7N8AWaQM6TODAjNPRZHA8LaQeGhKljc4pY4Y12wx
M3E33g4tHe9UB5ssEbpew6y2Pxz5QlG/0HGeFmtUfcQ50J2CO50MYRbnJUEeT91dsXBugELsY5mk
d9wOuJ3IKs1OFPsFUCWJGj4w38ZOXVGsdPp+JA94chCevQWLhWqNzJS0g3B3BEnQJfnD/lPlGjFf
Us+DkH/lWveunEXGV0ojas1EB80cl5EEf/awrGJRLWtSRSkuRtM9fGC0Xj2l2E0JuF6evASQ2yE5
x33RUdliB+snCuSoPwbEMMc/Sl/j4OxcSzvQDd2/nEUBrJJ+jxigrzgNv6EZO7Kxc7SdddFrIBIB
pXxmmI/0htagzpaLSHNcetJhba1ChKPBGz8ljDvBQjtkmIRBZ4oM6taWXI0Pq740/vmY1c8rijBn
fLeGhkLDpWYKaYJQi0bkXvj/LyMCIMvW4Rs/2zgXbr0/4YYaVw0lNFR8dBWVbUAB68A2+XSbqIO2
Cbfbnbm7J0Hvgjezgj0smgkVWBySgVzQNUF2ZOD74RlZC5Q/euvofMgOpR92UDu/m8g9QfpMTdv/
n8xNK9NmcZj5a/Pd8KpMvflpyhUS+f+CRhgc2KcRRGpZ+BQOvbonAeKiN+wm30nnSd4HBlb5+iMJ
8+2wvSaYN7paF5nqGy26oj3wXwyfUygVAuefexyrnI7sWkMvZQq/1lE3sc6Vw552+rOXHUTM+vyk
crdzw5AYnjXcSoQQJM4oh26SDDHbGnfLfIqcrPyrd5E8FM7UGESrECFvrNhQEyN3vNap8cHEh/Ha
6nmF4rmNO9kdvMl262N+73R6xHxvX88ttDAasyiwmg/b8AMW1Mly1rJ3f+FCASLmmqfQqwHBZdtb
RYOEnhufpZ0MKOWpyNff97VusCdEQQHDzNYsNPWNp4R14iXeTegP8+kWzWD2zTuoFI7BN2SnNrEa
RFHkMCH+yR0F99zA4gfVtD6iTKCkd+2BFnXRI1FkwQrPg0hww9XBaSEnEVf/A3L3RF3I1VyVd3Op
8yevXOikyxwhmCUWZsWFl9+/E+8oA/CASY9WBXy5Mta7cbrJGOUdBU/ot75x+xOYtMCsyzWHB2Ei
xKqW77BrH9MTNanbxSGXO1a8dMvQNktcbswH9HRO3LGnZX3mKVZhImedha5LBFMr2V80cTQPWvcw
RbZ5sTLp7WQMAd6vEu1sOr6kp201lM07yu6dYnVo7GrQV1WMHtZTyHF1CyLGsqnOjW5ncOWxuQIJ
+rcVIEAYEJfhVDz7t9Rr9N9M5vPuxAB2efJd3DduYcHccTF84ah6Xdf2tOAX1a8srNR0K4oD1xAS
tx3dQjEB3RTMZDsXEB5iiOvPCXGv0w2nyiaPq3LtQlOXUJXxcH94vk8Gk4JVcMf8asu/lgeSTGY6
fpHj7DS74bwlnm1/VkF/3OhCGnR+7X8XbDiygimo4EpLvH7d0NLTnLHHUHthE5SZGfklSPcIG8TM
szIos8Vswjw5gZ5QdDUb/A6LHXwj3rYu5KLEyE7CxaRNGMi8veujnIZCuac5/xnvv0JtQae7bXJS
QizeoYnwmqXX8Q0hwqPyuA0ByacLr1bdXBwwWjBQCPKssKuPXXdJawZ8LRKS3A3nRxHWWxkbv857
9VE1BDrZrBkUX5RLZ3RRidDxzpf0sNzHZyOsB6GO1hyumF/5Ms8nRSH4P3uMWpluH1evZnqeVLvW
bwT8Rbho31sIgrdoDQfGE4PjHlbsKL5F4ZQj/McnNTG70RqxLqPISt4oxYuJcHbxw2e0maNCVbz9
bUZQYSc74/v7sE9woAUrzPiHIm2ccarWvVutQmsEh0H48UUPBXitou5KlTsuwDJruuKbzEfcJPxo
xGdtjb7ndGVrjzz4TWATvBlVwG43+gY1sx2Fc8mUCLT8ONBdNbdRGrEq8QkOqHGROtYZPcbsO6zt
nYtObb4IewZ/cqLw+8puk4VXnLWf4vAx1jAgJy3wbneBdrzVoE9NIo8ZByK4CdEVK5pSFDkOY0wt
ql3HDR0fvB1fl4wLU8sWBPkNBV4qxp8+FNn/ZmR7YTWefXbtP4DzVxgyTiyBPq5hXpsr38osLeMA
Z8d9lfTwcTiJRrGxxITcGN5JLUB9U3S1Lv+R4ExNJJ3dUMiQvOyuyJDLjZbXKBJhT0EJ/DFMCsx2
xYjaoMo0s907pHhk0BMgDi1hTlm8Dc3qwNIaj3DR8R107OsMwUPb39DbO8qUF3M5UUFlksN71Gjf
qfd8T4dQTB1pi798ISCx6QWy7sTdEanJIT46JP1mRC736r20PxoVr8AOF2GMdPaGrOjHTN9pr/e0
FtnOCSL4M2Hzzo7nyVwyOVXfVAqipOpAxdCdjBlRjyir41CJ27M9feLR2akpw5XPyW9gfij0egtS
LuZ1lr2RambGVskqeJsalah13de0w8I6XhJ8EUksBJYgCTcWnxeAvz22eyMrjjZn6rpf7twd5NAw
6makQ6AqTHWFwvNGdlr/BEpBqLtecAKaa2VibuvsNfBWjGZXajoY8uD/GAr7+V2EBOqwnqpIowmM
XtDS+Wsv/MG8/HgmEokhTNplwNbTga3QHHRvjKzspr2DR+vBwJwWBXBR9ki9oLrDqHOvdZgYua0p
rIDqKQri6uS7YxuNKMhHpodZZ+em4pisAoXtcjzaEpBs50P/vNKOeoA+7N4bqL32p2B0Eo9UWoIJ
fkqAru8OhCh04xgY+f7U8Ui6bZWkOsnwlNXTdtr1hUbbKgzedJey7UZb+XGS9tgrg1COaCljGtr2
YVKAbs18AtFwx1nTJUlqY/GWlX6vfhgTjS3KW4rFGEqZ+HucOBQNvNJfhKJSSI5GS/mGsWSN8QAy
5TJx8y3PtSihUo5Te4rUiM8xMxd5bZtSWoL+NDudOg00c7tPNuT2dHWPqDnq8gUkdR98W/QoNDi/
u+J9+r+h7iXe+8UbgwMV3sWde60HpkoMVdfUOiJ2TMTV2lizUSeFrS4Yel6e8izxpJ+qxEE7Pa79
JP/1gxNZyfQjwD1uPyjtl0a2jEVtjLMIy9v6i6KewKyfsZ0ToZoLQjeWP8qdz9ji0HnEq2jfiUxB
3BSDVXkW6i4+j8lDCxrc7WFrPInld/9SC+K6IF07HMKP1pk8kHFprITkNr/6Poq4l+9HErf8Yff7
2m+tMscUEqpAiJJdVQxrEioI5bUnrcmo5OkQjeunzla0B+wAVffKzkumjn4nLk6RMNNZwXRcIL7J
rTGORpmotMOOa3MVJfChVSaFIbJtuYJNiskMBFSQESc4WZsjst0+CmGn9mqdD0QyklhnRggtZyi4
Q6k1/0VF7JVq5XkKt9gh+7UCUT8X2CrbcE2aqK9aShIqLRC4GKyeGrf9qqSWaUU/qtUeJ5B5osaB
JaDqyD+FDqmdydBGzh4JbksyUwiztYgXuFBd+z27ASxtg67AGxo6QqQJgPPKHmkQs+uiP2yoHeat
q8oKjRs+QBTN24pLtLZYkhqzuG3M+naCKJQpJOcDseO7Y5CVjsEfT4+QxIqgG4wCaPTod5nGWYLb
Tgd5QRTGHB3zOW2JGO8CQpZ2N50hBgWlccHfZEqyrlDptNbXV6AhHBXOMwMNEhaiKTGff4S4q/JA
zritxHD0mB5qSODFyy0GrkxBQ//qrrF+/GC453AUU/a6X4JKmxt1TQWqrOOrOhEXgwKFg5DCP59e
EMcI6qI6S4KCDVMJlaTbsQ5RkimYIjUafr4AyPrsil6cFuUHhXEH5zdDpEQABSUZI9nTkGrI8Ybn
9Sw6j8OG8b2RmDCvy2Z/jE6LxRYAxemZOTeprSSPhydM8UHe33aXh+N8PdgBOVrE6J0f9nu0zGjy
Hbm5JU/9Ydbph1WbLwDAxPW36k39Rkbv6ShrMTFzs39LMmd0yUyGrzV7FMG8I3RXG0Jg5XTnNWtk
Yd9bxIq2lFzoufj9Zxs8WwYs/250mOACnbJivx9+zpyxL4YvClsKklPF+iDK9YK1fVSifWS+Eyk7
GkxNI4hZBBr35OCHujMhXJDQHYud3i6nWK+haV+j9GI6Icrq5RgI4skxh3ZI0+ftQUxgdls8oPfR
qoItfBX0QONad/k9jcNnPlWw9y0faztPhnvH8wnaAp4iu+U4NVAk1y5zShrFtktV2hxlhAPCWKz3
augXkxfaOXGC4swZi/GH0shnC+NoifEiFSDfwL62cnRQ9qIvYliDP/M9WD3Cx2BA8jl8wXz/RjMX
tONPAGEPTJIl+Xq9glbt/SitkuBX4ZVODk5m186geGhALhPRFsdas+zdazW7nArSebIC0PaE0eqk
8BdTp1BxGT1Wrpb0oIXW87RwO1/6OagTUCGR8LsuY5rwh5nxwBUDL/mTwNVuUZB2dtR1U3uVqh59
sdPbNAigzyEiLPqo5NPq2itrbTkJPiyiMDeRMwrpFnl5f4LA8nFKLV1Kpq6ntqVpkp562FNK7S1i
//AFRikaQuuFYZ9CPtd7BFHbaaib1Z88KYxSU3EeEMD58g084f2KgNA2Xpm/zTFrmRDWTIWvERIa
clBcn199DcbkSypwUnEG3rjEqh584C9kGIifIVk61Y2xafE/WABjRsPlHwqPR5hb/wDuEWuQ3ND9
SMIwWTqSl4aFVc1QgDnnIIw3ZYEO0Dc6y/ebb5HJZZ5HlruqILsgBqLTZUPIHbUyaAxKHoo93Ptw
rIkZXcfsgxaaOft5O3Lbt7hiZNxY0iaDDxln8Whod+Ea1LshGmPDEhT1QSRZUriF+ZJrpD9C0VEZ
bLORugsWHIzRvZ3ZSOFoJyQgjCSEUC4g+Tmq3qvjCWzAIrYfqjjE1ecn9Ce4jU6DX3XEWn27E1s6
V+D75P9puG8F1UX2XXYzdx8oPVQXbDUiOUCOatK/+i+56WRNJD+dNw/4+YH1oElm/yIJvhHrDiAB
s+9kgYICZ+C0mIRNF0UNyhiiVUklH4kwjFIBAEgEGVQKDssJN4MxHayHbYHmaXskY8RBC0lUjm4J
D9KK5X2lhR7edxGtWD0D642XwWwNrzJulrrbLcIt/fSfwoGZUWT3zJku2I0VXpfRqKRmUyUtZ2k8
f7FIGAIcopHUbsseH/A0uZEwgCqm5IMOg4L8SpUgTFSxBNuqT2MOwL46ABdTMUjdK1sjkESxMzeS
nNw4FB+7ByVspIecZSiD5S0oxm+fkpX6Rc5Z4k36byD8KTk1HWVE8oDm7mNwTuKvZD2yu/aLfwmJ
GB/bzNRN9i9A87ro7Cu/+WPV7B+t05FqYzrs5kPk4kN/uht2os5XikSpPHjFKC+6cvXHI6tj25At
u4LEN4LYZ7m3s8k77hcx9lY0KXxRkIvJ0zrpchWYFRBEXrkwm5d+qo+D6I58CPIAdL87X0d0pZ92
PavjOz4KaIi/MpMllAhHL0+nfoCQWXv+6ZTg8kEOXKBkLX8sSSPD/IwDtoDQ4Q/QX9KZ92cTn2/9
absPfa+dZnl5qUUXpgD8RyBjUIYaNlZTlEmzR6/eDGRfzjrFv1IWNAEzxiL29t9AAI9D2Q9FYQd/
jCbnTgii+/eVD3KH03/unIoBoXbH1pLPQbzd++SFJqO3cBtC1hiq6INX7ouwG7UwEnMEWCO4IJM0
14oeSfyAxB9ckHsZDBKhRY15eddHi/eq1nhpRWU2t6Jie9f/2ANina1SyD2rH5vHdB42vPbI01JN
0rKQoEfS5+5gKIxFec7BS617wokCfrcXFpJILLY8m6J3Q3YLEjOBUulMHapzHDq7f+0tVCI8yB78
9zX0se5XDTDfzF5oHhBT+2qtaiTZuOpj48Qmvu/TWbgOLWNLCoBIyranNRt+qVYnpginUh4YqK/K
TlaD/TRCXsTQvJ18fdlr4cFZCqS2z7bP52S998c52Nk2gWDsJSJrPVeQ47TkqdgeI0DYcW3pwg9l
PLh+u4CDYxSIqD7RQ0d2NW85tLQwiVA8vTMUh+OHehF/S1NLySd2FfMJtHu7lz3ONSDVp0M9vIUB
ke7hPi+HSg25nnYFqy8RJE8W2J1SOAt/oTPJCa++PiG8R3s2XzeYlWtkHi7Nj/xgK+BMdX4heaKv
4wxQ33FO/dlmPqws7x5h0CFOVXJk+Qra2CXwNO8hlPtchHlaWfPmanwd6CuWB5SJ94ZcqfCR/kz4
x5YyxIUM30MOTme2QESYzi2Gb3xX82uaQyvAvQrE3ioPw8z4X8mkK9/IG0xnPiYHNhByO9PfMSAa
HQng2kPvQdci3yXjF1GIMrlh4T2pvGMiggUcWF7JB+tDwWQEaqQlO45+uGJEMGRvYOajhijBc1Lw
kEN5ziRctMIFQh7akEuu4OqPWRMwq7ONtprkQtf0AHCuirL0dSUFMVA8MTkSvP8v49J/br/1LgMC
BieAp9DbtBfG3pAv2G3hCkLHv9q0eiJMVLjQ7uEssx4nNKpAE1GWdLCm6/vTlFz6etjX54QiQE6A
j78QdHLfersaXxFpvEBj7OH/nkY6i4eox4EOj/sNC8pX7VWvmR1Nd3A0r9x4lslHQyL5au8fk67O
w5P3pYD5n57yl1R9sILsnhGiefozciqLVdeX4DpN4Sd0NeTZsw7WPLl8AxSwAnfgM18iwFbuaJ0l
XheMBo6vO33W3ERBuY2vwE4GEqifI3XasS1EGlW1wn/W8NcjHsZ8RPIderc0fdYLuvOTOBszVLsp
zJatToI32gP8noyuSFL6FHhS8r7CbWCweMywMFxLMqEXSNifgTFj1AoO24FH8UkQjHN7t5rKo3S3
B0Q2uEfrb9iRgQnGJgrrpcQY1XDMaUbXl88w72oWHt7eE+oZzoUgWzWLqMhIjd1CRKgqkket9YxA
HMJt33GEBzTriCX069YLV+//++v0zOPTUn2YWPPSnFMLMzRvjjdAtaOrWMBslOWrdUFc79sF/dYv
VcRkFV7A0IEN9CqLC1CKnjmRTmZbutSJJpntUGsq6XW3AInndgyRgxUIDdsPgmpy/wHKRzK+X4kk
RKxrNjN3KBo5lqsYLUf1c1T8xwbiwxGdNFtsET5hviVWmp32o1pLiujH+o8SYaVrfuWdvmayJm3l
khVmnLXenlp4IqofhYUTkBa/rnrnnN2qQ7FcVyyoXvORp/w7+8RO0NO/ZT9jhxaxmPbnHvR6KcVh
+EjoCchJ8Aeb5AS5y/h5fNf5m08dJuT4Xiu7xu1WW+JEhKSAIALSkjGE1/VOcg3/4z+a3ivRLIk5
cruleV//fW0m3Mu5gfaW8R1mYG8heNymOP/xgQjgPueJ7m49msV0zysA9x5C7GU4ys59JOn9Lp6b
zjZgxFU6lBAZbleHQr3KahmbScaqLORpROMfePUBnTYE7637WtW0OMVAoK+dBfsfcEeDI4Nesh4W
e3GdlDAf5FtUcReX4zJWSjbcYZ+cpStlHaotf9Vt/quRvmWNyXqalAAMAFRMosHcwCU65lKYf1UQ
jjTaolhDgO9ueA0vagciICNCwSrk2auwTRMDaQAx9HRp6zc7T43ufS4F6rKYSFgcrNrGq7ZEJsFG
krnSyT5Q1m5Orc2zfgHpuiOITAnuD7LR3qlV6497096ydLN0IC4Ob2sj1Rc7X2E7GA8C21BdHWLl
3nVyYtR3jTY34dKx+MgV7qIUZ7U6buQ98aQjcacEhoPzUz2A2ELzAMc7MiNhd2P8PUv3aaTAo/az
TkG7sxtFvsI1oRz0zC8GDV2BdCWLZN/bOSEFR84bToli/ikaQgPLHvEChb9YnaYIDbwLf3qwvOwu
biofs3wYwcPxwUeX+YIiwYlXJ0lSEiCdIMIlY4Pa39VrdDhsd8TgG3NmAqbl2v9tQtF6KX3cz7R/
voFsdxkhMFUH4tiHDhH4rW9SCqM+oC9pbm2W1eD65RIAWeJxcjmZE4KztGFZ8Av67vPL+dtnZ8zC
MnbFYkNSIp9NrbrGO98hTHhu3iMrbMBaKhlVAtdUwpodJ9QWGJ4c1NNjU94Xco+cb0Dg4ElvzJwR
pCr/FRnKvJ4kz2lEKiGuK+WmsvfxXvFV0X1TYiLT463sPKN4kS/mJrqdCAD4x9UsC0ux61au5Min
Ie+mD+Q2WM1JULiohiIiAb3dyGAIv33m5ZAdsyQ1fjd3qgOjSV5etdnPAmm0YQa+eNs4hGn7Tn0I
nBnHIFmBoPk9tCPHv+e7YWrwAXtWZ011TkznPf36J/gMC2rp1H6QXDh3rImvNHxzzu8OsnT/S3sZ
vNAXlHlA1omDeW8MdwMEfaZ+Cg1S0/cTyB2jfzHxhqXo6NSTiXDVbzJXkOsTYjbJ9b4TUk96hlXZ
FOw/QGYuFImfx3MtJSxIrxZh26/8m4KkPMxlkS2ykrPvbSCNxpNl7uUAaC8AROdvvXo2/vjwp/+k
mRV+IvZFzPUu/RNzW7qnBpozscuhVRYoOHt4H2CeKFaQrb2j9+r3Ftw12WWr3xgG1g19SUMGnz4O
3asgD4Xs4h89/ZjO5HBR1Pq1TmJsFSlhRKti9iIMfP++3TTcAAhBiK1QRNrZDubdZ4GMGW2YfthU
N/WCanm0MM1zBBcQhWAJBj7KK1+hKq128iZns9XrvIvpap7fPwVwODlqY68BbttAmm4fIzB5sL90
w2fUCErA5UydXbrkOziy1Om32z2fSzrYF3DSTF5IGUDkKdER/VOM5kvawAYgI4NLQE9vXsLpGXvI
URooEzYkT+MCQPwGH6xe3hWiz0JEf57JG8IKMO58o1LoMk7WHRgK4k1glMWVJkyOK/0e2ngt02hP
3k6/DxPJDxWNdocxoPjxtjCWiI9xET59Yqx1B/d7+AeHzU2ppufScNyTMfmFAbZT1O4mgBPN4qgm
AE+Jl+m7//RSWaENh0RWXmPbE5rVMpyO0OAZkHO+Ys1hxw1GZdaH+QWg9hswag/5XWB0fMl/sD3z
2QBs8L14dHOOEu3Wp4Cj0sWr91iwO6UDH3H6l6HM77CSTBllu7uXP3VimsK4z+bmYmkdEVDV9d95
34U9lwdalLWa7sfZgzG11S9EWb9u+I3xBkANxft4KUpN3NKTI2eth1BfstmVSTe5BuFOsdweFuEd
HMgvrQlOyWPrUKxZX0gh+atilWmzxQMs/eUEwaxaZwpgsDyCY3DGASYTmc7D6dPsVg8H4M/QixgQ
RMG+4hOh9Njzj3KwIjW3AXrsE3XeTj0H0h1ov6P0SZmcaeC0zItDY8lWFUt6IWIYGSualTW+T9Eu
Xh2uHz9J98a4ZYubHE6d6ko6pA1iXCGQXfMmQyr1YvM0bsLiYyk9byOfPWRdBiA921naxOQTKEFn
yCyt1c/OUs9NQJyVLJrs83IIeGMLhafdjuAMlBffFez0NaC+gjxUjm82EiWlCZuLUKnMMaQenOWc
Jcr4XDQ9UIBwR81AAAQBYVV0kHanICtBzDsiPE1mDcy3y5EfTrDl9AQZo/hbqONLkMa3RUhUt2l9
J+OaiplzNwlk5AVvb7xuePar+SJVtEBOCooSSm/XnCwo0ag0p12VoJns7YuCDOFi3BVVXxgs1OS3
VxWkOAjvnwz2Um0CB3gDd4ZJbZOQ1GjRnudzoyDHdWTAqXLPN4h+l24uBCre054kg+sx4Q+bKcQK
8SBgM0Nn96CsiEEzNLPSC2+drNkpMoB7sRmXGD/UuAi9xEzJtyPcki/P10ICqqcRf0km0f7fJbfm
4mdUfpOn1UtrwzA4lMWRqE4623z/9UZo7GbGdAG0vfswDEGvOhS7bahUJIUAw8hN7eIdrkuom7ay
ly7OPZTnDqxZ0iphWr9cNIaLW8RV1jP1bakEiP1sf3kcKBhiJw+hljbIecmu/UDJtuZMPE6A5fUz
9U6NLf0OaD/1zD22wINbA7FWLjqSON6CuF2bCJ+kmS4y2d+gMViKdNufkqJkpQ4f29udTArQo7eV
dRZAQfedJJuqhR+ZkEWoVKN7TUSxHJ1lqZyR8cOC7qJEi4KzJBIg2D6BSSWJwPoqSOrK4HQ2IzAB
E7nULlfoecHEvzD9Xq22k2rOwHfjhrYWJBApdU6Ea+jfzFk/QDtwFOFHPMBkpEMsfGEbaJzBkI9Z
ZIQiqhxKdZdVJrUMr4cUS0G7N/us6MmGEFZqneH78wzvmnKpZ8sFK9gMUtjGCGL7F9sHnelKz/ji
e0zDt7pf83EWT1j+9c3y7g99ROWzGNoyIOQRcKYK6oUz0lhEkN5OFbRwLKEYTlTNqJEgB62fPvqj
wvr2Fx/XXNHvQUGbeeQ6yFezjkojwL3rfF0jC/VeTyAJUYU5AS/ZtNubTmBhLyGB5icT9hJvPCth
RKwaYU5BJxH1BIuuP5CDM4rz52xOaRgCSnVOfJi2+2oUvQpj+OBMc6RTs3HnD0oG0gFdRfsnx1oL
QVv91GMwNfnCBFdvOlu2bf4PlNDQ+LhRxrSg57hu3elsCizf/YmG6KbCZr6CazNCybFTsfar1CHB
brMSqJjgFqFcCY2M4IjhIBEfVfsbqFuIKs9Ent9ZEhlbIvODlCwe+s68adiAmo+oERprqr47zKBO
QuD7C3bTistCA+EMcdJwjjqIKmWRDYpFCQgWBWnzLfBkLzulSmjgrmDzyniFRm6ViQVaya5nL1Yz
3LiU7ySNGVStGZvmJwmhSXrQOwhXX6vCBij0ITaBkaObpmOap8QvTnOkEI6vDVmBGnUHWis1Eln2
TyogGFHzZRERk8L6l5BPxgR3F6k3qMP6SyDjCwQmKMA8fBzkNGRzzA8YEz4ABqF8EShGrmLqjfIl
DKcIzPlNleU7RkSp5E4mEyuCF8N2XblONr5qDIgb0tn7bEtcg8zWYq5A+ehVTZ7zE8Y6/6hxeFYR
w7xky3Ih30VnL4egHNVnpWcm/AV5rtZF5ZtjzYOypJms92LM0Pi3NWl5PM5lMjKJnpqHoz014cGc
6hVXwWdUJFYFAdJLU/p0CSNTFTy8Bp0uUJr0bWg7DfzWn6xQpj3xYj5Tivb01PililnvP1K+98xF
00GcIhYAZZAugfQpV4w7/TvEOqzVrt3oJM7Mj9JLYWAOVbFmlT166XCqGOJvTOCdyKVtoZkNOx/2
YKoZLpgwdUkmLffhldSDeFRAL4wBnHiewIO992CMjR1Ddp90fheg4iAKNouaN/s9EkgRSOs3mk6h
Tz7f2EoaevSATgcbyDhlbazsNWawCQ8Bf1qrNZyM7Zs6PBRIWxJxH0jza9f6xW3Vao1OLFfccDxO
QFDo4fSg/Memtt+QmfK3huCLOZrK9JwQbAi55MZAJxZ1Rzud5RfYLF1iCljVeRKfFg+4b0vqiM06
R82tHmxq4Z9jb91TOYAdEB6iapGCeXO30XpH4OiOO1L5Zgja3lZPj8fB8o2T6kavGD24r1YOFSo5
JORpk4EFdJ4XNwNbLrBTc+dpHtiGa23OGdO9xYEJesb2cgFMfighgXCOGahIcBdbHxMRQI3nuDej
r2vdib11a2WdE0gCnKupSyaXpcjDG8zhgVht0rQDzKfmcnvQKsIu7OmAE80yzlRT/W5jpEAztmtL
XDSIW0WQG0lb6AIHcerRJkHdsirOZTXYQ3J/qB/UZodMxzBmEPzTcbW5FTuQXZ7+oSnYwkTUGZUm
tFfvwFPiVi5aeOMdSzbGxDQpx57oBE0MZmg2GHT8U0y9XVtnpM7FmxO/VgnyWPu4ss5x15JbXIiP
8lzqxwe4jeoHriOXYA3uG/xKVi1rljjMUkQxjY+jP1CxnT8VrLL6UESbgsG7Foc3gzEU+C81pAOL
JT2filrhQrWFpHN32K2kGVoozQRS3zHdmSERyKFouZ7jYr7eeUOSkL6S4vrwc++Tlow3fXknrCFV
QvQWEwaH1GjRRqJMT1JwZWDub8DhZVrETQ1Sct796iQNm0nHPWaGxtY0pTLsgubSqM1GV+8TmpK2
Mh3yH6tH4EhU7Ck9geoMl48zxMgUaTxiRmVq7PPA9JpVKfWVUvtqkVXWoG7h6DdAnyIJPK2sOGmJ
beBarxh92LLqvSEXUPyif1sPFggEpP+V3I664NyWqtXazMRDgn0rCd8NknnM2U6FQ04vFezIfAlq
id8JUxwNwrtqIUGIZq7x3fZEKQRmQBCRdy2hnZZ2yOSlrkPYWQyTHy/PUaNbycgnwbCYtz3Mq6V7
E3rAD5weR1a9+KFgQgnNuQH0ClhMoiXdUUlZLCOU/aXCZaQAdhXb3a671pNHOHV5j0l6osm0dpau
JAAZkLX1RvyTmfuOO0BF75MDXI9upW+wFMs543hLgJbghyr8EHskNSosNrWLXGe7tsfhoLZiYxXx
N1QVLEs484Isqzy8IOq36wIEZ6so6/9+j5+o46Eu0W5orSlqWvlemPml4wXa/cENx4c8TAKIb0rL
LAgs3OnemSTb9h58+gMSkrvHRYQthMuRSzgR5FWo/E7zkHsakxUlrVnpZosfk9wvk/tX6BKi9uwb
fxzVkJoCdV7/9Mtglkk+kYnJenuulnNCkdbSflGs0ULhtIv2awGsqguKzyouTz1s8EFXLzRBAWK8
c+ksc0ih0ViidPLWQxFYV3A5+iXuuD9LMSfmxwzDyAEj5//VGUNizTQFaNJkU5HGCDyEeQAN1TlJ
svEkiMBgstOViG+s26c32ZJpmrjkVNhH+Laem+kvJe+tuPPNqFdfmNHcR0FTHxAY+I15uE43+Wvc
8I4ALJycspCZpTFFs2kF6rqI/l5jIGvqfL+ZMdq1hX3/d/7W7nEEdzQahQy0QOmPwqcE7oolRTS7
xAgRYX/7Z4fnBDW2wsGQmNCxlV2IiE2magFPA4Rla6xu4NyilUn3Fp87VDslkOQIOe8CQM5qFYCA
zaBkDsj24ZXsjGGQmPOS/8P5UgWSmeahc/c0bo+SSFPs5D8QIDYYuDmHcDJiqaAW+SIfGKtNYV5Y
bRSzI9Jfr+2zxlLhMAXkPKtLniD7p+gr8A3M60+5neaYOGhbDukNJ0MuwfIKiQOyB8+04p/3XSzz
eBeCZZwT4nBTEtjBgMSWhdkKFsZfHwozH3ZMmiSty+6ubzYn6ibfpxJMbaxecu3vyRVQWOyZ2FnD
Q0oiJN48D6MPxLD670+UIs4yJDGgd7Z773sdpiQgvqQnUzOD8NypK9IbRHz9nbqTs1sc4LcgHyV2
gqmKWe7Ia+TIS3NVvGgrldLnB8VFt/BDmMTtWnWIsexjgtjl4eRV2o77ZuG2GBUBRJIO4I2adfX0
icxWIIs4sH5VcqfntWI/VBA2KY3zeI6zerLhxZrF2aYEYZ7Tn4RK2kcaUpSwX+JNRxHeew1Evsj4
8SG996n+g8WO4l8ZRQKlTbFqZFpTmr0+rsYakiQ9oh8LygHN2Z/A1C8OvLsPkQESzi2uhjW60o0C
m8gl+r067Fny1sHnPq5Qa+MzSzEgeS0IZUGRB1mGqdpr++G7gw9ulEFwjWkXaDmhC7sCQaAXE3ZN
dilAtT89835XUE0MQhJWHimezGwd8h8Go0wLz5+1KGIyPnhZgI+6t8Mjy1EoTCsnXqrsq/bqkKbn
F7vDzoYSQOwlLGcU65VnYacA3vqz1S93tV9p3qWf0FvrH4zwkFYpIND8+ftS27Mh9R8iPAPe9vjb
m9cG+5ZL4q/geJcj+y0ZXUQTpPu6LPdCOqEAja053LGiz5R+XaAuh2tmP+6tma2dz3H73i2rpYVv
h7myYm3o0M1X6wwwZnYI5djhEDG53fhgx4cQE/yYEJ85tQ0rhbHBUsKYAJMHsNf0KYgyqZK83hGv
ofmaIYY1ToTmVrBPILR8VhI2S4LE3+kqWIIPLDQiy3Cvl7zfr62c34GhjEqWwDU4XYYDi1jc1snb
PUQicOGPBdJZte/JYtX8GitQtUzquOTTk50aFFjrEbEiwtYu/qrMRqfgmyTcYGuuv7eLXM/o5Hpr
TchHl8CxGv8Z/Jq9qRJ0mAkp90glZmrfK1OeZvowKJ+PHUfusCyRjCdl2hHABwGYi0l8686SlzbD
c97jdORxF9AYV/4Wt0/nQ58foS2ajIx0R58OkDLpTnuTUSwiBrCBnAYADBbBFg0wILOryqj4FPaZ
eiMHc1iDqzy2xaniA/GgmfQmnSEUErVnvV5GaXb4LFq5eg0w2C9hUDWzkjB76eFdlWHvax+FERec
sg5v5OUxZVpSf9ZcXdM515LjEwZdVALA3xCAddu7LpgBsRFdCiyPkc/eOCapjwXbrxOLB7cO7G+q
GFdNolqDINaNs9ixSwCsU8M6K1QPhYl/FFODGnsAB5iZAaFV0Fbg9OBCZM98BnoeNewzDgLPYaoy
UcbaT4ED4ad2wZVcCjFi/vfLRDrw5wd45snDEG2oP5+gFN3zAsd7gBk3IQce6SCpwbJ9r8ZdmH8C
b9Tnk/cHgUpSdDu3bx7BxO/yBIEmBjW4cbY9fh/cXtB4xxZAHypCeJy52OA2jM44jXMBDnNHZ7Df
jshKn6dxYPuhZa4bDC/4hCLXa3hzoe6YbKyLdAQAPUWj8rA/FLFf7IfGy14gciSgqQJs56Cwac8I
8JBXYS6X4nCXU3CNkTk4+cltxM9RQDeZWLQN1eAaL4peSF5Y95Iqlt58LoFJsPvIM54fpb6pjs3b
bYO7kmZU0uOwWmQ0DKJiEzhXERPZTK5rzQ5oUOnWb5ANxed8n0HlWtC2M3SPgu903OkEfyr8EVG/
An+xteELJIoebyaVmnH4z72jCYWxitDqaxpd1mGQETw4E0a+xM0BFcZWVaIm8UVfS57lxbtGa53A
K5W8blA/5gYYQkJTUmvUJBQ4dGdE002ZTwUDJH2pJ2oJ7YTKDm4qM57fA8M3iriHzujtKuv5rUzb
a4a1EjfP8+Qf5Ym7D7L7Tsf1++Nj5PteA+PYuBBS1WwDkHwxUEYfTb60fQEMjwPwsvrOKxeE8N2A
lzfUaC8nFrY2splH8qNITjBaht2y2Y47s1bJ8UwhdacRXUshQBjE3gfnjqP2qPk3v2iqI8QS8ogd
1/wnBFTd5pUP6smda2JJXkpwfNbB2cVZG4h9oiXxHyKuNx91o5nC+5sFOq3C6Y441ZygkDo1BIow
9IB8kRlMD+HKte5PjnJ9Z4WTOPnLuSw6dj3vSeLd5fchBboDmvvUKvqdWpZQilmeywRjVZyEvWPC
vdcJo7Pz2PZQDk4dFYgvp4HIx0eEumdoMDnRc20GXZMFXhAvRcjlWXOE87u1VC48h+zGww3Y3XmI
Y2qkbL0JGnsQgwKQEgqewedFwAmBhpcWAc981p19uxoIZgEqkzV3VXnCWs4blEpTF8AMqup7KtRr
nqPXfQGNn8FhZRBh00YpTTD+v6fvooHgTH1NOp2T6J0CYdOXRoR5lEdisAbG17gI0QgBq0S2CAnj
k3MG2PZe6Su9hy4nctEEavlaGgRn2qs+BPsMoIt3D1LOVLq6qA+EUeeWNkHOatuvxXnEJH4Tvb77
RJb3z/fwZM2ejGRXCF9KT+YZFOkN1R0nLAe9+2ZGLQRCZGFuVD368AvG0K3ACzyap3710YKWlZG+
L3zXcODgqqgBna9/9OA0aFuLayI/FmZG9T7OvuhkwPCxrVqYO0T5k1v0aHYIlDlucxjyFgUZ0jPm
55sd09WAvIDyJ3Gk3QdnH1LnXc30oumWAqiv2ul5URZVfhna1k9pwSONLR2cxDzv7hCFL4L0aQ77
7659sWfsDZ9R6B/yF00aWqlZvUAk96TOtO6uVgVX2Tsi1sDkfhcPBehxpSWwaqEyUWv+amtmBZp4
Ri15MygdRtBuySVfr6ZeiZhA62+UzdbWuELazf6oHU7qX095RoMLjmx3o+pCLYJZEabIbFzq9NwI
O5fM8oOvkwIbnGpy635ghnhn9Pd/SqTrm4E3Q6bKS/Vhus+igk5/HIdZR9YxWlR3HzvIwuSRqHCt
945qWpigLCtXaB2MPmApShsf71j9Q/fA98n637rA19GLipnP1zBY5zRiz4tB2s8KgOF31ZCd9Dzn
mFvEobdNVrY7LV5lGLEobmhH4K4r6GD1mXVzzVxUA7IPOt3Me6mEFpVLWICZN46m5YqjIx5ajQAc
+0Nqysi6ZUYPlCNJANU/VImRlKkbz2eT0KGUg2r78vIRC7EloF6L/7fZKuwWOUJfZG41Phyhlso0
6edJVg/GX8npZjjSUZh0+FvPUVM+O62rzPbVQX4oAY8bbNH56JPs2eenERY0NMAzKI0qVjzIX33w
P4kBmZwxT6aZD1WX3zeM+2LmVRBiQ8K+AP26hH6f63aGMSbNYhzOGCePsDIie2FGJwLyBDhTiDM4
2N+bgOmyirHM0KxqccRrYt345RAEEsjFpERoXqK1MSrLEfmKUaVculbw4o33bObYUcw+eQ0AAOlu
3vklCdoCNEMPmuSZG3n5Hw3TinBS+zyyh1NwE4Sm/+TlgANB6sB4MijL8n+/kDs2a/A+5qH9sFh8
OLfyjRVISuDu37TvwcSeE076Te0wE6C2PLbkLKIJj7WwXfo0t/0K1MvJhU/Ou/em24IgU3P2LBtK
9zMFvI9fyn+HiTK3GUzrfsnikxvtFjCj0h2zHUOJrx7OA7pYsC5O2vIvtxLDOJIR7VEZJMNSeTdw
vACDc84LclkBRQ0MOD+ShtJWAJzLrCPWN65sYvL5SAi/wKlzwv9UQ/pL6KJwtD9BMUUdrTnt5aeN
lF8OIHDWhlCVJff2E0nMCL6uLU9UXa9nhSJ+1diEC0UbQjosnDS41ls1PUzvlc2Z1OXeHUnJFT+p
pQE9Qmi0uRJmsYNeXlIEUsjR1hvXNMJuEf702rpTMBZ5s+Xf1DPoafCY9T89qjxvK6AUTGk8S+0m
Qa1rcPB6R2+6R8NZ/fSDPfB0909uh07uaPb27PhW+8+obfpnzYbSAJq/Wu6udlz7iD9va0//1jZN
hwIGCnsWdHgFAih5SfZxTroccnFeeoMnAjThf0dwnvH+NtWS6zD2BNA3CKfq0crv3pRE5/g1XdNw
uzC+1ihveRKwDyQUA5FzWrIU7BzS7hND5WCSFoRtV4TFotW3MrYKInE8N5jmo62o38zYgactRoNk
S7XbA+nrKKVV5awr9tkxL4BzRBTSqNIz183LNknl3zurrjh6uzVUyGXauUyUCWKyudd2GZo2P13/
W2lB4/1Lf3714AEtIBW54qX5o154g2OuMW6lKLLOwAcwvxDM5JheE9zn/NZM5yjqws1LW0AFtvrp
QUepG+nnbgYOwyF0ZByFE5/0ZG4sP/Z/KYUeVYCb8nlv9EaSx80hWsab+CJeqAKzsslW2m2okl90
7Uky62ZsTnuzhm9jAKvWoUi03RAt9JR4+ncGCDVaKK1r3lLuOjAwCc9oG+OFtec8n+yx0rh4j9jJ
VXHV6uuKZbXIBk6JaUI2Oho00ySv+IUA+Apkbp76C9Ql4dB+GnIEJdpFVe45h5pwl2L2bYC5M7Wy
7EZdckRp23UiQcL5Gn7SD23KlfZTawxY80FBqRTOuU1rmpqas71tLrhrglxAEMIFvqhpNjW1DKBu
7N8OU/HRzBYjBQP4cLXPCH7vzaiGlGsCUSAtGMDhft9v+M937AKQG/KUpAc4IQySTRqP4ZLrgdIT
hLOHs+u4WBcGqkItsHk14ik0+ce6T/T9ARz92fqHsINiFw45seeiGDPKZDnD0Eg7wvg9yeuXU7uh
hbWgSkHEZkqEn4ojx55/5OhAwGfxbWtWl7OyagT0AvNgE7JI2ZiEFt/CUIol4a5p9/eVsbZG9QqL
WLYVa2uv4W99xOEjv924EvzkRg6jnLiqXuyKD1B6zYm3PjDXK8+HSCqHslbONElG7T+bvY1YnAxz
Nbofc491XPsb7XStUqpLT06d0pzVs2VoeFQXPfpEBlxHv2Lc4a9cILC5qep88tGmTLuLMg33yeXI
ONgpY6QWiAgkFY41OHgW63GSPZUY5nVCN90RJmCd9zmvHgGmtc16zuHhv2t1WasWZlBXd8qby6ZR
3Ja03NnRQiDpE1ewnlLmX55GHqU53exmWHlagU02xmdrpQNtPciELHZcKur1cl64wPyb7eL8HGQK
OT7B/c0P1L0ci2omi5OKf6bUumkFRurIB/f3DAxx4VPafJJeRHUPM3jXZGtn4YyY/huCMGyuleXK
SfE7zkndpU8OXKJI8qFWhyZ3r0Ja4xm9Q62/k1ZPiyZn7dXXWH5SSRdBjLeqsuqxlPmmbiQuAfPK
7eui4ztfmCJZWZnCG8koHJ/OAOwpTiMcPdWdeW0uz9NBs3m+3sb+LAdKbIR+I98OrMukninygP0v
WbREmINbyaR6Gwi7VgcNm0roTpGWFM3QrgI6Ul7XwxvM/UQZ0IzMjEFahVT6bDnTZiwdxGsOL0K+
kY//8IkBeXZsQ+EAAKSzydD7M3lYvOKc4nArCA1BMO6z/4PiGElu9EqWMufwyjaxJoBcVO/gSAs4
E6WdK9MaMMXkjTugv2hfMbg4CRGw/l1ZTHHP7t+XEh7DlISzy+PbsJAwGVRKfloIwvQ/InvPDAjj
oWQSUuB5qRfPaBW03ICktkCEwxDgU0mEqah5wUexRigpQczKvQ8Cod5Nt5MbUn1365H4vjofJD0I
spXT9xrgghI4KOGlTXKgROHu1ZUk23TgfZhGZVd98eGhspc65nmTJ2MwczLc/adxNyipNi0z1JTS
6AY8X+Xxl2kiRApOAIumzonz3Gr5sUjbOhnut/Hi5G7gVjd0KjLTO9XL+ASg163XcC5m88Gkq7kQ
ESJBf/+vnqZPjVil8U7znkDyq5aanmJGx83I/EoUIaTCOlonX9JeabktJ57Fxc9eAm3w+xrdAwAP
HnrOG6dt0MU1PwkJ9o6sge9hhS8OHdw7KnO2YaApyGzHlTOSqbpWlFYDqTXf4hu0W13fFQrms0Ob
Az7yEQQLNlcfaO2QoQ0awa9jS1JaRU2jdWlf95dxEtw+J0t2ll+laGN7j0FzbTMHTQVTG6VmCA7H
gWH+KJs8ErChVJ7/RJu5DXSJ4cg50V8oKK5Lhq5Gst6/NhLcA1h/8C4eg3bGpYRWFSRr8etytRz9
PmdcrLd7Rs4iZAb2RQ5fnEdtt70Zvxov+kNy3W5+h+oj4U7HY6sZSF0hXOFL9H0ixzVELCGYIGm7
I+RY0FhmyRaa0WENLpluWazFgT/C32FY6jltCZr/aMPse4zpV15f8Pcagg4oMo1U2pH+bdY7fxAq
LagM+MDJLUf/H/34qdOi7jFCIZy1oVJsumDu0hC++UhGU+YU/ALGXBwOF7XeViXRdKF4CzhFisxU
gNbYh4EW7AIPvzSydl1WRGhZ9mamM9W8U+iN69zR1wvnnvQoG8A9uXGXVShju+gvr1xWZ4MJDVVR
mV7zJqyHaQvfKZidgEvhPGk1THxKHY/HSuAQL5uBnqiR6EvKD4kW3D2NB871k+DwylxvXUfPP/o2
HxzYNKXZlcqh7led5AwTxzf6vQltNRZdip3odyNtXCO2B2zoUTJREUzkLDlQmTwNKEXtHyO61tvo
8XXkLQmdRUQay/wPn/89RDbyZ4upkVhjwMwvIZhOSYM1C7N3tQMyY+drDVKUGpK54IfM09DNCeAl
DW6oooPJ/iDewpnwbiY1aHIM1x/iC9PX64WH7TqHiR6ebw7Crojr9N6yu3cc+Z0WBiLeq38olHIQ
+/654DC+LjcN6KxXBZynWNWiPjxvgoQVsPOXAhV6mJDCb1uv3KbeXxHPkSg3c2UCVVv2oYC+4+O2
Mc4cS3iqjStBx92ANfb/D3Cybm7DK1zM8PaK4w8Bq8i5wk06rTQ8DuZ6GhWX1qiZbCNLRORtHcKY
dHUWHiib6kvO1YtgkXHdRW0vAgLSZlyLBmiJX7wwXiABgI0dZ4WuKMxi9OzIOdAk9+cNKKnIwlp1
QBbmHaMcFKzu/cAndtTO65RpIZ6Dj+dbynHEhisyRM1IK36HIy3wM4K0yuYT8qG5YHFOFXu31dhk
D5XSG9ixO4noBdzCnADkMc8+NkfZLSspZw3lyywLOnX/nkHepXcj68avErbdwnlbZTYR0bCX32y6
txHgl2nU7bdSrY8kkrnbGOYyfZRUCX2HdDhvesGbXd9ADdJDGzaVPHW5QsCAc2RaXuqBtSxIGsk6
VYKo/PRiP4HR/U9iP8Hknz/1XgSyAXrJ7vukgEtViOMYOfohBv4QUNyyY4F3gTj91CRjumckQKGg
8YtFXr7odEbB09AnpudOr1dwRv6tm9FAHkeJxZ8qJ5Q6rnz5gLST2gN1JK6Gtdv4KJDu15ehMDsy
0ltYW0vRQCbsiHfeJ2CI8aqHvoiSpWfujLpNYxI8rCKzaC5PBpXKEwp8MyPvCq8Ii+MqEsIwgLrN
A+TlDo5SNqNM9ZGcLbJcyG5aFDq7CcjJABjwAM1fSpK7XINhpz0NPW4yT0ufcus68rJGlnuARb7T
tKo8GlRdGUfC1L9MEg1Dl5a4wdSRwpMpuTT8+vdIWhhCboLw6Mos/0pmWUT2l5wqrxd8h2rifBus
UI2Y+stffdrr3DwaQBJSFXxVX0eMjMlZBX5lnxpNjVpB0V4v0g9DbSpnvfX6N0bzT+PCVMDgueM3
KZzvrthgrp8rV9f49UeW5B2jGMg3qcJyfGA3uu0nBX0DSEEY4XrdFwXrNrxebteoqDLCmTn4L7pg
dQPwN6H/7FwICQffY6vZZM9wYaEA6GTx5q0gv4RC7gIgEzFuW0XR+7GPLQM5TWB21loTsLgxrGa+
uWo2Tbfz9erfQ7PuyKyBAPTo4FAAEXTHUa1cngSrQ7JB8pgGnsTcQ572mCEfyZIXXuiFaEa4vW9x
JT2/V6jA2xbe1SjOkc0tcDGviIPxr9R8K4lQqUvA8YGG+WCtll0zY5zzEC4ZJ5NeA/5hnglto2nQ
xQobu90HU4Uu5cvuTm9Uko31flq4R/X5J39WE51t5zIoH/J6BMJP1PwMFfDlqb+RFiwjpCO1Q3/v
rxEQzNUpatKcwepkTI6RvSfB7IdfnZIarggZ1JH5wrYuBp4lIpSbdZGAIaiCmwSne7awxBZ7LBvl
JEm9Dkt9kTXxPykJz7/ATNdU4yOIUeCW8KGdvGQQVLbtjkRm2J7U2wekGPPQcYtW8Q6chff5ATmv
/ENqmpKeYvLwlVzIdtPJQvYIZYS5sxC6opQOeMEcArNUajkNaFEUGYTfbPlrP/SVPAOM95E8Udjx
WFQb3cfGgAwthygbt7IvVcVb12nVR5/F4wTx9eo7x4gkWDGfNTOIZCulM9UUCV044SthSy5SO9jY
sh/zm+Hlw6+sOaIRlS1zRZAfbSqHawNdN6x4L1q/eW2j61c8Th6nRHzH5DDnZTZD95CkTMArphSW
0QHIh9eaVWYmvW5uSIryutIOtAp98GLm49EDUIoYsTSe9Mesoxcl3yU1pwxzd885ldnZIKjJozNn
ig6qK+7qqgueYocpnX8NOD4FLkoEHe87eadZpkuppulAYYbZ50xTEZVJAHWXX2rGqii/9SE9klgq
Wo8/Dke/4mxr+suGVTwgcfYLiNZYsIqMkZvwHvbc0XMXTCSV8C2jX+yA8+A7hX1BJd8XI5KFlKu8
dwmz2RE8PmKZQmFknQDbWGW8nq/RG6y1uG8Z2KTdGxzU53sJNIK3nFHBiebN4n57PSF5XpBpDHry
QBDbyCvYRHr0yuki8KHIxeTD86LbApODZBu3QPzJdUSQB4mi0nCKOOhZWl/hbf3qzBU1ZHL21QZd
g7+5f9KbdFB1xXGUr6fvg8EgRbSpFu7e9ZgFgQ91qY97BSwHzLIT6rAxDkEr7r4fiV0IfE5+mE0i
m1DhQbzOPexuMrNueb3L8hCvfzVZ1VDXX52rMcBul2sIEwaY2CfLU0u+jVKCkoh+b/zCLqn3IZfx
jI2Oq1bUml1T+EAUWTjRcsaYRvdqCl/4MzOUnaRefBFUl3fIZjwHjF5yTGsIjj2g1ElVB+soSTXJ
3y+Sr+htgVGe5lpzaVzg0gjbSumoabKFN12+EzC5jvYAk2Upt9iaaSQvr5OkvbY7LuDVNT6v9rUj
Aa9pXkOp8Lr5K1hnzbwAONwSe5sIO+dNfvcGATDrLoqMM8Vm415CB7gUbJBLwlHB14k6WIvxDqQH
VE/TSv1ZnATqEEwmnZzqBKWMnZprDfAO7anoJRNmju8Y51/EiEYz46pxzy0e/eA+9DMqh/TabNml
bRmHga3y2z2V6Z/Li+hwfwgyCnTrSfjVeQfB5cC6sNZPnrsHtTcDO4hbWEIlr8K+6hkY9CjA34vU
MdXHB/RbJx9fttZlQpT/SOLZbjGFSsOHAhkxqEUM8JvcPmWubTUCj3/4Q+STl2/si0NX+oyGXAmZ
WOIG5GjrKK+5JNN5xVGtKwrEw182EpKfAh1TExlixE/229lTHkC9zfPDmbwEtaN+sZI+lGgxMYkO
RBuT7Iak+ZOFgwtVDUptDBPPqOCYpUZlySWKbqkYhaSoE56zgnkxIyq7subPvu1bTyAZe/4alf2y
AfdEXO4I+LkmQoT0hCBQ5os4LYhekE+HL2rFH7yJutn0gyWyAHpbM5xjejynrofIO2yO9eCzuYLM
KfRqGkAZJI+a750BX5hRU7cm/c2FM8wZT2MYWx0wgFW9Zezbdkp4tqCXTe+nMTIEetnJjkXUFf3M
OICyz4mMhroIK40XnR8Ln+iq90FfzuMHKp43t6SpjokB+ozV20djClPcYLDExCDNYh0UaqMa4IQx
YwJk08RXwqMbVFfltcOni7BMlQqBvynlQRgU5TNlAerk0fU6zRGHfFjUNpTfFl+c7Sy3piPnqTE9
ccbHxX+gJwTOuzEMekkr3xWS4W/IN0gU/y29+v+EA/MilgR+sHPgLWs2htLmNipQSG0vcUicN1yv
/EbZXfET360UWw87hUSZsChOjFqxaluuZk2tCM1X79pVrt0prYh5Ls9uOrjS20lSI/Evhzgz+jyw
P/iAsvBMEWZ9d2+qRvjGCcUXLlZR4HL63jkhuIv1/aHUOlCIuEe+zHE0MVpd76MtjXAmLlYokOda
ajnrZ1r3NkXNsQuvEDIVwWjZurBe9F7/RfttlzUDxChCrpHNnZeNW4pX93e+p+c2A2QqzB8HOUWF
ovAut9Yb3t/lUFPdjezdr4/G0Byhcuax8PeAv8G8h8UOZxHKVzdLPmJF/KwQG2+k5VSU86nXld4q
FcA/K2iMvFWUyyFC1FBiFZhs6sg3zWYhrcwtKvLSzNxtjqiwfKLqZM6JNt1qYOf1puibbZel6wNZ
e98kamcXiHEi8cy+UmKE2xj6wXZN4JUt2RN6zkCf2bt5bbwFlgl3P5yPXCrtQ075MPuP34kRtnJd
ntnQhdvl+NW37oACvnZOiAXPlBSy8JWqQFGpTp3ZJ6jwWeL+LXqaQeYkuwA9oW1VpX85feSEXwep
ZgMjt3Qz9obVhPEhhQ8gjUk9U+2gz3QhS7AxXVf77q3tiCeQo6MQkw+kd06k7IN16o8D8lml90t/
aexSuagUZj2zMOpPw08jgb6adri+km81hEeOH5B8REKWgBc2tdlfvKQOWFaPBtP6KiLDnCjTJtoY
bQ68q2oPoJV8K/rrUcdn4yt9stzSHcWsha6r34QUc5XSLEsy/Mpb7WW4/5u0VsyLs6KOnQw8lmrU
Uy+fcZg3b0D35ZIn2zdIgBtQy16haVQnac7Q9peWgVDiBcfyG8hcpc6PaH/0HoIuK6gmVuupm4n8
ks8UcOk6nFUNPO0v4aeFLDlWGAoLdpcH8ujJ0bJZFdmzA3r95Wrj2yr7XsdQeuyl/zpSZtgAiJa1
UFP7JbrDjbKujgSWNP6JmJh6rNobDiUPPQtH/+LNzP7vStRCNJnyPJ8qZ2y9Z+vPfJt6JvDzNsv2
0jqAvXCqohWjrAjrbOxNj42ulrmNLnwiDCbJXJ4KibxFvhUd2tZYHmeItpfguFqmW8XHhv7xDO9O
dS1nHRZ0q51T4Trv0YR8Bkr2P/hnm194IShBLaAR3xGaf2lEAb9DHsIZFYGuk3MjsmZX3oWC1P6E
NtVAO67wEHDYl2QNT3jN7Y1sdlwqVSqwKz9UfHVW18zs/U7qM+PElVQFLGDDkGsQepsXIkAiNOR3
b2NC+XwGt9lmkgLhjlEGc8uEhMyhNLmCspJf0chGTmftJLZWUo3ZvML7HPDyP4MD9qIIeEV06u35
mj26t/HbeGo5O06xKROdFd3vSOL88M92CSoRn7dXxiESJ6YqcssbKspaD3/EVQb4GEiCsqrAGJve
lFu9eE/YwUVJie/bzp1t0bylUT8LpcRY7lWCeGr1xR5lvWgdOpwlQ+o7pYge7dt7uqEALOBMxYuL
WwhMuTAzQEDW3WHwSTgcJ/s0s68UWnbaVf5sVIveLOMhFUwVU3WcSHanEYhLcUj1af5h9LYHKR5c
PttHuG4zRmfDK3Ze7oBx2XB50M1U6ISZSAFTqEvyB4TcSDT5u/bljWkeiA2ArzY8NYO0drZXHPUN
jYu9wWUhHc4DC5znS2KaeZXS1ab3RsUAHD9qUgBk07qevHj90lXLzlzppC1h8HGIOyAdc83Nt9py
x2zeyDGb4w+SCQmM94D4EDJMipNisn6bOPyjN+9xfvvd7Q0CmarwjBjaFf/E3Yjcyx/m6c+lKAzh
gZaqrIuB1Tni7vwPGvovusoRxnRS6iGm6wgmx+KjdWWat6+2bjbVYj/KJ3yljdZrFOhKyxMr0/Eq
cIx0VnGIhQjneder1r0wVsCi3sS1SW8cJwuayviHAC/VRg/rcYLQrkw1GBP00LVZtjOVvNwHdwYm
yuwfkCp1lJxlRPhTKXGQDw8ikdevI2G8EjHilfo4jiUkAkum8pWqrlSvSD/tcG7+WXWKVYk80DZ5
w0waYF2aTIIkuys+oSYO1Eb0/hvSItiLuTi49ELDR71u2cNYQcMnOagukzUu0CxbGtGFGxD50wBw
Y6cUxwPM33pVw0z/MFLexVaDsClJOCDz9W/dh2bruoxmqqzwhfrN9MVV9SduURGdWorNxgLAEGww
UqhQe4zhSdv84RWSqgvHvI4pbG/pPxBdgIF3ohuqqmHP+9g8xVPgU1sw5U4LzjfmmBQoZU80h2n4
DTEkTVbzrQmS/1YkTh1HIWfLfT67EIyT9YAvl63qu8sLcNrTTB0/ETUGZryU5tEwReyIm6J7Bn8R
TiODoG3n68BRvf2wYEAqzue884AD9BVTCP3gAOkNK7m/LGXiq+IaHPXcVKMUMXWnuEIloFzSgFHP
vBwe7Voy7iklQ4WdmrK4wbbqwXAbQgS+RV/VDy3w0j28D7BKIubEVikNd/hr3vCV5rAK0TDimLqa
vNuRpoGjvTOZqk5JX4mop2P3fz9EWusLkM/HSHAD7eBGGNQRJViwdHy3VJW1WCZrmTvfjtDt+VAD
Kh8WmJYS52xxyCtijg1chl6YjjOgj/OCb/8KsXRN0wB6Ju1CRxrJVVSU1DTp9QyYXtRRIqrPumdr
yl+q69YaehZ+7Gwv1+qxNtwDwdyHLwl7A+s9oHXzGQHBsvG9HAuOhgkfg6buuEK+5lceEmseGIqp
LNDJ/iXHwvmTeUUWRzA1I/ZAe3bku6G7oz4eodOfF6tLH2qel6hZnIfW7QXofr2XwGTlS8sgm02F
hyxS6HYT9cxBY3wCcHtKFXQWpvOacO6wej+6zn1eRnwvg0q+Lai7mqVA2JBhfL+jhwfjOlj+dA1U
oX3dEO/ifoL8xiLZGBIwGX3Lx+CexA8FBekNZpNa/QPmg90DLYilry0PVUDyt2wPUiKpTSOtfbCI
SwbACkAdrpSFHNSiGSO5m2dysvLI2zXcEvsLsHEpHL9vox6rj7EZiFoAd1NjLgrYnHkbs3kFqnuD
Coe56JedwqV/K9vk1YsID3gvybHhJfgTmkZUFzLgB7OWUC56vWATMHwcQSFle8BMzdmrZ1hewJ1h
3HgI/n/ipR0QA5TGztBkdLcobj3XR3QSPaUnZu9ZvGYYrs6Uc6QkKkEn75mdbOKYfGSwlKg2o8jB
PZw19wOWM2HMsYjc4l7kGzeoLUn1oKyW+L6hjmMLRceaXSyQgq2f92//0DEbP0LWCbyMxAH6osNV
2fWadsEjkpBYJX0TY2Lo3+5eppjEO3UORI/W3RvxnegGFeYnw4Xbzl9VfFJ0aWkwsP8FhfuhQYut
6hs+9AYKtTNCFTAuQrWG7Ft56lAsTEt/cPx5id0ImzyFfF/FPopUpkhKd/u9y1xLW14sIInjk9SI
zvFq9qfEokpujSovHDBHY77k2QsO+4A0XOY2AftorBWTx0YBacPKPxZvY2/N35sT0fwyk9lXB5xQ
GN/hkdqNZ4SFBE8+2vMqjkCY7DCVBCU2fIyJ1xKsC/S3VozWnynN1LkNc25XxSl2cVWKdirWadmw
rZf2e3FREB25er3BJHiVm+KiYFyAL7YbkBGvzCyzHzroI1/uScjlBrTs8/Vr2FAMcWcbEHfqtlN6
oc5dcZ3Xj+3BaDNOynsjHMG3C0vSSc6pck6alm1x//XwNZ7d0dpP8gLJDmouEkNrTIePccU1fMXj
/aQOG+VAY2L6vqLgHo32hBIOj5fT/Sa8BJDfKSZe03HkyBkz6Xg5ZZRNASxDtr7QNziRg4GXVFVy
4tvi42i16/ovAHCtW2dYKXr38nUZNJlaeZM1u/cyoy9oDgwpS0iEZBgtWtPZCzvViD9WiD+h3IVJ
KjbaDW2x/tZRZce/0Gr6dXuCezxsevxMeLApBKt1i3SDmI9dzbVv0rfEGNrccu5JQi3bif1mH5vu
jV69c+4vgk8ub7xyjwFJGRmnIZfyzvOTXkco1bu3betSeFF+eflx1oDVJjdqqKW86CuvqpNNA5Jt
slRAxX3eWwNcnzFGW/Ahr8R6KNm589q7/Tf+GZ/zrN3pw2fUrZ5Feoxznqb2+KgwkMBABcE+SiRr
blurnQLHm+mLWYawOTeHVDJKPld5yHhLnfmEj1WxZvgNkq/1FpZuMUnVbEUzdT1FjMpoZVVh7Kfp
GQvlz8dlCIRp1vQ1BAXbTJDYgfGR1wa1ubmsFzd4spD/9g5oy7ElA8gDE+YiLhPctHk2t5Bo9uRV
aoVutbA5kVXHgsYOdx+K2MHqecZFihaHXdO39kEnoD3TuIEO95rnol6/AcC92BliFkr3zN5v2Aum
21+QLhtaHEhbMPAMkiKBB+4FQVIinEUFb+IwU22mTqbA5tKXzemMPnxoYqCx5tXoi0iAUb3afkCE
u5nwzjh1FWoe7SNlOm2RhpPwB7qTWJS9n4ywvKYjTtbxc8+zhTV7DByQRgnHJNey2/wO4sYN4nnF
q6t9s9bRId87BLespRgrIbG6VNEHJXyGov1RVYuIjA0bIPnlH8eApRLOdIFRxRUf19IxK7cSao8F
gcjRaR2rvd7WbwTrOO61j7Nm7YhZkbypKGqVuEgZx2qro1gQMqiQTum8WyBaCleIJy0zKSTDC+H2
YxxWSuAPqCNCu7LdGJXIDuFVrribxhHAMyyyu2hklF5sT9zAeRHRrgFgELsZ8C6G0oRV8VRF5Vlk
/LW5bkJR9Lmb76oQ/KFdBPeJUkPliN3g27munbc0lCC0DWnZ6+LWn9gnE5RDLe71XWmdcCLShwBZ
QiLa6VL0ywJahyZf1EQSrhvl57kdVzsxZPCeg6dbj22S+AEf2LJS0bA9q8xaeYjqryP3v5xLo5ZG
thJWDlepUbUpevid9O4J7R4Ssxn0gQIIsS7bRjNDl4AjAMr1R5yuSnxmB66UiGGb+xbs+6KljTl9
Giyr4YYKo1XBDMa+EqYq0m+JCsy6PKX/KcSokU4h63XQBErdZtuhofIlvPUcZzaoz/UsklncxLph
Y26Y9QsppLUlERTdjdUFlKoAPt3HXqqO4TCsKu02k6JUphW1QqLmL7KL8gQTLy+/4Fl2kTcAMIzX
LRGiP7OTQ7YQazW5Dxy+ujfQuCQ9245HVgBl9same16Zn6GOv2dYWkP7tG50gpkHGuQFeXYuYrdi
zUxe/MWzAY+kdBXIC+ej1aWONbxxD/aXYr9qUtFu2b89Gr3D1nT4IUQnrdIyDuRZsDQLoUkVFLEj
VDYU9xIJbIDk/Rt1RS/HWsDuFuOWLIJWaIZb0dGEjM4n1zcebCZXIfwvF4uiMUCyCOtqZC6+pBFL
c1+Rrl8D0yNQSV4imhZk5Z8PE+S6Go2aEMo/erjOrp1MwQpwnAaLSFEM0iFu7bMC+wv26S5FU1k4
8CttnWdnW3h9YmwNALMxkMOxwB9tZ0C1Y+e1B8FI53f1Y/PgWq74AfZxflT2MLKOJgoDHaSfg+gh
vR2wNjN7dVkuyJoF1CJkzbRcWF87BLPlQuZDuckvtSrGy0esHG7tGJGUbeBvHXTYkxeSs/zsDSv7
bbRVxkpNpUdjGLzATEggbpb6rGv8UkZiutJNZ5yfsKn692ZgyVfAOYUz8hM1kjVGEAW2IW2sZPAF
+QAUw2nw87bFDuIJBC/0VtJ32lybbfezyS1XuVYMO0FhfNy1xr+8vWGcKU9WTdWa4nipJq+eM0St
QZFf142yCHk2Z6Bi0BAzy+Vl/R8/dqO+r6Wgr1kCSjyV0yo/4wQeUh8YEN04eHf0CZwtVqmrxXv0
DIozVe5pW4AgzAPQcwcc3y0hB12jdDhgMc2n/IeAAb11FHo7pXbs5bl1+SBScLhEvwBF9Faqt0Hm
RPa0ll6siEcX/T/DCLLZCNOuwzxG6lTtdcUm0EFY9SNIjW2uGuYskneqx1eUJQQ90SKvPyH+1pOT
2W4sOn7OxdL4Qm7MPyDpI9hl3LgBdSXl5Hn/uRggAMw8QF/WsaFYP0T63eKzPa3EIb7TeVM2RDSH
lh0I7SG+GhyiVRzv76yWVYflDoCCFblr+mG1F5qC2RSsCOB0KLVu6Fpn63oGNCy95KB/YecKwyZO
12rBbKKcp07Nj72eVXoe+CCbOv/K1MKKXZvMIJ+QXAGYSBfJjz2YFR6Qe1yIVqE0kWVmM6rls9RN
VAU1MbO6406sPJcCVKy+bj6mq/TH5r7W7lZoy5760b36L/zmcvf3u6ydkhV1k/7HNZnlVh6Az645
LFTTvNw8vf2rYe7UOZc22vEB49Oz+BMTHhNLgGidbuWHcUYTO1+i4J4H9AQAb7RyAX+H7G8O5bM/
mXRzXWhxXPolMY3PSFO5giDHBn3PcuuBBm82QxopHfvQPjcCtmknWixC/6nj7roBAe9ylxcbELXH
jVaFCb0JQrXSsNxzZUdklczoXzutO7bom88azJTAVbCzoMwFdkrRu0zPT+Cvjqmzmly/TUQmqfNl
2tTIttCWgpzOHshH7qymAsztmcfGLxir+7JG1jNYyhnsw94wPYOHBtFTSI8s8EHccP6qk8e+LgjM
buPsGFT6Ml3M8D8YWuD6oGiMVoWmbQrrXMENVGnCaLe5eGjhaylOZ0Qg/j88a8zfvt0F5m3eg+wy
o0Of1fnPir+fLxIjrwAuGXAJHzWm208b3LCMEEs3qPh/v1/6BlCSKyW2FpdjgGIFy8oo/BjAxFXa
tmWVoqZqdyznwOw5mGqJDI/xtxWaUZgQTRsbP5A00biCDo34rg1f2qN+b7E2JbW3mOrH/+T/znZ3
hH+GSUWh8xI58YtWnZYSoCIsrZoYcurxV5vRZx22HF0lOrv0d2mQ3jVlR2md+xyiZrA9ObSfL/hz
rwIbJZ4V8TaeyihG06t1/DvtRMIC1a103MJN1JaGySWff2O+MRauCvUtQm+6Go2BWtS4P6SCUjOY
gw2DF5W+AK3ZvyUropM99dI/T4IEzI5T3APN/GaPuebNEgty4Z89op2c/PuGBbVdocKUwg98YGt4
P+psZrSe/ZWPLwRIdc7b28hRHS9M+jbtlgtIHEk2zl3WmgGblV2nMI2hpsYzXy9o9l77uSIbLZ/Z
zYASn/zBrQLbqAqmlmD9z6P28Jb7mDHGBVsX1Ta9WU/GMw+xUWN4D/eSqP3BlYVKeE85N1rSbe44
RByH2bYXIXvuZJDveSYkf9hGJpVmj5XsKL8v2t/whRY3QEPuceqNVE57czK7tAS09LxZZ/pU/ePQ
uDyQ41925ezOUZxLhby0XYDkrFZutOfv8T0+dJO+QfyuKgS65m72Ma4QqDOFE1G/X9YvuqGhKZE5
4zbB7npJ1nWBkGSnRUFOgnWX87lrNIN7OaVfM6voUVpRpJRnndOtl4PAHQnUxwe0M9j6VlzAXkSZ
58zS0QZwpCvQO2PinkOJm3PmrZfl8049CJ2jcY7wk1x0y7/BkTZYlHcTEtnnk70N6P29CwFZarmo
ecGpbI8crB/TBUy0D9wi22RZgwlem0gZa6qogKqPLacMV8K8p04gfa2kGSE56x9nwIorEExpdy05
9zI2sUEiYCyPl/xBsFBI6wOEkjJb7O1Zs3kb7Xs0pnWmXalDVIJXWFkBS6hjY7ywkO/zEH5e/BfQ
dPPgaHx/bI0HqRldan5szIvWUsIdDIHQlyPYdAKHg/Bz2UABDGm5v7Wc6qIciifp9eyUpJnw9wT6
WwyEU3uBpXJwDwuhSZ2ERieQJNyMjWUK96m4b3EhMaklxnOOeRL56hzkBmJWJemaFgM0MJcE+98u
+aTt6s7QIyTcCbEeR1rygmaaG1vpylx9wWeMPTY+Wu+nz0VkUC67y/R1XCUFfK/B8lQ46PZn9XiN
rhFm9EFn0J3mSWnpxlfhFSeWcHvDghF45NquneE/mMEkVTqtAuAXduoChZbh0hxy12hjzEAyCyZz
Phxg43O8gxyT+a+OsBuyr04mkU/dJEYQ3qc2X5PyufsGN8njI+28UvcAmjLloCKinSFdKHmnbIPh
R65qAKdAv2Lmq/LE7xmg4RNi+5rjeOlJqxSgBkj36jZJ+jp2ARze40WuuVfnr4/HwChsD+fyUWpB
4E0BPMT9emOOhnTnoGHiPb0oH/ZOPEgKdS2DnMCGH29UyQwAeob7Mdc/5144/jfglsYpQ0PuwZS6
ls0fNYrrz/ww1giY0k/dLD/QIUO5m8t8LEnhirgCusqwc22iQ/mPrMpCht+gJBsWVREhVlMSBjJW
HpJRVip+n/fguRiQXhO/xM6ll51jTIHNc4Z0gPUah/smdxYDZj5FKM3sjr6J2mp3TCsOHhSDqUUu
DX/t8V+W7vZ7R4YQae2IE5Bt1oSipDhA1UZKFG1KXyz81k8mX3JIiO3nmo1ZYx26jKExAxvqVq+m
6qXdGY/eJks3YqYrNQRuJDhZPH/fCqBoyRCcboyD3bGogSGNru4GfUXLxcXq0mZJzrdbG7aRiuyA
sd0MGDRoL35e8NCBTz42hf67pLV9JH8UdhPx8OWgQ7Z39He8c5cuYYcN5/mi3Sy2AzHRfk8WB0O+
8ZvUtDyBS0Q5WauNr1qyrkJrygc3bB8UbjQU85AyPsepxNOn8h8tqxsv7+457g4lQG+Tr+vFSB94
LcwWpNxnc2S8/y2efSSeQyhF26KUJwhJXQhlN3ye88mkRCOYjq+adDJ1WEJHq7Ulf/JHfp2z31f5
K4zEVcEj5PXxMhArGkAHOAgyC6Tq7u0nC9yuzHeS1PtOVpR0wTsPuQ8BzyH+n7NzWV0xU6PSctlC
jW4sl9wsT0r17k0fXFf953A96Ff1b1bqnCLz0uer6OBn7u7m9nppUB1lbAb55jTPRv56SoEBnmGa
ukgVE9sDzCStP6CEfd4vqPQbSHtAvuwJknDtPpc1AUU0+ebKhk3hQpYjsbcW9YLaE9oOyJV8Rl2L
vtaG7YY8rc9lseHyv/ysBeE/NpRRqjt2zsWrpi+Abc/nlD3KDQGGv9355Hzj21cHTUO5jNvQ5MOt
BPnO+I3p4D+EpLXCGvLN65EsI9rUQ4CK1ELUR/oF44EejJ+N11HarsZkQTAovr1wy2qxeaGDwCTa
QrLtVsItZMhOurrdNOugTwGGVpUcoCZLIee2GnVtvn81SRueS2NNb/rqxuppS+xb87UMbb3Zszqb
26pZUGtiC2IK88yBgUI8tjp11y3uhx5bMFZDvsAU1CgjGGksnPBL91WKec33RQ0D9oSw1q2mpiVK
odp46Sj4gqntuwdNA20MxoELpwhH2pFIoi3SJxWbDgfCMGM4mEqvgHDpuCx6RKyaWp2Qwou2RXAV
7geTIMI72hw0KPfZGg3Y9UfJOdWWu0qLDCu6z9wz+DSB7/IIWb/VPSOSaZ4oqpK4UsOk1MjFo57n
nqkkAI0Yw/PSmafpQDv9vgV/Ol6VFbsDeF1AXfE3H9h0ju5iyeM2vawTA5VDHHne+wKhM6gn1tcd
2BMsvnAazbTf2O344RT3TsXBpxIzeOic1L/vEAH0aoZ4mWr9kySrt01Rz+u5hOnHaaP14Dk7awhT
wbuozqB2mjYh8DJetgFQsaInAwp6/VoTM+MHC9EsNG/BIcPGj0pUOvwAQhk6oD9qussH0be7GipM
NNC5PMj2O18aI3oNDTYdkBPB/2ku+6qESmE54CGezyU+lPQkH9D1fdv8xK+gOSk1blLxLTF5uDmT
iBSKisaTLayk+ru8qxosb4aWG6hRAajLiEPeBmSjNStcaKFpXyiiBvjladus4MnUBl5SfSZYvBNT
x36OTC2egtFBKUe8hiU1p9Vn8Fo8zkNZkay6+gjdIHad5SnzToAyFUexaZjVAm2RiGSoR3wLOaa2
rTgGJfv0Qyauw3lsMJmf+xAYfSLF8KBUyjT3xgmkGBq0iv4wji4jJyLxcBaHExtnb+QgOdn2zDTr
PJtZ2v1xs3nlXcn+nUltfyVrWxM66Z8RmAaX5Em+BhBGgmgRGPWCHX2lCPcDmjPyYqAOrt6wONPm
mNmyv0klBIrwvKudBVNSbAlwheklv3GVJv6PwHeB8Nuct8M7sDDGTcWPyggMRXAlwVbFcmb9OtD7
SRoBe59F8ArglCyrGOES7DMCDa2I8VjxtIkNn89pkHeXUMd82AJ9L/6ub0xIASPDb9aZayTRpu9z
shKN5s2LCQ2frcjtz6QIkeLdYqOyOPFWU9O6fvcY3YIdTnKUlY/Me8B6RvRINnysssfZEQQvM+AN
l/AqttB57TxPo/3Or/ixhAB23tWVPtPS5o5EJ3vcHGEcBtC0FB+D9BzeIui8hOsBTH/gd+6jEWCz
X3W000WTOkYns5itDI0qe25SlD2LEb1229bQVtPe/aaYIC6UdrSsH3dDObr21JHiNpvB0mG/z6vW
jNa+LGGBPT9+InOv/XgERiUNKKzAkbxqyess/iFYCdty8w5QcSCjZ6lTEJ62GV/FwDw/iQw383Ac
j6D7A86ZX1Gf4Zv8EWM2WYjoZeFAPNUf6TeI1GSOo59nsOpCQ9gUSdsfEfJ0Isb+ZN3bFioCKueg
xglLS6e+EDgbBz18clp2kD3BevzZQTKsNuZeEmTodJsM4ZOsU2SJApsZ+LpMtoOBOn/+qTA8lLt0
IQBCG8SX890h+27IVZYvUVRqUmh44zwqjMPDpWktLMoI4ZQunCvVj5W1D0YfTpN6hrVTRPpO2+Ch
yvA1a0uxsUVLL4vDlID9TgHDOh5uKTAMh9nOSnaaZvaFlyRRYbd9NCUaD3GYRZbpfOgI0LYCKQ18
SndQ31QvTKJHkV40KT1fRClQ6A36knHcN7ZUYTf83clV5Z2xNM7MeyJtdwU1r0lRC9JKX2ZC5SOs
p1LRVyjalS44065rpljjoGOb16bQ72mqP1mENmONTXzwodtdV1G/WBvg4AlHKPR3+3g7QJMf27MF
dvwd7LWx7ljAW6oypcahiXkugO7lOVL9LwF14muz1IwLxJTt0R2HyuhQiuUQHJsomT1csQ38jEV+
mqODVX7tansGV2j9U4mrAiDBoL4XOzkEVxJHaE1rdo99NjbAIWGeo8cVsBQU2LlKL73/HtMK5Yd/
UarLFM7MorFWFRQJeAXcUzuTWODcaIuFCdI9kywQZDi8MdfJ9Ev5Xadp0CnRraqTZPOeC2zIl403
yuyRaxv5HlwANuRx0AnvN2dY4lXks7QjMis34ONaNZZeXsdmmmMYBDVzW1Vp8gpIqk189eh6/7cA
g3ixH4Gg8GqERkDP0K7gVR+h/QgRXsXo9S0W+ODe2izwUwXMc1GHlzItZvDeL0jzg+fcwQpLOr5Y
BGnPVEoqx98HDuHlMi1ssYAdC9KspIRQZQ46vGpja7uf0PrJpZePlMIp3po1PVXZ4aog5SfgeYts
GlTWQYP9kcKBRLDLaaCCX4NgqL4jJyU0gQEmtG5FiLIy0mqIuHiNs+PLiS8pqMbrHyU94PY9IYnw
4ErXp+ZvnOnpD7w8XW4Mr8vCtAkUwnlWimk0UZ2BqjNMQygNgM6EEquMfi9OL0tVQC7bOeuPLNiG
9ezft4YYpxuy4i1eLj875T2GRGS1ncshMSE7ejo1J5anuo7Cr192hx0huLUeTqnopM8spCIhoKIg
D/dBjJE8UBXjq/1F8L3lyTPSRr92OgCdMgnLogcOWX4cnBk60EeXXdZl3hSdQetRZU/QTsYfzHd/
t7Vi800dBop+jmzJwRnFl99/kz7cVkBDVArXx4BF+8jOUHkHLisu3FS2/HvnfIHagN+iKMzSZ8hk
qaA8kqcT/9CY7XtLcmuog6GKSUNfwMBZ2BBzk6CEMvYxcy6fii5Kz0pmuDsV1yZNRneQSW+iHBYO
Jh9IvdLonBzy7ssj9bR4eLlEl16OvxQyvx+iFdwm1FjwqhmJ33F3Jvv3zKdQ3j+g0K7+QJZL7Y3P
DHmgw9J1OAYncT1oXmZ9RN6hNsTUILPNm1oj6jRLLt5fm+mo+EiaLoj04bDX6heoyARisRV+t1UW
ZXJXcMLRR5jwNVKdxQEE5ShfH1FDKiHCepgZs04HKMOxOD1WqSeOAEA2R/ZF0KS7QxTOgajaU4CF
0gV6Mdrgug6HWiEOFcf3njh8H/KtExtYLy8e/N9BtjFAVQ8hkK0UfLRsvybx4s+Tqz23Nes7lzvk
OgXwP/DST9qCQYh1Yk9DotZ6jTktZJ9cAMpWex59GstifVn2JRML8vou01Cc+4oP/PyxZBo8Ghbu
ABMcPbiA5OXtcTRoG/5+gRuKdbY60dj+VR0/VSPq+Pzfl8bkkUZwWVi0kLMyWjLpfBSsBQRFWN+U
ODnDMKfU/Sf8kNFjU1QKDalmt4+r3Hn3jSrxFCfjYIJuvUiH9GEHHj14DqDqlL7mxksOVGiL3q7D
IGtZQPvZlRRyADmA6oBBMuoJNCayMKxLp0E1Fsw6HOhOwVd6suBiJEp69kijNO15ygY4OQc45Tkf
gu+tVxqpEbdyBWeNTs8rpBfbeZIyFQS+qt0MgMitOul2dkvZASb90rwhQlJ+ytK/xuQt00AaxwiB
CGrh+250j1YT01IKwZ8Ie2X5GUyTr1bRQUGc1Vc0+nZdtCRkmaTp1wj8xGzpFgi+GuhS29F+PjOM
QDJLiU1wv1dFt0p9DQ/JN0UQ1k8lY0NkWRRwM8XFdKClwMzX84hPFQy/wfo1iElqqHomSTKuf6h/
TDfw3lSamNw1y4PZjl0EMDuRurjsepV0Ugl6YMm4iXyPmoui+u0bCbMaBYPQGoWsIxpP6KSI5Hn8
n6/5JVuleZ+Yzm/rhbowU84tNU0PZ3JOgXoyXzY0xTz7kh0dVqLmWmAycjuBpLOLd7UtBLd2CyFA
si6ntnJZoG0kqO/d3PM5C2yFDu2nDgnoDmbA3lmUKY9qNa4TXFQBPcKJVOKVHtRkHO8eVDzZsUlw
3CVfdSfHxyKNhtlGdwGjAY1BUq/JO0+RLgX3IPWNG/XO9VzXydcYfECD2rPjkj1BdizrRVtQRq/1
eo1JFYgpjPc91kRkDxqxv+KK7UXIVLcPseubIDO/ojmaiETLkSV5wWbEAyK8t99LczsheNXTTKS+
B+UmvXb4HbRrVi+yteTAi7SLiFvok/JEXI7NSJEyDYJBOO3c0apauk6u8m4G/DNncEF7wg6jw1wh
DhwRCY5y+TLsT7e6iC8qW+qjcRV3W+hSkL2a9buWvZ7LKWbHiSMk2EaBsJP5P7yqnq9eErbYfnZm
9FYyagb9xdBTpkNQXha5pVmxkyXY0uf/U9YERu10p5ZbTUdZYSekGo2nbRgzhlfUOvVOQuZjan4x
2m+XEbLSM8XxiVaTrpZNFRq6L321P/jsiuR21qxi+9JHRJ2SRlD2V4avhPqKHaMnkFyTs96oO+uC
8v7JBGZthJraRPssaOJ0aNBdOWSExflqwGxvw9aa3Yz0OZXIn3yHz+iEwz1aHJN9otRd9e2Fm0wk
qO2ToMyc6EGEKvJOrGgUNzB94Jimq3lxhmZsWykmHupl5imrSvN4Sj9+t1XgoHVOkT9TJJVFAofH
pZN5z/vakRioLq95yubjHe9g1lnDMUqbeH8s+UXmTcs3a5Yg2InP2Hfv822sUZpjGOY+5CxTx+e3
6xu/hlRn9ZfnKLWIDJ2tSFKZe3FcWi6XiUIpYHhfu5tytQ8YhZVcqEwybYbDYKCPsl/A5W+et8Rh
vFe5OI+MASzDpZIn5P75/XE/TkNmiAl3GiDrh80XG1SSjUDDwUfXtn2+J7+NIRlNrt7Bjkeq5aRD
ytCbfks5PX111hcU5+g9CBZ8zw+4yLuD4W2jEf4UduDiceSKxnY6B+xSy4+aXCJ5MQGvsJyGtS1u
jZMnFhHqrh+hu+QPefCyZbTqM1agU3LNQVGyJ2M+zPL0hHf8xkB0MBYMPiAHyJ/M2HOMpPbcJINu
SScDDAogY8QhxMaB1H4RIPQLTY7d4U5I98s68SS+Wlvh9lC5oMhREPMmNaNOmoHZmo1kG9QUF/uv
8sQudxKD/dJzEAGSLRohWn56B8sVOdzSxBTc+g4dLHr1k/Xd3vYZ35K8J+OUWEFrFTtmdkxbyFal
firIbBWrFmJlvNtYbDvInfdAFUm6fiuFG3KnV8zb8xlq/nGlloTACV4UHaWqwLb//8G1srJ448go
573cQuxd9mGHF2lXhbZAGRFE+H0YUWwjMYvOeEkFPlVWx9vASAcTZdSMt1eCoewnF8hxtW89ikT5
V/d/raDpJWFT3QFgekuLJ5xhR4tF1HaN/KjdqJhKP3EJAA3oZF3dWmLCf7Zzhw6IXo2U3Y8vgJvn
L3m77t0h07I0b3jPINxB2PQiH87vhDy+0CzgPidDzRXQOBw217r7am1LvSV2Jkeyk7MzCUUmJ0jG
YUfhFMcZxwFk2F21BNajEw587MmBxfIDdsyajimWz2egl0x07uGw13hwrK+6Dsf2VHpvFgKNnIMN
G68KzQDyuP3hBtlTy+f2nYL8pxqNfL8KgltW4cB/tjjUDUsCWNU491h20EQsg16daevejngMwYfb
ZIZBFYEOTxIa00vCneeXo0CIUz83LXriJmuaKmrnnII1dSJx66XBAszOKBrLJZLZOUSOWnlIF4FR
XHXojFi2J2ErwoEcSsCszelpzceATKsMxy8gFaJkZ0RJrFcCaolel60u82m5QCKqfuryNZ/5u75t
znew83Boi6tW8T5H/alGw1z3tBThRlzZtyBgnbhU2gZkUDOrjEfzusfaSc88La1V8Mlo4mDaH87r
PPKjRCsdlT70Nc48jRFgHBmZvkUSrUy7a59c9vKOyuUi7eLa2HGhqdyoivCBUiWdEJHF+RYMMi8r
GDdfvBFIQKLrzZw3SM9PgzRFontYb9Ct/lZNyNrJRVlLATEz+eTeY5ov9zTiNBFvLNpgVBGZybVY
OplcL1D2AMLmFqbBBPB2jMTiIqJRY4DpiMgBArfT3kPx3HrF9vn8sAbspgdPTuuJM+1DFwLGe5ho
5m46B2O80tQ5AA1/tz+DChxTvyHWDfxbOHjxVLWivMeU8ZSuD1Y35r9jAfp/puSH4rmS3howdN/S
y7iWJEeULamf6dyk/jeNgMaHQXsiRe3VhPT+cfWZlz8EJxa+avGz5/XU3SOXFNP+f6r57fwz0oax
VPCU+5Fu9PIxxSOtIVY22TlilhNLvrZ/tZwOQthJXsdz3dnsKFrBdIsVmDwQv4cs/2qdXpV+pPbF
x+EbwFHtx/LPFb/t7v9w6i1S2FPyCMqeObriizfoTUdDGnoTkwclNTlVp33lekadb0ITj3BZsZpb
HmZIR7b4r55uj04C361A9gvnl7nbddzuCsKAWlnflEwH/HxPvx0AeQWMRBxzZMojHUjX6bBz+s8w
tQePGCAjNHRA2q/0ZsTqMwM9A57Vmkc//QiwBYyeYZY4vqEfA2OQJUyeq/xaKaU6DpINHlAgP5t6
w6TLy3OosJyZQDVU7+Ijb9lfQkRnX9q6NzWCnQUjk8Vgpvw5pasBnlrLE3VeuVpa7m7mS2RN/pfC
fFPRZBSOiSkYiFMEA3ZGKbVG0CPncDtyC4Rr9HOpyqqJ2dUFxYupP2P4JLHYJpVxOYpT23dXWFPE
rL0LDhgm0VfLkp2jbfJdBNXZtn5s9L0ABKN4CmkMsJ6fNXe+1RCLdbPu+AlqpC3Zw4rUKOG7cLmm
3IzDYG7ECLBJzfMl7yVM4Kxe9aP/bKLPXS8F5+QB3i7qhUecKg7ellvEOQUR3bdHRdlTF8dYWSfx
yzHVrO4MV6CUTGyFFeBiboSdqXQR6CAZYi9xh8o87Dyr/HC2tv2M6Ov8Z0l2SkbRPmovZlhc6i1x
ggRjYPQR5iDuncff9cQwNS/HCiqqgmvjOCR5jQiPXrvLWwJX82iZaqAaEIwa3nt82jC2eKa/qGtt
mRhPUjsg7n4Xfm/jsRNQ+3qGVymJdA0RF+kYXD6ZdIslaRmMe5DvqurQ48yiExyW0YY/UR6NOb06
Xv4Alq8mRkdyMAekO4Z3Bu/Y3klcrvz67sYzJFs8XtLelzAAMykq448boFwmbvNN6kdfJEPux7Ju
5rdklVh6YwCPJyg718qqfPcX8vPyyJ5HLz+rLPFaUmdaVJlsCFsOGXH7C1WZI7dTSq7qzQSRSgEF
FbgD4lj4Nty42H6wTgr2s2Yx9LkmDSJJf6kBhV2pwCO0qyFaQJ5s2HkxGeTpYOZOse3QjJ6HFPhV
n65BjUnzRTOo0SyEtE+RujQzVmYPfwhzoFSm1jM5NaY8+mSeFaBVs4+4wYHo2Fjg+3W3fkZln+KS
Bxz7X4ND0XJ/+Yqt8hssmA4qPYY1kaSxArJsMThFKX8oQhsaoGr+ZVUaetX8QfKzBPSwUZbVwcDc
SreaowPmRYq+QIgyH1Jftgaav96m8dA+Lawl9AFbesm6Qiww/XnzTszCOqbztiOrjgz+w288I0D3
hxx1+13j2aQg0o/AosUaHhhepYUekLlXnHfpe6obbLYZxgaFPfxBIcrI7uRUq5aT41FIzzb8OL2A
eg6RbtX2IepKk5PIeEp3NUJPkEQOOSTUliIWpzIIQmV1aIjVpYRzWXgh+vK0g+V4px2Qk6K8+Ac0
L/xOkBYU0y5SOv69uGafRln6RAcA/aIQx/Gs/Rdrwq12pdD/jlfOBWDegvRFCM41RLulI8pRfHy2
bUrTmowJUgwENt4g756/IDrvifrs0pFvS4gvYXGyd3ZlcWpZ4NFK35tJ8hnpyVsC19CMIZhCOMV/
X1/awSDcXyPWD74myHv4EtinAVvTJjNFX439DSuvmBDr81V+gxqRJd7XywDndn/IjFAA52/iMeO4
3/rAKUocpem6p2JRtVf5YKWHHU8JDk6iyWO3W3cAhEBplVLe+kgYNKAytonaYwTyPGoNBQF1tN6s
ezt2CMbvu4cJJHhvFyX7pmfYip6/mcHTlX+joBaj6bMlWmtTnrlIpf52EBdIEeC6Fk20AtDBzvbZ
q3iwao3ISYSNmbUg6iPVWlz7HCWNuiv1eQJDYQ18f1ezigD7mLjs1g2UBPpdZ8FBRPI3QFU1OYiO
etqJsR4Pcu8voeSpLqfESJU9niVhDkwzsQXljnk13YJWcZgj6T9KZTUJEhm/0gUViP8pvNjDq6Bu
BMFYc/tXQrpsOqj63VToKD3l5CbQIl3ZF/Q8ALCdbMl/1AM3L0NIcQjwiO9gZsEnzEZqR5CiX0nC
IuB8MUUCw0Y/Zq9m56CioiJcWBPqADNewB+KoepXLCgCbLvj1W9TZTzAS+m5lsBm6+zc5y1pfGM1
rYkQ6Dq4SVQztoagBSOD7PzYozITisFdgo2PeSPeRE0Wcuy+vDlRK7gKb5s5go58ul0+PQZ8Y1xS
f0nEZW8NiljI6FxGSkjROp02CQezu57LujODoSw11jr9xZRaJ9OkHMdHlYXo4zP3p3uCslNCr7oM
RgRW5TXQmCGAuGfHCsihOSKG149o30EoK3tLoHAQGAw1VWJm4EQMb1yb5tfukVfiI61gF76BygUC
nuQYx7mzCkQhugtA/F1kue0hOZ3hzSpJPnx485PQ8S9xvUD25Ku8miZNZxLJVFUAhAeDqbfvgBLN
RAQTMbq8htvloE4x4peW+ag7IvBTiuXE7tYN38qFWwfgURAj1mp+6+11nRRU7fenuDqid25usw2P
GV60OQIttLS3bQqJi1VBjobTohH45wBtVtwV2rwxi6ORf8NCeN8i8OSZr63eznFHzDtOv4YXiqTm
2g2a22YoVq2JtxrRCXIfoOLQ8P7bQ5P5q76QwCNvrgpdMM0na2KnNv8DefCRRj144QEVZnCrgPVT
9QHtvQnX2zMkDi46Vjwc7bYROWT5s53T0C1S8Ef5+LP4TFclFDvVJupCuxCRcRXn7WE29mHaoXBj
ELF+w3VZYG4hWrt/EWZ1kguOCVbOwBbBk1kPNCjhontphRcCTJFj2Bop1eaDshEjbHvw6KeeIKOR
9juKDdXW3ef1wLGY5RdcpmJmNiAwLjarn3fqQESNOAIEuYr+M1+YAGXZR18j4DrtnNX9v1lsP22j
02cx3asQcGHyznedul2wwYjo9jYlDx576grAYtBPZAWkt21NOEyNQZoZR9ej0MPab8GevL4rvrIE
FiszsexU7UMrF6S+CRxQJdwLAvrYiwefq6kHJjEjC1wG09nb+j/tWnr/gCT8j0C8wHBohqPxDD3C
Jl4s3EEZFb7x7vv7rXcMWHncvaLTu4t/vnCHY4da1J9pOApR1u02WaTxKGVp60GcPV0sUMy0N/NI
rhby7tZhvgmPlKixa00yXih6+FgnOlkFCjnzE0XGQfsr/BV420bIBen9F6KnB3DEWIXXn/4Pe0Wv
+5kJL7BoSgyuwIL/kXVhIxI/u4+sQjo7NLXTwOLbaEHN9e1f6gg7h/NkmSK0SSWqL47tGi0ZEbK/
Z2lew7xmafk8yKFhk1Tmg42dPknx4idiu2/S+0ChLu9dt1/l21UtJV6+/S74ywx0pqAs0peC0NCH
yRnNzSLQrvsLgLWIxo4ka8MwoGFDypDa0TTmoKU+0yMzIEK4oStNSyUgVS5lSFb5ODKvZCLHNbRd
M8CXLykPsjNOfK4RqGIN7w305RSRAzPesUdBJqWarQNQk+uyc5/6lzwVDS5ow7BnoeGOGl+TWlA6
vGni+TTuin2Ae79+JGgTNiT3sZrxVoz5j/MtaRTriYTKBsS8tAZprMfgLXxAOt5s46j5P53FiaF+
KBpW7LlMXZi6V9vPaDBbg4JcZ3yJwtp3aT0Icu/nW3xMVXzFaAAtHrqF0cJR3GWHm/nEygO5u61Q
zDJ1ZxMK+EmeeQHp0S1mmr1FJ/EI7aaj8ssYnnsQFnikrOp/EFlW2CbTaqgcq3+JoO2tfJxT02Gx
RRhbE7qzBAiACNGhMTfrlgYUBGR5PYvMLpOZiG7fzyakWbXT7f7p0cI0TDZAAHfZzVjT+wWX9/Oy
RdkHRjxApmAwFV0orkZceRgz4ZwbgphK2sQrICohr0hsD7RM8O/JpREPp9/FYJBhmlNRS7YYPXmI
kBksw2YSQxnZJ+H+nZfbv6xoq9V3vXrNvHszhz7g+MRayCC7K6ZkGKGi/bAeF7sOoWWFfQ1vO0fz
jovKh3liHce3elXtyDMig9uhsUdT3APuoRYmneG/oqQMHvHWO6KStdYmik29EjauM7xGqZL5m7+L
8QmTt98o253ec9moTILsezr0z4v00bNtVSih2YtjsyX3JjZVgO3SRF3xSNVwvE7M+oQ6lHZlqK/t
AkOU36zE7qVh3K/nkniVQ1JYuWs/1a64wiyaTD/+jSL+yf88w9fVoLd9mSxKXwwoXaywHJhbTzlS
s2sSTLj5jldBbj0ukBWIixwk9+fZNp7OqWVAxI8s/2jbypfwan9eZTPkzbojvI7IZoM7ej1X99fz
ALgg2AbPj6aYtBjs7nvl7HpqRJjHLvNaeIQ/syCXRZYX0/7rpZgGvhU5Hb92Y/6GIMykJHeQCfuk
n8pdCYMzEy3rSj9Vd411qWf/vrnLIGGGAMoS7bTX5LdrnwgZr7GbFRvAKcsh/7w7r882Njt6NCyt
GKBigEJG0orsPl9b3gC8T5mMnjUzs/Zoc49nOIdHZm8P77GKpdUA66sJ7HhSItzCsZPAVzAf3ctp
ikU5O979NQDl4BiYiAmlV7p2r84p9nyY+yoFoQ2p0LY3r+u8yCbxasLNR1f71VwnUfihjn187aKP
qDw5daHujfM71vFwLIlq5gn+UhovC8CitiUmcSvtG/HJ2mVD87wBuJFBV8tAWGmN6C9KmnUfsRrF
MZd4gdwDN4QoN38zeXPouzUEv8MbMsX0RWUWZ1U8wAAyXsLqDxHqg7AsQacOmvNIVpZHZvNPO4Z+
HyT6AKUjAqIh+DKTZlmZfIq8d9lcd4yBNby6gnBTnGVpVr7UiV+SkKj37DdDYztFNZBpv1af2dS6
JouVtLLu881Il2Qouy70RLKw3UTZWyBZM1ylbpVcXMhPKjjgsIiczQDwGrDGTPx4I5aAmxfRRz8N
Y6P9A8NwcgKbEhKz1OLBdRiVBFg1/o00uO4uPARtl37NVvp7AH9V3uap++n2P5IBzQtyZoOn6mEQ
9esrA4I80b8wNaC96ik880d0t4cjZvfzYIQ5equ/ge0nQbFZN4a03Zcq7v12rdM8shJp5X2x0tEJ
3KGgAGabF9Rcuhun4P23ILsteHxjCbz8RSL+U4WHqDd2BH7Rvkc/KvKSB97Mp3oTIWK6Yi09RlVg
1HI2pCqyJUS9cFAvtnAgHvuQFnkfEr3FF9NMP4x0U/8c+hul/ysfhR5jpWUvtrTVeq73fnM3/51M
lD+o7lz9VH2xjYXgxyQLJpg5/iLoADvVq9uog0cWuLr9mEw4Uqm08Ge0LjajQj1ifTtx3v5d2eWB
bqSkEeVI8E6pJ3Mr+rHHqbz36nol24Smyo9r7D2FKk19N+3NVZ3qqJT6TTqDkttjyNOxHSyc7XDK
SRZG4267i1VxmxRTIK7PU4pG3NVBIDHKLLPriRHcnFpQcYiO0x3rP8dT3r9xzpJ+11zCB84hJ5JL
3mkKeY0lHYKwtwhPxPA2xMbwzRr0a2aeV8sQKizVs3wmRev42rWw8QVX5APFbxuEZly1k7abyXNz
mhHnXGqKTodYbJWS21uG1s7GBbirux36f+rHyT6jABpCCx+h/pgpRwJUr78ach/xoXLjv0sShMWY
JEK51FOkianBqK16GoTVTLghp6Iaumya7AR1833vb2R6NGHRrgyeLcxg9F6TwEpO0XlVTUyOcy+0
GeU/o0TMnq7pQoak3QcCpXhXIepyhTf2ZtPXhV947figxjmL9ZJHe9M3JyNg7dU0CuBVw6TSO7T/
uxungmAW9ReiQivBU4zOSvUZ1wlzxMUz6r1mrXwWjRIjIULd3byCbJwHmWXI1ftW/WMY1iITdrEU
CloOTCaBYhX7U3Y6tFc2IQKIJfq9m1QTWttA70Upmpw3o6FkoMICsr2pTQ5++HI7aO7kL22EQqw0
ybVvuDegzwqq4TC6Va3VQTnR/7Y8tScKhj5fXtubKI84Z8mxgDy7svl5vknL67kaxnpm+Tzl6OWO
s9hj9x50eNkgdV2UZqUJ6EyoipLV1Gn7wmy17OpoYTYzurJn/FEzC2ciZsHvNePC3H6BVoVFH8lu
OdTp0GJ4F8pAzrF9KNgzIBM+fgO0SfvKeKY/kZixdhC7AFZG/8tF2Fw8my97yJ28M7/x3F5+X751
SoDPBGOJw9IcaNeRzPh3ZU529tmRWmWveiHDd+tPmFwGvt6qm1r8OXWe1lCOTtVrga03VHRybm3L
Ey2ThrxXDzD+fgvg3/e0K3yWyz9UUBfxfyzk6WeTCnJotxGnEcLdGmvy2m5uoeKrYtOERD7o9BQ4
6VogaPwWC5wOhW1XDVruvX9xsJVKiR4I/MyQCKNbwwc4bFSzYp3jGjLqZFnmJzLNfhAjtBTLUuSZ
RKNeYeuoNgSuIKI/YI/C0V7MjypNVo8vySZhGfeiRuh2pygFD/itx4t942YXh6p33MBW5iFO8D7C
YMys1I543HLCrkyMSC7755mWtYK+9ByRFjanvMktyEWCSG57KNuCTyKFyEnUHwhpe9ypPoyMUKFh
Mff/DKb9cUQKsbIkd49lNxnYIH7b3ib+5pNk6OA+yKsLccFyu+z7HatBT6VcxIL0/iwk8JFmpqIn
7++Q2h2hTjahDywIN6p/AfB4+s62qAWD29fqqvM9s11Mouj6Cnc9OVYkySu8jhyWkhaheNQa1a8s
CrYmGff94N6GS0tWIMS8FKnCuJCQ10h/+Q4N6eZ738rCw9yul9aeSKzBgz8DxOLXF9lpn3iHki42
Ox/xsmVC1HtA8zs4DKZTxOl0bRnJtELKObmShAYtaDgiwIiQ1wMj8PeQ4KSAHB3urL4SYuLOKUO6
sOTNV/hRLybw14DwT3uYcND5ifTEMT0PFSJpx7HKHpIzBB0QG4lu4JZAdpnaCNdiG54A0h3jVH7f
DWd+iTGkXIjwtyVB01KWUCFW1Ps8DxqPht43zY3PReuukx/UI9ql+xU50qy8Tvy90nUwWCr6jkbh
4Vw91EgtfRhmB9mtECIBmT7YUeq+0EjVAI5rqex2kcsAtKtVqXdYzZH3D8Ee4T4B8Df+cD0FWzSN
r4P2NgH8LD19GQVqytCDiYG+TwkPNpOThI7fPRfL6LvdspLGqXgFeYiY64yhBmKk5rrl/jHs0PsN
h4+83GzC18Su5TsMWBkN+Fb6vWVTDVf73Hw+Nrilw16GQMTo29BIsAMpu/WDDXwgvfshzQOhlnid
RUJdCGNXxLBLLd4mwMjIpWy/5f3qOtWlWeJOOyMTL7jhdNu6qdocEzyLr1ktWbgfX755x91dXF9W
X4i++AnIf3ImVbHVqRAyjTLqchlxqtTBNCm0D6T01xjnq5E4Re37cRcSUz1jwHzEZbIir5KsB/3H
Cvrxrlqi9+JeGBltyeGe0HbohKqftUErrA6bjP1KqWpgpkaKdFFtmgbBtgxt0AckLOZlsWPHAfFB
9TewPOk6Alhj3beKeIWXZvg+HaP4iOwCxrnwUKR6/2wviB54ArKxVTbV9wLgSbm8EytVhieP1H1h
G00Djpj5EXMbHQs1YpTN7GQhcwnmqE2Lf15ZH+RpM24ONWRuN/Pp+Nov4vYP8nBoh8L/zTNoxiD/
cWMHR7xNNNMeHW5y8LXQn7FW2sb2yVOqZMYVtCC/zEDfv7kWEc+nFlxBJRlfC/qRA5kPLfHrzJE2
GmtqJFyKSUyH9+FJ1YzZSvJ91zaBfxozFcmdwa3+bdAccpWKS0WEKyfvOL9IadqNEWmrAgmWp01Y
QfI6aJ6zDYr+E4ymVg5+mQuQAYYbO458+WlCKZinw/+j19ZLbL6+jpfGWgircBZ628LHBGTh719G
X4+5/Aeh/CwrC7bBrE/dXA1ZrXEt6lvYSPh2gJ7/LRXyzPber+FuQojN/dCkn5hep4MOt8xOXzKF
M+uK5PnzcuiBKNB7BUJ55tHoV/HPDB8fWEy9T1kmv0icZQS+5B/FtHzbmd92nOiZb+fE/M6e03LQ
sqPG3h34P84eJJmsC2cWB311NH21qwP480xAtl/bcy5J1xwp4+eXErmcKcg1ADG4YcGqm4IAQmWY
+xLEvaKbZzKGvM/iNcyX9n8ClX3rB8Vo2tLBsVg2Hnde9HiRDelBwBCiXGttD27MRxslLI1X3oLY
QVj6M9qBq4EGh9HO67jY3axBlps+ChOnt3zuZFiF9SKRw5zRTXsztGfGOPg1tcZ4rJ4AueVWyyKu
Hny96YR0Rc5kF3zfXxZV7uqABsCmFFhKz4QNPa6ctcKPGmW2j0rP5eQFPYKtGszDjr6R6YJfXmVX
H5rTc8uHdhzYXZ113SoovHeDoCvmU6MHAq3c95u5E/vT2y+7pKnYuBci3I5N/2WjjvJDf01x+VEQ
nJyNClzJTp10M16mTOX/KZRWlNSkGbqyr813P1S0+3ntaQ7fCXpdblH7k8ts2ZiF8Pp4wsKKVX9+
V7rL2IeJsTRdktO2hZPqVM28T+el9rxTGZdsWGE3PxfQEgcwlLY7x45eta4jJQjJTI/SSs/Cx3IP
JBzFeDLhKew5GfHnslTRpd8zan92maQQ9W3mQgST2lw44OMV/dUuWv+KBvq+U896an7fmoRL4Akh
Adkq9EG37v7YRGiR5Rr4nAR4NXislRrMJeqDd0Bfxr3LucuyMPhAURew/VUnrZCidpk+H1G65aRU
ozcryDVvbKM09NcedtG+xJ82RUTXwiPG3Hmp8Hv6ES09rBnLZaYm3DZmRWLqkaFKgQXPS1GZau/H
GMT3RdL2NPLmlJMe5Bx4V2QQQ/pknPDQzqIJ73/jPA1X8dc9ttmqJXePRB26PMsILyJEsLpaTyF2
JYV0WuNofHpoEcmf7w7YbjmAeHhLykEdZ7rEHUDcaGlzn76AKhi9DBgQeeXfpyOngTWmwAFug5+K
Izhao38ym16aghlaOjzVvF3OTEKh+osJiJ9cvcTcZrQe7SN6LzCyTw7apP1miWcclZqxOk7hVwzU
sEhFT3JB0H2ETrWvSuU1dEtwKCCpwCsqnIwa7XvnBlYW45Fd97CnLOd4bBo4o9Z2K3hJXua6XEYe
LvJ+Ny7ImKe3f6nBEaasTx9KYx3z7Ezpd/YDikrrxQ6Bl0FhTUSVugmBXHwOMHY93SX8DtkuMzrY
/FNAK1Kp9u23j+HJCzr/f+rqargF6c1S/LRYpX635BN6pjnpI2GJxSBu5VRjW3peE4UV9zlCZ0sq
7qGgySHraoU6wAD5sVkXta0ITnTy+mkhqSJJIYvZVW8wFeIVEojCXmF/+z0/Uz0HPyeFP/OE9NwD
wQ3hY2iEcItWDS5JIRtaEVh+0GBu+w7hOm9OMw2iZJ5BRpQZq5ossi/4ZFPz6YDNaKh541yVTEpz
bQRCqIRz0smYixvr+lRLcp9bXXsGcGw7tW9aJ0tH6rHfSNt5NgejMKKTqI+LKX0F6AosGlBnLGcz
i2Y9eWG5zAC83BJhxJj8qry9D6Y90K6pWZpYcoL0IIUU72vqbMWzylMYX9rEvF8Gk6TJsVxFI2Cq
KvkHYEINYUDldxp34IbZzMrLNfHT0K5Lml8TGQDChRWV7svuPDL5fbruHdEsK0SmOrCw/oU4ZaPs
hLBYXDws91xy9vGftrfWK7ZiupETURcketmrKrDcnlQw02sGaILBBV19XiTL+aiB5kZSkTSimvXL
rjVUg6nlJ9WBOH0bV/7DCw4pe1fz0Wa/yI95hdApbYLLyi24/aacNVmlNLxsHP/e2XgQ1T2QhRce
eVEO+hRB3jI/v9cGPxQRHyK1r/TrUNkoOwmE/uPaMRQdPpMle/84AbT5eA40nBNk1s7JtozCUwE5
XQfXZ8mA7+FdlH5qHrDSehfeQtfFK742/+gNoWBCjkCekABNRhb2I/yszU9StDjbtXf7eXt2lzdn
fpQEMQe3ET7puozWIIULkpC1doD+4eHnPCRuMdRjumXl9Vs/xRVyphD6SxhbuI7O8C4eDhYLg76J
DN1kMCCUMuDz4Iv4fMRYWcQF6aKrggzv8BwSmdbRAmrzpTNJCMUJC0JLKKuNe0MQC62TJIiUPttZ
SQKWtVGmIzGejT/htXL+SnPeHGwWsutc9TZfa8by0pt5DCmFGOV9XIqDWmGCMWvZQ/xL5GlLPyv1
eVYIS2sRf4CpNKqxCRNOBKz0UZ1OP784tU/2HrnS2XO0ETtl5Wqtdu6tO2zvgZ+UCq2MNS/xqYjs
OqUIV8IjZjSEQ++jDWirF/NiDbziURHV6ay9NUaTgbhjaYtEHoyyn+7WTlv24eWzdZbma2XpVpcu
B7OCu5UCziR9onWLsrYQtiWwBGl+ai+WqtHDo/UPo4DsjM8TX0mPLH4mBteGNf/aSWIkc2Ls1jle
isMTbCHcvcIyg7hOnkjxmd3zE/zS+u3up6PFxj8qru3oH6sXpAvj+tXdyLCxb32cq35WAwE9rqV1
8K+IGiz/iBkVWT1K7Q0cQ9xHLdINhC7461k0YsdXpusxFZsMJ/Ytrk0US+SiXEnk1ed4NMGlNXD/
dJueqgwAUIn3bP9gszbVEiAMfKsU1qjiLLJH4uLTtXVH//woinl9Ccy5T8wWDTGiZltyNkfQaVMz
dE7vrjDCZXzq/stNYkwxjKrZWIMBArEykqmVLFKeLi74L13Mrtj8E3Srn83F663T29R+l3GWTX5w
d/SK0VhgmpRST2pRukSQSKF3jwvK8p9ACsY/kc0JV8oQUF0LZJPy11CDahhEPo1Bx7+BhGswnO4T
UnuAXVcpWwwQzpuLd4xM0amMT3tMihHCNwv4Y1pkx4v32gZU9cgwuzVR+oZsgjjZcv0ZrBp1bzMj
n23XUfnsHibwTSG0ff94wXsh9YS1plmZX9o0ehcCcUwQWRAV/p87mA2MNii0+eFbaMOg1Hb6h9uV
4RDoY8TQYiMFQx54aIwPVct1e5tF1bM7DBTGEwncUpMVdzr0rmUi44FD4WapgNtbcNQBDJvDx3ec
ETGd3QlMm4IayLYpgU55CqdbAw07jVNOXSwxesoLHPVxE9Ydj4Z103qGku4cQsbfJ/w9vzOaenZT
QzYXVAWEytedzeytUXvjcOVymsBPxhufE7timBOik1UW8p0ZTcG1PPV6JsYc22ez9lgruHYi+1S2
LQCvLrUbp6trYYqOhU6Fv/A3v++yKxhkb3H7+lB04naDhcxOCGrFTSBzCkGoRtGvTpIJXYTSD1D+
r+AGzjfnPHzCmHDM5kc1v9IXAKo1bEZdDaZp6EmkYiWicC6MRf7N2FA6atUNZNXQSyK8vqxRoNxg
lxslYNhdA/ApxuO/7dRSIMouHlXpc2dwubONKMZjDwjlPNRfk92Toosf12LiaWb+E5bZD+dguGrv
o2i4QOc/ysqxbURonc8mR1/UzdJGaTSEuuGbgWseN+bTxpoQUmhEcIS/dlzKpyOIV7dBrVjJrH1D
1j+vo0B/AFQZnEMCDZyvCR39SRbImiRcvECstQ34xyO/rqOZmblda+z9CZ/77QSYPCzLVx222wTa
KBDh3qvs5CAzgDryVnb1iVLMjow5/766+LAlHHSXXAxXnTe2GX1w6dngllZ/rjvo65IDyzDLE3ey
iksFgjCiDC//+V8yWMcWW507KaONyOlc+Q1VAzHRWh1H7uAbvnEEWT9B8N//q8m9wNgq8ir5s1fD
SF8eYrkxGoIssRPSlOfzRCNG1FmOAescEhlSj9sw4sRQkXePm/V7Jvf4onUDVeioGrWnMlqg+Kdh
+rCAxVWqCHqe3Ij6b1FXHpU3op0zlJMUyut3SBNiEU4UjWanTKvaWfw1anMm8O32aSqs1bjgxGCQ
Hng/6JlVPF4b4Fc4b3uLaGo+QjfgtB6HwLr1e7mFvrhQjmz1/4NS1VVdILtqOC8cB+mAg+0jh8a4
DYvE8E/NiNDmJn97WLJKisGUFusA1RBlv7/6BIPvRYTy+cSx1/Df74IUcDXPQNr/oWY22LetDGgC
TcDv7A+dAP2sxCpszwgrkAEI/MeZRe3rZyyQtaDmZ+RfL0OslOJebEeqPX70h8argrUxkL04JB3H
X32wJZNMjuAW1K1a80EfDWJqlfiljFEr1QbjAoO/5+9ohKlJpmU2AU3T3hSY5ct6qtq8oSMsVwZm
tblMnhB7L+UDo6d9Pfx2plmBFcuqgHs0bmFZWl0xLzwERH9D8ry8ILg8Coux3GogreT4Y/GriYNq
8QeV+HRojt77mVHEbqilko1f4DOwO4UfmHp4V+W+9dfpbLhemBiv0PTrDTx23zd99YRn9MWVN0UD
Fr4ZaeZUFAWZiP6SA6YvyK3+N4QPuWyA8yFdxTjSEZ8W3gzcDDZ3/tUN3KotqG4UqLf//jDhweaM
zQ0hSNdcc+3LxPIDNohDoEvYxEKPzBl95VG/p98BbodUtDtFx+NcWOmnbokezSRkAnfNfl706s7J
shM8IhhNVjxCn4/nX670Pl3vHMTICLJp0K9hj7+iw12q4IICzMqrlg0SqWmUpp5FiNhXh0v/rcxh
8pJS48kH67fVMT3V518dN0qd71PS5cvwzmSmbdFoBxV4o1qDAxeA3wiLtms9m+Dr8bxg0uw1Y1rR
cdOaZSTM2u5uwzkgMNmkiFBuMbGNoRgP2HkBrqHhiCbcTga25Sgw7b97UbBSGb5sMgAFrSgcEAFo
EsvLWnanav0ktzUSrdGU+K+IJ5tqq4lyKck0eX/X8nRvnUDiSXAe9HnU6Odj9viS6HEznIZp6E5m
BQQkywwhr66havL3HKPgtBUWLp63nF+UlKVoOUI/lKvk/FThJrthB0EN88QRm84IkBaU89kX3efU
ncm6+8A3+8urvkaFcDOW2+ekN6WnbpbfWVACM+cRDQlSHUioRW8CZ0/Bjn8nxauCLIRIVlV8L7Mf
6SrSIpDoS5/5bwiJPCKf6GmTywP88hSBW+WJPVXK0xJ/O2cL3+kpNCtHcK7/mK3m4nFVJYLB6WD8
zz4yFWgtFhtj/gq9Pl3/BhkhIzBrJe07g60t5yG3T1gUHd/kZhO6SGDZpVp0jj+4w7kP3+AaNr/p
YtpWqV6RstI0iSDfVdj2Td6jkQ8lz7taKBVpCxO2UWusCDADEyZDjHaCEpi5NyBEKdpHR4y/yuGe
yzVOH/oeh4udAhSQRPqJ1IXKmiR1qj9f+jqlWXIDjwUj5eW89eUgKf9IVHEfIf9QNhsDKaVlioqU
r/XoE1yGxHBoZ5VpnqhAqSdfb9n8YT0AYfCBmk9582BmaeOOsKTdsdmPDdMRthtpueEmWcPFkELe
QT+8pKQ2vRquxfTrJWqYhhH3aDVOrk4/10LaSqlearX2DZQBWpTmoBTO9qU1dOtc3ScK+tsGNY2+
IiHGKHeBCOR3pV+E0m9vmHke4HlDUlwu38WXQ7U8ZzD2WRlpufGiabRlMFrgE1oAJTRENvNFFF2r
uxbskrJ6QxQtK4hE0AQ7LLJXzlHnxJ0Dg3XiYr+01U53jYzOYyOIjwT2q75rkHRTbTSPKREzQHm4
DhhqoIVUHbTswQNZkuD6a56S4ofqS7VcS2FzNTGxxKlBo/PENf6O8YXZ+mIi0GNdKLNepJZLxOTJ
nsZY3A4rOI1OCLuIIMIqQmR2DUbYWMLjFJjfIvEaQNw+u2dlM9wi5E77pda79T2QQXOshr8ZMj2d
mHDsS5iVHPim6OUw3FZlNEz9yOwLSbDUw3f3NeebLL1yUbrCqOT5vkAS+fd13XoEOmSoKouGPu8f
4GcG9u91SGvcYaWEMAqGbiVwCENHVdw3NE2m5o18lw0sVn9m4yhl4sizudtTyyKd4xDKWkKz3mxB
mO9RPxA3uLL0i3SxldZ83odzDHtJgQNeZsTWJ7DU5m6naDScWDKNG8Hxr3fcpKRk72l9NyU+Eg3u
pTkZ0qiI5Rc1uJ4NzRoJxIjE1eH9OJSOOjEaeEnh3wmHRBqLLLRhIj5q0GFGWsU7rprDHmcs8LFE
cH9eQ00Bs+P5AMc8XwLLPZx39iTbERhzF9/INK60V+XxNizgD26AyeIOFcFho6BdrYkIcgTnkej1
nVY2Wig+OZnUNq553rIeZ+1DdxoKlxHSe95Psh/j4vFwrDg8CbCpnhli4C2angoEDR3IXF71AwDi
TZz+o+JIEfCVhrkqRY3aU5Sdserw9ETVMwlBZEMG84JeWDVnpeRY9bs2Yj8Z8oi/i/B2z7t4QFnf
HYTBwp3PcfkH8zj+ME6K32wLcIHQTsA5DVMK0Ok/Wi67lwqq6hLquMNtRvuK4/XLs9q2WyQyNNWC
t0FwHwydHFWMIAV36Wcsa/nNhJd02FtUIZcrLRjHOKaVpAZnhOsEqjn+zG1S6XdJxYk54CMfQRvj
jry3gdCNH/TnjNMv4JtgwfSIkbETY1iODusuO/5g/n31Eaa4qmmzlj57qd9NRFhm9L06SdcngvEm
9pVmqIrld57eYdBBu3zxUcaClYZq8gIFUkGM14WzRQ04Ozuc/vtduXDc1ze82y7E17q30ZodBLea
ogcNlxsh18Xe8gZM34tUIvxMkBjL1Szrn6Qm3wpYhRTyPbFgWrM+OWLc2uKBrXwe81nAdDCPt8QH
mAlyPwMvNZYbHG1UKR/EHY9oEN0GRcZKYduJqpTWMFzh11zuFhkHzwCBuzBBW4ay1xI/mpdWLrw/
TzC4dMf63ewVE48CzCyVzuf0uE8MRhTL+wHyHSBQUBF9yTSmgscVS9EZaOzNCBdt2uCsVi2bEHOV
9DK3wjyCT1MgZXKwyf3npOlN16Yys965bpHN+Dbua9C3HvYH71kvW3DtrU3I1F6OnMFfNBBnBxjR
GTOULpl9k2hXlsgPACObEMau2kzh/fg88bRTSIgY9VEFS2B0ycvhbVr3z1iLJ4thq5hLs+QY9cB7
C3i9Ocqu7C9Ob6tAU5ET8q3NC7wdkopDQZY46EQ2+S4Tlhjul9YZe0ucCSYNE5rjKxWxNpcB4nQY
9AGWACpUQxEKTwTBpVrgwdBFURQdTLjvxPpwpUlZ60Qrm1hRqW4pfw/lqfjgq+/8D1nEt3LIf60y
v0l7FCQ0Wfa3GDlZ3+5lOGTCxGEfsSWc6b8Gu4hxpMH2dDfiSjZ1mpUqQVkK4bmNZev/vw2sD6L/
1V0986R7AoPMCBd71O2TRkHFv9mQgadXRvq8HPX8H8ktKjCrGsC7QJqEtBJNcMI7+GGiAWd1aOXq
xQuzDJFCNGyAqzgv8qWHdZfyPjBD1TevmcRPtHuUxh9JlE9E5OQ4SZ4PBYY9DxFeV0qpB987XcQf
QqBLRrhRPpiE6Q2ANP765LFReGm14v6fZIYR0tbt/HQ8jZ0bAe1Blk9rnTbb9AYsxwU1LTr3DM+P
atzjawtfEVsjkv4EOgP8Pgp13HiFYT2g9+F8WndNMUkEgfBFTgjWg7oU4Qy5usn6yJ7W4iTEbtrq
s1RqN6TB+dGC2zolrloGfEfAmTQbWzj+gNkWzG2lmDLo1zzcgInQbnXF0rU8nC9X5/uUux6DU2Rz
OZejvho1DiJxMkLwcFhsNFEAK3LcXf620mdG4F6OjwMOTxganuBpp5SdsDV7YywasroxgxgBLE1Q
78CRQpK9qexNVweAcvMnn04GStYLAbgv8f7KE7BqXE3Sqp9kZhn7tjVCbomOQWYk1lN5NWUclCQr
zs27OPIkI67D37j3qJMBT0TVlNqg2qvW5g26V/HrhMO6cSAGOtRmsEE1K6qkAyn1azTBkt4pBBYz
e1mTX0coQMVAS7LH6KaHh1NTqKONErJtCLXZFf7lRKQXk6m+4yHTVsjjH44APeR6a+cRlsFL659Q
suiTwZfIWwcdf/OEwzRxwD0bIoeV/Wn/HWfNkgaoVbWkwffuuTSyuyq/0/R237whnUSEFuwLqFpi
fjLW+31q1DobcJGrrhZyRs6ohPZ1WNVmyvcdbzcidB41p3oiagN/ggesu1v5t1Z8J60banOFX/eX
Pi/+iKaUSsJCZG0eIcPvy+ea0y9qWeyo9YokMBqdB4fprPt+gL8NtjW4E4dkDEyJqKUUBN5mMt73
5xY+mIWQJ4b3dqMV9UmKOQTqJPT5wUdqjiyy/7VelKaNHeiXuHZFUMGn4cGMGSfdeq1cva+dt6Py
WNlWD7cDHF/7a8DUwPlbd9xiAHTI4Dxm6qpjNnS8QH0nNJ+PTpdT1lM60fejXbyLelT1pR042cs1
ItmgRa69OjbWI0vnQQyKZ+J2ZshlL3uEvLSNE6iwLYu5CQtl5tiC6qXezdNxi6MAQy0m9Mm9PDY5
qE1ECuyGhiOkofALZ/XQZr6+p5bRc2JWU2ecKGaccrd6mSzSpGupQsXM2qAjyTNpLq9uLwjn0+7t
23OD7ouFGeZGGIWgnI1xUfMxUUhIqM5QGFd2j7k4meDSKkdWs+hYtuT1ek7FYI0VEERiNAcbwkPj
GUPjce8TF5b3Jnd4lwu73MvdQJUesHRPb/TwgVp46KUTDouPhnmI1ldylSr+9XKMhBx4958p170A
PWM7lblMD2KBrEzrUts7KGf8S9AgbZd5UHIic4gcfb3dDTx/ZhR22B/N7Ndar1rzLfrrGzVHXacI
Ju2/ak1ZnknPTWaJiiPFTfI6PDDjWJpvq2Hltton9+FGTN3eaI9N4C8uYrqFzPRfvR3oyazf8GNm
kgFyPzhJQIiVOvWViNACfUGiafzdRLQm7Ie4VnGAGsD7v2O2IskJJh1CP3SEdBtcAY8SQI+GEHi9
NK3uylglodLPKhLsazuLL/bibby8WDHOasIHcxto1JRdbwFHhsZFYpuFq+srxACFQlJZB3p9jv6B
NAfWEpwPAInBX8hqzSZwjVEIwN59iiskiTryJ0ht0SN0tBsxMpXXGyGKqH/0fIoEAhTAPwpmWrmf
zzoNIt5fST8RA5nfhzSfpYo+z+M8I4kRL5TQ3qZFUn6BWq4rcHgqnyxqroUqSeDLx8rhPGR9cEhV
wKoGwr39zuQdoqyANAFqJZB59zH3HohgSdNH5m/dB5UGkgwyVwTpO2G6sq2iCV3hLrx4C0Fhb8Bw
/V3mUx5xCpKiKaQWa8aqAC36b1deiqhFUIj8Zf7YIBVi2NAspKyztfIXkRMkkfczg02XxQhHdG6m
wBtDAHXm//lmADSs4lAGDjlNrqgas6wiGjeiUXxuUMPAq7Ti1S0KIAehERju5mb1xo0Ma3Z2K9Tp
MIabWqd+e6est/wsWMg3ytPCcftwMjDu7uY/nTLV1yj8milrjj8QLEwqmf96/8SVWg0l+O7Gk4OB
A5+reuN6/2f5UUn5p1EK82tCimS8OSp2wJCToTFv2o3YtHUExaw6eHr+It7vQy5oNwnhlY4RevbJ
/Z3IsukXAQvCpfTW1kkMzgL3CY6i2V8ALZ2Pux+YtLweSJkpOER+kTr3m9j7psNpH2hBuxoqGidn
00Ce1RnqebGXj+7Ez/KaipuBbay2YdSvzmpDBWoOg4v0TWvRKUEJnFppKNmCKi3wFdMSc5zLKlPy
359DPS18aYKnYCDHbu0T8SdQk6Id0/4vPg0tIfjZMzZITiTWY3xZyjysKNo7khZO3enB0rkwrEFa
wiFqZ6eV0FnDzs2/mMsm9DBgicBi0pXGyU8DQC0AA8vtD4n7BKu3MQRMnfAzCnU/DrDw+wOqt1Hb
RYLGd7pOqL7Z5jL4twXR6D5STEahqOAITJomhpi27rILckRHtxllD56CrWuqsEdLtIyxZu/PYy6p
q5wQsy2dV1LLoc5UtM40xnfzKYi/L7r1hm2FRPXzULZoTH6et0zULqdQ+ce+D84WorggQUuLx4Yg
yqC7NZ0Y4YeKKBlH4uCWs353JZxkrXq/l085kzMuES2ufsfgUURBFXzc8MFRrRF720l0b/5sApBG
WH8EQQDJqrfRCmp6f9ztQoJuPtcO1xXYc3L4fdp8dvRgHKnfluBscwRBqTIhE/+vzg2+GcKLoOXZ
SQ7mJw2hjJRRhRPW3C3V1muFxuzpgBTD9UjDqkruugRoDzha9NDiHYBEpaZamIfnTsxz/k5u4vog
GVTcRq5u6CLCJOF4gNum4UVcvJJkgPgBHnDB9SF7tLsK8gTcsuYeCDYVlYGvwi4biREIB0U2tuBy
5Ju9K3OV/yrg/Oz9XVNAmv3SGkGIYHDJkxq2MjbQNIp7Lp1NjclK+RaKqn0pnM4ct7mv3PKmKW2Q
Gmduw4Ui0oOv1XiJ5FLfFqr84YG/VCm+qS5TgmvUHMgtbEPr+udRk3HXHkbq+1flJWTPYFGAgdAU
5qljvA2q9TuFOk/gVBclrFuzcZsd/ZWnEoYex8vvnteR9G78fjEV8CXf1yE5OJA25BEI6wmOv//7
2YQoEBIQWY/+BxVFZ5G1cV1osAX1hwsq7EwBKRBJ9kD2qrVI92lR0Pn/kGrcLml2r6olxceGuFrm
VtATgOwM9zdNsejBvUWrRPIGYiIbymXUWW8ZFjSkP6kJODOWNuUrkZiL2YfQTp6STAqGaLiK67kl
aTwmf/VraGiUFXOsTYsmH2I5fPzIR5/7z+dKMSXuqIXV6fGe+U0aBQZtYRdqY6/7Q9juzlxp/+PK
CsXMYu6qZRoyl11ds+KBTYHKfcQbtbxQ1T/W/grZDIhQBRerSZMaPk1fSbyHqYAkOvH5N/FEr7gD
ah8C14Y20HwOlHyH9Hx/NNxsh79U/wrRjsmBIxaxuMo+3T7kM1Pwzvn4mfCROItGR6LjfrVOgBY+
iLrJvg7fZbeB5ihRo40X7Jp1rv1QLJqNiHJlDgkmmsazR1xj7IV3pF7hwz87IHo68lfmRQrFrp6g
mX217emENqvxLkXc6NQxsoERwrq/GSwhoID/6RZwZVFfmJWKl4rQPU4l2AqvMQdUOJPtjoz9Zixk
v36J8kW9J63aVqdRTIUMp0a4S99Kes8lfw3Yy2M3A2gPHT+fJV3Rax3qzGJ8hcV2lNDOZcSHiDDi
+BPsljWnY70YGr4+GITDFjckgO31ivoYEiZKAsPz/xTtU+2fhhKJQV230gSWhVHORyzrwGm97d57
/yXaWhThtAwRnE3CBU+21YVscFyqh3XJngl2+2+6GrHbADPDuyZWpEUUZFydb81kjIdrY89O74xb
o6gwBEpZqwSAwDi1obw6y2lLIBYi3P9fp1kKPCjd9r6OD2sYx7lItUi6Tmmrmn0twGtV9s8YkuW3
0BSSmt6f+3llRtCzzdHHWNhfQIXlTmrR9+0WRe3//MyRwMq36fRrN+WblGVpwbqc44swF+Q0TY9w
rZ9ParcmdJdwewZqvHxqv5lLc5iQtthhx4o1k7npPJjOGufrr3YeAfHl6LOuO7Frcjm0A2S7hgI2
dK9M4L70tH+O9fWDWfj0xjyFal8xboKAMV+MGiYN7i0/QsuIkbdSBZygp2v+wgbTR7F6JyLjue+e
fYPo5CvSwASgjXDPudyHBrP4YqPkzfF5BMv8OzsJukBC4fGN/fvIw0weDSQMAthDurQj7bHXPj+9
2BVJvzzqmAfaF8f6WW4W5tdXJAoMkEaQbDhqE4LMFKgEyo6R4JojJMZ0g9BiIkfMDGsgMuu3yMkE
o5qdeX1lH3sGE0bC/49sSqgG7b3Sk5LORXMR4hcn8ElMuUWT70Y0v9Q2KeDDsQKUTbyHDg0FffKx
XBfLTfWcmU1sYNc5+WPR4dT2kEdXowbT9WYUj7IrrgvsDAIHqkk3LDWyKebm5mOjxfG0eer1FrHT
vwLS3HDOMTUO/AKXmGom6kgMTyqd0FM6KUoW2xnifKQMuO2MG6tinQzT7H5aH5kN+zpre//94E7n
1QHfR7TXK1H3/BUpkHDwhSE+EA9TD8jWuPr2IQX7UcDdm4wYQoopqL80SZE8pP4YedH6nAixiCYe
ziHuWYe6G20HpgAN4WnU1bwHQjm1Us4n0V/Dsu3xHJrypQyua5baMFoQpjLskWw1bDFzBqV6ax/t
PQs7oReiXrqNusx4CKDuxmeZ1nsX/ZIFie1w0ZEfNdO/HqrLbJu7P6NMVy1vy6h4cIBhumxPAkQR
HeoLUHWMM29myVBIwaspCxaZHboyIiBN0XKHF/0DzztQ/9BMQFBCzDZjlMm8BMbYIIzt7bEXaUxi
8lK6YbGrH1MazeWobA55OiV3b/DljRxcf5Ocp2Spaytb3m5Sz1YX1f+Bkzfc8l9ktiJaNb4BQy6L
QwdrBV46a92zyubkGpbF93Tfwi7iT6RT8JbJ62gxM5JjqOVxd4heuowfwj1PuuS3q2QXyFdJlaFJ
tUrPUIMHQjhHQf8xYVmz87YV4s+CjYApImY2P7xH4WNj8zXLld0LKnXEpddhx/Ju/wAh3DfkUFdv
Ej4X/AdIqsZNbqWFqI9Y1rWgr65oMBbYaQzlk2jsd0FKyK8HC+osztFhvFfR3lOkZfmrVPIEWx+K
2Hnm0laZwaImzrF4JKN5zpNE4wQF7LMZ/dW5ys9fzQUG6t4KK1cin7+9OGm2BfE7lP1RK2bzMZIV
Aq8np1vv8kFxhUXL4/zX65+FtaI+jjhK4YaWD4nwpvR2XxUP1Y6O8tm9OpVgSGsPFT2XFPKPkELW
jSD803xpTl/U2OZ3kcsH2I5MxAFSRDBEHHNsOuK0z7n6d5zKayDK6EL6OJXJexgG5DpVkeoFbBtF
KktqNdqT/7myzq/J0ORd5sJpDMueLGMjiOGWhFNXjgxICNlBd8Y9G/R5VIE5JzaHoM/nKgyioyz0
05aNeN0lAtPGsty0yzind8mlHVACh/QBrmzk2kUv2mt9QEwxhc52HAmREGmMardbxVFaDx3rywF/
eQaYTpm/Hd/+97Y0F8ofm9TXP2n+0XLQ47aQy17LvoR8agLL3+3TGJ92A8lT7SLG9psX7O3W30d5
yhWoZIjQKjeTNLOZbIB5VG86xgSCvgFYtTJ4d7yBhSXz6gS6n21siiq1ADReyPdnj7EELXo3Gir3
+kzOnCBllKyaCSEae7U0XcQb9Qs0tbhRYDueQw9tEbyPBj4RcFbsJIFNTomDtrbVjlIeLjEy6DJM
yM3u3brXPhlYM1kmb1IzzBYrOBBDlyu6dKXS327eVa8/tY48mwb+tU+RpVif7g3UAFEF6jPgsNhy
7E8BQDfWi1emAXxrbNIzAUuI0wBddt7lAFZGekNRtzCq3axEqKAUvq3y8ExaJT+JN0XqjUtm52rH
PTzMMR1R/BJBHUa5I4yyLlZUUl4Oj2J6h2OMaxiJCqtmzjSelo2lproRMJHNdpxC/rL4g6aLZI6O
NW2ENwQYNMSYboCSXIX/djY5n7K4UXVRvRf0zVkPaF+eT/Kwnzr5y+r/qj6KYZZyDVS1Bcj7dKTP
qtgeoahdRJQI/v8eXwdpjgy8y38PIH9JARMhLqtqIHm5XZuMkaQ/FvYZWO/H4Znxb6GcDT/spsEE
A7AHfWTFr5sGV/27B+aqcFSJcvJfos1StxdguPgroBVKqpnTKLDgQy1EQhFYOfhv9Gntyt7ZZzJg
BbmRDt8CPkW4yOBauAv0jFK/EPN8u68HhhAODiexHAiWi3bIMAhc/9LjEu61pvKlHQaBseHAE2Tl
i3Xu2AhjJQvhY446g834PRjC3HNwpXaNPcWpXS48+yqU5LWL71nXBSH4fqCwaqqZMcjpwAm2H63b
LexyEyLv2atay1OTirKC41lB1iGzUludHj7OAreUUofL1UCUH0X9CT6S/9jT0lnz5utmymDiN4it
V99osMBMbbqRuWxQqzo291NVL+BTErB3xUf+82gpJmT2NWzjOPh0XSR0ZEXCah16drvdM/DluaxM
lylghwuupBquFR9JMxGfi0AxUb1jVDs26vtt4DDLEJAVgIy41RJm86eVGRtTCCE6Eg4ZywddOUO2
2pjd2UswE6TUKoI7bh5dsxtmA8Ba/WYpvue2ZWsOwRo2IJdavxaRoIbycWIHRpOWRnyCYceFxfqg
agq0fKhRh6yXVX+fo/0044HMO6nuk5okP4FS31AuE080xnIPBZUw74QWf9gLQYeHL7R2mNkrq4fE
dkbXnWlwRmNZ3NfyBEJyewziZdJBltKtv2AFWAS3YYQI9LKeNxqDpF8qw+/4x/AhQ65yl1IVRZ9v
F7jcqw1fs9CNIYyexSiwvoqobmx+6GkGuxRKcshiyYp+hF44Gzu841d13IMbanZPEuQ60Y9Yt8xO
p+RCywFHUz9xNUBkOxSgCqF4fxEfgvr5DBe56iMT2kms5yz0mQ2amW9hkuQ6Matp26d9nZcjJ07h
MsyBPNDvjyvze53zjp4JvFibRAgZqeg2U1coSI13IdXydlvaH51MgWpZig6cWeOxwE7DYugGudzZ
H/qqIpoUc2LIKE5cusih+NQ+tpzjXTkg9b7IBKg0fm3tztjtJ/kCC3914lKRWHzr5lysEp9xcIV0
DPfxOxLgYCcVPmEJo+yt+FFB2ht5vkIwA9KaQa2OMHjVOL9KtHXrXp2L4JqDd3KzE1rZv5DHZTfU
hvDPeuCF4+tzQbEhUmT1fce4WDtzCqeSgxaPvpnDyEhd5FdRFk3kU7+7+B/AdXf4fDrabgAMCmSF
OnshL9jNihxVp3IvYsC++Fs2Svqc8WjB3bJ2uSHJQDLbNyVX/DYJ5ozDDFlJqxomeZOGSh1aBn7a
ER2Yq+6YjAb9LgVaftdrFEe/SUrkFM017zpwiRF89n830sTrDDGzUrrONGqAUaox1JQ1cqVtCeXh
Z1cQMitFB3bRQ+n7nPIpHa2PsOMclDLESVPc8fIEuFSByFCfiww9K1In2rfN61XAxL6EAlqB0k+e
/OZhDldMtC7s9L9h9mJCo7cAtnHbQi8Cbnahhujvots1yk+SREjkauSYk/nf/1I3yyNVFGyrPpLb
6muJ1shYN9KhsyHiDBVe+TaIRayNyWX2Dywx327R2/tgzRLUBhO45T/fx5wfc/yFQaS1ElRYnYKl
kL2SuyoVaTyw8ba/+eI7Am5JmB3ZIQf3ZoqB2QnllJz7qsyNL9SMZm+rgrRsXiUUSF+0P9StjWqi
Yt+NSPpiNdam9SSYxppcueGhre8TqX8bFqYMfZNVYkpQi1zxH92LXIsJqCpMPCwzEZznJB9+sWiF
nw/rl9rTSGBYuKwpPPt2zcTFknUbuR6N6TCoh31t1fiMxg7jN4aLgfaXY06CQg3a/387iDI5T9oC
hBoTVd7fkbUujagMB4DyhLikuP8r4jVDWSt261nrV5ukPjnNWPG72TwQza+6/gMlplmCiklSaUZD
szt7sLTb+iiATmjkQBic+7FFSjNwyr83K+fJGlNk2IelcJ+j9nayyQKgDEJi+YvZeyebLlX5v6Nl
sf/V30N62oMI/suIg6wskPPiV3GxRm98Sbn1orXYpT2LsP9jCxo+F8N1kqvhhGEhKLivoWTDL2L2
LuG+eSvswGaYilfP2qxV7CKrpK8DwIz0/GyFFqzDajk4kQbgX3YtNCglmNKHGgNbEZuW2IpLtyJS
jtj6ZpP9hnqGYrOEQXYtEdB0scW8+J9YpiDTgY5kTgl20LaDBfPeCRpDufueJOKjF195Oau8zmen
4SlBre6eKUFQoohl8HbMnGrEbE71G3+1EuQOz5+ahHrfrA5BjXb0UvZsnSTAHL2XiwSKQYfuvHzb
m9lHn33HM8otBHl/xuiz3zDmCR4glLZRhXa6v6UgXGp1JqhmJR6FcnQdBtP1glsjxLaXN764mwQF
mw0Cc18WjwE2FEh9xZyf5IpSlh8vTqlZ91gWr5gjwNedlM7+eITn0Gkz+9RLkWwr06AFeiGlwvEG
0FnpDOp33V/p4WShzUhXguTHvckyZGEXi8ABhs9fsYQgnrfiHMbzm/sVFTPK7LfNPZQ7RK+HSo/0
OnaFTUU7w/BLpfL1M8HxPKu45GVYrE22aclV5EKIA8jKzJ28r7o3eS77NADhNpzl4wtZyPpPPI/k
Xf+AMZ4DEWJ1d4kGTEO/YZH+Ouc3wBLAHCBG3/NVNtkhot/c5fdW6mcewN4Xz6k786olp+6ceBw1
vvxcd5WJ0MLDDz+eV3CqPGPFhmnJ9ro6zDQIxsRXlonkIl+pP9aOO8DB+pb3TjPThQPGdhmjFpoL
J24n2dHJalgYDSmu5i/LKDwM8OXJF5SFV5blhIfm6m3bKOEkeA4uTtkHawbRXq0lOkXsS0x9O3s0
wPvTljiKNH9zygG8pcnZR+cfzvp2bOgwsUlcz1zaoeC1S2Vs1nZuRVY7vzUFb9pQud5vdEphQtD+
OpDBoiBsTHlMlzDDLuLVTHXX+v5Ha93SE2bH/vyajGD8M6B+D+WrywdNRhDbJJSlHY5KEUx5rff1
YQ71qGRttzGVtfhACucWzkMFkHrQPfFueIyIxohU0t5ZFeI+bFcg8U1WMT1ADvrEhul6hykev/Vu
1WAIOcfS/n+TFhiO1RZS8NVMvPJg/E49fVJdIXerh3pxdIpf9MgNksvPr19Ipb5fghgzkuhp6/9s
shMGWCB2GwhBoa3PIky1c/ityYUctyIkYtnh1abwWs0Jjnxxa3K2z8eawUQGLs/AtsP3nF2gWhqq
C1OTXYLKDbjW5vOHDapdfnsAge5bdcP5G4qd4Cc0+7ES9VVhgcX+0xyM5jxXQMQIxG31+NhYeNbt
Tr4GGX25DadwnZj/X4X9KdMTAq7WeguStZ+Qc/QJCATY7RZe95/JwPQkcVVzD6RTZP/0gAoSjxgv
3RdRQYzfVParDirxz6jc8JJ7A17Y+oA13Lnw/Q28WWwa33UX2faoMNNvvPhdlOv/AMKY4kykiak1
EC/singSv8f8kUPoAgQZCSr4q7HXRuvgGkcxxMr7yuIZ0cI3gzviDds4QwZd4c510sU5ZXokYnib
K3fHGYXL5E1cO7PS/wVJgO9/qKmsVLqKNU0s8YhISIfW28HNnoPDsfmsJCyx27aPYJAYyvxjO4Pw
0fif2IgyGtBCv6E9j46Nt5CSVa4FMcVxdL83iwYrG/Y2EyhQpP28HOpFNpdevV9xzNaqAn2Eka3/
wQAPBPFaZD1B9Msi009rYBnt2Vw3E4MTOt+gVdHow0K6Tf0zQtA7qcoDRYqMXP5L0cuUnJNVnts8
yJgUAXHihpL9wG4dZ/IBVMh/PjV8g7SkpI5vGkJdCEY71BG8yIA86TJF8pA7E1WBGo1/EPCrSZLl
4TkPjWVF0RF8lQQP7G3kvxe12uw0yQ1fOO6sdl4UdqxLqVDrxeDGh60eMKNVP80SIhoSnMrO/Xnb
ibLmHbZXUeqmjnfJSYW1jvrVCBJ8xKLajEaPCK3/3QwAu5q72WOvk2rPFLRD5SX/2G2eG5Wemxng
Xo9AhHPzJB4meGgtI1rUBBiTU74sd7dGSGsStps2mbrxIk2C4JK9OR8q/+UDE/YCGJtVmwYtwJQD
3SR9XJuGmUkvTnkH857Zgq5lXeA93bewgVrNxOSHKIKLH80spGUCKPmzlBMM8Dlj8LjEOcbLzM1n
24EZHX1nn+GuU2GlgLE2gQxOOHeTQYeCnVtIbIp2XzS2KMtKreIqFpYUSITHfTT1LbQuSbDpynZC
gxTLiXrEJ4GW0kOAN97qP2MjG28ylzvYc2a0hJlJxHEQzJD+4bIbskYxrQGySQLh8njzIDQRAfCa
NK0i/NycKaCSfPWjwUbNbbsW92wTeUzJFSD5m/Q/157fWvR5v7fsfnlAkV6TRlObFqtoSBVb+iQQ
WmtmtVqEW6HFQrhmM4TaoxiLN2G2nKMPKvphzkgmvW9PnNFktA623HGwjNErbtXZso/WXqouGkV5
BYZTjV16Z+U3x5cY/z2RD4ueaeBiMPGuguKbog122ulQ0yXPMAME4HGkOiPSl+mCoOqJoLdIzlzM
Vkz9rq5y1eIFRL4AVAKwhkVKhfRQzveparKcurpotP+MawqgXqu3m75d6d5bzDI8iNDAJh1af7np
I8HbaijfC4JDdTsPWJ+oxSo3V8OZdRT8mUmHQUGo0+8O+bst3VsiTBBQJKGnW+4QpdFmEM2MSCvj
SKikqGwwtVZGmuVu4GuydJ3CcIIoXOU/ItbjxB6ZNmXHTO9l/JUYfNQRs7jDll9MePyhUSzOkLWf
Wg0xlnvYNd9Fq+6Y5YZ+Qt0wkSX1dm1AOeveFHg35cZicUR4BSaeURCJrkFX6wQOfztK+kxw8b8f
FfTgW3Qz2xI1dl3+G13Iowx+47QxNREpm0oDs1GsRUunkvrzjlB8iqXLuSc+iDmsGviNhkLqu5eH
lgFouHpbBkbd0MHslR/pDQX1EI2q3g6rBr3ndFWeJ7wSjquGYX+Y7zRqKLUj2tNPhQA5FIU5l2Nx
Cqhkp1f58FzYEDL6YZRKFkYMaD5RNCsnNhlelhM9CXKeA3CFxYqSREvBgYnX1rrOiRQrdcchrm34
pY6juoCRZH6ifyTPUfGZ3gsJHJ3bBGqoZ0/OX4eQQrvLVhBb47WA9/NIkI873TNGGvT26JV4yflt
gjo501r4YAS21SzyguXftFC33xjEPVZcdfn2gJAbIDNQaBvvwrzNHrWbNlJhJIsCpGa/KtHo414c
44tEcIBKxrv9Zw8nh8gerSELwzLAJbuneA0RknQvTKywy1DUg/sq0rFQdQTiHP7VpbHjGNyQRZo5
Hr1gifh2OSyU+whgaCezbBl04j+LPusXXt2nSqbtQjKuVCKKpUw7VT6xiYkMgYGk2BnR/uDOB+i8
6aU1C+BEDIJKf99axSrdkIS5FBHuQXf7kwXaeJdq2uFAFQ4cBkgCqKAdU6tY/pIdmCCrU09EMw3d
5Ju3XEp20kwzROrcsf6cIVxyNooKP2GbgeeCWBCQUe3pyXigbM+aizqTQ7kwXuEV/tNI/QJg4d+3
4IwG63g607Vt3+Xagp+wGNmtBbrFkrUWi3KqDhxoQe5XHTm4g0zmu3Y6N70QagvF0ZHFyrSwOt0a
0/TS8F21uv9kbvgn0n47LBrxAiPbXGhyf+fNiu8yOOzQhyWNTabLGl0KhNnU4QpinGPTYWBJ6xAs
KvqKOnVQb78+DJjz8n6tBj6SUf5f70472B6pAiji5StLaGIDcatBLEBiy/ZtyrKY/jVbw/zoHZs0
JpsiOmfXLFlerzE6aLtmLRpgSQjdePOVcny4fAy68Zpf8d+uup1D8bGCdf0sxlU2Nt2IPo4JDnsj
/BjxrZ3Hyq8B0k4hj95D910hIvELyPntHsdG1wwFbLaFMTZbI7C/d7Umyk3byF2bXGINMOiNE6bn
Nr3o4KQCgbHF5VDlaLEyiA85ZC5xf22BWfn3IeM+4NpECVbhyrqazmrzXzvDY69RjfJ6R3cBlV6E
JXQBmCPsvDvgpi5oELgf3VWjF8DCDE5roxeR2ctrpEsN4HtrAZV7WzUMeGCjH0Zlb2Vf8jowD4uw
Prm4Ue/L/IMBQHoCTfb0/+XZOCANGBwk42B0eI3Gbgjgh5v7v1IEwPqXAatSsK/1tafbNGUWRRU1
Qqwm+QjTzHUpbYbdPvJ/mQ4rJnP9gYUyUa6TMNGzwYroyFHhY9l93/FSfBQotuHRH0NFC7UzKhfm
oQrj8sH8MgREPC2GfQg3kUQKKwl/VN4HofKG1xs/mLWy1JbeajBHSSYyHFq/PNjYg86AUKqfGp7Y
O0wvoq0P1c2RToeQHwgcnR7ZE0645RrCkYaru2lxXZ5KBozf0lPoJBsQozdBr3Wz0jLp8MhoIca9
XQXWhHMUvfwIluPuVRrRMMV1PSsoWBZVM1+hbUjX/oVftTBcyO3P94lJ/sc4RBF/ZCG4uSR4n4j+
Qec1xw9DbsqLcc7g63cbBt9SNHysD2U0ui/DYat8V2JUAm2b9DnqJ/n0K2wX4N7I1wnTkyAjMeLt
QBuZVdH1DVXqPspyJpMkoZZhflhawXpQ4gS5/wgg8cu0o81ERmXNrl02k7Z0J5VIMxOUyZM+xRpr
vSmagVExty0xn2lg5iE1F/ErA3EhGDGmLCStZBAqNu3fgOVOZNGRE4pfXIJfiuvTLrGf2eHi+lam
alBNk0k3Ge9Cc+KccCbkYi6KHfgEi5dzNwcLglResHDOuZKFubAUIdvpxrsrPl6Zdpk00t5yyeJB
+uZYPU8ZcAMc5UMid8mO7HoF9rww9IaDn7+J7AmvrykjT6ELGQEuPhT9MX2I8KJsmDQIF71yT3RD
ZrPHq2RaMD8iQJ2bwlyFxZCpjoYWzR4crh9WbWMtIgkM5GHcleiutBT3rCJh1SirpxCY84yNaj0c
VPX1fL+1P4KJ4le3CSXH7iuX5aMdsTpeRKwDTrZRU+D1IRIgAE+U0T+6tCqvN0MQEpYEZGjNi5sF
7Wh+of4pguFQPrhvxgKezp26rOV67+9Oe8TCbH3WJ5kVWQompx+gaUDW1QSb+MDczwEmrkHqmDwl
Q5IdpnTObFSMLO+K8swlOOZgaj/mR3IaSbQ6nBaxFrFimuL3uUrq07U/dsIUoaN90hUJ/zgY7SQd
3Zwj68rw97Ag2KMPiVofn0oTckRl0nbJ4Rlq9EMcPjChtgPUpz4bAUReyGvjCY/Gii/Cspq6tsfU
34HOlIxveY/R5GO5MruGZocYmRW0LBJkJIZGV431SVrFsYU54oHgXqwKsGT4i6JvQ4PPx4d26Ox/
N/xjz+8D5MnrEndX6xtnEzG5r1he+Yg+7+Dc2tsDfHqPRqa6J41WJqVUL1DSlyUEwCDoPibRl2ys
qR6QrvIvkuTU0QFxzMWCWnM2SI3S8/B5I+SC9QYEg4YS0/g/OiXGnd1jCuQHJV4xHpqU7OONFgrI
hrfZdR8qxyY78cX7msgwzljiXplLIyilpf/ozogMp9vJz1tcL3lWdTxdl8NPRGBNzSqNoF4A/yy4
fx+RSX+JtXVr33G4tt+XNVK13dzqlEzcc7c1PbIKj874phPxEBASacoEjHTg7BHaem2et6I+/BZ0
bvOwj4pB5Fax++AKDCBHpAgD+GeMGGW9vxYXfTstIqXo2D3Xt1B0tD+zwRRbZc4GmjY5NPCpZqcw
shWA7gu8pCiLGiWPGGNeEpuulnXGx6MLCDtGGs3U2SaclrysWbFhMs9/0z0PK+vzIxE73UgP+Pyo
0dZ/fIboc4drTA0HRT/qbfqoZRTRYF/Asb0vp6h1J2wPpOXD76TL94DZK8wR3opiTTCKLBIUamYO
0cL7+x9VEnfs7Y4xbB+PhHBhVoEKE1LloH2vtgPdeeK7Gb5Oib2KXRQP+SGWJ6qyV2CDQSIqBNjH
N5RIjYUQf93mzCROLmtaU1srDzGFzG/CEzrQhXAs7JcbhUBxkvBL7X47ZN2S5hKx9vbTaRT8Ak0u
W8LOHZO1txu7Hbn59smkZKuTYLEgWuqIP40uicA2EhYlvq36FzhDFr8KPtHyg+bE646hAriYx+cx
I81YLN4lEjwuXdLht+W9sLDGKQRUbck9bysnuJiYrHRhsyLRpwzEifRjij4kPs63GrFPF0yG85Dq
I161ol/K3oYuM+PgNQP52+jBmYEz/GaNrMGev8yHnP7iwKj9qZhY2cHL1nd32fdw2FiW8yHDRQx4
xJWDH93PnaZ1An1qb1pFL/a2gojT65pMBJdHocjnO/1BC5bb94rb2c4DG5XAtICWtvAgRu8k+dS2
d8T9UK+IyqxljoHY8Lld+i7jG7rgXOay3/xRIdadoCT3XNj+WX+z5VfozPJxSzP6X1kneebf3rha
xzCGjiLurxwxpa35nPG3vMeSJRgeX21zI7Jp9AFH72VjmU78NkYfZMxfxsPwNamuHGLNprHbiG1Z
ei1JfiU6MA6CxUHYSJCWL8Fuf1t1AhT+6Ssn1JRzVyCz64u/zcTAnTrVO0V9TYZfnFr93hIf7cBT
jRrBzs6zBJN3Df4eOGOni6sZLCdLrzPT7B3/Tj4SBM6obG3EE9BFz2gSt+1wd3HG+rTIRM5P7eT8
7LAyBmtatRS4YIz2vUvHFETrysAUVqsnaNA7Vov+5nT3/MGj5T5HMD/7YyNTkqKGRiiiDzgUnz4e
NNBiZXB+wIAh9XLhs0HEQKZuF0mD8R1hRAgLEZDrclnLxWd9PDwI5aUksAiC1HS/JeHYnui+fe6n
PJOspKb2DqWOA0xteDm2ESIRGpAunzTyJvu0NpPGXeLZbXXpCaZL1FAixqCk3+nO2Dp44H42MO1E
ILr5VI77e10SKFS9jPwvTlLzydc2R4MxV5oSL8BVg6ZPe/A0PdmadZrq0N/ZxUQYlgPXLYZ4zwx9
v6P4HyB6slJ+QaT0xLYG+1n9L6bMtTdwIIA9bwMYMv7yPx1bFfnL5PI/L5f439bcDxfa2E50P2tJ
MG0sWWoZNyyP2DEi8LHaD0i7jlirgmVf4i+gL0arnkZH41cqqXtr4bKjD7wjiYCDPEbltjHpzfxl
6Hpubao6EApE961mYVIihRCrdbQpel3jWtadvXF/7i28971oPrWTe2nSHupBbbhFzWlH1ZGAe2EJ
RNp7PxZJoDmHUlQBEZHbyYs0M1nloyVq/xp6vNxGyP1tJlEhRrGFgZaeHUI3VwDIRP9OvMeByyvF
C4Lc3MMyMP/UTMx4UjGGQrBRN0N2OJvZpANNWfWowf9wHDxuA23U76EXsWKSncOB/x1if1P46cXH
Rln9j6vrn1wcJmvZxchhQ1eRwGkHvzSeWkPYwcyQUIsN410bBETTr6Nl5qz1RoPhhLVzRhFJu8Xl
Wm/Kz5Sbb+XzK8iwSNb2mlOxuwxNOQCoA8kmz/wQFOVi6dRm71KILA5kc3LWa1KjiIQTCn7RSLq2
YGfcSUDlRua4s8zEnUkUHNjOCYH5Hv89m5nws5E4YJ/1
`protect end_protected
