`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
oLXb6fg0L78vRlBlxm2zkS7OD1oK7GxcAvfMByiBB1qe/N7dPHSiCxLGqzqRREAuW2+jnt2pOwKO
Z4V4752I16jWwNOBPolGpf6WcrAUkFzQdRSa3D9OYSHbrwIthcf8grOhlTk7MMw/CBvVXmsyT7n8
Zeeq7kBjyQSLTruUrAxxCe46e+FpPu/ICA9w4n/f0Alj7IZzsKqSx1pDdwdGFGNdjj8lHX5p/iov
q2VNpJzyGdJ5+x186aTCNy+PzX7ldQr1enpoCTMIxHA8J+P/bZHNOL0fuc3XphsKRgdL4KtS28kB
wg48/Iz7IjDXr9mhBRuUCp+9fRsYv+GocMdwm/QGlfUDr7H50ymsZ8bj65ffv7XzANVbJxXuGsmq
ZLfMYf/WyPX/dWXzdMDvvNc5dkj/t47Cf7gTKV7Wo20xXSTznER2XFOVYsPDXToVQr0w8gpRK6pt
xSLrT8wDr4XXqquvm4BWtpdn4BgqDaQffGlRvQPqNs83rJ0oc/X/hc3lgbaur5/RyTaZds5n33MM
mn2QliABjsyAW0EunwF0Y1MW4DYOXdfayNVEjeaMZhLzUn5jSwASn2L4pA30MSK2TAC/zoCy9vbZ
L8o/XwlO/ckA/Wqvk1c2+0rwLoRXzhajBVoYsmCuH8B0uDlfZoE+tSAsCKP+zBT0a/2fVveZSYOV
zAS1REQumErzzD/5Q6iDbA6/Dfej56v3jT4WcXc+cEcgRIfaNZIT7kBUD3NzXaI38r9dftroTaPF
pAD/9UtsDvapxlD+ZqiAijhbYuLBTvamoLDaNhVxGqi1yWLNZQ84gjev3qE0DR/PhNjkjJ5E6dHK
U04sFr7RWmNpbO71O4t4pcNpUimQ8viswv1uUFyTC/WM6fS/Mz7MZ4+39ta67It1fHDGiFpsQYbw
OmaRSpSHVpILeFm8pSdYJ7C+w81YlnDQdE3ICVgQsRGv8vL6CBTM0OjhT2GhOg7QkoYH/mT2dMRk
SgzDL+lzir42s/GkDpyKTnbUi6AQgXe2XQCJB38oE9iz6TCKtQe3CDtRK0EnUWUMTg05apC5bnvA
ofU0zzGwCzsBFdAN4T6EvUwH1EwfFArZEQ61DvGcJFJxh9nrqOXHd9u11gk1e34AMdoAayLoLyCv
6F1hEn5JXMS/fas5U6jdvgtGGqePYrM4X9pZ+g/oiWUMx3HbXHSaCFeSmaKyhsCbvZjgQWn+OtOY
kE1YbBMxfiIjy5mjyw+T46VefgozWTaPhCrYsW+pt0Sxkv5QNU6QYqA6FAIk1yu1pF+Dx9cX6sq8
OdGXHjjh2E7VJFD58IOk+inFKox1U7cuO5zQAxFHcDiNEuo2vokUDklu/Pc6YzkcRS2taE+DKt9C
4/Z/PnWdbFXN3rxj1fZwXx1LxTnCeTeCYmIguJLs8RkKiR6ktka8HtqoBbKqts2H1oZQ1p5KZ2P6
5poQWz45LsnqiNiUBf6mxjqH3OAsRf1zUaxY0j/x3a2+aQnMbAjYQVB0W5uJys5Y+M12G9ib0gSq
CanpBrcl/tvpsxuR1pCNOUuSD0BuQfX/sZtP7D62CRpJ+T9oizSgrVZ3OSAMI7mmq11ldFcCiuDV
W7BzA86cq4ScS5BZAgFQCKFTz6DYMuZcZLGkDxTffFkMQq3Je0XcX3KOjYm9hQi9108sEgVv2RYg
7sE+f/oznHG8T4jPuDRWxxZXjN64sxQ2erumX1U6AohO61JFY0sTnHq12mSbpYDXudsSUM0DlyxA
IWC9Toi9uYrsAWPugxnKqs9tfseyYXL6H+URo6LT75u1/CUlgsVwkOsFS1RB28ruJE1dhZpS/55V
l/RpO9mPct6Viid+qh77GYfCR9/IQmbqqwPZnxBIhulEhmbOOhcaCwGCHHLSj4dvd9V6usyIu4xr
m6DuVvSjZUQisVdgYS8RvmVnpp6aHcKgYJsLDhb6G4q2C7EWLpItXjnVdPz42LqV8qcluhVK/PRn
TuCgLwOYKfjjoEwLW5HqCmZITu4ynX6AduIYGTd+0CSY40+bjuTNvZNiivsRORQkHfnh8fajArAK
vp+FhKgbJoEfvHKPcPysa//jlaFTwSqFMDxBxWTEJdTEGfM/QLgkW20xh8f1P1JlLQ4rdx0nvY01
7Oe2RY9iHlpeFEU+ji8boG/tzZPanMYE4GVQ40loqxW5pyhnvZkBJjM5rRpJO+JoRrrtSWTrDd5Q
twldpZ4vyriEznQe2mvKfH3CrXOjkKE/MsnrOt3MxRfhY9QHmzgz6+4I5qWhC2xk2lHc0/eUyAHc
45h4OvQN4UQzu516ODCNW1dUpDU0HEBrRBfrI6dtuetiEu8zk3cU96QjxpSDOcUppvBB6QkK4mfs
tT51pUT2lPLUSDHDgO+R8OuWsn8wnDuJPUC46YpApld2CjhH3+s85cB5Y50smCoDnG20M0btZQpQ
MpYyqa+rSZNyDG+1IrKHMSoJtE28kA2JUjI//xd52QYOGy+GxPlcSePB+oua39oePEj1G0igmXaJ
pmV8xjumDdDQ5G5BhycdTkTto+2tbeX7TfEB06lGOS3TM2uHFVR2/0MwaCGwZjUvwyzurj6RKFPl
q74dCJStvuB+h5vhAteIh42Yry9bGimtiuFMG3xX9oK8kqHLxl6QECwQ3AOFvqlCtqzIhkNJJdua
du2xbx3qDemCrA+HsCNa5bxNgvdwMVxfNdeFaYKvOAl6DHNU3+2uTsg1piTsUlHofLxzMUE+NZ3h
5dmBM7MydLvE/jstaEvFpuXD/eL5Jp2QK+WuuUX58/5GAHDpxYYR1mhJoE24hYeeuURCv4JhomKs
R1ufUigmfG2jamhhBKbpdwi+kLSIjW9hE+F722F7qTa5YhjG5925pTCyZLCAUnntsBdaN1wxME3O
Mzn+8mzA/AvZgRUIc7P71vLajuyIGncuDqdGLkIpXF6x9eFq2/X0DAdJ9NuDML6TY9pJrkm4omev
0ICqpa1D4PFnTN7CVqbA7XQqkEl2NBYqfPygV7FYMbFXqN9ITZngUT3QYGHwIkjP4tvnb0VImopA
vGE9PM5/u0R5VEmwXSGJ5fz5nRqUKZ+1fb9FEYuE80RhF64U00BOceYuHWEpNG0DRYzTBgJ0Y8Tp
el46eCq+mQkdVYNSxXShHLfOyuoDXcoMRHJbamBfnxB96OAk7MXmtcQoEfs3JXQcsgcIYnUDoBq9
qY3/5bK9FPtQEr5uvGaVnTu6mzHj6GOM321Bnm6fcP9DDMiMgvwfe9jxX+u3JlsK0UtlraQGKgL6
HNIuASXN98Z5Fq4bUBX733WWGAAYBs3Y+pvDeFEjCkX0Nj6ReszZNXAWdYKNTfJdAQ0ALqcPElXk
3kqUbdpIqAVIe3nfGCZ00EhrEJE87kqbpm0nVzrybgyNhfpNC7Rn0vVIsMUpkbblnpev3162TytE
/iBlCCGmxiW/XzZCC4McV8mWY/rrasVkFPTRvsjmMBGHwMuolB6oSvzOH3Wqx8EbhXo13O7PeNem
Je3l7sS1X/Ez1RlQbocyyj83h7MlM4ATi0xD3uIxiKWcVpqHdemZrV8aRCUkbrtd5whUXLrW4xT8
r1q111c/XkMhBxzEy+N+uk2/+8n+19HMRvJG8Rr3IsDJiWfFTpj5SDHV76mTJOrpU/ZBdFd759wi
i/jaXGupgF800C2IQs1ZWdi+G5Dlc47laYleK32zGHve+B8tuFD4u4D/IB9Qk9faBuQyWfTzhD8y
UsdLwNsthMJJp4LqkPX1UAumgFq6BqttVDrJZlunMOW8lT+4Peba8lWvmoEORBDSn4ygrp5GA92U
QZczdrdnrHkA4IZpU3Dmy3bp+CsjnX8j7pkbAFGnpSuuf80PvBAIx9JjaxRBq+W1XDaV3I2zMT3t
qtdLdjxgakwyhmjkS2q2UpTb3Mi8DwFJAyxQ/y0J6+0Jf0DihYLrg6MQA8ZF0lpc/xkEZEk2vuuP
g9bKd0wOiz9ryivlHVOIoQbn3HnurnFzUcGDLKzX6sXt5GwMJwvA+7M+P3pC+3HwxqHsy3BteeWj
obmLT/hVp3KFIS1eBgv6rE9ozcvWZz95JVhMfTOuYLoY75lyIQdLJnkHJ0mSF7E2UMZsUHulb/uf
bDr+6yPIOTSctKscAo+7EVnK7d9UVLQE+PELNrEH5tt20KZU87yox6LNxtcrquQFmD7kA1lvyro4
Lj8bcPrApECwMgRfJTTNxCKVWfwM7k7tyIxF2OA04qNy49FXnu4hQF5nyxJL2aXY62W8zc15SXxl
hr3OjWQanr9GrxGxV4usfz8NXxGjEPdaXAzX/zZQm1q7RX6c0Kxlfcn9T2cR/afGMAq8O2KJy5N+
WH5y6amm7xWMF4g7eZ129459jrdKzPjzd8cg5ucLNaDwJ8faaJpEHT0PP+5dOs02vTqj7bQDfMQO
KrfNMac8WBnO0I2v1xqxiocV0yb5D4MuJueIGNdGMOPrZUbN551u/l7bMqzzMphK/l5aDbPV5sYw
i4ACSVLJSQfR8XhkfM1TTs00Lf0gkpvdA3riCIdkzL4hoKboqaMz8CcITAqVDLTVs5xkpoP5uWtW
SCFRkTaqkzhKZl3zbYoOoS0wS/tShY5WTNjB6QBubIMAxjjF5aMx3lGujVcKDnLRdmyM47isZ/Ps
I4KFMuRWwN4YK33U6yDoGA9lqBqYEGpCn77xdVp6pN9iYOTLaH96oqxm5cUYaIiuD5RdoaEDoIOV
JOopS+F1XCGv6mLAcMW5KDJsBJn4l/xIr/FqgYs7mNSdjh72PhLrifE9VsBw6JMdjziQ9HS4w02I
wfkmlbXc3d3+rYy+sPJbVcsd8T6BXPsVu0jnbdLaKvNByCSEp+PUDCl71UmrySSH/HkKrElcTLre
mCLtQfE55Zl3G3g8lWMetQMnS2wRDP0d2XLFKMK+m8UznUmi6URfEkKxCTaLI8A4v1oWfcDSXRyG
0M5r+j/pWNsaLc6Sr7EgvwmwfYS2PJpKGze7ZjXiRVJ3MzH/4+4H/5/jxIofA+MpFWM6KagJyPr/
MqGBDy1D85fc7OVP/ZZt4jly1yox5SZkFfpJ2bERu+ntEmltXo9PoWUmBsWxVWFSLfLgjtmF58G0
lUIPvYrA+99cZFwzwe+bguAPE5wAkd1LAQSEFDMQxa5LPXrCucNFAXbGHi4oCKyv2MQBYoCGxnMl
hFzdoXvtBUFSf7xxxR1Z4nid2ouHPceC/6uG01lAiJv5u3pnFTrbdnGL5VFCHWfzWV2ZnOTTFMB9
ZOhDaRx3lnVgdJnLQpe0vYYhc6XXMGaJkqfOryqTVtQ1keJiQ19sPY6ovF/T1ZUXT8qjuiblBQiy
2DxjMtRysrXk3vy5edmFvqgaQUJU8kRwK8KFXmUZZwnzO6ICjTW5dnhvYkQdPP/VsdcUflfogP43
5YKDpkyQVA8TUBsLovR9w/WDkxNJECWO7RmpVXrHanYcsQzOFzwOwtCYXb06WK/fm18XbhboUmxP
UA8pxJHsut+Y8KlsFhBYkGVNvu03kPQJ6sYPqciLzNQFWmbUiAt2OyBZD9wx0QE9SmsqgZVs4QYE
eDDTtTeCpAwhoo95VCuehTHZ5wnOUGRLKduA4zuprdktAQPU53qRbOOalUKht7v7IF5OMSfa1Q0p
g9ZhpMTwsMG1hQ/e6JHGPuDUEdQ7JXXfuKz4gdI90+G7sAX8Vh5xQfeQxLr7F9wmn0LxjA7JZxy8
WCKO2yJe4mxGACHb1kAllPkRvWnjDWnRG5LfLx1hpy+9HLk/C/eg3diMK0TPhE11R3ZyrrhTkraL
tJMfOX3E3c8CQXGI+0Za2IYWT8AaeBJLr1tlTbLbVAIlaASTS3ZfkuGjCgoQc0VLgDpG9R/kIwAD
q3SHfbd4rqHh8UEe5w+N6CJTFDPBIskC1YIkujohZyoKFbjeXiFkI77n21ImLcBlaBWvJ2PTaR5A
Nzl68QisRgQvFMRZ763OkR6Z4JeENB6WbCACpMEv6k01xaFpWx0qVcYOWlAMaC1VamnVI8wtJeCV
88D9fJqV1SCQbN86fPoBkRv+XnlHIZhDjwtWy6p1q3IdT2iR1bbR1mcsWs/a6zBYtQijmZRATcYK
qCsuUEOzzmgAkYwZrHU7h76qG83BMCALCHTpYK7TYHR5ZdOsPeWxpDpogNllV7rJ/k+UHHzccLeh
xOd8z9H2UP1RZUejSf98u0xRD+FrUlPrqVfEI2BqlIidJldigLT6ciZZ+Tqka3ZA/PaTlSeWr1bp
TxIMsGCxKZQ/ijagDSfSdfQL+1bUXO8gfTCmQW9ScnM648y7Oi1fRxNOfDAAwIiRWwLV3/0JUWW4
lIYFt3kL8bCEQKl25+fguLPqS9+FSEjoUbiYBpgFMSj2sB8LZg62E0GcB+mKj4XECTuJCBCESGa3
2fs+u/NvU80OltH1T35a2s2povmmFNq59DNMLbUkxna2Bed9yAs7GpCdci2zaOfkHydAyPHPB62o
jDRER4Os4aExizxT88vpWO0xrQevGpAE5dpF4+67K4n9jKwK1jx1Ox1LPZqpSwciq0YoxN36/VS8
ctdp+KDl1OWtGdWrYKgATV0w+jdHAjrieG0BlmRfJ5r628sEp7pAviwCqUDMqO9KS+GwHVqopb2j
4kZMvAgozWMu0ek7lWETPNrd1/vDT+4NsJ+Sd9ZAWL6scwQkiwYEPk8NV/NB5EZKja7pZOToaEaK
L0nk1VRHk9kR8MhmvWZlirVZWszNm4xs0hr3YA5dnNs2vPbWVBI8W51jt0FToALGsYih+pAlwFuO
4ISYvFki2QQOANIJ19V/q3bQo6sZANV+qqfLdj8y9amYkDUPFVM8Zs5B2OFa6q0CQLdNb1WDcuSK
jBYouY0Nzmbm7Tvp8VckCrmSIseKEpZqCRFNUu3Q0qzMPaL3cZhuBsya/KQsD9OzG0IS2xNdxqdo
vk6WFTe8kfqRZIHNYDVimyFuOzJ3cl3LpQX43MUSqcL1AwJIISaJ8IVNfsTssAEBKkhPDg9vc4Cn
u5t1BfqTs76Qm/+HGhgplBxhyqB5KweO7hDD1d99BdhV1lRffLL0Mt+y8hAljiGq4CXYuZVoW9iQ
UZcfr1AqPISZ1JbUzcsqfwLKxM+jVUTvUewpv9t7dZk2MYLHxm7jvoVZN0UAmeYz8KxoMr7irgS4
WLyIdJMBqwX9uyVtLmJN2msDknT9ntKj216xE0q4hDAfSavqym87JqWl30mzqZTGIim4TOQcAa/A
OfvMTyuoXlj2e4mgY49oRVbUidzLjmP7V5SWErgUk3dEOLehhT1VCIx9PEUdZ3eef+LdoDp8E8dP
MF6ht68o+9lkxEq+efw2zIbbGmTBn4FXJQ0Jny6tIHNU4k7rxS81wHU/I4ye//XwQQSpyappAuCE
1RtKic7tU8RTVXJp5hqu/cUeBpGik4ltqzk0rK+xCAEcdyT3XmpBRWWLJbms4CjoexcGDF0nsaP3
OC75WE+WW51RaL7AP0CjwnsuxtJtOn20SOB2eHzWYC+1dn4Bb63tvO5gXk7aHl71rpS9ykETk6Xy
LTdOR0cf9jQ+JisJiXjktUlyv1HtoyxzqVv5lwCSChWP376lpXoW34uqdXmP6ZJSPkPx5kOSoBtC
NE/oAfvMCFA6jzVrs16QPqFGYBxYljdwqilwGTM0FTFEzSZt3J6q/oP/WkimoRMnRPtw5miYDRXO
yeftVxaBIYDe8PDLCwhQTmcOTc9iUnzWZ3LOd4lt3NZFczmBJlg62VfqB4Uuhz5spkxnrQiMywqS
yy0ly/CbmfhiHQfsZ4cUXHSTjvNz53oMITbQVv306SzgG5t3wrGnobKzMi1cnd6Sp5u7DSVSrtbK
YIx3PQRHTeUvw8yFx7hQVd5Aw6S5zh+aDnUwHwSkaRwXQl9EH/eCTOHCVcxCIBGGGOtfygXTMerM
fLjKLAaCNyHgkw7gOFDBL6HAaHI8ahOJXAVK9kaIm4IczGf+nivCVXEF53I9/CgHRrzVU7EvUlbK
XOxFM/2SVoo3cIuKJs9Vlrysj5lPfqr2R9TQSNEdazj8hSfTa4z+u8CpEQi5bVMEfcd9tgHSmMeC
8jb7BjF8tLHPQJpIV80qdHeUxgfX2SpdC5shUym43LOC2zA07jc81mAB3BXtH7fnarU8cxQ03OMx
WEuN0DDTxGiuzSEmDWdCnlbeo+LkMDylrdwfCKZhMbpZimqYE59sad6O4t+fSwyQq8Uq/Uqseonh
lfA53L2uTKwfYd6JNdhYyKOG4kVRlLeLMDsy9pvoI2P5UYxh1Ndku1SEjlEIp5ebBBrsb6k2Yg7Q
yzgq9h+oMJ7ZQcabhUq9Vmx6JVvNQ7NnTxg0viZtXrczYtYhtTGHw5KnvXjj9F/3yF6fHyYu7Woi
CLa6iUm4wbekStHQJWn4XhBYmNRRfRnz1CjxemwLaXNmvd7O9E8oZltEyj7F+ZuTtTt4reAyq+57
QQ24yqMjmJEmrYb0HWSvKpbT1dQwEC1mmsxEIgdM2szGq47U/qj9/SYY3R7f3LZsRA40bAsr1BmJ
XN2pTWYr43ctWlUm7OnqCtd7zdUjrUIUfGJSr0koEDgPA/FkGVpE23vL5I9OZHkiS1D8QR6ZGvnZ
CYYt6zmuydlNs4u6xH0dzzOdrZPl8JKH88wLRyIk+vyz4LObUYla7sZfiGQ0xXyP56jhbN0Bsqul
OOM8FZJdTWHZMjl6OicM1di1BJZtvYgJEJHJlsnooXgx1QwDipOLDbiSxNw++dyXGWortvhdfj/u
giHzFqlbVdYbxC705p5v7LNZIdT+GPcl6LXMJsE5Q/8kTpK1/G9gIl7gcOu2aTP8ViKkRFe3ozRD
Z2cQGJtYd5UaJ4TFn9kf6lckNT9q+nRqLP6ZkTSIWypKruLYcMSTCfOTQLdKkDdfTIRjM7J6WeSv
kvFsrdj19Uy+DYKyXPVdwvP1hY7NbnN2VhSFA2YrVdNktggfNJYX+qHaO+52PfVLJkzwvuQSggJr
9HrM8JGkpPiYdYtRs9EDcNwSq6UF7p4AQxch7siUgrJTrj78Ce8LxcQDfdkZbOPpuHjzZnBkX5zt
Xte28EgvVgQEDF9TsRoJMXSEc7bjZN6HIcPjyQ3d94rvYSV7Zjysihwrhp8HvZq5l3643oBIkKMT
NtKDyTI4NsogU7DRSug2c+RHKYSuWNZY7qOZZE+LsPC25un4BO2ImWFWw9f6ZdXcn5bgxc3TWUwq
sYy4nJ7uFam7rPxbttZ4GnT9EZiregv9tAXJxbpReUldZBpyoS4Frew7IU7l6KqKOnzWNiqTtpMN
fOSJhxZAv2XyjrHOooG8Carwi1VPXoT/eP6x8lOSyCGfuQON05pz3B0gtDagauZ7wG8wo5QRgA47
GqQy5s8+rod0wAr18a1iGhApQRHPOFTOG5pVYQroegEtA4VlIBg5QeHsgNPqbkF3i9uFmTb0DqoG
rNGrcm1Xx20l4AJaqH2UgqL1317suLCAo0ngmuTp8dVikfpTrPsTzCNMQf0fOX82N8upnmN2NySx
/pPTpWtKoPcfvRObPAmIBPSaflAkzY8L3FAcpvd8jKPmTYNgdvwKYTJZUQvcsWkotI8UKFcqBCaL
o4tY/ELSyrI6Tk1Ovui1J1RcgjfjGmjWLho0pUJ1GpkDLh9rNbzf1ZCbU4EqEeImbMxfWiT/zbrF
q3LW9LXs97PKUrguvA2Qdjzr7gi2qyPl5h5gk1WRQMmltski4t1Yo+Zn63r2TjM9Wtc1Pt9dX0ki
agcCxJm4XJ0GuRb4LhmaScOZBHSbXrn4fDJNoto3Cx6b/hBqLxgk5G1530tz8aA3Ucopc1Cg9hLV
2LyxdWnGCB4e5NYEOpkzu1MuxAG11Lm0IAce4RoL1aSnf5vZxAm84rJYmuRgJ0Xh5Rp+yenslxHP
Nn32C0DZJHJ6hTfP5GWNKnrpPIDccQXhJet/J5e27+2UQkl2PvtezwQMtQObtwlXjoA5MtlfE3hO
/7ngnbcuZj8v3AcBsGC4qZTXfMUaa92zDO2vGrySrZKs8CDpnNvNO6uj90u//UnhtDqm/laBInxm
AOHYaCj9pwOV58xD7AB+ES/56F3ru4xMS3NJ6jmjnwGRXqQtkauufwSvu+ncUaZZhLNVDKQycFnY
TqYvA+C4VzrxlZ3l6qZNGHpMZmMOumUou+sQeUbx9GZMSuc4hd+n2edmEDbwn/T71WAFVX8buWnj
a5OyYih/JMkmO4/aZYpo9z5wDKcCPQJepIKcaZZXmPEEK0oHrKjWO4vXMaf/Xu2pQEw1Kysp71VA
xqM9gRaUaCSrddR0nVk8l3a9qwYuHfdGcgKU7xic+fykgJSRvRhr6NBgOA2KA0TEqR3vN6myXBv8
EVFcxNwlixtnnjuCy/SImfeWplKkALkFeCgzen2VtcSj+XDlo2BJLgc9H9aJBjuxis0FPPwnOqDN
vPBwAFHphEOXFbg82gDPKxCzXBB+fV/dmATOR5Wdv5a/iIH1NeNadJpTHGkYDlVK0mCWjlASyEbv
TESmKsUI5VhmpvYhHuqiSGqhhLw5BIU7/HO/ZRESXpJ+eSsrvEb1C3V5fWVAtOwWFlAey7xf4Wvu
Nyu54OuAJFGZwpA9v3OhNxz39itCVemxTX12fPNCkw5cfrFksrhaalZlcf1qOUT7RQNEMCqzvjql
G00xqMI6tiHCS+Bzg6BnzBhHSWC8WtuSGQT1Wm0Zwc9t/34T6F7xJeyM8oUb9pyvGjKh1qRcno/t
OH9uRroDEGxuvmmIcPe7xBto3IYXbnKbEMZYFNU1bWAnYWTQx70VSUCquIGCBVOLeMZP/HWRWj3B
2PeUihCvHIpKKDgdF5MGeU5pHPd7LO4geLPN/tCB3RybKGMTf3g52IUE1thkvhJMINJjxQBH2b1V
AvQkTofNCVD63y3KTvu6OYpDIikQMcrUvCherOIQ7DwYb6YuKjt0+76GG9J08iZGziuxrfS00OrU
U8uj4KIpOqU5yL6xa4fMl2SJIAiBPcmq5jVYfQjKfUa3PlNl+0ojM+GIGeZdFyfX3equgYaIwz16
D5cqwI8F8gxF0pzkTa4kbigfe7e05/NNR2+1RbMSchgKuGPmZzaWVJMHKCcTxQCMLp33YXAWl+/+
KHWlR4/VQZv1w7iLUD+Mq5cdFuUHg4SsCLRUtZnCcOeIawoFwiLfcTOxpdHkkAYZeffoUJJgbKWC
rU0A3u1YhOahrOFG8hUTnJkU4toD5GoxPm+CEdEIvGOGeAINgI91L1eLkymyaZQfKMmtxOgcMhSW
JjB6qERg4bGr3U1QADQ/uwVRoel4q2SsEZl1YUptMmuRcvw665U7jWgCywg7lqLQGv4Dhlwz492C
GbuBylY28GIl6mjueSXyvaJtX9SA1bbPTgd0SILuLR2wSnsDvtXRc832xLyAUbZeyr4NEKbbZwGB
oiUF9HlyJ/pUwmdCw6ir9/ms0D03SbAQ6YggE4h55Ck3hTyZ/HLrlde2V+DbGYcHp0HD/UpHH4vQ
BuKAxlGGlPUfS1hJ+NuIyUEXkJgyRJ4GQuC2F3raqenQVhWgSuCTPDLCKLzGZ3Uc4/hSX9cJQcqG
NmBeJCDdJFxIOLxndaEtevhmf+mLBkIKpcUWDn9mjrVctOZSDr60j9fc7kasJt3qtmzTZFJ02u4y
izjK5mjQKfR4zN/DyS8Amjo8YWIbEPSlHFHuVAogRlJcYUJwrwTssiUydOdix3Y0hFkKKrvs1Iye
m83XoCb9ueSBW5URh5gSB6yI7U0ltEDB5eygu96dn9JrUu4P9mmqMjocxeOsOo++EUOoY8XATdHo
XRrBGkQ+HYpsEqGRpRz14WHYxcxNtZSa7K3AJPPU+8kHZOcH82HlIDsLW4kiaxzfkdDhxay4hgAR
x505/gXKsoldEmY+nCuuAW5M746JnIF3sJe71MeC4dR4PWO0MUScOF2lT/31yP/4i7ntlt3sJWWI
0PcW0+ROEIFZjZawRBPtv4OfZ7N5tLPpJQxhZx9hnt1PFZ3DOXconGa3Yjjok64ECo+yjrltiDfT
D1SI+xX18P4cgVUqQR0HjjnE4najP39diV5ke1MwQM9zU9e0AqTbMTrHOY+7uxW52AGzfI+zc/ng
ncV0dTN3sOsWsrpvNd2nCcq5hNEV7AV7FKu2OXRYeomtHFcm/+Fh5oK4zKk0EtMyeLUoEOj39cmt
R1fKSt32mJq/LS45SP1n7gNaTNjVoDvMknjqMNmBCbpVVabf4S59DsTAbni+SoHll0S80Rez8eGp
5eWE8tnCLCX6Ew2ZXMm4p+T+UHUxfiw8KtbPhlUAyZ8dUeeNFLxVG/69ME1jp0pF8RJvUlepwmFi
Z0y0Hoh+RcD9hgGjqSj2gO640u8C2DIoa/I+hPqlaVpnSA4DPHCf6sJihMTpDpZz8RmVJrP8gqnW
7yLkqW7s1tf7m0edD6aN8LpcB/+yEH1QZEUCqxVrinMKx8tpLyCJuS+KeL36LQi4h6NG7gp1Ne67
vNQUwyX3FBjoaw5cz0w/DjHbf3Z8B6rxKj5R/RBeGA0SppHmo1u6qRujO7EZtlqLhbQDWdtZNXHp
QypS3BsNVzjPVuUzDc9hsoi1RkHL64AT1t58QVPPaQA+3KvzA8VcFwAG2EfN4H5bLZw2UF7ol/b/
6+ah5NHI6UfYe0LPKGXU7y6VJ+G/nsPjUK7yCfywmnASIye+/jnT7hG51SEQYnl45y6IFeE+ViWw
T06gxi9ojzSM7u4uh4jkzIr0jByXWO8leo31ZA3x5/dh6kJSlDCtI2G68mPRhEFdhDUO0fI62Kf9
I9IOFfp6x26XAO0JobMNySAxZshrW6IMm0xgzFc4dOrghPFy78ZiU6PMBdMjIqfBWNkUNqrXf/HT
kMNHxAMSQG6uKo1AliSazRLgkrOsyGnmfZOnpOWDPAp+0ljtWqivJ+SJQVpsJYftD8KqaJpYsaUq
5PgGcSU0fLmrp0YBrV5fPuSqoUpM23rIGMU8d5UnWDzw7a1tguDkC6u6O3dIRu2RLNhp7QUTSjG9
gyOFMqvRmlaR0SlHz4vjOHo780If7lYQUQ7NL/+Kp17cYZtPsHUQL0B63tUx6tvBORck2CpLEV8h
fdKeODTjxWR6ocN0lnu5athtlbyvopjPmvjlb6+y5zUrd12wPrQRhLysk4ipG45SFIyLLwls7VYc
mEYxYQI+xg51a/lLi6QB/5hDLkG/XghkABdzzSgb25aUTehRMM9SZ3+V9ND6HHVYYYs6UCt208q9
gIyJUyIWvFDTF33updt0ZpB0YX7rjL/WcpRnVAzLoJ9ot41S++MQT3xgJcpSn+Gpq1UUmXYZafHt
0N7o1yIbARqz1nvjSzFdBQpdE7KnnM+SQ7qtsNSLp/wAwvHhr5wVDHnUCRqzLH9mkkVzuqixhWty
AwRJE5+QMWoBm+4vZAMERzVtCbFCzWrejCzVIwGMNROO6f+46nvFkeV5lN/ze4h9+0SBbqxlWtn4
gUP03jp44pwJTnP/I4ZdYKZfrQEPXvNPCjclZ7KZbnZPJjHmQem/uAreyF81WuWBp8Qa+fryAXM9
NFdVym2/9iev/abeOq6V/9NhLHJE70r+awoEjfCG/1uWSMBSVqcQP0Qh82NalotNXPUyeo2gXOM4
0YaIKtF7aFd+yaEUwyvDHU70746bSkWLTyuV1T2URIa9QYZe56tx8V4aMk/i98WE0mXrSa1k2aWJ
72bhyfwuzkABvNKKSoLqTaUDoVNgT264icjZGPMt2Rupxt43lL7H6Q7KtR9vO4Z1vg1kEKq8uir6
rWJ2ja5Qa8ntpOKBkUSRs1Zkkxzo0yKr1Z9tEqXyxcurPhkvQNskKYpjyTc7tBtcVrBlYUsXS6Jb
Kn8p1KNIcmAnwwagpnwlCzGX+xfazC4WR2YHHNt5RX/c5OO9mhwqW+pB5EE/qsGbaPSTE5kErrTq
GNZx/KKKw/DkGnk35w24nR2GTkIyRbgqhjUKgDbQfjKh+VQLTqoExpeo26k+oE/Pa6Vv9t4Kj/DG
w4sYTKVLYl7JIoncdSYm3c+d1nSU2MrtBaZ/PMe47lNflZZX6HDTVUf9RdeV5nKMYDirLFZO8idK
Zc2XrnWK/VmpDV4AUHd+d4/mYfut9twJcm+oBUW8AUoHGqwWamv4X5Gqdi5mwPaX5Wy0jsnjaHxj
RF6u2df2iv22xg2lpSpYM1/RBxpCQPhVNwtCBANOfK1hUSCS0vP5cAFHTgph2nCaIif3pEi7S6RA
s7V9JJlfwQ28gXN/d6zCOFIGry2qSeL3v3uMkTHrA9OnqrQY/W8p5UC/cdMJ9oTnSc+TsyiD0d52
VvtMoIt66k66WkagkAsW9R/9ZsfKFHbE/1REgGFfx3kQDRw26ZSaNAqbLb2SJ9Sokz0ki8650kyj
vL3+CBdzmc19Yi1OqTU3gLVweOig0or+L3SsGHJfMU9ePyt0uR+MmHXK2DR1LfGNQFeidJInOXhi
QsCHc+9fzIzVPOTGPSXnrTcY/WWMGRq4b3+SJeGOpRfG5242qMZI8YHkigH5nlfPY5ua6QuVlHix
/l5zFtC/E7gctb8CixWUB4XB8VmxnBCVTPPcltprFtx3pqimnEezpQAKGdPjX7iJ3MOfQoYGjH1h
T+EYYrz6o3efoZbmbD9AC5WAXX0+hdXlq9Uc03a7pNWlJPMVx6F0kurx9x019obHqhqaRUoYQWmv
8CMAXxO8zlh+zcxUHNHjGBEJXXrrF1ajdFDYK9oT6SKKip93D/6QS28TJXxYe23GkKnyT2ycTbdZ
f5aQnF4KiUmrj1bSVwNCZfCyeYjnf5/0JsWhMfrawI036JiIW4Wg+8XkveBzxOPzHV1GBCVGJwEf
xF6w31+Jwmd2R9e9LqsKTksx+9N9yzB73lrLukxMbCLBVvuSt2cuaFMtBltDbtEQRnyIEpyEF6Ul
8Pj5SsdmQcXqsRUGiROqVm1l8LXdcXWK8/SRsgSCDEzEjaBvZMDWjPsgNVtbpnT7lycDxV4QTyPS
rR8HXVjKZ44xqxPmMesLM/vh7psy0SKtgA0DXP6K4YiY/j19NOLbSYZTyQ6gsv9CTMf3CHxA9BEJ
uj7/n/OpRZeAGHD8uxOprsvTefOpoVyLo9ak7Rl+cWp6lxOQ+Iontlrs1+QLrxpKqlUt7QDW2koD
Q3ujJX+3JOA2WotxGnMgBLrcX8HexbPXxsDVRv/tPQbsU4bziqZH3pINDfNT03oZImctZ7yEOJBK
HU7pN8puhKoSPtvZU4Lb1LhWpWUB/0RpddyhuM1K4mOWfxM/1YHIzByRBS6uKtp8agf2aMeapVP0
LQtJYx0fbcdjtiHNr09KJem8Hj7qvC5ozrE3HlzNjfn9mvGAFqIGjhq0iZ25WnUpBA45CSsuYEO4
9LSCRrOtskCqXp9/NujkD1xaV5zd7WD3VG+9hJXBSGPvXsk8w5bBRKijtb41FjGawqAvcNPW1DnD
lRVZOiBhLrpM/kzBtxhMexw2mVU5NBZIskV7Q+uzYR/IE7ewxKXw/tc1kHRqsK/Mk2x898iPlbuh
xX03VnH1OsURHsuiupGDNAgS+mSk06m1CUo6Sby+5iQLO4iAFaSnATqJTw02wmzVoN5Tn+hFejQb
LGqdDzDtNxUX1TSzPyhHBARVP3mYTmoXEkibYBO2fWZC1AfUMjh3pvbO0yyc9Bpe8gme7VgcF5Ie
Nfij+meIakXu7+zMe/Z28Mmgfuq5mn439PAMARH6RzjsuaxYdKlOUnnVktd2V3XD31a92oCTvdnY
vyM+Ws4J8RIeEPEa3nuHdtp6D+8W+yoAyf0nKUDs4jZ7oqqkmqHK5PsxrW/3kDIySOw0R5xpR0qp
A0T+EtkF6fy3ggZCTmzGsrITeSKglrZQFJcMcx9QO5V3bgLDJORdB2plizGDgrk7VSsVd9fb/22C
20vVkayNT7YWq8L3ICj4cONfYzyeNxjSM5R0zEJWf90o+37rF7Rrzwo6Rj0uqyALv/2QkgkM99nY
PapVQOnIl7Nae8EC4hBhc3IbCR4Akh/MiyLz2axTYcQn2rAt+7hKzMK0F2X0AgYnK+F90Dla44RP
0z4wvaeIpBq8Kj/iZCtBaUanq/wY+fKj2MphwfQv0f6dN56XxjWkHt1LQ1ynq7bWM+GcD3tPLXJo
U6eMuf8h4LJ2mkyNzUyEJadGFbhIgEDAav8p51d61PZSZrXPx62zDZt+f5J1c0Cfx2AR/tDRWVip
10iAgNFz557uluoa4t/9S37jCB0EtQtv/zAmMQFNziZ5DIZ6M0fRFgTgWRN0UqPPK1An/qPWwYOc
Bi11I1Gqtoz5YQJ7j7sshKWRulfPA8EOrRDtx788bvvYg4LQjapUSu7E8tW7kMe4IWx244K7dYBD
Y3Jy7+nIBevI4khxN/juTU20mZFOBMS5Clyjwx67TqEtJ8kdOf/ZklP54jHjHxD7/AQwimVgl59T
gQpwM1WfibYNqu6FNln6EKko374uEziEoljFJMSX200sPK13lJzH+FfeM0TjaDxQBAk8p1VZDTgU
8arhEvaTX1Gh/APs8wXQUC3D0IkBicVNfU/vuMXYZmpQ6GMTKvyeGs5OUaVfUUwxqZh0IOlefPPc
GDZGpght2FgnboMhzvAbHeFpHQiAuMdG22XbRiYmjJnjILlFnMu2U7BXB8T+8RstGLRSgxGJdQIj
qL/kydvPQN15ChZwM282durzOTxz09ynGqAUMRYY5tK0YA5ANQlrm8RWaJeLWub8Z9UxFXTydVaU
DXAGZyofVGYsQseT5XT3jNXLRM/Jg9jygARNrx1k33I3VEpTnKO6xJI0Ww4K4W1a2FbUx7CSrTU1
+6WCjIJ9xLLUEhRGdqFvOLYjc6gRYrcGuQtpUEfX3Zny9xdXVV2TQ6mToTV9y7CEFa+KcIv2ICj6
UZKqrs1dpjoNTwKPBcyXNAOWBXWG6UXyVWwkwsId/fTs2cnUeKBvIjcHTFq71CpYg+ZZMKSsB/ID
QoMPKrxnK30cHKDZpUb8p5KE/+BPQrtfXV1fLzuQcKW7JdvRnDgYHd0l8Erd999BFHprgEI6Kwwh
XDhdStTDlhh85JqZBiIq4QVK2PhCMNJ4GAq9hglkyVZSF4jhuS2hIXWFQjC3jW3W5HPFhAEqPbHL
UNU6qeiuUn3SvYxNuEkzCOypZIefHSfxDSonTzJzQeTjih9LkE1SFpyOYfLL62u9yT+a2WEjtPUN
UhePjRfu4MqPpYEUUgzwt2tBSFatngHUh/MAvCm3iiUe5k04Y0fqmzogCwPMmB2LdsCpYImFZ22n
MiWLNFIpDwzwyBHdwh3wkGEMp7QbqB/8Z0nYtnVAfLT/gxInKBP9XoUJ9mgl/D8nmGgpykmfyBd/
Cf8tDgY+R3BU5anFFfTiqqfGhQWAXDlAiyxx9t/CdVo3IonbUU5eUa7q1kC5V9r9jUkY+x0UFacj
+4IfvyjWsW00DvDTVxRjowuoFUzKHiePaD7WKuBMeBKtTKsv/z3z+xrE1lLu/7j/u8VtWXBgnDVb
qWb9NHteIEZTXsWIJV4nQAV241LhrcMbqbua6UxGKrNc9GAB0CQWMnpIvmWGwV35Zuz140K3URuv
OGdfqYl9dpeeTJEIYYf34PZH1V81o+ASd//RxF42gCL2D7rJv/nNKZ7PcUifJnqU5lXUyrS5g/6c
JaZcO2vZOyzXtCXYNThwwjFtgmK/CQ+3PTpEMiItpOQCXfY/pGNJFsAnui7udaJ93lXtUt0rXhsy
2Y7gPn2QFshN6P6yslsfrGviMAlc8waY1FE3kLiBfwYnUJGydt1HRU5KOBxmDRfg2aEjvW8XODvB
6kkZeUl1lKUZlxWlW0EKG1Zp98mYN7WrbldSI3tP0/zLSH5Ae2F8JeeAuXM1WyKr8FDKKhjS7Jvg
mTpRMULZ5yjyW2JWrX7ivU0TyTcO95OPYpYltk2Bw56GMPoppLJB1ZWK3p8QkRNX3vdH631l0hDT
aUvbUdIsSneJfRkw8xqoEoZjja0nEvlytycJDpekXMhvJOjM0DdSI0VlsI9gxlG15lAeRadmgtKf
NsiYlEYeGtCnpOzAier8ViUmA3PHDUwVHC6oBG5zznJn3ogaKREg5dSmkY3ZkRQVAYhlz8dfMfwR
tMa38Uyss5M6xh4Gb7LGyq+eUGhQ/MLeOwgZLCyfPx/jSLVrwmazB4UVx+CBxModYUpm1YiqdDQ6
iiCd2efp7hnaqtvqnRu12wCAznQ/p9saZxjOZL0Z9SNn+gp6fpt24/IcSIT1CpdfTGamS3aylEzp
1dJnF+Reqw6FCT3adWBlf81M4sFm9FBk5PHe6EKzI3v0Y5Kr3A8K84rNax0AB2gppZacxJB0gwec
4U8jKN8d6cd0SXsuqytZ0O0tqt/ehgt7zkYBPg1qk2leQYpBO9lMRTOlpmcedOxDuC3A9/+s5MjK
0jtXJWFFoQ+QWqVUIL+ZxyHzvVfVcKFC/HHtnkkv9sN96xEwzNH7NVo19iesHC3R7eGuOcGgS7oD
kF4HyelfL4ESU9mKcOTzsiMSDa2WZNpzb1pvWGDgfNWzssMYbd/ttBuEvNgh9PiU9dH02Iu2owj8
QLlpK9TYDTCIjPVVuZ/CBLwvxlO9gsVCB+JTNuOqjEHC5X2inFhzFY2VkqM1TZzX10lNoo73vkgE
YXqGPqmMIMDVYQzxg3i0VC2T8g0L8+2yps2hBaoQ4yQn1v/wvU00gRQPeyoN7ZrJFB8lOHZgZD+R
Iy9Vu00Eyyfv748k5XY1vP7hfj5e9kVT0naQQkjUDnbXIQXkkJbjJhenQBJsR118kYLjjPaR1UVC
nzLhYlQV5O93HgaeqALjPgbtqHDEwuDUixcKpLT0DPCreqRkhpowsXOWAArMC6ROyi6TeoZ/9xM8
pwQb/DA3pBisUje+QmZdh3BZ9mVXPQHNgsrWwLdE8bIptPfSGmb84dKHTTLiHfBF62ECPeLBQpdg
A+qJ87BdKw6L++RksL5fxZjYAM4iqpoa+Oj1nmmdU4cXZ5tF4f72vw39wvroPMISUEM6oSb1/nGU
1CQMutHuhJxaFeSVVSAEAk2pquynSVYiF4bkj8GIX3MJlN/GZs0jdq00GgWW1p1hk789EUUoRLFR
habE9rtQUy5N3DEMnU9U+h4dP/dbGv6kgGivX/N3N6GjVXR0l5XxOFdWEA+nixB+mtv2a4Tx6Ig4
/bfjvldZPoeX3KWmm5/XxY4ewAX+yYiRovmzj1hlfOgGps7XqNccugyQ/2hp7iXMSIeURbO7y79E
9vyhRKoy7Bz8nc2QrRg420TD4xiyCaW3LeZKbxgR8DhPjYsjVsJn31chS0YLas5nGJo+0r0P8FQL
snQbuSLl2dez8y4Fcq/qj7CeghobVZOXNPRz5iAtmiaCvFsfE49nx+el8s0+6AjPRJ42T5BuW4xb
vSY78eFuey1flf1ScPCSmig2CUGANaujVrKpJEVZZJYcOOhgyV7Q0+iz681ptW2/9yfMc4y6Ci4E
SpBCSEOeO80x4xqGxQTR9HRAB97d6FjeTV93iqAeweNanEhPpMZviQ4Pk3Cm1FHj5EMGoXzS5mNX
afJHnhZNa4QT1VYSyLX5K1tKeVr9B8+z5sYngGhnkJhLpb9e33EYn60o9+SkeSG4GD84H46EouRd
5X6WzjL1uNBHF20qXWmMTTp63Mv6wq3O01qFxJC76GsWr0UwnLhDRdRKt5XifJu9lYju/Wy3zNuP
zFSwujge9XTYnlKmUJjWcqASxlXYJG9sHlMiNY5oEhSBrFBjtbawQBpPPqHh0cbO9qxupzu9Hwz+
saFkx3Lka/3Uy+OvPzTSut8W6YgCyIMGGbNE6KVZqQXsE1QCA9cPrIcIVkl14jTfWoAq/4I86h9K
FVVrn3inKGpB3JREM78sHFQK1YVWRTXH4L3zgD0AAlhNdWe/1zyp3/zqcTJJdbRdTIYqLDJcDK/I
TnKvoeegp5I04NnNlkvzSySMUyTKRLcjG4E1cMyJYtSmZfYXre9QUteB9CQ0PPVL7PTgpwOHBBo1
eldtFQ9iHeQc4U1L/RFw+agsPaiQHy33LhYuz+g6FG57FUHceRcOhWsDBaQeOSF7CV/Tfjcj0Psl
fX29l6RW3x1caaf0kSfdpiu9iPFf2HjbLbOpbIScQicmdiCaW7oyST/K80Ev5rxPYa9JeKjaDEFm
krbYk+c8Rzl6Dk3fzUWSmgbcg7Eicafsh3sAz9J9A+Dd1qgBG4jZlU2+vRPH7g0+Ye29YPFprv4L
p/zCUbQiO4/Ijvan4clb7+sjTEZLkT7s+JFhsBcDyuTcLs2L2HDonMATZrvdxPryPyBUp9D7kFdJ
7klyAiFV2BJt9pgKKylgsR76S4Fp21zWvtgD2tSOpaBoRYy39SqXtd0FFx+gUVuA567vfdMrfcA1
I8L3/w1YJ+tjjdntQSDZadwKFPcAW63y/36bbuZAA809OliIRKoGn0E/50GEar+bLJu/ZCfk/tiq
8v4tLhS+M7p9IsbEhfh3FMZqml/XUjU6oj53c8P5tFF2tdGTtGY4CbraWPErOh5f4t7KpSSA25CW
uBOOzceRzfZ3J3K+svLGTy4qCdoZw88jjtzvEoi99xJ8vWVmihslurKwrphGzji3+R5/YmBoRPe8
yVgttjhjP9P0ijQVhG95+Nqv3qveoOx+KDdotQIaHZFGycgkF+TbRPhZ71rgsCXsbci9ex4iHyIp
s+IhcMnN5EXIwNzmc8/zBW7uf9+8tIOxhdzXSSc3qNTMtGQVb/RNuxY1sZ3NyPFH0eU5ZTKTk3vu
0wgirYaJ4MuB8lG6zGPAHoJvEACh1+37d2Vu/f6l2dcA4wvr5yNLPliRd+QEbPKYgdWXX2HLD4Qv
bkk8LyqzgSxT7XsdVUHnadIfma5Kmlb9ok8zT+PX3B6HkQSS9D0PzHw8PXNKgLhey9rMsAv88Iat
jNImcWmfpcDqSkuGII+5Jb/LfyEBgf3tN2UoSsd0h1GzDlBbYH6qGGKPKw8QN/ayLMugaoeOjdhq
OWq5xbGcBV8hG7Yeb/1XU3XGsyTaVO9sCm3WwkXWcMiXHhBwMFxFbYzSvnrK9N/DEI+vyNUlGRRw
HwhFf+9WQUvmUXm7rEvcmwdBh8qG8VsRJb8GZrEnxH2V8KsHZnfgQyyCyxAdUdU8HLFvRa519XYY
DUuHvBkiTtWbTQwJLlQxTQO7U+MgLVsnxu9YfG3m1n28PmmRuwQzcKssHQcScqY7v31JVv+B0Tmj
RKXPFJRj7iQ9liNvBqD5PyVdSERcshTWmyVXXXIaqarbgGcrq/1+UXlqZ2ylcXQCTar6mNxzAmKJ
eJ2axcZYYd44KMUfxnVNfVnyedTWyL3+MKDMPajD2hFq/SxYuxPDTOYx2a0ilTPLqH9Gnv9v+P1n
kAD/orYG5WAtYnXPl/fk36nJEKuqIdf3hDuD2J20Ig+GeYUa790bI1rYi8f7TpWe2y7k0sfwViTm
JXWg09/2SofOIRexaXQURU828PfvuBdTSGAUO+xeoHXyyP4oLa9NPYOR0vE9J20Gzx7ufJ+JEoog
k1TjWdlHcckjBWU0bmGaG/Xj8VSabvblQ2D5E+dVNaEK8SMaLHm5IbdnTpQzf9TMNAgcU0DIU/T/
z6voyOMz7Uoyee5Z04zoxLrq4RVIl/UY1ZI3lW/QfsGoOAU/CfCCK2INpNBAZbSI0woo/y/e0B5N
FvWoChgyOKOLmJ8oK1eroXGw/kga7ce0bJ9unEPTiVXUwBKCmmr3mBb9nTAquy9+dySkZ3XBTRes
WtNb3+fWQeHv1btOIej8lPfu5dqH6qCdg37FYLe49KWIBe0z1z49bXIFLx/XNoXICSgJ2NcJecTz
mwbdCA79avqSK5e+q56CcaSQQPkQMlmQnj2g/cxb1+zci0EQb+QGanYbf4IFJqEiSVP2OumKJ2nI
/Co7JsYre4RA20/hr7f/m2GmX271wjJU91RNFuz5/J0CSiAUByVxEUXyUuwlTEoxlVmZN9OxXgfd
mN9OwkJu2M3bjOr0xMmEmUUUKc4XMg0hoSv1bbR+uc7g0BIMVWSl3ldl5t7GFANofZX4OLpaDeLt
+qegX91iUnjeZkcpm6r58YZKsHjqOYj2y7rr0RlbdhD9hjIP1j8m7GgP4BUDNFe+eL2dvo0LhAkv
d42jlXtH5xUAOBaZJHLSHfnRGjF8100emcr6wzD2so4WNathHQSD0JK9Ydekd+572PCFowSnM6So
ba1dMm+zgOYHPTFsChSPkn7bv0hKUNWoPf2C49WVz7066fyOyY0A+CBmr5VuEIwBrAOHf9MJxpfD
zBbJ7gZYrn98LcvF+6Akc21v0E5R0U2enJA99SXy9TDvIL6nNEOb50F/z+GIJwruptMLzyHCaeX1
9XLL4ps8cuYYuS5GUmHcySq3CFTmzHqDLBhZTkOD7CTc1lUAW1KLQqNoCZp6qSgQ18FNmnnfB7sM
ojRiUpdhoaau8V4N+z2/iK6tXD8YZtnq7oUPdPRVrZdmvyGqsPq5sus2FRBvRBP1LB4pJzWw7GlM
kJ5PfkBA3QkQ75dU+Eq6vWiNMsNfvCGj1HfJYAyszBz62P4617GCMGcMmYi8UwTQy7u2HzCUCK50
K7dowIdQn/lou1sATqHFyH3Ddq5CVIg86gX6OGnmz1XW9ZQblcMUeMzVj7wy+cFHJnzsT2JRLil4
e0puOclfQ0E4BLec1sR6NmGzfBPohifm5p1YuUExzW9T5ZxTNh73Ge7rFoJ/nh0Hl4ezaKC3V0dJ
umJsjNHqFezoBoIvnryfoYAa/IvmiViksKXuCvcwfFO52muv2Nw25goWGL8LAfbEWFq6u3PIwqM7
4jOYU+Q0Xtw8uP7lcB+reDIp4zXvdg3hnKFt/aZrJwXaLrXyWijVHgpzvFcOkFu+h4Jmpe23qiI9
PLjxKkdMf9BU1MfqTyVQfrFG7/H3+sLnX4omVK16hQsqNve+6GK45zIY6qxBWA9aOyKnOP8Yp+5C
6DP/IR5XH1O5IptSro0JVC0a6DzWyFN41F6plSjfywRxA6moHhp04RRdnwm/nl3zcp5Kt0SLBdfp
33480Jwsi+sNXI/yhQs7biWiHIqmiMYzcWDNrYuZq2IVJ/1yUXZ80B47IvMq4uCKTVBsPIfmRgnZ
aYOR2s535jD40QMGNu7wyD9n+gz52srsWyZmhWUWCk71ZC2ZyQSyggM0QuSbnKyOcJi7j6cyCbyw
vAI/0XxhZX5oSUnm/vTlR2MgFinaic506aTcIDwZP3vE3nRhBlqvMm87hdM1bvBC5tsmvHjXQBJN
TVsZq5Rlu5Zx/RIj6smPL8AGaGRPr5r5nbqI2zaZJoCysj9XStUm04mFQzd5YLxnNM9z0Z/a9O6n
cdOvoisjJxxfophJ2AdT+ziw71F70INePwK+TK/6FqxovLjVd9Cnpda1qfsVSS3ijI3y0icEgyYc
fvfuo7ZKQCSjNPWigDi1RoFAIbK9qeAkMnQX6QpHsqs3W9IktmRgLjCl5f/fhMQGSoF1DqIfLavB
Okv65Y9BSaA5s9kC1ki948452HOAQVDnpgOv7i5I0eLCuP7jBNZf5tckxn8lli72bf1VILpndCf8
4u5PAr1UQfh+kzGpflFf04yvRVYB5vUQi+wT/TwvMZP4eJSJHEIKOJQsHttmOroHYv4YifbkK8gR
VCFXN5Oa3H2puTn68uIeNr4lrbTG+2UH7OUCQmOU7nCUTgtvKVidSYS60Hkr375uiLsf8bXbbhnB
RGTvXBG9C7jWxaTowULbT4qG37ARCdWbUAoZgsr/iaFgc5cQzcrSRpo9ZcQ5mq7COJhgS+IY7xYi
614FStLOeNQdfgobUgVRmUdS4aF+D3dud0dyaPUeZS+8KNPE2dmbuJiaLUThd23Et4RMrldxO9Oi
8iXbn5tfNna9aZVQroqdLGVuJAjeoqcV3WLpAVZaeoGn4LBP7tHYUjnfcnK2WlFxTel5Lyk/ptLF
okL9EG5fWyKMqtBZPE8LyMl60RnawJ2r6fqOaLUi/AM4SYZIvcVahf1sQmyRlVxGM0DBsOqvjMMD
h8GNKGJKiIPi+X+VA2Pwvxj1pMrj/bYSHjsk8yKkxFv8p+h9qVE4o1YwYWFOPUk55YgNkUcBL54M
XcNdaKXmQ+Z4K/woDOJEoeJ0sKK8RH1bOQ1DFeZUTjQDFre3Pi84kiHzl9SVlCmEFoL9DHbuyDii
BZGwmt53yJ1u5tSwWTSawqnCX5xExET0ffeCQkkJ93ke3qHwj6y1p9VC8n7xQabQ9eFW6bGpS2xD
tzdpbNsk0kf3HHaQWA/nW6r3XvwWpuDjknB/FdM2BhquXs4ZkzdHJeteJ6Vnk2ihS+mKEdPeYea1
bZPsqY8ePxThrpVbxZIAbvB08ygHRXrpSacYP+Pewwq1CIUdE2y3U2KHdwWE9SmMubntOU3Xr0F4
A08+wtY9GygxXarg/kXYkNGl1yN3fXJeP8BMMObxvOlykeuN+MLIzAD3lyoJaKnbM/GESlx+yld9
aysy1KcYwoshSF4WiV91MOye+iAcD6/nRcDdkBlmWEqu4/EIIPpqwWxmMTbWR+QMo4Md1aIhG2Ig
tUM6s0AiXhfIyrNXRum9mn7f3KPQbqBA+YqyXZqRr+4DSQY/dtw3vY54IXQGQbdAYXIXRHHIz4I0
+oFvIwFW9pucT7cYdMzGuIoxFHPfFJiU0Ud9CBBObF/Qr23rXzR/RxtTmQcq+/A0ajH0xbIqXH63
0DhP301937kwPcOrazF/IslHswbZ/Pnummi/TNNSTLt2sqTjnrNQfGOOlwsWhHRY/C8+P9NTQ6JG
OgJqdHYn+P+2+GsJPalFBIgtqQxq414zCGJsI/6iyOy1xQfahL6atugY0NlZhYFheDmgmsInJtgv
rGEaoy+GiAeaHVyD6eNYwzrXOXYsSHz7FK6Gyd5KtjxPcI7H3rRpTctoB7fJsd16KxgBm+wYkhuh
69YetTin38W7TESbVcW4JtOavBetc2BeCL7IZg3kxAyy5PoMjYYzIPPqUj9rTNbmhW7M0wMrAjF+
HeIkPrAl79VvzfMmP116EsQPkfAqHIXiNxby99rAmNyEpRDMpxkNFWwmjtPIeqQgJEkXYK2CB+F2
C4+N1s7/NmxFtnXkiHypnVwplPWPxX6UWk0exrQcRH6w6pkHg5/qT2eXUexvZkgL7xRLYxFEZj+N
awTC9HxScw0nPFlGGzkYWEiai5rVUrRNHX+QWYMap7BNPITAW2MMLrdL8acMqq+VfLNEcckhk+z3
9urn3MOZU786AzmZCKcfEXj2OkYqFcVOR5PtnFLNOFLFdrbj+Tp0/7IIrggV8MeURbtKut/Q8lU4
7vFeinhbvMGSM0/dO1emc82o5B42sSSGALMHZREtwotyRY9qxXYou3SgltiTUX5oHWgRTHUaTwQY
iy1jxss+ZWHcyioelo8VsAxAVJSjk+UqKwc8iq5BdtN9CsDLyRTn46JudC9HK+tFp7S3uKh79Dat
7aEo7mHmEEvel+Xt/k+evJcJ3cQun+kOoAynabTmflIoyjoLXX6nKBE94OQVdxHwcoVxhww1H2a2
an+7Nd6Wm1OP/0s13KCRG9Cfuwe/JVnzU78bys6MG4dh8NfwM/CEMHClvcwG/6PLKktjdQ4vRZaJ
V5vfA4dUFxQorQ7beHCcocklLxJ27P57i+tK0ozvJ56KQBxWHtU052ZLBBJDCyXVLLVbb4lSDnr4
irQ15H2Hz3VylIUCuZUVkA6aC3P27diIjS0chU9RCoDiJrnXb9AYt47Sa3ucX6FYCNY/L67nAvti
eGcx/IWom2/nui4T/zRGj+nFTYEmXINm3onW7Yq2sFNh7M5oWSdtmZW3ahKiOddKZRXDkuIrawYO
ZfDikKhuz9jNuafTnEmOkzJmjVVvJbnHvdqRzAAHMsTUbMGLt9T1rcMht5cWpewySPbGoNEeH2jS
r0AqnFsXuZNBWSTwS5Qd42OvLgpZzinX4vPCv3t+ljsAsZVO4fBWueFozMmHk3SQrwoUCOiADL9E
PDDmPd6dhMQOCqQhxPMk5vvJcJJuTW3l7RKpMyhwY2XIhdezQu4l5nreussjHMoPUMBSr+5gZvWl
M5ZVCi4ftKVncPloj36FuPyCsKulJhOHzJJGOcb8JLFtpJZSU6sLHKtoPtaIrmU3FGEeTmoQwS/n
nrcpLLZot5gNmGZCVD+F8L00Jeg8SBV15BgYSJiAKDiIrZKLKd/XOrwcOGuybvdqxI1YubwbSVFM
4qrzdZZVK0Re9Xa6NRab1rsf2l269mZtZTZHqcCpdvHYu5BhvwNM9FWoRSObntM4eWzwbI+FVQ2V
C1yyiCmMZg4nmCkziF9nZ88ohFyrXGbg6H69urcXcz8/LqI/DDxhKnOYsYkqgnH9N2+m/mPRhCEw
lSDRZ2vWqIsSXNK8KhRTzHw16Rv/e8eCmvX8D4tuI5hG4lPEDBtqldrJFSfiv5JGtKj9Ha89RbuG
lKRofjMihvubFqpjj4MnbJCwDL3caYogY7Y2bKkZf0f7IcjyS/+cRRGTkuZxXV5iAIER7TungWj5
BDA+skpvjLQjwZU+w+qQqwrwT6ndXvuLB+igFuzpGeWD9xzsLpm5H1M6QnGVyX8RG3n2tdALERgB
BPpZ3qe2Kd436LO1ETTPv2f4FSgV6QXW0S/Pm+Ax0T9UI06owg7la3Upr2xEzfR2lIL9U5d0NTeh
zaDj0DDLo0vSY3cfDdu2gl42psoo9B46MHhkhsUAi7uJJoMYDGmSDwXCZx+rmHibbomgU0vcy7Ny
8plXLVPztxV5oUrZKwh2IEqT7qXmXtTC1LAWk9VfSrDxmpOTl/ZSwVCHB8Q9ZUSOtXSFtEG3jicR
33wW4WukUjqsoSP2pX2E0YHXR9mVH8iyHtaUtTSZTiLK++QJRoCHUgkcbnueIX7g2sjKdS49QFsd
F5jzbN1/0GaV3UuAsERTwQdnNgYUmVl87NMk/IMBZ8ysqvNpDtGBPVYezRZYNodcOSlH8V5EuRT6
FjHM0Qca+7KV3h+PXejzSMD2wsYHCrk3hxsRPQA75qZIjDskpVZtbyff55ncpKAi0oBSLD3JewaF
Vnjuio+lutRcePhwojYj0Z8MCZb4BxX7/DQU7KRcNSJzBRJted7Pe5AIPMWs7lJj6Zjp4jcO9Xyv
1iW5ilJgjcZhQVSLMnMfAhyd/IHTkmAVU6p30CJkImBa4lqe8kN7lMFbJuhI9Gpl6PzqsaACmeI2
kI6uD++6G+13gybPSWdMb2rkpVcPxWenanb4JBwMlOPMksclqjP5kIcxEngnDyX+d+gtAxB4nizU
Ozd3xhFU0r6kM8WYyZf549y4u9Pt0oGxDP7LYm8g6ZTbqBHHNtJF1t9at4qHATr8vKzSkD+jT+uU
OYFR34CHMTwqAh9HBBdpiXphAWmNdpKIO7Z+nntWyaMiRZh4wOs6pWj20XB8tG4dHtcaTq1Vbxt2
iCeJ1C0cuvRpPMNnB5nfJ+sqltIxKG6iy8/icLWaSIZC0CFUgXqzmYd/ZaEYN8SQPnTA2ctYBSQ+
3pUpjYP7y/GgGCav8W8H4dGq4pdEKEAcvzfgYD2H9tpfGn/jzeZRTiD2ALWDQ3dd5wscCAP/So9F
jGU4G8JUuXzwtBmcxfmaFSpwS1tmCWGBXpAIagjxcSKTmmw5wu94i1N1uVVocYLxW4Jw5NNh3e8q
vclE9V+zTgxVjqTDDpKxCE34MPAiJkKioR7D+yLWRBQxwrEEHZtZHx8iEBXUNRXMfrAQsRRapUtT
ilEi8TmJwK60zK8IXNLFWK+SGfYLX7Bn5XFi29a69+dFZfAAfhQ91Li6gn2RKuMYql8VL/yGdgKT
KvvGdGXbxV/rtx6sCQ6FX4O+/Hfj1sKgdZ/tATzNbrFVItQ2mnMJIkzJ+Kuzsz8hCfO0ugcy/3uH
/wMa82Wi2Um3aUwcUuAbH80mxY8L3QkqO4IE5EO/ueOhJmjHc7wYu0wwOnUnPxIZgdgnA1DzGe/K
95t0co+dgc7gvr1GbfevfQvXFlUo57u4Yp6uqKHo/hqEGTC0Oxm8Tr3FDrHgeSDKdvAEXuNDw8qW
DTlCW+IStqOPEDdAlHRUHzEyg+E/RvfwH4C3pBbfBoisD7iMzGqcIOZCs9pFlmOU+e6eS3TdU3vg
yJ194eQ4+adol0jXxz2Qp0B6OwSJCEYS5BgLIZ6kykUB0IY5KILrMln89Uk2Mnb2O2pdQbGa51Fd
YeAZJGDczF14EM7CJokig//vkfp8wxd3EfDVCPpcRuAzN+ItBuS1250Ex+lOWDfffJV7MADJ+77J
ZtMPHdF3ujGEh8Bio8qkR2z/X1lZMundIiiFwFmXoBaJ8nSZTBgow1WNOMQ/6iBha3rnTqAWdqa7
Zn6WFJy1EEvC2W7pB0B3lACJ0uZ+YfCGNSUf9tKdtSTqk3CQ7SiM2wMs6DQ9QWR6EJARnqlexPO1
X5jiinja/QshsmlG7gKLD3yVNhdcaKnjTNNq7+6O96HaRhfiw/UGF0cKyfn/OAjCBo5aCLn15dYf
BnxF75Pl18VdeKD0vLEEzVpSc1y1Pmcqd2p9ufidnwb2JP6CaeCqseu4naUMLXmVooZTO3CTJtiu
QAGepHzIQ4dpjc1ryqU6tTWRPgLkIrAHWH4jzU1yx6IJVyrk/Ajwzt4k45X8oFpA0kIFb6cEJD+0
LIQbnGY0VVY4ojyDV3dwZijW3T7TTexk0hQRvE8zI9qB81svG6cZR+3YTqOcwug0rnwt9L0ZmqSZ
Yt7mlIlDHpKz1rvUBeN+YdiCDP1so7AYzII0cp8xZoG/+CEBTWK62yoMrFDJcLcl0BYVhnUiVlRq
9CkBAj9SAi2kHXhhtJRDOeup2awH5GdR9yfMmXESqVEk3LXhQuL+Ov3MKYHSLShX7pifiBB6/Mw7
WMDmHUyBMakjSHi10s2kt5uR5b8kFy4zYvpEOQuLwwJbPum4M/PHXLqgNY3pf9fnCle6mJ39LGuo
Av0jeZZF6wwnFd/kxWTzEs0RAipjnu0T2uj1hR7mPSGid+snjnDDZ3ScVejcyFDVwPEOSU70j2Nl
C59KskqTERJo6Z5kyayZeSFP3rgd90IopmALuYctm3opcdeRdNzhf/zX2cAMV6Nh3BaVr/VLSm05
co42CIjcbEp9SCNAAimt/vCqUUae2nvgRnY9/HnE2OU8RnQOS3KKFYnIAOvbmIedIOmUQiHYfyIT
ggCnIaxHgTcpbYKaxuksEo1NP2NdEYw8C3O4cs5VgFg04kjdQDm+Bf4o0qZajQCRexxt1uwPR/qx
f5UStTkYq0YuweLYK8ObGNq/WQj9EDDV/At3YfQZzkjgB/oA9DRqC+ESyyO+FmsiwoATU/BKaEjg
Pfidt1CWr6uzM9s7m64/MPDRvKGi1bEfO+IRF/81H7j/EVkrJ+9Xxj+xkoxNPZwWDhqRvuU+JQnw
si4uFJQBc3CM0Mnf8bJOohx2J7ut1nBEFzQIA9yklfkfdoV5rky3MbTmbGOANtVL967+lbcao3L9
PRFlBkP+p65nmhbM7cakH+ej6t1aKFne7KOhC7TUNwBxbtb5soqTThlcT/zegTb7xGv5cDyvCZo4
Y28Lhn05FmjKjw1qVsRJpUtAEDcIKXOId4+szbwekWhg+Q8DYaxy8GBQo0SLvD7UdmVhcPLvJJ/2
Uk7uFZZ9FVLM9A2JahyLGqMdbGlqPvjJm33bEu6Gws9SpyqcVBpESmsQ3mlAR3d9xn0zyKteQcYu
bTYe5TqN6CJz4e9QbhkJYirp5R1OC6SPt41ghgA6lI41HJa1McdOxtuQzMgHYcL8IK/Ufull46Yx
zQAZUiIt3BsvNaTQMcmamJy9+23FFCmfA7QmQxdboba436LMpF5I2pssByXksinFczt1gwNaH6iF
m/bxjuagL/pLeHcXiu4KbE/ZeFXw/0jPKlOeJS3XPCABnwXqk3OeAL2ReTHF5l2mP409CO2VJJ8D
H3P7RN7RY1YMWmrc8n7AJVpMVRNskS81GTw8cKniYoww2riMGuKGY2f4BsoSAGz9ne2yoxVH+7a/
vz9qZNfIEbRYLFZKLoFUFd2yQiT0KNphQGsfTgyNv6Xb/3UbWcJKElWmL6Pv5kqIkN33JP9S7eL3
LE85ZQT+0Y3YBzNFPqsUie7nJ6U7JHOFLEDPE30JadfC60maVxv2oPAdp5autBVXyfcFOAeCjr1n
JlDQ3QI7cL5VYfM1qHaIY/E5QfxfdHIlFhSQRDWFfI8lkrWn9rD3abenv9KTdHfjMKTJXffy7nnL
UskrcCBUJeB8lumCMO/dus+evLiA7YIgul/62FmihvmINxoTGlJs+VWr8WWErRhb4B00TSdFf6PN
D2IFN+n7ROK/yMhZTPTxJ4To7XJ+JpQz+IrhqKgttijGyj0SClkSzg8zu4qnOmw0EWKp1OTNe6jl
rTN3UHa0hHOWr7C+9Zar2cCcbyBXPOjhFRrbH699KnjXBtwHCv0EDXTzkQCxlEiowNr0trY4lje2
r0mR9QLpszfJuR4JJPlALwjmkkUglgD9du8KfXzG9QCThSiWg6iZHTj/s31m95YmBJwkygwFSo96
quk//ueg8XYcrVKsHW4iM1YOGhHMsRcm5Nd1TCBzCPnLGqy3n4tXNKzgPfjq/j80Y9n+yqUXdQGG
bym7xIPYO7c9Ja9pwqEZSNER2/lIQAC+sihyj6wTJjf0FUDGg0Y1UMgA70tHHSt95X5KHzd07X+r
BsbgSP4OZBh9W+cYndn40I0IXDy4zQR3KqGtFsufRa3zTTeOLCu59SW/oLUMTZsjtsHN+oLxfbpJ
Tkk6wIu0u3P4On6XEojb0hXEmnojsStkYPyNEuIvzlQIewYh++xNx6cDqeU1133iNMZWghG2LEWD
G/9EI2x1vhpwnzA7Rvi0p9htk6Sl8siJ3fCKNEgFebGVv5rHFFl4EFPUuDp2UiCx2Qfm1tW258dg
NAPgqLPZXWzGl/EcCJ/QaoL4juH5W0urQJFMLM1cbGwa233CAF50oJCnHsHYCTZnU6qhES/F17td
Pqn7JOqK35YTMa25AM7+B5Pj53aWwXFey113HZt4uARSkudRKSP4DJaIb2uoaL3sgr5UqamaxdOi
INQERegJsfLJtqUEb5pEzvBPQjZiMAit4to3/uKyLHhmGpElWLM/RMfP7xbZWtOikCAX/BZmk0+D
pUZaVd90fZQKn4hjGM9PGhM9zD4G7lLzA/UUujRVpLySbT+gG4gKLp1fQegJe1iXAWN0U4Rw4J0W
QOm1IL6FFFb22MazxbhH+NsKFBSpPWPrxyh4JqsmGgXNil02a02Urp/YtS0PzjYiHvANTde1W0bj
77r5mKjoWLm1o/3lduAws+QAqOELFbRbVuTDAh02A8UqE/f5m9Zfa5lcaWHMv9lu3VDS0e2cH45Z
qbUBbGzNMHJCijbzDfQkJCluICxEX7oCysEheyNXpeXFYXfGdt/lwGh9pZ81cNCqOtMCeM8726l0
CJGQ7Vv10SB3qGEacd6qjvREjIF0jh6g90Daitvka6nbswuUbPnHxBNisVn+S+oa3LyI06RbT52m
mmPw65Oz79B4AmVD7pUBqgOr9olO2pFm4Ar6dzEGBpzbD4S6xceAgpkEgjbfMH/SthDUR3XyRahS
jpcMgxoxpMjcU0WAh1UmGHw1HcIeMdPgSLE+fkIY9OHYNbBm6x7CrSocgYDnlcRAXLR1NkjrRscX
W43UV0SpMIqrj8ZJVkvlwM/ywNQ3jut+KJqAd5Hbn6p/YRrhZZzhhy+QxDVya9iba+qjWEfrGZic
PVX5OWOTJnA0sXcWLqNGA3HoOb8SeNPDxD1V6VDH1gubWYCSDmdlKKb8STSedk5bBnA7arzli6HL
LJ6tvssZP//w8MldDwW+7d2f7KOxCiNRgzpQDoBAyKwdy3gkOm5P5kev9PZULpyVT1bkhFj+8z/U
n8KybUfexIuZ6qjRMSd9K0D7WUAHge6Z5SVEc/Sg3TgZIVbSJToL0gh3KWKKbsgSh6HCVwcaUGbU
PH5ecL0qBp5NhL/ir2bd4r6bVJgJJOvGK75jkKC+EZ7IBl/4G1Q0Mcvjb6msBlhBvqOuCGzwKgCa
2lTjnLNZn0jG+LNhuf5Xzm0JoakQ5MBer8hhZ5HKy3sKXY0JkHJ7M29u1GmbkjLxqYI0BmzUIdzg
nRj7mI/4V/5h966Syz/yABq+ht29GkBBTeSuhHs503L99XRroReECkoYSyICcB1QLBywbdHwYcnv
YTX6dAFvjT+BHRoJGabZ9n9tkDg/PukSXZMwP0eD33FkizP9lGRQQxVQw3/UxswkBnLBmj7uKmqW
C4IU8qzsViMgGw67n32moiJ3g6fS841XdWR4ZrJf4Ruw8ex6XKFmPmtpZR/9NpDZZ9QmpuR7KWlE
WMWyagIlF/756jkwFPzDcHaxoWkYXiElpPDKGpRY6EtlHJzeZfsHsI4hcNUvmNcFeV4EO/2YBaCZ
6ao+oEtxhO+x6hilm62ej6QgGMcmo4Itpe3aDlvxnqbFzxe/JnuX86dqdqpHkgkkQwj3zCtU/H82
5TmTsIRhKM+YiWmbN6uR0yetZl0z4uGydwYfkD5CDcwKIpwmBXSOa8pdoFGtwuSg/o1Zk2vpkSPz
VcOknFYfq7p37k/8fNWcDTbV0BAwTYXJO8YMgYQmbgd6xUByYNOsJ7oYgab2XSbfSbIOwTtlvj7B
9kDxAGJqbtf0mjtGDKo3qS+EIMZpoC82Zx/WTuOjUSLtM7wtMQd+MVMnL5QTsXBYIZHbOfQasM7u
RPpF92dUQbJCegFiHU6OIpA9S77uModNhF7Bu5a3+Wx6n0ve2OAdCFby2jlalLyV+XIinn9+lTvi
vdkTr+1XHBkeOMx94tbsm0/hmg2wZgNMAWATws4URcbX6Mm1qMWlNPHvvrQqlWZ9D4k37ltBXEfg
d0r91dUpwtCChGXUr0kSTM8u6OAgRZp9kUZYJKPHHoIP3/emfhfmx2CaRqJGlvvZO6h6ouN2+Ui+
4jH9GK7grX+pdkQqCze3W/RoVTL5v7Ph6ZeWlGJ25f3Ugo1TIhP3z6m0l7SeFy1t/MxOoxqgKXs1
UBd6Wq0NIbTBU0G0BuQ6cZMZTOQx3CGeinWjBqYyyLdiLxYgL52Ia9goENL/4qDaCZKv9MjnGYmM
NBaYnX3eUh284jAmy2ohHmGol9WHF7yrQncOVvYOJZNi6RnKfauSgT7iaHUUpEHVIhlZqGFRpW0V
jn8/cHCOqnJOQiEr2abNJH6TwzMSujCXTfR9adz4xWPy729LkzoVeDMqH6EYwSSEmBd71rcC+b/p
2DVjP9vhx/wCDrDeM2oJDfoJVIjQzfgdJkg/uPSoLP5jwFb00GyCHtN5sIZ5mhII2dq095SGw0MO
zjuBMwJNMqa9IH4dWahJmiNXq1dzpl3Ct+ganlmdg6F85IFjki66thYiHmJECuPMpdFCKy9pHFMm
Gd+d9HOBCQeOm9cmqcdCr4kMJQVhzkmA18VEhVan9TpGcIQa5Bvr5y0KFGdYWogXNIFFni9VfQhX
0pfdiXvxoI79JQK5h9dtpGAu2Qp3tjo+MPU2sjthLwGoD7g+0h70Y89GeV3Aw2PuPWBeQBCq/HIc
e529OjDrdbSywbAhPh+AEjOHvt+3b7MVzmiUlzLguDSYxaMmAnG6HIkYK5dqD0aOswVaOn0bjOhM
/VXQ63DCzyf/DoLgsqA6h4DwW6L+RzM6rTnJgxRstZvfVT/s5eDWed+Y4laEtQK54IhUxROX0FM3
MrIctp8RrghLxGO30RImN3JXx1JXifp3NTR24jqyrxscaO8/Ne2ICz9AoflfhNNMvABwPDxX5O7p
1TC/aPzKizKG8btY0Ri4L4IFC7NLFieZRM2Rcm/yYKYhW+oipA8yEoVJendmW95NIWRlZZJ0wrMY
FMX4fSYuZ+LaSiUMTsD1cAvIIWxGlOKaOizOeGkyKp4XQY+ms+DPnWbb9I8G32TintgqklFXcLqb
TOSgJLAC71ociQUHMU7653a+viP0Gc3WqnZdzvZ45wjoqy3JPAeW9A9NLwkzG9Z3H0Fi312cCgsH
JVmFc4RuK0Z2Je7/YVQiABCD4qezT2sOVMD9ejDU3k+//uLUzS40aWjuYh6nx67YMKpR+UJNycV3
jVBSt87PLpfg+GhMGZw3wg52xOUsEcDlKHoyzwxZVIcBwQ6C4ndc5r9MWQ9wtOZqcw3iOXGLHH3b
SiFLypJho1+gTJPrh8J2FiTX0zc+7+4J9rXCwXVN0TMMjQM56UWFj+qhEWa+VBidY1L/cDwdl3Io
xd3Pcm3SnDVKaocLjd+p9DeiSsqmyl4WLibkrZdbXc1PlaZd2nWEesqJXx6uAvkyMXuWStlqtXVt
c/OxWbt8TIc4MDhpmhYauen2ToMjiFuPO2td63YQErhQyL9qas75NCdCPHz3xy9hElBn1Uk0k+Wm
IHeYzTRVaKFIJNk1qGIcmxLLtvZgXffH31mUNfXMIa5CXhU8mXU274sp8eaPKMLT7SSjiPTbqRVF
dvFAWV3RbOEy1xmGXpi/Jwc8GID+YPLcKcl8+QVqXNVqQdlGHrtPdOojj8LXlhoEwyt0eHw8Z5sj
Tu42YthI9UhhTGpE9AKM3ZxunprQrJjneb/b41QlJYKXP59fjjPddaeBAzWmaknWZBniO2S8gK+5
bwFL+szgmxr/FENraZpYWIP0kT48a6slBQO6iwdlq5nFzY6VeZ78yLjRhT2pA8F/EQxZMW301Aid
0YYYoCr/V8p5XYK6rWkcG6kwT4o/exyGO/EFruplChrFcAfDl9rbI9k3mmvGueyq77M/uHrNf5P0
RpazWzbSez8xOYTlaBJp/mkUsSHft4/645KqkY9PXeCm+h5bBiPtdCSycdQDj1jx+T53Z2d3fKDv
Nxos6mQX/5jED0vEjEuq0QIte5tM8ok5NC2WXgaxfrlXXxaYvkFakyBVrG1Z4zIGpDjchC/A+EJz
oj8kfS1VxqjKdeAi11JlTOaHbfxISsz+FvVGvefwSIJIbuCA47cMXMXa96e0KzEYxUIAK7oGJ1Ll
ALY2uA3n/eYBp/rThamsvli1UyvcKL6bDh+BUHZX5epE0sFVdHTygKHyb+npHkaX9H1epEOjGLIY
G0M1qzqvaO+8VPdRnhsTDDhLoHWO2gzd5i2hrSqOomjtzLa3TxqwghTDNYIeUvLmKbKvZDbFfP+2
yO21xvzFk/weBsbR/PhRMJYat0aK0fqml/YzdyuzkSwAM4OFYY3clkrullt1KZnExFnZ9Eg10sUm
IatRHIY9Ib7cDGtBgGBIGEqb2tjsvwByKFAnppwWRvQsH30T6kDv81Su1OdxQWPMbG6MikWIo6d6
FpT+qdHU2RnumQy3yjtoduxU5SybU4LSeO8K+ZxtSUBrsEo+DKiKG1Zvu2HKnzn78Vd9AcOL61fe
Veiey4/c5V8IsuwOJtWKMjTPfFGn/cALDf6xDKWDZTJrRyU+8bIW896rod7Uosld5pDH2vSlBvFR
0buNmHw1B2Y7Luf2sKUwcDmkdro7s2Hq6OFHmNxFLsG59CRvq5CIdpStYac3X1luoC580O14t7p+
KCApy7b2OwX9nPvEQxrSEfgqbORQ1tC95zI2dIm3VklnzB5WRHnI0r8bSviV83akkgOGBlaxVc36
yhBJQaJtf1/JGl8Nh3j7mvodpciDvtRsJgEd0UhtwWFruWV+ixaElwZUIgCtZI0azZJG/LQ3tcTv
3IpAiKDV2msk78G5bAqzYvbjYyRuZI+75VNUDmSH/GZHnufSPr0g/uhebYHBf43CxoE6bSZ5JBWG
K4q5QFYEeY9fiXhXKYlXa7DXTAv2JJY7kZI3cWJxf7zbxXJ2nLC+VyZWkzapRLaciI7KqFgZf7vo
l5Sdq64V0kEIXvCcRp6syJU5XI0sx923OoXPa6+DBKoXpHGacXU1BA+ZAt7UXapUYmtyt/XQspTT
5EJiCH8cPacxQXpsFLl7RC09aLu/10VY1sxpBmKjCuBkgRG8Q3DMNp/yn8IuxPclSde/XjOYVgEG
F9BOXfu5TaT1TsjT7DG4qC3Tw+/YzJShFIXZ9Ttt6CAsmRQ6YxZNQ2wCwYA60gBaYaAKOaJQGWuZ
5IS6Rv5mtM+maSJ0gBxALWzVX4DbfwMeKvluFLbZ8T1Tjyl3J5imzrSB3qH5n6eE4YlQg9ioH5Jw
Hw/mkdqVRgFUyldeGarcRiOfOvHvdhBFpsLsaXKXYFeEdB17AjIfxH8sY80PbF21WiHRbqhy4bou
mMXWdZbl/jR+O9sW0q9zrl7YibZpdpUpuOTlCGkM8vJlbe4nA3jFHODQwlzUFbrZgXmjb8tso4cR
1VjuISvj5TSG/7kesljeKNqKJwEGMYDS6fjWx2vwNh2FUBsCv1Dl6dU8Bv+333Iyae5lXZSCPLaH
9LJuatccp6Pij2tURTCapMkwNCi7DqN7A5oMt7TPum8jM4MxUNNctNUIkqzoc/xo+5SZewcZXbs3
e/jf6MftoLPLHfEvPsTPSJ07YciWRiiBaEgDdDHATLZ+nP+sF23FuUrqK9GVWi+RWDcqZNEZ1UVg
Eyn2Qb83Qa3IvHEMkGrhAoD5S33kbLaXaeqZLiVghxbxYOCUumNTa4iWC++SmfGyH9qdXhkoqzxU
vYC0czSimivzfDwHlPYbA3OoojfnetPEiME5kJwOlkLp7E0Pi2iDOQ5HQtO2ZaAHve5i/z8OOTar
mqEg4azm66EfV9uF16NGqBC50Jwuu7GyI5nLiTmapUfg5o2KXMGL/2HTrXl+ITUawUNl/2CqZ5ON
sp54lFgV7cA/W82Ofo6NjYYTM+F4f54Ak0VUjhr2jYFBFOJtwBWTyeAI5u3lU/yFrvLsxcIo9nKT
PfJq7hEOtZmL+V4ftH+lARiBZZR1wA6qWJR0aWvRh7QgJ9xhGCrYgGCaYNqpLBxYyWSCcLHiqz4F
J8U1gIlv+EldOvwjak82mjIMaEFR0FyXMCWK4XbViIBe0FnL6qRzK5LHVU3LZis5l9vzZoZZTS7z
YOophcT8XXNgKLS20+D6jH6hGrNT6XOu74XyXyr3EGKj4WEYLBK7M6QhnhZd0BGmCgEg7uiBUqGe
WMKUI08bwku/ocl5hovpIyykZ700nrYsM1iymW2J1RUWvTqGd86ayXbxHWulokkqIeOwtIvrf7Z1
9HF8N4UEt6mnEfIzuzQad8vc36MoQlO80bRPffw1E4sEiYjcTlaJKlCTnMtqVJ9JfsekQauRekF0
b5qj9FYovDd/kjPK0j/6fq4xtsvIJe5vr1mP0Ul7blWT5h2ZndQ7FlIa/UIIr0MlOlcvROrkCqF9
GP1ig1f4RlIHdrf7cYGXzplcClD4QjAIpnrG6Q/OCdmj9yYMD12JlNrfXZrNYJMW5+oW17iYDj6c
O5x2XXv/aO7a1mF6gk7FqDUo40w5CTQ+v2Kk9xB26HsiOEHYkLDj8QVG5CeiNLmmibqpzOXqVilA
Gowi+JN9n/8Yu/7WG079a6y+nu6thqYL+sfamIY03uD9FieBPK+SzbjVGHNErGqdxXezhg18h0Fa
QPDvRLvNvpdCaYFcek3rpP4idLXmkAiekf95JWqV2wCL7M6jnqhJt5zh8OWEyFYwcYq6rKDKU+c9
NJ1ZdKUMNWHhy7n2JtT4Dt0U/CnukxM0NUOOKGMCyNqCcfBd0G9TdU5ersPQlG5g6RHXRQpvYtI4
rvzHHL2WWLlq/bpYB7xW71UBmIXB+fMPrLXF0fkyeEyG0JyQb9NuS351PgtA4QbEqQbX1XGn71DN
foHj7TlZUxSJs7WKOLz/g6EK4BfPKv0sdxjSLeh7SkA/H0OEvog8x5omQQpgSC+fyKqkmBjzuLE2
pvZon82VzI1EM4Th8H7w8VOrwZ18Gxm4RWzNvyCMASmmwKYUx09ykanTQE8UlugiOShfNUU8vZgN
RkxJYbAKKAmGn1yf5ru92RZ8eIV55PLIXfSClUxy9jCKMosVmMddl9V/L2QEsp+EeuwEempnjcnp
/eXDtpDCJS176Yapca45OMcC1uSZra3p4LRz4rgAJu4PIBWGhAJHhujvyzRMrBMLqOT7nkgqjOpm
DZNY5boiyEYzhFkYCZkJBZB3zLKNn//FUkciSCAZVDiJh51Aiz8swPl6BZCzmOOxCRgDcZbPVXYA
mhvuHG6ErhGP+nmbdrQ9I6UxCpBy7AyV6xvHC5Cy0rwBnFtZd4FyYJtJ6O2cvt9+HRRvQ/yvDnjH
lXWNPb80tRAinyGPSlvgJAdPkGn70AwQ3jn9IqsgoxZ5Czzd6lk+TLly4j9HZ+oI8RQsl472/anD
cjrL8sW9wqqPmdA6a1MGoIVOI6/pkCWhwXqCD8h9lTT/A9xXHp1tXJIUJVPc6CQDh/nUGTtRLJep
VXWI3f7Y2J2CapLvZ10J5YTc6/LfydunoamjULysAnpGhXYSvsFZPBl1YRyCjFDFriT4vofiebhM
YWeSEa0Zh9YzGNfm/djgTmq9G8+IW1afucjlFLz6ygKwcathRluKmIzdR9+eB56UXoWipfuULFOO
rXkgfNFRIp5ozIzteHKb2c8yQnwA49hnzFBg1gzF9n5SJvGdmf8XO4ycsdhzusB/l8pZQjnXLjLi
fiwdl1PFmAz6EVpVgO/MSJd5K27ea/1sgHvt/Y/tArkD2Q8cOB5RoIp5IagPEfRvI281tsWCIyVX
nux171/lQ9kBX/PlP7RheYNOQuEu9up/W5Ly/7yweVKxB8zQhgYOXzBf9xvnk80i07ArnA1HLCMP
kUb6bn2GcDkVlrFUnntmDX6161yY9g02mZ3NsuwcFzYHtqcHlU38b56avdByvjxRBiKw7s0WxNsV
vmGtC1MG4DnqB1zFx6iet/wd9UlKI+XHfsw4CVBXAPzlEOHUvcWGth94Y8QtlJab3B20jYsqq8ke
/rCnyi5EjmEWhKv0exWXXDI1T5BWwAGX/zss/dW//lP1W9XhZshsojSTDY+zqNA1LzvlILRUyupH
wiLwwVMRsaEkUEiLpot9dZ17kDixNS0wpaTCWVieI6aoFOuCcIm63bMEpo68lqOD56o1VvaVEGKC
McnjGfvAmaPDJwfpJ20J3Na1jhavwP2v/m4UjTDe/ONaQ6Ha8N5QWu6ZvZoTln4wUuLnID2NinrN
SKiSVKVG1KQItaQoYFqsm56n+L/QRFz8v0yU9u3LxGhN5mxJj5Xlb4n+8H87yS+1s64AhXU9G0d1
kDiq5Fgp0cZ97YoyFZM2i64U7ar0OApIB4/a6b6YoZ737dGAec0XO2wdkTjE9eCCqXmiRDWwMOTp
qKDf1UA/lSiVuEUKhvdRQbafWFYn+RresZsnvU4ByJ40CvLhBkNnSeAgL6V/OC3VlY0JdN9725V+
6aoIIbt9IyB0+tu2WmCilw/8wFP+aexU2KYaNStUwQIzpbQaYyhui/4EZCfETL9I6k8isE5pbV1I
vGMidGU3bFk42jW1VpB+MK6MOtBjA/tX5EH5ZOfwferAeWsDaQN5zKNHv4hLqKa+GtUvBVNRFtST
ZwXnS28x/T/nxgg1cK/ZLccd+mNNQ1mUwpgPmGwnEIvs/6tQKKLWfJd0TJdLkRAqmP0DU4Mbw6MP
hMt9JiYCUktFBOj/Hq4b6/rhB+pljN2WJxbr0E2AywEBdQhI70HJ0S/qWrgUm7GcUOOO1oUblbjv
5Fv3TqUdp4KBEa38EB1hhe/Fz+W2j5z0OAQXgRHpO5aL2Qrd47e4u/SUnsezyTSrsnOKVs8PfnGx
XhrIk/hSlLzcf7MahCk8Ny55fADq2gm7zDdkdHdHHNAL6P8c4f6mwfXnS2A7QV6jIyH1Hx5odSuO
QqWR9k1niyVuialAv2b/IBUHiLx1u12hElvDilfMyxTSaU40n0hohETI/UhHJoald6JW9jZTAUd8
D/1DFLxZLnEHWUPM7sAXqCRKvLLojwC2Clrb0ueLBxVpwyWixE2moGVPPl55XWWB4EncNSAIm0pQ
qZQLYUKfxxLBeibqSZfLs6pNeUbz9b5miHYyNpkVxLej5zcw/h1TRWuuN53b/rEG/g3bFKjQz/NG
gOmVofulfw86p0g7K+HE/ngt4f+Qlgb+Ev6vom7I1+CTWBLKVxnFR+8cWhCu5W0cppZN4elaELx8
YK8T0j36oU+4tXjl1j+UXqO5vrbaBh1T3HZay2SzIlCqZ6M+SeQF3ut6MSh7IzGvUE4Wcq0ZV4Z4
YQsAY/Z3jAjeDoK6XA1N20yCCLjn/q0h5cgHSDGR/A+OO8CUWvfmqtFwn28dXu7G2UzQyR48XfTn
Bs3prfjvphCmG0BtfR3N7l3QIz74lHSpbA85pZ47mYneijfWcnw6xuYHP3zv429kVuLtbb4S8526
HGz5ow/CD9ZRTDSNJyh1iVBqAWGl932Rtzi2BCc0UX5gG3twtCNCpOSMO9uC61oNxZiheoA15FJi
E5DIA8XdTP9zyFavJjCDuXGjGB28M6ga3YIpaSHne9XGeJ6asWCWoElpaFWIaqTifPLptRwfK6JY
bXD+cFyRo6mxC6JAgRJBkNvx6TAeivstDbu08Ji6Wx8EPh2c6iAUn1A4xploEK85TqWGREG89SKF
PKcFFKaPbmY5XJgT/op5cAII49h8Nb+SzOPSOCptHxczEDyL2anrRqzOUKzkjdxP1ehWig12snXW
6CwXSAb79+gw9HC5ZuMmsszmzAiL7PrbDQTSbX+2EFQyFoe9zAF3S+RsHWs17oeJgeQaMIt86034
jvxQvB08ZmQdA1GW7PPYkU5e8uYLDHSDT5d+baycWZJC2GN/I3ubiZQFIBnzEDjIoGoBawHud3lP
oSCNoD9LWCZjCX8Ubz6CtdiLka/KdKX5gEKNdsmkkwYG+WPF3fyhIL/jUVbVQRpM7m1WV+Ji7ZUL
AagNmQmXIeFeiFNg3TtWYJDqVf9u3JXlsVHJMXeorXKMqW+IG+wc5JAi6lDPdyGsW8wdrOiOs+K0
9vWq2I5keg7TvvVJLx4qXQVgt/XOTvRBkL+fC3r0kWdSNLqmGaq5s4wmgMY0UhtAD19WJ7hg8bnH
wCIldugOIvnxPkqabV6nv+cWm3D3fjHOO/Xo7Dy6+99T0S0NaDwC1Oez6P6DrMwUr87txlMoM0YG
jf/paMkw83ncgHO7473ohvW+AkMOD331qj+Pn2rAJW0Yf0hWX4DTrEfW+nO4m9MCs+K2aeUOjrpG
J+LQMpfnFTmMSWqEEi87jxB4c9EFgfaAu2kdR7TEGVPiLH7ZjUgaQH3+iTC6vPOyaCx56q7aj7oh
g47o3oJRqJ+t/B/mccOeYmGr6VpYHH9FgyIYRdaCJAhNmRAYhBcvvZyyjR7e3jcfi7W8YBIvaZ8b
nh38VMbJzPb6qQ62KVaY9XcwpiWoVnZ5yYlB1mmOrYpkAw+soguewRyBaW9kEdlp7RO8TWxDkBol
I792zAiQjLZ8Y8qBA08+sUJwhrLuz+ae6pcBdpWN75M5iFynP7jlISUSgYpjVKgKFIiXK/rLVf2d
yzRw7JWu9y2v7FR3MtR/TLfGbTVBo5aP2bZM+HLLqXniYyErh/p8Wi4NIL+sqjNRb9YOkSiKSvuv
5EBqOorzHFGPczxBYK9P1Ga6JDUahB+2ovvslQq1hkbfUx0I9/SSuLscf9sBG7PfWDTFZDGaFP41
daPAbpswxkRpY5IMz8yWTU+GkTPkvBN293cyCbZ2aewwra4xu336k4L/27lAek8SCcyc6Q5A4lrK
Lwhy/yKXE4Fo3LlGCPRU7nPdbNKjNVMaIAmmVCet3+pQQoFKp8+VkGws4x7RXy0qxmvUtuBKd3gk
IyKY1Ml7jUp7CrIrREOCi2YHB7D0ebMFW+xQr5RMUCsgZ+IKV/xkt1cO2kpwAnqARsCRbRSAClov
kLiNGef9HXutTSNyKFFC40fhJSqZdE2tPqfKbHxuP1GGE/e9gnW5gmtr43yEglUkH/gSNZd/YLpr
5eV1s5R3U5b5J1ZXILW95Ys8OkFuCTCn5xofJmsbDU8F7JjekPOPY068WsxZPCcD3ytKhQ653z0o
xLUrg+7jeqTj8xbkyhqUS3njtjmpE8tPl2Pq5Jas2+xOSFfSn0FdnOtnG0+QVlAiWUX4DPQ9nKEo
LEIeMqZClCxAAX9M5J3CcsTYOOSp0KmNBv6K0E8mO8mHLOj9c2+xVGDaOuUFTu0LZyy0wzibxFX4
c8pcIC/VhWGNx8lbo+PbG9ye1tGMm+LrzBWuOtb0Y8ULYAwUAEsKJZZtEBi6tLoUmBva/sioUeXY
XsPG9D+7RT2Y68b/3FgqVI2emNoCBe4T6wsDDxFWo1c3dwKIdWQOI9WSYb3P+9+/lCGF2rKRhNZ+
c7HYWCak3W8qzXDWnzev4/Qe57Fmykx/t1d6cVrrxXiyJ3Z9HFbs6+VonWHs+LeRnAm5rIWW5wNG
+0j0Nb7HzBINbyNjS+utmgU4FPPpshHgy1OKqx+jGcoDyqNYlBasXDUENxeOmOmPtoZ33wYH6nrY
wrJL9EP1SFJyjwOVuqWatc73eANLtkkgFA7GryK++pOwHqp3c9r8QhwfAutRF6FK2ghbMWZxV/x2
4zkUm6dw73UqYvZRsBUqy4b7dQs/N6OpVTBQkvdnFVZrDR5u1Gth/SxpYZQbpuC5K/IaX0NXduQV
GxNMAnEr9FYhRueBOo6Bq2E4x7m5mlW+nrO5Mp3IsO+CjXhcf6wTSyjputs75q61ujkvSAUQmnOg
wFoSwLpmZQOCoXbLNLEfbYB/WAFUVdhMrBi6UqWN239sB0lNtd9Mqv5vX3fjuhPE3IX8ZGyCIeOU
OWHauIom+W03NToqTSw0L15m3rMhJjJ6kVfSL4nicISBQSSyRZe0sJCWbtYQ6sFSoke0ViCap3xW
kxz5CiyQ9YnHJpR/8hIYt0CjyqAh9IR11fS5UepJeEqmEjQNLOZfoo5g7NxdpN3wv5cIcFzQH/ff
bLy/rSbkbi0yI841WIp5iOMdmCuS18WITNTQHX/UiNl0Rlv3pRRDPA3hHszUW+uGeYgjfFc81fIV
xC1jAY5YYdvjYsTeN7e5zY2AYIUmex/d9CdljIMcpD7yWWDiSYklV4K4wQe7Dov9uDzsZ+D6bFhy
I+lX68MrtS90TKbZJDn30Ch0EtpHvvfMcDRgfo9GDQOsGe5u6bwM32nhP4FQnDpTEnyHdDcs0xjw
EajPHNvDmC7SVvK9col6p93RjCwqIizSd8r+/mKI5BUrtCjYpJ30DJLY0VYsXl5aF6pda4/zFmby
Mx57lAJ2SxkTTxCtEJYhxcc7uIQyjJoD/VVzqdrQUZpt/aek5nsa8XlVCQ+h1vLOw9b5leocqw2S
0Q+J1aZjg4PSWCskQjKHNCIiS5T/263Nxwztm8/0zZleyqFWRnz0upltjczLt4M0ah4i5Crpxppc
n8ucVHsvwPT84nnWcobRIo+gAm3TNjtGIQlsdAkgfzWB0u0W7SdTL4XJpd1GpZXZt1VRsna3qxF0
ZieZ6RgrznGizVyXLuirBPVbbyCgjznr68Q9GyfgDxB9g8WNbMRsjWQ41zPy7rwYZUmQlTlGbTU5
B/Cj4Rpcogzgc/cnQVi5ir0n7DZHb9uwhf0Uac5RNuyh3EW6uv7ti3DCjo65g8CHn8Z4/KkH7MTk
lyvfUc/8mazEY/XVrLkXvIEyiOxG5tISOgIa5AUh0ePYqJf8LD8FwgMG66VCHHEVTUhMFr4owzE+
FVYWTWVpU7chvD/h5rlIjbl7pZGgkwhU27YLmCks7PNHhYnrd+Qir1gSePIMAGwCtmyWQ+1ppK2D
1hOO3IbDIgitqWERv1eKycOd41tW4olmMXyjjl6FU1xZETnuusAw0AcvPynxV1RIfD5U1hp7BprS
mYpqjA7Vrmy0MaHF8wCwdSrB1oEp5Pe7l9W7zaZx675u80ZNqoQze+UvysBkyvRp2yjkzk+6pCbx
hSydyrl0AzqmH9WKCxZfjhyBRbn7q8baUbeOKK5MYbcGocZg71kQzCu+kAaXtXG2fOWMiXFs4Knp
KsGjPQCY9EPJzwvrFfkl2cA6M9Q5EumwRdSK89sUGnSLMFGuDJmokEORSRrVHK02Kw6zYnvqvmba
8cLUND/s3JC25nMUu5O6pua8u24cStMM1QOSN6hB73F1mRUAN/cUatf3pjJp1Rb9RFOPnzJwj7r0
XJ6ZeLDfwEQcJ7rSm373dcODnYzHydom4k4Q1eyqRc5SwMRdzmCeSE7GsjfhBZ9r1VeSzjcU+joY
lw2lO0IWThhwz00OxVKfUdsb0GDz+IZ85FCeflVYdb8tmpZ6GIz1YnlBvPYQFDpae6NaBTt9Ach3
GP8vmsO2Wi4F/m1FsmRBGINjS3JZvMwoGPtL0NbUV+e8xZjmDK56NxPf6+9b6NhN3QDhAipechZH
QRgOLRyHVv1CSoBZkx1br1kyvsTYgiYE9JcTwZill8GQ0CMh8SZybbDgAQLiSaLZRGVNpLZLHPeV
msXlIdYzdP7oChYACwAVLzfw/th5Sy8kGQsbANWP/lvxbMZHIlKlMntBDXFDpaX5jHfnkO2B1xUQ
f7by0vHXjU7A9JX/r2gqEf+8mU2eIJACW8Bgi8G6odhxlANUEf1lnilIyC2rgNZm9l4StXexTbkU
2aFwhsGI1DZMGSOyId9RXdYMa7Isc0PeqLpT5cS9XUUJeOLuYHQrhuNq86lcCVI09huXzS5tUWZV
KX5s5bcaaf5QXL1syWsBqCxRMslGky/DxNB7LKK766UyeQ2uGRgkWf2HwDqhf8HL2TMsT2HbcHgv
4Y/wGnhNLSLxC1Rqsdk22RMXxdfcZOlaGSKL48VXWayHq0WoOSk/jpx6jQlASjUWemC8EcMNsxG7
4si47ikYSLvQZEb2yFp5Vj4vjcNSrjkI/VLqyUVE00qCWfq6+Cw85+8/vptOtHyQxdkifH9jon2i
pNSbkdLypX1aw3gt+vlqaR7pCTgUsCEURTl+OY3zTjEUmeWRWJr76aEnLXHNxZYj1DRV2Mxj9dl3
I1/IMnxKx0NTsFhF4uM6pf8J8nKmShpqEyP8SD/psGincSqqMubE4FT1t8zGGPCoFk8yywhmKuly
AS8FEW3bahe3EXeNikZbD6t1nPyNREnIVBc62qn7zc2ijssdXMSSWwEhMKQ6rC3LsQOZuoELaRpU
mlpkvdESPz3AdLDT5qnapshBW5Jzsta1TreUOVB543yT5aoetT4NO1GddACB0q+msWS1OpM2waeU
iXgdvvPT2oeVP/zE7tLRNnqkczDbg4bv4mSD592yl6x4oWKNBjeTh7b/ZJQ+P2EEWtRvNHyezzXW
I7gqY/hffNeuKlI1Ic1B6+igcvMIeX3mHGGOPUXVxuY+mBm7r3pYIR3vwgREWM8/HByPTRLgrhf/
8oxgQKqrBpFyulM08XyBxn0PZaCSuv2j5gX03wM1isp5NGoApfpPke4zzmFdIURYxn1xUxVcbVEM
54mT38m/A23JvfI4Iy7EPnGxXdRdy8EN8HZ9YZrJBWKn0+PxJosY7xbHnvu3Tpv1Kc0pw6UGl1UG
lKIG/4abpC105Qcn8PagA/DkRcaPIhlyYsVW5/Hz6Xns6DnpkGLRwWzSkrSjxkhexir7o8aOAb5N
z3zut0j3hWoBTd0jU+L2r7IbYrz3apKbACQzKCrj9vomPav8o1z7hNV/LekAqIT8QYVBxxKOUF2N
W/q98PV6qNwg9yA/ih5UEbhkAymPuHc6mdLfYPb4/nZFa8ELiB7vwy/EUWq/Uy/zqp82/uF5XpPK
6VBXryRlSabwVVYilMNpvQH9yt4P11EsmEwMt8y8FOrP2Tkz8MCfRS3FEWuixk1EoI1oat9k8jUt
YcRTXEk5hTDHw3Pgbo9pLxAdOAbp08eac8Tqb954uFBr1YJaaaJvn8DDOW6AVIfGI28TLhGAybvA
OdzEGirRagc9GF0hQMGKfg/rndHAF7D/LjG773fsM3yLOXRO5wKWk4tecfFqIh3JKLEXg8EL5gmL
yOVUZfw16Z9i8zflSFGcGPszxJw7kr33XhoUKaG1fs+Fim6EEdegklXnDyaQQgVql4phJQXZCzEQ
mT1FjOUyV0wy2zTx42OXUOsKPPCziriEt9/1xfAZPwksTF8dEumRLew3JKyAqz4BsNWWPmwsf0Ba
hWKPprVk/WnxuWkB/8WyUVP/ovUASmGEnXK+uT6YRNasj6akFtrbVaeS1dZIm3XHj1kffsWGvKoH
DueZXYzwFvgpMg/IUVeIBkNxKN5XA7OCgiYHaz76jWKkEZ47FDuqcAyTrxs9gjmLzAkbEExuOG2u
W13bPy3WfJeSEDPbJ6RIaKd7GmEY9r6I4w11anyGArMJOREibjJMVdIDQL0GQ8gW7d/fKFbJIhJB
XPAdR4oME13VnAi8oIrngINztfiz8X/wZcI/kZLDZHW5OiXoKso1sj0Qh3AS6P1zcv//88czbVfc
Ln8uOxudx9ZTlGWycQ+K3wjBRGcf97ERPJ8wJ5mhRVXLYW1iB7nYS6O+RaKaxP5j918nRblZDoEc
NHSP/F/wLJg+XpRAeNy2paFlv1WC766QKMrJUJwErn45thxtLvxKRXKIQ7drOG6kVy/bDJT4zt0I
F2IYkbh6jzwhq+C7F96n4ru4uYhx5M6NYmdxEWpeNYPrvp7xXKGjzNF3deBkvxjT0Kd9VAOFsTCb
AD5VpV/TMtJSo1ktqPsy10JFZmmgv4Eies5fx59lTXhmRaNFueCIi63bAXm6Sr/T993Eu2FTpxF4
lh6Ktq9I2ZM93R899zWX6Aqfrfacvzyia8HPnQCE5ft0HhGd8K0dmjg3rmu+a26FXnLvoTOgtaOs
BTqnShBQRsFePnmNgYdpaYxnQ34yUEB0y3EikHImY+zveP0kohHrHOH/ygTpTpLPCCiOfipBn0te
ozT8BuHVZTHRUETPs0oF9WMXQ5CIzXAKEmKdsc1g5L6QPeZg8zZTo9+g79wNlgcNt7MObY9501ZW
eKfZF0LjpfQICvwqX3+EtMwpezuYyM70xuGRR4ssBoE4MGJRrD+d5enRA1NRSzo/SR0qCUAZkeXm
V4K8Fs2cWtGp0iuDPsPFaGbbxProETP2Qy8NyyT/fmvsbGqdDJUpoDl7aIf8vpS7PLMUFLcdp7SD
TXfp6uEQzfeM+u7L7rjZZ1D0D9l+js8dPcOOSOuIygFfEOhVSgugub/H2s/r45Bi1Qsp57qhXVBf
7TauWaU6iJ317u4HflxNyohIPNeBGuBWtGOX4Smz/+5W5oXGLveXeI6+1hAYkFuFrkiJFppS6ccm
noLDpt63LgN9ePz5jQ+HF7M6UQ77Xg95sb5fiBGbKu5HVokrgckmgtkO0sWzQkLD1mYMyHbbG1Q9
54ioQU38CZF247mc8znIyKILnw5bayEgb2yYzB542EiaHfCQ7Us0DQHIdEzpGFD7a78ltN6aN/xp
xFQ+bO+lBP7VcGOwuRXe/XUlBtkK7XCOtxwbvMj5mY4Ss1MZ7n8+YSODjutwBS4HvImopooE98m9
LDxMQS7p61JmJWVDeRX9D/uty+orFTViggYNxHw1FpC5Au6Zm0EkGOgz0DL01LvlgJmoeIYKKFwW
je9BoBWF8IfV9EsvCENi6bSv9qOWg5Z9ep83E4mdEZeK09KKM4ht1DSA5od6jEzVuj5sn4v+0qj3
WU/f3asDTyb9ml8OqHf6YbGvJU3Q3/NNgGFuTPNb7oxXQWh8w7hdDIJO+OY4NELXcKQ5AN6n0mne
nAO5BQ6ikgNxlZa+D7Xz9MHmm9aBWPwBI2K4f5bYuocLSXJeBGuafGoh+UYX7zv7f3M+aBM2IOGr
ArCN4VtZsz45MCoaLS4JMiE/MeVoYC0uFOex5768CC7Ilp7aXMAqszJz6XULIe/wFAujVHhyrUX3
0ZAhU1Jd6OXL2buECpqm5ywPeTh4U47nEuV85m5u6Snd3+FFyVyeH5fv1wLIi/GWfM9iagDtgtGA
X45gUdJfxvINOm6umvhI6l85R1TwoZ4W0BXqNUVEe/h9LtsuADjcu2T/j6hA/BtCCBrmDxPHoP/a
X0Rbw7zlT9Yi0798dNjlspVhV8rwCWhWQe5pwSC6IXgPSNd3MhSON4ZkprKdHrFf9x8ZFb+BZWNy
sgVwyEmbyJxGe5WLTtmMjSu39voocZioymRORTDeFPlPv/XxBjjtzbpv+YiMul7OJjMpSO7VvyAw
tb+6pEC2nugxk+gsOjDy8pvnAFyssKonOURHlqE6Ed+S2HYWEolfA64uOppdRTHH8hiZcCso3uZR
vGb7M9ggw21xj/Qc+0gdoagxQYP9fabVLPvIiuKtZUUT3iCo2eT4tyQMQcOMDYclVBdb4g944tiU
++xC28TCfw9tZtEYGufTSyYW9hRCTfb6ez40yHhEaT+QyR9dFa21dQ4AEhROVd0k3Ol8Jz7dOb/t
qGMJvvp1/qq66SIaIplc8/Mtc8+36IqYpEr4xlLjaJd9ygIcAlp5tW8wfz4xuQpyWBVg5akj99s/
jf++wGkQVV6rCMmZhUE5skIS5B3Vkyu3O/CVOOjVcBLHZuDv5enNGNKWjx1O6mZhK5dgjQBEyEZn
pC3g8Pj5njB3H/JzJNCjLJDc0A6DwaF/a8WjwJ3hEJ51N6g9FFkbClB5FPNzhvcQ0/211mIIzlRb
oRqSRaMMdGCRpY3jJcepOSS2sUBOPPnL7a3U8QJTUIicBaLBlCer9kcq8UpAK45PJIUHzHFV0BgO
cUQ6MFaBbzln0/+GTALWdcEFGkfBmSR7Sg3uojNS7+04SLqSglLD2h6uh20lLXHECpmjgerjSq8X
WEKhs0+/1a4DMEOLoS3GKYWSYUPowsYNTp91Y26isNOqUOd501UiJau6jY02gdPK4chf2rfSVnL+
5+/YohSq7pkPiNsMS2NKxC2yPbMrc/krTcCR7nN1NOepMOa2XD1ELwcZ8Sl8I9NxQEV42v8MueHw
v9S2UBIlaMW1fqkdOUfieGBztdkvX79Sco7bc1fWME1d+M+FBJZKUTmSwjKlQfJzC3yhCVAPAyNX
KcKy9u9MvPUrev+hUZcMzLVRdfPZttHgy3VjTZpKig8qMvTKR/sHt5x59fnbHDvxC6wprRf26Zoy
Z/d7tXI50zOBhgbAqx/1vvOz5VjJD5Npf3g3pziko+FHY3R0tcDqDYavK5+0M7V5rDEBefGbUHzm
oXzx2FzkDxO3uopxV5xYc/2sXAxE4bWtZubgh/lZvjmYPseSej1VtJoY34W/WNG4qM5yJJG2YMIZ
IoOk8/C6qe0hbbYQ19a6eE7O6e5P94jBeykIpx2E4tXtXp4+7myE/ubzEJFSMy0g85japnog7iQi
m3uMK7CBvDlmHMYmM0akKmaMG6DkRrsNKusnyShvsEj1XnwLInkXN24m55Mo5SWLEMasCL6G9Wjl
4DHlwxt+/QfKjhQ4Cj9tgwrjdjmgmpyXlIM57RtRJn8Fhid5jYA9qr4TBsUcixj5pz7ft4p+ev4A
iz6qfgtcTEwMj6kJUumJ+MGHf8oVzrwPWoHyCC/cA2Iep9msGYw2pEWKmrmPmDr37rCnKKYxAhme
hLn1xNIFRhYLL3t4R9lbbrY9AkSYqvdtCW225If95TyGi7ddd53R3PgX0CXTdMyFzxRhyycYyYJc
yrDqUxrqv6vg/nYQBSf8Lu6E9kVvzfd1w8HlkDSS+Z6pblYvEQEl/k13ZJzFQK2NbLyZU5ccL1hy
CnxY3/OdJvXt+KxyHQc37prxTdvXlWn1C+aYB8nvqEltja94I8S9hGEvqWY1YX4VhZHGsRBePXnA
+5tIRVipxzq2LTB4zw3RQYkq6QAOQrJetIlFZk7AkILq6kANeXuBR4GHaiKQlyf+IELvBFgEKdUL
aCtprCZmE90bGNm4FCI9ncK/ZiSETbdVrhKqTJxM9SwwcGexmMjFEVKhgI+z5cyz/imFDI6fe9yX
l/oEwuQZ/yxchcZI/ovEM1zUC7PVx5CLwhAXoty/mTQnRJgX3YEHdUlH2myFV6QSTxTQNUCcOokV
+qzYzDiYSlktmqMV0CNTMwR7BeONA0dqp4UY+XKfSM5O1JWuntXWo+AXayEhklO+gtof0vVRhp1T
Y0uzE1EQKKELCCPYb92a6SXgF+m1qj3q4hjIKGaxI6o0e3FPUFjymLNGpL9lCAd4jtuJNsyBFIBV
Yz2MffOmq+QO2RmglXmj2JFy7kM0J94MZ/IEw6ltMU2D/9c0evNINWJMBSds/C5/tVVHVxEHic8B
77kE0RW9LgHFcYnB9WnDVVvb7cT2hKyq3SMxekzPcyuBsbKJenlN95EBTctmqrMb+r1mZakMtSuA
53EEMZVetk5viZRtFdiKk6Pn81duiKF87aN+lgqhWUptziokKo8EbedWR4rhvOShVHmTJS/+c78w
APnSz88tpnhmGUjkz2G0mOQJgUkFqMUygqLIgfnYN9Kv2H7UaAJ3xb+W8HUpBV/xq1h3ApTqLoRs
fX+ClqA+m846Kmplt4JZXb1ciHMIT1Xw536jymkkcaEgc3lWlUOu/o8cOx9BZ27jiSRuc7t+LTPi
jjOvGZ8qRfDxq7OibPH4K/qP5KHAwZ5jyOr0xYd4qd9mEumRm52CMlNQqU1MtAI3SQMG7jaKgTxg
V0qXk1NbgrkIhr6h3gw2amSn7MHcCRvgPd8faApRcZnHE1j2wGmTgmtwSg+zDq728NrJMeu1RIi9
muJwTEn4M0ndeCXupXZtCbqUzDyj5YXTr7AhUw7HY+UKwQQBgbrGYKXbDyc5SSqKncy96ITHoX8x
2Qe9vbDZQAN3BH6bsLmbout5a1MtjH2OTm5ypJglr24OifdpurIbpKyBYRSBLGbzK5ru0S2/fOH1
0d6Z/p4HS4UAoADS+uUfLhqbi3hvd9z4+d2GQRlLKMJGO+SPdkHewX7GviGmcu8AhNVBi1mORNgM
BRstJ/IM3q9yOMOsDVSwXuwZkYpCHRH1qylHw3DOntLsQ4MkrrqhsdABnE0uccBB+ItzKMD5pjV7
7wH9vqc75+YtnCCt8ADJswetk1iOtZke4b15t4w5R5AhbFiNoSuDNDrJLYMc1NpVdOiSoRjOPJiY
IGlKv/htcapkQuL/rmMbgZ/54Had4E7aqdE/BkRe2+c8QYG0bubql2OElMNUZlpL+I4BatxRPF4z
6lFTMcmbNY9IZFnGm1cLf6UvPKaxO9MCObugNssvgCOuXjVlkI/5af0mWOjBhmm4UGhDNetN/ZmC
rCi62b7zwowTP7Chnd7fgBlHkWfY5FBgEll1vDcVQrTv9VnfOd5FHwnWUWYUduBAygaAvmSOpBsJ
db3wXWZWnWfiUedXHn8WTyJFzzQJd3r6qJiEAiZsfWK9uSV455dpjNDz1IsvY8VvfkW+248Erj5p
P8ghqFZPd/BD5UcxwUgML7To9nTWKMzZYVolWvLhFfhaXtGYPtPq+mAynrF2PP9WfYdg/V85VRZ/
c999lzwat82FS95nHbzH5DKkX9GokMGjwpyTobFN4z3eC5RWPvvmDTe3x+wE0IggpnE+UwNjYjuw
lIyvWFQQ1pAPKmXL2poxQDf62ciEvV+FUwTk4y0crIHQAlnNxEXWtH4doJFpGdIdHJ5Z2WYwOUyI
S4OUi0mK4dSM3kh1GobIX5IuZrsnuTCewn4jcv1kNLru/qnjx/hz+bpq57GEWD+WxjhI3OFUbboX
5kaDdH2xdZ5eHhIGSNk1aAlrCvqR6+b1MApaSSGvDQKmCrN/SpwQmqf8sp0IN943hZbKLLWOl/mm
6onYwiuKFfclYdGG6dwLR6+q9q4e2KP6azu3HZ7mRQvXhgL/OQtWp2PsJqD751rzGTCxYDlYc5Ak
NUQrUGk+nkirEXNrXngiQoZdZvGGLea+Lc3g5J3/asrEdP+C0i5Nnji0C8GCf5s35zorxiwmdyIg
vPa+kA8sNqjzoUzgrEeXFAXb9sv+0TT8AD522GY5dD1nFR1vJU/unqDGlTNt2P+NlcycUcpJOXme
TA8In744zNpkYKngSjKETqKJGb1Gl/ALnSE/pqHa3ms8euKC6aUv+bQLvzH2nK9tYSLnZ6GKhO1A
5X+xcNN+uMVn4GrpUhhouSw5z2x6qFjh6almCSqoy8r8RZDp1A1JRjrCL+9vYOjhOhaf+8dMhBVK
6wc+UN+XCe8Tqa463NpsJKj/wKeAOvsRf2HMz1gf3Ee88pwZqsENv95aokFJopwrOh55kitQCKP4
QkiAqr3/efz08CE6Kwmha/wna1WSKSKg+jPmyBgMfrg/wf1YaQK1QbBarZfgN/yj/V0pGSY4gPQ+
fCnp2Svh7LJcSaAhDAuA/FRW4Hn7ZBS+hACypiHfAk452nV1b5pXuplzHw+vAOgv1T36k7JnpmVH
CAwXHTumaPaQ+0etr+XWtRWhu8y977uvk4Z86MV+vde9Hx6Bt7dz/R0D+yBXZlqE9kEpnxCFH2b3
ZW+P9ufGZ6UNk7kwImgcJ4GC4xgC74kKKGKarXv/Ia35BfqVZQGRhpeMD+eYoeeJICtOx9NDqK8l
1NtvYNrAZHU8BanzkTbGVQVd8CsiCjQonhsdsAb4qsMF3fXZEBWB6BRSGjE/pAC7L7qMtVg+g1QQ
sF5Co+yBH8WOiivridNfvPvwtTS98oqVFaroitL1BSXSZLiO3uHQBnLbnQ3pBIVB9nstZsPZzAtn
93Ur+LxBLM56w9OQ0JfIRoq60mvdK9JtZfFvj5Y/p6DAfHHxwM/2ON8jyaNeJkXDEI3PJMpUpPTq
l0iN8WC0w2D1UtHcRA1VO1BfVINFCL276KTIMXHAEEX3xZh1qVzWGBTbu+COsE3XIV4VcXV57r8F
CvzzgP8L5XAQgMxk6XXiOR5RB2ZuskYdc2mY4A8xJeyj4f1UvvdGtahnu3f2BWPQj9PA5P4ja2za
GGeoH/oX+XmJVaOyYf+aKQZS3bRaHqZxE8prwKhd64ySrMzoIZtTQhAAyu4u29rm6RUqnLJnDngO
0BO/9o7/txyVR9lDN/cl6WnrXrbBsK/+PHNVheaTsdsLnIgKP0flLjwV0emHB5/YurOOl7ERLepO
b6bPq5whkNUklNjLgXXO1WB7kxlKzdt5wtU90mu+beX3OOxlnKGVnmUReRso3frJPAAxcGPi7Ifd
75B1gYUBVPavv/spPN6fly1//RCbgTMqIfDY0mg2cVf+0xq9DBIHOCJPnW/ZGplcKEd1CclOxkPW
ztcX+mBF2l7bB3+itA6orFJzzL+ajRIxrGsrw0V9qepRNCMNkPsHee8ugnfVu/1NlD9BPBDgVur4
yJKNtGCgNzdEMdBJ8Ld0aQHs7a7QRinl5MNtg9xvBWKZ77cb0Rv0r6jlNbs8hlYiOgyGURbH7152
gHvPRiUrj/IVQvZewcxEKCnv/Wm4sqp/4x5Heg1bszKIqMgzPka0U3NT6TvnfDMVik+4C94T/k5W
yWA4XK0AeOI/+kizuXzRbuiOZeCw6fsBE5nQWKfjC3cYYFEouKE15LSronEqG+/sPZfoXZjPE68h
BK4wUWvZBMmOZdo0no624oTinncSOM2ETmSerD5ZS+EuXP2dWpmtPOWOIhwqCrfzyaN229LRaKEZ
jHCwW9txz3DRtpTgZH/Aeg2s+zrUx/0TiEieDoYkplKvubAzgnWVF2TAIcUglT0ouVYPQV+DTlBT
MBOKlx641zebm9MzYss3pj4r/Ac5RTQ62sH3+n+oHAKe5kyJtYmd/pzpEZemajsvTCiPJ14y2/NV
XnBHZvSgF+BfVpLTK16mzvZ1G0aaL+q1GSgNXRy6B8dlcQVPhKD2vpq5RFdO1ufAmuwFDYOmLdcB
u/FkqJhL1SIaAWNN5xf4QpzprQPQPo8mkgkRZiPiyWI7a1J1dWxF51ED5EUMci8yUREOilhrxGy9
EIi7PWPoD+EQqFL6iqa0dE3wUEdfyWYKPNoriaWydgX9pdP0z6Bqi0SUY+HLRPKGeoANqybJnC1M
1YTYBaOPgxuyH7F/lc5DHoq9ip4EsXqkoYqnJPXu/e6mFEwkpRrgMlCFZ2mGMwg3ud1G7xrh5eP3
0+SE+gljBtTE+1BBf5hJjBPWsYA0lgGtoOf8knVTDUNRf4/UIRixm62CU3/w7+OEN+CdpCxzyAB5
krEjUVmH2nqLWOyMkJJCle91ZBD/Js1AiX8cGmZRzm3hk2M/lYvPFe5xTO/sXVUiH818yOBaE+Is
LGVpdZoXKYQeVGne0tMhhYGO2edTyaFuef1fOwVCW8AgnxqocDSiVXjQOodNG1dyie+RqohaReNb
JCnblDOOvWKKLTgFR7OP2Bxsts65RKxMxluA6n25nMxFg/krYlOHgXK0QdnLg+sJelrK7gmZGw6Z
/VSfvrl+OYEylzRhYCITPnv1vNrN7oolWa2mK6Z1a9giawWwPWnSoDo/p9YWSj7kOf7U0vy3a8PD
5tfCkyohSXnnm7HvPpDCLhom/2enOAHnJXBBUCXbHXPwouVIHR5ajJGyD4L6pD237Ob3MCgUW/as
OsuC+oZM73uyGorVdqlEPvGGLCeJtj3O3hiMZ4CpS/PMmFPVf3x1u5bMMo7oUq6T0lWvMtMkWjoW
YiLopOvFAiA4KFPWe84RtLd/jUwQ2p9WWhMxvYrcweshcSmiIJvXqNbys2n98nT3rJOXeyZWWfRK
5p3iVCmNz1ZpyUBPydcSQzR/eAViuhF3v8E2OpexA46AphREyuA2Gwet4/HK3gmbHFpifDmnqGAt
YOji31T+t0qsCjBWze6HiXuzXGZ8qa4VsRJjuoZ2oHyrajFcPfX7xiaGtnJuPtRlEUIl7rFVvhvW
MuSqQbEzwsBvi6ZJl8JW8PzOadRjErdYUwf6jFXfuUPefypkiEf3sgCGMJPkILRRNI7gmX6gU8SS
TJ4ntorRiM/r+y7k1Dwb4hNiIFdU8KkAqij4XqgYIIe4axj6HvZXc9CQSwY2ZFY1zN3jN1AGTJRW
EQ7Ijd31FonuwDZGxKe/03toMz7sMkWuKNsjDoHOabw8YJIFUuqhYUUBjcxRz3UM9WEFe4z9QX3f
RO2ntNO723PbAW8FBTat9/KTSvJ4Qi9kCeb7QBsySQ11DQsYFNNINN4C2bWHoNC87zWtbivNz1n8
Ln0DK2qRxuPlf7Dvkvsi2/PsNo2W3JntKajE0H1R3ny+JVtcDnBDTubgE6Gm22WZZZeZtqbH4tPc
nFRvc/KEFQR5fX4NlJwW/WyVglyiAQmx4O4lRe3k/B4gpybsZZLfJdxkI6zVllEyjL/zYPOk8Tr1
Wu49l2aPxv+Y1ntfpWEE2n4P1d/cAhPIeel2+GcpDfQZBYhj8dd4VCITGJ/7bvZxGzh9mg4Rj255
V28yfAYwDlZCw5p/EHM2l+ZpmP11tKZILJH1PBGTlZMPmZ4kjC0jBMrsJ5GjGZRYy4SItAOk9Shb
ZePUvRChb8+oxqNFqgBips/Yo/TGDJ4FZ7XX2IuBe9vg4/upL6STBfHQbey/OIcWCcjaM71H4zX+
YD20nIOGStaGSiAdwYFYdi+PrKSFLCrWvBqd5lEORDLeorEJJry97567Q638spnTmwQ3Dt+JwX2H
E/nVV9+UvucvSslAWCK5FZvcEVntqP/GWRYqUGzPSAdp7IpX+ieRxKl+3TuuxkqNXE5xk6sxOO9h
V0Gl1dmj3/xgOvSoYVEDIhGFDdXRjU9vYLBcSHBZwOq1AxgcEpUO6zoWFga4epXUBWBXftiiTJ9e
YuLpAOeW0Bpo+7IL4u1EsIWZggtaZkPEq0NZPTgzQk6RfEobL9kewsLh1xGUuI1b+r4SpW+l2ppq
pfZ44adoR9iP4kio3nrB5RU8TnK/fVZS6SPB4OltowUbGi4xlvWkmhrMFjHCDyNVjSivYj+lXqcc
aTxCGp90KIYRQzRbvA3rJmriVl6PrKKe+YTnyTtM///vUAt1j8T+TCCXH4AzTzjzqMvstmjN0H8a
P9w50qgHYFs/3+KwHLyI+tmvbl9P6RJNAS+B2lEOoi4q40mX6cMfphjK83MiBBB3EiOSUXmC2ww3
jrrphqJX7DMQ49gcKuzgFhrCkY3HAmcK5HxbQOKtwUmviP/E5DssENWZ9TyOTQWq4iZo/HPsgcZZ
dMkcYhppa7r3EPYhfcDqwfjcNGNX9iquTNVFykOnUEGlbpM0RlhBtGEw1Rzk3I0cvaYuGW44+sxQ
Ey1Ytt0JocLQ+qhod7x4g2pnBX3YKtPpS5fHpMSL/0ZGnqNNC5EUFDWuxRHoakBjvumVKUQqPToM
qvGu5ETDs2YQdRSy/8FxGzq2lmcevwKFF9u6Od4cHQPsvz4wfOfbwJ1mPcvKD+XUVVa4sozhbP+q
RFqTcMtRj57hPgZg24ifR5eBqvAbnf0Ai6sXjif0uiMzLTLb9Mf4X7hj1r7EbXiKD57EjA4cNvxO
uxLOanbW2euUkaQviha8Ql/XWx3k9a4jCJuyjoOPKCDwIN2+FifosZ67uhpoTRPX/TAz8hBeavGX
xiu4kVrOC2Q5kXngkl8ijw2VdToUAd4hatli8REYElQ1Yv+J6ivypwlMvWPDvUXe/rFEZa0fKLTY
SGeWSxRH8ERGZ2U1zPNxDYZaXmYPSiDQmTTUb3aQvZv3wpOuYlHxgPBscCUBSpznfKpHzQJ0U2qT
3tAH+2xzVxTTM9NLUGVNVNz0ZwyLLprPWohHcKtmv/TRgeb1YLCbhfDrk+AwRWoeAs1ZcsPjJ7E1
2yoGgVvTTkrMTejXPSSp7nxEYsSbXBE7IcjjzkbJn5cPz0sCsqOKziEBtp3cMwgCkZBdc3RC+y9J
4/Y+HrYn5OB3IlySqxZP5WxL3XmnJqGJ03WEDW9vu/9HnDrfPV+bqiXwmvHnveyHkx1snqqDQvyE
99pdKhsSPP9eAwYLTnog+qR4uaesPSr5fedVb5l4lBqO5GRqSmrUnh+zzR+VB5lclvjUWg7wj0JZ
32xXHAhrGSLdPunUxpyowRuTb23+GL3MJPUgsuu99HhWfluWW9/8uCK01bq3b5HTdYpIcLEcbx5Q
xxVBHLnCi50BLefBMhtR4t7khlfRNiGbsrtR9+Nq0vu6oGoOkzOThuAVhoyigT0BWkdl0Kb/9wc0
Q5UsrVHpNBR80hwfZKIO5N6hsb8LNaiD2PtJZWWSzMk6iISuVEvgeDIcDt7D4iIvj8t6uolo8Tk0
93jYEZkyxiXjdrgq79w5ilZBdhGsOBJip71JgYlfMSh9y/Bay3MTIdiijxc/d1m4MLwmQOWBLyfT
UJW4EH4DVIMdxR+V5Z3xUxi7PX1Fb6Ws2HJgiowuFF5BVThLfh1AfMbjUraUGyi1Yg2umLTr28xD
EeglZnrynfxpE8uOQ+fphSFzctQR+mhuS8yNKjBohUyijq6/nNZlGhILvXiMT8WDPOkal/oh4ykj
ZW0NVhYo/CIncRXvOPZH9EN6jQDUG3weumO9oXU1lU6ohus9L09V2jv+izwjN57RmTxm1FeDCYFX
9LAKA561OFHa1xskxLfOuDjBIXWDxyDuj8/AUWf1lTH93DkDgoSK6s2TnDjC1QDVS4CdmDzAHuVj
qY935fp+hjLuMEx5vNG8NB8hBQwnkmaKSqMCFVGGb9xAd3ll8T7twH9AhTaXJ2yzvJltniC5a792
3+7y0y64W/A8n1eMki1IAq+spO4eOOhMYABGpjHmKOvj8hUxCJ8ya0UIWisW+VjZREwvbaonU5kT
FN5ti6qCsmkG2oHH86CfTtgAA2LJCCqFD1z/skdNr5iculubxyNLiUYuONKT0tAs/ZUXM26w4vBL
w5IymfiOLnCWNql3xn3qIlzbP6GYvkN3VyJwBsEbBqmj+Rd8FJlNOPX3BFGcl0kkQhaVqjRtAkGW
nr/iYTCVKHhUXZbsL8ez3TvH6QKy/a2BlcQxEN4iLNlQhmQrv/iyZSZxVjlsikvrN8JhbYhggGNH
B4UbIqc8YOxASLCMkhCHFgMCXp+Sxgu1r6QR16o0697xG7rIaq86cjQHisaF/acIVU0bxpDnUpTu
3UfYLG0hD5EJxr7uEnuJPzwO+/4tZVhOft9379PmQW1TuL36RtfzE5k1/nsIZjOsorjYRExIG+tV
mlFQ4sAfpPfYxigco1PrI3OqM/XIRFyRagqtJmcNDkqRh2GpXywwDEBrZIyQzFcvuLlvLiv4ir0Z
xSqkWWglx9D5k4ZbtUnFbd8rcTEKJ9W1QO83uWkGpNW5g4Irft9gJIRpXgkMnK+IGaPE9Ct+bU3y
vMGsC4bqwdzVCB0GQb6pT5Y4MZCRQ5hUD9OZg/eaAmTad5OBDYxOTMa+9hWhgLuZm7sceificyBj
5wQZYd7B3Me+4hXvGwrzOoJuqJkGXrr1x693zxCcFocc7/YJtcgnX1vwJzblX9DOi+P3xWC+wSzT
snd5TUhptA+OBljYR9swW9W3GJXWW4KzlcikpZu4e6PJqezwZJ7mPg/fhmx+FADyYgl2atVabRZ+
ZTIVas9m13f8HzSwGoE3/l9knQHSpkd7hQBqnzl/M/XSlQsaCEcBOZ41eES+cDZMduo20B7SNY73
alV7WbwBAS0ggxAyfgfBxkxyM0YwwvKs+1S5IbaX1eOB0noZkqHDn9R/ug8R7D4WUSuChDsa2fMY
xxPGSXvhlDg47/gka6nSKac6YfF81y7FkO9qNfsjgSQ/MOP1WHW8B7wXQpIUzxuRB/q0Sxt7K4EO
3t1AglGOA2qtMA7a7GT2hVsABnFkmoEHXTr4prLC421U9NPXAQN4R9rhB85iPnPYltDCtHKuRcrk
gufTk7lYLjADhuzLgTlxlSINFAZ8xKZ3xVt9rd8FZlQh1H/fppcvpgeKp8w4cpAl7pwuiQu4CuMw
UY8H3MxQL9K2N7w3fOlh5mbG9vL7nKwu+Ag3P4ndmtT3yF7wkzUskzBlYwydBxTwMWnJc1b9ib2O
54twceY5mbMJo0Y3HCmcCmVGjaj4Tq52eqwPkZ6A0IrLMWRzKFYVx26ImQYHHZOnSnQg7l9HS3Nj
ZQTpJ7XzVqvrSA4SAC/Bpe51TE8LiVixnJ4YdaRI4+P7J15LYiKZD9Lowqkm/OaYPBw0h9XpZbAZ
8uz6emg+cpl0Tmt1ZWXdT0H5H/L62JF/49UUZGQ3Uec5IkKhoywbp10laa0kVNr5PG7yb1sF9vFz
i1UDnb3pVvnPyOuEvCb2ovPjd5mcWpjcCuoWHiMEdkF6F6u1iMjUjLBsZN+/PDLYqkS0zQi3Wou+
ERwQXlggo+cpIJrIH4//E51K09tSc+fH+J5oeLasPe5Sj8v5P37wTOvHN7ma4hoOB9XdTnBOY72W
ofsu2gAJLw8vb2XTPUZwZ7c5W6s+nlINXLjoBx7oE6jP0Rstw5t8AgiVjJx1p7EG+tp9L0XMljqI
TrGoLLp5M2QfjCQhBYX2WRMxPJMov0bUulkJM6CDzK510I6CwkTjbEhLiXRJBTCnGm9V89P+/7Gg
cNVZVHrMd+i9SH1qN5dYjzfhdewXh2z9YGgrXSlflq0Q94xOdjdIibskvhCN5/8jg866ckA6KYg7
W1zz+2kKeOiLemSo6dgjaJkFYQ06e5uCkJI1Hw1p+ImzI6y0OkQwDVJwOIEsBte6eP5npl4w5YZz
07wCY0G6BUrZNavDd2JvgSzn3xizrNKe2q/MWkSXy57YQhRM/wKFSIg2lKzUdSG2TY9fXoLgpvMx
wcQ3VSSEHH4DMmwSrqLJ6SgF3VH+pdbZQq6VO1aANP9aFnvhFkRNDh4vWGD9FpX0rE6SMhQE1xM8
lnCckjHmSqB7Uecpfh0ylK1R1uCDDjDOav1RPYJrlw3T/jtgBRlG2upXovFAYJmTE3eMdO4FnppZ
7zWRadWjB/mGJ6n/TeTtStolaL01Bodx9CAzU8B3Xz0f3Ejn4ZLpsgQZUBS38jhILJfSapYf14yc
JyBA3nZououz+iNagfDDLwof4dg/3fu0quJn9ixKWOjb8zjHJOahx7zpmw6FXR9dGpmcEyf5tGy8
AIUJRhAIwmk3vU1LYKkZxlSQMZcPKRyfkX2I9w4JSzVynB6s2bR14vfS3hN/1Bp0q8tKP/2VgGYZ
a/xP3Wih1WaT3yqXQpfXb3Bl1gWSGMfXyBkKke/bja9ixNLFt8NpTfnLSBSurh0CPNAvzy05nM+E
MpLBpXiD2uAlXDAFY2PD7LquD98YKOK6Y68RyscTp9qAtPDajYVCIgNpc/PTvpdPDoxPTq3atiye
Vcq4p+2ok++1UxbzRwq9hH7UbdEWapeTxkOebc6tvmt3Yyq4dgqfDpe5pbIVrSbXS15VFmYwIHpO
8Rd4YCZpHfxBmV1H4RygLcGxhy41J7HbJgb/3X0gCmjGLq6e3VhRUjH/6+W2h0GKnATIkeHMlkrN
BXfSQSrNWby287PQ87Dd23MhgYCqL4mPWl4EWBiO+vsy3qJcDu8uLXJ/nimJl4FKDgh/Ehtmtxd4
IhOpm0qkqdOmErg2b6HRoNSKv0UnU+Y/06Su3u8aYBR2yvBEdHftNh4OZJZINc7IoRSrbdKKQl6U
9ZI+myCDQji1Qkc699xxIVtrXO9KP5+ZfBfcBq5mx6YK07tqEnpND+QF43JBYrJI7C7f+uQibHWX
szAuWauIac6Mb09czeVrRf/1d8zcErx5w93B2XtV7Qsn0Rwn2o4CcCHFm96kCIJr6Yp2LnCT7NTm
Tdi7IC93N8HIDLu0qkiV8/kUosr20EonLcAyLdeTy+zgFfGSDvSufBe1zaGRnd5o7KA6dJc78abp
l9S4UfI2OnNm/ziyreHErvh3qUKibRQr2OY1od6zZsvWphQQQafRi4RQk/nlm4roxg3VGGE4y11K
Tm5cRbxugRBrpn0KOPVSn/LhBDKejUVRrM00Dtwv8ZwAlQHmlVv8TyLe5apvmbnGd2IHLfvORgvv
xyNPr7NM0ShyGV2+SN1Np4SadxarUzZyBlGJHxSOiJzX5tg/kMNbtgjobjix7QszZU8dtUtBhExp
IyhWr2i7ljITHMmSpBmRTwHuWzKBH6RYQ0qoaWIb6wjWey7oSRggngn6cCXEqNtrnXqY3pN5Bq/x
WJF9yTmVJPL+8y/T30IfCpsp2EX5KCvpVd58b3xPbgOzBz3kFV/K941RzAc6Ud4NzoavWHopCYrq
JtYfkbrsojmQtA3/RkLrYyGYelSmG/nGIHAYAtQb1C6W3YbTX85ivgBGDKNZZvfqEDWZK5G5+iiN
tQQnXU+Wap/u8XYj9psDFV6bn9I6uTwrrHprDg/BAZKzxEfkOckSiB7Zf8qVtlMOROjCsBhKXMIF
MQPSyJ988BV86qU7AFZEh3Eu4YTIhqH6j+uCO+hRbjZdDZZcwL2XmvIAvUJ+2eXpjborSfb//1XZ
KqpjVv5TuYyTUSFZBHMYGka3DL4ZLUHeDyNnpFOKC0z3WRisQw3L8/H4ajXxby/L0aoOv62H9oTC
xXhbIbtDNNc4HqL+PB1kPP/Stdl5MyBsW3TIUgnkg644059Ww3R5ydM/pvKxgeLaXVg0wiOeeUGr
se3PEJ3pzlhwWW83XcYUY5jzm25mlxj3abjI9miTtxrXptLoC3fKQ5a+sOiwm/nPSoXYw3jg75XW
2JEaeGGbF2iLb3eEq0jOJ+XfTZYRTkgGO0axYuEK1s+DHw7MbFCdqs2BIHpQBXCilPmyy2axX9bI
cZiTEn2gS11pGhBWk07zbJhgzlsQVGW78FEnnJCDtdaVkCxY9QlviwhAfJ48jQ4gbcVo10vkH8qf
zR26hOXqJCsIVCHGY9k1o7nb7YhrhVe+cKxYTpTctKnzhCpg4QimPFxvQuaFE5Xd5I/S/6A1EjyG
+QQ2KV+p9+YLUjNIdo9bfibnfo/hEKCkUtXUHPNAwjBdzOEcicZl1HoVKyF3XAguCPyzmz9VbROM
k+BPlsgW+EdULfPFZvISASQgI3vnJe4goBKUMWjV3kP6OkXbVnDgaOlt5p/pKMXsixhNyBiEv7pi
OkEYzqaLd92XiMfuPE/lr+uE07Rqly8XBopz8/x9gLeNmdJvTLFu0iuHxTs9NtYkwFFK0//e9oiG
uHJ1dEi/Z+4PT5EoZkj2+BzTHuxpt5vPtf/16e4pEGxyKgtz/QocUWbaNgGXck4Q7P5NxbpDhma9
Z0VfSLH322E5EIvzhdtLgTsg0ZcQXHWloiXmDkL8HS3q2EyqrIIRrk50dd9lodOz0MwJBZJGfAJM
CamLS5ATFPo90KE0G/CYojexBWMi6zAPmJ/yGRXEKTJvM2rEZed1LNTzvmKc3430IrACWbNZXgXs
0Odec7LQl1YbdUfE1utYjR98qg0ERgxFdQ/UMsqyc5E0IvgaR8RsxD4DX9v5ILIxjOsERVWWj9Yu
Nv3PV9bCBytRYl3aMKWUQE2u1YhO4j5OQ6bYSVHTIpm83etGOlmHaX6Q612Kq0r4877K/rlvI7RD
MpwTofCOTM3RmymPYpviaI8FSFDK4uvvLnS5Mm/eW0nXZtTa1KtfdPFt/M0wKO5Vbrmri0buMXcq
gdEBl8mIOajZ+a7fhiICzc3pTMbmvAWwIPE5jmnjJSnPv3+ZyBSUG3026VX33yCEZJOV7apH+vJs
6jxStckJ2mP133VIQlEEPuPEXor3ye943rUZocPQRN1NRnMqJrkVAuR49RqNjUUHWgP5rHAUa/Xy
wEWAOhVB4pjnlz4UH2NY6XV/hkwUSnFCg91285ERxdMYzlKJmVxWk1L/JCeVA1SXwYjWx5N/cURU
mEgPxGjd3YhWHejiFz39YOqJZwuYI2uP95lUQUdeh06rxYNj4CILnRlcFU2D+iP2XW+X7zv/1hlb
Dp53cmNH91kC12Ocd9Y61+Y1K6ImQ9utEx/HD8e+4h4H9naGtm2Ep+lA7Ke4VurDAw/G+dL0Brmz
nbSCM3hFHC9oBD2YABWs/yHWDSINgTlsf9gYooxKOesle15jwyhHFhdDy7uSvM6K8QCD9cf5mOpU
23Kt1jBm9uIudNf6YBstFCk17zeB2uOSxjAkzKxd/E5xzvUoWexLW/ecVQT2lDkSNg45Ygb3OP+4
bM175m18o0oiA/7pBVx2JbTNDx7zvIt6pV/mrkbfj68qrmbz6i7EmMsaco0XeQsnOdghnf8hKLaZ
2jzk7gF9uqbtnXixHMH9PfdRe4yRq2VTpkj/Hkw1lYDknhposfIrq6lURMiCyNpLhMfHDBnyqzZ6
RcC5nA0wnzma6p5CXfjjlYeyKnThd57VIMi3Mvx1faxvmkOmqWwbJrewxqUvndYUcr2UJy8otmo5
v8Sw7ay6SH0H0hh8hOHbo7mmmfYq4qxWX6JCOoCad+5jy3T2QzCElTxSoUHXEYrXijEF9t9gYoGC
/HttYouTcmNtPym9jMYaoKCY7O1kHeJoG2nNB4yyOu9SZ+ZbvK7SaFVbpq2azW06g1gkNSm7S+w7
Xz9Gk6zruqGoXHZl+2HBn0kJLTx7cjDbFiFz3jjSnIKusDpt+J4jxxBIJm+fyGMWNPWA8a2LgVJg
4lErxf/QR8dbjSe0GFtbgBQGCjGXGDha1jxkmalgqs+55S+xxiqLr5IYTtMsy3HEo5wDYefWEbn+
JPh4whBwHy3iBDL8cN6NSJY9PJFuddDyGluDmePI6Wia6M1oLAmpGtRbL8SeWggqYp0/PvPDIlTl
RGx3teIjWB8HFM3jKDC5VqezLNWY+Ckx+lT2hmcDWF9TzwbtvhXufd5x7KTUK7G5Ovvnoj272tP2
l6hCrmaDiSYrozjqJDtQ+ls9iadEzhSs7k9x0Wp3hCr0o87L+TYGwwzkKn6W1DG/A/ZcS0BZwTCK
llahDmToCx4qS4kw7aWc4BRHavzH6tnG45CV2yFhaAUpNZK69xfqkbNmWMre2qemIIl1vYZotj0k
Vqfd9s1H86pknm0ySf6tUrwj2rqlbU6lCjarVkZexj3xEMNdMcMC+QWMh6+3GpMqI3pQEpQLsP4n
mv2XlmxMQ9funC/SXth3ON4mUTAWQ+ywYl61HGJy+fEZCWIvNeRpkBxl9FUGYQaGhp8oS77j0wpD
mMnWWnCl/pBXbxuR/ke056CcWco4bp1xAKluaUVbne2nSOoJzgSF7xLK3nxW8oXJQ/yVp5mg0oXD
eE81H7OE9h0o7LGfyyeh9ubseUXm2TwKjMt7fVVrgmhRYIer/d4Lwa2CzdphWiUqOojfwq5YlGNP
qNn1lUWjlT6VIf4lybmUMkfFNh31A78jxpw3YQrUffVSYMjbhbAopXl4K3TEJWKt8fGCJNFmX7YP
mvRDSsEwiKmUU2FUnW0B0nmxBlP13H7YLBJpaq46yc+MJrYL/fJGeeSGaFY8KHMZCyzUno1Ld5tG
c9GXhfwlRAfiaPg8LMAh4EnCNOVMmW4VTt+v2mBkp0XkVeY87l4JeY1bTN+7e71NvAjNJFMI4boH
mjSh3DoNhlNNCk/IzBkj4FXaip1ZfstO3JAwo9bfK+QWVaz9yj13V8nD5zlmWnBrk1orC2COUkid
dN4BcAodUMbCT+K8au6f6fSvoojuHfDa275yLcKs2CevCyBT2IFEYjfRAwLamAd0qBtPgFIw572R
aRWEhDjq8xtUKpdCChbxa9iV6b7SPLOnbtHxHOP/4A2n6zwUNuuqNLUVbzu1YoBkUQLV3mDCcHb7
xKYNWulnpgtvMnMqWnX03uAA8IeZ65E7gIZtMFjD7OhAFMMiCMKpOYVjzS4OTyT6Jx2Kadmyhdhz
o8ZsNmuXnzaopi65ZEXBq/jVr4ooXZPTN7JQrkO/sJto16Xc7ojpZCh0wz4288RULwwGgVf+kvsv
F3utBLkm/kCQORhVpoVITq23jb0oxJhD24owyRRMSU1Vj0MPH2PwsXUPvgN+Yg2rhlyFlKtBbmzm
vDEYsEYe9wtG/AHtLhZUAuhWtgcaSKFNrGwW0dUeee5BpmdhTkEkpDOUP/RfLXG9/zE5l6kRiWQV
QvSEI+LM9XRv5xZ0gjuHB5yWWShkZJUGYCIY5Jqvk90MqSETwTTTHZsmChCpqABWx84sBevLLuP8
Vk4Gys3LH6vo3N9ZxzCpd+t5rtvETDE9NDLY7sVPiALQJUxkwgLfCBkbtgYhXsGFZh6vpYTiaboT
5Q6exalgJS4w4Nax030pe5ul/9eUgwcuWZpGSJrADnaMG1agPrYdpTHntaJeNUxapCiSMkvyCShL
Y0A/cpA82VzR9/M9bbvCDGQiOIOh1ErJjTNCGkaDqYLV4nSqRMEBn4jlxgS/LYlWTSYYRomoYhfm
NkLOA6HD3ify01iqvrXqitffYqr2uQB4Sp9WQWbFRV2U+h+ZdY/+GLiyF6fRb5sB45ApukF6xub6
s+hZk7W2+kBRbiSHy76D90t4U1/Nr8WzI4hNpKwdbpqKKDs/v7A7R6pMeTEPR6bo/DqEIBuZEx7e
TZKIL5WQbKd18rjCU29YfhltOiLMVpaRyj7Yhz99crF45fKt9sZj8DHZCPOZFNr3c3dmBVanhqhY
nDx3czP7vaymvZYUBGA0qMebSzZEi5vSaN0bvqxRHuZO7Ia+gtDsS7SsCNR6EUG9fSV4m42XI5uD
8lntCEsFy3Zw+nbX2CKP31ZKmCsFigsEcG9kRXmb3bt/hEM8vfslteYkB2QXKqHd9fO3AdMO4u4w
VwR7COCkpN30BI1vEsJXPzh1oMJQqlCeMeNB1Y2ngoYMv0rLOoS7qZfT7EnBJUKNJkFppvk3pzYl
+Np3c/zch65iGOYJpVLL5ahL0ouSIWTlQjfwc9W0evMcAR4caV95KEP85gngqDJHDaRhkN9M/c5A
XsFmpNAnz/CKkZ9/3C+fOwGcN22BmLo/EGHM5weOyTsSQNMxgQvk6u5Y1qF7cx51ZR9o7iPbvxoF
w8himXbgpGISjS0E6767qyjW+2nOLgpbf/9HphBdW7Q0EFYZ9r9gdCZObWobyRtUU89HxhYjiSkm
t4RLghBWxRUnGP/lG6hAdiwqg9Jqp6r4sXu/2M0jQ3FptuFW3F9Kw4wmPxbotltg9x8A4SGC6ebO
2DfBxaPcgIlhq/uxoduf6KFDJMlc5W+0oRzITj48laKZAkhhnUaM1Y8CJu5EzZCZtgrJrgUakRXx
RWS6W9OSSstTOcnTRhCW9Ykv6vEboe5KkQSU1s5losKQPaEYg5pl/urO3mEhp8+336H8W1sWM3Fg
8KaFitnLZLwslXLq1L3yD+YLBL5H1ZJdR3d+LOjuOArfknkayT3yNVYp0648352p4KBjMtA4kYjP
Q40T2DeYDQzfN2wFb1Yqz/qPEMKw+2RLAePBw7ILy7ILXiGil7PzSPrXje+d2l5vMKi4QgOgbtxr
U20H7hGCBwjgl+B+22UNjVIqknTmkWGAiYDdBZzzvjLEV+/Uk+iMzMlKrYeLqkgM+LWKk/4d2oYT
JMtqO1PrninATS4G8ylG70K7Tze6vcpo0SHn4CLVnNDCTkuAvTaU/2ivh9aHd2mC8s8fUIRSbIWl
Wg3flXIqCK1CGz28oXxeI4CcvQbt5eOuFpv+ZnCgLcRZEFVC3+MhGnLTyleZmIm831OakkGbaF5s
jrmdXS+EoHVx6swsYkUyMCEfwgQjoO4ViBBziVk41EjFuwtd5RpNdKu1BlCSL3GPvqwywn7C5zN2
/Ege/Y56JpMYDBZ9zg8/CM3bllBNZeO/dgxhTo53iSjaMQw1en01wUcIQJjhEC7/MY1RPhoQXSVP
FFxeJuds1e66wd07Tddef/pMVMnSSf83XrkpBu8W1WmhdQVBc8GHRPXc3CjB3AfjcBL9xJx8UcOL
6+bjZP0qBb9liJ0MY+qTc5JXxSfNuSg/oaPZH9/LDRfZAc1GHPsjOWFJ2pQlRvWZZq6JcXCZSKvi
T8J8VTEBGsw73JjIjSO4xCFAnvDKgaeo6bFTnTlusDqCXgnvrBhkx5yOG2A96RoNlwiIpyVmAeR4
EGh6lY/yTBF+eIhQQZMjIwGpRmhPgaHjsnBUbi5AaQLiyaSYWzXL7h6y4AF27qWQ/jdTivdm3J9r
lRRI1QLqWclbgHAQyjO7a6DaB3IN7N7MbFTKaPQrSey+KLoqgPSVc0opYBVJa3uiGL8HTg1LpDw8
0w0v1mif0APLvRc/NnSRP0TAkd7jOGCj+Xv5f5HM91UzB3DtfqPLwfP7sgMuwBmW91ecwb1Qq9Od
wJtMcNcML9HzDgTFfGBChN+jMWXrUXNeeGj1EMpVu7YpAuOebCnWZCPzoHEzDceRN+RzIfEqizPV
zUu2FRL7MNyCFdCFl6uvaQUooeiAWpZ2z6108mDc3LurwJZjWC6K70rIl7SkB4NxFjtV63JQmJlH
hJSRmtGDRsU0EPhWWE1f3TX9aGaylbdC/Zi8LmBTQxf7vIBKEwNrImaRQH+BjhgBimLfkkGp3567
B0TmKhGoonGchyXIKAZ2+LRQM2bYEl6ZL3AkGt5tiLtd0jd2QV7nOPSF0fZCAi29vUPPYU2jSWaf
mi7rhZQpmViWfHoAXqZqwEmk01DGmGlj+cJ3v/1AsjiTr77CtWUC9uUJkeFlW0gob4qMWeF5vIIh
3gt5D/UR0vo0FlEIAr8Z4ausB8Yq+yr5Til+maGwfs1HGcEt0WQZc/RtBVdihop8rnvus5luekM3
AtOw9dFWIfZcyWPtdiXMBE3tq+iPj0qOr68FA0SymSJL3PWkLgN9a2fmz2eNu8VJe9u29hreI9xa
eygRJi18i4drMDUMtLRkWiaydFEgekjzw+OTnZxYqZ5kvIBYCuMYV+F+2tX1wRzXGKFmQey6vlXy
ZwU0L6j99gOUrpfA2289j5WWu/ijHU5lb28KyhhTPn0LhAwOHAaRGhGtyZvn7XmbmvjSN3YgltoQ
z5tZ0O+vGp1g4XHHXo60cHHj1t54rZhU/5c5Nzzy7hbnhxDVwVWSbf+ZcHG9xZPM2Z9ZYdrmDujP
LrsPxGy+jItSEb6/V6nnFCh4FULSVu+vBXLbxQG6DwOWPhWHcLpYgl+ovemClgbn7hH852WINQl7
A4mH+NbL0zmzcW9j9akKGahcY17rDWvbpBJpQb96ojy/l+Z3CTQz5K/Dzgs9Mfn9QAw33o1+gCWP
eFrpT4juTi2tR0ERMnHRWm9/op82Xklavb2ZKEQm4LKHfx0IRFRs2enPWwDDCy1jHqz3l/8sxB79
6zheJ8lVuxr5ikaI5eD6yG2op8O0+bezIqCEPmOHfkmtCTr1rFdFZuAHivii+JUrNBrC5EUcPRfq
qjDMJ/4AAqsTY/ym0MMqRH+mmMSx3YejYeA9QUwSJ2fNUCxogpwqR0zzet16p3YcKwFM++hPmLsd
vvf8jPcNwflK5+CA3zOlEgtIrK6xMv7rWQSxHVBh4DNoEyjuItsIELhjOEL1UBfl2vGQrjsoBp6U
SeSqfDlvsG4sY6sKPuAotMGz95t/l/DSLWVPViMtK2YofMYhfz67VclP19nnd71LU8xW1Xsr8TsU
TE5ZBR+FJCdg6EvNv0APZooaDjPBbDJFJaL8UIwMfh1U0tvhFcuZzvvYvNz3EAfAfXaFm8BUofZ4
mbp66yGt1j0tuTyzDU82SlCGbRsqW95nfUsUZMjgfBTw3NU6F5fNJ8+GFKrBbOSTyIj9guiK4yKV
RNAjT3IIxdi+7Z3dhyRU6JmkBgbHpT5+QyLQy/V9lZDlSfJXYDHRWZFbYR8qK/TiyVRfO/rQPu/r
QeQ4U2m72tpWQU+5yVUTp/AkehuJPXIGeWFY4fYOV4U6jzr6ET4VdAwyHqjxwcbjDE/ZqSf9PJJ5
aBb16u9Bnc14BDTVzn83kVK3esqwm93OLDr5m7AAOpYl65bySU1/n0KdwstysFlJmV51acfynYMu
yrWwv+3dwwybMx+YfG6ZKZMbMZA53+EtNCy0jIouY2fgDi3riR8/4IaN2+AMMxsnczZCKDYxzrZY
qI1Liq/8R2vGQ0tOdaK4On1uFjNd7cPR7ynSOoIH8Tcx/ykz7ny0ZJAF3qdKlN3C+xXsJsS7KjQF
mNcALPSSbsLhkbVLIEO8cqpM+QmuXqLQEOqa8gl0t9AdSOdSI4ROn6lIE+UiqTF9HuaLRYZ0Bq3V
taPoxeHf03xk9BijxxuycPPSJ0+zpzOzBdt+kuAeOfoala6+ZbDZcOpwQW/KZwY6FCrbkD8nT5jf
i+GbvIjOhQ/Ti5fuRz4mxW4OKQCKw0P+C+Wq4/SMf3jhNDNZCC0DiLlcsVsnb7VeNFjiQjlYrsXE
GBjMjMhiDzebbyWVvoCW/2WW0i8KhmCJESB/p2Ip50j6rfDqmnliTMlIYTO6iPsOwkRIhiS7xkKW
1yVg02sPJMgsc0C/QQH9Ios5ZEZXzvGi0QN4aHmY0bmkgERksQftjXv/tJm2HHdl0w1WrJhGNcug
uadyUD9rwY+46i3fASuvosniphOdxgBQvYvkU0gHgodenH+c7MZj6c805VaGwbQKqRhEWK3178NT
9XC2KMtFVajBqxrwvWZwyxPn+9TrN8P6Am3DxAFo5rHGQpng1NvaAfFGFBdIjL9DwSkwypIJFM/w
Be9qHdsmUEAYiom/da3Wx1M+j4Iz/l4T9pdkN99qJBwtdkvZ2nNW2hoHpXFEaILI/Z2PAccgymSj
ZbNfODGuf6j3DfGa5VnNjyvRbqf4hHxPnSk+JRY/7uyRSTvarQFwbNUO+gQ0W1nwdHmuBTZe43vF
+NZwY42uKrF5KbYkd7IAUVGibVugIdIdC81XSBfB0jU6PUzMiSCOP9BbytJo+qCDp2Um5C6VVhbm
vX8P9noVxEcTqbiJLpEIcT23rWAdkU9OpABtFVPd7GyBX0TMYQStTRVKkfBqDqiderxa0Q7+KexE
VH1XOKUPJKaSlZBcCyXKMTc4Atek8a87JeHh+zPoxqKhS9Q+WAqk4YJc1eDOrJWBgWYpqVu14iHO
c58R+T/XSsOzPSCjQsIIHaDcGy4KKuZoX/XcvJGhcAdus+irnBVPSuFWAuFfkRtb6fsXDUrquasc
JlO5XkWtJOVwa4ZzRdQyHuFg9JV4h2on8WS6wDBD40ap551K5hE9Eou2T5W1zte6AhexKEdMsyvo
/19qj6cfKHeDaE4uXWh4T1xAovkxdJTBAvFkWIpuonhr34AqROjwWiM0uOXh/UN8+rZ9xFIjTUnC
gMCi5LUYBIBVyw2tUbLGrrSRiqG5S5/bMHhnotg5H1dAOAV7nSr3Vq0Y+4+E5qmBuMYDfU2Lp6qN
Vd5UsPnBBFG2mS0SQLHJoP3zkWDuUYxGNGljwzjgT1mh26DaueA58mnOwZWG3fKm4E6rVjBZGI0M
uT9Drv+fO5/mNbk2yvRhRqALAJHTz09RPQNcPL1GzttvrF2IenMIiXKZ6FcQfEjnEtZjs6ZSHIV0
uFtiWKLORr/ntBYtyx/EKPrjDqFyNX4Cv/i3uYdYwz4BXQRZEsVDhojMS60gQc1o6spPWD8kn0qk
jKfRp83H8zbYbfQJxYqjPS0/gTsHV8EvhA/tts5vggHsFqBPKaECHO56DouEt9yFWVZrlY7El91a
MlMp27chvW6z5Q4AZ8hz84rR/E83Zv0s9x0KQJh9bMo3iW4/DYfsDOKBn8+k5YD90lNrWJk62Hfp
3cRjqwpIVkFaHusgzrBFNowaxy82/egGmm3RbH7jI5rBEPvF7Vk3bioS7uz0xqGQp9Pgscj0aGor
qwvIhtnZM94MQAQZCcl4bfPcPZ0GdR94O0STTS1EtL1qTBIiLcxoNBkbfZ01QL+pEvptWnnRG0vD
soQaWxkNddznMIFl2Ix95SOXnIfeoi5n1B97ioESg0X+C34kY3/BdW2paO9X0suS3DXjNhYXnam4
4j2Fqb5Nzs1TtfctGlghxZSznQPQQSH9k/qsT+Zr0JSz/LBhooaFa32oHifTWV+PiewmjjkI9wh9
WH/uVUftAzNRWkUtheMSA6mM7YP2nEJM4oldmHVQe3Iv3t8bK8DupjaU+02HC3zoD0G8lCVHRsIN
eUkPTUCUPrYMN5I3Kw45ktjjJ/Ul7HWKNa4SOjsdz6XW0z+8rIFmfiNM/S0/YklwBDTEv5yLbo3z
1ZTlAe1dBAUaqQ0lVxld3+/TxiONtVQvm2KQONmLYYu8OVJyjojQxl9JqMzUSh8g/wG12TLV+u9r
w2NaC2sjZz2lStSCjVDLQmnuWDG+g3YJeBiMklPxt+7+DAbs2cWO/zQswjWpPD7xzNPCtZTK4okJ
4Ov+P4UClxxdo4hmfT1smg7x/zBR8h2Zrb0+BbC3tTMWgfWjcsCjYq3ao9ssqJENrUTyC6OQdAD8
TJDDFe7Y9Hw/cY+MDEZyTC/MYQflQco9x60nmUQ1ogDYQBJMewteJ+fbPaeBRZyIrFWFvohJIhb4
4o+N4sG9ZojCjdwJdgWv5l7Ce/PXnP0FQ/CsEXyAgzJdjPbcX+mLJukcugQsa1Hdav6ZTySmGQI7
r5VScV5KLpH9r4Phr6pWfPZCIJkgrF8H80zaLSmhdSnPnGgcZGYKa6XxoptWd9OGCpKEZ4/0ibIc
CCwXuoJpCHuTenXLQJcz6h7DjdqNoVvXrX0ikJpmHfMNVF+Nj1D8WoY74fZSvhpEHR9/d8MnFmNl
BQhdmkzZsk097OjNQQvFqyhphulu70vApUKJ+R4bQXkU8SdcGoEKM1mJJ+fvz/0MtYELtnMbi4fI
MQYFtBTdDU5Uyrzl0QoZFWgWGCgfkT1c7dBMvBK4yEs/tf9cSsA9lFC0fio/sqGRClft7plqX0ys
hk1l8DhAChWI2LihBUI9OS4/+UDQyYLCA5/WOjFQnjEXxraRVYokWtLp8orDJ/OaEv6z2vaDntOz
Y/fxUAWZI7CNbqnySy7b2gkhja4SAgKVBfapaE7q6Fts0mvLy63YXMAbMycSgll0752Qwq/S9G1z
qsRQfqB3jbsph/yYMLZUslRRLRpyFHoFrVWYVQktxBsyIADX8IrKdsMOnwBgeF1mNZH+707M+mEI
UgpF6sogbLPTasz5zZJtg98E6iNs9PJjBt/wo/TJ91Tb5LhOHg/BZHpZO/vo/atyLnuQa/NItNqr
26EWTOqR+smXG+azScxIMPuYIIWMckTM51EB1EI84MWPYfGNAlqjhD1vQqRhhqagdgcdB4nOuY8d
x5bj2K+dQ7N5Rx5guQlgyUlr3RHjp37URA1E3l6CIvhpiOL9U/rTrv4aPyJ6qZlYWvogP6/Al//N
RwSDiEvDsbXqedd1SakZMxFhmD56eVoogfbaJZXx5u2BMy3frtnE77UwdUBKzSdCBEhS02NQzlOW
Y4HVekdLWDAgYrTtz+ZozOtF0+0TDXzVigeVYCFbo+blPmOWZKy6IxAUeXJoKK0EXzETyIt4uNDS
hol/gScS5l1QkKONM9WPeuDQEZQ8hXc8Rf2vdLgARd8X2Ip2ILV2z+6IbmMw0yadZmAmE95bgzBT
5iZzlHilA3uaZS6WYdBrlih+DtP0ZY0gNZggK9xwC23HnDMxo7gX523LYtLwnNNe3yBNPTQnJHDV
lVz6IPfqFZQwe0g6OAFkVDdRVbgDFa5+CWS48DpgBNCVQxUelltHtDBM1N1L6utPEjxRSDwQSfNK
ybHXgsSPiB9et8jaIoUXkIF13eNLdKULbTQ35mqd2+d2Y6VwBiugzCZOsI0y67FcQEAi7PXyTDhW
ooKYMF2okoeG/NYBnEnvj99bugyNQm1RZJmZXiwikIMiI0aZIpx/tbaAuwq45T4S6UAiykKJudqR
6g7e6+mIbweHOMW6hqQhT0VhEVUmBUYWDAmdjMXpDfw2tSyCY4eMuThraunFqUtCeUlq6egornGv
5K7L/o/nFvxiNAjMwCCrGGqjvHSoKtzzJugNC+/oHlrju5oAbYwqRRZYbRlH/oErhjL1+L1GW68+
fvmmxWeE81WHqafALo2OeiuflycRt1nmgOnzs2HWBOCaO8jKD/2jvtjBaT7bYMePCezNGxanc4mu
BGcCL9B0A6Fs52oxC1ukiuDJv3JdgMWuGHXzURGf8Kvx42F5yumskkYB747VKuZ6hy5DhiUAAMnB
GvJm0HySrUv5z6+bmTj/tGRNcObDwTccJ84HKlMHbH/T99RNrEMgUDkTth806BWTnvsGNhn9VCGG
YSintstUHsdBJgIWNT1+cCtjZ8r1hv7hcBcpHiJoUaDaOBMugeNZ9Jw2tLc8Mk6GGkqoFXEis/nf
Gu03WJxHTbGqH4UNTY90AJpZg4TlFOUjk4ebr7jM/zX2+hS+IDrbZbjKwi+lgw3IXp03j9iQkOBj
FscQY7V37AWeu+CYPy9NFrYJqXwu36XXpxqCDOlJ/klEOqk1extlOMeDuO9PdqVjiPSwUbtFC+eK
f8iCAlfNghjyRkk/V+WDJECNHx9QwjJu0Q5Ji1WQ4yYs0H9+Q4BYkgcS7QUEVj+sa/CN283a45uB
LabpYRciV6RQ1Vm4vxg6ujlj94T0zFrL3ppU2IsfOVeGBQRC0VB1St6Oly07sKKYnE4+6KCtxHik
IbFCPNWGlhhmiv0av1yxN6+yKVpcsapS6aQLaHmM7ZmlOOZiX5SPWy2ZekEzyGzvzNTdTq05sG3J
mkklWvSICrhsugVlNw4ZYmvWQcU4NMMn8+d7c6NFAKVTtnhWJVnq0lRLm2HZVPw5IQX23KQ1v0Ge
xQJFDfgpgO9a1B3i4b5cl14YwPVj5HMPqLSsQ30QOHtKCgYJF7xzQJ8bWSzuKr9unopLIrNsxiS/
rowzeGZBbYniJ5s2ij/m6oKZ8TqXi7ImxQa6Ha2MgOlYr937frh0ACGj0qzY4vkvTVz3ASkMaa+1
thXtiUvwoicR4zVt+a78lXabCfD3cDOwS9FOD1iDEUociwb2tjdZ/33tQ7WlEst/iz0cf+39fesj
k3C/g8DCehkFHxxJfDIPR2d+Ta8ZrFTjDNMj9dN8A+/d4M4TjYjDtDxfKYskVJBpY5q9Ym107wcd
0Ib4hDtYmTwqh7J0mOAMO1i+1rro2gaojma/1WII1Zz/HtUKSl50NV+5MzGR4O1SJbwlrqPv0RqA
X9mclbX5GgV0qGCRqMChGsk+X6ZRvMe4WHN1t7W9mNzgONoSjyUlkORoVg5hFAoA9zfLJ0BlhvwA
IhhZoQ2U65mgOI9anTm7DuGtcM7rDo+claM2L7gMdFiTnyrmjeCxAi2dlcMllktZLqDTP9bv0ABb
kBWoNZIUDIGNJ0kptTLgmcD8lPO1hQNdVjbx7e3n+FudJtOnlGzXmiz8jxXnx88eSP9wNG7dbfjB
KwUzPKH4tiWQRoZOmSVKtZo2PjdWkEukB8ZGx4Mvo8/6fJ8NnqPgg99nBPqJpHVWg3m6zE8KEBT+
asGppmI8iIF9dfNDsuWXejxHE4wgekWWorQpVuKrEiKN5OUfejdMAWNfhxYoJxH6TNoms8tvfnzk
8Kd4KvDkyozjyael4ABzfDYxnbS4qkJQEi9qU9bJBBqlV2X5pErSyrHGAT4tDVDIXeAcfPwBfPpE
XT8LG/uDrGagNjNCsHmvornH0tIwpRrFXVOH4uHjqDo2+jDG5mK3zA5Er/KVi2SvhdbFIZ5W9rbg
OoMXZNM/z3vfCg1DE5rHc+gh7tg0tYopbYE5e7QHodG1TiBMpNi3qyOrAKqyNyPpWWVwFNnHDgKp
efM14I4a0KWzp1DoO7LQEgcknfGTdeNdMaRAr4HvKVtj9gsrvK59Q3mOR3Ha+tslpwMYMu5LlKlv
GLsAnIpcp4t64yDWFviP8eVx0mILyq+cOqmFi7sc6KuYyNkVN+ttWD3ehA+k6P2s1vmVd8JuUqmM
kUYpM8rLemP9ErMdBbxrxRVn6GESJp1uxgPGr1mn8ioNGzan+MLUJSE8HR57ISa5vlAiX+CIss0X
X+bMs1wUNqRxpnZoM6ze5RuQkgprY7515jTH23dVbBvRARPZ8jmBNzSUnAzZhIzGryYLk/+oduGx
QGIr+plD03ChyFyhpH3DSEmVBHq7KgAsvMYpJpXJbJh0X3KExf/3vbUO7+bTTszvF49O2j7ztk+a
nyG4oU/MgFs8bYhwPdYL0jRVy+aQKiZnPzPhspn7KlJhqV9bJbWuJySHvpHP9ajg/f0dN5vqxx3q
fTJBrapuJeUocIec1BYODTH8F+HPRTvNjuWQEgkxWhMdqaBqaqMn6KebKXIav4ca6KZLbYHPH0qD
KxcZRozEs8Ta4M/Hp6Rn68Pg7Im8TEAMTjXBeuAPA1XqMVgXzKyb7us2K4xlAVFZubmFBN4/vou1
xboolKiKk53BBD+RZ5zqE/KoVBG/7eirSjO38ohFSbnstFi6QWVbUWDppRD+he+IxzeGo8Muw0sb
RjlSDiVFVgTNT785L9lJYDZnsZ+Jf9OkBJgzdml/gDKJ419fERul1UzLWCG2YbuwvKSUoi/yt+gf
yHWsm/8JOJgnHyUBqgI8yg2ht2IDESZDVuOTR5RFxwdxU3UrCGEuweoPqRutg17h4dloBHtzZ8Qw
qIxGCc4/p6xKU735vgf/r5tVUuonfqtpRwWyfG2HzwDPjdY9uhaktKMPiHRbt+jGhwH64Y60yoJy
e68Y2AL4RRcxh9SILBAD7oiK6lJtJ8sJasivvvDwSZcAo9J7L0Lkua+MT3bsh5rtepMfgPk+WyXY
cRPyxwf8o310LZuoqdwARIfc0Ah5GJGvqVxBQxPQs7C7KTAap+MnJtQwuD75adLRSTJfTO8oO4iG
0qba+giS2tnkW5QnNT72HHPXSiKye/f8uKsoMWgQ8tAGHCpbkJqFj15Dk3qFHrwwHtc9hR46SYT7
MqA9rCU2aIwSZ1tL7mKjIvX04jHU0shku/wInrkqw5177tJe0SGF9cGrT7IQvDwZgHEJkkwfTdT7
HIoB7Qh7ItlgSTJP3MzFbVpdAlbg3ftSffdk5r31B8+YI4+VGupLa7lZxq9aNxFpLnB1ZzPB0I0q
G1zLeAsq/JJdxm55H9LT+Km/IynDf6PrEb2jF2WzVPsbZCRFC1ERhppa2R8+wbKNTUUna7Ylatx+
G12e9/VEbBOK0oN+ajJpfGgp/EZodotlEscx5ALQP6iY+A1XLJ9H0IXQtufu5DNmlfBBEIFR9zY/
If6mqNIXIfZEmTCcLdoeMtFm5Fr9mytuQQWETdiuYVMTMrvFJ1DExjZplhFCj3JIHthMUy8/1lh7
GYqn6MV5XMcqax+h34J+gKxosCGolp0pKDSSy3XElNVM1YqvlykBIqxXWLJtVYrQ3g59hkGorCNj
ig3XdieVUZUPRtT8gPllAkY9UPG9s11WUV2DsBHBClzfJD7vLHDtdChJ28aCqFetGNjZUtxCxUlN
VfCW7iEhmpURqB5bpqW0srMZknzbOkRzSCEMzzF0kfdXYzBgJkWyoB9THxB4Q77gFdDbzFWv82by
NG1sfQZFpCe2xyFKLMBrTK9eNQiWvlaBPxNXFeFEMi+mWE3HoZvxVAeG0oFK8QT50hjNXLckOuaG
xiCqLtpcZyFAb64JtKMAp1fi1W3uqlZz1fO5Nn15JLvOvbixDjaI9h/rHLlsXKTs2Mza77Ve/y68
loOWQXNuRJaNY9vqjG1CcvVzs/p60D5cRJBTKBWJ4wKrbQunIIIISxEh05TnCCFICiwB/k8/pfoo
cgIZ2/JRARuYpXworkF5idpvHsKvWRSWibW9FmBSr6UzjM/r1EpTJ34EwzG/CMRqmi10rAht7mbx
DhWdJtB4ZfHItTt+9V7q7w4FXS7SRxcC7b9aIl5K+mVjvPdqnFF9qt7P/qmpAIyn2dQaR1M8+NIc
6+JqBgy3pHrlDFU/RifAl/key65HsZMHXbW29aKJpKjhu8Kxoui68qdXPXitjn/osMI9SwP0O9GK
bORcgfyB9clpnpvXOBuGe17fg45fsFtC8tIgJ5++IUAe8sPzDAQ/Ykc/9xOmJJ0YLLt7FGd/SXF8
rbPzRTYnqOjCTMCQMbQD7ZUdsXkQti/P110aRfMUv+N4FyffeNfaWLdMxZovHEKu8xCMui6ohoZ8
32y9fmgRDMvPcZI6YiWrX3PYqxyiV/X5Fr19UoOvaAMfv6Q/E3nb+0x4b/fsISxZQLA0oOXtybCk
yzEKOBG7oMwCgoD1FAsNT0e2XuLUR2c2pzqyrVP7HjP8HeakfXPoTtX7z2JtjgRXr8ekeJ5BMR6D
vR9jAfaTwkw7gQb2/YzAk0jRFM6O4LImc6NLHXvI5CIN6zXpHSouiE14ft5ExnZmDEOnb6ygL75b
y/SMz+fCJmHH5dCxMBSXWUPToKpzMnp8H7qDJ0uWZKxtunI4YZf/oWnAntREiU2uTfIPHZg/6xGr
Wx1JwxnoYYe765uT9DlT7ssjC3eWTt2YWS0w125zltrqL6atfXfrOR67qD2cFn81gHtqlX9an85s
5rjnsWmDScKfW/cyyzWxF7ZZTQ8OQEodsOV69YnXevYUjKCrZz71B34rME+tOc+F62Ma17C3I4Uo
TLBtkVQXcmcb89w57jniEm+18PyocYsfi++J9ndGZ3RRo2aJyj481/cC5N/Nyl5+KnC5PQJrbpSF
fwAurKpf2066sY+dgu1zfXgO1Py+bEnQE5MQqwySznYOKZ8MQd3vv4DmkVEzMrZh1sAEou879SGt
H9QnrDmqIeEzhVn8WDflCIks+HQlL0S4790nfxrdMbgw/C+GoFEZDE11E6MFTmFE+sqJW/9E7DX5
+vf007hkoZtjArBCuh2VKog/f6bzbUlwiBD+UHuoQ8a6TNK/JsuHAg8O72xFXjWaNvlJicTPWz04
BE00mVJoiOWlnGzQy0I/fUFPC6+rly0ZlxbaaAxdqLlzwJ6dXzA17iRgdkZbbDs+zhwK6TGXVuqq
JIHSNhT6zgtYHiSCOfoq2E7W/QInEkyZ0byD8EZFPpcMwHY+1kS7NwQY80taUZcQfVXhkHuBqPtw
l0Ct7DjDP0vkFyoKQmvtpsulDInIkAxkbMFPAiHOiEL3B7eKDVFG0RuJyTYew//P+Ej/04F7IpUY
6niOb6yMP/O48byQdf1pZYsu0oH00e4d3VUz2I0NfTRCGQa67oPuMUgyX4uJh0oxvJzXmg9diS0q
RCZoQvEhJLMemO4mKdHbZSGNwM8OglT7qH7wMp/5QDHkedkQrenl+1+vJfa90GKt9IqN35ZlaoPs
gX2twrHo/FPkxmPHto2hnBYtjBKXzFMoC+/PafEmTNk6ILpQxeXRPl94C2onb/jf0rTsgbYElsnM
attmv8pzKt5OAqF2P8CAECKO8OOPJ/cPxvQduVTrPm2FhPtFpc8wIYHFuF8rXX8wVvBzZBBEwtpl
K8PrHkcIJZVbLBip0l1heljwF3m4l5mPUZwAQeMcDKIFm/rW+ipFSErAmXqG8s96WmEAzT3kwfSu
/14CRdW+i335c0SWG75LFIXBq5+SSunOF9QyZbVodCNQiNWwYXPSJeVHlyY08fyZePQ5wGVT873P
xmyf9+PYKjX9R3h/BfyE5TccZXnpJKn5VnbdeJGkQkVK/4x990IpQXwFdfg3Cl56HjNBh9f/hpgN
YEu4uL2GM8Y+H6tR6UhpJ1Y4baaGco5UTMcT5Z1rPcsy1s58z7tSMo2/W34L3CA4Sr8D4uzTG0MD
Siz5xcvlMGZB2doyn7GOrjHkEhuHdk64x/tRgo5ugLaPDgRg7Nh+Q9UA2frc00/28Nv3OrGn5ePp
4mLZpsFpbhGPwcww07AdqnNq2+2TO0ROl/xzXzRyoj+KbnucfDvw4GgLImSEqMDuaTMtM6Bbxt27
IyHHBzFfuvVDx/G4qE607eXBJxnmt+sQuvoplMRoh+xHlGHJm82KPdfxNR8GKgZT2Y0gdYgJ52Kd
nbu2bF0dpB5UZibbnoeBJMqQBH3QkNYWgp5+vkwP1mOe7w+0AtFbSKT1qi6e52XyEuP602Sle9A/
5irkRX11FsEaZcxOfxmlMknfd/EmNgnlYZ/q+WgWAgI7Vvc0oJXOCfJGnBMJ2Qd6evnDRZMxTIaA
l2UqKPqZgROCpHZy5MeBYsuDgFLho9T1QZTpSxKWV8fbPk/fq8G+S4LljNeFFKO9H1VKXKlRV3LO
K3ujqNBPdjgsDTdFAMjapxdE9SV0BtxbmVHvgFK77E/duIDXRBS0gBHjOkewAydXcKCtgH/gviGQ
14g+BKGab5d8RPDhCMq3xqyRAWpx49Psb3dgZ/CaVWpIwgQDASLAytyECVYEmbHHzRy5hf/PFwa4
UcKvuPurlX+CGetzjsbWyXxW4mbQrPSfmRUoJ7D86PYnB7Yy1qoUFXNnUcHkz3pxVFcpSlXn6DGV
qsuYZcqF8j0LYVv7M61xNp/RCd4cGS/vDnBSWLFg+4wsVbjV5jhxNAS9LG4gEMEYJbgl9vRYMDcU
aUzfUQ4yN/CUlMZ+YjGsln3vMKBD18WiqtOcdYzZ/r1TPRKU3IOQaV85etOhdyRZMSLzC9c+YSje
FIiGO9pVhQ4Zif/QntMP170RxEQJ65peIj4Wjyzp0bpKQrZj4caAnG/Zaw3ffwQqZHxByGskatih
+8Vzrdop/+O6FveHum76x9XzIh1qWLyka3b4z7VjPunH0iCok18c5Lp/cJiRinbtLPKjaWA7o9DQ
MGT5q3ogGepwK3CVlebFTmQUNzscJ99X/HevmOpipnerjon/S01V4MQfmOuG+zO6mP2NkgUKWRHy
PNbVGtKDVhfVZoDrFIatVHXMXNLFzYnKqnXPOE6bKNqT9Baf36x7n5wRKiYNFzJjqhKs56hHfUU0
gLJyJs2g6Wn+o+U9uSsMLX/N6hbSEdI2NfWphA3777JghCsymZVKTTP5Et1SHXt1HAg68isZ8WLP
knr8JEmBnINEiNBSO2ic9d5dWI4Z4Lp5tqIdy5a4fR8gRWfQqmBrWFlxgV8+QirKY83dIKrFenBU
BHR6XSMi6zbXhHLUpN+OD4zdX/QsdGXItYug3Xzv+8j2m3NkCanQhw85Zana81fPnZfa17juxQPI
eyNee+Rs1hlMUK9bh2UPC82qF/K9NCvOQJrBDbcDQ8A04H203je7zpWU2VZchI06M888aUsaEVW+
kN8W3dd1gEvsYCE3nsZcYG5NkFvgXcOYcIzHhrW9k9eRfwB2ODxbETCv4qSXH3XFcOI/l2HyeTor
VYzPR7odOLLT6p7roAFYOmMRFYCSyDdtRFcf0TsbtaTIDhkYWB5mpkrw/qdKnN0XPSNcbkPoEWob
GCDpCNp9AXX/2KuQz29eNeg6RptM6e2s0oryhrTClGQrHRtiNY/Lhztd9QY5cpkzmYgXhWAssx93
pkqPI3OZSkUxBG4Fj/gKwaus6OAyiEwrN8/Gb1MqmIZK97LjpKfUGTU1E1dSz4L556lZdOvAP15Z
CTizJQ5nTzehd2TqGIg5W753//6Rc5CcVMD608cXeOrtHiw8MecQFFuTbAuPyNzouOBQG70+LMUs
MUqFNGV+ek92s6cPMy69+NWCLZ+QeFsBria5tVoGf8MHGzRmJiWMQjSRWYUFjOV6NFVm3OQCI0iZ
OIF1bet7FNu1wJLOWhtSdnr/uAM8jtmBf5/Etkd88HEqK3XTSB2s4+q0+qSNgsxbC7SC1QnYdWEs
CWXsxNcek+4TMvxv6S6UpR+M54KU+4Frt+IVYtiphJjjxaM7LaTNQet3kYZFnuy4EqD7SDES1XPX
D38wY2pc0fSezuCeRfB0BQx/RJPsAz40JEWELS6qbqNULUs8VHWUTMwVSHSloH+tKhstV9YUeidx
C/osoACc/ccVwDrmIIkH2ilwFHVAaQf+W+4n9VIg7dNxSGdHVu5G3PlbjAQg5+6/TweFZeyoRoXp
CuMR/tAZizpd0/4uNmOH9DzB5VLuaJ+KIQMP6t9SebGy3bpaWGg1wyMn0pr1rPyy4KyrSWlLIfV/
7pu7uIalsmW+rN+naB0yuGzrYprvHr8L55za7Cls2IILBa3ccHT6KQGoyQkGgghyNQ7mi9NmB8TF
WMiKs9ATmpn4cLucQAnjG9GekXZnBghoCClx4Bo4z1ULw9X9w5ke7tgjDrdDSd7WwNxxuswHu99t
5hXGJJpMw4X42j/Nr4saffolsDi1/IXBJZhoiAohuCvo7AvhciiTr13YkT091aHxhcB9UOG88+wV
uN9bkAlmU/yIDT61TRIclnt/KHlS1TCvqQDhj5GLT1kEFuONF/wqIqYow02efAetrRu8ESXiSdDJ
BGa+0vpvoleCfJFGz/2XSiEh8Nv7Ixzfkzo66naVZ7X+tEVNnPaKYKRRlJBkV4O6d1hLIVBuDNBA
6wdvc4oNf2Wf1TVM8TQAnCv160BVxrHPvp96zCOQmLc5+wShwbHKQwW9EfjLe0/D2m1OntDWjeDI
g2vjKi2klSGlwqdhymPtcAVddtC98sHJEwjR2YGgiF1vr9r0x4WJI3q5amlrw3T3alhhkq6CTCEb
onjxUYyDzNzTmtN+x8N7IHF+GGbmfFK4n2RR9EnBvIWc7N5G3bvUZCevDuouLQHmIY2P+Hg5HpFx
n/HRWgVInepx8uKtcAdOo1vDiClDTr7hNS2hyfa5eTZSgxyiQwpQNBF3MVDQygcgwhFn5ehUZfQA
hPqYsPKkcFSiIXFiOISAusO+X1a276T/TUI9xUrSJ05f6D1o1GIi3UQkYnRWM9UpoFUCWn2/ahxO
FDYADg9qfL4I3JH4OvjsTYFfdiiNZ/0tx/WdKVPsWpn1VNzsTJhiYIFKTBUriF+x4ah+jWYQSI1S
XL96julOq6ZmXukCWkK5N7RIu9STzfeW0cNmHKQpvNxBnlcxw1dLVdolJMAqNVT0tnB1PWw1C8JM
Ttyu2c7iIxAlP6+S3skl78b8LpTMcuitncfQtd/9vG+oTboGwD9E/Xt+/k4GxnkJDjUxJyuZJYcy
R5Xdh6JeI3W/dd7gs3Sw0E+TsBQKxgilDON3y9ZAasdXMurDjjPz1O40ShW2duEEd9j66XB+CCvQ
wOiDsnokh7/XfTPri6P/Ljdv+8urCU097xi9fldEBkgXg7Dkr7SLbxJPfnq31cpIgJhGqiF2faX4
NKf75rQ9LakKwEosIIXeOcQ6x/qsd5iCM+VQrwbO1rJ1khnJQHxtIwIia5GjlRPBf38VtnrfU/05
jPQBFscUTQ9sfemfk0trlCPP5Qlw0n/SzHTKWSNLDFYdWbWb+syCkuOO80mxt5tJDTcdl36GlqdI
JmhBBfBy05Ql1zhxCQX/+0aK4YShaH/TbyeeUHEdO5ukru0fs+8zsVqMlwS4wim+A9UIfd2wNboc
CqPo95bMSXxSTrrgl1Ez6cvv1X2PJdjsNPWTH9DBH0znCNqdLEyUnHn6M+F23Uwx3OwHRwr2Mu+B
GTA++MKeAlf3jGXXjhzXoyA660JKXNRPY0YuaxuBUIrDOiOu3rlE9j6qD/gprfnfyyHvdpjhlljU
yDtehGdwHFfgdktO1G55xRc9hsWsFVqItyL609HCEQYHrKnyni4g38QofoBiZq7ZArPGYhpCBY/d
pfYr0b0bHb37GGpkiU/MWXW5KnAK3R9Ezo3k032sqdTX7cPVENE4HaFJpDqJHdWZRwZWqnDQHE7K
4nVRC++R8oULuXZOsUuz6sAxyDdQE6s+XHSHxlcYVa3CLDjdW2pFBaT0jPkZPR7UZJ+TqARAwah3
yO1Hv0Fe5rfmuZoEdjsNrQiME7Q6Oy0JwG1cbbjE9q4wNe1xiQdLo9/dJrqepK7hslFLeVVxPxaj
qxMPpMH2Q4Ejfla/smPU/5/KJIeUaH7guvQHc5lpFJxBiCIa22OqMCv8NM28j7hK/go8Ut2f7M45
P2BtSQccoqQt/HL7/hA1MtMeTIJcCLV2Q28N8KkXPXSXeLJH45Cz7VrAKMNZdoxdfoLlvKPlflfL
b0zsT+eL7nk0VkCupJA0BUnfeLbraUuh2mUZGbAq2zYPlP+kQ8Buo0yHUSGy2G+1C7ucnfYYAe3T
d2Qf4dEdhr0UDoEMjkGGyrhYFGzigaWPi3pbj09S+k1T+bBLJt9Yi8tNGN/7eLoZMQFzEsnPm4BQ
+6IJbH2C14RmrMFNw9jZKka0C4V5a6C0AL4PCCB7JZHr9ApwNm60OvRkCQGNeJMH2I7vUp3Hd7SC
cqVhiPHZGvD9x8V6Fg5Vwi37bCdeeiNlwMH06+n6+bWvl0QzfC7oVSzKuDY+2o2LPLvG1v4PYuyB
QnMUn9nIW3I7sLBnA8/5xuQrJO9mwGg+gHwK+ABukAnxrVKaLZUtJljRGgv6xUOnBKfE5y73BFcm
MMzpbMf8THR5Z3PwwkyfY8pn7R8kn1lv6twM9ONczxZMNNwT2YqQLImMkYn9gCK190K6jxkLmSE4
MaAOfWf1O25+UCFh7MPm+K+xlGSlbe95qP0ltaUOU4HJoWjWRvVz8r7OJAHypu4hitoBZu3orz9j
iqLoWkkfmkL01pTXbATKDKKXKbLfD0nWoPp7W7z5bXiNnCGg6BN79jAC2rHw5V/i6p/fp5Y1zfDB
QysfkzXfH3heRKnFm7XkrjQgsZQGsA0ryXUe2ReF/AMRW870Wwn8j74ljzQX/RIeJuuU39KAZJoo
oWum5o5tq+8KvrT5z5N5ZYNoXP4XsrEkK0et9AYV/jFzSFPi6AXpCWlUU2ezgJYDCxc0voA1DZFC
W+Pn+dUOsSJ6I6vrTvzVFLYW/RJdZSagpnR0Smtk0Tg75gEDzdf4StxReoL7jKxOZ1K6KYQR+8Mr
cg2dY4SMKmq+REvu2WY3vhqDZo6f5fzFFqZY1P+ZZywehTXSB4zHkXwPhO+8U9fI4pmm1hRB4iIw
j9NzYTt5KFpouQfF6pbJiZ7+x74EAH9D6XVDgSdiX1lUsLdQCHyUg3/Pylf5AnNXQfSoJh50bfQI
pOal9hKlUVvQnNSoEr30ZJZNeUpdTCqfWGRrYYGgj/YDfdbf5F6Pzxgd3uvogoHf5tMmM/OCgnl9
N3cjE/ZaViOlS5c/z8s6CNRLEyhlQjZJHOhU0DKxULMYF88QyI1M/tszYzcNEjG+COp10ILeKUNx
83tTe04WOAL6lX1xGGfLp0Ots2XZRdnB6XrukRNl/TEe1ygeMd81gm8A3m7KfAu3n1Nv33flxjcg
w2ntULSbRZx2AR9mOraHrunaJp8t9q11uupJBUgWp1gS0/DwwLucHvv4zhOxdgtLQWwIAv7ITdER
8Hr5AK+M9AL4IoSkV9Cbls62eO6NiyxjjTqQdqKdqBMB0enfCFCoab+T7SJFRM2uXJ6s2h9DeQtN
ufkMmi8VXBazpGa2XGZrc7nHdVSh44zzmBYY1QVOdFHpKv2FyBimZN4JYwYsQaK1Mn4NeOH2dG+1
mbI3sqdAcF99iqColdTus1VbElhhYM987GKn1fbvTalQ5zDX+TI+gajMjUc1fEALD6E+1KYtws83
9YOWuE8TGY9hRdYzX3CrJ3Ul4dO8O0M+W6FZZ7BRklaGMYY68aVgdfbLAGCCTQXW6qnqVpCpqbS5
pENG+lMQrMJeg/0i/xk4O1B5xnD1lAV4IkKO2+8abrbxtXEUBVpjR088XLhF3w4ENzpI+B34wmHC
1wJOeOEAd9bZOqxVsx80M9aW/u5ETVp37pQUz027WeLHE9/VwWbf48PPu7y1R9iH9JgDINfHhjWS
OqHyVDG9pmVjXyz4HvtE2Ftq3AXxHY12uGcKmu2fSr9xRVS1Opdxlr43CllM5HsW365XwWvgoTYb
9fbdPmH7x6keTxmmfstlLWceNgoFbeJ2pORr9k6sm1uFqkUO5NbwCeNYWsmCgUa1/8ga7uqQ5GoA
n0n9hMaSFsj4jvmG7RdCUaCs5NDmg//5+StlY9HybWz13v9FIlMX8s4BMSXQlGRSMFHpTNlSL5hu
/IPAM8hZ91YYM/CSevOl0JMWWLR1QVwop1STNQGqxwWecI1ppsU+Gh5XH84xdEQkx+NMo/tH3NRc
45E2rC1hWNsLkwGkfwVom3EscHruL3Vs5ql5nP98ximPqQHkLuTOHC9mLXIRbVCBbSKQi9IdK4Ts
tEassNtKtM+G4xFwNRTrDP7tzEtwvtNg5vH1Cef/mB37LS8XP9uKoiNqXR3UHvCl8E0I5lzj+CB3
Pqbdo6W8/LGxurzk8YjLcZH1oIAgqqo7osppYh3+mFKw42mubsXN+kiwkyCi/0S/uI5I8rXX5eHd
2MdNxnKywQb+ayC4KV0oCqZ846+9sMeVzd7IlKNEeUUI7ZCC4tIEgIzHuQs4zMcqsSxf7qXhva6p
xhIXmnPiWoRDXnTvv8tvDS3BGXwud3J4H/dkZi3qjwMd0Ydb9MZvXrbPtWhQuuDug1nL7l3OjuSu
Dqx3eLynT4XpWvQf2bWq5Gs3QhpmZpONspNyipGg7BqzfZKZMNvQ4qblP1lsLu+mJvGP/BUCJgmL
5mbXPTgT7i3joZ5TsIMEbG7SXtohcsM5pZGqpxz3wLeMTLD3UDXAXGT0P6Os53cW6UQqU//fvyN9
YrRsF++Hnzu6wYp30OaPhdm0RFWy+Lthnc4OOebYSceLcpWGIFuyUlcq1EmlGbweDLIgzAns/IAK
+fR2psqOwcsZHCUvaGXYWzQIathK81m5ADWYjw5+yhsqCpj+34UiTIqrdogcmTZ4JhdzSX9D6voN
jqTLEMme3P0dvrEKjZ8rogGPxtWSnZ9IjcqCVA2SFjjlW3GR8Feh/4EbzI98oi9Dk9ujcUos6vxg
Mt0n80SdFRrAW7lPZ/UqxifACaEIoXDdvKfqqxiJFv9EoM9+gN0MCS1BKkcMbI3AcBGimwGqUbUy
Oi3f9F6JhzhPs6U8qdWnPxeZsoubBRHw8bKqHQydx4K594JKC6xzOEwNAJkHB8p4BCF0mZsbEFzk
1omWosQMmWAq/CeikTOvkSw1dfNxQTnWkMLGHkzYyYOz8mTB/DZcTejnJ/34CImNw7tE06GAaeyp
e6lYYM3ee/4dRrjEPzkpIm2jZL+aG6SjgqjdOe4X/InzyJqY5o/7bEa4sUN0WVsvi9d/hWiuQsh+
L+YorGFV4swcp0h1dPp7xkqNR8Enhaq7PRRBV84vngZSy/Z5mBAVDF9T76Gz2KKMf0efUQGTTyeJ
lmdwDcAUmWyxpoETw5CoVQPIOtdOVYiY7dACWWee2Ai18zOI5S2EPEoZkjl9lSpTCEVl444JGSgy
SYDT431ZdFbdVk3b19D0PjKkU3pncekMunvbYjt7/jcyuVaa7Pp2dlXBxGrbyGNtoRJvmPyrXe6L
vNlZ4M8ddgezJM+KH47KwAIY5aJBb/E6A1h1E7KMOjLdl2SbscvrxWU2uXL8aYKzRP+7nMK41ke7
yTKpB2H6cECZz/0UO++bEEfYmO42U4d2e2waYT56MJhRkTK95HT0vqT1QfCJGFpLfdyKyKGMA8zC
9gbEYWiL4QHTGn16Pv8372LyhTbD3mb8aeLHAFE0FgeopCx8z3cPlLjY1P392ScOifJBcZ8Wwu0x
du6v6Jaw1o9Bzt1vUaKOQrYSqVg81jCPzReBG4hRbnMoUJtAypbgIeKjYpYj7C1zT20LLyvskxZR
6+mgeP09kChpSf0YttwYEDcWXriGhxCreGM/AvOqDx5BjehC8Zl/Pz5CGnitYQM1PbPmFN3PB3j/
9rD4eKKf7vgqS+PchnM7/dY9E9UaxYnExpLgTUJBrm9U5CCv0Cj6gXcjgCX8X7z47wQR8lcLo6hm
0aVhZxbHCNeS5460PihnazczspRPTtQOUqkLTmvu2ysyQv1pGPltvxJpp6F17lMj1MTy2FSGqNzj
+KinIX+g4k/DphmQXeRkPrQCe4f4jrEZF8LJyYzza4AuoiGlO87TcOBrYyDV1TKbFt75kDDLURAQ
LNOkDZzQrLcyx3DFmSc3UnY1QabApF0JMtRRgFZnW3WdezT3chu7rHimipFYW67t67PPWEoFVGoS
O3l/zBkxzIBWxLSESI1jicehhwgGhgvwyipLnitKmOicE9KOdzGO65wE9B/+aIjivFtp44Mv/0ed
XVZH2OEcQfu3VWLIZHSuMeGOaw1zLS5lGj9maS6K5bzGDf26ulzxOM3+Ab8sGqLvGXB2dyMcbj5Z
qhjyQigpw8AID8cpoHDvfwJyq2exFEnUfP6v3+jC0+yrF+nHbZFwVlR7VwUELzX/Z426Y0p6CpPP
Io0BI+5GuOxR9Fy3d7E+vPGXqMz/PfUTr79uE3aJEvMYhw6IhEZOrGQyAy8ThtmfJGcLdawoVh73
ZYZmVCpbxm6oSujKcyve3rYEKMnUFuOAYzhtQ/S+yYwjlfJdLBrsZ6urMGDCg0TeUERP3q2awdsh
Bbu+cHYj5gDN88qzLtpEYQ5vX6etwFglpxqpq8yUSY3scDesOvNjo4wvontaQmDdByd2Ok8i858D
1Rg7lEvi2fh6bmsGUyEequ5VBg2Pbt0TxrzZnH/palQIjzr0KTpuDfpxa4S8WY6vsntxC8o5F+RB
5GY8MPArLH88yrRzdR2caqFTRSwy94pU4PmtFhk/ifVVCrSs2jpg5Je8JmXLCX1otqPywWWwLPxm
e3tKQMGjVIa9NiHbrVKix9fqLkS0jQ7uk+HL443ns0y9/RcIO449krc+h3T/AKGDxyyVlGNJFtx+
O77G3Tf0sVRal4kpYaz/nCGsQVMqYZKjkBAlrFuUZxrHid+yY3fkbvuk7XwF3tsdLseqPTzcbWkY
vuJ/zhfAKfUW54EnzRpXdIairdTgL/XtXjbwbJHM1l1oguKQFWE3KYmFoxBNvTm7r1dS2of2Fk0V
oXaBMTwvJ9Kq4+8eDuEphXbLt9SWgZDlzrbuybapz/W+AWx5+60wIR2YjGq3YL+bTOTPf4eAc2e+
WXKjiWCw29fwO/JTgnZq3913JibqG2rj/NKESLI4L5HtNSii2FpS9ZKQo+vACE1qYSobt/8+i+xe
UTEPIjK41wyMb+sT7oUxdI7+6ne0c3nOyU1JiWKhrD6RztjfjDJyFgEPtXeFhI06IJuJ3q2H+101
TNymbTka+OtkWx1HBnXYRNpKJKQXzyn1MLJc2qS0WCw/mlLkCPJwoSJ/c7/TClRzSKiJGyfmIlf4
Rm5eRryTeG6ZNXOfNEj0n9Vobr2gMg4dEAgrTuZdfAw8PF9k41Uh2mqHesIbUx3m0ikKPkeUpYKk
GvXgcRHVKe6IY7y7uIBvKEHW5YukeglO3nUy/9R1g1poMr0zfEdNLSq/Y7Kc13dS8kKHXw7Y0+aR
kF3pJiBbE7QnmI2k0rKqtB6NiOqhpZaBMYccL/ijugQe8WqhV+WAVExtIx9xuQbnqKc9SLIktlb7
8AJbgiGX0sRwQSObrZ1ZljtVU2kGKXw4kYIwKR60zErnLIUBd6HDziqhl0yFASpK8CEX6IA2/pPr
xIfYMzTTbLyo6MG4Yj6TpBm3MDIyj79iED6p1eXf0YdtBuTj4rfAdlaaUap0IugABmFrGSGzH0+5
lT/5lmsQLTY0Gcqt+Hk7IJWE7zoFqtQX1MrXIsapYu5IzummoKPcSXHZwhe3r7dcX8Y8qxatLYU/
yY/ibcXjVauDMTjKz75yc8IOgtv4AW7XjkN9B25FRql5W1hUixrPtnuokOk1M7oYGSDrb8+P2Ev4
nYQxr6LZV8rBHcn1k/PEb1fLUX5j6IdR2L77aWx5sIlQFOiazkISo45Ga127fGo1f4ZpxNNN+Ocy
BYClqOgPIW01XQPQg5Tk/nwKHaliJ6ew6D06OqrGR/CqpHccsA+d/YDB+MRSN2f5nuJKsDMjyYqH
vdguxZcJHZAsk5KoztDoUCNY/sPaGAbXYUleV/wNi+XYSARepI0iukHkXPm4x0d6fzu5R8Uc8HVw
7s8D+IHl/kasQGKGr5LknbEBOXDvNHFo+yTqKowr2fsTO5QXDVw5W44Z4D0DIsu7AH1PbmTUXmyW
4FRa8ylIxJoMaMaSx7TbnZmCj2MfB99QlQipFvbsBqo5E6UQGMND2FB5DqY0kYzNsXxVa4xPW0vK
hDJA4Ck+/fBNzxutV+63zgaUgkB69crPpV2O/WIemjbOBtmQQExGsTQEbdtbYGF94CILyLfVAysD
3q7wJb7NnOT1nN8HFIh0Pb36jxCgvxpHBDhIbmQZXVxpKgpy8pd89G1OnCQgUx3vpTO+w/g2qUdg
ELyHjK8SLIvD3mwoeNYM/C4ohEKTxidIyAw+VKQ98gyD6nPKFzVHfqNub+qfwjr0b6cBL2d1XDDa
30SS4DEWULkUJGr27txmOJFyCQvl01uqXjCRSv/jXL9/nY2eiZzv5/ciq669KXRWgdGlJgavgu4k
/hyTRNXaFteqnFP6YTOPuaykumVqtV/abfy8M94QcoGqcrU8afK5ec6YjwiXY9uNggRiSA3aEVy/
UwX9z++Cb0g9pIjDHLmxaFpaZgBo4fZiRBUgiF44rqsXP10YVlNyTg17WP2sDxuaKjlITrqStzNb
LrPmIHFtiZfTJIPDuoWqEuKeZDhaPMzUiF59QX8E9IoNkbt0+nixiViUG5CiogFlajrnEUKrR23Y
KW9GRRMQAtefUtlEGzeZWqTo/oGl29X8z6pjO9QDUA2SKfwxaGMGERAbMpn5Y9UUFHgN7A+iHzoL
fPfulPDT6RplhSK9Axn8PokFY1eYLzQW+XEPx0vBsUz/R0Lh/48U+DM7V9rqCpVWe6vdPkGvP4RL
JcFM/PDpR5vp5OeTtu0JeBoQ1r+NkHgDRYaSMS+tcZ+NJM1nAWe0T3SlVQB2aD8/iBu/blfqjjRk
RchnRnqk5Ft7yS7pdqW7Qbv39+tvtv0bInf1zLCVm05X4Ok/ePi7JytjbUfdKKxqIs7gRwf93D8K
98I+EmR6bV+HtvbCEc5+ciqao0z22Uudt49QfgCWM6C8uLpfGEjSUQH7ypeinmGj+tg5Z4HM5Udo
QLaHj+YMnnRuF1gukrqR0xKogOdSzjsmsfUy4nmJTEtIJzr6Fln/5yJSbUphcyhHZr5q+uJ3+oxL
gcggM/Ig83M/eodFXGiZk4geUedBQntOdZIm3ILEb2cjOi/F4SECBqxrnJ7klMr8TM2586QEGkWq
do3PpvB/py7ch/E3v7G1xpOTNB+R/EobRYGDec1Inkma3+LJjKA5g4VM58fvRL0v00MbYqNTu86Y
kgDbqPBDP4L7PzYRtMmuFlpUzmETCzsu+wBb5auAuT9VPx6GK+TPhE0oyWJ82OlIghcQzgsfQeEl
JuQUA1npt6CMslAtfBBYKRodMd9Us+g3StJMIWw3E535Sd8xDpNOapiGJ5GQ+a0bfUGkBIgTejO8
Zd84GtBJOTCn8wNduCZGWVSzcCHXv9Taii1vJHc1b40+CA3b5T3wMy5uxyS2JgSs+Dt2snQoyInX
TjtzF6Ds2/JmIyMAK+a1OpRWiCSBBFUTv5YKQMUJxfdZ3v4U7a9g67RZsxYh+c4CUpWY1k3zWlNI
uPo26qTvH/xksn3TEwUswZKZsvHURslJTwKCyEujGaJ1/vW385Oy4/laCNXiMbZ9QAJt/xys3HWO
EwkeCrS56RGgb8+Hwp53bhz74p+jAnY5bhSy+Dz+i21zjrQNjiFBd7ya+V6D7NTRi7ojPcOM6u1N
V03ptqwEDlQAAu7wg4t+dltXlHz140wQOay/FrnB6rokdrylzFUZIuD6R+PzTmC1iGC5A2p5zJqF
yE5Rk1EDhx/saP9gDUjYvuOOE+E1uGzKmeTcXaBc3nBWUV/jfww1vxBuREdL4zyuTyMO0j+Te1du
X6Du+8JDHwtaBrMVAkZtzl/L+UsKf+BEYPijaruIZBDq6z/FfoiSkL0m01dCPUZgiXJ7LUSEKqdY
0xyUBXS0MOMf7rwU2BgyGd9Uq0Sv8SiCG3gvbu12GlFAefM2KL+brq8zTe34H783a1xZpUfq5sys
4AzQBoUQehflv4BnXQjkk8GoeCrp45hk/63KuStfqltVThaGpsNLNyAeez2S2p0yLL+30wEmDopf
eI+nsKwuYQkGgMwUP5jIF5c9jfEWOfNvtFbLjqp5lsLffgX3C+gzbAKQByx84o5oRHofDOkUOny3
7J7+ttwEWFcjHcCr4xCx/jVOOsZqwOHk/UiOBpTP29ZtS+GylueLsVgr0+exY3Ns9Gq1XPnTuTMe
PnFOlzbD0diMPwSkCwT6JhJfO6TPlab2vsV6ePC1Bn8gJLFnip8RQU7ifM5TMpeSpFO5Rqj4IAx2
6IHdRAoDMPRwldIfRnJQPiqTfNF1bp+wILoggb00heEc9652hrPHD+HDkM97eECbLDoEkEnUJfts
wSV5blnGXM5UougF55b1dh+4ZfHPeXk/NpDJdqLt22ALEAS157/p84Jy9Epi2YXm6NnKyIDUtSx+
vcWcz6CLxiiv5TNm62Jw4WOcAaMjhaLVz+wvaKTxMDMruIvYfjlcA9+f6WVkS61YxnaYMNXEos6e
YRba8qIJm0BWrTu2hIe4f//BIQEffC8qD7ht/Qsi+x7BYkbOgU1wWEJiK4YRnixRZ4fIe6uMtYxj
WTzC72BgR9RE0QPvx1vyl4bmo6pUlrcJhsUd5Hj8NnX9j30jtp585lIBjcJzUFwEoVyrfIcxX2xo
OuAkbeCUK75EyWGwIMIFp37CU/WS8ooYrwaFBXYRlJGJMamfpeBJy8gzxMK4+4BJacs2qCfWl9Io
PQR3gAVdaFBYe88eNchkIna+HWICU9lclAREiarlM53il5mkHHRwDGo86HaLvEt+akqzqMYZF+15
p5pRIoLiU0WufhW7silv6NCwC5uY+E0fJ8KnBP0Dl134aZsj2w5mn2SjSdtx4S7fZR5B7W+AgV3Y
06Mxk9pm8roqZIxPm1O28B1g2pmeIcnSQg2HZx6GpwTii8t5CQ3z9CacBlQ58HdwU44gOmDQKmWZ
2qHN2mtfg9OmE6iqCBy4a/Tg5qXV30iF8XOTU/nB62SBBQWXEV4QojJf6YDKypT9dlvF2My+J3fG
qQQEz0UbWJF5lYehC7VQ43psCr49lCB+sPKk4JFOwg5qner9Sikc1sanKZG81XDkotyhyo0npLjo
iBHM0FlOKjt0R6ojZY4wVCh+9kcYjefqLi5tD1oXNlo0HnjwUNi+Jxu81xlezGNRCpKGwroS9iwu
ZjFjIX++bFiFrSc44ZMfBdjwy5ebjsmRK8JRGXg96yPZHIvxpQPkjzvX3nxTlI8KUz5e/cc4ADUE
vsI661/HDmEVTUr1n1IDxnRgu1DaTSGLwOQpg0adqeOnODFlWVgn6H+BNa+5TPBkgWf41FvWlncx
r8OPMrVUTlo5qC5udv6HzhTfqxuFSLv/C084rbrtKvBKZDHVcFPH3PhLQznvR1pas/TXYnS/JCZC
wfiVVGw1LkQ4rIXgAE7dgkPoyCTYbahF4ujFdrWj9cgjoMHxf0ZNX4Bx5mKbXu87+wW9EPi1aENX
O4U9i/cCoFpOACTLpZbvad6noBtoPDRL5ICXDtXWiQxDN59xgibBbm2KfPCzWbA8I8JMlVMCrttp
/XYHh1pJzz6NldtS84hb/A+RWZpUN8nRrOaKoBwTpRRz9Iu2HIdcL+enYMn5UUCRd6+HhmqPYWHM
3TQ+nORLMs1nc4c7BY6WnRnrvvAQekw9EmaDxieNzntYRJXW/Lw4g+EHJunPUzMjHCIHeNqvVEhs
gcdVjvtzK4EV36dcOZ8Lo7WVj6soONK7NMmT7d3VN3Cke2v4FgKYWT+dzAvjFOXAjRYcQRAySdPl
K74ipEghXpTkj8mMACL6AgJQxZDiFUTobWhus3KbHwwDeZe+avhueSdoB5lz8YaJKfCayPnkRwLu
/468XuFTzAmveYXocc9hhTvFFhSQjcVc7ZJkY6JY6nMYUZQtExn0KLY0JUo8gR3ZXlQ8FXSDYrep
0s8V1xNUVkB4vVMlhmH+A5q3+4YX3YHkJbz0iZMMr4G+p7dCvmfiVJ71efHlfh4eMLoia9dUNfj4
Pi7yf8I9K3aFifHlZeftpRWE9V4G4T3iTXeE5Y2u/cwcmfdiTJH8WmxAQNB+vmttomXd5TJsU6s/
/Cvj1nR8K5gu/UOj4280Tq6MNX08DVuab0r1Bb1WP/R+DAsYxFOz3O00Awkrd//uuF5CNNI8/SoG
eiZcI2Orygt13Ru2QcOMhkrrphv0KKecsoTcjS6mhh458SXt7e0Ck05Q+tWxjjDs4eeCiaJTKgSn
un9FOI73Ci6HfUNA63tYOL0NB9SLAEJ4VKeGpue0Pdog9cLgUvs12MQi4Wtxogspe9Iwuq3UX2fG
kYeWtCjvQDz1gNT+L33p7C9ObAkyxWiFsPvbAULX9B8CVxc8qzC/OvxVZE4iYkEcxcrujYQBy/O+
yuQnAop+gc9KN4irxa304Um61mdB1te0850pgnL/rGItFy0GKJx4Urj4gnWEvQNBS8/18WS+yc1V
osWn3bgQM6R4Zz5A/PJrgpFpOurpHWUP5kh6dZ2MIVaJ7ofG6ZoKvJJsMeduZ+3KMtrRGuttQbUx
cl4vjWMOTAXAOU1mhNmeCLIS8IEq3QXDY2X0ACL2KAR51SZeqel72mSwNEC6NSKilwSiYPWTsoAt
7RAPHQbbsiDwi2vuiygZNUHKU3WhRg8QD+fYDv/6fnoCp4+9+xSy/6pc+l47DhOQfKP22zn25a6W
+G36Qgq/6LRsaO6LopH1CbLcmXddrStRnmD0A39ufNq46G6x3Zkf2up84HvlxoPj3k9Y6SxaL5oa
vpjCvaK/VmVZftPz9Gc+yrcQIOu6rwPX257xmix1Buvk2YX/hFR7+KOh/ooJ+t0+kFcghJIWdaUZ
/cIH/RsE25YeKofnLEbKzZKR23dhynC+9oVecS+Zqesm+jbhv47s3cFEmci1SCXlOVIaoke8aG2i
dtdBnofqO3iwp+5iUyu43lMEZQ1BapYccvsWZhaoVVNncxwnS5FawzGLJLoY0D9CMfzvVoogXpkE
7PpVZ+WnYsI2l61SEIdxJ+/2vQjI42lysCDnhVAN3tHf1uUrjBEpzrFMRfXV+/WEe93W/bcXfJ4C
H61ag3RudDNvk3imjom3dAsUSvd6IrFsVpVgdkhJpN+F25SvR+6YJ3/RHjIBLq6O/furoV8RwewM
VbSnpeCyxGitDKKpOWcVyDEHCNmOCHf18VMUq8GWlrLQYv12ReDLkpo45GAZGO4CDPTiPDBkl/sZ
k4SyFpZhQiyuODiGMb+QRlKc97VuyIXGnNlhkABEF1GWjo+1q9s5vgGMOOKH7arFrNEvRCnWstwJ
cNkpTzKSJ1Nb2FlLz9MwP+oLKqB3ePezCPDwHupvjVBgqGBm/N1pHWSKaHZO/DoGWASF/lFWKzgY
RosIw6Io3ZFQz2koYm6FzExM9sM9ueaby0x5STVJeUXKsAFe/M5SZa7NovvPkqoYyyhCyDgXQUos
wEVq8+xzqj/EvyY7KsgjZeaCxUsTUdUe7MKD6iyunv1ZXOlKetRi+mR4flf5hCYxqMYJ3XSmmels
KXbDIo3rx9/3aCC4Q9JGHSToe6OP7MPMnq4kVwJCLLMvyU1bHRpfAK/0bEL25ZeM3Z1ppc6PxgFn
K3Cop2JEjTuvL2W0PyaeQm+y9oFlps7nVNhLh4nQceQms4pLsbUolHTKBgvr0IoONGR7uYoCClpn
N9gpyBNh7NAvz3S5Wsn/mfQAg5BZcQ9bxNmqtZgS7JljP7X9QflTvH7xBPM5tJST/HzeL1117Buf
27SeprnEgOK+NEtZSwS2yuoSangPqWo66Ks5FMjHVq3F7Wrd5btJhM+o+IAMBQ+Na8SAvi1NSN1w
nfkK+MA9OSRySjHb7tN5+XWxC6+OEb1wzjcKF5qkVe7XGHC0jAqbQ2vBPsJyInsKdHB+Xx4NcUqA
8Xn3nRYYM6Zh8f600DLMCbdNqScZKIxHUBjpEk8Ex4wXDqk755g9N9JlWA5Kz3/rUeBvYiW2DlkU
GWzp2X1S0oM79JlLB4Ei34CY0xQTVr9d/uGhT0Oa0J3/ZhTQcdngzrVSuwSdq2cqUHh05Lbfww0+
1uEelV3y/fO7g9z/8EZ1kOW4HZpLllWLBRhjqtzuN6x0lhtbvJTJe9nfwnvu62EltaBv9r7IQt9n
pN5SNuf8eznIdCAyV/yfSjMeCmqYatLepcHoeAyG7rUkS/CqlQT+R3RYjcst2yk2lTVorvnuZ9Og
BiSLW00qw6pXUK32Q5msLP0mRwpEdr88wn8m9NdudawTtAxvI8E3onV2cxUe1M6i47myQdk6lW9b
XBH7dcqOkRAhBDJ1Pz9Zrhuzx//gvkhl8B3eHv/j12JCA0YeHJ8z8bGZsqyjV/JP7aC+wOuCIuBA
nMJybVJd7Cr+6CFCEOWpkxFhxKdcNRxr18HIPtd5VW1Z1/nHnq4heL7LyzpD0c5KZTr8iLVf+JCH
RxMMqd1iKh7SWHOuNv3O7oAEvikT/DYlQykdmRAH1BBQxYQmFHz5pODjpu3hwutzVKOnv1gP56pL
SXoAenl5o+TtOC64XnpFSjhGaNJYqBx355Y1AUvJEDLoXku2pjN+a/UaNbv1gX/Xojqwbo4FtOAR
G02VNUU1xP2bEtmHw3sy8HOVvgvjGT4/HDJbvQTCpoyX3akUuecdDq65uXEW+vMHpPRnhllJkNO9
95cXjgpNr/nxLTW8JxhkiFCYEm+B64mrSxrfD7QO6Wak6JZezavbu+MWqC8zOhy5MSW/hnl64XJL
Ut+00cg5L+8FHF3ahSQR/scFuw8RQmgO/3nf287kEgKgPwnLGD65hOLIb7rDUtN61CoBDhQzLJXV
jfLNoDnwWUSU0PTy/sARDNXZlquRMR4FKmFw5E//QRM/bCjPi5LS8GbuOLj4F4YLgvW/6AvesRvU
RdZx4OQTs4jL6rXRAsC2n8+TYotMNZT6lzxQ4r8J2NoUS64+sn5RpHDuZYMmtxdyopcmUIy/HW23
im60D+byiJ9poDe1jaL7BOgd0FaYZlhvxmJoZeAgUeQPBGYUnO4jqc4smfVFXD/SsP4E5FYgAOIa
fSlkRk8uMliIbNNKDlUp0Vz7iklvdGinVXPcUp9vlFnnooA6cbHlniB9TbFEA7jFVE1PydzUZQg1
JaSwCwgJSOR3pJXyOHXhLa5TznJj46evWDNn0EeBaIDtBsB/BhTq9kwRNCRvtgR/EzaeM0nCpz4l
k8gZzo2Sy/lRBWmIxL9Wh8Wv2FmrLTrLfmgV3KGg2GW0EfGM0m6/a1xnYkpTRGm91NK+Mx6k3z5l
Z2GQzUUTgwKqJPfUp6W2qfZukSCfeCGosRSCmvTIVtx10MNlJD3wjd+KtHKqaqjXSRGSiFa31DBx
XpRTwMHZCPFCC9BtlQEl2WLP/G6rA8YxE43LN/SEYugcveiMEBMsn4og5Fxe/INuf2kTf0CEvACu
cJ6zFAFXQEPXfBA+AApl9ut0FC5vKCN3NOie7NyC/oIuIi2EFvRLqQJ7qWrWte8NbpAVSjVngzdB
/jRqDgXyCWg4gj3nS44B10uzUs8DCJAt4xfOgmQbHWJqnJDG8Kv8Mt7VMU9V1GmDxAdG1kYi1jCc
z2XXXJoXYpSicFaorU84tOBZL9iImzevcbTohSzHUJkCM3yFWqSFd6f/wG3/sxYACL2krPg1wnd9
bkVS0YChX3ONb2Egxii18Cv0GO/dzYJMvRLwERMuPzbNHq6soxOwS/7/oXvJMjQvFDc+X8jHrp1N
2EBnY2kWHAiw2eSOs9egmRoOjJIHCQucCZ2BHJXYVj85gT6E9Ri6LS012pJB9ecNCUsdVPyZNJt+
DceTL5MBi5QUjYceugN4DUquJQjLu8UkZo89KfNR9OJ4YmiSMg3P76ejuyXQMQa/cWZ4Jzr384Gg
XKj0o7s2vxyYC3nQrUjEO9nURtrdXjfNFWN45FV7sucMv0aLD+WK2NywCCSt/R+gFSNdXyv4Mgnd
vSy7Mbs4HjE+H4PB6BeAFSdfcb5UkBcRuVoyudF2Pgd3EpNUntJTT1imKJyqQL34sUBTcUyByXKY
XplDlP3yD1pfXz72faeYTnLkLD+1mRoOJFJ9bbbjUrBFSENTxLjldulOpARoPXf1OAmN5kDv3opP
K+fJ8DxSfzwd7VEKkTdLBXj9CwdGbd3q7M36M6to2m3vFTDg1JH9t4etnCpT5s2Rt3KXFhHH+gR2
ixFwAD9b4MIM234Ce8VqMlwM/xUaUK/+l/E/WzgJbZuK9sLCkl/ULu99dZhkrxfQ03ewANDBl7WK
u+zXsnekMYonTcvZGx85tzccsBKxpphG1017s2hJOEzz49crGwCMBG7y3AU2ioTgHzCzrMP+tDqe
6iWGNFItUhEg6Y1+ti2Ajk2DsUXQheLYX9cnaEKIHT89x/GKS774e9c8bdMVhUy1fEmOsj7UOhf2
sBLPkrBR8cPchLDJvOE/rnPNQzO0fjjuKk/YGUgGffaf6we8OOQF19SCfZIG9+kzNQVnN58PRZ9d
2AwUudgjQBVcE5H/29uc4XoLnZB8oLW8BLzdd0ES7EuRwsBBoCnpktExPXnSUfYgGP020F3rKbIH
vdF3rc4PAP7F+n9fTqGaa4L6gkMtXbZ4iOYF8HZI6MaO8PTMrZeqjDY4T3QBHXBFOsmV2iQLn/4G
8KqXE0oslE8egSFbWcJe3/eOIg/mFJ3TLZnDbY0RZDiXwrcIzmEKh1LdN2WLFTVzD1RajS5PKG9L
Av7yw5hOb1tpYewsYI+ncqALc4E8RcAujnsvnE84EI1paDICjXxmecySWQczTeNBc+XORS2guHse
layD5lsoNhk3o+gEzOg68ssq4Ee24OD4X04y0G3I2c18SAXW+PYLsLSjcB0xAc2WmBoZ0eXAmS8W
QCClNx4o3FnQCruFKIF9XZsTp1kIg05d3QkOfevTkRePbel3VdBHg5RE8fI6tnn9u+dSY9rLmeFB
BatHUYoH9dnzlPPWxlcmpIuouVcHDmRoxu0acre2TsNwXvQnqXdpGsDjr44CIEiAcHdm6oEcFacU
NcwJ/Iw/mD1bFVL8TOO5n/3onE9CYK8wh8JYuAjFE7RzMQgG94dyuy00c5AT1FvOE6CV/KIu8U4j
MyhEXlaVKf7Z4K80kGz8D7iQcstXV9E7jm3UjZi3Oo2tA+ez9gk+ygCUWBYyebJ1XqvTs+ujaP6o
SPnjwNfKaKb/Bi38tlK2Ra6w3jBPvYl8Op8CiN7bPgnCt0N8c0fX8IQGBzhfTVBVNMEEFra0OK+Y
zP3BmKFi/QdIaNmAxIkAruahdvA0Jovb/lLhMJf8VzMai8S2w+55HfLTPMxldktz78QF11OtHvqf
G6NjlMdLw8lf5cBd7zYMlQJ9PSrIEWGYcPDTfqzWvQSg0XM0TAuoxg2Gsc08WHzOi1fYuSq6cZ9m
wbJk2umaB1Bmf0EoyjU4g+q2cisJUiNGOcQOLM+zR5QHqTjoBB+ZPdU41OUtlgTZpN0FQf8uhTCI
lQBojagBVwjj85c6pTZX9hdZNgGpYR4dVdrReM/ad/hB11+Y7gILYx92FNnc8tsrcF2PYs/ZM66a
KgK6yPAZKgNply1S1sUtmZN5RHser5AkPFVy8rmQ++RU5juJH8ETlzLMTOOelEngybv2Db4Wx4Kq
iWyUVNePZuIxvbiGOeKE4Hn2K5iqGN1QdSVVWZ74ZKjbUOG33QE5AmCVX3RrmFUDwbW1o6BPbv4O
dO2V2YoMes4JF7IPMaIkrAu48GMWVUJgVWv5eY3rcHs=
`protect end_protected
