XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Un��H)�!R%�>�^b�{?��U��
�[�[��v6���_eJ�\��'z������#:��1��D'G����/R�xjI�����oC�/��M�m�͍��a5��2,���[|�2��2��۫���g&����=���g�mY���`jǺW��j9��(*:91��Q�/�<-��o��Ճ��;�؂�>������Foꩴ�C,�I
GMc�\������|��vp��b�*�8)�O�O�0��.�J�]�eQ��ۙ. f�l�xX�m�9*}�e>w�[�=s`�=�Kޒ�t�M���)�!m��`KK��#���j?�2����Vj�s�'$rc��*�Cnz6X�{��{�� G��]�^ul>�i�^d�;�F�.���a��̃����:%p-�[
��vd��d�O�z���{��4�k�;P�ʃyN�eݪ��.��m��I6��+��7��b��5�]\�3w[�ʵ�8�u����/�$4��[�L2�>Ñ<������jF�]�}t�v7�5dy 0�u�0�_<5�щڭ�0�{X�z:'�N�c.ET�+��櫺�v�g
X{�Kb"�v�1`�%A��[�:>�_Zg1���V=]'XfW/R��a��LS�����s߯4�S�����K��|��)�bg>g9���K��X7���t5i�p7_�e�\�C�~�Ŵ|,xJ�xC����8�j��Q����]o�te�X�y���tK/	]���֩WwF�mj�H;��B)p:�ӻ��ԛ��)���S��XlxVHYEB     400     1d0�G���������=0y�?��g�ت�5����	�����Q�� n\�v:�\=�G"n�i}��$-��9f�	]�ГU�Wz*�$?J-��D�j�@g�����D6��U���u(|Z�S�ꗂ���mCka�1nda�>�^�����S��5s�e��(,Rڏ�L;�e憫n��I�4xl����D�ҏE���oBA� �u���7s,�5��?�F��#˧��f��G�\Z�dK�J#����p�w\���/�(�A�{�\0��-*뀵��	崹0��s��5r*��Ry�T��ƱK�䛂��u��Ŭq�R��,������j�8�X������T\%��U�����T�֋=�:N�>qY�ί�%4Z�S����~���Bc��i�5t��98b�,5���ܢ鬜+��AuJ#�P\�R�[vQK�Y�p�"�����|���t/j��.���~�O�XlxVHYEB     400     110���c�X�A� �c�6j]��v����������AA�����Z�ެꀖ������G$oϔ��C���ʱ�ŏT�ӗ�w���'��a���Z��c&�G�f-$� �4|q$��X����;aXc�t�vx�Z�̕f�K5�Ź�G�Q~�c�b��h�):��~ȳ��.��G%�E?u�&���Z �y<w�l��>��hg췰&	��|�����L��F�lm�'5����%���Z	Rϻ5����u,�ȗ�k&D�K�XlxVHYEB     400      f0JuU�ۥ�?¢�W)��4��D��":xS���QEGQ�P��rF|��=��`�ssV/��ɾw���M�e�hu�h��G��ʒ�i�Va���s������LQ��Ѽ��t#�_��|�E��1��P(��=8W[p.���eHr n�6s$���ûHźw��P��|
i���
v�	`�uj�@��"��#�9�hA�S�z� ��wUzC����ҡ8/��
W����}D�I����qw97p�XlxVHYEB     400      b0�/ǅ.��[��x�X=�h��'ҏ?PT��\���[�g�A�m~g�@%�1v��o��[�f2���*�.X��SU{i7���3E����Rq���Д�NL'y%�?p.�)��k���Q��.�	��9do'iB5]�����YA��e^io�����Nj�	h#�� ajXlxVHYEB     400      d0�X��m�N>(�(̴�Y�2�e{^���`����I�O#�u�s�����F���G����xʨ����r {F���]���E�&;�
'l'� ҧ���  �-bR�l���q���R!��ٳ�n�l�� �O�J�<�^�K��e���O�'����e��:�bY��2��?�~W�ߐs�F�4#�ڨ.�&Rxh]Rs6׵�~1�q\�?�XlxVHYEB     400      d0��b����-���O��2Ε\P7(���,���[�\�5��#W�W/�0l�ǬD�V䱭3�|��*egR��L]��v��=�.�+9-�#N�D��nQ�Kd�@��N�D�+��7
)���Yd��Ў�aBe	�����5d���KMa�D]�N�xg߽�Y;�t�UZiBuk��so��U���ȑ<�� e,9���GuO�����m�z?D��U�XlxVHYEB     400     120�UB1*i]zα6���9����݅p8� �������7r�p���_׼`E?f�+�|ċ�j3i������C	���'[B���M��!
#����7R�=c7��`�[{k�L�[��R��c1jS�B�P��vD�~6�q�G��Ϧ�Xcȭ62��K������gX/̚�V��(ɏ�h`N�>��}]������j�!l��(j���96\睃]��]o�E�N�H"D��!VT���c�J�e<u�S:���-�M�g�S�O�!�'�,g�]6�M7�E3fFL�=�a��D`XlxVHYEB     400      b0��|��q����Z��#J�A�I2�E���i1�`��#mp~�|���Io-`�%K[JN���f� %��䒛����=�O�Å����)(	�p��g��:t��4�ͼ9T.>*xd
�[ �<���;-r�u���\$�BSo�R�\�߳3-��4K���^qB��z�߬�#�XlxVHYEB     400      a0LJ�kVふ�k!��a2�mڧ'p����q2P�t�r�>��B���:3� V4Qj�2-G+�+ݺ.~��rec�>�,�w��1��/nl$� ���:+����n�ho|���t� �}͂V�^`��/�[�b�ݒ}��٨��3�C�i�M:��n�+F�XlxVHYEB     400      d0���!�/��"){$!b ��B��R4R��mvu�dMx
��c��s0�nW�E(��HS/$t��$aڂ������+�ɔI�T�m��o�����Ǿ��:�_��r�6��ѧUB+?z@f�l�{5(���d��煃�Gc��X���t,��m+[ޅ�bAA��}
q	��0��Ǒz���&��Y�wv*���>:���R�бy ���� �XlxVHYEB     400     180D��lloI3�w�e����)��p�wU[������Ri*O�Nb 
F7�@풴1ޖ��VY"t'��liX�Uy�Bu�Z�D�����9�'�C,�~S��z�qӆbs�G��u���e����ʠ�h���+�4;�`$3Z���Ȋ˫��]�XՍ﷼��c��Yc��������#��^���/�yl)S�1^�~dqhݬʰ���Zq>j��b#W3��	C�ަ)���v�qQj�;���~Yuʺ�&\Z�kI, k�\�{�K�~A�'�x\Lض�����$���i�����8Co���}�S�`�Au�,��6�S��3}z��+ڐ�C�f,v�E`�S]�/�]��T�F<m���KR�t�g�[�{�'�XlxVHYEB     400     130�����Ţ�AY�!��8��,(�Fu-V|E.���?�WG�>��l�ڛ�Ũub>�G3'��ɼ��u|�D%�F��Ĺ���!���\ ��; �~0�.��y������EF�ìY�*J�7�t��C~��6�WQ�\�LmHƍ��uY����({��M�z6��fj�Db���܃^_Ckeb^6��%-�">Rp~�[��׵��[�$~	��F�Ǩ���,WR�]�Խ���1��}��}z�޻C�wzJ�G�b���&��1�f3ȱCdf7���V�#Wږ�\1ե������h��n8��XlxVHYEB     400     110���ɥ�w0q�(͝u�(v'LF�Z\״�
\Nw
����E�|�z�G7t|��A^��S��85�4��7���3��F�hI��` La��~�|:ԁ��ā��$U0D>��(�&A�!e�Jo&�P�<	a)L���e6B��x�fu��]�^�cʺ�Y�����M��߱4��+#��&�G
*��OX_:L�N����J�������K|�u@�]���W�t�H����p�c�� >���g޼�쑣$�ȪO{.���M}7;$.q�uwpXlxVHYEB     400     190����[�/�K@О��9�[MDC@o�����|�����ƫ����CP�ldϜ\�	�<(�v�x�[��~ܥ�
�k���4 �b�2�0�9��?^��s-ғ��Pɂ��*�\��E{k!M�L�W1�S;�p���K��u8_D����!̟e������鮭�og;x���I�ވ(cHt-֍&g�+>:9�v��..�͌��e�f�g�z��f4�7���#�s�L����+���XvrC�Qr�����Ѯ�; ^.�A�ռgx���ڵ����ӝ�2�?�=��9��N����#w>�{޲�Ѹ㋤��HF}��yp�D/�[�9
��pz�W���ҭ �� �`[4����#�eo����m��A�s��q~�و��B�A�=��XlxVHYEB     400     110��dl�{Y���e/ؐO��~eU@�6G�qg��9Q|�Qb=��Өy��D��:	���qY�1g?2tS���A��V�<������ɸ��)�������U��Ǘ�::Jf��LlD� ���2x�Ka\!�~	3��7t�ķ�W����"�%�gX�v��)�㼫�������iaZ�y�e��^lK��F�?b�0�~o����{�f��ϫ~��I��2���Q4��;�����ZՈ���e��,�&*����ks�XlxVHYEB     400     110�9q�n#�����>��cD9�B��L�Jfhu~�O��96n'Bj�aY:���`*����y�3���@\!H!�Kѧ�Â���_�����I�Ĵ�P��7�?6J�ߎ�7��lZö9[�/�_o��f��l�s���=��'�%�^�X�w���G/6�X�����,�à�jA���Zz	��}�&p�������l�Vv��s�$��t%�RX#byGxPm����2�>'�c�O��f�	�?Qwu.!����/�qL>�O1��XlxVHYEB     400     110]޼�W�����}(ey�G=�<`b`�8}7i�A�t���<f�0�i�ɮk�
S��'g�B�Q ���	��Iv��)�1�Ѭ�}��-L��P��n�������</+�������o��Uz�t����sHޢ�pBts,���#yy�W���
�I׌���%����aX�[<[)r ⠐C�*�IM3p2����p�����J=!x��hti��U��P�:�$xx�9�K�(�� ���]Y9�Jk^$�����]C~d��XlxVHYEB     400     100݆�w�`�K��I���c���bg��J>��m�҃�]�؇H��1�G���1*�h����s�'K1�,`r_dv�P�)�	��gBrܪ��.�3�/ID���I��$�wy� �tU�*z.�-�
<0Y8�.0睔d2�[љ�)�9iV�ւ>�J|?�ꂄ����'L*kïwC�7�UbBwߨs}3j'������n#"D^���M� �F��q������AP|��tj�U0I6޶�d�?�X��l���XlxVHYEB     400      d0j� 0�=�@��Tg%+{~���  ���Ԃ�����FL�&�<F�������b�GݱN�M��}s�S��{�܅�R���jZ��Q�{-�/�+�a�UȲ�l��aS�$',�Qcu��[:VKw&t�"J�����.��v�M��,&�O������a�ʢsY�[�v�"�B��!g������K�4+���zg�P
������EtXlxVHYEB     400      d0���C�>�۬ŘE c�s��5Ź!pd����9&.�n�BI�M�D�{p����/qR3fL���Y/ڽtc��HN�@�M�md�F�C�`7XU̧���pf+���PE�����x���p*��і>ȃ�N���v�jz�䩎�\{�-j�jU�2j�u7%L�l�@mB�?�_��d�>��4�eY�,�a)��Y��XlxVHYEB     400      f0hԨ'ܓ�"ȍ*�oWn	.�@f����O�e�QQ�Y��<�Ć��]ґX��[��i��>�?}7Ϥ����d���A�} "q�)F�͜W9~�-�j5��{K���SF%����OF
�K�@3�'!�.�݉��Y����j|��l��A_�ͩ�!��p�Y�c�҈g��]ѕ�q���<N�>\Gi�:�z��/�$��V�����e�tY�a���Y��Ц�.��7yh7>�XlxVHYEB     400     160�_Hf�A*)�3	�F���R���v��Y#��E�/�V�[J*�#hi�:�A7]���	#����N�k$g	�!��\J�v�s+	�])bkO�3��Ϲ#��=�-��nr�E>��O"{�O|l��?U���f��P�� ���!�f�u�^�Cߵ�������|A'V���^:��Hxw�$����~D����3�C�^�D���z�����>tWr^1]ߦL�`Y�'�%�P�P]\WB�5�V(��;�kH̒�����x����s������s��G7��������Lt�9�e�*�3�;o}Y�_R,�I�A��wX-bY�h�!�p�I����!��[�l�IU��5XlxVHYEB     400     150|3��l�J\�*�8O(�Gq��a�p�R�,go�HW�k�-4���v�]օ��qK�p|=]�Q�Y�GKi,pK�	��T�a�����H��ӿ7�+d.��0L�&�W��Wj73s��'��b��uՓ�Ku�r��2hrAL�Y�3Ƽ���n82�0��]���9��4lD<�/\|@@P�(�5�'�q���K�S���+�"���5��DQ�*N�$\�օ�|�6��Fid7A�+�x(t�ͫ3D����E�!dc�K���
�SZ���DvY�!�ږ?�:�&��gG�o�8��+�[���'�Z�U:�n�=�4��m�G��@|�XlxVHYEB     400     100���d�g4��v��`FEw�S�2j���ivр�V�&��dT��}�Q�W��:�k�)A��g�L�����.Kt�����!_/��:��K�Z�F��*��%���|`'|������#����-ׄ���k��z�����KP���GLX�z��a���O{���/�@�l�w���f+��m�5�L����a��m�l�*�=̪fٺ>��'	b������K�i�8C+�>i��"��Ҝ����]U�8���XlxVHYEB     400     140ne�i,���-���z��1�rS��*:���P�_�Q�6��)�0�5�¼h%��eOej���,�]��rب�m�6���J.�ZF�#�i�$D��Ͷ��^�Ӡ��OR������և.��W-.���~�D..�=g����
e8&ơO}�S�בw�IvIƘ�a�^��i��1v�񢂋z�:��T�D�?  �͵�;v2觀P�..W<��GN5� �D����m̱:�0}=����7L,�?<3�����ی~i2V$�]��*+�=Դ����� Hu���M4��fPj�%0W�lؘ�Mkx~�$N�d���*��u�їhXlxVHYEB     400     140�ݔ�9|+|���S=ϐeo[���]m�n���?��p�a�E��؋���#���ſ�W�'�NB#��������P�,�H`�V�݇5�]���c��H�#�Z��f��3���RI�>a�n����)�f`�8�B��4���d��]Z](&�3��{4�炍�m[1��8t1I#5L4"��K���=˸����u�[�?K��������R���&�6+�O��������(�y�3�&Dǡ��֝p�m��_����'��{��	QvxO�����MXۤ@f]}͊��]�$i��O:�PW��Ҟ��XlxVHYEB     400     130�G5��aD���&���J�H�Zw:���o�%����·1J9x������s�t�%݋�S�8c��D���*?���1�$ͩ�_n�����>�W)m�KF���5�ʷ
��@�l2%qV��k�2K�
�e�����@.K�;��{nS_+�^ ����2w懭ݤ�_�!�՟W|y89�:�Į)���V>O8�H�l�sg���N+�s���JF�~P�����01ئ��k�׎�Dd�/����JEi�������?�@\|�������m��,��"P�l(��hXlxVHYEB     400     120�s��*�.(��4�k�F-Isp&\�ת�O��/3rA;6[A�O����l��pC-'�o>	T��݋.���Y)ay�� `��؉kY0��i)q倓_m����>b8�ԧb���~3"�=;�"߲`����q�{E��S���a�����-\���Ҝ�p��"m��1�1D�8�{�+�6� �݋S��7��h��j<��.���'�l IV�h��C�%���У�o�>'�'&,���>���&�tk���\~�i#7;���������r���GXlxVHYEB     400      c0q�B�����1��-�VE���7�S�YN����:�5��h�F��]���B�V0s<{|x�9���b��WJ5�bi�l�������������h)(��fe�U~��qU�h��M1P�����C؎� tzQ�G�H��o��) ������q廒b��AI��#q�'rP������]OE����K����XlxVHYEB     400     120�� �63�"�:��k�$Υ�m�����l5|�i���EUݐh�\h�R���+���*5�<�m.Gҩ�Q�ƕ�Ek�5=n���g�'M��O�)7 LV|$����^	�u�P��� ��ϔb6�5��'�}��j��BS���7T�@W�b��iB-��e]�F{�#~+Ʀ��\�0���#�4�,.'4�"Sq�,��]c>z:G ���o[�n~�T0��'5����4Y���r�|��l�K��9��Y[����Rd�f����*�-a�wH<�
���b�JXJ�XlxVHYEB     400     120���@^�t�=)�Z_¿`ꓹI��b]u�)�~���ԇ��m w��v镝s�:q��7{�����t'ϫc"4)�n��6߹� ��B��j�����u�Hg��iX��
��Z;�^؁��B�GѼrgÆf�\��v��"��0�U��(6"ꁱ؞�,@�H�PsWd��^%�Vd�o��\d�?h�������k�R����M�,倾��
V%pK�r�W��£��"���G_�1(5���D��pʔ��NY�dљ��p�'�%5ѥ@�@�A�@���\�E��c�XlxVHYEB     400      c0CX2F*@jL�oKc�����$/`�Rp#Q�l�k�\R[�N���5w����1S,MJ[ȏ���o��?��`���$���@J^�8�UI���M�FJ:��Kn�7=�@�?��6��T@�,�#�Ií��1&m)7���j`����$a���2^l��#̥
r��	��*o1�
���`���",q�t�ƹXlxVHYEB     400     120Z(�9P ��%ȏ0�C��|yh(U��^����ǀ"u0j��ވV���,5�Ӯ\<#	�<S-�Ξ�3WPS�����,��6��J�|�q͍$���o�ij�X��ښxI��ֱo�]ձ���Q��@�xg� ��)���ћ:G �S^QأDNxeՔsdr��)��'\������r$wA���%���q��;�.�P����VD�<~!s�)� ��`���ǲa�h��o��^J�}���2{rWKF��b{[ܗ徴�o|Y�E���O���V*�Ju���1���_���YXlxVHYEB     400      f0�L�D|�*��2>ܖZBF�I���i�/Z�L���@���|ok��חe��F�\�p�-��R���ȯ�C�
	
U�)�k}E���Ef8񊏾���^;Ɣگ�-6l�}S}�`���j��y�l��sd�k��J�du�hGW��5�:��(�)_84��S� L��j�V1�#q#�@���
�$�7�V�U��SO�46�;Gy�zjQJ��h�(R��1�wK�����~[����4kXlxVHYEB     400     110������h��C�Ĭ�������Iҵ�P���0�{1��hX7#<A"u���N]���q���i��&�>�7\K��r
c�<��m?���*<��`x��:.�vG\3����n)�!f@����O��x�܄9�K���B48��X�=�G��Orw�k�J���`�M6��fe\�e�
������J�!�'��=u�� ��o�x��+���tL�0�l ������t�JK>Vl>RE��8�d"O2�����Fja�U�7ޤ<)�0�"^LXlxVHYEB     400     120e��8�*�l菾Gp���+c8�� ���ѵ� Ŕox�BX��-����9�Ya2���J|)S���P)���%^���ۭ�Y�N��������">|�}F:;-M8�</V��]��|BZ���6%\�v��J���s!+J4#a�8��Ty�nh%�n`�`�{�j�o���Gm!�S�ܤ+���/����,:� F�w��z3�D���1+�C�u��"G�A�MؔpB�}�`)KC��{�D��%h�	 �����Q֯�9)��l*��#� ��L2�s�O�XlxVHYEB     400     120�nR���gd�u��K�t�@0���J�\�$c�
��j��o�0��3�fc���y�X]�)v��9����¬������d�-�cN�
��4�џ� u���[��@:�Q�_I�x#�y�a�9�����7ߏ��5�9Ռ ������,��@�}��9Q^֜y�Y�r��"x�A�	�Z�&��:��{}VBQ�?	���^�:_c=��̗��b�m�
i���-|24IVfU�z���pe1� ���﫛�.���Ԋ��g݆��a]��������y!�Yt�'k���XlxVHYEB     400      f0�{������M�W�U��W��v�""a��=�	MM�Y�&.�S����c����\�:4����%1cX�J[Ol6���b���u=﬐��9(m�s���f4Pr��}v+��K��2Cd3 �5CK=�%��+4��n5����U��խИ�Tt��8�?/����8*�����[�81������+Hlr/;��@�KR���"��D��5�h� �+���v�����M�.�XlxVHYEB     400     130�4�cD��Q&_1$��@iԽ����E$�5��C~��-y�`���K{68<z�͐��ړ��g�,�li�r�o��Mt�������	�c�>�&�n��}X�:(!sk�����,����b�� d]��Ga�}���O�7Ѥ|�����I\��:"�Uo��ǅ�+#�+RO�g,&�w��~�$j�ʡ�[-����"����I�S�vn�m�5az��aC@�,j���κ��0
;��۟��8��B�����o�@e��0Fwr�,�a�Tԇ.�Mc*~��#(�Qu��1��V<��$lư�]$�XlxVHYEB     400      f0�5�q�0�:ǲ*Y2�1��p��h3s���B�N'�E6=����4TUB�������oTxo7.ٗ�?ӅT�"����N�:�p5�>㠎2M7^C�JC�����6$*�ɹ�M��Ž������?��]��d�R7.'��U��J�ȱI�)P��&� ��Zsm��^w�		�y�� ����}=��,s
ԓ�\NJ��_�T#B\ ��M��79�:_�0�B����+�o����/XlxVHYEB     400     150��b���9�tA��-�	�8S��1�:zkp=��i)���8b]��	�*�3Zl���%���e���RY D cW��q�ovx~�ʥr�R2z�&YE���`�pqow�|bN�*ʢ}8�{��K;����%�;c�(&�9P�eU��j*���G3iS^C��^!k&��^�Jď)O,~�Lk� l[���D&�|�<kC	�SA5C,L��o�ry^��tu�u3����f��\9j�F�#�����6Y��agM/Z49�}L�fC��	ަ�K6�o��0�4��>�D:$f��h��"�����kR��p�p����e���6 XlxVHYEB     400      c02����'֛�y߽�H�F�㫭���� <IVO�3�I��=��v�����¦kt�e�H����E�Ѓ
SZK�"���nw5���|i�q�{�����^}��)?ٱ�\�X:*(c�Ia{��A����zY���D��bM��+I�!%!�o��$��nΤ� ����\��C�q�nH	���м|�`>�t�XlxVHYEB     400     150����	$��B�M�Dz����I�x��Hp�������t8��>��Og�<�~�0�r���=���E���C�B&���=���ߗ�ئ���n��J���
߈6��}YӤبҐ�C^ޟ��Y�x�b��a�FEx��}#�0�k��� � ]�Bdlmz�d�2%�XE'����LF*Da�z�Z;���W�&��E���j}�G*bIv�����V_'	�|�s1	�!�Z�]Sh����w�M{�J<,��}���
�iye���5�T�v7��0֐��=ؿ�5�*�L$)ژB�:kMG񛎤 -�F�B�(X |��vX�H,������CXlxVHYEB     400     140ܙ��O�m��r&o��*�M�1��M�1�,��y@��	c�b�͖�v�`�Z�X���$҂��ȐÙ��[�πG��{uy�P���5���Ě�+�<��zŬ�o�'˨��"���u�`�^|�7�����~��NA�I!I�z� �zO�t��\l`n[���k�I���z�І}�77�F�[����}qʮպ�Uş�����d fb�������"�Y�vr�v��/����Q�?=SΦ�W(HEJDf�v��\|bq�:�;�	R�͹�Hg�Ik��f��_��u��H�x��9
������hz��8�T�px�!��;XlxVHYEB     400     100B�\�=~a��FU&��y,g���(	�ٿ���
Ux�V��ԇ%��c���i�0�d ,�	�W��hs �P䪏����
!�j�r_)(�KUG�aY��H6�Yh�e����/p��2̒ޡ��iH�en�u�(��$k-��hI5�'T ��/"ÜA��Q�q�� �I������PA}᠛&�-
�s�{��{�_���2�ZP#G�~d��~haT�V�7�1U�����% ��b���0?���tJ,�S�PHXlxVHYEB     400      c0 ��A�p�WG���p��%�$��M(!0�+E���JR�Q�?iZ�'��_�E`�ME�@��4ی)`���̍�#���m����F}�����.:�[�����En̡BK�\`�l.7?N�B�� �~ Eުped'�Қ�U$'�ZQku�3�$Hl�(0��$cH5*�w�M�ǭ����f�grg��XlxVHYEB     400     100b���1~:2�8Ɯa֢��]����{nҏ��7��7�3�Q)��II/,�s�Âȏ˙r�}7e����*QQ���v:2�Co|	פ�`�?�� #��M/�s��Nt�+v5��0p��)2� �+��nupȧ��#V}�'��k/br��D0�6�*ic���6&c�	�@��W(RnԳ�P������=i����߹Rx��h'��X�����\�`�p��QVx~����O�PѮ��g#��f�s&XlxVHYEB     400     110�c9�VV��&���Y�6Ӈr�\s��()�#�{��{���#�I�����Z��%�&��@mVݶ&�1QΉ�1Q�D�3<F�W��D��|�C���_V�ۂ"��ƀ'[M%V3f��'sY�Y�Mq������Dsφb=��c+�����D}<�h:��/޳l9�4�y=��U�+|��~*�C�j���(�6ܑġ�ZE��K�ܓ ��K�{��2�1��B{�'�[����u�X��Gڿm��7y䋁[�2����%X9Ta.��XlxVHYEB     400      a0I&�<�Xf�eX�X��Y��~ �$���W���⺺24E�+�1�c�������-��4��괏�gW�X3"���wG��`{'	v{��V��"#tIg��� '����Y���VX/�y�QZS�'��f� �̰�`yN!���
C�Ơ��Ӡ�a��XlxVHYEB     400      e0�.��Y'j  )W
=yy�����^⁪-ί�Bzݛ��[O�s��m�ž��8�tl����Vo)��!O��4�%���o����)yƓ�Q��têa���j�6������ie�{��10��n-�`�cs���^��(3���ы ل���
c�A����r׻q�D�djZY Kw/���[UǏ���P�g{�	F���is��i�S�HXlxVHYEB     400     1a0���XXb�!&�G'|z�恆���LǷw
h�j����/��+�Dmc��<�<��q�I����>�Ph�?�� ��9������$r9���(%|D]#�?d�_�<��3�y�����ߩXM�{��
�sܪ�x<���"gܯG���l�.
�J�H�=׈:�Z��ql����=[�X��@�~U޴�(��9�B���5#�F�H�]K��Ȫփ��Ɗ�����Չ't�Z�����!e8_�ޫ�mg	�F���Uh4�Bԩd��Y����_�YZ�lzy�����e
��Yg{M��6����Hkx;�^HGCqy����4���,% �1�W��zv����������°�Hw=C_�"zY��O�Hj3'�Zz���xF
+��^���c-�q>�q�Fl�XlxVHYEB     400     150���6G�V(�
���/^��2dӯa���Ð�'_GAʐr��$4ۍG)	n�
�_|B�ǌ&p�Zʻ�z�FfuN�1���S.��b��=5��)��4z��J邹�Z8���"��$�qy	�0�c��06(9�G��5�?R�+,6+;\��6���
@*-XrP�7=�R�7A]��T�ן�m�p�<�Y�0�v%���͇�����>:��!��3%��U>����uy�~d3Ϝcնk*ᔧO�>�-�v���S.��_�����P��vz��X�}~�r֪3/�H�c�ɶ�|%F"p�.��mއj�q�~�Ә~�x�*+��)�XlxVHYEB     400     120��g�u���u��/�w9�.+�b������Vx5l|ȟ���g�s����L��>Ċ����a��}�)��XN���c�����D���e��q��\EƧSRP삙Ļ�J�Y��%y6��Oʒ3�����>
a`kUlq)��)H'�M�MR��������3�T|�Øq�Ϩ��:{o�#!0��Y��9=�5���?���%��RcV�u�$8X��	�xE������%�v�%^J n�����5�e�����<3����+�fv^vfл<T�D�ǅ����XlxVHYEB     400     1d0�:XB��Q.�#����8�-Ё�\��-�Հ��V��w|5e~�EM�!�K�yY=B`b�o�[k��*1�LMb��H��O��p]�J��4�WJvt��7}6�' >Eąr&h :ꊶ{����y\d�3��d�uD3�bC�w��f}��þ�k��uq���\U���J�Q���u}I0��6%e��w
�'b=�����01�LKh�� |<ٵl�ى*Ho����7�H�W]����T��b�~'�{��s��������!~"NQ���(nq��Q�j+���u��魶��>�Z�k�Eҕ[�=C�߼�~͈�a8V�BN����Vg׳ך�a�u�r���7C�MHX= �U��[,�e�!��̨@Hp��K�oK��$D?��ቫ���f�%���c��X 8���;�ݧ>g�=��'�'>j2��n<� JG/NM�M��r������@{0����D�ːnXlxVHYEB     400     120yQHj��Q���Ch��.*D�Fh[��F�~����eN�������{�x�	�kl�CRl�߫���%1Vc.�<:���ށY����Mg~�;���7�Sۗ�Z<A{B ��I"� ��n�e9�����H`�z�Y���(7���2�m�]�Jz�����|���������S�L4�/(�?�����z���>��NZ���[�������l:(ds��ڴ(!�%3�U�#�ı�9a���n\{DG]�G\��9���N�td��L�*�L?g�eL�XlxVHYEB     400     100�(����)J##��_%v�}x6����Li�g�u�#D�֫�'�$j$!�G�լ&ٶ9��̫�@D��&�*V��fl����դ�2���-z^�	�fSx�{wa�D�욈�>�C��Fm��a����kv��[�=�D.�ǀKz䮔�L�s�Xt��@ �@�{�;o8�'�m��;cl���E�r�B�Ҽ2LYSО��ѸFR/OY/ ��0�%�fW�K�d���\M�m��^b��$Q��}���V��j�`����=XlxVHYEB     400     110�t�F�P��7��jz��=�d-��E��@���:%Ks��ڔ�$~����M�J!4���g�C0q�4l�ߕ����F�(_���އ��Ff���j�͌����k��I�-�5-m?Ͻ�
�Fh0x,�P�)+\�;-��d���x�K�	��E~*�MR���ʠ�[Nr�S�����5p.i����O>�Y#�^��~?��'G��
 �Uu`�"�/�:{�	�x����bi3"�ܙw!��Q��{��v���^ɛ���XlxVHYEB     400      d0�V�(��TϤ��<���"����ZeG�����g��Z%�y�X����7D�|�""m�Bq�b��Sɘ	�S�B�̓,& D0=��#�����H�{ES�*;����g�<���X���� �e���S�ʅkD]r:��Nǁ6��8̽�y$S�f � GQ�
1���y�.��1D��~�R,���k���)ڪޟW�:OT���������XlxVHYEB     400     100��2L�&�(R�eq>���S�×�]00-,Z��)�y���e))�Ƣڋέ�Ԩ�`��ny�I2p�K%�޻
�ј���fv6D�CcơD��X�,���W6�FN��	��&h�R�0�����;5��,='fnfd��4�S)zNJF�f��,{��g:�X�8��7lv�ӝ1��+qʇӒ�.�';�fZt)x���NoȒ�tgf�R��T��y2iw�X]g鬪c�k�=z�ہ��!`�S-��+.�:	�XlxVHYEB     400     130�t�%첖��eÕ�"��o�l�Zx�X9�N�Y��`�|��#���������C���ȣ��u�=R/�����	̎b�	i<�ݣ/�t`�w�ip�!����I���u�*k�K��7)��=��.f_l�m7,,=N�-��m�^D��D�?��yl7���[�e��K$+_�'��;��e��vU�����$驪ι~�����BL�����Z�A�e�s�bqd.Dc�7@I(J �z	�j�iB��s���� dKc���C�
��x5� �յ�}�	FV�0�NM�:	�19����ɍXlxVHYEB     400     120�T���TT��\�GԢ�-���?�<��D+fW�{W2�%�<ru,?��k�r�A�f��[=P�/�3�B]�B/ R%`���l?iJ�����cF���C<D��Ì��bU��Ro�WsR�8��>8�R.hb����2��+q�����ަ�� �6Qb�#}�V=��A�6�͕@�y_+�|��'��J�[�e�X���Ɠ׻��zAa��o���E���ѥ��qg��-/��1�� Gn���p�Ψ��~���i63
�H����j��j��XlxVHYEB     400     150"���ţ�f�!dh+b��a9f�(��!�Ǥ���%E�Y|\�1ْ����!��\)�I�F��W���h�X�Μ�֝3�xv$I��u݁$%,ͽn)ݡ"� �7�Ď9H��F�8��>�l�(�H�bH���+���>>�9*{���G���_��AI)�]�\wWY�Z�_�ꠢ�ؓ7��M����9���+UN�,��`��a�\��l\q�`���&���!��Sϒn!�~"�1�t'������P�����V0���6��ڣLD���	��P�	th,�_y"F���f�!!+���H��šv@)���4��rt�i��VrW���	�rXlxVHYEB     400     110�ң��!N��
:�Xs�|�,,��pg��ܦP,Lac}8��BfI7h��-/���KT�b5����Ȑ�}�l d�m�p2�_�GU8�L�3Ul,�y�M�+� �W��8.�޺�`Z8�n�1���J��lJҌ�#ai�ZCWf��-8u��¿Lj���uC�^޸'V@�!���:��o����k	{y�ʾ �t��^L���V��m�Q��}#5V�yL��5,W�]ʈVZPO��I�8*�pǊUb/y�����r�}�>A5XlxVHYEB     400     110Q;�9kk���[���h,p��rq_��8���w#D�~u�,�#ok��U^ڞ.��6�@��v��ʹ�+JoJ��8�RDm��ȃ�6���S�,-�VT��YāR���s1}�9U�d�H�RF���	R���-o���w���W���5�t}/1�,㎉��	�(Y|	�c)1��"X�F�i��8��ۦF�v���G���8�e�<���ݸ�.�n�𠧦XJp��ǐ􏱅�*���x<��1Ǡ��6���Ⱦg!^G�;��Z�1>���<�P��Y�h�XlxVHYEB     400     120�9��=�u�׬���z�鸖��1�iI�'/�~?�=��v�QvnL�yQ����"
��R��x]Yxf�����p3}3{���>�o�V����n����ܲ��JXP#d�Y��~r��D:X���T7c�kw �Pkfz����k��,E<��X.-�54�F��)"xZ
j���0�z��9�$g'�{,w���v��J�k
�_��fpj\����-�=�Ow�6��@�8`p�	e�VT�J��!;��% ��5@H����� �}�S*�హRn@ɑXlxVHYEB     400     100�ٚ� �v�X����%2��ߠ��"���`9A����Ӫqt���d�L��J���-==Q,E�X$�Mb�;��3!pP�U�𒍬��5�6��h�~&��1�l�o>o�ηo{��H���>�z\���Ԣe�X6D;P�68k2T����Y*��x�V��="A�ݬtD���7�_Po#g���ҥ=Fb�\���/�[wߒ�(��2fv��C��c����Rs����b��*�` J�T=����9P~�2K ~XlxVHYEB     400      f0���
�0�)��O�t/Mk��R�#P���>+�ȢcG�%�����8��טgKۿ3W��M�e+Vs�z��/�0�o?'��mV���M���>���;�}�+L��nBAW���Y���՛��ma���,��D�>����*Ikb���o��� SX!)��~��x�4z�Z�C�9S�UEɻy!���H���������C��J�~�f�_}ʍ�8�G�k�OGB���7i�/��[�XlxVHYEB     400     120`]A�����6yt���|:u�E�*����9�3��6Q�ߩi�3%�q�Tv��]	��/
����t>�*O��24��	���m�Od��ף �d9��<B��k�Hn�d1giU�(�^�c��T"�^��sB����Lݦ�'�V;D,%���K��������V.{h�v�F��Ձ��?�/+����X�+?,�O����_�5-!TG���EX�L%S3����\��O$��@l����:��	��ϡ��An�ӳM��XNw�Kt-��d��[Xy@�A��␰���U��XlxVHYEB     400     110���)��T�{�3�F����c�dI�2إA>�,gO�#��^[� b(Uz5�qLٙ=��8������P{�ި��=p��F�6��w�zb�^��}�*Na�Ꙭ�~�d��F�k����-��8}Z�H
�l��1�K5�_؋��#�)�l�,ɾ��k��]�s��������1�յ_Y�*<A�ޣ ���$%����u,�*{�^�u�c=�;1Q^��6Y����M�BJ�t�.����H
P�$v��n^��ܔd��Ms�$ǔ�r��fdMXlxVHYEB     400     120v��s�9H���F�����b�B/���ъ��m��Ri�܌�7�g��a���_;���30*:��O�s�swi�K;�7���2by�pty��4����#�;,���Z!��fY;YR�22ZdA�M��x����l�*��S�7d �ꟍe������R���Qa���I�M�\|ۮŗw���j�E,�3H���י�ή�����f���Ԓ)�z�5k�+>h�)&}�Y��Z�.���р �9"^A%�����'���{��s3�[��Fg�R�0�5��hXlxVHYEB     400     140�a��ktavd}���5�M6�/�����<�T�<)�pB0n-���3�?�z-X��S�-�V�K�Q*�m�Z��>c��@�b���Q��-9;k(�i�[n��J��/QJ�7���z��|>N;㣪ȁTŉU�2�
��Xn6�W@>i�}�Q}�g�H{��H?J�Mrt��a�X�����@d�$/{tw-�&�Xƛ�7��A�0���8?ϕ[��@���F��o��ɧx�ԚRq�`)��	�J��`
��"����b����_ �w�/���s�����̈��)E\7��=h���B�v�@�KXlxVHYEB     400     140�3�
�����`l����_*X%j@��}VH�Y��XjP�7�����J���x���z[����'DD�0Ea1G���u'�i���q�C�!Vh\ �U�+���C
dePS��Ř�=��4x�0d��x���}6�ަ��;T�e���@T
� t�\��T93ħ9��$�9����Ъ�1q�G������룦�'�G��;Y��"��f�=�Da���q��L����Y�^ؓ+!��A�|�"⢢�L�QC{W���*��CԥP�������1�YƩ�.@�9�g�O۫�8��?.�b�&�XlxVHYEB     400      e0}��`8���
���a+M%��6k`;�3A
���ha��A~���m�z:8��~,�����9 {_9����R� �»}�a�A
S�I��xs_�؄�f���'K����9^%9�D����r�����za��U��X�QP��B��G����	Q�3�/-�!&q�:���iy6����o��N߬����,Y�S��ډ�\7�~��u���`N����<9!��XlxVHYEB     400     140��:���,<���^9�۱� ���&u���L�� �����e*�<��E5j[��xk��j�K����z��Y��2��:�^s�ׅ�1:l�J&������G��D�mM�B�>4�mK��6T���;TQSII)M=i���,��-�<�G;�}}�%��<^)3��d����&�\)y��|����姭�8*������O����x�)I�Q�l ���
*�QHR�Y�h�sd1
e�?7.-R���M$,	N��t���T"p��j��Aӷb���j�1t�
~ь��d)R�&�,��B��]h|XlxVHYEB     400      e0�)�h ��^�;v6\p�#����n$��ؘ D_�3;��Q�<���F�3���lFH >�D��L��Z�$�Q��/$ ʗV�]|�`��0�i߃gZF�P��0Nz{��F����>+S�O�l&����~Gr���U�Ǧ=1&H��0i(�B汤�I��;�F�.�t�7dU�)*Q]�^�&nZ1AԌwhͻ�d��ӑ��rE�O���bA�k+���XlxVHYEB     400     190���Kc�י��4�G�xn��k XR�S��_� sJv�"�����c��"��6���6�*%h���)�Wp����5�2¶�]+���2��✽�ot�6r�"�Lƙ�{�x��}�V+b~g|�6&0bU��,������95ŏ��	�A�T�מ'��h��q/�ۻ�9 �^�Qw��:����J���h�a ����
F��s��2�^��x��+<i#)��?���Zڜ�tL�m1Hv�ﰅ�p���y?��4{�"b�U��	���+©R���W*f�z}+�����,��-����";$y�4��@��|�����d�H�
���ul�O&(���)_���t�S���ʪ��n�f��>K��v0u�������C)7��XlxVHYEB     400      f0�g/��OM,Io�7>�����6��1HL��)�/W�0��6ρ�:�%��u��{E~��3��6[-�
�&����ׄ�X �9�1�h6J��3�e�ê�����!,�!K������t�u�<A�.����g4�i�u,H?�葉`��F�\���u�m
�(�⸃^v��N_��-�ErubbB=��.�X�9���-BX��5	b ��" ^;`��Z�@��IDKNq:XlxVHYEB     400     120=�MJD3t��8� I�w��/4^V�2�z�c�g��T��m/Qjc�bk��SPy�y��d��j�v�̖XJ��� z��g��^߱j�Fn(D]I�a�Y T[XШaV���~?� �t܋>��u���'����xU��7mݕֵ�'����>�\�;GSv=F=M�d�wE�h��y������$d��4/�ozR���[�L�YZ�0���m:�B��`�K�鷻˽�Y�$�K�Y�O/�V�_�k�� �c�^� �}aʸi5���-"i��35���=�x�r�&�XlxVHYEB     400      d0��7A�(����y�����Z����P[m�o�Ǩ�td��q����<�J��N-Sp�����oE�[ ��%s\�1�f��M���q�n�"n���Xd�^��p�8����x��襶bm�.-�`z���2�@�d����}Utڦ�dD��Z��?�����BTʕ�m{�`�ZD&�p��SS7���^6�j�}L��y՞�K�XlxVHYEB     400     150��2�gE�|�X��5��n�(��>�"��ʏ�Y��ɇ�z�,r䙨��3 C��>N2@�1#֩B�<��vg[�Z��_�WV�����k�q�\�7j�Y1���|�/�ͶZo=�o+}�Za��3�G~�`@b��,,dG3�� ��^��.k��ѧH:�����J�61������dU	���st�鹨��s��u{(�1"�o0˧t��}����5�b� ��us���Cx��1�`�JR���&pmEEa=�J��ab�G�p'�Gs9VԒF5Uԁ�q�H�B|��(���j��Ca.��m��RLSPi��\�wXlxVHYEB     400     180�By"sﶓ-���2�3����ÛY$.Df(/�xܖz�t,��'m����s?a9�����Ē��9N	�r�h�G�iI�v+\E])�A dQǠ�B�W�iav~7G��uȸ�r�?�!�:$��C�4u^�?�D+	����j�ݵ�P�.^3�S��lw].�usNF�#�b���YU�\�Zo�%��P��3UNXχ�(�F����ܚ���Ҿ�K�O#5�6t���!�I�G�k\�3��[�b�iߤ�����C�m&iP��<�ƚ����Սw{��䵀�zjVP���(-����'$�����$ߠ��fB��L�qve���C��Ï�#����| ��rJ��a�弶��R�P���Xtœ�k1�J�mXlxVHYEB     400     120�l��A�x#K�K^����Ϗ�䐅��� �P���  ��AC	M�@qÙ-j�e���2��M#L�g@�b�k�A���o�Y����`��9̇X=��z �5v����u8��sv�#f��6Y����f�N]Z[<���U��ez���LH�E�i*�5h�y!���j ���p���H�ɧ���㏪�:�l��:0�<�����Qv���BBE�^��8�g�ڙq�M��aJVV��%��xL(����G�/�OU��9�ފ^/��t�����2�Җ�eXlxVHYEB     400     180A]E�*=�-�y]�q�Jy�J�ayWo�I� �+vI��D�<�<�UDfmq�^��_�_�]�v�JPHY��}zd�p��YX4��]�h/a�zk`��2�%��Y�GCcP0��j�|5���ș� (�{���c��T��c�e��j�Ν�a������;m�4��jώH�D[��D/Ҩ�RiD���ӵI�mM�M+���+o������~��H�{��H�(�lUi���F(�����g-�<]z����K9]�a��c����)��
����JC�I֫_Ws�i��s���V;��l�T��^�5	=���~��7��-��X�)�e�(Ăz$:��M�M�������A5ub�>$����b.�SO[�����߅/���d;�κ��XlxVHYEB     400     120)}6�L5b�-��d�j�*�A���#v�v��.�I2�3�I���PR/w�rS�;�$��*���?:�J�Q��(J��t����p�<��$�T�J_�kJ����r���7S٢0�6��B�(�K���N���aR3�>dW�ұ�Ϻ��o�����gU�[����Q_��v;G�?����Pc�[�94�d��_m
~���)���2���
�mU[��[/�~��9��g���?���j�z�h^��l,����f��x:=կ�2�l���7�AN&���rXlxVHYEB     400      f0���]�ܼ�$�����m�!��S�����V���F�9����v꼆�>WXy����	@O��5�ޒ����j�j6)N6��s��Y�o���a?=����A�u�
xa�>�O�]L�f���퉻�e�[�vėp��L���'��2���$�O &�ݩp������t��Ҁ3���Y��b�9Ȅ.����d��T�}	��M2s����tXh��z���0�:�Uf<�qo�P�2NXlxVHYEB     400     130F���D�����A4�A�zv��h��ٕ!~s�V��M�b�<A��I:`j���9$G�B;��x�@x��=빿}�����'s�v�rX����a�u�_{�h���i��\!�$袘���u�p�n? !̴=_d����z�-�\��`���.O�"��ވ�!1�Fm�������E��ܣH��䥒�^�\L��������|��d�n�HZ�F�4��D�?y�-��Ķ/B9��M6�S
���>"y�K)�3&Z�@]W��>�YT�5�w�Y�P�+�9?-X7Ve�&��fmY�{c�\�8XlxVHYEB     400     140��Jh���SMGu���`���׏��,a��:Ս�7A�$�23zzܐ�t�	�IƮ�׈:�mm�ld�������w�ß�Dk�T1�Vj�wTM�Klg�P���V�5QzcR��&1E˻3ݪ�d�'�<�GA����d����B��1���yH�J�pѵ���s��m�ī��H�n�[}�m��v�1��IX��,��pz�-�ؑ��V� �U�B�d�������A�M(�4������k��z���r���{Mĵ0;E���vU�^�K�4,)D���M�k�u���D���7� K'Nt�i����9��Y��w��s�XlxVHYEB     400     140%CfP ���r�g�R��j�����IMG���O�b� ��1掠��%���������PqƢ}Z? s�K�ϒ(��Q/pX!D^=��"��"�fzi�/����΋UB�@�,j�F��F������a�$�u#'��⛹8\�%J�H�Yiv�����S�Q�?�x�����\�$^�jj��D�㆖���d��2�$_�����5]Ґ�����_���_��M"͹��۵�f��'���BZ(����4� 3@�q��lg��U�?�:V�� �U�n�
��*�����Q�9���y�XAO�XlxVHYEB     400      f0�r�6>*��*Q���ʏ�;��p��>�-�n�v]_,�֬��ג3��!�*>�� M�Ed�ΕxzބOq�������Q�K��Q>���,b�U������I�f�{�V ��;t��"O(^,k�n6�XZ!���8ul�hQ�0V�t����Zm�U����]yQ_���p��V�/Z�x9��#L	�����E�!G����;��Q� �Nn�[I�����]����J��&~��LWY�XlxVHYEB     400     140���)���g�e��%H�Z�}�*�/�fKC=�,$+C	v�ᱼI�x�����5*=a�8W����s�+���bL�"7���x߸�$���~	r<;���7Bi��N�GY����<&$��v��$¨�����b�p��$E��A7��4�hV��\l��k^�G]�e);�U�X��q�מ�E��TŽ������;���3c]�KEM�{߾�^��\DI}æ�֯E�b�ѢK�������fC��I��ɜқ���J�?��xet�Ms�K����-�z~��\�5yE����a�<w�6q��{���H`����� @�zXlxVHYEB     400     120��ւ:�F��pj��}XVC0�ߑ���m+<�nf�� 4�����Pz�T���"J��o3-����47d>���C2p��8j!��I��/�9�B3�3�µr�?#K.�1�&=Ҧp�gk<sA�6l[6:!O��q
m�O�^��Жfow��`���W��"��ߎ��9.���*	��C�׀EX��Pr�^��b��{����V$�&�G��N��q�ҥ�5��2�Ȋ�D�}�,#��Vk��0#E���}w���Z9�J�ȅ�����<ޢ�A7��4��'>YY]�XlxVHYEB     400     120�O����#�a<��� B�[�ny�-��*r�P6(�_��x�x�Z�Nd���"���E�3���PB���>y�aS4��Z�#A�=��G���Li������
��ls�q��U�N9�4�;޹� }�@š3��GdB:V��j�y�����^Ձ�uy����2��&�9�˃�]�ۅ~�2.^ F#������J1��4��E9rL�{�����XUޜ�<�9˸�;����&���/h�������U?$� Zp@B�Y53�6��U'�XlxVHYEB     400     110�q�H�"aR�J�d�Y��L��`jޫ�an�bj9���H��ܭE�Έ�)�c�9l�dU�xչ<��@'����ڔ�y��20�����i�n������,��&L�a�y�8E�{���m���8!/�t�"�+],�%���e������x�G�>��*�@����h�`�\8��[~��s%�����Z(�M`����J�n'F�ʎ{C�'���5�� ecӚ�����
O�
1:���UM'���J����	l���RkOf}k�;�XlxVHYEB     400     1608y��o4J��5�b��a��0�?�0S���f���P>)�.|�Cz��c�7��Rmh���c���Y�Qe�NDh���6g��8<��E��ms���YC��u��������{A�������o���7�?I^��؝X��Y��pg�(I-B?	]����f�#P��=���-Y��6�kaj����?.��{If�d36�}F�Jk��0�,6����iF#b�.�m�6cIeGJLp/���f@]ƶcK=hj)���7�!��l\�����rU�J0�crQŤ���H�Q��Y@�⨇G�2ep;x��	�!�ͩslx�"�Q�Ji�H��Duy4xۉ��E� ���`9_HIXlxVHYEB     400     130~֐�~��<�8��\?���H�\��l�;Lj/t|�-H�W�6��j��>���6��V��nه+�b)�&E�)v��8>Zpss�.��+���[�h�C�|"'������h�tb'� �����Zb�F�7i�Xh�Y�`�nh��e�_��(.x�Ẇ
e�!�0��m;ޣ5
=���a� L��W6!��OU�Җ����4��P��֨�TZ<�CAnm��
�d\��*�~J��0�?j!/}}S�@avL�g�w	g%�H�Z��N�أ���O�~J�nD�fp֨s�S�v����XlxVHYEB     400      c0m����@hQ�Tz�b�WN�8;����mU��܈5�>TQF��
~��F{i��wv��aC���q�Jy�p��/u���?X����%�$'=��kS�*�������$��a��w[җ!}�=�v1�l�M&'�JmJ�U�\�B]�<ML�ӭn�S� 4Dɥw"0�~��&O<�
T��i�{�L��XlxVHYEB     400     1403胀-$��i���6ZP)5��l���쑬;�Np��
�f��*dv�!+L�'��蚆 �i�pcNco�DZ�{ł�a.���YX/zf�ݩ���tCޥkn����o�dgg��j�M���|��U$�Y����֦��}�����dvT���^{W�Yv��wCp羓n�y4B�7��{X�q�p��y~�d�S��@}X��̖v��6��K����i��/�D1���xw޸���[�̊	��_K��޽��&�a�l1Ї@��'�K���a��@S����!�OR.�'�Bu��bb�c�\�B��������XlxVHYEB     338     100�+�GƮ����S��R�hbj$�&7� ���=ItPV6H���6�l����f>��@a���cҼ4-!De�&�U�WD�M3.*S����\A�8��Х�O��˱�U�P�[�p��S���3ZY)ܵL@��Ʊ41��� ��]	)`���ci��j�_�(�%��˲�%�{Z�<u����-�8�m��H-���6�J����+j�lm��v�d�Tߎ����)f`s}��2,����}�e���~����.� v��4�N�r