`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
YrGiVW9flYyYKUVn3d7U3eHEEKckzXT7S/Yi/ZiXCkjjUT13VieUOcsWBHolfHeP5wAcXY50cY1o
+2Ih9/QinQ3o14KNebrU5YXaNuRGziBY111ZOsZD4JYPbaYKhw57D1DagFrRvln0mT7uqQhLnvWg
89E2YJXqe0Axnb2UwPgwI2iosqlFENoW3F6ZPu1XIRfaqs87CcTw6CdClcLiiqmDey1FVE7/9n1B
5wgFy4usEURXEDUmwHpS0skMAlTm0tqj8B8pJ2J93QV7ZWhYas2tTUJxzb63PI6okP1vqAv/mIfb
5gYNh1RVqc9faIPeHC5odMY0UPIKeha7Al7Xdg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="lNVoUPF6pphH9WbRZu3JJSA+iOG4r1TyCPOA4UFd6rA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9328)
`protect data_block
Vg4R8qdbP1UwtbDgKP/4UjtAAxwRY9hiLoytwCjtKHQDROY2w/KFGM8h9OYjFIK79iePqqvrW94T
W0hMfKcjDJjDvBQnnHQxSdPvF0OCI2mH+3PqJcg7Bh8hvT77iGJYzYh9qryxd8kKkSebIrgv39aO
XIwB4S80lrLLqDKbBEP6OlzEpsS7EWJuAC42s9udGK1ZLzAJRf34Y+BO3pA1Bqx+zphU2P9/AttB
WfhvmdJt+0VWzcrH3ZNRWQ+Uo+Q7xP16HLXwlkNjsNLZ61SdRe8EJDDzh1emy8SIZwAtVkd7TRVd
iAC71YxV36LZ+5IMhy5V+QEISiJVyxcL+qtyx6XHvRZP8CYztRP9UnBlCzvKPhyuOpf46fzMPlDF
U7rcnEMB8D4g+UOxBFzo7p/oG0lfmTnLt711v513oz8JWRDXuLTXZUdQ3sqr5LDvdVBWjsMDBalu
LGeweXIlhY/z+qF0io5IIkCUnX9VhY0hYOnryHhw4RG2At7wOTjQV81jpmG7PwPCHf5Y/f4LyGYT
TChrsLGrC8DjxoeAxdu7SAVAJKtTKpYbSfbuziRteUzmFlhFBrKb2Ya1ai6if/XrGoLbz0MQEBrw
TOv0QTYBcYHC9pTOLcvBTz7CuOLT+r9HDEier3ZT/GkqRPPA459D2jS9DZPi0dJpmcNc+DIFGQ2O
MtQSju2AQUOnmdrpJcmXd/WFqsR2Fd2/TsTzemXS0y1khbvppBCpurPnl1oQCuMYCQjijBYQXg8W
VNEF6A2bJeK/ssa/4J7XDUjUMolP1XLHh4A6TdB3MI7J9WruS4mYywL5mqg6aU8XZ++OzyPiFu2B
wo5Eepi7QkPv63xjaB1mSCCcVDJrgKr7PaA5bC7aEP5dad6B2CUfv7V/wD4nbo24rkCXBBVq5n6d
XfAHVOub31pX8AfnSx3XsgtOJt4XoljK3KFZU7tbAD7DSBmXiNJxbXwMax06UyIVrZhlGf7Jv5Ny
yaS+ydMe+DVoIOTFPfF1Qfrh6zFHkl2o6Vaii0qxmdYm1BnWfHAMI27p+jvvNPnfXKAh/issTxtO
fYJuvC8T01AzVqOBmL1no9YlAsrAaDsXlczBFg16uChM4poxUlPKuNutIC6BV2w4/y+2sjR7nTD/
xU+Fl3WdMtlFYBmPJb+bW7r76dBui1fHwP8e+sMKIxVYvSOf0zJjtXBv1t9nCdr3nl4C3+ew/0dm
zsZX7FjhcTSLvprj5IRIKYGtw/C2PksvobuGa1FoejVAITIfuOH7Hq6Q54uZnL32aN3Fa1SEXl/u
thGblRXpcuLlfD8Gm0YdksOwaNWCJSfmeHP4h6fwaVEQLAwHgq5i2AiiW+vRnR3E3T2bL3j38l3r
xr7FTTBtdx09XsE4pQtl2xj96MchgdgSlzJPbofb9IEstmthdlyS5TN7qATA1Kp3lmSfhtvSQhft
ypIx1H2uODIPWLvBswCAfJR3YGxJIf5j9qILcC1dfc1icfMAURYh5J54kwSjDi5go0EVwbSc4hOq
kPJ6mrYi9gbhrQZfQ/c8ujOjkE1ejsXGM6T3YxRvfw9b5MBGlCWH4ynGX0H572EwrKTOO7nlLK9x
jRvCgNAElMkMljldc3ar9ABEILEOQz3RfQHrsUVMB7Lro4CQvGRXi+UM2tiwsSraSfHKZcNi3z6f
L/2Syr6gjpjqC2c6Pexx+n/I5uHmZoTvWNHjZVGUa1PDtn4N+l+CHblzFSdyWhDDwrIFjAc2xBHl
0a1ld1MkZFihvwms6m+5ATIrOJXk8tTCJwBHRyxh31UBMAJj5OADoboOY7Gar8PRPACPDVPD2RLR
OC1R/9h2ONXtFZeESWuzAtWIdhhzQwMaY+neQqez4/cJkbTzoFW2KBFWi7WyFQFjlAEXSGX9XFnx
29J+hrtYy4lF7GdAnMaXUI2nfe9l5qdUw9YWwEKYSRbdv3ZehSN5ZltoTaY9jbEOz2cUir512emi
MFfLbdClQjSF72GwiUV2pk+MDXuPcS03cMHhAnlxYGfxoVzVUB0ixsMx8expyiOTJgqab5TqvADr
YnKSZm6QChCnbeCI1Q+Ug+FVN5LVRD6uRpw0wy4038rdzjOwuOzgaY8ZCBiDdTEFBoR72qeavz4o
4uAuvmuhBarG1L/3pAFmV3XFm9UCOfOvWOB5Xni2c0A7dJAUE9WnxulCVpaGLbBZVQvKdbEprxcA
4axglRFysMv7woYehS0tOR7fQG+xeJ/hyIrN3U9FSjU4lFJ56FTvsDia1gaJHa2qA/OxiWuUPFta
gcgZtAPb/o0+rf3Q9LjipVAvpHxHTyCmh+owMYAUZgVI40TFW/paEoxiXdxv3H3jq8mkz93DBmVa
UAZk9tILTVMnGDCqVW0DzKAP0lM7hRbXf6cxKZUD0rPXGdAB5dDwNV0fat8Zg2R11g1adSRf1WjU
9JuQRsvj4Ud0yqaS7BtxxT7qWiojxWoZVcKcwhdY2njyeHgv7Z3VjZIh1sPtvDtCKSrjw6xzt0Uq
bFl44Gr7Ik+oq03D/hMhJZdCKywXd4vWGhB4MvJK2s700iXYQC5Y9MFUXRThAy3F/J/HRXo/Eohx
t9y1T4RSgMOhDa2Qt0CX+Z3YT1M2IsLNl/iYIYtXOoIJQtqj0yhlq5+7gPXxHY/k7cn6oC5ICtRI
pukKogRw035R8Z0NdwhXnyjF0W7iyL0+MEgOgkZlq3EdgojxhXYmaMM1BtVpyj5h5ucwriM7WFWU
Lk6znZfX4QMYJL4W2Su0IhBiReT8p2/7QN2NPw0OAqGti1rJlzbTWPT/rjjYhnLERM2TinCC4pXf
Kz2YG0OVO3pMWcNONxXl95XhFia5yHCn481P5DPmJBT0tWfiqjiik1qWYlpqJUrSkXhKKI+qpT2j
8cTx2xjlISyVDUrAfmJ0cwZH292Mk2zvRpje4T3L5GT7X8FJ1jy5RIdGItTfm9PF9HVaOKQX7dzj
foykBiqHTYGG2rZErL6MAv1pniRW3FLNkfh3htD0OegZaZw14xDyq1Qn3cwuhYmfw+ZlEQEPt21U
T6pRFOgo5XppdmrKVU/APepMrSejsAl5oEl9/WjvjP4CxFeuSLPAzGU3faQd3yFjB0/TxIvSb3+P
N8m/ejXZ+m3gBNmguE959C8PXnChqG1ZHhxVW9yRZ6AtfKhmsDO+V8/TxGvMq/gKSbN4qvK/VOsv
TqVolTHFsyd8s83fzLm2O/5NB7wR9hd28wMg9MUxn5aWqN/U1+8b0MKQ/nIYEhZ61bP2cUqKgd/J
D14THCE3zfMbF24BXTX193aWCfKQ68m9OJInKzDcJkuDyXNNam7dNIb49Qw+DP2E+uWZnqapas9d
NqeqmKv94ifeAW1znFy9GJWSDj5u3PANX/6dYp1MxBpyBbICzhYCHr5kHWh15Gy8AumWtbZGdd1/
N5nGSyVMIUl8PFhzbFg/P8KDd6oFnF9ATVjxzouEsajfq1T2Lq0GvTPngbkF0W9kvxQ7ZEZpDbu0
OIWHG32KHDUrKsxKXZNJIbHFutYIv76m69rXvTBWXpl/SxXlZ5ID//7kU0UBwsDpq+uknKIp/45P
l3zp4UuMVDuR08AzZ54VC7vxtmVJn1U6sGbmWsV0wdtThAQPv4Nar2eiPrvR6TPReMXdTgTx2LAc
6iiidkGg1uu22UQvdUdQun2t3tA3E5h+8ZDRM+a24GlwQZ3HW/BATkZA5gnb7Abfp3CtitZGHkbp
Z/SQdJ52KsXzMpepn7a0LgKzqsnfo7ZYsQpwSmyOMuHf30ltcF93FwBfyqy3J9K3AM5A4D4ZIZHv
jBUpLQ4jviDdflz8sMpRoE3QBKyAw7aUs0Vh1tqmv03Cba/hn1Fltj1RTSeK2JawquDERUmx/XRC
0Hlv7dbhFtzsGWKbp+ZPUf+33umPaAOdcMZncdb0coCPKnSeRpuXyNRTQk62P3GbFFQN9h3adI50
Sj1syReSzNwYNp6D/Lnt0lBgifkO+SxsoDBjh05/HlOabZT7eIeHu5uxT40rT/6cxxAuC2EAbxZY
7p99nVwm8c8FmbF3p8jcly/JHN1Fu+2r+OIc753QxASq5flt9Kjk/fRkLFulSeRSA/52nY7qDUMT
DvTloSet4pzYMi0AQjuVbrrql7hG3v5ndnTbu+dW3wNTKLVfb3X5s1SCceoA6ag2PaE5hSmhqpON
m/xRIT6UfaI9abWKY2BtivPvuDYtwVtxwiwegYOMmXs2plWGC3Mrb/A4hf9owJrW3C6PV+fzu2Gx
Gz1/rjy5IYSp6vXq7Ps0REV6En4YFqdyxGuUp6qGfvq5yC+yrq7x/KpzxsqDEkm2eThF3U6TMcTB
bNHAvWKbMlgeGtvWYF5AfJQSXztfJD64fQNTXJYLPRxXv/+bI3DFdBAMvVMWroZcjVuTZD0g1R2e
Y7VS7qRUaZZxG5eMIvSQDOEIKaZrkR3HHYAsVPM7vF6+0HIhwl1OpFb3AnGOShsD4uz6HiauqOuo
J+YCL/e/ynZKJmJvs5d8qBIeIQG3fGiLtwAHH3M7NR4vFK3rPwdJvbzFCHGLMFos/BjWHMInazjp
+bQYx35GKCxtkWhpekv5XfNB0jaVQLGuhHBQf08BbehvU7ITN0UVtm6lGVSWry9G9Cbt/4EzaLdc
F2mZaupo/WWE/iRNQdQCSMPM280Nst1OMOkgVJuj5CfSD/A+WQkxSHPaEENwmfcMPQA6MbDZlrEP
5fw3fYRMmL7tq2+VFEkorm3m8GknyxXXdo5hPbtnKi5nu4d48/NqJ4VemTlJx6SBPSgII/Ryzqcu
eJVH2NwQ6c99dVA19jSnDAQ8zsQy0Y64nk+r3CSM5oDO/Fexq8lzs10k3VWnoKOFinc0tV3lCes6
iwradDTpxjuS561E0xlVbP5A8n8XrnNvGepo1srlc42Wxc7u4fnS2hN3FSM3aV8oLUQUHzwzdqvh
ljB8uPIT5vUK1Wv+WDiT9dDQvfkjDGi2IDWlKnMlDeyvk+lhUjfdX6/CiA5G0HsgNLAt2sbQNRGH
Vo56TtHfENUQskSh+4ILU9nGXGaq5DxhD8klUR4q3bnGm4BUowr883Eph9eBZRxwu52QChN62iQp
WGKPTm9dqAY4QuiPtzeae8BBecp+iEIXZ1vNRRPUHe4yWnrfvUmhs40Ixkuj/AqeQj3/hyT/rBgp
y0wp6+XxPV82oeOfy0lpnMogMmUHkl6zjvsj6TGUOAqvyMYt1rYpDZbs/GjnLPjWDTrIIdZyb5VP
5D0gMZyYPklsgN+bCFNzcwg7laIFSilQO+niUgKHlScCgxEPsY/Imze7e/8VBI1cHYOYBS8ekMer
GsxxzdtGUs2JgazJbPagfqDEZM+7MvCMGQJE/3IMUBFPL/MPKw34qWtfV7n8Iv6s6dPjaZlunjzG
SP1D5tQYzmPczrm1RPopBjozI0nTNel9cpT288dLg7yvmq+vF09/iPbsnRuVwKenwLUOjSRZu5o5
Z6P5HMlGbpbgrr6F+mIxd60Qc28V7bDRr/ee7zYkp4ibJKjsCI1/4SpPf+ZiCaERJO1yc9zUCpoD
lVuaT5fG7rQOVTkEMkO1xgVaZsMhjlrbx/ba1v8PFOPeXHEPJBMYfyIAKXIosgd4CbE2mjQlT7OG
M7qzMJ0qVGt+QPSuk0DIkrFfq7f5cEXrSFgg+p1bqQR0KG+MG1F1SzgLnR+0/vWyALaZ950EWcwO
9ky6VQE5T2Qndt8FtfMPkPQXab/4L46ZRfdNU6jpJ/Q8mEsOrWiM2GqamuGzeOLvkhpTUc6BcKCq
+4JinAdtpHvL4Xrguo1CF3cHIy3MurVrzG+h14R+jYlw7cx3JHJTnZIGB0prB7de5NEC3bh9EQJP
yoO/TGZ3nZchMIpxxDhqyPYziiTZndJ9bXni2rUjSA2WZS38VovlDjuK2wyog1wvBmzVipk+F6T6
rzTONc7rvDQi5ogqTUPSiqbXlnuFUzbDiKJP2g1WoaMhEqmmFuN0z/6V1CAK1lubEm5+fG4WovLP
4UcpCPX1hkbdPPE6i8q4JN/undeQfELY5XgAD/RWl8GhbvPZYT3so3N+U7ZtA//jU2dbpX7QJVQ5
GjPOxei08jMEP7PBNAx+JkrurWytnA+v97Ayze/18CWa85jfruKtvqqw6NMBrGe2nEMj5RLgeRVe
gT3Qpfk+XJutAXAoqpiqCLuzcH5F+9t3twLj1MMgyOP5scwvW1V3yxiu/gV/ZDuSYY98RPJKPohK
D4rpH46iP+hSNb1fHEDNxJAlAVJvdqpCe5AhkOgDMNyGAaDyhbJzjySNnI0r/iF0D5bm7Q5IY5/h
Lv2fHqh5zbdMJFdDJLOe9y9J1Mx1zlTtPw7I4QDuwhERYiYdm02ZN1jeN+yBOEkN8rRVplmhS32f
je6n/3goKI3+Su2/WmWf5TQXdXOfPzB2LlhKbkO9kFYakMLPva6l0DdlrEqJJXZb9J9F+y2Y8gC6
bvD3rUpV+aO1UHbH5SorwhdmOkMm2pI+oVdlVjOeRRSwJeNlc866vlz2VJ9JS9oreHOfXKt7ObhX
TFWE85ewZkjc4ukbqoaU66MCGiioFfpN+2Vy06Sqv7jZj+0AyHjnTSlzwPct7/ccoyIECNIdfuTJ
DFykMgalPOrvlPbMHZVN/340F2dCpFxgq/qX3nYRR+yE+vcvkF/qk+cJCWg5ol8VC9rYJCzV5m92
sfXhBG5MzuPdbI/GHWIhPWQDuZBQz15ZXq3z2Cy0wqTnaml5xnAfa8aZFiVDK279leYbp3Dka3cT
t5C6BvLKvajnH4snp89JH75M0mlNDztmGAwIVzqWN+56sExyKkj8hxEiqZMItFqqqndFaTC3ukkx
Sbp3EMv6PmZxpl2PabczDGTu7ohpLC+/blssX8G+qhYbJ+Y7MtN4l/LkzRlPgs3iblBaQ+5egI42
b46QNtL+fTUSQo/xrkkBkeVQ6JVY1RPGTvIPzboEN30Vn8OfbeJJjrWMkhyCk7lPwpXyZYeLpAA7
wAroG7USl/MFDv5r6nwqbiAlNOQapY6umT6xI6CVSjP7FduBXkAcep9WU68XG6XScJD+GijYAlGL
o65irGlPa/reyplYknYkXwR8eW2I/uV8Wph1PqL6g/oaU1ltEUmOzdAEMQenPIweVZ3d8yb8lSsI
Tka/DK9q1cCzLzUlnZqcqK2GxORvZKgFZd/WD3iAz6miOT3Oilg0JeOYX6uMmMImFfWH2YkfHIZi
NsbunDZrHYV9pIhRunY7Yc9nr+VkICfmIyo4hGDh6zYf9KJc4diaWoAx4xZR06iqWkL2KMr0kEOg
SK3aRlPFWTns8S03Kk6jYzy49KaAthkkSQBd/hJwxMY8LP+BprTl8LPNIwrCmz9OI8dqBwmynQvo
Y7JGOilXampGidt6jXp20kTGK90cJINs2PRp8k7bJJvoVRPUaQSykJOP6Ep8jv5fDweSBRLknQvU
cDXvrt02Jfh+HGIB5KPlwkyQs9Pd7Z0WIDz8tT8dDX6GqOEVH6OTUmCDwcLYEvo13WM/e4zF1SzK
ei+BqumBmd8R16MuInEtmNpcUHXJbl+GDrw7rottAVty+fVtGJh+C91kAbAgNi3k2s3pb2DnOVTh
+YLeFHu751UYxc6df5YIILMbHG4Hq/xvNyEE5QINsk/y0ymroQWQvqSG/9UdWHEKBZUZ6g8Zrr91
9oCXMFrURfFUnx7ux+/1P8OcWojP3jCKPpGUfydCtglDG3/wptfnRpUvZiHKHcQzdJr6Mv3MQzcp
b69+NqY47hd4Ouk+K/LoHrwWmLlGM7QuBPXnl9fPXyPmXwy8waGNKuySNkZdwviYcJOO8+romzau
vm4b2jQIsXMaVH+OVa/KsZHJIANwyVJD6foEwsFbJlJVFsTDn1JCidFeWGd8E7tEWir9vdxcB+sI
RlPWkDieWHVkaq9eEo2tECHaywCTAaioS0dVzdP1r0LcI1cjpz5hIMsd/MZjIV+CNDC+JG1vKz0g
y4+Wf/zi1XM5uLAXq6YZaADYHv1JFSC2a7qWBp1SnCAprbfjcp2O0EuXL78kNsZK+JcIsktpgsMJ
CoV35yMe1NukGEGDQmh7WUxn5dVJvNSEpIF8YqCp/e7yRxnuQqynNa6Cc7vJAdzulmB2/hQyllYz
YbdFwzMOYyzPAE+3zVWw1XMufDaaOmSkx0xHch+I03pu5oo5Ble79hMl8bDJATHc9JQw0sUN4KL/
ZIB4zPDehaPAdoWA+n7VNquOI9A+dy/xIhML52W9w67KyI5wy+x38yWlzc+pUK97oPcoAt8DaYBt
YUjQEIibMmd0pA14Fo2Z3AKMJWbFxJXwoknyY7mB+knhCokl4lgAq3DiPJYoku9J7tKSFzwfbXsn
AXsomu4df1nqebRU5hnlYHx3im+ynYuHZwUxry4zyIUNPAaudIWeJfNfPSOMPMgi80/lL5PKKggV
B65FHBrAPHVBpOxtGBGWNMUty4D1/JnvOZvBvkdn4JbjPXz8L5MXDiPNeu+7ewduZ6vR71831kit
kk+lbXWGJtJWK82PcB6GKDqOzqDtcIiAUgzex2Rhio1UZdhGWqBs9S/Xa26B3yHl3e7a3GrIJKHz
Dh9G8t4M4T+BACT3FRsx96c/Y+a4wicxgoXIuIwNNYL1UirScRSfBAqLIhQymuP8ibMOjJxt49YI
QxxMpqxqZVwXEbPIhubbz9U/pE7puBt60Am6H5418Z/TZJ46aFwvecyMOT/gOYNq48lYjyEn9HKs
vvivqR/MC8VurZRtR8xFX+k0FCz93hPiwuxYIsaD4ywJo301I7q7JCoe+2OnI6lvBh7HRr4dC65q
gIiC4tWtKDGBHIg4NN8B7tPrY3efDXIXsI8xa101K+KQC3eOGj9FRSoh5EKn0Oiizhu7cBBbsT6C
Uq4ckP8GP9wmogyZEog5/uh1pLzliJQ6V6iGZSFv5+mgbhsmJ8GugxPS1qZ5gzvPg2RhHWchrQCR
JEOJ6DiZs08fJSerMq+s40wMd6nX0/FvWJ7y+QWthSWHfL91xjVVvodJiVvdCl8hnCaC1v1rtfvL
pEVojGmws+d8hmgvb5R/KLq8MTvx4ekA6wn212JBDQETEPXq5jAMjviXSWJgWlv7mfPikmh6OVBR
da9JpNhZt3QEYmi4Eey11O1CM8AMStuI3HyRSwsF6wxWXYjsTrDGOtH/a1oa3Af5IKLZ43rWugKN
HHt9lyuuRiMRIcQ9WPrsYfMKRlXqdZwTEGUf06UDtryPn7J9wEswYvZFwtl15ZN00WIxgyppKy+E
teNZiz/irxNsEkLBGxHo0yUkTL/w+Rbu5IAa8qfcbQ495aiA3BXfXj5G+d75o1dK4Q9l/4P82m25
DjkJ6/z6CtZlWUPeXcAtDIdyqSyQuKjCJP8iyEjohrDQ7Ysxo7rm0u3WLMvE2Gv6nQgwB7EQPGbV
vlFePD6GZvhwGfRqZ0soj9hv9xoYjHICFBPamfrAJAwLmavKNHTxFayFek0fZftrCvAJ2RhxK80I
zNSG776A5nCzz9bJ0aEUvZ5OUg7tQMzPeCAhV6sWH0NoTdWpl0UWY5oOD4yxzt5uG/SSXMbsw0nP
k+QI7sWZ2VJQCmzEF9iVG/wMoecA7aGTDYCgEE4WCYfMUVdgWQcuqh0zHFEa4TG/IP6pQRwGT2aF
LcFbFxYz9ZoH7jAEd0ZSgri6IvAcEl9P9S92jwYVzAaytFi+21CAMUXMT1uvKWVQJNh9oe1kYH0W
XzxZaw98Lcb4DtGECRvQciTkKh2pb9VzIDXDYSPcKykjJAISdxIW0We5c+Qg0ivV+E6Da8sabWdC
6ticz/X2vq9LtRcbnbcRrx5vgOrHDTZF5YKMPY0f7VSq0yaD3ZjRZT/HdEnv2ne6nFl3gisvww1j
vF94VWdssLqEuJMR8nOo1Uul314qiV1wLAm08Z26DfD5JQq2KAKwBMjEEiK88s4TJ5uXIrrY+glp
ia9Vjgz+1/230S+M4ZEM+V2BXqbdwkttRNp9zz3yurPADeBzHu6XxMBUkR8724CYhoVmfi6kQasG
aBQ5exxcY7Db8la2PM1YwdEIHWA+6Cgfpig7OjUyZAYIjIOUqlUrXMfcRkkhmGrkC8Re12U1fMxN
WSMZAsiSsrWuOpg42sr9c2U2yhkjVm2OaFtBOYWxRAivxLiWXfz3JZjYZbhwVL6EVzg8VDDd2SKG
hG6TxN2bkbZS4L6qEtqUMPm+zCfzSjJzE6C9xM8e/w9dlbT0iamX9s0K7DmkZc7CBSz4e8XnQ8ES
Dpokyb2fO0qwOiH4ZweVeefyq6SKp6e3nngczvNshuwuFBpJVakd1vAV6nl7TsZM6jRDnFOyS2Bd
ixAYflAteynZJWiSqJr3mWKsYeOGZi3bjExkvTLGUhoa9VqC3xZs6wpozYJflV3IGc9PzlEazf0I
d0B22ryZ59/1YWPfYUK24gyvkr+E2ZUMZMG3ECBFpo+d0s/wYDGR1Eav/ZaQ7FvGxRwmpR1Qf+ns
GCbvmVkPXhq/f0Qkk137XiRh2sA8QmWfUzj0jKhYBbcrKob7Frqbi3PqXgPVIwVp28fepj24IK21
zE5+5lgFH4koOf2Lot5XE20XFJ1LLz+ThpM1k5BnAB70i9GqQ79mxeq0AjQpt4vd0J7B6OinujDE
s2xn34MQaoEp7oCisg+Ap06UWZYGtRwhAUMuvpXaRyv1N48pOJ66YlRr17Liczq0HmN27QLgXrcm
g30qXhnUPqrW5vt0wSOs9KGdE1ZuMuY+WjQGgcCeZTmi+XJ4XISyZ4cjnPMOpPE+7sVS9JdClpaA
2PgRyB1yLRtBC0CCq0y8Ob8w8wljfVx83Mokbc23Jv8tGFdkrB554imqSDxF4bXA0JcN88azWsGi
I9YEkMVdUrcRcjtDxK+FCNaxXoGm6ND3HejcJrs2fY0Que3uBoF6HjswNm/qeSyvHI486tPwcycr
YI+hAlgSzf8e6oyrgz2BE/BS71da7gD1NwDHCK9kK6OyNtqQwQp4yQ9UaosETDd7YEnnkStzv7yG
wpxy0gmKGuSEkFOi+//uHS2bLiLrex0Ijw8k2gNjuGCe8vwTj6Gp/Tk3jL1UyTXqdru3nGm1HESc
eAkNsNw7SywVptpnh7N6KR2qwzn9iS0pJznvIkHJHcH53Wzxm2NN+koYB1Yr2Kcy64DIHidaRdJ8
BcX45GfKI0Rgh7EJxF78jO/G2zuUbyk6ifJykLNwiyrCEzHXrDg8SL33yviq7jly2hKLzVJtSu6T
dYF2GoUMcHnOrdiSwkQT5oHrKbsoTMGIVzhx2zblz+Y9/QN4BqFRI2TnhRhCeRZXPgh/okwTYZgt
qDbxLxxeQbG0iLThGeaHqoMBKR28ob+oUfvqezySR43IGr7TctTIAI6Le0JZoODF82ZQF6ysP34U
YpMfAW2UidSTNUKRt9TI8uGsVA34kNay1W4V5iGGp1begUFUmWhGOqD0/TZC/y/NRzh4+S2If8E6
qyFPdxiIFoA1npDrCO0Waw6i/iPr9RO/pvjKBbV/BPBtx7E+OiZwW1S8RQ4tY0EfDPAVc8y6rWy2
PkvMT0ESsjqj11lpH7U150x/v9hKIicFvc/fbeEkHYfrZVNE+pJSf4AF0vqjLEtCZ3YbKaJJvHl2
NJKb34b93t2ctySkiuqKZa1cgUMcz6R3VP/eQOZ8O9ILyiY1XF2i3IeFsIRBd7LDG15iXaANPT41
efVurULCXrXpq9vPl5Q+k4l3HiQEfwidxAzDfQOWKZ7VgEplOrT/AiofHCmeey4zj4iapb5FfX69
sG75vDjlyNwbDGa53BcNUr5N2SknaXmLOVIfERcApkPZ86iAHhABawDGk+4N553BEagxsjBPoJKI
5r6SaZIgOtjndGQYPEkpbn4G6/nN3RtR2xLrbyMgQqVil1Zph7B56s3vN80Kz07N+/rgdDel2Nwo
lOP5UBf2ELKDnjWwrJLpKc+eOyVx5tuPHR9Gb7+4kAVgeDw/qU4BkPD+KqwYhgujlG2QArVpdxdq
UqB78rQZxTbbyVXvruy3y9FFIij7YSX/6bg1nk5iD+/6Si92oyGGbIWSSfYBBrPKWhbjA9Ae5smP
alGzfVf7mzU9O3A3mCc7xw+Hzz3ErP73UEaFRV8KG6MiwSH1mpDaxcEGgO8ID9vPlHDNqHq3tD43
zXYlFwG5m/5ltcyj/lWDIASARlc2RDJvV0yOIkdBfQXU+giodIgAXB0tVZmVy5PYHqVmSBDp3JbV
w5japiXFd2z5/Mtexlz9n/kuUhrTwOFMtzzZAcEEtKuFgfYKVmke3uFozpkVUEW24dnT0jrHzS8N
BEg7CM58MxowvPABtiZSJJYzrqx6CtyWWDNMrgBmw8MitZkK29JUSTfgCLi1x3fbRxVrZxH9KgDW
otHWfSKDVNIiB2Cfn+siZsIJSgnshGPsAEGVyEMNfyejUPvO3g==
`protect end_protected
