XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=&���3С�ťif����͊�lӊ���e�H��=�Α�@MS@�������%�=�PT��F�̫/�����d����po�T=+��0w|�'u����UH'w��-���Nh�>2Nf�Nz/�̽�l_F�ܒ��:Ϝ���t�Й�x��:1}�Ⱦ�5w(8j�ۍ��)�?5�.oRC�Z�߾��5;�v	I�L�� �֪��k k ���k?���*�P�i�Y��U����R��s�V�1`r����ޜ��Ć���֓�]�
x�sDAn��9���w�k��m~:G��qoە�s��f�Y�a>)�ъ�������y������b5�5�vX\�R�({t�꘯^��9!F�V�>��К�H (���`��Ͼ�w�}>/�m���nȸ�yn�"+��L�*� �x���Y'P�R<�HR}I-H����w>�S�Y-���Զ����[�p��O��d"�
~6/�����N�k�=��o@fPʋ�N9?Nd�����ٞD�����:�5���O��A|KTu���}�:2�:�s
��dP:�L��6a\��ί�l��� Xu�� 	�UB�I����U_�No���L��ܫEr�:�}0e��5��=2�|��˗l�z�3��!O��E�(^`�%�R,%�T�U�m�x�d�~�Ȍ~Bm,�O8\3���Q�z�o�Z}�!�R��t4��a!����ad.��A�`ﷆr8��B��0m�r��zz3�ݣ�
^���x3bHl�(��XlxVHYEB     400     1d0g�����q�e]Q�������Z��Ճ�۷�=L�k��`�`�sз��eq�C��d����[6N�ӯ�l��=���눳�S9*d�(\1`��l�ȗp��[	>��e7�	F�UGg�1唥��� ��L�iZp u%�?��O�bЃvY5s�C{�}_���A�"(�����=)�#>������dYp���f1�d0��4��~��0=�-Q��>H�Yw#�T^E��̖�O��DI����.������e"�px#�u��4.� ylQ'�9v*�����nAE)ՔD����� [����`$�z럊���<�����1�}�P�4V�[�Ҥk?�UZ3��!����������	�(��v�;�*�'ZT@ZU�W���m疘-�hV��ȧ�|�2�Е��z���C�_%5̛��7�K��}��dL���������E�0fk�ae�XlxVHYEB     400     1304���^��>�w����]5������&���n�*��T|9�V�1�z��E�٘XY�[ӹ�s�O��Q�Sz�yVC�w|Z#�{�y��m�f��6]��PiI7V q�B{
D���ca�[��x�x!�E����Ѷ���J�)�,�|�Sg���9~,��T�����U^�7|~��\�^Dę:�a��Uf��'�x+L�f�����{����rۻ�i��(���қmuoy2t<�Z(��kMo���♛e�^P�ڋ����X�Ï$E�Zkf���@HZ��Sr'"�}����"�hXlxVHYEB     121      90�\}���D�>K�S����:�1U��HY��}�#q�9
��Tzh�������	!3xNB�2ǁt�V��b�2l]8�?��F߲aZ�A�ꗱ�L�[A�[Y=������K�0B��ї�ѷ����[�b7�����:��,7�w�