`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69168)
`protect data_block
0USWSUGxovGsyBJteYpEoa+uZS0xhIrRdED5syosToVbIcMvx834OaTrFby0EpL42KTILaX49Yxl
bvhohfseTX4qERDtwqzKWN5aB7AAKbsIlIaS6GtXsfjJoBWZYF9a6csbqmu35Sre0WaTfw+9KA9W
31TbmjPTFuAQKWuv6zvtrjH+dYhAH5kJMc2BKNFvAUvEinH6yNY040QiWmeeOiLHwJlX32Tel6gh
XXWgWWLCBDvW2J/A6no8TkrOA1tLAUtntmOaZTSBuK7yAqYDCO5vAG9B0pY5EzjyKNpB1WYYvR9U
HpGwyLvYGXt21uhhlepH+wbXBZnQYyyIFeG13srRGz6MS0yd1tBuXkcfAggxrmQvHAznm/nCKcw+
JR8FnU61KfAfAzvAhxxI8TSa3O6EB18HyDL6545uOKSW7gcgXNw8J2M2HfE6pzx4jz1zeVqw630D
rUuVnAOAmrZCNw96L1z/YyL1SoiVG2djyb2Va5TPOahTJojBi2Wg1sxaikNYDydn/92QzG+uXAh/
jggG8b7yHpM2g5dxq4hiOk5UMcNeiQgaWOjhPgCgsLrvDCzuCHHBnpfaf4SCTehOTgHqCxPwenOE
ZM4pLbbcTMrySSF1jdU28FBjtbpgmC6ZNBxWxvX8XZGq/ILc3I3nMsLTFiettXRWSsF3MtFaXQvh
8/weez2zDXdebIyox5Oo7Fz9Bw4F40xIGioDjIKc8Db7aO8WpaHP6P2G61ppM8SsDaHsypac7sZs
XFAkHVhq+SLuGzxDxJcCKiUnkVQbNOWgNvnfVzDRqf8Pz1UReBUJLDRxoIjRAf6ROcHhAFYaSHKM
88/DW1usbGS1cgko4i9VBsE39gBh195xICxxZy0HPDa5HUwkyC+7u6980jvsOv0Zr6m9URXIeUlY
73BCuiLTlVqr5ipz7vw/rmvzZeSJazW/f1UID0ZStz4bngJ2w/wguOuCMST5N6AagUzM5eVRII3i
eYHQKhbHsS2N5TPuC8y6babk5+szC9eBuv7VnR1rfzT3Ft9pcJIPAPVBJegq0Yj/sHF7mcPHrg3C
J/QDVBOLPRiYY3X50ET0n22nhqYAiDn8F4qR3sMoXE1D3dX1Xr3xYbdu3gWOMYL2oJar0i+xsZ1o
3QZ4S9EeiHYiLOJiFmRHO7+W0X/MjTtOTqs0+vqSE0LUlTw0wsrkA3a3v9oTbC+HZpy/BUHM9dQS
7dX2k+nU4tuZz3jHQWga8YDK28Ltw1FIDDdExndh4Tsrb9Jqw3iC2TU12nyG/WkrviELXGP51jfc
M6WYJR7xZ/M/zx9E2VwBBNrpVivJpGyJd534Hh60/8Yr24HKXUQcF959HqkU4ud7sxUVuvAbufDl
GzF5gpJ7YaoQnULSyAhThYQ+KivVuFtjRLn4MdB/8dLkHlUadao16BNn80JG6YzR4VnyX5t1Yj38
73YvhI+qSnNj+Ll7cD1Fj3Ylvv0kO7n/FWaEz6hF4E+bGA+L/ENN8GQq5C1BmXnVSPANw0Kl/QfF
HEPuFtxW5iXHYWY1epOT/snfLCJM1nk966bea5wcgN4VKiELhd295TWd8irZaeI4mVEksEv5EPkU
mJngXVi1uIAgyt7CLrF8MAgB8hZoDmAF7TJACRJyxinrIdp90VNt1Lf1WmpRlaDHx6wxeSCXkAwc
2I1FkHMPBgeesUC1gff8JgDIrNielhTfn8wqTcVNPMDw1VkFujPLWD9ohI4BXi59LlWImL/TbvvP
Rcjkgs4+1T8e3QvEXFXsV32PqeUbznC/cXMklhXo8+maGQKmiEan285c9mkKzk/txmN5gpYuub3B
T3YX1WwYZ9spj7otGjV8gGxP1qI2rckoBi8znA37sVLGpdg9IsjBma2Catj7lzNW63CEXGMRCpHn
fgAIdrDphysBezKoa89UQakpQXun2GO1bdVTIdreaAZvGVU2d2yUa7ZyliKVMNyi/Py0yuI5nzPL
1swHMbK5xinN+9C9K6GppZs/OwRSt01kd4lMrfbBEmcW+FxaNVlz+8DAX6xP6AAvUeV3GW8noPO5
Wmuek4dne4c2ztRDtYM69piUAe1obS3oJiK9i6Tdx3HpxP1GFxAMpfmFN93dOzwZVhFjRUSj1ohP
nO2A1eQpQ4duz9HX1ACCuQ8A5lpEdtUTu5svlEGXb1r2dhfCTomq5yWdIUNQ22jiW4acKRH9rXwX
6x+Wm5v+vpEGJVw80msrSyQ5tvoRugmqx8nhmg6hZYiYfG1kD9OX4lZZw3z1J6/rErRhffnMHed7
JBOGslSdwEbqmta5ElrHuRiyUpRkPS8PPaBJMMq5CKDY0TKEvQJnh/u418YgezCnnxnoRv6XqFb7
8uSC/CvqfWCkSTtGbFg1OwJjlWMZ4ehNYWXDJoFWyuYS7JFtMIexy2zYrR5YMTHXClyn3s6OSBNN
cS/1fQ3ca4X8+sJCerWm/KUpUxeXh7AMTjsdfi5s+XkrMqyDqFqaO9ZiyeIDf7QeNNU2hXSjrHsR
8aeq0yzmMpOcGk2s5xGrynRz181DcO76WdCurwte+mTxD5q6Mtwe0LHt2fcJ7iTf0keGohnDoEbk
Y/VPTweIaRm3yRHk9TVDErUe5v8hfqMSEnHNS5HhJyltUdxScGVEkM3eGn6lFO93Y3kQBWQxbjN8
I0R2k+Rbt3NFI2qd02bZ/6FKnQA4lFI6MNyFugmQ88nlGPmNkYq0opLQmepFAkH0j9oMEwhK0bWL
ymXfcyPYlxzAx4BZIP4CLLNbP5MdOjhs+lIE4nwQD+pppPrCrSq8upP1sJN15q8tMnBwk/sMUibR
Q0h6Iu7fkQRKmtzcYi10j0nfTFYWZqDqOMfJtivnW36p3TOQu6/VAUBTKlSlC1q0KHVZAuejTbW/
UOrw4dFqlaB/XOm3wYGFpUEa+PuuBSFJVl82BRS6OI3IFST0Kwnee3NcdF0L1l+24OC9C3FmhM1A
kPIwW41fANiVjA3FWdzeqJXGk3WhtKETNQEaRg4pgYieFSWS+M4SbLjcSnQRTyg4aKFtHkmfapNo
osDDT+HOZNRiuf+Wc92iyVcXLwxDIc8gVi2W5FxNs5J21Ov1ngCtgBHf9sd2OENdifwnzirzVA6w
0upHTgfZ8Z2t5RCFUrt5bvHko7N17J87OVmjxHja+gJ56QUydtD/qA/wQw9XLfkiHrzglqfxqkO+
P/w4BxeExhdJxtK4aSKlqxoFEKf6vWcdoOb2wLZCLCo2w3cZm35VExwGVSuZUiWaqUqA4Rnk6UGn
NhsdawiTU+TAEUNjV358D5OY6r5DspTDabSyYqupRrG+ucam9JKlAe1lf2dkVRdwXEnypaDcUPJr
KL7VkQbwuCshFbJa/8lZ4W7xr/DahILHgH0QnypKQP48SMmMuKF5xgWyGJzz7z+d9ZTcl1ALrHdi
2070lTiqeMzYt+f4P1ZDDA+blvq0O/JI3YZ7HqSaV9SPJflPd59jt9JTZucCzVFuoOU+oLr6vfP9
UWPk7SgO1+RgKon9snOmVUTPiWaUNHJazTzEDx5iZzpufYCWbgTpiipllzq0BDIzxd83vM8xCAL0
m+iS9/1/NlL+SvD+MMcpOJAyR0ky72XtTJOEpbDhZmrFyYGH+o+BTXcPXS61unAnBhcdkE3Q4iYH
v84iMaLVx1IqZCykISbfs60XJHmZIhY5pA4VhfgfG+OF8tl1dT/zcoOEC1RC+ApNpB3c4nukNMfV
BKIgIdJW4V+1ri9AIfPHxEdVK8uW776PbYj+rcB3sDd+KiRv+CWnybACvU69o2wJO2VF6yMFz4/Q
eKYfPRjShB06bBgdhZ8UQe1LOB5al4rV313xvZuJ6+klZBx5m+Wb3IrQoXeiTSEag83QzWZVrSXZ
5sxnR6NoLZPWeHvqmMDILWCrHYRdvNdJ0Eh7nR9tm55YXlMWaIqqXCWRFGPZJoOhC771m3kZO13A
jzmPSzXmzHy2U8IMKDGjRrrX2EUXYPU1v4KzOMZK15BGbD4iYbn+ubc+hA8HxiIxMaXF6sYvXFiR
r2L0Jvk9OiuDkJmTrMzv0DqWsPKQgCNrMmIYbsXaytYljmry+/+qD7HHil8aarFmSUqIlc86SEH5
bJMJqKIc1InUvG1doihLihGuQNjWX9nb8LmDThg0LET15dU8fL5wfU3KytEMDWGCPJc+78XwuWLY
2aI1sQhlxbU6Ml2b8gX0wqv1fZ6Jk3cYTtj3/DQWSdtfJErPOk56EfHFl8RCMcWKvI7Dvs0620+/
/NdFJS1U67QYUDC7Rkq+S1f3OtSWLKfQ0ZDkc7Fw/GqnFHX5Z9iAVMfctTbztLOHFcv+MK1dU8U/
6gTqyzW624DnpDBb2rUugXrtaWQoZdpBiaF2iLR1yunyFhVcrc+hnyu/Rest+5RDhYR7J19aMUoM
NidhbyTbvyMWEWSzsZ5OxK7UtP2arHn/jrLi4MQNN8ynL5AEXkJwQ/TQpki/nY064VdFVBwMYRUg
+J+Zr5OyctzS0CIHLWFnKeUdsWTtqjVHJ63plkWGGUVY70Zpa8gG3r6oiHUAoa6UTsZbSU5NW5BB
bmeUq4eBijEAMBMoi9KLcHwfutaYqbLwm2GUxrAXwrlA+GmUfysLD6UZcF4afhOJ8pDsuT2JgSHu
VQ5S3cHrVyPXKKe/WBwfQKU3ku+BRq6idXNxvz13UcBMJLjeyyghfXH/Lo0xQz44QRTsL9EXxdgy
UcUCuYj4aByygxsgCes6H1As51cq7sbi02m2/uqR3nJ4d8yuXPoXYwv9UtzU7fECufQRdaHqkLoC
teqFnYYeL3D614lJUYRF3xTy5dYPZPT3ZUTNxv0ZOzHJOl6TfmE5EM29VV/sYgXnsnbqVqyMzsAI
a/7U7XjdvYy9RJ61ihufyHtpjx768EP0+PW9nLOJ2mG2qPbOQRboDHy5FaCRtnY2zOtyj1UJj4fU
OGgOFReVGxymSbTYPdSOGwNUVTqNI6X9xlrlT3ObjSWnhsn7/GEbJP1E81fYwSnXH6XYS/+h3UNh
6qjbY1sEmb8/HcTTwLYHlzbrY45z1qbxSGUfRUAj4E1y/KqBvdVNTnoOW1beQIYBNO7G0BI+utE4
czWaMsd/7YBzWQjuyG2Eub/Z2n+UDwFwdkg6w8znERiH7h5IxxUTWk9VTnmTUK+ktlKPrE8pl4dN
z8C2IvI5DE31uJ8yglldoDUPHVNxRkMnplzZmJiuxBbOjG+97pmiJKxicY13F52oX1iPMx/VBpfN
KDk2bC69NZepu4129FJfyor48MuGyes3NjTBqlCNxneXOBqehLvEEU+Vkf1wxmWmRoMmVhDEjme/
xFGv9efrHbodrjzL2ofnwB/d5QFSh5sCJIa1tzUWRhYMsEbDlLWTkp6oVB08yPaLfMQdgKIuM0ZD
x1ytDcJA15l2mZdm3GWb0eHmHur59RiAzLEOYIZZuOFXkipbBMqruf+NVaNeaOvnqI993k4FCulw
/G7Rco5Nn7FVmME5lQ6C1myfwBfiHGCZdPL+Gn9nsgONCLlssxRY/Zb8HoeCKBzMGshtntnQ7ZqK
GG0JVPXP0jooDvG1gZYfv/kivVzutYdxhaBkLPdTc9at6+pB+Nn7GOBXMFFrQHnC6p21QYhuKN2e
qaDhKPIv+bIvvOQVWHRSqZ1ffpJ7Ym+NWz1iYrKnIuXMXxIAcuLfqhS0J4wegHG/pdCJIljsqvTQ
alHYOLP/Eoy96X04o0tV3jpP0SicNIkjVJXeeum9oWdwzsbxLB+F97sDERJNhcfyhdyW9EGn6mWN
jJtiDC2363vAmCqtHx1NhclM+RolWtsfyVIf8ZgefESuFuEkYuwqj6CGkvzOrbg0TL8t/ODNtDXV
L7tKmPeNWbgzHxm7/9/kLEvtvrFozQ90Se2EYOtYKoLHQFCoYnTyqTTWaE7OL50WEV+UDR3NrQdk
2addfyyFGO3oy5dKrQzd5z9r7zuppX2end+D/AdiDO/XGTOr+ubWWWQ5JYN2DrLQu0LfdaKzWpz/
TPEHhRWj6TfP3hwcBFV1EBGyTQ12LKx5VvAWnUvKIqG3NYcKyHqzmbZavMXxyiosPQMSkm5C7lx1
jXtkyJcGzzL/9VNcDOYYoD9B7Xky6ZrRRyovEwV+GV2N0UZxrED0fvIKVQ5yyAhdgEYeKF2HIt3W
H3caONjbJxuRRlXQpkxBUvcSsyDY/FysAvhP5jegllOhioASgiiCwMzSRcE0Jyo7ec0IUAo3YdBV
4JbCNXyZBnIPVMHsIXUsrcTwLV8QQF3FYZBsSnFNKOeGjQ75g5vT6C2b1BeQMDjCrMDdqUm/CCIy
rfPLospOBXrRN868wYjdHaBhX3/ALIblEr9bEokmb64kcN+ve9S4zVNspTSqdMe0p1cYPjfX8gf3
YCqsyewkTcJ8mzRN+ulCOUP1574Iq9o2b3pDxH1yxEx/3UJsXzCS4n1eVC0wVJuUFhGtVTfGwBhj
GSXwjQGDTr8ZD5FDQz374tBKsXhV71ITrfTzXPynDsqHQvsUlN1QpeH2swxl3umK/JYrtHTNRNv4
mfF9Clw6Vq+GcW8fo9n2aLeeJyYxxZ4q8+Jd6FZp53AcPWAPZwsgLbJzX5QVj2fNgWQcos7Xn+ZK
d7C4gUQs9MAPAfwN67/nK9AZrrK0ugY3IpEX+ZWxQ65WFK/2dcNbmBsuLrNuF7NZF2hZj9fqs3At
IvWHpw+/wL5REKuffxw1CdcfoNRuTBgQgrPd8Ir3xpcq4zJG7mZt7Cef0SaOTkXWfQ6+7ivtXLPl
faCf9rY4Zp2jwkbQ+dFHnVjNbWTSuyC1f97ksJ7DnGoWfUxzxCrIV6j00kXuw/fqLPEuqJ7eVgXV
NGeXzHZNjy9vJLDuO0lnWFSFwu47cs3LGdvEZP2GPLEga4jw9srC8jhm9IQt8Xts/48/2tmvPh9L
4ExV3MCYndCOEawlADsNqo3Vo78di1VXa2goyS1dAWk9CY4N5JwdnL1hY6fPJUeojZUCfWhbKPff
Qk864doMNAM4o3Z5/Uxq+RqKEt/XrkdGxxhh2V9ah9XrR7/17sSXZXGGqfvEx5o9pMqQSj4JtxFw
zFOyKXswbloHc0FCKmiPL2dOVSscZsozEzW0TfxgT5P47yA/WQeRnwHqNsRhNfXaTRrw57jhOhLC
YCpQ9VP8m73Wpqul3FelLIKkvfzA1OpB4l7aQLYuZRnWyZ/kcEH54/HXzxK1b06WAStM/25uRp4x
2mGLTB9Xuiz0Kg1zFIShFw1oUL8jxDb31Ko5AOFsRwsTXXMjWz0SJdhN9c3muSt517RhxN19XFyf
iHt395xpW1qcZ6gbkmmdpsh0iDbxaE3n0AwoBSpkbfRPNCxoUoZpp+Pqn/B9sHfSfsBQw+Qo1+15
pPsT63b/fRKTLLrVq5ObpAk2FQane+SMvEn7cuUatEYRm7YQayEBtbmb3oh7uhFQ/gsUAa0+GIaW
YD+hrq/ZFlcmnY9nhfl/RM77Nys3Ywhtl8D80sNvLwDkq7ELW/SRUUAiz3A01g3t78lgEGnorqr4
sUF4Rapps3Mt+9y8b+eC/iDCOZWogpR1juO0YtCs3ylv/XfncQ86W3Xy0POURGWQA1nLT7VScMa1
Iy2oznIwmo+gwYjrgXeXknWdNC64TgYHjg1dWirU1RfLa6l84pjUUQC9n2KJ4ez9WcM3xS201OkK
PpF3QoxhIcTechoOz8YMvnOm2/ESnuMFIToK1SFggJBW3wMKIQOpCx+gP/MAFZsjKNiNfGddPjbS
dDiqxuSqSmMVBS5s22ZfHVUycYCnsk1n6NL4GxNTIKP8o1FxQC0IM+7IxaMTmxZ7hqoIl/mkmfz+
lEOu0TIWRj4G1S1SoxEQ8umLyTUU9Y9ZsFIJC5g6YSCcMSmZeRrPvsvW8gSFeWepTxv/TjdJlDks
Foqp50ztr95PJ6cBxZRfbgHKurYFqkaGNxUes16zxPnKM3Ah7BKrL3g54HwbOqGT8bSx4BCEM8iQ
QvVVylA3Z/zaIMhsPKrND97NhG4nVRT+sgnIwcPSpRXlg6NRHd65XULj7Ogp154oL+x8HYzVK6L8
fe2dYpcEDwjbbhLXRm3AbVAByphGBMnW0rtb0GQD48npPissK76p7rA0sOESXLWb1MLcTxI+ODm1
UqymQ1WiZJS1dC+BNrvSLjuJU4sYui1yZ1hPaupFgr0YChS+N4dtZr+FuJ+lZZhJn0O+UmU+OsI0
W5gIgDSBDYFd+9JVGoRraB2sa9oHEtXUkIloIvYJUVSUc6295c26aQ2D/UBmSzKr2nLL+Nshq1cI
VHp5Xu/28ds5s9fZBX9iLJXavexztEorgzCFIfTQlPzMfXiCvKjr2cyNT5oA5jQhlPa+lmq1NFnU
rJqhyUDim3OqfkaIn18E7+d2cTT7ShFrLLATuYn16xkKZRBB3sADLQ1OFgRJmRBf/E7yddA3r3Bb
ccdHZZogpzfDC0Z7nml9WwDbtt7JI1n4haE2C0BeSYBP/KAZBy8I28oLX4zxHDtNPfqwJ9kIHW5Y
IGZlhJbxIA3QyDJOd2P8k5RS4s5hFMHIVjApfKULeWOpj00/8C5Ihnwy9Q0kX7tWPHN+F9TpTF6b
hxWdk6XElgtpAGBzVLwLhJt8paByAIU0SnKI3PEIh7qH5uenePpREHTD/3HYG4gbvRRJO2rubW2x
ZYUqv5LMO302+0SsN4Bs1NEW+tR4InBcUc+7ihZnCor2ojCfgGVolQd4WBSU8BYFyCMVHuWFEQPz
S2ryYqz11oQB6O2hNzzU1rultvt5JnvEomZBksK5Ugr3yemgNPa4QR3mHNfpP4FZ8mFkwQdxIRDS
CJjcTU0RpFfEGAjcuTeWUDdKoj+yogc/DGkEq6ZcjIEEvwC0vkN0KczWHAL/l5Nu2WabMLCeVs/i
p42AyFjMjPICGiaQR54/6VSZClFJKHHXZEJF8OzO2kjECyvaijsxARkzcIrPObocp5N9Op5LYwft
w1gwvLWxYbh5330Mklv7GTyIE3zDzS3ozUlEav9tCmqyKggbFdLJTd5DDsdUyBpt7+gHzrXF5Lvw
QVHik65qq7pJL4b5xb9eIfXtV06teFdzf+ZUAuc8RNafWToVKdjBPqLCgXu4qfM9CwhlFYoombY2
5hwQw5ViIs8lDc/j8dP90MweSoHy3c0zsIRiDUtdNEpxzFzWyDmhohYnhxepfePw4p40ARG3fWPh
cViNZ/ViZ0PWmfqKNF4C95gppI1QgZexI2pvWBvRjpdyobP0poXot9p9nMx4UOkE11LXYLLXGXlP
CupaQc6Nv/CK938OuaRP1F0tnJGTeuBuUKuZWjqqbh7skTzCjo3Nb+tngR83HnBpUeFvC1NV6esG
aST+1Yf13NWUHzcYiaxFLzTQf3D/2/rc3zRkjf2dfNOL8EprzOH/7zdrLhXvG5AoRSFVI1lu+4JB
mVHqjvzSL0dC3KHom0EtTtm/uTIIWqP4v/0SBmAXnX0Ru/MsCWUpaPeRdMIPoUV3ItxmhJ7mfWOK
rx3K6YAJLJpAaZ/K0IRfsHM/0E5ov8935G5lcKIvnZFSs9F03aerxqxovu9JlTxhmkbUQnPrICw4
X3m2+jJo3J48yRUSDekKDoSYhawX2b4aJizbW3diEv0pA7J0Feoqtwm0OkJVH5iN6wSbTjD51jhI
L+s2sGZ5B1G/dNHtjGNbAXJ6M9qGZz7ZnlQUbSdz0AsGNN7AZIZBzUy0p41CVQobrMfBbdFJLGj5
3kilLt3MrCghJB8MnkBqz5Rh0zB05DWvxlsl8m8dbsuJOKwU2mkwJx/xIBlYT4s7LPt17s0HrEGt
18XmICGGHcHBPzk569y8yzd9cSSpweW8amtLhArP2/W5Mo+QS9B/sGt4gHJbP1geYgirhykeuBId
LohtAr/OaxE06638ZgeP+qqvBSPB/AT/oQMy5ml19etchAaUFT4d9dN821DtZC8qWiBK4f9+n/gP
0k3eAh+AVoHtEnFpqyYDJ804yHUOxJ7CPPzZpMt3QEj44m79MUxlCV8mH07uOYqO7IRFAa6JxBFq
kMoGac4TUr5AtbFFtytMnZB7ir/6k7a6rdeaGeJ2mQDynzlZtzCjB/JKY+fu7NkXNMYEaLOeDiHw
xo7W4n4yW9wEOtGfSRgODD3c5DzEE8tXZ6MeXFPK8lW4rIZbySUf9pUel1MHBqWaXwr6T7Y7XhDh
Oxl2n9s1jU9jPO6C2Jxf6WrYOIyGy3PL/Tx6To8GuTGybXpRQAY1p9ivK5EDJQznFocl/BbG95J9
zNQEWXsrLNrtbAXx7SykFS4eqIiiLyshoYIeME8sor/KPw8tvecsEaHLuLXAEy2CbBkKPn4OMDnD
Gfd7r2Ks8LGin/F3ovMjurN8AsnfIbbdDC+gvtG1uA1WY3y1mHE1F++cKnOpVHKD1u8UGP0XW3FF
XeWosH1jo8rrQO2Fg1WKBzkP3XQR1qL0TQ1FrfDWZ3FMZZ5xl+xtrUBQjLlcr37gbXpD2x10w2tS
b7NjkcQOvLdJnt5Pi2ZhXWFUuAKKbSu4XsbdykeoItTnbzOzJZ+fkhUmmT9sC5t7J5tzZMa8J9sv
Ytcb3sWgU/YK4WdltQdyZ30aDxD1CwrRTeQIfa4TBqDH87ptTKZ8Mh94GoMmt3+FuhHkDQEYDCr8
KaFV/YXC2qirXBw9GHJk3eraMPByEVjwaZIdkkqNVWFDPe/MTjIkxgS/Is3o3GZHaIFarSIFumrR
+dgsPTLTsCPiWXTzL1gCRjt7Vr5LyW0/JOJJTFsc0eXPcekbHQbMkf3qerojHOiqkaxzoBganGBI
UrHtDjn60RCehB5asfs1A5gk+SmJdyghqMfaUYW63DSK0wY3kyo/JdqXMbN38VT9WZ9i99r+oI+i
dXgW0UFb3Qsm28kpjrht+4v+nnbwiXYZRTEJ9tdqSV28LnczPxr9pG9OUbBm/8Y9hRpDgG/bKn85
Is2oOctXRC/jkH6GcxIUze+N/nu40r5OYuBX5x3N4ZvLq4VomZA2ojBxb3/5EZ6LNPTbVJkRYXyl
kVsue8bL/innK3pPq0jdVijJqLti+gFXUobiCP13QZZ8tTKOOelsUSepHE9gg6tk3pok5CvewH97
prWsPH5MihsSFldctIMQp6IAl9Ety4bFC0G5wQ5J8fdIpufcJ9JQGPlqPqWHuANnNbA5o8154qnE
ZRyybLWjZkLvRU9PuxJ2ihGauF/qQytp0oRjhKtYZmxuy63WVLCNZ1J/7MIvU2YGOOyvKv22BNN7
82d9b20MCPmet6PscQYVjVtCSmHT/PSxvZlR7gETUK4zkjbPyzFscwE1aL64PiWRh8czIZBzkkD4
czou+5duyqnyWTuv8vmeaIxhW9zOEgN8X8s8xJg65C+dRokazBQJO7Rxwx3wsDZKsCqghBswRGWQ
eVGrxkL0M+kPSXgAtAL+zSa8lm/lL996JFBn5jOrBcP/bqEYOmXxcytaZcF0nArGXHUZkhU9zo6h
7XLicm7F/OiFmBC0wLfn5s8ZuN6BXxD/3DoDjTjt5BgcR1/ARRj1+0/0ntU3xypVUm6sbUXoqiX9
IYRfXEqZWq/gFSdtdlep5mkqbNjONAV3aNpKOvdbMms6DA50TtKItAbc2adqeVKPzqL3CsGgaeNb
M5m9GfI68qjF2PvZvJinwHZTc+HPgGvJxRlO0qoj9bkaMR1rAfmOlGFRO6DiUFthc80nptYeada6
k6ztXArwEBluCrf0QE9zpwdPiBKSbQ71cb0iwG62JBVGGDNw+nG4S1YB5cq43xQKXAXCfikeiwwl
AvU63SMvTWATMwkuF7KV1eGHRZHQV72gohwZMtKK8plSBpIfIiMZ/x6n/jHdp2fBLCALpsvT3n0U
uwmhXTja0InQ07INqVA4HxmfQwXCQQLaOlMdBOHQ0G0bJRik9hg5s1XGeDxSyA92OkahIRoGc79i
zD2uGcMv6jzxgDMNu9OFH4/9WcYa2tVUdc4ryq6QhCL4LUuwVyvCchYf72lxhsBA0bJoslKW3EEM
s+/Way3clJRUy8RhC3rdCf9HrB4mS7JHd7KEB+nz0PiRa1hmYL89D4/ya/5qu8foHpY6DVwjq/E/
2eNedeKfwwLMzZyPc3BCTGCfhW2DlrRY7q3z8mF5xlzsdNqYNSqvJqWXdNnbb6UOyZG4ZGDMYIeQ
zieVeqdSWx1IIPxK/7oP37WTIgyxv75GIJRC76C64EqZ1PsOW62XGksGjZQ+j1lTxk/y0Yw7u9gr
HCKFDUr+UW2MhGawfE7yj8kMGpIzhPulMEjY5PAGUeLwOe2OFV0qiyAoQFf3JyVAq1prvjxKW83R
HoUNlO6y6nLcRUPF1MLm/lOdBQLzEQYEAy/CyPfIMKgl5OGEpwRdZkEA7pqQ5SlS7Zr3hMBnAf6W
rFOOpRpsfJ89GyaxJ6Ufv45h1cczW8bJ7x8GM7tlEuaWEb0iOccefcB6RUyd0MwyR1XJuD/IAXhL
v70+NuV8JBt7HtYrJmv6XE6rIEZz9H4JrzcTiv2WUjVdl8ehU9wFLAs36SY4bxcfik/PRimpsv0N
LtlKp6O5PSWwSlDg4WQPiUz9ZH2cBD0SPgx5yaAIiyoBRp5l2fkIQ+6t3mf6nHQ3mR4z3vTwfO9V
dielkapTOIHlm91oDqD9M7TsqwkfZzd0LD+eUKSMqJXKcO8hkrSa/6xtgr4VJb4eQi/vSAxs4Kr0
eqjJoUYof6HlBYO/VhsuRxjfwyut+bpoEUkeYuxpcjbGF0KzU2sL/LAdmPPx5Wp77dJskzz36iAu
pWTsu6NShJOnFoAPUq6NzrATKOGUiXphJW6BGzzqG0NmN5a2EIdYzO5IchSzvmdvuY4fgRR0uUdS
05CescVPLoWuBP94JtY3u7fe0Sj89FMgmXFBRRHhWSr3flzBNMmndU1R/qqICA1otO7jO0vOX+f8
e2Jp8TzeW4yPmOM/wugyvaFzRO6k0vtBOZL/FUJ6EOCu4NY1qFF1n5Uqt5JUMM74rVVGjWLNoRA0
ywUVHKdRZh/cCUApmQ+zW0eHdOcfMsgSRAiGFzw/pVXHjhcxqeoCNt5xvGpineq3Ck9O9hhcymz5
TaQaKLjfH0GUTb+O5MGWuMgHHunTJejwlVm/0XR9YVP07g/g9kCEQDBRCRkxr9IKM/JnJSbv8o6u
7GPqrf8qwopqOwhW5jCMluZ5Jc6SCFUE7eZZ+uk3bhvVwm9TKgpUbdVONq+TbduSxNw392lyLMEW
f2FY2EwaOjZ9rgOZmMvaJZMSoenzFGx6A1DoWh8BOl4f4qtutqwhotRVMGaF7miFcYSzpHhwxuZP
FcbD7on8sgcy2qb2P8HudtR5xBtEPy5LnU3uzz/LSbzi6Ko7Y4s1A73BBDUvfo/oDsMadxZax2c7
wSVr7vkYOSgMfAGkRe/R/L4YBFeo87ORb4kIl4yj9vQ/mqqmjkL5rLtRgJUY7+BMGVaPf+mF+0J9
tnabSXr5+9YfILSir6m1Wv71GXRbxSM2/gGaQMfUJ74SAsDQjQtNZClz49K68HseC8/5IJgAeoTu
at6taEi8xX12m2wnzRj4FOFb7Ytgg7OQYhqLApwSt1PXyj0kVLmkD9GDVXkTqQ6nZyvHAuMC/TuD
Wp7eZFwJvzw6oVR7U6ctjbRwYlmDAtgj0f4fL5cALKwymivf5gTzyCQiFdblvXzO3LRke7J641o/
8NKPonuDuRgTs1VjKBtnIzuCBWE9xbDTDUfi2gYgds5cY5bfRuaFeHZbmHQBbr6AYuyzp/YayaSc
rBEEnY280BUAhAAEbv4i/NMAXXnavRCL8463E9i3zOwSnSq1BSzi0kNzFT5CbfzCM0IonM/4AXqp
69w3QKaDkq69RQkQM40dBh3lEuW6SFp62lFarQHzQQlloWRn7OqM7cd7fgakLUGIKOc60vSir24X
70mOXO4G9jJG0zuoySlAbWOoeMQAuikagKm1L7DFUsjREoxPrgtPvqmB810ABkjZVrT/qaa9FSUY
8Iyt1h01UcySr4zUuyENYxWRESTJj6teeYcSSitfY2x+uUZ5wYp7rwvE3zCOAZPX3iY7avin7ur0
F+hc7pzeiHTnleKBQ4IMlLRnJL/2ZiiK7wanZSqayeB8g5DQZ4cLO6Q+Y9jmhBBZ4TcBd+/5/VAi
YqNM2iU1JsWmHKH/MrHMVi/WKYbUsSY6bh9m313pxvJg5fi0qQuiEPyvi6UWW+92kkAp02CNS2sB
SmgKD3ZqQqcSuatfjsFZGMm5+bTBa+/YrVx0z2TrZMj1+lQjpm8LNiNaOQNfgQ93dkH4Y0fXKPD2
rBTIs78foxVeKmy0Kbgm9OilQLkrgmVwajWWJ5foxzDVtXY94rQ+ApWhY+2lWDIN7vYjxTBgiyau
WTnz5JglJyQ9Vsn4p94JVCH1W+ch3Qd1gELq6MbUKus6h8L5b1V7+cEYzZjXogmUZzvJ6wqEw462
1SJLwtK4aRiVuGB2YpSHmkek3DZKil8SkQr+oWOrM/q4cEFcQQYRgQkswTFV/grZy1uVxKow6y4P
bykkDlpZjQmh9PqexrQyu20fqZeKBYVlwkUMW6wvsRWlVpvhZd0pVibvPh9cJJ6s8MYNUstoa3VN
3gzxC8iiA5zvJ7/L4HO1Ie9sA8kLubEO8brjQExJj6wgdOuynCgRUEFFTBeo9YUZBkPy2ijXD9r4
pqMfzWXiJ8uPiGeXpNQY9TJAuimtq38NZeeG+c8fE5jZ3ZK5gQe3K+uyLGvnf/onjya+1CBAfJ20
CezRGS8DJjy4YTJC+Vhdv7y9Nnk6eKQaZVOuz7dsLK4g8NaAocIUlpQBrHsx4SyniKuWw1fw8LFz
F5lL6p+yzQXdw/+8jcYUxSoy6H3l/d3HSvObhdYvEV+tCFLntF5c1fDJjB7FJ+NvNNtcdAgMqgx/
u7p21iIUF2E/Ju9HSnrgL15b2pgSizN3OUJhw/WXLjGfcafrTkb8UpibsIzH/qh7TJt8E69DBJ5d
InUc/FlLbafwgU1ee/PzENcxiEgcXhIotp3wBEzwpj76o4qVqOYF0ipz4E//xbgC++q+yw5WMiWz
Fa/CUT6qHqnZX0Z+ePO25Z7ZIwp65LoFTlRjJ6L5Q3/zr2LcQJb0FB2dL7HPD5qlDTAb/qTAmUUq
yviT7VKJ02GnmmM4/INtoz+OGIG2BwFcG2JG6M08z8HY8Urn1hb2c8IvFKnA8ahvRlx1IcW5Q2gA
aOE4Lk+DcAuZck6skOYmSsIVEqA6OStgGEQqzmI5j+pve7Pf3m4ThXk463Uuz8GAHvrXRFpOzc22
x4K6TumXEHoVWc9C82WTQGJpj24iR5mk9P8MexKCZRyo7+IpzCGd/Kave5jh3QrN83Rlvulx1Z7B
malYULl4VQe4VVkyqf1VINvXaF1u1ZwOg/bh+WSu77uVUUZOq5tn40j+hPdJmdES7qpdna2gJ9Nm
eVbQycAzKx+ihf2nWDbVq2XTfx9L9HprI032LGR9UZTXEKy7rn2vjiiI7R05Oh1+wN2RuYxu8C4Q
AvrboThTl4BpUnWsgERDRr6hxrMDY83iQip0IevNf6hOBvxMS4iy2KK/iQZX/tMiC7alLKWD2f2Z
IHfEDkP/+ka1yLUJBnSXdKawRFo6Zanfrl+Y8Ut6LdXjvkxHWiaU0toTrmk/MV9IGRfMu1Rk8hmh
ZFo3WaZp3x/Tq8kAYws66tDRzaBucWhelueBoJ36DBTUWYcixbTlg7fFQxqVrb6f72DVXW/fqhtE
ZlWndl3poQT8lOGSWgkirahROwy0uOWEUJrn7+ffudepSuz1GkbvbgqcM/TLHjzmJJoeRaIAuLFg
UEWNyr9lZsZXTHrx9A9baDSh8jOjjPNCgA//lCqcPlpVfa5wZdyFWbuIr+SVwpOaJPjVHDpUlmc4
gJqonCowcNfcGbWaujkX43kqt6hG18pnevWrpFkmXyuTLomuKf2Pba1pJ8d40KnTYz3Dw1c89IK0
DUGeAq4kQSv5U1Uyq8KpQBuV+4z045IVsyUmfg493RfZmPNwaReqiK/GnGHdg2BvIN/LzGfNl3P6
vvyBg0GyxRAfcg2g/u5+d0B0p6YEikaIvs+pRRtqi+1WuqoP3TFJYXalxN24WoKGcMwvTUahHHyI
OWdo2V10rkfSlq+dlFa9zSB3BJVYqn/Vve6c4paFtrkwPLVGkhdvrZelqKE0HNqCZsgrd1dHWgo1
Vhf9L4WMdGHj5VZO/fnMPHoVatBiKhDtfAHqACqXnVF7B0yvRqe6JJN3XNtp450MPFn9ZdZ7WKLU
ukkq5e8sBhv5F+SDs/YMKuhYQ55zC90unlIAF9WDXwJlNPrC9elr6N8D20dLq68SDYZqa6NtvmAk
mZ20mgoFXp4Gh5kyhG2hlzzfQoeQAN9fkOTxgMax3OHAUbFvF5bthwWCFqYv0PPoFQVlSFlMWJCu
iI4M0IMO6vOpdbrMyrf5Fc5FMwGMAe0OgoTlU/MTGrv/dCxzW02oUqqY5n+GMEvAsWxlt3C6aPym
ta18FZ2vmesJh9VsB2c3sew5NoA2blKpZ+PCi9THVmZ0qJ7+Z57Pmlq3d3vb9zmjNMheYPMqbuVT
pAJEuckEEC9lI8GZF2x8B/TguPKTS6Zc9bPPKkKCl/xLfzgdVYhgdBYrfMGAzCyiTrge8ZnNMaxX
2AJTxA0bf1uoX4pH15TaANS+M/L+oaH19XVMnlZV4puZTqlvIIXV2R8oZVh1xRAvZogLozefc/I0
GQDjwBq+WPEqc5VPMch0HqL1XmLa6eG2s9jtmlFTNKUgaGxn6viCjeaSt5Ndea5aCq3Mr6Aul6gc
6VZ8RUpgV1iWl+BXjUBx6gLNKEXYt4g2kAduRs29Gzc4m/XHpwXRKvW3DBA8JmfsJ85cOVwZ9/Td
KlhkHgo/meuxSsiBIwX4i1AhgxCGUJYofIdAJMXzkCMiBoUK/zhJLB9K2Z5RCCWh79Q5Q6KgOHcu
YONHLgbJzqAGomIAnIXvl3FUALbpjeq8QBaQq/9pnUnyIogxSTOwwp74NdfgUXpB2uUZePk+RWMd
rJ2UR5QyrCunG73TamnIYn/HCwo5wmA5q0du9+87iELGITJkXmvAb/0UgrFoHLQ+3xemUwG4/TWg
t42KDewgnGkou9TJRl4fK4S0trepJLkIN5wnWvGAMS4uKlMj8+0pAwfbiYvyggILi7JBWQbmj9Sa
iThqc3+ZywluORuRw4DH84tySFBnJEdxoeDNAjb1OwzDTIUTZI39dm4ytZne63QpdRQs3YCOgkNE
WcJaoS2FU+G0y52+7IY/07J/gNXrf0cgseHwMB3s2WJJT5WivSwCJDY6eZ1boELj9JZus2WBN9bS
yYg1ZjIF0NJ5PCcKzWcOou84bO1KRAZbccarPyW0GsVfNz30aEV+gXOrEaiK8axAPf9ZbjrbYWHs
pQrgRYqaCvZMQno6WhZx1cz3u4IbejRcTE9yKoC86+GHvpRYzdDN1QkiFnTK2CL+wds1FgioH3jF
hPnV+QSE1ULbQi3KOftwfzw1pyN0hJ5wnJMQwWBhEXI5yuVpYUXfsWHQcRjvM4nWO/f+Q77kcVq9
ue9eACU3Z77QJi1TtqSb3PFii2t8/JYMHI74hQr/D6dXCxMtP/wSm/fDmBeOCtMysbIW02ezx7fu
QNLLDiVVJo5KMHg2Bpwj5YZMGLBQ21kyZvCkcE2mBcESSVRCztIyeNbx9/cgYnFM5ufkr/Kqr6lj
Th5qLEgfGVOEJjUTfY0OB+jZvqMWDtcjNToF+047IAFtGMyHOP1EKUJ3XrGlOsn+sKW2HmHfjATt
nnwFeTJH4GfSp2LGCMW6QG3YEsUyokHchobw4UzbXX4y3P/e53ZVJfn2dI1uFdt4+kuZB/SmY05V
tDfZ2w9lOMqsuNXjTVebJjoOFk5rkS0swUKfv5fC1q8TJiGLaEHhsRvap5ZxZnbYiDaROAT9Wpyx
obGkQ7eKqjTHwZr6esyS8lrF4d97RvtuEK8s4A9nFw0sKfcAAMxwiErvCka3qMWtRc/EQ7+UL5go
FJNsjvXFm5haegt/bxZZFJGqNL96IQrTVJgnDI3d8EZFPKO8LdxCBP9nhlHcqRUc9CujqGaPRjAt
PdKzIvZxa21c8+Jrtr2uK8vKvcas4PbQSnwIPrMNIcwvb58OiawRlo3XM5kU7kRpJVm3Huq7Trhr
qiZyA4pEsGmfazqtKBMgSoDL3Mocd0N/0byknBPNtfw1AyA7tmHVs24v5RUh09MFmBNZqqa/aecR
LgB3At331TtxHRqCuzLQVyDJRwzvGE+WZ1orIiY18MzlMhomO3GjrIM5ubWO0lTRb4WYDjMjU+eO
YaHHnloWwOBgNv8aLgQlT0oyjvfmYCzg+VNX0iRgnzSul2TeNi9eKS3XNmmJAmO226P8sbAPlb1n
bYuWgr5LtQQuzh5uTBTXKBzzw83uO0yS9sIMVlYnTt2fFA4jqI/W1X/1gJ6O7pkxpcW2e/O6ZzJH
HLnbQcEhnnb15V34KVv5mA19LSLXVDSCjneE1uSqpVw8G8HFMh4thXkjSYlGw14TMExgVnojA4jn
D1TGagHGrqa96+tRbY3BuA3XNhgUG4Y5iNQqloE5wkG54ChpcjBnPWyLFeEchJGPpGZvPDmcFo/9
OT7JIgSkB33gHqOqDuPwQjr6ZHqm+kLgbZ7EkAK/RY1tSuw59TBT9+nULcXdENv0B09YqTRjCpQa
ZFUgpKoZtPtOG49QWpp/I8VbmJk7NTdHy2RrujDqZ68OUhOX10FIURODYQCgBCJSGsAA3x6libxF
fdCcEUjitcJYNsnhrnZ45ELCEBkZmyegUf8IxVqgVSm+W75h3cqqzDLsUFjgJyWjqE8dmO2RXBx3
99A5inEldICRl785zEHIRg+6MXEtoh7HOQgGXK7X6Dr9aRgWG9dD2TenH/hL3CixLmRb4CL4Mz7e
LCEW945BGd8Q8NR3ZMcDpLkSpP37lax66w2qYPK2gqz42pAJ0NWkdlvYlSwmEMPBZyC9E3CgauWN
+dfjtv+bhV5KrfIeQ2GcpBhQHcDbCvLyoA0ZO/wpPfi/CBCEp/JlPpIqi3ueUOc4fWvwaK6M+OY4
j59pq76pu7naiiYnAr3LtQYk8QBUIohVzrpSNwfQ9IJssBFnGFo4U1DwE94pn1tTA/3re2DBVabr
M7ZxJjYCWvZjas1ptGloMhDn/a/hNIWh9RaHUJ2rSr+S1Su6kk4EJ1JXfsPZp42nbAnrAbSA/V1y
lXY2+pEZCmRKn1fsrtn1qEotI+eNJzZh4hRti6SNttllghN5kONDm5Miot00i1e9jpwSlSiaqm63
mCB3W03kN+/z3OVsvehB984GaQ97wREppu15pH8NOd6uLWnFwmkxO9uFyCBT4UDY2xDwy6q650Dq
iGYte9rINzUBvvSQSRmXKxUgDjwTDwYbMIAjbkjYyXMTMO31eGvLtviY+MwXH+Av2DfmRFgVXtEx
L33QXABHgceXro7eDxCtZhXvdnn8mhdS9lIMoeYfsOUxdN3XlJbyCa+0I1Z7IPYMeLgiW+lHppzr
8ymlbDk0pw6RCpnaf3J8TO7YggBo4u6mLzGfG4FLO+kVMZVzZV+OeCRU5Lw5XnXzUPkrC5SHbyLj
bCBHg0PcNIZ1fjGqsC2Zo4QZhSxvrUBpN3ANw1wi2HVibGCcMziFdmUbbNIOpYAlRkfn+o3TjUu5
/6WZVO9Lt0tijxGvJJXEewy6c5qyITg1Cz2l1pHtPRMgaPGF0Jf06t95A6+xx2veO+aS8SG37bXQ
uaxIdtvpkV6kCF9dXjTq9MCci2aphfDzAvhOTTCkXdVS4j9RgKqE2UI5jUzxUrjJk0kwr+CJbEZR
yuYUUcE5BwASvFV+2yHJdRC+TSd57z/QqUGa+zfXhC2/VoLtie4AA470TwbS3ibUwAxamJEzI0hR
9K4LJz7IH/7XWgYdAV5vCkKYsVk1KSiao9W0fG615r3wEuojgiW2omwSMZh28mNrMrNlsF93117I
3CTSGZbtBiXraLy8OkkLW4omh0YUkKUQtPxkcAp+MGrV43rMbLBtkjw41l19sZVoOZREtHsscVsX
fNbzPC2BHXpDfSYq+ktRmcZFOTwu+kaBIjkIdNbm4356K1gWOafontrvoFqyMMEHrFe1zDyPyZqX
zM9ATdw2QgLJCbppVZ0gsly0XbA3Yl1u7isCOflA16YV1KH3B0F6cmJRP6Bt3tgVn9VwONdBUPdB
43y4jolnBuu7xrLZo05yNUB74QmBaqAHloVZTMQtiLheiq/yy+kJomMlZD1efgk2jdV8WrVFRjg9
wC97G/d9yoJvOcC0gMZ0tX3lkdbO7OFRtFowUlMR9CpTvtiYrVlA3FSvv/7vvAEVHHT1uoDpQIIG
V9Q1VNLyE5q3WCIc4KQ86EPb90/liZNwCWEsOjRJSdIPvvzxPqgJV+Rd2Ds0TWuGt/M/0rmOap4r
GJy0jUGoDcLauM63FbnzO4n1rD3zROm4I0O8l/p+yXT7Kaa2EECBkEJMUvRYt8PkTppjSYZnFPNs
a5BOT7KNn6BWU0cxK86xSuu6BDaIE1+vDEJVZBllokrgboHbRRaFeQP9JinpmFGMM2upPdIu2BF2
4t3zZzVDjBWfPeZjGX8zAZdLJo9qEh7aFQE6b/TR7v40H2xxwDFZRlzO8AA8L0VrVjOmg8l9kPWm
n3fOUUUErOuSaHUOeWoZbfkE8l6tSwQ+iRgSEwSQ2/dnnzZIGlg5XuxAvs2WMbA09QAYOoV6xjfy
Mit/Eh3L8nmP0viuuReipYuXIoJLpMxTmDHAMCwKGHfHZW5Q5FCe6/lhIYaN8pxN/SjEVyE9+tVI
heTNa/lUmUmUCO/bDtcVX8dav5PBUlEYfukCqnnJIyZZN633Xef2Cdtkdaz/wSzZjJoIOcO0fzi1
kFHbrlSlTCxY8/kbO6sR8IT03q0/Xcp4qw9aShBevXAh310siVB8jjOhti1pFqGcGzG+Vj9vTxoK
yAHUGv0qpI5enNdzgpoL7RXHiVnoWyp8u9IEIBHHrBILT2vmcrqdVJAX0O6cBiMnotbZdDAl1DEM
O+Io36y+e4t6ioFWas+VmFOfI84uUNSn6EFDwIyxmrvk7aI7Ov+8rCyWClY9mrVHXMZhJ5O8M8ws
+a0OMB8V53l3TXWDLTRFg95+S6U15xdeZPkOU+m4L63JQW7J7UMwZGHBsabZS5uDuUNFUGVbY87A
/bpnsTbCYMvgkWjhmc2axF0uPZx7KlMhHcb6clfdq71rSQAFng13qUAaoc5wGyBOd+f5RtSf2Vyc
1d5RFCIZSOcnle+TIXLuPGnZIIo8qmz5/B8cwQOMbvsc638kssPeJHHDXzsPbLxsTX/LzA6mHhzt
WZ1rS3mxHAK6EqlZKkcswoBWHH7u4szBVpxYs0603DCM+lSAFvuyF3Dn7C0G30KG5QtuFMP+ZEZO
5mSGKknQZB8bYS6V1knBOUSLM2oSG0X80eU7DdnDw/7EkHN2V1C7yFXxXfpAph/Fid2iO2IUujFd
Om0RYRpNac9BSubCydNnJpXV8dnLcQ/D2ACRx1WrFRxKWfI57MuxH598TeS+a4gWNt/H9d1sDAtf
rtPcs0bwa1QC1ZX83A26j2K8I+JYAwu0HIkVk9RmLQm70IslRzUYd6CtTb9mnEreO3I/7bgPuQIh
UF8+ke1u4Gvi4CrPH0kScyIjsxC/5GU/qPl42+CLYbKlCOvV0l6OFbJdfWnX2gLDJuPGoEdlOPZg
2kDY07Y+HlzmttakXQWQBtkYBlUaKiYoYBmh08ang2HDbJXKDUNCdMH5y0memSR4uf3lEorYGN60
jQN4LNJ5M8/9QTBYlYZzjGR0P0v+hAES31fGZeKeNq5kHDtp9he+nOOtH+vNE8NE9wXGrcpIz2oT
CusDB5DsZDqcgMSqzeAD2dGXy9bnQzcHue0E3G/caM88Z67l0pIYdwXp4+JiyEdT01u5qWwRKFoD
9V/FasJqR4RWFK7S1cSD4bujOvVHyXq7+i7Asu3CuIGno2YiW9HwmyLbRNkOckaDyhGH+qDPL+BA
TRV9asb8GYDPqZFlHBax6SItZU02jjO6CyjV1MtdBauoTSJeHOfcgHREYoGkAT9/uoEUJXrHyOqA
o0QpHTV3SlzaNdMv8F7zw8yLPQUNqE8rrzAz2mHlidn3op97hf++CKgmSVIaBheNnJn+xyaoM5+C
RMaoLdaOdVbMjia+PB+g7TRgrRIRtpj+it0evSMrrdDMLaDNe0/JKhYCVlhOMRZis5fMKdqTHOBx
d1BKK/YzODz5ETBdLt5N3CpH36ff4G+uLpSm19V2JKyinGqa2XvQY0SkVl/KELtJfHRVh2T5nG+p
eUEzLfxuuc+Z/8capzHyqQDrUerbqzOQDYrBDeznIZOgusHm/5B7meO1A1gKmkA5Sa/F0JEhBHeq
Hg4uigfe1WXdP3k/+tZVt104fCAADJXsbWcWp190v6M0oQcOyiWHo3XITsC9EvN1rLu4ENqOaOFK
WW3A3liXBBTVuY/EKEr6UjV63SqTLKmyabUJOrHM8/xCznP31Go8/IJ9iX6W9o88AZ1+GHcNRVKi
fPo/d5HMLcNlZeHQDFmiYz35Ak+SBxmWFSxylG5pZjOx/aLlt01CTPDo/qoIG/pTSLXvqO7Q39J9
1PmXZvSckl8cvIMcoACb7dV5sO9gUsZLegjiROP0xoE0INzPLOewoc/WPJkDa8NalIWAI0Zqi4RB
6QDisatoPi8yw240Ufr7CawdCURk2OpjCBWMp9r4lORQl5cVA35HYWwaCWK0OmGc4ojp8RstJeuL
KgZwbJRIuIs3MgSnHYrH+1pU/p7hcz8NedJIuByv0wF+DHn3mbbaE7OewR0Z68x6AIUcNFstYbqZ
93CW3Fm5kECp71Jz+CQkJG0/kbmXtzgYg61YQVUG+UHt2v/6a/qxX3vwN2kvlewNh778x2PdhvMg
3f9kA60y9axbfySVKfpKDisBmpuVq0pz84lbreXrCqDVDnxovndczCUcBd4VRlY9FwD9CzLMd8k+
8zWawNJwTEPfgtNyEmqZkzpaLdI5gk110/xSdhnyoZK3ojfB9Rsujm/rC5iY6Weo4ZfhPuF95L97
BsNt22tAKmcjdFSko7jyP6DEWrJXeAcfeg/tnAkWQ/0T+7vmNCPj/BkqE5EorWiLqzrbPjkZHGAk
2E26s0vbGzxbMJ2JOst+qQ4nYhzvKGXy2gd1FLhyKDRaZQlj1wXHuGxw+jqLffiX6F73Kml76mQl
gJZhIjxTzMqFEkXrGnKat/12SxziCT7vqcf044TRDzyYEo7aK//6CslrfK5qU/sK7fq3oBSzpgF1
M5Cvhu9wf/njiPkyyXqqdcZNBgV37VqXv4i80DqdybiV0GIy1DtTTyWZ11uZP7rl50FGJc9EjnR0
32O/VDx2sahobMyXHTyiRKEnkdX0uWjcY81qEZi+I5wicyJrvuGAPPmtEAR/0zmvDmuPdqFp2htf
wLIAcIqNlGcm7b0ZswjDTeD3b84w6MqpLR6gHVu6zqNN2LLbpA5quq4tZwIby9EXMGrBobJ+V0AT
mr/rxXPSzy6Yw6lbdm179pupR4aCUxSlAIY1CO7DBsGhXnZkAkQHjbBtsnenjIGZ4GxfCXriCkUV
zU5z5KT4gu8zS283EF9j2IymCZ5FDYcDGr7fXhw0ucJVQHkbHoSX0+14NtDNXH+QZKFXuDyPxYm9
RRWi0oN2Sggle462z1fQ+ueXfLhBcgQY04Y7nOuvrmGNCRLv7wDRgO1vEN/OPPgbakYPRHQfXHOV
xwYsyIJmzaqhgLATyHjyFFjdraQcDVnx3kNJn7rSNTHv+C8xOcVSgiTTReGyXRYPfwQAxExj2/++
oUzz68vpYYnIxLpqRABOikX33HZXtnnv8+X7hqkWpLihDhRkuNNjG19RGuBaF8DytIn4LKYVSowl
fyLJF/xy/ohABM6RkE7A+RcG6TpVi3dun3FFaRDODhdUdMEBbo58UATls6fbYCfiYvgP18WdzHVo
mFE5/mBS2RgkjexpDuBFnwds/AAXrh44quKnOzQ0EyhkRtCTEPdUWC/oWSOpwLvmWPJbPUxvnKLf
zQ8+PWmTeAIoSCJ37ZBKR4Z7j4xK79yXTdAhwNUFf06JlFFJGR0s71/YrafO3TCvoci6r6KccPCL
4uGU5oD3KBfsVkbz8gjExXE5eSEJjd6BeBgLCZQz8yUdI1aQKnD68h0KTg0IftTET3U9eFurMpBW
OBCdgEb3bMRdFO6DKh/qL/yuzX/SKFREy+Z8270mBjGnZBpqAgZvKfcmHHI1leosiZh6HVhmycAu
LpKhj6JXliJ+F3+nW6paiT4WXhgT0RN4MvtrppK1CqTp8D9VVe9KO/gUzet2PqTeoHlbp0QMiDhh
mvEnbyVr1sfoUFivkAd/cV2k0zmYimIu0Sm+T7FFN//XqyJV3bKfQgm7SeMjEgYXKMuvrIpql3je
92FLVXFym1iNkRWUBcDy0nYDhehPqp7laDfPO49gRRcdzW3sn7B3MQh+3iOFywCmMeOWjQAqGvKY
xiHf5BqV0/GWAhZkm2vpbAb4bjDXEk03KTXwRe3ss2c8yXz5TEMzEp4Uv4L7c8f6hrpqoCZZghej
0zMovyDxiJvmehq7/Bm+8UKh3y1lmqNvYZ8VrxwdSxLY5ZeD2HGDsOVTyYt7pSyOEQ3vN+WxgQMr
G10Ek1QewgOxRrPwKXR0u4iXQyJE2SI+RgZSOwr0FR4upk8OTtjWu/YpAju4HVaHfkWDsN+YZ98z
CRCYtnIo75PtWEGQdt9jS4exS/b6Cu+cx1ggKZXg0j8J0VgEBGOVfq4BIU/Tz+9BP0j28AbRyvgw
EJXyuO1Dr0Lzv6Gw47+5RrQlXZnjOfNT+I1Q5CoB1+SzDLYZTxYiDvh6INpZwfM6tNq8b+R5Z+gc
2NJs+AYIMsFJLMekue1zFpdFjWqt95SPtHckq05H2mZnA9UmhBFxCV0GEGNJ5hXwz9qZmv0Q+iQu
LEOvZYP3qLZZP+pcUPZHdSncqLe6NdbPV25w4Ot/xQf304E8j1M4IgKLmLcX6aHgswPGyhmSVzev
Tsjl3ZY+A2d6ZBODZIasMBxEJzKkut1OD+pvTi5ko4NJYtrR7vaEyU1mre5Nw34s35n2c+nAfXf/
zPad7DCD4ZjTSW5F9zFqT0LanCh0C/kyaPEyuhZI0iIfie5qKIzUEt8+3FMR0/ZL9HY3ITxQu44u
rzigL7Xrmkv4h4GO4fO6YlEexXJH34oz0CtsI/lOImjruBtfMtZJrwObKojR0PKSxypf6t+uOEE+
oCAiu457Nq9KzybKx3RRztZKEHR2Bo52MV7xEMmokUlcrKq5PajkO12jr+CYO6Q+CdOC/rvLuUpL
OpeqHpB/8iUl8SUG8OeRfmcYvyfMoFcpxQqVx81bMz/SYIhtPner75QO23eLuFTTU73EjAR31JEA
hpLIB7A7pTyOxZJe4koZeo/BFI2qgc237p7bfWp5e2rni8p3gD9bIFmpMg7J/zgCy7uiQkNozcd1
KLQbRudPbLtcH6zJUc8HKEKFUr1pbWz0l6bvBmrXpK16OJsJkerV/wi7Jp8iE2bo+tM6GoEpGlpC
jojnGfM3R+XEATdCTTCzl0OdjdOWRT0s7R96n3MV+I2VUX5tVfve2t8Ivl5FFSIaLvp0r1IXw9i5
OW0P5GHBpSypXwkNfxp4k4HafUOrv5CeIGtFjImgCgD1SLxdyS3qbUnEfzH0vFDjUkAqlgoVlrGi
vvPqPyfi2it2nkvZ8pJvSXvuzjmbA6O/g1fTFH8X1peaKxiZ8ZP4lgXxTusHpBGaJE51PFlKYVBD
6/iMZr8hlsiPejAdD6Afz0bzJLsQUyDX1iDuZVC9PIqlBV8pSY9sZiADQWyKnreb/asWdP2md/df
y2OzLm5RW/qsdzQRUifhj2hGYdCXD1wpS/fSkwRJ1qureerSAYfPiW3yC7amuqRdgGiZ0M7lI1Pc
wGU9WQ8JpJqG/0M3ghMWUnPj9T9mXBcHzVOF1MxCX8P3IJr/wbagi9XXk3vwfE8R9eZ4liOzk2nQ
rArSBoS+1wxNXWqQvw+Ll7Zn5EbQDpAysTkbC57u4bMCGv6YsY+E14A7Jl4Lw9gzgMS5LIm0n1R0
8ty95QuHeRuGjiBSVxoPfVhgPkIUpLda3JamOBWkQmgvBuHrBlRfYWyQSK8wcppbplzCxhf1k31L
vr0RooGC14o/ybMrMQA9ZuZerVbM5stNPlMZtuL+vX6M47TGpnesv/rWMel4nDcwh+AlizGZe4rP
zwh+vf6JPTtFSROOwdC+Z3N/L5nMySd/os+7rh0KS68tdpjyzMJFOPA9DwjX0CG5RTA76T9pgmoW
SErAC/ncayEBum1sR90Vue6euMR+OhxdcKcLzZ59ytCWv1yuaG6Kq3I2xk2L6vmsENIfNhDleLnM
yy77nSri7Tcd0xxsSeQT97jO1FKpD2GaMRjbXqBQu7wctgXc01b6Syg90LEm2E+Q+MhEXfI9so/d
54ciVWnwUjkQ63eXi9zntSBrjNVwWu7f5tfjIuvrpmI4aCFOmmLhUwgXLcFzvAILGK1E/Etl78db
3uWUFZwYkLovjxWtH6pdnrmcLdeWfp5Mc/RgWXnki6WSjDrM35hloKtML6glcDbr57iPq1jYIvdz
CAEXQmjGfJRM7zbWDmeth+b7Gori2on4O+zL1ixXDMwmUUUfiaYZz+y3ZaI3q8XlVmOQAgjnDq5F
Omgbu8hfu0HLb+EhR8aaHzYVocUobu2xfbdHKflE5lZTsFTTH1c5fGXJ+vdoBHYHyVqfXbp6culF
FgvOG1VX8CXcWL9SGF15EON0LBps8LUexBJEu8QxFCcjcFoAVfPgQXiSg+4Go6yz/9PqLaFa+50a
sFR/KDPMedl51Ru9ieWUjq/BFtw8jXolbjQktEJ3eeCkCGEl8NPBbuthM6HbFfZ2d2Xoni9Myz1h
0pu1T/m+JIcMRSHF9XOtoJsCk3NxymUrDSOi4AcgvuIxzpRIQik52KSbJssqUK0mj2ZkoH1reUv6
uIwVwThbKb8c6Ad7YJZRJdOWxSkxRFH3lbedLDypkCNHHYyyR4WlSGDhIWDMCYBnUe0GJsEoNlHR
aBN8h+rGlb9Za0ZNvZhw7aTs4K9K5idFMLzCySfxjodV9lO/+/EOkVD/jOMLViQ0QqlEt5aFpVEx
/271JY9DtB5INkzxlAPz8Mjdf/KQEacSDplGo9wrbNObSUXGhfXONnK4kcF9OPVdUm9oafO+Fx+c
Cst/nauM9LuydoDMyDjH4O4uJTIxQeiNxiiytCUm0bsCUWPLAk/Ec+O6Whgnb5cUfalovoQ7vLKJ
fse+L2BPswXdaQ5LWNr6imIV48kEbfBZAn7Bg7g+HzwYGhKCVJUFq/0ZzyW/kDLLVtILsxA+brxS
aybHKcAj5MQJUTH1qArD1sVwR8l4UM4UtOOYL56Fzc+O2c3PD2Rt7US0iYN+396KnZO7+7LfYaR8
VgRX7TR+1EgX5s4xc71bBtE5oGW+okULWLz6qUUewS1nEWfiCRri4Ckw2kfBQrxD1utlgPi1j8Lh
bXrMX6/P86GXeXV2Q7MI2w4uG4aRlnyv8/gzEYQ6OIa5jJDHjtqlZuNN2KBJGCD8AWtHF8nT0RuF
yEkYG++yIRFzN9mb3sV/Mh0SKOKnasRoHGpN/TLp6NVkApg4w9dmD88/GU0n6HdzmyaA5mhthQnP
D/WWwz5ycnDcgwatAuBsk1aOY4Mst5sXT0ggXrGnVHCc6R6D/R/G3h2jphLpxIlD0WKKvMK7Dxkr
GczMPczwXZgX8RyZ6snDxB4WvWFVlwlb0K2k9EIxjyolU9u08qfAqY3yFOLnbJBz3+r5iH7YV61t
e5PKW1hoRm8Ewm/xD6l9YkqP3VjXebxFibyNv/IzezO63szQHLNOJs0NwoFhafyZM/OibfbEO5/x
6IKRPtrMhO/Jo9LMgEyz+z+uYjpkw0TN2lyfG623jyiWyU2AGwfj1BJh2VW0mPPClrpAuXhu1L0v
KxztF2b7+95RYdBAJswjkG/v9rJV7zkOyohrbvbILnnM96+RBIIt9R8t4xFNNn/TuwGqZZe7ucOU
QcoLJkzz91OLIoPBTh9YZ2s5eZDTBW3D7A7YCpPqH2x2Tot1vitTigckKGVd1K3FlsYe/76B1orb
sMCo5hKADue9kLpLjTOYzho6I/+XtSSfEZGnm8H5geuzjLXli7ZmOmXuZVGdowzSdZ7oFm45v5VP
+QBfukqUGc5qg3EQNZ1l8EmZfO1DB9KbM+s75Yy98C1lNzLXy47AWD7fCyqFT+ltxNw44NiV2QYX
52hAkmRBWBp50HhiPPXTrWtcBZLBDL/2uMyqJOC7ZMPiGIrNF7fBWfJ4E9j555I1VkTLOUc0gksp
lUSlG5rpay/2KTu+uXWxma03C9eBt0i4odaqbIdRnLNdwBUYGqMzdchPXL8fJA/sdOBOBbvjRr9+
0gMalLqfqYOAGh0R3tiX35UqQ3Cn1WRGDLQvI7pbxONV/MapfUU8bGoOl5pmnCUG/leibfVxFe1o
jiXNAwJRI7X6Tsx2CN/cOXEG5WTkrUsHj7UC3CPU56cQw4ddJUy9PT+hby/VZeIibMjaIcUDE5r8
JU++qYRoMjg56F4q91Ww8OydOANrr2EpZC4qWvC0u6yJapO1v6PiTyKVdUWG+QXejZ7oplWjuLfO
up9pMPG6ZbtKQJDDJ1w/3p42sIBgkky3zc1jr2GgjJY88+xlOnAk8CROTfjLQg2eRcCHhM4Tvfzn
Z5irgTEgBW7eozbQTxWwvCriLE+C1vIdxERSkXe/HHHa/QIBBznKKixWPU8cxDhq/hDrEI+Zr6R/
Gz/JUWc8y33Luzg6TiBYg9LyxnIJj6V1iCc4Ob426JZtx+Tet//g1gFOwtC6GKcPUH1igP6crxqt
lXqcU29XJSc9oM7MDnsjsd+1dCZp9JbUn7eJvIlDxu9u8T1mJooz/Pvj53UgiZ69dygWVTtscyo6
k2Byg6p3e6FztAx2W3bLvIGat76SjLfL0Ms89CF/TgDe1WYyGEMys6YHqtPSxHmeUPkCpSyN94d6
PIZ67wEsOLGBRlczb8YO7yk0xtK9jL6bb9fAsVAlU/cLE+Nc5jNuDNG+6HifWMGQKL+HfoVjc6fR
Rs265bfGTe7emmJhBHcSR9B+5+qrfHFL7UBBx3j7YOk4Eiq7u//cBJxn7bHyTiQfoz3KuhsVWjFS
bN2Q+c1jmv4RzPE131KURKs/zW250HSMLBzQFZfHjf9B/brPPGpIk8pqLjI1EPPpR+0HHzNU6eUZ
nhRWIOSRuNmTt8XDDQMNmZZr2/EwtpUkEXZJ3aPpawPEcBswzHTbWyVaUugvFmMiyxsBWwsaefLw
mdmKyd877T1jrtNVCjscrlfje4XfEtuxdGjMQ82rH9ZnBhvR5JPCAg1fVYW6By6VO4yW9w7SZcLx
cUFMmjSdKb5SNcExSzegycfR+2q3q0y+grsGh4MJcZxAuXCp/4CxLhwJlPylqZxuGg/gJNgpvAJJ
MEQQsctiPMyo75UAyV/GWZnTx0nM0jxOv+OtywiKevDdMYdDQc8PqTSRFslTqqkl5NS1ZT4wka5X
RgMYCVyantji3Cbv2DNbON86FfUWeyWnhBq5GjWrvEsao4RgJC5odcpmDzTE7Zpav9Pk9hG9PEkp
+/CjEE2a1qPMzkLc2neCYBUrEtcwJrHQl8aIko4Fk3V+jESm58OhsUTo0uAnX0iwkG6YZTgdrU+Z
hSqvB4A2aRh3xbfGOiYzCfs7H/fUhFEthqCR5HcYHtNQXNgyj5HkwKL9DziKTUtKOQ+wfBBKQRqi
yyOcB6gheakbhqlAgpH+A8RxvdLebNku3VlHHcy8qF0CVYJV4eoW2iU4wBuxuExEW0BShE+BAI9F
zs25IVYEusYreUjm7HPACCSUR7zwhfZuNVYTQD0E77MkEurHWQqj/B77cJUEeFZdezyV88gJrjy0
pBl79mn8MHgeTsFuO6/SWu2zUtSOnn12P9TVN3fe2sZKpLhzixcUWiBcBae0bQ9mlv4bq7FEJPfQ
0nMo7wPTRuaXKjX6XO1sD3I3R852XBUm2dWabaG5ais3y0BOvqCt09VZTXblecxqLKJdNOVvdz2/
qr2Eoj7YRuWAqOOYkkTFuy5CWngCkBLdDvLQrtSaU5T24HsTwIIwcI/HaVkWPz41Ad0Cuddw1Oou
DMztLB5TyTLv7bn8pJ+aYxWz4SPxX43+dpypGWniy1Ob0hZkGRs7Brwtm2kzw9ZXnNmeg97/jygt
Cj5CSDrJXas66A+44TvFISgEn0G031wrPAxd4S9OYx0ccFKuu9a7t838QXcoUNQ4nUTLh3xL++pe
yv/kLQ65XEsYWy8NeNoh2POacwN1aYU4yIrxQ0cB7EyEqS8QbOpCu7fM6CFiTIF6JOAUoSIUyX8J
97IrRG0/V1DIi7BgKSVy+o0/JWPoteSlmNKKu3JXwLPAOuOv6yA9Ngkj69Qzpw76BL/8ACxipPqo
ZF+RaWg0sBWJJk+5573pnilyCviCINOUERaFTHJ7BeMfsreyDTaSQx+5OhG+I6Vc3LY+0l/nIalH
W1jXiCMyXcASBdkAKvg6ieyl9T7zjANpP4r+A4mR6ds6HbjfBRBZdDmiynyguJATThJ6A3Ob0S89
j74DFrfoSuR4Srhzg+ocWqgAh4QlwQDu9lDXycMHqVwTNZkAplPVKP966feTD5vufg9udEqAcaGe
R3D0Tmvc/i7O417rW107+2H/T9Bb41vTzBzrgHz+NxsQCTtQ8TMrVfduGpy0CBbPOGBilaqvp+GI
YnFhzNprMtn99EjOyuL5zn2uE4v8l14fRox8HjCD8xMjUvw0co68OGQRaHqvwGcOKj1UQAHoMaZi
lR4bOWc6QLOPPC+DYGfESntj0Mnd2ztB4dKcdEky15mKqF6UawO7mYa0OBJfdfADyXfgWhDPkuKi
Hvhq+XZ/pHTustzUsWyVTHPBuN/6QxmyZzg94rtAhDlgkdhvp0OnxSfJsgrH644fbpNwrcA2hNIA
s1F5nXLRjhETcpdb7fwxKdWG0znwZ2Hg0+v3fVRZ3wfx0UREYa9qOosI5cjyN5EF/Ib4CCIFLjIW
PKd0xqaBK3oAgOd5Z1IJXu/YtU7QoMqDCoERfI4N7W34e4PwVMauWxwro2b5M3MZbFK7O/B3kKkJ
BKfZOoomxasIBE525HDCIvxy0JzC5AH28jTjhRktFtZusE+qq/wE2zP8WrnAKkMiyy2TzyFicaML
lPvNGV/hLOGxyAean2qHK313hwUoapsQlzX4SIyQ6NCdgy35nUh/NhXld2l3s6mmhpK4tB0E79pv
C0qiXilhPz5F1CDezFGn31v0Sv4QR/gwVbVFCYoV2WIl1K96Vt6UeNzlot3p2dcNe7jzLjnw9ZoS
/EiTuriJ/drRvMmikGtlSDzRBsqJlBqYNwL4sDCJqsoOdnLv82XVl1IMRtp1emwbdxfkKQ7zMpvh
yfekmu3GPCaC1zPaG4h7ip/w+IcpVvNXF8WdgPfnxLk+cuUH9vB+IgHgsuT//B7PeUOGIkcT63WQ
SPYWX5rD8DlPMLKJieEB6Dp9V1PI+pSqpknntL/mtcUhN59dqaYMIhTAbQf+MXlap19F9RYV6wUr
YVHwqSWgWc9rUfgZxZsvjzpWVwBrO4Xv/DqrHLe4CTcPXt1IrP60MNj1knp3txbTQWuo6ZlCH9cl
7AHELg8L5oNK2+X7YCc+7ZJtwWz1EIZuL43brnURXhvXq1SO2MShgTjdBarLRfZME2VSv3c6+IvA
Mu0gtiE/zxBNETkNu5ZKKs1r/wI+FYhOCWgr2P0so0xzyatA2LoFUy+K8/svymlu4q1YKBmaaQyq
kwanNTIqOS+LEjMqUckpwEVRe1IFjP5Fb15MItZ1fLIhG+hTnY/VaOBb2vtmkk3GV2CQB+CbAQH1
k1HACgRZOMDp55+oiwUAYp0P64B4D+zcNCQZOm8hn2iRVvmNRhwDJo7TIuRbs693RAd0JBnSBOKJ
Nb66V8FYw/zvZ9hDTfnAeZPlBXbW0CygTwL0ozXdXVMDjlG/ktfRUwUbmZDs85mrgjQ3dUVOSO3U
CODpuR6VhDoYT9sDN0nx3qhZcNJCbNzxFAAqZpxRgrLpoMb3kxzLBz+djFOJBh1Oblbsjuui3P94
6g5pMMr0YGynORMMKpFgGT14g18oWgR6ocCpBz8YZrp3dQY9blQq8zxey2aTow/+nACSE1450ARa
qEwtU7Di5+rIJuvyZVdGzuW8JfUn7l+nWPhTupCE/K6bJY9AsZotAaGX9tBj62hxYqJb0UchS6KB
Bc0R8E7AaUySCaqHe+goMMqHxV5e6cgJNFjG55OtuWELBd+7j8sR1Go4jasJSGuSsczePM8BWudu
+nL4dZGHgtL0kZ75WGfQi38LX7vQGGkOqW1bEaegayOzQikzH8YdoYSZ3KS43UQdKYDoyGgFsof2
3l6ATD5E6333thCsNyethxDP00qeMlQh+khmklfZkovX+FGNtmcz4EevkqqnwnonXYAl3xR5O9Yu
EoKHCBt4f9EJvJ40W1vGc+BUU9HH+pSzWiWZzKfenEMhVWYqIg8jgL4EalJilZDgtlFZ6EGvc42r
FrwrTS9A8R8gQnahZ4+6yluy7G9IG6lscQEPh0cmxOQ+k5XawbZkXknM0MOIzuznr1+6k2QaVUWY
Af4Vv7C+uCoCsOMNLjuROjqWWJjUnsKlue+bsvkFWY+oGd0yx4/FqlasNdsZhYYEgWDmRFDMZXnz
Ws27QdjwxqY2269UL6jfG63ihCOmeu7lDEFeFbbKeeq6piTrzZ1KzifIufVzjBQExGFEnOqwyJKK
jAL0V1FbLS5IvsSJwwfpI0Ocvn/pfo8DY6ju6Juaj8adCj4u6+oXbkttzLgc4eJ2DL3JucitB4BW
EgkQoqysNcfSACQhPij/PXMcpvSVY5EMsVVpq4JNuXTPBpOj8v/Q+78yhD8CGMUeHuNDA5jWSN19
O9LCsCzLRQCT9E8e7PKyGfQ774MUGdDKR8enR0POoPx4LkZLwreSduCzad1PL1wIuk/owTJ+SzL4
y0wUqjbkIuIVUsvL6Ebb03m1T045YwPWCJTRW7jl8CMgZUX6+U5vjULf5j9F70HtUyiVw9NwTDMy
xLzZzFaZ9jQxlfVajb/R58JfCJb4Rrr66UEueYlISedkR+lXI7c3OZeV/3T9HuEREZ6mcrmaHF/E
MJMtbU0kcvhEfKmLpNX7C1kzcHy+wskYSiuxHAuXmOLCbtZA9pQFHZE+aWizACkwlNKlJ66xlb22
bUSXyzhqavSGgD5ZJXg9iWB7Ann3wrFXPqKTjft9Sv+caAJgUr8coTV5E9zAzYrtNb3j4gZJNXgW
Lyt9wNunY6P2I89ow65866x8CJjdV0jx2KsxUJtg5XKCCPtVcr3Ei1HhR3RvsUTXjRPfsb1Pe+5n
FF8UxvwNcHNQkMOdcOLwt84WyMvpioOy8QAH9XCvsOAnedGrsvaiUf6WsY9Am0uZRhON2Zmfw3NO
5eh2ZyhjSlHE72DWJwf5NysMTSnldBhby1BmAmIkDhwHBNjbmiVUhS3JrCB37lOyDlJ2kPNfXNdF
PwGiBPFoKfw27E0AsLSPxxbuVbF2qPWd75rEa0FYwo/SnnzLy/4YGHCG4YPckCMK4xOPwOjiAVc1
4mHi9HaUej/So2kgvYftAq7lLVJ/+kOXTG5aOnES9uMqUfUvDY9JQ8M0pW4H9yTG/MPl8cyA4zIg
Q5MISAcYgPl4Jpf3zZkTq5V/jtj5RsfPFOHjn3kLjZupt1t1d+7ocC81MiMy8y7hGsCUC1RJNxCX
o8puDDCKrJamkhd/u2lTdsMJZ6236Pg4m5pJVI0DDPrm2RC1l39EOwlahLwOuQZflutuDvq5TvgU
fg9hPSxlf602sAV7wy6S0BX9bXBzcjYoNrWj1ya2fOJXW/UqPtOHoIDqgC1U1TB/T9IcT5MCLirB
KtE71En+22a5kYLWRF8Eoyl4utMrKRuHx9mliz9P1JuDRlbI5EUV/RopVY67Td0CXKsG8CHS65VP
7ZR8hNRFyL2abaYXZJgKC63/XXmCx+NZptoAgzytA+CClfBArbxdlvJHvkIcU9gX+JFTKJQbC2Gx
aXD+xQt9elTTdT36VuZwybWDas2uzQxYt44kQJ7Gp++qgx87DjRzjL/Iv/PKPOx5IUkyXbXgy2m6
u/G4JyfgwPnD+eK6GTYCauL/Yee3+rHCZYvGOeM4AW0/rw5pU0Tugm07h8VFIOaac8NLBaTq4QDI
0egspo3lbi/BmoNgPo9yGHWYG+xja23RGWoWFctr/Y6K8TlgxtQpaBPvTlYILHd9K/vLnuHRi9KX
ZIP825F7isQiUQsJKYoU8w22AceEylDYivQmvCQtQoTj/Xz0GLKUzjv9+X+5dx2TG8s5d7QgafHj
6LumZUoqH5bo5UjCGIKb54NbOkwrErYWlbkCDO7HvaFODmTQW2ME7pM8Ofb/Pn2X1+C3n1utyRWW
6+AzTn7VnMpwkZd++5Hso2vDhjjmlwcXpOwJW+rmQm43RvuEQEY3R704aRAz0kWUo5012K4DpKwu
HdUD+YezPzDOPCmRMuhYI2k2Iac/TmCcyBALhJce8Uv7varB3FAh+xN4+PUorkDmE8UBzJELMDFB
Te4VrhG6OcRUKiFj4Gz2UA+xChfySa+1d5Tp5wUOiBEt26My+oMJNI+ELqIzMIriS7ThIi3wced4
ZAJPkBG0kQFsRHN3C87zAM4dZvydJ4IYTybsZO8ZZk6RB++mwz/zUxu1mag5k/+3pj0w1aWzucQ3
BqwPErtVUCvJZG6NvzRZBcSLsnnC4d01F+zennlgVFG6cn1VQvnaO4rTgUhxcEyWWtFFGdUIcs7N
f0ZUAj9lbLH04Crtj5wJB0aDDQw+WvQtcI9aIaXFveEaBjEie/WANqsYLBlQtCmGFvubB+GvaxGm
ZLhh6ukEQFL1WrL8dR9tx/04/5kFbIS90DL/naagOJltUb0SObuhu4tNwi31O7ZOZ/lUkK1e4/ap
uG27ih3GKl7wsQzjP1cfTJl6fbLclDTFMy8SPrClDpVRUxe7rPLvItyUnLVzfYsnyihAJa69Kou6
kCG0eYtoGAEEq2ullMJSm0PhZus+glK5dVuZDuUpZCP6VaqWUAfUlf3GQn9oRYtqm/vNFoHCOaXT
ylo/8QXSEHr4MAIoxbaKDiAuPVXueqzh2Bv3bgb06C+shsUrpo0uFZtazf4KtNdRWItsalf/cq4O
+hDl8gcrLczyanmDGSfCucCjWvWWlGGVYxV8HOxtSQNrpZ8ms2ZUkCIhzfMHYMY/sJY3eH19NNRx
IYT8m0oJvvBu096NiWn7GpkeqTEZ118oRFeVW1HGD/46kjYQMWI9uxy8CLs0Zahra6bCbcOi/9OK
4+PyRBmTtilzSSc6TziexOfqkMFm4o2MiELIpD08Ho7HQwl2GWO8RNl2gONQ17rypz/MQzNVEo5m
SYb35B+NOhSvFjxlvcGCaWUFPbPLt8QembIfDIAw/2KDs1xxuZtjnk4rxKKNncoCOJm22B892BUk
e7fCrfybvw7DUo1zg6QBVJZn+XJyUyeXcNq1zcC1D2d7OXRXFhTULwvrxNSJ+Ne2EBvX928gMHh3
eL3QMnggOO++6EFd8J/h8dQw8bqmRpwSzTJ9ifgr1Snm+xiYrjPzJob5Sk+eW31JwA4PHgQsjaoq
PrdB4FOBnOg6Olk2S49jTkUlbBOfxTnc+7zWAdILKkNpHh7DK1u1GGo61Isd4Kpe7SKJR1PdD7y+
ADlP7jtW3ocypeYVwuholG7SGDfUY74wznCAKn+KYIg1Gt1nQIfWjASgnrv2BYR+Z4bTGJM4Ccs2
buKf78BkawYMZ0NEI8utmbDZloR/ZjYylDM0RhxsqkTmI8M+yr41i6DApYilTaGuJqoFGlLpgxhx
nzh6XL9b48lTSLQVfEWR8m2gjGyY981FK4NKZ8Z/8WNTort6yh44nj6VARl7kBFz+wXew5aFSIiw
Tyx12gCegvPY6h7a92oEsWKMWZce6LfclFLmMPZHlZstziopZW4tRkL/1T9QPNEcUbPG6l30fNAP
9gDTU6Vw5YECKVIjlVihwKTF0Lom27d0qT3Wrvnq0HClgN2MkIK+JYecW6ZJZyYGLAlDYjSFew0i
wY2i35jIUindTIJBjGiU3fxHNyKn0zkVR0j5GZ24MucmYJP0oDOJj7fjBlszXyGWTmY5Ld7APABE
hThiPUP+kGuPcfSt2myaHAL9a2UEuG9jKrWkvA/IAYPSyHP78lxNlLrKrF0ACOcEXb/WQjoUU166
xNV7lha+6yEM5uO4KLBQQfUAhzPxeuIUANiV9Uh+fAglcU3y2nQk4/t4iSphDNIP8uUt9QiEi3YT
AkRf6w1txSspB2csoNhcQAs3XWRmmlprUJJlwFOkWN9GkUlXFOqihMNi2yemtb4QiM2VScchdUqm
OW9iV1QGZBQziFLmHMLRSI5ivzqumXx9IANqn5Ng2b3fhaTUCOFn8nmMUgJhmMrjMFHTYsPKdbXe
JXdYwaJTY9meA4CuKgUEo+56WDUIUwtX9dRGsuG++Gv8EJ4RPntmXbyj1Tc+kNJmfud1h1B1qzdV
lKTYzUTO83sQq49TADgO3cXhdkeCWEaRnxgRSnTDHUojbYK6Cp1NWMVYVAOOskzKIIQh323lrUw0
d1H7PiHUq4+Q/4rRlxDRPisbPOvsTvBXHL9PpctEbipnm+7dtuaQcXE7T8onW2fqJxK4Edc/Lom5
wCC3NX0DvaVYsHTK7AUNo+wt5Ng5I59L1+EjahiUakyilFykFsQAD496+jCCwx0l2uFINKewfNNQ
YsuZY8Qko4NOlWyQ+BBiSr+jxVD9vFcNsfFbuXu9qnNkAoDSAt2l7gR9QUatRPtMgo4Tp9GJAy02
uu/iV6T2xvd0TMzDTRg7z6ll7QHMtSFPVG7h6SQuJzkY74x2im2BVNaO1fWpT+UhbVEGCbrR7KhR
Y/qgEaIXXlaFNhiql3qu5D4uia27ZWtkQlGAUBS/azxY7Ne5zvy0KsD5rfgFAc31R7J/CIFDHdZt
plbGpfWdmscZDRgrr6Igxd6wlzzbp0ci0XpWS8iv3fu31W/gteJYum4FRu9kZAZWn3LXBEH0BEMe
DTRaF9qvN14vxIo4n1rf8g7RuwIg2RpV/sIRd41uce2S1HIf2Vsz67b0gXbv9llVe2sAhQLl4kQl
kCsMSiyTT1o6ZdvMGUdO0DdRdQ/XCD6F3tnKUUXh0x9bBINkcZnsiRKjxqZTZIBAx2MgQJ7hxS80
19D4X6XOLYnaJ8fVqsmGu2zN24+xNs6gexvkIiZ00DQ+BvSmI4yF5NOyQ1S7yoBkWP6UiZIALq/a
kEIOWp4tRFTTE3McJgbc3temnaoXmSj0xAeEfhkr2sXCsN5ew6rFA/YlNptZaMPPTSFgKvIzkTpp
b3ocPSNp22n8Prny6M2dOkZPR8mXKLGqraZVzTWuSOwT1A43Usj/0d7IG/l3BsB91kML22CHfMQo
M+BJoBwf23AQOtSWDeAKXp1hJp58f1yMjDg4PU3v9n5eOBKAwD2Y032XiwUhKtwaAT1k2WZR19zA
LeynYEWciTHRng+JulShtiMVGsNmSdX0wq51XAnxG5Fpto3NrR08s08mf2k7JkR4J1WLjSxmuSKG
jEFbYuFTzTSiwBAwcegZBGDa9YHHG9XLNARJWr3YbmGTN6pgYnswbU4eMabLDpWJfnd5ULVS7iTG
Ik1v6eMVYsV57QXikshnITV7/5GNYmNCn/SR+irsDLJ+lS3KtTYukjepmMRmRtBCgis6m8R4JEGW
mMxUdYIw/U0Y6q/yTmwLRDiYKL3FplP6/b/998a8NxX8GGr//QIB6MIfDqcrIvp+T1pqijA9fgU3
9i7cVB5DpoqGOL3OELkoQqAzMsAKSf6PEZKoEiIyP/r290vwzNAi7D7PpgKSyQIt3UJ8BEc70eAs
jdrBV3Ltt5bmzLL0HBMp73zRh+pI/0YxjvX+ZOQuYYTV/vPQJXw/sTX3oDX9O29R3U2I2pmmzvVp
O7qNonIhsNGpzw7SuwWP4eU4H6ipb+NJRtUiKva+IHT2fBy3RdEei7QkbggMT9skR5UL0Jr+GCNC
WI/EG6zcJTcbjWx3CTvQb9YxdV+167h8sjj6JKm21yUU7Vjky+dPEILdvUj2gvDjCW92upCbaTYU
FDawT3DyCCnelLRKDsonqjpNIuKnW2k+hhWKJDeR0vZDO+WvSVHHMM/OZVo6PEJc8Kf/db3BXhKY
eof1cGge2XsELzW0X/FqPjzsXpL/RlKOykqQDjj4+GpdJKw7QbsosAZ2/olB7l2EHkN9Zvc/9MTT
x7rnv5D/b0pExbRmZcxppyICu51EGWrCHyDwbk9YGN3dZdic8Va+ehpcw1bZQ+5/Y1f9itxbAeKL
UOSh81Cc8FeTlNtmOVxtnFFL3npoUrf4TL4Gsdl74DbkmHEFgQWkopMCYiIaiZqRfxtMR7h0nGOm
7i8xCjLctGwOEmgUyVUbvDZKhf74sM4H6dUpNglMfP+GpK8EZnIi43/coWJJz26viVvOxLVGL/Sf
7vsqxLXsw/40g755Ad60j+64U4MeIJQPASw2Mum5vrZRXOtwzJE1bW4wRSaI0+zidSzsZiAbWDAN
V9GA2ewNBxQVkA/bR6LSyQPa3XpXbHcCIUnj+S+5jGv2x0VyN4/GXq47wjFg1Zk75YpzsZWCz0yw
3bRxgvffJhnEHsCgVcV3uFaXcMqpNMF+KHLiKlGQMnL5QDTW1dAeZ63jI2qzOyVfHOtBpId7mja6
7UBlc1tQpHwmynwqE1VsncJoUXD4eaGdhbVihg8sSSINEnRJVeTShSs3IscmpN9mkdZKRORblGbB
puH70zousZk2hxh/ecoT9QimrJ0TbuKx6jQEKRLgSktiMPTSGd2FVuPAUkmrdwgss/CHt8cK7ial
jZGLpp5kaCsSZH2uXuKTYuYhEwtnQDhRd2eouSJoX25/p3py3iOfwuYtHycvHVabOyl1diujtEMX
09OByWRAZGjfq5vbpDMmpMH2cYAy69bN3it6vkE+zIgr/cW7jIapfXtDE/mOSF3LgNfG/LuKVwq3
LjtmzXyETOY+bikL7ZXVZK2+JwWR3ricQT1jT64/sOg5SLKdAcj5fYKSk2MqK4UnRu5Y4LQDX5at
XH9AYExWB6X0dnPwMjss3EeD3Nq+YK0mQU3/JT/qJPQkwkK9LsPISm+lOp0zQ8om+hrh0fjFaGSQ
JcaW941+f5vPuDzxEuMzlS50rstFBCwkGHV53VTLdw7RuCPCdmJAC+eyaEUqofcG5pUbmwyK8vh5
h6JWYRlyt7W1FvAevedRfaRw38kmBoppaBsM/f4ez2cqJJHjbRiakyHbVwCpoCEAWk9udfWQTJMu
m+AleID1Q4T9RGJDaCIbvlMa3OBuQHlbeEugcO/bikv3xRO3Ebj9IFqjjFdGYneZUTXoOEA3S5xe
Z0vE5AbCxKQ3P+aIBjVuiYTbEvT0XWxI1OYAwHc+jK9Js6FE1gbYG50oKpR54yQQAo9+xfqSQKEX
YXtRtGpN2x++ECuuyCQ6l1w0KCXkIV20pcL8bh62cedU7Y+NvB37IYwTuciUtOXCsbLA8M9hwd2a
z+3D74bPE9SO7mGF2w5v+Njv3LxwMu2NlN3eJ0EriuX/+PggRczZlbMzyFVszUVIu1ca0q57rjO1
8JnHYO0PiWtqMMTo6DDeyiRf09TilBdKeyzF/FjrzRYUb0ndozQXYK2Q14Qqj9pCFO2UhGyxhIO8
S5/xEZPUojkFWRpu+UFSkoxOlURgyg/inCalBoN2lygEWJ06NO1Y2iVXUDVRrvUSxwgJu1LI+Uv9
S/Ou2L23klgswpjbLZvn9vhT4xogQ7kt7AycOgjMsUhAd0RLFBuZ9KEuc3aDdWHywV6vh8Zha2Dn
O4WskSFmtP0i5cZnCDl9SSLUSzAxZvTHDxovN7FRgafnPOp1jA1uJ5G/lt/GdfGd82z7KyoWRCU5
5qtyMFTxInp/JYhweG7BGYjAbuQWMMkT/mpLEfClcpk2d7UrljWJNJHK6YKf7qdkk0BTj6ZX4wLe
JzItKcunDfeS/Xoocpi+qPg/menmvbCzpv7Gw0VdfyIMOPswdM7/PmjF8CJQaTuyBYReB1R7UuQa
+fBMTAkp4zCy/n+Je6JYZrITTRoDWW/DwaTS8RPB6kRGUPBUXXuuFttHWSsHMjEmRkBFD87Y2c9M
3viu2KXeIZ0MkR9MdBNuJivgdO/j/rug8HTIjdyTK6MbM/s/sGI2cjwPNU+1rnbSuEvJVt6IfEeo
h+n3InnJe6IqJIEnbdeddUC8dj/uvYFfG9loyWYRzUYsprF5cQ9c384Pow/uaguGjTnV4nkYnNMi
aWXEOUJROkI7tar92lYIOpRAbmcgRWt+jzvQSxhTHLCCjlwZhMdHraAaXFq6Avaswg2VH11vXmRd
sEwHN2qlyhaalH2iUUtb6zrzcBXxJWV2rMBGgfkNxnTu9w2/W7MVbjKTX1kRhwVe00lsz67tKHgN
L3PKjlTFhNTS/om7mZE2g0GZZ9vy+KYQCmq4rHdVUvW0FZ3MYCTJ8eDGbhCSyheEEKRbw/1JJ4R7
l6wCxFrVREU6rpi1Tf1MXhJIG7eH19S5fyJO8J10RRZygiIwQePzjuDsSwfMahXYnMg1gSiOuD9E
+4LF3yW5HEyw3jPJBXH6TOYnkmByckOYxpaPXFP+J0ApwhxoG7pIhzI32DCnP3DZ/o3Bv7o2tK7+
mtc3AOdwe+uneGkYhOKrTm1RHm56nowgCcdy+PmfP85jUZsLxGXpTToSafMv8gOaeA3gcEIllpuG
ezgDbB/Ct8da5a76hPVvxaT0iBwm0uQXACh4F4taqj0D+UMEj/FZKxo07Qd8P6mn+i6Nz1ShrlRH
SColUa4xGOdCq8O9O262qYFr1SleaQnPu+zq2yaHKJJooTYIKj6czUujOUsZ5EMNHGzTufl8MPH1
NVcJTNF6qtVvlNlaDPM2ni7YfP5waLg4nKlG8aY3/7oTfqcOVaicW+uodBPvWmroVYKSozgPxTrz
5fyY0r+PC3S7K/6E6SvLe3fu7Ou+Xt9fEfS+vk4RfZhHK/efcKjWZ4iTHMvKsgl+HfuG2PpyJQMJ
94ODyDbh7WZqj/FXXI9CgjPm/JYm7P/pI0GdOPz7ssrUGNer/gZVo1eduBeSt+ahPaZEhff1WeE8
AQLjlsvW+Od3pL0dycG3uHgkl54JbtIpw8SDhoVpD3kPh/JCCHCNFgKly/gcbsKStM/5f2YTcoXS
/28iBG7kwqKWJUV99ReSfuKeZKduGDq95dU4lR1SOqG9JWPlf+8VLsKfOFEhjQoTt6c6I/ryYHdB
DZUntPDqC3MSrTg9uT1u+M/qSmigV/qlDmoG0/NdQCZ9Z9UjYPkOOHvLAgG01cOSpD0A7QkBEztU
vMaCszLpZNSgZR8HfQbx2U2i1arv0ECv5xgnU02o9jczq5fieJ/G6+NlEYnohXP4jv3cKnH+JJj7
biXu26Po7iYJsOMM1Fz9jCGllr9pUbeLMJ72TlMzmHSDZ8um/ByKGo06h7LqYzfHoDQcPsX62CfE
xcXz+QM8x8vv1eG2SwdToN/eCJ4/ewJy4Z/2DtSfi3Pqu4w+7WmKtoR347uc4+u3oA5V5iXwMY6X
celeFV+5jV3t3BlEUWp5ExMl4OV57kejWsM61dCxBxApb1W6tA4/VURLlBZOFa0jHHZ3o6WjtSBm
NT9t/agoVeCkxRhLeLbSfahy9MeLoWaKbr1qS3AO6ZBaD/7bwoLR0JlJ6C87vXAsvBc9hqUVUYTs
7BR2TzfF2dGz/0F9LEA1SeuOGmLVymMukmXx2mVyvgS5N3z2FlRyZBISeW+0j3DgUgqt8bViz0ze
KjDpU4G/0UEbgs01vJ9yUTTu/X642bmxEukZKPLNGMFzZwvz6JDO/WlzlggsV+ts8YdtRkH1TEl/
pVL0xiJlCiigp2bLUu7GdVdjghYmL/7BeSRHf9Y97UQ7qPU12/E3ntITn2R7BC9kFS4817sPozpn
cEHbDNuP+H4oyosCx/hs5AwDBw2/Qzv9KHj1AUUI0uINinMyxl0hrLSdP3UsCd/Sg4+n4QR/wdIF
F3Wa4fAPTle7Ngab0zWL8V7g5xfFyFnviXXZRtUvZFp3IAjCMdDR+2/RcywpyeOmiuIXKQgeAAqK
jqh+KfOdrYRBONRw+5YQu6OexpSTPm7oaTkeF0pCWDhAG0Q2QMrwnkoEzMkvmMyw4O2/YYFikF7N
CEE6BN+crvfKjDHw+UDmM0clvYBsQcGCBZapIlCTeThdaf5t/QUbyifTk2oCSeE6Y5m089o9Xhhw
it2kBJXUS32IUxzShCGtRBHeLeSkTTTgXhr7qox0pdOos4hi11sg0q2+9ppWfzSiGAjh9XJmgqmK
RLcHyNobXEPKxhuprLxxZSxWQ9itox8pAeYzf/vXzPyiXkITQ4bZ7lHq+5rvyjQWythhDmx2EzeR
/tiU7p3+tKnVllhuffx8kNnN60/V72LKAV1BKeKh363bjvo3FxVPIE+wYmXrG7ad3Tlh3pwW/llx
CZSrzhdJt1hvMETZAyLFQMQBpSWxwTSIaBl9XPSvzg9+3LTv4u6I+Zvllnpm33fnZ8RxoG4wnCr/
cpP6dhltLdpjImum7iJKxL3QOASkBoamkEIA+uTbmwQlmEblH2q65NXbiw2paR9zZCFXf12aCkuj
DElElnCJsM117OtE7WSICgmjcbNSV+GD8XlSL3Oqb70dnxj0nNGXAl8syPxtSuFlTM/8LHX7b3c7
7I8bLqvUbpMWr5DII/Gm/Lu+SayasS7PdWawRM5hQF8z07C5gCopKhfEEPKM/Axcv7e7moykolbk
RdTgnGqFv2QCl8Yim3M/XkEeLQ6HQgfAW2pp0x7zAazl3VJgm6fNJyzN1vI3wKA/Yw6nwiV4GTD3
7SIleD/4UKvtY9wLoGFl0/Nt2J4yM2BKLDKU7cvsKqLk3n0QtlIBz/EwwuKcTu5iC/MrDcTLPp5Q
5P8OvcQEOL5m7Cs4X6JPY9PSWWuGUyTdZB+kO7oaGzK1Vh3bn6u+3IhrTiSUIXhjtSNSC2OJNwTF
mI27eUnua8DcWlSAnvnaRGktU8VA5dcCFbokfUCrlk3cv9nMEZnMJ6d7YmI0InLaFSXnk+bqzg2g
pqrZWScgwDNaGNX5LohbW5TBTJOuq4GAG8Cmq+UcdJQjkKjHOg92q47CRQbDSavYo1jCYQ7zIKSW
YvR9laX5pQsfhDfDv77vb6q0VhfJTFld8Fh2s9dUy3U7riE8cT3Ug6leGWdnkBz+Zje70q81lW7m
wHm82c+NfTncwYha/iMMJ+fn+gQ+MU+amSJJvufuc0K/nOEEktfQNDHMzJkYb4BeQICKW9Otwq4G
vpbwYoQYPsYflnIyTQnndG+mpmVJinktB+6txadfaCDfvD9EZxVPqW55it1HH2tXcb8FxU+fcBT6
oUAe+qQd6JXgjGoCBmu9twgxIInnitOMw+OUHjG3J6ZImMTxxVkeoeL0qBGsB2qqXRWMeNt7WwOJ
SiVqc8iYF37JPvCDGKBcIervWRfjQJQljXpuovbj0C5HyExoHndS5tNDV+YUe9XzTdrellWAZlQC
z5puAysLnxNlY+vGmOL/LickCxGObImX0IZfjWwGSYuQRPS8OFq9g7inBlQV4V9Dlkrjml7u7m3z
DbcC9WRv6CQEEY3dyf0FF/m/FkZAYuOeUntRTfTV38akg3/UDfs9o2Uv0gOgO0k2Hrzy6RzOJKHb
SCICAvmYPBTOalLV5NqC3HgVJGdKwjmvPnHaMWRT1oYnQLvB/V88/9K7ZUvyFLbHe73/IBStuaNs
a3x3I4qzMLFZj0KUGerXWj1AGc7LHO91Oe5YRJwW6gFcsWcm0D3N9OF5ppYvw5X4jIR8HWiUEtYG
IjnLXVxVOWhrl7VLGAfFwSnqcHqgy+k3vWBx+VRCdXtqEJugd8I2VzCvM+WRT8Hd9Lu24npZH89U
JWxlmLeuD+b/QQ+IfX2bLYat8B7UFpfK9QMGmb7dU9Rfov5+s7hFQ1BqIZw53MGgxUHBzZ3eENXU
BMiQAhjJzZYypgdmTWiRHIOv2uXlrgZyO3jal84ZeMQZujD8CV8o1eUP26Af5SrQkO97d1ZO3Exn
SM+ImDs3lWfofRYpxS3xjmP8f9SCXltRX81fAy78mzqPxT2wdpRhh2t3c3LDKHgG0sG0mGTm8wMi
TE9kf0ZnGPzix+ACAAb9/Uw4zgLKilrpMpKPNvN9R2bgdwPztQxvf9JtAkX1i3icY13jA6BLgF/9
o1+5i3X4Y1Dk/vZnRRSbuKNM2jSB5PlswsH6RPlp742rZncqz0nMd6Txeu0N5SXH7VBUzKza6BIi
9LqgCm2ix/5CvQKcjUICTwm7kZqeVFeQxDfSrrRkw5dh0UEdJ4rDGQXTbiNjzPAQNh9HHtEgcjx6
SiV+aMIo0atpGVlPYHPJ/v85nN/hVwAin1wRXNZKzbWkrcuuyvA7YPpXS8aIWER9dxOSiqjfjVie
Y+mK72SVdtEnSTDAj0S2j72i18AoGOiE/gxxc4DbWj918JOTMpQvgMhvKzCcfiC3u+dFIfhJ+BBm
yrJQsPGiXoDL5NtyOMldKp9Rt1BDxjpNP3oP8E0ayRnXeAmF+SQPs880fW+faduJAqLNu7WJTmJc
WD2cmUS76ol7XhPI+vKgzT0zUjWo2HIGWEJfeM+7CHTE3vBQ1wzoANER9dJ6DF5NHefE83XOd0g2
hdgDE2ba9EMh8oPmCKp6nArCNIGGKuoJ3E+8KxMVGZVaZyL5f6xMPyH6FD/fdAqojtDpdg0Rf+gG
QWYTL/eXWFyZlOy+bNyK4VpFB5sslvqtxOwT7Xp1GcwU2Oy3g71O2wqLp7IweEUPDk49nYiSOWoT
1MlIQiAinUxgyiSlhGM/Zw3MK8lgvKZF0PUhSwksicfUKW5OJantyHiJaZNwm+9Atyj5IFDd2Xku
VodPywLH3anQOwuzHWGNJIdhuir81GUVJjmAk6MLuShODQQ+pM+SI1VA0us+8GRv8xVOAX8n1WyD
I3jRmO5dAC5JC/yslr/0GS2FFQP2WVTbE62ueEvqus1tVhwJbEU3/BjVE0TV/Xq4UMx91zoH6EaH
7bO7rwg45cjuCrIzziuNivt+i4zOADSx0oGyCRQvMvNEPxhZKIBDD0sAh4tcpoT4mpotqPm2/qcD
G9J1fJqNeNA3/qrLJjX5RKHHzRC9pujHYHExRdY75QikAeKNKsUOWgrQe5HVmGqaQCZFVIxZoxWl
zMtybpNj0Hu73/ClMeh6XBfvuKL3nbnib8lpqOIEorx+mhjI8zhF84GWRkm0zwmQ6qAzQg926Inw
7OHpgbmDq3b9/5CMXbUFmaqQ5cGQdesSah5b7icjIRvv/YhI2EiSmFjZZM5OBFAaiXOhV8EyuHMq
/YJExDg5EQd3IiS4UVSZrnfFFZx25FzzIqX3WwpiYgBTAz12iSqcC0w7FcJ0CQRvsY7whso+z+Wx
+jfb/pxzFU201hs/QY0G/KeYuRkVvPQYDqNMg76TFqwJSUVPhfSG5B+Hf6kbPvovx63fpHp9nAn5
MP7lwKtwdpufCG50GGxYgSPbbhU2N0FpJw6pK/aaaQXQvOvjpYIcMGLbEcFLcLLTrfdH9qofT7tf
P266QRTasCB3cWriSYuDDkibgPhOmjlhmEL18gIfHzD93qqeMqr7DV3/G+rIXylGWYoU/gtmUacM
RmaUhsASen1Zh5V8VBTsaPwaYhNMb1N1dfYgHo9L7s+JnYrGas2HC1cQpoNucU/4RSHNKnM60X84
5GD6SLSvuXOb1Z7mG5DLaMPjLJwmJrIdF2UEpahXG6747rxhZf3Xw6WrJ/gvnZ/3DQ0Em3o1rww3
WpkSOI3CGLcQH0TNCkJSmAccKs7JPfLc0pPG0HospaK6EdqhXh4KDiRBV3cFauW3yxSxK/1oMn9f
3Aj7e8qszobYXF8cUJw/hlplQRKGbgeB5FTZqFmGUeftb4Kc9EnG8LCXUYsbppE3nxaryYk4w3v+
rkMUE1d8pLRjuM2lB4b21TivjBs7iWZf7KqcftODBOzIIP3/g+NGSNNwTlHsTq1SHxAsRAaT2Mx7
uCuI3zd25KUBp6hC/499cNdEZrxwao2UgfcrG4Uni7ofa4IdnqUBpC255MrewOB7boldqObSUmcX
/Ad7ORQpKFJHWyc7fdQqUswyowihwLbJS1cdWQ8DNUSX4/VerSY3xu6OpY+t6Fa5sA+S6Pccy8h3
3ei1Jmpt9lviOfzl8O1xQTbmFyvcDepvlH/MnJmGs3RU0AaDzUJBc6k5b9/kBwZe9dogwJK+L8Zs
JQm+1kYLNovH6G9uI0TtgxaYvJn+Cyhyhfpy9gv/ybKkUfTwGXG92CaM1wCmis9m+ZqfbcskRJFC
y9GqCWALTgTAaCqEGqf+2x9ZXO1yd9dl+WHDIrD+7NKoDmfzeRHXArayavt+V+LLmaZUelwHNbP+
r78zdsTN48hdFfTnzZOqRKrYvCXrNnJTZwlQd47xhlPyNn9j9dTYQ7GKxjAU+HxMerBwbqKc/axx
bcy5c/Tz277mnbUSXwEE3cj1Fkya1EQt3o6dgTojmAg1wY0J9tEFFVqYZVUOdAVq9at8x2Hy7drU
tN/8fyJWKfwWw4EMip5YfmG5Noiwj+4ikygn6oeQsd3hqxu0INXD52gCkQRYeFuR2Kz5uj44oSGM
qc2sU7Rai93ToWQZb5kwc36wpae2UOx8bttqDxKE6q+vGC3yfDmH6DpqJv1+gF2JtbnZnjZJQ0My
P3il+vqFtbzWnT/aR40crOyWF+FJLO/7eU4XMX8KKF02Dm9pHD9ecGEAiXG+tmRqCbKNcvOb6pMb
TefrIfM7lJdLorWDAvrDVAVmnw7y1WIsy39SC70cYKLyS7K1WALjddLIm3kLxiEl7Nt6su+EmCl8
b+P6Hr9b8HvMjDJO4QLwVqQpsGACE0Rx4U1K9PFtk4K5IYMyvNURgC/pE2E7EAml/Rk8ieAnKj51
7htisbJNMN91McVqWy7W0hk+QNYw6nAuxflgpM63YEXnQkmj1gMIfyHGM65XcK3Q+yug9qNrW9D/
xUWzcr3sPmxf4Y9h9OF7325/H/YN8fXJ4xzQ5URPROhXwqSOzqwiJy118c9l1ZOU6ztLku7nLlxX
ULtov70WgqV7uzVeX8E99KKL8e5LiGNsdFvakCTP+tdX72aR86M9E/QNZBNbkgkMLluUyJnAmm+5
2hOMcmkj18NM8D1LAeenRAyj524/pnrUrF7Ea0dYGKA7XorHWrt+A9pHaFAqueWYJD43x6CPBKzs
+Y1L4gJ/Xv2O4FyhRW57jxwErtVeRTY72TQ9n8lnepj5tASG67W2u+3adoKY1CPMv52JlRQpU9UK
YLd+rSXVnBHkgdT9xD3dGZGD/NMU911yeH3XjUmRhdoPdMko3bNwQ1bOnw0Xm9hwZTUW7w1Q/n7v
CjSE2CXPzIULKnOmLRjpgm/qnn+aZzXYnnit6I5DaHUPnlF/VfQTsXqXzqSrxIOsFD+XnkFShdW3
9iJ8dFUBHN2nhNDsBBO4zwf3CnD6GmL+ibmX14j1xGEV/gikF2XM5nWb+UByioNnwy1KjR1u4OZu
J2shpgABPrZ6xIGh98y2kX0trU13cFkki/ID0mh3eqRfA500gg0RDPXYe/TxlO25+M0Lm5JAGmEW
mu6pQz7voHtrSjYHVO8o8iCixubt1gfxge4zg9WCHVvsuRyoRXfVOOnI09SS3lFHz8lbRc1qhqTA
56sOJ46kh3139ryjVu6XeClMkk7s5uvQ7WrMuyaiW5YLG3NWUUpeMLcnO0/gVS7GNEwip3VBTND/
0g6T88ljMU52VZ0ABvbfAZdzooKNR7RUJOIaAsqdNV/tOKJ9wHRzKWFgOT7s7Ejz2kP2H3y9pgib
sp0G1S7AtRlO12rDHVKDTrhL08FThliTMXwSWEGtL9BOwl9DV5G7l6obclOqAhFhCqjnk3z0fbKh
k4d5l4IIqVWUQAgiP0MKDuDzT1ZtrR4jwD9Gc3hrzUJuVsAVs+xW6vaptkVzCwKVnMbZvOOWUaMg
+Gme1iyMP+Jf23rS9C5AiCM2/2WNAAN1MF5X5be2vj8Y/KvoScxdKAYYLRNpn0MOL0Zy1Oi2vuR5
PN8bSN9F0sp+FnICZqcNCDgJKqUT6tnP9u3exxFXEUwvuldHWwaj+HHvirw92Z4Ts8nb3Dq/p3Y1
a4Ty9Orwwg/KisS6GiR/18PjzBd4/l0Nck/Cn9zRYzbKyXFZcoef843c5q7wKCO/oN6xlbHabwyN
dquwwAny+yJ3eiKlcItCX4oGpq30thRtqsCFjU0CwTQOLsiB8CdeZ9rzb+Lg1hAgti6DNJulgaH9
uFsN5YD/8NKmJhP8dSdJEqGqXi3VyW/0LKerCSnz1mtnw1rhWVmkXi7b2ISTFN4LnCazrh1FyKI+
KW63QEzjroRKPjVWtrlInJqSoBMAYcC4NiXX8DoMRgfbH98izEBS6RAxnvFrv5VN9RFAJFfbZrwl
9TsD1FrNzF9++4NfiAMWh1HTVAsqfrUd2vuENyzDSnftlQ095Y5qGT3Y3gXbX2uDNXvoO4K7jmW3
QkRw+Zu7CcdyEDaE+rLRdWkljBm8CruSjOB1A6JWTk6+bi62DCA4dobW/nWirr8w85LX2hC1Md4T
UXge/y59bCBwJSQ6Vb7E6JqBQdyKwxmRiX/XKGmqhocb/hI+BHEok/8GpNDd+Ww+o6ldB76oRTe0
jsdU5NTzh3pic4A80eXhRPxnNEss7MO7RrJFahVFjHKnoxIKMfN+MAi0La4S8er3CxPSHc0P3/mM
WsTCAUd6T6bSB5jgrCOvE9UXpQGJqKoVlrxC68RGjJmsHtigFAox0YS/yolSGdSxMAAB1Axh8E9f
inyLlZamohvDOa+VqBQEDFnaZn4/a/QvP2d05EYWwptd9rUQAb+aDSlcfGxwd+575RgJEshjgz93
I8yff6toUX8QpcdCgXmETWNp8MGQ0rxrLBwRluM5YNPpqJSsxZ34hYWKeGDGRrpmYq1jXbrWjItp
tnAbBCJS5c+2Zy8lEY9Y3jLzEWqRSA8speGkXkasL2PERDbZNX6G/iRtTWIgt/HwuwW8FueMfy5u
m7znlPlKBGDB/P4zmJkZPy0AdVGpITiYzj5c/kVA+uKSCnJEF1UjV/dlalXtZtuw7OS7M2NLH7BO
87Np7Yv0zLTnsyA/j8J14XSq9Ul3VqPw5SYnRVq+XKmUMudvord4X6JYBdiviZKTtftc5EgMHHr4
UyNxtD9v3p13tVxuz6iBx2K+xzBXdZXAy0RwMzJ4R7I/lm/uIDKSoTiiXJ1s6M0jCO1HitvCdM4M
oZLMRHhChC6fyK338VwB1A0QVsoASzURP35FzS2m7+UjMg2vZ7KlOzlomGMf9WWf3HNWjgULl25T
gFp7rEwLFirxqGEMEMwH/l3A6nOKs1uIBF+gYSgbObJVuFDTdlm05Sa3xCQTEcEs4PUk18E2uEc4
tuq4vs1AHlrbSYlxYY3OYsPQk26NVzCn30uVnrRA9xJmqFMTwuHr694z+Ch0Mr+uP65OtC3xa2Pg
PUl6BmW0c3xniO+Ic5+qNiJidQqx6b7jOundKeO+nuubSd3J09fgFenXbrBl1OpXVewT+zBqH3B/
kfZZlLaQQDudwyT2KgUzvhr+x8At5lXM1AjStin55Z3fm32VGXUerq7HCB+7d8fqhfgacEAcwIEE
KwkcT1RqjbIar+mUtGvSuj+wK5p1lrL9PbfQB2EGky56tSWHvMLUI8ImnyQMrxz+pX9vObXuQki4
b5HTdsaAAJfvL+BtDachL/WSUhp67JNDiu75sIt8rv+WD7izBj4Zze3zWveewmojjgkpOhyyKGZd
s67HzpLwmBHF0Ec4eMyMNJquUg1mOnjhhiA9gr0zv45d6yZg6xpDp53LmUvdMlv5P1j2U2CgaiPR
3ro9a0LEOhAFWKPoNddCI+tVSJpdacluejSqvgxlv5fRP1Ogjsv/9OYdHoj5S4UtUHrxm/roHT4c
+z7OD/E2KvooNGiqknZ5Uau+oUCivOGS1/qWKrnElXFs5w/UI1bah+pi+YyKdSjBTzonpGHtDoQj
9dPw/aIkuIhra79BX7DpfWJfwNfCVWOiTRU+9ssLPbcIlppTOrY2JF5ljXChEfywIfV3gV6mVT3w
jng0UgM/UaTDqPEO8S4p69CB8Ksf/dTfn+ifqhAsAf6LJV0JBcEx/QCWgzXWfSNoYd8P2jXxMSlj
AM+aof6ooNlkhgGPAVnlDV9913OFZ/GkQA/W5RrBCEIG7ixq2yjkeIe9A1bfmFHyPzJOwadLyhWw
FWUqBfVsDE9zqs6Bli5Qwz8V/E55mCxmuqpyl7l4skrVDQPQT8YVo7kkFubD8n7G0fvA1sfQRkB9
+4dRTnbLQ3rS2Sz/vDoguDYzOrWD4icHjOsJxBVUd+b4ayMiF73s1soFz3PIr1KoJpHvHRAflumI
kKPdjIEoOLDVEbzA0Tmk982xpUX1TDsuSKgxDXtG0AG8AubzG9bh0GEU7FsRm/aEJZOsWogQMk3m
W0cRDDkoZH5cnqz+Y4MlKwgFitGF+xoAswukazAYVYr6wIDT6GF8GUcJ7KuZviynpMNhEQQeCFnk
rTaOfm0MKtJXwUZ304IvHT+ziPE6VAQGILKN+XrNlb1qshPU+SAsJ2m6nCy5Iom1pH2VUAcdG//s
TTuwei0tmRcXtuoSsXJnIK6JFR6KqTOQpDev6vO/kWQP5EbY2kBHNWRp/n2BY1w7F/FUPqGX6OWU
x5LV+eS53+kd2DQGRZSzjD42TbY4iOb9GSZ+/sLGO+oUsEXJxiECPB5Up88aW+OYnsL899bJrV3d
r5finai2DxZbvua1hczY+ax+bKP2f+dZiAoiRticA6TD33Cw5HALqiQliiCiywncitcEcB6uUanR
5EjMHiyXXayHk4y9p/JNT3F4zcO8WhnObe/CXADzh0o5yTwlMa/4B1MWL56bTZ71rGgJIcn2tWyO
fTR0VWm6oIsWmP7tVtoE0+RVmZ3BIP9Lpxt/W8UNRmxVKVGoID7tZ3oD+feFSdJoSkHEk2A6iEIQ
9BbCCrvZQKE5caKA0cAu5HmSwlYxkrdE3ZZMj76cvJiB1lNDD7yJu9pf06zUxsELNz670x6+lo5e
3jBtkyxysBAFKeoJr1ceW85VJBY2xbG+ZIHzXbr6zf/Q1SX6vvodr2LiLphiLLXIEspgWAgPIyU0
iLIf/wUPU0Tx1P4OHsQoQ6BEblTc/vqbRNfdT4Mo1JseXb2dYSlcwLeq2nVo4cSuy9tUcaQWu8q+
EhAxFmKcSVmkd9CwcoN/m1iPvR9vMbKZ6T049LX4JTgKvO9QaH2EY4f26ZBwL4kHFzv1R8gCgIj5
IzFrGtea2lSx6XSxeoj8uOW3404VcqcHoO/JFDYBby0mrEGsrmqu6/n4A/GQ+dichHyUI2ZxLEyZ
k7V+sRLo2zdfKMTW8qQ8Yp1S6L3rCIiWMnFvkxqGSPzSZAiUpLrBjkfs8dobWG4Wl2RkI3TiHGVC
88VHLvi12A2Xn6YQFnQFm2xEcPdk7N/azYuIBFEbBRnxqaBil6e32gEC2T9Ddjep8WvbMRZOYGq8
RGAhTL2DmyfyPn0u72+vMPdACL7Yt/8I2C8JwqVsg8VuJ5rpLOzpVpboidYIynoxM39/0jt+0PnJ
+AzzVSuJXE0PImjWMXQTXH1MDCVcowSVrUKZHRaFflHFGQre5gRaAB9diCC114VDNdwON1p/Rqiz
4x32E+XrRJHIaJ0BnLKQyrYizshlcjEo6eR4ObXLvMZPyBXD7QmBGfQIaE0ZyHWYJmRIo+vqkYzn
M/gpGtgDVyud6gTXPRooyvGsFFTOUKmUaEzZPaUOX5qOcv1hP5rBMWOEwx2LgzHzqVh9GIfL1joc
Ys9fE5PKo7rYqJMdHET5suQphcKlMiA3T0evLE3pSX6bDh359XTXyJDInAj5x+B7x45EPTc4Aslz
f0dmA3OmmbBa9vRDyPAxtGSte1csbHrE6RKLJpOvWa2e9oCqUMMGWABFr5jeBMJJkwH97X47FCin
jIqTLT+0pmcIXM8agOohMdUpmAXajuhmjZ83epV2kjhAQE60A5zd40k1e+fxSePlj0QiouqFNKYr
te/yP+UyuAj5EhBO6QNILI6cYquJiYQj86wkCN2NFMU5HFYNn1OMQBdthMM5q3PCRhEDxAMYruch
tqdOiqAi4h35Mpdxd/Dt/bp6yskTjUdf4KEpmncrNoIXAFq1AcXwNTcGyCxmc3UZou65f7LJlI66
944UGgmbrA3iNtfR1LpJeGwLqIGmBT/dvvN19TLdU55LL5ufifcdhkzS+Fh0VtA6HYPauNnIRgqu
2Hy+D5FSkcysquGQ/TRSNPrEENQsJjI/wUn6gp3Q+VqH9YnPnxrI75obZRpSib3teMkvF0nheTX5
Pjk7HXYJ6hSzFPE5eQAmKAEmiTBSErHN7YFTYQc70bY52Ulz79/cipzopZxi3ymOZmz+0Dm3vvMs
GrUL0awn4P5CnZA/bJ4/O+2VbWmz4CcPBILBO7Vb4IBrhdoCIOhv81Bi1QZze417iVsltUXhDOmq
6wts9hoy0Hh5wNTYmGCQBvxxnkRzgqwlFDzGgKBojRGvgEe5wEzfQupVJsSPb68CKCH15Sgf5AlI
VEYiNka94oB0vgkVzkUfF+3xpXPErcp3HjekqyejhXih4Q6gD4ZhaO9e9JT9dl6p8EB2LwfQGPsQ
Ro6Vr93TWAAMebiWFjpHaMEefTp88pWEntqsg52ivjGNbE/oOW9QYmE3hcMnzZTmID2ddaCO+mqg
S//g8SeoV6g1uko6ItvPkeBqYrx/tylD3qkr+qnuflpgW7hIMmPGVOMhCv51s8lNuPETUPPAiRXm
FEh09XengPMg1oHOudVflXN77hh8ibwZthvnr079lIu/QdyjZthFRxrIi6IOF/aDx9xka6wUpFhS
gadm4MYX9F5vwMANCGBMzzRkcLTj5Tt0GsslP41A+HcITyeqsdqCKyvEUof+qyBxejxLbUNj8+W4
MiaZViARdbyzWkaJZKAuaex7GTyUfMgR/nSNRxMUbAHQpqgIPK/KcpP1OLus1cbmtFC8ja9GijqN
LklUFgSMEiXrAgiAHIPNlb3cQIZid8oIGWA5K04laEVXV8FUBEtxL11hWO4mU86duFMm6+KfaSC4
jMhSpEs3sieDfrbSG3jYC6ZSmF3D6BD/iU2AM0Sv5pbUdV3IiPslrmukFHa11ONzh8Ay/aRB/NmM
6LCD1iNwc5tH9WlUYROQ/bSVlezV34k58iG1IhPMDHyhGTRWFLUGWz7aaBCE2IgrT213wPp8KRwN
5Wq9u03Ti+Ja4hthkgxRARLwyiM4K9xdHL8Zeg9qmwcLsi+wy6f/TdkaTlW/Sx4IhPrb2S1HsCAT
86tsNJxbyrlmeph0kEmWLl6DzADImUg7O+TaN3svFHZYgEMkUT3VMNClQs8QF0qNo+0Pu9p36RtF
qH2Y4rSdJ44xPyKgwaY/qcfBQFMin9T+8FtUwH83b0csQwqMyVumugenJMOJW9q6rHVUNKYrBsNo
c8/0ZyG2FLMtvfRcMP+TxCXk6nZ+KImnkyKpPYBrH1WDmg0eymAKgM4rCsrzR/VdphXg8XHCBjEI
DINcDBGsz/D2UKvzcfmgkdqGTlrBwdAaosDdQjypQI5Yp0g8sTixwjoeO2miFT0nlIrWNfbz54kK
fPZKn/RdQvJDm0sVlvV5p9mI2ysBufCWvOsbRZU7CiQEdE83wg6UnRAKlVPoPzZZFi/YLHAYJhGp
IaA+wqUw2V7K9ITBEttGPQfXbBKgwi3Aqd1MjHunDsSNa68+1FhppAB8sQaSTxQOESOM0oWviv/r
g53/uh7hNLFxP1R4ZyrUIFH+WDCYtsbV4ENM3hxIxzWve47kf8+11kiurydY3TGmSoHRWpfZTDh1
ukqTSDXer6H+G1p3Sk07j7PzwQS1NsLYfyuIG3EdRiVDHBHbCS3pPvAYf77dtt3BnEBrb/46vStj
FKBs0IScERsrVVFjIPdmrybYCKqoKux29IN+hzrThd7zndXSM+OkTNIGCCfsx8eTI6TZ8JMW9O9E
JE+TASBrOCHhIDQQprMGN4qeoLNjRb+C+HavOT7NKKt7bufCMmAq3uY4FEXe1rF+GY8B+Tp4qh8w
TtMUJQuQw2CWA4HJYklx5CbP/mwhHYSVDHvRyAlr9uGjLye1iSYvX+EmIhIoqnC2Iqp2xRV/VCbo
1BjZ/mqYEqybh/iGewfdbdHliHM0Aq6QiGtTUDdFs7r79qc1JaXjBlfGZGUlDJcmnZpwL/sePcIG
PpDS7FXScCHvte9FQ1mP09QLXFlNUrTxORh5Z3Kg8p2DR1Mk8PoHv3asWRd8TreXkK6hMpxx4+A3
PUC1NNH4KUpgM62UyVsildZ/j3/r98RkNPWJTCebJtimA5viSgFF7dh2ginIzpKytzUn6od4/OX/
yTf+OEeRrIMX1uV5P5sBvuSE2EIID0tcBD9vBzlTgfqMRweNIsA5iq/T9RAC0lqwSgb8JInJ7c4r
l88h/7uUM7CTQPhKe4zKIYQ+K0fxI/Ypg+9MmEGoflwoPcqE0jt6z6xxe9iQoDKxiMmVO5clsbNm
/n21sd1nCKYV86+MUQkQ38D7F36Gye+rw3w8tmhRqdf41eTa4sfooYJ8FHip3tzlTwAUEoPOiOLT
TGb5X1H9RPUgOYnSVghzefHLpRrFWeL7iPW8g+Fo9RJ6OIZVMoTKZiVl61OBwBo38VaH10e7oepO
7KeA+l2aeHcxutkaWzzaJTXEtCwfMLY4JF/tX+wjUkl0hymneAgYpSFqEUKbPobRQT2a7QPMKbRF
SbJWAyVmTl88hPmzKUOUJk/BSAP7CqJLZtdEg54kmDvQninB4ylfEhTxRRyeJIyoNr+rzUxIW/4d
SoclOpTM6mWI2Zy5umG3DAp+I7Cg8JIfGojrMXFRwFJzRgtx9yvW+Y7zOugPQNDaOYuQKURoi/IQ
M2vZCP9XJJm7qnTCK4lEP4KdybQ/Z/UaWTEkuX+Mr6vTC6thzFpDTv+YZaTiP6yX4DgMvqEpeG/a
7xeRN/Xx1/Rq1sTQhncsrNKPS4BTayLmi2hUJA6+OUHtZ2+yp8YPQ/psx4r/OnXgTxbIu6L/3vWH
cFgKsPFW0kdWQEkAtlCf7sCc76hWwd7Yhco2Zqxp2f5XNUhnYTWCYAQPYh1UIHxC+0dTZNVURAE8
5e94/9v8rEmDZN1o4BWzTK+tDMP7ZrCADV8kaX3JWCj/wHu96cfJFHvgN/yIpcfK2Qdz1V/YRtaN
/T+jOHsPK43C440S1u23yez7PESI/UT2bMijigxriDrJKilwhJbp7jui53qKTUuFJXYP6BiRtPFB
wHr9FsgT6uUrMTmlG7tKT4MhhM/Zcc+FnBOrDxVah3xBSHqrlqatSUjWtLt9/NAh/YcNKKfTADmr
92eQ1n7aOfNKQbtHk0DJ8iLLelgqmAMIb8GKQSYZAzGu75Fl2lHM8EtocRw5Ka3cmb2U1BR4f3vO
4AJpqbmFCIuHqdP1gK4qBoLOVzj4uQiR593Do19iQd1V9AzNS3jmRfFI4gAMyGi4RvCkfGFA5z7S
pZdrkixGaFJD/7s9tMSS0FiU3A8z2SNZFvnMjXLFL5ODWBHfPDucJEXz1VcBuzoBIT3+JEcAaADC
aN2cWTmGg/k410P+pClGGZ/40MJtblXhCzaO6qSpXytYnsXBxq1KnXoNzVrmxhMnmdm4B0HmrEyj
GN9DyFP3fR39G+ow3jplus9RewGfji/09N9ih8wlSJV9Ua0AchEvOtgV5YQiZYwdXuhJ/xuRjNrG
khI9D8q6gy/DfYkcWSmhGynEuT/+zNITE+OGd16xwA1HGRd7E6oo+Hq5D7JuBivSzlvBBKwKBj6n
9BOwBIDXrLpt4rQDK6OHgCrYnC9lhTRXuir7tfUGENECkL2ymtSKud+DWG0LxilhdIQA/WcJHbaL
VJDpOpFGLDGLmIJSCqy4xVUeXycxi1zrbJV5f0Qb7jGxL1MAvmGciiuOtuuwTCOMLSn9sh+Mep3u
wKoFlNP2PkyIMuWjfWH4iI3x38PCxFyYVpyWwjwt1DFZ0EAIO+j8N07cVSabbkVgyjYUvi6qYkLK
nizYjA5lX/BeCpEqtMMkmaODhrIuYc5/1y1aiL93e6nFVzoK73gGFyaOeeicfCdiIKoP2t8m0bx4
EpOrHeSUA36dM+eNE5nKMegccE7SA6VXec8yjlv5FGRuOCYHYfK+yJsrcr5Tkw+GJslF90mWhQuL
U9dTFCfy/K1aId5ZviYcd7bPxdbg2HFGkYfkbuZH0dkqGZUBeebW7UGmvoOSLbMwsCgK2peQO10E
waftw95ZHNUJElg3UYWBy5PFZa5fSLXFIKOmGuGBtZbmzMLB+9xag3xWWsFqDtUiR+rIsuAvzGFM
pHJvd2mKZ06U9R83z8MGePltIQt0Jr/KY8iZoz0ZAUpop3LxunThl3zK/O4GIMNculn6C+0jfkOt
Jpqmfro9qvbGMWJOCdVcYhxuo7KIh/SOlm2KbfbXoyDcmCeT85mdKgsvsnWH8yIJ09nJ+0fPSR4J
HXbA7QfHOYLUi/5M5/OnY61qoTPVFHmIqzEjY5N+X/vO3WGp7/voT9zqsZzoP97G/XT0zAVcm7tm
zZ+NwRIa2P1in+P8KdgPSmfBN/YnBVV22Cmtt9zZoVpPN3QCexvpUAqwwSjECXQbfC23l9iR+t4V
puR7EAq1J2FweuOgs11oMTAZw+g1UWdzwoxe7axZLC6YecPz6HzxcZJdCp+cIqA4VSoq5ugwa9M3
Rb7JabTxo/9Bv539q5zwPXa98pCX/VlYbTIQIikXBxOchTaFEhJ0747NcJ88wtOz+ZYhefY5RqHi
6aRlxLIyXEwc0EqrbFmhB60jVMxr4iXHiKfWjAA4im8mmVvHKn/suRMb8+4ItVXKfNE4yx9fpjdF
AlHOWjwjYuyHb0e975s+0+DyFRpyK3XgAQcPGKkJfeY0agoBJKiXngceo6xX/i7R2WcslcPFP8Nj
0sWhF0ntfe8+IDuc2jGnYXapSASj9Cpt8Z2Jed3C4S/kpExZiNQZEc6194CQEikokfjNy+37uAwb
0v9U+zN+mrBOAlJ3c7UpfGeuddiWgcpyMvAU9WqrY6SnsjxtMShnID7bDtIl9ZQTjOwgkYcHb8fn
YgKC9TbBWs0g8x1+S+M1l/W+eFtQeHwu2rooEHhr8mhVN3LLCsE3qNFfWh3c0znwRWlD9/UyB2dZ
VuK9N7sUVbKunMqCTz0yeIJ9jS26KpTBUcooI0RmUIbSrMQzZkoCR6HU3OTU494xRwg4M5i1GeVn
qJSYgkkxzOwXUDXRIflftdujXuXQQ8xLXhXqQd2ulb3eo662WuuJlK0K3ym+CQeOfZjN1dVj8XLi
D/QEqzaHTBAK1V9pwIxqqjdkCs6rAXLEMDxRTipVZ2MtYH5p5LyIx9c5Tb4+N8gc7HjIlgbosa1N
PgrZ50G4klnKJGz4Wyyv2GBHAZmgtbwUXS4LSz0geEnIHyXITFMgbNEdJN0YIFhwVyzFbnaECopv
0+uMrqu4hAE0FKs/f3AA4VfQBi/cwOjIPmEez+LTbjO8ayBuID2SKP0C5rJ71ulmW/fXA4dR/otN
lMOVu+t4YVv6XqTmY3xJDHIEDUTtBlCWddI+YG5xW8SL3qxJUUkpfs9URjQ7JndbF1GCHqlUNbBo
kv44E42mtK4Bm7XmWscHab6mX7VRm0KGG4ZSRBxORLRUHIfrzQW9EfYgt8f/mQ50WxzXvmzekHqz
C+/DIgNe0dacnSbKNbwQ0lFco+A4hKqdUCKXmd5CkTtqHGD3KjM2U82n858n/U974hliR8X8rSwD
CFm1WyUPSK/j4Hm092/ZiIiNiZBtBba1onSbKtoYHaXN+naEchNFD5QpeTgWUiKDdIlszslb2cxe
uspRRo9Jc7qHn+Nfq66Sp5sABgeYMeqmoogSAfiG1qp1boHN8YZXbUfDhRGkzCXZpj9N5kjPe1AI
LC5R57mOsNxLGYMlJxYqLqPh4Iy7P4q1gSbmnkqtnZBmb8903Y9FFs4EDEStOgdsMYxJTLeiOHYO
nCefA3daYBNSgHCd5pDpZJd0t1PVEDnwFEGOD5fImR6zYDaGgCf/AEd6OqzpAOLO18Iwh/BCFGhu
uptWAnC4E7UqQMmJEcfwykavQUHJNqjt6U0ZLzjfTGUF+ukSIrv3+9QSdS6U/43ayZ+RPspmaldR
jfTCgiqGbdIkuOUDwz9ri0hv2gsUANV63Htub67GP6Vb/ylzAaZk6M8L4JnLSjvABZEtHlDHx2WG
IMjgtKnBX2hZjadsLNKENONS+t7+XTXalf8YuYFkUMFxuXcT3sRnRexrZd395xiQTUyHmEbotmmi
JcJ5uHcS8/EZ0rgIUpfRgeVnWoXwWNgieFXzhN9zWiLbfRPBUvvw7QyQ0J7Ei3rG6F0ksvMl5Z04
llYEZvFmWeRzpQ7b5xZFoS6X/0GmlrBvMwIlEAJMcxIbkfkCCPATNYU/ehlwVPH1D7gzb6VfZVfk
ibkb1MG61lMM/CwAdrn6IrmdPbrs5GOJYf2bDRqPx93Y+WgOhL6TEnsISRVm8p8nFc05+6KEP506
eHui6ZpPgF54EXLu9NRATot2oZnSobMey7jmd9dkzxUzZMvQQCoQ+n2LK/VQhBldAdp6alQjsomg
gsv1i+B8t5UlbfmPryzdCqzTtEzSkfA3423LyxeQWmXm4qC1qhn/SdPt3EsWVPJW+X8jPyrcmPEr
YTArYybGaJ9dEIgsoHVA/rE0io7QfmB9l6fo+N1QlFfPCH4IS/TNVExsGsz2EbQ8o3lBgaURI36q
IfMoKZJmNuxjJxvUH4DvejSqFVTY89GDQlV2lKThmbm54GDG8kBMJu+VsleXteSNurocfyTBEbl4
/y+htLOhOW/XRXCTU5D6buEBqwld4FRDEJPEkE4sPluhAStvLLz46ciKSh84+NdYxNHiMjIrMl7r
WY4V8hOBsA11znYYfigBo5sIrMAuTav3EYrq7hc7dFb27KNpTsQ/Zon2T2bIXRELfqs8MvTn9O+G
vinZJs/MCtqxCa9OZIJKR62UA5gQOpxhRRIdSRwA1XASLUG/Io0wfnJ+gmzbD6PGwyHbEnbYfgnR
jP1RxthN9e3WjkTpCDk9j8c39rOSeVf7JnGuL9C3GoSo7yLVngLCc2qiepLfFJuU4HCOLh32U+Cc
h5pCtXBfhLUqWdqtc+S6NyxkwwDP/zpyx/i/1P7tBtXsqefuh5TyOR6xg6byJFRGOpNCAr6VUqqL
PgGx4XhUlrhSIpRcSfrvzzyr8Fm7wOEYUx8Dkr1upDDTR3zsWtEcZTpDoxDp7jWr/cw2Y8IIiLD8
IHpySKcavePw5Y3q4/JVnRjCvm56Z40CGW9iuvJmjFn2oyFUL7XkoNFVpuf9IiXMVtElTj4VhITk
KhIvKMDrsOsxtGrLIr/6XAT31PvKEJ98B6cnL5lhjwQGb2GX+8vn855zvYqj8vfAgO2X6NoXGjB+
K3Heb4Uu315/d9EyoCX6H4nPLQCzPYemFOoo5k0YIwaiOfX410jmkTQrdPiazEl33/Q4Ly4gO2/d
jlcE0k2gUoblGfYGr7tM+Eqax9wqbUG8BxwZhgPXFoMYqJBPDpVZyxs9cRI7CWakNsXUroM8W9x8
BIjNlhfjaB4bqX6Nzg1s/GY5akxVApga0wXb5PmcBYDCMUyJZfbUAmy2n+6Yszb5THofozwJJX4/
GeJSMUvOEJ9edHUSTXU9OpXT5Wdc0pTa1T7a2r+HPIo0nM3TQiI8a4pAzY5etdP57gT9KCWXWwvI
W8LHUtp68W89EdKm76pYoTMp0B5Vo7GpJelOgEatFFUKSkDrXZ3rRgjlmi9zOuNKe93fYZdceqRK
SLv1s5jLWrxFbDdwGccgtPPaveZ4uiUiFppmE/gpgy/yrUtxbB1COe5Wl/iZPGNX92dIPt55zG/K
fu5OvyRtwZg4s5olmWyd46LbTXYWxh6UIgUOj+yzmOfKgyWOj+EKo0rOCeixbU7AgyZqsaSyJcnv
y/oHUcFfxOENkJYd1ijrnl74fqFSecOyWjRCygfvKL2r1x5jJdrl61Xk9n8zpkQU5GY7rglhLKuJ
MzBR56EzpTLGu4u3AmpkL0/MbJs6rYpVkBKiN24M/CRZXfXzbBG1E+TEiBOS1SIWQxbD2/21rsJr
iyqLyZ7a/RmLKX5cSu2IZGqTAaU2JDBx3TioEo7I9gVTkaMkz+vylbj2g7nsMfAvo8TFAtRpmCnS
Xva7FjWKMbJJw9Djww26NJTkqNSgaKwdNx8jwcxfQQY8M+3pS0JocB0tEe2M5DYKYlys2nfj83lI
ZdGIuU/6wcBSzStYZ1AZZMqdQv71P+8V6NrhfuWKFXfH1I/RcrT16w08gJX0AimL+o3xUu+2Ee9n
8DylMaPMi4uWg5FOo51UyiZvZfMC92451GgWMvNd5oJSuB+7m5C4tThzsyEaqiH93ELNIdE7ISko
jq3hu1qlx+vptiFbWxj6hZcoTvOom7Vn4DE2e2KqadOpWsUJQy0jq4v78ACE57j16Exg+axUQYvO
mAHEKoBWaRAmDvCj5vgSwvUOsvTS22vgkqt4k7lcqqWd15MkcLrh96CvDNWnIWlzovnhYtRgfItC
r8EExoU8p4dOL7kcWeThWJ5cEqWduKYLrYGTRJN4WWbIE7dWROqJAk0jm+nk2oyQs11NJ/UDbr/A
2pVk8uvgw8AQXKmp/yjGNBUTaM3lFlH1hmdFnWysZGUsE6pFmtKRK85emEcisF9FPd5D8SFK8kOa
07rqMiTPEwWeGHfNGTVOt4sTzTDdTKDs9lMAJfNq8DVnGj9OAaxCMIz6AHI3+XkOahdGWWG3iaUX
gVloU1ZFTcA1oMINyoJOmgpCAWIeHtAzS5WaE3Bbal7lGDb1hXaDqkMKm6oUk58KFLnFuRx+Gtkk
cRwiC06JWKhb8+CASDXkFr12D0WGqLCLUS5R+X2XZ4Rz0QZs8WJeoiFPnLXhdE4G7+t4aOpMdiJP
O6UVT3NfGusdkLdv6tR6X5d/AMV47jJ2EjlZpoStOVYcsS9qt3c3jBpz6A0Jm/LXN9J/6MfqSmSf
huvzUpwxYX1DS35QHm3Oz8X0nsM4Kp/tCEJRPh7/XLV8+KfRBchrFoYGmZd5KXR1+L4AiRWqQtlC
5v3V1POcfDLeIePbW+nZbCuvzc1dcAt64UNf5dfcGpimjG/+FO9MUFiScXPKIREmmVLlGoSTDGcT
ckoeVWu3A1UYCA/xaNtCoGSW3amr6LIzq26DfuXaESmqve0/KdhdzNyoIwa0M4C3gpuvH1EdwOzU
c/d3N058zNkMXtjjSiPtOzU9lScBWP+K7YXq0xZpHHPG79OTnHEQlMBBo0PduB/AS72n0bxWVFio
1OSB1JOhILlOXYM/4ck9hRvhLdBlXfOjjsvwuCkXwAh30/jolDB40/8a3QoGtMAksSm4yn2nOJeO
pIfN/Ky0aU5ito13Xf2eJdAG0v0id+lTpeLP45EIpodUHrWoAUExb0Mty4zj5/FwKBLVjaXCSyPF
1rYHbM9s3w+RqRWxrDcSI+ugYAbq9bIs203ylq+YnN/UiyIkyBxsgKn00jZHxhxVAQfgv439qFRh
fFP2uUCvm+HRjqedLWaxx+nrpaQifIq2MIwrRfS8pNQvNgfHll/+kosg9grYbKi84siBd5R4yJU5
z+Tp52ZzmKusOBoTS/hpP6OIrBH+fvA8ITQ+YyRxJ+TPVPhxcF7HiLqantECrm0NQmRsIGfpoCou
d853gOSffMWQ89UcCvoZAV9ghs3XJasR181zWflgPSs2lGbh+9uvSiv4Rk8r4mF7q4Db0jWpkgyt
KxFASOKDUgaJR799hfqlj45AcrWqB+RDh1O+XnHzrKX31IllU6ml7gpOOoBC3doB7wHwUrmkdBW1
aG7Ce2bWUFpcRa12BTtk10BF1WLC74TcuIEco7iGwZZ8ZokX9Wu3MPbz74NS4PDvnYG9rSgmlEQm
yNZu8MHRLv8AUMbX+WqdynUqblwcbwz2qGIsLfAJegW0MDU6/qT0zhOkJgqZv3vFZfwzUn8Eto59
wSZn8BtBQylDgeTt3hXq8nCM9PMzExahADGJVbrCGhi884Ue5Y+qeR0omU0b0VIPwDt1LYmx9R76
4+kntbZHmgnf+MdxCqN0JjfWiKlEhcNraR8UDMovkefFgt8Nz3obcM1fEWWfyhRVEcfCrSuK3M1h
U8YJe50TUWEXqO7EHQOwIySRyzvjlGXThGuCGQxF+KrZ5u3t15ETvCMK525Tvd51NQTdiDRs/+jS
b8MPrdzpI3/1HGzw6PC7lq1UCk8dcUGFo3VSyXHn/cmbBJnF16eH/6/e+Tkp/QfNJsmj0bCl8z5q
cyxm5zn0AlQyYi/4i+RHqj8BR7r5s0iYrsfiz7WAMesgh0QPvbfp4DcBL0HtQpSHemZXG2QIzdJe
U9nuq2bgCkUZJaB5DAUd+/ernskXO6tAEFnCo4HqFWe1mWFkfsjiArM2vwpVLFsLR0MhwP1vAkKv
2edXQdP2i5Dq5pmRV0acb4F/5k9T7dfP+n4k+7exzQ8J8u1Mh/MbfQaMFzsVCSb2RNHNnM8fpR3U
vbrn88CGp1cX+7KiZo+RRnSRyxyrg68Hdz6SOWoxhzhrQHm5vIg8xYMi3XXGlxayTNH4QDLHu0vJ
pfT+dkHRYr0hqsMTQL4feVlUuQBDlloNr/+FdZISxNvSsK4YVsobPfe11Nht3q8gRwLDQfXvyYGN
zdChCuvbkefr+ET6hw7Gg2XHat/uQNEy3BTP4zbx5UIxFLAazaeSfwBnJTIvHwwirY8bNmDnJoR9
BBFQWMxwzAIbItEEv1mEel3Wp0NkRAIXpDZszR5ebeLI6qiOft7w/5EjTyd2X13rVAnCkQqklSU1
ZUtzjnW7etTPWMrJlPyxHxkdCtyp85JwTi8jiV7AGi3vl65Ur1n7yJ8TClEL1fgo3M34zg2OIen3
lnyhQEEzsX0TDW/PCDDf9/NkxDf+BVOaxaf2Qb3tiE1TJa+1/XU7122qpQcVSCCVD9P/zUmd0ZwA
U90UuxDzsdqtgqpXAWUzdme3fos71NVxchfh093TqCyxI4E085+qwDzdQ7Hda4UtMoiUS2eziAKb
nQriDBY7SI00bk1XS6OsnrnT5I4KDflOrwtHgZmYVRa1fG4NG+LaVcDCOiUwAmlq3gVeAZV49FXz
R/S9Kn5iE23+aC63g+Cvp42Y8t3xr+Y9S7aDB+fsY0lsdrTTvNWSwNpPkRE+nM/NfNxLt1T9rjfM
HN+EBl/Fj+7mvLwW898IN7GEw3/XOcD7oQ6IvjI6clL69xT/hnhI/9DOZrhy3kZnxV91+VMqPXFn
ll9HVjL03Z0f2y2/xrn14exclNCfZaPErqENBZuL+0B0+ip6CYl54wmJuvcqNCpbxUbx6qPOrzDe
8IGCQRj3CP5c0i8Zq4PXaVfY930ACW/3PlxDV/j6RmXObJRUKFZmwSCLZ9OKQoayZPs3NCD0t0ED
Nrr0+4KXh3Ug+lcqx02QEprUmtIdckOrJnLSNuuovK0a6BGUWo0/CX1LSnax/bE2ZsDLwv0xtcts
eDIVPhJwzX+H7ZPYZzKJzKMC3UnhgXqqhmIKG3yiv0td1l46Po6a3frbMzUCOK8ZGTq4q9nwHY9G
zkOq9V4jtZUbC8kiuPuTFlXzZYvVd7lM07kZRu+tkRi/nXKwB1jL6TSCP5P10i/vGS8UK7ckkWUN
lRpIGl7h5KFpU2DiVMvIhSjeEtjmisU3tJlOR1A6gjuCOhMWGr/Jyk3O4P4RWTmNoi2H0cQ0W06U
rFYLydhw4AStARLfgTGenY2swlkL+JF+kH9IF6393bkNIhZ1FSLOssdY7yeuLo6weFBKIdeEodEC
+mQpUi2Y8ZBeeYEkoY7BkzXC5eWEVhe+uscOOCSBH783FgtGnOntjFt9eAPP7cDIY2FByJPQDEnA
DMROFZZ99JsUehFsDHXme+t+g3euq6Ae9USBYMJbKUrBb9agCzvd7tzqJg4CMSzlUhyNoj8iKfpY
veJ9BRiI9jiJB54eMTsYlP5VlH5lBAv6pa+jT6h7hlvu2znKhoNBpHD3sGWHyx/7xnx5D6CJ617h
n9UnexToJaZ4ReBrCh936ZqeZVnCHLbXzwnN8e7i1+k1z4ZkZ7x1NoMSginLfTcAfttQeNAUKJsi
JuAuU7MqD+ms1MW9V5dCWTZudQlan1cIp4K009/48j0NrQgdfujArVToQoWuCJOVOBLv8+KgNcf3
hTBF5QVrpqdDcNceLFrS+p4iFKd9DMfuVjvWNsgMF3sZmPv5afI+SYAiTEl84+wbqOggBPpW+C+n
kod6Sw1EfySv6ZcJqY+qBA/a3tDKUiSUsm6dn1TqWzbwiPsfaxguQAnRkQv0KD5aE+0fqNJfHJ/i
bCOSMLoZMk8IyWGJYxF59BptejyXoZVrEp9a0NVSIbUcMt8ETCfLoGsaY8rpRGR0PN0G421iLNfP
QMe33I3GgwqQo2GpCHL4jv2Cd2mIvQKIWideSfh5AxdTxZ6ldmMnRNrslwgrvMUYUvRUsyOUlxMv
oZg4SdJ3Jr2HPrBHhXlXQs0mAxbsHweobCpqdtPMp6WPv9SVXzv4ktup0pHaYGVvxWN1jISZYus+
t+OUKzem/lAlDs6y7MIKMtG9qNwI0OIjymOLUJEx3fIqWIg3tpk3CtkBkU+jkBHM3q5zp4aUbnS3
jVHo1OTrYq+uOwztilkp61PzEt1nVLKa9nWkx+r94L0R/BNfI1W0WZnzjuFLZ5KhFlJZz2hSirDz
KTJ8Zb9nR22xIhpWr06WIh1hm5SF5D7LcFUeVHFzoeUrn5MexUqPxdbevYDS5Yx1fZLebw+fMVMW
Vvk/YvP7RdnvBxZ01O36tBe+zSLNaN3XQH7EXaWiyNrsdQJuw+1/USjUXVVC8HUtq05uGoyziWsT
tapvkd4By0t2dXGriPBtsZYJfjaq1ZhxqoKPlOl58IogvMvOwENEMVIBvbR08L1UA/4mWHIS2jS4
MOrRZvzGYfPALJ1xUafkBlWgiH5OsuJl8a+cHfLCYG/rOrTD7u2Lxz5ZUmq7ByzCDsLqsVPfSi07
hqErrztauVcI3S3v5QEXfk+EpPaLVPcIJ7d2f/iMXrpkmK2evqqYZlak31DHniYSni7DsSwCwD2d
LQQh9S2leGJRm+ayUIWXnWaY2cV9iHnILoFUDT1mtsyDtY8dLRgmkGwjOhLPv63u4r1cJ9Lzecw1
vnPeFpGseIyTY3ylFJmRggb8vvK4ihjovreGetzmbaGEti9YMUOHDcdoMauUM4Lwy5wwpyMsIIcO
B2O3efTt6/4ZhJH+RGNvJCgTWEA/CTNqjB3+ff5075eTeXLmJURVTLfXE7egtxz+QxvYiXBq15Rf
ZLn5zwNCN5pTD53zvzYnByAKemSnkAzDfpY4A2V1wHZy+ZIe+6hjP6Xh9NgBnD4zDOzU1E9dg+V0
Zvn5DzhnYLz00PjvD8jQnZ9MaSUtWOjhnWNJWV7hKb/NIPCniflhhUbRPla6gdg9Ybr1XQJq6sUe
HYblllWnyWguE7vYfD6oDNloDZsAOSsvshfhu/GvoeuK4Jl7Q8LmoSzbFuCr9JWE9z+e9Wu/DbCT
pPz8XNEP2Bl9Voud/su41hRUuvaqlrNxcKlrtSc2eW56JSzzIy2F+/jLDdtlP2CQdrMSZvc7j5Oy
NRS8Hc9dfR4eqBtAh+56t2hcQ15RY+6XFo1CT249QJRDm7o4acdntxhhpdf9ONtLArb5XK/Eu9He
+oo18wxIMu+qUglcd2PWCSZkXtaveLatrtimtC+dcUzgI7R8LjhSDT+Py1wmN1TOSNHzc/lSghSE
sbcGEYTSxWnSQ7DJagqTOyC4efFnwCCO96VO5MNvO8PSu2p5gaoAE/284Sm7+SOp2bvjQgCfZrD8
EDQO0RkBxhQLPaeiKMTvMWUAK7uMrZyg98kFXuE0K++MHuWrGje/3D8IpyJQO92KgqaBWnf39buG
FA7aU58SA2mq22jjCymIEUOOB/R3Ji4TSDHngFLTvnTRmnT1v4yvOcQY5SvBnVJjzq0SZpJfXjQj
RwbN6hkQiEGcYfBBhVcXwuaTg48LYJYZajM1pA7S8Z9QkRlML8RrgxWDZWMkp0Hd/o86LQ8WpwjM
uWUbrY+h47hWILHHm5P/VstZRUL+mpaQTK7qYATIpjuDmYQ81YHxNNCy9VKyGzIicsMhJVedwSC6
JYOci0dTLT7k+vStJ3GqqZ8Y1o7hw4T9zgSioemABPDN6csDniGT2MhqCA5KILVpQdcXLyXJpMZE
6qyetnzFTzSDD8TuN/yXhXiqKTJ68uxZzzGtaijQsTLycAcl2Rensi9lzuLxOpXonTZiOV8NGN2r
3AltJtRlNE8js1Gzf9ICvJJC1BamcwTHuX2gXU9p34orElkjNAencZb3YKfXSZcmOCSegzX6VcHG
8o4DmdaTf120kFp/CwC1L2IOB1cDCjLKAwVodmfz6CMJhxt3K87WSC48cNpwyeahNt47PYgjsJ16
2tzszW/MjuONG/kxifOz1wyW2YbAB3vQrD2f+8E262Ge+ILbFlZYUYKG7TPbyTTKYg5r9quj2FJD
asEXEKqjT3ihPnTqHhDqUv1aHzOYoJdeFZ1UgaEsK74LCcLpdJZcAnISughXKjEXcURcpv2PIbDI
TE8qNiuRGFZuwNWuJw3yptYjSAofA+LfL5GDIG32bHwBoBeKCAKAxPj0gN+8HR4yYl05MpodPf6+
C7pveYmKzuVExiBvPzMx05xCPQGS9GGORx3q64+2KVKtkyZNM2u0yeX3LtZi53TXfAWmmxWiHjj/
k5eDrD1nD2dlONdS5Dd3HjU1Iy+rG+xe1lsZChW+QQKe5vI93v7ADaABNdEEr9vNkShYkEiaRW8o
9rpllZUMuPYTcTI7tbQ0ane3FgKl1mV/5eH5PA559penhCA2dhkF5bqYEsOkEBdiWIlwoCJYK2/x
ZEvdJMMOTYRH/+gi1Z7nyhhKtgTizgpkHRnowcn/1H4CUXtMHos5hxaD+pSitk3NCtrRlrgywdmm
U12ZqFhwDN9oGNbWnWm7k2OalLyzSJXi1pPzf96wwhPi5RU3fYLpUM0baZ4IZ1wOgJkhys95d/td
wW1Jt3SQqF1m8/dQ0KxiN+bTuCvx9s3bf+ObFqOany/EV2xmXELhesJbuxMaBWhETGe+sqLHDZYR
ABltIJp302k7cSXltfZ0PuVkhBEpxmPcAnaf2tDIt+HtwkpVS8gDnspKM7qyyHvqbXeB98sKnxXx
T9zGeb3BRRT7YSyiZEKcl2spVOJCNTwkXjdG6Beuecf1tU880ZcMdw7rX2nSh3M2N1ZMKEYXh2KW
0DBpHbOWIiQoVJKi6hyd2UEcGbQI6lM8hiQyJX9zqUomDEAkKHSxgeWw3DwLVylQYG27I/cIPEzB
27Q0BivMV3EigE7KUmAwJzrTnhchNaRMxsuf3uctRBEXihjotyO9T7HS59Z3K5K0TwKlcFmMj2Cn
l5KD6wQlpdiIB6h9gOmcmWKGcGlQ0XQxK5FewFnMBQ1Sn+QwwXDXn/0csI3pBEIqOqwcdXQ+Gu4H
sJWg9+k9sPF1dsIcADIuGmiz+4OCprP2VrhhzIvRgrvWaOIwwRhpqsTNeMWW4K3W8/kMDpkXwID4
zD41lXaUh1cfTcWQ+fX+RKPLx8ZI32stjZ3l+sHGeysdxwywsUOZ9IcNcZPlL0G7SX6xFcgaUVbo
vbsoK9lYaXCLAl6S6RIm0JwIB7ZhC/yqkMstqQp+/3T52ktOZr0DKX2QwuIsiQ+Nian3gzyr51Fu
ImUD5NicivUkc/O/SU8DkCXnn1gcc6qWTLYjYbaIxKRDPIeHnXnuaCn1VBiNdcR/VRcm0kJE8Sfe
LEeX/eePnZ5F5ViV50HOdEkbCbAR5GTuSlnn+roZqniVqD8MLFqCLeWbIGSfThkXXlBS6VQsWoi4
Bhf8LBd0Y2JZUh83AcNYSUI+h6LE7lddl5vILwRZTDRORGqB//qON4DG88TJ1w/Vr+fb06fir0oq
8WEXeruXwC0KUy9Mu5rVEiolFlyLGs18vOJkIiQZCyvXPuvsc5Y2826OwIJOgwthbqJ+pO19+zo/
z7Y99bU0IvojQZ7yViscCACOfk6+mrhF0F9dLcpGMK27yju5dGCEvbnSZiR563WwUmuO18E3MzWN
9RgV8adkwQnpkzKaVXUWWuKN0nlwxMLLqPKq2Tn+tnwA/T7t1/mD2wofJj3isQAiCs53Rh3pLbc1
T57VNVWe8vXR4jSgTs27248sKi+LMhTsVP4FEBQ3TWaY/2EnpOD8i++2fqXa6fnyXzUw7OiTwV7O
7e4Z1G9t47z/UdNXoGYEeXd9omVzsznNUIolxfbz5ev9sqwMYQiBF0hENllVwCYJRD3Z65quf7jp
euPKrZNO9FUWvRzCeb1nUOc0tSTRp2Nz1AnkRIaqB0Rv4X0DhLr2M4TuRpbVSHAVTr8eChEfh4gi
arsM7Y7abeG7jE4NxfiLSz0MQCuI+up+q8YbBL/rpzoArQI/7kUiJoevE8IPfwwLgLoGtrTkIrIZ
8rnPivEYtsG6MUQvkIpicy2d3FqiLwr9yh4iVN3DgxOwrJk26nOeqUjOyvET5iUIK0+c8VqzaIas
vxY4jFrwSTGDKroq4PNUDk7ZorV/T9tc05PgmUOmMVz78dHe1M3kYxUAi5Io4qNiPDYhQ7IcRk4H
7F31dddQyPZVslm6lkaeZDHK9dwLYKXMAoAG9qNAkA9z9Un9NFquniRZrq2Dqif+2PJgxpKUpqTM
9tckj9Cyo3UJCHM5BvlcHhZOZ2+p983juCQdu7nRUtdrG5mtPM2LUTsnjgOtDUcA/aaEhjCEhrFq
AU13rVk7ectdkN5goNAehIG59f/999z9CUUQhqUlHVCNdgAM1mCwhdORJQl/SuNsN875lTU5wPrq
JskigAT844KcDbiIEOoal8p0k6rUP99Hbraw/x37hcMVTWzZw+a1Wvn6B5oj95vFHQl2Cskv1KVZ
hZvLA0C34iVr0cjkG4FX7QhjkdtGfKU6yHXc5lgPCGassYBZP/JFtNw0T8o6SP+z1XFakUDWvnFf
6SfW1xgd00Ldee/kWSs/O45c0AOZ7eLYjMBjoCHoUnCm+7PKzwcoDHQiL4xR/hk8AXAXDwtKysST
99uqIVtxT3gwk7yN9VAxGrHinNeNdsveMmZwLJ7vF0lyWme/CdJ0zj5QIA2+uBImmCUPnc2Bs3Ld
S0SAGdbg/5W4NrhApPLq7/HqtCvdNJwN2TiHNhjWbxDnQJy//dE/1kpCVsuIx3EnnZeaajZYEide
Xadu6fDU7SJJv+IyxpTJYT/hqg3LQBJcn3+QdfoccFGmv7iO9Xggq/MIPJlg8vC7KsqesRMdhgyo
OrsSRi1ge/RaEhjxcLiknbpOZh+vSgKStGDUGbA76e07qHXzgRnX9A6SAuzz9qZPWcaGJ9pTyRG0
LVKN2EgmO0PVJx6C5oO1ngG3DJA/REeG/9Ml/6aQhUHM869EheQV877PIrSumtt9Z0CidFvnJSrQ
j0/23LBPgnPL2KA3kotLDWyrWpdTbmO9Auz0SyBQ7wu96yLbcZBVPyl2LK/GUxoMbRes9QC11Awj
0IWqCRiINyMdcg9ab2cZK57I0dQd5x+3YdquIz3H4Vg7276KIJjwTxRYWk3G1JqWd8YmMt7dAqE1
d8toQwbflhz7YE/MXDCWsB7yJ5q1x0uHAG0A2dKHdkJStTAX/LEgDQP294vlBMfuyfhcm/0Cktad
o4etxNkR2DWPnTJaH7F35jfHlglO7EYvyF397m6pYvYz8Bb3lsN0bWeXkGZEVjG7VN7qfUrU2iLW
i4TagM0cFt1fB6dnpbu/MnsThNS6aUC1k/eDeg1VGldTIygA/8JyalBVTVRyWT54GjdX5J64Wn17
CvWBtl1MVB3piNwfnYC0j26qgfDtIQKxA7e62iaHI36caA+RAmgti187XDzd0AXleF3VHoHtCI2i
01f/nHkbomOw5UtUnq7jw7vLk3192pB6UqmmqhGqykcmQ7EcAFb/6v7T6JeRUEQSPzeXmgEtFxWF
5URrb15pQqoLMAR5zEMoxmxhKbcQsnUD3qYOK7Y3+b+Wzjta7Y7eC+ckxR2YbNO0DZpzlJYKbr6n
MGM+ycV15V9vT24Eg73H5gTaMYD5ziF4BRHnQSIckKMSlX/X7cNhbDCPBHOsxUTtI7CvOFapLSbI
FgiWkcnhMtUv3a0q7eDrSx63Hs+p2Y971kMNMBWi7zakH5AH+376fI+AQ0pE/hzxOWnsisDBlxbo
hZR4WRjnCqAO+suQvebKXYpWaXOgjNectr3hp/rC87J9Gb4xgI6A+tPBt21qAzqPdEZYz4JAYpa0
33zBekwrFgvFUrB3NDmjTXmIvpsypEryfSGm2IndOF39h/6c2yfljilLLXuT3NDNY5mlZGpaXD6E
D2NxmL9yUZhnLIwTejAa28jsr4994MKrIUGEUrG/WbalecqYiaukudvPko27l/+RgyoRRO2vIe7O
T7ZSoj5KVWa5MYJIWJ06SNG7kkb1BWVNLThLZNjQU581Y4MU8dfSeWc04syeANbArCtRNkJF40aW
U5FHnEj14S5xFnqYOZ5wtY0UOL6DHQT6+LEPcnyWE7uRJ6zIreVi5aBgmwRtDHiw9eJF9x/RNC6X
CBr4NYV8lzrkPwVP+jgQ/2jQp1Eqsh3Lt2K00bL+YBWCIWY4+pT3l5PKjOFdizJM3z6/iTQya5E9
4IAJxn4KmR7/x5kmHx3ER3dopYtcMydAvrsGvG0NrS0TzHg9XSUsqy2m88PuXpyz6Wi1gVG6mdcg
kH3NV5YEGtB+m07uaitfua3fnn7w6nfZ9n9/du00LS5M6HIsoq9H63fJaaHTNFuui59pcS1tA51t
i1r9w2afwerDCBUlDAZ6H4YB1fhHwbHtIXQ8Du6zKHAGRrRKK3dttqWqap+aUDxQTOP3lh4+c9q0
imM+Jz99Ck1goCC7EqGuYG/EBD4bq1o0c/u3PM6WhYbIbdB0zmecpre+3yr3Uv3de/0lMP2OxYJp
aEzlh63rE/fzOpEMEYxPlje1Y/GW0SotiOZ9VKyeISB1nhGInM0SM8gIuAM7LHjuJEhMeObaoRIh
T5TfV5Qzaq0S5WqPJbtYM2okenMT/UWmaSY5gkFp+Ymv+6KTIaiDFjjG6HveF0EEC+b2S2HrFLq/
3gy+kWBqJQsZf8oLLi2Y/B6hbszl5NDY7X4a1lKt1NQeDefBZXu+PBDoLz4SjEHMSS6XWCbkr3T+
gk8+22pLhjBUP1iMriU2Rb0+9j0Xvfq7PraVhCOE/AkAH3DDD/hTfYSUks1OkztoiMlSqQAJLcbm
Br0YRrYI98quJjGvyb5FYmLQ7LifZxGvD6/1HXo2+2VXSJpRmFvzGCAp+7izdngmxArgqIQy9Knx
eBzX71PkhvlC2ZP9jL95uXMXzpK6EJNalm9tTHTd3hMkNQcXgFkZQvwNAguHn15W9UeFRIHXowzO
7Pb6wiBoB6NIk5+ROzIWUfWQWh2nMULDW3OO2jWsJvdbZ7/qrqttlSGrCnTcl5Xq6b0bea/+pwJt
P63QaKbOBWrph7nAQHdkQP/DDomcH1kgn/OjghS7Ux4acSo1Wnna/ztrPZ+UGsIiZeclfjaJy4Xa
FMu43B4pgJm65GqpyJaDfbjzGMOMvj0yQsIm3R6TcREV2wo72G4ZhZr3N/hS4LvMJHsWpeavJ+Zt
qLYkgz1TqU2X7Tb864wpc6/ZWe/evZY3lZDvidStbrMpsMVhLDGNwgYg7ugUIK6NfUtkqbSPgRNS
RYWQjisJKI+Q7t8zljqmCwgZzB2tQxOeqxwAaX9Lt+WPKNKcmiFetajho3RnLj7hiLN0Nx8FlBh3
u8Hydbfy+ggRRDyV/ROOU7r54Z8qwBSePb8Dje0dd4rcSloa3V/s89/8t0DGvBtDhLWifE3oQ933
RpQQuhsavo+kteLw09moWGivtsie1zg+TG6rsm6JOlVNkFSXskXhJkHl4zx9N6g5olXqTCROH6w6
E6OGOSnjI/B3OXMJwkYreBjfU/9+eKRQf+0LoVe/OTbD8KsmxYYSqhLzQ0+FDp9wRe2lIVSuG6oT
Zvu60EB1txqae4owBTBgXhQSZC14vxAWHi6K0Lrbx+DTS7JAL6bS0Opuk99KODp2nrq6fDMRE0DF
6I0dob2N+Ozr1vstpag/4ARqxePQOIPd++k8n4JgJypOXIHcxrSnPuH7oOjTBblVsdIKZEFhdm07
bGwU/Quwsbp6Y1MrUbc1U9JMP7gxt14uWqVrpssJ8VQc68AC4FJZQHr2fXqR8DMXKHCYtYvrrLNe
pOwl+Qu2UFe7nzV7EwlfffcQl5eRMW9crBIhHwZar5VQWRquBUjXNGzaBd3fPoNt1cLdieSoqJjI
HDlIX5bDgoDTX4ccyq0jHX8tww7lokY0PcaXf7NRCiirLSl3Jl6byaMT8KMXc70wn8tICr2B7/zZ
LLPAfOKm0fv+CT9F4F8JLrVow2KENl6Epvy9zWzp4LSge/pYZidIfrddq5uTQaJv2wRmwaF858uY
B7jv68Iem8YZmMc+lvkzOHnidRzrX92hZfPxeYA2UdKDxBSw0OToWHskcImPRFuyBYLDv+bqXTfa
2m+EgJbg+cXi98SDI6xyS0NxoPH6LA/tjt1sX449ISEcs3d1HUsPtI1oxhWe9BOfyiGyNUjnPfxD
EGqALbqKGoArjDU5NihZbSy/IhNRbuDoOrtzpiTYEBupkaJ00kiLLg4+WjJ7utQUfWJAUHQiZuwz
ChZBfcTB8hK+2j2ttXkvAaGjYy9ofm2QxOaMaB9SA0ubqVRzGUgvEVJT2mVQXvhoBt7vEP9gz1V+
xWxbnGZbakvg5pheDfziailz2Ugf1e2Y+Gn3/ZNCWzDKFaQDuOn2GRP4zBd5NJAGGXpQ+oxWMkjZ
2s3Qhf4VNiFAxH4qMK0rPdni3A6Dm6zoCYuJZtjTTvCt2QlBur68lD2v/bnAsxxKZ3NkgKTie9V9
ulMLxQZOzblkpZ7y18QCcRB+v133sRe46GFnzVE1TFWFNwPTJ9nLGN94cSskqf2/A397nksvgeax
IVGA+BwzxFv0VEGxTChza744FRJqUFxpbRfplD/vWNQwVg8ypvT/0+4MkfXXVBT1Ax/tejGwQ/mX
nWWt9bGq0Fj6HJ7NqniYEM2Q3kesSEr6ORCy1jbCGQmBEuJaQvSCLiHz/FzMq37e+AucoRgLpLEx
JL/JZAohosDCFnysBNJvkXLOL3eVbiu6HsgNjrzWoYjDL3g4ukryrbWnMs0l5LMejU9pq1HXAO3h
5xAnfrKP1AeWaMzW3K8QrxAvbnJiuiPZGtJxVbnlDUtE09LeTqSIVZp2ICBDwGu6V5C5+tx4myvc
3gVngu8wHp22VybNFj7WEs18UVjzwrKSb7KwaUjUAt4eLokBvfexOrue99wzD/3QCRuc85efRPwD
ql+vcAeQ+DiidlbTUCCFkpqSXLHqn9415gmQZ5d/QDiDe7amEJz2R7eqQQ7WmfsGbc0vRIB43vsN
lQwEEHuDLyETOZCy1l6+h+P902geTI/OYGczM1ts8nOkP8GTJddRPBCuxYF2cCBpHBOmuud8hbeT
K6zGBgYkcsAfgdFTGcRhrzntsRhpVLtSGVkmV1qimwwBf0T7zeKWF1fiplDrNB3PMkKzqvUWU/1v
27oc1JS6WYNNHmSWbq73/+lUTjgzlU2uqKHQSzeWMKB0B9xW6fxT/Q/AHv6X0IZ4ZLh4BQUdbHFv
jJIOdzK9aVjDQXb7wRRFnF7kDHsv1hxXVD4j4ImKzGylofAGNe8evEZu0E0Nx2hIgFWHVEEDa/m2
AiFy98fIAQNu9uTJCRiJQ0St/LMmdFXNEwvUQiAFG+xece3WqWaaSU8q9WrCedpuCAsTs3ZIzOLq
UraB6QBsaLGa9h0z6MCVPyrg5aUSNm87xFJQJyZdsSMhEDgC1XtbC7xHKUrcxdzPoUVjdWupAVi6
umfwyaF28A6am4PWxpW2ATeMGn2uapeikOOZZqsddTSvtNAGOD07vE5OQn6CzHXcbC0DthfxDCU2
wFzH+M9b7LoU325jDbIsxOwEh3E5b2Pyi6gjk/GXON9oHaY6R0WDn3QJlErYFjwLGcox8WOQkpxm
ztJfRMI1MTl4wEFYDFMN0qgwXGuUE2LUFQbNHo1mQaCs5WSohmng+ku+J8G7vnjx2hnxiqzKQkn3
Vm+ElXdlt7+mTfS0wmQIHPwlDxFc+5s89ewRYKh44q1yfuka+cjtVUHMEDtvgUsJPUdIzTEf8Daz
iuxt/izLCVnWW2+oZodUoYAlMJ76KjTSU0RDav0oeZrL7AVXVbTAVCbLb0x+1TkaTjG5H1gbqbvU
XXhG2DJbTaiU6Vt78hgjGvr//8nwPCsBxmd5gHle28FXIShI5bSx0NHE/YKbjyYGs5K+xRNzqKWS
ZQfMSYRF1DjTlndvxidjb1cw5LdrRyAcNgp9U5kYWYsvNMm87SQI+6XjF+CD4ccq1pvqpl96ht3e
ds8JhYBOZOJc1KqVXwXFm0mP8X5iIr0MSaaEOLdmkhzabhi1nvKuDZrneQlcmxSSQVWk9tmZfFXf
54zpl4/kxVpdVY/i7uAn+Vp4ZdzTmN6R6z7hsm6HamwDmW6psBTASX9y5inrpKI9P+8f3+txJjlj
jxRB4wqAQq/XlaVk8kWpdRBE8oCIEfA2qdpq30ikVLnvMrUuJFZt0G2mEgKiROikdqjVP608ITOT
JNL72fMgVkIQwPXfZdJjy/rtOfnsj4AhCq0s38jpEFPmhbObOcnq7N8BzryHRLHW/SEC6nzzLb6S
68IfPBqGzL78jpRyNJJLaM+1EKOMxg2B9WBu93bkoLcDKXDARVWrpua1wEhOfToCgFQvdSrHMfXT
I6kxEQLACCWaucEfDzvgfVFIP0tKf5GgO8FVTF6EJ/x82k/Xq4/Jafa8W+76//WUfLR9sN5HFR0i
whZFlEc/WPbFXtEVymARbdKdjlpLogMnk3dnrNdE7HTCk0UldHKV2yqiIw/GzlVmE0jmIKQNfMXo
/0yRzDAhjOJiUjzZT0z7RPNtexf+UC2WCaFlwT6F1ydaic/RsRBFDB9gCobNS65dX/ZYx8HC3ri+
SnYkTpCd86L5GLdEmedQFdCo3xjbdEqLdc52e0ne9F4TAYfW2/rDTVLqK+mslLis9VWq2YN6jXCX
qQrlU8Tz5TfK+7u5rribM4YbYZZhuhK+Qo4dbSOmp/UbGyNO/DEVTlMvjEGSBntlLUR+U6Zr0/WZ
JTZYxwK7KV8uTSNDHuxoB8jZfvw2HKScXwFKW833RXk4Id9/ejLwG+bclNjWYy/Zh5PTJJJV23C/
TJN/oOECuSrXEVfYjikMPtV5uzDGmQhPR7LUDxnzVS1eQ33KzH+72u6qGzY6qOxVFVV8+hT7K2d5
cBnu2ioQCOcZHafh7mdNweYkpwvxJ3R4QU/tad/kqAjG21z18ulSqRY4IVeW14s/D4uFvmRk2w2H
KORcJThaRcgOMcuJxsEYfY0yIyMq/ESZgUslj0YjKLw3Fy9x7wjm2dVMflbq66QtrGoPH6UbNkz9
DaFayddu/s4m5soU0pnNk/PYtGbxE0dzF6VJ4z3yFQzcv0l0p0hSj0MLjHdNVVhUkZhTqu4WaLvK
tXDpqjezG7FJpEoZ00P4sOACc+7tWhwDwaKX+Fp3Z6eRntgPL8X1882716eJJXoD/gR241EQHv+Y
ICdc05/J1vwGpGCn1gu+6y149DljKZszQWMNhRoqlvPp34S/Qyd0jw0YRnocs6DrLRQ69NxpPdsl
sWmEnJbkij68AUH4nnofNrmrLkY1Dk33XBeRukm0v2sJyZa0yqMYKyf7CPNnGxbodLA/0RUrgLp+
3MFT2RtjBxsWmk802nBoJXNJGv/SAR1FR+Do5w7QGkrKJIq+u6CIBUOvWfbZCYLV1PcReWMd7Tj6
dXQ6hUqdLXGN/0MpMNNnwHlOZjDaBs3J09OyFd2GQW/e5ocmBMJb3GGhvAGx1RBZev1p9rZWC+wW
4/v6Ji7Tx6PqSG08rbVlHUaEW0TVAU3quWecVUuN0qe/s4VquI3rR/I4MsYisblI1J5hWBYGobeA
gH3S5kCrUT75c0VcImonbvxnsu1AhiRNsUnYttugZfZERHeNGq85kuDE4CNrQvTyHnlspBlEPyue
lnAoHdSm9FRy+Ws1a7a1H8I3O7vm2yNKI9nUm9flVHr1PvB21Z3xjbnU6ahumcU8KSindWm0yLEz
5o8qLzwmzZ1X0JHSRB8EuLj7VLsRYWXC+WI9qJ8DxPvkvm9SsWE770Obj3ZVJ5N0Jcy/cjmYgNCd
Dm+rEURQn0IITh+Iy+4Tl7aqFfOoOP7YHYLRpqYkfgkz484vwzdHZib6Vd6t3ij6Z/rcs5SJ/Goe
39EW3xh7cTMrr5hmbmXQXZgk+dm5OjyNDGBjw/fvf0TO4AdgMO3z2b81zK9m3L9J7ijBSRZvjD+j
fx2rFayXRrIcmW/2+HoH04j2HgCBoDf7I3IhtcQx77x3Pa5HX2HmHPtUI9quHmvjQCLJHpoJu+0M
uEUlhpVF+GnVw/85DCdZar8aiQzw8ZYIqgrt0JZkWbCOBvQxTEZsvobNxCJgHwF3RGCOlPvf9HHh
iXo/4dB0r3TG7pe/Y/A13UqA+H5OKQOrlwTlR0LamZqOzObLGfhIB9XQCtTkTgjSiSNxkGgrjdJj
jhhC98ixFUPSTAMqknd7L3L+eQmNgvguIW9eOtEbUXaX1v75IkqZnFrv0LgGTPhhTGVGT47e3gzT
GzddLPkXooyLzgxvY9xSYBilUEunr85WaIXosBtjFzu5/66+Sdpv/FcTQThSb31uOGWfrIrFsgk5
POYeY5oGWBGsYtKtR0xcyLoWLsz72t4XdLKdUPgwOaaLjxVplZrQvhFw+CjZ1asSaF5xGoABQLyb
mPlqbdzvxC0rUwVAaz40rn6x0DPDsGmA17PlpYisZVvv7UCX3jQe+ESGuwJi0Pkkm0FG3QqaTCmu
YMqm/ljvAZIH6LkyZ4KATOTkH/csCCPhVjTyimZFm7pCRILwyva6JDGwgwoqk2JQ8XaW9yIO+7qO
ZYMQIh+q65sfNVXTMEEX1PVWIz6SlEwHJYpsjTp6ONGdGIRp92O06RC6KpEOtVyetN3bAS+tttmg
FAmuMMt6BEun2YpVifwqS1Au4ZCXuFQiqW8OQYShf679dfjyhn9i1lxr/nLEkpkSblL16D94vD79
srLzNleWtDZLoynaKhS+sOjxN/rx01t2+vlHS2c/eTi7rTWqy4LB3/yXatgbPrgkwdPanngKOyLG
qkRde2yKbt8OiX93E0XgtyRsmDtIMErejrWV+2sMuUoCD0fXCgCcS2WBPhLxHch4qyBEnbUAyTCu
t/++ElMSOHb3KqCUzcOTyF2LhVjtgAxAl81oVlkPvDQJYcK73jrUqx70ZrfjIoax481vZzG/R2ga
dXfq6WbLHFl/LqvMWToYU1824QPomyFbt7rpr4rQhNrFGg9q+sFFbv0msyM+4nYqkHkhy2V+Dni9
IEmkC6q0CCT95cLySq7CKhy3Amo9jsV3M8ueyfl68zO+BsHnyeGtH3CLI7nQn6fW6W4xc4iQTN9Y
aGTdQ0To/xclPDpY6wuqpWvMhEBUA3xDsgvmhkQe1h4zeskG1FauIxdaP4PWEUj85qut/m+XVO63
bEekt88zU5lTAVV7vo81q9+O8tZwvNBmFrAHPMD5zX4br3lXcTWt8IqFAhHRAoe76mC5zLzl4+/i
AifBBCYMEwHFRA3jH4hObcXdJRv12LtmF0WGLO9gidjH2HcM2rhKFCbeVztz2hw/66Vzio141ljn
xOCLUJB3xUylYDv8GJXYR4HLlqy47EalKNNaqG8u74x5E+U/FJ+HOHDEwJSqhcBKn6B/ZGa9JMzM
iTi2J6zTr77XbnZoKMAv3FPpdIJlyeKWRkfvNo7hXveN40mxk4unihFzyM8/Kc/+tCp7iJO5CW1S
ef4Ik3AP7Ru7feIlSBMhAyOawd9XWDHxwvOmPOte3FlDIrB+7YuPYjhbYfV4Jc5kxfVjYcCGVvNe
qgqrSeU+eYlO+JYix8A3g0+xjTi0uV8hq784mhMvo2+181SMYhAgPdgBgpzadUH6DOCvIeCREAdt
OKuzAMT5JykxK+yJCJXEUDliDZ/pnhOmnGN+1tJBwGHLGlgk5K3lDg04cI3vy+6h7WDD9gmsESGY
iQTJZ99c6o3rpyfQyUiQyeUm05fXOTrNTew2SF6MoHuVLi99bjU7l01+7WsHp8phEH0lwfns4d18
gcVEe/84zJFq5nvDzd2ZmiFUakKcV40FbKuObFO/xahUUCEr0QwLy5m7eEDLZD/ewdZJVbYtOdaz
oT9TCNzGcgMzhC4U5idfo6GMXQdBPsjgZEF4ZRpOjGx8qH5d2sbn7/+4iu15Qvv6h2CMKR301ywy
xHj03ssE4kd39Fyz52XAbmBwCdEB9d3V9+6BXVWDqf8T8eLhA8BrlBZuyHNo7c3K7GgJIiU8+/h2
6Ft68Q3Pdl5bSAXnluGuq/fRG0jiAryAhr5QptqrO7VjnZKqBHu/tRyIy2kLOdBPykXX8cFkV3LN
r/u3m5t5uJcT0dt7+QQBtWmX35ld40rgTPF9VH8JoYuniMI2vyq3qaXNfyDtOhNwvGll8a9L01mX
vDnr8qpzJECZKKsXmHvj2GOhXCbhdiRsmPRaNvIKspqwQJzr+iTifmkBvJzOLwJqZzykZzdOPFph
Bqh1/Z30xSB4/xOa/sl5HMS/yEutcEWAVTvn6HulxW4wVeYZuUAE/1tUBmgsC8ThSL9K1jIqDkWc
g/pPG/rE6X3gPq/fdkUxmjtARlyhkElzR2yREyPjvQx0YT2EM8ia/i1rkHTqMdZXXDRCBVLRU8hq
cZG/EmUfBzqSdet7i1HB/P81Wdh7vZtSBexdFpm6AcrUiVBDm1Pa0fd6zH67AfiOTok8R1ApBVd7
dUtUoR/ejseAvwJePg889X0mwF6pN07adXiS8qCBKr5dKpvX+525c+NwgrJgA/Ll8yTU7EF6cvmU
O8pHYOjMtUdcVf+TF8lO9ZRN2u67/UTQTiniTBoaA86h8bqA0xVeOffTtwjdBJBcgy9NUSIIwYbe
DIASsDCTH6lV2kuQKKQY7pO67mEf9LX4md6I+/OybZDv560Zw8Q2rTAuPJHLwIh8ffl3RCriPHWY
HgkIlGPkSUkrn/+jLuboSoHzLOn24lXmFQm1BU1yXVyxsdJI0UMgsB3sfrprQ2yA+rhSqNfz/tNe
eKlWbdtxZs8cWY0kRg2o1DoDQN0/6rbIy3LAegQvKE/wjWTRUtAkKjuBRRGXTW62B6dcBDgUBzB2
CduvTV9QvrYKPO0qPC1zP5kKBhpN8vcSpz2ZOLH4RJwzUTD8RzBOZIkU40/frxDa/aPON22wRJR+
ftXWe2DyhZZm55zWtE9w78soY1HF9gS6nXNjVtwchHqFOvrcTHHgEPEojZ8zOBUrGhSuhRK5x3it
HEHsxQ1ByeT+BWzjjlAa27Brlp55uCsfLddaBULC+xYT+09BSYzmB31mGu5DhE9n+c32MmvnGrAH
PFQk3IYvwOYCi/ayRrMu5fmiuvfFGu5dUbgnKCQCalM9/uOeM6C2qtiRV/j50n6MO4Ni7gRSkHW0
WWB18d5WL6h/+oXq7RDEW+sFu+d/9hjTgX+pC4q1HePJvbmcd83xvxFWVkRfC66KhFG8KYoaKxrJ
xXxlryL2PMrBHsEvQ50p/33VylXbQwjufNOZ0bLUcjmimUJia9rlIgn9JPWscVIRrwbJ0m6roJ7/
16bW+naydj+U91mRp4yiImtlxAdBqzE68pT+FDN+/Kv13EKMwCKHc/3GQ3Xix2+Mv43+nqT3opwz
FaO94kzLwlIzLGRQChDlEzPrsTTLLe3gLSlFR4m52fFKYwn77INKUW4Ijd/bgBU5OXrg1iI1WvsU
I9xtOlo9IZmq9eIslJKJgGFTnIB7YYGauxpsJ2jUMJmeiF0qfDyPcaWdgxDv8N52gzwiD2lVxxkg
HJrH5Ec9TKlx5MpyEXKQfeKM27DMAPz9bC1MrYcKbtS/ab4BfxUFzXJEwgORQzljwwD6RufFqe4L
bGQyysimuPnIJXlIbLPAZblMYnl6QA1CnCDtwqLYOJEvf7w3DMvTOfbOAlOvQ39wy4yO+sZ6n8CF
uk1wZy6GEzRDHQAwGIzqRprUQriaUtAFtVXZsHb3m3sz/Yw/6Lx7a/ZCgFSO8/sjjQ9CeMIWLwDA
ryoYuWlloDxwqhgL27ZA5gqJY6Bidq66Xj9MHzy05YuPxZHZP4/NLYrCRLGIN4hZpbechWFxsT1B
wF4vl9HATDHwf6U5DcSg/9GFWD4uSdiysvKic5M5obgpX7ZYIjWmWWhFSQ8qP7R3WTt/w382FE/9
6f28uk278DZw63eiPzDiKvMUb550vOkNCFhKIebmwbqAnVu9uQdptnAWem8hc99/X7mXR1wev7Xc
DUcqKmtFK31KdogHSsy3UZrJ2CugANi9gTyqRBPFRGR9RFhw/c9QS+T81Ewr/dIgIjJ9RCavi+q/
+pOxZ02rESH6e0flyAQMSBvdXlVzZ4qg1+3jxDedmjiArbtePN0p3I3A+YwhyyVB6V0VdF5rwvPk
Z4fnHLNQdjxfSX5PsnEocRiHRwptdU+7MBDqqHbK8evl05TAcryCFX//yLH7SORAxSm87pkje9+h
fiW1FQJ0iddCk1Tk7UX8ebhDCw4K1AqzjQntJgH+vsBNUaWX7qVqSeFuZRM8LeYX0ByCfcUmZSkg
FBp7lh5d7lf9g89hML3UrYxa/m/JzTb7wV1gg8K06LlNALtZkrM0SwYIruu7X7aEsCapFu3UiczT
OiWQQ8rcqGvuwlRSkNXJQCg4w5GLnlw0jQqySn15oKyka337X/l/XNjO41fpXvfB9fXbT2hQiYYD
Kxyyr6uCZ7jiNrQ1zKBRKi1JXDk30ZMcwGx5iKEhyjyNKKMIMaHjREkTx625PvtipVh6DQsvz+qm
6K9s7FkI3DZjxSrgbWWsdw5YSAXb+KvII2DhYJo9BJw56E/d8J9pYG4lVAk++PNzeLhaQXMUSH7E
phQGxuODhRMABJYSl0rbbxkxIgNrqTTUgxbyTzrEfavWUnSNvak7rXLz7i0c30XToQdvgMg4Sx0z
PvLVoME4egRBOeOKCVUm8w/QM9uBENBmxykoyHWU/79HtTMtq3badY1qaa2rqjtd7muDYm4hIwG6
kZ0u/OfeW44xyIH0YOsUOdL343SfFXA4pKhFVZKH/rO9Bultsu+GWmR009cxgJVNxvEMOlBXyHtH
6LglpUSgNisv5AHL5KTva4+oaClISCST7A4eHro3Xqcrbgo6tY8OTL9bGz7PyniNM8RSHFv+Qdgp
ZrKSHETNUaeClq8ingViGOGJQTIGlWmwT2v3Nx2ub4v/1agobFQuRgLWYQDOoE47kODmQsxoAgdg
CF3WZosPC93IPlgHaBSaCeD68vi6E3u7+KPlgE7FUYA3s5n81t/sTS0GJNyLbY3SNbnn1TZLr1cB
b7OGg/Ci4i6KB9C+ZupsBFZyEj/VN6Zi857amaswDjujTNFWM8HJA5sW7BCbMOl3OniQ0v9H1z4p
uNf5eXHCnadouTqwwIBP55u5IW8r4pWVcmTtBlRnMaFMtB9V/fu6PtNXzP+vk0cg92hYWd4/Y19y
qDgq6Njd22nW8/bak9pHRN6tzGwXxZ6e2kXIU/1L4CmJFH69nt/iuYLF7quC6SQR7Lo3V8fKTs3y
NunpaPmySRoZkioYyyAhHMAo7hctl9onMKPm0DKfNVWJcYy4OS1rhmMh38vE/u0h4562A75n1Ok/
AGtGADR1lCj0G2eZbHyoNckonwYsR9g0t8N9uUKE8XquzFp6zYSgalfYf9AWGGxqg3Rj9WsOeRyf
QaSfEtbTBbFQU940MER/3gwSfzn9vRmggQokuVft8Lqu/z1jSecIT09CjEM7Xe4C92SnRr3oKZWU
Zr9ElkqY5m4L7YtGGGTvQAvesGe/rLETJ+CyBvV44tQNp0inrRSiKnSwR+2l9krDwjrmFF4YyyE7
lPZhv98WR/GBnAkwS7io5dNt4zv7hLgX/2r++jjNqRaHfp5auPysOdOBjgwsx0JEsQDYggfuhf0j
+c2utq+ITqIiQC8koI1yDTb91ktlDeQ6v8nxUbj18F1JWrSl05IrW513Xamf57+QzFtIs9h5LF6p
hweglysSUeJejplsTaQRbDA3PS8ikjRBLD8wJsGuGwSJ9EJ3qvJ5xc9Z+U+nVsG2grrdCIQW5o4c
0+S+qwxA0MRwzJCnHOxtZOQ3qd4OQJPHV3PKBqbCe/8hb1iA82p9+xTUc4ufDIWQHP6G0mHMiQ2+
O9fM+/0qbHePsdBIwQ2g8QeHK/3G6+ZkCatrdhZ/VISGyJwDuH29oRn/YFq9mwa9VsxreUEk3O59
r/7rWbn6WbzClu8y4kf002dlKCkTVaOvXWLopdyTePZD8aRkkqo6dcRSFt5832LyDtI5mddF8ZsH
ir/k2MzRiUUYi5FVYM3oKVkPlyy7DzNF+xYOElxHGiCA+lN8EMirM8d/V/2/pS7v2bPcRJyy5NUR
4uvFIB2qFJWx5ysSWMPREha8o5OpmkbUo2wp1Tkr2vKhYWjEtxGJZ2ACmpZrfYm9lWpYX3obbZWm
5Vi2JX+a1D0sAiX6Qu0Sc6EIBhn1SI8+QAGzzv4r8p6UWjX6OKu6ZdkWVCum0qdrkiT6hknHUyln
exjeNAYNDaOAKu3qHsR1YKv2QnKXKXUd9OYFdm0JJW/GHOGONj/ROBB66MLei+hGsMZg2BdJH1H1
fM3/kUnTJA1692munFxYUpGs5T5JMiIasGPHkSJdnH3GQBPNbA4QepZYozezByJ3uQrPPjQu/luA
ZsPmqDflqrCVgJDJvRAHbdZlglr9ENIYBfHSYEjt0i8cnWwXZUCjnn0UcOZFu3h82jG3us86gAq0
2tn3HdLXh3JoJa0FpKWtUeGOa/hlNz4iGlnSC/op6r1HRKwvCNrqffnnluE3dhIbrqG2T0A8ysTY
0QPEuUKMMDYJHC+fGg1LILK8K1pwY+6u494oMX7QE8bKJefHdAOzNZlUXt25xT0Cc9FUa6bpgbc3
CB+mx7lgpKsFgNEmJXrJb5ImZpTaT8PatKzYgVbXKdMMYd8yxaI225OzjIn81wg6qm1NDgRq/1TQ
acLPHUtzhl6e9Z4VXoN7k+ljRi4jcVQjwc18w9yX9IsfeDC1yjnrH2rtlE1yAhj6nk3FE9xF5IUd
IDtQpJfjVKQ2FB4iWLnPmF+Qh0lRnU3qX+dkDpbdqzDG0PwffX065soIMGFc3mUU5wC6YIXiJ56R
8JHYUW3d8Duoet18RDIEdsf8l1zij4mwPv7/qOzqgtzPk3yv/5q0h5kA3Hc4uG1SjHxkUHyS9INW
vr/e+DxLbcNaOmgIDMQFieStBeuTZZ9KCjPxdYaQTvX9RDTN3BAxfFao6VIjfyAf522KfbrvvYST
Z/b3n03yWCMMS1txKzR8RhwByrFb0H1ej0eETOeClRShofZEb7017OprHTEv3JbVZ6oDGx8GmO7q
7cvmub3/ZBC1pcguCj9udJmtM8fWFc88Ux9a+SYUrl2GshjZ0dEY96JsKfLgyk9XOweyF63ps6lf
TCH1iDFVyPUzy4+h+4oR5WitDXHwl2aqznKOabjgvVA3NeCuYQji1Ky0TQCRlvF8dQHZopsm/lU9
gayRZ8Qh4g5/gLJS07D3mxtZFGEB57j4mxobqQQ3KeLkbzdHU7gfJ/S9J1IJRbPkJUwTJ6Y4sL2P
sC7URcFSHMYlsCGwbEn4eeCPuXAoZGmTVDA3A/omagmMV47//mqRBRtszZlCmW90tRZ1gTQB/qrt
JTeKmaj0HovBCL/tfdyxka9uBAWVt4Mcfmx8+J4PumYvb9Ss5grTfhhP38EMjutNlES4QZK/tZGO
ssdfz5tQNUWH0DzesgzjDxT3kTbmMfddwSX8XMWWFggEzNAnRRVsm7bMmhl6eqyMbrMsrZQmRp+q
/nyUopUilbFvkSWQ1MEMIhmSaPfQalB3MEwFNRmOnMGk0f/Cprq6bJZue3bPhY4HFMr9EgnmbhaH
f2COKXqihWwXuWFqVmTL1VTaM9kBF7RM+ZO03ukLV7r0hkV7t9JLWdXHnwDWTD+bdUVxyN5D+wfH
gnw21OoRhcORTd6+OrLexBmtb4PgTJ/Z59oAoPv2+2wzX3oQNmDiFV+iGrmngycR1F4J4IjYGI6n
3wceY6IR9Fb13UMCYpQX+zUvwu5TZRp4lXE9/R8Okmqez6dXvVCeiQd8uESIZxnh7Gue0oik2JbS
/4qOV69Co3A9sKU0z7caZQEW37NrxxA8wqIGS8aqrP1TQeKocUGO761UCRwKJ7F2JhvHBgGV784N
nGfz+x2e1h1eSJYEXhwBXqdyAOWUYH7jJkmZgl+SDn19Lt1/x1gLf43Io7t746y/Ycloxgs7VG47
kFfnvEE2sIX/TQR/tiNN4FgZrVy8gBpKX2Dbmf1KKyCwifzJCL+DTalxzHgbghXYnKglW1trvy2x
Da1RJAHlK2ZYY+sOnYjNnxNeyCgIRGtPILWJSrIrQup5X9SqQotUzyJMTpabO6Vf/p9ouMthhnlF
uZ+wlAWmqjwJyYziPM1BdHgEhfr1jzfIaj9ofSmrcG26kpkgBOHOzvqVKklruDlwwPpzk/H9PpdS
fVCDcb2gAi9TcK84NMI8TFobu0PfwyBB4yLNMFe1/+lyqEoovWbcwMlXydfMBJj8m3k4CNZTvhCv
e5vm4qLcbvvebLRGhPO3s1jUq10RrjDaml2S9Kzb4tDT/gTXqnAvlaCzhz58Mqy5h0bhAhcAiNZA
np1suq9HdJvb8HTv4vO6+4OanWSpr+F0BAhyJ3xWV9zJLXHrDB3UAnyHmcAks/ISOp6Yivwo1ceD
VuNZwKVLPwDimRK5NstbsexQPa7DWUrJTDJ15WsomR++UtD34MOWzLEdbGq6OPI9pbc0kGifYIiA
TupcBPFbF21o/c3RxB67ZeOmWRJHecWxkoRXUnM129i/eeaEbIQXlygMqBT9gLGFo6AUP0j7aciZ
ohM+sA3Sy+7PrDrXNftwpEKDVtzwbLbPX8MNEOEwdKkXZkdRMf+UrOxbDwzvTlZkThjG1a7T5hkO
r2reX/ECJ3i+gS9emmaIIMG8HgplsRoiDuFnUH7BOV6Wq4RQnGvABLfDa8ODLp+w3yrsvvYsEj6i
SovG0fy9P4VVvaR3sPdKmyxGaoy9NCd/W+thA19zGkdcBqwsrV1piwVYAzD0HO1lk/FChu5UJSe8
1DRTk/yzF4UBMh6Bj+b9BVekgf0H0U5v3367+vsSdsZM5GCZSuIbH9ZomEe9TVO7bJozEB14QGXg
p17ikrTpWXiU8dtW7TMKEFucjaysl2wpP2Y2ubkOHbNETXFHVTb0u+L8F/6FdzY7qhswVH8g7SKJ
ZlxIkcPvXiQgvtqrqLzhlaeqMqqr6ipgs+brhG0ETcl+WPy5ww9C7B0JZKF6Lc4QcmD2DM/gveNl
enwOjDJpEDEub2Mx6YLgKryEIBKU+Myr1AEf8ZzdloGG2NdFszaAKThdCxz4r3HA99Pg11esF/lD
mqE6wC6OPTdNnLWnqNktlnKeXnBdI0LgsoGL+BEClTGVesvMJaB7pfMsqmA0ky/uWeD1qxEKRvwj
2BQe+3dBn9U9UjvKhPzRKHZcNQBOa6DkuwgQLVbIypzu/IU7QpBRl6wYq2/g7MvE4/kb8+3v4jBM
Yh4YUIebZZQPpDjy+5QhsMePPXTxPCKivwKiJkf2d+mu9vWnXNQ0q+UIy5IaVUrD9/W/sPUJtMFI
JVNFWJhLmY9/ygH0aZzeWnYhHZs63Az0bbItQZL8pVB7gr08796lFFlxxObCQHfjoPwGiIWMSYnS
jU2TrQIblcXyudBbwIrz/l4lqHBagZVtccCbYc1XwzgWlUrHEhffgxc370L1tm/PoOgGy3WSJZuD
IZuP/nhkSiRwEyvSm72VdXB3kkzKvcxXUxdh0qPqe5TdjRDAMa/aOs10/ycDDkBcIz8YlNQgzzJa
EDTe/HoiEgfK+1+aSltC6Q/+DB87j4fczDxWWkouAkjK8oeCyppX7aM1Kve6kuhz+6iXsPVVU3Zp
XzN7rECy9VvPGa8oNXMWhnv0xGflPQi2H757IidTqjS7O27dT3IexvrOm0N9yTGWdnyC4o7x6jgZ
00QYwoUhCTm4n5bhMzRYgqsRUlhsnz4+gOMM2EsmMpUoaUfwRVq5kg5aMGefs6Ckd77lgAdEssx9
qEFGPavnpqXgSfa0whZP7MsSpHECjL+eAI4R1iH1MUMOYeAjJqTAhuLDBEXCqw5L/e2lO3xD1X+U
KfX3BjPSh1B0ABwQLPeWetL4exi6DMYjDgxk13mzCOPuA0OVWEkjHudgNL3k8/7FBqF9YLNL3VPS
wPV5P5d3IrRBY5fwHv2Yp72RyPtaCoeeBft2ro4FHmG5bl3SFCw9Fv8KjmefEmesapQhyY67jEf5
gq/EM7YUbPyb7HwjbN9CGZYHrOvPiYBGFsSKkdK1TU5SkBCYB65q+62vGKrAHEUkdDfypsmhtTbp
ZvaQ+tzyKR/zsBh+K0b98NJCfCbdp/mEEgT9PIxMT6YTDsLomh1N/eI2avt/0saAJb41YmTDCayM
alvoYUEW4DOlIS3v7Qc4XJhnTeG+gFbpBx9VFAnkQRt5ydbeq5aIGrIA7btvU+84SlUNEVE2Os7I
KccCNiZ7wbnlWvGiMYxJZsoym1WlbJjBqw5P181RBIeKF5LkszpALnK95QPgGwv1rpw/njXlE7QC
lnxcwHOuAip9yJ4OVq7gsUO32erqMxQd9A4tBUOsNsyUrPz9GFOurHSuXQMzyX4WVCayhkHYcLyp
KwYQMAKFB7/PclG3TiLNmsoyrV0uyqJOzSNvg/3xUNcXzF7FpT7QxdTERGMghFru/nTatSDZMwae
PY6PLHDBcOXP30r9XC+PNnnmfRz1n4wZOOPtLoc6+fciMRA194PJFxjfjMCrSu2SpOkPc39mvi/9
4eyR/3OoMSUxbMJOfjSegY74eo9/UAjFbyGCBh/vIkM66YSgXfpVQvSmtsWfCAdRWoxKbhNnsZSd
aPWEvrVf9vxAoYDcbgy6l54h4fYB3efxser3A2I6a5rj7AhzA+NQ+Pi7ugWwLaZKBnrzaieuQyja
XFaipt7HPbdzjm5tDktzhYiesTloTanjovwNVZRLbn2SICe2wwOt9FqnuwJYt/iZ00TaZ5vlXvX/
bJpX5OzsR1uLPwhy8Ee+CYtjROboKG8gMP02ECoh4yUDbX+LmXF66gLV7e7X2doU0+5VeEcKeshW
23Bl0FjBsdKNqSdi08k0dbZ+lNKFR5A+NILmh5sLoFzkLWJWuPR4/gA7ScgdbBHI5SecKPxSeA3M
hR3d+IGLDO5bun2Iyv9ISdjTbdOEuQYorAeSbUU59XOyqgUuHzB6PQ0Dl+sMzvJc5VJunu8Xz6Lr
y10gAnmyGTGGmsyCb8y9ahWPrRxXwh6DNRDlpLzaTI0EDx8019eqb/n2u5IFwpMHu0pIvi7a0IwJ
hsW0D8JdtBi97ucljQcLDke19ciJoV3rTeRSH2QsEx115+7T+DwbG9QEg31N0514eStenvOqoVoO
7a8mBPFPcY1vSvIpFQerJ/E+S2baK+XcszV3txPZgaH5H/tSP1jt6RzqA5kCSWQIjSSIWn6P5WEz
255l/93dJflrTgd5ELwqJHzzR6Z0mZZlo7UHd0tgjWhUzxY2UwV/iJ4BPhtujRhYs65y9OhULWHC
ityyh5YFqWnqO3jP+zM6Yf1bWX78gPPdsASubyY22AJyMQZ3z+6H17LHqKl3gI67JEncdrEcqv8u
WiGgB+/HBwzc83NrkyISt16sqmpVoEN9e5nxcE21P+DCrNszzB7W8iSpEiqnqKGzbNX/mMJWTD6w
xwBJqQ/JM//kse9VNng7z3DUVEjK8N6vKxo3w+hKY9tsRLoN4G916lyEwGkoWnGqLNoT1BT+Jx05
I/DkD9CFEx1B2M4EQ99AqsOTYOWgcbExJMMF5SysiGFxcnO6sQC4doYI7iVBKcmlyjeT65AgkQll
ObO2fmstNzerc2+fEtw1ZxnEZT64mGefbxOsFCdcP6R8IctEYF0HnjfrrSKbusnKLGaaPeAi1mp7
KQxGuCKmy6TXefzHCsVNGgF/QhpGoPOiY7znsNQd/QlokBpApolWMFNfFNZe5cy3RvYefXI4U3nH
CYApQVBUPxY2ancUG7L2Bt1g8tbdDpFKkt50wtWQcKMRuQ+kZVN3Hgl+rtK6eiDIIrcbqONY9xUS
fiWwkSExzFfyCRGixhYHHgd4SuGDRctLU7/8vTyJCAB5cJMSeDDiWlnt/OqCavXsodbt1R0qx1h1
GaSoSoxoyNXJjO5aOPXhgcV4n4XLqvoRTwwhkhfkXJhHwwXh6Qjf6HNx1PgeaD2IRzluJ4VETIFW
K96CGslsJRsvgJ7VlcYGxK6TX44Zj1SH+pb4xeNZNJsg5/pdI/rS14/V3/oD/IzYfjEWm7XIyXP4
khmialKvgPx5eEVo+IuLQRSH4Cc3IwOvMopvhdNrAqj+G35eNhucQVOtFGgxdW/aDf0pXNhksNQJ
bncaBsmXby0i+baYND3a/KaBCBK5oPDpAjO9RFMihUTQWYlnapBvgLSRAuF8thtZihlpFtc72t3j
dWMXaSwuy5PTZj6eONZhitkPEHf6FcFHw2ubCKE93v6rdsQq5izDUyIZEnTnKvp3tSI3SECSgSkJ
6oIWW4L+Ja6tYY4gX7LVs3w/iqO/Qwjaq9XY+DDEYnq8XCy04Xgys07qUFBhq9VYpuigO8+Ljdm+
P8XyI36XIg5ie85i71TBFeoCEskpRDk9l03m57S4I3wGyNkWN2wnoUALXXPbpXf5wXdtWP5u2H4h
aJAxYqIMWd0JLxe7SUP9tPTXvzHbSzdySP6XH62MXlOuChNZSy34P9b1gJE43dyOwaFVIS1VQobv
bjyJANkhJ8FGJ8HZQeIaElMVT0QHoXvXfJHPAzeFrzXWz3FwrH/US4QLLdsPUm6xhZ1MSevvvqlO
/hHHSsaKfpgvyBN2GM1ddJyEHXhSzwfGT6Ce5k0mWj1LqNPH7V2haQe902BJN1vrXlixkW8EmJ2n
TJ4q+4Lcpoc4DQT619rzlnh6/EXsDdYw+BtPSYxrP0jOxjQwVGzgVQO6ycUDb5bM2QGhrPf7dga2
uF73KbhDmveecATRWbPByxoM50HZUo+1ThUZKQDQJTdnaz8nQLrRUcslHV6q6KkEm79Q/vGWE4dw
ZtxnJgs7EjRThB9yfoPf06SlipqFuPiapNcIveniPxajvQfHHW8w57GCX4TKyGUvVBIXMvpnU0U2
3QeVTH1C+olpEr7jTwKPgZ8l5OXub/4KzmVVx2UMcLqeowDU/Bc6VPKKAt2W5R3BLp84DlvxOEbf
dpeno1zLf5TiiUtYd9BkmylEk6MMUoGwLN+GHyhDV/LzdMmOephqhkplJKSi71htmgSG74U9i4+U
hdUVXDo3EcNADuwkNKMv2tlY8hLDUsUBWRszbQM6IqrYMlEgpIh2weIPdYvQ2IrM375nqtGrKJp7
utUyVS0aW/qQc77FXup5IJwdYEeWD+Qp/9IqUiDRpY4+/DpZ80kTjjtEuXUSdoHvjCiSA7+UeVoA
hVeDFM6J/+6Gpd76znmbySdo5hzhajLWQN+oWkiMcR6PwpDbiizFK6DvZtkqwviSjiFPZMNmHQWJ
brAAxNDDjQm/JjgwE8IqVGzGeIBxHNQUgkd+aZXKdBCXNWAaDm0GaOQkVLGv4D7Eh4VrkXF5OzDx
j+os/VXN5aVsFNxatTrT/6vNQEfmHPt5zgq3iNcuMgC+S6f5IyHJg/3ogwmg4g2uJeS/fkqE2+bq
5f2D42Ws4aC1JgJ7tNsT+mukLboG1mbsq3u2rML8h8d0UCoYCvzKzpKb4Rl1bUnAIrkayaSaMhDX
CQPHdhhyJd9LJkhhwkbPBneHoeDWhDRVJD0LYcuqpd6I8kObm4nXS2/W9zICgL/EGubNCuLtkMsD
j1xW5F312VwuchzjxL7E1DN/fJGIr1lmNo/SrHtXq3k+ioxDJcTLGF7fxtle3GbJN7Yv4buiLXUu
E/r7oGNUDc/C0kNs3COGblbRKsRhaqh/t+i2JorBFX3dTRrE4+n80mZ5v6XvXE/yuHgxOribmzso
+u+9+ke1lhgt+hi9Zy6CGodGeGrXLgUdYrbBsRMqDWZnZuwCSd8tuC95+PL29bLkAUgMg0uqtqHw
P8NVOJO2lk6a87+MhRvC7UvOZsBgrZyi6g3Ci2pZPTdLV99SfYPUPKI52yqRvYh4jw8B92xjw+0T
lb5knL/vLNPuI/B0lTMy4Yygs1Y14pUTdT9vDZxMINFOOaNbl6ODpkRY0FvDdVpJ4NQvD1sFKGdq
fgO7ISnupTN6gBjg76JVmh/EdfZrRI1B6WQVrCPeuCPPg2N3RYkultW8/DtnEYgGYky15zPzhYDI
Sg3kfHDgOt2ykzPMrXlCGimsvbqmbLJE2jfpG0jAN5I29s5c1XBhmTnzHsZGy8i07oXhbd9i3ot5
dgG+WZFpTWPzxmXl7z4mkZJCjbZ2YRN8/CQJ9yrY0aW9cSdGUE7cGltk+mlsuYn5CPPhIXOQ+0eX
95gHMKj7qJXiy3ab2M1s1kzU58jNo7bYS3emyZ9QeDqx7H97Nz8xvMqPPKStU2BdD4FmElBSltU6
U2EHPBzfnXCu0//UDgACQUY9syLDYamy4LIcNlvbxnYR6K/UaemAXBFtqI2nKtyAZeqeOG4sSTWl
gyEJnRKn2qG9wolz/gJNlmL8IZGUBZ0alPfIGBVTsw4AZnW2xnWjqMMgBccbU/Z+I7SDyHY9EMJH
17nNpjh+ReB3waFCTYP67Pf50to0cbUuKztli1BA49T44xplSiV6SrfB1eRoAwDxs8DNk7b/tn/R
4aP6EFT4OayKw9ny9j74YGkwWB4w+hEk3IwxJJDTaePkEOwtINiYytnxpjfCx+clHEJEgz+jcoGv
oBIDSmiLS3clA9DtMN2kGxNNuFiWfaSmWnxJQlYm4ni+e5ixD3t/dBQ2lwHE+q+mfuOylogG3CJY
pDU5lW20GPzcp0Rd/YP0lWPdmUy3kNBkcj8QjJnVwgMzG28s7v0zjaj98Kip1Mv/AoiWdLtyGfKI
VUxVbjNE8WnTBMcJgPeddF395qDxgQBS0Okz3R58IqNXg3HYzUzy+ZnI9f6OxFFYfzVUwx8qsSa1
KxAR3X2HJLT6t4FTeEMP8jwR9rzYiFZDh2amOxic0zRxMWfiffGYRqUI+xuFlpDnfKfpvVUAdpOr
C10mgb3gTwdgpsJ/KepE+H0umkYN6Hzb93K0PHvGjgsFr3Q9gqH8/LdvJeaXxpWE9Y/w0U0oVTb9
ZwGRqWxiGi/n61veZsYo/G/hVTvnr1SQmpv5oRXHIwH7LvVrAR07St0KytM5L3484YcAz4gUlYz2
/M8pZdiIiqwrnRNEA7VKlCc+Y3MGVFSxjlPaF9FyyQMYvvatnN+mouBZbYJp4VVN57g5c7Jmyjma
Zo0E5iITW2XDJVJEgFwtjUbVaTE7Nx8uxMN8t2V6vr9cq8EuWuQqZQ8jw+UPUKMZUNX2ViYqIk0M
KF8weNQEeJUrvQLFF6kzJBlofJsP+CMXWI9d
`protect end_protected
