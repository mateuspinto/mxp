XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}L�g���ۨ�z��ѠQ��,����r(��3Ml,8z���z�������ȳb�����B���Qg+\�K]�J��~�|��;Vt���<J�q�H0m	ϴ�>g�Cg�S@�L�)UҧH��"�_,������QE�����c�����v-��G���z�����ۺW�0a6��ӳ�����!�,#�5����IeZ���F�6Ib�w�rd�� ���z��v�0�9R��,P�b��H]�[8�_h@WO��M�)�K�*����x��5�=���A�w�i~ߨ��&���J�bed��'��r頸�z�����K΃k�h]�W���c��;Oy�T��to�I&�8+O:���k]1�I�|���e�1A�����7�$����)�Чa�1��_��0����ߥ�ЪL������� ��%K���p9��v�K�aA`�R��{�p>2�䩀L�m�ێ�	�/������n�V��"e��45�h�$6�+<%��UdY��l��OXU8��T��6%���	|�����C�� ���Ї\R�V�����x
{����-�3��0����C�?��}.i�Z��D,2��9�OTw�)R;
���_J�����e�W�U���
��e�uI�"TN�D��))N�d�F_쯾�h=�A��rd?QLq84�9H��}�ʮ]RFTO����B؉�'8yL�����D/�t���9�6Nq����H�)����z����$�Zybl�XlxVHYEB     400     1d0Q�!�ƅg�&������8r,�I,5�#�B���
�t�R+��Hm>!��/�r4�?C�;ķ���z)��k��c�%
*F�������R�1�n��P��.]��!]D����!���1��y~���Ϲ��t�S�AQ��$X�k��W��P��P;Ģ�F�r(R!��I��N%ދ��=u�d:J����v��k��k��+�1��G�7��˦ޕK�OA&a0����A������Y>H���D!@s旁Y�?��B&mu�"�$-���r��f>Pl���0&�������
�eu31��$�Hܽz��\��&U��h�-����7a��yB�S�:k%����4);D�eg>�=g�F�;�u���%���x��ڂs+;Ld7uX$�vae�Jâ����}5I97�w��3U�@��4$���߉ ן�W��K
�c�%i�M�Ijh�xP8@ ca�XlxVHYEB     400     170S� �׋�s�\T&՚��Z:m'����{��A�$�w�N$�Gx`�1��S;������Ux ^�%��lw���d]p����W����WP��G����(l�5��:�u��74�HӶI��9���g�j+������v��cb� } /*�O�-�X�����~ͳc�<fr
)��u
E�<����šs� ��O�M�2b� p����n��Eg-��ZX�{�i}G��%���[6��90���Y���-U,�ۄ��ʧ+�X���9��\��I%[�rU�F��l��Gx^ʀ��vy,��'�D��W�U�j���%��|ѓ�p^��M��4c���SvG)�#�ꤊ�l���pS�$6^qT��XlxVHYEB     400     120��r��B\��JS�y��6�p��N���$zZ��6�	ȼ�E�7��Krhїu�$���#�����X䅹�dTQ%"<xώ�M��駓�m�A+��W�yUY ��z�|�ya3���o�KĀ-V,�z橆a�M�����q�Haq��p+FJ��#�K*i��sߓ�`�00e��������ÉHC����!A�u;&P/�;n�h��Ԣ���89 ��]�QQ�NͰ\�>'K��r�L�wf ^���F�o�z%U���9n?Q!��whM:����kt�l�o��XlxVHYEB     400     170'�7V&��|-��Z̥�
k/
���%�'���1�|��R.[8a(����E��9�&<EX�:�Pl�rh
y�i��{S�A/���wM ��ei<����>��`��-g�[TjSV7x`k>9H��c�]���{A�R�|�H�wڮ�¤C	Z�(�(O�ɟ��K����R�'r&�@Cbw�dc.�М��ڢ��w.ܑ�Y��.R�z�nh�a���G����Jm�����z�>�q��q�3�o-��j��`s���יF�HAw���^��I�e� ����w��l�q�#�b�PE:6D�����'�"���	>n�l�f���#���Î��w��L�?X*�B
f	=r]�XlxVHYEB     400     170"� y����P�+�ҳ%���]������IR�_���)��7�R�����L��lK�n�f�Q吷��Q\
/�^���yp�����[��H�A�B�e�Y(=E��F�Յ�v���(��������:��P�ZHT1�[��VН��>�	Gs1��V�Í�?�'(ǒ�Ŭ�?G>���E7�/
��z�|Ǔd=1��A��-:QO@�*����p�;P�����d��6��]�͚�(|}k�D���c�"�8������J�sD�g$���_q�)
�B�1jb�����Bc�A`�F�]�G��y��K�m�b��M�T�x��ŀ�e����U�o�Ǩf��Ws��z�y=>�MjF&�BL:iGv�_<kXlxVHYEB     400     140\���%�.�����u4�V���&�aj7R_Y�Qܵ�ݦ�~d�(�ŷ���O�P*Y�L��u���t���%M�_!I�c �ش�7���dy�PZ�Y����cj@~c�0�K��P�$�������7���7yn�Ų������� �����*��ԖAS���4�& �nD�/>1jf�����8���ӗ^��Ec��"�)"�>�Pl ]$;uY�jH��4
�Sܞ*���}�$�~(��X�N���ibt�R���veR:�����iu�r�#��{�� ͟�g�]��c-)FN.���w3�B�H*p���XlxVHYEB     400     100�9%��Hl�Bx^+#�R��/�WP˟�۰�Q ��n������|��C��pղ�� �a���q�S�נ������8�RI:��E5>�?�AP�ƻ��e��iG��N.�;��36Z��D�RY��V��̠��X��L���	��M�Ӈ]�$(��b�7����;�[Ƥ7�XJ`���I�㾲2x���� oM(�Ͱi�zcH-0āy�]�;�|W:_�Hk�:�hO9�v���w��TY);[%k�']�XlxVHYEB     400     170�v��̉Ũ��:.�k�۶��J��('�فN�V������[��cщ�R���':����:\g����Ӓ&�*�%8wG��W;����sڧ�7|Dj��N�3V��Am�6u�X�AA �񡼄�!���U�3�(
�	iW1���K+����	#&��.N���b�,bv�t9�+������Ҳ���B'&׹c�m�����*Ɣ ���hLU�S�y�`l�")�@���;�e`(����~:��f��`��D�:�������D#	�n+<塕V<	��$i��d�~*p�.t�m�T/	6?cG*Δ?�Lw!K�
��n�'Qv��m�`E�٭��5'�szV�En��dw�P�XlxVHYEB     400     1b0^��)3��Z����Q�o���|Q�s�\PVq5+[��+G�Kї��:�<U��u��;���l7���Ķ=.n��V�V=]-�|��11�Hٜ6��t�7.J^(G�bQc΍��Y�ˋAT"�l�$���˨� 97�8��������f�7�d�^�G� 	�\.�BqԎE@�w견^���|#���zS*8���N:�_ֱ�w#-#p�s`�O��y$v��PL�����kFՌ`�I��CO����-�+}���G������u�J߲�����`�b��5�P��.2�и	�G+�,ƫ��S�M튘 � �ə��������h�qC[��%@.p���V��;�h��:��Jy@��+���!olPxoK2�M�4vś����̫íG�#`�Z*NF�?�
�m������n�����"�U��XlxVHYEB     400     160�u��jb���x�*a+��`Kfr�'���Sf̫(���}��F%��[e�I�G�Q�����~�s��+�;�9fY����0�#ցeRa9��dy�+�(<m\�l1�G�^uK�1e�s8�ߡ����'��������<��N����p�#alIGwi�
N$7\��_������%�Wk"��w�� �����ݰe%�� 8�W#��NN�Pu���W�_�hGj �����Pi�K�#�j�MeR����V�U����p�|�s}�ͻg�3Mގ�6Vh�|���Qs�v}�<��IJO}��tx�{f��p�*9�:"�G�5�?%���)�����Z���@^���z�yQ��JXlxVHYEB     400     1d0�L ����F�M�~l��)�D�+�	�a́��M�ؔOWY@mM>��fHw3���4!WG=����;&	�R]�[��Z�_¬ZM��:�i�y߿P>����&E�	� ��@�[nն�`N�χ�o�ոj����[�������PC�y��F���v{�c!'�,���=�>l2ǭ�O�1-�?�1�gT��
u�h���d����O��o�P��&��͍��A�s=��XtS�58ݺՔ�.6 ������}T���ı��`)�����-�V4NGTz�^jQ�R���h�@��v��¼����)�/��Bc�E��h�j���_�^HF2dlC/yzQ�.�7 �ɣ� �Qf���!ېU���('=qX���<���z0�{Ӓ�eː���»��ˠ�^&`P����a"��ҵ���G��������z����&�^�UXlxVHYEB     400     170|�5v	=�%`OJQ��_�����\��[=t���,���/�N� ���#3��t��'�,YoP�>* 7n���8��ű/�n�HX�qph�H�3T�h}��݂%T&�e���H������J��M�����]�%k--�#��O�F�������i�����z�)mM����!�AoR9��TS�������A�[�O��O�ߺ�		�]y���A�%Y Tݓ��@	}���e���& ���Y���nŴ�?!�p#S���g/1x�0�n�Cj�
�Ky�$h[id6���|���,>��D��tlo@������	t-�UDD�g����Bj&�U���D$� h ����b4�t'�	�6XlxVHYEB     400     160��{@�-K�\&���C"��kc���
"�eF# *��n4���o��\�H���z[�&v+gv��?�	?Eѷ���D�k2�פ��?��Q��j��XjX2����vh12��k��>�ÚB�|Ŭm�3�����*U3%�a`�۵�6]�a�b�ֹ�ƻgrgٜ��C6:7�����L��B%�Z#������1U��zzsޏ.��!�Ns���e�����[[ʋ\N����(���E����?��b��ݜ�k�.`�g �����W�;�l4��{�^���?i@b8�3�6��z͡�4��G���Ec{�]�W���.������z|P!�v���_m!Q6c:�A�H%XlxVHYEB     400     180� g�L�z�(IN�:̩ቿ:�e��	1������u��}?<�X9��~Y�};>HoȀ�����&*@����`������E����X~����ۈ��p�=��k	�c��4�)ѐ�O`���lF�$h���4�I`v1��(�|S�U�=&�������%��=��6񓍕��C���Z������nvt��x
�ߖ+e�І�x!�9���BR^wf�� u��=�}ө�k�������`��ls��}��v!cm�$�}��u��3�>l+����e~a*�>.b�U۶��K�~�Y�\7O��ʣ�b�߭(�G�ōW���l��=�|5�|�x0Gq�L笱/vmu'��&b��Y�W����#]�XlxVHYEB     400     130��i|�VWP�s0Фm������F������A���ߖUv0�#�`��tu1�� v�l���N�݅"=� �0%�3
D�a �t�8�m*��0ȋ��E�2��X@���T�[��*�SÖ�a��.C�!ԝ��� e��c��,�R/���&�ޅ���uN��nA0C/��p���p�|a>c9��E��~�:{Z�4$�
[����¼�e]@��$�c�c�NG�y��E��Dh���kSB4��Ĺ.BH�u6I�������tn%�l��ڙ�*?��Ç�R���u�XlxVHYEB     400     160J*��8�Yq<��y�#e�F���r1���q�7�Щ;m�S �񥻪@��D�q�L�M���:��8�mX]��)��Av���Ჹ��0%U�_�zˊ]�%�~����Đ�&T�5m�g0q#��(�עVU�_�!�������,���4>n97z�u�^���~fT�3.�.w��=~�	� 8_]��=p7F�>�Ǝ�m��ʂf6�������9�%C'�i��m'5�~����:�!�>�M�8	�f!�����?x�	�W�>�a��� o��*�f':~؝|TC`���	pl��zAal�e�ԯ`+�Ie�Xk�����5y5^��GU*�XlxVHYEB     287     130�f����Ü����|�x�R�T"r'��k�=��sǰ	=%�X(��l'��Ǟ9Հ��.�����V�$H�!�
P����{r�IOف#��}��D53��K!�A�*�b�`Tı��H:�.��k��������=p}YP���˔`�_l��,�ڠef?x޹58�� C]qX�-�5�Kzv��y�����*��:b�=�}K��� 4/֍+.���'�Xs�j���tlӨ���;�E�q#�R���YdW2�f��T�����{�)Z�����r���7{��`