XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o!*7@�$q��X��K&b`�{,5�1�ȃ�%fA���S8a�pE��Dq٢�Z��'�sv���<7G�\ �0xaI2'��i�\H�H0������sX���qjWtq�|���\֪����uB����|����J�cz����~��g�Ηã����'�"���;=C�p�䉄��X<�k�/�o��]�$�^_� �IH���(�����B�%̐�ڿ��H��F:�F�!Q���|��Sj�rI@�:[J� � /J\I�aɅ���?�:�|��H.��B�9ڟb1�}��	4�@�AQ=-lWvei�}Ǽ�qG��q�,��2�x��XL��=�â�v53�	�ͽ�;od��\�����C�H���|pА�݋<��t[i�� �_�\8���KEN ��GX ����^
��B3S��ѧG��?ea��@���XI����`��I��g-ݍ�����O��Yt��h����l�A�k��$ɥ��q���i�y��&ٻ����3
�?��>_٘Ц٫�oZ5F7��U(갠R�iSD��2�n�x�X^��5[!�K��6+��c5��1�໮J�m} T+8~-�&�t�7 fA;y���]|��Gs֮�h-	7��VBU}�Rw&��+�?!�S����:��8���Jj�2�Y�ʞ��cŞ��]a��P��.�P뚌Y	����NЋ�G6�,���V*�M����?�D�m4N�"�L�!l�c�j:����G�k���XlxVHYEB     400     230(n%�a��O	/"�6�6���@a���d��A���e�NFB�)��È;���%���3j<���T�A��F�nx��7{q}�
{$�ܱd������u�tʮ��r��z�,K
�`]8z�2��D����E$�?_V�t}A�yOϚ�X���V��M�yF3Lnβ��mT���O=D�6=-����Z̎�ﳐQ\f�X�� 5*��)O�6I�wң_$�G%�4C�7�_�$3���ܢ�� U����M �3�4�1+B`��Eu�r���u����H2�]�~rZ�uu]��j]��y���D��[�$`��RkT��K{OC�cTY>�u|��ٝq�� �eD��U�oٿ�6*��?w<`�Ph��
#�
��vGX0�h9��~������Q�b/KW��u�˿�zC�',��C����f��7٤<�AI�>�D�>6�
"i�����F�QdNi���1���^"u�%��,w���𓥥4�n�2���
�b�m�(O	�Pf��HtZB�kn\ҝ�}�l}�a���P�C�׌|��Z�X$�e�#A��ՀK5�t��XlxVHYEB     400     1f0<7bVD��D\+Ӱ�id��qW)_kD5���Oߑ(�נF��vT����� �hh��"�
�ה���W_��]G*�9��	�����hSr�,Z�_�'ŢfY��pm������3|�����$���.j��{��j�E}���ϳJ}Ӓ9�ӏ@:;���}�yai�#����� ���/��B]�
Qa��i���:`ϸ����s.	��1ծ{�
I^Zɍ�ި�$��M�r����j��	��T���X\kjG��f���E�;���	ƻ��7u.Nˣ�.Ebu�+H,	����m�)`@ſ�� ����$�5��J1�M���*��*ҩ�풀Q?=G���	q��+��V�G�!���rQ���\��D���g�oه�țΑ���E%j�z�z+��+��2{�@L_v����tP(<�':1*�j)ǁ������q�-�,B[�[d׿P�y�О,m`Wp8W�(ڢ��o���L��}f-��9rqXlxVHYEB     400     1b0h�VU����{~���� Kuo��4b�j��6v�p��¤Ӡ�hWq�SǮ�w��΋���7��_���p�cщ?J-���vI�|>��.� ���
����eS��a�\P���`��~�煷5��h�$ ���@u��,)�{*d�Gv��M)2��A�����uEF�����htT*�4�F���C�WP��n		�m.FI�6B�u�������۸��-�>��O��S��N)r����{w
�Y_;�����t�`N^�eb D�����X�.]c�a�"A#��T�p��[4��	h7U��ה�	g��K&�JEg��_6ծ��T���
�wݻ��9@)ˈ,�*��՜�܃��7B�dF"0��A={ou�F(Bԏ���0kp8k���m7\����wZn�䦈��1ŏ�a���XlxVHYEB     186      b0F���վ°m#��=�BP#<�\��������v�u[��v�0u_�M7��$��O )9ӭ!V���y'�՛4<�c!hӦT0�8N|�؇ ��e�m>�;�nTz�G��8�ٞ�h���ًbl��ᬎ� 2��	�s���h�'��7���>�e�0���%�q�C�=��