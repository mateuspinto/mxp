`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
DhPUZ8DVIj6wFyLePkJfRvNSfKIjOm2LujTHigK8UMzODKbK1yXY3juhQ8FzaP0wGw5Ket17r1o8
9jtb+PjR5p+GNCMPQOFbidMwLHzB7mM57I0t8y9F6rIvX4lju6IdaHKGY0Eju/ijC6s47gEI9KVp
tHjYOf8hxVncUjYeURp0qy3s8GF79KjvauI7W7/hesvVGDWa2LaTpsU9+4nzzL7WC+rgjeZHjguO
Xtw27dL4iep8OIwA1TJxAfTmo6WUflM/db7EddCyhLXn68oglqqr1Qxtqze4gIFNI3PWxdogfadr
Hcrdw6oG2Z4WuAu5qvHs4XH+pyDkgAuWTe9nexp0pRDnxz5pvWX6Zz9h30G5yVyOyctM3ieVBa3O
lITGbko75VvmQaF9WYxuu4o2MsjBUGeMqapARXE9H08pRgn3VkLauiTzadnqnUkI20LKkFWHSDT/
HtRb4IlKt5hMkywJrmQCkl8KeYrrKeXKay3yzBFOcynfBIPfAVg2jP/rR7tiQgbLprXJJzfu2who
CT08XWM2bc7NFTRWpGzcs7rl8p88iN+I/dEUn3Axg0OdI9nxDHA4Piu3XKtcgE4odHV9H/EsUEte
dA/J+33GB3E1xP7cKcNzbF4eqwZpv0dKbSwnt29n6kB6Qxc3dAoqn5Ew/akomOT1ap2De0zU6CE8
NOuoKohx+xzRFW1UotF0SYEsjWHWU+vaWLtodabm0zELxbX504dkCMtWc/V9VMAtiiJzfF8jCSJT
HO6WKyomXtJAhcvR4mDifuI7WHigkIGakatUJasXJrQBZFoC2ykpCbmF7lVBWBMN/QHi86FtS+wG
8P5ZBoNgqfvRn5mLJNA1jyJ2JpqSr30WQG1a5wR3a1Wd7omiKMmCAWYsZroR6STWHvrafl8vWc77
8z5Vx7Ta02vcrSdhzm5Dz10ta3SGfa357qW4bbYuFZRj3QlWO0M7UM/qmu9ci/UU1KCbsv0tf93X
kFKQadWlcNBcvH2MWzBiEzIeH6mkHforE56Y3hJf/iK7ChlbP4m3DWlW4aotQnU0dD6nbd5Zpsr9
qJQSJ5idR8hgMxMCNcYa0Qe8SJKGa4x9T4yDdMXtUSB3TW9DZj5ReH2rdUmOppD+pRr2ypD2w3GR
NYmOkCnZZqa42OeKE1zszytaPN/YEx6NA8wsnczLQeBIfJ68lrRJzAWWao9j1B+XV6GqBCoZUNjq
bqC4oxfddlYtX8rr3j1Wnt5NHjXxx4luiYaH9GLywi5O/chWTXuKIQQs37xHbDES1ATegFe3ziEi
Ef/9TLq/LvpXIM2ZD8C7m6gwb8ch/ZhA2Xl8u+5Gd+O9SRJu/yG6gComK5iEynDGBXIcMlajFGU5
zncCuuhGsSmYGBaUN5Gyem4dwWqfWJny90pLBCaiegdpMq4N4DsoZ0b82IbbmPLekMoLHKRXifik
/gIfqNvgw0PO5IASp0zy9db78001wQ+8hPOs2zdKLj0V6BOSg/LuJJaKcQECmXMS5X5IvsRIFcJb
m6zMkkX/l9PsdUoGLydJjz/pUKvpzJMOig44+rqmUxs1B6O5f3cwJFufqibk1wKYDcN+Fzt6s7t0
+wHgMbv4CvTks7Gg77HHsVchK2ZtgzZsYUlGD/yAqb9OrBlfKVkw33FwSasXkjY4+HavuPow+J7O
7sadyl6q2w8wYi/+vJwJBXNt57R2Om6SfTqSxhEHcfiZ5GNJH8vGOJ/ZYcOPZbQ/q8Q++bpkhBLb
a5HVAjdOuCN3uRTI0wzZcKUVF5PoIRwbu1GpsAkHC/1EdiQdM4LDqZAyIMF/jky3vFU2U7xFw2SI
bbdZraTWQWFXdCjcVkIXa3weNgUf8WNwblls41Utmh82lvVbyMMw9PSiPKrFDdWR0jMTPLi3ZbW8
N3/bptDkxMCGDHBS6n6UcR3LnBR7wtUFE7RvoqFoa54iIj1ZBK2b9bYg6f6e0BvYdB/ogviThpsm
r3AtnKv0wBzK+PK6fu9oG6Uv9DcC9szwE1iHXlagL9q7xP75QhkNi02vVevj/quAWnfUl3wUzRhI
6AlIu8YlvLssF8ApI+5ATaFJAfDKT/NlxylVjrjGiYm8wZUAwtp2n4D8DX9m7/bVl0+pR//1CBOy
DL+sc5ZFCJOXRES2/dkyb7Sv/+tAlevow7j6x90MHyT9q4J2kqE61kFWrH5zltzpeA69K6wtX24M
GxR7MU43NTt5PU4CWJcsWbKH7HlGFWxKKU2Fo9BTOxfPbjS6Rsp8DOwCwE9y85DT5NBemNJctJKE
QfIjxxUTZHjctGpDKTLGQJ2T7q8K6S0wLXvTjYAQddJXLGeFD1/7c3PLo3NmA68py/ncT2PlqKen
vdRjmJp2Viai5YLM31M5Z7+wjss1YuG+Ualu6zscr7MSpO5MBcwhCcvEzWd1w3S2D3bK6J/IX9qc
c6nLVeqqL8ugtvEgUhBfletOTWTtpJkkZ9v8Ptxwyz915LEJFASwpGfdv43Ez+cT5whsvlvHG0C8
dwhTgvSBH28yJ0yFx9GqDd8EpKTJAJDDe7rl4G+t9TDtuYp3u8JmQwcrjSBOYK912S9ME1Cbqj5K
juK/MrxBWOhDPENUvdKVUjtVhP3d07aSk1fQJh4R1ca7MZOdqcPq5e+Na3StkQOPgbGb2TYWS5l/
E984TSxkSblJ17lxLDkXwo7lQHB1UxkYTK4qvNHvHEsIV//PWupqI5nUKTHn8xGMPWhPc6m7Ebvc
21QGE7tKqEJS46yixB/5isgJmcw3wKWZWTaWX3nvg4M/Z3KO6ry8XFlE2py208dgk+r9jI09zVDk
9Ykc5O2XNBuECU/y0gCR7V00mtuha3Bh3GWKp0Ov+CCzFaR614jBwnsUdEue1hVCH+ODVZl7T7f8
SiBzQS/eeSY6DudY5WOaLnhiyGyqgfVyWFNZkYIsp/ofzowpju9ldtMuBYl06kRWFveAACL59Crl
xc30ybs1VwjKjITt6Sm1dhNazxUG9NFTfVOidbMR4wK9bEOe220H5heJPW7+rKUj0KA0eEOSZ84q
BieG76r9ZWzmwON2BxRA//yz+uOEPgVHIH9PKoTLjSwaZuRdeSNnQBH7n6qJJ9pHwb62TVf5ZiIZ
1QXbEw3BiytTBE4vvLkXQnueM1EqjFskODr6p158DfeMc8nD/ZbmExVPrbHkkkb/fshMBQppYPal
6GSK+AfbwgWvB7xeNTbZGS1U+RxrhTaS5Ck8Ptufw8ZLNiWQbHoYK5qeDTgBixxmyj/5eNibFSoa
MLJ1ZE0n90mD36iAcxGAzfizd16ozLQrT+PHa3NnxhXtnrdjid3YR9XAzJVsD37vbDaFd8z4NTUZ
PICG6ZrZeixBcrBWNkCWWeRDAWID+4zfC49bluSA5OYae4RYSmaFcXROmAUXPKm6p9vO35c2X854
2IKjJnrsEuBLMM5inwZ6SY/JwStUximeILMqRdIpvfb5XQ12ZfL3zhWt7Vg1JVWAVYIuAh/H39tf
WKRJb8GDA4doz/wrYZjoc8gfFQQ1OFGyJal1F7tIXcRNcQJs7SX13ISQOC/4FWvcYEyAhI2jEqWj
ZT0H/19dt4GWiIjZepmZGYmkm495iAze4Xr8AbAB0G1Ce2j+g98pWkK0dG31EkJPPtqkHaNr2FuJ
OZjKNz3SAdKYUJhGoPQ/D4rnVJxR8KQeOHYfN+Y5U5chgSEd3bdcwinWAyMdUgc2T5NJj0JU5XcD
UQWN3vW0hwlAwhdmJLHjt0BR/CofDCiaEGyhboaW84JzlnhCqUM9nwYtk04K9UFa9ZxQF10W5Pk4
abtiUnMry7yAGRRd3OYEoCwLO08gbHDNbya/Q581b3Li5i/t7BIj3rA8612iIzIxCzAiE9ftD2qf
OsTmoggK++j0+HBHIiySFWEEx5o5BCqTqgr2hUDz0NYl+XJd5S0G4xsnCDC7WvSmQ2spqNMe1uhy
ToOOKDJjMV3WxMOEwc37DqlY8s7c05lCncftrFkxWeK8Vzx+g8uZrIBpe+cOgEon4yy7+y+HFams
/CuoXBX06r+ZcBGRoMaQCYTr/Lcp+2NHpP7WInuYneYugPAYK98LUzffObWgI7RvKMDHCXg57V04
ybU05N+RVV2TCd3WzLfVekuJ6Rhw0xCxl9sWq13mRdeXVYdg0bHXoQfGlroy++73H/tzCMMt3sdg
jrO+dnLX3wO1SpJEasoXqhDZLjZe5ScYWi93950ZANMw/5NO2BGiRVAfa5XpG25vz20LskSubaT/
H7vRCGVV99O+TXol5Sl8BTwm4tdepI+B6DJpgkpgfJfRZDjnF4dQToTnEg0tGzzEF1dKhblS+pqF
zwrQ/xCGq/h+am7STMyHwfezZ5v2uyGPr8Hq/Z4fMBh8VexKXIWEIR3WQ+0xBAoNSqkGOWxFhIxD
ETIyhxN+Ut/YJZI4isKlg6AUYa+IkT4v+JhAjZVyoeG0Xen5Sx1iaQdD3zKSNf4f5QyOjABQimA2
GX4rqgxPsD/bCXP7zCTopb3OthIdhiaxll7f/uSXuyQGyN6ds2l1aIkCzulLPItmahBWPytnfoQu
jZ2SjsSSs9Cf0o7oQmGiI5LAQgCeSRwoIECWPNaD7YZ4ZzSLs5YLwszNAWlUJG036XXDd5L0yxh5
t3VmHaGN7DMQbsF0a9XWmgqRA5p+rprkb/DN+uEFAz53i1UH8CL3TrxShE1g21X4GcmWjTqJuTo6
sXQEEAh+6uMHQRCobIEXzTkw5XUdj8dznWEXVQMGPCZriggn5bUuSTRnc5G8Petz66JF7JIQ1ifw
6Yfk5Nw2OgrlF2AXZCUMwwCz3cBdzMWY46AWHaHHlKnBqX0jY3fiaJdgFcBKzsENuZ8AosQ2boSJ
ED8eoIDy9oNMiBU1OgWD9jFEsnO58IZsxFcqWOD9iNus/9PL/94IduaF/dNdFzvAS16Sj4VHXzNo
RrnqQnnSsz8+b/UZzfAzic0416U81Bk0QMnS6A1pfI7cAX6d+9iW6g0dIAWb8D6d/g2jQDz0Mjta
CDZ7UjiOO3548Mxi4gsChx4BpdCF6L678ZjNFT+ilpWc/IgLXrEv7kcDh7fCQFQgF/u+W3gJt1NR
eXHLjbiytVxGapITqfHIVvafuFvMvR/O1tpzvpwWrdmeGCMaNkHthffRg1sXd5qrzA52YlelQmR9
1OCUG7ouGWV63P2+PN3LQRoBgdJxU4aA+i49IMfQ9CGusmPF87mF6EwDSdztg339cwpWpcu1r8d+
CQV1RQcd6nEoPyTjPFUsZwjEsm3GpxnjqQXv8fqe/96bbPAZqJWy4ycobz9sHFCRY9w7ae3c3Qwg
WVX9LnpOoQteBoVyRQTaCtvd3yqRY2XGdZL6SGI+n8R0xbFsGfIjpb+FUgPhIbrUM+BPAhTDD83R
YmdTuIthzvgQwq/5SfCMjkS03xSJO1asAPNlAlHuYVM6FKI+7Tx9WRdV2KYrz7mz/QeL+bRXYi3m
CiGVMFEOA7aQ/R0J9ZtYWzTXqVY1zxLUfvUP2+6nehx/MWOy1kEeq70xoLNQGvfrAJ/BJzK900Tz
sGT5356IELVRBTE6hYTUpkS9uGysA8Vi5BzlzDa9lMR3XTt4M+Q1sGdeSAvptBBgGsHfLYGpeDVd
DAdTYjEsV5+2f0JSe9RT/osM9FPdroj9+nRmwv6K+VGBLw/yzVXDacd4RddpSmNg4U5HifOKN61R
1crU5eRcbw37ByIiKTvkhR4Q6zzxXcar+ByyHyTFJ7ztuQUXhQGwA1HXJfXlXNfUrOPCHGpEFhDT
7yifyR6s/v3+cSR+5wwS7O8ITWBY2BZANn7fseWA5itdK1kItguKb5K3fDb2n8lMvVx6G3QIcObA
0q2+9KSibi6JxJyiw/Cr6hxlDeyaAL1wDt25NEZ8ZbVGko5o53tWN0bpQ97ERfkD9zJUCAn2C4UW
GTGn3zb/c+GPHgtkECkB/h9JE237kIhTJoR9niIWRGygiI88go00DQ5rnYjvuL2YQkMS8CxufixB
YzjWJvNlkaxJaGvoAtU44E/EX+VVsIjsm0OwHkyPkmYnHcYGGBko0/97vKNFtXOhuLb5uLJavaDh
znC/oPRwhMDQMqbfb9zHGQfG9thYH5xQVbIL9XpZiAJARKwG86yQ5RGvCAZKXDPcjKYp0xSIbO4q
6lr5JJyR1B7+ymeVPu+hraefH8WC0hE9pJJHoYXF7ZBZvGc1q83oqfzzt1CYNfiLM48xhCRiqdVf
44M/SomegXAWHWhcpj9RUwzCsygreIz03wzEiZUUOoTmX2+kXCDxMYS9QmkvNqswvl9y/pAv9wrT
X87G2D9NI5Z4TL+jrJYkLbCJ0t6MNFM13I5dk/bgNSXDSQa9nYRLMVrADbUr/aGQ18UO4PDaPCPT
a5ZRhIyz5OOvTGuwUy4P4pbxh57NMlg75YU5hQBPOo16+LYtO7b5zA5fAmjzBKYZFFHdMtLbuUDh
jcSbPOR5ejQOxA3KU0vInd02NvZLwNKxT50XCfBQb2AxQGa0nyPzHhRnVo+P9r0IEJqG1Sym2/0H
ZGNogB3reyZ2eVSbzk+qLwbppHNKZmka+PcCJEMKKryhuhULrL+PfXzgKEBL5xr/E161EPKe1OjL
KPLzHhpEWZXiAwyv7k9PyaZKmqHW4y7yB04In6DpQdRmShV0NcjszIV4pUrh72RgGauyGZjdNhar
IpffeMm2JJ2OhczkJIWMrWulSZN6MRW01yWqpcxsxH/JtjZmljg4sJuvuQMVGt13GDF9DKEA2LuA
7iattewQK/cAkmYkhDA6y7bBJVsT1UJTkCg6AIpKlm4f1OLMEkWWteqvenXQxplNEvCpejLASIYi
arKVr++3R89CiN+sZhwflbl2V+uBECWrKx+Y01RqZ954VBrF8L0601RS3xndEXLGI8o8pA4zSz01
2nLL2jUzcs6hbZEl/bcz0cImqSnoVZQ5Y0ZHniLlipu2ukt1BhxwrUWw6cK8kZNWQQ3oNY75vm+C
hpKGfxAX0AtKPgFNOOCgIkaeysMxYgV0dHhqBHBPLS3Sgr4B3LSu8NT/GgpLYQJmEBQ/3frnmStq
2clSrF+AwiIsTigE0RYYugno8OW/rIhQNG44dfOPwuvaIEK5aOzrlNgrsSxARMCYtpDimkMBo54P
WLQQaTwZA7xMyobe4LnbpJUPlO+sTffyDdXBlchvq+QROduOQaByDTbiC6f8lp7CUVit8jH3bVtK
WqY4ls9LUu91O/YlTj0L9ZCTbXNn9nVdNuBkxPGMbmycjGS6r+aaUOWDzUFFfnzzQ+sq1OVvjfWW
ekj6rm6vBbUFeBRiFwJOILMCzS3wkOzkEsDmAOpJY7TzwLT5VPlyo7vO6b0QNUmtbEhMUy79SbRe
bwcF30ElaZO2Ozz/NkKltTyzPlyfIWqvKV1MB2xGs2EP65R0iIFqUTE1Gycx4SpbJopi2eJ5uJwi
vBBReB/vA4CMHy28C0dGPrrSS9zVTwMU3QqVK8zozZ04pWok7P41AXosPh+PKOGhZNGc/RIWfK5v
SMS9S6629d5Ktb94ZcmNjNyog11j0FZeAmYY4wPDw6BvU4qdvolbDpKasfW+shJqYtnYVOpXat9T
5xw32mAbIziyQ431ZKXTckmozrlUuLSfn26aHBP0FIkWf03Sl1ojT2MCOdXwjWPLFRbCd1mDwSgZ
hkpoDSDpVw9vEZjmH14iItj57Z0jH90cvxnaRE41UhPZihmm0G3OwUpyz9a/C4tytur883hYDUUX
pNq53tHLYSoU+4eAfx/9iZSVFVfpYP3AAddOiw7MQ/uapcSEr71mFT5VnhsqSOMS69NUdn+PjVfb
k58tOND0e2wpbOT4fheyoXU2+csUKngwhn3K0jEBghe72oU33tECTRCdAlGNWwXRHYh3HMqNyo5Q
b2gzH23o9neNmKDjj+3kJ0fxiQ/pX8QFW42eSTLoGJr7KogKpfXoVFas/AQd4v5mvVTD76GGvpiv
ByYVOQEvkLPOzG01kwac8MPMWVc1oyvDGJ4i+WfJWXJ7+Ho2Y4UIf1jCKYnVvlYFHTS5QiqalzbG
mAbkKnn3AZe1Kn2f9Qf/HNburE95hTAf7CDRtoiBfpkYUkLAPSH9b22K/pjZ6FM0AOMTzzM17hHF
FKlPng1LPsL9/V3KDzv6Sjb52EUjIAGIp8g+xSkLY9AVmPdpF75kJJ8mvtgOTTl9Pdj94kOF/aRm
UceG8P5Q6k5gG/6EHXGOJy1aU0RoLiJfVwbLEkX9Xpl8GtLuMbn6B5sGV4vv08nNnbGKLWJlJu8J
dwBj1fekcjkg4RdD4PES4juO97yi1+kTgnk4A7Nquh6RX8S8C+dDRob39D9Efc1TCAoYqb/G6oea
HE22wB+CIKZrJ6IZx4SqAju9+BFbPbO+LpqEBfS0XEbHc4eqdrsqV91TqVNB/blo2Ix3SerZTQ/t
rSzCYL4CrV5y7NHb1YVZaqB/2mkg1yenSaywJPTYbvVd++RpXMbpYnK/gv8L4yBJaBpAEnCgYWZe
NWXzH6+/0Af7YoOwhjJL7A6eZcL9KwSq9nQJDHNQq5x8UCPycuufXTr6UcCRKkNe4UbrM4AbWkUX
a7EudiaR7YZvMIm1k/IVDzgb3E+zQaE1SZA9Ma6Wb74Gwk3t1ehhCxYPUw99fOHcsD4jgZcBaaIf
bEPpuh3B6ZEHzcdbidw4yQYIzG0k3TwQUwlGmL1U8osJUn6v9Ao8QpF4X7aLSXUBRIJRPMGDSac4
VV519tEKqzzoNkcCpOGrOLua87JsevpawZXjINBJzTqJGeEab1DrLBXACgUAa5gbwAMdSwRsEmUa
M9/GKGObZg0Lok3n9xSWfLAMvAJfUprIl20fy4Dh3/7VTbX6oXeO4eCR/cpm9bFVswh50Fu30cDt
8k0jhD2xnbRLdILZ5T2SxOIcKiPybOpCiHN1WToA1AYXqVxvbToO4ucqeFJQ1OSLD+2LkKWvP8KK
v1/jOhn3MYvnF1z+ZlLOf5eFeb4DR9JTcUQtXcNvmamm8e3fIQjihlfw4RVuru3Ryam9ZjTJS70o
HsCynNkihALT74+ohvfTHuXWLQJcBwUB0vduvY0TgwJvTucLSK98GAZMQdggKDBGgw6QL9ecRFGF
pQvWPVmpxHVyd5l4vt/0+KJQbhogIvpBnDKDv0Is0yA9K+33yg2AtZRqb1RKEJZyivyxbWiIaxrI
51fp31KNAFO/HaJGsY3FgHO0ihdLtkscXicy561Q6BmulImf2fAaOQuUInYbmX59rnGohT6mthI8
llJifyB2FcP8r8u800pILd2J2pi9fOMtIlQTMOyXSual+SMb7rkoR9SKJpRtgsTLWdQEttLKa2a/
8ZxxAV6jJpja3EOkq92nGVFdrELCTT5UujLjLc2GV9YbIGuYC241BN4JHO4notI3NVMuVH8mTAUi
WNF3mniVzPhecy8WRXK36KKFBr7isIsVFGogqP9fbY2GC5M5c7J0F/CXs/GggjObFA92B1L8SubJ
ytcJd5PwX/+Y/O7e40J9B26xc6skWemrT1Eijf+6NK9ajZ5THveJWCp9BlYpZZhSkZVdCtZ1gcwh
dD90RA6wEYf1N+UXbqZrLAGcwZKKUxIz5CSZsixcowUWjnqDCuB2fHrIWsITPNFDm7He9TgozgeZ
fwAaTGy0RSUGFARhYZrBuIsSc0gfvLMYRtKIlWiFsu4CS+n4nqo+GM35elTzhR6DRMCbhk0bnIp2
MmQAG/364TFfDbQBeoyK8u7nDhVj3JhMhpQORvK13lE37+emdTcw5tGFhxHK5xv2aX+OQRHrbaNS
+Fg2ScA2Chr6RdoDSdKVai+IO1i2qhvcpxtNH0JO3qeEaWVVs66dH3KBQykhD6hdgD7Ws7+wFU/B
CUbDAOTcJ0SEzKMRdo9pD2PbN7sHUHdVWXWe4QJJCHdWCmyUffwnYeUtW03ZWux5xXtokEkTNwSV
3uWMvNUfNZYn39WdkcTy2FwvLSoDLXhMxwniU0lJlxKHxhS5k/UP/cD/2vprlVpnQjWvawJnhCGt
GrL4CPcabYbrZk7h50lVUf4vSNxRHOHHDyv06g6ma2cj3/ch4S+BMgLRHB+LQWswrs2jJvtnFRUJ
cMIXbK7STJtpxETAtW1tG3UhF8Htd9mJr+AcPv9qK2g0Fm9Y8uHJpbm8LJx/gesWZDxngRfaA/1E
WYOk9HS+rEkh0o1tAIiwrMLlnXVj3XKNcJPq0BFcYbrbuy/s1TajB5mOtlS3NHpNYM8nhoDRUWm/
vFSLU1nqv7bvMmP16N40T54HvasKrg08rdAF/7XOO/3TdedYWDD4Zo3rWtBwx5tllkhTN9fT1jIo
UcEQohiTKtAxO19soivTwvCTtu9+/jH8qqPuYToaUX2HC00+TKGE32VsxmhIAphads7hY96RNPvz
636cSMyVuvhXXWYMKPsYz+uWQeUi8CISIquESyflW9ybNz5eTn0e/A84mSVLlLM2XBSmG/rLIl1T
XUZMHAGFCPBcshNv1USamoTqq9Q4zgfC4FSfs97Xc1tTP/gmsIQSMhyc3yDUEjsJkjrVojIj/vTN
4kCSK0VonkTm+VMPLefJy8PPtF7QkP66YT28upPegecoGf8Ps2pRA1x7KBWn/UTtW+Rb6mYaTG7L
fyJlhUNAC/CE8qu8bCGguz3LTC21Q1Rf2Sovmt6nSU/GwaDY0rm3Ty7kMUr47I3j3GYYfOv97Mmn
n13DpXn6jGHO3wkHNg5J1G4+yeXlc8eJauEu7gSdNtuhWNRtRAsPyZVNj5f+bvP+DucJCo/8T3ji
2QoPAzvxDoJAxjbA26Iheu6KxIdOMp2jJQxuzvwdMT0XJ89+t6YCgLXGsO+Azb25VzMwMgWtyoCu
HHX98olgaaxgWfZt5T/NocUlYRZpnAkaRGoXSdECHaSSpCSxcNWbTwjHVM/0OQYTCCAJvTGi9yI7
62JO+hO3WQGUw/RBHnZ5FIEf0ZODP5LZXVm6Gan7GSmoiru+nJp9LPpTpXFaJsfrgFBKBlguUzbL
BKqtafqg5hYAjIRAPOCIkRNsFEZELzn8RKai/1R/2U336ZfxdqFlGBKfccFB5ozX5UWem/RdwL6h
v46UA6cmA9kUtceUoyZU+ytrkTr6bOKt5YHBnJ3iQZUtqv+rmFsRNKoGcrdgAz8ShuTl862gWwvG
BRxno2dprya+E7fuVI/DwH5MEAx5LSa4Hj3BiJznKIhQ1eFiuZCRgZHiLUlELkXka4wMBy44IRlW
6VEA4gEEdHNMQ7s+uY94BMyxMvjTmO3b8jjDpBaANi7zitdofVFHg8i0VINHxBFAqLDVrGlm14zb
OLDO0uDJquANM1NrnZOuBNeTGbprEjq0BKmLXj0+mM4TMll9eKfV4uJXKmMcGDkx0M9bdM7nac8t
EwGtr9liOHTb+N0EpVZ1mAAt42PsMFuaWWiLBkjOim3daxBzdXq6ilNKnsU8I5Tgm11rQTETUeGv
ioxdQDgyZvf5HpORGnmBdH6ntq40a7S0u0s5NUWQp1I/svVuVtsGubh2s1hUjZvDsz7WTg+TCfIb
nOxwim/k3Bkrt/vjpmndQjdLGUezsXYM1Vt6b/6/PC/VB7UWh9z8sBQR/emHUp+I1AptF8JUTPsw
KhklvtxNIIft8vFH5VazzoYc9bySmXkWdeMpVvp8lOV95C+oLm6JN88TjwNWWtgzD+MY9mzEOlNS
kDnibB9y3vvPPNW1yhs0IOuUr/rowbfaS0U2t79zp9ZxkcbkW50mvJrPwO98xvVkcybB0l0ZOQsA
mEpTvLQ8XSJoLYGKzk2D1a3wkKM3+X5fTO1agTUHDtF0tNHibwj79RsC5iSUd1Ip9fpTwJmi3DyR
QOaWtxmc/zHgvWjHQr0U+3fYU9cFed+7l19QPsBZbcjVtdAdp1bqhcHvTA8/A1MMd8/rkL8avdsr
MySQm7U1JphhJrZVXbKU3FlQ+mAgpiQ4zashjsD1QrtMbxNoYEdvFfPBUo9XBhDr4UalWAy8B+c9
7IZyOsPJ0R5nLtQ60mReuP2upCfY0b/dE/slU2mtIZWy4cVQAMG98+3x6nk44HqlVdxRfGKfMXXr
qImYX4bf6NSbBB5wrZ3TbC8vtl1w8F7BNPebsABXRHu/FqPcTbEcLiCTjxcUYoqMY1JaBmKlYvZP
3x+VFwqhi+viy7GQVgjiIlaZZVQjWRXDh8IijqV1GDvwnDa8NuMw8p0BHWAOHUn2jljmuELiHwq6
dW4+q4Cqs9B61rDlZGkMFUuo/2irp4rRXTWFrOzpGisYefKyXSqchvxSKoEU2INSHNwSzvQLGMHL
NPZiIBtu4RhoDqyv+ILGdKfH7hxOzWXzcUKCFFV+qgozlPJ3l/hjFibEMhzSV9thiempnCUxYLqv
jPpKHhQddovtFpb4PGjZtN+r5ZCAbLRItq1oJlF+msRm7x6bOLolzpFFUKENx2p23047P/+YVUVE
p3gie7wRI60Xtr7QLaEdAZb7q1z9KeofrMqKU5xhu8hlQ3ar03F8LyLiItZkaYFopw+X6RlnFQC8
BQGNA0jWyJXMLxN9oGXbf6lCNrilgIL4KIdUjD1gyHjpaMmbSYbqm+Z45dBLFRUwdYu8E08XLK5u
4U4IV9K7m4Wk65EiBPi4/LMXaqFOooPWVvuXMt5TPE6JdFEBnGjLRKjYt6sd3Nk9pg2If9GH/+EB
30kRTiXAqlCatKTh8DLZHi6L3kL08YozkGUUWGGnn0wMVgjkPIev0R/TPtijGYApZHqO5Zteht8Y
+47xn0Wh34YD3mFmqFBWoOi7W/2dx67tKNHjOlmWWEzn5h90Yxk3L4Fsr3nzEaDobHn7fOt41fjp
iN82kO5qMkZNDiBm6P04PiYHYuQa/+THg7Um8YRI+RziNe1KHgc8ze6c65N64yMjv15YsaGbUU4c
KSyNIr7UxFSM9Gv6rBW4oEI9lkhtY3Kf+GoucPnQPNkpsS5U5iUtAXLbpJe26GdJbR+24C8zv9ty
sFxqmnKkxpKeeKRdkxYYdg1hvBA8LPvhhSN15kL0ypqFv1fFyg+aJtk55Kz60otBJ3Dhwlb7a8VS
wxyn6Ar061yAXWOKJGrpn7ipzlLOVVSnx6QIGLsq7KOsGpoVHUbYKMfiA2pPRx+inWfCIb7vUMhZ
L8z0sHrWIpAe8B6BaHqZ7GwStjSt96tpkM1gcKattOfBzF7P37ZoacZVQOEBCC3r2EkQOs9YkksE
YKvfVAtdAP8+ib9FAeGG9be41CxFebEbBkbm2+ohSC2KFEccWf46aj9YGYsgIYyeb1MwUdpx2M5F
BnK/ImZNdqe5djrMYwLBRVedu9zfH7fR0ZzIzpf5NMH1lOb4vwKMMM0jxbR6NZJNsKXsQ5twL5XT
aq5VHbzZJoV2PziPijhtj8CEnZ4QVx+/MwSPwFO1h3fTZo2L/b7rCjHPOqJn27e0lPdtHlrEDjYY
RfvhwbWndUWDucVH7DNOldpEcoFvqoKyygtkzbSJ/ZO51tzmMQEikrnsnxD5dmFhscul9FHMby/a
kqM1h5OZ2nJIH9o0navY+wjw0I3EqjcxByQsA+0tRd+ABv7AeO+5juZDDO34CcZDvHJPEZgiMiwk
OTS/OAGwYfa/2TwtKhORo8pbnpM6bqMoM3adCkt/XCckPcxDVXgTpOu68qOgxtvY3g4ZaFt+o6Ic
8RlmBpvTbDHeelx+P45c9l33eqrSpF/V85tHPvdrrplQwJEH62pWpn+vbKPTEQKKRCGtMJGbJyCZ
IGV019hYUOy1FW7Wgcl+Bbl6U4AEioilbnru1KtqNbPkvxcHb7M4DoLjqW8oEhNte5J/7FB9pg9i
Z6kKF4FuDe5siWF5gd++2saF8bcQx1AYKu6BbFt5bj0CzWtV2hH2KTHnnYEX50rlXa0cFJAJU5dG
PndNvXhPh/Kd1g55zj0yRcaN3lqtgNLOSYQNNV3QOUHIlQPsQLWPk8d555VmP0zDQmy8A6JerZro
NMsPHKVlFa3qM4I88oXMTULq4BzqM2ALlZQ1OGVyyjoQvczhJXuUm8qjGbUCfepFCjq1czY/e3tR
Het4fYb5ukYknutKPuQ5ofazssAVJPJtu5C83sXydEpUDtuCbnISkQM4L7qviDI6sXR78ehjDkjB
y3UxayM4A9JMMWqErNiyG0npb9Ttdkr5JVzALYDiyW5LSjo+TO1VWvvfYtSJIfud6pBlF/clNo8o
8llGZD6qGCjZ7usveH6EUPVfZ4r1LVmqV4CnLvuLWLaGMs9eFgJ2B8NN/8vq6wETfUfAWLEw+bKn
5eEbRQxhW8r7gM1OcswV1dcwnmrZ7QG2TI5A6tu4z/c4y0t2qIrwlXmfmO6VkVcmqVMKOwhzlvHD
7SgRtMPQ+OpKUwHIpltSqOk+XJgTBZecaT17aW0oGihA+66d8AitXTaFypbmJ/8ubnUupCjWuCDB
dqZAsJK18/WT0XNWLmKlSL4tXM6zXVb/nAZhP7m0E6lEkKCYYuyIzvw1Dhcn65yYyP3EsmSyLFez
ZvHEPciw+t6Wd7sVKjhlez6xGu7ju0/3I7GBRiZKk89MTRvcS58a3TVBZ4MauVbOSNcRmdwljA8M
d/B6t4sJhDKs1r/gfz6DSQ+JFoInlg9bkWljPLq057nOc5Qu1Lb66eYOnxJYuVWMUfNCn4EjbJJ/
LyiveBb584gxHr9EjGKSB40b2B25W1Qj6qV3BYRvXE5FxXmjUx3Oja5gJq+f2w1OabQ4K5xyHqIE
t/FPbQVNa1sxVnL3vLkKTBInsTwt61v0MoLW/51umd4YGzQRu6Usd0Mm37EB7vVKKpSle7XfUjkF
UC6OrVItTLxOerc6XXsMaDg8qvwUNlLAakPVnf/gnh2m+3EashJKXhreE6CZlqf2feq5Ehxhzx0t
iDRtoqkfQ3qwUGcQMnlhatcbKTDp+R1nEL1GVsIw3+Cpadp428Q3C9VJn0aRbzWNXthNZQQcadFf
sK8lpn/C6A8kgrMMmSVtzg3pKcSAaBdv8YBeOL6UmWdXK6Rvh3fAUNa8nVvGcHGcGYKj8Jd5hi5T
ldrQn1GXfyeE30zJPwmukXn7VnLDx2TJaNRxVhzH7O9avyABGyZdSTom3IM70dWgHssKXaoovB91
/bBpFH3jeirtojt1ZcIfYRbuOq9u4M7RWLKQWSref3sFOjCcO3iNd5JOQxsRdcbUtJapYbCdTA9W
oxXbw/YPtcxv8AT62gAgA+PR8KkJI6H4jed1AELaQCZ6iqptgQqmlYbkjAgG4jZHvIyses09vhAC
JMOzSXpqM9Oc72+XPE3PABYTCUqDOwnVlJWHXZeJ59J0pBw7M5Qv7wb/zdGOtKZjdlbUIrHOzRKk
pH7HVAlvQmHlMH9njCAaDoz5nsPvb10q523HuGmwqFqv8jJh6BRsn9JCdjtFAYEQxoaKsSQ0OT0z
sGsLeVdpsfCunKtqolKOXh/arJgZVDMbmdaUx+L/2Z2OBWBsY/LwVZEvdO/3b17wE2r6Jjpo8GGr
BhMOm4nJ+iT3pi0lka/wq10lJq0PuOQ1yU4H0StYd7xingvPaEl2YDgLQLw4tn7K98Qbag0ZA+2r
b99krp/A2xXXEgSGRH7CN5MHYMiEcO5j51Ip/t3zDDfrxNNvDbxDbd7N6140kG+iEt5rns4xjGT4
ADOfhxrH9zmCj08gUu6we3uxDC5Wa9RB+0XvSRvO/lQsl1N5OK+sSsG1NGHy7y8AwFgLSs9PUsBK
K2YdZL6l9iXYtHVWsLCP81CFgu2IftzDQOsCFr87pL5gMg4NCqmzugLR3Tq8dWkT4zBLp7U/jsZ/
PgeF/9czfpO+ffdjyK5Lu2zd802thbaM4RYsI4q9QHPhlCoyOQy1iNFDtB8uJDiNPcW2WuvW6KSZ
HJdAx6qWLBybaJZqLu1cdCTCDxzvcfifuJvrjSK/oq1W5xustgrTvqJWvdIFOt1kDgzHeL+BoFLL
3+n2fw4T0aM04vYXuxQcwF14ri2GY4EjWVvYtIqaK3LHD0zFRdqqCzOLJ3M2jka1GZQ9JYeGP74K
xmyCDOrZuMrdiTYJvz2axvUf4jPKDdqAlxrHxwpUhZgSy1UH+s2ljbBWLQ7XBQHZ3XMxOLigpfNS
3S2IEeRpq4xtsd5bSM0edBjo3eNrFIS2Jy4+8Ib9LQi5DYPc1pCyy5fgQ4mO0bjv5C78st7KOEVz
WXiwrEjjKYL54ctyzm6Iedu1UKhy5mXkk5TJw50Bs2wb/gSpaLgm+YlN5RvUHP8p6gZv1H+3W437
3z2DsBSMrcT9T2nkSngZOuoIrj1P1pN58dbHpDkSSVeHNtsY2rWGqQRHCTB1ejzH6n/rhYNJtHTG
cUxDYpzVFVw60TRaJv39Ha1Na7QtEyJCNgp1T1hTxS6bXPx7eFPVSirghIoUDIeTKGvbHjFkLyRN
wQVLc+riKrfSb/7FYGdwjk/pZ1IHxxS62B15YakOWr7vi6RIV2BbNRH2ry+xQ2l/VawgdOryWg3f
9bfsAbi3fKchr7tEGwbMla3mgNIriLyQJUoElLlkgPhMfEUNe23AM/cPgY8DUOsHpFF1JRasvC5f
E4Aj9zPNhehrg9b1l2DispItE/ue/LYC2l67chgaVKFU0SxaUuHm4DrdnkAX0jV4Dul/TzMpy28G
6LumxdN7k6lNfr6O/KCVcEd4/5qZyxHKDGuMoUU0SdVwNUtTZtPh8nq4wYQU0tFEFToaTJaZH8pc
VY9SSb0lTCruq2mV13/Cbn4teC+vQKmgtU3gAlkmWkXGq8Mvzv2VISvhzlvf5ZS7+lARGOJoofH9
x8jEgzr6g9Ru6e2zCDFyjl++jUM2GtKRRAovC0SfRP+0JNYqiLf2CJQBTkG3x8kLU6PaGNRGHFk5
rxakNLKT/XBlU5DpJ6xkntomfspY9NyUer5OUhmzct4eihDx9DLSQc2I1kxNlmBxQLtHGCH5A1R/
axQ7lU0g8Ob4oJhOGAC6BP4Kihtxzj5nPTFWUewDqKDzUiBDHjf1IVRZMUWFGLtsVF2Z5SPPvvBc
Iz/hZaXf8QMLypFZSFxk/Ru/j8OOT0hZIwGpVyJpfH/l7eR9gECYU1UPhR8BnEH+mh1NegE0U1YH
tS2YHyKJAmJxLsIpkEYX8OGD240xbXHTXena4CXPLZt4XnavLERQUvDp4hAID3llKzJqlg8tq7js
KnJN28recDWXImm1ZWmPO8S/1Tm7WhZHdEDiUyf+mL/0QNFRX6tX9I0IHv8rsO1JaI2W7AW2leiC
25LdgRmOJw24lccnQ81o7fTaPETj/HbuCiIXXlgmVuLR2hEEKeoVsr7jCr5hRnXFsVu0gv15qlid
wpohPeBoUloXt/4vNQOsugIiV4EgB2K23Z89DyDtMVpVu4dZtjPW8sDv2/i+D5H1vtcaSyMvYBRc
v1fLngLFdz4hwjReWbBJOEsMStN5RwHsulATaR84IlTRDXfQWvR5j4iNEaaPS9OCDUpCvF6yLyBA
ATLfG+oZ/Irfijqx2u44GUzkDdmbNaTFepRnlGfDHSsDD6jIfXiSmY20/67RC9QMKLu/Q3dhqaeE
bgMiiLqYRpqlnOPgw/gjPYB9g1J+mIFaIlltbINUvkkD8fB1gNc7bDSG5TkxFoyvsP0tcRqJvYMv
SzJeSiZnYFFj8B8K2PkVKthJCxDZNXZ34k2CVFgw37v+3QlErPQ0kYxYaQ1wyCAIWn+E3rsxlLv8
dtcXEo4W7IxykhUtHOyAlvxp5DFn9s9nLp0jhxwjCtFJSpjxnXztavkwsCc5Ab4a/AhWwQLRxZmU
qDXoYEoQZ2+CMttBdf2JFzuDnDkOQTU9rwVMfCqP/mgSkf6JWzHITkQNG7byPbTRPyV3RA0LK4Kz
tc7bDALPF73DrkBnk7YHlPi52dVHyxDL4hTBuD6j+0fVZlYlbE6d6qKj26Uxa2Tjulao6pA+pVYK
9xzcmWJIstS2Vm4YfsCoiER8HHQ+0DQ68buLtA7VDsqgpKwoPOsjSmPVAs7Y70I+xM3nO6uQJX8n
XmMn+/fV6nTwDCiqaLH87XElLC29kw+dlH4Kazpn7TPHkH/rUYxjk8WcK9FPho4wKnVIz0xclG+0
6sywvM7O7wkWIlh1SY0yAq7fiQhEdkRNIZgAXTd5lsb07xgILJxV7rpGtYQWTOg+cMGGPqLJTA1R
sVnEs5R+ox3df40D0sb4wDA8RIv7cBqpHCYX0L0N7MFOdI/fIzDb61+nUcFStnkeDDorcOHXJTi4
HGGw6RkOAbJRcBWNwPjTkatvm6dbJWcfRFIzgOxmsNlSV+1FSfQg/J1CkctGBBZPtwnXl52YltO6
7HniX+FwhomCy0+5T20sCXoy3mdXszFIn9WD9uj8cv9YRHFNnFbavdWm1T/S9CcnQH3uMuEdJhtq
GpmTQKYkx2IvM0kD3mD9NWk1oS2Dl2uVT+l36gD5zgUrikjqthrTJabUxb/r2ljEDaFR2KWNp3wf
h0/QC0ibfFdrEUdcUMbM1pJO8fSoOrK9LVlAEgnuXE9R1thSvthkfAYViw/aNqcKF9v4roiVrrEj
V7rSC5Df8U8NRYOZ+ro5NOiq4LLgBUZcKBGg2lAv92mn0dMMPJUYLQUI0jmzIIYjqiWl938OQO2L
nWCcF/8kLmPBUZv7AREw1J/MV5CGZAp48LDem+OHosESnhehw89QG+hFXELWXO1+G1e4OvF9NR0R
/lPa3zZpfTpiU86/gN6TeiRB9rC9d58wpNL4qY/MjPiigAzRpjd4FFhRKOcK5To8pJX1riMltxl+
xT97s069YEXu2XHZQjdV9u3dplQbGOZXWSn4U+XCqHg7a83coo+PCuYtCGp1N+ICGtTbDcJPv5mo
jdluElyCEZs/oX9mxJjEzSBTFNUV1L1+0l2pEre+8VOPXWZGmP5zBrD7W+HJYl4qN7dRQh1qxSK5
nppwTK6rAXAlatRZpCivJabdm7XpNP/bHcjMkw/bm8iPVl6PPGnTTTIVnALz6mQsB97M3SfPraGk
kZYY09wJjFXWERqWSzcqc9gxMJJxv19mKK5fr2FkpND5sJw8UxCwHwfOqkW1BZDr64ELwVWMTNtN
RrbddnRadku+A5q0g+OZxVz0yBwXXlZ1JFZam9SKRRy6V0GLkDRQ5a/3kr9JOpIjsa3dB3PZi5me
29mT2dRo84TVxEGxgHKdn1jH6budATBmbwqCMDN3w8yHsIlTE+atJHCT/34nsA7mCqa5D/OtRrjo
JcmXHv1kDsEUVJVOYeDIxXVygIygn3jk1eOSSmVCFWBGhzjq+WLnbAHlI+1drY+z9S9frbeI6AdO
WOY2zvDzxeEk485X+eCpJbx8iruccksiEqjz/Rxt6KQQwwYmkJ10qU8cx6vOn7+PApsCVkN9zdHk
wJ86F5H/l8LjXM/ha1w/dxrhTnb8wCpodsmClTpbatmPAeYvSfQOFcWBYLKQ46KXRAxb+5EARTAp
kgzwo5hVhjcFwTVfUQzaclpInQijtePg+FCN1vYNm5NBPQQV1kzmUeDhQFWdr5WeAby4aOEVG4sM
1nYYdaNS1mVgD9cIue3bj/U9yDA1C+i14eVVQ0Lnh8Bw8RS3sa2gNVcQC3HobtpV4A9QKfP9r4OV
6FcRyiCmnF8UIjmQOGldcgRZpB6niaFkTxZpqjY1XqQ/dl5/R9ir9Dde5IzT+eHTLQgzdsLJ+pfu
iT3gt5ljQDaDKcrpNsp/uPgAL97i+xSJdIoeIz0OgeLDWkBz9MZupWn2npoXKNKpTZCADLPWfYo4
ID8YK+bdAxiRoI0SxVe/oKgYwhbbI475LOrsvx9lLWSJkq0xP9hr3GYadclsr/7kM0xMVOnEPUyx
hUdGW5yNkcnPBV6JYu2Q5dZg4iBCHix/vs1zji6miHYVywHJhDs0F58JMt8buszZuFH715k0p8gI
kORaDHjDpkODbAXKr1++PzVADgWQl5MgRe5v0Wp5LmcZgVdGUcjguOZ79C/a1Vk8IlBR1WBUvtZI
4S3a2MvV7bEz3JfTeB4x7R7DpONUU84nnrKARN1XdpgTD16YrVcZouugdUrNx5ivaJAd0n1MM9NJ
YMa9cMEdYPUu4tiWqwhtokXNYMRaY708ducWTDpEHaF45l1+xhBz9LpsPkaYcqZyj9Op4XpKkVo3
DHXXfR++CRxcd5wKbPdOMHJMmqXKhlCJ9GJIi7FsW23rjis2NwVNQvC6j4ywSWbrYLpBRowowpNh
mnS2nqHn0jt5h5MGDMA0+mU5pZ+UdyAEmBHJW3UjhK6ykyvKrhySRYoj+UfqUhgjF9gdwKrUc/lj
ji3dq1t7/6GwshnuMf9z6DGkrNx9BbVaGCYmsobk+m4s5JxVrFFXfB4XxtMCzeVWsGrCegxVF2VS
BsWGaI5VrcNP83KVuT/EY1NepeEZ6W6rF72hjWbMxno2XIfc1FOe4N3/7A0wUbZUHwYhaailHvEV
LTFVMu61C/bB7zJTDulATdnOetUEuHxxA3gBCkaBDPIPpOSSUv+8LkxdQUbCGKiHGVRMZpvTFqzK
g5G1Q5OWJdsC/jqg6/UOWhm3wuVOSB5DmwKpEvmRPoVXkTRw820+o+1IfS4g6ARyrLUmloGviQVC
L209xW9Rp9Mtwh26I7I29b8ZhdBiG7jrwU8m/PBN4cnWawh/mpnpZSxqGKBpFjCvXw3B14aVEKpp
tVbewV4a/khED/4jt7ijCJsp7YP1jDRqrmQdE8PNHh0P5+z1nWtDiy7BvxU9rOQeuB8vPPfoErvq
ozQGp9lBTEHssz+ZupVdEkitIUSA4eHlQt5A5XfZu//jNue39G3k8DY9V6OVVYUWmPSroxZsDnbo
YJQ8TxaT9+gRYgduUTGU4PaPCd7irPggWw2dysHrlEB9mwL4ynPftVw59oWUV8cnCes3ymdFIx/q
IKPS+FV0qQgITdHPKgzpSrMdXg36hycQrM6KnCZE4rJmSvTSPu2r1R6oP0KCavfyaXNvG8XnDCLT
uOhkc8GwSvlKfOKT0qtmYXgDYZ47HpA/QD8S7iuy5xuMV+eYrwSOh4KOdCoIEcjsqXmjWpW2NizB
vZ5xs7HUqiaZG2arfR5gsTvpnENMbXFl6fPwrzvrEMaHAIgrF1sgbZTgt5cx3tL5ofSmfz99DLp8
K5mYSYAbpxWphZooxVvt0VSLr/HQ/tGtIxtol7xC4kaULdfkLD8J5WqWYiBagJFmQgejIztNJRfu
hAA//mEw5d1eUH/IQBPwv1rkJE4PKe8smYTs6alb+vNMRBtb7K04LAp7i80+gehcXUjJQ2QlI9l2
MIofvHA/5ba67eJZKCZo8jOMioSKxU9ROmYr6zOTGP1IyEoePbWhO3W+KGzUUuigYLtAjLGAHwnW
0R0VBwMGeNrUlTRSsJQDz342UdvgGZ4qrUxkVfvzXUpyDeaotSImfZtYZx9RWEVoICDlqGjRQdvB
CaZzZ+UgpCIC92ZxIIiDVmA8OMzIZkvsZy7DILrua+VR/EJvj8evDAy6QiM5uaY4SCFPdV7RsjhP
sDDfVNTG48012roXy48GrEghonPvqe8t3TvTdkbXH6poMF5kRbgAb6hT1FAZgTu+Z6TcDzVCWEOS
enLiOKp4aHA9LMvk+Rm2GUrPsiFyivi7/qxJ4IO+7Gr1lg0yxQbA3mWBreeMtgwbH9m0OcSW0Zgg
A7Qt/XEuEDg6duqLsIrGH/NhWGvWkVlBtNrR3LeVGhcP3FeorEaNac0AE6haBb2Y42c6yWriEHaL
jrEWgyNI9oiWMhF7HxkW0lwZ1f3WnZvbQtoPx9Hh+/AxEhgfJbi+fQRYVCOXwqpfMXS8QlXk/xbv
1idwCh/ZeWi5ioyTwD3GzmA9Ek9tBQz9pyGhD6st77Q59M85p+8KquxysyewB4t3G8egjw9xPZmu
cUwMbnlkd+uLe44YAhKMZxCVKogyMmDI3L554MG5tJ4IuTD82tGI5QQv6+DGf1lwKr1CWs1fNbpO
tJ1tOPATlbKjxSuY+9iq+EnmbYZzAz/dCxvibgM+IHBG+fUqA0gDcC5CUGPMtE9NeNmQKccgKaGy
/aDTsnsxBEOzMtJn0/PmesXvkrD0maqGN4QmcooysVs16w7a1W8hhzcqPZlLKWlgJ2D2MgdcghKc
QhN0UVVXmHUipmK876m+oHvNpaQcToqBG66bQzLreW2saluF4eWPRyEzQmWuM7AjgW8o/OZ8SS0w
ovepZ8izbkSDrwYNtS7TZxlj3G0cH8uEt1G9rgX3HRKh2f3+V/t7+fUqD/GN0l5RasCej9J6YvH5
vFrj2unMEFiOWjY5DgvGIK4aJmAMgQReKnT/700keB3B9DkZHjuWOQ7AYnTnhsmujKow/y82QaWy
kTr7n4rlrAhXG1jRD/8Zbdqr5dL6yhQVJuP0lwMNRyemdoVeamkqOsOnAm0Y5q3Nw2rUGRtqTb+H
YbF4Oo+fZ+jxtP8R/dry2aCk6K/eTgMHJrtRwnLHIG16+VT/Ww2Qtfi94c6ifqeb5moQxvfoSJ9A
MGG1Q4TXccY3jarm5DOGsC3aipJbrjtH5zpxVoOB4stuJvWXKTVB43+xH/Cj9hnuhdm2PsRYRYfz
zuqPXwBIGa/SKcPNksEAONTcOu7KVR5q9e3IOW9gPAC4i/USysyj7dr2a08LpFSzhtaRyCqKwe/z
fQF+FuxbRH0mpvgBXl8RmVdvoH2fYa5zFt7cqEe08VPPktDGKDUqxCHnhWve4j3N4j8WOaEdyiVr
+1IsfZCbV7Dq5qe1L1s8YU1XNemukzlwCnNo6ynAnQT5l8irrW3+/YAR6N79p5k5fhwaM7mof+IC
MFi9EKBu+fwsPIaDUzeYPvX8cVDsEc4AdDofpSfxOsxB9OIuy6WbJ1jzNU/JW8YHulYa6GGomtwW
oiAW+SKlwB3owBpQgEuvqTIVE16E2rQGuuX5l9AqX0g0Zd+T5OM5uGLEKqz+BkkPLi5Zo+csHfhd
jIO6u/ltl4GBXvmNwc83J2VqsoJ+UaUo2zuFRUtGIiyYdMBlBwnUUodyWvNTdMWyN8X+Pp5ohAGl
hpqdkPSE5mVEHEi2YB6ky7krRTtkE1AiMnu+hM+efULwD9cusggOVMlA+PHaBQJJWtQVPTVyzcop
njFQKBK7td88nLEBIzUjA61SMMBSlZfy+iINvjh0u93ZO6i0+o1PrAycvrQu+f1XNw2rrqQcB6CJ
z74FnOCacXLY2DBKDH/HurlHc8ba1LjHtS9Q2dWxdsCkodqBSeVrbYfmKUdUw5vPSBrmQPbK9d+Y
3vSnOao2HSnBhZziYKiyOpPzZQisGbyUgOHauhL0goODgekfiH8euFQhWOs+KY3V7ZurPJdomi6d
BCGAjXMldB0SY+ZCgLwFhYxxWjsUyJ/TBLdxO9ssdzDdOMHRb+68Qb1JaJ7mgn97KB9A7UsQOFw4
5O41ZVuJomnch/1i1qZzXLmcMp+xrv5bDKnOmhnxTmIxBgPE+cDiqk79cbXS360YBzR+TAYOQM3O
wybINohYL7z6d06WAbvmQa8UcztY8O3LQlFw2mHtp7chy/lXF742HyXe3bEH6F14zuBixZP5t/XX
MiXcfrEikGSWJBc7D/SN/t35MYruWdMTGTKzGR/bXqBmTfmgAFk4inZDYUhk8r5qnHqAMWp3yrts
OENiGhA0yTGzKy2VHKQatGxUjXLryj0MsXwTxT6jFZHUMWeXEXhXvtXvOwplheQwTjXuWqXN3xH2
yMdkR69K3F8f+O2m+n+cDQ6ZATZr2I7+6DOxE1Wxm85FG76UneI6gjHDvJpFAUYYjqbgOU8yra1w
CQaHwz2fB6TSsJOft0o9BBgpDap0LpfvSgLyas2fV8sR8ttKXIV5qLFSdDrCPe9NQVtV5mpDzKie
/ouXbVwq8U+XzsVLQitNSqf0Fi3g76KKKaOa/xVWoTfUPonWoH+QSZCU8KQVwQ6NduDnYRHzppur
LY6termbOyf8Gy0aYLo1gTho9f2Tkg599H1STthCfWXfFhbaacjc78IqBtswrWvC+F3MUEWUEYG7
P2zWMSyH6IFXN75xwhWCVvBWGZOs2esiiG5gCzNSuiiY9ZCljtlxZfB11TQgnnSGXnqMTpubZo7I
Ju0i2+CzQWFjGKR0x9QTCGi5g1Gjfha+GeqPMWQPmRJXtRqmbC24BJ7gS3T2ImuOf6PtyqhYV2+Q
QBR/ThN0mG43jw0hHdVbzEIol7ET1YVedPG4jE54TZsYYv2so9w0QxmB16311moV0NQ7Q3NPVN0x
3kAVuzeQ8n/aaUgEnCTzvMgWYv+eZvvGWgX9pEYQYck/Sa+CpwnEaWIlNfrzT2o0P0gdK563/jc3
nJF/bNHevHbOuidIPkd5VGvLyUI9cCCwtTl+ur7iMRqoAx5pTvzxEAwihcgifJ93OgYwRk9hr/A4
iWN70ehcpk0lU67Ma8fQp3wckAdZr2F5Kera/rMSHbQ6AQsv0Kkcu3wtjxtJ8hHvYzSjQQC1m+xI
LkQpuuTfFDzisp7SZL3+TzuBZtJJPDVaPjJcUliUXkRWvvLs7uOLMssRGlwjIVKrDpGQApvKjl3w
d528PEPEcMo746EpXQIY+DeNeqe1OfR8+mdheWHC8V+CUw98hQmmSMuz/yY2p0gcIbQyqMNHCZsS
L9GXcniSoHhFziz4+v0Blg5NYyLRAsUMxjzTUMyw7+O3vTtrRGF2w6ZfgOLL0nKvBwvDXh+q3J1N
Cco/neP7Fl2k1hlFTvePArrxC4xMbxCWWaaX0DT/RTXng8v+rMowE1rTjZ1mfL+KDYo1oEQt1lHB
aztVloY1G5zz7Yqhu+R/K1tdkyeT6Duar3EmjkVDTIyYQxyF+Z291d+Hu/Ow6lpTCjXpR8i//TSm
CAaiMFmItzZ31zES+jIuKXCP5gHN52mf6zQ8/Go3AMT2BVvjBT9rU4SMc2g2edw9GW0JDfCv7SOV
k2gfxg4Qrkvp0r1syuG521jfgXed3u9zXoMM0jUxCWyPsGm04mYSgkipAE59qMedP6g6kSQ5R55P
FgTrDvc6iiyh0K91yCorU9b5IOJ0ycYoOvAoj7poCMEmAdxZ5tbREZXV3IW4k7ozRyEKoc85VE16
rFQfDXF+BjPc5izqsVuBheWuqZ8zj/Y9lKqNQwQZ2LMCZmiIpRZ/mML+uVenkA+8eeEZtOOiwJ0C
LNDaVTVG4y4fjYPtN6a7PUkeBGho3iLd8jXGrHTuHdLJxH486CHm1TI3VDHY+GWhUmmG9XNjs7fY
uDLInrlh8h9Z0GVLR2uLO206y48/hQTwSm7qNg2Et85VEc+prMAnVGc4oR+lezTOPK3BlQWnJuVT
MEn5JfllkFqIsRtogx+f546ofSz5zcpBuvyeMMSXonOFJdtMxdF8oCqrfGK2Yc7kscdjxiZc1SBn
xTz7Gx8xNc62UC94A4XCFmQMoKHel34SoKFED6Ea9u4cZG2DVx//3kYUpKZhVQRQny/A7PptjGzQ
zKlB30aQHOcLrzZiWlfvOAU6mvivX6Ccxc+98q5NSGIJhFX+YYXjPwWQM/WlIAuIuOOzE/Kd1Nhr
c0/E56C3G6NHWIZOE/dfRQnF1rDqCG1x9IHkqYIr46vHYEHCXiWqgW7FOvZ+sZEJatPXlhq5ybxB
Te+q5XuRUurX/h+HGeSZgf8yPpulMCx3mb9w3SxaMnwbav3nbZ93qXCZRcFCX/mSJ0sCA4fL7xlK
OR/3Lcy1VMUtKjIhLGtHevgxZyYg+6Rrbxsw49GBR9BPScZrAaHeV40sWZM8/TTDFHtNVbpwt6Ez
RwcaALDDJpWEELfUyux8gsbe8Bdov5jpD2nzhidQSgNhgxHxftn9dyuy0J1iP4Z8oW1Nc7H+JlnN
Y7Ruujft5GKh6cd0+jejpp9DMWctqjkWVIQqHxcHv7lpxo+5H85ZVN9NKqHxlIs/DHS5Jb+kxvwk
afihWR4U4xxPNpAo2Q56hiuaraKBHov02sNqxfy/HVveqhP+4dEuAz1fp4oMIFE2NAKnifKZ9QbJ
V+0wMPhSEM/N5gzseHfCsJT2aaByrWEfke64zxV6PdKjGts6vv52OKtYmy41lBMtqLVruxRJUYhh
vp7iXTOyeWUH5rmBvO003EKVaAv4T+yC5iT02Nc4jAfoVRRvwy3coB90f0uhH79G2Dgry7ovU6be
FdjMRB/0R1lbAD4FODsmSF3EuuqZYBwpQuxin/fOCHzbL7RhhuZtfbkpuQK9Jne+it2wmpql2MPR
o41zPuitbd74UmrSFS0+VvGGrAUXaVv4KGfyzIXcyF9oYKujOiWn6JYicV2cRP9SUb6Iz5UU9Lge
D+IKAq/lTKUlUCGeaut+vHcl5qxgYOZyTpEy3qEBvOr9eW4JO8YVtFmdimGkDHzqbfUMt55tEjVQ
KdDhb8+zoMBtTgS4R8ADTYWhUGuWtqxvPYq+mImUe4cZpiSEmYoG4dJzkS7iqgvR/Lx4W9/Pnw4B
9g6U8AphhmJc5oDEoJ61egafOJvf1NrF2puUVGLOnappf54/DL2Rq6FLcCDJl/Vc6S1/9RAEVHPX
xhqiAnhfefB4a6JPlZrpBUsDuhp5rq5S0+dR4R1rB/GlTo/zRDtb5q1h4adYRAZwEV51OzQMki9D
yoGRlrbCwPxWtvpZvHeiizlXmGqxBnbepKoK8jFtulq/jiAwBFsxnZi4VamdxqX7+pdIxDgScnI1
tYpfXaJ5SpWSuKJNcxxKmBYCcopkuAKorViJPZZydQ+G05AzcMvwgqNWMiFnsA5tnuN3kRsSnc9b
PYmfnW6mJNzl/h5H9uEIzS0TDVRtWK6iPBAocy9r0ECHsNmKUMYLkjgTslSnlwmIKlUuomcD+AX2
VzySjpZxak3tWBmCwqMLF3FGuGVUxKhsB9PVtnM5lVxkxC4OXLEHXb3E3TxB2waU2nLG4Smw0iiu
E2kBRzm7UM1a56glL+l8pviTyvXc283+frktVPJhZCmDslf+KnZkRcMvxzecfw4bJXQhnVMG7831
VLpYxJiYg4hs4jnx6+rJJlSW1UEj3fyHsOqdh5nXELwoTO1qR3T4sEH37xVf4aVZYrOvqnKrNKgM
kPY/dbEQjbyPKy/AXe5yVkCRr+a6BJs0GGobe6Q9y9fKJ1xgEZT8JNlu4vUxXvf5IBURFAi2oH7y
X96vYQSxZKzKeRtLwXPQaPfoMLB9Y0EJ/xK029lk86hxDDqxsLpRamuZg7OeUejGWCjjyeONeS6Z
izTeapfo6ynSVNZg5F8ltwCrHDVVHnS1d1ryHP+zj7B0yovjhUeMEzVh/H40khEZHQP6v0axgAE9
F2MpWchO8sCzz2588Sf7XoRk+Q3cm3PRJg6YxjIz64rLyemXu8BNOqHMeGzft75qDir207R6Nn3P
egzUkJAOJ0v/2QUw7D+5QzQZ6oJ4EGqruE1oXlh+aIAgVD4BtD6H/sUrSqNZoAB2IL/jw6ES/7Dm
pCV1JdYZr5mFbbNyOQYqQOChxEc7Ww1e/11gMIADj6p4B98fRESZG4pfTxkDw3JqyMs+LMKj7UUI
9K2/kXuHu39BGneqS89Sl7T+rywJPaxtOegeu13YUakM+BCHvEEF03eoRhWs2KCQYtfzDSiw07hF
LZbksYbJlkMp9l1HcVuXCeftV+xawRoy96zwh/gcX3iCkm66ivmiRZ5ABMy0f5HB7ZLJiIL+JwHv
27Jh7Hg6Ww9VF82STRJxGYY47L/YFYRyravOqqTD5Wu0yKX5zAvuFbkcBe6PYmZ82dEJ6BQRiczr
srwf5cesrHbVSIrVcb+HuDUn5Yz9+EAkMIoTiBLkEuRD8/c+RDN3aHSyv69kPwdiJW29phwi8Ltx
9C/e7AUurhnCLpa+ywGvd+kAHneHDeGFHmllzVD+/BeAmSkQstMnpyJAEXNc7qEC9MfSZ2I4cT55
SClXDAzb7bUjfZweTcyMEnnFEGiKyp225mMGzc0JIlTQrPdtY4XA3FIO9ORFtfzlhPSGozcWezMj
SgnDN6AsU2XHIgH7OoSdWqyl7Z3gJA9S7+Jc9u8TzCpYjd0xtzZDnaCs1Rf4yV5kR/Sm5m+QaQeM
Qosqn1/y0wf+J0KSi173R8dMtBFrkRuTtrkpFWB2U5ebL0iQnOQGeoBcZwG+6gL5G9D87zqSi3RD
nB4/8nlaz/e1nU9n09hm5Tsg+ibvDbHRJfuawDD/J9Qn4T10BYGdCFPWNFuK/FP1PYpx+P1eTWTP
+6I2MeD1MVWy2A97Qq6MbkxRNOVR9zwrWhuD31WKZ+l0ktGPwWSWWD1Z3dhbI1idlNAtJfuCzQKs
iYBN21nbY5dQWmlbHQjRMVNdh9qWH28m9hpKTGlH0CnYtkSgc3OQ/daYHPBZ/i9luy/FLyUS7Ah9
6SNNplF51y4rnxuEfkzh4urYNboLUK5WvnH7LV9wQ0mL9iRe0o+sklA5YbX4XfZNZLTj5AsO/QmS
pAD4wzipH3T+ijdLYqyE+0rjSaBx0F6AWZ38ZMsIEqucZI6TV6uXaHhRUpMDKdei28Td+O17AZQh
lPQ8dFKqrKgLewjlwwnfSNEan+z7lPysJE88G3/VJa+foulugrnKgCelItF4Lfys4G/cjlP7VT+9
ANz5IP4UmeswN+7USUHoKzcJQHjX04jcu+AEjEAuCPUeq0BPMYSaBDtUeXKcflOUp3G4SL21kkIv
as/ipysPkGHRn2/vvVKRg+4lg+jB8XSQD+qC69xf59AsIq9TJ6hXIfJRTFkxfiR4PYbAovcQq8Ss
R2PIGA6f4ep0gwFpfOFvzRiC47PBuW2hetYhtv8Lwg6d5F8FwMbHYpmgsXq7mVLTRqoAY/nBzGbR
4j7G0m2nfi7vpCo3G9/UtgXb9REST+1374HlD/eh1bLICdCpenf3JuvTAFgk8s3KKgaGEcHx4NZC
nW8BJOHZpOuVlgGJ4FeDETbpDo2Im5V8pmihn93Oep4zsDovJjPZkUea7WBeqR5MTiazUpNjKNMN
grp0luNBJqEzi7HWzSQB9bs3COm5wf6Q2xAQDI/0IjbJEAgxK+whQwXQYVOJY2Lkg8lToIrLl87C
AeCPirUImBNjzsOoFSIPtW6RZZod9Bb1ljrw0DMnCddtzQ8VRxD3hXaPVgOKFuZjojA7hgpNFnZG
irSDArLqTfRvNu9pBbiPnYYeHaPpKBaGgW4lVhnZGigw8LJE4+Wt5uGb36LRVYKsnqYzYioG72MK
rS/NvpS3cXk6Xn3u89kXztH8CFtJBo9ULWk+eWGbl7nln9XI7fqMOaoLBFbdaRnNP0dlXiOoTsRA
YrJCM5hkyila0BdA3x07Pod0dtV2xq/Me96EeLI3YCoKoqE/2Gjq9yLmv7OWdVFEnVq9cePxJmDW
02eHyjNVAbyCap7tTKxn/k4+WPp/SNVk1t58HMo2FNJrmKr0cqHRBgIfxtz0KbqSrt7KNZQTN6Qe
6eyDH3cn8aYTHteTsedrXupt2KtPZBgabdenY1ERY0VrGZhvoDAvEVL1TPEt1GkmacDzvxwFoTup
AEPrX/R1AIfmTlmxdV2R7yNb4Pg0zJmR6THKSXb8VbO/uxKk3IEL3F8DVEh+yhdMR1oVtVlYUFcn
XfZ8SWBluSZZwzWRmu3rxiapQKSc4tUVq6l9SoC7Kjajb7R0C9qjXJtstqCLvVjnajkFaLAsVuau
TI72NiWkS4Bs4M6lmkKywuFnwX/jJKWMOQ0HFqFbuWQz9/QXvEjl/50GgScK4Vgn2qZI6vzJ/evk
x+CwG8947UB1aDLIcKATiUefEBIRM1L6rhkSQeInu0/FDXoU4sIXgQN+51+olVwJ3VovDn8t1uiS
S0F1WRTAb/TawUt0jM+bz8WfuysjGnlB6H9qyeQ9Jwby5PfBKhP2auExRmaCRswkf3DDG0wr6XtK
WjrHtexo7ZOWcr5PrSdqMr9PgNiAANpwXgyKeVaC8Ne1FR1vv2M8FUGorEnqWlm19Q1mI7420GuM
neRbzEs4+Oltyame2FwzWuQnceK2trA1gEqSFNI1uOMNht8ORMM6rmSSDnS/IONaTfXVRMb7gUkc
tsR2WmrVJLGTx96US1zdlyFZQCHhPQx7VZJAPDFJc4KlHJ9h6LhrI+oA0Yspt1pEhrig4qR235+x
EMKrkBgVbw5h7FwBObar6vN7X2WVUmhhiLjGpNdmVB9aLwNS/pPfwb7A4UUpLUgPmy6GT0bEv85P
rvwYzwdw+2iKTwlzvxtZgRjA9r/VNChCcKjBG97WZSUul3tjTRcTuXWxpoCSGtcFis6Ww9pWxtrS
BaVnhDB6vL8nDliqlg+RC99KnnlT7yqdIgpSAOjrYwuEBlr6OoIQVTXDCSjQp/XDAAgvcztHrIwz
z0FjOBH2zEdo5MMAtB+T3UwByHooeBOsb0xYBK/38PIjWIK5rDCle79CC+qRSSUr2wdC5QtHwT4t
mX5iPeD3szXpv+3iUEwye28rbvy+wF6KjNdR9hzHOe9WOCV7HB05hStfB/fDwL1S+PojyivQaPgu
9LG5pYo2qexY8dzxK8EPM3nB6io6n+X7EIM9kFprMbq31D2AtcPCvuJ+TvppY6DPsQfl9D23Fmeo
pivtraILFaXX2eWt5tE1L0W8h5ECRU/22kt95OQiZA6Xt9ID/w3UtP1UBGjGl5+mlzprplApxaq4
4eUH1kmgaN7MuPm6QqwP5RShxcKIge3FedLEN9EOu28b1iVldE+XZ+J4tNYH+ZgVClJaa8REQpaL
rcGqtKKLox2RN1rpuACt/2NKZmdtT17I2Opf9Zx31NylBv62BIxIKWZCVZHUxGhnLpH5IGJTpXU9
rDoU5mhAiJ5Ir1P9pQJBnYANRtFpzStMcI0qxfMvrRWzp24sY/9E4OTe7sc6tr0PP0T6xrAoAZps
Fg6Z5cEygdKef4AS5lXteeJFQ5eFzA/2gWUAmsJ5nOXF2p7AYRyJKcAFpLfbQtpfxOiiB1qFf8iW
3irbSra+Gxz936YEbTUciamuqutmM95wljEDI8OvwnXHGzbn6enQoCRPPYS2caRljmAU9sHwCWiH
7pKE8SvVPrbltsVl5FayETr0NNfRdhYF5hU1Ce0Xb9ihl9vFs3433aOHbI0nJTHjQQS78oTbMTco
K0GR5TwWAZCXaAyg8oDtc+9JyJIGrydrwUBmTLcBN63l+HvTuCvpE4FZWlM3LGAQ4x7LRlJBOQtv
7zbZIGxmQFzZyUZ5FwteneHJbwhSP0BuxUoKoyWtFAmn7jhMZRCVDNFts5O+xAHRR+12lKziJMWj
lrrd0bgU/kiUsEAw/UjVqNarFK0IpLfQSwtmewoVX6pWfhiAnL21qhuk2HxW5aJeMl/ngGDfpFil
hCueEsD49k2GfYvErwMyHMDsvGK/sBQ/+2uUEzA1ng9YXhhZoSI+iqBMrtoNOR4NNEDdiPWkSUjO
ooRXKUCuIHb5X3qS2IEZJtOQZ86yZkZmfus9ZKF7u770siU6kubnivptWfHOfQlbdHt3YOxOY409
2Pw+cScMVvVmeEb6JleprZdQoiNrt67EDPCoT3rKyUhPMzohvM3Bfg8rhyq3yaNnKllYjEeJMQ1Y
O/mXfKbOP6vM6O4r2X0Q129HLTyFeW2qgAlAQOMcmvm8CXo3Ot4Cqsi2gsfUZEFx4RU9gJW4W7B5
PVXb+W/SR7suc9o5ddhE4FEHeVLhN3iNwSED/2gPw+YEVkmO7F1TOwVnutayxcVDAoT5m486o5Om
TWQLISWAhWUW4EQ6Gwx846kCgjqASF1n/E18JMotV9EMGPYoQmr1cFffLSdC4eSwq+fCXJ4eSxMH
Xck2uz9ZxtyN6FS7PCIc7jWcFgUV3O23YrGX7hAXufHwlPs1efssVwYImS/ILx8MgWpGVLSuN7ah
7zPOhNcswBqs3zR1Kng/mzYMmqzJWK+DLTW+3ZHAaiM6QZ6er2+hplmId6QXn3LlahXcj9NafGkR
VMXh2Fynwba2+YjUkpehoYzwlsuUvtZhlw6UkF81NmCH9IH/qYHYXMZzpK18fhCZAiSY1VS9S0Qp
TIHmJ+s4IgV8p1yZj1kCkHGqic18srkLZKy4w42kB3F3izz0zsHPeTcnGl+OIDB3altipSZAcIIx
QKJVvwg5OVJILFvysPNkJJBjW8eaMFH255WY0Qj7284ybMkZ5F5ZF1Y7kHYJwmGeEQuo91brEYQp
uu2mfl48bK3HzR30ZTnH1rVZwKS7+8AJVLy/ff/JhppMImotUHnlQ2yfNhmL3VneDoHbr3rVsehh
81KG9GzPwVBNekBUeMSMfv3yl1uhcHjlgTAkxcxD6c1802FLu9sdnkl5x15ySXhcWtviLDlM3iHF
ap8AH+cfC18cXBc3sOMSy02DUV2kflJRFFONYrHSpDGuuiu0aUHK3dxjyFS4k0DeGWBicMzRsSbJ
epG2UuIgTY3SP5ZZJv2aYNcgZKRmIybdj0Cz4isKr4UwAdCM9NHAMXXrwMg0e7vSy22eNNrLyuFm
x6Wks9WRRuu0vntRmvKeL8iU33/DYa3DH4aXdTvf2gPrkOjGk05jBswT984iHQr/rW+3OLS71P3W
4Z/2gwZwKPWZFPDGvnxHKub6FZwz2YbcMJFkDi8YLgubgkD5mRiNsDdbmoKL2TlPqZr3JyfwXH9X
jj0xUt4Jw/3+1ABiC1a2IGVoVyz2JRD3THqUAqWMEJac0BnL3JR1W55xr1k4pd3aufm+GzQ97NXr
edg8WmyNCaQpauwgeEI/xcGLg1e7tB2ItVBBnHacHgZ9ult+uNORiM+qvllTs/LHLQ1mWZr5D42b
mumZP7K33aS2xDrTvLmwZ16oXt72tJ0T+k774yxwnrOzjWjv4mJzPBGuYPyt4xlyE+qN8whc8l2r
XqB+KM2w6VRviiMdLggV3Em5Lbde4GRN8U8TJkYdx1xMa+jB2yfs6LZEiU/XzTZlBa1/RjKG/ZYD
l2vQyxqblcbHWmdumTivlQsrds+aRxd7HKDF/NHJFr+x4ldYLOgPgGGQyKY6leLUj3Se42ChDnXe
fXC880aCn+AOICgwe2cHeOkb0f3M5M7/hjzlBhpEbIVQDPTBzumnPhuTeWvaBuAuoHeuIYmAaLVg
/Tbq4qldxyr9o/zigbgBO2kbMZyS1F6lBgBiyW/SUtWL1bbOxyJq3HmS8yFGRZe+Q2WUzP9v0Cox
HQnNF8ShX737EU9BXaHYjNjBAeM0LsexbIXErlPsx2l3l9y8rj33SqLVl8sHKCaaSCqd9XixBcn2
/6zTedZ/UiegSd4pqNkjQl69vrgGZIpw2g5fnLJpO3LcnO3H8gurl1PrnUM6ubPw7KsKRuhFTzQ3
khgR1foLJ9US2gaoG965Frl7O93MnB2lM0GjufBB7D/Jk5DoBkbPAqJtUrOqwDuRLa0pNz/aJbji
w6y20ix1bi9GybetOArI2DjHIUX5K4h3ASbt8yZcvvd5g+boSFV1QIFt5bvsFqrfq7Eg8Gh+MuCR
jfXI4ABjxFPOKXTPbc24C9j8+P+0/y1o4RhPv1bzS/q8agKpXYNAg/MBexXndynuSXKJIcwqu4Zr
VT3o96QW6D385qI3UI61uHZ3cGQYZoSqLPAifcgCQfXh4Igc8FMb2ore2wyU8cW/zUyPlHzUapA3
dXoP8XAHUJDMH5VA0W1TDYopvQjmyzOviUV/A06bBB5KpQsq2jXNu9AdUQaRtWbPhauFU3TKSbqO
g7auwAyXW8fkOEzmyiddaqePFlJprgMGEtBbL8M3PmgMqy/d8uvOQAYJOVJ9NgZd2xwzepNTMo3Q
AVgPoXWq5ROz8cXnmMlLrHwfkh8/XJoNlPx000NLm7tx8qCjslEauwCmV7Y1F3rw4+Hh3SfvqC4v
TGdS3crlmGSm7+aIo8kY1PWjUpCaEUFCqnnrfprz3REvwYfCf15zgF8aME+yywr+Wfguq/DVWhfk
jWFG10QU4ktVdxnAef+/HlnEXpOQjq/CD684QsyhXRzRx28BGn1NZLzvoMqpUpiyaD8z6IcbeUTa
J1w7Ktvw75m1RLVqcyWtKB4Al4q7UlMKXg0jILJQxYuIuFcJKZEXS8bqaowu7Qi3c2z8C4tPMeT+
l5sAMm24OvQrj2M7UnoJHP5oAvOHOjwkJIIvZSOJi0Ct7f+zeb/iTvMGytG/JTTnjwKg7ST687oe
OESGUOKpjT4RZD8bjJ6HqxQnsueHRtFQtUGSQbZcWU2cVojXaSFzsRPYKI/25KMH/E4bpVb6utZs
5kHbjntOJdCavM0pZH55inlGjxTzC5IlSu6d30QY6Nk9OAT5XgQPx6IiNdZZ0YD77YzZVfvDecPv
kwmrd6wvvL3DFp6ITnwHKRPQdiCXLUnPvrTc+AYIMtD8iyXVXfQTxJ+/U685zeQlkuNuJk+Lu7Vl
Ms88/eAATXSVZjsDfRfydmZ2ZS9q00PgVtIFNUg3LhnLOJcct3iabmrjHA6yxUD2av3XI0xHDZ3s
0HSazB4+mqsr0GqdVq0Y8gCedVOadJPszooPUgvrjsLPQphfCCzsSwSUha21esiK2QG9QhHpuPG7
OvrGNxiP0iKX5O9j7TMw/IoQmoghzun1Q0E/ShjEPvC0K0fu1cFQpJNug9iRmY+HspcFvKObT9uh
R6WVm4SPUbxq8S6ds6qFPJSPCEFobytvzcGE/odcGuYiQv9UhT4PeSoLZWnc2H8dlAh9WTjvYXf6
zlGkgkv9VR+5GSCtHMa6QbHjAfksYIisDvJmgLOIJLd3dRA/gqMpmYCoMqf1bmb2Y0bvaqIgZFGP
het/gP+h1JX0KkcZ6KY54sZGcTWSlDVokPrFvPEqgy3z+au0slDwq+vSs0Biqy6EgQ7alwx5HTBo
HshJMuVuxjBI2pSD5AH49emvl6tbceO4W+bFiTRAOTJVAs8qAGoM9Gz3EpfWe+Chcki8fvBwLMk/
u0EzGQJyf8cJ16rjaliWOsoURlrQMzeDPS7+e81pEAmzUy1ZsKVFcfP+Ov3nXeLL8wiK+Ben+FUj
ABs4fNqT3K2yGO4Z3y6pq4+vwKM+1JnCUtrfHFOY/lEk1PDd4LUGEpf7odvA9XC17PInhjJ/UOK6
9XyZ3C0U9qoEJmkTUhG0jkST8DD4rJFsQE7R0rcafhekgYG5GbEBlMRMpP6TdNL9KqgeTgSO6As5
Vy6/jxeIhYuVHPPjB2FRLWajB9HDDIZ2TxC4TtPTJqbl84+iN+DAzbWNJsetLoLf2K0SVTX+33En
oBiwlTDtbE7FLGz/6tl0/WQu9ruH0/au9XqUv7Ko5Dt3b7gk6qrxBEkNSMI+CmWVZPTBSJJbXWCG
7uSsL+CYFPF2OClRiTm3z5BH9PfT2A+CwkYJzbeJNXPCZ//EL2HPXPUupeKMfaXKjYEGHWiKm4CB
Ha1MjDV3SUNlyJIo8mbEf86NLvFCQrO2BKMTzuFfcSBaCjZY1gkFHsMhQ7kzq1BuH2imoVBSpgbz
kaeNDmzFr12kIzTh1Cwq97ehu1bn8Kulo0UI5+mxFPozTX2b9Q/jBoC8FLockrCy7QTYB7t+Npd6
9llZqozYutFXa2u7c/4WIqO8pVqqVRHuPGJIkVrTH0hD3Ce7e3H+Lz8VIkz+V94iYKrfBV4Jxh5d
mRrHFl+QKRckhrum56r/E2oy9H7d9MwJB2QBx4vd93PMf46gcA1rag9GB6zEXVwFpgT98SHyHOoD
Vm7UjRBRV5XvxoIN3RJVyR6/YGS0BjXPaqe/xuAnUjQuxSmFDj3p3kjp5mHcEImBpX5o/4BunchG
qlorqVQ/Fm9J+mSIMBvCb0Qa9skLTiVzwxCdn7E3lBzY8zkU3rbHcQRDkNSDNqoDpxA0/tWap38X
3AHNIopxkVzienzAPvd4RlECY+tVHdCvbPQ47HKbwZZQ5iPgsbz7Aoc9EO4V9aykghhCdp8vGqDh
R1sGGG5uDw28EtRfZUOvKlR+Ufq+L1sYUAbXhhoRkrElId/LMEune1OQ13EkYMmaoxGDNJZAQQSa
F/iFh9BaOAcZzQ7l5ehAPx957s+oxxwTfxdFBbpIAF/bTm26LAyNrseK3TnvsO6sQLn5ZiyhrbwG
3N72WYRmbPZsVNPdFZlTUihx9RBcL5M9ONaZmtWCPGvAW9e2vQa7Ub785uroA3T3OEJtB+NOzevw
B8SFb28cLeDaWgU9gNCf1z2b04Izu9+29DnFWLeoblDmmYqEb8OdCF8zFRpprCVc9egi/OavFAF6
/fcoHYRu5pfG3fz1r8TYCmUue+ZtUpBmjNcssH7LJA0wP2ki3rjqtILvZ0GkTOaoDY5heolSuc0u
t715mVeuWD7qrmqZ6/29PpszMCa9ZPolaQEmV2qKqt5BStbcup8R7p2vCxl+W9mpfEoQLW7u2hbk
2TAODOmYj/AvM//A8fbASd+b/+NA/Lw3wztGSL8zUff7I44GurfdmBfxfCz3/dNQFZ68De8Jag95
D0WJaXwcf6opjnLocCYHc915DhV0a6A9EzoEfR7w28plDNH5DOGQQ8SX9rP1kpChbRvINSp1GBJe
Uig4aaHWexQvSFcmIUsOAsd5FcP3lrltkwbCjuOJyfLNk4j0a6r3rPUSqcvFYvfFWTQVzDDiaEg1
YUx6gwaQ8mhqF23Z3xq0HqkwciMOJwVKaynuO93g2sBEtLkfCaWrSHUkZDkfXHYwXVWrswNeHOrq
vbUm2puNu3K9BPMkyiDxpjyDIWEJjHMhL7No0e7lhT7aZf7V/Q+w2Xs10FcooCCfDQfhcvkpNmpy
GBrXHdI7PAesYnrB6QefCeLhG1bBYdNKtlJhct53Y4aJu8fJKqFYIGT0y1fJm/Pf9lPlPHIX42eM
RXJYk05MXLZT5V2V2B0IFLmi6cQqLTiOay60EJM6CG/egQGdEk5o4Ylw+roLcdPRbEBS2P+sUjgq
tKLgvz5hfGv5xGih7ISXsw93zFCmmeDBnW8RswINbozSfxWbmrMRjCzfJxaQ/MazuoCdDKEgjTDa
5ddEdfGE0x82aIYqZYbQcpjLAT8nchP7p7ownUMq7hhqliduqZAvZc6j+3ERFMtp3GPLQ96dbiZ2
fVkPmsIVFV+UDm34+xcJiRtyj7L7Yh8S0exRmqO3hYwAzrQ7Fp5YHhz0yLlr+imNPZBbvMtVuMGn
STYz4RzSI4DIbO5UDZZ98JnXCShYJ4FqJOHoiZCiXE3wAoZukdhJliEGm6W5MavsJxJW2JOzV1vb
EkBYrERx0oGEy70LRJmip02JTrzFZ9VQ7xNv2Sc9GP6w3dSJl5Npf4BHlyN0zH0ClpuijYzIOdc2
0nN9QuJ1773aaYhh7oUHGAcfi3m0lxfyqrkewiFYzEVMDQTBrOUDPe+uf769nZrR+yuRpwN/Q3cF
p8HZOXsG9MOLDdNCq6+uBksLhUZ1G8T1ndmTaQ9o9CHmwkkYlQHfhkcTFEnOkPalwmUY4SrL9ZMs
lC5Frl3jSrZv1vKoctL6g4kbnRdks552SF6krRf+Ruioap8DL/Ei1Sepr+CWba5aFR47jWVxkgTW
F93H3gWOvNn2d6k67/3dXjvHNM2zftfjdKp8THnogUruH8tMmwCY9Ocb8RyPc/c9/fMiGGhQDJ/W
eon+X5BW/cEMomh9GGsOqmiaoV90s7CRaE/r90VGrGqi5eEOzJdf76dmNRM9fY8o3vsWg1Vppgfi
wuB86AK2rvzW7Oq5o8PfvtTnNc9sZJe9Xwh1zw345oGUGtgng01x+5i7RZyQWQOUmcQvkc82iq+y
ZKaYoP5zHFY7k6iPdRvMF8ClGFbxe8piJ0TPj1eHITLib8+VGmeFDFj0HzxkQ6GOeh+w9iHId+Sp
H7/I+I8Jma8uTQQ2aw+is3JLXsatgfJ4+mhWAUsH62MlVNk8tplyOvmGi2NzKiEvxYcTjSOJ1wS8
4ElTS2IMmOHhIraEVR/FqgRzJa1P5UbSMqz08eqXM721Ka0xR1sKfxayp5CJNRmY9DAKHN/c9bLF
1UWNDi3FHoGNuOu4YpAx4F2weRN6jqTCN5Sx6UbmkcDO91B0+H9+IUKL5mPDPGL/XnOZT92qwIZ5
GesCkWPaJ9vGij1e4V9T9/cjo+cP7EyzJ9tlk22HUA9TQibiFriRgCdA6K18ihBcYgGvSBVsYOV5
g6eXex5vattYprLqULsxRj7Pttk9oDnJJX/XA1pD53zcQHjrzmtJlLi54K5z1NyZ9pNKgX+dY4sI
vlWXpsUZBLVFezD4649M0iRjHJzAIWSRU2islSAyOc1PfRMP9rI/u52Xn3S+EBsGnSBv++qsGekz
2Ghg9R+NFWg3ZCYHS338IG2Sow/SjHiUy9ODQR+AHY6HalsV21uz20BX/DuDDhDvhTzpgFZPsSIX
TRuZSMgk/fyS1kPWtGI2lNJrFrIhrB/mj1sCMXebtyvZ3XyMmOOtk8KCNiLb2EpWNi6x3CHWQSd2
pHH6EkQCICv1SDY07EoHLl8q0Lppqj6be8keikpQHZ2oOew8xZr1WbYk8LeeO7QSUuRx010wx/t2
Pq9RlhmK1lK48JIl87nSVkrdyZCl1mKbRO90wjsNJu/HC8GyqIWlMeeRNQ5DG5q+xaLM5emR5Q/f
P5nE+7IjbO99zf+IG0dAo3puopZf5M5JsfmWptpvkd8/pL6F73bk2GlWLP1ngYU8/u7vZGDGy3j1
3RJVP71ydi16Rv9fSqQqzSHtEd42amPGeJRZpvMMRs04EEetsIvlptPKwYvEatNGrikuB+NQelq+
aup4WMEYtH0KYWwHr2hynjB0GB0T0qR76gEFpouZHl5QILoRgEvpKtKruHJn8Imjl2x1HVn2tNes
uSxaAsMR2Ujyyknm2qKqeKsDUu3MVC9xntvRxwPXGoc3TnBCwIeV/2YT1ibT4WcMNAJBM6vYZ7dH
SgdlV3hKm54S34FfiaDWt1SQhBxr4zx70lsFK/gycF+JswNLVTtDm550BFnYPkQEjCygIGb1kVoM
UzsoEjk6srnX4XiHuT27X6tAwVhvoAjERrSMGxUSwT4dH3fWDEtQoAg4X3SqgW+GapokeTEX4S5t
lFSFnTcG4h71w5ucCo0OU5qi9Uk9ylsleF4FO6pgUh2+Jv40ocFshFvxdgt+ukuAlSSfjEZNFVgH
DSUndrGMHX8CH09qOuvhFrRY9ktfGrmMHml4vNjlazdBmSIzEJPelGq1crWOwCx2/zGhnLAgzHd+
eO0MjjG96pxI8IELaKtU+u770mMSO9dV0c0aopEoL2nhzzyPuPUQyPr6DzwHThH1xmVaGbatwoGi
EoUuTXKjnOzPwUJvkks0xUZG30Blg+RoTEvuIzj9ycpG2cSgeuun69KYGeN8EiBZjLsjPxHMOpTa
yfHDmg3FQAFz7qjadeDVOUG77onOAjfPRLAZaWKH6Kv3mrOO73IAhnkFGNb09vWgXRuVuKaOzk3V
yNH23sNbk78GKG4ICll9rrib6Wb215SdYqQVYQTQ1v4FxS2geJ9KJ0dTHjXnjag/KlM5EdxlswyM
EBev2PnfSU+XHdju8MUyLyPN38lt/FvPHh0J9vPJHC7K4nMkKAvxsuaPzHMvaA72w+bJzyzjS6YJ
Jr7+6A4Q+uPaADGvom6+oFFYiexmiNdJvoGyq4moLdFhbq1NsWrrOdG0PZw8TDU/HqYCUxO1Y0/d
+y+ZnyW0EBE0iyea6CezNd3M2xEb00N/AGHKN7HscKiG5DbJA5btKRrnKDRPLipRrGL8rBIBRLxd
utER5kV94yyC+ukgD6I0CNjZoA0EYvRnRogQYKIlcqz7sR/Mh/Hu4rZ40KRExmtdrPM3ok+GcjHt
huJIk+PdXpsewzv7EtN/vxz2qmFVNvANmxDfrNNx8pAv0azTgjpkmO0gNsK2h6ZxVE8Vc/uFjtNc
UqaegX0J/SEvNyZTegQYv00YXH0WlGvtKx/sHZINCj1GnQFtLH57x+t2CUsX4xkPI7ov66kJavX2
1K8grQGBlKqUl4WHCd7VpsqPVIEtCQgaiQpQrO94ywalJH8q0IefRWOaZ1gdoMvmOvgWng8EJIRy
5eQoh8vV1YJiedKYnbtFTbo6Eg6CyJ2IfrvMe6Yi0ue8b40j9nD8JW81GSoogzmpapuSqTv5dqC1
o9vG4m/M+FFVm/uYCY7RuTH5d7mfHMLF7/ann2H5tLVZOcziT+0c5z7izlXqSr3/CvMfuiuXqsYx
9C7b8NQ1ToZulPUdUV7Iyog2OH5BN0OsRRU1EwfRcHRrUFm+CsnZ/69mQRdmxkAocLbTD6+/giBQ
GwmNIEVsQtUe5q+rAOE8WWp1AEwUBWFuygb08MDyQp6C4L9uJOlzsUgm4N+L34mReYF9O7akG+4t
fTAeC2sjCP9D/iM5oeP0gfwbxN9CdCefE5IAZks1H9HA6rNiEPGCGHN8mjecICbczEPfrCIEQvnl
rrFJvdnloem6Uq2nVmEapkJIT78hbuL76wr1TDm2e4EHIjLpaO2LFZAZW3yImiPULQbppqrelzfZ
koWhGqY6rvXZkf7Xc0iHvym2HKlVXhVCDGiTekoUfL8cwKQy34riqjmmDKejJV1p5Nl/Mcg2+ACK
yFBGQen31U+D40U8M3Iw30Y/KDPq1C/mYlX2+quvJrp3qlKxbxL+aEEx/CKPYuS/+7id3TdwLDFr
gpnw4ueylf8dSWoxTmjyMzgWSFXMvjYgqIyFnYtOQmG6BRQp9Ukh5zCz/2N0TVpP/LS4AyqW+q8J
R7Bedh8ztSPEv/fi++SRwWrPS9SmH72v8K91kQsK7I+mxgMncpklsSyBWrG5+S3SlFfhqa+hkg8G
mIVvuHgjVWC37xeswAd5H5gOC/h9v/i7kvkXASxZ+1W2uYC3g+BX9p6qxuiMpBrYvKvDNzM+FIoG
n5DhKvAgolEE88X2jzFxyejsq1xTZoiRLQr5rw8dJC1nlmpPDO1rpK5aR0LnjtcmDqjCLGbwOKE0
ZOg0MSDQDP92q7Jfxn1teIJ0YEgKun+mAnvz1ZT0h/JVw/KT/Be+FpHaqVhqUt+bwEbXhyHymKEl
OkbEcWfKMF5G41YtySxMLw17hlpYBbLzFMIkbrCQikNJ90evKArz4luuZJ4apHaKsI8vn/U7WP/j
S0jWN2upg06dBygrSC95GAdNYwutje4dZ380OcjsLUgxOJMOJadsSOlN1mpEqozq24ak/265f/JM
Heewi/ZJnXfLuOYsN8S/Vkg1RUMozV4rMrVV7WFaqeXVHwworWGGj+uFeqE2V/x87Dab9s9pqUhp
/iDiWtYpuDMhCfqUHTucjZsH7LV7Xww20CKnIPeyVkAeVzmQfqWhRoPDYjMySt3kyD7e6nsR3sxn
Qa6AoDuQMQY0xYnHUxtTFAuglU9ye+o4QK6kCMF5wBCuoI8UWqtAbUIIWk1r/Wb9d2vbjeUxY6jE
kOissyOIL7GuLI6KDNPVnhSvsoAohY29qkod/AWdECAF0Zi2LUzPkF6cclvv3UhVoiImQClSPo9r
BNA6Q11Gm4zeTXyHK/6wGm7xhNV4MjXk9KubJ9/Ej+q0GwqlrZSDw/lAnrmwu+2BFegZfsxVn4Pt
naS56idbM6E9no8PCtQXLade6rMqSMl65wtE/g9W5TmdE6rXXcIsIQuHdbA2sKB2W56VvFVJy0fb
s1YKg5X6rfZ9mZaUKrkI9L8BvGhQTt1mkukNxhv1X+bk0tdPdFNmwDZIoquCTsMyL0eIFaUOXtIu
SEhh7YGHep5Zc+O4nyCMyevN5ciyBiIV1IOLpOWu6MXxv3ZA/S0KvueCq0y4OZJi+IUFPIJm3QtM
4dJ7ejQq4eZHpb1UIKx/1w6Av3u/lbCCJiw2UfG/F/+ttmA7rivJpFhWrVQW4gYcHZqGOXtQHAPS
cHz2hbzC5jTVnqm1rjTpOnX2do0UY6UMNg66TuTf+VelHgBgKL9NHwFlMGm7yV48JnpQ4hcNESoc
nSJ12Qvt1a0/GNW2IQfywLXHvlqEyOsJtdXhWUgyxjeMsM2B3YGZKNWZyJSM0f5qgAB4qHEDw6y4
AVIKGpWNqvavyeZ09glLbSPGF3EnJX65ct5pavRkmJwVfjtTNYTUHGQSHnBmTAjSV6z+WqOrIyZy
pmJhi0xP8bsRkkbmyiuw52e4CN1tFYnJ9dFti2FXz6uAYZhkyhukWJ1yGEMpD6Qz1a2HNHfW749w
sr6fgXqvLZKMQ4w1zYZvSaJ21u/7Weyx5fWoTeP2+RDsmwC/kN5adQCsYQnl2cYLrcJP7jw3T9MP
ZwEKqrriVHrTYL5dTpbcBxd/Wr4cEY5FPwkBdD78jXQo3HFyDOdXY4MMMehH49usJgGa9V69fzuJ
S8d8vfVuPdE6JT9cXq3MaUqRW6H4lefWXPex5TSr5HJ3+mY3UIWRFmba+SX9Sh9V+uHJ4yh7YP06
db2EsA2rQ/oTeaGGPaETzP8XKat2sKv7qjQqEit/Ovi+zoCqVt4JbmzKlKKMyRMXuHWogXkUV+Lz
E0jf7eNBtymrhYqDBu/EmCmpKMka3u2l+7zeKkW+3vW8zW2f1Ogt7NK0GhIMwo7M6baD6CzB2Ekh
RvKtXng8MjgQ7OHNNhirpgqZU0UeE26F6OBvKDPFpmtSvq5Msqufi01/fI8J2EMmEeRCjzHLBR35
1HgzVr9/U1sG8HvzSQduuZNXMwtw2RuT19tHK5AEYJ4hDAW7KpwjjnUm/JpcKa9Pxdg0pUnxGRBt
3AHWuUq2rccfIMm+RdukR8EYpaRb+ZUKIaAHoJ9xnODSxJ2ek2HGtRQCYBsQUe95S8M2l7lQOfOt
Cpdc22Tn6RJHRaqJUei5NerL33BekY7TtST63uEEGcbb9KRR/Q2woU7NvYIezuBu0Ex91TsdNQJ7
nwndfiMd6S/ygtDL6f6JqTgK7JuxfsH4i2pKvHGewIrIJntOQh50VbZa/2EYPT0v6IBuq2hl28Jr
5L74gLFBEKSRGHRtoROPC3reEN2QzkxSiAkym7hJmzJ0vwoCokSlsug/TwQA0+m6Kr+WQW7j5C1u
zmf+55o0/ALeIFNTXlIlvfwuGiMcYcEovcEJ/0qrLu1o2zpZ4akveqpwBFuUiyyfKPEv7EfOpGN8
gxmjtkHnJz+cDkITsjlNuFsOyefY7Yc/MWqA5GyHsToxPD3AVtM3lDcz1/Yk1KWdJa0mHuKc76dT
NqNi3lLk52ltJOzT3doymiAkAfarbaHmVwo1w3maH2oKiMajxPG/13qvOJSgFU/rthO2liL/8DDV
j2Cm16Yco1eLMTivgwRB+MspYD5ZEyE70t66n2brt/vpF3dBZTar271yrjdtKe6o0ZkuOxVVDNQd
7K0qr4rbYwS7BNe5M4P7JiDKfkk6D3g2lrx3IfQuN30wk2v/KkXsEGL5cii17ioRM0PShT84OfOB
R53ixQWaInlo56RLzgp6PHidPLp321EyYawLZA4C57wGicUsMNAg1W5qJN0xnKZKh5gx5L5gA/Dm
QdCOolbGWndA8yQBEkfGk88u2G0oHy2OIM21biyE0i22UgqJ15zOH9iVT5BaoJrZQuyUNJyBLFyC
5aQouTp6DkwEkt3fbgT7D9FtQQUnRblQofr/SFzg+sOuwBe18X440f727FvQBVoAU5uTeaTxx3cz
sHs4+R67GC/tud2Gb3ZpmhEVHjdiAXPt8SH174rnTbOpnCexmoXMEhg5iDud8Z8MUBR2wIyaixnl
iAJweRhn9IMUKVgENHb9IE2hQQ71FCIkOPyE+Lv+xCqiAWO65oLWefnniAvh2dZaRbYAN11WlFWr
nI7RsV9m4oWg+yYdB/zhWNG3Fvl1qNj6p65V/9N1iKz/golbfEsVtnh4i9d0ti9OJPUhwFbrfTXY
W7lJUeLVEqEZBxd/e3uaSG6caX8UFOv53YkB1IEiQFW/hNLpXd98xhviXsHyu0Xj/I1CK5PnHtBH
GurxWbtx48qrppJUjfzG8M2Rbz8IcJY3b8uPSrPe0PXjCxGvFX6VI5It1V2HK+FY7eO28MFWC2Uv
e2siGkqj//mAflDsNc0tZa8q4aPkofgj0JxmrGS1q7gKnBCJK9JrdfE3Q5HosKxovyTYNv1hCj7e
FE0xq2dMAlmoxtaPLVkpwC5OC+EtkIAdS3glbTx4xYkM3EShb/4OPmYlfR8s9Q8MaksR5kriYCs8
RTicsen5RVePXXcxXrH9HBx0NHNZUD3uju7Mt+y2U5jECieMzTOfjHftbyhTk2k6rmAXogmRURK0
TK6vpCa+UOrjkaIEXrNGnAlfV5jlSRFG/ZNn2c6A/P8IfmVYaMjXto4VisS35taMddQDt3uQvqVQ
RzfK9WLh47fTu6DUGOJgW5+83Iat0hrqKYNiICWAeEOl1G2iBrEckCsSQs5aEre/TVGlytHJRhl4
ob1ay4XFemg1BpRi65XpjzH6uX7ixZMP0tW9C6lqUIyRuxPV4I78dq8l8sgqnnKVi3wbcj60WFKd
pYnkA1E1+V7d7QWNHLVcSHY7zG61CF7FJ+0dPyvm0QeT6sdolf1svjNntMVmKCK38FV/sZcB3ZZd
lez88/JJ2nqxgiy6toYm3ISiqjyymgFSQUtLS+VwXnt7ASTeMfGhM0dYdxIFp2PbCRvA/x9dktpA
ZFixG4lxXZnD6jdLPyWVL3Zx/8JbbBPlGzO3rpTkxX6he5XzLHyDHxiYYShpzmyWy0rFXFuBNJ5i
3yR4aMWU5IkFHIVyrgK7HbyQdfbXd60qKyjfbDvN9xQS9wsYHdIW1/eLckbgwIBWlLf4qwllLVny
pAFi2JF4BidOiVCpzebY0Kd8IVTcD4unoU3PtAd/8Ho2bct4PEyjmTpXHYHa6m1Gp/e7zMAmzxzI
aYXDUcPmSJ2z6NimgdU5zEzTdBRzFHKADN77Hkt0WjOpbmW2rDDF39E9nkY7vcIGCWr/8nyIRnor
8RueftX2+60eUzaPp3SXgb4Xj8iQEUvi/W/dXgTHtlmf/YqCeBTeZvxZNNS3Ure6nlFOg/RyXTzW
5SDevQMD63C/QI9Sbo6LPS/TQxWdlP41B9hcaw4l5HCGJspUkUUOY4Alb8XmVEtDxUM/iNaPZooV
4MGCYVAlbo1cSbm/Ebfl7kBNTJgs5wN8dw3I92DwWqym4GoJNF9JzxRaio+ZKV3PtHnZN7O9sLti
mHDCjpdfRIq0mEf1KWxSbMjkQ+cN1KVs6jcrIQI9zOMPj8F+g+7XQN/MGQ+A8iiImNzoU9m+ib4E
11z2Tag1WFESC4WBRiuqq82m1k69Vu8jAy6iXndC2pR+sojw5aGcnv27N6rVf/hvDV78oX19+GID
86IbVlY+LdHeHdt/WqSCwIYUweEeUdUDMmsmj/k7cJcvuzJNmiF2eHjg68SzDO1Nw+I6EnNDdLis
wTezSBY58MsDsv5Pljkq69FV/ttDgWiYGFP9ni9MAw28teNqCbqxem82rDxTdth4cYUmt/LmLcAL
6V1RnCydWAFH/nePDLH1nEJGfPJTAv7Y5pLOTd4UhnnwyZNqZ6vBWDKjS/1JdFn4TAOopcpVvppG
wsLwsyg3igq9TY9jUyNHaXGIxsqx+YZHnJyaJwwh79TD8MYYsYeqZYU/w8VPlaqzToMS0rq7ygm/
/JY465loq7UC9FB0BxBc5/qghkcisj6B+DYszO2zozMDRYMVJVf7FTt6fv6hOeNTkox9jXSKD+Ln
SSVvxsipXF9UyJ7rR1AU8u+V8DxfEtt8bi1dGui1G9wCmlv4sK4mZV7yQcyU7h8/b4/Mk4nZVWya
g4QW3l6c7TomwLFrs8U1yRfvLdSnKgk6WZDOVV7cr3azsfYy6S5IG0F21bZe1Oi8hfANWeV11lyL
po9L0n4uT57KEy/rsQ2nh6SU3HY/86UBDVQsz5cjFR/d6vA2hoctJb5g/+I/s4Hw6zdJR4itH5Wx
Z+9KXAqzmy+1cQkIRaXXwx1hY+qozBvC62whdlQWawXWEnZdDNdTIsvxckdEbw4l6P48Mr8NkDLd
oDNPb9i5+zAlETTdMx2jVvvUmGmZVYCcqD8oQJ9IE8cslrRUe6GKlOF+JmQTWH3WB93pmNhaSJ62
YjsTev5geRZEkBaAy1OntsE2zsSLjMrIJLpmQH1YS2XwwlWbGYRM+6iTF5DXiZeIDghThVvyTC09
1NfjFWY2yt+KuCzht13FtrG1ZKlTG94RQ8V0NZpSz9PHH+ihHQPcWxok7H8CXn7UqpMrlSM82F17
At+VyN1bA5o6Zwux6Xk8vy/Pjs/77sh2JtePhcMP0oomJtyvkuHJbDUcjsORjVvQjvzScjy2Ce1F
ui7OT2mbAu/QbKD8bIx+fTts+WnMPfKXNNw+S5ek6F4qfBVLSxg66ll2fJxz2oSEaPebobD733bt
iEJhKL64/NkbA4ATzdW5ObzgbkYyAXe/ngLVp4KlIQySxgy1DZ69+fM7j5HiPNdUwSEJNCRfR8sH
bP0Zq4ExbGPLYDIcLTvSo8EpfJoCPy7DAR2R3auzpAq/ggr8b2OXz6tZz+YOWsJt2yCVFYJzsYmu
6+YXgYgjUPtDqH+6GXm5Xu7E4VrqNSdLoeZp8zy6Ect36McJAjZukg9oo6ARXp06NUtBbvD0VIB/
I8OFmBsbXW2fKjBwM7V6yI9tWrrqKKc0Il26JGqpnlC/nYEebXijyem3LYbQAPcNuuuElyyhMynT
cdYJc6wW1yQ617oh+RI5LCtYV+E6ehB6byd98h3ldESDQc134ehlpLW7xQ4dvga1T+hmG2f1Q0Yw
kIa0bff+80yyczkitlYNiIm30Dnt+GarOBu7Olz5rBve+1F47noFaElq5BuNsQqINU04Jh9tLjtw
EETiH441GnLf+DaOGE7Rce2aKDfeSjbilHwDY1gft6q76eJashHIyIHtW0Z7D+DYrCmXA9pXHNJM
gRzpWhFLrAALx6MRT3SMUqTqto80d6BPrD1Q/Wdy4r5P7ibYUFnZcJiGkTvn+o5+4kbsdAO64rkb
g4dJeJJoHOpS5cYeZyH+BdD7I8VBBqFOZ+oo1eQu67sG84Ffbf2mgo8alpqgX/3vxxiIUaHJ5oti
KvcQlz/9zs6rfspuUwKzbh6s8TPO2/v8jnYWzw+tO68nQ0F1Rlvvi1kGSyidetq8SsQYecRJylIu
ZZ1UflFNwQYLueBZHduw3LuMyCwyzvnQT75sSTLgpGXrZ+UPQHbIxuyGdEQUFMvYRNAQkPSIVIpW
+GiBuAQs99Zrza7LXMOqqoLDYZ5Yu9dxV6WOi9k5kQUF2WI0HUefzHLMbVmfj2p6//Sxnp3v1KUJ
a95v2bzAQ15Ayrb++y4h+tdvk3RtqNO6oE+AOHlcSOw6tTqMIz2uhenTWPjvWmUBNpqBY4d8Tjig
ZFEQKxbXUsNGPKO3yAl81Z0dC/fyRu5FagKtmjrE5Qx3vln4EsU/U4iuNrCzSVdPfyqcLhqUPYZC
F+446Kctru2m7CawHO4SQrN/K7oorvcx6MMexfcDdpxVcOkplUGioM5yY4t8zG2cUg4RhTKi4ea9
+2GHBHWSRTp1p7yy+RsFUEKzXYS6duHGcR5a4a2V7fg0dYUbHU2wYFXctHPkz9rlxI6a9Pqd9KWP
sEqGy/2z2v6Vr9JXl+HyeZF6wFAcu5O/kJONZWgmtPIAl3YsjexpHR7dokZAUiAWXdwH9PFmdB2g
lvXq4dAlMtS3HCm3mfhIIgE+Js+z0Cgeus7TiaoWK4Oc3RyguQP/hty8rWMCI+xsPGJZ9uTNei6K
r2CqqHRPs5WIn9nOZHYbEYB6oWRpFibEyj0dEUz6IVGK7Epyn1fIJw98dsQNM1b55siPmtnenkPZ
M16DzKWDmko632c8x1igbCDaqsv/mgEnpMgIIek+hFpsCRZxvG0vfClaZeSndA9ggoIHA1ztkC1B
2c4p17WzEp495MZcPyvDjetNn7G6H6ehSXTeV4+VDxh6rYhnB42dtveUctG2NV8tInXVqxtL0MsZ
kPtiiSh3xdKMfsah1x9j/MFxTstMfoRln2DVmB5gwxarUNFoKT55qYYueZMHEXbpj2qsiMho/xpt
NO4UN3HTIMUg1UQ89phzCHJyD5SOhneNMiEMAUOUapGXLIVVc7CPRkaVi4bj6YUlmRbJztAbQBG2
cDXQu9W/hL8kWmha3FV/NyezgRG2kv9o3WH6HpNtAit2BSZaa5r8pMEhNZXoiclyvqBn8MpMOTuV
6aKd9iK9tIwwCUrGmIjMrjVv2ZAsKBLf/onB+2eePLyDcPVlx3h+wFYH7helL7ziCY1eWHn0lK9j
Wbtd0dtsUEdUAIhuEkrQRsMVkldORljwX+Kq14l6CUnXUwg5sF957MXOaetKPUnEChmBX3q3uFA3
/L6r0y05Eqwn1AtDIDnxqsJLrj6i8iI6/15WrizKzgUC/lTjqRUgEBuUVfU9UO82lKDNk9x3Cs0J
0jJ9Sr76F1gDKP8y3pn3DUdMrs6H0uY/ZjHSRrhS/IFOkdJ+SdFniCqQX7jWPR5G0Cp29u7h51Qh
x3f6fRjJCWy3wYiHZaHPDCc1F8hDWtadQPSY/RuLriHgXCNEjwim05NVeq8mMgtLchf+r4fRMwom
kzJF3A3BPQ6dHJINYnZhjeKJlEyD7J7HSSP8WsE4Dz8fGcaaZS3/pbH5jdJOn7IXl2YNILxONr35
Vz3Uay54lNdRntGw3oM6G/GD8Ib29d4r+kmqhL8fUWo1R1oiwK7fa60SQyOoyA+1PlbTtUEMTM/0
V/XK05m0mXXjygsb7NZnZROdQBHko+XcCJHRteV1XyPAiXpWjSi1q6Voo44w6p+Cv/xHOInkq7gq
8q9ZKoEy2ViRSbUyjdyMpNpQPQ168c7ZIcq1GEGx+1XUDqVXHPTlMVU7YvIsE/wytz1sYCxAJPfI
g0Ygx3/HqfykCjuAPVGgqyCXo/G5pnfMcL83EU147bYMrZruDC4zMeu3x+w755kZ/yvCvT67Hedp
/ThlKdWmFNc11kjHl7pWVhwha9J/n7Un/dhuSl4AFt04k2CTr6AdS12doo6jVF7pt9CP6gXrD40E
QfOIfsv3LQTN4mhaA+ciC2RFW4SX/RJ0tlrqqMEXaeRahyc0RYRJtizihOovBYyc4eRqggfVfD5H
MHYKtTyPdVl7zJXTefQgFFnYv3zXX9GcwrQcoKBTVEeRQPSCBasd1GiKxccpgCQhZuPfX0Mp9ny3
tqcSDevQ0QfaLXCwysLS8qR1MSBeDtPmm34fCkb0fRKaq5kMlJNvzVXjRNySWL37etN4CNQVv2cu
88CklgogQFB9XrbYCXikzZBEGID1vEa8Dk67NlfFEhq9hA1h2BOIPA+Y05DvWha4EGXP0ptE90jR
+bE3X3MODfMgDtChYqE0E4xBEwgxPvKzt32QBZIaxF7Np/WxbzNzAIcukjPc/sa5lWSiv1gd4lk8
E0Aeb9JWNNCXLoiSDIj+WDm3boNI/wKvmdPeGHSf5K66zHBiC+rdQnJ+PUO0OLDIP44VMwLDKSn7
lGaheMckOMAyYLcBzamOOEYvOpB011crHmVQaAvYhARYcauVhi0ByI2WJsJL7xO/seYJolcrqXtr
CWj4hHCZUUbNQIXNQsHyHw17gA8wwYOe6WrrD2RNrZqm+NmWWsQtFtyIPlyeimhezwoGeWq9N2CH
kMi5ZV0zWHg9KjNG6w5lA2NwmteURo7yh91DZUnXmmbr81j4M17GzbJ4tRVRGpfPpQitvGYuh0Uz
8Y4qu6sYHdDfgxwRxzGSK1HRXZESEN10PoPaNZg7SSaNI709Be2G5PP06Bh/wZNYQd9qT79AZkJZ
s4TqSac+RJ00HJt2gkwbmSN8oI5XZV5A42fppOf8PVnByEjwEhc0GIQ7ZP1pmLFr9hKWOgNod/gK
TaLEKMaFFFK+fi72LvctKRG+5wcVl74JyhzIdSJw/tMtHUwa3chbowEoC0dXQMx8xTO7CiusR23e
IitXQcCCdp26Vn5uBWkgAocQSiWK1ZeHuvqtwDbHUqPIc3bfEClt4B0tV7/NXtYL8e+TuY8pnEtv
wZgXMs/qndhRYCrJvKEmnnxY9W0mtahohkf9+UhEm9tPllqwpE6mnUnhWPzifiRgzTZk9SLnwFSC
q0osDhYevIeio4CuoUjmRT36q7XhgfQqtseJ4YlAhtyv9imBe4RLWjKV8Os/yUChrjpCDOQU4Jxx
KrC7/Y7EqYMxyT+ONJccGWhDVR9Unbr/pIJPhsA0YeH2J8ZIAKMJ8gF5dU9bFKnfyRWC8TUfKW9v
X+yntZoxEIPgYCkq/7gLlKQfXfp5ASjQUPuWYwcM7hIRLE7H9Nm4HPkzFeoEUidxKJ8RtUQPB2U9
PlGyhziHjVjw75VuoVr69JhM+rVLkUNOLmasP5b9w4GPvjX8lkky7hPgBUPOVMRQSuh3+QhzGo2N
6Evo1pqGd9/9Gzp03SfrPqzx18HJqx4dn+ROekI1p/NztKUf8bhDlGROuHVQfb1V3q0YQbpjoYxd
SzGt7OgjS2EtXfR2bQYz6U9pGcnOEuQWa1iuUIfTMzGjhg4ed4PWRX4jCNtAzUyECxaMrcgvw0Ti
DD/Zjz9+bk3TPyYycvP7IwRzZMtyD8uAIi3EwAkhoW6hwfJ5vGiCmg3B1VZoq1Z/Y5w7ENwHx2U+
azjiNs2eUZvFUXbOy+dTp+KSTXDIiuE63PHSjrdmZE5QJbYHlAykScHuKfDrjVSRTiKk7hcCmk4b
MZHlodsBfmqRgNbfZGl1vxUBrnB1fS8XB7Q4KTPk44Vakd8jcpt1AkE8kvBYE4EUoBzIHuokFZWB
7mj0P033Kr9pvKOelaaOq5yIHwNXpWEkBQBCFej4zTUwShjc2u0JNNtQdZFsBp17apCJ+ipZT8gP
FGIGBmeFjX7Os8+5liRo7YXTfWM/aTkIb8aC5/aP+x0ySGw2lcihtjbpVCgqrK7x7OMDcEIi6ntJ
6+U4GpoBvaZF0eCYCPTm8iMRu6mbYpxiL+ewN38KruKk9ZueuEp2F1HVF+SJNnm48RUv/WN4+u3M
dxo3PnZReTpdNU/kDcr2tJkE9MZ3sLgNoRYa8POUR/gCaDiqLRD6e/FWUgVmn51I4A0nLzUIfWcm
GvBl2A8a6LgC8C+Ym/KFIRLONLvxfTq30h9B7ks6dW9RNhblAleF03frYyZqm8NB1gSeUfE2kEjT
e1SvYGzkpPcFpd/tV4zKsIFpuenAWA7ZjMOtB6xUxuK6rp3cYFdjzeOn87Ie4l1lq6M3YUrPre4E
pOX2F5Ekf5locXaAZXW9Q/ZB2t4mW3f3D60MNIyjDLYPmV8WkPcCfSHuGNwrFsdVYv8I0s2i2ZEl
LbA265HSSkHmt2x52JR/OglsRgSOgtiLrXz1+DdfCfkayHozXot7pr6nQm7a4Gob0pRsPRuPBKMf
q3cbr3PUgkbCcww30llngLUGT7dKIBMouzgSR79o4rXHdVvJU+3oJ8dS2pkaOwanffceoRXvkaVK
FnY+9UTq8IMiwU5pNu388q9dKwa0I37+AP6oUTL11n/4TOrhdTheo2EiEUFhSzhVT3qLtQ18iz1U
QcEGE6pxSHRrXGItI7p/c7Z42Ist+7VSunnAlFWQQRzwZ3iW8fxLdpQHWpmRQ/nQwmgf6cJI5xHO
hTEZaFIiOBpOqxNLBie14fG4xO6kc/Up8QCN8ojIv4zpnDwldyQaPvJVDmMXKn5vPkTkWxFAtAF3
XfMVrndj3CJKQ1TlP7m6ZBM1Yli+zGZfP9z3+Q4BvqkUbkwW3he1bon0SYoqoDqwacpy5DRdBbUk
TUvF2B4eu3FXBDCBmQodc4MOSERreeO+WjYDicki60yxYIh5FhubH/LRIXjL/r7yHI7QXgastPRE
sjteIbQIpGr5wcNgg9qOwgqg4pr7j0l5pQPs/n7pRm3xHJOstnaNJPTLD+wdmy3P7MSk7kOr32Mn
MBtNm8IxYPDReAFv/Yttm26+pevsTCnwCIcRNVOiyc0yjTzmxj5baKLIkwotep9ty3ExBFSXLO2p
i2maVSJQSVbCck9hyHAwjkk33wZHhI2+CKQckCduWoG0TubMH45Ba7JaAOwREe44B0L4BgGxUEo3
RuwjeHQdG+TfUewF+YuovqjW3bBkBgtDyOat+TX8YWbQHCaPUHhuElvvlA/C0/yDuqyksNF/QUXc
es5mZ2mnIPAypj/BBNawbU832+Cy6LAteNBa3IfPYvbdF3iQg/KUDnc9byTGGeragHtQT6Fl1qxl
VtTG52wUvBHEWq05WZQWLB67IopCFB2Tu06rB1VRLzXYt59OwUoLkxAH+YWn0cgayVlbj4K1o+c3
e0t7Vo5KYLr1+OFYGWS9X4evd3ETZUk8vhErdgJEcxTzTf/NzOLvbhmWDFUWfa9ZNm2Xckb0Occf
Sjc53A5WH2QiyOBgw1GOasWKR+0oy8cAEJYi81xbRXyl5Ccv7XX0JytvBMCKn9BjK42e/Ikra6E1
GhiML+qcZvOXnv+9Sg0N35zmUFC3GnHVfcLsXNmbgzvW8HZ4fWxTmkK9d1iZesheLWaVwMDmAxAd
1hnNkYQKD1Z4jfjX9bp9+ltYJWVRX7WcVU/mSSUw8d5mivgA/GMINn0Jtqd75ZSCTADrR9dXaYmY
tLwnxNKSKRZXzGiHS9oZS84vTcKISXh1D3BQoePgqFNEgqHMvKI07rHyc14KXzPu7NDLJN6btodd
SLqteWQncvTKrOwXOy7DpGKVBN0yq+Dbb5jO66ObYdRGFUZccZookKbPMA4VKN8dpxg4XXQLml0X
Pywx5UPcbCTuQdOb+2NmT0XBORWo9x8NnsEPpZaAuFRGF4s2g+OvreRxC7sqidNRN2SmpZYlAVoK
clXzEPhqoZq1UsUo4D/W6FLWSn8H1S8ZwicJLJCcmBz3SY7S/MSHyNsuaK/Bq5SKa4wDsr6AYqYe
evWEHirUfthR5JBjsOaLUjRvaW4+w1u2pnp03syuJ+n8swHfADbQrqfNDmH2fhJYrQArjD95IP+o
HxDP4OW63ln0r2hj/bHjUQqSfpIXgPasY4rriGQTzwXujrcv75PrYnOyTrTie2GXhctG8HfLLV9u
avpbsm8UOJhqzMZIpvx5XGO7lNTRHbAJswxIO/y3kBZz75swLBbm+5ysrX/hjETU/3/Hx6fgLqwS
jhTKy6TmblGs3u+Jlj54S0qqRjcPD7XWq7zGSpWO3tBibGIBzVe3g/m1Q0de3yacNEWRugZCzElu
KgEp3rokneVn1xU4eH2QYx7gDxB248RQZNYPIORuz6yfM/1pDECzPSldBrIHi04u+tVj6JIqkfLE
iwlhd0qr2y9d46V05maXmR0nNy3Tk70ZLeKlzuCMeFpvyYrqfbBd+BG7ONfTCi1vhSjzMgvd9X41
SUPT9050TnxI0Oq5dPEN3/WxXMFBYCrX5DCKYFV5f9ZQea40Oj+9r21oscXIc+I3rPK4l+FXjpBp
7jGbi9nuDbg5+SPGX78CgFsVQGOby0SEiuNqfEP65Kf5X/sJgc5EgEwAJOn1MCTdJPhwbPNXir/I
yAEtAIvGYtcRvMz0qTmSnqNXEgfXYx4THOupdMj5p+xy4w3n3BpyaGepr+JHiAj5tMhjiOuGfFeP
hz2GFR/KnvsEuE4GbeuGoQmlGyPLfeWYinMk6MZc3yQvhcrNkZPAGad70pXKCrNY1PcojEVO8EGr
ciyisQETUAHjdVolUkbvyMTpL6eph19PU2Jb3TPFG1sY72cOxvx8/xxFFsXi5CrbPRXbRZN5qSEO
dJgHBw0ZZB0Hba4k3eLaiI9DpgPYk8CpknRXK5/gslXYvhetJJuz6l6jpDGGJikj6DfnoSIG18l2
BQsYFgWKpNX+42Rvzw34LEyIExk+qXuzc6mv/b2fTBIihbypNdNaIgEqKAvF0a6GJOnKLfhsVYdu
FHC6fpggFvmJbJyyc03PEUCPjDK2BnriowSlG4e9IsbUuNhF8jQOitbWLQp6XiHCchT7PUo+irbX
P5r4/cJ9IKQt/G9JLZS9YmjuJflIQPF6y8w+IJyqtaXG6/ycUQs2Bv8Zw7FbANdhOZkfn+451aPv
5RefXJu0GjHFaIETgOKOx+kk3o8hJBA9Xu7nH1tljqrcousvXsNB93LnduQTHJEzuKrqxQuGzRc9
seUms1jU4+E7zPviPB7EW07gBUEdFaCch+y/SoKGIKTuYrhMMD73LwYBGUfgCClszcWkXtdiIokr
AukAcI4zdQX8yClz6CXdEcQZNM3aa1elbbtSnlWREM4CQAOqNcfxhUSoOu3zCYransAkBqhq4Fza
P2uysXtxIqvA6uALqhbEBJPQvW5TK+45V4xO5/FW2bCN2oYpJO9Ti3CEQQWzivHxqF/xr+z3+Jem
wP/v9XCB7DJZOf1H/RSrNG7O8Q7guHyqQfIEXQ7AoKIfP3I8S/IKLGc9JZ4Jz9+rmVXeTAJRzT3s
oQClYhngaIXIWHAFX+sL8+y1rv/0adP6tsoO6N/WWd7qcazVxjgXFSi0EEeggRUFbTcFC3rVOHsl
nBlAmIyF0BkdQIae0zToWlbRtGcmMarOtbjS7f8wcaoE/2yO76OltjTAevCvucXJ/db2TGvTx619
ig9cDa9Oepn8IS+TucQJtFR3YMYkakdaQ35+E1O2nHR+v29kI7cMdKHfX84WxnL2ehG89eZZhIvx
sg8XwYH3fbHo+oq+t8r6Hz64JZdRus+TJxesVMxxi11TcWJqUVrgMvkTZUIu7kI6yMykHWgYearv
0qUsX4YICNoib5cwGxuXVrg1d8HLTRrECh/2iQXLG6LSItDEBOcs7RnJ8YnhFBsongjGuIAv2QrQ
4pl0eOh3GkPK613LRt/u8UDdBm5MXyqS1fMgEilrCkVTnTPdpBgQz1kRblJ2cZJTJuee4m2SewRE
9VCbhX0WafZQrDijWi3prBtIKt5IgOE2rzyUU14KVOEKVv6LyKucfXOSFT/WJByY2DdF0NF0N1Xu
Mvv2E1T2GZxxRTdFb+PQnvSfBRG0RCrsyoQFMtJZUL8M50fXNErlzu51Xofd2ghqeZj3P/u3/dPB
/MwCl+GL5bbYHlxhW1o2vNK7F5bH9TAD+MGXhMFsoqbNgU2Q56WKq9effoVCCyG2IMiSHW70o2nK
/O1mu45CylWT1+l89ek0QzliLDb2f0RlS2ACiz0n2+s0A2EXldMCRWxLIrv59Cjvp5HkwJC08i+K
b/ZJKG5aVaZhSIrSOWIjj/8HrlE3fL37OcZEUheDwcgYhCme2cRGTok/JMKGAxZa7z/Q/m5N8tRj
tO38+iZEyntplt/woiRRSyyK3Qjs/CgK/Il2TJ6lIiNsx18CVV7eXYWHG49bF0zbssh4NxeFIKyz
JwvT3QC6i43hraucQ0UUpIJoENf1FG+VzUhWXeyHSp6FUn9nPWshmdU0KSBcCcRCNh62egkY66SX
t5mP3ffn2wXr5exVD2NiR2EUmbElSRW/QV+tMe5R7VGT6amUqAr2vPUJH1DmESUcemua5hoKJI0v
/T4PJJj8PBP69enWEI2OVbRYNu4SXI81yVFWmPK4a98ZwzVvNIDhoLqSB/Y3egBEM3mEnkqJuq0b
WUubF2c7qwXx7ZgtaqcoB/tGOoxdSCwg+nVBFxMnuf9BYa2NA9O07b8d3ni8fvDyb3XsbyvSkqxF
CScbMjYUcuxXyXTM+fMRiFZRuHylHKxPJOLlTf1A90m6+49C2QcgWQsjq7JxaB1B73RtzBDu4kIA
NBtTRZgv6ViB6PYVGZI1NUd0jQT8ycH6AypyLrTxhdVd3WgI5deLioxHDYBoQjrD2e1eWbVvjxZh
7ylFHmLDwnm6lqCCykfWqvBgKjEo7uE2wPVmDs0rJ/CXsj/NKFDcdDZkp7ooATXryZz+F887p+hS
lp/gZll1gs1UKCFs2GCjhaFNwJUH2+3ULF0IUCxvLEgiA9z9+byDU/YWCF0PyzNJ/kK/UUFlqmUF
urS/UV3AOhFziXg4wkrzXt38E0biyPAVFf4XoaKeCftgyUjD0GuEi/npQmOJ80I9+pfAnEPg9dio
InVsjmORHogZ5R4Zhz+/nQX0Pz6t1P1fx1JpNHObKsP/kMc1uMThpUE7snQZa3Y/cyjA793BHvuP
DRQWe9LYFPXBeuKShdby3braIbQEbF5/CUTgm/OlNOdBsvUjzFXVcdMLYnHSC7NE7wr+BpYPyVct
ZGcJBT6n0tnheBJFXtXPEJlNhquMoFs9lUgLTXK/Jw+rToKCEJqVq1UmA/JU1oqH6pi3dI6DyBwo
+RG8ET2f4OTxRu2OAMhebj2+HSoka9nb5FTSALgszilgJa5Z1qBKcDocMi7n2ZjbEtGvOhoszb3M
2l493q5cXiMIjOUgqMJvwrRSaG6eSu8n9lr6LUT/ySnc/xMDrRunN4K8MBEnNzB7jyNlT1TiufcL
yUQ4d4wZIlBLy+kVd6c3B1fOUY1f3BR47NvpWfHUOagGcRcJEWeKIJnOcFqpT5gggeo25IoOlgDA
ou92XYj5bU8EKlfsZN6jZWMB78yKecWrBEOLU70WfQZMh+YPqWiFKY953zOwxvPNz66PCaOVAsN5
HVGIJdECvU/svoEjpC19LSXEP04w82eZZ1vco9EuhEXBjkD7bw/ZQpp3x7RT80fI1FtxOjsQI7cx
qeUQzcwKY4NaDdyZz57iMA9NQhA4QDsgj6lkRe4bEMlmYYWrZKQ52zqeDWiybM2b81WopqSLp5xF
3F5u2ZAzkSv0JPODlkvKCeQmvQwDi2aGujX25iC7lbJg3lF4TeL4WKDxxGGDjxT+D1Gs0V2/5RCi
h/dS4Hw44WbaBJ7gulX6mLuP6c7cfxzvj6EaVRY74J2pUvzTUnTJOyX2i9C7TcPPhfavm1028hP5
9z04xYmF9G7Ma1SXWEJoa08MZ4IhB4SFdQcyyvQXw1GWo1E25mhi7W6PWHdsabroaH90DoO+e6HZ
trQi/bNUewTOCmbE1fRuPTdPQ7xkm0EsfMHK3jy4fAY5HvkWuPJMujvLIw23kkcwfPiCkIomebjY
0TguZDMZTRsF6uWTJJ77iwHxY+7ciBHr/NVZ3Y9/ZVezT+6xo5PtfZFF9N05o8K83IWp5RXTVxA4
OQM/v5rIsoD+Dkfx58d+EmhnwaPokFofZzkXBnuVkMSZGXf76sAi5S9tfD10qAH8F/3GXu3SJACQ
OmDXloFoBXeRgzIHX8zqmVCNjUTY30rViWVhJMbIE6YQkuDb51j/QLLr6aQrtVdlSSkr7aEJtqDK
z4VTPrSmcvcPSmNV6pZlEI+3I81Vw/HPduXti5gDllm2KP7LqkCzc8n82ro8XmCjKMzAtU53MLWE
VmihCh3gteyUkiRatFLYPWml4SDCD5dNk4dV/gYtECgMaXT8+mCHgKWAc+fay7QfTvssqOMnC75y
OlLuk6DHoHXkegHR3hOjHt/2APEmf/O9kt1LbRPE+Y8TagWkjzjr4j4ld1/XY623wtzvRdoFwpFl
JulmGkN+mVCxSlnJiJm6dK4GajbdxLcRgpQ6CYNYt0R2GS0RmO9UnsL3glZEXtoKqxuMxTaspOqP
24C//K38BHhS36HEXX3w3LXY39cWr49Jutfw/G3E3UEBox7xe5N9GT/UQxzDvFWM+UPeDZ9tt4cM
DAQftGaPRIZwGCVuwxEye3qciSEZ8A4JqSj9j9QPZvoq1kbpsUsUcLe8MpNTGn5xiw3ImmdDXE+Q
76A8eJ37OK4Gydg5I1vaZNz9of2XVFrKoo+cRew1UacL9+mR/e8ouIVRZMk3hhBRlZO/4O9rsO6r
ARjiqPOgnuGBrrmWy1vyuyzO2fZksfYq4Lgc9Ws+dzJL+4A3bR25UTgn03Qh4sdJZvGo0tmN2rkv
wFUv8CsvBZegbqdLCV1CsVIPuX3VA5DesLWmPTkUgz2zjkLqWFbsN0pET+EWqxQ9NdmcPWNwhRGX
UKsT9/nXIpz3TdX82ohDr6CqrQiHqbug8XLZtpGljnCghVMcxJxvry68Iisf5Nf0tbMGo9nf0jMZ
Noou8pOvzAkTUooQYW4QpRXaHSOKU4NxQ2HardOObWWMFV5cBnN54Xy1duuyEMpzhgkTXHq7wU0F
OLyYGL7KFTs3skYjNQSEm8U+/rO2Wn/m+z/7oVD4ErWuyjQ9qBS716APM5XMcXmeQdj35FXKzSK8
SddNsrwvi3JhndQtTNfNjkrlwPiE8IsUA7BLMdWw/I1HQC9HCzivyuGI2mA73igMnh8W6FzpM0oB
mWyDGZ3S0WXHY3W0uVdUDWJyboV6cUobNu2SWa79dMu1DOsP4XB0/FQzKWQxmtYl/qpkoJRJXGjR
IN7M/N/tkUDTN5Wzxh5N1KL9a8ztn2EipzxpszmdYoraXjxv/xhi+/rrUEVWm4t0z0VTQILO6jJ2
RdMhkb+fnLHwzLd4MYgLXhaxYoWXhmR5N1RVYS2k9bO9quxr496Ruj3wxAXD0XI816pj1yDbUumN
lAsFb8N+kymHsyE71sM6wsr0ZGmoxfT1QouRATwpL6pmYb2XAss8JbKqEshxM3LEK1rU2AaZ4HCK
GkCq27EUNMOkGNQjPwu7GMywC4dnpWTnsrz1lmcG/KQ3iO7n1goLLz/YABlZlT9HaiVATGuYQc8V
4RhbQ3APywmc+7eqOpKk/LYRRWa7HTw3vjrrKuUzbRWDXZL/XUkk7kOWqIJHlWcs6jjWaEEVfUqg
b5FPGjz4+FLcJf8CD8U2owamhuQjfzMRqUO5kf/QutIZmu6enPKK+5FMM09tRDwMIzECmE20Gzdu
BggKmjilAIHcpIIxuKZ+UHTWZmAUPefszRd7N8JwuS6l5FCQk3VQmsS98D7f402f5U5dXfAYQNVa
bsrmm3zB2GejqT36if6awA2L72y36OE0K2QXuRelstd8lRTX+mUPjK6nyf1zY1pAXJo9Wd23C026
IFG/h/BgoebxkIybaDNBtgdbAtdVk7hgCz/nXdvXnL5yCF6Ot9pwiCt5giuJTTLXVxMLljjQIX4s
Fw+Rdb6+tL36o4GipB09DYD3lV8ndd2oVvlnGQ0CwtwmcrjZHsP+ZPySuz5icoBFzhLsEDFXK7s2
6k+/UdhBZkSsrTjT+cZOVXMBE7w350grPjnpnUWkCZjAtRPugfShvwmjBNMvonPa/YmQl2znWOPZ
9/nrMXyxOZ/GjRIjPWs8UVnVZ9csCfDGd+6iCkVdByoHSu97P0r2HDmoyZfzb3Q3kGV47xWTSwO1
d5gRt3VADrYVlp1iZgYaZR8EcpvNFJi6e8O//aYROtTsPOZShv6bAVIHSj2Hx/80Bu07lEnFERH+
HGEwcSTChpK6AEXfb8f+mkwihcDTxyikCZVbvT6aAvyVL+MYAp4SHEiT8Ma8YK89V2EnqYTNxwJP
Hki2qzVcaSK7u4W+VddZvE2vwIp3hvHf7eAEg7ziFNEk11067nMC9wOkB1zadmVrkykZ4iPOEVG7
oI4LUtUkcVbCRsOkmsI8hcIB8vXqv+SvqRQLQmKhxvHfanVKf4bd40M5gMBvpwnCENL32ufYA9Oq
2H47tM8LlEZr+4BNi8AuhO28fNE8dQjOvWvzFSm8Tf08bJE8KuyTAdjFZmcNg+pzsSa3f6j5xHGc
nTrEJgTg/FAv3qO8Ou+R+X/Gx1tYWS7NUgFUYbxps8JTsjyuih0vVL7klXRDC25QzF+mCLO4S4Ws
ei0WD17YmP+vxGGgrdUE3T18e53uOPLpyyifAjxVdI6+/ZerAvoTbfDSJrQQ6G1q80TfQ5Pe+WDP
VfcLK9Mg2XRGjKt/3cEXoj9jF8Db9Kp3TlRzwiIIcq1LeUW0CZkjbWldRAS/o0g6IfITTBvFSygP
i6A/47LrW1cYoxSLT69U+Ch73rBxjFuclHSVeRPhgz7m1DUSNhoYGDUcQ0fQpiKkOrl3Gfbipioj
UG6AAjdpOqWWaNCjCO54m8oj3WvlHCryMpqWWEAA2PNO83ouN+uUxiDH/OLljV+P3x3biASVBQyE
QhSzMX+lbkKMtfpsfB3L2w+XaGjGzta+d17r95lt4i2MsNKDBun31UETPpHf1L+vhe+99s9OGa4N
pcFNYGorzn4mwRp56TWF0xzHhRbDGM+EA7IdoyL7cu277NCtUX16ONYJoeBBS0NoLv3kGXeo7IbI
7kuSIkX4uiN3VEekLaNC1K7fjTnUnWZigwfd3Q6SW0dT1E+GLC9oop8Z3y4n2qiKLerJvt/DEger
0v/JEOfc7F8I5Aa+47VSdyxiS7RS1oBPL4OvNJw9x1WQuOEpb3b7tEfND8A97oFsMMkTO3NMvAtI
o/Z9l+wT14N83/aFFGzB4n7TB7AhXIQI9e5CmEKTFz6zWuSV1cGXsCMD0P8hxsN5DEz9y+frG2iV
Rua7ydIQs5piD46fVVyFODTMkFvW4SKc98EgGRYPaMEAMTOg0nx+Xk13dWSGMMzmg2ZOSElDpxIP
aqDIgg9WIB5kDwdrpbscBIbiMONA34Ahc/Zp2Fip8mAmZ9OFX2fKYzwSpmjq/EAUknCrV0kCL7UG
DbqXytx4vmXksuWv/RpVWuOs+zxPjLKvvVBKHys2chWPUNpNiDdQe4btitBv1PnIu7hPF0PPls+B
yLssYdWSt32ddMB7HjNwKkmBUkCq+3t2JYPONpbYO3VoKie2g0OQ9A4NlxZIyqd7MRVsyUFwaR5+
mstWedj1fxgSPEfCPcNDBnrB0iA1fynMw63Sod4pMvHlXfmH6sZnxIS8ux1vHrKwMcL4xmucUxpq
u1k9rDlWnOZCvwlj5zUTIIby9hrT4JvzIpeyh2sCdVgtDZBBEf59VvImmPf5Br9N0ZfIZvikAJTR
Os/bbEq8KeLvknidz3B8spkG29HpSoGBX69nbTDhEw6letLZI4pEKc/PSCalJnNrfrfXiKI+aYds
nE/55hJA2rpwo5DOt7X7GXQIY6F/OcigHPcVHhmBpaT+Y/NWjc51Clqbs+ZYYw1i0NTa6NsAewPq
gfR7w1QZwYkmKLJf5ivV7zHaWd3HEbo079rjUTKRf7r6GsR5b8IqPTnFazkrpJJv/bRFNBz9Gl73
RHb1TyPXE7/OgW5nG0fq1S7O7cjGhXHybYxX6JOrLKoZKl9auNd5cl/NqfeC4jREZLPA0VR+DNW7
t3Y0aUrSoCizUrTVrGbeBwW/cs8fN/bZajfPxkYSmUzqLbb5e2zPt8YxpUMiOfNDf9l5tX5EFkkS
VPoM2z1j9bl9Nr3ZdtSQIY24P9TaYLhmQ2Jp3dRVLjFIHLWA9D0TX92HYeeTc2odhRsXdan/qPdn
sepQodIAXp8w3pzV75P+9Rhh2mAVTVVrDrUlq82UpUS+F+BsWx+d3ExbSAqE7NBNiDiepbvZjWfY
DfdK+T4yZZTWay0jNxzTXzOfzbDhLNfe2e+Z4dBgZcnfCF+PM1na4fpmrEwe3c/SSDgOqAEd+qLi
S6jmWbJ/RvDmKdW+dz7D7NC0xWRWn/IWoY+o8O+LwcLjrx9LuEy4xLRBq0qTyygrclF2pgjVnLLU
XWD8gwOnMN30hZbQgAVuI8ICUroyG+SGgK+KVTECoRacedWK3W+AhPPFTZg+Xftfq7/pxz8Pd1qc
E8NOX1dZyLgPRPqmoPY6TXK0lHz5WY0epfnHzT0n0fw9KhwLl85ThWHJ7qlitdtzh7DeJKSDqNtZ
KTv0G1XtlNWMeOqWpqt90hIk99zyRqRHilaRaUfJypTwauRvKfXx4AEyPtRVQ6jUHXZ04Zyb5QND
mtCsq8c46+cLa6JJOuHbIYr3kZRXkmZqjrTiBLbBt2tUEqZzYZZ4C/UfK6VJNYkzMs3MOHRzmU9P
jRHLSkLo5rvp++B9TIFTFtSVGEw8RRAvtT7f6mkijTSUG1Nc5yU/suBmUuRNYe7xa/Yq8Fo3UO9p
186sYNnc+VbZAjlva2ioD3dCVH1wHxUJptIchUCMqzBxiynwdewW9Xoj+RZLOCauFzzoUuvHzUwr
UvOse04u+roO06VNADDAYBX3I4JN9mK9mnuv4VtD1rDZaU2V7zl77zTAxB5RvuWUGkU4ls+MjKKO
QnMUkYANl9Ii2bwfx1JATmXCRRCIrhB9ql5oiwd9YOHUHryGz5KkMffnpZqUWZw/8qa9OuXUEuBH
SovM3IEoXCIs1Afzjk8h4Fc4MAfn96eb7eVYLwBRp9CJNBTx/oNlksMj3lYwhJ9Yxq1E9eOR77CI
JD7O1WqyjYMbWk6A9xQ5E6klo7k+EndL0fuLsH22HDrUZ0ITvwj/rgGib+FSC7j2a7iO8V8bRz+j
8StzQqQLDPpIeqjVwSBbK9AGxrG2r6gt+fEL7IbKZQtvzsSAZoYnn4CHkCMVtyn9t2EfQkCkjypk
mV6c5eH9nEmZhGnHNjxreNxunZoLP9RCZdF58mo3o2rb4fgjDdMDSoAyJzH9twByNLkHb1ZIR3eu
BA8SMu88xicD8qobG3Y2xI+oAOa12OVDzRi2ii+8IZBE239W9LuP2Abebp/fiWitPlEBRmxgZyI7
m68hH3mqKZj0KXm3AxeIbIgg40PWdg3LYHPQIbK2n+wA91I88cfAMzcvjdW/HCs/jVHoal93cQsS
ztL4TvRdGlqi/NW3XGhxL3Yn5MvhITBoByBa6f24u5b7ysKVYRefMX8OPfbT3lNx8GKvB1PQN1ou
BF0/8IILDJNnVAIZAEHDS3/lNcqMNtMLKdJ1succqqInrfPJWYCGlJRZC3w7vwJaPgn3U0N1A25I
MGXQZoQCbtvuv1W53Vw2r27Owp+OdpK+SlFt0qgAFuN0j+QBKwwZRPUC/paOvjAjNSbQOqggV1y1
AN50nP839NLavSrcn8P8/astS50uA1OlKlE03IbZRfhy8IXEthcx0VLSNEh4xfYszP0D4/VBBimW
K4BoSuy/hH+RbJOwQis/gX76dxUS9NUiDdXE8mfhHTvDOlwOXRTdRV9EwldHpe53SN1GgRpnfWcG
qZLpo1Jfu3UyZaZ/H8U0tpOxvheo18+DmOoOnis2jcr880ehrjaOcZ2qzmGEXwGn8DuFz3LI9WKR
41rJbgaxfL5bYkudoaoIVL/XoCOcPW25ETliRvcoaGWorYb3Wp80PjRlzesje2QfApVpu+PFrRAR
PJHAbRT/F9uwp02E6ZXzXryN7X7wwdcMpFGSrrx6s5vtbP9kG2lNX+ZcRonT2Ig98zTauhIAiPd5
8zLqdJBDDO8HRhhpEDQy8A9KQglSP+uCPWGrQKAnpaFYIGHHQaLXtMktBvExLb/Kwk5sf3PObz4b
MZFyY6khC7ZtmYzvkmbHX8gNYPSp0d7WaN0MmptyYBl0cKJjstN5aFwu/u2lf9OSIUuu02VCdLka
OyV+mJkloz+AEzhAe1zJAnH5OHJmziYwd86n/inwg+68NH6DURu9fDDmXK2EobCi6Z7/xwTsFbYN
xijFBwfLqNlkbK6NUrd0o8rmVSaxeUmV1hNdsMHrqerOe6Pry6HOJnEaeIKMsDG20ha3GFjO7TKy
vUdTXwFp5qkJ39jyCU8RMBKWxGzbKmRQtWwP3kMJgZ+cqsAn0txxmFriYwTx2P5F4FyAARiKNp+d
ln4ibVOv3W0NkKVYWL4ALyJSXxt2o+Ou4gMmz16rOeyryRPodgB7XMNoOCTICQaynoj0zYRsJa9c
wEuKstyu7olR9TzCrQkUJpZRerzN5sz/nOlLAwW+vZanOXwjl/x6cCkIQfdJNpmMRgzskBMQCGXG
B3qEKgldwunAnutVkbUNviqmhC/5rQ0jrfnO3jzD7ZxwPbRdNmZ/v03H3l16FnGf5CJxlYStoTgo
YbtU8akUSEa/R+yeFeZw/Ch91hknxwmH4Cn2jrA0urTaMQ8nx/1MOLln4mZayyMhTh8bicjds7mN
qSWu2vYWy/17Ts5LDSsHMMiJ0bmXq86vxVjmCjAaOmeTEs7DR/Hbbjl6ub/WpHTuanfyLJiP//PG
xgLw5vVExfKxetD+3z9is9WLDGMVUf5fCRq6Co6cMZGFxbMSCT24s3WeB/NvbzTsyiEpgAHUG9y9
v5EODqLW8K5HrHFaAj0Z4O7w5FgVVvCti986Ggv6YzbSnKPNSum7g52NwMgbWvlIPI29iG4jJEof
peNDN5ISYU1coIt3hjh+SOKsFVAN9Ix5P3NFNLxAADKpoMd2GTpBJDs3Jovd856+PDc9CgmmrT6p
TFT813u5Ox9aqlohubwezNSBPBJsJiWTgsXzj8/VV/uTvCd0zNI1gyInNvGhfbwIr2UiYh0yxD8g
vKVFgDhJ+iaMAskNPB0kT/u6lLUWHHZn/bRo0F1uHJbzfYFxczZJHFWOnw/Ebbu6l/05/FKUpm6O
KIVafEgnY4KqDPLr4BGfeBDgwQzRqr6lY1fxpjJV+xf6Co2IhyFd1zkAcKgnGN+U/DG8YQ82yEZ4
V+77X7smA2ouoPzxI7d+DEmxbSa7Sv9kXIGa76n57hklGfeRIeY6T2FYDVJxz57t84qXGhN5aQ4P
3F6TqDppiXvq8sLgsQu08PgrQSCBP8WKnrOBUxwAaKC36S/R7Fu7LbXdl11w87HshGM+EM49/ORg
pr7yaTwZSZrJev954GaFmBCWEx46kvvtuq8bpP1islDg/+Q6hHmqn3cCWFGOcWaQo/tAeHmlVOPh
2AKjegzrVD900FUvoSLIUUsae45xsk8on//tT4N2U2nLffN52WnMUNl52YhluGGNXqsJ72p3XbHF
N3WnPDZCS5Yo29kKiaKG47ih+iXQRUeUZ18kA60GiHnZCUBPPMCdbADivtlDMVc90dGqvQiVSWGy
ydTy1zA2c1pm5bhMPnrOxH/b1NhvjMPGhzsQdhdp4TfX+TCOwzr30Wteh8u3Bm9ejE+0eWW9+cXF
CSx4jj0Dk+MH9lWaBK2dmBJC6GMqMUaxMpr44wGldzolBuMZhn+v5VQ9k14QnSe8rk3SfiSFcBu6
VFL/6Ld5LlBVer10GsNBD4zTAr8kXBySD9hJ3bUFYIsRPQsybQEV7G/a3C4Ii9hDL9mndsVRM+3W
kUL5fOj5a8FUHdphxKG6oaIw9U9Y1t1pN1k3PoWA5/s9nuEBCLUGn4wmdhQg96ACyBQXv9aciCjP
/XjpI3DSfJqk/TNkHGOySiU4xgywEiOEFptL2pQmMuRIb10agnPXnjxO0upVpnqIQ7nt7rZml9WG
YD0Koin+DCKYODNoOnZ+5cYm9YMoeYF4Zker4bhYodsgulf9c1215otEQYsSeyH3z3kFArXDcANi
gp3YDZDv/laAwDv0+xnxaoFC6U3QIDQIe8IovhElclVCMyNhEjsRaE6QBX5pkMHt613IDMTP64LI
pdYmvYsI0GFZYVMJ/rPMFaHUifuAFCvBvGvOamrUZtPfSj6GwfdHttq1JEFoqX9xumYvrVgpVenv
29yY1iWvH2yhXD5RT4tf7sLGH+eyisOUqjPKlFzMFtJbFe3TPFY2GTfGJXn/IkSLzgzFTn3T+SGV
piIWeCopukewLqKgiIa0rX5GBJ8JRKk9ONAQb0c9o/FjB4z5zpg9AwSuAY+yjddqrY5fX8Te1gE8
TYj5lCbTMoiarLEFTYIq//yjBUWzJq4gPVaCLmGBQYykUI+nzRGoE0Fp/AHLE56vvrAAdSBg0HMx
CN6FTEauRsZkiJWpX3vrtYSOhH0XB7bJTdcBARIdG/Q0zzsvG0FCC4hg2MJwUcFlx+XcDooxI/Xn
JihYsAa3Jj5lEp6adLjE6SUW0JHoX7BO03VKm7qsK0HOZnfTkAQbtvBKyfPGebq1VdcvQMlF0ZfS
h40WM5QhlOpTa6ztq4AaAgao62V995cRz/AcqOpATRA3Bg76UwlO7PLLpJg9HeN64HRwEsD7c6Xz
A8xlcry8x/7HiD4tezUmtJ5TG++sy6r21q3aglK74oLqtDsvAsMUyDxfd+rAHxCOMX9/X+/bYuzj
IMKURGMl1PpUGS3k3N85lemlVVFbT60+K3Lleq3Q39uTGUK9tJINGvqMu21PLw8FtmF8LjfStCdx
WjpLajtfUl7vJIRXS0Rz3QgiKhkEXinrfoUoLD2DNOyhIC76iyTlh77VaDfqxcVWwu2NxyZaGacR
h02uOeaSSW3J+gmBSFeuLUhsff/2PY59KxxJI8xmWah3cq+EZRH0EOi+0XBARuDRpIKHJRr1f8RD
SBpog8QAyG3yWVgRvAv3E55870egTGHj7GpKSdcnpnA7Y8tB07lchvnfjGHxDv9zfOtWHr0J7/h6
yKdYw6BYFFU1g3/ucF7aXhbo76dTKFUNvoJc0ANb1JBqZ617oO9Epibt2FAmOD9D68QWXGVHGrzr
2t/0BfMfdQ1U8Ksr77Ie+BXKJw+Y5SbWYRKckNgGsL51E+HDUoUrf+jJcH8FLB0wS4U/A7L4njKO
gY0gf00pxMmhpM+d0RiwZ+ytNCgVr9Ivem5vjbib/UDOTh2jH8DQuoa/irTfVmlbd8SjDxJElfh1
EGzQ3Yenyg8rZnuyl8aAR3BFpwXvenoR8jySN9/AnQtigfBVY7R3tFApDLZ/jvNk2xwgi3hNnwLp
5edXzXw/dze9nYyxBHvsYPWq/pK0el8OK1YMyZ/1hKgFuFmOhnIgnY6q63Zngy+vfyRZOpz3Ve09
aD63Wj+byE5scJW25jjMk68KNo/0/9Gq9F70UovSNoAnHxnM5FkccWTwdTf7lwT5FJikIBQY3usC
96R75ZRC0ww5EkUMBz3N6ZEoQwt19zJTHNqiYYvOFmFWyn0rGOD+uN8GFYsfgHVu0M4/ROXJDkVg
jw3KdT2FK+NcOLEZtAHQV3RYcbiEr0tw7hjgW+XCwe+cr/WHKaFyi6X/NuHYtqItIu67ilGj9KtE
d/4f9k3M5hprqaPoqAwPu25Y6QClcQdmy3s9Ty2rLVXg0cJz8waLX+VZX++5ujrkqAvMiIVwEzNp
t4mjpm/UwQPEVbB2gXcMGr1zdrn9vlW5dMos4g3ehE+GoPDmJXYRMEWVWjfF2+ag3NXt+07Nooue
kHG3WSKxQJuVGNbuTh/U3EnOk9WEeCKXxLfxHIOSkCaush6mICeJRW9lF+iwn7xzY0OkOEDpFv2o
NLt7k8senFaa6nl5eBaLg/qTLnnko/5PmwPzs3qBmElQ6C3VJQNz+gO+lerBo2hgvuz6ngvx3RYj
TllFZdBKbZZiQN4A1pcv1W85vVl8XktYYkCVJoF0i7j0PSMV4ZNDGx9PXqGPHqcWA8bGEcQKxyud
Iv33fSfm2IVU+KBHSrt0i3i9j3ArrMe6kvItS/wfEORpCIRhWvOuuhBbY0mt/M/Am3jDhN4AoNc/
vtgYf7SldB+DlVZUSfWSYbpcpBgztCsWMGhBkQWb2XQ8piYDXYhE+wMh371LDSugYNtT2zZmnFia
/8Kx1qyEjzzlVVG8ee90+zrE1V6uFa8LKDbM0ZYk72brr2EBPqKjvJ3l4v2IOwnBVE+VhlIuVmxL
j2XhvZ7Ls0bqtPOnBRSjNj7cGUP+n/fQTAwtyHQeUa5Mulzn+zNw/YCuMKBoWCOCGITXYxJ5uQkY
b9AFvLThoPRsGLnAGhUh/VAw1A9FWgfwTo8pB8sAaMHx55ROgtRqTNfMtnNCTuRR5EmyeznyN/Ix
5w8D6ubybmKjR5hUcLUMFKaqUmCLfUwUDxK5QETHS6gnB8CMNMe3IspVDk6f2bclMFLK4HDZRcgP
Na1gT6nOvTdwaWBB6ljfjJypysqiG8+i0MKuHdxEtK/CfCeSJB4DS7GGahxHEHv70BV8GgjfiC3K
3acRih2QbrPYQNox1HDoYQpAEtF7XKnFig5EXFUAyASGVKkCz8NEUVU66tGB1Q4oJVGfjFlU/Pj1
tUInF6gTlr9fCaWuLI5liQntfE+aGFaS0VUsu46Hi0C7e1C4lwu+3RWwg9q0yonKz8LqX3P4Lph6
M11HWx2poiHC7VxhnPgEDNLFfunyOlgRu260J/JThySOGjo0B0D/PW+S58H90/lMEMDxDuZSDsPD
SMbPthz82Me8qS8++3d5kd76tPKaLCzAwNDNhZHLVhLtrjrE42115tzD+5fFZL7hksZbBiFkQrq/
mxb0rYyNpDUAhdS+kOJsQL0E0xwyfN+Mf/72oHB9Lq8cfW04dLL3j/AsmHlJLskonvw4CcjnpMei
E9qJyw0cQFQGsqdPrhUNak+m7EUeetmpTk88y3l76fkrrrirlZDyEIqT2n/Bat4KYZ12sfsKMbDH
J45XVOM3nzkZbhQoCR6VNRrnVMxuFXsS4WuN9E6MQzvotbsB1iyq8bKlkjdWJbPTa8995lnBgKxT
qJsVrEtcxY0IzwfImXrHuoHdXGbyAxTVUBC4Vl0O/F9JEHiIXmt+lB//mxhCtdO9TLskjuatBPWc
t3qv8M619Nbz6gO0gtVVyROqv4Zpg/Kn1qX6K7NCvTgcMA32HljhlGVCpD4yaIvtntdXL56d9xS4
cvwBNoqW2rRKLBt8BpO17FfphjTQ8VN6xRpOgojpwUh93jJw6/dgr5VhD1LP2Mfv+RODDQF40Yzj
ZqWlQFLxYPPXBBRBUDvwxbvwCquJXOXI2hi6fdeoWbHrzFmDvAbWdZ3FLKMpMj7/6jR4KBR9qxEt
hQy6P4yMqAFtWr6/pvr0OgmCmeJrBaFxFlDJEvEtSibiLuNrF2cCpqRCy1OzfZy6yKmPQlrd5CfD
BxDp12obo0xh/QQNJFTbsyVt5Lss7RLEG1yppI/rTjdoWOmkYA33ER07e5RDBS1zoo/dOPqXkmWd
E2gAXJcAsVkXI+JWNLt2YL0vLR7nKzR2jihQnG4JPekCVTsrXZCwPjcXfwkC8D92vH9SvR9RXyZn
t2LxuKRcV7r5oxtXVebL0+YCAavWWYnWZh89zg+QUlKoiHkOR9/puM2KeHN75iMlb5tOagTOLTw1
7Ly9RWjqvdtWyUO3AJC3ShiZrJdxt4DLsT0oLbrL12XOW7jvoiWEm9SkDyppQF47ALJS7jBqqgVz
iHU8LjxD7AL8pCIBhlZEUMR8Zm5ZcxTssDbU9p6b86crF2P03d11sX1Suf3giStX7MavbK/fhQ63
dQdlGL2EkgnpZEAx3Hm9FnT3bzzI9XJFlBjNGqNHBjFVwA2fu9el5opDZyH4Im1Aj84qw/XhOzjT
dUcEk7YiEWNFK23TotnevPhlUXQUYMmUR8CgkLJuJpPD1R9wDKYWPUJ+e/W7oQVbkEyrk0aaQWT2
eno7OgOSLO6OuVSoMMWd8ZfOQ2k1Lc21g74EyM/YA0shiUOs/N5IssbEeVU0lply5/P9zF7MMDYt
M1y/IO5sv5uMYlPCqGB7WEyN5zCqdlmG+dwHWaRJxkTyVqlGmlzfiS+z40olH9VuTc5cDnHkq4LA
pLyeYoyKsKFzA3iOEmK6+llPVVRropw91d1ipr2Ey/R1aQQ0mZcXfIjiLEY6FaoOzXGuiiblZa6B
acVtfaUjmex8cMd3o899goqWiTvEA2+KrGo6TFVNDC5HHs7mU6DgcJEWFnvT+frgpKlIbRtJyI9m
RJsctxjCG2NkmWt/VllGE5rJ/Z64IUhm/qhYfTRpD9KIt9dK6d/fmR7rtpfOUpbw6WxqXc59qfer
E4W2gpGiu/xJ9VQSZ38JS8kzLdzoVP6xrYNYI/f7KvRkpR8DZAI+QMtifi9gTmnusW+twI+bprwB
/HQpxeMesa1q6UCvIwtlJoQYRGbpYAzlOCssfGFwfEL+gFRfuEBYlE0CpTVjV92Ob1JR2v0u2lzy
UNDu/KcD8ZGzN/t31DG21y9u+ybTckGmyrd5ok+sj3uJYR/zmENIhPHNwqAMxkVVd3e5qZOJsBoU
uT/3ckMMirlIlRfMxfZWSlKpFENITZ6spslwcejB26eRjAIlJ0xHgZDYZNudOo9Ve2C9POaYlmW1
tQFbvjGcVZ7Aqe7z8eS3di1sy1xhMxMyYg//ISnZRFFRqgvEldmLUlQQEMAunt498ayonceay9fu
VLo3P1p9RKCquMhLrLCQfxDu0aFM2zAGNidmj0ckcZ8gcrPzRtU4rsEnYuYZjoNOK4teL+qpSVK8
pZPKRgvXqEnsykGaXrir6nuHXfClszBl16PKU5oGM1v7PRRdJV7gXe6e5bPoR02vfEIQ19qrqNtr
aDdjmKPN9bXfACpnWQ9Ei+of74zLc3S5Y+MtOQalO4HeZJJFeUY1xUCtHKCTfBzfSMX6/uPaE+lQ
itbbR3CFU1j4RynIlzNwSs2KTXbPQcrrhIJvsBJ6B1f1x++C1clesfnsl87Eiol06oc9fBGC5An6
06noQLOOeezwld4AxIUa7wzv+vhibKqKJLeLA0Df4ey62sa8yGWaWZKSw8R6D5LXgghaUnqODoTs
sXfSEeBjMAuxfeD6/2inUPmYzeyBn36mUa/IYeiPAV2fTFKexnBBi/D53Mht2orY3LEMGpTnka0A
7iKAeoTr9mNWz3BTfH5GWRlYCeSVU//Hxu2zWIgyjex4h/p5siX1aqpWrEah5r9nD7EPrpwdCsqq
WptmJ3GvuQaebkx/lVCTW2d1hpoprIoT+7h5zne+IazfBR1mTOurW7R3geFlL+gSOSPJjhsb0eiZ
sh7PAq7UGbSxF6rZQEeTcYeRjobqDzKpxxetqo5/9jHjayr36ijIeJdQVR67kZzEp6lu3VaLsBwc
nv/jnFeAy6kuf/htvcIGxmrtQxhhCVP3SPR4lXsCW8rQ7cCS4o0LfHtyaXiAqmj8vkPgcktMF31Q
WQ8RfPRstW7JrDEhxryL90HDi6F+xUtjtVoPrZZdKiv7wM5SbfuDZ0jmpDdxqFvXoxVRK3+L1aX2
Co+ZiqC7uIQqTaWRxVaFjqBKD/MAXaI0EkiywXVnLIl2ivJBArHv9sKlnrkKHibRyBC0c7lg3Pcs
RT6FcZycmxq8ynfvkvXuWq4FXSqc4FRGpFSnjXWMq66fQnsmUyaXuTcFdgy9GzbHyNuKF7apnG1+
jpHK+Td2SxjNDQwdkt/YXYy+XojVyyUK7PzWOYaZA1+dsxlxJNXU2V1ef7Ecc1gPNNxqhrtywKZs
yrg2Vno4P5ENgnMrtKXUkiGyXUCRjdZYMjltQVACNUbPgTn2UJeRYr8QEuFMyIDVtqi3X6U9/fr6
C9UTxThNOtxAXTee6L6Zf8FrOuZwU/W9CADX8TYov5QSzaBRf/l5uKqyuA7XmV6XrJpz+m8nAk5y
46PcMz5Q/aq1pMAw+/UNtDd7gW0nXWOV2xubw84w7cacUKl7eb8l7Ij99gJPq3POj9uAgJUb6bdn
hLj/jEJwTs/ox9CWe4dUTsdi0qoOClYv9hHfQlUIlQDus8RKrIrI6BD1qQeYQoEmeQEJ1L78b2ti
1FtC36w3N2eA147TYtgFzlS8ZRgJ9spJz03/jc+KHn7RLfLz6kWEwJiu+iDMrxPHA0AD2DCC1ce6
k4p/cMqX+KsU9dgQvGe4rFDFtVwtzjm9jGLkB0A+AQlOxKjtGKggzagEy6nyptYyLOwRa7E06E4s
KTXnx0sdHRR1DDU3Z8BsPMOfdDp9yImo5T5rOSXzxpEqLyWYMqN1GHUEw4GtYZUOBvhPkiZj/dO9
6dOUyuo6whvRQ6G1xgAbIVa/YlP1bM16PtVHeBIZu5mz8WxzuxhTrjuiyPfI9EzxKtgN26OlyPJg
IE4LPJKEvQU0Id5yq7yFgJcbkptf1fB0v9eqxAugW7jU1/vfB6CLe+ESNrDrKoFbi8cSppI4LMBH
/V8Z3BTPFpS5XUNbeHPZwwGhRioAeOY943miqUpnwHgYd49aKWMNSqtOmjNuUyhSvEjMejW5UEk6
t+cQ6WxyQVCc4ZpfFhtOrAMGnoNsahxLcVZ46Xnfjq6WcxzLSNuXgcuHPNHbiZ4zTSf2630GXgeG
BM2jh+tezHahz2BbcVkSoHk48ui2xQOX81+jFpVsDYeutMej6C9DJF/MhMKDZtvsprO0tHWy6OS9
o1nvy3JfyJHJD1bt/vXAsXjI8x87+K1E0ux+JPhxt2H+BDZbRRfBzGyidryAkdreoMFAn5YNXrys
8QrvHENH7sdRlyIkeJn/i1Cx98nBcsybz8E+QimBvHCNNI6X9eFUTAOopPcUCJuiVpqZNgSblL+3
2+ABk/rI7EVBD+T5BxdxDlI9YEkXGa6//rzsoL0JheCuAWCs2Swymu+6LbyZlNM3t79NnTrV+6TH
NrN6FrUTlMxH0TOUoZ072Lx0SuHcZfZDpWc6B1pyFA9M/BcuVI4X0uvRafXRbCDQUtwCE1r5ruwJ
IBmVOxvco3o1jbBfzv2aTYY/MhwmyBli5xphGItpHEz8dRQqKWM13N97Q880bHVWHkARpOBUolBc
MXXQ3xgzp3LQg/ou4tuY6wNfESYpe4HG7huhsZYqcO6PwQLfxFkfQyPsNAu76GtcUf6YDlFz7Xm8
bCuCEbHSV/Kmqn2vuwFI6hXkF+WB16WCMkEdPuVQxHaYb58eGWBSWehuPh71SUgGA02bon+GPFPQ
ECP/Xq3YrsmwmWCy3D64RV3ZVLmc3PwuXjPR/8cgvwFq0YFJ5XCHZA+5ev8EJj4d6k9SdGTY5lLi
WyLsUrt2svQ50gdGiXCFspC0btKqlMALorRKYkkqJeAXwVP8KmDmRYoe1Hv7cNDLNNWvQUh1MwxD
UOvV6wNU+BUl8MuOfSDXPX9446K4HsuXu6ShsIF2kX9K9XLpJmyzrvjYVKAFV3snvAm3jQjV6S4V
WtL84IyBqix7E4Ko6BAv9+QJP9tyRGvJCKp3Pap0uiRYbbrWc+Rt2/VMKSTAPQnMVkgBhBGrFH42
RVCVtanGdiXuYhBbFVxJ1b89HxbsX4LCG8RdqC/brTsIcsiizAsyt55nMTcKX2X5b9oV4uVjcwQQ
IFp3R/yUK/e8iQ2+Yv+f68gcu7XQXz93VDPgW+AGpCrZkn7RpLwxMs7LMSj+H+Ay5nJlr/iu+uh/
g5sktfIqqTYNHGN21VMtOE42jNQ2X98wT6DGcLI/6tzL24wHM5ppMDpdrmiqhtkIJ8xMsXVvLtBD
qQlfg+ux7xq6pQQpvVLx4yMPE5xHQ+RCCnkCmZq1byfdkrhjFtrVVE+K3Pm6gtVK+cFD//vVCRJd
Cdn0lsuXB+oLHcdk2MGR2UdUrSzMRneXDK79hO1bnjsfBT+iBYtaJCvktMUDoJ/pr/iJUXZ/A4pa
WolRvCA5MXvb6dmp/KOfVE1A3pZ7GrUv0rkgCoz7s/3nd0e6ymgehlTfw4t+v3rbAMpzyCOOu6Zl
VUZXFPPpWOyLA469RcRWKAz8hYnQpNQBuVFCnlNZCc2VK3MCCwDMhV1Po0jyYpV+61pnnPO/KvDm
oCG3MUS0CEPya2+vHr7/mzC5ezqEx6Q/XZaJRGfo9gPv5w5NA5KVpFlOGuuQLMSluadmkDygThVD
ZNoL0Xf5NexEubLyBYWT+g4TvAUALe0CjTL3++ZLT+oPRM5e78ZB0o+lDdk5jDZre5G+W78IJkzo
WqnZiFp7qHaiWd5TKRFlhTmdUv/fYsmRhMpIo1YJ33BaQ4tYB0dIhoVnrL8Sf+du+0lWDuPE+95c
Swmr6AaG4u8xR8gtOV772VkKaEgUB93a4Wp9ASMedViAbCBVWcgSNsy8gfN2svOoa7d9RYCL6qYT
hXJCQmQu8U9n8uMi2lftjhiLnCHplRG3oj4HrC2Nw4AYrTGZwW2mmEmAN6Lp6XJ+ggS2O5YPuszY
5hGpGUY0z3QdoN+KD9Hwr7VGVsAErWgAdE6xicQQMDRjijfamfdoBI9rJ2MqHozFjqmzXGaUwiz+
JC4Z81QRP8H6dbYyMosfHo/pgnNk6bkvjhJcltq8/Zsg/p/iYSbyRwBGnQqWd6Q5zUIQIA3lLvmW
+d6BXAOxj3kVFXKnb5ZvVgMDANMl3uyDuEkE5GsTq8dCGyMX8bkQri5gyjLgWTWUPUov38nCUeJL
1CijEDeGrYlumNdQ6BaknkQs464ztVvrowa+dp8RgOKSNkG1O+w14ah5/VoMR0ThWED7jhzoX9rK
oXaemDLJDJ9OHjKS3PXxsCGjPBOU0wTcPRL10uPaD/YN2MlGe4zpL6gyFDNW8N7ykQsqlOcmRp4A
58g2eCxi8mJ4A5wE/cHMr3VUe1bcqNDLbQnctzLguk7qitLKsxhosbEQU1VTsZbGBgLOaKKzXn8e
kZEVHsqvpt38pybeA6434tnl9ZiX3M5796uSBeWLRfZ+30PfiQe5EjPOGGb5K/f+u8d+TMr2SxTh
iQPAjGjl1MUzU6To/oc9AXuyIGWxg6Ro+B8GKsLj4diyOsS8DAJrUMRFLNBhFfxyAFy4SYYAYr+6
+T1Cr9TiKJ4RkwUQTUyfeXwLARcXW5Zq2fawUptFXDgmTA9l4Vsptcmc+MkYrTCJYXAsPZB3DS95
lMZquqHgjsI1veQQHksRQ/L3PScIVFqrM5ffBMwhd6r407z4ITptYTi24QxdxmEB3ZgJq5QkmVEl
VPWWGUy1rCqGouAvFX/2GCO91HqJqHyQFz8J9Rih2+oHGkkCF//LoP2ROzbfhNchQ/Z0sSaC4tfA
HZK2kQ6nIwuaycu4Zg0vCB3lrm1sX5elmAuaNgqRLoqPdMHTMs4Hi3GqdEBpr6mTI1acOIVe0CPk
ZOGgEWU0JNuncsP1NrQ8hbXYbd39MtZ5cCP8ZA3R8aAO3zOgF6ug6Ox1cxQgQl4OJ54Mp7h7ha85
Z1ZFPiAPXyUj3Qdj8yfG2lEcjkSJ9XSNKdPebV/UrWGggWJZx6kWILX2DjDvS8838PR4PvFEkgt7
nhleXQJXTbiFF6Pu8bE62Yedt0g342huJhADziDY7YvCmiwC22dhNkwkHUQSajK/pJzUpiS042KF
1QSebqhasKIqgym1b2YMpMC9ycAd6wv/MaxB4AIUUkQ7kaOond9cbX2s1UtNO0By6H90nZ25U9Ir
sKudlp5SvMB1QyUTwy7Ngw8RgIqicqpGYjtl0fShevkIMtP8htRLC6O6ht8VuPm+F6fpbmNq03W7
V3yOOdVyM8vrSE49K8PCD4pYl3fbViSIwP0tFdoDRosZs4yupHBfN0a/0z8f5lnHzDXA0+sx8BTC
MTito10/VyUxAgs2YihfaCMlOC1Nf0VhHMWc6eDA9S8l6rAXXiwy6M/BLR+kdKL4W0rCWbpe9GYq
v39iAWWUG9c1uh/SoSL5236uB0QkDyKMuD9Sdyhd3Ic5HjTz8T6FY6ojZul4MS7I4U6XY0x270bt
8AbGhlGf53cGZnUbNa5hgYdGVexr7VlzZ9ogzPA6tNo74n4RFtBODQkaYJJqxj//zRrhKKlFAY8r
QXkw0NnUPzAXcDpxaW6wGLBrjtt5aMld1fEI244joOD6oMCkeOSaCC7LscdnFdxXziVxmZ/RtoCr
4OdzErzudR3/N9SpcQLao2NISI7vQMJteeA7ouCk6Wpdw4qs0+D2kmhQyjInv7Sx57NUFavJPLOI
d9B/WVqeGemw9r7NNJSwbpN2AG7UHR0z8RcEXVrOivzdMH4qi88IKRaomJa0NxXDHCe/4VhoCfPJ
OSaTN2021gCF+Mi7hQ5AaZUwQsSK6oDArMMigStKfKq+KJN8mMcbOzqMbHVDk4DhAHVwVKUSFEK6
NA/qxJlPEhI2MBYQPj9YeHAEbMJLnPc4cmrFYgGMzGUbL+QJ6Xh44in56IKRquuBykaSdIM3kOJq
5BxxcORnlAxrEtNSpFBSQNEl2IXDC++N9AaDupShPT9IR6OB79tRD4qgRT9F4zNtw4h6UtFfTR5v
YH3yDCdnc1D5LPbSG8OHBxNzyGGydNg6Xa/ObbhImWk4hPH0TbdUDfh+2oCiB7/VY/6qfN+/Fxzr
ZByavlx1BBTl5wU9RIhy/p1inrhfmL6MdDza21HWrKmxMVJRuiHozaLktjWncQz4FLzG0ePnapWx
gaQeiXay5vSiA2mxjUfVp5VV6Nv4MWtgJjq7+iC8DfQ+eixabMJa508cdPjSe4YfDf2cfRc4JQ7u
OsL1Dum2R9l8z+bmBdDJ2HYdF82C8j4XisshBoYf8l61yTX+6mFh+AeHOvEFnl9JMMKxeeM965Mx
uZzDfkv1sWWS5S/BXw8D1CpNMe0EZVUtVWVYRv1CHaf+UUpOWMw+VDPQj28h9wM4HWArLw5AibY/
pWwCjtppDaRDu77SkUZ0UowXF42f+TeLeOzkcnXdWfGrKmdFaZDqh7gv5oNJmFOaSnfCQAgF2h3q
Y3yrIQlQORyTUKoZr+L1YDQ/cerAxhVYLtaZXLw7BpKnf1hsGT0GuQp+W86boSZdbnMeYdWgL3yM
9ILJjtOdAN/s9Z2+Z8rM5td8Slr8ofjpwh3AR6FAmG1lobVBFhQF2ZochvzF502L1Hu9rI1/IcRg
a2TLgA5ePydMPIrjScWO3uVEQCn5Ng6FN6Bojhd0qBdRfFZdyjF7KkNGtPH2oUFVwTrFTDovYyay
hmCcuT2t4Xgv9EPndzFcXf4aemwwXl2me3dGnhAyuwuN4zpvurk2RFABBKJdpviFvLkBx5W5ALai
MgOeOGZA9F+0nA9hdpKqPOj1Be9PPmgvL3IeEZ7DYgIT5XbY/fVQzV0ppyDIgg6e26d6LW1avz9k
sMy7rSnTdFmFvd3Hk8SsW2hlyK0p8BbKtYFKz5GsvNUvFQCBUkads5Ald0nRpF4YCx2fK3WvLxx4
NqRWUfmlOdf6vj+jZ2Euj5U2zaI6/3SMEyP6CV8QRjqWkw7chY1s1vrVPiTi3sXCnOAqAfRwsaW2
xYe4kIv63XxqoXgHpM4GDY0MJ+p1XVP+4lt+Eapk8/4mVgwMBP7WuxsdUygoLeaQrkxkfWBVpBU3
bVyDgiJYc4qluU9ZzYVdVHu+KpdpkFYtg0/AKYLR685+6GZZJ7/NF2vZBuQoxk0YB+WYRIinrUZn
oOUj7A3iSbPbvXCwbKwNNPfDow+98P75vL7tmTnNTaEm57FD5YyOMvoj/nDlUKdtrhnJzwc4OM3U
eUw5QwKtt/+IGWFg9cXJEpnzKDKIp2ezGyuuiHpENA849BeQb+nO0aCeXyRP9d4jbGLISzRRqP9/
fhTMsh7LYvTUU8ZKeeuUW3iF5WxNmMHZ6mlKO/gDmeMe+F2eeU6ITqNTQflX48CBBw5c4ne37x3Z
X35UIitifdrtsBB3wfU8Lr7P2fDXx92hXD2tTv6V9FPOLawdprtzxW/5wB+H5Ec7FD4O/jITvDz8
wjrsuLsYQ5DE9V2qcWkY7sCDGqFr9QUdqLPQ7UO1cRE/uMgcKXepgCbbctwzD0NMOcdMYyLTltEh
uCO2IZDCGzemdcz2aS/8QZfe+SvqZQDufegiKqoHiWLOal7XyWIuoolORXcmR7jl+0EIYTGXhA9B
lRrLuagFj1jJOter/3Rih95t/DE/apfIh0zqc4IsmuPh5zqWM8V6aYGBJvHaK0/GL992ohezayud
eefPbnSoMA+crhefOdpak5ttdyr/AijB5nQKbLIJaCDZ6P97GzvrFz48y7ebqtFcXRgrzN1drUW2
6FKCQXIUyOU0zgK/q4elTjFh0MdOK8AH7YR0wRo6bXUqGJ/1zPR1sHV1lffqTiIJzf6u7XgJTGb6
pYzVQWgSDvq7eKOP/VA6k1E+PoN3dPXsVHzijshtykyu2Rw3ZCuKbqFC7CD2IY+jqtdobRgVbblG
PDmfjW+taRjNj8TRzKNX2BejthZ5XoUy4w/SfROy5KPwTATb09f2BqgpSihwbQr1E4D2Ueem0g1p
HNi07xNX1d2jgqKIJoqcBFfNRDTWH0RRVvvmjkshANykq+jwRfe/TG2HENWt2TNQ7sEzDtY7/VVE
7O2mAE5/G7AzXRghSLAipjafrElQKKN+p5UrW0z5pFrbyguOeJ/7Ad5/azmCkaKf8ZA9humwL6OU
uWS+vNb9Qv63QE1bhea98U+Q3QXiLdCtuNS3YJrvJNA1hEraBQibhpsFeGso9RQ59a0RjRBruDbM
2c/Adl1x8kqFxP1VyZrMmk5zqqsNoqUuYObva1t2n8lswCVRubTzPafihQdhAdv9uNpkUe3MjBZ/
suOe96howbBvlZOPTxUyCGmQTalqUKeKxBRK2J7xjqXfxvBIjedU4FSPDk6lT3fpTTwEtLeUObcm
A1R81QPRsjYNQHt1ikVHzRJdh5g/j9tjQpNzYf+rO5SpZZ3friMtZ/ahJzwkRzCsF07mMshxOhFg
0iXZL4BDvsrAZ1Y7qfYa85U3NAe89GT1KswRERpsnfyY0POoAW6+S1ZqIQWCYI0LqB2mPKmHVh1E
+cnYe0X6rMJaTUEHG5f60xxABNjFf+y0F54Ybnn9WHR2cZQDu3N4V9xpZg8HosGuQwUIYvnesBPA
sR5KVNEnQuRjSsRaTDRmZ6tZSaTN9gakzLonOmoD+bKq0RuRyVKN/As2K7AWq8V3AYUMGV5rG8/X
3vqgYpll6XDb2j6GEtVSJKppZwJwsyRTOFaFvpOIyjk+YEUyI1fIHoLr+YaMEZKE/GIDnw5mT64F
D8EemwXdIkEkSYQHw68FVck1SUV+gaUnajEHi1ETjFTM53l66sTUROjs0XucX0Xbdw9+ucj2g0yC
B4mJLRV3V5Pk79N2zu6+UXQvqLTNUB9kQAc4GDsn0ty8XKMigEQ5cG0fruJpT7i+XhyVvDJ+4sFF
I9E5sc5zuq39HUPGvPhUhMjwIGEk6IXPM2fHfdZ/OE1wk2zxxq3QGYpEoCGBlKlX7cLuRQB5eYir
ocZS7x4HCX1Ev+RViI8ZB4zD6/bMxB6ED8e/C/BFjFimTW1ZXLX2nZiBH3oH+sJh34dtgPZCxtLS
BSsQ8d9jQPt7zgV1eagGcJZ3wXBkKLbj5j4cO4V+2h5bYQFj4Xi7vLdT8CuZft22jMSTHUBxr81z
jocBvRLpNHzXiaF0vNFlWoHp9WxY0W2djrODzbKcCL6/pmvRz74FHCt1r2GyScS78+7rOgKn1l1q
5FCEe+asEY9sBUUY+gqfAW/KkCICD92ZCzAdJMRobUueEKc415ns1C2uaJohk5xc9wkQdzuY+TK3
SEJcQpaXH8GjVj0K2UQU6qULyTSbmI126T9lTMoLdseOyp9YjvI9S5jXTXfpbxnUqAQ7TY0Tjbox
7yeXUVVtcxFQC42NUB4lT9qyP2ewyk1jbwbqaABEYG8fCncE3TIb9unneemJMCcRPbwupwRE0BvQ
Ztlo9gBoooNjsktfT3MFJuZVNER8JM3dgfl89YgQwPE5jHxxDSbn0SZATkdWSu6zQjgJsbT9kEtb
RHTV9dqmYenWZKoXB4CNDwcPxXTQnH6wtn1LTEMlNZFabwrXpz2n6OD+rql5cmzDtt42mJbwiI0D
4zbJ6wYrSeC9VnZm7ZhZwyHR41QXgpe/8zyn++xq9Lpkv37hSo/Ko9yUzczNaB1LbROnf2UGjq0f
HzOlGLKq5EQxZ/V40mu98lU35doH7pu/uO1SdF0iJhVCqgt20IMP9XnuMnviLxSTa1LbuTuq5/rj
x20J3jfDaiHCW8c8RI/hWjYldmJESlZYWqEb1AvXLGW4T97InAaxP5HA/m6F6aUy11T9uXBFTdIv
LALuYusMrz9KqcRq/Djz9RVeJd07lTCsPF27Zr0wzysOWPscDb5h4Rf7nTxv3q6iSz9NDXVm/81Y
ZDiLLnfnJ9MnzO5EhlmxC1h9NLDOKoIbSHq36iM+9sONZNN14QOFE05r6LjO+UQ2wx8Mlj1yqgSq
0kMJyFcWxdK13JTuGV+Lv5qjxBTOMOwiJN/uYV06lUJvVZWn8+xA2QAZNMwRJ4r/tbJ0wiBz/nPh
rWn47EFjexBon6aW8UvkYr4pdTGKt99b0t0Qkx6r2yb/smg+XGp5BINT0NqA5RJ8YGTDWNmoVG09
8E+N2dxoVqNLWTK5rDtDi1ZjGly6vEyOHF0QtFvsRgKP68K6EtToCKKg6i8ZOOjFJNHO1PYvKa+f
5gAeoUpxCKdXnQLpw8a6aCS2xJImbJi1101whFr3oMkCNMjbLw8RS3iCdyboCEbj/e1gtW2N7g9v
DY7uM0yrnzGjr0YkHVOxHGDFbLWFqwsZIctBykeeMgJpO3qwczA8yPLPfQbIwq5CZ2jvytQ4KKyM
wqUo7LWs7LuINctyK77HZe0vj3cZLCNsGpU3Y52inOeXdD6jH8TcAmvqvRlEAv12fDU5efwbgC8t
ffUU5mnI9RwnLhErnUSouC2YQnr5H38B7ntRwDYt49O5gvwwulCwTXu6MQpFPIbgMCoCBbDU3Vuh
7oNtyktQMffM6AnavQjlEDqubpWEK0gTQt8QxOes3cBcaqEFAS20UQMxR79w9tDdolTfFvvZMEV7
8+WJl8j8HanptVvZ8kydz6mFxNEq1eAst/F6X0Jo4WYLsYtYCs7cTmVSxngcoT7uHBXhaZBiGjBE
U4cdLrUbtL/gkLwzWoWTE+jBOeM5nYAJPq6ZSE6MkwMLyPvvU1MQD6jnV/0PhJITOjVruH6V4XeI
p4OV42WU7Fq7wp2In4sS/A7prsbjUgc9z5ayekYeYA3xgC/3JDr49kU35wAJpe8jGubKTqYpokot
2uZrN9jtOBbayFrzjIlRR/bksEHZohJtHjTu1bOguaCH0JGxkMpuYwr7jUZvPkfYok9cSscyC8/v
AWPiJSxY8ecyx8OSt8HW3uMWBnHHR4Lks0Mic4aCY6T+ne8ltreV5yuD/toy+JVbQYJr1JzfIzhh
vwvJtig3YbdFrVMlYrsdawbksiHdEYpFPPI2SJiRS738CPuEhHRT9AVf3DUvds7e+7mD9ZiDaXaG
UBfh/bjk2s7sKIM0yzH8kTjGOcNeGXTZ4PN3wpmamaGU5/kf1+YQR07p4EXnGEouq8T0Fq7Qjg6p
0FffF2xyoq4ysvARkDKt8NdXcdAxN7Hrh9BSZequr6bNAdQ95IB0lCGrV5KMkXOwx5D+JC0P8a/G
3RiqFiPhpbPILA8Hf5PJbPvQxZYQg3/Q7I7yU7ioHMr371bSvR9isDZIJbaKkmAPr0LU0yCtd2nd
ecYi8eWsm1UAmM+WsCvcWGmntGcEpHez5o3Y3aDW/8JQTSE4zHWRtrH//xp+R0fMjZ4Yb9IHe9cT
z9kb3O6XY5NGOraFtzZUXJVLiAzj3pYt5b8zlB2ZME+UlusQWm8Bzo/JJdhZ3vv/5TD/hAGrodP4
ZqYSdmS+BtONAnsHYkR9yZJgQtXNPxX644k4QeCHvbVPUFUigwwkkwZpZEzLWJxbMssKLkC1NY3J
eOfkpfCRHrM+jIJe4187Wm5ZFpPSQqhd1pCTK5nH9VpW1+yC1Lniv01EO3QRUZZdkr86t7YamlV0
Dk7DQXzZ90Pp9+HBo88+q7yHeAXmrcNGS41Ax4B0i14kE9X13JBSgIdsDnxDjr4v5uZhoBXvUCld
cI/yVjfLdIKlgSu1Vn+vTkq7sQ55S4P7ZGW+ADhEoNtbzphgVG5fmOLuFhKsFTJYndDW/TZzwB8A
9HrLNDdQvwA7lOCh/5z65UJh3lL9XCSxOt8LlgwVyDzu/yl5CZruhI6ysiBGcodYHagsQRb18sg7
jABQx5V1qq68cBGXMu4S9sd2tLcuhIkBKy9FKPEAkPNY1zpqwvhmr+ZRho/Mm135AHRaKi8/q1IS
tl9jt9lOYGc9AJjYSTPEHbzCdFrQfr7iRHDi3r2cMrw1yhkWl7FPftGeW8EZ42Wmw2wczzYf/FUr
v4OmDNpWgz2AqGxn6KPhJCFJEwYCB6lTOtBg/S7wWtIYavG34w8xaKBjQh4K5OFU7WSJXXvRIQ8W
XC2nRJFJ9qzLotAPSBfcXZdMqbXF6AypzYXEr2mzLZWe+5GCKJdZlepc4eT2bSiXBFyFCkvb1ekp
xdx2uKPdIvVl/D9H0JZIAOFvVRZwXYaa/NurNOmiAWw6oK5dB+4/fAnSreGv5WBNk2SC+/pjTDvV
Wcu2aQBpGsSf5vneoDX+A0dkr3nUAPHQyxLYxFBlq4R9fWKqNj41bsvqCNtm2LHFh7ooOEPqUU/x
7HewQ9v2KwwZDAijgxMYH50EPslbgCT/MP9hIi2z2mn7q06w8Plzs/4341BMCSsYLOPSYlKqOeBn
VjyUdIvxOyhJZ5VjU+EW3DetuYAPRgIHRIF5vlmGZGwL9kp/g0bC1w2I65EXYc0gUk3HyhGCF/IM
EyLnyAviDiMrmadk81dmD4r7uHywk8phcVxRJ0m9zfBZqlhaWUAL9n/yV8zlIN+fUE12YbJXqttk
x+GSYdbVTEbJB08L73drKlp8y+daoPqXzd2kvPZZWgxyInd6Zv/RXstDFKSAmt0cIWvqiHuur6MY
jEa0Nt59SnT3nlsy0Y3y/wVT4jttrQ2yre30FrweT6h57xRrFfPhhb98fLYMyF8GjI0cAdLh31KY
qok2ITu16zTZtTq96yXi33JZzXUsVH4n6quUb+jlg0yAeNCxSJjDPCxuroYEDej8hUVrDGklTsM8
Tk1hDQp5GjTtbD3aAsWC2RfsyF7lMgJlUvIXMmeoXQTB1Bm7c4qIf8At4aSz2MrsNdetLPQYuod7
qU5vOKM+Ojor47MjOkO/M7+beuIQEdBHCLpglb7TH0LufQB5uV3Fl5pdtTzg6BghtwBYBlT4yFQY
Phs0jxCN8k50qSiDPtSqQlg9Yc49n0Wx2npe7xdAvSJvROWokRBUMnyxXDFDsy4csJNTrBoQdG0H
Snd77ZhtXAC83btY/jzE+tJ3a1H3d8BTl2B7tUC3KFawn/f5pVU5qrrUoN/vD4svF1dqrXV+4oYA
FEGiK31wVQXmUfPK9+gJQsL5aJkp4tkwdfistlRINVZ2OtW7cubBEd5om+KlooHKZpBaB7KHVuJr
wjdYCmi5/eebYk3VHotA8dF3aOhz1/gWdts7GE5swG6fHtF+54wugnEGgwTwp0MuEkaMyP8B9cfl
ASWAHFcC2qWNgmesoYDIns0DmFVCOL0LDtwpKGTRIWvFWirHS9x4lu0klUflkhTYRUeL9ju17J6k
EzcQQyYJwgRO14g/69A8j5eGvWmYp+8NDivcmQmn6QMUZRAUNThnWeR+f8grvpizaBInca6ywIm2
yhDpiUWy7ST2cVIzaNp/+u6qBbbAZw4pubEzWUjlN6+Lo0go48JUT7IsOSWn0u/gJLbV4I+C5tid
242/7GrWF1Rdgq7hXWmbmIpJDEVh+YRivUS5Q033x1+5htmgSP/nvrknGR5rtNRRaaYyD5OBqZsa
JR5csXPgDrwtYtdwbh/XopZeelBFPYbo5Kw7NbGMqtxmEpNH7apd3SWlWdJl1eKjjd5k7vFw4p+K
LL5gS0bzpL07hCmLqiwMjVFciWWj/UpuuqWgvQoMSFBBNWFP2JMDgrrljtLYxj+mf+qC8Hhym6IV
YHbotvaa5yWoKsgHnct6DpWnqV8oAuIEs51qZ1sWWyHOx7zOpFRVSiV0L21bPGzJTqkb9A18an0U
vvMYB+FDoeWqBG1RYpfGRxj/ftflp5dxJK96r5iy+gTw5VE+gSZ7Xp6Zylf3drQ9nryXZlbuJJmi
/WguThaFpRQw7IwZbPnBqpjVVb2f5YZon+NVzGGIG7rF3f4eij7O5tywLlKCzOjZ1/P7hS0Om3n3
YOpF6frR43jEXBaqgM2yVzO+pmxZE5Ode8wX6K4SSIfzNgPWzczlm17iJDQrVWbkWkKnmBRB7tOR
AyNZuA8A/2HU3EHvY+8i2W+rJsVCgowUuanUQTzKIMFvpsU2Na2kz4eumIztsgeKINq6uIhf+KHb
UIKDn65jab5+V8AuXKeYW4FhxzN/ECzX5JJEK1iglWmnn+ZsWGFwN9zVLcqrgy4BOJE1gsEw+qDb
GC4cA9bztEG59iIiMmNraQzuyzbbbtDhRviNh0XYxruCGpB7cLoZC6hRkjKRGtmOLq6l8DA1bLhk
l3iPGXcu8t5GNqPrqg4b+T9K5QyJTHEAvvwc5yl4sKJfvFnbEuxy4RDOeVBGsGL+3GElglEWGbRo
nnoOGcSZFcZDVhq008wppTMlI0xsLJ1w4Q0Y/xd8mUS6kKsz8zZpxzl1/9aZpuy3hOmlesBRY6Ai
6TwD5LYqIry7tiJAMBQkRSDChADs1hcPzDogXCtXckkNsrGDCS0pneWPZL9fGVO1Vqz4zck+jnO6
hZJaRwyb2SdzapJvJTmNHCiaZ4eA+1j/FmtbrXr9dVWUoVzDRXhuphOKzaZCPZX0ywgLsrL0R1Ps
Ze19RMiojov7t3t+PEMpEZ/H83n5aVi5vs4EkorFtXW6h9xsc/kBTDK6rNtDbQaSoikuD/N+JRYZ
0929/IOYf/qEk+uNtLX2Qzd21GOux/XngXLqXQ9xfsAdWmthCMmzQgn2G2N3GZkjG5M8eSkqBQdV
QL1R+6BP6Dpo/8ALsp1CTCJDY+L7FqVlT144E82E28Dg5bnij5QykII6nCRJerhHMQ3iZpRJ2Eb4
4pkNZNY51x3CKcIkmnJSJGU/r1HD9HONKAfdVgKf2wmzj8+geP8T8givaCwluFeW0c6jDaWtDkpp
Dw/UGPV0jrDuDChSEFD2BxYGiHcLoTR3/iqjM9KSceOf4dFyKT4bRutKXVycqOp3qnWMBcskxxph
Tg2vkHujCLDwr7GtqpVxq80Pm6PVSCaYbYIlZKCBeuKTS3jHXLU8rVhbtlENJPHREcj4yC6mSetJ
+6zU5hqlrDy3xrx7A6fFwgiTeWPLNOqAd7D/ljKWMMS/MrPaXA7XCTS5Mw0PXyyi3TRECCwVO88r
QP2bF0lQ6Wcnf+NdG9z0Xr3koDyadSjo6Pc/Q16DT0JhgVOKhqz/mKpiaJAJQlU6MD7xB4Jrh0lv
F5BMYVqFd1iA0+WhVC83fPl9NzSqGxFbPoMqiKP4X6bwTp6GIlPEzpnOIoI8I7XE8r0Ik9xRwr82
uglST+58dYd/9latscfkx/LDWjpa97WxAxckDTcS86yPAPglLAsrgK67ewgQps6cw9THiEx3wA2H
d6Xd70Yu0lME39J2atTmB7oQXKa7bmsloLYrw98suKbawmv50jwT9enxZbikaHcM19W+ksuYKpZ+
kWQfBDQLWyUUl1DoyVYlUSzoSsFz0QVCFG9SixpY7PakOy9G+VieMkQTk+NUMtGJ9XTrV5+SdrUn
KyWjfW359k5w9lDksZRBIs5cXJXzclCcPDM30kmdYuk0L1Rogrez8F6RFatbNUH+9pv4xK8gDNqp
yHl6boI6j7qrQX3KBCptottWcnld1dGB1BKBhiHSoHP3XVwQEacpeKpikq/9Ou6HIu9ya39h/pzL
bRMVBeTwIz6+EDyR+Z7MyAx/6Gh56wegiYknGUEEJZsnzHmqvOn3jpvJ3yCnPSL0jCHOqvEFg/6x
zD9Kj/qBcvM2+FFg65cMVZAf28Uk61BQlbPzM5Gj5LFbPRQ9wUKcoCk88PU5X4nz0pzLbQqp/u20
FQwdFp8yfe4gGC3hZoY6BZQVi7Fpg6NGAfpaFf5iO8pNd0gApaTj69tZ7avUOkd0hnKUDPu/FTAQ
sewYdUz6FSH3jp9dWLBOdJQatUcfwc3I3Se1OaKQvQ6Dc+1/GXHMaIcXQwgy+Un1NND505BRnfIL
MUGu9W0UGJ67Sasd6ppypOkWvSZ7BxR/Y1Q9X+25m8HBrOPGAXiJ7nrpW5dkmlKG5s987qKNmU98
B7T/VwHrQo5lvsliMlyy++j+kJy+QXqJDPq7d7gYnabJapCxEf4lixaTiU4cUQp5EYzdtTKwm8Op
v9Brcg4irRi14vcVgANbC+GFSPV8PUbDNUkQjsBE8/1x3lSitsbf/EmrANRptJFLZtmm5jHNl+/A
Xq7UXOnbc5AmWY7gWsovn9MWzZ9dFkW9PuCqo/UO56vYF/1Ht38EO4hrdypgPYG84v8E4mO7xpMb
gMPdEzW8WodDfu3oaV9avJyM8CIexLm1hVQ1AHzYl5SUJ5LNTrYQG1TzEinc4L1JTbZY3Jp6pAOL
d5YZvweN+RWDfGL8un58jmTlSmVAuE5pdOmAhNHMfGpcYvAuQzlr2EpOf7MX9q/ThoERH1QlyJua
nxV/iOOMJ8xpjk8v+SJKsEhm+aslP6Myx5nj2Y5nyUK+S+99NRN7L+eNQ44MKQcoDZvBIviBKC+5
TfWgdWAh/0DK+SfsWVpciT1AWI3p9S8D1k1o5rXo9vK1sfX5uezBKK1srXf+u63JJ1W26D6W4v1K
6T36dRUE/GZ56MWHtWMLWd+wQ78GMuRx6PlVmvPzB9v/YEs4uWuQaFbTeZdHMwkwv6mWPFzSBH/V
+br3nHKMjJ5jZPe+Ys/kSweasRsSnwbmemTxF/QmUQfJMIM6fLLUFvzxIvXpKeKAadBNWaw5TaKm
i3X8wZ3gJNL9sLX+/2yZd6alynpFa4ZiAHJbEccyId5W/rgrvL+pt7D4x+sK2pizolijHB7Ic+L/
XDE9ePNmpViK/3/FZ4uKz5W5M/kxlDEi3dNsTQYHm1FjexYKOSYKz6F1b6qBkQNCa4e6eHJid2O0
Opcq98b7a/1syez6+PwNmKudGUjXpYSn6Xabh7Nyn76C3dz1UYK65ZX+RWps5ed7PbsiUHuqwuzr
TyzD89AIJTopPBP15LRS/Oq8o/hrRYyfg4my7HMnNDPd3zeWmbQv5ORJQ1245KLIQvC5FKaWWDVs
7zVnJJQo/SWTL7QUp7XdgZQQP8aPbgLuOUU4ZmGhVT/pEOoOuqgb4njgYDtV6N5/EiP207cEVlY5
N+L1csLesrc1EOowNCWwMg1nGJSPDyI+DXTqp3Wt0X0bV9n1ZTokPm2cdNQjfe0mc4U5RhQXq4r8
4MAt2iJf/EtCSBRx2lHV4gV2M4PTHPWjWCfOZhN48QA7C0NjiirX1CkydFlzq6y/jJ4PivwugdHp
ICQlS2pDrNdF5dc7IOUVjEyvzcKdxO/bQIHFUaFLX/URdYagEZZ9gpZzuM5z5muceHKCmD9CBL3h
1rTzuMeTss8CUAxZjL91UHAU81wsrhdJeWgx4HRj6dckwsgP+ytzDhtZ0rHPyNZ4SQOIeU8TwGiW
l3y7PagAfk1yYrJyA1m0cEYDGnMq0iGx3mggzOfbIWFAog70aNP2VU/5V9XrYvjDq0dBfWhGdq9G
riMzB9wex1gplYvIJMRwO8nCMev0GRoTWNSszq0V1lJsouy/bf4FYk/o0NqOjsR5CH7hyV/d4VHH
MCx+ySYOafTv1Fmk5tG4alyxO6MG21l+r/2NucHgP0SqFwUmE65M7TX/O83z0BWYXlX6NC8ca0LW
HDVFpunLftVoydnBERRei2Lbh55nKavYh3JXV1agPsZuKAA8mJTgY1tOulDYHUPjkoFpuprZIZXF
PpMV0pSm9GHawyBmKVIOjx095HJ58eVAXUmt7d/E8nHK95RORnGGbFSXF7fbEpJiQ+GlNJ2pbmTx
gq62KKK5YEjuxv/oXRj4bsaINBSEvgelR4aSidoYtTRGJ2w5awbVjpVNPP6wwpnLNn00TdUsggod
vxqs4ENqrCA7nJoXXmJnrjVv4V8veXhj9JPySmEXoFbYKVi9UNn3lLT1gjEguJOodP2/4J8+AFJB
TtOqEWjxTmRTaODjqwPSsWPJBKzatndtbLbwhhGIr2fLZgqX4dvM217wKvm5tVMkPShpxAabfqd/
uzz2Fd1nU8V4kYKTkrdOB21MsQIpPf7TKt6yDpyXW/i2j6yRvWNXREly2qLxV98cxVWhYeC4p2NF
9iIN8VarUheHm5jlJ2maLz73Wj52ZV9EyRkfy40rmwD3QXnjdhtDskPWqoPKpFwyYW9tsUqDuIb1
E+jV8/t++l0/T2mJ3AQjcymVRGOEk8P7tVj0kX4HgpHhHZsALfFdFqXffYhjT6QLJAjrO+IsNoTP
Y4MltjeIFWNVW9R9Ax/jhe2BtrUcPJfjUFLHtWMU9pBCq6coeNq7Q1oAoey6RhyB/QSP02wFt4hY
nLx7OXJTxV4GpbNXgbRgDQhjK7rZYwFo6ptiSL/+ggnZlnKhygpXR4NVb1tyYRNZ8toIEhJZmrlv
g5ncLZRR4L649RVrDwc48N52ZIJB+wDGc2LA4NYJvvvC5C5R5tVLw9SCKVOi4AXZTgTOd0oaul1l
TUaFMU3nDxZOHHPyafFQ2L+RXAZnhsCd7QzOWtMAUXpXHo2CL1/Ob8N9pIN/a0/Y/DhhrtHP0eEk
NtE7BxyG1/IgsTA5nc1F1mWk8GOo+y7hAYl6geCkqqxRjCSz1H60BJjtkN1RIYBL7UYdaViiFOU2
mIBr43ZeRqu1T2DeA6dLaoxade4hfeml3l8UURFf/Lx/UqIzlJYYXnCFULEFEcM2mLMN+Fa55Ayf
r790szZMBJbPqUUPG1IMeILJ/fMPanw65/cUeEzun/TvEhcssFgafoVtQyjh0BILNjQ3p8SrLC/Y
vqBS1MV0K7f/omLR9Wl1WGn8sroAZ41K6igvWPuzNKPsRui62QVC4pKjTJY6YMZDa8Br1KgSBL25
aC+mjIUKJRpuHlKI2Tls0Uqsre4F9LXThx/U8mnd3AXaUb7ZpfuO5HRwQ/K3Og453RZRMGySIcd6
92qpOc0PcLbfvGiEUObVBwYZjU115Uxni0vKupXSZh3S0Bvtb7rCeJmHKavjlDTkG/5UFiAM/4PK
e6K/P2zWtMRQxaMPX2TVMpejMuhMUzjGhy6jIbpNMgNxjnt4W81diOdixZ2ftsYarWAvwAAdgVs6
pAKdwy6ZQh9yCVuZgRHBmZvu2JmxehpMMsCDk7hhMJgurd1z86Nf2DOhEP6BbEu7rqUJijOhQHSF
F/WFdt7YOjl4GHmAOaaFTfvyT9PW7VY62UMRKP5/bJNaBLCpEzZOCyrCYMTzvg6YbWtYJ3eds2AF
Agy3PvFFi5gyn9Zl6+PaAhS7p1RcSW2Sv/c09v62UmiKXPIxTWyBxK/4WCKZ3tGG93jFaFJ2ypAZ
iN+u4DLWuMLlsOSs46Z346RcelMGqjXZ6Lz+7qRDsULlOTuIjH5AzPSok45FT3tA+GkekWPXW02T
j1n7OpjjASzFtEMi7UmhziT9bM7WdU4++zVTCEt7j1VaGG0q5It0kN9XRYE6mEBUY1p57gjDEbs4
Ub0/UI05olFBCOVFPPmqrSTrRXc2e8uH6b0vpZP4ONfMNiYqDXwHFBmwhqMQoyvOvWJRQURifQv9
zmw+5Ubk97xelsnp6hsm6HeL5rq+jAmQq6fGdRi49cP3/CvmZSmkOKel81RBRcBbBzNPcmPW77M3
xIAoCR/xs0FfJUKwZhvseN8PlE8wQskjs8tbIkoXyUGVvVyNm14wZLCP4nQTOLqOlp08RDGLMjpB
8o/DaopJHTBT3uztVkN9je0LX0BtRdjXOFTAq6uWxO+t+TvUFymS2w6+B2iwAEmzVMUI/1/fJlkC
PFC3EnH3z4METL/JuWwsoWymJa7U9I2e1a0BGJx5oVjH5+4Un+1r9DH6ceuR85pgApMv5bBiTc+9
BKGQOIbX1hUpx/3ntLVAIO2qDGxkiHMZvrG4TuMIkRIyrIY6lOkx61UOBEj95c3kwEea6+Zr+iPM
MwEZld3qVrG5mD//YHSdlP20htRnnyuErnD74JZqxKh6ibW8SzKDeI5NVgBwdL1iNWGMmUH0IlI7
O4Ftc5rshmpD/fe/PGR7oWwZzPBgaYvVAsf/l2q1AI8B0n3iaY/cd6NTYVWHcVJikrIwNfBl3d+n
nLDSoZOhdOCdmvHVPVGgzRUOGxxJO8yQ/mNhoBJi0o2XwxEArLj+g7khTeroQIUS+TEvtS90+k4W
TD4xJbXP67Xfa3/OMk0RTe9e7fZYCDqKJxIfvJkKi9V/UB7MjKAUj9jQ9QxST0dtQvuJoSFe4jjm
xgzFoeQndLJyZu8yrxVh0W+S7601e0H/GX03YQfraB3Lsgdg1ZInW/Cvsamh9+zKtUxBgO9+smEz
H18cy9sCaoCoGMxc7tbR0FsaFKjkQ9eY4aJpKOdDrlNJjY1QIBqAZYWx41Wx9w7VborXc5zM3LZX
gotBYRnQk0PMoeK3SPhZkFO7eR7AVAN4z7uMqwhj2KCrT3ldj4PeTISR/Qgz38ffgaM9KzV/QEZg
RX3gexe+MSaOWT2ZoBKUfHHP+Lbyg5Nyqfmv4pzBnwSpIDRyfvkucdHnjG7DRLAKQHKEjq32ZUZg
BogS4kT9EMZxMQjBxB2kXS57RM6YlBQjRrJsbQLqWP0afDgBPaJKaWj6wDfwrhaVjxVyj656F08U
c/Yrv4AcbeeWkNjCig+VVmCSE2wvyAyJ+Yijyx5C68+LEfdf3pjmbX+LRQLi4tzIlJuFuT+gKaWw
riog6nruvZXy++QWlte6na91aL2/4HKA0RzXIRg8ncx/fpjunvWc12jtgWatRfo7G9AvylM1HMSj
qyY90fc6jGWyOYOC6NWVVbcDVDf/Gq2/Wh0c4uqlLbfhRbHsSdKo+Efy7p3k2kxDHDcBYwqejZ7d
ffIdlXEE8scjEpKswmPCbXZhvSlkDWmy7EF8h5MaOivV4VojPDuOYLb/XN9sLogoDKi593H3JyEx
3yVJmiswazfhTOaCkEcpeg4oy6R1YXffr2IYfd83Q7J/tjGFDMS29ZoYmqSrOsfLL8SnSXO9gRnu
ZyJnNkrvczh5VcVNvH5LgmXUqGjzNqJ8A7eHfEjfK81WBl0zA8dV3n4OyJClqZQmxk0z72yF/WwD
MDWxvPH2LbAtTm/0HG9zW5W9edWeUVIMcBFCHb4jQGUsApPqiy18AQ0BNoEQbWpaw1VazYd8RscT
98EeK7aXLpyzezVvViIp4Ra9o3FrBEyZ7O0DwGzNv3dsxPPn3Rz+syh2iWhqqbwBb4ULBZIQGu7T
qM++SM1nPUTUmNoHJ+VcvHx9IdxXfOmnRATl05t01XnMEGUREmbLUVa86NIxOEbjcM1w77zV4w5H
szUvNpz72GooKEx8PcRuLQ2gDu/AC6zfQXDBD/EohIpL5/Z3k8QnBhkPn/YCBB0bzWGcCRejdyXy
ryW5fIE6AtSdpeC0D1fUCXKMIVqPEwnXlpnHeZsaUS3/4vB8rfmvH+G6RcjSl+CIVViWktJrlQ6g
fEUg6X3ex1vETh5EbY8cpIuNfIN4+kK6nhgTCb9t1VM1040P7uB9ZfJK25ymQwQRqlIXL/gm36xR
j7Sr5D0Z5b4y1oAO4UapHNPvPfpMuAvFHmltD+2AeuSHYc2fSXQ8LFNirVIYo74cT0g6u/DBgtMY
gbl+nH7GMJjfM4I649LcCAgDB04u2+agSG1APBs7HMSXp+YwcI/LtRFhffyL4gro0vVC68+uIhUh
/QC2aoDKgGRYGDL3mPy/jm81QldP+WFZPBXS1j/tzVkxk3vMr+5EfFLKcjhm7iCc/7Ls1O/dmyjR
no1nWJwwWQkFQEmfxpGrvOSUisXuMBL3QHHtmDGbQa+aululfdwS5FOaCvR0JCSAEPx6+SBeZJmu
AcKDo/VpnoK/3CgeeaIjbQewVBKPCjsk2WQHFfl9dTKt2iNEbS8mEZp0vSChSWComkbmZEn6rp17
NzpmzqFq4PATqZJpkwqW+3Ew4d6EbL8OJEmiyjyuZ/FPyue7HkPh24Xnn2Ai0ZfJ4nVNzxKFEyuH
jhyf+r5Ke7QHCmkofB5WSdmTqaVi0eqQ9tLzmBephWDPV+N0ksNzcitYpWacK+HhzOldTlgxAgNA
lnGXLycKqaAsx4K0FfViWG4Ce03zmwzJZXvH0bQRRL784o6VCKjPniGg2qpe1ixyE8uuDcTkhR6k
XY2NpWGYpIO4X9HRTTLiGgd23cXRcfyq8UM73oJzWPrPbrKNOv9htvC6kIZQfwPRVLUjOobKAeZb
mAv87GrdTbjBsmZ9WO9bkrbpfSG7abaSua+KTtsnESPrDxyiDfJDN71rNt2JTjczfH2UQx7U6+z6
RQ3IjBYTt1LX1//pIa85zhvGtjOs9wj19U+I/wa9G5QcvKkep2XIWALzh28KgnzHX7QfD/NqEcbI
X4Iv4/r0kGmj/4IYvzns5YiS3Lbe4oCFW/6KnDrPc8C2+Dh2/6pUErPV0qUfkQitk7yvy+gUvH8x
FagH0KbGNSzW2VW6C749BZ4bU0JKOATVVtWR+eZ51VhCU3KQxOzZ9n4V17YP/YWoaFH6jEu+JA97
dvgTM4pLg22GgjTHzgYNLYiaRpk/fj6t+udPqzn0i5z9hu3UbsNpidLUx7KPRIZ/15eO0HP61q+j
ViU2wsmTLS/bkye0Xs7x48lFmb8WCWjsVijlC0Kbmosusge7FXut39Ijjosl
`protect end_protected
