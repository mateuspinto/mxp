`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
FpqRCKMTdCLa22tqzbUMJenDLiKaFUxqLdYtuHi2RkGY1+92xTnRfQPh7i6K3rJBnmpRKA45/nhB
HbOo0q1ubdPzlKbM33FddEbGDc+3DgVlS+yX/uGbum1QbkZMm7cK/nxAHzF6OS9jHj7UIvVMSIY0
GIyc+BCkRQp6UXAdG1B+FHRH9XloI2m4vQ/VQh04TQPyygwYLLjdmh9xmn/WLrz8p0xCTdvk+sUJ
BAH8odFLqsVHz5k0mZ2yBPssxudf3bypFvCNlVaSiAsxnOgvc5VNr18fKg50vkVnGFs1FX4DgM64
Fz3nvcp2dZCRcO0KmeTg8KAil0is9p5TxBjw4Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="w4VyBNHaStS4q/IccoC7sPqKAB2WD2o3GQPHDY/fyNQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`protect data_block
J/myB+54pYEkGo5GIbKnQeNCxlQRreeM4/LFh7zjBs6HzLGwhXXP5KZrzY+SRKttLaoa/XouZTvh
ZQIkrbwGjc/KCdZBH1KySiAK1eXddnUgU98OfbdJNHAxMcGdo2/FO37HiVPih31YaxUtmrNV4UFE
Ot2xwR+5wCghoHzCEK8EKyPyPZRKDRidTInnpwnkiDTov9/khvCd2ULk95d6ni1RxeME6+RuT4Vf
/bJ2/twbpGlPx7+TFUt9d23m7KYDaBrTZU4Ei/GCmtjtsDFlJ/f1qC35g6Xc3oQU0fmNdbS5UHWb
WzGufh1Jgmh48VUUaxn8vp4J49AIF+3SoOg4k/DCRvSuZoGqE/xW3JxTDAHdjcUjhWfdrWHRDYcX
FgjEkruAaV0Qbe+wTdhYOJhzTSSlqxqe2LoEZrxPTTGxMM1lGzj+tvhKI7aTQLTNx6PYmiR6Szg2
HFmp5dqXSIQ9pxhaSo169nDs3S0K90l1SG+3tLwVHV672/SaOlb3vQXB3AThz/5MiHwG0GWNG27J
/Z4Jddw1JIXo+5yIVvoudW+BMVD778p8Ob2n5Vo3e5COhXJbFjGF7f03pcVSJOF6sp1BID1dgiqs
pWq4GhrKqWotYQ7VjPKzcEroRLlj8rPwe/qaSQBGycdTYYufIzRHJRjd4BgEJhyOgd+RZMvpKAeC
aiXzUsHL5JM4dSKhR2xNbbO/UCBBkTgUYAlQHkj3nIBibo3qZyASRSA8NB7Ctd4eFr9wXhL316jQ
7ueVCk7Rq4wFya/kCOXMsBsoFzAoOudFvhzEnYk3HpLSK2BCX+i61kKlVOnA1NSk5psN+uhdeVRJ
SF1XYoVKEOLUCr/QPqCk9WpbNWiUeWD4mokt303KTP4zh6/70Oz9P785Tmfc2eB2M/JloYg2JI5O
BFBQX/+1sEHJfaZ/VMg381JNMfH4od3Phr+zMCfDLSX9Ta/7rteJvTKTWCXsZmJmvOY/TC+QItoc
TWgcXlXJwJ5Zw4411YN9Um5o5dbc27RG+HLsMPCw9NlAFTyzVmHB/M/KDuwglaVp6UGNHnCFxegr
X1EomgM7HI3Tx0NzYetsCxVpAIFbWxRRZSILs4NLbag3QfZmbJSrzLKWM1RmHNXwzDBnzD9XJzZn
4s9iElI8ERWTuv/bhq3KtMqKT5mgtiLRnYiq5mMAyjZsQAcLLOZ2PEp4sWWw7soE9UuVnBzDSKIl
/2ew0xhnu/Ro0YrCeEcem54m6vZlyR/cZcru+PEg0/dJwqj8TA7h/R/mcoGGkUyxDNgtJRzOksCl
taRUv8EVLnBhzVVsiW2TFDP4C2BUmITiIydHNhiBNrHFDZSXKcHcjLU4kHxocKvvmtqOV9ojDjp7
1GzrAfm8yOgSIN+IV4azf1A/yzK45FOv9c9N+jUssBR5lhnCMWdezB5BTZDzRvItNfj/zc0RHo9X
4JMktMFvsgnORpfq9t2pZJjXKOuianWhwoDFMEBJT0bs+TBsinnfaBZZXXJiorD9oT3iywkiDjO3
/UsZrusUA4WjWPpHj4icEIOH8k+42V+dXVEv3QmXrj4QbID0eaXbjGHHhkFDE2iKj/CGzXPuJuVu
KMR0sjRgfRpT244QXKbebxhIe6nSUw4qd2XmfR1LQ00SW5pS64OR4H7bwcoQQFZ3/pWo+B0Mr4hD
TuN6xCjN2BMmlcMjp2VNr9bBLvDzi81F1kQ2HraqqaFzntH8+7ibY//QL+87GTzxsIbC8FutCB5a
XPDuvMbXuFut5sghULFTri8ZQJLPBYctERO5fh+jQiNJO0WGVlByiqIy8kBGBu3v11cHPz8ZpfD1
DJY2EMY9E307JQveCcYai90zhonWrOzUdK7Pb1ofk1m+F+PwKAKlueKsm5ycJDMOEq1jnr/NpUBJ
6sJZAek0MV6fNc6XodaGX2ShAgi4TqhmgjvhhR8ETy/QxbVKZeO/mbhWrPGpVDvkCtDsgTyA2kSk
TuIb4QMAqel87k0bORsgQnKz9wKbx0esfmrc5KnoR4MVuR38PUfaArWpgfQskYYYJEO371vjc92z
Ai2IVg2yl/gObX8KoAkqIyCkVlz7NEFtkwUqkmuWuSH5dqeoqZg0v1bEo4TgrWHnBasdgJAKTNFl
jMVVqtmHRPiJpil14UsAXM1DE7hbgbHvmKrAbcenrvg6VxWtzOI0Blrn0/wutVcXu/BT7FVKKVq5
AjyXGrpfpOUoaDM/rIfMvNI1ESN6PDmlVpEnFQzAkSC1gDhMYYYBXC20TUFGcVayAPbBz2Y2b77j
+e3JNevc+LLb0FHn+R9k53dpm6dEHtBjR99Hgt7l5bkxn3QxQRywHtKpdhEvATT5VzQlv6WjrFsT
9OnsJtfNPVtMBt+FO3KR4TkecpKT400vEEn63Xs0/ZpQLBSvK9gedCvngj0NlJS/rN6kQSdBfppT
oA+hBCgeSzPnpavD2mSw0RLdh2V/KmF9xcB/2igcKMf9Re0ms2gWS9Fz2IrIqGE3iUPM3tv10iNH
XLXNScz/p/aOIliejxr37TniDKh0t5PPnP3/J3TWbZesxuIPqOuVyLc44FVUvAX0j11tSftQwBJw
GY1vGCdnnQm5VWwya95M5pdzP9ObfNFxb0hWrv9xdETDxjnj8IhgGooXPlsXFnmCn71BtJbmkTPw
amtoMGHCE3yJ5ibBbS9wXXj3ezseH3mrigCSZY1ViHGV38ybdXQd88AbgARkdNHHE50BWOUk11Za
88Asdjj0Cjsu981enJ0Hzin3Jdn38IwVGbclJk+IHS1AcQ12AU+TGCjj1BV307GfGvp/s59EQxtT
H3ckQuHYD7BPgFE5mEEO8EN5Ljfb0qPoXsqP2TKpsBYFLo0jusCfu17V47riAhFQ6Jt1tNcMfqqF
A9W3M490lg+W6/n9LQf9xjsVCbiNTxUOTvGH/vZ4O0LiZZUx7efs46owi0eZNzqbWc1nT48s82Ga
fbEl7eO/iOSLH2dQQmBijKPcO8nCWk+bJ2KhANE98F8t4p6uMIKGx4lS9mUlarorA9S0GZLcxaK2
z2Nf3XFZjVIFvboB6rjwxDIy71iDuxcQe6eDgpHL824KkIzHuyxYk1mSkw3YSWG3p40dfM1CenFE
UGievPpi6JabQRN7OkaSj0qjCYa1w5DZnkEmYKtf3AyALXiRiSnBB8k6AkEul9NNutvolkAs1rhY
YykUGTJ+2tqhA/luwpEkflP94UqldMH+WXqqujnwL8EnV9y8l5oY65TtPzqtZJ8DEpuBh3HXuafr
H/o+ThJjxDUR5I1z+0k5Aesmjx2B3r1U8Giv7VfV+ldvxJ2U25HwJ5VGmugESidzXJl4mN0OtDJ6
iyEw/yDUqdtfM2HorNarucxQ1xev5bP1tw3hv/aPevmoVKLzSRfZX9WFTjDGE5z0dBGrEqIbidyj
VetzjReH7qY1OEZDRXo9/q9a/uI8CfiK8D1ig6RN6OZx9Fm8YYP5He5GOiKmK4Y03meMVDA9apvP
tP48nT7hWDvs53EtJqchTNyFUm+Q/O7dh5LkxTjOa90499KIDWHDOIdia597dVxiAZGRe9nHglnv
wNymj6yB2MZj78Ym9JY1dt6MFXCg52ouQenUHZQwGyB6YCJAtwYFrqUdjT6DZpAkiR9ifZyjaeuq
Ndb9cQ4OpSRrVpWwoelVFWLIfFmYcxIawTC1IreNyBovo6ymrZrj/lpzwQ1HDLTxnawttRxOAAks
LvmxPz059xWg8+tbZvbVS5/5b3Q5xD7lQmrvnsPx8Kkz7m3Lf7PzhdQPPfraIiJFIX8d4sDxGucr
kejxQPF7JNWhJgZcg5BwDpqfmd0UUeM2WdSH0SyVeyM+GrJ59y80lv0wof+d122gWF2zoEHfgzXj
FXkWPSEyv+PwrwVKYofcaR6tH3CbO+oqPluNX3S6ZncxO6MhexGHh6NTADEARdjhXYpWpveXeeBp
Vn4IM+8qx45fjEFOdukeFgo+WigKrkQWTT3dmfMARAXx8QZbjMtzoRmX9lKtGnUIbrQyOob5aGo/
/XkArbR2DWJke1hr9XaP/Qr3VWTO7IjQP1ABPTMRo+ACCtrsukpsvEuGlOqfeGgnv1ng0vh0wb94
9RsjIJZ9eCOEUNaJpjqQQSU+AUhhTmdUhN4qqCv5/rqQxFW/thGkNnY37mLWx3xUTOBnp+Mkdb0v
KpucIv8f+23fox8dNqfojRPhsmCd560yJil/0xFO8d02k8tvkwBEd3fhrP2RNWON8QXZEWWmI03Z
gUo5O+ZNf9mhxWjX6QwGaQsLiFOUtLFLFXlVIl93qd3++6Dw3TV2Q7MN0qpPkoqfGX3Z7jn0IJgK
9jigvJ5qQpf7UO2l2c49ylttQABwtfx8TWHZ2Rkdf+6RhV2QSrNZHcc7E4OWaajciI1/dZtr/Sma
VRC21NDzF/WNxhOsfCgU5LMjMk8V+N4TIN4TS0ZozI+prcj2+TXzKsMV9WdZgMKgKmQixnilTRwD
j1UtWji1kiyUc0wkry/DFLA5MbI2hQH9ow4ZbObfa973AehnHdf5BzlBeNkrQEpGIrxLwZxElrbJ
jJuo8kwxKT2IepU0/1om8Za/miOslMhZ04wAarLIHmwAVGwB9HgVNXhL2SierQrrffYsfej97Vmt
IzkFTy84axFFlmTuuCTMETyPSTBy8FqEPUm0wYmz3sV3+V5srUDLeaeXZUUN8ly2KA73Akbcm6w1
T6d+TT2qq1DWCdkmMz8ER1yVZ0OV18IzKDC2FAKU8WlUGRhICtT2lFbNsbsKryyaO5u0jOON8zOZ
QvTESMF4nUq0K+Fw81QLzVdZtx0wPqWC0V8eAwyKtWgL+yYXyIN+udgPSexKYRuaSxZueZ//9d/c
Jrg1aP8/bT6X7ZkpN406ugBH+mzuP1CvDKbL89sMRAXxniPeh4Kme9XsRdk14iMfbzWuIQWIMZtP
akd8UOS5bNNGeastra3Q3a9SSoGHrpJiKvD5caTdiaAoO+s9AN3qqxjm6GvRxMbGPMzr9JIEsmJX
5GTSggU6Al5FGBxbFsdPHSyfoFHh0ER/Bwav/clpnh0vEE5IB2+bQoj24+qx5IMyrZToDqKzuniE
kmxGxUan4cnI8/yym0yBCqdmIHgli35aJyvH+QiTLhFlZesVayw2AO1ngzeBUuNhlCMlSZ3U3Jlu
URN7yqnctcoSdPaAWHkyttCSsjQIcDXKltoaqiW96f1nfWm5T1XWS/iXjpzD7XUb6Hjx3ADykt2v
w4RbzCFrQLj+/dvq4cjZTy1qGt7TWyB665XdL/pDNKQjvpmRBz6jk+A3DQ7JoRQNPdfAsntHNuwt
T/bnPUHvdbKesGfS2QLy9DwrIY6eaTHrw8H3krpAoJ/7/1f/7t3W/UhG7oqgkese6Svl39fg1AT+
WsYhRXsu44SsNROlucQj1fvl8m/Wch/YMCCTICEMf2mKVkzzr8wPBuaJRRUnX8thQYsbN13HQLso
fF9dMXzYC4TNPsS5dEYnveukDk067dFczGytA6nnkD6z0B4PGUrH8QhBH/n0Q4D9cVZ52ZAkq9gn
UWocg951AJQ0k14GgA81GfJNBNQhRsW9fHyGmgLoAqpJMWKUvXmkJ3O/1XXKO1G4k/9F7wRCnDLj
x5XQgxiZIb1ceS/ivnUc09J6T+fsap3w/ZeItAg7wkUgZy2TCamjxovR6bZPoEmSLuxmf+TFJkzn
KY8uFYSy2q6/JbP+/KVfmllB+rv9ww+7E2Sc9Z48OLS4uAVdLPh6k1/mYtJpN4Ww0+a2hYiOSCyp
L7xkyQ5+0kIrLcVXIwiszDEJjuFPkOHe1nXTA92+3KwyRGHqliQUlbrEfVWD5sCZHcHQlPIyhk3C
qypvcAiSy4Z2abnrVIBE6Vaa/aVVt4eViQweepoydWvbuYHlJiCuNvq66rKOzRwCQWtnOYx+7SA2
mXwChnmYVHsYISV61pdCat/tZqeCMCeL7ldyeIun5xABcD6I+7QLyFx9LbWYvYgg3HZUSa6T/OAv
92mOEVvtrlh3OfQBr4TCFwrbYpe48Mst5FlR04gXCGaFCBrF8Wu1BCXSCEJefis4fA6DGeJ2e4XY
TadhgOmnwoo7lPHR4YdgGn6nJtxeV9OgLDWZO2LAbIsFQwgUel/AvqLyyHCKbzXY/1u7ciEkVDyq
Q3Rk45SN4CEtC47+TZKGfiZA6g5MAWzYyRrXP9sebpfacRJijZITZziC+ozYVhzgj8Ny2fVoqTSb
FdMhIZO57rNwJC0KByPXWSg9MJV04G4Pe6aQ4RGqR1yozmDnQyJMggBAspHLw+ILrDTc09YQdk6l
YTRi1+HPgM/Z3B1hp7Fe2T/9JaNGbF8h4KEbTKdcYFEQQn10aYMKSczoZSya3CnTvoehT48tHtKF
B8wGPsDTae2RjT7hkktn9ScdZjqkZewrGCms8bUWCQ0PywLfE0pcFm5oUz/kMAC9L710zriM0euQ
e0iZP3/W9hEWTsInClhV76B05E6oQ7DJvaiMS5J8q+HBgFWFgKXO5ulKE4YVnv47HocCxKQz5u+u
51+VPD2jt8XB8PNvV985tXy26mYlFYd7V0mk85qJS5OvptaC/nWMx0k7qOt9ustguSaJgOF3Lkyu
gAJF1vp8UzVNj8XzcSCiOkmss4d9FLwxg3UXytERNwAs9Q8MWvNz6VCUa0wSwZoFJg3ZAEjksxx/
Ksw1ccy5DE2FiSCrocrsO6YkYdsauaZfYBHzdKeLzy4wGqrqGvSTvqiHj3x1yEL9OC3yMSoo+58Z
0gXYNsOEjXN7u39KIh70UDsRMv7V/i5fiooau94Vysw64DgV6kL7S/aCpjfYBUFSIiUO4Uxzk/9j
HAeklfF12Q42UWrJxfpGRhdpDcHMKWIkG0485uOmHy1g5O0QtdwdjmbiBx8bkuCJmEvbUiQkr4KX
VFUqIYDQaLc4cLs7QcOpSva14OH+U9CcLBqyFfIBkAaYexkIniDIrKrIq3M3ooG2+ch3Tr/XFwmq
UVMYMSlPshXgO8eU/DjacYMyh6C/jrpNnT01qeMNblDAntGo35LJZXspN8lI0b9XxgrxTFV09pl9
J81Fx02iADvwJyA3Lr404ELI0wZM1/jM+eRRvH492yGXDQo4KAYmaZnM9cAzEOIMA5tmeVx9259l
OjxjkqxvRztEbGp74wylYs6blbJNFxpYMBI/9cBe6QZpU0L9cgxFoCFAdgba91qEpkyNakrXlLTH
QBx9AlH1rPpOvxygijfRGluvOrNepD/aKIRlWH0RkZyzATLjHJuRjaCTp82ZV9/vi1L+GAPp867R
iG9U/ecyhG5glMoZ7M6qZjdTnU2Fn8qXSLF3DijPe6wbYo2DSUpFSxki5qRGchXjPHD1/3M6snJc
ayDX0qo5W0IMdD+WOa9q+RNGd2kgxatKdcWNoWJwdy2q6tsa8rQf+wEOXKLmU8FwwColWCQmd/pl
S1/lS4z7oAPoSBpUmV6HNCyf+KIDOWryPC0lhnXsHnJ3+brO92l3WPa5Zysmo1Mqp8JbdUsqvPq3
HKfgCGZklHY9R+pdWCdSbguUp6HP+Sqn+A+z0vAxfLzKYm20oGeXxf2I0mYq3UZxwVa4KnPSqSUf
zube4kRfNJDcyFjIQXAlL+oH/bDjvW1jAySuoXSUrhPDx2mrnJdQrVzQ2u3gBBvTLEmBJgoi5b4T
9BNeH+ZaYmwUgVdpYndblL0q/L6gFqzqgdbb1Ireullildg0XIwd/7OmVGm/0Yd6Fcm1dZ+xSYyP
2mBjW/AuSgSJUMbNoQqU9VIORVZt6IO1m87gwyV8T/k6KsKstvTmm3vVCqRRlvWYrI8KWDAOEsPj
MxJ4KLcMbmaZVTG4ee3YHKLt+108BTPWIwl5qV824SAuKpNLi9WtwA9McB45oVm/kWejXZpCb30A
0/9OFiG1XgPRXbdo4LK/ecrfsZqV6PNzfHBqC73ywQfNSgS6WTc9g/SmzwzavI2SeXCd+xf3zouM
kJ974Jc63IUqAl9yM8XsB6pZARF2YmKO/3m8MKv3GsgmvBe5Q97c9i/JcChDF86Hnlc7HUKObuQa
1kuvjT74bMSeU1gVIn4eZPM0jI87IkAQs6456U00qTxM2k9lQwWE4kErHLgDMez/JA+K3/By5eic
sNwIKXvbGsWmW1yGo7VCHQTa7pO8npodbrUbOr05EQt67OWSA6uqW3RBzs+YCxsiRnEqtmoN4bEB
2wyUGhJMJh/HFdhYZ13hkDartZsCwSJJf1ZYVd8I5/8ncp1GNGFNjver2D++mkC5Sgk3a0nwzMmk
SY3dSC1bCVQ8E6kZBELPgrDqTI/01FM6bh2Lb2POsgX69mIAVk8uqU5ItMMSj1s6/50Xk5WuqCj4
HfDhLqKkrhp+HqqZvaWa2tnUfhwQ6QEYo1OC5QuFJKa5dZQm2+J5Af+jtNuSU//VzmwUceSar+aG
3JeadNPiSfY2mOifNVbala2juYN3sqc4Vxd3L/wWPQJ5nViehLzQnx5mX3m7yzCbBY6BNDSmJ/N4
tspabmMUK54r8XcerWrBq9Dz6uwYdebQsDv+YbmQzlNIKz9yE76Nk9TvaW9ujYucCil/AEKyngr5
Z/UuAW5c2g1qsrS09CrSGa7hsMTb+Cr5Taf6dgkdQ3hvaXY4hziaT47Q2gaQVAizmV/gB5tz8z4F
ivJ96wfa+ZBbmRy/y0y0D4xyvHqMhIfNRtHoKX1ITv+1d01Fn+vL+NRkbBrK/6RrAq1kvdFQerdt
ModIqMjNGI5geZGzumTp5oRyovwt9I1KW1BEsUqCLBEcNHXK7nD2lyZZ3KEdG0J5x/Dn/d+DdVUf
Dw2+inTVWnzcbAV7n3USnSm+CprUGNsAOQALYSU+7nv/SX+HbpM9abAuGdSLeOKE4Qc2DICG2Uf8
OH+Qo9DqIenCLSgYINRef4ysJlXr8Zkvzq2KVE6E88SgMPdZ5oyHaPHiqfU1eVwwBCySBbS/9zjI
T0C6u+tb0UA6o5wi78ru8lu8hUKqOCrCNlDpkhRFyeTF+QrX6ckZ/c/AqZAYT3pJWIiqd/cYvbUd
ijngSPnsuJMFqPScqrmz62/c/I/QvG1Smup+J5qrnSSzV844Ol/n2+DM4kb96bgMZSpqprpDkXip
gLzT+3sCIqNnDGyl+8lx48kRrBDhHIiaP6kdfXppIJS+zxbm779qhwzR1kuPkjUJNT+UwyZM96JP
R53UxmycEYGGZtXBkOhs+KfQ6AvUHWwz/Ll6BmcDOF1tpvHZvPGjnRG8lXZy0VGYr0YmqJot6PkZ
9ppdMvywvYlrUnbvXSSWUdYEU6TvKwxjwDd16L8DL/aWxMhNWs8IRumVRZNJDsMMOZhBuQCmGnr7
RSHRCleTs0o4b15jk0l9FxtIXhbT2ojEh5/0FYCqub1gcfM+3JZ9CapYAPPDRq+ih4QW/1SeMsVK
F9PG0SeJLppNG6uxm/y9Th5+zGdjD4GTiTrd9C4SzDJsmbFVmJUEtWr8+euQ0RJntimuNtjUPGYk
/3a5bfOB7dOP0QPK8NBoAgXXvK3gHULD5Cn2d+mar2mZ/b/RmyQKbv069MrZ2RebSUAyvzX/6/wK
lxEguXNl3WlecnQuJdusFK/AjpMVxmf7S3eLO/zTUBhQ61vCObr9+y1BVKhFLnLvInZC7uTHNpVH
4AOp0yzvhAB7lKNYG6qNVug3zG01hK8ylomng5h8CwTO+2YhlsS0wUmSx1rGJTgksbXnk4+Q14IK
Vx+wrh2mMLd8ReOUvhWSxXTKQRV6FV3KH1a8zkQS3c+5IlgP53OZdEh5vpLUXXuQgJTws6Uogx3+
NC1f4x2V92iRUrKofUmjx6Jyd4Ey+/E5EEf6rT5+4ntIpLIvGPFvGRtka13wbDhqpUcGHDt2lFVA
xUd8MNYIybu8rLFduGDW4XEc+FkbDFkOG7sI1ntTv8AOLILXexLro4HKVC2cQa9pG6B7EzQ9kGVi
59yNadzsRsSDxC6aanZX/RItn/9q/vaaScTljvXbPWCm30D45TXZIGBnUkNYS0tcNiYBEiqYcvfY
b2o3rigJIAHWhVYylZgD2OcwVYOkTEAzXBObXFL8Wll5NupPg0b39+KLYjxV/HlR5n/Mci6F5pf+
Y3xZ28t6/i4MXwFaPxmMhxsdwgF/A4PY7cV7p3cLXBwDDqYEUE4BnnweerHeuzZ8WRBcJK3NQGzQ
8Ic0LCNud/C0KTjxmCg5NpkeqKA5RNY0/Lfta28A1vZkshbKuEmZgObewGRCTyRh4v1LrjuDR+tm
ZskvJjPCXXpIxuxrNz59Zgky4hjYx5Tc5+TuyGwt0G69SI4miOtctnhD7g4UOcZunV1T1q5+fPCy
o7gamZ+T7COKXL92HJe4scz6LKfqPS4f9qrY0WiRQ8uKkzSE/cNfgxUn6ljBzHMpICA395yDga85
t7AaQoUMCql9aFzVqq3IImMgssAJrl8DZdyEJ5cdW60qyJNWuXlEy0zdh8e2Er2z0RB9C0aAEGFP
jJnz5BKPQTvVJA8E6C6QjcsxzY3beIF6UImiDmM7rAcLn2XPs+e7ol57iHrllfjwunAmzF4N93Eg
hcviuRB65zpwdr+5dYDx8T0mnBsh4ShrNo9KXHRTk9LyVXhs25nVOgCNwH5y+JC1OCywBKn4cN4Z
A+UDWkjfxzItnkaTD3zKgBiVV22tM7XlXKCzW/4ZesfCoPugQydCTtN75+hBlXMIvNKjc+ApfL7i
dgA5fjjOUEjeDn8x96jStOje3/va5+807FngsdRlmPjEYA4pql2m7KukhHOBDxKBp16Q2S9E0EJg
FiXzbOLf4I64rDEaKom1vpuA+E7nBf9b5zWcpccRecRtFpzZ0gl1Q+Ssv10FWsQcnmMD384gLZ4g
826zZepmy8GP30zTH/7MAyxkQP7MXE3hxOQlLDLeMgcxSq71H+n0vS1G977Cbcw/5Wm5oeh7p1xU
ks4CDxZPN73ZS27LwmJXPRxLMD7V/jnTnl3pvrBU7z6YWtpiuGgMEUsj+A1t/QUVxQVxWs/rXnjY
9TyATPLqoNNxH2v7to6mvFjF412Abl5+KBhxBzK1cd2nUW9GJYXIN+wsHh8fyZ/lgFRFfK4Qh2wm
rFh8Qn3t78CYytgYlGZ4+aQJTD5urxa1EWQGBr5f1QrnKLiAm5w4YNItriXcRiCtEOgS3y0V7BSX
nEtbviBuE5W5fvDAs0NHVHnDUOZw8ApSWs7R6T/oI12wOUHyNVfxXsj2HMrL5eDaEmVn+NbleXrh
/Rrayir51u9Q6p1NPo6soObhU0ID4RxF24pKavIDbp2peO/sosZgXoezsQgIaY/+Ugkw++M9vxsQ
rNWbQ10CsQ5l5LUuqxfwEO01nWSRXb0p82DcY9CLoi1b3wwAVuEbRLm5rb/Jt9dIeBOlEvHVL5pW
V+hU2mIkykYbuFMmFio3c9EdEv0ejXV1DpXQESoi3+z7IiWdbWEszr9IveHYvzWZEwwjsraqVrUv
IZgUaIPhnn4+dWxEe5AVaXiet1VKdpyzZoH7dh7ejagWZFVfaBX8YlcOPLTeuk9xs1t0lXnTtHXB
6wv0zuNI9oJvL1xm1KQHokKApVB8vhZxGldKE3fQvjx45MP9cnRC1YuPygMto/hQAkLOI+tUv0UL
aaSBC1Ewp5CXThpJZgvIXXGZEn8kTDPbuZnM6kbASwslTAydLeOSv03QoLaYzN0PhcCpuL8jZfla
z54HjKVinS0r6nEvegObTWnHCNmrvIykRoh2Q1cKqNrvgroGKK/N6a5u5ODcBUrc5lg5VgnvoDue
BXWSHhCkSJ4OkzqZNXiPbIUluGSgh77X1t25fXAQ4H0+GBVegi72sHkkFEYqqd36ly7Y3r1jRPAJ
rynh4IIykC9CT8/bgN0+jAmWGeQGWTfAFfYbfUpmtLjw+/x+cx/BMWRMkz7NxvgalSJrE9Y9QrDU
biW7X96a/Kuxl6icC4MEtpBvu6mH/nBw5nMKIBerRNoPR8vNf11/kye2KKACLtgs0BCLtv1/vfh8
PqAiKcCC3MtuHE0gIeOZD1pWBLyZJxMn4zUFmmn5RNf60EljjRPYqU0KDsruF83WT9fDmhmOuMYD
sI2jIbkeiaL2JGqk6xJ0nHkySR3/iSSXOnBUh2SQAEbehw2QgbyjAy0ojMu0NY1xR1WFqAZCmMwr
EF1xx+w75rxNHOeTYDcO6CMLESTJCXPhMAn2QVzbBlwHfxPsqzPcUeQojcu4ub6j0xpVA+PjS91p
aoTlLxklIeXsw9fVt6uU8yjbLDdiWNIhfuYuzCPb2RgeTPhJHGWDXeE0Pr5HeYFK4vrsYfl2rve2
FKYx25NfuUtk+V3/pTDrbfKxI5wFUOGkNTqka1dKbG1ef5kdxT/+qJEj9d+d+rlLwbExydcTtnQw
WI/oZ4yIPpaFAAK/xznZSR+JnBlYoEKjGBDq+AkCdjEOUbbpIwacFNuSQvLddVURU8sMlHqHqFc7
eKnUCD0iwWGa1DWUevFuXegLxecwe1yonKUyn0Na9oHW8HPi1pQUuOPc33+rC7pWEVRG36IwM3u7
dEjDH/4YZla8OUfIBTZuj0oOVnZ4KxCQZgGnh3JdNmlHaGOEbOiVGTLRnKOFLoTeEKi6fRANlA92
B7xxY3ISugEUcErbfWG7P8qSBxVgEUxzP16cUerOIebfPkuar4gRfdYXSTUDbUO2umBFvfHy9OzZ
V/YybXEwHzIWJxjNkbVebjYgtRqeG+EXevcuuaVmgwuS/532FVo2yJOszB3JoRg/YOgDebQUhLK7
jetBsn/YWDez66i0/fB46jRHG/x57bcB9bF6nKL6P9Vp9TaAOxfaKU0o0+wfItTuHqk5CVa26Pip
/WZRv2cAmOkOl56wIsSRoxvokH/crdOrflgCKALKkHNCEpkTWI/n7ztsJ9xSkLWNUuqrraNyZNRa
f+LBLyVoMpaWLDEkwxJXvbSRfYqvXkoCUt6GKvPuZ1oT67BVNOmmXpOXjxsgWXeySe7t3qIU2AGk
yMRYfeed9JtgNMUHSz+WhjKQcaPjHv6Txp0U+1QEYFoB1FKV3qqwZCSVTQPyD19ohFYqJcwgstfV
pqkOReK4wRZ86Jz52vM/zchMfUnDiM4EmUYQi+ary8IMHOHxtAeZYyBctko4lV+C9OUOyXnxR6AT
Zr8mKMZvbErg+vOLZFQgRKX3hujG1X5aGLpj5pZw3JpkqBBhB/uBMm127fbQnAg7WSez+eWtpoaB
YIkqGPjuygnY4MaSmAN1Hw2no5hMsJasYqP/mz3bjQHNA4QpnkMR3jUS7trjRmcSLZUcjdjFkoCt
HW9XO0DN60U419G8CyyYbNqDIdkg6SvP0Ld2Vqf5uCQ2poHewe9wvKgbZvuSIWOp9nkdVgz06dwx
jfZ2bFuUPWFV5sSZR3X072seHmyfSbnZES85Fo7ldHK295Fwr4VWPm7YlGNPItKTO9x55VcPtqAN
ToomTxq8Lmg+XG9jEeOalpeW2QYtl+8v6eqh62zpZDG9l1+JvZPEE1rMqekUGrq0kOqn+PgJMQhf
3P3OFluH3+QJqsZUUQxRdTSARnFNq+Df6nFt9MbUmPFq1oPtfYqPU+48DRwkD0N3B9vcZEgx+5ps
upUch5TkqH52kVButO3+UQnAJu2+Hg4TxafnJTll2q2IZczvVblLw0mwiA1bTjsfTUAIDm0zBB4O
7CKZ3ghmJB8fd6RexOu8VNbkG5iDKIFRUy5LjJEsu3VbhNCc+uumKwEhVIH3AM4tpWr7omUqknvj
Gp60Mlj2CZ3dt7YyXF5lCU90zEffZXPGQFXaLhMBagcpR3U8Mk5t9H/cso1vLXuuscHuauptvN0x
0fIxykq/9DvDLsb/9mOPE1Yw5sS35KOEA4Ukw+/2xdYPKZjRqJHvK0cYtGK6jj9OY8kmzrmVzpvY
3w3C9C4L2vLk9Z6w88ROOE0d73dUkmNMw5Y2uTggDs0sFUCr7GkDArRDe9hRW5DQYxAna5tss+Nu
QaZElmV6SBd7kEMe1DgA6gCBbH4xfvW8f3RKINjiTVMq+ZlcGN1J1bg9XLpWDkvFKOA9jkQ+e/kE
bvO/n0aloy1haoSP+vBPecCyB8mUQVQECSxEpfVSUriLUWI/EprbelpbsYlkG+vjc0/r9PgeOw2q
t8ub6FAUO2gBt/RwrMHSWINHFrJTT5cKe6EPJxpwMltzTkoqJfoGqprQphNRNSfXLZFuKjNkXalj
Cy5CSmm0aTXwtDqvQ5b1dDMXwNGc0Q8ITySjbPnLxxj83b4ZLHp/ALTTDyIS3NkHA298199bKknG
Y9NOg5sB3Azz8P/KGVnl89U3+BoebGeJOxMjLMS6d9f1slACbJfm80trLxvpGtJPvdvpEss1Ropf
zcbbmJpD4L0MbTYdQPUMRXrSJ7D+GQdaiAHpVZKHoRM4eeAojt7E43kGwp90fvf44EheHZQ1lFux
v74gC7rKKqyxYO18aA8X+xbuf/kBRiaCuFtDCF34brohu7kIe2Q2tzd/QRHjphEzaAd4Nau4Uuo7
It91V7H9YGle1hMniccGbsFLKa0oshcVMXYSDN0fj3hUY9EsIFLiXANdrv36nubnwLpWhgYTkGJ1
YSwo54vf/P/c7ypeQUFTtMhqJRjabFIrrvuEcE6eP5dmLx1dZS19nvM+y+bx+O5IB6kh0uMw7TZC
5BHB4BORTSctKQPQmVxkwLcRSWqbrzmqurF9WAQMYfbiv2mbAHlj+Z6JozvMKgTrI8B64ro4FiDW
Vb7yxGWONxG+pR0VrMnv1Kx27NLY2V7VpfMjpZ8pDsXJIW8iepXtgRcX2doKwS+peiLppnzUXdIk
pmh0Dh/biUOKt8ktc0ac43gfF0Tz8HG19eOYAgn3AZPPZrDIPEd3F1XvqjySF3pKA8a0XX12fGWj
rOeZFUEwD6RIBd+GWTRBkU+gSvwENiQF2DzL/2wFaFVzbIxeR7X+5NhRLOGJducl40bDP+jW6AHx
GWhtSiAzn5eO6zaWb5joYSJT3q8Tk+OJVxzr8qmrI0RMvT94gkUu2cybXer2Sy61kvGsRSnmtndS
V6hWYwFGZ05qvlw8Gk4XtrPzkY22E+8Hca1h8qi0p316bPPhvdZaIMFFqhadC1bLkFPjb12tdgE3
JnbJOnBvkdIzL+Fik2z8B4bG18/YuP6+DyJhZkPGYyjZZBmUEI7gGgEcJYGjkzNFvppMg2yDMOEJ
avebcG8M/bBzQ9YBbAbRkaAHC47tmn2fmLQe1mc31SIKxeA2JurnIKM8wXAOAgQVWnsZNw3rf7Td
zkiCqkqRiONHE4MjZMpKP9fmyxFnBrFJbm2Ero8TUm5pSkJa1Hkr5w8qUHZBXEx5Bwpcu4TpFA6z
E6SUl1Qpqh32QJT6XXvA7YHVI0MCDvLoiPP6q2NZtX0xzcZeHIOlr1z3gIVVUn4ROjJozUab5/H4
le/06A4G3YV7O+x/F9Mj9cBmN/2HuAfG7ndSfs7e6st1CH6LNsyJU7qLgHuKJHPXpG16O5k9Yvzo
C8A6wRBjeDyFvvIJmu+7+DLPjf2G4utYMAHS5USdx9z8yemO126IHS6DIe6my6cqfG702n6y2mzp
lVdoIG7ZS/yKKlCOFhRgsAfWJFls2vw8YUwl3og+lGUklQn4BBjsJIJZ4y4A23Qj/IZN0yevuFJe
CYsXFtuJ31A5NaG7Kjfsq5FUD5ciYhQTo7+tuwHN+JN8MatTNkORD0WTLm6b+LC0xVJSb7/1bmdg
8ReSSMGfW03o8iExqVwHjb8cPuAGjFESWFtIn5O0ckdGBh+ZZnxSRPXEMrIsBQOIVCyiA6xlj0Dv
rI3/Fjr1qZKe0/iWJA0Hur9Myhwhb2lJEDTv++zLdKuwzSE5M3H4rBaGzvDkh31/cRgE+Eh4IwvE
TxRmYs2t4OPpv5ckZ5Z+U4X7D9deW4o1yelb1lsPH94N5h4o04ryPgzxpZzQbosVqpcCQWKkVs/1
tMmuBE7bMobkUULzUOk=
`protect end_protected
