XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ih�}����J�a�n�1��NB,�N�g���Ħ�x:8~�����~� :��2^X����s�T��m=��tg'��܂
��;��i��PĒo�{NU�x�i/��}t��r���D�'�<g^:(�Ǻ$�b+É�
U�n�c��Y`�a���N[�)���?fC鷻���-�t��r$�c��Q�����D/\��8|!�e�y���RP�Ū\�B�h��9��v1���<� �7�a�MSoª	��U�����B o/ܫ��ݤ�r�#W��vY�Ocx �f1�uj'v��qJg)��n�n�$^�؛�(�%��o5v	6M���"�,�ͯ��앦\�L��]2�h��v��rn9U�V5����$����5��2�I?ogˈD�Ӝ�;:��'RQ'��y�0�A�Qq�K�%�{߶�H+��!�)�/�8`�'�(#*������}l��lq�I��hE*J�+��wJ�K%��(ݽ��i?J�ܖ��� ����d6�o2��!K��0����d^�v�VY�GIB��Gj��
��4�s��u���݋��!<��F�U�����p�|���Ֆ�i�<w�%\$P\��r8��7ZJGY6��%me�A�m��&�����RCs@/�'�+!�{�`���y�Y;�9Ը�l������k�.47fv(K����\�����*�iN;ը.���_��^��~ӟD
K���5bQ���.�<!�����v&I�8u�(ɱ�P+=��jB[5���9paXlxVHYEB     400     190��Sy�S� a?���C��p��>M�^4�r��A5I�M\�:������<Ã�=��y1E��&����1���NP��z�/e4
;��J8���K;-F`zY����é4�|;{�=�q(QkA�~�G��~����n^'֐�,���&R!Z�&!<$�ks��m�W����2+3v�J��b�J��5L�E���k)���ޚ1�&Fԇ1��	��g[ �ʵ�Z�|C�Ep�%[�G�~g�3�Ǖ_7�z�v���K�ݞ>�|���vo����A�ȫ��5�WD�r�pޙ�����9�ݶ�y �I�.J5&�>5���w7��/����^
qb�G˦k��1�\�9v'?CC���|��-��~�0��L�R���,��ϝ�lŐ��n��B�i� XlxVHYEB     400     1f0�ׄ��,39k�m/�����ȭ�Pnʮ�<�pG��o`t����d��WH�LL\�=\-Y���^I��r��wte��S<f��WǱ�AEƸ��	�����-��q�p�*�~m͵*��?�.�gi���$u�i���oX���V�r!�I�6n������&
��1 ĳ��#�w*��!@-��O"�=5Q���f3;5R�+�ߤ��������l�Te��2�cDT�jk7�Ԅ�k���-H�ۮ�!�!�d�i?ǕGSgW1��ܼ���SqU�Pm��J�ٳ��a`�c�{s���į�����li\R�|�I�rw����?�~>i��饺J}j�;11��*j����� e����W�Y�
!X�?թs���E�r"����(z~�A�b\�]�\�q�����k�kT02|
�[B�v�(�C�]��>�bȵ����Ӿ�j��lGb<�W�~��*8���� �+� Z�XlxVHYEB     400     200P���YËm0������|�6�q���]�|��R�-vx0�f�����8r����Ў����q(���p�㇣�rW+�%��K�$��*�3�2�Nc>%R��D� ��N��o+�y��V�,�k�yl7���k��)�'�D[��ͳ兽����x���L����ͥ7�M��T�əKӡ�BDN�W�{u�p]�'G?&�)�p\�JN����9@�B�=�x3b`!Z�"�{Z�Ӡ�qg\ҍ�x�}�zz�\�d�5%�x�T���5B�D]��!a��Ն4BLr�,Q�J�=9TH'��)����4�������\~@���6篗_ ���(��&����|8~����C�Ē�~�Yc�n���U�T0�}��Oc�p!i�s����y��(Ë?G*�	tȼI�Ɨʹ,W��sDj���/��e&!���= P\�S�W~q�b��K�`#g��.4m���!���ߺ�x�@\W6�]ŏ�ۢPyXlxVHYEB     197      f0�Pӯ+U|��{�	QN2d�B�S敌��F~ _i.����z��Ќ����b�^���1@�G�$$�F����%M�PS�?hJ�H����.b����~�mϩk�D���e-z�KUW)��d�d���e3"D�þ��U�g^�H�`�H���U�xƅ4����l�|rz��?Bi�K��/�:��{�x��q��{G��NG�ެ�h������l������1��?-|��1	ʂE(
+����Z�