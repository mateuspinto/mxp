��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Г8u7�~!K�e!8:���O��>w*~I�\z�XوV͚�i$�5Q�����̞�@��>����)��f���t@�@@���ӄ����sq�(����_��UH��ұ�b4���2��r#=�)�+Z��:�a)�����B��;\'5�bH�0}�H'��Z�q�"p�jz�k��.^�#�)��R�}�GΒ�� Q�[�:�&�g-}�d��"�8pL:�����a�}>S� `(�u �I�-~��c_�Ҟ_���"���S�=}]�`-#��,s��[����5��W�<8��
���=��4��V���>��ulI5�˾-!$�4t��������L�ݔ'x��z 8şذ�U�ȑAu��Ce��a�I�=�Vf�\H�vfi���b��v�6�
� ��һde$ڑM�� (p}��p.q�u����#�W0���Z���6�}�Cy�t��W��,Y)�p�H��]~��M_u�[�G�������⏅|n�87�ӺC6�:��,�R:J�
i�TX�IR<?� ����Y[��bo�]l�������W�^�Ж�[%��G��b��
��.%|��ʙve�t~��w�������{@��冒A��X����W�y׫X�t���R	���q�q<"�w&<C�1С�(��w�Մ��o����&�E7Lx�}v�e��,i�T8�2T󉀶L�W�R�;:E��P�^�8>�03��A��zyD;vZ�H�ׄ�Nة��%UF\���N��`�̠��,���
���M�4�1�,E�["�$2L����gWga���o�:Ǉ�����Ѻi���Vu�c���*S�$��H��pL&��7�I��U ��nۤ��*�{`�M��5��ʶ�B���k�B�6_�`���tvM�ȉ��7�`��=)vt�g���m�{���y������	� �'������p�'	�;���Ĕ��p�g���W e^{=KT����8�0f)#��ʸ!ȷ���T�\����3��1L��f@�4�BPFH�mؑ܇N=8�o������lǲ{�u�e�%�O(s-�����ՙ�Wgyz+��2��ߔ}���cmX��ͨ�~�:GѸ��J��MRh71�M��x�t��S�ӬiRo8y�xS]�t;&P��6��g��+�����Q)�f���]�Df���a��> �51ϧ�b�$ �Qb�+咺=es����py�o��_x��m��!\�-	L�&R)*��8�Wr�	Ywe&��c���Q�F���/�г �.�5"��u=r�V���bh�I��q�>z�X���_s�K���
=h�H΂<'�I�)2XȀ��K��n��U.��F���2
����K-�{����Rq�w�洞:��#�$�^���'(r�</���f���\��5��2������C8�=�F�ٵ�2��?�<=��y�������J���(��}��K�'�߈�'bpDv��_!�à`O�����Cyl�k�ad��Z�D����$��6�On�����У����+���]c�O�?�]�]�m���|s������
#	�{���D��7۱IbT����*���]���m�{*��H5ZB!��[\�ҷؾ�T��2C�� +�2����+�r�����2���J�~�P��{v�Qz�AĠV�]�5D������¼Z2��#����+{y��;���Ld:�l�kRK��H츊ꥃ���W�O]܎ًx�x���c��K�([-bI�D�V�*	l
��A�D��0�^H���CI�-)��L����v���02�M�,��9��r�G�x>9x�1�4G����H��.�-�����tyU��=��ec]}O�� �w:�k>Pw�0���g��KK'���k*�d�1&����-�TY��)�>cC�mQ�lYT;�K�e27�M�m��13��3('�E�T��w:gb=P� ˻Z�F��<�d���4a�Ѻ-ȗ��Ȱ�]��������_�N�9@�B���P���m-�߻�Z��I*ƙ�fbKƛA�.fg�R�������h�Owc�⤡�迆`Ǭx'4�߀��0�������+�ѡ
6��A��wj�m�
�,,R8�[�ޮ�n�tu�?����x�L`�z��{s�=l�V�O�(��#3;��Q2X�%Z?|�.Uj�P/����M�6F���!'A���e7T�P��P��}�s����HZB�oozS^���T@����R�7�~�7v�]���)b�5<qZys�b[+�=�;(/�cx� ��U�0{_��]�+^��H��	"��] u���J�i<�kRM$rbA�U�����0�Ө��Ĺ}&��Ui
.g�\7�)J��5����ݶ���>C`�Ѹw:�}5x�J�nfW�5�<�{p���;p`D6�J�4�rZp��f ��3����*�k@ ��?e<R���iOT�
Q�����h&�(���nii���T���/��Q�pl�Ӣƶ��˵�܁Ȯ��SM�S���Z����̢�Uɲ��j�pϯiE�a{�7��N�b'h��I�/�3T4D�9�4��ͼ���X�_���!��Y1��B��t8�u�?ݵ��
�s0��F�L3�pr���m��8rh͓�h����\�fs����L��n�W���)n�2�D�����8va;��yV����.���5H�,����Ϟ�" ������@�Ῑ�^�T�jZ��7����0��X�x��U�"]�'
<�!�&�N��2<Hs�x]~qf;�O���L>QqԲ�&��K���[Q`�4%���Yp �^�T_3pL�]e��/w�Cٺe�i�M���Px%IME����&b���܂G<��{;�����\�)R$`c�����Bb��V��92��^�#8'�Sgd��d�u�<�X%� �i�8~���2���8%�	��T�m@4~{Q�p���%����O���C�_�Fqx��3��]�+�S����4����6An���n`�2Uӹ4�J@��mmL<,�c���C)Ǐު�.?���=H9�f��[�c�� ������š3c'��F�P�p��UV.�Łx�f(Yw�bP�=7g��[y�j�ױ�:���rJf \������GJJ��(X��}�V�s��	��%�SЯ��a��l�y�S���\F�FM���Pd��]C�?\Zٻ2b$bͦf�<;��G��"�y?��Cw��B�8�?<A��SD�����<��쀩����魿�"��xsb� ��w�Aw���4�M!l.�N�o���D��������~����#��	��c����%�!�^�\bR��{A�i�$V���)k.~<0�\M�M3W>����mt�gV��Ig�ǲ������髋(�#�u����q'ҡ3X�s���EX�d��!��*��A�Hh�Yۋ!z��$y[[���l��$N��>���{P&�!=*\F{b��?��E]u��aXBĥ<�كփ�z�N٦Y X厒Ea��ň������.O]�p#�}1\�z�숼�d���/ bs}������f��H�>e�Xb��⻸ވ?i"�D��`��LV�QSy� �a��d�P����l��n���YE��.U�ҹ�5���ŀsY����D~�v�`= 	�DQ}�8,~�9�4}��L�؅��~��F[%�y�~�2�X1�S}m�5��ů� i�R=_��'0���L�����W��l��x�	N�F�-�]y��r���	����x��;��/�Ǿ����m���Ѻ��&��
��� �g���Z,\~_����86N+@� ���Z����V��;Տ�y:�р�i!]q���m\���0�^��u���)�K`BL�d J�7%�}��u>J���Ζ�֊Igod�Vް�%h�Y�e�"�38������G<��O�.�ͧR/RT�x��R�_��?�zm=� �4)k*һm���+ 	�3\]�4K�D� �a�L�`uչ6��w"���lD���3�	<J�^S,��s䥀�.���x�~`9���n��&��Գ֫+�},�Ox�
�d��E��2�mm�t�=IF�x�p�������v�#e�~�N4u|cdڼ&�ڠݾB1�K!��Z7�8���R�q�9�PP��1#�ݫLg�;R�O6|b�Mp��(�6����)��*�:ҽ"� A��2W�{��
�pJނ�#�U����M��x���z��Zz�@�������.�c
�:��O(]�
����޿/.�����]6
���w�v�!/���tt�Z���x���G�HN��-M����G���`������bnEE��T4*�EN��bh��jz��C}_�i#*F}��W�i��8���!չ6yS��/4�̮�	Tz/*�������tGk�7�m��V��S5 F����镊l��,yd�Y�	1�C�ښ7n��-s:�@��J1��~$�?B7��D�be1{�x9���Q:��[z�t���L�<�Ug����cNc�|~7ƭ�;fxl�"��H�8��8S�u*�⪖5_������ۊF��~x@���Hg�ƃ$��0�{�NT�6K�b��{��`�}���������&{��.�̽�(�IJW_�!�(�&�o��yHȏ@�����v���$�8�b��pѨ�t�l�Ɲ��ˣ��fgl�p�ݾ��
�#�׮@(vRq���ag�����=�F�OG����G��#�cz|Ln�ZR� ���()૝����T �J!�ּ��-Ӷ��O>W7���J��E�2_3����A�?����Z��_�S�i��_�_"S{�"����;���KC�Y*��b��ܵ��"�N���9j��$B!2tRV9T�L-�C��~���N��B�0F���]�Y&�ï:�/�BtF`r���i�pm�4�=��2�H
P'�5��̈�7�Y�"��Y�z�o�Ѯ�툹�����o�e��-�1�}p�T�p*v���`tڧ����)��A?���3B˾e��b���b��{�,�'ZE�Q�����%��$KVQ����?�WLS�K��$�|1ճL�X���{F:���P�R��S=�F��~GX�����uۓ��_J����Oe�0nD0|z`�o��FC��L�HA�ce-�V�D�p�h�<K�i�98���}-����c��̍vU��M��8�ɣ(.͢M� ����q7}��|�	p���-:|uTُ���L�6mv�&��5��c��R-k�m zn�I<���ȓ&�~| �ڢy��y�i�����˛K���t8�V�Z��L&\񦒟5�0d]�=>>K6[��:�	V}p��*Յ�L�c���z�7����&Y�!C�B$�u-�{y����#�̙����Rd�L�q�xƨ��x�^|��d#��U��Q2�9�b:}�	6���X�R߸�3�`�)z�<���_�x����<����7~0���9�:��W�W�]��3�M�@�e���2�V��0��(�KǚT�
�v�A5\I�]_��;e	W7O�*�!'k$y]l��g�;�v�J������,�M�mc�]���hl@�*E������{݄'k$�:N����R�
��VnE&�h��V�#�׺�>C���4\���zu>�µe$���(����dv���Q]6=&�����.
�f/�ea�ǌ>l��Z�O��\}8�"H.b�'�,���:WF��MՖ7�&���)�&���M�;q���Dp_p?2��d��0I�	�97��&���������&��Zx,��]u�/+绸&��UP� Z���J����c`(]��h���S^,Q{�s�b�p&�8�f�)�&S)O��$<�7���ߊ�Q�{��+�z>M&cb�a+�S�S�r�k�	�@��6[�Ю�:�R��7��+7}t�^��P�'�d�=l�d�����mPM�������g�����k��GQ�[Wn��Pl_��0��c1�?A��	_L,��2�d�f�!�[k	�C匎��b|�}��'�-ZJ�	�J���nw�Nk���9�#���n��:��|�4�K�����W�V�Yvjn����es��ϱ�[�����t.�g��e�ցT��;Kt�܃�y��Q����so~���]��ժ���s)�O��'����c��l;�6}O�(�Q��E�+ȹk���N�+���N�b·ks��*�5��=��Ȳ���{4��v'I]H*�>y��������d�=���{�l�I:���(�>뺺�Uz8�����^��иh(W����߃)0qj���%�Ϙ�eL�W`�o��NDd��~�u��d+��i����\�Y [�5 ��x	^G�E�N�X��. ��.����%Z:����R_�ܯ�n�觝��b�}uI<@���3U��vH��Ƹ�yX��F��r���}�Pו�&�`p՟����F��?�p�Ҭ�C˼�<��<��׮:��O(�ŋ9x�0>:
��Y�"�=E�)��?ha WICo�ȑ�x��*�c"��{�ب�y���T]L-��H��	Xы�(A8.��ٕ�J�6����g�<�+cV�|��L
���id�}��6\y��Y������b[���,Ct�P�N���]�km��<��Ւ�v0m]&D���� �@ȉ��G�mm��a*��T�Y��rkۗP�T�?����îߔ^�(7������cޚ�ֵ�ٓ<>i�d'�g֦i� ��en�+���h7"����ռxx��L��p�Y���2O��b0�zCm��!+�}<Y����C�_'����A~P�"m�%OA^w[t� �[����\y"�7�O�&戬~�h�|�t�s�4��Ңs��xgԙ�$f���К�I*�q}�_�w=,���v]����i'4i7�<�q``�X':_lM��5������P��5' ���^�-n���^4�:[<x���e�x�����3&�d�$35�ղ�`���Ӵ��7�?��7�BV9%
{q��[Km݇���e(��җ��@qt�j�]�ѽVl�z��$�V��:h9���z�N�lMgU�i���n�OLq��V\r�7�`1Q'���|�6\p��:$�j�+6j���C�^B�t�BW�mZ[����p��vc�>�k5S����I�kd�A�,���\��v/攎�% ��c���B %�.�삠��ƶ�t�+{����ͯ��y�V��|����j��&qsN\ed����U�aP����ǳ���{�1e���ݻz�����?Ï ��	�$.�N��5�Ѭ