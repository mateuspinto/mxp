`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
soBBE7wsixi4zPh/I/gWv0dIOkqie88R2iPXy1c6N31ZTDS8AzKMgamwyf2MgXN0+R9HTlbPUl8j
sc2RLBAV1nM4KyX93xa6hcoHI8LPohMW2YcwKPe9qDnr6cczQzdGe1FF/Cl/DPaNlnfLiYPp1CW6
pE7i7VQnrGkJlwepbWeYwLOlIzETn1502vhCl9gvIPokbqQF3j+iR7CM5SrQBV2cHbtSjCK1vW7R
LdbZ+xAAiXahaDZDSNOaJNKoG65l/FQxQHXHn3oLVZkGSUhK7QRYEsgxG3esrdQtM2vrV1hKK+jo
MHehG2NTq+UmiViG1aKDSwXgHyxWay6dvbHtY+KMXCJKsSz5/SNZpzPa2IQgEq4af0FZZQ6g8s7N
9+tRJbrKX/4KB/medMxa3eDKIx3bJC55c8f26IEgtD8dkPLoxvZh9SKkSEfdRN3vh/RfXy3xIAqc
uWqiomiEe9UKh2QTx/IdsYQ289gdC2LtPGqpFEBcZ8kB2OAP8URxR3CYk75weV1Uog65JmFdHTbj
RpO5bfL17dvHo8MOzhXlrxQrLuXxBqKSDE53n6Rb51LRPncsCJZs/myk1RADDQ/BjWzwRVpAz1Wp
eDQ9hlj1RXrnPf8OAtcaleI8rxiDmeen+5JDPWspsb5dSOSwBM6mjEOjmup2o21jDA8vlrtfND7g
3QOMU5lWMVJl7oATHcatBHKEOwAw+aUJ96VEhH8EqoJaBUKzHQN4YvnotW9fCvtKvBjOxrwOEZRj
I7TA0znMt6pt9deCw9SkM3ffW4FPXDEkqIiyXOoo+qRQOnvmKMxPir6l4RrPEt4X6Sz28ErVIwRW
zJfyeW08RYuPffniwDglv/dI7h7VUh0yIOrGOvbFs8+kUHhFp4B/BbSUAVCpO/+YDf4fkNVD+u+1
M3I2EVOCBR5VyGtl3GI9HY9Mp3ONr1Yk6iO503ixNmSQ0CIBC3mEDlsfflQkBbPzsRGr8WsXK/C5
5P9D9DUE+cY0s1QT0v1KfbUTEMBPDFWeCvcBejLBrigOPwNMY5ufDSQQ858V3nHELHKupx8JVwkQ
11t0MxUnAWn5cpcjMBaeUFqbMVqDyYdQQahaZL5GssqGna/eKbkhYvcDcxw7G5y/6ZiwNry1W467
qH0jRYSIwwp3mhlk+ar0tpRiTOrMbjZjj2J+i0AOlJSHhyH9fp6YckTf43mMxPF9300Rzo9LbRf8
TWgS+7CKZpjXLreKz0m1/es9kiJg8kRFw5t4iMJYl25BmvdebikQGIBoEH1kUuOypxBgJ3QKEv74
pqCykgSEZvnJNRqhXfpFPl4BILrpWh5Zg1RldkQqOARta7UOFTjE72kQhDLonjj3fhagIWlzshtV
YHPWUjkfpaOS/7Milh3RVlNgtLTo6mqUHNCzVzN3iN51vcNaU1zuGnJLMeanmm63HoAMVEpM7EPg
En2LGVLx+6ZlNwQzTv9q6sDZtwkKhCYYu26G5CG6SJI4uuaWG24188T+5cjKTNv9QtxsGAmURUlZ
YkrZa2vQpoJBAoHhjeiJVoZA4AyDrsYEkaeeZMqcXtFtBCOIKFM/syuqbZoXuoqmMJveCt+/oqYa
Lqfm9pZMmonzNblXI7ZL6ldg77Gb8Bt7CFUA/B1EzW9mixA19z4IHJqsXrc3hzy0o18P1JzpM7WY
AfBXbD+zI0wl4gpM1QUiCCwRpYXHuDSB9uMzY2/XpJGkI+on5I9gl7D4Rb1lAJSGHacmXZ5Ek3YI
BwOlHLA7XFR6CPkxDwOPlGPoP5RS9mF7nOVD8UvotWZJyu9cx9ZwJ4GZxdipFebi8x2NYrQBK+8U
alK8nWdacwNOs1OOz/cwfIgtJQzYjmAdfeev6yLlYaEvA5JCWr4ixGsnnDQD0yapcG2MNH9+hOHd
8eqXevHyEpVjEerEEFXrGMYlfnC7aWxNM76A3IiM7K3d8Cuyi1TScv3VXuWCVH7WA3f40Xl8jB6t
lsdmbDd28HmthXnbfXnq3dgKohNt5vh6LVgfElWgp6SWg/sWm/hsj/2cCsUwHB1/GqqFxFCFknyw
z3U1J8stJsJF8uEB0ZJ/f+hcL4GpVUOg3ww7cyqBwpX7a3TjeoxyJo9MvdCthmBXf4UXjGieu1RU
C5G0ihibMs2yThDBZZUddLpf6onu5y4olYC4jatHPETHcqNEgAS+IQR+hmVOrrGLoVXKaotkK/jf
6oUlMi3OtGGclFz9X+LvTEhH8TnGmHReGb6P6NP5jo4go880pAMfm6bNK2PWurS2et649SOM6n22
rlTzVHZTJVwGp3kxlhBXX9ydaLfuPUpC3e4Ag/dRDAjjruNB5Kwc33dbo1egDA1U1sj3u9puqnqI
NL95NRJiSb/fLb2Z8Q6/BgQBszJFdH2KgbjaZd/kmj0Pwj1q3YCdDdbutj8SNMSYjtIy417L0mcO
l7vt1o8/KaHdzR6aaiKzRjs/AUK1p8zkieP/UYJBJZWrKu1BLiab1FX7KiAzwb85dZ6mo0fuyBph
iJOX9A/szOz5I0cRaFopMXjYzC6JJLbOVtrzigtROo4C/NikH+82z7fsTlpRI4YxgzBS1NYeMIjA
pgkBjCHAwYIJK3IIdTI0fhjwGp7Z4LzYz9H/ph42AOz9CIf90c3gpiGQx/eICv/hP6+TFZNsDXCm
OWe84mdKaWF+ofuj3rtQ7NqCoOQSQNaOuUT6pdiNUg24pNQJjoCyeMRq9Pq6kfEfxOsLmLny3YcA
gYlgAsuP7BsdYRzc3XLzwJXE81W76OblcMSwfIXcuW2xSllYVL3vjr7YXFaACNMVhnAah98geF3V
nh2UI5KEOecyeKpTfGNVG2JlgKPsaKSYqk0wo9SAsQcpO8/tPEYMkj33W87a/0bj8VAWrPVE/q+M
pQ4O2UKTHwMNJH+8xy7xNOFKcFOVOAv0EDxkqiC5FtR/IbUoREhmk1atpDTpTsh2fy0EAGkajPlf
fQ4cLzgdwPxh4ufKBgZXHaBLfZVb05tKNzuCtKYPcXFL0DVSO1R0VQjgEgIWkum93xe2PTH8Ip7o
QsRr2VJA5uKxcgGGFkITxjeJaNVc2pJ2yPS+Lyv1IU2cu7Ox1fJwXuVJx4b5KnOzEK999nsXgPYW
SQd1n7sLD6u4cXVm/Z/rIho1DBkOre4Ntu2n9S/k4SlEOXbwLmanmx9YHkcjMgjZO9vSvif4bytS
Ws23nSFHrouXIMd9CmBVgndBZDu54RnIHdthO3oB1w924j9SrRsD2YOhpUXqaLgptUIdDMkrqvrN
rKog2uaxJrYe6VMWIsb1Xt2wuJFucZBgaOKcDVxfAjunDfc6kvm9drXk/X2JCMxpJveABS5ZCpO2
J02jMSQ1IaphBK0oydL96GbTKSrHaQsyh9laMNQaA8yTJ0qfKVD7q1LJjLUlBnTm7/JRrmjBM9C2
uRpO1m8wCJTYvEBShO93gBIxkri045Qb6gtTC8tz6vVjgLwbH9T5SfaV86ZJ9KC6/1Bqe0vF9BWY
FlwMMnd68WgACclNS7AEXAOqr/lO7HjiK4WPTneWnxc2S3RCSsnZw1Pu1YF03P2uF+dgxteonN7I
oCcztIRvAOm5bHho6ROumr35NIUjrpYDO3LDVWbJsqxwOmK3On1OTE8Br55zH0KYmJ6cX6mBWHJz
RK9HUGM4xlx4HMoBns1jbhhYYlbdC/6LL/2DdEGEubob3K4UM+b2AC02yzlIv/EGQNABD9OCPnzv
CQ2GuJn3rGGNK/9FTh9snjKdUcWQvWR2t6go0QOTgxZ+RPNU38hBK+sEkPVSf6YptbT5TJ5B+ACp
IIyNOwEKQwBeNwVQrkQMXmZQqtrkR0Xzldn+d0pPWDqVldQ/doIVdnj1H1C8J5B4nzbiYELLLxDo
yaLlbwYlMh5a3uWG6f7smHaYKmjrCoEIspRiAMGFGFA7i6DRP9Guy89e0Xkb+dtTjm+Uj5p7scRI
C2UPtqHK4fHm1pVA2vPEdNcNGFSMzjP7I3wkbGD8PN5wn4u20NgshcEUJnJJNRcvYGRdTOjEyZcU
00XSYUWSZopE1sKqayyCiWyhfV81bfk3nr2RgBnU+8Fotb8ZhO3bH3KNffy59RNFVl3nFG3Se5T5
fO2x+VQmXA1txxYbUjNH2QVCQKP5GxuNLTQ/OZw5NDhBNJ/e4oLKwKg4yRwmVL56zA4/WxHG1+9E
9qkTFK2DOFQumVtZs6eXHW0g2ZamZKXbbnrzA8gM7SdRZIkkByDfLB7PAjnm5x25Rc9BXOZH5Iqm
4Gxzcqhr1GBXc+EwG1a1kfx8FMmZvmuQpNEwadzDAsixjlGHNcL0C6dViLwAulqqvcjzywlxzdfW
k41eZYndMCJmhoJfWd9m58Qr+ZspWwUDzH272VDq8sYuYUG11lkQZP+x1OvSzENg+QeG6HpSAPE4
pomBesnVGvjUKsZI9ZsaIX314FFqUXr+fNi3sf5lltnXtvIF1KIRMLsSc6WQIwzxrcSDPSZOUNPQ
TPX/B+1GpAUgfT9ec2tU3HUmqaDaW5ifdl1GMx4TQ1E3JykiGA1hyLQgzI3Y+y2eXR6FCCZlHu4x
DBuHjkTd7S0HSZspJRchOoOtJ2ljdloMbNTP1IYLZelIIOq/bRbPwr/2BGt1Q0WitCojxwQwc2sF
vpAs7dI/grfeKybBAHOw68iMOewzlwk7ItUuD2Otos9SC7bGpkC8hutqO25v/Bs744a8sPhROYWD
83zF2T//W27B/xB27h+H3sW4ozBjBsacFKMmg1kLw0nT3rsFAS2NdiIib5SYiYABeVFBRJmSP2Wa
OtMUoVa+RvFPRGjmf6v9VWcbbpTUMHxZUIHEvIJvmrKnQHNy0ElxK7XQKk4G/veDuZITbsB06QVT
GuGq4V+HP6jZ4hRh2xNf1Gx++Fjcp9/Qu3bgRQhBgIfIKWg0xezFgEpVbrRMKhH+16uSSg8BmI+d
kCBqnt9lMbqGv4tTgp44aKbAXQ8QSAuAxFVFwwbUdliPquShro46DKh32NEbAlQlODpdEyGQ+js6
qGMZ9hYEd+1l0zWLfAHtP3g+IWy+DkIvZur4s5GdquDMCmMZAB7nPn6Bugimb265eoXiPD3FJXnX
zOE5RHtZ6ldCEl2oy010+VWzIGvgzX9m0jtc5eW8s/VyVZTFoadczIYDitZ3MGxiNUsxHN+uC0lG
pVOLv2oNRCPX1f2sfNGLKquzyrBF1DXBX4ZpNh2kIGegxEnK73Msst9epm4O1c6/Zm/K57auEF9J
Hpqx/i/8hegiENmyu+1DUzi8u0egoM2/0FNM0CeQS99lDpA6CFiLRHLJbgDI4Fe2ucKx9z9EATpG
jsIQfsDZMDAdkmjkwZxSdlXXoPMWtpZTOtn1SPsF2RVg9Ia5gID1nf/zS34/XrMh1gk6TPn2KVRp
/27CNuAK7KZnq1fQJzT4L6XG1O9dJ9jUBT4OnR+uMuYIIrlKYK7xGHqt4PtBssQPygN5+ZOSuMzT
BXguNB1QRP3gyfmedlmMym3Luzz1IAPrffO1b/mgdVJcmcQmNrR9WfEm+VvrcFDD+AN6pZji5CcS
Id4jscPv+WNrxGzAvZjxA/Iytn5mmQDRaZweNYN0BcCUL4DrlhAfAzamhI/Dahqn4osRlvTbHDto
ys7nGv0IH0/teNI0TA0UdsqdOKfR1m7wXq2/gfF67EPZbLnyN9W3gcPjiB4R2Mfr3xezRf4ypEq8
0y90aHKxVDlnVVZCONUSd/Ahl01PquIlbfdC5mqjqmcxeW8un6cgzc5oXtcjuDQCi+a2kxBSsvT6
/fx4gxl+ZR+mQEL3/UJiewi+N4ZH+Q4WEFHKKrTKBHpsgLo7o5YRizEUX4EfVTNd5UY7pjH1RSEJ
Xr3o8xFx1aoi9TLos0ZBxpny7U3Q9JurlQPydPjDdWyY2E0EAQyCncx5wKzgP+JyRv4GY4k3mjXo
dlTOt+fcB/LCr7QPMIFy2rChdzEm1e35tg5wxYPWCFvJNSD7ipYzMYW1KVFWP8RXI72Y23GtwDfA
urgtpibwhjFW90+bdwNS0dGAUGDjYQgDdPGHa59P3zenLjZT8veWYcUA7HgzeykZk8pd+Cx7QQTD
Uqd8pmQVOo0GsC5sZfK8pnvcRViyafkTjcs/VIpwvNZowD4sHEVkiCdbTmIitAJSK6ao0LLkLUOV
tfTeGWVKaDtYmU84PSwr8NX+EF7xvGNVxKYwQLjPC+a/iApgzTgJjH1K+ZMRSQ0gpZLBsJJjWJbY
P40CBLWrQyTRD4AaTv4UlLrL9SD6c1BqxdI332bE4hPesu2eZAWlWRiH3XJA4D+w8nNKdho+xhge
ElmBVr/Vf+PDv3zg8/JXm3+hd8yW8XFntpxtREeDPCm3QaTRDjTPhXkojq08z7SeTazmPHobcelH
91m/wNE8QCwZSZ0xYfsegMP+cG9COSrIPT5Rm3VABwKzbGckYzbrZHU6f9kCEDhWZOaXlvbSK7nB
dSnaKomrXAKbH0jS8dtXNdaDCXm7k6ogoMU7FLStOvbSZVeL8Wwi58RKkuJFt9Xu99S996VkqlhE
0p9Tf8CmiYBJVhVT6KL7J70yb6DjgnuYEYMtIQwdQoDUZ8YRRILBKq3qygWhTgDr/7BR2sAUWSE3
hxIXU4CFqRT8Tv79e9s8WjexlYRY9BY0k4jSLwMElKvI/AZ7B1lvhj2azH+g/rmDIiFB/13IvmmM
7QjY2gcPvIuXY2UOyQe2xV7p1VFLA9tzpBKcnDnJuEsVHWIsN+Zh1encIG8exYf1ESPCEv0t1TaP
pIfrVMvDPBgdfHjko5PWqgg5YeIMSl4Dbyks4H0csuSJwLTZaCiug6TtIv84Cgvk2Sv64VQW6qsz
9OOJZf9G0qL1CZ06vnUXVT8W8XNuHT+/lGkhu1+f1daJ0vrjBfQMHadfOjH7Qqv35mNSY90m3oOx
FPiF01fMxPz6gCrmxpuZvN3IocCqndWlSoU1W2FqJjgtKEsiUYxfv4/VI645gPiC0myTvEQQiIvr
pkRHyRVY0grpq4oubL2RGPBpl0hDa+JyC8xgvy2beoHDSNB6icTDAOqz1XNsqBq2b4UlGT9v8BlA
OKSsLpCMx9o/zMj5IwtGkmdAypA7L3HnXNRj1t+zYIn7qVIelTLXiq2hTIWJyfuhmrYqxh3EFzAE
gka2ormxdbD89jV0VkuUfjDXj16EOmD5iNLqlSHiF/iHuJAmWGm4UQa1pzTiiVgxQzqOWz0SWvWH
I/BXJCkVk53ZqUmFGu2+N4nRRbGWy5as5SdLemP+8n96xCoUYV7p9vFoQp7bLq9IADJ7Lsyjn3u/
7WxDIeK6XXijNC2xT7F0C6MEiXM1Fs83NauMJghBv7XX2tlHRXiRwNMP8KN5Z3j/dWU/9g1CzTA4
gj/787C7KE85uCqxM2UYxuAxamyc8Wx9fyGcw3KUjVhgqKAxWc/DQ1j8kI0f/KEqz8KpWaffZJDJ
XprZMxtpX0Aab5sFvaBqpRVKx8OyLAcqXmzMtllm2mNn9BewJJaFRcjD9zxbeoOMY8rS9Kc/Y3s2
nXQp7ov9DgHD/I/HPNb/J4QVRnMeClHU8RR6AHoZvuJltIuaPyy3dS/me1Rr5lga7AU2RspP/yuj
j2rxAYkGknDqxnbOIudkJgDR50ew9llLmWW0mtCfUciWODNbgeegBlbmTPZkTgFkSrdR6+FLQvpf
B8OHUPqG4NChxF6mH33Vro+4z4r0z5S+wt1fU0cKDwZS/uLQdjVW3mwkXysmuj2iAi5Th6gNFGD4
1VC5pUUcIjqFhaOA4dZbmZI1hV0oTwP3ZWtC/LO7inJAKCR5/4Ew6HsXsco17/gCgcX3X4kz5URz
CFI9m8TQVIG1/6fxXfU21SS1msr9X3K3CI/i+dZOiU2UOuFbjcV6WeClfEhGvEBvy6cAK5NSRbnv
b+BXvnggfyPXqFG94OdBBDNl3T7OOQej/GhStq2sTufqiSn0Q7pu5mPJ/p6uNu2TzD1yNb6K9WpX
k8W8WFDG/AyqPQ+rOx1D822e3VPFfPQvW2+JgTeJvrB3GO5csyzztaltTtQpoN/AKnGh7X3Bm5Lu
z71xBSwV6RTHcK2U6xuKy6VCu5Z6GWy+3+gXHR0eF/jLDPinq8xSW8Npwtr9kl25R0WpOz3XnpGN
JUk7fzUkIHXk2RKSjOoOrswjgemOjyl8e1UshNnTLOtK78DQq2Y1nofHkEDsCHk/uz8LzExjKu8P
jy8k1NypHTH/n/qnr/VIRIQQFODho5pu/DON5ju9MrzlF+U9uYWaunRuXnkFC915PO5TsBjNJZxp
IovpxRNwxbyUoO8PUZyPBLnLUUewEdIC25hji10nj5cxh/D5iad2xYvBy52w7oT2fqSk672Gk9GN
5xpmgW9spf6m860+qseJ8afeW8nMc3B5jFclswscfkzFf7u6KfnZtIpbCuWJYArKdpDJBQbtwEdA
AP9ib/TaNpR4b7hoiu42QBLMijCRFsnIcHcvscYyiJvf/u3uA75FPW2OOFqKn+y32yxBY7XGFOyM
a4tEICtJbWM4o63TmOl+HssCz50bXteuB6qKjuUEVQR64mlVvutf4j35kwY+z8p0Zo4hL1RWGkRQ
w/b50Gvf4IEcO51PEPM47iRrBFOqiuk+ecHn9JJPFj986YQEVowxVs3NlP3EVTcb56MQM7vALE1i
Eewdghpbssbaqnpd37unmAXVau/fUVeFZln49PSUpyW5Bsc5h8OSujV8YGTcaadPGO36T7RkyFQ2
m2JAgcPOABOaiPJdwQiBGMsa0Hz+123T+I4qqvovoHL83keDbEFaDsUvdcFYPa9cuVmZRyqZiclG
bP+T86SuUXL2AqnJmQPpQ+PiaFhAF575cm7EKd0uCfs8vNoW7jfAD2+oO3VBArQfn2WR4NNSz422
i8M5fuutQKyAjlPeHbCsj1fJ6qp/N2pkfVxjjicNZbEuSC0bQNmLSIK3hfLPqGNcH5G0sMAUQC9/
c/1MxQRudl0WEDug1R2szTn4CtN2D6MbRE+A3qfzSJ5Aw4MZ5KOCTqs4MAwpkuJfkSU3gCJgHn9l
mFhThlvX1F1E4yfQ2dhAxqVxwNAWCO4+LrmKxUdUEy/Pf+I8C+mb0DvqlTbdMRSY02BZEDoN7YmH
EVf9OCNJULqpQ3D/2H1A+LwuGsuTgZ9YDVQm5jJazwT3Y+Ow7gGiUcV2+xD8ijyxj4xrzOjSSUJS
zFINz3tq8VT+0mVFYU+zbGlXt/NYxATN2+F9LgivpKUn+WWx2IVfmHj1y2ZOMIXDVCj0MegwImvk
FHkw7O+2zuvubAUrQ4FC53mronb0G/JjrzKvHNKpd8/PD9RrRTOF73tJglNLWBJxYAUoSWH3pSmW
KlBuWDkbPON7ZEmHwuwMEmjTg6XWNXHJIM2pl517dwxBHBz2hVD+AXaKRCh3oBCCkodF6/6tOhfE
Lh3LHXfZ49V09srtxKnZEsUDCsXU/usd4lu0rBHOqSIx9N138n1hwoLRWMucybb6Vs1foeT9IP69
6Yum4gZyxILdIggThmSghRAh35r05gyMk5DbgDtApNUjqCNzCTfc3FwmAbOxx9ExHtvxxbqplkzi
ZnR2aV0tK+hQfycmk8GFQMY/mpM1MYyyPk5qwJAvBC0yDcENN1qJjiCW7ngDNpMtp7aDXNFg0caK
ALqWB8+acw6dweGwhFewVCctjp2B1MoLgutjb5MiFFe7izHVcA0qFKfWQ/+QlQbqUUY0s0C/RcKK
81qax1FIiK9YGulxMWuytfo1pHfw+BO/qnIaj41kQQKZXa1CwlJ9KJr43fAe0SmfRYOx1zQB55mJ
xfMl7CD/u7M+NzUWNWiXoCrENj1CyMOFmu9NRLoULXuaIlcAzwJoFJS9YiW/cxmXiWh24FSUQV1Z
SPwE+6j9KdoXaHTpY4IPJcnxDna3GePGlc+qrc1xX73gekrBys23hTTftwZe7cwm3a1Kb0Qlmqfc
Q4zq4Hc0t2ix+H4LvTLz53PPJd0OTfoLkyT+lXsY2MsSsiODpcD+ZmD5SCwaun1Uh86S83fbPqxR
enyJcpFsWYaJZa2QlY/EkCS+5yG5CiWURrJuEE9+Y1NhZES/a+5e9Kb2AfARDG77kaZB19e4U/lN
Jha3gexB+Ob6EsqmUZ0heK7GBJE1Bp0MGH71bPaGCvZWBfcJAydlEKl6I4W72X+EXK8ttOSwQfzr
MjR0OD3AP5N40d7/ZN96g641R4gOLE0VOhczCvY2W5o1XjAAbc2FOZX2xRztQ4C384nR2kt2jMCy
FPxeUR1QUPTTdcpGDEy0MT6pVN9SBvuIp/NZIaiBFpTu+t0qUGj4wUOuP/rSOe8EU24ywv5b1gef
bXyiPMyckuNR9WA1tSA095T1KZZUvY88RH6/bj8iYKDcjilNhbiCubz3V5GSb2KriJRec2UKdzgc
xGBvCUu0p81/7KhgadV64eJSZ9dqP3zB8CPRhJgVnN6vsbU9kgsB9fPJJanskzIwCAS3wlgN0ht7
a+z9HrrD3Y28DUwLXeKNLeWTjqouQj3JOXM3HVVx3cHSmQA928oPzauWOE+5n5lvXnQLhfAymUfE
/yhesqlzPtBe53WXFEQKob2daKK3mFy2SlISQldjN7CM95KnQoNK7ojQaZkkVgyLGdDHF+eSOJDT
7SlbhsAIMtdr/x/Cez31YOHHH0f00j4Nrt52zViGfm6iXl3hdmoZnSCqd7IAlUnoHhJpKgbvcdQ+
nO2lc0CHajMDFrSHdo/QVZaqPVxqugHTPzPSmnwquRIjGbzL3EOhzUsOir3LO8DonmW3BaAyRVSf
ia3sYyREN/FO25ZEvJ962oZ6x/eDdyq4FGjDgetLgSVu/IYug48zcavWGFnzbPfzgXpD3leenscz
DRj7kzcYOkBvtZspgIYAdhP2IIpVBjxcV6xrTBB21idCcG15Fhiko0oiampt0xaWlFldRVmYTmZJ
Ivd92HXiXPDnFijYCixw1JzVDP7009kz6gq2g1KqEe5AEpMDLUUoh+qPGVOijq2L//8xI5q8+9T2
SirrxPzJWuCxa5miDS46jcpqMr5+AUZZoys9vYR8uSFxLdVYf4OAss8MoaLm1RXySJoDDp+r6MsA
7EpRbaU2NDsJ6USD4UAGcR+rYa75kH4FdADokgQdrkcqv7kCHIDhXItEmJapAV8BrcsfzLRtobhh
UdssBxcO7YHmtvLWjhj9/7seHqdN6rC4eymhH3TB2Opfh1VOVtBCcJNeLOum9RE+OKNNISoZ8KOg
/shH+lIEgir9u75HUg/9x7CY7piHKYoCML8dwSnaNawfkCD6suyhl7rIUDaWzk/nLUIEGyVU51Rp
PwOT2CH1aSNK2oWql67y2VchoNKnK5eNrPxG0+tgQT2Nfka/TO6cAvrduSKftW+VmfFcLPC1yIBO
UpA9e1dChZydi0IkIs41tE95s72uuNJ7tPIHOUZszsenA0QT7Y6UwamB0vwVwuna7T82lmZ6NJnx
sCOmKPfBUt/m0guubu/HqQQkrBxlIdGbUn9GKW2FarO4EMABv08beRwU3QYK5O63Nv97svpNBtGh
Fx+Fuk5ShVwlEhTkK+mXeVPVX67hrfshUvQDlx3Gs3Rsh7TzSULIBV0jXxi44S9zA2IVTd1CqYVl
PV9lWLKoeksI0CEerXZt5hRR1VhFLphVwLH1HyZ5t9x2/YXLy4hJwTgb6MUrnmlTa6ZxhcwdZlGG
taU/OGQd+rp9N9JUB5BnM86yk1T1CDVSXFigCA1iT13TY98ew9xpKpnrieKFQ2hBXao1dUPF40EF
bypuuxMbONT5Pz4cMzGBX7Ma/fORlWTakDAHm04PuMhXHqlehOBdL3fJj65kWAkIufNIXEnJuM/P
vr94KZY1pvTDas0wD4svCY3cDR3fufGlc7Sz1/YmRLa0UWQtUU/A+zrpwTiOTvkzXowRN/dc6j0x
ssOvLz7fUntMNZ5Uu+RaVB8AP5wX4hZHsP5GPbEWPER5QkCxYiHtOJYSV6Fh2EZrBMVmB2kue0U2
2Zat8sJk7Y27qyKrfuKFmnnTdxIq5vNXhsoAmD/B/vGnUE+zrfX0+c/CTYqsTXxk5qss9ehWa9Fj
vEZDrB8g8bInYuEYchAvLmTW7wQAIUYljBbk0l/Yc3ZXVdszGZ3Ai0KLXukHFvq0Zsz/cBqyeJF/
DBRRp1PB47kA4x0H8gx9+8VmSVXL2HFiXoRp7sZcdAVetRH0uywc5ylrUpF7hhhaWhFOByiqAApy
nPsppj2QMS71hW8CxqjcXQ/sq8jcLSVbfcbX00hsIXONCGJtU3nPLq+pDe0zSkQLIA0IEYIQQbsl
FS30hvfkbp5a2l3n0NosWgemmmhVw+YZc28+I3b/xvJWCAlcdZv5/loeBLnQzYhy5GQiXsHbPtgD
E8Ywj5cksTFw48R4jWDp9/YnfWvVF1bnyxZu3XJiIpEGSZpIkmgxwXy6k91JdTxTm7aHhqNpVCiH
gCvkhMFQEwF7cVH+foubMkbMDHXKn1SXB0m/P5vEQ7w9kfmPU9TOZcwOYx26211Da6XxwZDsPnnz
h426dIS4ksDHp1E736qBn4tdwN/Omfi4iOYQkT4db9hCBvbmWRmEn05YJ7vsBczOy6tLQYtbJf3v
/U0qwn7Myzh8fEvSw067rGm+3BW3xDxDxcMhBYgmBqvMwkMJ+J+7W2Nte05wcG9vH3ov9d+cRvFF
BCsTAlJ7LeAhlN9D0jfjbES4b2PGYauNHVvRFLWeBKIOrsPoRGeGPXHuME9q7iA6x4uZsfWDaZ4k
pIDzhMwzFuy+XWlAD5vkbbX+6YTEkv5FrHh3d2jxrrTRJWQLeCdldQnct0BuNReRKWHYJkiWlwjV
bd6E5yB9xQgVYPxmYH9ffO6jhoMd5TIGQNvlh/90ZYA70GgvRB2lvHe8A6J0a/XOH/zKT2m8ujQl
2bnsREEIhq7L1at7RRGfi5UtWk4gpfzWvXKDyJMy6nUOwpjz9qokNngBcKiHTY4ewZeYf8v1qkdJ
+UuYV0sRoYvYdS3fnI1C0K7M/K93fMUY7JW/FnZ9GHiUjdQpREwKfVV8Eih4eIXlncvz/NuEqF4t
o/Wk9LSrM3s610Ud2xfe1R8NazpysVFdluu3amjruqIaVEpfDpC7WuvcEu0VV23m5AjBAzLgNTyw
5+0gTQQF9vdfH8MbmvEmF4ZzGt7E5iksj5ARaFc9hvuTT/JTr7k7MYY84EOIMRVSt5sjMwfkUTG0
aI2rj5rH69zfWKZQqwCA8mPTbd9Yz6pCxXp+/M5+o+mwpXdqZWKxbWguplbPrL+VkOXgSPzS3Rew
mOmE9E9VFpD7kQ74tCIMrJINzsu6SeEn6P/XI2PlT70qK/1nFj3KLaUs1Tvjc81kS4AfHcweinN3
pNJ2e8bFEY9v1SelzHkeRCr2MlYqv/2Ij58XDBf4sm+tfa8/d5lsFjDw/V7N3e18Mfg05MX/Bcx2
Q+NO+TEAr4nmC7EvCJ8gqxfVwW+n8nkeiE6y4oBQbhCaioOI4RQKUauAKTJvotZvmtyoQg/qCUUp
lfadT8/BlUp3/EoI2VlXCzmN9k/aVouXwqnvuv0LpHW2SKwJDE/DUTXbHiq7qP+wJ9GQiHVDva0H
omfFQwyrSMFuwoxj3isLbV9o6G1QC9K7AoGV+oBd0IlumIYGZ9xLoYpdVEzdemVsk1sDrP+017Lm
hNC/1OmZKhmSEQ3MFdUOGEWRwhrr44Ti0hKszqWNLi4QqlaVPAFQ7GqI/rA1SSmWA392LTV0AgRC
rrMRDyldWAoBhXnjGwhi9FRg+exXMsSD/P5LNkldwO0UNtI7QxJm+boqLEdfuuYUFc+WfkJu7SX1
1ANH7qAXe/vPxK9Ld/9C95vL4Nk9AvE7YB7PM94U160H64tHbhc0Mplns1kPSjvh7+X23Hdk9aEB
pzTl+zuOcpniTTRzTRsWu4Hzl9GrlqRNk9D6NrpvlVi8OGlmUivdb04qoat1MFDJZMhAPxf7p3g7
xHWYqRqjrbrzsC+HxTiMKOS1bB/re8TzJi/kBEGTDIX99uT5yKBwH6Hz35aHkntj5Nusfiri1vOK
DiY6nqPWqncKjCfqPHuPq3i4zPoODRrVizsIeIqG12hdWVZxJD//7njOsr7XDs3XwIaP+MTBktcj
JfL3VD1UW+6hjfIAI2JZ0B0MxC2JOttI3rEH282FQZ3rZNvR4IFha0RNfB0xm36LYrG+6yrbw34S
tmNDVpzvbvul8jQ1tds4415NYF1qNKyxrRGXE6zUATwFHHKbCyY3F0cOsp77hAzqBb8nb9wyY7OF
5uyIka4NiO7kfD6wX6gONTBOFbnRSW+rzZsD0JYibbEPmQHCLpdy2leQHOBif/HIbaCL/4DPcrTx
TfZSkTq8880RrflMPTN0rkJL0cfgM+1XYRIs7Ovj9Tr5Nasx8CMJF6srX7FRui7OhLLE1f35pGe8
MA6SwDYC/i5p04c0TEsUXI4Bn6NJinXHzmWJbMkiRME5+QymkCiOlr7ovCdO1hfjSIG/sZpS9+Tp
IYKVCh0twQasiCkC2mep5go3WEPOtv32Y1rIQIii9v8l8LmObQJmklSnweUNdZDPHzKBsgLBAfjh
sDrxlk0NS+NdIbbv2kZZe4M2MAzrzJlqAi9x2TAxCgj1OMC7PJIbYHdFJlR7Mep10pjxCimHw9Om
QwlgLbbcc071thg8wHf1PkySE9IM31eoAfe0LQFYM+BCl7Z1ZlSZ1bWzglrbINuAlCGHGBuak5PG
ka6X0/f+/Cg1pjXTcHypl7pbTvCGy/6FZHu1wiODgHSz/MN92jsPEbcuwVgJUiZ358LjbduFevnX
YUFoExiVykr0uFyg1elGU8e4hH+IxlQjsG9UgSNJG8NuGOmVJpUu9W6bLiEFOruQc9C9oGx0zvCK
JF+J7+6GLrv47yt1p17v1UR7EMKo1rxTpc0LZuxA6013d9l4DFGdpJgV3j2B7ROLhpfrnm0IQ8b/
Y/2o9MMYRFIXz16pZ1cv064cg2GUcluI5HxeW5ZfUmDV1OB9/K0rCEl1GKA0OT6XeEKw5VJwlcGx
nsuXnt24MRgNEqL95tbvtxSmag9JCY8+iwwVYLj5KWigOTdxABkOBqPZT6uc75XgTMjth2hm1BQf
+sZpkS7JNooLXRDgjQsL5i06wUt9SvtjdALyINFIR82gfITbJ2d3/MJAsjo6jyUMipuiurVTR4pH
45f7Zz2tKP0HiagTRkDK9ACTSIs/7xCOpc6Ynt4J3y18em5Qw9vVKVDpqERrlBgaONI2MMM+IeRZ
I/Zwkt+qtVoixL4L1E3uj1HXrDlWv4ASVXIi9DS1/a/Mv25kClF0lFIsVkbgJbj8fx01vgGr46Yj
wRsrQwt1sqVkH+p1vDvB1GH0mzvcAOCCmGUgG253DU2Sz5kgvfxgbzQju8K7hKPiGZeMhOQeLhfh
L4j3rREihyLDr5sX4wNSbn/wPyn8U4nKlHmerMa87kusREiplwwz73oqbsqGggUGpeC4KH7+tuFf
YFLuvJVRf6DJWP61eDdIgW2ib7VxhCthCPSx+NRwSY1cjuiZFpJBfHz9HHIidywM5J6BQ0Q2U/XQ
VE5kcQCuJmQPqn20KCLPFaAT2y6J/1luJoH8swA4nFVfyGJpYnxgmdXYzmzNxm29qF70ruMmAiJh
teRtXuqwgn0tVmR0F8W5IFK+l2ylWymJ09c/TOA1O3wCdkjvhSMuw4Dq9w/5zIcUFEZjzViPIpjU
6usJ9cuPKVBtB04jBunaGl78hGFh68cI+VqbZobI2e2d3zRiD5Ex9fa2A3mYuk2Tslt468e6g+5u
aNiEhd3xWUmEskw48wmwzwDXqduqEZetT22OSl+SiKEbsweCH48RSaAMeXWLxGZ8G5L9BdGfeV2+
24GVOuo6rapFh1sEja4SEICqqj8N6bD3tKSNI6AFlQk5/OV6TSTp7ywdqpItVuqkcBaiGorJT8es
mjDb2DkqCoLanxXQ85gEj4gZlNxNSrssffjEwkni6O0PbaVdelB71cTTXDZ5tMnoWtUm6QUY2eWC
SDABROX8e94ebfC/R5VouAuyxABhHq37ZATzoBoeWXhu+rYeOfKOB1xjWNO6LWcYsqQ+GVANhe5t
SsY/NpmQqMKxrF2/YYhx273CQJebbmPp1BSsPIpNoZIeZI4tAnkKeREoZbW+s60G8znOF5iIcIUi
Di+Uh7TM40EZfruMxkv65E3ob4tYgIWDNqVb0xcek4mHAXzB2dJ6ELP2COIWJ/ehr2qVVU6syuil
KlvqzKEJbvrNEpKXBU1hk9eAri9osVrVVIoQGyQv7a4RmFPqPE725eFQRzrIDeXlIgrw+hhtYx+c
n8Wl9+yxmwkcgrY4LmbcDLor+vtQGLKlW8F6VGBJGU1rxbQyRqEIMGXTxiK82YLbxlgfS6uolw6u
obKryZcWH7Sz2Io9uXxG4/xhQ6MfGPbnZ/VyRXtZrwr6Ab2VOCsolkatm84yDiTwfU+HQ/q96qnB
kF/E2+oFzWKewkR8G2crb8d7MgWtvVUn4IlmOrp7Q7e1fFE+TOfi+Qe5P7Rb9H9M57tfIyseLYrw
SEV2oZW+kflOziiuU23rBQwtn8Nug5ur6tNkFj49CPEuN9/v6sNfe3sNMzCVit7fNuhxa9YhB8zO
NhvEwOTPaf3somyWHw5RWAZbHdgCy0N0KWtVtWbqrpoWjZjK5LUI+N2ezlbezxd6QDP2glKSgaMX
wLG/SpP92zK922HqoiwZRmQgTgqdZQE6086WbykXqtrQwoDgoj0GT34aC5a1or0neDwb3GWzdktf
7USMeXK2SXl3qMsIIrcd3vxBv3g1+tiSPU34AzbtZ9tiWX/VHWdyCuc2NW2d/u4gXblf6xSEIk/l
kHFHpGVHvkXaDS/OnoHcttk3364d8mGueOHQhE+5IYUtdOQh0urqUXXJjAbOup0uUqMSyIdqXWTy
oWcD3tv241mfQMHvU6DV1rURuItuJC3O6ChHEjKsOuzf7JGO6l9OajN1WW2Vh5FC8pZrIp74KJ1i
WpRLKJjiW9ufT1FPtsp+hCNIaYDsvkhpCSfBMLn4cV6qp8KWan23wMfLMgaNSVAW2aZuHzklZTmj
sBaLMH9hSLn5HgJ8WHcGSedUtSVsk5scocEoSwhef51aWEenAUi2ncqY6C3cgiUzbfm5qew+okpl
I52jvr0SePRSguE/BCPCeGlTDpH75eCSPoJnAqm1KF5sL6GuaqedmSD1EwkTHBySG9nm2o9dnCH1
KDyU26vmOZA6h6DJKb7hzJ03DWj0gpfgq3fxcOcjsxt61kohHBaokskxXMTdbgR+pts2ZPJMcSu9
mw4mjQj6/RbHG8mmqxDtSGBGvge2RlW/i8I8nHd9sYav0Rl5Bg7xYeKqtHMGxJ0DIdeO/i3RwQ74
+lImzzcZU10/5DBIJZFTMTM73+qaEf9TfafGPL0oumy4iop9wwTRS3hYR6tb/EZkYigl+Ky+rI3+
XjSCT5GsA3ZbLC6RtXZvygBOSl0xJzvKvXMH/JTny3RNVxXXaHgQWPSKEq61emabRfQjnSEF0Hxa
clRNBnACsTZZ+wRjuYWQbdAr0LQYI6UjHxZonA6zUC3bpalPNVDZbGZTtgYZqlZNijoCUgFF4dqW
NAk0Bz7ena+YmA6cYjxkP50hPbGKjyRKKOWMDXVFERQ3wfWNgDua+Q1FuseThcCiDY+RDSnYFrD+
8MIMzp0BnfHCo14DyB5Ebv4VM4xwIFx/AK+AYf1814QQ1e8GYUhvkc0hTv27FXpVtYsh5yvtwfce
g646DjxhnFSthgh55Sahjh3NscEeX2u2L4z0rVpDT9BvR3lplOJoUxp/NwQX0uC0Qfwl73IAb0YK
lmA6m9Df71qBlhG8tZyoybmXOfQ6Mj/dKQY7rDCux4XgoWwN8WHHSB1cSV4C2/mrhbA1TniSLqAM
NG2zKCnH3Rlawff7MXawm2l4AMvOQJ3ySCGxk2IZ01q5tUFZ2F+Sqdxh5YL07j50XiPz4Lrw4zUk
zYwuokaPhPV4AbB+viIsECGBGfjI/AW4NCMlLa2K0ucice/TBSRAS4j8buJpYxnOTgVjd7lKaIPX
uycCmN2EUQR9GsIP2kdle2ni0Qn/CfUmqHQQvCT5tNjarY5u8EPQOwteu2B54BjSrRzzaMK5WZah
30rOgtLuifgnsjh4tRsnjawGu+LEFEfv8NZF8DYNNL0wR222xVCr3BxS9C4eiSM+QRS8OGgX6M3z
G0wbaFXZX6dCvyFu7tfES/c6vYG2MBlcm4oUnPyIhfjuFHAgxOlFCC6HEZglZq6VF/Fj+NGMkvEI
7/TMdAvZItEbMSq1iragCP39bFFuUGmLuJnfK/G5f2OED50QOe+Qt1srr9RJLdOhZKAU/3rjbza5
jYoqk/k0N04sGj8RPQL5UDLH1xBMaDVDP9cdUw7+eaCXsJpjIEqe5OJQedmoHl6XGhVXc89QZnLc
2L3YcRnwDLe44rE9c0XY/RQRjZVEy8upMPqw9L7elAkH7pAAKsDgWtw8cVD9yo3rXfhO+0r/VR0+
/EZdALASp7NBzYYl4g9tlNahOzNZpt5cxYYipQ89pnHxD0fOh/jlxCwH7yUt8QjeBZgJDHaPhXk7
svVPZhAVUPx+bi2tS2WVOooLWaQm21vpL+WFjlMwSluE9UgWyjMAI8jd0ukKed0ZaH5snqdNHhlv
FhlZH/WBLORc5/Pz7CTl3PgMDZscM4rW4rCUanyzAX4xMzYlBcLt9Akkk4bqNlUfshbquZxuEbhw
AKM4j/qLe1qsWOfgDcJr7G1kVt937+UFgqp/8euQKT4OfWACZFeiKxtEGs+YQOMmxVg2zCOCVhUK
W+lquy7MH/tmkcgGPVjQUwYEbmt/qD0+xeLCKhVfKOxKM71zgicjWqSHT0gTAORTwozQtcqh2Y+p
UKoCgZkkrMj73Jm59gGPdQA54/lSdWTLIR223aMZUfMg4y8JE5f///oPYLQ7BMezJ+ChNJ0A1ZmR
33YQRVXxY4CnMw8hW+xiEGekNyXSGIm2vDn02s5KoXNBYeFidj/fsRbLmHnNmcw3p4Ct/1CDVv0K
v0lsYWm2558cADw0zP+ETMBs4S7TfoFyRMN3sC5Ymyl+6hVabHzcIGEE2POKyDcLZWw5WpRWRQPp
ltnMFk60vPfVOwEspcPmd5PitaHhJ7/Jyjrj/Me1fmL8C9BfzZjYU/RM3nKK/vyp1xPk6VVxDIE0
o8d8PvbJJpmSWftV3yn62DdqYSkCQ6vS2wvtHSnYpzEYJxjRLJpw7pfUsKYuprh5X3GS89Uth3im
fHdLW6tm/BLIqd/MdPSaZjMkIIGeMn47MusPVX/vVfCCYLRlqD2eqwcqxpWCkuGk57KM7lL9rXzM
9tkN3rkqX5O/JDJuEDYY/EswYTKNu7AWYLPJPJ6zHUYCRXpD/iJD3C0RofSXK8+577fd+f2DIdob
H8Dedk5N5g/CaTgDW7Xu+LkiX3jDouU7dTgJD2fUKKeDTrbNpCGYbAVDwXARXflGV+XQpva4ogiz
IEKfWUVjPzbS4NxOotPb5o1r1mj1710BM+SgSHQHYgiLRAw9D81WKi7WEqYm/dfvd4DTPFayHgDG
vGEUalrhOFoWD/DF32d58MuUbwgjVlEphQaULc6xce8czjzMHRuAkxKHubyZgopm2xC4cod9muUe
vL4sTYhvDrU/UEVXy+MfKJ2JUe+jrUHhTiglLXJm6lLYl1foqZ4rKYnXIONK1YuI+GIYOV+nm1/E
4+r7PZkkFMgKOxxzeFFJ+j235PCCgPibVISnhevp80w1yHwqNqt1N33y4WHEhv4MFfix3Rnk+G2d
03nL+66ZM4Jy0SQJ6zUkakl3sYqZyz66cj7NedVaM/viENw=
`protect end_protected
