`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
b4rlueON2ifxN6m+LYz/MELu3hp2W3E67rTm82KSBw1VCs5NcwSWMMSaMcXfbCl5H836YLXMVv7T
HBpZXuokndDCBjRSjpTHj3iEnYfDcHf+CqiHj0cQXovazprQIB4oMWmaj3X9U7f4zxOvZNm2Jw5E
zt9PVJ9Al3ImkqYI2BMS8dVYBQGYEuDpzAdjivD6xKPYhm2ofK+ZuccjFA4EFjYAIaWykQqJOkhu
YXCqgdI30Dr1qrYan5rAteGUoYaQnXmwrBCraI7XzUwq6lgkjTApBBE4he8TmR28VkE/GdGPzaKp
MSh653MtVZdwpSPMfOzcOcJ0gT3n46IgO/hXsA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="OeJrprTHc6QbsipkKraSqa6XNDw/ZJVZz2d68vYLbFI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12736)
`protect data_block
Uq7IY6x8PEDYeq1JDCfFeaNbLbY7AIl+2zJju5J+ofu8c9bKxN7K6NhZs5WSN2lXUd+vm2leiwdv
BrpPvV8eRNCmlXXyb5U9P0BtaI4358fRaoFfNOGrZONV6jSKBDk1C9u+xLTsg3WdnWEujkH+tOc/
hPJxHfp5qPtcSKadE64ZR44wV8bFpkQF5QkpeeuO0QK3G7JYiQbM5oZIzbaLRIuiBSDflxrPB/OS
ScIwZoQ64r6QdKQO9xYvX/fYh9h9nn86DwHNNBd5smuYiYGWXUuOS3moadZQj7U7nG4NeT3OmIO/
OBzqBzCAiwa5LwTlUInmBPONDVKoAw9zneBPvZIXIkP3ns7/j9SNv8CfCrpy/lBZ5fLevW3vKh9d
I/nuh64D+jUescmHskxhg7ey6ys5b4zJgciwFVGIvXUVGTbfCYx+m1L0t/ucf/q+OIB1/CMkoNiT
bBnhIJ1GxqcnVDzpeEI0qVBlb1ZNwzE/AAY38rQL8+FhRFqgFLHJbjpi/uD0oJ9+m1FZvC0x7qSy
yylpthhqfgoT7w60qnUh2sWqGEMvPHgu+R0i/Sc82Obdj9ZMog/b+pYz6HyuLyjlXnbT5NI70cWZ
yTyZ4kswZwHlWpbEz8YXvtZevZ/02S2lTqlgRG53zt9McNaVZ3iqjRJXEKv3viSkdy/WXbdC+Yxp
vOEmys4M9XAisnOjdl+PGYdSs8GJHmq+bC2qldqEbz8gTSt1BcN8MSzuLH+e1MmQ7AhTQ8eeWsLK
8U2fTrWd1izDalczgPtIh4ke0BIV5Wy0DtBdDfqAX/g7Rkrw780Dh6Jh/Uxyy+37ZhiueUGlUzOY
oci1ooOJbStZHzQb4wp+tpgtn/3QHbhuPZuwahcHP886uanNAwoVxVrzKJ0pk4jQhV1z7CIISXDl
HyKaMZyzm9P9pCNEJx5RO9vVVesLloyWU9s8eFG++vRuhLPwtyMGw/lr6WuNX0oscxSti6mYRlUc
ZAqSodcgbYP7m1jW31M7qagUXuZ57OlaDsKRa3yDWsKFWldcPc9K0WqQ6tc9UNFOl+Yr4Nx4WHGT
MfxUwR3mXYXWOBbzI7PSOWD1HmfSeOHs+YwSbJ8pz27zrBoxCaTAG0pd+WY/lOjw96tnoLQhZ+cU
g4Y9gYo5gF+BysGMZKYuSx0FWot/nCyBREGsrLkeKR60F3SaZGC5S9FCo61qutHhBCQ1QqdTBQEA
yoJ4iaYgygdngFVgr/GAKmSiINqTVXsk/s1ZMcRJ1ovufeWeNrUESQTxNIpvqm7hBe60BQpi9DYK
2h8pnQROORFKTRtO735TTVJKFPjebjBiu2eVY8wrOyEsdHVKpCBY1lR5t1T0olXJ0ETGT/HePVIA
Fnvssu74kor5E1p9hPGiyNcTvgLLt2VAiJWZdHI9jnfbuazjxYQJXf0gMl3lndhWgpuofrqGrmIx
aRkSvH2MsoCyy0uIc+mnpLTgzzznJdk5okTzI8lHwl5q/xQNeNze0tOz4qXXGNP0xgKLXMa+5ZHS
o4QpG3cegHtefUmreEBL8agIYiSMXEJUqC8s2Vu4vSSPAnGodh4p/EGJKA3SJLVifUQQ10EAe2LL
nUHrCsHzbCI6YvkPt6WAQ9eikTabvOqRFHFynaZXGMvOBesnm9zECXABUdwY2V81liD6HgJ3DAwp
7iznqwWdvG4j8ZzsvpID4fbNb3roWhh/GgzRrCGNVw1JFY6Jei04tBj60T6R8UNdhechO8MtTHIW
QDPOCak2KNF5i4jjxj00+SMhPS+iBpCS+ZLS0cO+YtoyHK+YT5MmLIEtefDM6uwx6n0P7IZVP1ug
ltt75FZ6G4C6YEB9Sm5UKthFU0k7T+7mfiTeIIOTRwiP4oM4jrmDWj0aKFH5MrsEdui5Sl9vlWQ/
bGCXkVqtc83NMEDmjHaKF+r0/QePWnzxqoaPDZLAq+ca9L2Dh6Q9VVqDHudS03EpurWtI8+8VhIS
XVVICJgL5LRdqDPBGah4mGroQ1RO+BE8tcq3OGgXIutO6LQ9K482CSWcENykP/4NETxJC9Zbe3lP
81b96am4IU3+pmJMRVGQ0koZTMPWVKK3xDGSFP4IKlDeL8pDNBYT+9iZLL2FMhq7wiDmgvr0aSsM
IvHyZCLCLjAAsT22rR12rJmAqQfcDnvUSoduqYVTOKxlZsgM/gVWnDKhYjSzlySuyJzFC2l0Ux+c
tUZY8C/2WGqdNEow8LYbmKrbbqorsFyH5+7bSNyR0Ljn466NxZIjrDcTDy8wHSbdfj/oFGuk+PYd
y9Vq3Qfa+kWYHbtVkTJi2I50TBYdpP79nzfrNx1CO5u6V6f6NVIetl0wk0zS+JlKP14iOGpoUVpa
JPb0FMWJTzwQ3HwhKafFcE0uI+T5K5L5OO08L3dtQhECvedxnLVWmiWXPTb7DCBPn12f8AieR2Tg
TJIOH2YDm+WFxjO/bSiC9I9rNg4Pzt6erIeuf6hoFjihnpdDCzvWwhu3BjKqS8z5X2k4OY0NpH4C
ayYxrP/+qj+jCm2EP0COwYER7Ly8o57sC3neQHUIblxQyE4qF9OkuTZvP4bIZWBn3Iq33wYRLF4Z
ZPed235eh87f44qgaMiI0thUQc0cQ/JN+KLZCDyyLbCq/z94mUJ09k/nwAaCjD8hGTI74VefCHPh
Mla2lZb27l1Ik37G5lfxSLof9g24BtFFb1i3k/hnq7+MZDYHMbIXHS0lIso+yGyONBsGi6ZEsfuF
Nj8s4C2I2rR68W5nEzzePS6Pky+hMtHlx5MiQAe+Y7IKGlscX2XJVwM7QndDxhulDIqEvahzxg4e
LKIvJ6kHeo2PcLUbjwhebMAFaG4qpIde3sfSaIJJK7lRwb9NfX6olOGBkau+QT9peuP4RBp398XF
paqxGoqXXvd3wB0LiqLrP3tW760QjEnbtN8XBYdwsItthP2VFwL5lx8m7Y8wGX9ufl8gBFAKRQ6k
iyFJmuKSpeB8qKSHKg7NfTEf/dQHcrjKfk59EctvRRH0o+oHfN+Zu3oByu57PXb5xPhthvdROt2G
aAn9pyGml1/OZTUXM2MWbsB8TBzeMhx9hSwz1MncSunzEakZ/6qb0IBSL0pvk3lSv6k15PonCQMj
S6p6OgdbU59ND6bTEwfBzJbfBuvUAWKJN6t2grBNEtmzdQNgwr0Cf9wnDEg4rtp1eVZ+PqXP6z3k
GxHyA6BFSN4TNSvy/c7Z3UWZERi1naF2n6UbELAuaAiW9tw3r5vDUxvFh4uvyF8RUoWMN3QDIh5m
yxLOSnzpXn9bZD8VYzff1RpQz6eNnX5eJ1SQvdZzy1pkZ4gok5juCqvg1aOhcKnabTcUkkBPHZAm
5ceMy7jOQlKsjt5KU2BLzZUjyxQ0+Gqx7myWaPnel4V24jokROyNqIWjKcgQsFoZAxiHHW6+RAB2
SKeEWHHwOOeEzBcW0qNj3CZ/PspXUgrRKA8+iLvE6abNpUjKXku3lkuK+MibdEd5kGKhuY6uYcrb
xm87MpavgETos3gkdvWbzCTHduHtvQF78lHhx5FXjJ8GDi1QVrepJLSxBzq36IdKpUY8JXeDJjfz
dNsRd1ctIzb5TEnE1kDiN0DVJj4JSo4Dd2EeOstGsmvr4XBUETqb+qfKan4549CmvoWueqHfUrUd
elH/eUqIKiRplGRMm8j/6JK15BC4Jxn6Svv1mKW3aF9ZdbDWTRuztfpsgRlaPSD/dGDBkISGsdNm
EZTD5+7pvaK3zvQgDZ6/TGfbb+42UIdDJFQ4F6pJKolkDy3jsjOPyCfUkEld1pqcjyKhimbjZ64T
aRgRaWazc62ERaaU9ggWI59qFrgcN+IM8ZbPW4Bo0RzRf03P/8lKuNIXndoFp/f2sC1U2rA+K4Qq
GzDsPdezqwh0XUs2t9StqADWmWsClP805zlX1GO1jurgWFIvAI0kNi0Q85xe/KwKoFcJCrTxavJs
pYLSvTnHqi0wUncy063/qUFo85FfL+Fg2g2X0V4K/HEsrTHOpL5mHxbUvygVuKyxw07tO/EEr7ek
MjIvNCRTrLpSfj0mHUND+2iEcDsa6kdnCcNdgZxsqeqHVzLzNtH091cty9luWUa6FNRNdDKfjHYg
3nj1mIEZvCAQKSDIR/NrGuVByzQQetPvjYExTdr9NQGvnGo8kl+Eb5JnR93ytThhDgkvOEabVpIM
xqs9FIwLHGeLrHqRMk0YSX+IvUNVfxYUqrYDyKWxBbtZeKeSzj/QtRJ8Hlcjj2dBwc5fyIqEJFaG
KTtyxK28nqhlioL4Jt81T14vvP+pIv14Bb+NhvqaJKdr1fspZtrfUT0kLs8wYl5KdhE6986KG4eM
FYU3UXDM6cyaM4U7GGF9RPYF1IDEdfG5mksVPzaY0I92O0cLbqT8ZrblY1+WDpB1D8UNoPEJh229
IvspqCTVb6HWAdBmQOrOXENqHPc699aoIeNQCOsDq/Wee5Wch2ob1mAv3+mXvVHV5At6AxT1sveQ
ACYANFL0nZgsTNIcudmzY7wjcxK7LnQODqKn6oF6sI6PSSJW0O9BWXkJlcjts5MHK59ZUQCoSDj8
hvZ1z6gK+lL3PVeLam7EaOSjXU257qk7AZgtsD1KEasw1rR50zQSHFSCF9m3nIlp8wKfkJsR5T2O
d02WECM7QAUBHi2Rvj6ytd8n00gzoKTWYwBJiXIgNWwhlMEDc4aoyuQpXTUh3WHzF3z3LXY70yVc
8Dt3xaFVZyemeMjEpeTzyQgfspNM1WVEXkZKds3B9bGIHiUqU9ryt5ip9U8Evw9WSDeRy6RqJT9g
gl+az3Gg04QO/jkS6UZoK+QdycAAznz8kwgLlKNlkx9+ZW0snN9VCC85ctXA6Ovg5kco0Zu2zSik
yiP9Zsge+HO5OI3pNmHJT9Q0jjGoGW49SXD9Qqh5GEhv0lhznV4O4kYfSB51m/p3uud7OhtJ97jX
FF+N1FvbzF2AXUwI6SRkCyHP/bh1dm2lEQ2xTRc0uwzeXm1G99gcmfgBzpUctrKOUmciNFiURxsp
glhGxFudw2zKzKLZCKTtdpGrKv+BEcN2hMLHa8coXHE4HgOtLldKUTLpo6Bsdpvytl3d6LHXbk+B
6DDlyjNOl971rKArWdtipoOt74Jn7Ld4oz6z5pc6fltYKg3GIf5A++E3eLb/bedT3byGhRSdZCM2
Z7LbNGhsaLeO90l4W1B/l6JYblFEktZQyLEhvZFiqIP1D3bCZM9nE7kFLjYJZWu530buSwGnyDmh
rb5LikyjbTX+Vs62fPYxx056ihPSGMSyP2Jb3W2M4HiFegD3J2EIMeUV20bKY+TW5K2jLHMshS15
uMJVacGPYR3AtKWEu+1VaJLfKGxp0A75DRfoR9dbvy6QCb+ZScb/BEUOu9AtIe4GPlZpLVDupw+6
6Vr8q5FLtszgOAHHYPygUW/lO6++fq1t5vCWF46f7eaI3FBoCkaRq8cqLZ2k1awTsg9VGUfigVc0
2Lf05T31k3sgVe0KRthiUl9Svf5mTDaHYm4gyCkEtXuOS7Cpip7EnSArTNaIxeVFS6ODoYzI6A/D
I2BH2qOi8jqdr7CJEf1Neo1ScDUktELMkQd9xQ9HTmZHI/PRRTS01ZL1fbN5COX58jx0L2n7mR8f
S2rvbrqI1Z3HuhxTckUFEpAsh9JL7Sds6vPE95KjLh2vgz0cBB2Zwae47B/2zhCbwAOu4iENlbQM
kcmmkzb5Sc5wbDvZsEjNUW82YVlJrQRRRrLkNNNV99d4hc84spf2hMYi9vASq91FXy+8DVKfUlKb
46yzgoCEVf/SI6bi8T/F8BlTmavYPrz9eS/4+ccbvsyAMWDb4yZJBxEyMsM2dq3zvYgO3vbqpnx6
gZ3KkiLYgqLKzF/lHFMKc5vnM0DxI8G1qWKY5hLk2bZ9hDmgHMl7SJdwIJ0vpr+Bn01toOaM/NyA
1J1zVHWVFdsa7a06j0ByWf+sxxKmhb/VOQOscYsOKB+pxq6+NRlT6y4+PV003Ulxdz2q9AkSE4Q8
I9V+qJYUmrwO3YrlgRC/pxRJhzd9A5j8Ru3ubCz8Me9cvHQjWQdIk2JnDhiztHkZUMMa+MgG5D6a
ZljOJFg9dN/vYda2Ocqnp7AuQNEW5NlBp5h+cqDmgKT8iO7RAgkkMuUgmMJfBvS/tiWsRPjptAD1
JkB2cS8Er+wO0+nEf0xlsBJMED3TM5sCwVkN0vtNvW0KY0kXJOq/QD/n7kPJh63IVPYfyXJH/xkz
w3iT8sNvOX6OpLGsVRxW4Ch1KrMmfhfbm3gJujlJo0z1JJiXNIxK7CSKdtHeJ/OOhuO+7fTkgqU+
E7zhX8klhnJMD464OP/Ff7POf+HT7xT+F5hleKMtYkL5x96lWNccCHPVfk+bNDb2svgtzL6/DCcr
79tLZ2DWWkfmv4Iv9eJlV/PfgJmypI6WYzRU1egKiCD11+kUt1iCSwDyMnlvVI9UakezuwPS3qte
1JjBR2HaCc3IppBtZwgOhgGQ6tnSsMZwEvKd1UIm8yjAfvaPPmjyu8nxvMXVtSbiRkXio+m4r2/B
VCRBerEu2r1b2MEiM2mNdbrLWeMm6dWYdaCLq37UyBNGlbBBV6SpUzyC7JCPZL3V6SUvXXWw7Hc2
/icTN7Ld4bpYw9sUvVFj3aRvXDaAYbEVYEjWarry36PMg7/tOMGYSf+jP3VpJfPIfCi7isdjoYnc
XBqOJeo3oujR7hvAu9TMCO1pkR/MEwDIP4taM7zw6EeHVIZt/kRY579Yiqh0hV3pWQV0+HmUYLNp
h8CTaUOTlixtuy/y4BeOsu2fLhaZwjCbVRybGiGzKCTkEJt22z7zVxlmZ5CsIzsNSVGGsjNDKLM1
5XgneU+m8dqYLIhefWNTNRkP0wrZJqQP78lWwlwmMgRK4JBubPCtPoLFv5Zf01DNgb5yANg3CCIo
yyS9oR21IWU6ExZjbyQnFSEqbrQx5r5H6QgXukW9Eg6i/qpwT0Xx33Y3FmSHaHou5wQVwPz/M4Qj
2nI6dM+oNCXeSAYAGlajpT96JWp3x92+M07wQhfaAgbhzDB5/UG2NZ0yLtr2hYFrluS/AGRddgk7
+amMVtsx9fnslBvlqNXxmlOKPzBei6/nQrBvQOc3CqfaWclgML5hcN3016h2uhexh+Z3o3TwJzMS
4SnCGy226sLeWKi8fCkHxMUY5IP61vmgqNSDX1O87YmZaFEpu7nyOQwE4Yan2vv8ugFDs0XgqPdx
oo6puY38T/Zar502HfFKUu6fILYpKE7/qR9fCVeZL2tjJgw3CxbfCB6Bex5Jj0k1vG3aMAOQQJ0U
VwJ5XHRtJ1q5T5yNmwFq6nuv9D6QXE87tSS2gDe2trHF8hvjiQzvsSWNtbU39nn2uA7QIXS1Ca+2
jGbZ8THIVcCvJK3Exb41fQmNib4ioT8HcoY01CUJsq5+4hF5NKX1WGOfPru5/CrSnez9NfD3Gzjn
dEEFwgCo/fRyO8+rP/RD/NAULTPKx86v/3wAXdR7fWw6dE1cVijYHAOq01DtZUht87CYS8EukIk6
3yge1vwSJSnad9DH7ofWIWJ1AW4LjkbaXiMww+etqJYhGg8WuVKWw5EN8JXsskCQhPqcMeyUDTQp
BopQNVb42fVkcWPyEcfHz57SWchPvFlgs+xhQlHMKPlwASpGoHmsgl/pbOFjPZrBjPp9YbFPZE/E
EMfr4d0xt06n3dBnwaCCdWQgLmlL8BPpqZzuZiY1RfeMm/VmtAWocrlR+OXKFJcZzQOyX40s3F49
FcZHwBnuQjhLJBwOiiN05yQ08LO8cSAcaBlba6YK2WaciSgk7ev2Wfct/SWhHoccWscwd2RWIuV5
t7CpfUEkKF+nDUWRRKtu2rE2MMris6XLIBfsWiBeDBT8pTbatzMNx/TtizMnkRwVaOwq/gK/JNSE
Z6XfRvC62Vyvj/mVbMgk8Qc/Unmlp6Xx67WFRVpWYDhwQ1PyRrKKGRIqQNVypGcgh4VvRRZ6+jpa
vdEKqR1KgNWXj8JMwi4CpdAZ1E91WiUWuQCNojLzKG8Lxv1tg42HzMoWRujGKx1trf8zEJrMnkPX
82CR3iohI0vrWPTlKpxrsafLQgcu87Z2bLnK1FhUHmPuldtNZFPUwnZ5vYGejEusbhFwP2aNpWuF
u+f4SpVPu7XItbTzeN9QIcTgtffpFnOq/oFUnHoJ7vmxQxhyVw3oSYPZK/rwIMFOOzBbTTkCohW0
RaTUR0nibpJQDYtwdhT9Fai9NBudKBRHmR4zj5BwfhxjOiwbYDkE/hKzOIJJY4fUsxEyjvzpVlhf
jLVQPITc++wLP7V3RQnTygTPZziKavHy55OVs4CeOwm1ltznM9XhwuGwWNrKKi34wqD0Cm/CNnPB
hJhnDsiaP0Wb+dU5TOjn7QxAGoAogdLfEYeeWaMyvs+47gNpPTRTavVITrrxu8dCoHbvaWzFaIoh
/ebrc0D2N2bZ2STSwkxeTuS9eQyMVR97YMUVEvxY+lyPovA5f2TAZQEyZZeUGg4EqYoTVGx0OUZb
b278FfhUg/22JfM0gQAePzOYbBWdpM1UKG7X/0in1XtdK4Kj8SIKt/L0vIpkAxYsLKVN41rWN5up
w+7xlTnto+G4BaphzX9OiVGvtLVJGClXLk/Ril2nuQRucGhb0uVg2QUyL89BdGC1JgElK/Bk9xZZ
wEXo0o/ymd/5BQq6b7m9J+DSu1QfFu0E1aBI8oz7VXSlRKSEFPrlV460JMTXtJXkEvHkDaPzHEzf
EJs4oDpdhE5dsM5670k4gZUw1PPgGGbNGRGVCu6Ibmd0xLNMt+uKzgAblPh0tnQXARxk0HQHK+jY
/rS3fH5diSF36lveckZNJZkvaTtQUr4nZqUTP1GN2wlnlBkZDv8oYoJKOuv93BwktOw9DSHqehwG
DdqlvV6xEaIzAuIqlzLrW1Sxsy0YNzpcGPTG2EQCNef/5YPN3cIX7HAy2Gtb/chIRix7SyTJyGrH
jopjji8qiKCK/FjX3tGQvsAh6j26O8+M6ofHPm9UvGRBYBbqtL5obptTkKsKhsS8sFKOgnudh4Yb
jbjgnKsu5xyIgGeOcp9fV+RbQGp20fTiRAPEBv4xqB0fP8+jdvIKHSbz48jJMhBCyzYKbqT9I34c
jbjMYfOK9v2lX+l9GzRzPtdWGYwf2mmI/RlEs8+kkdlMMW61uQYl9PKFIfbE/1fOoYukGldic4kN
eo+n0Dqw9A2sf3RHU93zgM+ObF+6M9GlknHZ/b7VeYS/ACvVwilGzBk66aA+X6dOzavXOWfYiv/y
RURiSTVe98KGkqcJppmGhK3OdZzT8Up2JumK8KpIyqheAoFOyRI27gzLqsPWyowrKeUAWyTdTxR6
ASOwp/Gf9BDpPjpLJMorb07defpLV+7oPmhMxmWwMXkCSkuZH/IZMQaLpvP/Uqav5m4rIpwpqHYh
+O9+TRp8JWXNWqCvZsGVNuKGbc2ybzb+HxKOTpRXMvlhA0XzVHtJOC5V8eBWxKDhRvzKAhudOPO/
MEd/EqwbJjZNMtVDAs9MGt7Vp4ZALwoVSgG48/TFRnVX34fpkz7uKQNDHrcPAZAMN5OE1p9tnQEZ
xV+Cr3GxhlGZnvTZYHgAowgA9pwJ3C5Kxgwosg6WzAOX9LmKhQfZJSmNxSa6sxThiDx8kXOQsyWo
cdPApgl6gUg9q96u8cpi+ZgecTNiygY50Q5srvlyaSniSsQ8q8EF2t62Zlnw6Kumohikg/hEFZ9Y
rf6LTE2cwLy6ZnpL76nh6lul8IFB2fLEkCPElaOPhS5tUB0QIzWCggoILv0MbO9REWgc2Ed56lSF
ERSSe4n6mzFNylEwfIgVfK2nNLO1mrGaH6IfjjgNbWMlq9rgfnMitG4mFlOoOGEfBxxYa5uqJnwc
MpkwEjIIKl3Pue79YqgFvtN4lc5NUVR5QFn2Uqy5HRiTWPEnfEGeN0WuBJwSP52UZN0WFMzK4agF
5EcNrDsEoKfieQ3VOx6+U3IBvTLl/+sJii419bzcsR3zf8jsO7UwngvFJxlsl7DtRA1e6IROf7qI
mOak33Chq36OkB5UGF8ku2cLR/1pDeTmLaa3lTIsUerzdACh7W8e2Wd7+ChgqkDesAivx9XIF8B5
gjIaRbmsU7d72rRoXvAsfgXu7vt9mPXBGbS0Sp6/gbf1SeN9pYH4Tjp7uSxo8k1zXaHiIf1pA/9H
kO474LcBCcUfC5YciQeeX+1f8TUtk61uw1D5yqIItWPSTY16JYvO1BdY6gP5znD1syqot7eC/y/V
KrAnBVxTmi+TSJPO98C3VohCs5Ak/9bV4dwHKwr2zmSvYp4vYln5gm7JkckJbnuMXgGhMzsUaVE0
X1bjIwOD2CuZrIDDRyBtnrb4oORJhL+H+LZjywIBDNKtp8R9D0QaCIWZKNR1n1sfiC6YebWSwu4X
ZOlFm+Fz3amaFdcyAiL9c/R/EOGrR+KA37Iv6SdNZd5gFcH6BekH7WWyXgo+KpLD4KezdeRY+Uel
F7/XZVu2iMfJ46mT9HskX7m0/9YwqSg73lJAgepqChD4+nzTQWPC155EPPRdk/acohJF8vv/Ez4a
8lb5ti4pNyPhT44zZNJ30BtClbsgJN50D5akV7WwcjaDRQJYey7qZ4lmudgT7PL+qcuxz4xut7NT
3VrAKaI1MC7KlRS9cHxevTxVJqqASqjI1o6qGAsEGMXdZhHq7d8VSk3TFHgP4IXRf8qQuhxFhbg6
j8pwHhjnPElKEaWy2B8J27UA6o1kYCJaIsNXn5/XrOcVn+QeEn1joe8QvJ2NUwJpBm6N+gmesrgA
qONzU8Uw4OebGjfAeUnQFKXO9yiyzCjfHqqMPGMX/RCmWJUfQwDZAF1KzA+DOHDJwt8ocl6V1kPi
DQGKMnWQKmoF1MKx9ZhmtsyslY7TBQ6lImeIZDz/UhC17l/0n4A83TIawsPZGNuaZrv/kZ5i8Mgy
wq6GclZNdX+2UogegEsqa2er0SoBao0A6vvPsc/Os30M0Zy/WN8lGo4zH2PUPVXlicQ5IIwTM8Tk
wmnYguuHEXoZxUmvsfGIKMyOnyVoa/QVdhkqDL+gC5ZLUw9333Ggz9BT6amzMzswZNtB3s8OMZTS
frOtsLvZcBOBKLV5Uy9SS+kXdCPeBx1y64eh7zK2DFT/y2qU8fI1uM888cgZl6uUYP/Dc+y49KPm
L54SNWKrT7pPnWbFykf3VG6BKiT8V3xEnchW0HhYA/brw1E1fLbNkpYnqJeg4Cr6cVCF+N7ryXhL
yDy/+NbRltemudvsd1//GYv86r9pE634PW9NXigbUBvO4oLZPsBi0/l1wicuJ/gKCnOyxulG/Wlc
+jPNFIu8Byd0u073/Gydmb5yj+XYwaPvZgixdj1SKdXmL/MYsTNXTlMtepjOXac9hCndg4tz4Q7N
Lni0zUPWpDXdO06OJY7UAN5uz37nwgzjnVEnM4t9lNHs9//0RUhb+lWUmFxrk00RQmgxMm6AhdFg
JxNCrqwpj9Mr6/Izxttli72rlQpGiwwk6xjEB7rp+kw0/19YXj3nE55Xlfhsu6zZfTFJMs3UVBD1
G/50GvLM9pT495LIBq81+XF9SygQp+4Y3Obr2XIqaY/mrN+y0jaYzhuZrmYFV9gB3apQDj2WFc0r
usYZ2+BLnvXSr1OdbpfKd44I4iim/HZUh5D/heExmH5DFWlbYRtSDws2QK5KUo6L2TP+acidqQ/L
n3usL4SG1d8k1+TvzgjmayvKM0+RjEUfMO6sfEouXT8sinlQFFaK5WEg4wcgD/fOZyjFd+0ubSpl
hPBrPRdwpBYd0SSSYitUY3pkNDyQofu5ZXCcH8YHqCBdHeawssO7nUfbolWMUUetLL/hj6lyyAkc
9Tqqv/g80z2iJmJEmIqVvYdqS9jxv6PvVyMuTESZS9rTTjkG82V9XLW8V8SrABcDH5IYiO0crWiv
Dhy/hN4K1sufjHPC0PpN3H5dImG2TtsZf9sxRZ3Vl0SUMk81X3NxTF/TYRBibztiB3BaQBB856QV
Kt3LOUtw42wcwwS4h82JphBNpDfuFE6jdH+OMdUotbGj8YGk0cKOJQcDN6K+8gO3MFtUSxO0tJ2n
T0nsgFGqavEAFMgajyLAO79fRLGNeJNR6dqH+8OaAYn78k4c0gwJtHH/Z5W/RbSnBlNdDVxQghE1
BxCp01WzI1RSuOixRkcy+D6RmgTgOmDshFgm+OLzC8Wp0KscSRfy1n+u3a2v/8JQ11NoEf8xOnjv
Zbi89ue5DBANL/M2XJEM7FbgXBUnqmMTbdma2CTbYyw9e1bpK6X3NnMFMHJEmm1IuzZ4yZnDBFvO
pXz+nE/5oScXRpMKe8ENjkbVSo5r/NQlJ74uyus85xFMWbEjWZprkpcHoyrEUD9x/excjM6tUU7O
sFJ7WZfDuMAb8UPRMEYHaBvJWYxURgNJfChLqeIHso8vn/4RCtZmXFx06C3+WKyfb/C4PHlPvy3O
JaEppv2Q7ZEFGvRz3VSNKsmP0mq0Zzo8EDhQnN19m+WDq4b9uqyrNPRyI1SbUYJsCdUIxAJQTMYj
KdGRMYxSFd9aMVn4Y4wrCB1JXLXRVjIWtVc1Bn9klRQsiKwzdkmLNZpr6NDXF63CTiIuVlR3Nkym
gAiEQp5f8Ur+ECz3P5UGqDX8/JhCzT15zmSddyINaWaXDqB44jlRQ2ggGVXQPaCk5rlqU1qH3iJ+
pcp9Oj9w4K7s00T3TyfWXEzp9Nxc5RzFs3f5Xdq2ZrVev4VM6EEzcWfgBcSa1JfY82Iri3SWn+aY
lqGIg5WkT0UXoqhQK+AsYDxDjOFE+KbW/mGqtTo54DbCyQptBzcEoBnBNNRUCbQ1POIk1968iBNq
jy3TrU7iEb3IwmyasHScb7RVAzfErN8qW/jbhhuwOISFvYEePYhvt2jGPj8C10y2inoAG8zNC9Sj
NQddc2wQy1JZ38Cvsefjpm30IRylrhnXc7nFlgUlvJRXnxk2mdmqzB1PxiAJr6Xd76BWxUzNigf4
tAd7hM3Dd+092SQ6HEgS7JMdJgDDp2/6ZbdaHEz+BcQUA65FmXnyZLeZgKPsxPnr28EzzFjScqVQ
XLK/PnKaeZv6Fh/mMOxToMZI++WF9L/opwKo3jl8QeeZ+sECMeTnH6PqrJp59D/ghV4081w1GYvU
0rEr3HUcOn9g3Lkby0Y75GXTeV1xk7bSCXo6fakv2a5fcBoK28Qs6SPRlCN3edcqp7kSWZSUzr6m
3r9Z9Tn+GLc7wgVEkbdIKtYKmAjoE0NtlcMvhbCuyRG7M1VHLvp6EZplmPTRTpY3tXNGH9f/EtbI
vF44HDjjOH6e/07TH/Zie9FVGm9KvEhJdajtw3lPSGnvGjdJuuXaMsOjHNS4aPQ9EV7tg1xCIQ0x
xxKqxgKg7cLqvd5+7Og+R4EOvpfEVI/dIwfyLugEP5s+CBAX8PdhrIVvEuD19XBuvuyMa0p01AH8
clOvlfTiCbExVSHSvS4Kdnm5OyROeL9dppsqM0VtHXRaS/RfcLK+RNM9H+yaMo5HGdox0z+3K9Hd
6iLNiSdPTt8aFvZ/z+CKUTNGxQrBtHy5zlj5ADq7tbAlvmusZwqqBVHaEkyRtZW1d2nsLplEskOA
CwWEjjNJv4B6eWOG/e0vsDZhIlIikPTAd2mE+jpZlU1XKwCn2SXwl2hLtyOXTGdJ791qezhwTFlX
yGynPJsJF1A4Wmc0TrPJQcMpgi9zRqcCXy5Y2mannMERkeHHofhF4NANTcrTtyVS2Kxivq8tSRF+
iSzj1BQeMkA++nUCOKFpYqkLEP8Y5B10jh7M5iSrdBJ04NmeuCLUmCfU4tlf3KBljJ97ecCdyKoJ
PPaOENG8m0DkNlrndwdrGZJRfw9LFdE5ZDKnuD8U0YLWYT5EHuDGRjZKHJ29PE1vPCx9LPfjf3JF
FA9wi/WdjgnV2hvQhAN6t2zN457n67ckSSk0v0irIjNOrFAoSvMB2nF6pbER2gBKnRndgPjVpmWb
zoFDWyfQRhPU6h7o0KgDeEoSosOkI+bwnuURnJGDZV6QdML8DhFnrtDYxTI+zdAVaKzGU5tA9XoA
toUdHw1YREljfDaap9010FPZDbpDj/jwnG455wsSn30JrqI1ZA8xq5zryOMfFKrFpPORDPEky6CP
GAtI8/uSq9g+fQK7ZZWNI6he6CecqdeOvbnSF+Ubn9XMZblBfP4q0SG9Dm7T2PL7tMEvjON54l78
GZqqwVK2+zp1RaM62E9g1GlLFa2NZC2wlxTL+VMnSeHA5FBIpiyShSFoyGCVxCRx6ZisIkWV0NPT
sxgtJibWhOMC+0HXihgPMlDqcP3ufZ7U8l3wnNlS+fvmWWrA/6cb+mNxONlVM2oNXDNrnwi5mqRy
HtB7XQQ0y1t+KAU6v+5egSkh3OV+rCX2LsB387mDxlJt9VkxpuCVg22cKasqR4ep083lk36yrUqM
BJFavbup0gAnqOmoSwBurLBYYk/IvwsAW8rA8weaaS+FEReCS+jk0cgn4xGPILinJYntR7jeX/QY
vq9LaHzd8GLUiqvxObKs1AVMaiZ5lTkZcJ3BZ7fl/fwAfFXu+MMt2CVvGtnrKZg+WcPTaZGZIDIa
NQD/zI/UOnsNYU8PY/mE4yxlC4IZsnWBdwUIfGbFEqz4HLyNHgLSf6R+RilQmll8lUyu2QdqQMD7
CNSppRbmjq0OXW+A0KSy1aYgnT5WeVs/1glB4HdKhlVHIi8zNSFp89Y0Z9NNgegN3jt8XMUhAzCn
kEpytVbi2BjY+2UX+Bh0A2bC45LdvNxFA49mP7EAcqs5CWP4yZXw/hDdWehl51BDAYjAWviGdHAy
S+XVOXVnljp4VPqpmnDNaGzFpl33VbZxlCNWAq64TF0fvidFNUHgYWWcb3y7zOsmvsBzY3YEtnWY
jd3ynMdf+v6Rwkbf1etNXdvKI5G0kuZL3HiTut00/3n9oBBSjrWyBVVMa+9qll+Y8cceZfTok1YE
/iaoEB3aYQ8ySUtLtA/0LkFd3xqDAJYTeAPHWsi4xttx1+Rp8ZHVOheDEQtVN57kJiFAAN3058we
nzD6a3PvheWhJj6xl9HranmNg2AU+nZuHhmc533czOnnAuo5fYXWkbX6N76kZkB5C2cDSF/0dZMF
nOZ7HxRthVsi8ttwcbvUy0qcHHR+C8FPJzuIsToPaY7O8J6nOJQvNGBjIwnshKIqXzB1LhlDLvZB
9wRKXGfkoXcwXO+Bp7FZRokd/tGT44zKBEcg5oeixJ7KThtbhc2xdh7LBP/836+iNW6AiTOB5RLV
c2ZUdUu9X1EsuYE5sGE9TVzGrrwiBY1h78oTwiAWlrhz4RpimIKwE8ub8h5pfOtGlMm3RRQPHU11
a9cUzLjxP0N+0IUoeHU8+i1xN3R0LsZXvttq5mXMeZroc4ZLDxLs68jU0jan4l9dBG/OE9PhvWYi
EVZrfV0haA06AgPKcS1dPkiknOxXO5oy/PM6mVNlSo1GTys2Q0YXt0D1bpor6p64BAqlRghNzPh2
pdn9GqmAYSror6QZd5ghJz9089fO76SkD0p7KLORrmQmY3xsrgsPnW0ci6Hq3arpdP6/go2AIfqq
zFJM1yHTe2mpT3+hYlGtKzroRFNl4QQQOwGzadohaZRqfFBmaR/qq7mxOdwTeVN6iOvnkX2q3uIi
2yK7+IKEaBwpRObNKk0AoH2cZybb/gLlxOs/K07rKgdvOBTosqgCbqwSc1DkHlFpsXc3cRgIL7aN
gxfFiZBfmKZdMa/GgwBI8iliybcFnFCVwo8mdsAbwSpbdvupD+tg8QXJ2OzE9dhza2b7pG5oLAax
5thlpDGWbWJYNtexwd6H04LnSNUqhUuYefEu0E2SEYAhtZmdhPlxHZcvWo6vZGcvTge+kHzyUidS
CQZXe87eE7HhKgvv4fLARLq+Ky553Bj6wkLN59eb+uQdnJeR7wa2pWfNxTqdtue/6viAzcB3sh4F
GHZ3fpKCz+Q6pG6FBSoKKwSJXSm1UORWT/iUSxGlLeGm5GcMOhtU3OQ6DVg/+2psB39L43UOTt/R
4TrIvSnGA+K24p7aHBtis4+bZaJcexI3RX10T0Prd1F7ZBChaSqUMNAns5Myx+2kNEtruVwA9dx4
AIOdgVr+YrBe275X2P+iH5Ib79nDXllwHuoZf37z+ao08aBaqlLnL7bLMHboabnSuqRu8o84vHNO
3UmSYI5Ci76XoI6MJ98A5DUbI9tZV73dD/SQ5edoctTBWkFqbQV3Lj9hnSqLbwttwE9b18QsBel3
kv+CtgcKqWIdMmTn7PyaHpo1DT/H0zIUmphxOrZOzQNRdfghuYqczvF/NF7bue8N3hUmQGNrfP2L
gQIUVaCufmIAMTNrB2HPWiXwtqfgfDR8VvV1wtYp5C8SaollHfl2VuHIO5Ivob1eTcrdKQmK8SPQ
03nwM4Yp7DuiSQhKofjL5yripMPnvlJIcVynjv8aZ596pbpZ3k5sOoVYqaoXLGlfm2BuKXBdD7UP
j5ybh5Io9hpELKbdpp2e1detlRID+adZcs3VN60IelihUNOa4/isbw5LOBRBloMneMPVGHrdlx13
vrbFVfBprnAA1aKZNjFhAt+xREh4Uq83FrECrh0MN0Q2jXbbMjqBdn/WfNakfwru65ZE3MxHZhu0
ZM7JtVBHh7V7JVstV6D4GNAHRQjg+1AtGGFm2mwR4GVwoNPYxd6onasMFeRmwya0F0h7VTj7qz3D
3X3P9JYLgh1EQzTTEhW4qHqpBeub3DoCcP+M1LKLmIU5VIRPdqikAdLEccNUnWiXOAiL5AzaZGmg
+Bln4x5sxqXKmfXKB+vqHtnzc5n+0vM7TMEzr/Wwt8vINz9K2K4zjr9TLbv6M0CvQ/cBpwgFMMXq
gb/yA4Wcs61bDzwcpqYrF0ogSOGiEpMNI7VCv41nUvQkx9IjFPMl5RuDG3mwiH+lELK6fp4GZHNS
fJ4HNbzPt3EteuePH+HastGfENQtAPcDsg==
`protect end_protected
