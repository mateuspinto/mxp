��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���莑3ːz~�H�{j8���_L���-Z�|S)�\Ί�8Nz#=O�etU��̍��k���y^$,�0[�i��GtT�,e�՜��f��f�nT&Ձ����~�c���{&︹�OkZ�@��"oc�m]�j�N��2k����	�Ԯ�Cx��M���;)d�¦'U�~wӑt�2'�J�C(t�U��u`�K�H�|.�E��D�t��]����YA2cf��84B��j˷\�3�����?�V�^�uj�	<qs
��ȶ}�<^�#�`����qt�ר�X�頼
S��(�L�:��[N��mA��=>YM�Z��S�sݏ@U*X�upO��幤���)4��:Ek$��m��V�b�N�M:^�vk�Eg)�aN�(u��3���B��ŷx
����~��Q�9�FM�y���f�b�`�Z� �I\�8'���C:�j���.�T+Z��e��Ѐ�OƸ��x�xK���������F�+F׹��Ync�i�B��k���\���c[���;����j�Ii�:H�f���1q���LGء��|��-��ǡϏ�U�i�=h��dɧH�Q�dH9
Ɩ(���*E+�MP�0�Y�_�h^:;ћ���P���Ӄ>���ܨ�
[rHT�"i� ��(uW	!��5J|�]���[)8��e��َhh� VB`i�t�"O�����p��[R�.\�i��Z,\�rW8X��l!�n Y�P-�⺌]L�PQ�����WX Wz��
֖�춵A�[D˗���w��+�_,�ʙf���H����kt��-`�l�m&�b��}.��d(�_�:��������<\��t��쫊�o-Фj��cՔi2q�z���'
@�8�a�q7��퇣�d�������v�͘����1"a,-<Q��N7X+��_GGl��m�b��3��7ے����l�A�^b�z/C�׌��	���]$�cm��-߹�}}�&��gM=�[�]�m�a~��K]_ΆSSYd,|�n�a	�RSޗnYT���"�Z/h<^�t�2J�7z��U�=�IU/������Iخ$4�A�I�I`M�:�%=N�Z�7m��d�$e3O�ũ	�S�h� �6'3�K�t��C�C��)��,������8�:\��'W�l�.;Z�/S01�I�8�	^.eՋI�Pyv�E��=�%G�,i���J���qac~P]sɑ]�!i�����s)�c �'�We,�R"_{,�N�l��T��<���<���F�Y Yi�Vj�/��4��aW}ʧ�g�����;awo㘤��0�M ��(zz�nJ�0��Y��cL뾩��.��U�H�z����m��þ�����Ϥ�%.:y��r�Srl[�����bgG������'�LD�i�v�%�ׅg�������c�¿P��,,j"Ypr�&7�XRKq�'�- ��F�X⋿�n�\�H~*>�[�/�[�N�b.���Sj����y�$����%�՟��L����5�\�u��n]��n�	g�<�G�<p��������JH^��9|���e��K��v2w�F��_ّ���G�VM�F�*�Ɖ�,"�?k��ҵ�y0~g�J)L�h��"�f�\��E-�b�nQ���@2N�l �T�@�v9`
�%����%�� ���\����QnD�.�2@t�Qh��t���_l��YU�3��`rnJC�{s�t�yuLa�U�������u8<P��|kM�G�B�K�� �[��83w�t�V�Z'C�C��RT1��F��ue���_unRQ�Q`�g��-t�f\�@W�ֻ�szO3�0����R��@Đ7pO3�G��� ��V�s�*!ș*�:���3�AJ�zlA��#��7�	Kg��ih�C����6>��sG����J]���~��6�l,�������n��(JnF޼�����L���<c��V�?��I-����0�bU��i�8y���>�4�Ü�8�ҏ����DBjQy��F
�|Օ�<�׷�;�q��iiafJ+�޶L/�~� YgF��"	��]��'�C�X:�jݝ��<��G�Ƈ�h� ��0^�fC���F�C��.恽�'))X�v�yqӎ��[{��^\��l!��a[P8�fRt���ȩջ3vk*y�y|�)��kmJW6�/Wɮ��}�M��9�wK����GpsQ�ɷ�t�ǻ������*U��:�����$�]�s��5ޱ3F��gL�?���W�U�:�����TV�P��ů���7B���ȟ��۝���:d�G��G�\����+K$_.sG֭�<���1���9����ͬ��Su�7]���t���bvK��ƣJ"�ib�C"�F:&�o��0��|d����I`���LeU�y-��؜��
O[8�3���� �4b��boP�J5�a����������n��{���af���j!u�����a�4��kR2�P"t,��E���SO����>�E�v�%-�K3�����j�MQ<��ց�=�zL
��,�!t����U�,;|=���+\Z����4  A���S/����[��}�.�2I�v=t��Ckz'Q���[ɽ,�L��Q�αg��]�~�ȱ��8D�h��ej�os��xN珅�g>ø�@E=^����rD,߰0g��\`(sOʑ���4<��1��}["�g���-�	����C��gƊ�)�a�'Gɺ��y}tO�6�~��Ӏ�1��5Z�����4[F�	�n9d��'��y�.��~c�c�,�٢��Jl��墤n�������ڝ:A)���%$�B���r(��Y�!!(�����{����������M��g��7���gW��1��ש�§�}a��{�w�eXe�������<�̤K���so��D|��m��6�/o�L�������s{ �>���}N(TC ���(!�6�l��S[���o�yD��,�!�u>j4�@P�����	P�Y�V7��2��"�c���Tg	n��H:x�+2�:Ll��'	�����@%4�Z���������a QK� !_T�)�:X�tݙ���vڅc�j���8������V9�J}�����.��z:�����4{2_&U�
"u#�ی���%����'�B'�t�vv>�����&Ae����p���b)pvcu�o%�E]�����X�	Ê=W(zp|p<xWrچ�������#��'������9��{Qּ��1�LM�\TX2Q��j^�=P��oBV/%U�l㑸Z�(y��'���Y��@�5'8��D��F} - K֋7����t�i�7+�O�73:|����3_���Tפ�1����񱐛il:��G[D�$(�@ D�N����}��AX��jn$A�kN�c1A�Al�'hҒ�[��{��W�Yc6��	�LP��k'�ě���7\v@��"x-��t��SH����2-�p�%�dM)m���7H*M郱�o�y��t!4Q�� Qpu�+7p����G�P�}���>�ua�g��ID�_D��
�0 ##�h����W�)|�����'���D�&�c�w��T�
��`��Sޮ��z������D�7�������p!�|*��{�R�޴۫υFX�z��s�>��)���VH�d��.���w�6����ģzi]�mh'�f�㛤�ү�����cpo{f�3s�Bs�̛�:.��:K�&��4s~�M�{e��Rv��Q�ĕ9w��/����p�B����/D!��]i�v0�d{�I��Ze!5'd�L8��b��gQ�k��<|pݲ�9Z��FV���6�qm<������E�lh� ��(����-�q���J��e�=/(>7Jy�'-9����Z���QNfۘ�&�E��m��ӎ�͓�#�^������1���/���1�X���c���v��X�".zot��ހ�U�i.o1`���w����V<}��`��씉��o#5Gf��g^�Vog�������tE������5���ζ?vY�_J�ɒ�s+�7�٘�r	�7ߴ���\�uL�4�Z��2,4������Y��<��L��mRA�o�����ł�����qi���}N�v(_�����x��:�kTn�`��jE7�-��U�?у����m��έ�FQ���n\\h��G��ڄ��~B~�� W»^����n~2E#/zQ�Z�eV��z�oʺdq���%�#��-�hMf��4>���t^H���}���4�
�e>nz�>˅��gΤ��Xb�.f"����g��nTg�F�G8l��މ�i.��g�l�.z��E�Eъ�v\Y�^�w@�y��9L=Mk�BlE9��J,�
X\�[S�)������BCc�#Ÿ�Q����PV�%����][�n��큾�NPٵ�5��o��^�����
/
3���v΢�����>G%2�/ab�89��#h���Pvb���Cz~����b��3
nn�V�N)V����(�l�b'
e �MZ,Ym9qb&,0zD�����r>���m�p�$6��[�X��u�d6�!?AjS�P���wPd,�ŏG�G�ۦ$����D��fF*��l'0�o����Vu����.� �7 �9r�e�:
��@��]'�m4L��J�s��G��7�ҴH�� � ~�/ui�8#��$���a�)>�(+���)*�����K�Q����h��]��)?Zx�^ˌ}k�4�X{��P��e���U*����G��W1�l����PI�3RF��yټ\�R�� y��1~�n�[I�W���i`�?:��Y[�%�Un`$h������y�×��dD�����,�TN�@� /�$��C����-G���>�F��SkYg�Ei|5������(�b���WR��t��l�(�[ԉ��G:A��	tX/��'ܺYQ�TK+���
�+��cp�@�"��~}v��B+�!�]|�_W�q����T���dz�F�uY�Q����`������& �c�W��9�h�ABb�.����Z��! 2R���rp �\ˬTq$�BL�E}G㿅6�RE��
�-�r�4���ח_Hp��̉~{Y,g�	��Q_�Ϸ���+�kAUb��e�YSܱ�{�,-Y�:����e�ry��*�.y-e�Yp�yt�A���;��@e��'��������_�a֭x���0U��Q�:8��ȋ*x�dX.6�L�fz�el
=� x{��[��"� ���(�^.��Yn�NOk�_p,5N�q�"v��'*|�/c���;e���`�pp��K:��[���#F��<9�^`�?�\�S���[�6�a�HT��s;[�3H��R��d�J%ԑ?��߳I6�,�<T�?/W򩍤7��Ӄ�Rr9¼�QEW'�".J�Xr�#L����UH}�Cqj�Q=j�C ��%�Fax��2p{_\gwN3������,9b�0�[Q*W6�<7���e��8Z �ʏ�io�{��P����֌���]�����I��B]�Ϳ_���{��?m�n�$h�\u�����NW�>����w 0�����P��wq1�5�f��Of�QKV���y�H�`�jr<��B��]�����#)�k3z��M�O'��p�l~�|�%�^'���"�P��z>KNE.k��,�������S�U%�E�2�mG��>)$�����C��H1��������@��]N�(1�Q`EFv�Gd����.�M;���������qKo�A�� �dͧI���q�;l��(-}�>��f���j6��[��!���#J�|{z��3�7�IUM��E���X;#�J<���f��5���%�cr0�8��I։`t�e��Z)9-�%]��^�V;v��1���[L �C���_'vY�y�
�dĜ��Ϗ�j
��oLhs�5���*�,Q��{��¢��AP�5�dr��LХu�q�zB�9�5�Xg �J[Sx,��I�&q2c�.'Z��~�onh=0�c�V�Ii��h��%���+.�?��^�@+>^`�<(�Y���`�[���'�8h�̝���5���Z�H	_�5-�a|V;w�6�'j 4�26��y��J�-#{��ZU�A�5�Z��f�s��z�v98A���0QJ�ש:��0�x�^��ym�QG���Fp���o����jsU�!�<���,X��(�Hoh`�_��%2}���xu�Ҹ2����ꕅ��ދa}��ӗܱ���$A	y)���:~]�A��?D������.�N��)�>�()���xH5R�Ϟ;YQz�<v�Z7f{��#�u��SWv5������st	�� �bL4�r���g���Ltkm��)�K�g�z 8�dnT.J��j=��ŶԠf������,��w�6G�G�j1��W�E�L�VK�����;��9�����`���UMx��ZyA  I��p��!����� >��s�-T/���^'�5������nVt�l�5���V��S�0�þP.Y]5�;cպȭ��OX��6��������}@�S��Gp�������ҜX���J��2-Yb� nd_o%���7B8^��daK%���a�˖7s�k��_xY�ʆFZExͥ����܊��V���\��0��[u�G
�EϱpU]��o��1ԏ�Sl��/��<�6��9�Uߓ�a�E�������0��sB� �����XѦ<�ލ�Q
��U1'Cd2*w�C>`]g�T��h��L�7OPM�T�v4�(5C��Vle��glfK��d��1����L?Ɏvn7����14��+��ْ���J�!��j�O�������V���Y��E#����.}��t�n*�ʠ;SZ �~m�t�=Zd������\` ��w��l�!��:���,�`��+�'BE�?�	��E.&p�h��t%tP�T�K�N܅����D+{�g.f���1Q���q�4/2�U����Ҽ6"4�U;�	�>�=��P3+����:�����KE=���ucZ��Dszl~eBV��%x�Tw&IN�uox?��� �J6��FY~%�t����[��9<4�a�ȴy�6x��Zл��h@]"��c@����m�m�HD"���ŧ걫�%�!H,F%���QUC��e0�_�
�k�͈�� M�I*B=�;C@M���(cy������ǲ�H�&�W$[s	�h9C}��~��㮮�~���V���Dݔ�Oc�,�b��,bKh��+n��H�U�M�r]�.p�O��l��0z��n�
�|�,R��3���4����}fvnP+��pfU�/5�#B�O�1�;޽�^g>���N�P����2��N�{f%�T��1�ȧQ!	*�mx�b8f���F�����]�ݟ��g�m���<����������9�+|߾�9��#ͧ/up�+4��K��&�k�g
�`�h�Q3����趢S�%��L��`�����s�$�Tr.�FaF���>�nStY[�?��Lb���))s�t\���eG��AKO��@���I��?�C�]U���ה"�p���1zE0�%j�f��F�LfDW�'Ԇ"��Axz�GD���1�ޯ9���.d�-+OH���9��� \�������,E���ʺ�nCk<t��=<�r8��CT��)��	ڇ�Btϟ�K���LKU���<�U�d��c��Ts��q���X 2�d�7ZXx��-�0�BOYQ&�/^���f+��l�I��k4�#���?��A�2�4�n��,h \�c"� �0�8�0N<h��pV_^�NKv3���m������σ�=�G���>ͦK/�╪\�����*�U�o���F��Z�![R}��g�X閻���́��.�^]�������� 9�Ȗ����1�:ڙA�r/����2�F�R5���ݣ��U~/)�^��H�B�V	|��&M@aA�����,����Bu����/�LF�X�u�������	UHЃ�-9MTb$<�����{L�f+f�e��idP@���p����5�%��	�Y{���I�s*���<Jot���S�%�u����cM�F��r~|o �s��?�����G�/���#�(�\����ΦE�✃hT��sw'4*�F�i����lӾ�8�7�v���b�d��.@���l�>���)[9�7Z�)��=N���������L��w��s�G��)����@{J�j �cuֵx�3�r��Ij���,XA��������n�CO��>�54���ϰFȸ�	�R宝��|�mJ}Rú��b���3����2�[.�&��}��Fgl�k��6��p�s8x�d�ӚfK���*�K�l�5]��^KOĔ��~=���n�}�m���������A�\��/J�I���@��P_T�y���a��ߙ��D~�Ilqf^7�td���뀴4�Cz3����CQ�}!V���s���á�`s�B����.<!_-�:�)�B& ����Ɗ���7m]m��q�P�B�R;��׿���y[�������AU_�ܽ��XbV~m�QP֙6lEP��+��n�nQ|=mY`Ǣ��B��w2ӕG��SR=ߵ��; 7yV��T���c.xE�ZA��"���n.ŗ�~A�>ea[�4�ڜ�!O�	Ċ-���y��܁J"X�Va�af��c��h�"��*�c'LO�|�*����.�4V��K��Tt��8JE�7�2��#���A�-@Q_m;�!bsJ�x�ۍ�=���^�����(��;ySٓ��J�	Ϳ�Y�7��
)�6<�Y�θ� -����u3Q1�����y��
�qP��������9W�I��,\ӫ�ݥ��+�T��f���1�-t�(c��K�YN�{�C},���FL�Y�Ƥ.c�n���y����G`��a���o�U8LC�%��^��r3OJ6�����I�51�~��]�@�a޲S+���3����t%���3Ʊԫ콈y� KB�YJ��vOʿ�=\dQ�J6/K�n7�_��u_��&=Q�]+���A>ժ�Ԣ�fy!��~�$8ٛ�W��w�-�h.���3׏��#�#7A��1�B'��%��c"�����dd��g�'�_zm�q)ty4N�]u�5N��^�c�7�+����ҵ��3Z@ӭ��߻���uϚ�ڎ�U	�L�Զ�rUM�B+��}Rbs�p���=�a�&�s(VD�^����� D�Q¬?��_�Tu�/d��be?O��0O�]�$�h�A������_jU}�Ĭ��w�c���JU�M���\q4�x*	������߳��0�:�@z&��n��S��"���Jap;�D����G�.���o4U����RC�=�s�
��,��`Z��l��lN��ޞ%	�Mlq�9穨6��p�u���Q�6����p��uA+����I���^)�K������E�p6_�-"qOD9�� 7Ju%V��r��؀O��1|`v��j�7�{$J���>�e�d���
�u�a��+m�`5D?,C��Z�m��5Cw���О��Η��g�"!k��mX��b+x��`$B�'nMk(0t�;W՝5<Q�g�J�������D�v~sX��٫�=~����唰 9(7G�-��e��%<�%�m���6H̔�돔��|C1遞���4~E� �����$�Ի�`�_����锪�Uc&�ˎ�6]D��Ӱ�6˽�t��(iH34��Q�'몔��(_[��Fڑ�LJ�@yif:3K`�u�L�'+���q���σ˜D� Ƙ��I
J(Q��:���8x�����	���]�`M�T��N�
`c�b�Sm#]��<,p��҅�o��x�H���ZV���.�<۬|�cI�c��ė9��l�o�
s�:b',.v�?�W
"���u���7f\���?��
�������/@b˓�.4F�h�:t����4����%�"�Δ��y_���跓�Ʒd�~1dK�����?R��p���w���P��8�v����g	������W-jg޽��/�Dٞ���\{g������ەˣc�՛ "=bw���G��`0�Ѿ�j�[e�_啹OP$N��l�N�I�J��Uַ~�w�yщ�yY�Y���k|���P�v�����D����jS�K]>Ȩ��?,[թͫ��A�}�}��NΑm��9ŗL��IJRӶ}�P F�ha\�x_�ݡ���G5��Q5���n(9W�w=�H��ٻ��	��ag��׌%K
�yc�y%����n0k�Pmɜ���G�N����=��\F��y�o�Ot��-�Tڅ!in��5��(<�q�S�����'8��P�n�A������	t��rM��=�s�����X�p�%6�]j��8f}���sa �7w����U�Q�`�C�&e�4h�u���L>�Ț�t�v�&�,g4����L�߲����5��$>�y�,��b�̀���D��zi�Mo>�XY��}��"�>�o#�1�R�}3��h'l��[��Ϙ�5�p
�/Sk��~h����`���29�{�N�0��]tJE�m�[Zݯ0��L��Wݾ{�3� �A�p���M�	�W�[��F��p�5�}���YQ�3�;D'���9&i�����Ϝd�Ts�oXA�`��O[5@�5L�$5~:<>M�L��4�^�y*�Ę�L+�~�(�-4Ӊ4�ѫK�h�����wۻ���CR���@�����*��7�R�f�3��C1���H@�Ad�`�a�&��S�C�S5M+��1�K�#T;����lӆk����]�_H�.��=�z,�fڶ����̉��<���ĎaK���j���<x_բ�݉C/B3<�Z�W��b��6�Fjax7@2��.�,��w��(�U���S7�^��#���_���p����+S���T�w�`���ڝg&�=,����}2��\�u:'w��4�@�����S��5o%�iJc��LO]������(��7�ZJ�@m$]�R����C��x1,�������xʓ0]�3b%��k� ��)������G��Ss�������l
�ZlΞ���S��-���!��zb�eB��+��:^HX�j���8�	���lX`�g'݃-B��X����S��/z	��d�ak��T�&���w�(������c��W�6��g�~�k�E�:����7�~ɠ7��o���c������)��i/>8dm8�J��X �}�;H$D��><��l`��-/������8����\'�N~O�&��?�h<ח� k1��b�[�\@Oc�Y4i�f]Y2�2�V�$���!����;�^��a>�T�:v��M�S�2jG$!mƘٛ\\/\�M������)��~�w��	��i-�&��,��ds�lZ��^�Y��I6t�������G�OK�`�Y��.�`�GZ��ɣ~w��+&m^��F-9p:\4[Ҿ���PߒG�O���(o�,P��p��l�	�,F�c�	��~K{�s��)J���(�bb��3��rcE�����. ���5G<DQ��s<��p���K�[
�q{3��*���Ue�37lڈ*33l3��q���E�}��;���L=%lVZӲ�������Q ��|
jn!�7�����U&��(9g�]�i}.i4O�4^�ĳ�����_p^��8�Un�r4O|}�#�K���S>Qk_4���T�G�,���(Z��Z������9i_m��р
�:	���D!�d��!p�m}�-���d8���*ً�ZG��}���Ё��������^qCɜ��%.t�����E<_�f�8�~خ�p�����[Oq(Ͳ�9��	��$��f�?����Q��1Zc���Hi,6y>�����P��V`
�i�vZD��o�g��i]I�y�j��
:��T@�ץ"��|֪ؼ�dBo	f����	!D���[C�¬�N^��J�!TRC|��{�a�bf���\�B��͊cč�z[Ь;^�ƮEb�B�M�W֟z��;��R�+��k��~0��U�pb�� 㰕�( 6D�|�l�e���`_"�S��1��K�hDW�[�"m!p]���W�g��(��P,��q�q��S���1�JD�".�{�^������AR?U���g�_�H�_P�A�t/x �0����7�'�hfi�t7F�����I%9[S�����Z}{�Wt�x����r�s:o�Y	(S��W��KM���)������ٝR� |/�8Y$�P�u�[`6���L��%�Tmil;�[[��Oeo޵OnU�2�J�OL�V��@|[���0����K+����|��r�u��<z�<�^[G"��q��	Ñ�&�,::}\Ȗf3Ms�^Q{�Z|���?�X�V��4���6*�Ȕ�������/�ha:��A�g2���t3
V�
�!��IO}D������b6�$�}���y������u�={��˚%.����fR��'KB(�_����2�ma��c˺5�nh2S���_�n5�ɽdٺ���`Z�0��z1ً��x��+:��(�z��DR���Ho|�0�n�Bc�b��L�_�dN׌�[��#�A">��UB!�;�׹D���d&p�]sz�r�I�Q?�!�a$���l�)^��[������	�Y��3 �K�d��~q��˲�����oŽ4'�J�ԊM5�R۲Ca؝��@x%RF����� [�4������g]����p�9�<ݺ�3Pڨ��A��e����c�_+yφq*����A��MQ�^���nv,}��Ž�������m.�^�*ш7��+j�Y�����c#�n˵��%�Xdڅ>��%_m �q����'݃n�J�E)���s����O�ᬤp#)�;���{�c�%����B��V�R,�v�2��l%��?}��c��z��$��ɻVH�u�CVQb�.��w����(�<ZCL�����Gd�*� r�;�k���I9�r�j�
1ʓ�P�r��_��M��t
���W���k���x�B��%�����V\������SŞ<A�7y>����xc�����C���B�S8��?�О��>���=��NKFG�<I89 b�e>���������u<�-��0`����KQ�L��)�j����5Qjqc��M�^B�c=��2���lhP2�_ 3r�w��1?�y
��e�T^���̥�#n<O�&8�m�>o`k�m~��x˂(-�^�e�£�c�8,3�����tsqA�E�"��u���I+9��v.}�����r���kX�&S ��y�:�p#��}c'���^fj��P�j��A���T��n��>�S�p�$0qJRt�� 0��y�����Xl8��u86�/��RCh�����W�>������X�쮱����-��K�F`a��U�����!6[����)U�$��}�}r1W<��a�Թq���E+:�Z� �if����Z �i0,oV�9�*q��f/{�ؓ�$�$\��zsl�Y��Ջ?dsƏ�&��7���Yc�����Qr��$@=)��@�%}k�	|�M�SJ>f��T*_ _�!n�RM��@��P���O�T�j�.V�"ڕ���$O"vT���9�ȓ��� �G�A��)��8h:�ϖrT�ujB1a�6���8?,+��6���hO7�UG�ޖ+�����gf�e �l��5��Dz� {��6�aNV"��}����Cu�6��+*$z{�p��\����u�W+6�Z�4{<�/fF��FbV��&�}z�I�?��rL��OU�tͨ�K2#lM}����uA�!�z����i�f.uUd��Gp
75��,�B�����'qˆ��'�sC��W�0�f�[3����`s�_`A5��"9՟�۠q��;���&����yc��SlQ'��`L�!\m�$mmp��e��h\�ۙ���qb�5V�i
z��3�+��I��l?�ƌ�����Ɩɭ�Rr�3N�1��g'�6�G ���~W�V����=���	�r@�}��9�l��b#�}G2����O�O��qo<��t��~\%*\e	���]e�Ꙡ»y�<MIơ2��2Q�`�΂Ptb)!�'to�eod�~nu�����Vŏ�x�f'a�?OY(Jd��ƘI�� �P�l����U�&�s��ڇk�� �F����أД1�y4�7V+�2l��z}Z
��I������Z$���y�.V6���U&[��H�_B�\/y��׫�D���7QٮW?�dg��Y�̗��V!��D�g5���_�w�C1�����2�Mz�����S�0`�����d*���2��g��Z�t�="\Y��� �T���J�z�?f�,�b����p�T�
�~�ה�P>��*��r�d�\�"�X
�3��+9t�a�����Fu�bΠs��+" ��#��`^|ݸި�d�SH�Q��)���βr�* 3U76	�p�/v�c{��+��g�ǰrG��~'�[Ŧ"kX��ų�-������= ش-[9Uzz��Er�t�$�����;� [*M砝x����[WPO���7���x���t�@�3e���e�rr�#SӁ�%}#U%�-Q.��om04�� g���6,��\E���Y
����#���ZD��d;�Z'�ގ������g5�o��!�������M���X.��n�?&�&�L]�Q�?bS"Ci��'���a��x<rm���@^�����*��\��.[�a`u!넔�NHY.4eb�j:���xi�P��ӊj����Sކ=2C�1�r�b�e6���y��~m"��O{��k�	��[���4+��F�z���b��)U��o����E�ث	��tJm�O�y�12T`��%�vcJ�����]j_�2��6I�칝����06@�/������]wWR܈d'��kJ�C(\������!Kq�d8l��;s/��#\� ����@�j:��:Z�s��\���Wtɰ��̢��#n�Fc�E��ֺ���cHE�	��*6L�ف~���3	!2\��Q�<����a^�#،��� <DNI/�Y�#��4�'�!$_���^ۦ0(|� ѴN�� ��r�[*�X�&9���m+�@�t�!FN�1f�ǻ,���Ґ��{O���f ���<���Aw* �
�ϤAO
#@ɭ焉aÚ��d9���o��*���6�%�_��j����>��c��#��!׃���{|��e�@�6zv�^��m`��_"H���w��_}��X�)q�N�B!����d��?~��-�dYN]�dsg���&��O�yx��Ń��Eqx5���3d�Χn�P`�T�q���^q}��ބ�R!sۄ�l��E�����o��`\7�^�k�VeP�Pj1|�rj���[�9��ya��,'���p\ݢ��:3a��6���W�VHDS��˩��W��(�jJJd�@�'������V�x�@��ATF���|�3�:1���qcw뭋�v��-���3�=�&C� �f������9{9�c�%�p�3,�I�0w�4�"n�L�xév�"�r'���_�!-���"V+���&`�h�:+"�Ţ�rp�1m��	�l�e���䘜�te���5��sE�������E�4�֓�/N�	���Ѭ�$[=�{1{,��ܗ�w+���If|Fh��$jl�7�~M������-�v�+� I	��ki����|��W�K)���S�}�qG�&��k� z����[>3�(a�� �
	���C̝��(~������_V�]ka�H)>k�0.����a--���b���~Rܞv@؂�7�`�c4�����G)dh@���N	Y�f����>��6Y��},����?�2r���ӧ7ٔ���$�p�_��3�j���;�_pb������A��ۨ9r�l~�.�'����s��q�e+�T$��<l��Y���^>� /Uw�<��q�xPJ��r{Y	�%�;v�������[���8���M�'�Q�a�������J೫��5~�UO�v*N�L�9*n �Z�)(i�>�]��gi�es����	=ߔ�B,n�m[9��Y���\��")P�8�PL�r�ލ�C���E����6׀qskit��8���ƶ6�K���?�at0��WShK�����.��MӬETͰ�c�@a�Ң&��W%�B����E>����@F����>f鸖dL3隢GF!"���8
�P�����$ӯRÅ����%���[�&������K1kPm��E/���G�1�H/�&���u��Ɋ�����#,��Ȧ���S9(���Gtx}��Dw9��J�ί�y8w��a.!!��&���Tӕ�֡��!^�X_�	Fi.��<��kN�B��e�%-�/g��T�z�ښr�i14�Ŏdg����}B���><���RE�j3�gc׾7�zєȯ۫S���z�TҩAO|��T����;�MmHc�ד�-L�Gv��Jצ٤R�!�W�W�[��>���y��͑=p���u	��-��{�	͇���Mc��l0
�q�У{TdD$��ЖN!dl��+�͛��Ds#ڭ1_fݾ��i;�_S�4��:Kʳ!����Ջ|u�H���@>��{Ƭ!�XU;�K���gs8�h]͑�y��  �m��]�c��K�������-��d���8�遨����HN��|�_(ۇ�*Q�l��w"!,��RZ��L~��l�j�7�,�j�JG،BJ�&�m�8���������6o�f���=��n(A���/�����P,,�a�_Яp6�#���C����@s/s�oPuv�NÅ/S?��/���tq;-�S���(D����! Fp�X��w���Sџ4��(��M�P�W���7P��X�;^��I���q4\�ZW[g�"	���ڷ�[����=� [����Ʊ�{P	z�$��H0�.�w�/{�e�7�P��*w<�/�9J�``�͝0"äYd_��� �PqJ�7�nn���Ax��B|l�`X������u�u<��އH��9(�KgU�N��B�o���4%���iW�mx���]<���O~��&BZj��>yg�rF��ݶ�ߌ7��½(�cF�y _�&JZjZ�	��bQF��X#z��%Z2��c�\��b�h9a�L&��{��_*���+w��ӆ3m`⤓�֖&1,�5;���L�w��3���]-�,�
+b�+s�hd&�p��`8�qO�e! ��6�*K���������Y�}���٢�M*zO�\��J(c�C�a']��N���N*�H�S;V9V��2��vߞO�X��%&6D�zB=�� [�!Œ����Az\��H� H<OG/�fm�o,�|"/]�?����4��8�♢2h�$b#�����~�����y��Bz:pd$�:�ƥ+̐��q�t\6.��]�4? W��:�0��F!V��������:1���������:`��󟩢f8{=�w����	n��� ���: N$�aX��ή6��WE��;��܋yA&9�-d�Lcۤ\�L68��B������M����C���q���[�H��Uf���Kn�e�������L�q5?F�k��%"�V?��J(�gO'}m�K��6 	P�|pRN�#d�K;L��!�7�qp$�߄3��y�y�n��[�[�&�[��3 ��w���1&#�������CI;4}/JsW2�7O*i�V����䀯@��|H@9sT��x~�9;sүd1�R	3<�R	�����it�q�+�&�D��h��]?+:Rm=�s�1�5/DO�N�B�v���e�
�!+t+��뼆�F�IꏖD�-� ��H���n^�%�^I�Q[�6���QH$�0� ���IE���x��Fs�c�Mj����Z�lc��^�x{�h.Y~�ұqAM�E��<�SK��~	�d1v`�"����y4H��}��YLڰznFV=73ͬ��-�x>y'<��T(��Y�b"h����Y��Q�5�WS6Fqy�G��׿��#:�;�Y�}��Q��\�R0����Z�'Oo�a�8@���rD�P�^�RaG�96��j�k%���,$&�R u�U�3L#� 9�3�ԟSE�Ɲ����>t�M���g��ǰ�cƯ��^�&F�zĊ!ȶa��vi3j@����O�e?O�-�<��A�wifRȻК�;�_���V�ے��}8��]�@����B�{wG�\���mB�I�A29�	�
P[��S1,��;�/n�y#$΢
��p[1�]��T,�&��X�Z�5ui�(g�����������1N��Cυ2�{�a����
�-���i�W\�tb.��!{�R�֍Ѽ#���6�Ɠ#�6Q)B�0��Ļ[��Y���7��L�� ��|Q�����9D+ \^�4��(P�'}��2�w-~:e@���R�[�#S(�=6�Kk�5�Xj0��vd��`��
4!;?�V-�9j%g��Cr�_��5Z�ᩆ��V���H��ƈq��46Yإ��!Yu�TG�zH��K�lFu3�n'>��?r_��P�����_�P ��S>y�kϙk
������*@��������vs{��Ά�77fF�р�.��5�����Y��!
�����d2S�B�3�^3)٪��W$�jWN^e��˚�@����yz��C�h�^�#���9p�d�˨�����tw�e��q����Ŗx�֠��-[�穽r�C����y�����
�k��b���"��$3V		������������{KI����{�vDuk�%B�T�W6"驙Y;���4g.Xr�� �e�Ҧղ}�C��׷X=<W�B۟CG�9=�:ϥ�j�%7=�כS{�$�<[�x���j�������>�|�&�G)��Y��!��nòjs��o ;�t{.8�<��CQ?@�p�Sv���$]�&M�7�-jq4��;�$�N1��AѼ��Ezʅ0��;yŧ��:�H԰�)KZ�ٱ�;v��
��~�(�.�l�eu��)xhg�Yp�L��/T� =ᅀ��Oz�������h� ���z���EG�Q����G�q�}`�S�k��R?��ܭY�Am���Q����l�/�'P1��Ͼ��\��;���KA�2�\�*~�C�K����d	��5���A��?�JE���#ԙ����Ar,����ة�<�.µ���U[��۬�|5]�:��6�0 ��X� �C��c?P����U�y�Zg��5��	�Vɐ�8�1�/k��L�����L,<.WVQn��ֲfCE3� (dN�R�z�Ү����2�i�Z���_SNi�;��l�l�5�х>��.���R�B���^���0���;l	Nl�6��a�]	�E]\��b*H�����X���y@�?���"7����r54�Mm�_�|���B��?�����v�����g��ZA刓?�8N�*r<�[]�ŏ[����T/9�4JAH)x_�T�L��o�}�&#��p���nؖO��.�)/�}���ߚ��t"�n�x��8���.VOl��@/j�,\Ւͅ��=��e����9�;�A~�S>4?uI���خ�'������PV>&�e�OjL�����{,�:���w�u�I���S_�"��S�ގ��2�Fd�,�m �P$�u/�5�S���$Ъ��%CK�+�Y�4��2zPҒt;z��v�!�8KLp�����c�:qs���O����e��#�	p���%�u+٨z� Ԩ�k��y���ړ-T�k�T�U=�q?!�e{�m��i�iA�Ȍ%�#�r�4�������Q�%x6� wj���?9��t��e���������i I,�s��W+�E�t���/>���T�^��}��;��I����G�����ҹ	5{
��l���_�K	��,�g�e9�6�҃Ͳ# ��̥�������y�Ѳ��=�G��q�(����qm�����׳`�^��`��L�ȃ(F|zt�j�X����C��wy��En�P�~ׯ^�႖<7�*��a9%�Aگ�$`�J�ÐU�q��k�9&��]�6����J�Ȝ,��L('qd@���/N�;_��X�*^s���׈��g����ی��2�;^�Y[�_�/�ZR�B~(�c3�mZ�^�/;���T��9�Zø]4�+��~1���S������ ����W����B	��7YN�����-t�$�`r�L��H^��0)5x{�Z:�����Џ]�'w�=��>�����/�<��^��:'���ȷ6�\�E��7SP� #�f�U�Y����*����X�o������Q�H'�-���1�I!���Ww�1#M�
������O�`&��PX����ݝ�҈u����k���,���ĪHH��[�鼪�3�3�w�3��&��b��I�x$RGٞ;���:d�3bB�˧� ���	��B;�	�����\���[Ը.��ra��dO�g�A
$�)�{���}y��(�DRX��y�wZ�f��8(j�̌��.�W���f؁��O�>#�j�CB�Ȉ4?U2����`���
�K���A����E�t���,�/�~�AZ�_�іW�S� C�-����*��B�{�?��``�w�gu1ɤ��jl�kI.�0�9<g�M���O�R8C�Hb�S�f ���Vf�h�ca���^N��7<C��}6���k~���XEB�J�ɋ��g�zՕ��玔�ݵ@��|L��G�f��u�3�#n�C<�|����/��Qp	Bu����2��R	��_�<��7I:�+x0�K.��v�M)1�8H�0�ɭK����� �
e,y��d�iO(�Ɵl*xu�ж��������>?��r>���d}K���2����'"��"�i%�{����k��$bI!�5�BU��L����E�S�m��@ʉ�m�Ԍj�E�raku�n��>��O��}����'8�.��Hn{�Rm�ʍ�&,����CO�,b�@��[\<.`���)�^Ŭ��.\��2���PI4"
Jo���%"r?f��2�i�Ī�����m�g��~�I�5���mx���}�$ݶ�p
�1� n�I��)��$�K^�Vd�By�r�/6���6"�q��X��pr��n�\(7:��r��qj>r�dX�H@���P/�+!����*��OV�m^��e	��H�w�Rp�*�C0q���7������T���0w��"�4�8�1�����ʤ�=,��%[H�y>
0����t���BW%!�$c�ѯ�/�n����Z�)�wM���/����5�!��d���� �Bg6&����+C{�3��9W���� ��@s������'�H�9}�)\_�[ٞK0ZO�uaN#}Q�O6.Eޞ�<�}����������	s��u�plq���[ �!"
Ŝ�	�� o�1ͽ�T�Z���rq�&���y�E��P٩Y�p�����3����:�"(�ZR�1�Sk5)������1��*E�/�P�JJg�4b�(7�[LK�s�+�t
O5��L�Z�ﰓW���Ap(�ܘ�g��*Y��g�[ܞ�D�m �ީh���Ô5�Q]s�	5e���X��Om������,a#	�ZN�J3���� ��Q�8RI����I\��?�yk���l�Pʒ�~�(Vt�#�ؿ���9lҳ�ڐr�J)o��:V�������Q�o�PF��Q; fRT���G1JbF��a��R��2�W�(�}�꼞�H۴ҳ���ށ4��QǀεV��b�+=��'}btW���~>��1B[�
@��U�3zt�wlҶӾ��Zkތt����̭r����ikBD���-a��m���ǖ�(��z����S�������O.`�n��~Ř��a����q�c@�YQ8ygVp-0�`en:�4��fZ���A�y�3�H�di���d<Ծ߇Џ\��'w���2���V�B9eY)ܶ�hϷ��]�z��oKz�Z\�Z=:��W�d��}���� �cY�
�moQ���.�̓_��yu��J|!|�э5�P�rҕ�G�r�z�WBÂ?-*��c�e������r�L�{{��!�85�o���xE�1�,���(����佄�I����o?r6�K��=�[~��7�:h���� ��¶?S�c��m$���2g�=;S��>��U,=-�]iB��0Ұ9[TKbb�����a��7T!�O���D�:΃T�#���q�~ft!ڰh	�J���$0��Gy���7��6� Ëj:	U�l�CCĨ�Ax4QIǡ/�9��|㋓��ذ����s�J8=�/�߶AER�o�����s�OJSۏ��j���2���))(7Q��"��U+�pt���	�`��/��o��L�zwğ~�!yΉ��!�#*`�U�&y��t�N�pb&��l��J�B/�寣�g���=�}L�w�aU$�Fvڭ�^��['�R����S�xu�sY����~��	\�my�N���DC��B �|�袾��azv�<�0��恅L�AV�~t���q4�_�q���~!���yw����I����$�{2�2����L���1 �g������#�) ڏ�L4��DXf$l)#��r_}t�,��Yd�nG%{W6��T��4��K��`J7Ä��<\���y7�8�d�̤H�Ҩ���"�Yѐ��I����tL�S��#�%w��j۬im�ӛ�<�L��G�y*哜QǀSLo*}o^����e!�$��$d�Vb,��'����v�� eF��w)kޖ}`t��DR��Z�	,I*?g�K>D�au���p�9	]SD�����/������O�7�ɞ��p;s3n3���Y����!ndJ�F���Z�}���x�*r��]eP۵� �
��!�X*?���&l}�nP�ڧ$:�ג�Hr����*��}���^Bd�X�`B���n���u��Q��?���0�L:۪E�4c,���D7�kK�Ɗ�v�����P�L�۴EQ2y�פ��y�n3"����s2Wo�[��	���*_Í�MjX)�?�n�v��
ݖ�KD�Pv���%Mj&;@U���Mg��H(�P�ɟ�q����3ar/w�67d� 8���8F��E2]�٤��N[�QW	���˪{k��� �<�B�b���o����r�bX��u�������aV����Z�/�"5#���=��[��J�9��E}����+�Z��k��"��r�HV{	� ҵ�$��j:�x�J ��{�x�
�����ƛa�1{4�� ���!�x���t����fh��nun%��V/��ҵ�n��ZSϠ�a(p�����U�:�*��ŷ�����YP* ���L�o1����?w~�l��g�_�������Oҽ��J��64}Hי=�2Ne�?@���,f��J����b-&��3`�e|"���x���$�hŜ��0��5�11�/E�a�cj�AH�0�� 5;jbm-���uVae Q M� >m�S��c���o`��N��*Mla)��
Ky&Ȁ�M��p�����|�XS��� �.���V�	y,�v^�����DeG@�l�L-
�2@x=����R�sl��N�e�����o�JDlэt���N�{z ��%WB�'���+�AX��.I95���r����,a������r1*$�s��`�(̇�L�(���I�~c�m�����ȼ��%N�E�m�p�Ǽ��r'�u ����VՂ�&�n[!���ߔ�N���I�DM�
�"�!�������F�N�M�ϩlD�$�1� n�N��w�|�������M���(�W�fq��>�%,��M<3�1hW��O˾���5sNͣ�+S;����ӫut�2	��	+F֥���հM��|�f�ïnl]�P��.d�!�&��3J%��'�i��&l�������L!n��q�X�9^�ʵ�&�N�|"bbkǪ�EI��K����|�?�1�����v1%�$gˑ�l��$���ɪ0���G^F��1��("$+��nz8��/|\)�RKFx�z��7�u�B�c�P|�+����:c�`8��n@�E��������Ӓ� U�!E�3���W���]Փ����qAO��RT���>�XY�U�r�ўq{�VQ.׊8���Bl�?��2�#ۈ;�D���+���Z�C�7�*$�+�w�w%�W���g21�^I�1Gp�^�|�%`��:�-Ŷ�����*7.��P/�܎���yFC^g���c&ݩ�KSEx��{��0I{K)��$�.���t�7���%��[g�
6=���syeY�h�N5�O��!�_ps�^@�����aE���r����.G�+�T�ŝ��Y��#D�3h�(=E��� ^l���L�-
ra�XB^�1�6��#X��L�U�8UjW��C�+J+�la���k���j�1�9,�z�12͎�C�P�$ dA���k�{�&���������H�>{�,K���߅����g�}�ǩ�-�~oo��a�[�&t���5�C��Þ���$ 5u�k`#{���g�OS����,f��\|{�^7]�UkZ{N[*I�����qyn����
���f���P�MF�~m@Z+����Qs�M�dSm�	���Ba��Fw@Rb��1L��b�@�x�L��.2�K�K�E90�o�ܐ|N�W���p@�i(P�i�L����(iJ�ޤf������d��Q-zX�KKo��E�kR=j��� ��+��"E}�	Z��qk�j�� eJK#��gN�]���@���e� S>b/�N�z&�F�4�g٪��KH�e��Ȇk��ί]��X��_��� D�t0�-.>>�V�;;8�|�#�n|ࣃd�ІL]��k�,��������񐖐��K�f�[B)qj�>ş�v�,9�q��l��-����F�$b�I����R���q�]$qj]%0�(d�=^NN�klN)�Wں���7	a��9i��O��C5��tה��<���2�Qs�������.7��E'��3�Dn��_���N ��+ા1�맜��Z�q��S^��8�Ixu_ϝ^�g�~���ױd�@DO�]F�W������ז v+5��ԕq�ڴ�d/w��=�O%�7�����z��؟��%a_n�ڝp'*q6zߨ�j~Zq��!W͂OkR⚚��;��BCϥÿq���\Z�xU8jQ7(�w ���>�B��e�Z7 ������/çI��"����Bb�>@�+�&�u�P*#G"��B�mV �5>�<��*���&�b8'�vA��q�I*l6ieA]�������IT��:�'fD�v�K��ݧ k8o֙C}u&��$2�+�yd���tӃ�d��`�L�%$�GM�������+ å}%�U� ��¿�������?�	��zZ�Z�r?@@e�9����D��8�Oc8��w�n⨉g�zI�&q�����]��݈� ��#�������<Ge�����g�ީ�������Rvcc��b���)�+/���������I��	��鋲��e��F8;L�h���c�jG�4O~��^���З%a�M�3� �]��夽kc��c��{�����'=Q+�h������+*p��9%��)E+%ʺ>�ˊ�'��.�[c�D��� @ӛG��1^��v�B�g��8�cjM���`q�ł{䯢Dǭʽ)�r��L�?86�L��H/NM)|,`:��0���b;�Pk��m���:a 䄉s�j��w��^�����U�,p�
�&�a�ZM6�%�����D�A��{��4K�kHi0� C/h�I:HnX���4�*�o
����=!$�J'�MQ�1��铧6���%��l}:�CE�v�	��j�^�/���ۆ^��{�W%��v��[��(r�CxvmLg�UUP[��uc�9w��e��\__�E�0�P٭�Ke;SQ�����^�:�֘��v��l����'l=�Y�sä��<V���J��f�O�y����z�f
��|t��hV�B��<�T��o>i�����y�i�t����23�<��I�a�m?n\��$Ȇ���\.�pl�쯤�e�t�{�Ȃ�)��l��s;e��	"b�PH8��9��h�5Bi	r7������<-��Qr�d���^�D�{�E�_�"Mb�=�R͛�ͦ�e|�~n�V��lȸT�����b���2����!hd��'ڍV��ҍe`+�	z�˸��Ȫ){���xD��0ǛK��XV��g҇�x��T �6'��8��Ve�ծ<�����P"�?���I��:l+fH��B��j��O�tI1�_3�8L���U��v��w�����RSV{���Pt��7~�5~p)�I�i���X���)�3Zڽ����|iBA���)�y����f���u����}��8%�X��c��P4j��$_X4]hԆ�"���]��#?ڽ��/˲����z���%&�&�G�Z-����������4u�K�+z<���lf��,Ct]�h+S��ȣ�i<! bU@��1<G7��wO3rbtỷ���iȬ؀��4�0��E�o
V�	8�a�[����j���d�E1�	+�Q����C��������_]0�΋c=7?)
���)�%ۙ^�A��v��\,�ZG�+h�ϚU3ܹ�������Qp�gwc��Z�ɻg,?��xG��k)t��/��֖%��������*��mkӔ�·h��zf�� �R��=�F��F��Fn�et*YԭO�cy2Dka���y���)����$M���gl��3�;~��%gD)�N��  ��2ϩb&��T��b��lH�!෈��\6���:�u���mI-c�WY"��d�[�]�1�K�C���F�������7���VnI�*|�:�G�U0m^��ۛ�k2Q�n�$^iَ��m�1�dDO/����Y6��oh��ۀ���DX��/��G�73r#n����:���<�N�:���a��;��?��s��G[�>���m��7R�r���%W�A�!B�$��C��"<�L8L#v�GCP���~Hq��{�|%ĺf��B`�߉�p)_>dc��x���9z��̠�&�I})C��̢!�Nj�T�	���AX��G�"�2����ww �.���z���m�
M,����(�����`X���
G��S�N��Q�#�9ߩo����B�J��AA����R<��5��_4_�	�v���T�iI9��X�y�>�K���b�b�#&�� �8�D_�eO�ǃ�>�N��1�/�%�ë��sVF�ɜ2�Ov�T-�p���ֻ�!{f���{"N�'2ZXQ���/KC.s��|"к3n�T��"�t������n�2k�]�R�]�8n��{��ި��-��ƹ�dSoI[�n'�y/��V�6{wW��%_�S2$/!Tԓſ\8{#-�&P�	wj=nh��KU�`��*��"�K��
�Z��ֲvsW
��ŋՖ����Fzʼ@��ǀ�E zN��ޢ�S�ZzP���uf��_�$���9�e��>00���a_&�7�+�>t�`#��K�5330�V�:O��La��Sf��朵A��Ζ�_^�C��m�5�l�yZ͞�h�<�t�����En�yʽ6���M��T[�>bx3(;T��$�6����I	�<��_���F_�|�u�0禎��KcIKpM��o�V'٬V�c����ڦA*:��PRle��>i$Q�^�U�� �\$�`�eN��=��*�%\_��޻+"z��7)��ʈ���3X-�R��ބEC�͘J|�9Dsկ���Ȃҳ^^�)D�%z�؄V�^�#Y*GY�:����z.M�^��X�&ڱ4���)����eo�st�:�Nl��r?N��\m�8T�:��/W9%58�݇�tﭕ�UX�Hx_B���q
e��'�g\H��8��)���l��X9,^7Z<حqBK�Ee2�$'�)�������"�������7��O����!HX|��l���}�_0.<>�<��)�����忁`�M�1{��Z\�5�Sf��p�eKBu��7|��$����1�y$�#G��F�wD�s&�~a�T$���hJ��W���r�dTU��L��W�k/a詢���C��!��Q�����t{$���ʠS�L�~��m�Ш#�$о;�ת���:�C��}/y����©��=a��:�K�X�ʸrg�d�e{��qTe����F��xh@k�3�_���g$�`�֖�F�5���N�h����)���u�ZB�P���&�+���WJ�'1��]�����m��l��UxZ�"��A����(, YzF!_�#�g?2UY�38:J	�F-�*[Ƹ-�F9s^�~#7~ˁ�E%����v��,�WQ�R�ڞ4��b�	���99r�M��s�.�a4��=�^)Ũre�:��M���f����m�yE���B�[�6��ǎ�C[w���S��&����HbL��;�ڭ��K6�w���������+ ����y�o�iw�fx�l��lA�;�L-
�j��u�|�N||�+�Kl׷�^�P��jnBIr)LWr���,����d����a2�hǻ�!d����bF��'Uc�K9��5������U��dKUC�&������^���Z�����p��u��.ؒ��h9{D*��lˊJ * z�OA�z����	��Rq/y�� l�����^�^�D�<����d���3QZB\���8��`��mA�e����\��Zh���Ic����CK��	�!�4�Q��V����V��>�/��/ɵ�i��]_�F�A�3ϊv�c�_��&3~�l@���+xǦ���.w�3����&�eq u{�8a03B^�SQ|Y���ߩhB�(+��J:x��
�cx�jH��e�F�Q4��g�u�o�?�؛6�,�1u����w�	��)��|�tl9�u��þF�|)pG�����k���>��>�R^��9�5�S�|<��u%nt�c������j��[m�M�Ł�aq�qE/JD�y�l��`|wt���S<rQ@�6�Y����2�u*�?�XgT�� 7�S����) ��g󴃿�fq��L�<�zj�AG��&��Ԝ�N%�e|
MQ��9��HE�e�m�����,-\v����5��Y+���J���3�T��Sbq���t�c��ﺠ��U&���� S�t�͒$��
Oi?Ǝ��
�H�����%Gڷ�u�w�d����Og��ԇ���P>�����.���y���0ݐr+ȮKH�~��P��W��ٍ�04�H���:���k�m 0�?�����m�(����ϾM���?�ɷ�� �pତ��Ո��D�A���8�*��/ds���	������<ˏn�J���:����ջ���t�P)��]�6��wg��7�)�.]͟��pދ��S��eˋ�KKMW��4wE&
&���>��)^��5�~���t2���*�Ec�:�'��ugIR=�z���g<���r�����;ܼ��=���\f���ؒ,*��_ɄJ��FDm��x�6Qe~a�eajS �U�;��w���v�6Z҈���Uu;�i�AU$[n�-sp{��(��%[	�������#���q��j��\�>�\(?�ϥ�5��q�n*�]¬S���"]D��"���(�c1\��3�}uw5��]�>9f?f�N氃Tlʠ�����xRPdϴK*�B�X�@
�z�KO	�0x�
K����*g��a�����.���ИR!�^��)�ůu?c����W$U�KO�G�}d:'��|����AJ}���z��\�O�;��~(^"	����ز�/?Y;��b���Z�2�[�b܀�J5+�f�������JY�h�T
%�I��NE%I��oZ�M7�1g��~k3X�\QƔ�L1�Ԁ�|�qDu���CR� R5�ٵz#܎�d��?�����~G�@K�B�6O�,ax�4g/T��H_B��Q_�A�]�<� 3���l-�Z��3&��������8J���۫��o�m:؍)�hb�˓��z� ��N7gb-�J���ф�������YXN 	PIV���܎y:Z��an� �*��_� �6#�U�wو���Y\�g��g�G9_���W���=\��$��]���(4P�B��+{��V����E��D��f�B�_����+�B�����O-F�V�a����P6���GH\��cp�²9s����x��$i6q�b���L�*���M-�WZ�"�Qa�:J/z��tV�#㌗,=�w3c�Ǹ:�8��Jԙ �	�.5��.������M^;�p}���a3կq��̺)*��Ju�	�Qs�yEoXҫjk�j�����ޟ�J���].I��!����T�Ňw�A\�U#=�;�I�����yEZ1#�V��6R�F& ݜyq�S,��,#�x�a�Ɛ����]����������o:��~*M.����ܱ-�?�̈́�s�H�c�SNy���b��J<����K�b�'D�iޅ���Cl�8r�XJ��D��,E6�ڝ��	75�$����	q�;ʳ��ҏ�6��>�i� ��7J^t��9ȔuM��A�>3�͵hm��5P��y.�Iv���7�t�2u������Ҧc+o�O*�z  r�~_��,�=�`|�'#���M��zx%���
���G�Ըk\o:�]h��Ze���DW��'�{?��x�t[um_��F^���4���<+˯j�K��0��?D�p,*�	�k�=.��_і�b�Z�|��W��[!��U
s�L��Vߢ���������j�c��{� ��O���^v�C�|���y�[�rx�OI���NHV�ƣQK����7�Z����U�
�x�i�u��j"��k�Z���5�:�4�ߣ%.��zY��$�HR���ܞI�z`p���J�j܃_���)3�EE�`�F��g3!���rM�Ѫ�;ӧ�d�kQ����8,����	޹Ԙ<Y6�ͣt�j�'���$q���4��y��sd�K0*�ch����d�A�K:�S|��}Z|�T�c��nz��k�B�e3&A��ȡ�%��M��#��6���]2�͘��N�FM"��S�a�6p��������x�R�	�'4ԗ.��95�	Q�τaNB�X?8���l�>D��e|W�	y�I����f�B܄��u?L��zsT$��_Ǒ(9��h��U1¼"J�k�s/�(t�(g�˥��J�c뼲)��:i����ӆ��$9��ѯ����$�aP���2��6m�7Q�m)���	�2,x"x��V*�'~����� �ʟ�Μ�2�Vmj)����L�[c#���BbwQ�����ߪ�ms1B{$�%��y��;��a�3Al��͐1���[{؂�v~��g��$�+n�0WC�.ō�]E�2�[���8(�`r�5�'�/��U��mbč�BBTY��4Ր��t�f��-gJX)�d܁m�a�=���y��};�)0��	�+�d����=]+U�7�<P�T>���Q�<w���z Z�P-�0�i�J�eRK�K�����LW֝��1zT��l;�,���/��l�����{N�0�$Ҁx�b����T O1'R�^�=|e�zi�xzz�y��(3:�(���1t��a�>��,��B�O>�g~��� �R;C�:f�����٪a�*]���ق $)�z�p6Ol��a��x�R
�-�(35I|�<�T����x-E.S��G�v_{�|�A� ���<��ha��[�����+س���B{?�IIE3E�hV�֘�ܯ�z>=��]�]󾜶��������z��c̓p}�g�K�� Lz�H��jE��	`��ŝć��CBp5����S��	j(f.%O�1.�JżK��X�c[��\���f��n �.�����6c\��|�f��,�C0�����wF�V��3_�����O��@4��5�v�L'��������B_��q�!��lG�a�!��,󜠺*n��%�j:3J+��Re�����$�y�3������.��^�-3dF�e;Vc����Ч�<|�/Sy�)��ǐ%��c>�:U�;r��>,�'&�����ox�������e����O3�� ��a���eH>�i��V>o�3=�F�"�?��;[���5��F~MG5J
��o>��\#�W�y�[��7�!z%�+&�cx;��˃}!����Х�?�e����?b֭��?RYn��ܼL�y�F.��2�zQרLg����qA�aA�������	�C�����z�l��iS��ũ���*�<����f�E_�0 �ۄ�w�t1��Ew�>0�7F�E6��ȧ����G�rK4BT�^�7�dd*�5�9�%�u��l�����ʞ��>0�
�����=~�	 !?N�M����)9$f���c{��r��;�X��1��]����kBTq^� �4W��=�"�B/�!��	-*��Ǯ(�1��4^?�ib5��4���I�TP'��E��չX�m#�!�	�)6�Wv���Ԥ�:�cqL�b :�b\�g��.�_,3�S���N7<��7�u��ב���c$
F�wqCn���5�p�����'�ٓH�/��c7������7)�_�O`�{��h�N�%.�g�C����P�d;��[�P��j]�=��	&����qv&G��)�ϛ�E��l��.�\�K�\��4��4ἩF=7JT�I���ǜ�*>@/ɓ�?�P��~���q�EV�5,�jf"�����8Ķ�o�U��+�	�C�x}�Ts6;�%0�����Ы�����#ٸ2��a��ox`�/s�RFy�P�o���N�O��!����	ծ~�b�T�����d��\;���!k9�������f�T��u�Ԋ�8����K�)�nk�>��[���'J��庈 BV$F�����2���o�����v}�~��DB���0��um��CO�81C���g���|SM�u���9��J
b��{�k����놾 \	R��'��"�iܕ�|�&����$f�#�j5�rG�@]ïב��'��u�O\��}����d�C���xP��<�#o�H��4�dFڣׄ��~��kԉ=쑌���Y
՘)�~���.Qoo����|���b"��8�`�n��y�p�@��ű���+�D���󁯳C�%Us��!�E+�3��oM�	��P?�k���)�
Z�3+,Y�|�($�B5Ȟ��;����5Da9��P���*�m��B�E��I�2:�n�eϲ5�f�G��>�K��:;.~�¿�1�Ǧ�6_l&�OJ�!�WF�*ԣ��O��+#Ǵ���f�6�|Sh������c'�>6�'��~ȯ/�w��GZyU��*D�tGo�u��jk8�y�����+ޥ�MFkk��)
*� T8C��FH�UՋEV53u*]��F-��k�O:�E��Gw;��9ϥ�e���F&���m�����ed��*�AY0Puf%@S�1τxT�s������~�Y�7�Mff��ί5��:��ҳ��Fv�;��-��+�j�X6�Ͼ�@eereIF.�=������J���RZ0t/W�
��֖(�h�ĳڻ���`���*Cj�\�r�^9�B���]�@浴���\���b����}���恠���=G0'��ֆ�)��ѡo.r��;���/�	up�i��F�+���?��E%1CX6��%I����x����5t����O�����u�9��1�'{�����|eC,}Ш���R[�X���&{�cNa9��^�{(No�]�_}�+ڦ�ʽ�Hb�+z�v�Ozޢ��+g�8���r��I�Cx`G�a��֊	w���l���!F,Dp<�❈�I_MA�|���N��1
�SJ�m)��O�G(]��k d1���BH��z��Ѭ¸�FUVOZ��Bd�f�av/��\HE�f�c���s�R��z,�P���5��W��NC"%1~�Ɛ�1g�=}TJ��jV�H�̶Ԯ&.���L����8��@��V��*���R��X�����,a���#�����϶�x�I��∬fhn���ؕ� 7k2��`+%. � ��v�,P�G��П� [J�G+���&3�N�Z�s���V�����?D�S��hM�h:�a�U׊3����#�5���,���6���1���iq?20�h ���L���2I/� \o�`�x5@H\YY�{���GZx�U��J_L�)fI}+B��X�A`�(뉄8&Z���2��MX�g]��Uӳ���/�����7Rd._:�qqX�l�C��<��6�bG���.դ�g��u�%�+��??
G�O�����p\�P�3׻e0�=3�&Wj���̑ZS�F�{z���;.���'l�N6���wz �bʹ_���V�~���#�Z{[���<��o�F�Q�>��i���>�I�U��:Ƕ�6�������d
��#U7��2/��/�Q������������IG7xU� ��H��Bt�-z2m���_G�eD��Y��?��so�B����#����38�9iڇWM�b�տ��*�m|֐u�mҝ!5F[Y#�  ����� eAaՀ�KkJߝ���N�p��Wꏪk�*����	�@��\�CMr�Kt��vϳ�/��ǘ���?���M^ck�������	�V������ߧFRa�>B:��]�+q�&��U�}�U5� ۡ���ZX"�h�V��Աؐ֝�W����'�A��/l�i%���nrPt;�閬[\+�2A�H��r����A�,7~7�D�s/�������bb�:�{@ˠ��k��<�X��"�|to,���J���q=�(5��ߑ�Պ�{~�8<�{l9��������
3dY����l��0]�����Ǐ��؇|�"n�$�m��[����O�Z��Q�g[O��+�ƥDVRo�_vW������>'h�֋�=�v*w�#[��\�7�\�XL�����QI��̓���w\�H��T�	�W�jj�� ������Ȭ�&\e�a�G�������Ǒ,s,J$����V�\�JD
��=��?@B�-���Dv��?-;��|�乄Z������|yU4�^c������������7bXi,������W�&BL�Đ�[�����E�����fq:]%a�A+�W�cs_H�kfp�Ire��P@��`m[�gQd�*>�x$�����]8�B㥚�e��I��Ցޙ�,�˰����0�T���a��E�CH'G⊵���!�vb�ś���T\A# �!)U�*�u�\��x��\ߴ������������:�n���"V��4zr{Ay��~]�G�-��>�FN5U�I��1cF�:��$���KYdŏ�	��Եt�[��LU%�_�Y�r�+�B�7!F�Xjv��+V}*�^<�9ݸ�I�)qZ�̿эڹ�阣�NA3�6�����!�ᐎ��^3�<K	m���&���؈��o'P�о�"��Wk��V�u�%ᚚמ���dތ�����IH�3hE�����2{�tt�7��@�۳�C&�r˵�~)���}�i��PR�w���Ké ��T&b&��.N�m�����B�ܼ�wSHZ<[IsT�-.��u2���y��XB����L�*;_[.��@B�5�e0*��B�i��;_SQ�w�Fj+��m�S}b�k�>��۹Z��@a2V4\�/,)G嵩�_V�%&�m��K�w�)�'K���l=�H�r	f����g�;��Xk"ez�_>>"c��3	G�u>m���1�AA3�g�!��V���䗙�EjF�%Q�<(��2����B�������7Sj�+�PA9Pj�N�uR5֮(�cՇ�b˒��~I���`9<2����;�b ����ڇ�)K�X�r� ��k,�$W�Hw��s�#a�עn[�X�ڗڞ���+W�b�9A�V?��`z�&ӽȽ�I�t��yZ	My��c۵��@���Wi��7(h�<�}�ӑ;5��J?�~"����s�1��#�\q���\�D�IB_��毉ӧ	3�Y	1�J$�@9��a��#2�VP!��Bv�̫&���6$���~����|#�x)���c��ym+���]O��<%�� ��Nn���Y��Yu9��J��)��G�~	k�"hg�섦�]�Xg"���]ޒ���u���B���n;�'�q!U��!�<�/�$3��E��V�����tMm�:�)���c"O�+`��ea��)�aܟWy�,�ex�}�v��( �1qò�i��(h�t萢Ȫ]jiӣB]n�U{�Y���h���������rpKކ��P[@)�u�I6ʤX%��Y���'�$C9N��6)�ƒ/�סzG�Pjz���hd2��{�jtT?`�ݳ��^;�*zv5 t�lߒ���TݤvG8���Q�?qfgm�ѿ��h�o�Ե�s-���yB��|�ʃ~O3�&_''���nD	E��J�5�E�ΐ7�y7o�UԖ�
-z<VA4�O5d1�t���������W�UN�3�W拄��!�H�o�x��D�4#����'&־K;VV���d���5��5����a���)�f�w�1WZn$�©����i�Tx*��O~2q�� nb؝��)?����Ԏ�S;�H��5�1�Ʈ!�#K��脗�1�r�bn��g��1��_v�����l��b�[g' �>rԼIϛdw������oʕ�b�a)�}���'��Dn?�[�<�0�����,���{:��m][�q�ob��m�?uq땄��ȣ�e��:]r���B�� �=�ZV�Cbu��� �][`lo�VNl��T�'khL����"NSZ7�˷Ů�9��3C����l(?qU�-?���J�˪v���1����11���[��F� }�a�����n�z9��r�I+뿨��T����M��XAYK�a-�]�h���:�i �({�J�|G�G���8������}=Vq�w�7*��c��ԗ�^1 敎_�A����AFLr��,+fqك�m٭��Z]?�t���$��Pi�7p
��T��I_�C��m_mO�>^��J�
/)X�x��U��\S$t�eY;g�0Z�|͹��[�2)��?}W�]1�[x�ߙ�[c)���	z��Ŏ���'�5Uh��t�ng3�i��P쎇����r{J�l���A݃�$+i�O�_��^�+���1�M�l݇a��VE$�P1f��z3Y{����X�&@S��][�� ����>#_�t��8r�H�Ylq}�h�#�q7#P��ޭ������}�;<�W�fn�r4���x���#�j��5��V�k�~�9`�"�h?������?�LS�u�V���R��j��p���٬-%)�K(�T��U��&�V�����#6S�8<��a,�7l��/�4�A��u{�@Dx�o��L��׹���'��Ob)(�:]�m��|��c��~�E�^ο�7�i�~��|F���~�8K;�eB��p�%֔�w9�Ϯ 3\�R�`����W{$�ǹ�-&�(�"�Z�9��{���M�L��D����a_��#ω�zg��l�����Ol1Y�9�k,���O��Ze�lH���ܼ�p6�.����/><�?�4xYu��A��*�$��c8��03
�QH#I��ރA�g~d� |lJ�<�~T���,����z[wO�o��K��9������YY��'S��:�O�y(Ӆ=}�k��]`�x8&��8�����<�	O	���2���J��Cy-���9���w�g�V���̫:n�k���jW�6��'�_7we@l9[�����{Y���P{k��J�~4��g����xS�F�E�8L������}*�K,�yvof����[Q�
���(c* *�l�
�W|||���K^�WR�ɍg�C�U��ݺ4r�p������@����6j�Q�1]^C^���䇥��Β��p(Img�?�t����8�������4�%Ö��=m�g��NJ��V�A�f���b(�����z�W$��5��z�����r�<�d��9XƶZW�C5D[?S�֝����M	�����Ͳ_Q⌤,�0���鿥~<��p���!�'Z�p�w�,+����dQ�%�uŖ(-@\�A���%��t���ИS1	���v�	����ee����##�mǂ��nOU�"�'���]T��O/f���R\tn�C�fA�4����������U�7u�'�eS�v]pfa(9�J|T�m�����=��D�b|����a#���{�Im-ľn������
��"A٦�����N�T�U�δ���_�@M�Y���}b�Ȃp���D���y+U�9���-e$ �2fF�!}̛B�S�@ᕬo�XRC%7�U"y@��J�T�����0��܍=�nD?�(m�a�_p���r<-����S���o#���g&�c����O^�[�
*�z�"bf���ʹdA�k��LƝܘXʷ(�-�)衽�>A铒�� �O�u(���t�����0�Q�j�AZ�<ڹ�ӚxZ.O��R��~���l=�Cl0P�/�}�Čf ̐��/#��(��܊w.��Px�`�b�ً(�)v�D���d��S�	�,%��5I@N�N����O �hu�a�0��Zw��`۳~2{���'nC��,��0^J�-�J���L��T�b���g-p}mD�j4l�G޺I���g�X�6_�p�x�E`7�J��	�L�
��=�~���_�b�o��ג�x9��վe�*�����ş����v�Y��vԵ��^�}9|q�i�^LpfT����g,@���l��h�1�G�#�J�v'	�S���>C�z�żO7�=q�~R&�	���Si�	���qQ��!�n� �� �����#���4g.��e�h1Ɛ�,xҾ�*� *һ�\�Ԟ��%1���y�ߢ	<.~ ȒˠK��L��H2��pJ	 Kg(���:���ec�\C��]�
�nm:�1�ZM�o^B�NX�_�k��Je��R((+�)'\h�y�;��ً2�MO�Â�NbMH������ɤ*�q�!���Pd=����"��;��9f����BFM8:�����%os��#+�d��_?P��G������m�ݳz�3�����Ow�S�i(��o����e	�Ks�#�!g~)厶���n(Y���r���g#\X#���?��@�FC]�V�v$����6/�͢C���k���ڕ[����u�H�-UVҀ���O��_���[���Y�z��eo(%��p�I�z��}�ۅ�sX������"4�%:"|%�2?b�)��y�ߋ~M�"�h�����.�t�"�>I�R6�p��3�R�����p��Hi��y)Y���'n�!z/������l��>�tꈇ�xW��4u�F��7����]z,爃�CIy�f_p�Q����A����`���7�"#��:*צX�8��m�;�P�j��
QRbzC9[�Ƴ��7/Gʅb�fp�o2��͔9븏p��>�5C�'t+_��-CPs���R�8[hz��@ۦ|�b��(o�G���c�8�i*�'�7�it_����G
�w��R�w��e+��ғ�q�-R*��4	翯i�ZO,<�Rx�8jOLJ�ܰb�S.X
S���T��X(x�]�)�A��`�'g!��l���B5��.e�G��(0�5��K����ň���Ykz�}���a89$���Ç"�j��{}%���ʧ8i!C*4��"I�oN�ӡXxb�'��I_\獮�1�@�
��;*��:�|���>�W  ��ws�8�4�(-���8���L�E�ߠ�tk�!���z��t��A,���d�]3d�Q��*?{�o��1���O���V�vV���6+8|Y��aZ����c����<��=��-|���U5<���7Sl�_N|=�f�F�*���x N��<�V�A	4�G]��ێ�{�@��o�f��f�s>0�o[P��.�r3�gy�3���v$����ԝe���+R������U���9�V߆̼n�Y�#���;�"�i�W1��W�D���&�41-��r3�S�y���b������KVa>|���M�`�f�2_9>�U�屑����E���?Z��T��TXqk��/^[������.\m¿��%Z$U	�9E�80d^Z�JѼ��jb�`�����=�d�AW��OQ�L� �U�cy&���SH���� ������,����*��w[���6�z0f"�q�0�':�to��o����(#��m���aN�2^�(�0���+J�KP��X��Z��x��*8t����WB��:�y̬ 3^:�Ո'�0؇�s����,iv¹��k��3�%��]K��v��˨/��Q	�U���W-<���W����QO�`���B��ЬS�ݑ�9h�j��r�]3�gi�l.[�5I�է�ː��%���m��m�,�6�L�31�v4.@��x͹v�!�?*'(��ث�Ux~ϚAˈ�l !�r��kV�2ūEM��By�����^�C�>j�t_>uF�rC�f����ĳ$`F�_��(�Àkt)F���]����{�!_���ݭu��tB_#v��x��̲E�e�t��|1��G��~1uN���4F6����˕�l2ý���8 ���d:}\cfZ�K��H\w	ܶ*Z~�HȫA�T�-�5Wʤr���0H�v�b�]سUa�lg�|&���һ ����
cy���:S��r�S�˩W:ȟ�%�z������g���`o��2`�	|�6��3����Z@�U"F�G��z��Ϡ3�t	�����C@RoQ���[�3��!v�Xx���ɶ��`��@<��Uy�i]�M�;ػů��b�Lbד(�F\��a܉�� w-�o&Q��2��{�
q��w�q�D8���1���E�lj�¥,"��E�%.�����	
��&�T(��8~�����O	2i[�L���M��l��$�s|��"��JgS ������$0�LO1�w���Q���*����)�A�����q���Y��%�j]��L�;1�L��40'�]�У��ͭ}�K�1�W��g[T]�xeG�y�Z&�hD�?��t�p�t�pr������?�����'$Z".��*z������/6�L>�B���#��*�*��:���F�d$ه6��M�!�����D�A�bQv�0d�m��m@��M���������0�p6~ԥS��,��`NhU�y�7�,���φ-�N�5W�%���<-�B�O���
U�JV|�ӥVW�؞d�n;�
V����gѱ�C6ĸ};cl�V�Y$�6W�3�9ֈRG�����	g,y̔�Eϥ8�0���11&�n�;ν�-����j�����h���b���J��f��A�az��\�le*%��jψ���ئ���
Kb��C�O+�T���=b)Q�j��'CQ��Q���C6�]L y�'}S�"<xY�Y^���0�'.Ci�d�8�׉9�|\�k5�^��i*�Md�X������mX�q�g���>��8B\����gn��zp�d���s���c�=�-�2�k���΂�US��	�(�Š��l��U�(I3������Ip�TS��] RH��f��-�A�?>	��9�/��OG�40\�UW2ѯz��T���{��	~<-^?�i�3��B1Yh�D�ߐ+>�_��mwӜ��Sc��)��J��<B��0�3�,zsd��F��}��!�">w9�[1�]���p�%�������{�WwsS��]T��]���^�%��ŷ\�,-�����ܺl�T��6y��̌J`����*h�!��D�{Ĕ��)�i�Bʯ�6y��K�V�@�
����d�߹o.�����	��U=�*�3<8�������V,��|��c����[V�s�WT܍���40�6�LyP`|H�Q��W�;��JXmCvk&ɦD����G��PzJn㰮�R�#���{�a� �$���nN� ��C��2����� ̑V�֢:��"Z��hK�,���b�2��\E�Ȣ��U��'�����C���C%v5뾰L�<�B������-@��#��nB�ќ�xx0����ε# �Y�Ǔ}D1��4�Yx������9J���F�9/���2��(8�����i�\�RR�.~y�b9�
�ǐ@^9B:G�hXP�M9��르o�%�o����&ӌ���B#4�R�=��K!���.��F�+H��_�c�Q[?����?�@�ν򐴽���UVNn�P,���*�=���L��&���gH�Nʻ��-�9�b$��=ƿu7o���N4[�Έ%o/��������Ϛ���S\"2���thc�"�]r�	NC>|�nZH�Z��5w�/"��c��ɈOlg���z����Q��ퟓ\��eIu�FgF����C��&�ff�`�< n�8�"�����8M��&&w��%bqH?7"����qŪa����d�\�7Tщ�E���R���e(�C��_�p��v�E���P���L�w�.�_�V��P���v�q8S/Eq-��X�&�΁fHe}6*�{�bf���Eᯁ4�f���b�����&I_��C0�mW�m�I5U`��l�
Ce��x/͗(�Q�����#5��ɗ�}R`�u�A��sm�����X���3$�M�.ր��;��lJ���p%�ߥ���;�׸�E���As8������$1e��k$��������I��Dv|��1����V�j��9x��z0E��?Q�z~����f��FرT���~�~ޏ΢%4N	�$&�u[.ĝl�����VS�>t�%���B��c}�׼%MA�V
M��G����l�����$C�!��G�5VWLA�����i��~V�&F����+If[W�v�U��RW^��;����,���U�s\ػ�  P�gv�^��W�_1#�\2�8W�1�W�$���x��N�	�V�Zv�j���Y���p�ϺtDG,y�w8�;7(+{�x��W#�eK�2U3�#:�T�_r[���/am�|>_���^�|Y#��{xH��<0���q��.56e~
�$θ��m�d�x	ufS����Y \P��o���6�=u_�h�������{���3������[���ވ�Q�w��ȅ㼁p��#q(D�n��GCr�|s�,I�V�J (�tn��-Dq9�H،S�k
��ò�Jk�{A!��O�3�4c>�\(��'IX(������(�z�����l�+ť#��dT����qr��!D6�iU���en��W(d������-05A������f�A�=¢2�)�odgd8��ÞM�Ž
����w�f|+
ZU�'�Ђҳ��u+C��'�:w�p��&��ӏF���)ھ{b�G&�I������W���⏁���z"���)�_ք\�ˮu�{4'�Ww��0��*r���e.D�����Ru[�9@5�E�p���6\ڊ��*4XV)w�������F�_u97ӽ#^�˪H�=��	+�d�ڀ.B�S/yg`t���k�&��VV�D.)��s͍�F2���S���>x�v��_�kDK�v�j�ؕc$R��J8l�qcf�͘��B�8�0>Bs�>�Ho� /BȚ����"~G�E���0+��q^����=e�O�>����1t�V���ro�JQ������f����|��D�_d IH���oU,�d4㐙�?��h{Em�����8"a�=:�=&��4��C$M�]��Yl��W&7���0 �vS�Т�[2Tn��p7��!�X)�ź�X�G�Q�H	��J|3�j/Yڢ�֚�?w�U���[�����<�=M�f������T`���X& ��c'�Q�uǱ1^y��
޶qk�"Qg^)(���:��t�V�&T��F}	�����m���(�v�8܊9S�Kg��;����L �Na��v���bhtB_�Q�bz��D���1�A�}\�k�'���C�k"0�"�����5�3�+G͉��[n���x�ɧ��K��e�h�W|3�L>��������,�C}��6�c���X�h(
<��������I=�{>"��q�Z� W����ɔ��8���5<8��ov���i~�	f��_����kv��sW���^� V"/�_dAEw፴������j�C��Z��->,��'HzwQ����������`�c�6鵡̾����(�tLH��N4�쟒�rI"���s����^bIJ�5r
Ĳ<?ם�2}�=�=`�u��4��T70���C���m�:��]I-�� /[i_�s7�Sv�wձ�69E_f7�S�ٽ�__��pc�kU�>�-���������A{K����!ʑ��5\�'J�����q��TaN�{�+��]v��ݾ˶g�B^��l���}�;�;|�Y5�i�Z��ף�,!��=1ڑ��[,%�e����-�I~1�,��1�3+���!�jS9.l*�6>d�8��3����KR�@q9-y^�|8th�T�J�TWɂ	u F�!��$�� �v!�N�j)��'�כw���s����xS��e@bn��,��`P��w}A|X!���0��?�]mN;��|��bV�+ �B)�E�Ɉ���M�8
�V�I��C�^Ls@!w11eESJ?}W7�!�{���VF����)�����U��=[)��!��������!�q��.���@K"��r���_�j�5
�Wj�D�taB���>�9H�5 �h��u���3�)��k���6b��f	c����Zw�)̆�SQ�Ӯ�@6���q�U������'��/`R~CQ���^s-?�+�(z3w�������տ�d�2���r��o��C����\([?d0�(=��7�V��Y5���p�V� �-��
ʾ,�9��Dg(J�-�ME�)�$1�]� iiӬ��Kv��Ia����	�����OEC9x�ЏN	.A夳�=�1_�M��>[Ƣݬ&d�  ����~����6�t���=`��)ц���ޠ�q�ar�����4�wa��J��W}bff�H��uSE����K�EZ7�Fpˊ��N:Ρ_����
�Цj�(M A��`i����G�<)����5����ّuU�4��Vg�]<C���.(HJf`��.M�� ����DǏ��I��*$��G�O;��Zm&s��k�ST���A"b�z�����T3O�5xZ=I�K���L����p�o�a�O.�K���l_VRy_u��{c���)m������.�x��F7~C�r�3Z�e�-�8�}3筌�=��Ϧ�u��V�+��A}/�ZV��t� ����}�H��j�����Wߋ� +@�͒��>�L7��s�uO59�����W=��*��N�V�q��G#���h�?�ؒNr� � S+�C����;ّ�,���`�筋�'�kE�R�m��S�N��63������*�٢��3W?l����-@�Ą�r:���7�T�@�;�,^ԣ��-9z��̪V+?�p�8�mj,�D(?�D���﫹y�}�	�I��@�?p9	����E��)�������{�@w��X5�:�L��y�?]mB6�����:�2-�?�ևJ(�S8;��{���v�)��C��8*�a[����}��؝琮s�9�1T�E{�z�IBpJ9��T&�N���Hվ+��Q��a4�b�l]�����YǄ�u�%���r��g>����.�U�