`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
jzHT+BvcTiKVHAlJPKFpJsrZFwpSChz95iSL9by6F/lMHDUDm3easqKGmahcILh7yeIj/QECslv7
4sW10r/nOs+1U1pCCpIk40BcjHnONxPeH5FdIX/y/DUqbiLoRmxnSyXnx8gt2oe05kVfJHFOfo97
EOv7W1FYDcerYSXk53qRlX2eKC5Dt7t9qAMdpHGL3Y6efg/wLNPS3jrC88mE1ajzlnmSM7U1/yAH
iFdEzNgbXUEsqFzNrmvrxgcLyD+anojfDQDE2LH0zaIdwvVf0+uSU6WuOZXysF28hbVAWsdeavHN
oxIy8ayHKz0TQ6SvRjEIUVkNTM0nkd6DyPfIUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="6CI7pN7zuEKK94Xv1e9JddDMCKRSOPWwlcOmaeXgy4c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
QxYu7/+r/Kgg4FTSrnwFR1xaMaFGpY/Q/wLaI8CEANxN+Vpq2WHi4XpO+IT4SRrWKhL5U9RSxMbR
clD5RxK/Dk8cPUgd5oAgplL91SRScRVU/Qq5QHsTXRoRdGlwimYQEcaEiSCZYk5Xo5X42Kpcw+98
DNz1jnoRDZm9U3WENuD0xAvhmeeKCYj6BDEoKAxratvoMuzaHS7SsF35vRgTMOsGbvOLQTTD+I8Y
kql/0YiSwYmZp8cytTcrSeCtiW/3MflJKVnYR4K2t0er4XKQ8WNGhOnmXIfOIsHXi4/wplj1Rlxr
NcxLeYF8H8JDyWjblTHUN3l6nq1+3QvRRqJMsQZ0w2ZVfTqxTu/8cwBL5CXPf0xz3LY2CWO+wNXX
ZpElxB1yQw52hJbgyL/LvoqD90jAPCA2KqYXgHoVIBhEms1dJ/5rcyIyvfuAaY/Ohn5K4XF3NQpG
RJMhoviCwAHBHkf1ooiVXgW0dMSM+nK3I194d7zqtl8lWHHXVeDy6oSGuBhx/mv1jfNywJ2rIb0a
qKuBeVdAVhSWBcDZCkV+3RIcuZi550ju0zqD8M1oEik1f07YxiyKNKzPpjvduNoKmW5gOjbvfa3N
D1exHqdplqw6OIKBrVbwZ15jzOC13zGZUFZdnJ8RE003DaeqBrhrz8D12dxfqzY1zuzrcN0BJbqU
1Tet8UIjquz80hC7K+pc8txC+WPJY85aZTDAhDM65buMPy0DbEKoyutKuVEW3+jcrhX4TGOeb8t7
2IKsT6vagUcdx+7SqtPMNFuFmJ4Ces1/Vs+MfyUnJsKuXExqH0AhiZPkilqhgqe4te/RueDXe9t/
k+slT1ybpQhVCIVt94E9uItUHWwVzxIkX3XUf6yqOgUoLxResYtAsVcF0yqxgFhGVrxS4RgqldBA
uwslc/KTBD7+Pt1yGEE8qH2qw+848rM+zB1JTnV7voWw79KOyUqkfqmJ2PqlwH66bXY25ohE983M
6d0/aD7aPasWSSTehB0IgrxkfuOPv0f5OmxzGfVrsLuy8uAGd+R+L3IswRDsswhuzIAy/VUPsTGl
4bAWw6Tl/fpnV/pG/D8UryzN36cqwwoacANw2mbMgAHEMsRVyd6kqptnlfNbR31cHZH6O0GXNBGu
S6dv5pGfEnCMBvnbFAgF7BVYXSALe+VDjGqlSbYkckeLhcTheT1RjHNa0NzYIBifFFe+E73Jh6a2
dsRj3UdOPJrkg/0eUuxksml/ttmvgQVx8HnxPKBVaDZMOp9gBrUmvZ9sH5jlFjbFVh0IT1YBOAdf
ChyRWEiv9A/fJuYXbggXZoGq6iphwNiEf3pRfi2mEMRkBczCftHLMgoj4Ra4ZupIWRQK3ydJGELY
uRNQiLPRjzZT4M0QJfzZ3NrtZUpDlAi6BrsEzIbKZ1tyjUVRZnyyUFiMObbLlnvZ26ZdKzR3L3Cj
HBHTPmI4HK+WUwZPI2mNCySLaQX4+7VnEbQj8V2Fnlr8Hfoqnd08GqwyuOai7BiTR7FI570gZNEq
Hk2JKumcnnwtk03oLAiT+ziYZ9lX81pOHJHaM0cFWjy0fXFfuSzOBOYbnVIS3jPZT7ULFqLTPsOJ
xVxnGPZE7vmuvPIfIjU7u33AVcsqOQu2u9P+RearaxUMZjMc6D2KlNxVkwmjZRYdqJewkz1e2+bF
iOfBi0N++U4zIs8M1i+ArEGzVHtk9Cb86zasB3u5Q8u1WkXPIoX9aDDnSUFLpdaXOgjsVzme/yHu
xczinTKJiJCks49HIc4ztznJDWAOUK16YFRBfExP0TrZYhKLfe8pDpYpQVVUglhIevExx/KAjz7t
xg0RjoUg0Ju4tAqZtS8Z3be5J3WkZ1bcrOV+/mqwOfDVORFM1hRvbP9AOfNB+JnK5mj2EQ4gdTs4
r908hLj+sejfg3RfMOLijXOeDbIogCylouoK+XpvA/5gHRX/XsHcbcRSBWc327hPIbt4anA/wh3G
IEtKbZNFVDWtIxIKwSgrDw/A3DZldLdREA3SzcRShwIUsjzae3Oh6qUYXsHl3mILXjdil/royWgg
2aFEbmEm86U/OcIbMmoiv72JCxBmuMHBsx6xspd89jDABFxOPni8pbgJ32KmCEqlulp6qLVzX0TR
XP4sHbi8aM5JM0nsr9yPm4RqAKDJ9HUXOScKYbFTU0c9afmFNtHgNVJ2oXKXHt2SppyKSIILKKAh
zQf1oF8nbeLdHcInXrz8btJE5TC1KL0LpXpfI3Q//1sDSKF4a8lVBaqy/8fW6E+NrcskEAe7ULdo
8DMGpBCY3aQfw9RRoc8isAWhLdP4Aa+cqhqH5WPMrCyZVCAks2mYbiOEsvg8YyRj+pPZWHByP8V5
4QNRrc4otPOieTsTBRLbr1/DMBDAV2/PZy0tCsABsxHIW2gi0/FE4i5+n2nezDjkAWuZRUtHKr8J
GQ8tQchs2IHPUCXCpRKjxq+V8kDSvk51bhVStq2eFXWW5qREn4xT3J39egvplVMPc8oss97Q9euA
4QJIq9je6PCfR1eXOFuHxbWE1IRQxipL6IDB5Un9VorEWFxhFmnZe8Q5G2U742ts6lhXjAUYXfcB
XTqVvK6xCdSWpGSKM2+h9WaDAHLmqfgRhgn5Ubv4AP6GLGavQ9UnzJ9PBUb9IACgaUV1ubBUw1zO
q9KL9h6nUxuAD3A1EaiCW/7zJhGCK6NtU5bUjtvXdRZDlhIRvaFqY3DbcDLIFjcI+hTxy0HeVNKJ
qj2sBn4nHfqjqSLBN2oAvW6W6vLnPRXpJxNwnTW+umFeMDQZRdxp72YuKjiG3ovunb7IV7iWhV3W
xEESZHrb2Hw4Kw4MMLX6bkg6T0EO+Hoio4g1OkMBy6suseTiTqbjuEIIBdDDUjrQZ5WDSJW5Q0Gf
YHVR5ug5h8EqYuijSB6pfIdRykJ7e/9yJZYOwA89LlzcLEzq8ifgYdMXMW3t/A2K6xnbTJvoQ6OZ
nYYmNFyVQV21SlUSgYgz60F6qkXrLVPiWZCtTPRLwO4OkU4MeCA7AU3ZECwle8FTzHLBvvGCcZOi
Z2HGxEeZD+I687B/sCz3KaEKVxNXMxYfVl+vf4LKt6yVacqmsakQilSTOkPIuk9sfP+Cd99hEqt9
JSd8xzHo5MtJAhTr5xRh+nWQ7eF5LLKdJSW2ce37OwLqvVTGpLANLnmx7d6BzhOIic5AFNI7/zOu
IIaVA9ptam/vH2wWFkFHwm7qgr+XhMRbRPTH3Zac0adL9z57TXvPGZeI+Ws05N3hlNsMTrlgGFEm
L+wlcY71OnGir5I64a15sf8CIM+QvexFGJHriDBqvhBOoLyLJ1jy5uEPxXgDTCWimrTNQAdVlEYz
3ykiFhq0Wl8hDOCgOY6JCLNgKI0c8f/unSXZViVhi/4/V9lTEupj+WbXpsk32SC2BQ4hg8hr8I54
yZ9pMUDtewAxjI+rSrh19+Hm/EHfq5yAddDNilqXy1Xsfxy+62f1/PeHVp4KfHtgPQLvv2yBkKdb
hAOTncpzYi9sU+JreLz2FRiEU/lNOxSL+BPF/YmHrXfTWFqqctdXsd1tCDhZWTBs2T3kZMBzyJCr
UtymzVl4WIQIu7Q5Mffrf28z8GskntSQWwycLMPTeVY3yDTQTfKFgK+BJb7FZ6tPKm5FrQjItGeF
gCEZFQSevgvZhaKtwT7JNtx8z346yXpzBJFD/spRukR8PpoPFRxVgcAkQr+k8AOV/879gYF6qQCp
789/GxkPKFsRpNwLQLzMlfc4bSn2yBiG3O1whBjv74Zljmr/jy3/PduYYq80t4R+lFDtn5Zy1uW6
D2G9wMpbM/nyOViSPxVEOeZnQ7W8xbGVzQ49dUIXFKk1G9ODw1ys84S17Pof7fnQpRAMVHemYxI/
z/NM1GA2/TGSPznQRXwIxl7ecPffr97g7Drmv+8KgRZuKP9hEe3VYTdyqVM2UHHPaBGRI72Xap83
1eJ6HM6aZhteliDu+/KXFPlTfnSFodFsswthvaI+qEcGGh0hST5sXfbT5q/yVCLvvp9VoCuK4Rvx
zYuoZcB3zKLH4S76nvoKLDGGnBdDwB9HvnPVLd+i4MA3M3lmBphpY7YJo0hQgJx0RG8ygadgQfG4
IAIbkmnytp2VlcXrWgKAjfNW49sp1BqTQlHVeiyivk9vFgyKrcdNAI/197LVDD/Q73yaz4uDPy8z
QqYskHYchCnAdbO7waL/7iuJezk+QdvjSGlVIK+ccOi0zD+19Z0pJtxhd9qLLljPWacxI9eRWdAI
QgwQ7+Gh3XWV97RR9nu+JeN+4rxMXV+xoibH48ri1fdShS1x+xfTDLEZdyEuwEwzcI3gtmusCaX+
vlqvCJdsGsQMHPh+iBSbpob/Cu7QupghIi8MbLcL0kDe2FusPSrbDxanwsuIo7JTDbU/9JxfteZE
tY00t60aTZLlzPKpNt9aYwrEU16Jm85+2JTNwJXxQGjM4wvdV6jb01EEq/b68f83GviKDxnpK5hp
xttH6giLgoyHhEARC1bDBooNsZ78ffeoWitCmrJdzFO5B2f1gAc6+p8L/NtWn6nbe6Q+YmmAeAw5
asngbvmWSENzi7X0zn+LngEh+gkRlZ71y3jfxGWYCW6L97PGYvA6cnhEOpk6h0jNxT6ohrEVDUu7
ZesjaWR83g1PpPN4oGE+YSID6w7dkrsFLLdDpPNU1SFIxhRY5+jbY829c7jPR/RX4bWlya0qjjnP
s0TQqDdAcIh79AyGepotGA/CBHy4klDefuipobNyShyc7ZSYjfAerZodr2niXvbVgMQa0LnXhZY4
njlhUuUxbyuSiPkK1t69MYwdxJZ8PJB/uWc8/apLrxeGofc81WqNuB+DuQGC9lQu/WpFHOwPJ570
HSLStu14Gmwh9voIjgulUOUxOQeLe8DrKrh7c7b6nr7bck21ZunYv1IP+5zNfgUG+ZXEe9l+kB1s
aBbPCgLQdBEJNxcEqh0jIwX0mXch1JrVqPZG7A1u/a6BAhucHDEFOIOibqQz32vlIavzafnNAb3q
YxnqRv/APU12enqThiHrL+5XXmTUFLPspPkYYE6jM8eHwjk28qAPakYLXMFahS4qu26lPiKzJZo4
Na3e+45JAl8Go3dn3E5bBrvQgsXC
`protect end_protected
