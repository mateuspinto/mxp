XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�R��9�
�%mzi���v��aO,�wl�bV45�`��*p�Kil�6/�L�����������a_W.G�6�@�,��<�J�^�q)�W��v�4��]) �!��B�������n��0�3�7�$���k���݃��yH���g�=�d1c����̃��L�ղ]�e�e�t�����k�Rp���̷����kR�Jo�������&5��ʡ�hGg�9���ݓ/Q:f�H{G�{�jERC��cA�|�g�c��%�b.�a:��.�X�/�
�aϙ�}ЗMp)9� ��*�P�aU�àRT��n[���r�ޓ6Q���VUl�r���{jzƠ*�d�ؑ3���T��g�������f�Y%�D� ���q[2�Hk{p�"���,���O�E��#>]���M e��$c�����yVg���tخ�)PP�Uz	e��)�j��3��k��S���b�Q��K�ō�����0*F�_yd)l�V�b�e��H&�%O&����(s�GЇ�3��Wn OB�J>�s"s���c?zF~3B�O����k�I��CZ{�E3�E*�2[*��n�Q�y��:I�}җJ�kTa f�=�'��׮,h�F�m5 �����a󲉜�^!�d�yW!��"X��������E���}�
R*.������uA�.C\k)	� �^��.'ab�`���'��/q8�]!s8e.����٥�,�u������M*��O�xv���zBR�g��iF5��tցw�e�_�yJXlxVHYEB     400     1d0����x&����w��`E?�>�Tzsmz)_RL������KF�*���5�!%�ش�H���1)0�g��	�E�ZbcY���]m�p舧��"�C6_�"�ژ��} (�i9lN��KFI���4�v��H��H;B ��b�X֦�6۠;�U��+�WW8	��j�b�}��5GFDV.gn=��-�]��3v}K��lʈ�H*�l)�q��6R���@5��0�|�>*{?���cf#P���/`৙D�p��;/��H��-==��nyل��a��'ڞ ejJ<廐���������ʭ�S�l\ ʭ�oFs���I��u�齡��wT�q..t��y��u}�?V�܄���s2���jE 7�
��w!�4.^HU&�W���&�E���i��蛕������;W���_�,tj��j�IF��G4�ڡ�!I% �i���Fs^��"v�hǼXlxVHYEB     400     170��o$���"��x�<5Ǐ���)X�-[2�)r�Bx���w�r���D#ۻ��ݽ�3%�˯��K��hf)��Y���Cc��cn�q���u��\��U%���
G�����)e�v�!�űA�z	��~����,0'�vv��8��P���tҝ��NΟ�?J�.Tı�:3Ny|�/rWK��~��"��~��T�MM]g)�F��H.�]��ӄ�$�L	�?!^~4��(t��G:���*�֓��Z��1���5m���ȘnY��~�-0m�"���:��omf�Z]4�Ơ'}5�@�UD�qǮm�JzJo� 5�j!����O���M0�����̪s��>�%���Q%=e�H��<XlxVHYEB     400     120罘�tŹ�<��rM��$2�H�D�B0g��0EoN}������nW�dwlv�p?��bAT��eZJ�)���W?�j�{9�/=��晱xSxhB�4ж�:�Ju�|#���6>�H!�5�*O���=w�T�s]�D��i�E�C�e�]<�C�uj�a�Nl�Ng�z6"4�I߫�ù�2�~�=�-�O���tHX��pOQ��F�/�W�t@=�>j��0uD�I(��:�GKHB9����fo$�����9c[aFs4GG�{F����c��OO?���!F��XlxVHYEB     400     170�MG�&���bDe�.��_Y��:�������>�U�9.�o������_�,�.&<��$���s�b]�7D1��3,S65:��'
�9���~����
����N�pz�x���!H�3LZb�G�{�D ,�����g�6q�5� f�[��]ZT�Z�d����2����?n����A*��2���J��A��><P/�d"��3e{�n��hUq~����`�Xu���D*:�E�3`s1����	+ӣ32]�; �i��Z��Vj4w'�-�5�Ӛ��7����)
���;z��z�~_��Ua�T
 ���5��p%j�9OY,i��N!Bro��:�P�T�G=��,���Bˀ���zԤ)��
XlxVHYEB     400     170HVJ+3�l'��1PЗ���ׯ#�GvM�lJF`d���c�h��?������u���H̒�T��_���ߐ�FM�*�ԯ9�_H��!scNv�L�c���lh�4��逸
�M�-�e�wF���vG(Zk��F���J��ۃ�K��HF��>���D�CG&ҝI�D��P6�K��h��ڨv�;�0���o�Kсu��$���>��9,��-�9���1�Q� �Ο�_?��C��}��N^,ޭ#Z��TU�~?��[�j7 �oR���s�M�X�'���%K�Q��P��#����)j�������cĶ�ă���}Yo̅��Oqv��#������(��q|3��H��$x{��b�XlxVHYEB     400     140=\JRu��\4�9�����WTdx��y����m���U�L< �9�� r�9�5O��9�������B;���}�H��بB�t��GB�s�с�\�:r>I�?+c;=��#lC����$�
~� �Ji'
f��(�)`�%�s����03��S.�,�=,֭�Ҭi���+8�ηq	��pz1�B�#׋�黩��>Q\r��{?ѡ���nB�����n��`��A�D)QB3�Ēa�g����@�ǔ�i��Q�7I>S�>0�_C�σ�a"�n]M0��u�ssZ�����x��/����ȉ|��Լ�f
��m�١�XlxVHYEB     400     100��]��h��jNR��S��G�a���?�Y�~fi�Ci�|��M:��|��Ĉ�F�qP���i�b�����G�b�g�e]����r�gy���q؉��b�xÃ�<�J�ۅ��2P6��x#^e<����ީ�ǹ�Dѣ��PS�gB\VB��To�^�9�3}-Ѣ#���[�O���Ox��S+v=�C�PڂB$)Ez=N�^4��B+[�F����g����CKe��Ws�uu��?�i7^Vf�ⴃ.H�x��)>XlxVHYEB     400     170$�j᪈�������	�)�$:����"�ܩ�� �G�@"Z��m����o+�;V�k�3�c-�F\&�O����p$6{��lkd��|Ԁgm�X� lJ�p��+�o���UL��?T�����O��+8+�����c�����l�6\sQ$6�>˪�[
+�I�O���~����9�g�'�@w���G���"��؍_�3�;�-u��i��1�'l8�P/u�$��z����& ��A��X6j95�f�jhS��*�%;�_/�3�-v�+ӎ�M�zp�H����r���V�ś�e���V/Zy�"��j�<Yv4I�k��Ǫ��R�cV�}�%�ҷ�v`�#��(��p�AȄB�.ӕ��XlxVHYEB     400     1b0oE�8M�]+Z�TG�1*~�yӔ�~�'�X����;y�(}9fm��{�!ouY�r6^Y�˭�L�+�oƝK]q=�������A�8Z���Y��|��
���d~��2w��]��V�oԯ6��S&����x.T�����0U`+�<���Y�A������F|�l4�����IaH@�H���:#�RB$D�b���qr ���Ѿ�I�Vv�$��ޅr`=�)�֢�Pu��'�&4�ʧ���Hiu�BDɟV��X7��i�Ӿ��Ov[޳�Cj���|{�tu:H(���6R*�m8�qI��Y���1M�14����gO�B���S����c�L8�Yu�ju�*y��7/ԥ�Hb44�T �jh�5E_)ե��/�>UN�g�8�'�^�4rN����p��m[��D��?;���/irXlxVHYEB     400     160��<LV���l���{�܃��F�(�?�m��˳�C�
<P���NCp��P%��\1{�~G=�e=�,�KwѪ>~bx� jI�4�� �<슊�?Ff~r��Jn����"�#
�|�_����,��|�����ͯD��ԍˬ�uQ���-]�K9��I���f�)Hm�6���Fxzߌ�ԝ,�#��}}�A�?}�ZWھ%f��164L9�������߈!���T@F���v��Pk;�$�b��!��w�d���̴2�Y�
�Z$>O~~���6���������|5P��	�����n�]�s^ܸ��������5��8R��]��"���Χ��8�{����+�x��-�XlxVHYEB     400     1d0~T�6p�n��R�o�<�!�����Ō���Ev���G�X�B�������� }i��Ps8j�j�Ɇ��	(ӧa��Z����mW�+%��(��?��@�`��s�0b���h�G����GV����w�Mq*�5g��R�d�.)Y��G��	E���A���4�/�BѸ�c��&�*U0��tf�%׵��'c�T&
O�w>���'�����8���E���e@Lo�F���F�#�����Z������>yLC����L�Kq�F�i��S{�KI��fE3@������m��9�Tzd�u@�cx0��vĚեmF�d��%A(�_!ީ�J������D��o����_����f��*N3�ˈ6��`�g��`d
L�2ƍ ��`��̾��J�K����B�X7k"��V�Ħ�'*���<�GK"�����.��IGNH�v���XlxVHYEB     400     170�»-��7/�g�O��)�(��oK9�����_@��0_VN�^�GΫ��=Q��N%Ԕ�$.(ƠDks�0A+l#z��y�g 5V�U`0�YLH��j'b�Es�xyE��
���ߑ�����o��Fꅭ��d%��T�o�u*�a,�T�mw,������ǟo��]ŭ�Fk��*8�QXpq,����J��["�ݦ�u�mr�fuM�T�� ,�&���4�:��*��;�f��I:�ga)c�܋TEvKB��v&җ%X/���Y��v�֍jo1����D}1&B��j��8�������ٕ�	ؗ@\qho��ǏvO�&Lq�n�T���̯.I��+N)V��W_�6��d3fh XlxVHYEB     400     160m��G��Z�t);���j�IDdj�723�D��$ �a�/U�p�Dl
�M�9! A�!��h5���>W��;��{f��;^��J��Z�%_�i�w^��ɪ�������&���v;��i/_�����w���z��@h�}K��+���Z��R�ZՎ�I��A� �!���An!��:�f��Ы��]�C�[���,FG�f4����=�f����_QqM�`d�,I����g�JNHGr�,�c(De����޸0������A�=iQ�~%@�V��z=�sv1��K��nJ��$���r�&�\cbH�3��t`�)�Rd3��q�,��U)��9�_��k�m����P_XlxVHYEB     400     180&%0�!�,�D��0��l�<5ȝ a]P��p�+¢����;���2���b�^�-��jTʾ(��-�Y�C%i��!J�����J�0�Lѧ�v�U1/�^�3ש�6A4�O�E/�b��Uε~��bFP'�� �b�}խ�����J�U�<��d9�yR�ǻ&+t��j[X�хb=J��M���]߾����ߍ��	�V;N&>�w^���%k8�%uk���}��?}~	��]i��H~�fJ5��_t�n<����������ͭc��嚀�ֲV@_�4~t��r���,{e��c�0�R���\_O��y3��'[����*�����M<p����q�A�d�-�=������\�r#�k�F�x�0�XH��Ӈ�o�7���XlxVHYEB     400     130ެ�]J���܇a{m��i�xj�;�S�btW5:�>bb&�!���@��B�+J��������e�"��36xH�'��r$�9�C�E�R���}B���C���yXp�U9+]/�y��AsL�r��IN�(���
�n�Ro�4*�b	�쩸��DR��G
yת~b$�rM��@_^��-I����-3��fTF��B4.��G�S�3�VOw!�6��_�^��kR�`������l��ק�7Ŋm���\�丵����d�yJ�e�uvm�阢�Պ���BA�N|����#���G=�XlxVHYEB     400     160�j����q��ͧ�UN���TÕY���yC���7��5fG����Y�q��*,0�#�H<�zu����-F\��Ҫ������L�ix46
�	7�[�����CV��*>i7[zI�����7�]Yy��X�}�n�r��s�>���E��y��\���I�R�0\������ ��z�C(�j�K��v��JY��#s\;0<%N����uȨ�j�>@�F���(��@�_cA�9[�� ��K?�@��cy��S�Y�s��6�d;|�xf���O���k3�Xޖ�B�9��)Ýw3(��-��7|<
F�+�����g�^ f0u���k'��r!F�]����=�|S��*�-]�XlxVHYEB     287     130�AJ}Ld�j��,�d9�p���l��+^���W��w�ZFQ�J��aN�47�8i ��6��������O�A�GD.���ԋ�jU�G�+�_x"aϓt��R#|*_��F�N����ʾ-��V���۲��NƱ���փ�r;FP&y���avɦ4W�Yl�Y�ΖOC�Q'F7k��(*=�a������]����"+j#(�f�D��[��	�2��zf�,�D�G�AT1�`�a�)�ڊ��r��������O%;��ץ���b�Z�C�*�\K��Lf�,�
����)�^�