`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
LmnYEHHWvRT7HgYUNNBw8JEYUJ3OhpYXVikkC5rzj3WPNJCSn0a6BWJvbYOlEWCbLNPfWkMcReRk
COmXeAjRdyZHrBJk3HRq4lmZ2fXKELjhtKmgBLXklsn47UUTCgGMV3wMjWzojqbEALfRZCsuouQA
lhF/vyk3/LKzUQbweRL8shHUGVYD6mosOGsiTexOKSwPL+5vMuXATG0EnNF+A8zNp4d6zWJ8S22/
0tVB0uMvRHYk1v5h4DuSt3xMs+xD36FpMMwHmsAIrqiRuwI6EuL3wnex3EhOkdWJ7oo7rXMCHfBW
CHD2FqLR34iu/uKCFyFNhv3l8P2uW0xThmOPRg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="IIgooRMswM8ATFOIUIKtEocz7SUPa9NMsDW0RUFQbUI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
G7SRqa0nhV8L9PcXtLu8/hcQCiULNG4ljtl+aLD+z8JcsCdA2olkqBRhkDrxL091CmkiHIGgbYOY
oDvOS3Z3rPE4qGgX+vGHkVc8KA2p9Ac1S86q+MKq5DGK3b5DUKmR6mrL6Tlxqa4veAdrzzHJJaxv
R3LWkD9kXaH3C60MZhH3i6bP8GZqFIwEwpP4fOu/2eIPQGfNNXTwvNwpejjain5VSsrNJOewbk43
gEx9P9X9YKM+6UllVGLYQxioCfZI3/F2pAa6sM8i4oXV0I+rd7gpy7KkoiAIq61lSDNctV/Wrp/c
6yVnUk00q9aSt0Z2VG+v7F8X6rSREaFMem7nldS1Eg3iuzsJnVmILqjjbS/XJ9VRm/+TNls+JGt/
YxggKm4xcNl7LxH/cG+PXnqMxXQp7Tb+3jbGV3nWmQbTWGQTOCGktnL9olcZB3bsTw7vJD3OTvFi
+DZuKeCcUoquYKJzZU/E7c/QMtilvFamxUutrMOGomwAwQtMG7m2LYS1fkPnBbRCQtWfI7MJcD1j
XEcTqDrXyaUnQXhRazKq/4QCteppAeBenhVOoHKcCZYEKVRI6bbzCWWmQTiidgPi2qSW+q31LhpB
H2tUfUl0ss1LpLJNgC4WNL7rWbwrwBDzPRNTOdRP6GYbTONkml/BS9N7icmtGyDLseoUL7VkFdA9
JVwrhRe0rZWEowXyFz3Icrm1sEYvzBiRTOoAx5ck76bbrcG5OtDXgkgnYOsz94N4x+QshPwoBLWm
lKa3ou1+2SHgtukv0PzbKVDOaMupXqHBhw0SHUqatII805rf0d7RSPKejbyY7oa2D5a1jGgJLhjF
Fv891r1JF/LANuAY4OXqWMQbgJ8JqBESgpx5mz3/08zIq649xUmM7/JYJrA+Gp7Y+9edwpRVh9L/
0d2sZQ3SUiZqTRw2+22CP8fjm4s+RgaPsFM/NvvjSflX9RfzBF8xP6e86ew+rqLU188+hb3M7eMq
cRciPobnZ0HXzKuAriAIq/0ac+qsRQLtYZ1tX0QGG5r+sHmMqa9OZ2MIwFVCgT6Cqs2WW+oEZX8J
maQLgOLR616R+1/3aIjkroRwkoFh67YR+QlWw0Hi1Xkl+g1iaTVGOlZefWh0d9S6lyF+KCQvDmsU
5O/ijBGYoZmKJK1VWVstjyWyF8yZ1ItvcO3rSNmNDFJXj3oqgYGKwa5QTp5Av/Ecic4NeWIC7SAn
JdLdABbOYurHOSVi19FKSg==
`protect end_protected
