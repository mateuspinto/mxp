XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@"�4�w��2���-�o���79y�d���y��hS�Jd�����~^�m�������}�򞈂�wS/�K�k�Ff+�u�m<����'�e6
ڨr���_^)2 �D���>�$��5�2��|.󜾠x�K�5(c�1P �㢓�\��p�b�Z$��DpʷݙI��:��hz"	�(���KuO^��j���U����Z-X�$��dpc֭M��:�?k)5_��PZŕ�pBȌN�q�L�Q��]�k�{Z��2�5�\�] �x��ɭ?e�0[~Ӵ�G'�6���f��;m1�����<rW���]�`������J�y���,��u�[J�$�����2V?���eH/p7q�Q��,��h7R4/�?��]ɏW����HpPؑ�J|F\�B�!2�֗�N~�x/���������~�j1��(��Ja����׉����/��A�X��u���-��M~V	"�	m4+4�F��$�|�!Vo�T��Q����V��;<�i�!�Ω̃y30Yq�j����x,�G���)"�[�;����m�g]��_j��a{�%���
M=#����H����iHsE0�,�c�T�QzJ��G�������@ga��s�qfϠ����D���R؏b�@�r-�y��~ t�|��OJ�h�R��p��vs1���D��H`��-����5�rFBi\G��&��M�<��f!��5��NF�ڀH[h�wM����vAJ<�i�Z��S{�XlxVHYEB     400     190�:K��p�z�yΉò�-�2JU{��[��3k�澯�* �8́!<�Qζq��xq�<���o	t��m��T��O��}e�\m�?���J�4�	I�ѣ���W�aP?�S}������/ƕ

�Cb~�ui٨g8�CN�o�4�������l�aH���%x��&�A�M8�+��N~�}܌��"0��*K-��H�$V�!�x,~Ι\u.��q�<e��Jݒ�1��O�L��c�?ՆW�1V/����8XQ���[�(ĆH@߉3�\�-�3��|g�x�Ji�TWv+�x�S �B|Mx�H0����/O��zμK�Y�)������O��/i��l5k��z��A�Z�Ɇ< v�=M��'Pi����{��H{0�x ����p�����ӎ�XlxVHYEB     400     140�{��oG8�'�p]^II{��?�]&��ϊQؔ���4r�]�|�T����L���A�s@]�=�?x��{����痩���f֡�Ήj�c��g1,��L���e���P�ր ��Ӵ����i�ñl;pEM���JC�'J�B.ie��X�#׋� ��o˷�����o^�d+�(���[���!���t�C�~L�V� ���ͽӮ����(F����Ti����C-��7)ph�I-����8�����!�?{Q�钌�Y����R�x������>��!�ǮB�jP�dݩb��͞�zE�}]-�/8�Y<xg��"3�&�BXlxVHYEB     400     130���=�.����^��P#�*�َ��p�I���_�<�3L۳~�!~U򖱮�֍/����*9�N�t�~.K���k.2--�Ӥ�3̨_kɵԲ�[2���;l�q5&���>�`�Õ�\]a����q�b�L/��f�B�_��9�#B��bM��	�[�x�v�n��3i�t��ۭ���Í�X}���-�C�J��d���(��xۭ�Ѷ0�sĠm��FI�tda�5�TVB�/O`SM�6�(���#�^���'Ӕ&�C�t���~���:[9�˾�����*1I6MBKߞ�m��=H�XlxVHYEB     232     110侱@�\߽:�0R�����1S����(��l�p�����Ǵ�
����9y�Y7�xc1��i��}W��{MȎ�ܳ��Sd[��y�F�q�k�	 ��	�&?򡭞 x(&�~���n�*���
"v�.,������_-l���p��@���AՃU�N��Ҡ ��@W��-�ꨩ3�1��.�
�z�wM.���A�P���-�6����<m8�bf�n��h�/1�F?��-�(��X�z�ţ��La�(���2\Y0�P%&r�[���/�