XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$F+�>�)@�R���f;/��X��$	^�⺦�
�y]밇�=�����~�����Rc^��?�8s�ȴ(�����p(��`�n������Q(���#��O��`(�4Ö�@�򡪉��Ics2��~���85U���]��t��z�n��ED����v|�M��]=!����IȆ��Ȅs�*�#$<
P����O�Me�[�x�(E�]�����P6C躨k1r���H�}JL��?:Kt�b��C3��T���u�F��H�Z�ڡFd�'�gh\��J��^�z��l��E��:�"�C�MP��\��_^TL�"pXsG�PJ�O�@�F��6�����Jѿ,���mH��������~��f|�������@5��UY��΁Q�3�sO>�[�n��:%'ᚰP���n��'�U�T�R��u� p�ě$Ń���e~"�b�!��[C����i�9~Gs�`����4�,1�3U�P��f�fpF��9K�O�F~K�r<5��V�9���`��N��rR1>�rU�F��2#�EU��Ad�ȩ�"���iٻ�͕:,�57��%:����JhZ���<�����B�˃����U3�������`$BȅLb1ׅ��8rTg���b$
f��դ�B(y����[��������� ��V������C��c�KL��2�ҕ��5���	����ף
^�{���%������W8��$U�l�` ��hU�>mF�
�V��XlxVHYEB     400     220J��G`��õ�2�`�9���ҡ���u�w//����O����a��M� U �Ғf�s*� Ok�����X@8�D�o�F�ë���8n L�#ɞ�N��:Z�Gx�J�f�@��Dgt4�{��J���{
m~A�I�̂�u��z��L�y�"��;��L��/}�h�5�v�����zuO�=K��9�K��p[�ɥ/�/�!�����i�������lq%̩K|��!��>vG�\ԭ��0���-�]D��du�p��`�4�]nG���q�uq��0E�0F#�/�=�M� Ӛ�$�Vu5������,�9%+oQ��y�:�(}#6�&0/
QJw8��a|ԾsN��4C�H9gd0�S߄]���ke�v�{Z�ǅ��aa�T��m������L����
t�G�F��H�z�t�v��S�rC9Õ)"7.@X@j@`��+P�*f	,�#�4���1s�\m�T��E�"�����b�BrIԀ��8����<��*GЫ���bH͘����R�2g'׊�!|�J1	 XlxVHYEB     400     220(a-F���W�K��iټ�x�)r�~�w8A��S >��xQS`ı\�/�h��E{�����ߎ�yFu��&�2��^"��Or�K1��r��p�6�7k���t	wڢ�Ί�2�
Sڽ�	����S�ows{��<\��1-�pqa��c�z4�� �����?���v6��������c��E�-ChҼ�{�Ѣ���3N�����
`>���i���J���$_�M�k.�Ϥ
8E[���/U}bl���O:�:�x&���/�C�N͋�2-�7'oY�S�l:���U��� �
��]R&�rX�t��u�b&L��ْ=�JEJ ����H��� |d��[��_\�c�?�6헨���o��ax�G� &�!	�p@��t����X�3������O�z�M��؝�1��&4I�O%jO��w��R���d�|��[���(��j����N���ˡë9������"L�-�Ć�4H#�� �� ���ᤫ���q��2�z?58���0��vGg��jvb+'�WBU̫��M�7��JݱEXlxVHYEB     400     1a0}!b��Uu}̨��S����F��lsR�ơ
�S�K���hO�.��ص��(���u{���sT �u���	M�o�/
���_>�h}ާ;��rT!߳�1�dS�n8�������j�������rep�#�bGݙ��FЦy�ٽ�-���J��e�C�1���S�2hٖBJ�K�7"2l
�e(�:��څF|��vx(�UJ��6?�����]!����@Nr\~�A�U}�:g��G�@p�:��ҹa���]���^��	���u#U�6�6e6��$E+�qv�(�}�C1z5�]GQ��/a�J�N���O�u�������D�����������6{��q�[���Y�`�kb����@i���Q�M����}���*�TƸr���<�2&G
�ʰ��>� ��XlxVHYEB     400     130������=D�2�̡��!`�c���8�%ĩz ��Ĥ�O2�|�B#�r�o���>6i��S_R�k�~/��nW @����
4ߌ��L���`��Q�Ϳ���Z�f�9�Q��P����G��G�g�?�"e[+���&�eӼ��xx�s�Έ���l^��k���m�@�~��dɫ�j�;��:���z�<
غ�m/AQ5��Τ��;���� T��e�t�pU�+lן,��T|v�<�b�����l]A	����}�u�Q|*�C]xD�ԲA(�ś�k�����ng���P)]�	��XlxVHYEB     400     140�zMO�[b
����[	*�C�D�����	+՚.���� ����2�@���r��;�:����)F��P���Hiip#����.�;�ȑ�o����\?��>�h>.������>HɁ��?��t����s�tlC|�V�.�ٞC�'���]���k�m�*'�,Y˳L�3�J?��)���P0��:�s��ո�Y�ͣv�� 1)P�mgً���<?����Bs�(ع��:��-���(\��	��;�3<��:�����ODɞG�播(c� ��[I��� ��+�٠j�=C{;\��d
�/۾�q�%߃vʡ�XlxVHYEB     400     1c0�����|Ǣt�>b�Wq�7u8	X*�.�s�Vfe�W�Zya�>�ᰎ3��"��V�@U&����*�jV9ˁ�Uy�ň��ٲf:��ޙb�[>�U�j*	$���0��p�'�Vu�q'�VU�©��]^]����s�
  ����5��K�V��[�%����Z�oF��!A�ڰ�U�/20b��I���L{4��`��`B��[%����u%V'"��H�?��@?��N$�BMCm�j��I��M������r��Ty��6Y�)�Γ�Z�.[p�t.+aPӰ�8�2e?�/��i�4̆��E]��5n�@������9(���#c׶#��S�(��	UȤD��Q&��C�|+b�*��9*��-�f S�f�f�8m��f�QR��U���|�M-(��h��S=�c[�T���7��<i��� �K�XlxVHYEB     400     200�	�(�`��� �.�[���׺ҁq�/A�-G�&�7?��h��uY�ڭ@Y���0��c�� 5����던0�l .1�13��'2���j��ͽ�i#Ӵ7'z��^+���t�~c��(���t@ �K�$�#�F?����3�X Ok*�1{�g��`�����X�SF ��0}(X��9;�)��ׂ� �U��$+>�O��/�(/������>�Yw��goq�	��|�Wb�ԉ���K��S����aWz�LR�{�ֹ+��^���!<�k(�5B���@�r�}1�Dm��T\�Ǎz�������3�$WA=������ ���tJ�T.�iq���v$�}}�1I�Gw�F=�,	��uj�H2�8>�TJ4�#2[m�s�$��_oT���Ǉ�vL��V�G8/�X8?���M�jCTK����E��T걣8y"���6su�����s@
�7������ph��~��8Td�Z�7"���%�a�r�骠��)-Qڽb"�&XlxVHYEB     400     1f0[x,���U�WdC<X�]LL�;���8�����t�^4x�W��I��<c�{��)[�Bs��� kd'=xM�QIzցn��201(�R̓*�B>�_����5�B vZ����Y.� ��v�`x4���eR������:-�*����TB� /߶�,�QD���:���Q�<@�A�z~7ڥ**���Z탷�c0䏞�N��;F��]��xCB)��%��y���f0����1��n6��G�A��gI�������}Yw�a_-��M�����Bi[��E��~�nk�<�_g���eRHmQn�-���UDkM=�I����q�[Qek��$��R��~��e �t��(�ճl�t��ӁN�޽��&�fz�!׎֦��`�5o`�b���s��!�-���',��@ކu6sd��I�6���V�y�|�����%�[�W��]�t+�!�4�4�����'u�΃�sAY����́�S����W��l�=���`�i wt�_XlxVHYEB     400     1e0�2R嘫4�?1��d��O,"{-r`���9)���f���L���8Lv+�
�	�,�]@�zG�����W��RHxi�7�2ٙ���;�����l�33��s�zT��"�M�����{!���!�*�m-0+�ޕ,&IV?՟܊��"/w3�jC[��a��Y�R�'i�/%E�)�?x��SP�]��������$S�K���{MJ��Ÿ� ��F��l6��5��-�kW�iU%�;F��Ɲ����x(c�H��(�A�%�a�d?�� 9bC�+8��r�˘�ݍ�Qm��jFk���6��6Gv��á�X[��ŧ�<��E8�[����}��"����ĥ������(2��H^`RZ<��@yĶdYlw���Ls��jj#�
O=Z�4����=�T��Q�i�K_�s-%���.J�>z8@��őń��߻����T������%�(g�X�=�K��/ym�׳QXlxVHYEB     400     1c0	��IK0�C�]��]��Լ��m� b�̠S��b*��PGp�)V���vI}bk2P_�o�QP^tn��VT.��9O�/Sc�f�\����~m��d_o9MA�+0d?V��Y��?��#TC���b�å:���֢�˱�Dpidh-��gXbs�a� pa)��,����#9E��φ��ǩ�ʍ�k|��x*CrV�f�`4�]��{N{I8�M����hC�~?�Al<��l�2q`�)=h~�`�z�����"y��8�˳�~��u��/�K��kt�I�MT�,d��:q9�e*��v��P���I`�:2��qU�D���w|��@8�!���EywD��z��_m�-���t��oީ�*u�}�i��o$bq���q�c+������J{��By�k����r����C�-�9� �cA ���6���v� �RXlxVHYEB     400     130��|g��O~��Uf�a�hG�kx�N�o����u����x�FO�:}��s+w�tb��"�����:��|���fs�/������v�ӑ��O��
��A�	�tww�xު�7��˔�^��E�OH�_$|��Z��J���	$�߬��0�aE9Z%����,��O�=�#i@rh�^9gJ�����Q���0$&�[��$��I�795d�1:�W�h���*��+Y(�/��y�n�Jj?謑 YԪ�a�_O�Q��|.ĵ���`��l�r��#��D8ZDx���Θr�RZ��XlxVHYEB     400     170�WU��[��9��g'���M���f���YqS�th^%��Z���1��/��<JН�Ց�ߛh���T� ���@��$tm�)g��"�2�hwM `Hg͔ �_�'$.��Bw r���طϲT�i/��<�v����}n�PcJ\u�U$wU�#l��f���9v�ЀX5�y/Ə�`�H/� y��n({�4t����a̺�f���~ONn��%Ѿ��S=�<8�Y�>�L��a�*�C��%n?�%��`s�Ʈ`Ҷ���Wl�Ev�j�j�b��?73��H���8?�� 	�"i��.:G�׊)Lg����0�G��66-���*��]��M%��2�̳�F�WIk��WY挮�%��XlxVHYEB     400     110a�ܹ �J����!��q�&�xŸ �u&�GN�ۍ�����rV�.�2�BoW���Ae��;�� ؙ7��/�@2�gv�3�����a{�/;�SػsX0�+-&�MI�7�U�� ��ˎB�U�Zx�z��Q/�nʢ�!��P�̀vZ�քv
��&�;�h���ܼ� *�j��7���+X�������8�;UH��.���̷���Rm�0����ߛ�����I���o�s��Ge0�ׇ'�SV������-��w�F�5q[|���XlxVHYEB     400     1407L���ĄU�z1����p����k��"y�,��$�Q�×�C;E��tҸ^�G�w,<,�lV�2O��z�<��z%!۝V?>��ݝw����~�G�WŇ�
J�,pĦ�r�e{����h�[]9��:��r��<
��Cs��Ӏp�ʈ^,2�UOe�Z�X��g��zylr�+��h��Yn�X�\���	��F)1���ad�Q�O-��8�XȊ�����dB'��	����Q��M�W`��ؕ�nC���G�������D��s�c&�]��6�*ڐ���~� �a���D�(��&�����XlxVHYEB     400     130���P�ޏ�s�� ~%�G?�#w��R�V���x���x����l����O�ƴ��si��Y�'8�h���m�zG�h����j�Q�{8�����q��!��@��1��@�����[��JQ�(TR�ӮA*Q��T��f ̀��(r�rJ�܏d�9Nܑ}�R��O�L��{�IF��{"�\bL��?a�:��u��/*2+A�D���J��-^d�1�����~�hu|���X1�s����z�,V^�08���%
�.��ߩ?����f���D)/��B�
���(j�:x��^�XlxVHYEB     400     130���do镏��0�s���%�,0K�m�+L��Ec���ɘ�8f�F��JEe�oa�4��U�p"�_�o�y^H5�މ�g��$����P��q�[pS�vz zPr0��Z´�� �m���5�/��ͼ���3��9r�D�՟e����=s�9=@���R�&1. jY=��{���`Km��� ��
xF�N��V�ٵ�c�pL ��X��H��=d�ۂ;4ړe���>���k�[g�I8~M�d��x)�HsJ�E�f�8��*r��tYͥ����׊r/�	w��#�>��l����QaT`�XlxVHYEB     400     150H���d�5��9s������t�L��ږ�!��؛w-����mC���o��r�w�֯����@lŇ�ߓ���R�vm\��H��$�+�S�f�h�7�Db����-1"�ª{��+Y��,V���d
��u�}��������h��&QDa隭���gCeïm������z�x���9S[ኀ�Q�Z���e�Y������ 1�d1E<��1�����G��BqW�Ϛ�k�e��G4`�ؒ	��l�����VE��^W �Ƥ%(GO?"����ĩ�UkN+�D��iQo5q���$�F��ns��0H�w!�h:�ɽC;;9�9�XlxVHYEB     400     180�^�����59D� �b�i�5��?��M�Lz��H��&�G�������K2t;�U".?!t8�b��@��=��̓�@�����C#Uܼ#�:�);%�E�M�h[$k9\��l³Ɍ���O���:�"�̄c@	�2|5���'�����Ra�U���Lq�SgekK����Y���1�VFq� �կ
�s��J�"���S�Q�P��{�x���Q:����Sp��F��_�j͙Q���.���Z���s&��B=M|�Z+��N���׏��9�f�c�<��������7 ������7�E9)�tЗͳ�ˣ�����ho�Y�Qϭ�Zp9癃{�����se�Y$K�&6 G���=�����I��сs��0�V)�XlxVHYEB     400     1d0+8�>�֓ů��P��3#~J��Â���}�a��[�8,C�����5���MF�u��Ȅ�������2fNԀ�,��~�fa6��D�[1�I����G�~��W����]I1	�{�Vy�c����Q�X���e.��;��^��G�E�$S�d���A��џ�8�H.�-���&��ve�&ۡc9r�lɉi�.z���W�����9g������+%/5��U���w�`��T|���g���
k�'�v������b!?a��8^/\>9IE�aCq���ۇ�1�G��!�-�,�M2��}]��=ST�+���0hH����$��Oe,��vƜ�!0t���R�/W>��j����v���-���3���������8�M��@��M�a�<a�r���d(���3��S��jT8镭�˱?hd�/7t��cȳ��hX?H~~6�2�.�$��Ɩ��PUXlxVHYEB     400     180�p�j��P��U3ͦ��Ɣ��d��#��Rw#�fw"��)�o�_���~�cn�c����˃@���wC\㩛9���hN =A����`.��]a���@��G[���YO�sD�o$�N����/��j� ��{ɩY)��t���N��ux�p�Uv��+$|6|g�K�1�S,�~?5{�X��و�4�+)��9��j�UH�2�C������.���M���ˡ���y���=���6�&`E�=��9��A�������{��>h��=�`'���BO��.{M2�Y��ѽ��1X$w��zv,�E�o�� 'ݞY�:�+l���3��a�k�wyS"�B�L������/}����:��-��� V�0�u�O����ic��᷿XlxVHYEB     400     150m��+���L���9��]w�m�[Ў�u�w��#sƀa��SB�;��t��`��yˌ���hWd�3��幀���*�7�9�A��ޤq&́�����Y�5o��?H�M�Ra�i�pTh�L������΍��>�3�����$�����"�D��ƈ�i�g��?M��V�mg�<N"���,����|�7�� V 
�QZR��&J�8�����d�;a	Wzp \�\�)B]*�(�Ʒ��5��N�5ԫAL[H���E@���$(Ž��ض���=�T�8�Zcj�C]�;dr�%����@���$��Ke������XqN���ҐXlxVHYEB     400     1f08�E���L2��1�D���� rfk�V:�h���ID�܇FE{to��0҅C͜��!�5�ƿ|l�{%=2\f���Y['6|������3W������U7$c]f�o/C��'?�m4+qq`H8�QQd	Ԑs��-F8�c1���}˨��\�UY���j3NqS�7���Ip���$k-��/@��F��N�h��?��$8��J3����,e�-�J�#\�l|@e�d��M{��)[���_7T���rS貤g�m� wNS����,�4��"x$L՘�^�����>k�C�����9�O��K�b+k�y
D������
����&[��:rC{v�[�,��w�|5=1ӑ!$}}�-R٥��C�uA��K�Izhid�vy�@e�i����aq��@X��J���̝h����4䘉����aI����f.J��V�`�m�a�$g|�R-.�м��p�~�Ə�B�S`;����
c��M��Խv�n�ᓬXlxVHYEB     400     190��~A�r�Ҡ�W�8`VW���ca֊"�4�8f5��H�l19>�e�J%<��
�{��^�	d$4�TX�6g�_�g$����zJI`�
�\=˪Q��4�$���o�ű"�hF��bW��κ	 Ԡa����(pO����Ң��m�vq3���ݢ��1=L��)��j�mh9�_m���-���]����W��S3�j/�ѥ;q��ޚV��I����3��ނ��ڂl2��>OD��!ވڑ�����s"���Z@��M���%l���^���?<;�����Ou��w�y<��S�}���)9AZ8g�E'z�~��
^�w�sF�|�)�kGj��GW�2pl�U�J�e�z�����숽���5�Q�sZ6;�T�����U@�U��X�F�	cXlxVHYEB     400     1701=�T	7�9��
�4�[����+_��'��9fK!�v�7�1c9��`�A��Vma��}�圣[O.AcA��!�D��u2$��U��?l�{�c��)),�	f��#R\��RY�F��K���e��i%�h�B^�t��IՓ��C����¡k�z�v+�������~�g\W�^�<*����p�А�u{6�,�v�F�H�r�)��O��d���v�K�u����T !�����>���d�����Qr������JȰ�x1��}���e�gZ��GbtO/���qhH�Ѷ��iG��_E��Z�=���h�T�a,T�Ο�uĖe������8���7ղ�ߧ/�C�A2	٢ �g\TsXlxVHYEB     400     170�<z��h{.e$ā��8Q���&F%��/�R��.	W�]6��ԗd&�y!�����9;��D��3k���u�v����h�ո�6�Ax�z�;�QBrM��¯�P������5�R�^g�-sO�9y��k�TY~V�
 r�e[]T�e��v4�Y	��`�����n��������W\���������덺�S�����Κ�>�k��i�c	��8Ҟ�����4k���	��V��tF��t�^*��a91"T���S�^1��P|���Ä'A���e O��K����/L0d�O���_Aͻ��)w���f�"ZI��c��.�P��!�S�B�v~8��Z�}:���*,�;�v�ɻ']#�BXlxVHYEB     400     110~�P~�oe��<�K�Ɠ(�[��d��N��B8��"P㗭�
M(�]t�>��T�6	����&�.���#��}�����pҥ��9�q�����6GD|��5lش �DX�h'd��WX��"�a�/;�Xw�k'���0Q_4���'�=���DyO���N�����'��sn���39r{6��&��>�P�3N���U*���MW�x�EF�!VRB�1h�K��z�N�v��"��錱)(90N��%�͆�Ubc;C�N��3EXlxVHYEB     400     120`;�*���sr�X-�Ư��x�z2���	����{��{bѥ^j�S��k)Cn�E�s, ��%(�;����!�Y�� �����dc�>ݦ�
b��A�L8Tș/Z{��~Ц"�|rsHNQ��/��A���CO��^�┄G&��n���f�>|�\DsM���Ŗ�^�:ۗE?���2]�M=��]&ؚ�}r8��-�{��}:�G^����8!+#�6`3L��Ԁ� D( ���L����[����q�} ǋ </�5g��I[ᨑ��g��q�r*XlxVHYEB     400      d0�c(������콂ju{,a'��$@�K�%;>
��n.D�]>��(�
"���f��9K��@>(w�V�9x�ǈA6�z�S������b~�<��O�\�ۣf�QN�H�BGn�6�_nݞ�2+��=L�p���=�~5*7�<=����D�|F3˕yI��)[A��5��O)��G�)A�]p�8� ���S$���SR͘�XlxVHYEB     400     140c}~������i��VEj�P�	k��V�aĴ_��-x=z,w�*t��i�]���@��OG2
�G�c3�h-���[bȌ�Ϥ	(J���g����rH
CF=ٖI'c�0��p�;��!�g|�.��'��:F׬j�g8�M鈈��w,��nL�nQ)?A�B�Ɵ@Iq9��t[8[8��&~��g"��������sy.���O����u�}�D���Z��~�ч�Y��gq�(�S)/�����ʱ�e����ap-s���рǺ0�V��d��%j�5�,�9�\zUdo�l��Ga�?�sN̲�գ��������}��}Q��XlxVHYEB     400     1406U�$z̺@y��? ����	�xP�^��I�,�?gu�۞$E�&PM�D4/�y�LZH��G��ʜ��R�ͯ�<�"���6� b���f��f%�tt�[�a�ނ����}�I���U����0\��F6��`��m�m��q��+ҥ��`F����X!�Ƞ1s����W&y����	2-��m;B�d�I�&���`A����$�^�M��)
V
����>_~T�d�n\��V��F��[oE���#p�A��TXZ,[�Z��*39� ��J�'c@&�V�&���䤁���n�m;x��1�K7�2�d�;C�|�2�c��XlxVHYEB     400     120B�\�ï��D���1@s%��/�X���� l��`�2��G;��B��;};�11G3�>P�p�8^��^�IF��ڥ�`#<<V%���zTK������Ҋ�Z2|W�OR����_�,��`�+�=���J4��o�C���HJ�zt���1h���'�
��y����h�4E�D�!���sȿ� ΰ_�i�K�w>d>�� 3{�w��˩�L�@�s�$��7�o��5��X�5z[�psx���@�tǃH_rs�K��/�%���`�c�c��1\XlxVHYEB     400     1a0����I�z�cj����K�I`���u����A��	
j\�tо]?HѿW���:��:/��Iyg��kkr��?v�!	]��D�6#��4��7�t̤p�Y��I�~�����@��B(��80�0*�#ז>:�`M��"� uTd��y����1��q�"	�qw��DS�[囨i���R���;Y �) ���A�V��t��<�T��< �gF�a��� H�YH�]ܣ���S�z�y��b�͐����z ����ǘ�d��a����l+5��/��Q�1PVx�Ձ���
�"N�N�>�wܿl�[�+�[�'�|���e2�K�������`�a߶�e�p�{�uQ��	p^췳��ː�w�J��c�m�^�,:`�W�Ob	77\Q#Q�e)�]�2��΁���j�XlxVHYEB     400     1200�F�ڗU'�F$��h� \��%F��Q�*ǌ�.�
X��zB�K��ũ�m�ӈ T �Vp�>7�t�d�����|8��eg��F��i_�H�v��N�������C�`�$7pݨ�* �I�Q/��ᔊaŁێ-m��F�WZlp��AoY�I�CK ��E��ܵ͞�*L3
�e�ϣ<_M��뫻G��[��߮�gE��I�߂g\18����Wޥq��.�W?$���Q]ib�ޏ�),��sJ9��z/*�upNQ�G���Ni�:�,��J&GFw���XlxVHYEB     400     180��%��H��Ț�i�Qۖs�~��u�V����%��.�}d {/2�{�G���� z�Ӵk�C'�[�\����U07�6u����yV2��p�d�
�<KJ��CZgYd�� �����.��.Ԋ��OmZ�`�A��`!-4h��X�kD��ӓ_����!Ǔ��.w/p����%��Z�N*��[��T�8��'3�]X�%�s'�"���&��5�������k�[䧡���T�3�d^x��Jw_,����x)� 1#�p�ģpH ��@
&O�,ΥGΞA���1�P����w]���佒kZ��,��P�U� _'1:*M�{� �����G7�Ǣ[���ڕ�oi�b(�n�q}(���p��XlxVHYEB     400     170p�Z6�e�Ճ��ġ;>ꀘ�����z�H̞�)^,4���n���b��{Hw^��l܁���x�̋�CU|3�9�J��mV`H7��MQ{iW�*�'�i�hO��+�����vS5��aq��(�D�7��Y�u�r2�(����������rh~��Z��1�3%�%��a�>��6�i<h��7��Ȳ
�=f���Ŕ�=.^(۠#|�i�i���w�3�H�$��h�{�q"\����%�Vb��� V��9��X�f�����d��+���[�>�%|��
An:�Y�=7.k�zsZ7u^E刪�i���tk�;�i~������f�A�H��"� &4�.���nB��\(�:���XlxVHYEB     400     1c0��2�e78���E*P��+�R��Z����b���K��7.� �)�kM��=�[kסX��ZA;�S린���?�o�y�0�ci*���ݑl�<A���~�`����"Y ��O�0��p��s�|�����7���ԅ���s/����r�\��,������H�s�^�H/u��d���(�W�	2O3�ؖ��@1ߵq3OǑ��?3��L=*��v1D�t����/j�@	[O��;g�p����B>v�U�&Gq��Hտ7t�3���L���8E<0^�t��O��	��̚aH0�̂C�k����7�*�3L�W�������l�6s�	Eo=kfl1���H3���֍��(��Fm��ߢ8dӖF��j��rK(��HU&��1*��u<��j��4��#<MW.9Z�,��Z�Z;	S;o��rEw�e�XlxVHYEB     400     110��+;�Yg&i�i$۷)��x�f�_����x��t��Jbו�床�O�-JCޠ��N�;�6�A�? {��*�"�4��K�<�����Bs�YO8%bH�?�eE+�`�*@����X?��vc 
����-�*�x����b������k�Z�}�|�g��;{���(zS<�B{x��{�Z���k�G]�����|w��<��w�&Ww$�7x�3�&A�h���yx2Ͽ��1 d\m�m�Po[vH� "F�Ԁ�PV���*$%�BXlxVHYEB     400     170O��+�-��_ܭ�ZM8d����T"���m%� �-��}�8�1���|���ck|�>lYp� �~��Gx�4��[ě�f�o�a�%ai�D��L�%h�p�'5���V���`:� �N��ǵ�F�b����.��:��H&~�$`��B�6��e�
frt�ͷ���c��vI�b��$&^�w��:��;�l��ʙ����Z���C:jw�u�:ר��V�d%VQ�[�����sg��wg]��.G�Y$w*?�K��X�1�y�©xL�	��u�;�(�.mf~1E͏g�x\�ڧ�3��f'u����4שb���C�3mLQ%	:m�]	!�n3u��~�Ֆ"cAz��(~��;Jk1m��h��LXlxVHYEB     400     170n(��%��7K�؜f���j�İWV������wf���EK��^�gSC����k��כ*)I�ޓ�Z(^�?2*��f�g��y�����OOf0&�2�uӕ��}�k�V}���8��)Ief�ۼs�8Gb�����4U�f���FW�:7� �Ԛ���Z��?�F.Ģ;z��j��ӗJ�S%�`i;K�A�)�c����f�����*����_�:�NGLW!���D��?��p�<0��)&c�	�6N�Q\�)' �LҖ ���Ki�A$?���>~f ��J���\�B���M5���T���/`�v!�R*���_��&(�/�^+�yX,JzN�gUj
O���j,t�a���(-�AԊx�G|�XlxVHYEB     400     190���g�6��P���ܲO�]�f3���N�n޿���I�̇~�/�viL���u��]:�Ή�xW�&�E��-۽`�9��{����>��d`P��r�c�c֝e��'�DG2��thI�roWD@�(# �b�~�b���j�Дt.��ʠ�G���,��v0E�n0�ZS
��Qvg�i��n���͌�<)o�xQ+�@
{+�٢�|.J���/�{�[�����5U�K�g�FvN���G�yS�N�!�z,�&�*6@�o�W�mi�J��]_������4�²L�W�7��ȕaH�������:&^
T���ُ*OO���8,�5ǧO�GYk�i�����̬ר�ZWݾ7;��Vw�
�ԋ�$ć�եh�nC ����V��u�XlxVHYEB     400     1b0�:s�~>�� �>=Qd|2?���)ʔ�ڲ��syO̖��g��gE_{	b�cn^���pWa���zn=Ǽ����>w|�Dl9*�/�Ӡ"X�Y��E<��F/�cP��c���y6%���R4�9�^%i�Ќ*<����ʉ�r����nfy.�k)�W���aT�n��d-�r"�N��6���;�CO���<��Q��O�I��A:\.�.kZ�<م��V��!NR�o���� D����	�ȵ6D��S��ꪲ�߽_P��V?�(ع���Y���,Bza��G�����X�>�^q�N�b�Ԇ9��!/��Z�@�X+ڨN�|���B�\[�C:��W��D��A$�u�Q��\:Ş��H���\Td�ϊ(_���}�]��^f����)�s�N�u�ux�/b�Kh0�� $�8��D0CY~XlxVHYEB     400     1b0�~�/i�:ǡ�l61jWϷ�sI�
��(nʈ��,�
s�p�D��oa��Ԭ��V�o����Æ�Y�h��KRן���(��{���Bh��#U���旷z%��ғ|��~4��
c��2����L��$��\��wg�w���wp ��P�ɁӉ��s�=��HEPy/�lӈ�����^��P ��4�j�p�}��n��{��b�ǵ���b��GW�|<���"�%֏����8�f���Km���(�BΟ�B��z�Z��*Ӓ�E�\I<��t���{e.��O�����	����\ �(�����X~�l�k 0d��L��(���S�i���� �Z��oLK���vg�ۊY&����,b��"�0�YW]��!��7�j��o�=r��/���v�D�i�
Q���G�8�+kG1�y�uUXlxVHYEB     400     1c0���&/��f)���"^KA��{�h��6���I�b�����+�)ty݀�te.M��~d ��(4KM ���q[v$�aS�w��}zs�}9p)�P�L�Ol��X=��fr�떾N��pj�e)���az�M�9ۃ��ʠ�r��$u.Ź 5S8:�ʗ(hϼ�7��i(Zo�?@�q��u�_���cxGV�tj]��f�� eof����{��9�o���ዖ6�r��[H�>H-'J� ]a�8jOy��ۂ8��2mO��M�)�xa�O{������H[�\?�U��)no*ws�i3K⛺�x:LGd ^�;�Hb�/����(�i�h��	qAR ��ĺO/��^әR�𜨁M��O������z2�}� ����\o\�Xn5�,!h�L6�MP�7��0��N(�Fh%/ڱ�le[y������*�Y�XlxVHYEB     400     140Z����H���%Ȭ��`;��9���#zZ��_b��g5>����J�r��ZB	�x���7,f�8�*�V2I�.�^4q7��װ�(�YšXe��?I��sB5N�j.�����8�o�̕B'm "fG��(�&�Nemm�)��@��j4���R��4�崞���?�Z������|UFdӶ�0
�`��hXZ��Ȓ�̜4��4{r&�hD�؞���_��c�-�����faS�΂��JN�~>[(�41���lm�t9�e+Z���b��Q�d���P�&���t�c�R8o�1ⷈ��`N��L$�z�����R��XlxVHYEB     400     190�%ڸg[�+W3�X�o�3�=@}����0rj��e�*��L���2T`�a�h��̋)��ڕiHg~��>�������fu�ڥW�V��F[�3�(rx�L�k�TD�+�CMJtZ���P*�����aͲS�WSC��������)�`TGQ�0�j�d��;l�`��L)k*���_!a��<�m���P����/w�D��w&�+�!2�$�Do���h�*Ϫ�(��W(��kZ�5��5�*H��`\��8�O�k�jߴ�/�e���Q�zms+��ys���e~�t���#����}��)?V4�l*��U�V�dẽS4�g�,�>����{M��JB�#�+�SR�N������,�
��B�=�7-c�·`ڟq�XlxVHYEB     400     130�#��5��m5U��L�ګ��AN��6��7�G�gb�U���h	��1�^��:r�l�f�q�2����\�K$�$�Bj�xz>]Y����t+C��E�Ǣ6����0�\�h����"��x��<���s�,a/���Y����9S���Jb�T��֮�����*b��ڪ��,� G�V#��Yќ]k��̭׉vQ��ս�0�ʨ���f�z�L�F��v)`8y�a=K�)�#��	�����w�Fxy2�$M�EY��4�� ��Z�Ot}".����W�6�w�e��;*QJ5�#oCXlxVHYEB     400     150����E$�����$l/f���F��p�h�L�	V0*p�hi����h������ۜȻ�mj��fJobk-������-�T�j,�-�ץ���3]7�\�3�
>az�9�A)\c^X����ѩ��Uuh2i� �7�M��E��_����u}88U�����o{�5�x��51��X�I�i"J�ѓ�3t
���1
RM=�(mf S��}�r�A�^���=$�� P� ��[�~ ���3���J�l��w��H�Y�ّr��}V�?Ƃ+h9�7k��+����ZݻRj��Z��� r<I�Xts=�Y+G�WȮ��7�"
_XlxVHYEB     400     190��(�p3DX��=�x:к:[߂PAvr��/�_��޳����BϏ2*J��e����U���v�]I�k��5�XT�O�ҿ(��If�쑵)\���M��S̛[�e�b�cO����~�z��ȵ��Ī�*�&^���s"	Ŵ ���j�{*���_�pn�+�����t�>E�Lz�w2ԸI֨�y���Sz���������5�7c/��2�}�mI����qI8,-������ܹ93L��B+��G4S�S�E����=Fy��>eu��*�1X�d^1.�n(��n9��MR[�P�Q.�djM��l�[Բ\P���˙o�qQ�[Tqq�0v�-�u7��'����<-wFv��$��0!</N�S[%�`�`�xֽP�F�e�"�[f`Z��XlxVHYEB     400     130[mF��ӳ�`ҵ�|���@�A@(d� ��N��L�u.4���^<'�	���9Dj�i]o����9��;�+��"a qsYj�A�Q�x�z�⣙��*3��\��
=�0$���N5^W��p:�IA���jj�D�
R'����Ot�2���� �6�q<10!���O����N2aC��4^��cΈiS=Ʉ��i6�����̉Q���NP،\	���Ņ`I8BE�� r�f܅)�K7��6֫��1�2�����{��?2���6����-��fOvp�]~%�д]��XlxVHYEB     400     150EO��b	پN��ۗ�(�K��=o�c�jxp�x�2~�2]� ȵ�PP�x�i�s2t�P/������T-C!3�h�6�W���f܂��N�����`(�4�v�8A�?��+ڲZT��8��j�B����7���ދW���E[2oW�z5~�n/�r��U�X�*�r��X�e��m���ZT����uf�������ޢ���)|��QxP^~�qG|��7�/\�ag�&��+���}q}$A�&�����7mx�I�i�J�u\���T �&�`y��x8됫��Q؂f��Fc���\WIk�籃R��Z�O�o�m<f�?� ���aF#AlXlxVHYEB     400     1b0}��&��J�V�G��>)[�V����~N̐� ��WYa�n5׏Z��=# ्7f}�:K�x���/�cr��Hg��oY���G��$|���s���2=w��uk����Լ~Ts����*�Ȗ��n�P�n@�7NT4-�{x�Kr�Z�P���,)P$�J�I�mQ���A����oM-��]DEv~����?^�9�I��þ�С@!�Fߎ�s06���	��H �\��g�t�\��hK����4��b�+;���Q�TґEu��7��ts��J�a��F$�	X�lgN��l���8�%�#�`L�/�g��eR?�j�%Z;��;Rl.5�0�;@�5�,-G���XMZ,WZ����c�����}˛O?��8��6;���0S	�y����� 2#�C����F}8'r��2ueQ�XlxVHYEB     400     1b0E}�K�)�8�������mu��X�1Ҵ{'�^_�Ol��ˏlz�<(�X��g��D��t�c5{!�<��(w�Jm"!�
���,�w���\�T�+M�iYtG�&�Vt��KP������g�޺�F�m-�1v�����Lm7ڌB�[	��A+2��ӣ��}��&[ Wsnk�#�j�����;��㧹��mp>@,ۡ�OC�X��ޕC$�nO��ݐ�mԬ�d��9���(E�F�#n����E�Όl�͂�>��I>@r˕y�BY��,����
�<��6BZ��kJ>�&{�Y�+�JBs����f��_���/���y��넠����ۗ�S��S�v�����e=�3�a�x��$SXI�׌�҇���jk��:T�p�R^��)�l'|y�2n��#����b�7|q��Wo�8�XlxVHYEB     400     170$N���+Z
����uf'Pd�5���P���=`1�ӗ�����������h5��-�F�9�mF_�ٌJ���M
�'�g�Ç�sL8��{�*����)[�V~ohsA%�5X 	�}��PU�N�b����3Lm��Ԇr�4����P���U"F>�U�m;z�H$Q�Y
\�����f3���̃VW�O����'J]�07�9"P�_��Z0�p�k�9yG(|���uwT=�H
���}:�h�����%i�2�j�g�Ru�]Y?b5s�2;��*��*_��AFcLJ���������~�a@���D�]�,r��i��.�/3�y���b�����O�a?�aD^�Ϗ6�	�[��:� ������(�XlxVHYEB     400     1f0�d����QH�(�rJ|�����/n�[�|L��`�J�J��w��k~���+ڣ.z�_k3b�l���EN˨��ɔ��"J�WR� )���<����b�1+��	g>�]E�`z����^���,ܨ���ccy�ݽ�n�ok�5_�'f����V���A�;��g�x5w�U�E�vs�>m����3ڼ�����v�:�On�����(A|���jp�J41���h y(��\��~��=.�@O1����ۭ�� �#�5��֤T���T�F�j޵<FP�)�� ��8ﱽ� �}�]/e��)���ӯM��"�_�K6���X 	���٨9�D�԰OV�.�z��il?`��Ȫ(O�mC^/��c��y���e?X��e�(66�S�8|��3hh��v4O9���rk��/.�6�dh�L^����PL����&��̐o��	�&]}�%�ghcAj�)�AS0��U]����'��C�kXlxVHYEB     400     130�3�d&�&l���P?Q0�(e��ӭ�'"OxRbv�����DO@�c�Á�,d�}_?Ͻ8%��,�~�f��������Hhf$���{ ��lf��kXm�ܷ���O-�)�$3Rߗ�?�����?���j��s����'�T�nS⬺�.�>�ijֶ/,���I�!�BH�-���y�Pd��@S�j�� ̂�<$ø�A9��ε�<�!�y-��C|^���RE��W��YN�PE��a�Yw�1�
z�9�Zd�㑹"r2�L�J0�L(��!W�Q��h����g�H&�q4XlxVHYEB     400     190��+J�q��V�Cv F���L2+�Ǻ\E���roQ�+�jU���/qi_�}���wo��!7Jv�ރ> � �?��}���oSU	h��wt'S+S�,�4��Jt�� ���*�$M�z�w����sz�U�{v���D��͍�>�_�)E
�"�`��4��*UV �����u��AkY��� ��d�:o�f��V�D�2��݃�;V����8B����/�,�����I� 
R�r-�g��H�כ��>kG�RB|��v�5**<����DN�1^�֗N�9X�����@oc���Q�<4�P��Ҽ�����ٍ��#ٔ��GF�_�N�Ĳ���Oy�7O�V�Hu	���"��?�C�SR�R�_�H��[�[�9F����)}�ٓs@JZ�XlxVHYEB     400     190#�.k]�r��ӾCS������C�� ���*Y]1����C�����"��C�0e
e�^<�m����QuX��օs�ɛ6�4�3e��!�$���nٹ�%�jD	��{���*�5�ܡ���6�;֍$�6��������a��d��jJ��x�0�Zg�m�[	Yf��0�~�H��Q��[�6���4M)�o��ӰT��q�yM�Q}���6��d��[�\����n-|$�4>�������N��`�:�0"5���[��y��Uǲ6@`��@�Y�_������#����W\��Tg�`�5�!G��8ʿ�/�� _��KX��I`�[�OEZHJ�*h�ߦ�u�
�_���k�t�A�H�~��=7����%��<�1r@��ݔ5��RXlxVHYEB     400     120j8�H�ЪL=\J��}ts���Zq�|�n˲-�b�4��
�3%�d�ȧ�oD!̤��U����L@�d�RB�Y�'��-%Ǹ�z����s�cɩ�l	�D�pC���y1;ظ>hZ�Zͮ�ʽ/���C��)�WMc�ѽ����>xL����A���U�TkyR��;�H��6 �*Y�����1+�K�x8��%^xR����|���N������F���#\sW�ZAPj2b�\̩�9A��C�8n*�"��R��!�[L;�og�ex��Գ�/A�!�|��M�8�XlxVHYEB     400     170���Q���˂�wu�4yJ�ތY���X�����떪�'�J������{A𾄝4mU��e��$�:У?�6��������!��Vl��U2�j	��ƌ�Ƕ���'e��U)!��x(A3�A+)]v�Њ2�W�R��*OY�`Xm�FxUz��ίm�\�޵xa^��/1�,#�v/��Ϸi�/H8=�;:[���e�B�K������bi'�����:�I!�ߊ�b�^��,���.2��=b�ۇt�>�"yN+|Y����c���w���v���F���kH��>�D	����Ou6I�U�>�Xz�E� [�ȵʵ���(�����~O G�k�d�ۣT�tc���p�K� �tXlxVHYEB     400     170ug}�\d�d�rȗES�EU�y��e*�e���;�=; :dfc�@���MG�����BD����0���2N��d<7��������Lc��|�h��W�m��@�w�V|�>&����0�o�-�z����ׂ����u�ȭDC�{N���rQs	cʂ!�C�T4`|��\�jO;��m������^��'����|���0 �1�Y>Z�pC�ˡlp	b�53���ٙ*2�Lv��p9٨��\�lZc3<��=Q��J�:Ð�o���s�u��c)�Ǭ5�*�h:G���L9^="����\�)���8K�*m�Jg�O�vt.�r"��2>gY`J �Ѥ�k��6����9�P��� G")u�wXlxVHYEB     400     180�q8� �t��ehSH_�&v9���B(����*��S&�Xo�(R"�ʹ_��w��ٌ�����a�x�;�N����,���FW0��I\�\�ʇM#Y�`�����ܯ_�� !��m�۳�x|�J�U�pB�!ɼ�	�o��Z�4o�P+h����+x8��\��%���ф#�Bǟ�R�
�}�Ӣ�`��2�h<���<�a<���8�^5'�ݛ��j�W(O�Xy�Q��e�ד�y��I���ܠlA��}6N��t�/}�C0R��h�ov4�x��C��vQ�l+lK7�{q��wz�k}��fa��Y2�ܷ��H�(�&�@s$�0�3��������Qo"��1��2k�WӵX�`\���9�\gR}�%��g�ԉ+XlxVHYEB     400     100V�������t`���/���M��<ب}g_,�썓_��Lr� ?���ݤ,�ķ`4�Ӌ�Hu�һl#	�"֗(?���U�<6"Y�
/����	[�<4t1�$�.���!�K�J�7���}�uk�U����=RP+��@+�t��(��i���|�a�L\8��6(��֞��2�;:ӏ��)K�']0&w�Y�P��L���aR��ɢYe��H����,2�D$o�M��}�5.���Py��XlxVHYEB     400     150f���+b�&�Z%wW�!%�DI/$5D������pw5��ٟ��ݡ8k4�+Ksv�-�\�1A�j�]Yč>��k��P'�|&��L+~�
�Ҹg�&B;���Q
p&n �gh$�6�6y��JYkg��]��E��u��;��|���E�(:X�1&��fҪ�ߢ�On���MϦ*#��?1}�<�U�b�y�t=�:]���
�:�BI^�2�ͭd��Ȉ�/�y�iYf�#�2 d��^K2ᬭ`���ե�$��L���]�q(�r���}޳��\���p��zdK��+`U��l[�,O��G�9ka���|�L��^vv� XlxVHYEB     400     150�}`����������"b�O���;S^�.���R���������4��y�n�X3<:{p(�r��f��]Ѻ����廹�2
wݽ8K��=��%�d���Bn^�Yj�eA�R1�DӴ
����P�$v�I�6���3K{�&�A���C<��.nR��n������L�S7���d?��'��W!���	3��;[��؉��Ve-@@ZI)�'�������=�!s��;��FF��!@�ԧ5ޯ��\���:|�t���N�yht�ե�S����pb�3I{��{����Y����Z�46���8-I�K�$�}N��H�W 
[��^���l��MyXlxVHYEB     400     150��cf��iٕW�ݏ��O��iQ4�Z �M�+f$H���(k�m)�#D�*h�2�;���n��|�yXZ�_���]�)
�*ݛֹl�9��Zd��6±�5#��4��Š��J��U8�^
�M�NJ����-l�t:b�qڲ�h0�
��>s��f]�>|)b[j���+��*/_��'��ۮd�+*�� �Dn�mW!]9��)���#����:��~�ٔ[7/�\S��_Q
��(��;S�OG�<Y2��V�Y�O��z+w��5/Jk!9�FՃ��k�牛����@q� ��ȯ�<`�͹�Q���;�	�2	m��=uXlxVHYEB     400     180�/c��X�*��.;�Kb�xx�ߓ<�(��Ƚޛŗi�ͷEHH�",�(}~�ލ^�N�l	�������h +�����]2�I�EO�L̔��5���fc�	I��U�>̷� ���Q!`kH���ky�9�hU��M�%r#SN�:��0��w��� �OY�JCM^Vx>�������-I�zy�oV�&ɣ��1��O)�"��lҘ����+c��f����0�xy����Nb 'ou�%K���G׮�ovw~ܦ�xo�b�t��g䊳�x?P�6*�No�&UǉW&��^1L
�5gl��f&E�zʴ�8�ph�sec�c�A'��s��yq��t�Yx?��6�f��pJ�y#���XlxVHYEB     400     160/Ѳ�a��Y�1�V�`%>�������V>���h���E��Ĕ:�t��9/!?��8��/ ���	V1��N�wc�#~�"<什H�oN��zA�&��vVϲ��;��I����s�e�7���m������X�#�9B��# �_��V�
�����ߚWu�V�?`��M{0�$�p`^�=r�-	h���ܥ^��$�tѡ��[G��n�:����l�k�d�#�ώ��C6�R���oM��>��@˼"�K?���1g���)�'9�\k��tM'����Y�tߗ
P�	��Z�`ׂ�X���1�j�U�S��
�qjcv�m?��VXd�B_�RQ��k��AS�����eXlxVHYEB     400     1a0sB�,��6û��R:�r�&ى׾W5���`�_��)ɐ�3���-�s��N4��g��㩡	S\=s���~��bT5�ա�~�m�V�jb�b�w{4�n��HH�YV����]��H��
o!K�X�����fԊ���gY��=ݵ@�6��Q2;#pӍ�E�k)}�Pf�����'�I�����m1���ȣ�!22�� AJ�F�^���;1N�M��+T �_ulg��m�6���5=�rC��jrq[��ݔ�P�`��\ת���V~�����������]*�-V����J
>7���B�Y���7�n�}˽���-c3����a
I~��js��80`�¢V�������)��T����z�&Yv�.�O@�KE��^�Lq��1l�X=��͝���5%�*�ӷK5�XlxVHYEB     400     1f0���KaG�����'ڠvT>���I�����oZ�{g����!ҝuJ@-LI��cơ�.q�O��9A���D��aܜ��:��)��/���l/F����l���Qv4�����J���m3t�0�O'�IG�5SG�ye��=�v$bI�=��8�U��L1�R'��NTD,? cZ������R��1;��G�����ނ��HOYـ�z�]U���3�wP��!C��1�g��BS��^m�_#�ܙIuZ�E��N�g�����uEN���K0SG��BV�p��6�r�,�ˏDшv���(i��eV����EA��t�&I��=�J�;cǝ���(�Ô��JG��%P� T#�C3PH�$��iorυ��FkyOH ��D���[ha�85s;��.V���.)QM��߯?-}�T�F�������J����>���xn�_jL�K4�����sn�9}=�������/p�s*`c�>85ɽْ�������(RXlxVHYEB     400     140���Q����%���q��\%д,䦋.����D��̵&���{FJy�����<z<&/���H��d�"{*���k����z*�y�;���[�U轎�6J��)&}�)��&���K�6�ߚ�d���0���Z�?��@YE8��h*�m��P{��E8�!�`�dq��A���d�G$����q�`���;�|1��Cv�QL ��U������Y/�<�y@<��Z%s���SvTs�z=-l7:��@��=�>�o���� �r!���F�{�&� �dV�p�$�`a9*��wƶ~�Q�n�ATod~pXlxVHYEB     400     140�q7bTc�5��X�/)o�5Y��B4�4^̤�q�e)GLKf��T&@�׈���f�Wz!��	��u2��f��sH@���}H��1C>c��b�u7�g��ۅ���
s�4���)�4��[�������i���"�M-Υ��T�O���c뼂C*��"��ͫ�Gw����ý ��HsH��3��	Ӥ9^?����u>F�%x��K���SCAi�[$$����Eh֕{l��
3�To�@�.G���p��˝�<l�k۫��Ɠ	�n�8t�Dw:�cP/)!
��Z�e>E߃}z�w��E�Wm�XlxVHYEB     400     1e0rG���7B��U�84
��?0�6�����1�T~H��,��y�-�9�(�{R���5sCPS���c���t�v�/��N��Q�X�J�����-h�b�z�-���Q�N@f��Ρuvם�ix�_)Y�N��ۅ�L��^mEJ�Rl���� ���c�e� E���L3�&.�i}/7����g"(��:�1vl��K�b�U7���KG��1�b�I��w�W��!_��_�A����Ue�p]F_��z����o����a���5�5wCs������Ek9�|�Ce�B��{�r<=��W�H�ͦ�)p�XÅ��P4�r�#�滳��*�<F� �D��4�Pq���)b�t������%���F0=ߊ�~�8� �`$u�:�և?! d�.-r�,%�?��2Tp[)����� "��7�����\t�11���_����J��h{�%ȗ���r��WaX}%XlxVHYEB      90      90�玄�s/��������`<
k�9,�L�H�%6��>`8��%�$��&2��1EK����S�[�	>*���"s�'��(t�e�8����_�˂����)��jg��<�����b۫�뱉x��Z}'���`��ʥ�
���a