`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
+PjWzNHoyzrEj359FVFV3hwN6NWEbHpPxhiH+0g+0tIotf+NDRMGXx9OU36uQnB4wL6Ou/6TEnfS
9YK2nkdq97D3c+m5Gp0enKNY/ftTkdSCJLJSi5d6AAVQbBrZU86ZjAU6jd2arPb1aK1sYosWDrls
JhvqKi0p3cTzr7IHcNSEKzbqpZyb9JRzf78nz3hKfY7W5z95OO67oEaMUTbW6TIfhN6tuxdecBms
P+cENlnvIb3t3Y3uOhnttbwe3bLl4dQe99vhi4Aamy4vlyRTKyaed5TdPo9Z3kPH7Zwk9JavVrMD
em1zvCSAGEunRyqgAa5CQDgqLJZxVu+C39cuC11TBA34WAfdABdWFQ1D8oujtVMAeRXpgWx08eQu
U1/J589TCW3l1Q/wJ/eilaowT63XHnXV7pmvn+4j64Yi71+VpFLhG0ebYz4IiaJiGbh0rec+Uc1p
LNIu1Epv1vreqdO0NVG4YdFHgp2YvtAJv950EZa3E2IOWeUDAeQCpFDhTOyVjrs6TfccbQk3xJtf
13K/0t7XMkaA0PLIUUh6WsKK6uvFLsp0si2JnRy30u5b3+zSdBaj6CG+BZX7WVkc7YI/0EGEZhlB
PwzV5+zNOojfElTs/p18ujYd9taRftlG/4YKjPgelybNHwrc2VDb0tw3I3oPCZtIswkjtEr0/6dt
jdl+5F54BVF5h41uNE84IjxNTDh08v8VyZ5xEpzm0RKEr+Pb+FyZtIfAiGUi3BhlBCARxBKEQ1eO
OX0u+FoQ6jhBStScFbw54c8R1/HHTZpdYiLuPN+uv1Rrxjn8oSLkyBERX5CDXc4m660+XSqR0VfS
khpr+lGRn1C2UC/LVtrd68KF8oY7P1eKsHHmf1OCOPbt2q2ngA2RuXc3HrCV3kW/ImN7HAtcSA8B
AxgIvggYGWL1WrCgX7lLqJqVsBAq0KKJpgFUD2xZUyviMmExJF22pkmuNqbmBn6zzi01ECC35l0Y
UAkisVTSEuoe7kqpZCZ7iYkEitsUoaps1nFH3ZMoVwMzEEXz/+FX8Ro8UOkeiF8zvortsC5tcKZc
D0CI+gQjXapt17Kle2F8y3pbgooW0kO6UGDD0Pn+cHPwIb7AZKfn6GyAYBuT4hZ/77CUcELzV3SY
NSYlR5Vhth3qtMQxqZ8poTFitcgQ/W8gqltmoUq0Lh5/YWOFPaq5I2n5xXVw3tU6euuat72StMEh
OA7P/7fi1IowsOKDjdafDcs/TTVLksvGWPxCKmRVpmTOQ4EbW2wdXrqr3PNPCFhR3qHJfiFIYnJ7
GJTdX5+Vl3JTEkV/TbmK+RSMK2ZAWfc8Bu3bPrUbzhhXI8n3WWxP4M/rIHM0a5OYPcBTr+lWDSCb
4+x7E5nCTex8ZhahuW01CIlrCh2sjwNzIEF05WsD5mh3f56iWm+2R8In8t8wB9c8btbGaOmg9PRp
g3dCm1sk34MQTVjMrWwAi/rGOmbV1aaqgl+GapadCoIKhd9m377rTByMcsK896FteCqzTW2J/GEo
paVfyNzwkhnHyaVtrBYefwZoCDxCsrfzlIb+clsQs1KJf22WI1tuTn80AFTzHUetjRofjymZ1/Sp
at1hGDQZW8Ruxp2h37nJROxw9o11sSkV1mlPrlaUyICIO6GxuQQFd1ZR0Zp0u6u2PZWDqOFxjYyy
+3GVZ8+aBLUG2fqKLnx/ASbPsblPPvg8Sbud/tw00YgMy+1aUKxrSCijNJr9f+r3/olCfUwydMij
sdWHQ1Ia5JREe0vijPj8Zw3w5J8RPLhRHXNRu2kYz+Q4CK29TXhmbfpLTPWrxuPrcG3k9ADSwxeq
qzIAUc/vC6KZ464PB1TU3LUk1rKEzJ6FJXkxyanfu6pbQL0jzzm7k9PZA7LqivkTmZSzy9E+1RTD
kq45wnbs8ihdbbLlUjDG5YdmQLDrPwirU8Dl16QtZnA7s4vpKgUR2qrPwNJ21GtdzgBzIx93Dlnv
jUqYRmyd4Y8nLRaK4OSfzrmbVhlIdkDwB0P+6Hw1UAXjoHgV4DymFXd2tjg1KR6kjVkIcbrMh/17
ArR7jju+83c3AXcZEsohQJoGgegZT/JrcsXng80ewQJJNYpRtK+VZNcvePWYhzRQe6zg3IFK/Bc3
8Q5sEY1KYcC3H3lGcaKNls4W+PSWLoYVD9bnBGa1tCCr/2dgptgWtPLdR5FbA7ybJGHWJtsMn08N
FxhdWmnaKhZCbLmWxWEpZ3Y7cqn/b3NRctM6FCK3TDtJi/08XLWJNzZBq9Gpd4b9I4sCkT6Jim0D
pGCZpcipPNTUwXxbGT+GfM/WqW9Vv14WjEHYZJcYdT4h0AgPEeQ1mfxitqvmknSc1304bQ0T4Ny8
M6NNYnRQmE2h9asTBCjlsEzQJUhXn0kGKdl612A14rLChQ93zrA6MLpze0e2ZIdFkxARWshOgRsy
BJSuSNcsbv3gEo492PhhNmeuY7Nz/fSEASAi7FqDLgpmx3RbXDBK3JG1/fM3UrQ+V/eEOYBgpk1l
bi8+OQIUUP/pHEGoKap2XznbtRLjCu1VXsu6PCEGqxM44+B+vu+3RRHqJ9oity4wF6VP0nk9bvL0
AFZGd9MdpnRdp70LuCxmCy3d1EgUNkpEDclds2scGRmzBHogyBplt+678ONJF9NRJoIqQiv0FWqC
NMFFX1SvWMAMMvJtyPgd11DCZo3kMlwKv3y260ABEChcvJNDUPFccFxFHRSGvwt9D5R8Sr61WtJj
eQF+wRYMlRFKsEY5+1kjDnVkAuDPHjOstOHSUPGZ4GgerQSoeQr8XxsVoMIJvcfJ/LXajzGdcDn1
jvHJctG0KbXAF1WGz8KJHtlyYjthYCryBsU50YMLFGOfwDU91We3jYZUXG5xMAifXygI9fejgS6h
KqCjsnF4XLsgSxq/X4bioniY5awcWffHOcAHyvRASYglT2jO/Vg4AiVljL4bEaoWQXf0M8a5tcuw
AICvZGypkvWZEguevny1Bx3CG5XgNF1Z7aEGEidIgqA9fk2K2pRSHW0O0+AK7O9w2PqQty2ZQWfN
reNIn4m9VQrT05p6lXPS0NE7S+OWovp9syeZ6tIr6J1bcw/BqcTcSGA+gNG/VpGl+qyZTL3EpXtB
hMcQgKJROX8IHHpj5xHNI1ojtCND01t0K7R67Icbe2KZ220y3xI2aDtTsCUrtAe3G3yv8WBHyEEO
ZmDneT4ZNJKz7j9e/AABT8wh9DAjDLc4geaKUnFaXzsh7xhvFs7MeLwdc4ZPxIMcOGV1pPD8ZsIg
evwp45StguToU62U/QGUCGDJxlo+BJxQEjXRLL1w56eI6OhJ7+YGYBlCcwfOouj46ujn4YcbXrMM
XtLncr8uIvw1pxzL/OovWG16oJaK9TV/bs/MJ0E+DxNNiGM2rGw+gGothcHvgZfHAVO91D10+RP1
K+/jHVCurm5ElO1PPhzpQFS1ijPQhzc/qM1uxffkTZOKtjgJ24gcNJstTPmkiVqTj2w25gZ+Das6
sfzFdpXiOofXslBaHoX1dCG6Itt69j+9Q4xaqfQTEEIE7nrgxT0KVVlRhEaEVQB4lt0gY74rQmR7
rNkabQjSkLao5wQ7lUYfjaYmRE66P0fzoTWkIYFvHjdjPTYJG76OhtkGkXKUjlxoGjMp9WJXi2qz
YlVvIk8h5al8wwKzzkOsKcbMw3iDU5N9OcDbXtMd+8qEZt8IUSEPPN9rf4/9RL7+kZLOiHp1jiQE
nVYqehfL9vYN/dnqOA/qKwv1PWaJkNu+AjWfFsfQSZ42AaV12TL1O1BQFk8CtADqicTNAF/8IbyT
k6XkYN6sKNqeJ+f6N9xH9sWhiecMs/C1LvosraZlEciVRJ4m3yGmpOzOPBOG7w0STGsr5a8lL3ee
X+YgnIGhj3TNXPjHZggpD+IFerViVJuH/yp7CAvETtYUkps6dsFIH7HmNR389EmYRlqYKI4yz1tN
br1yBShF+8N2JgYzG2epGdozjw+1knRlZTjvKHncYn5ssvlMn2/WxUgvJ1Neu8IqbZ36cj5uS3MQ
c9N9m96UkEMnUIxJqSW08Llz8aZm8RocJbMHjmUl4puQs4ZnuekcaIgJe04UiC8agkaZa6Bwm6xm
TXxvH9KV+EDpqy6WQvc7ZIsUQYXzJMXrBEnQkrNjiv/4X4f4rMytb5GqU8IDF+P6+FLEM2ExZJOL
LfkfBadgp4oYedFnMHMWurAWcpiHug4DDBf2hePUJhxq7hWh+yhotXklIlIA/Ipp3uamKMMA1IF1
fZXkaeWogMf9U9LtbGRZH+oI3dzNaBc6+MN5jamlhvmLRX/qk4WW9Bbfl64cDhAFDebJUtKu1KCP
4tsuRPN+7767X8kdrQMi6NoVoeKDU4GpvbQG14oypYBmEBqkUmuVqHWuoqaUqbiLe1XA2Pojsk2P
/ISQipbLXSwqnNxI9Plsj1Ttl+XerBK2fKfxpKusWSTvuVnEzLsCzZYXNZ/Psan+2EdXBg/D1BXF
Y/S9brYgbqkbOPwmhDui8VFWwd9/TvCTvng77lCvz6ys4FNtUzE0Fc+qxmrQmyAUs68yfj9swI28
9467CJJyCt5tFmuNxZI+Lh0ChAkNFQ0sD29j2CRlWApPRzG19AhYWgzprsfIG1eetYk3hRoUNKup
H1Ch2WvgravbmTVnylaxIMtg2OSZhsbTxEtAKTkf2a27JbHtcjpL6UgzVjIAn9gb91FwdFpor/Y3
y574lSqJ6KPeudxAHab/o9bR3gOe7Kjcc7hhXF7+Fc6gOPmF61xUHWfRT+BanUJYCOgXSTlciD9L
ZMmxEKtYNOhhzknqTPEkApG2/b3MQS5AI8TMuavj//PhGdDFoAhGAV6y3tGiWzsFQfUyBV8l2P5w
ocdZ3aw8gnmNfA6crH7BU9kIcmriuybVNscig8b1fdg3/heIfOyya2IwoZcK6xB7Cr4/+8H0W+jT
f0jINfZFR1God1VJQKcsAbIXEgOxly40X8aKfIkNotQM/C5U+YOxn5h6k9tcNNylCyTyUdj8jIit
5/zHrahtnkjCyYglzejTAZkxdI1jaNFN/uJtLdJ39Z2xOEMz56k8oizkoISVdpjH9UNyIcBvV+bB
ftUP0UPOc2unlJLV5NiLzRZOJAzH53MBknxI9Ib4zUGA1CAQh95PdO856VssMZaiaIuwIf0VNfmZ
/3RLryZBuU+SsHywUt/UExNunXSHOKqSPvcpWxBb+XvCDphSbVuKRd/3xStIjVdoqtFo5Oxp4NRx
QQh/Fw8mObly1vqf/xIG99xT1Mat1Hnf4wQ3jt8JTTG+QZs2g9qLefU74KXmPnEAQxj3Tf364Ey0
ahZ+6d2fkV06VPhK5nz8BCAhR6cXwfnTaBVt1q9LfvTjbgTR3HGO1CO0Hu0mIhdOymMfOvcCCJ2Y
RvEDyE873NoyKmFws2JeQU7dv/5EgDaGZwAdlZfa7emHZTqGPq9MdbLfimKPAEb0s0B26RxVUqV/
Af8dY+KwMdsRU4aJHmyUt3SmAAruvDntV56ZoqVn5Kqo4fuEn51NCE5MTWdBRXaHM1NtuTd+IzKO
GU4Po89oHNjcRxGe0TVy0KHh8xNCMoA/wkzprcoeizAXEkg7HQXrbXoIWaDELyBjjqODjN2WsXs2
4H4PGqpg/xlNviB0XEKRbGS6QWPMYJpzV88uiH6U+rfhYj1FhxQZ66bCfFCf62WHeQuVXakrGPkf
hNGS5W75M8KFnmVDoQwzV8JMTc15Wq2wHtjcRBhA/R7fobHGW5183ox09DPTW3aprqCz4CEOzKo/
LLQPJFVcmKzRwA+zPcb5kxosZheY9uxcAsk9zaCSiG7aiJG1wiZKkxfIeAzPT7ohfp2Ezv+0yN09
5kCsuqaGn4+q61SlerozRxPiM4mW8R5Un+BqcObU5N/bZD0sKWEgnqPvL5Vnmow74EjEmfgenolp
bz/hs8KY396EzNoml1cYfwt0w0MQ+Btmkjf9Hz2h4rdWf/VWEJwmH5z9WBXDJ2q8niXows9YfWQ2
7WMoOq8Y/BpsbcBaQZS4C9grRsv0wp2AIlr5RxYJ+FYqK0YJSU5a0ldCDWg9NG+aVBY6HuZFiZqT
kCuPUyj7SshfiudFju7Y3AJH3X/fde1uYqcteNMDCXYU34WdDMMBmfLDn/1iWpS63YbVWepY/YGe
oMiXJX+G5BddD/2Y//VzkYH0mQ/ipdH6JCDgMdnMrVRF8354jEP54r2X7bL0+P/d6f8ETRIa3m/M
aFAAmNpixsC6cOx5Jz4HmG4PR7YERoS76lQZ2oXYwAxT7D/n36kgYekLNJzWbsgKZVi2PyXF0gxT
ZA6anHPIOPg/ZOFVu5GKDLpOmJyyOAY75EE/0G5KOx/KcnvU/JmJp9jSfpI0T7RUncfnRznLl6ul
/gAkOVe9EBfwtuN0LDUiZhWDujIDVmitMy9PVcu2hhkyxmImcZB4Mi12UhXxHTLeGzVjx2OzHEX9
RWZSU81ht9z4wF4GAlS9uqk7OvDcke5hB4s6BnebA6hmeZ/CukEPeAWbH59iR/X/AvC2U1tXliRt
vr1VzrJ34TupElwag1jIFdldLN6I6zDnUVQMIMHCsnfaXVz8jH0mfDvBH+Y7eLUPn36mKm9Dj/Yd
Rp/o4YJ6iw44aXDZEjEgclor3Oge2I2ehbGQ/CP7HvPN3YdGToN9ESqVc4Uds+HNk/dNnIo4HUY0
vAbI86HEPNkG0p4qKKS0S9372N9wq83PG0XpgiTaMI31T8lMBcNhvmb9ohpGJh5AmpHv+YOlSPok
wLtOiE+mPzCbLS2LwehcBSfub4G9qUj6cM2Dwj+iuH0r52kLpAkltqrWzuC+M8qRbqdxlXk8atu5
hDEOh7+zOKy+4Nn/O/vrEa8STt9R0WeAVXgLvIIFJKWjG9sxPfgIrADf9CyJgz4Z+nvhIY8wYHII
G16UwYiEP5tTzZaruD76/CyL4h55ZiVDKbFxRCYo9rXKXhiFykHswbDr1yjdY0ABPQkW7D0A2+gf
ujInNyGGoayUGMceS+SYLUV8hgY1Jt983OnImoHxc7NPcQs11eogeDf6E+HNUcFCKYT9IQVAM4vm
Gf6WF542nV9DZCv4+F/QWSPeo0fMbYYwDM/NGRSj7YeieGslE9i1qc8eiHIkvWIRDEsvZjqoQSac
w8B68hTjjPzG05X6lhC7d2Nw2JaImw+RE6C5uF8yMdVsbXcXWUmHG/TZH3igB570dJPTRI0LEZU9
TE5ZE/QdgkgRvVlX6vitVmDXKwwz26EQWVIEOUYwDIkmE7iNpUJ0bwoz0B/GedEpb1r4KMsgYu5h
7Iz1LD0I+Hbr1a3q6aCUQugao0Q9fSoxFUYjf/OhioCHsEmxRCn/UbgZNLqRenYkamAU8KzQPCzq
Bdsyl9kRw045vHsgbZN5q+i4FoFlXQHcRe1YeVeBPnJuvat0LP9HTOPwamCZusSvKkSeR/hxRQEv
IYZvivGtr3W34ubk90JE/ZmgvNpECucV0+vmPTBNBz151wCUPds9lYmIzC/A5Ls6ftB7+dwvnOOX
tNiUdOUiBNHklPYJrYkkRw/+RPGMR7QNDGVYIJ36y0CdZzv1WfBK46Rouu9vSpylgNZHHNdO74lV
+2AePpcHzhKU+03l6gfpFXn1jYq0H5P07hNPn/0AsBjQcyQDhR/sm6VmSsKzeAKpA7d2wLnuHQ9q
P+NXYQhMDTm0fN075xjj/WSVFCf+4wpR/xyBR+k2R270OvsokplSEBqzLJp5Ivi1hfbY4HwJiIGx
ISAja/KUsLpePV37Jd5Up6/9AtQn1ZG/7aiC198JmF4mCZYDL+VogApiAF9Fe2Kx/5MU6hHaCuO0
odHKtQ8dici366WD/+5U0NPwjnhxf3Kf7XisdeHb2rbPE3ED2kJI43j3TuvK0BKfjQGhPT9OM1ad
LZVxvLrqrIRAB5HwzHxp3erqJiK7U+H/KP/OeAk8uRC/Zvt1Z9uPVv91A6mlPbh2Mtdi8UlE/Rx0
HdGA7ec2XTAju6j14Y4UEKjbAvjAoBmBvyNzgXdR0NK33aYHcVIoWWVy/Eb7GjdnrpezPjYS3p+h
AQtQMKuxsCBkZUdY1nrWWBhb7WCRI8LM4vFhYr6lwk8z40la/CV7/a7ky1EJbl2yqMiGsXGJglQL
X+7Y/ILAjXin/hJFG80sxBF6qfKH2mSG5QUCokXBGl/Iw7Hk207m5JY3EHSeUZ4rfRP9RAOMLz1z
48ZACsqPPiLU1wXnToMbeX+So/uBxwWwiO0KNILgFxvabOII4oHlSF7YuNiG+l5Pnb0nDRmJQ7h4
3d/xeHZCIUCwh1bRZDREeGvvHpr9/o94GbEoAHVHxMf9SYMTTBLnSDXWdMYgUJI4qWpSDVsk+nOj
QlSbHe80T1Ct3dA7+WMB34W+AXvxn3At0KimqSmkmR/e+eHQSvBxNo77wu1JnpbkdppSrhP0AWte
R8pnGlrqQkk6yz+Ei+OluxbCtbWH386KNokVetuzBv+1S86CFjbI5CqRBrok1FanJLAs5/XQZpNQ
Sa2QySqjuTKH75tuIyaguA==
`protect end_protected
