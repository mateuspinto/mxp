XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��HLM}|���ȿE8h�
���C�U�ٌE
;G<COU^�C��'��.xH�\�8^��9��Qb�8eAJ��@J3�'�U�
��1i\�pկ�oe�x�}u�l��-�q^�Y��l/�;_-G�%�=�I
�]�K����h�g ��B�9�^�E�̘u��{Gw�V,G�B�F��C��8ꃩ/��Q���Dt�����]�8'6�����i}C�̢Vn�'h �,�Gіt{�H���������-Y��`,5X�z�i[Ćr�,�f��M�CJTh9�-�Aޢ����Y�^+|`�{2�Lxg�GF�7�-�WM�h��+�If�@L�&@�8p�u����}��s���dr�U0����r��p���qi���Q��<�&r��MO8�@�awn���l1��7}Db+f��<�/���s9��Yl�\�X�۵���/0`CJ9ov�t��^B�(8�u�M��qB	�׋�3���"��:l~nDLu��`�ʠP�̤b�d���лL���4"������u�!��(`� ħ#|W2�H�N;��U����%�.����8�v�I�`OI�@+)��i1��:^�����k0L\z���%H$��W�2��F5Z7��I�(u'���̍�vI�䀠ʒ`x�DWj�b �1���;Y�كJ�M�zģ?i/��;[��N��^g׮ G�2�	0nW��W�Q!{x;��zm/;�;L�[B*��
��:A���.@Rb�@���N��t0�ȥ�W'�hUc�lDc�XlxVHYEB     400     230�H�iUT��`2����Vf�%*��6��8.�[��v�x�I}��5��ݍ؁@�z������g�����<$�s��|���Π&�6ctXYHO�m�����|���"��I��|��KK0-�� �j��]����wR�I��P�(Ҽ�ȿ��?���]_����E��MTN↎�m4���U��*��XB~ų�L�+t*ҙ���2q��6X�׸C��5��Zw
mwqc�1��� �-�x+#0�?~"��8�$~�p��gH�X������K�9a��>�v�ڤ�)�[�ʯT�"��je젓൭a��|NH�r"���W�zlr�I>W�`��8L��$j��������1��y/�+Qr��^ G����`0 N�Ag+ՙ�\mz���E���R�ό[�l4�-��a����[��f�5M��ͶT�s�����O�W@���*���-Y���y����&����k�y���2��$V��M�=�g����d"Z���"�T>�;{�o ]�UQ7���^���	�٣q�U��6�z�&���8w�x�_3�XlxVHYEB     400     1f0����B��R�}�������y�z��A/~�\�̏�u�	�&�:�b����P�j<e���8*��އ�~�����|�(�"�iK'ƾ�	L���tɣ������N�8��f�`X���!���Y��=3�݀��H�1�`���M �E�R�f��S�@啠&'E��y��\�`�`�(C��6J��\����ʼ�f����������q�Ƿ�`!���Y��̿�p# \����C�K��/�;Nҝ��������p��7X�t>��H�8����md�f���v�O�Ƚ����׌p�iE9�j��_��|�|�a4RC�5z�0��k�_d�i��7l��Y�N[(�x2%�<4f�5�ڕ���%�������;"R���KU<���j��j�6�E�j��m@�A�O��n�"�o���έ`6Ǔ!�E�A���;3��C��ju�6u�(�ۿR5 �eM�������C3
���W���@XlxVHYEB     400     1b0�% ]�q��i�o�!m����I-�~�٭�fV׼Ȟ�GJ���W��|j+q��I#��귞����|B��t�,7����j�_�]��,.
���jg��qA�~'�-��^��Ę^^H��)�Q�[���ArEB��������T6��=?����z��\<s��.���n����k���Y�r\�o�&��ۅ�vW��d�:�Pt-����hp�ڨ�S$X�F!����>�[��8��Ju2K���A��`�J����oַ�Ø�,UiU:����Dm�n8AZC���˷kI)��h�'�9V`�H6ǸusG��o:���2��>ao�{w�lx@���]qj�}�T�`�[�xp�k)��^����ڹ���P�2M:�S�)3�en��C�V+)I{��\"��U�GV욒���D>|A�{hɠ��|XlxVHYEB     186      b0;�))Xid��+�U_�
1`�8A(�M*Ѯ$��!�z@	��L�J�`p Q�����T<tA �b7��6���3��/����<��Ҿ8Gگ�����p["��ux1ͬ���2+Y�P}6fP�n�ʈ��M�1��ַ��Q�:���e�{�N�:���RȂ��R���%&�27ry�A��%e4