XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����V��>s� ��{��ѡ��u�p[�EP-�:U)�)��w��=��3`����t�����%�+=ߟ�9ls��R�ܟՑ>{��nL�la������NQJQ�D�`U��6#���2BM7�tU�aS�]$8�:�E4��]�t��2��4"����n9j���*���%�co�#��3���<�w!�$}��s���p����s�T��6�I5-Z�g�L�m��1�
�&/�iϥ��H{�,��M	�H�z��h����OR��V���T�j{��q4�opf%T����u�܎�e�̈́��O����5���I�a<������:��h��1^5G9�r�"%�^s)�� n3��1U@0�n�Ǆ��E2�L8xI�2��H�2@�49�0��NW���k�\�V82)!����}�9��c�A?7q@DЇ���[{c�g�,�U-���/o�d��d��_�O$H{ј�ڀ��t�wn�)v}XхB���"�L����2\���ٮ�
�ؘĶ�v�����m�w����ܸO%J��+��#��:n'��j9�}�9h����k&���U/��ٳ9Vr˾wH2Edm�M�&���$o˼jd��]�ϖ�(����lņVlA�Tpz�u��0V�x/��µ�HR�l���e��x?b"2���"�*�u�R	aŏ��'�{T��n�.D��砟GO�۵Qڿ\P��M��w�D�#�P`x05	��p��D�07}4@�//�=����pB�ñ/5Q���>}���XlxVHYEB     400     1e0��qB�\�M�nYҒ���D�m�{� �U(Xh��7㐳%����`` �4��cV>b�AI��ͻR%@&�P/6ɀG�Ā����"�L�-���"��.�Vi҅��=��B�7����`"/dK�qFF"ϙ_����7���N/&��+!,3���.���宝������c�@;�C�8=}6�J���M�Ϙ���u�z7�o�;&�4�O�S(��b\����̧�`m�)��s_V	��SD��{�z� ������-�c��z����Hxq)�a�;��HC[S����̞�V˓)�^�w��
���������K�Be{�c4B��;��!�h��C�'e)}'-/��<~W�Y�߀�>}�$��0Xa�P��"F�O@(A�)��6�i�䓏�K0�R6�u��5��j��	��5�^���FVQ����pA�(�MP���=��&˂�������}�a��V���ŷ����`XlxVHYEB     400     140&PR���Ή
&3\��+A8��B��%]�X�b�:�6ja.;*�a�h/9����V%��X����1���H	>�p�c�����R2�槃m���[k�����i��(�R;du�m#]E�)�h��w�a��y�����% �C@�L>JӰ�\�q=<��s^bj��)Ί���pk:K�~��!��+W�~�Ow��2L��~Z�*�a��9�ԃ�p<X�eaef����P��X�!�?Vݷ��Guqd���4w��]�/���ݣ�c����@�5H$X߯��t��~u�Hml�Ky�P��e��d��3�W$�0���tXlxVHYEB     400     140|�3�\E������	�1��YV5��(Քt�2<~2�D������~}fw���Č.���Z}E��/��s;S�^�E�Yi- �È�R���fNL�21�(�a� nRr�0*��/xj5|���K�_$>�2��T�f?H��J]�p:���*��p况Z�y�*S�?�ֳ���곋#`�Z�Y{��fz�Ӡ�e�-4x��,�W��UUx�pc�)�%�{lܴЊPJo�@T�G� �-�6��;~�U��¶�37�R-8��ߢ�����6w�D��8�T�%���]ıl��\�l܍zi#Da�*�><XlxVHYEB     400     1a0��Zã*��u{��|��'8���0!ݻ�Q7��RP��*��E*`���h|��#)Y(��F��҃1���r�=�cE嬸�Zgs�G���Գ�ˤ�+��6���X+o�q)�>�&���@��&�巪����`�A�����
���0�^�� �=�	�S�K���os�GA}���ȥ�\T�
�O��Xu��Fi��6�n[��:��a���[�DH�^]��0�W��C�Q�/�O ��5����bb���6��R5='��:��\7�ɜ��m['sT��7�5ע������G�s{��Bxݮ�)9�V��ο���R�z��iDL^���q�J���j�{K� RV�(f;�� �/�1��<�f(��h���0�H�ERL�O6te������yz�{"��T/�;c}�XlxVHYEB     400     130z;�s$G�d|��R�})e
h!Y=
#�I��qTe�y\>���!���҆�� �r��������=W�����x�X�t%���d����j�T�� 6
f����!���(]��2���GU��'��o�D<���^�omK3��v���g��䧫~ŞA��&�T�&�F��->�<M�AB�)̥��X��l�Ž�od�PLLj�\�������d7��W�S>�!����S x��tB8�����ځ�Ğ��VI��3@��A��Z��&�uR�؈K@�Fż�U�+c��&Ɂc���d=9?L���8��XlxVHYEB     400     190���̔�H�J]��@T&r��_���u&�gC�3"�5�_��� �T{�K0~$�$͌���na6��m���1ђ��s�l���^��Dz�D>"�I�qnx����=1J�)u�r�r��K���,���Yr���á�������t`%	-)b�azv*\j^��Ә���b�Yy�b�k#{��&ܘ�)KI<D�K��0�����I-�9z�+�N�W˚�μ��zS��a)4ũcΊ����(����L�y>F.M�>�-WE�_���1�T���g!A�
S�~�+���3Y$t<�+I7o�sI����<�ճ/�&���$�,U�~�_RW�p�F�x�� �|`~:���t| ۺ��k�t��d���"�����Q�A�o���̸F �XlxVHYEB     400     160��/����)hP�臲����w��(���0�P�κj�ڳ&1+�%*U?���`|��P��5���:u�������?���u�j`�
��YW[ey=�P�|�ף&��~��:4L?��!1(�s��?X<Bw����j`'��QIF�pc���#���Tf륋$�x�q�߂�x�M2+:����^�{�"U��2��%�+b��k�Rj ��$�q$ �C�*�S��ֳ�4��h���Dܲ�pZC\�B.	%��~�q(��sF�)�uW3�[<s��G&osE������jDi�7Ӌf$n�IR��eqCV�o��M���J�����{�+D����.�[��4��˒|�a�48�XlxVHYEB     400     150B�k�}G�\�f��r�����^ �򄢵����КX��/�Zȑ�6�����$�5�)+�"����6H���[ܲn�i�s����4&���*3TX�P�.��Yc<�P9�R���F2��jf����;z1	;#Aq��6WtҴ	��6H�v�G�����ީ7�̘�����A�^!h>D��P��h͗�C��Z�������C����"����~Lv�&����-���=��:�57�LO���c	���^�\�^�W�"��:�O�0�!�Z����]װ�ß�U��يH��r�ޛ���SB�gM\؈5��>�Q72l��&5�I��XlxVHYEB     400     1b0���U�@��E_7oP�mG��O��Di���G�0v� A<-zzUv^��,��p��|9�\��Q��_���&���`�U^�lo�k������}�x/dʈ^�/(3[Ѱ4�n��������O�[Jjzm���]5��M*Ic�uxF>.J�K��Js�5�(��29�"8䛲+b�R�|p����F�-!����jkɯ"yp�̚30$�ʬ����-��!H�YJX�n�+<[��r���I�	���Z�z���_V��r���^��2�b� T���]���OS�9��k"A@0����X�Q�%gƐ~�k��9R�L
�Yo9��dH��֖�4�y�BÁ A�n(�2�f�I%�Ѝ'���{�Pł�M��U�X;��m'h�����Y_��wT}�	U��g�\�XlxVHYEB     400     1d0&� �8G�
(~ڭ$�p7$�2���
e�vԘVY��8�ф�`	s5i�DCZ�%�]���0�Z�z�TM.��� ��{��EsF�*{ɧ=ZGB9���X#B~�����]�[��韩L�*���p@�hZ"������q���zI�G0�O�B�36�|W��Y5*?fM�8tωl�s��Q��j��W�̨7�״�*0�י*F�^Z�pIq+��0�<�uz��<J�$d��i�Hi]Z�e�6C��s� 6����Ney<j�6!ܵkP�yP��w߽BA��?�	�;L�ò��cR��u��v���E�c��s4T�r �ל��'�	�|zj�e�W��]=���[���aH?t�[PU�<x���R���9�j�&�̼b�2Ql�=^+�L�W����=1N�����.-Hp�@�����Qys�0�+�_Dx[w7GA�e�o�0Hm��7��>M$���.��AtXlxVHYEB     400     160����j�K���ؙ!,��w��,J<�f�BM���"3�'D����?E��}���Y�j�w���0tԎf�7t,8�f�&4���VQ��Զ�?���u�!G_�hF�_f����|�{�Tq8�E7&|]T��ʘ)�2탁������[���OW����;-�tEYPo�L��:)���fͯ)c��
;��?��k��*:�ڇ�ݿ���`♾��7
�a��Dx�bF�i��LFo����ˏ`���qZ>��sS�\��<G �d&��E"��UP6�Q�[ ^���_;86V-CB��`��(q�!�qm��Q-Y�k�X��"��Lv�կڹ��p~����7tca�/�XlxVHYEB     400     130@R6��^{E�L�AU;��U��U���lv����a�]il��[ �hG7�uӥoL�Ә�1$��]�D3m�֍d{�k��k�gm���Iu~�<FH�6���1!H,~��%��
N��y@z��d��c�j�_�pJ������዁�F�����U�4�@v*�د��k"�Rh�'h`>���#J�
�`���ehT�&2��m"��[�<�o8��~��"}=�8�0K!)��5
�T���
�Coq�f���ͦ\�N(Я����m�6���y�m�{��8�=,F�S���XlxVHYEB     400     180��ª��"9�������������9�b8B����9?<��(�����fX�Z PSk@C����x3Kt��x^�[�Q�|k2� �q�����xo�qy�rQz��(��b���A����|�����q��B1I���5�!֭f*�^�)��?�%�I��9L�Hڄ�=I+T�!m&O	�cd#gK���r=���C/��Pn?a<�f4�τsFm��`���0&P�g�7�kn��"�d�����?yDt���n�[�r�JU���n����Qo�$l��3��8E�Ֆ�k.DE�)���yH�u_���̈́�avjS��v�z�)Ǯp" ������Ә�]])�}�K!Kѐ�]�>XlxVHYEB     400     150x0p&Ȏ��!.-�t�Y�����B�㙁���*"q��b���%�~y�9��ƿ4������FT(ʰ+;F �&ݴ�xbt"1�����'�n�qD��S]]Ӵ�O��	����A؃9re��x�LRof=��ؠ��Ǽ�?P��ě_ KȐ8�����L�����/���je�	<,���ƹ������7�-����c�����(Z�D�K	���A�|�8i�4�;I���6)�����ygD�����2��n���O%��HRB^�����J����kƼ����1�a�0��??5��mױ�-7�卬MvXlxVHYEB     400     120p��[�dA���(��
bo��De��qŷQ@!�h�]����.�S��K�)?0�"b���>��t�N�x��%� ݂��п������^���j��)�\��OE�ѵ	�L�?���]�Ӷ֢'���&��s�|!&�餞�����R�@�b}߉}FZ���]/�@�>P긽ҕ7>|����u�S�"�x��(�`[(�E��<�'uY��w�T�s?���_�6ńۖ�)1β���X<tY����O֟$�<��$��t.j�.�'덓��l�^W��.m�%�'XlxVHYEB     400     100����̸����?�*����yL����4
�p:�����J�s~4\���U��%�4���&��� �n?[��"FN���*bl���Bh�eYkf�P���� �S�`�S���W�W�Z�Q���Zӟ�3���{q�4��Rf���ju&��L�a9�]����(�3����x�fX�8ş"�t�q[���q8�����p�>Ff���(�[�,9�q(��_?��u]k�v(yyS�T:�����bXlxVHYEB     400     1a0���dh�aǎ�gz��'ǵ��'����|�Y�	�>�gH?�݋�j<�I��Ry�U#���>�  �w�9�D\��:�C_�ښ���G��b����`Pc�	)̉���H��n�CJ�V`��Y'<ni��kN+��+dl�A���/jn������t�f�����S���7
[yz�|�f���)����3�xl1NSI���M ���ٔ��q���_���'��%)��v����a擷�x�ē�>;|�������4���2�!�� �+Ǟ���i�$W_������p�)��{u�n�	��xr����V�w��̊5��Z��J5�_��	A)Y��؍�>1��_���GS��9�3��$K� ŕ�!T(J@�.o�K?�S�W��ױ �>�~%�
zYؓ�������[�ͪ��XlxVHYEB      27      30}��Ѫr����!F^�iU����n� �`K�;�*H��r�V㽭