`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9312)
`protect data_block
0USWSUGxovGsyBJteYpEocBaTuqHqJcy1VH3NR59Ys7iRy4WfzJwTo7aqwNOOF7eGddiQ8fOdJIi
tA+QzbBlxy5KvYB0YbVBHOKFqm2bwBZ9xfngqyYW5Z4kE8vnT5FtUilTuAqUvn6be5iTfInRCWGn
NHwJ/v0KZNQ64zJLheiZJoL7GvUJH6seWoPzHmhFoV24sOnyFEkdAWVB7robfokoV6+VCk5591Nd
fVKGaq9J62/6toi/4BvMfLYXorFiv7s6jza0kp+dh8hDkBfHnyk0gIhi7uI7NMknTnP33/Aq61V2
i5cxN+g5AaCz9KpOegPRr+vrOwA92mhNs49wxhzL726m+fqPh7HUo7EUHBflSVymie0zGe7kOssU
Fp4DpgVxmrUa+4Ft6z8WcoH7uV38DqwXi1n9n5VRGR4eKmDUiwUt9dkuAjwDZyri/JSpVF5YdI8/
U8H2W6zELZ++H5MapwqOE2yJ2UiXrQ/leCnH6P0yX22h2pg4zFm2Kh8+WPevqbSI56mw1Yp+mSZz
gFRpyIbkQie1tJJ1Eqqber9PR+IoML968eEFwoCjZ9gpPlvMafx6c397L53IbPZ9elHSr8xxw0pZ
bcDglvfDgghcTftwYttiP3L4PblHqgrkwy6V6mvnXhsOEDeS8N2pzVrYpKBx4/zO73zT0llQXf9k
a1UX4QabgKhOP6sLa2EKU6vk2pn3afJiECiKPaENoi8KQ8aq9iccp0wFxj5AiLwrg63jUXh6ohZf
h7p/ebgQoQub0WKw7tyHREGUoJ73q22HTGrqZ7dVXD0gpqZvyxziqWiK68p8S/cA7IRVUTC/ij5l
hN1PwqMixvCj4ao2YQ8lojVMyP8IWpZZSa21TK82wIHWq4H+I4Jmx6eZdnmuyy289v9MlsiM7WQj
T4lJXgggAJstSk5tzXK7D2c2ovzAZuCULz+CU7B7v3Ua6Kav6jD6dBXq/V4nfFcDcWmLrmMAsKmo
7MpjXmbbzODZYJK9ouvHN0HmwcuSzKr7VDqkki441eCno7W8qE1UuMBB2xzN0zZVhi2CrNBjhMq6
BC1FrIAJkZku0AkhxOQrkWoqC7oOm10LI//GxbjUD/4xMxISyWC3R+JiAGro532AopQStyr2eW81
9YAtROZa01xC66GZfr0YlQC7Aos6R0sIYc6529G2LooiLsLgohDPczzVqbLEbUWLCbY9kcw6tnHb
KobZsbALty8TrnI2JfElQzEc9ywVwW/CP0DwvOSy/ys40qPLujB6q+6IFsftLV6X/9+wngj6yTRm
rVA6Nhe/uKSTJ1AmxVjzq89b/g2oN3FCe483uji8ESk3RmIQM7f11D9oI9p3nraoyxeDj6lHDdqO
8+Hr3MEya2rRgUi/EARgfBc7fb8wBTgzqEqSa6Ghk/sTzCW1KNWV6X03MPBgtH/wt+bDTngAf0hv
IcjkPm5wX/pH5ozRvh9t+leo+b4mCYrOAaH0TFDHrPTc4cgEwcNpMAPcrgnGJ7T+lEdN4S5CU/ZE
WYeK6mLGRLE8AyaGzgWLGp3B68Z+K2JUhDAiBA6FFHkZNqdkhh6oX+8qNDvIZENUjWtmcEq+sGvV
chpnGJXjd7Q1znX7jHtuzqaNHB0Ulx4fLZBX0Yoseh9RjmWfLf2NFX1rRqNri/X+5n958YI1DL3A
3QLVlXxUxd7PXFzQDUF/jyQOm8fg85wAoWrn/U6g1pnIMK51WXlEYzQwU1JZlB9UYm8EnH5UpZ2T
z0CWL/Ec/8/YfppXtLZDb3cm5POGi01y7Nr5yoQgDtJluJBpatPh2uKdBQ9Ox/muVEnFjAIrTE4W
IPFNLwDXFKzcT47T9hD9xg1ImumT18ef+4eFmvQQKyCiG5yWIVbBgD9APyJdK11RZi+TmX9WAXe/
vX9X/SLfj2oVeNBcNyoouelk7CMFar86No3hBMDI8rdw3IO4gXABvOk/cOnK3ShOInz1xupp+en0
dhmlekZqAL6b4XnV9PRoU0v6gBTZ/JFSWn0amV0QAGvfrd/KVCCi87ZJXqedHrtpUVTnxvrmMkuX
mGfi91xJOu3JIMfQ/VWXVFOy/r+RtQk6LnkaKBh0lJMTHDt9c5NF5+VlMOwzV/A5PPyCqG8l1H+R
gH9mOAs6JAqw4qCSVlXA05AxsKFJ7qQbYIF8bS8IFn8oluDVPC7lgOFBMTvL8LCT8/UbRrha+Hi2
Iec43zXIIZkj0wKIFgAyRcxBD1JtDojUmASZcz5ipP+RNuRzAGAh1qjf5wBhIQO4xZozMHMvd3P+
1nY/0N2xE0CCJ5DRR/EnNq651uXFM7dsXXFI9pyzaqPyGIWQmz7WZWu4EcqmoE8n8PliP2jq6HZo
4WclsIRp8YNt3JaEpRFeplQP5tPTH/2d7zXiJV0CJ6/av9EoohgNDzdtSSUEFqEBuJw51d5SqnNW
yebSOOG6Msolu9qSapOQh+w1PLlhFqrnIA7r/EnkncJTrSea+Wi8JXELj1sKx4+kO+2EoCgxgEGJ
jwVmkD/9xMCmFlfHQ6QWeCPgA2e4ALKwMQj5/mnaj15+GVMNoFqAKX984dWv71jWV7dhEFxq5v3C
FxSFpk1O+/R2zzrV/OTY47iu5xc7H88CZ/Urs4P0WgBhwZ2oGxbaIbd2/Eq1t6ZS2vQEapO/hspg
SfUPjuGGQliZ/1X1VbPMxU0q8GTufya1r5ZLdAKO3BBmxZxRbpRdGYq1imJ7u3FjWqbcj9YLfq8k
VcMBOwl1Wf+qi/zPtjwizGjhx/iVmLUAXBfpy4fd3h2/F/WHitU5H3c8Q55FowGdI7njiwPVE/PL
twBVAsIX5qqwL7wy6I7RKNDe1iw0h8Vef4yWwIasrZbJeR+shTOLU0iiUVeMlTrXeqvA9Zc5RBA2
YzQe0r1UTXbYfv/P4g24vWz9xu2NXR5rTtTjrEwlYP2yTmYhyXSvxNCzQEXxraZJpeM1H4cY8j4v
FeYSoJPrdr8vqf/G50DMNkhehS+BE7or8v1Qos5kEd5o2HLkNypvLZpP02+QW6du0N/WEC2o+pIj
Hzdm+674QPhndpjnFcI0h8anz9k8Rk+BSXm4JTPb7dpD7H4sZpF5JaP7UoDsHD7GG23cIukzkkQe
Hz7rtBnnEs+OQT3ecrlwzbvyYovEmi03JKuAViSDdjd2Vuk6USh89k5NTPDWIgfFXwFFU+2ubdKW
yBUJYz4FFMhpUCvaGBRFewYYOX23ojsaw0dWaUaKuB0S3zmLIXO6NRiPSid/8hBy28k33KNFCho/
1iTg4GKHDiRSShebpGp6UKvAFT8QzZtad0qfo65P5v5p05AdeJ6fAFbBUmcSMPIx8J6tDOQnoTdD
QzMiPnMt6ZaWX67tTv3/y2z/rkZPlGaLWX1ws3873VucOccsWVwZUAd+9EWSWymFHOxNVZaOROeZ
CmXlLWK0aFNKVowNQY56R5GeRNkVmaP4CSe3z6zEiTsjpwj2liP9uAudu5oH4IC7SZgM43uOQ103
IKbpOIKEkoMY0LfrJ7rF2eJGas722YJGhF1g2nhWfnnZA2RGI2PO/LhQG9Dql4VCtzv+nPFf+3uM
VetjQba06e8PU4PTkGzAOKM/Em+Nca/Awx+9yrBmtcrKi3C2Vfpq/hNx5s0wRIOK9v4nn5Y3GL6g
eoOzzNTcxlBMjKu679xK6oKONoetSIIL84Pw+j/M1H1vdhMge4AUg3qRBimR8E6Ad7EfYirzO5Is
auifA0BO3nQDJOoGIMTiB6Wr5nMUA+H6jBzoyXlA5oxLwMOMJUBAXt9SskaPEeLX3FzFLGUvWYd9
TG/Yd06r8kFc2PvRGLAkoR2QLV1yfh+5OTGXc8XYM9snFbp75eCEOQx5E1l3y/iRMXewnWRg8QPw
2MpBRAr5Ud2hFdNYrniatWurT1qKQrTwJuGHS5hoU8nF+ZFZPQ1PTwZ8m7gMZW57u+LHm3aNS2rk
x/Fb+tjRvTQZAFF6/6IHSVqdf5q72YcxkZGrkblP4+ikZ3Pty3GQwt2RG/v7j8v2pIdMEVGj8lFS
PFtB8wv13L/vGuroILAnFpa+f5iZWeAk7bDTDpQMjoj33VqAEXoovP2Csk8m3y1j9n+dvoBBYZ0u
PdtVXqYcSHWxKXQplR4rVwX16IQZxm2InzQKtl4Z7gJzN7R+a0R4crzyp8yi5f5dNdB/iG67xFqB
C98Jz8z0CaO7ML5xoXn9A/mD36lNuvcha48ysRgIAGePRpAhighw/lVdLbEphOSCkRM8d/XeyyUf
yjRyqUUuMiUu2BeyCSqQQGVnKc90YGEpecayRnXFQDKsMEnbJrl/mf2HaBSyNfw7BAnAyjcpyIEb
WAc05C9JWqx8X7a6Wc5YOIBuSdWC0DJRh7SQdxXKlHdtzRJ/0luj0BKzZ5UpikTzpckmD9JQco8f
bIjf+I0f6V2PnehMpR5vBM0+QJ7dPbRI68HI0HqYk+SjqLQqJLvOTNFf/Y0W5peX6ZO9xYMtPFvx
4JPtDh9HQlCn12O1cmVTRWdSQGE8Umvx/7y7DqV6cwbOPkOcekIfSiblrHEXVtAgN0aSPopP7LJq
vuqvakFQwSXp9Smpc6egerX6p2eOAIAkjpHxKSZGQDf/QKGktayYnHOCXKZzqcCqLwy9vHTxlfs/
Hp+qqqvuJJtnbfsJlsabl1OFd67xkV9vGu3JCcnkPt3DHz9R1FKIT9JM1ew6LQ7znndbZUP8tdqn
XZiUiu5MA1ZTh5v4InqnM+4/DOARZUuSvDL4pUY4cgGxQKQr0XCgtweicoQP1F1IQ/BtYc7kTM47
aAlTbXxV3B/Tl0Col2RxVU6g/tVDan0QHvuLjdOD3zVJ3PPrr2q/KoGhqGyBnap5LDn92eIoBpDj
6XCrQXGWJQEFE/dNFtzXkmUwk5N3OtVrOuIeqgvtipfj0cx+mZ/VKAUr33iNH9uBg4KZUyr5B8yO
MC+33PAnkpPJguxurUHO6kPtOCTeeWWRYju/7hCJZfz1Ir6YXVKl4sGuBSj+JhazVaeqdhFBFBWk
a/zzcIQDjr0Wh9qGyrBE6JGEelZVBLGI5rn7X6Eix180TSoP/QpBtMS96cqncNFIZDsrc0px/Xdl
KfV6bNWmfYfvhgRUIh0cn3d1UqXw/LfyYjOImoi+jcQL890qq0vM0KDRyCorxVJZv1sYPdBgU510
SLuGYVAB1Dhlhtb0aMjtqVdh+Ti3cGcTCK3Xk/pGGIvKaYmszQCU2fLA5PTJJbdJViSQg17WLGUV
jiicjSnatokzEH1iLSBggLAMmj9nKRJzbwq9KpGoeB7+577M1lbyGULaADz1m0KFjSRGu65YitSy
6Rwec0PFQwYjW0iU+2TOEhUIVB60s7Wjd2NcCCaIfYCk7W9ljSrwQImsIqP9FwHQ7s00VjrkNy2C
TtQ+X8aQ07l/d4n9MMnkCLdW43R0g9wuq2ds+zpfh9dGehsytGpYlZkdGE5m/KBEd0S8VC47jmbt
HVP606yz/798Nb7wIwB4i9AyxdAxeu+ihsTuV1MAccCAtvurjwXUQq1Tgnlvd/T+zh7cp/q5yTWV
xSRDd5l71r8sgI8jeFU4toppQoD0OPrP/eo376YXSihbHGf4P+vfdvV8pJXLgbB0T0RcES4IyLuw
x8Ka0djx9Du7/Q0s+0YSqaJtD8PKx3AiDhHdXSpE6jkxlX/JovSwsevboRUnqVeoPwNoPU0g133f
hzy+W7rkjF46/ffk3lp0R0L7bBDkhzy8KVFZoOTuHlysBtbE1Wx0cYN1xjJgDrpMjSmZtyX4KySP
YW+hXM6D9166dBQ57eZy0AurZqqONCknsEYgYum7zFK/70mnnU9C4W8o0C3rqeG1t4HgsnZlAZ6c
inyYsozEN7p6z5B5n4ShCRZ7GcIajrUE17yef/b6Hi7zBHLdswG7vdZVeSPUawYmEl3reaziXA9B
w6RTcwh4c4wcWTCcsdG7Q3d+YmtxfavsFo+7tAD9gNKXCiuG2V/IizV+5cBYqLE/itmYEg8h0peh
2Pk4mZJ2IvEY4AG0yWN4dN5gK/UNIPWn/x3SDxmU3YS6bB7VGWU3AVNCiOenYALHgXYlQlF8v3P7
CEty/SOc4aOSe6uwMlFULoFkcP/mt+5Ria+UJhvLkBd7Lci1TCDxYtIDD2O/hsnwZ6Shs/gan//7
QVvbV3FJOLBQvUUVJQj+udlMkJTm+1E4qFN/0sYDw7L73YWiX200Oiq/M+iXz/zLVqEVrQPLaUnH
uccDWGuYtuvbPj3eAeFI/JOMU76SUqfaUdGjXf/R3W0F9S0uA5UBmcDXvu2T/g86ZuC2zW+mAfb9
d4R6g7gBwNyzmqzxM44TA//zvCU8gEzw3W95r5/vZogSGABI/8rTyoAgJywjU8t+RT7uRlRGRvHD
jgjGBQpITWqiIPUKU1fg7QFqb4QT+7kqInxU/dJs0L+mqbY25BOO8PZrSRK3kJYR0uJ2btUbaTRe
DV6DP9XZmFt9kVlzIwSjKMY6llGODrg45+JKpxoeH86RrFRZS9Vx2BZ6i9iBjWyJ1ByNwlNFQKdg
3oTn1hxDGHdA6oPDN6yQlZguTxFIgFKQlyM5T2DIm/ba1T+yNU4Q03XXN4Sa7JKD9Do1JN3ox5aS
/kV9qQClQ8dY+XjIuWnoG9fPNiqqYWHsfmyA8m27OISwTRTxmFFof59OfjwPquug85o+U6A/0y2E
a2eX3zkUYlrwsKpmxOhziC3ahtgHpp4bBlRg+aQdG7C9YFZ28F6g59+2STeJ/g5P14/OrkX+pad3
+zo2reoxtM/ih+D5D472KDJIqLgzmru8YwCzV1ooYNcU7KUGVgEo9z8LEmRy3BfXYFL9kQrOBtwc
1ayLZ+I/6hlGH8NhaCaCz5uvqECWFqenHuBRWvzKLV45algD5HljQFFj+Z+SAG8HqxNp1f9MCBYR
ReWxPSG3W8xDYu6MSOSb0ynGsZSWxwMzraLRcPilxtFfCT0sSzz+1MbwWF7B0fmdO3H6WBpjHZNr
UYSobCEv6BuhdmR6Hg75oim7Iwu8t60tQWWXINjaVyADXHNL+FbfdoSBHUBBJvokhid2YReWBxln
35r6Cc4igmESE+3sdumN1kARGwnpS33kDyvCm7dRbSjvCGJQIch9M0chXxDZDYypl2+1Qwwy9SV2
Cl+50H12/0QdDNovJSPsqrxEagrEecCqT3+rHIDrn9ETnbI/WPtykfv1s4JyHZYcCDeV3KnDBf4o
CiLWonfNINw5HvtMkd5aYsz3S1AA/vy9mVk6vEL4wcBNsHfo9bEqNm5cmAYhbyZ3/2qgGsKGAVYs
q+cvOox6H9rqCxbyqKM1hzFuAlIpvIcK9Tf5dM+Tw5uFU8bXHv9yj2Y/0r8Dxi25tS+av+5JmbCP
m5cKpfasLZlt+iEe56xw+FHRXxAlHNOO85Nbf64BP3b746ogTi9OeTPD7mi0lPT0s0/sLzIe3Rc2
DM7nwyEBZe/0lfnx8bp+DmAuTmpnBsqfzDW9mLZiaOz4EK1CP+uxUOVw+L5961nPZ1Fjd/C1Aq9N
PvQPsna2VQZJb6aasTzFs9dg8slnZ67hR3o8wJ3IWBE4ciBDwkXKLFVMyGMgRmFPtFQP/KdPQO/a
EjtpcyxUhPpV5joO2CWgzuAkQuT12sthnu5h9KYR/naoVxd76MCUe31AluxKq42NdNunnoqfvECd
fXcWIdWbYt2k1KQKp7ro3xbQAvaceKr2u6EM6RF/CEKc+EoYQxU7eoDpRFJRHEX3Xi0WyUJJIsK7
TWKw4i+RJtGW9/KMNNGW5XDnGiK2+roypoM8hb/7VQcbD2EbcCSN/MqQydpJL2kQ1SYw9xDrXyD7
cRzw2m63rqusKxNUYQqIulElID0pjG3HLyvV88Rsa/x52w/E7R1fcHOvOBGWGouB7ANqoyGLESPI
8Z9iCH7M7TTpqHdRletYxvECttITH9gMg34kK32nHTZNOs68iyItlzdw3rAesuNUCMR3qp/q2pi5
/+sDpfY+POCDVA6XPbU9UvwIEQ69ITEHVJxXBoENt1aUKU/2Jqxiu/0nZehvJR8lsQYc7jFIOhLi
sI/dz63m8wbv+F3/XXKLjggHLgjYBcB6UKcRbcLi/B/ioy3/f7VHOQsuU2zmT59NTGYAMnarn2zh
mZ1MoFvW98cLxI1C53V31f9Jc4YhJOtkVhDcqLehP/CjL5ivMWW7/Ddi1AaKSi1TzdtJmpZtOqKZ
Qz6yZAi4vJwFnTZ2FYnbn32lyRIMPc0sSAgwznCGxQR++PLd/NdSfsAOAcA4ymchpaUV9390qEhT
TsmKgxzvm2u+TYzBtTTco5kXmNMAZfPtRz8TyiPcLPW4YS71tS9lO5cv/9WemHMCJF43zJ1SFQWP
31nU3FZldTOvRGIyIhJ2WxtMG0lcKlSnIssLcL5E/arPOSGgl1FyIAiDoAmH7opE9f11mt23Iyvx
ply5+6Osay8kiGzigL6S+YGiYxqnYa7/xcgaC1KQAUEvub1Mb7hOnygrDNsBqZ2aWX961J2mwE7h
5LVLQaanaJA0sKN4emBtl06MS3DODOJ0ZkTo9HWpGRbY0NywTzg7Rw/z21UXN/df52hxB1Y8HdH4
3La2m/c+EDvZCigcYWxSDS23WhrtgznFf/IewcagUCnk02ql3kXUjosQdnVa8wD8TSfnE1/zMw8i
dNV6W9VTSGsa5GF1kIxHNU0B3nBH/uJajyLF1GDNMxKXr9DE/kfUhWz9YvowAWN/kwwHzVe8yQeY
o92lw9mzye1qGxjoSCPbA7NJwPxorCizpkkUQPMSnRsZ6R21hH8eiBzn3A3i8lXjyYQhMblctJ/Y
Es2PG9fxi44n0ImzM133WjKmqK7nw4U0Xj34EMmc+iFHJLgh18MbMIySQ8VAOe8UGItLt5HJWsVf
Bone2cWi42bIi/Yq3QB7+mN4a18jvJ/wCl59qLAQrMkrHFcTtVlHegRGh+ZMhniOfrR8S0nvoCws
GOSPecYR4oEqkCBWGTbwY/90c3ER+zFiay8sooMIVfpXSh0VEYk7n85325eyCxDjTvkcIq7cTDiH
+1A7Cp3Xw7Bie12np14k4FvcphQK6twxbnpT0mgXcTjzVHB36IssfgoHIDs8xfUHfjKKxfjGCRHU
gxWMDOApDxBKOQxv1IaTYdDS30n9tBskuvLUAP6ncef79+Zj6NCgG/9kjR3WzmIprsg9cCqkmCuh
rmOykDzCOmE3iIl0XvASoCOt7DZ7w+2yjQVKvl/9x12VwKZ0+zyFJrh1/ihtS6JJmnm+CfTAEYjd
yProT3u6IISxfPaibvVqi4tTSHqiC7dYIPrAULL/hyf9q1NCsQtCj9jbzT7cOBLdusJr9ky5Koj8
zfpe+XRt+Z7hPhQ2n0AF2kUQMjb0G87HGcsWHZ6mhEY85e99pxQQ9FT7ub+HW4jPu1WeLj2DaxIL
JapMOHmF3Ic9Tfghnrr9PP21N8sXKVIswJ9y/t1490PNoYt80Q/7f8CqIXDyEzH79sTekXMPPqBp
WwCjbzB8d9zplig9UPCJesWVZ0yH+Jvp0KZyk8iUK3VWzjiUnz2VjKrjkjUj3DU6goJGdxu3cTPK
qzPxkxGLblWmRYVjDPy8Ec7VS69yYHNcKXmp6zmQPhSk2e7E9vFQBkn1F6MBOZ7tx5qDItzYoqfd
RhZA6G+wEXbQcIalk8Z9jF4RFPn2rQqtf+9kjhLRvesJftoLy99iIQx4IS6I2GwdTUzbP14qaOT5
wQ9b9X8kFaQqnUgEUGEy/1NsetviaxReAee6CJWf6lQ0Dfvv+bpjGdHQ67ol89/5W23BKLnGjXqm
pI8+MaYlQDUaYQaXCJiiMyfFeQxa08hwI8pV6eODbv51ZCBeRWhu2nHbLqA6+fsoi/uwpGE/9YlL
mpP1XyrsyPto/YfeD0ToGm2x6Id1pQUDj4eDX3NPWO7dbZgRPIltoB7g0VGhP2ksdlB2S1fvR5do
JFcSC9NvHRlLDb8vrDJu58glaRr3e61nYcZExcu/HJonjdfd3umovf5lGdEk6suQibJswoUekFRn
LKTs/yinEw/IOlvt7jThI6fl8w7fQLTeX8AXvhM9oV0SIdIzY13U4go3zMPE7s6UMoRecD+koqIe
HHf7w2WMNRnH9JDv3EH/frFnhrQDPczbqKeeHcD39QeJi6wkH6daBgIGbT8y+4FfiZUp1zVwFbVn
+UJuYIj59pTvFFoG8SeX9nAunqdEq0klZ63MGvOAATHzL2H3Lekcduurk+zyfySZ4zU8KL497JFU
zl+f5oB3swptsOi7GcTV10pi0mR7+H2jFsBKiD9hKRtMC1m86e7Ht7y4NIT0s4MF0mvTnuRnFpv9
eDcAagVBrLlVRC1kc0OWwpjoOBKf7h2vsZy2E30NG8AuKS9WAn74G2r+S5KBJivPsPNFlUrlygOU
CKJQqDewzvDp5QQpJgyfryX7ThJooOeKnHiS1dwcj0mWW2/eI2YlQ6lsguUZtu/Hq0cui84+U8JS
gAH0bp8vVbjg59/wuMYxF3EQwy+6PjS0O+z3HEYc0CVCnAKnV0NgAMBI44ID6fdFl+L14AjQvPot
W97ggtkAX05itYbvZVZSD2/OlUZ26a6SwEH6g5y7qQrSku9U7FoHrHElTpMOUxjbwOkqzs/XlTaS
Wici+NxTTO6xa+LjVWURu2sSt0gUwM5NFtv0PHYxJ5pNT/q/BxupzGDyHePV7EYFgEzgD90iAXTc
BlkqTN3mRGmGRQME6V4DiX2GVLg4Aq+GeiMDQtf/iUK9FowwaRDFWOkHE27sd6VKJaKzioiIno4v
2p+jV0yW8TunEeBAfvaR9oCweLLnzyq/3RCnwFEdoshi21wSzuJ9z+xY9qZ6rI2bv45dmuMLYj3R
d8ZPVf/d84Fs8+iWEeX/N9NueMSthdHhCdvVcKldNg5h0WV2/qdgInzhALX+LlHTaQLCAOpQBW9D
L2wRxwv+5OPED3ZMPiQPniqtXEnx7/2Q0QyEymFaM6G1Imz2yJ/I8BwsUmO1g86GHhhzd7OWa/Tn
HJgnkA2BMOINleLM0Q5L68vm56zZFbt4hdGdFsey8KuFJ5ymoEdmhMWtYiRMNaeVEA+PQwfQ5bDn
Mgk3YdU9Fu0wxmOKmZE95eTzJk06+nE5kTRPgJdokE8ImfNDf6IGsWUlpjC2QISrOJ8fEPbML3Zn
DR3yaQY/rmAAwwIB6/CU/jkacR4ccQz1hquPnhDYSiekq/88ghA6iMsXqKuaSR45B7UEa1gyCQZg
ED7H9dav3o5S/LxGKLp+qwhvh4K7YyyO2qcGfUUqIj8WpoICJOlEJj4Wzfx2M5Yzhor7eIHP7AgF
l1zsukthdm7SZcS5QlUpiXectks6ojFTcbo64Lig7cy0vKYKJM7bFqj+ThiSO1eGble0twOVHDoI
Ztycf+q413KH3u8m0P+8QIv6sFqqefej1Nw52rs1DdiG1lsEEIi/efJHotg7Z9OK8RUgVa5Xj6uy
vbhjBX1FeebZpJpC5gRjLdJ/MmpKVB1KvZFew5vfa/wji28ta6GPSz52KIcarzwDqdm8LZpCh1KM
pPj3kWbEoeqVHPsffZDmURXeNP6plrQejBSVMOXYi7ZwwB/JxDcK3S0/ch/IhBJw1AlXOqNKxDpE
hlFDeg0D04XUPz8gTvcsv0oHjpy+PtllRxeN4nse9FdJhZRkZy5xv/cUXHSm21JxW0oolqmuGcs4
2cRpcn/PI/zruc0MapWuz3lwUwbkJRDlx7FOXPlKVbKdjzS4KzyeytBs6yYleVru/sqAbk3qOXT1
7BjCfaYdR0z8hPagrN/4DfLvI8ZWOfdavJ7mv7JH/8ujIpkJlWKqJ8hU8P3isHPoe3cayRjCo5ti
ihdKvyyaJOdJ1BA1xYcFCLJ5129nxGWjKp+/J0sHVbUsHbRFPvloMdTQnYNO5tySlsUKRbCj7L+h
GVG0MLVFWE48tD3VNKq4GNlNWX6PM4yScT+AVUWQa0Kflz9dzcfDrHZ5rcbOAL6YgmypKfMXt5ns
Bp0WyygzJFO5hHBpZuJVD7u7eyUfIb+aq9kArEeRR2AIcLfi06LA+ptfRCxpe/3LfTKR5c3bv/uJ
rG2VrJ6hp6AZjKuaYI9S96wMGHdq0Nta8qjGRDR1c5TA82n4Cb43/DxLs21BW8Q+CZNzawoW6smv
PzPQeqiqCyx0gd7rZeuonHhLvZ/jlPfXuAxC00oDMTx43qAS4HAeRIFWZjt8h8I5HX+ArhjUwXu4
Zq0GdBrmCCNd5v9T4/SZ7qAQ2wFaDJOHwboo4X43GzguzHucu6ZoFuZUtw29RwP/sSoNGEu9oRMu
e6c47VnX69yt/WHmqk4v3/EotoTUlEhEBiyFFDL/35RzfIwtixGpV+tP2hAAgyutMLWjbRPOEnZO
q3IyQwmmQEr2OTWpJwnUSj8zbtdo
`protect end_protected
