`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
ss3ZswDUBY0yh18xLHs+sIhuu++XCYgTS06lqqDyDckoK9jtW02IwwoPQd84FdIPXqqRBzHsujra
EC9eks4Pf+GPJTcQIwx17bpVyffueh6LS9or+rktRX4sEQoTkQu3rFbFzs19DhCJD3CO9/3X5/tZ
UFY9HmEZ1Kzdt8SeruqFy5P135EYBrzFtFZ8YgDW3E2V+MrzvM3MRmIyupyFQX+vFsOKogIZFTTn
rHj4udkkVUTXamOBVOIMi+R3DMwyZYUAI6B3OLF2T294GRbYJFYDIsPSGI5erz8z8XLNfqx45Ra1
Vgu6MLlWYrxmpZxWS50QZaR/En2R8F13zi01f704jDHFX/Wyujy0g89AA1m6v/wFEPeHyjjuiUB/
8N1qNR9PxmYhfoHyEMEeaGnKyvHZjJcuvItvYHSeh20AOJV8WwUsgE5ztvDZdoeNzH6CAPP17Ua7
0dcO1UepLMEu8Ffcpz7ftlQg+iz3D+sioBF2ZSwcK5n4BNiZs91/+auIhrmZPNJVX/DseOUoYDEo
DnM2dRk622MfH8up3mT6HIuuW09k3nQ6YROPHxuoF2s2QCQdEu8le0B8YQXAwE6ldqlOv0xZShvK
BeRLbyUrKqqkKVOhSK7oooX5Yfe03ohymiBbBojWWqxcG+a0LG48tZc/fou/upYJm2COMFk9Q/MW
GYNurmurWxUpkSBA067bD/XFW/08aDFNYc+lxw5YgNR/KSvYLfIiohKLoO2Gm/f5yGg8DWjs48Ja
PN7pQooLMC1z3rp3HcEJNc6UhFWhexLWQB3Xvc3Xn3seYQKiy96rzaRExVPbQFRsr0zbwhXFcqvK
m2gR1B9AJQo2rBQSufoKSKMQ6dSeQjr+SkC4nByCrsqYCtN+RRx2HfXosVhaHhfyOI6vlIz9ioW6
u6bO+QIJse2KSs9SL2esfZb/iNLKnqNSs2VaGmFwY06SA12oF7zoc8n5EX8qRRSL7Q+B3PrlBExL
zd0PUQKIAXR3mDe/Qd9cVyqQMeM/6ZVwFxXdM2nV8FNfV//UK1FeCCzzT1z6vMJrAlM0pX50JWAM
YIcD6RYMltJSylpFcG2pNxU9sgnpHGWEX0NWXKh6BMv3THy14v/J1Zey1dOkUx0x8BCwx8n3IDX7
zUCy2EGYq5Oi3/TZGRazcg5s6Hh7u5iyb4rvzdbqkDBGYNVrqqqlEOwR/NgapnOAWucFuDWzd59Y
wH9mwW6TsyZ0ZuCKArsYpHZw5BBFdvoP3a/3tD+tYg313H33nHCHRPKx1JEHx2erWW6FHKqdrwUQ
vLKIoOSJgexgBVJaATHfX7+5hvIo4epPim/IkfRYTKbXCkmONvsjEaGcVF5v8dijeDSZOzNgCRgZ
CVyF8lqy71mUY8tAuC4zyc70OrTdEw9x+Q/5hDItIQOOfyF3HyH3tG+tmxbTfCR6gi76eIr8eruD
8wzYkuU7Sy3J8rwjYGnjXpvXR8npxiESJ3HGJr/ySHj8wpBuCQ==
`protect end_protected
