`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17632)
`protect data_block
0USWSUGxovGsyBJteYpEofLk33WgRZd4r/RSvYrUFPROS7zPz1BMnmh6kdjwjvgF0c2tUZJPEd+b
zFhhxJjbgScPihaNi63cJQVBC+vniYp8fdIPk3CqZRPiLtq8mMN6OaUjYaeZQLflUFAlmsgUXvAu
Iko7IyfKltSQjUMpPfpYpfvBlO9Exmac2OdPogq+WET0s/B2uBwi+T6LjVMqnyY/3GPngvxwwLkU
axzwuz/u1Gm1XlomaDqa4HQX+CbuDZ2uJV6fTomU1zwvzjH8BlLQZNrhvyobzClyc8YyegxjKYbg
INgQJHpmvTFRj7skIZKb6fDz3bILuAFeLUxaBhfCmZUEjEp1xFouyC2nYMKwBFprBK+SbEv7uPSu
aUWlNHaDn4oyTRncKCmYlpfWGodlHmqpH6j1ggKfnqKWgfFXQ/p8SuNVuba8ak9Z5iU6ZJbjOrgl
O5JkxYPuFiE+mMwqst/KgJGQz2pVo1ANeCwJq5VDiXbMJ6LAySKKj91AAGNZFWJrc6edXyMrgA27
w+Dzg+DQ+nbLM/TMS8H1l4KE9ih44S7ZP7+hE6/zSr7ryHKHwn9hZw+KW46IZgR6IYvDqTE3i334
XJLJBlHiY/prhREGss7vBwP4R36XZEK1rFmpYNm8puNzHyrkvSNiGIi5zxCLUSGWe+MCE2vk3uUD
sSsgP/vIs0cgBAXWxUTUJRsw5NsjtkP76URyxwFILvKLAhG+IJDFw/palJgoAaa6fn8eWVYLWPjR
3qgeN/75NPPLFbxh1mx+CbpY4ELHok1ANPaOCL4Dt12y7MUj6/N3/Cg9kUW3vCGJCbRdUywgyehP
YISc4N31GIOsEg9y9bp3tZhg8UznP3RMe/f8gZE/ur0VyGYck9Re2VAEyF/X9LVz2xjeLPnrlNyc
p8inczCPfNcyNuDKSK8Wrm8Np4cJ2W1Ztk4t4wFzPVJbIXnaC5VbOIX81szvJxEPwyv1gvRIq53J
FmngovStPTF5opOjkMl/lABhgsQDZG3tfX7ivGXefW5KettW4+YuKs0Jd56AfIwUfBRtVf5epBn4
LWvDKOCSkrw3l3Xc8kx4vuXfgUxK6DxEVXCP6cgvoaMZrFEp5qmgDm0QFLGq1yeW9+uq/auKqO2r
+bYzqk9At1c4vISyIBmVbWDk0gX1zkrcDVc5tlhVHxUK6Y/UXbkDnXQs0OAfMlwzos4CrVNS2BzU
cMHU5IrU0HUU3yln9NZkQozgE2vrbNhevqaURClRngVZLJjOO8ZetNqZmbyEZWFBXkSYBOjQAz3Z
MMf9y0lapqDYMI3Kj9eTsDc2xLjh5onmPGGS7cvcM6gqYUsZkuujF9i3g2IkNfJvQ5ZNwURdh/c3
PgKaJaRTwFIDwqxZFh2wrb6G0kjcVDzsKiwpXlPDUCWrcsbgXiFtq2Otg6f16h5KDz0GhSU63wiN
FMtjUhREoy/ZZu11Wr3hYtBH0ZIBnMTlsyORxS6xSnq9xiNRUbLstu64o2O1UZq8E5nCpeI6y4Mi
WRyb+ZFNFlJX750ttg7T4Xc3ZSkT661Sp0lOR8eSWbkRYk8xRCVl0fO47AAZ0xUjd7pqxmiQMWFh
y/8uv2sS4zyA+QP8upFgz7gY/+yBGNDLoQZuoEX17Hkrcu/QX5UzEH1Nuz0WK+m6i54ULWBp730q
/GqCk9c7C4lHS63FMi/QiK5FVnyHYPzJCwu5CkuKsscIU4addEcgedTCtYQQKAfys9bf+5eBqVEW
C0Sn89+AGpJ56VwRoLa60V1ji+fet1e2aNqM+IY7OZZsyq1wMQiaYeEr0NanUsysYypFbH3LxZ4c
0Sp3EhlaXER1L/K1uEWTjZCSAnoxTIlKZmXhMwnxk9jLjJtZiXFC+++n+7vriVRKfYS8DFP2aQPg
PL011j8pMl3LQcTJSGq1fIMGI41wOm06Fd9iJ4cxSQnYhRCDUKUvjmaKgZUdCy0l2Ccb1xewKRRO
pn47swixuQRRAN+ndw7js+5KxA9wFepfq0IwZicv/M5FL/guvk2RjRJm7OAx3PApGPb6nf2/sCrS
VLrU2zVuoUWTF2+9lYoxp63+nV+N6afBfR9tMHbnsJB7mZGbNRUD9QC8He4tSp8ZWREYKU/pOl5m
vKLm/D1/HXe0jAw8nY9DZIEEupSSBL6Cl6Zh73itChRqAW3evHPrjn2DkWnwDIFf1ckVWhKLJk5R
LfLQ74B8PJ2Icn6DsvQEzaHXh4EBJTFi92cCoo16PW1150MaT2gdoloFvDcz2kNdmfItrZavIEUj
gM0B1IQrncEiQHyIic2wOh2nFwsBQD1md0C+LdD2jlpj8Y+j4jBTGFEM4WMqD2sKfU++f3XPGwBN
tYBJIiSwT9CTnnMXHUHO+9czrHUgpaENRuRJ3b9BONStDnBUcEXjO0kvV4smyzZQd9IXLlu6175S
BZRpoKn01myQoJBfhG2h6JN4spzLiwa0wg9zljU4oKGOx0ZPdE05e0jpGRCIIKTn/JEQ4LfBKMNQ
AnNLBSLe2WhupOAlNvY67WgrOm+MLgsHQjPME0BaAHi5ZsVHLOQmj12xSsHdiFomQ1aMaflJo4y2
qPITXZh/mPfxOLhAuvREI3VpSlvaTRCwngJbsfRK5Mqe1fuC6TdJLG472COzqy3V/8FZFa1SqmZK
l3urultREgjxd5wYukNEHUMPmz9Mpjtydw+nVd95+L6HxePEVRyWhZybQbbkw2vjFsRK6t5MHyU7
0cG/pU8L/7EY2sMqmWbCINvwtuNXSZh3UJQ5CQx19GOLE4Yve9Hk1ofyN5y2+ZtUDXrSaFYVmQbI
RTFGuhzHFJmdgI2gHRv86sBr0AF+qYBwHOeLVoXRSBfdXpH5G2jOLC99bSTQkotcUNYBcqxAaciy
pinziSVVt5bCcSHvH5Ln8UcWBJc6/9ltF+QpRr8CRCLfNNiTl7Bcmy9dLOUmFb8W8P2aflDs445s
uKfVbS16pAT6Y93lfJKwzzFo8C0N4Dmj1CmGzi2/dQ5oKjtL0tjoKlqDojnZ8FJ4D5VkH386l2xq
cnHtfIcdYfjGb5I+52mt6p5lhHEyjLXm/srRD4nqPM7HvSMUU4I1yHFOZ1oAZHIJ1D7g92WX7FDE
jmNFDUgyD6q0cZYyyQbjbPgVMmbpGUEYmVF8cgEYn5rQE0TnZS+z9QmhTNevdGHeZRsOFn3uZLdd
oCJnyKTy9kOurPFv5nOLhp+6A3YeigQXyVBo5Sb2z+8vF3z6TINIix4kaUE3ILKQ4q5xHzGnr32U
2mslmmY4/6mWEeE/Iau10KOqPL2WgeWkSf2IN6sK5Au5+qybEokjPNMEexqzgS14ONywxoygRkJf
UddxanluGSaipLcodT5Xr5dOGZDx4DJQ8UI5yV/w5EfNURkR/BZ5v4Fd9IpY6llyiZIxO97T2OLG
ZKZsxclq9Gy5V9Vj4PFMTFNAaa78+RcA4+jGtuVytGMach1vU5L/giqtMqYrj9Y2FGIshgS52LTq
vrx6kd2Yg3CRD4xLU9NLFegNyynbDFtvc3uX7lfsuVa6Zsh0RdaAj9pOYKBdX+tCbjXw88RceXr1
5NiPUK8I/YmVCZJ4FSGVbh3nNaImFIRG+t0WjuyQg/FXXMrH4iUJn2oqJ76lZ8FfuR0qpArCCRlP
cygztT5WuA3ybMUjhcFYUjlTeNIXfmuvX2l7lA+HJGNhefeVOGBDnI0686bnHeiRqnBIQJcDBS3D
2UG0NZ0SOrTnNU+Wrwze/GFRSfGzaWmQImDrWUeX98/ujYcSLof16rZzpda0pHbkOIjlCiPpeZfS
ZsVk7YrK6HLmSI8fNzOeOPbKhrUgcGPvdDuPO9IEVU/Rvj/zjBBNiFprM/ppF1XijAiidvT4pVTh
3lOBJg5IQqN0ALrdX8D3jgKaKsXvvAoQRaRxNKabI1GuArARMrVhPMlRMQx02f4KI5dI6qkN+cst
NWjon7zDe5L/TnmU6TxMooVBH3+YPOTZ8jqoGSoMmxPgJH8GaLAzR5NCWCNX8/7uQMpN7Pk6HDNR
R8I83fXpHd48IPDniV6iK/2kNgWHQ6886bNHn2g8W6ZupcP5qi3qO1QGo9Zf9FsNK7KXGK4qrIh+
C8V1LFx9jhNguxwPjmGUk/1tJq7jMQVSWtulcAzIaWvdY843qgBKnhYG8nWe7RSoPQTzSxfad61p
f2JmSldLLU9mTr6butn7qa3WDbXIoGGYvYtWecOL3t9sXUfCE1e+FGi4RYtpFpe4jpD5wkTb9TnL
VdoSA/xt8Wwoh06ZmsaYDABZkYKbDcay0alBjSSXeHHzzU3hl3QaGa8yY11e0B9zmABS/pnbCf3h
HP5GigrN8l8Dje/u/R7JygQf0cy5XSu5vILjRdtopkJff9Z4B9HyOqTgrowBLSAPF51Qjkc8ETSP
5ia1gCJo9feLUq+3xKgzzQsitYSij5BV5WPM988wYS6OiQ/+j/MApwqgPQmdKsVUQVuU1WqoQ6Y8
6BHjPHJCfRBbuOLcvv6AW+4DsfuCyEo9S5HQSEtjWmQwNWwA/r6l1lvjZBTnKmqJWeLXIWkARO8Q
cFJKayfpbcnG+dlOPLYvkZV6l8bRAQpu1wgJXdKcXAfd4ofiqmTdudU/NF3hTcVkeaC+ykf2+kLj
Q6TEg+Paz7ee5FEnHURl5Otn8VjocQnPauBj/yMJPzH9YpRyj+eN1PPSrqpZFT+LLdTiHck7xyZj
sboRJEokUdJSya9SVlY6JQiseazIRQgOEkx12jvA3aiBr7q1Hm0slvLSLJPEHrf8t/Bs7cjEf0vG
SFTbPuZEsjBOZYeeMdf+pK89cxz1q6rp9bimvs7A9p4k/yq/Jbb8Uv4P1kNXB6GZADfAGjZPP3ev
JkpHDrywhawuUN9PYmyN/NNwo63ALCMEISTxxR4uji4vqjddWAlV9Q63WCiJJhbCdODB9BlWlLVU
/InX90dGcDeiOoJ7zD+FAFmeYP06lJ6yb4nb7KDLTF/rD/Q8+vlhWsKGAj7e8gVGAnlXfEwAFph4
fLU5M3ReC8/Es/kbP1V8SYAtHUPu7pmLVJQBkKjSIN8l0aP4vg3Kb7rP80xTOSJkkTD+LVEliaCC
nJBcFZlhEUQ6Vs6L/e1JwewdUaQt5Bw08CJsUgsl1SAfTg9a05IyEVDVdwrpZ0gL+wOAvA2bhBZc
30unevazP7phpR2FAsm2cLv/F8/LDqVUoz6hXbw4Cl3xTgkt/DlBZa2acgD4lEnemH/8fZIMN4XJ
zDxnPHiw1eW9HpKQ8QyaUDEMcqvRJ0S/wsuCrNP4T4YjduElI45UiTFcz29+bh9T+ngXpaa3yxif
AcS7wUTj8IxW/jQ3r/cASHWsA9HOKJvJJaBeiGi6zFZzgV11AcXLgEfeAF91vkNHLk4/nr5PUewt
IFp999+iOJIXJfmjX30ZTS99RnPRXTcbUVVBBSnI8G1GIJ5nRHYpAWPdhgeY0uy4O2aO0J57XKHs
PXMdbZVychOT7nbU2gGGptgofVAgUQtKkizy43BYT4VNDdG/xX1wuBAkdP0j5rowRh3dXbxYBz4G
IzwLAa5rf3mX/KLKMLJYDBaWnT12m6+btlfAMqN+wsM9FeuSN7ZbNp8ksNxYlojPcAmFjo3P/pBk
dyAKXDCkJGPlaJE/vkpL/NFXmBL3nhLgRusqDjP3LCvowUw8g8BV8xii92AtbCep8TRaOV4c8yLl
CyYnuAyy1Aq6r8Kz4n50J6IL0lGTML3Wzl5ATjh+WPu8fLwuDEHMC8LirT3J0TJULbglvmbhFDNs
vabcxmwFEfxvCTHCOAgenrNv3wpr4w2qu3vmbCiMNLkBnLDXONyTueNMBfRpTwCHXdgiDl3RVkgg
G2mBer5qPURvnjPmFniWhMMvPIiIogGpbDtb0mEbRh13QdjsZVTwBk/76Wp0dI0SHho89egwBvFf
14zijKGpCl4BeY0JRHB6Nxx+0hcNQKRvmLb6YEOfaBTCWMzT+JGZwp5D2+xb2EZVZKGrISvAAJDr
mG//dGDyafC7ZXzZtszEIkXD8+6xMXSQ5vEe+EgBAczSal3B12XbPsMnCtLxQ6cRCPpKsCZtWV3c
rsAdqgHdBnqC8nqPR+e/3nQpgy0WLZN10xlYFc/4stnBTNovrpzkdKfu3FIJ9vH/nBBb+lbPOPXW
MVbHxKyexxbB1/lHaMmAVIkHE1pHurStXoUuxyH6a2xnfPVs0LFxLRLAqntUjomTZRd6KxfTCqZ5
nTwURUx9Zo0/UZcpPqGuFmY4Om8YABU4P3xmdjqd5UeiL1t3ivnmritRLeQx/Hr+P4kUB5zPeUKQ
mMsTWm5vrlsKK/UGO8qpDoGy8cF9RDpzZc0wI6IYKvMzpQ9BZILdKi3aFhHYUdd4noQG7Gk7fkj3
RkrDrDRPN8cCuB2TITvRppnruCv0jbZtA5Ovb5Gekh/umVDm1HcFiAHwiGAVEElVtkF2g5zJY1fw
gUtiMosCINAPG5PJUDDJ7ti3RL6tNu7aSlkZX3qVYkWhjz/uPlWqfi52brH2Zi7IxyrjL27cnxhF
g8BWw2DrTSt5ECnzZhPJlBhbapCtw9swx5MlIgXbVrQHgwg6Sqg2gPLwoCEDDuZAiE9agA3BP1qz
0LFLbwfWexNJ4YdaAgia1X7ClFYZrVjJOyk3OVKY+eJ5AcmljlmcUnHK4CBtpc9uVNXe0mUpP5YB
BsSZOrQn3ngPeSYXHhRmKcFRm+sCmmqJ+3DrCjw5pYZoAKzKtnKLBnDk+A0PmGnSSurb+FbxnIB9
ZALYbDICt5TCRG715LMA9Agm5YMyEYPR2msNGLAbk0umu2HcfSJHU9xNbSvs0pihMA9jDXBoDxc5
o4g5STCkAs9LWCsVvEwAx+r/6EsuF+LfZPa+cBty84pZLtztP45bTpKriPb0PyjqX0tE4KRzYCiO
9atiJQ9+mid07bnn2qIdhVD1Q+xq+xBulGIu0GV0HkqLJnQAtAWlXODip/JVr+s/LZFISVv2sxyH
jC36SOcrCarH6kSHIWsS90wAZnkv6e/3E67je2xAttDV7FcwUxTnL1vp1vbNZ21qxPh/ayc9sXr+
EERKP1/I3yuowp6ZkMlWO4XjrGf0jnw1T6A9a1V0fEJN4IL1AYRMkougo1J9D7PYOTVmKYVdTPZz
fzPwl5Oy+OuuopBtskaoINbXukws1Hip5Ly/blFiOpYxACA/I6bJI2mW9H9HcuwyYNdQ6Q7+7YSr
CSYlttTjYvEwM9k3SaaGmKTEvaJ04yI25lZm4+kQgafK2imVi07WyK4HSP8QBad+Jh0hO73sGbNW
u2fbKxwVHkPmMLn8W+AVijyMSuBnFVpoW5FFgvbs1YcBhqWhEbZLEnbA16ajaMFa/xaAxsg5bjKZ
gwPaKfnm8aT6LudsIJz2NW6ejnQvgfP9KAX3/QboUFYk5WAaJ50/kfmG14w7xrBJEaHN5F1DShq7
FJI158iW9FuDmjnZxGSD75YCOR0CGtYNPih0a8kZyYBIoK/FowRHBuIlzvSHQHnXrEu+9/oIBdPI
qlxje0OVt3Y9zy85D66cPpiwigic+zHUewSXScrH+HzvfN73P9G/6ZaVyeqtaSFwlgQ5qaREwcv/
4jLrweYSgRjGPkT5AMszZkH3jKfIlN32pWP4uVtTxGhv3WhfIoAP+pjqnMM+h/5/A6+0GzymENFS
68elKPSHeK5q9GEngI80uozWp34OV24utlyYnZxprquygwRDREY5/GtjX0mgHH7EYKLoMpicyrxI
IzExisEBGFqExn6LAD6OQJhFv8HWqdJYqngQ30OxxYh9iVSkXK08+7zjzLrSm7d3/+nsqti6BIyq
L4XUKyoB3PeqUMLL6jRTO8S53GrO5lii/ZeZ9hLiDIcqh07AWNhHnoPmj+atGT+7E452Q2Uabcsx
T5gx6hBMPBKXSQODBzkmznGiw5XYfS1llGlk8qH4JKyJ3MRKhk6dJuVORgc0c5VOi9QXlBffrvPf
lJTZB7miItQTNhTA8hl1CeVuQEJiWJ1tShTmCJ6Wuaup/Ab2vtlQQMi5b3v8zF03LVhW/Ks63cH5
oujE3CXwAzq9L9z0R6sKmSlWRMING9L221iD/Cpzt/KYz3uJnNgN7z3j8uwMK3Ate5H2QkDcUmUt
YTochsVQ+c3NIN1HPU27N2jAMbw8t60XlMk3Pjq1N+XldVeukk7szEo3W0xnMqK0omkaM9PIStmx
ovCYBpL4RkDu8qi+cR3/9/GCyv6K4Le7lEXOKlmy/mpPk40hDf/vPcYcPfLQh5SGjcISEDXkCXI1
SoAlLTRYWPLzMCoBAkUJzE91gS72sXrdFq0McRGa0LQ5HV/N053u4/+c2ME17Yn1Uh7cNZB76Yr9
msiwTYZrB9cjNDHLiD9h9g/gHRU4GnILhTUN9YRz8SKWh4Y2e4GCXkG39lS7nC0Olb5cbPnEwjre
6W+R0CyE7eAqNRytLwv1itPVzdNccvFmeIrVWJsrHGZstoBDMWOMBacoDk2zPc1kc/lhrHTLzysa
G9O5mHWtQ2BuM0LoYY1CfzpcR70ViCSAbkEDkE1OrzNwaVvLqBKnor1V/dTPDkRN2SO3vSMjTno5
dRN0+LE7317a4/YZyc4C4mr1z9HWnw+x/nkVIhHGtloAxtwmlLsJN9Rj+LcrAXv1003SD+phaAVd
X9e0BaHCq0dY7WVn2+knetK+kYB5cHmser01dnfhSqvulxwqpJkjpdI5QqS/Fy5cWnQwc/yMCdA6
w2wMmfih4lfaD4/uJCGPgjMcDzX3ORTJUsPCLLaO8UseNsoGT6iM3o2lVDOuilAbg4GMjqVwFTAB
frXfGCSyxFkqx6khyq1pza27yCv/ThTkUg+Je8NHuyY2bH6yqAHluU1Th31UJXj3GaLNR+2i5qRy
5LnvdyjSEDcL5Lik0/wd1vcmhY2LqnsdXI+f4sIdlRxs/m+TmdhW/yMzlh4BZInWKdBZVfjbw2Ib
nOVLUSUYRdYKsWOQ7pBu8VttNizKdUyDFuGZ3NxM1daOvP0bevVOk0O4xybkWlmYDc7AYDrn2a55
tRx9+kbqGtjH3JK3RjrpHrwlhWqKCd+YfxTjnuNQH5NSg4UOsGCo8y4Po/wAdPuE0uPkVjq9iwpQ
6PdYxrudJtm0HTadxs8mel9GT/53jCbqVsX4xM+1PGsvga4cjcynen+aQ2MJ93v5WJAtznAuV93G
QMDWd8GJARqvFFja9QUhOh62INjOpyQcSOm+3wzyc/IEh0Kdx9gK42hXoBY3wuugomd/MqNGEC6i
MH4/LoGdLX3ZKlWivYsVRfO4Ucfpfj0Hzx10xfH41WtKv8mNi35FMhkizGGhJfZaQKWlClL+sIx2
sj2wBAGV9Vi6dKsi520WHJ1/BahRAuiv0FtzoQKMjZY/0EFOVnkkKInF0YxJKKqYqCcyl9MwDifp
K8ytLiY/moAf7idE/85dEJXKwsgavE2EHMtdYPx8L+RYwHskpoG6zvOv/TobHR3PYDWADuIXFiye
swjgGEp+IykoJVOhUARtXe7ULenaZ29mgaPWHyIxPQfCxcd2vc+0YBnTP7UlGaoSrl5Zh+z1f/ym
LUJ89xMEn8TT60gPAWc0g03eiJRUucl+edG2M3Tq/IA7ecpG2xHfHocBQx390DYA6ggOrkmTfBA2
r4/+o0Nwbw4d+7aYq1CfmtdyNbJZcAi3pnigR4TCVoW4Kmeb/1xjBn+DMtlW7NCb8F5C76U4cCdV
aLbi0CKLxuT49tlPM7eiA4HJTKa3r7w5tlqS0VecgsGmQzs9+mes3D1BMNBbTZUyNAlkn/SnaTcI
lovgnyLgDcc4Ae7Q39XQudIQJSvLu59bSE8wQgpHofHyqivXjAzGzljUyGdXlPwPlbwMJulnnJbE
OeMlGA0GNYFr1kbLg7Kph1fNC/5p9PUbXcv41qqsVOIHxb0nJ/Y0Ot5Bj4GGEGDiDoRkM/Ace2bB
V6tZIu72onQ+rqs5cRoX+8aOZkmQqVRduJpaz7OJxiWebFSlpIhQkc6PGa5lQG/t4MgLNLjIVupL
iPNRd0u3sIr9xFtLyt+zqLFe7chQPt7mtaith8sD3YdYO7ZKLnNUy0KUv2Gx2JkVFUIz0eNV64aU
oUllUc9Va+gvWrdr0+sJR7xOMWBKNSHuQ0qqP8FHqtIyiVWNkONDD0hp//iJUY0dw/2mFTALBJO1
9lWt6dxkts6vF0mswn0jN00jnxLzIrg70+8lY/zeO7QvU7cKT5oKDjwnQw2c1hX8tW/FZKC8qEc6
v0We9DLflCtY5tlbbk/AaDz+JyBf8QkPJg5u05d+JOcrWxx4I+dzx6khk1pxMywAZQxw09n12R7I
KukCrqW3FbLNOnbvNmaxMjyU7WMvB+kRzKluRlWh4oXAVwqst2VwEMeamb2kLDwSoew//tt96x3N
QbA3sLZ0I3xP7AAE922C49N+UNPrJ/Qf2uf46n/GMT5727fYyrFJETq9yrYvTFUHNH2W29ye+ZvX
Ec4EiIaJz2fpkfwm9H6IypDiKQZXrFxhtCXU8t1swY6T/U2raAZVYnV7P7CgiZOTRR8pOU0MzLOg
9tv428HSNtU+bdCgqwssJuR9HjlptDWXu79umGUFAfTad7zD6F6zfEeoRc7fuNjkJCOTLEgNyoqc
kKYaQg8Ixp6bnP+kxYqBeocSw2XaVWytuLZhTxL28S/Jcs/euSNXNX/9nE9H5aRh+NEDxVlM4d9J
h77Vc1ddp+x0SUDjkE32a6ZnnUck3XZAGK9q9a9FmnoLailIdLD35wwkZSWNDfo6ptAxZpbsM2jv
SktAVbI6t2/+M1iI+Mqlx4mwV8+KsWA3nEKddmKrG30yXMjarV9EjJfe2hb1ov0iMgLDa2X/MD9J
dOBCwTLvYNq0t7IIoZJNREReKIlUlpMHZNvElz+XiwWBum9Rn7BUHbjd8E98Uxdh34A6YICJ6j5j
XeJWcv5MErQFcbiixqFqdyUJfO2Wlr3iErMnimHH97EM6NjwC9KmyNBTlz+HDDUP1CSRY1hb0tC2
VH5TsS2w5rmVSb+Yr9+yC81Q3/I3IFcjue3jVSXyCTl3g4ZpUinIYbrcxH8W9vUPil/CvAajcX5k
F7cLtvNfR8Q4EMGztAS3n7ja1dDYcI/urMXL62Q1F4SpkFW5H/qblPOZwjlW13GXkgjCtqFtb0A8
7MLB4EQbaRO29t9xf4HZ6v6TjFov04iN1WCbJR7gLz9cgTHHwkJtBkC5fg9C1XMFSNnqPR9kfjAx
QInnD0gOWaIGQe8eUEuRNt+e1ky88WdAt6YBaqJwuO1f0LU168kVdIlE3cK9uYPEt6K1Swv+sqW9
Y1TRj7HrQporsN3VyE3kA1hKa+M9robAkTd43VydvtjMjm0XThA03BTHlY9u5g1bf+PwADzJnQ7e
ereY30EAtNkocDVwZcFvw30ge5/a7hFQr7X0QLopo3TSjC6vN5s6ZWzwSELCop/PMylOF4n6+/2A
U1tlBByyyFOEd9MBNpC+Pmn0EWBc0fKsDqg+33oXYiz9r/nCNpV5sgdj40sE4LEdKZgWvLx2A7OB
4vA2S/HpljTepvN06lMQZ/jywM3IugTaK0NA/xfuy6ZLKflHUsS0OdAgHQcvechVeXJNprAkNgTj
5xoUTM/syr9iinRmk0+iCQNkddF39d01u7gAh97C8y/WfwIvmyDQGJuKRCIXUgraehRPqigLw/ov
CyEOHem0nLBT2pLJTo1DkN5M/ZRkjzdyRmT/p3OE1SbnIDyN3jgLBzpr2SNpHsirv1eygsEZFF3Y
KttSvcT/gWZ7mb6zDBCKzIO6iO4tQFog2I6n0MIzocRQF1dDb3jRgXNze60uYm/Y9FgBCsVcWZjO
9/o75RhlC4VlUomJPXnCGmG9fhHWvfVW3t3yU56IjBJRh+lcp1Xb8nKQD6voS5/V3sGfhnGVeYsL
nUdjuxXA2CrAtXls9PfCsPH39vYwY4PlVa/64ddYEdg5TksOmjAb3ZJIVD9IOi4omshP1NsW3/HB
rTbgCTK0Yh2XXUuPcONpdpMgr5zrAbhG9GXp2v7XrGN9SP9Zk4cLo/YqSX31njUQZ2vYBbl9wPE1
SfrBGhw0cFCnArzFbE6cTujgfapzcnEKF8ctUkEo2THi12q6Zv7bun4IZVK7uau7qwR1AqfM1dQk
0D1+kxFg4cdrdFZZ4Dbg4W/e0db7qMD/pqGxufeQ9NzdaDj1eBfXJ02KwzkM5Q3ezx5GUB2JN1nN
B9cVmBF7FWLuCNCQJslpqlDMVxmGTIIr1PSrGw9Paf3cF6TAAqUB/FYz32sK37dpUSRSI/ERr/F3
HcfVW+Trp0yhdhAJCEimEPsYU7WNAK0P8Y+qxerSPvq3p1KuFXZ5o22r/YSOhcTl/JjAEemcNGyC
vSA6+5gcq3uQ1/qkzImTLknCtjt/KzQdVZ2fNjogGGKRQzcHEBgTtycBL/sq1q5iqPNp1jmzUBpL
I8wYmQMaIDvj7kHquAkX65BmvlOncrfxS77Wh/+VbZQlGGVrEwUMq86Wa+L9MHa9NmKlDBY2Bou1
fTm9dCsqzrBSuTO9WjyFW5Ad/6HsqrwDgPLg1dS2jIm4seK5D3jjsHFdL7il2FP6On/YqLNwVcw4
XdHu4zKYf38BrX0xhLHwq0QpfPlWwxPdlvR6h4EkpRYuhElJ9gFuncq5hplnRDsNAFSLMpouDVXz
PxWb0nmoE+p9etqKuTArLOCpTpxr+BsYNVW+xPJc1TxgY4FFgKzLHGZwtN2GexYDgzp0DZol7H8U
Xo057sTiRWuahXE1c0k8vuoHmzAcJ+x3ML0vj22THd3SVihf0dN0RYKcoeovsOwF+1V2puGh3Tay
fLUEmFoaEHcegHZA8S1HhLaavy1oGuMvpKUp6R6hue6owrpSE7UBFiawp3ksDkgdwVeuH/J1CDdQ
QZ02soOhGwhb8yGzLIUgeDu7QvOy83DSu4T3syT5pUy8+5eVH08I0Z2ilke8Swo89o8CylajpmPu
mvmMsgipR6kLLaLEhKqsGUgk2/uby0ORE/jitRwYUmMTW93CF4ZqLGLOPlLOlCPl6EaDzfjagfET
EG9ELNDK7zszT6UuqzGoL8fjqmHFMiiE0hKXHXfOjcfjBacPHql2gTnSgqgC25i8c7KznFmezWvd
4+BHxcsZk1jnMFRIvnBiLK10O2dNTnPE5EL98ZpXLxDm87NX/V1WkPY72CQODDBgMS9/znoC/HO4
dhfTqU+L47Abmi2Zyfcaq1ie9UtkEnPMnPzEUIaB7WzuZPDbc+DmL5sp0bjFFKA5SLfRHurPWS3C
mmahhhiG8EamKYapE5tCBJatRAbZDHTYZFChJYjtU7K66VJYIKjCaMiJEZvGWvfovyqjmY5NYMP3
KJbrppIKQ1s/+iiLf9geCXbkwDowrC/JsPfuR8jw0Pilabwyt53MGbXKaVWPQrUcVQLY5aeYjcRd
TPHkyo7Kwzl1jox78uD2ouEssg2iTEBMPWiFnCF3ekDJghNBZ/PV9uBYrLoNh/5f31KVzuwXmB0r
CWcISPPAexcH+hulWNcGbbCiE4oOPrPzRaOnEOW+oo7ZbcyvLAh4im6ZAQRalwGtxvr63aG4lo1c
WNwD7qpvI7gwKWq+bww3OzaR/34DqUni34QDmQzXl6dTrKZD6vmppj27/O2/HQvaHTrTYnV4VP+k
BBffUGEI7hQuDOLSekbnXXAF/LyI+nenL9pDlKNkexcJROh5RWCOGVzNQIu9xMmfSZH7/NU5jr0b
GIakBqkb36f7o737MvGQEVZJICNTLQ5VfW/Cl8YBKIjt1aprGwWH3dD/pmzzn0Bv4vzcHPx4OfLJ
wAqOIqj/NO89wwhbFq2oi7x/2Jk4AxFr4kLEH4AG1n73qT5C7poMkU63pACzqrhueTemdeYGCvIS
7wjsOsGSLAwVYlZQUCr1y/KYlBxK8F1bU6cvuAXTTdzjKH7jvjrZDX/2q8dQxNLy6fJuXTyqZBOD
0cg76+Vymoz2dUu9UpVUZBQunECw0RObnrDOc6HYeluA4c47muAmXME1auByiiLEh0p5bmpIGYBS
J0OQx32FkF7J655Q+/gQo09b3BHDiNwHFmwqgDvOw+MUlLRZaFCTqCkeEDLjgSPwpc11qN50zPut
A6ZlPVhug/krW1JVuI9+wzhXa2c6z8N4QYsYwwls99BLDWqZIH1HeI4gJ9to1I5Mk9nQhuBWLDH1
AfU+gpwzw1iAseafwLH8WdZRmBO8gi4aaYpv+a/z36xmuKefUeEwHbfFm8BnDp7E200RqjGV0d8H
AQBcNXxV6NE0sRR0IdNCDWrfnzN7CN3JqYLl6eG8ovJIErc48HnZeK91Ntly4JolnH/oOu2HvwzT
nlcQzAByJONXnXYQA4QcP3is8JHy12VH7s2SIez5/N6tzoHEqhEK2vCqKN+OTwyvUmt/WvNehnwX
GW8b4Q8lnM2G9r2VGRh8Hsq1TxrBuh+05FPZqnx4JV35OkkXSEp6XEdlZvWDquwgz5WoNChCpYfY
Ful3/andYuXLz0We/XPNs4w8MWITCtsgHQHLh5vJUJuVnXGjcNkCNvCgELlJ7iKJ55bnl4yxNc3d
Oyi1muV2pb321uiupYfArD9vJmp54jCb6B7DLexwPHx7OQbp4a9WnjjIvporj+FY4s42LUWDhcot
FOdXYdVIWN4gBoFyc3wPLGiEH/GKe4liiAiz29XGHu1PwvlWv18F8ygfrGC5Hv1Zmklh5fkAftF0
WGfNN8ARR8SiqYmh842f3j4qA/IjQT/bov8cnv5LUKXQDukF/pwFsnwgYr7bdO4ERgwVtqqyTh1P
s/aNphtfPKOKvzvaV/Y/tKQOfvOP+GHIxVNuzUytrBSfkix96CDTtUbLjA3qbK1Bnf1qNPy/Jz7Q
gDHOJuywk8quu5sb2lUU++tgoYp4soZSqhg70py+3J42qDuEDRParuBjSzrurAJIrf5KSEeWemTp
jvzkfFsuds3K4etgvrgbGsCdhAZpggblLD+jB9j1DH1QMGnYBcKTA2OM8JODf3oTn9HfKt3uCxr9
4BnTRyuga2GahWsDJdzPZIRy8zRjsWp1B8gPbIEvbponnalqffg2b8djMz3IyfSTqnPk6ao9xRcl
3eCiERkH3ZdNQXcTHaGLEjCWzVD860D6d3OgJQBbibD3nn3AMO+R/y1CBHRA+SPxhUa6b756z/QX
bDBmUNmUtYZ9oXa0izkkd9H5Po4cK1DOFpaN09tvOxV1inDp9wImSPl/WTdAr/2ODJ6LYhxEc0iE
VHiQN2Uf8OEhCmjE8XYY5dmpgK/7aa7vrXJwn7e6Mk/ViUduo+5h4JBd0I+x3tP/2PE01gAA5oOv
R9lYaB1yTdCxLyrE08cbqMTITnGXueKXdNp77muAK3My7B71/oaRbawUS7jO3Z7QN8wJiUw+V25C
2xkEZTwJFmO31tBmI5h/ZjGDbu8VzeI9nuNlC9uAGZsVtkkeBPrzsxL90ed0uTJ8ipYdrKAarE7l
+ZWMJCBhQl/+oCBI6xAsougc9ikFFXoGXYvLeB27bQTaFDw4zLT5Xuyowf2VDFUSb7CgaSN0vnZe
Tf63cjZPxCh9angNDMhzVZhGS0PyzDWUCsiQuLT72TFCXllAHOGfeJIQ/xO+PAdB0eWKfVk69/8w
sCXyV8kVWMToocy4HyNNA0t4bnXSDea1tW4VdVTPCJOErAr8Vwe/Da4Xvcv1htgm6lrqrh6ykljA
aeifBIH3ADv+WZhob7/wNSzg5u3imwoz5rqnAXTh8UyZblY5lvfkFjjncnlEy5Fq6BQpnmeuOPev
I45lgExu6+DHogHPQ0YEOyl7d752i2xSW6V7DDYGaR1P5QTy/WkOj66uqYS3PGKwSNiQaSteAP7L
S5oAxI00FLvCvG3HbP2uJvx/BnULFu4ecpSDe6ymhT1wsgomJrXgkRG8aGqOuj3DwfgtTeyIFNc1
6iKFLqLLPN+QBY+Rfzj06M8mF/5Tu87uAq441j4NJxxQAd+63N+bLCZGGChKjKfO5EwKwb0G9DDu
ZhvzFcQ3ePAPOc0/bnQEvsguO9cSCzxGhKEdY8FVIr/+zHzoadrdSm40NLznjYMjt6j9R88ECTMd
ZOnN16hv+srLZagmatJ1UH5XQPP2bjaF0DZ1hM3sYW7DkrpMVd59uNxoeqRNPIVE9Qqs0wwRJtKz
l3Z37LJo5XstB+askx03o6Zw/atQgwY80CpjAyN+n+ftKl2Ds9R3hay+7JyWeWAbeMCSik6kMaC+
Pe832LIghZIV62CD0N4KSjcUFDM5RWsaheLJFlwyqa5SQudGubF1c1LwXZ9ZV5ztQzwH2v7ie4YQ
jwW58b7Ryd7dx+m/wewVLAUB1LEkKcMTw6cBvUPlZ/LZGEs/40NJCsv6Fsnor3+MXY47cyrYH6Sx
KdovYwdlw2DORYL3tLM0ZFs1qqOPvZJtMAHENQoJdurFNxPUQ6IHVu71MMpNDCqXF/ViDNYpj53G
aCa+fRM5ZZsYq6qqKLdtfs32M2+zZTuNPFszYq0MJ4s8hvtO62jJCtplWakTZHbkQyQVt8j4LEE7
/cvRnxuX3+PT4iUIP8C6/twwEXF8eltghvt5B0QWzDOjLwpuFC2CxS2lsl0p0Pl5l5d/XKCKRcuQ
LVf67Z1XSUbCjavT5nWaSzAunkQgkAr1105sFE7tmH8/gcYWISXnEkB+Cf/SL8T3ejmTANSHoPPS
LIrQNTInF+p4pde8zU4iqrmvWpddhc+eBQfuvYqWXkEsupaJyt2+lTVC5aPKktGmdH32fCvubC8J
En0rAge23D+/GVU89umPlsa8JEbkA9KvmOnNoqEBM9Bk/r2h9K40KYMw8HRJ9uz5rDoi/3hvkEs9
ufOUpYLNp/7S24W/xQE2D08YCQt1Zaj9L/JzmLud+bZ5xaItzZVEwqBvIMck1UnRdvFco6VJvmzT
Qtj7zg7WOvtSGMmhfAGXaSkcH221+sKL7Cypm7TV0Uw4pIM4FvvDiHkWtswwdp5DyhZIAzHV2N64
TTpIJ8Mpvhsw2AqBTnfyZ3d3vEonE/gOKaiwCmwOmh3gtnPe+HPOVkFZFjtqmZrMiYAxUzRbdLwg
4FB9RwRFecBrjfYoY4Mv1Zc8IbYuYQrnDcR/CZG//JwE1ehRF99/5IPDK2sLOytnQKikg/wuxN92
DBUL45VMuRddnQVHSxe9ROtNs6xvmHBeyScZ39pqjH2Aemrt63B6g0d0/uKF2lasQX/FXmXvXpiL
iIQx0kg0dtl+T7Yh6PSQsyG1Ha7vTzCxtHDTbRJnZwfEVjp+w3NVnKXR+QkjuYx5WuZlTC2Ifoxt
H3y2ItYgC/okr2wjChJiu86A3x/ODx/G+udcG5Q4vxwLggaOAFqy3Gr63NSl1zvKYIVxRGfC8+4A
GRSKJ89wphG4V51LmIoszXEBhRkhk7Lx/jb/2T8o6Id3J5V7o2YeiIijgc+BVUDNHnyC40j0GCCH
vMD+MFeNF/QcerbTxsCMfkYe53w0NFDPOqYmzIvzSUhsc50/7oyFVopMo59EGqmtZ/lhQigLUWGt
g0zB+gC0kklNPtU1LtoImTZfQ6yjo4hjP9ERKjVlDqiUTeRfN7rNPb8r2jNCy9BlV6MD2e2pS9wl
zkbkl342VQVIw6CrmduLt1ZC67t9KmnswEqFHPdu0FW2YTyKhIvSL+L9GcTuAeLbxTMm6VQdtWUD
/S2MJQV+OACWlrkLIj43eYnx0YezsJXbroI5Z66oM36FwHOlVIir+8Y1Vh01R+TGSumka2FXIEgj
Gy4SNuBPvVqjAx6m4NgkGgdD81hRRyETlgQMd1PFs9N2zdBf4L82ofwC402jAkkNgG+T4MruinIs
vYEYrhyFv9QQcAXHvsp4g1pI4lR8yn7EGzOtSrWSxThJucSfrHiFnvsYEvjfrlYO8aYq+3sVZv2+
JYGqMaOeEYYuz9IZ7hAgI2UZCkQRNBlG+viQnSkpkm1W90NQsHgovVZ64rb84dPjHZ2/pz8EPMUk
RqJWb2TKTEqogZWB9CBTtaD2liHggTBqEJntSqYuTRxG2T/OT+5RvvK7ErU++8or3PtmlQHGuvDc
K9Kth1xWLOYYW7W0MUDZWyGkq1mCARaSSyvxkIR7Lcq8XZuEjFke+gN1vOSv8dSTHTXAkGojITPC
5gZb+2x6yTZRSQT4FSd35NW3qQswhapmjH5qzUE0HWOX+htG4z5cX4mLFBxkuj9caZHaD/jp2DUl
pxuB4DkLm1NkjNE5p48e1WezlorR2pdjHKnrITmwGKwK9rvjJpqHCSgcBc5NSw7pjZlY2kV+QE3s
WjgTMMQ1+1xsYb9ECZi5Qdhq+cHP3MmE43US+wcuGodtzXtC7GPAu1R6Yi5ICvK/Huk2pMnnblpn
k5zNTEQL8VfFWzdrosjxMPEE4ucwgBnJaKPhkUZdPr6sQ9ZIqzkYhRefQ9enb3T0mrQUhQVzkeeT
5qdG1/g3tM+myD2LSe5Hhmz+uzfP+klQEMlxd56fdii/VTyKnyJ0jDL0UcdT8xZRYZNUwrFuNkWH
80bmriZZpfNMOPVT8nDVBMEBjU/bp3nPGqQB7LOH307ZMhszYJjyQ2TrGVYEGfH9qBo+v6Z4NbVN
kzjVDA9EUDlpfZbAJsFHE7sG1jPBWZyw/wRE9c1vQ/SBTZr3+Hfl4ECcTPZ0Wt+dwRUEaZRsDrlx
I5jenpxaR2tSvlb36LzTWK1jt58wpFbCGrIoUOplBddn7+tuFJARKPhK0yaNZMRJpVV/pmqbumL5
WiUPtXGhI2v6AyhA6Ej8ybhZxDSCefgZZOLGL/3VgsrCJHyEhGkfICddUXLuMIp6CTizmzznS3sx
Liktruwe4unc0TZbZcNffCzF9hobM2cvZAt2tWHMZalM+Mz47/Qtsh077DCvxTMBq8s13ttT9cpo
GuiaoBewaP7YI7toXN7gSB6Hjh0Jz0VeZY45nNdsQW2fFgZ/0qNG/YQ6fUkbGM9rBfBo32sY/7ZL
xm0djzwKo+PQ+I4shIDZf4hb/QimGikbn4ifMD0vOMmnC3W/SibP5MpY89fjh2pMSocXjCm4amgZ
IHkI+9ln/5qkL5PWmOZ1XX1e/AhOGDt7aTOGr+rJhJiC3kUAdralbvsL2AIJ6Qrzpe5ZLaemAgTq
O/p7AJ9gkkzb1SCdQEbTdt9eeN04AFDHrl18O9KeJ8/f5CNYxB5RSGNG+YRERFj1i2YL/eIQLeTS
N7wCzbDZA5ya5w4MEBrSZ+f4gvTY0V4QnIaRs+0bn3VSZ91eNOhokO2gcy9omPXeji7e3ytXOFh4
oCK/zcPxanOrTb0W+atx6h8VZjzbbbkzXu+dG2sLAeAhV1LWABB1IGVss3VQ9/o/AJJyJUEHfyAg
sYL77KNbky6svrcyJeTa0Okaw1rDDMTIEvYQaYMOaRbZNrVcdSkdNqE/QiBmyJlpoxALt4ltHFlN
Pu15CrVK3n4z4hfJ0VKeuXiM/vh3CQom1mgYWeABzJ9XJllUPtojWQSIMC7v1E7WkW3iuFMc4Fpe
k5PglGOuVrqM6+djvDnhJ7UUUoMVS8qNScvEIdpRdNtQRcrmh554RVvReIh6ALsCHUE/51wRlb/2
lflBhqeODeo0+JG2unOE7nPlkxrc2SQgdGrgfqH0/flwbdWOXT6xsxB7veZl+dVaKEukfdGSv3VU
PViKJ+I6rVnuwolI737pNj7ncjUaVRBNiu066MKFaKCI7llveYC2S7YvhSKNzK7EH+rv1kUzTBy6
Dev9MWQykbVC95eo6rUdknme3T/5jFH5YhrOlz5bb/K4Kosy7I4F9NALd8zGH8D8YOqd8232FoNd
aqvFrirL0FcyrKoPPX1ZetEuj+6xhq/u+OABqzxp8yrLGS6Aagq+s9bkzpxP8s5GE4DG59iUqxFU
lpk1eY2xeDRJZG8Rq8G2THvc7LGegAI7gCaFd9x9GweB33jjmaLsjV4/fM9KNvykLlSg+dJm6Ziv
vxuTaxttL0/ufSnJmXnYypNY6NDFPU5ecLuiUJyLPLzDeHZ1b6O7fb1OUFEtuq1BgVwngYVp60Ws
4xYuQXCVGRfDMj0vhyFBoH6uq5N2sMMHN0DBTDNqal2coT+zaZmSkMTbqHU0UwyEhihsgZvcAdt4
yIdBvI66xY5FdqtRqnVGHA09lJR/P/0w9CdtDDfzefp4vIBK5VB0d+jcO0w2KQtrVgzQMB3Be/oC
93HjAYw9n7MLMqrceSAHd4wAeSOhw076MUvAqdBcS6E51Bdrt2lXO8mVRCA+5q9Z5/DQ1M7BOAk2
b7mzQLQM6Xs9ezbYfOTm5tHOgSDBPxELDR5r/OnIZBebOCnyGe6ibhhLtxdsW67nQuBUMBBaBdYC
pY7ZqyIk7a6Y2gdcT3QmLJ/10tH6WhDHs5JRO+WNGVjvvG5gU94RQ9os1oT95wE9KZm86M5V7xgM
NA32i4UsyOxWSknFAZTIX8bg084nl8KIhw7yH7J4zxN/FsG+DB9JVxBxwWMPr0x1A9JfpRiPAYB0
cX0YabfX8BAjrHhhc/Zl9UAocGYiE2iZVKygTJ76AaI/tMyaeESlqaTc6EG26WSjEFD+19PRMlUg
lny8zXn0/khqqIVL4vkwQvoLuqpOonzWMZf4IBiZWPjXj8ES1ivogRibolAYazevi/G4DvoWEtG1
f2nTLWog0RItctsaQIG3sdrgB1Km6AioSYPgvfq5TojwqVEYbq1dpwAwn0/2dveV6DSPVtuTnIMa
u1fST4aJXybCGQaNoBTfJoz1PiIQZwZqqeL1ZYLYi29mxTs2kbrLGDEnKEVK0LJvOiWGKmQ8rEPY
+KnAbFqxdP3sqtXgrqv7Ic9NP3CWk4u1zte9KV8h+7MnIhx62wvb7o1rDgcf+md/CzANhmDoBdcB
yq/9yPYykWBJ3tydFWIgjSD93vAcxXNmC+hT9aZvI5GGA2bOAWuHQdl0s3Mlt+3iJFMMlVFk0VcP
3r0ltxBC4t/GmNCSs/53xdkCarksoKDfIpNZSO5M0EZiq6kOWdf//IBES+KxbmHIMYiS2p8kkwsP
HySA4XGsF6idOf9ZqMMlad2gsw5TdSGGqc0emgTb51kv22FzZ6yQgw2vcmqimgxhHOGE5Da5iM+3
rnsXeaS0mrsyToEYLXhsQHC+8IcPQO0RxcpI1XM40sdbevYf13EIukFiG+L7pBI0oy0SRHr54caG
6vdrjE2kDn55NoPqMCrEPHYI+U1GlbRrbxg2Z8gASCuF4c3x2X61GZLNCMBhaRqrUALrJ/a85PE1
f/H8BbJTeuTd342guFMCObxFcOOoM6I7uDl+KI4va2JVIvp78/SVzip7i2f0iFKH7MJGhhOVkAoY
We7pICKUk6gKpZy1iogHJxtMlO+mwUXl4VoZcJ+bXC89qulmN8dKXVQv2RZNC+4BPe2cJ10A2QQd
UB6SEyDi01IC2IMD9Q/JN/bbLRPA1sobZNznn/25ukCtdOT1Vp71/6cgp/Q2GfshAdrNdB6BYUnA
wZllXAPDMNbzCQ4LdbWQhDBlcry1dgPati3Ob0YJoLQYm9bat8zbZw9p2L3iLHxmhdOJvueuUcdY
pCMRh2kcENSph4mJVOS/wACTmUL5FOslWgtu3XxkV9VTXTsQfDFLXxwA0f1totxoa6nokE9ES0Zt
6LfWehuse+aeyJUvr70PUPpYybCcpUjgz/IDNIK/8KzM9Jfkp64Ov6ktymiDJSIfkF/ZfnW5+enO
uudBj0YBRlIAUXGY84FrhBXclFVkyljm+JPxoK8v8dyTAZX0UPxmeX7HeO2mNDTE+sKYAc7NVxiV
q0/RoqMyQKh1yPuaoy1yEeO1HLqMEuBoaKfq7aUvgzklIfsbdvIBWwrIdNJQF6pL4CcwL5PV4Yqj
n8hpcUQK5/9u8vBjAKkBJaYGTFea1Gg4Ay44z9Q5Om6+o7C/PnAG7ChJToAhuBEIVBqdxH7vi9Ak
lOQGsP3VAnyTbySklFkxm3b+mENKuIjqdVPIFnOToef+qX3iHynvVs2nASi7GEQuFSJU++KdaHkK
Q48qKJqNs25iNdfQJY5M211z1+m54v1GbMvNAsgKhhcJoZlcWAkKjZ/l9mm7B3sp+YbLe6etn0hd
TPraY+2090j0FbHovfaDxqlkUDDHJnmWjd+nJB+IZNIi5h8L8wxpz5pUDqHAt15GY0EPaAX49Uvo
TBXF1cxQw1Zl9D33sZ4JkU38fh+j5OqsExUdsE12flOzRZKIw0BhCZ4k7s1zFf7Yo7PeXlhIRw3I
tcdRfYGg3+5AFHjf3+vwhbay7c2n/VOLdylztgB4LNixdwu4Zb66a1c4YZe8T2Hnn41lClKpYh0I
wIbVqjugymcuFSB91yTKyiDXeatNUX+czlZgB3jhksLYSFbzxYdXROG1L96opRK5fXLenSfDTrSm
7jt+AzWmGgCWrickl0yjZuN8sh/qWsu56I/YQDUButBiDJrL4s8uEDe3WR40OCmt32DuhPkY47xJ
Rrxp5q4dcbp4lC9frIkHVjkPGZgvUkgvMUZsmcE6cEKu72Cy2QozTKkURHdF6RoM2Uy8btMbkqOw
DuqAtR7c7/RbAvrxK7w5KUBozMMToR4kaohbyJpA58sMl8KM1GQMRO5ouza/xZ486W/C9T/5a2fd
cGPj4ieGXzo0/bJIUYkX//EzEOyz6F6X1YZRqMpaaTy73x9JRNTWosUyEBadKtCvKSjTy+8o+5UH
NfT4nF7+QkJwkZ+l2ACNLUtxwjVwACmErcCg2gsVhre2aTkoct/zkGx1pFtgsexXh+EnuKYxT7EK
PyzcF41dJGA7W0uA7kNd1LNwrOfVO0DtAOeUU1LSoAXcnh4b/LJ7745t2a1ddwCIvQbP1JqCDAX0
ClyiUZg/5iXSlQqbr9gdCLiKW/n+zjmTOL54LDvZSf+wpXYBTO3xwotut9TtFgEiEkrqLrDrF8B9
Xq+gZfnv4q5p72s7X+3PtUsT7KZx02pm6s9PZUysUH70xna+YaZ+Nh4dfPfIwVA7SNCC9rS38pRW
CFaRATy8lAS6vfuZX1Vm4sWSx8u6oNIU+kAbDzov9bsXBUMWet0yLsXx6N3nxRO+t352xs60a/lO
kqOAx26nigqm1c3+Kx502kynVIII0UclzWBt3t+qn0zMLhX5Jw7fhyyqPFQOb57yS1xQM5YGzY3h
18aBNOYvo3lvXUdoeY1DZ5PorH0sT33e5MAWOQhelQIdr6epITUMrTgWF3wa354p9FQBwpuOoFdJ
BR0jd5INsjlWKJHxiyPUwD7mxflEt1pzgS2sIN3gNC2JlxMe08s3sRQZZlf8SU9JB2Bg72Kfcc/n
jKRGd9rFg93Vq1CCnVTXLvWq0nDlXBOO1AJhE8NXJVK7h2cT4zfrkenzCQDX1Ef6eRnR6U/Sem6+
ZvlxWwt8EcSi0TJgNpZdfUsWRxw7uun0C8mTTqbTOvwlVIzameznsdJ5p2TTFaUQyZg5EmyxOtcw
ZGCetyvjkOLU7Q9k+TY1OA5uaQ==
`protect end_protected
