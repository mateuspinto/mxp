`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
al37gd+7NYpTOfccKnsyCv7cEdXBFDpJ19yVFBG+xBdLE5n8iJisG9CfA0MXRp0gFqWmpEhcYtzP
5N7VLM9qu3FU7mVHg9zIXiL24qiPuV5guB863HeDG+cdydHiyqlMslGncvrjkHRjcI7nn0amKWRi
c1JWslsLS+kqhJfQAmQipFDeQiN30n3c6ZBljdl7l8u8hYIOjXlXincFPwg98lzXiVR+yeZjcdVa
iB14D1d9M7Snp5gd3M0B7Cmp8T2fteH7Po2craNjJ89xD6YAs7Mr0nAkJ8TRtqg+nJ8Kmu2BWw6h
rJctSmzwFXuU238YoRmCP2K5vugJnXtNbn4ftQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="iGiHbfO5+Odkx/0x1Iru5I83vOhoxa3j5ac5DXNZY0s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9456)
`protect data_block
eSHRWHSBa8iZewtWb3z+rt2uFHOHzLXCH4YrxUFW8A5xMivX5QF4520+3MFyhYIcqV+T2MIJ0iAR
LMGi0lmWI2yx13c4zSUXeng8j99UBW+erIjwm5LeIYawIGwmOul8jA/lwcsOISNVGFw9uz/u5RJZ
7vbcdKDlS3E7OeK2BKJa/IbsbTVVOc43Jbz5b98+AEUybc2QrfkB3/gzOI+HWF0rZP17cw1+UIdg
OtThT6RiUb/fdUXI39po0JlgkZkm6ox2RCf9GJeguKENC1Uoe2GoA7h5dMZLE3ZX0yit4tbrWKup
AX6GsTjq5B/zIYQOJqNcy9L6tDttdCt62EYJau/NCCqnO4LomXUBy39lot/xUagEBJigAsk6YIBy
MArKIItyFgY71+RiR+6WkXXvTxjOQPhJC3vUEuZn7BHzspdYrA3xOpIDR/iSq4J7fHeHZFumPtBV
edoP4pMZm7SzSEwedXn+JEPh43x6sVG7VyCdRMFOYwnW+jm+7Uug3vpjGa2phCa3PHVFU8NbHeiw
Y2OA7ow8JiGHGtc49RARakn3LaDXkkroUt3FMaNTvoG7ET+2qKsfjhJDXr8rap/PrOKQWCDr1TSk
zhGNbAFFvhjUOKb02zyZC45plQ8SJopVoCp01+lVJRiPpkfruQfdM8Sp83YqiSEhtzWwGMZylfht
OVu0lKVyVw72FovdWbv8AuzZwvh1H8Lmvnzf+mNqVI0zIZXcw/7u3yP67G88bcejFH3THaYmALNj
S4umEZav+aZwr6hYZERxORqOZFnqWkMXScTBxvDQh3kvKRVYNYLcaGWh3LdzdMQf2U1XLOtDot+M
bXowY77pNf8F9GrTUQQlSssCLlwBO6MNkKZVjXKGNXtziem3FOsi3x0ByHQzcGQjraKXdFOkJOIv
SS7BGHnu+9pNrUHtua1Auvsd/KUkS3M6UjoRmpdbHq7rBCJ/AHR2c5MVIgmqtu8QZkjm6JCzgCf3
b0y60UJLeTKtOQPVwS5mLNG33eotX/sZTsDUksKQOdg559hBN/vIN0s9cjgn1GLksGEyPoq8h4qI
rjeOcdTAwcTMhxQOpg0t3qeUKkh2hbC/qYYjOL7//QuVFaf7BqeRqOcBvmfKfgSSgE/Zv6xk5/1N
Do4xDEY35N8yZT1icxLjcrmsS8dnJLopMDS+/khlIz8rZ3nQZI3Cw6ygUDlwSKU76sPMXeUd2Oc/
AjWeCll+xlxAFszMP8FSHkbjSIzBE4wrpMWIIRJhMgYMPechydwl0xrgCrGFxNYZkjTa5VUd196v
gEYVaS35KywI1Qus4wMvyubAPyzjfay69nIURRlhFL0A8lwd5UAMvU4Gt8VN1XVhp8tUhKBcsJlV
gsmx7r6cohjs5E+rRYTuqEBcAWhUWW49mgqXOKPxcWX98b+HdE9pownqjTByjqUANqh3rzm+6cQk
ReB2XNCNpmjoYQJUyCYkFJhis9JWyDde7nnvFNJwDlWprb5vCA4il9RoL6MjmJtRgHWWFwLIs7Tf
6lEf6NMrtHsP8ZjXcwCVGT98lyvr127Oihy4EAIEHkeQSetw8XppDbA2rCSaBVUln1EkmJdUyXMB
TihF3cadUxG0iGKHQuo1tksbQb5F2JlQZzL2cnA0zIlSYchFgZijZsLXcIakS4ZWlryaPwjEx0og
KefEk9VyRmXHJU0MX+KUXNqFJvSiMENZwjSJQluyRbwPIeI1L3pURAk1k+EKHeN+ZwnNhVClpCIf
W0DF1n7QHszwWHm3ks0Cr3H8TGPOoLyMGYsfGyjEDr0WHzG2twyyIGaWRk9zNEnBuYMoTdWV3EvK
KWZ/cZ+Yjg3OfLQoQJBzDXoIePT9cGWQYh/Fy66A2jC/fmXeRKHAxuFW2ts0uLWEZx1G07Xsm7ul
EUSGtQWT/bbPdGLd+/wWB1IeRheo+hdsnersmF3qkrM3ecLRdEbLVDa0ksUsjKRVFyaW7MoKbC8d
b2FQCCarHwfvz6hZ07bR4hti1ABsSZMwRiwEHwt/iu2DXEaz77r8UZ4jrzI2qFrJA0wSzQ5ciGef
ak1K4AxBABYsqUz8T77wLBjrxncCVPDwZPQqa9y8ohr1xiwqgTJhIFQ8/IUZra1uohgleh85an7b
c23fzKvQkPYUXt+eztlbUqhwLxmSI9UWWfNV03DV5PtMlHFSjxf8QIANu3LJ3PkmpM0iJqBnbsWr
PZ/3z6xpYFn/2NmzuhvVa8CcFyNbGGy68lvllZpHdBFLaVp35fdjdeRlrbSSd6/mG/V+rIaolrcY
O527jGW58XxZUxV/vLCknoupaoN1PdCsX7FrBMnjM5roPo0g9oC8oxqDcFEAdkkJwY/cxRosL2PZ
oT0CNm/+1JdtQrnEKGk+CaB4JJFGXXLDuIeGQhEuq1iyAfM7bhqJnZdLkvFb9ZZdR5/C88BhObMS
AQKczAIm4rrJ5fyM/F6f38FP3ytJzgZw2zYcz6Qjy1ZNjzpnmpFQ4MgzCzhiJ+eGS4m5VOm9QX7m
C5cnHfwMtIvkAjM2SspXzj7Ypr2/1nN5vjwUbh3V+8AAs2DZhPiN0GppXM6zYiCG+4Jk48tbSYcL
thSUG8dWyTqBis++bz+oDtcHCoVS2iVtVn+iZd03XDQttdf0sdp+LyQ2Z8DPxNlaN3bkd/5P8Hhc
tz3NKwx9fvvvHxMy6JXPigWl4PF5gE8U6ZN60cDQGUBDrXeUSfIrwTLdDwYXVshMLWKQ5oztlFBX
7GQWVRgV8q0Jny4MUtbmeNzLEzfj6CD7yT90t3p+d23PCLeh+OSljC6GOeR5h2Osxmpp82C8eWyY
OoW6cabgdtos50zW83GDrM68ct7jl5e2CL+rQ9EiXkaxSVLURwKFfX7bjFPLTPb3kP+2hw0ax4Zl
JBGm7aNlbge6DxMJLJcXm5XonIlSYQKPeNLSOR369c5dHce18syHEx/ZHa0I4C/weJGP7+P/+ibI
GGRzPwWpSjmHT37cgYp51NkmeWxQ5EWRZrpW/3GZ/ezlXARyWqAKsZVr2ZxNT3jQZJqdvvLVG8jq
lAlOX4cWJBGtNcHCRUKBjQtQRptmWN60dgSWQIDbJvQNmZWI8Qhda1ayOFE5Au5BQcaJFp71OwxV
sgM+3++Nm6e737EDs6pmAhSgjNo4c1ghjIQIGXSalpK7OBq/vbyl4CSDdTqId3wTqIXb1lXFB5wU
8XQbQ1jQT3CN0MxgIUN+jvo4SdO993ukkZdHlKMWJ/1NTrjGzevb+X9VYI9At8ZU4bNpdtofBOpE
AvPqXEhvk31DNqTyXqgZhdiX1vMYS/SBo6CgfZD+8t/uySWLIBXcfHxj9jc30r6Seg+BJOYgCrL3
a9Vlc3238w0MmW0f9IITIduHqwhG5ZPlkDclbqSmJydRKpGN9yEd7GR0XU78wtrZavHnwhuhHVdb
T8QLA4g3SCRJnLsK0wtJvBzpxOBm3gD7hae/5HO6TPB549hv7dOg3JQxxDG3KjIlAArCUWVGwCAl
r8L2vLK9+CR6tVtWfvfUVM1SzNXC8TYtftcGfv34aEnpu03+KVMd2Oo8sjb/qr9lB9VZgq1C85h8
I9vP0NCVl3Bnf7nz9f0aTbifQoqwHZU/UVTJz4fZulucxpbyqs2qY3Nu068dyaEbnueKyYxBrFms
gHbfAkomQtxTm9v2/EsgPp3XpGEZZRI/O6Y/hUUoNc6ERXOcWPdEuC8yQ5Jewc4yr1qlamt9MFXa
A9KUEYr6TdtHAfcjZwWlP7VPcbRboYNJPAxzZV84s2FNBTFApjX+ENY1ofwIdZ86eo44SMTT4p8r
cISZnW2eAMthhANWIVT4FDR/udo28bvacifRsHSulwQiIVm6KtnAOwYkEtQCaCOJ0dRTdVdyGtOx
TrNDjn+dH+VoU9Ft1KmdAqpgC07zWyl9QGM5cLMQD+8kM3v+c3Yrvmx8+ZFGNvvB8HoXZtG0DaF6
OwkjkYTeQxFBO0IPmmqeCX9cxQjFW5962hjfgkalqtYeAxCtYWX0iz7bUx6F+/JRkjge27B5bOI2
HSjCoNDfxvCFLDyIaM7q0QF+ZNaHer9a+Y6wkO2uX3sOndHHwPI3TKlmWVcB3dVFG3mZkGjNVP1c
4wUY/hXeWxrwO3RzBy9393+eu46NqfEmb0nFXq0bDxcZpTAcrFq+drYOFt6y9O8KWJ+iywzX7V8I
PmqEwmTYdHcSOXdxZS0A6ASS9Lunx8+aiUET4Sj+auGt8UcPGfM3mUhEPXw8WV3wrZ+tIUvlXsf0
qk+jM+MoSAbboaX7oCO8REaqDtiDsJhyfD+sig/7xj0b/qhh91nWivxIRgFXlat9d+n9fUt6hF8E
oS1rjqi3KqSNJZU1iqogR3I1T6yejsNsOZcVTCuWiCHFWLcrSPUqYrLWCpneWSuAteAEd+of89LF
HtqsAoVEMU7QZN2Eeolad1kvRjWis5yOLc1r7Q9xPal2a14qyI8X4viTjSArzxgMpi/E5XY1qB+o
EujknQ6MLN9aTwhX1+bZyWax5/ktJM/ZsfmTcgignVzD2BIK9PJ689ZwpUcuLfutgFxDWBvaeKrg
BahEOZ8T/UQ3NduL4KYPci6D1shrSiBKNC3IVtHipoSawnGaHh2ATt9Pfb4zPa8YKOqaxZIFvaaI
7jBxGaJ57dUaXJR/KLuly2g1vA4qG9B0lvQUhpZ7dZjjsi00P6zXjFJWbr+CXOMyXdsQsOfRLtVx
zJLDbS8mcMhjdASbcuWXjgCUVimML1LYiGK3IZoDA9UoOrybg8eS1YA9PFrrc+nf0Un6ldEse839
qAqzvcXa4C3eNfmwHYkr4TlBlGbH62oHnxs2NBxSbofeLp+bFbndAepBedn4Y6/+jiH1wd8Lbol0
VLJpE/ff8GmFEMRyvsCU5Zm63zZAxtkfTqIKdIOCB3YhP/fdY1lo+bz0hi4ycRWNCyT5i5RZfUA9
m9xlwBz66ZxVaRp5ekvL0s0a0o11zNs8ia88lYXlSrlKNAfXDSwYxeA65wjiUydbkDFQWZ/y6+2R
l9mEySXJU+bgpsoXNDniVrjPZuDOIJPdkMCVj4LQPcPhoIo4MFahDVXa30hNserxQZsTppwFHUpg
kzz5G/c+45+sGA13yRE9BuLlbABfSPOkEuLbMAGaK5KF9FKlDI7vZoJjlpH+J+hR5Jl9TQ9VX5t6
si4tGi1Vtin+nOK5vry6L+m/9+KLY4sbUtdIf1K883nvphF5JF6OkEl5shjUjUTQkAl5+RavR3/Q
OCAH8u75VKPH4jyhAa/jFCfQZiXorj9OL9AgMHZ7fsq4bV0/Qb/yYGZHJkBYBTFqh2Cldw+S6f6S
eyyCLv5vMt1vMy2KZeWlSHXTl5s6GJHgZPu7IMRunMpp8rsn+gYnQngoGEbaOF+kqRewRgHhf3AC
EcSmEX9y8S4q2QNO/hcpqAO7OILRZn6YIivsGi9wdDp6PTOL21qyOmQHNKkfsab9OK4eDL7U5Hge
0hAHn42sRErzbewV1qfJwpNno74Zw+0NjCu63cRu1W9bjlN3gkt3dX/RMUt1IHUVt6GLaXfiew3T
lqnRgEQkYCxPvJtW78b5NyzKtyYIJ2DSucIEaAAuydIR05yh6sCcdQEho2b4u13r3QAshxTO2C/N
NaWNzM51wvUh36rp988Pe6jt+f3KEm0d9vc5kOR1TS+2dmbKUF9qipiM5z9ODVaJXDiLfs6EkfHm
sJ6mZw0IY3awqLfnBRAgU4eNN/16Bj5w8/Yc/PExGPhm9jB0jivVFPru0F67nXfpJW1JN4dg9c2p
nJ7FAE3KrF6Tihg7u7rQKY2P4VZ7rWVdXfDQcFiGxBWYwXsxpCbVGX66ye+ZAbILL/g9SHuU8VKi
9GQ/upSOE67Y/wxs7dt4hqDYTKDYGsGBdwV9jR1nBY4ykjnN/rNipSNlyuV7Pl7RsV1ZWvCrOGmT
O2rf1iQJyFhB86T4jfzmfKyHjqeVyK0+RD5M6T/uKKDqpWax0u8xNdr3YZ5tKshQUVTsaA2siDty
tFcJvOs8aMErgFzxomaX4wzHK9VqkxLWbEwvW3hUPpgJrdCvJIj6ZTYR8bWvvufgONW2qfXz7Ax/
bn6uAy/48dPB20BqTxnnEl417PB0C8xgxMkswWkBCPwWmXNsKYkyZ+74I1v2IQfKI4U3bDsr2hQp
JfDFABi8j05SP8MAeha7nDpkR5wNwqeEyIEUubvpFn9DHsxhum0Zewk7i+7+P+R8po8tXtf2L0Uu
HK1RR6zIif5LILmJHcI6+JAU6k1EJuLnAPjbwaBbBnVWRVgddeHRCcTQF7MzA2fB5Qqy88vFEYxq
mW1gRv5CVkg3ICxHaD3/F5njUmg9US5bDgqZh3JGhTa8viLN6a27KeEA0xafizgyRFuz/sV09Qv0
G2RMoDdc8mELI8ButPoIMM0VHAry9oSb7UZp5QPDlBw5eIeRDe062b1cc1rbJRrhECQ5YdYBk02x
z/3nKihX1ddIKO1gq7lU8cAn4XZ0ZPpKXnVIZJ21zi8gASZVP4D8cxwZCiTBfA8Ab6YxdpkOwZOS
bmpVoK3pYu9RYk8/MUkRMEswW9ksNppn5YR3Rz0ClIxpDRkL/OATwoiNXsMlfL2p28aX28u1X1te
WCRi6mwkO0yqmwpKzRUIWHJCMjm8KKP1WeoknrjCrCHwDtbxoobUQoJ5jA5hV3NQ5h0KlkVgxJNl
5a1TGnazjuoeDhjcvWYRzBXtpHqdvE6WdYmeT1/lHCW+6iwn1EhTRdwtoiBktfW8NO+6rX/4GNIz
TzYvZ6Ffhy+ZA1BIPpE4jx92ZayvtUuq2epbwAGYoOT39/MUktNl0K6PRKauhnCSuMZg8vuwWw/V
2q68VJVCZFdWxKjLXjW1RC9ZE5yoCGCBM4A0vG5PnmF+IQs47g4x2vGjpgK1DkOmiNLAW37RV+8f
aApmyVRbFIvtC6jw1v5buftQBlTK0E4GW2JJ0/ak5FVuhFWLmX6Padak8LvRopwfoxP7E3UyROxa
QmShrlhnQadclUbhYaCPZFJz1TRxUwyY8j6B1a8JfM02o3lWmFPycbMmDZvnEUmbsKrf8WYT5kQM
dkwPrLfdMjoZvL1Bhm43TARYouvEwjB2zxeOmQmZx1jtjWFElM2u8D7+GfQ6MlWjj26FhaX37XxG
Kvf+2w7uYwUHyMNkQWxoNaroNN6sYupywyBDtCjxkbiM6X8BgQ8ZZMvTqJE+VoyKQfMhbYDVNPC9
wyDbCrQ1IjUrJRPCQhGF6EDelAmG/d1iZJyIWActqeWTslgMFasNgGGLH+G4pwhyoH8bHQHV9DyH
fNfJEQetRjdssqf7ZDV08zQpeQljh5m3I/vOW9yE8X5XtgXlhPz7iX4M9ITKiULqQVzwWABaOguk
ph+xCclF0mdLQ9ftX13yfUQ3S1KsYfiDd8REtZPgBkPcfDuMn+P4qg/l2p5VewKAtMSiJ/qdA6pQ
YbBNfFsg5nxOXBFYPhJOHDXYIGas3IhUTmdImm27Wv0V/JGj6V04/rADg2mLLUyWHCGsftkbcRg1
MfuMwoYlItttKZAmf+iylutiyO5iXJgX5299t9PfjVjfN9RQB6vc5W4BxomWyl6Gyhti+vbn87I2
Iy4GWVws4ZLfv7f0VZTyAoVOKqMmID+CvacbTkb1K4isW8F0x8oMrBXK+2oK0XyfaC2sAhmwgIbZ
hAAWlM8l9H3agT2zEMgtJtJnSrymOzcxqrsiW+nwEZktTWyM4Y/3jNmaDIlLJeydrT/7ESto9yqc
lkBhxFcbroWE1lUGbeKMXicDk8+/HgRhls1qJQSSc1nKLVg5X+ewy2oqdSxoQ9+xTbj34jL3T21w
YC36hDD8/7hyG4XDerzMAcxhauxug+o9L8e7NVgoWxEK3tO2H2GjfhoOv1KVOImwyVWuIOhcRZWk
WvMPodDR640wvsQ+GUjLphC2HqdWMMRYNfz2UElvukL8w1TgWcsmI2G6dBn/diuFhoP7+PS2nRym
Whz79h/DMAYRiVg6SsMApqU7C3WDrv5ymxHemEXQ3QlHHhk3Psij+4gSirnockp9sMcjKLnHClqS
UfmdS82K8RHzCiUh/LPyO4niBNU7h8ESIOO97AdVFhONojggzD0+8+wWIaKcXB2JYpnJgJgJ4Zcw
9lOnSsXTSv7FeGlM4qm2tLAcyzul+vIyNS3o2MM+t9+3kkYGYaRzCz7k9KmAcwasxX2qYlfdiAua
AzjV5fd4t4T5bZn3MpZPYogTcbDnq9e7TsTjZZjKvWX9EohleXnLgAkdjw0XbRK3rPiUV+yWMK81
6Y39eC2YiCHhdaHo2ALbqIoDlypidHDeUGaJOW4bvO5OAlMddvrof6VSeUW1W5yIMW6oPQKK0Dm/
796wPkDDGr/U5bmu3iQz2k5xlXkS40t7WJOHP7J+Avdgz8/NSEis7J5NbP3o9QdokCMuEY6AbsuR
BwtyKDaGJlQIf4D4at6oTIuM/YjDKP44RjSXy1xJRLPjogAZJ2B4Gkxj+u97NBQPIHrhhtedMSH+
AYVDHgzh/RjfqyTcl6f+PEiuh/bXUX6kgaGWFkghpoEcA+EHiItxKHBAKwpmUrP7j6SKBCkN0JoW
EMLmpS+J8/RqGornRnkzbEOkeL02ly/f5DyjsNJQ8XYJpBBUsJPhpJdKKc1af/llb28pZRKnjGhR
HP90D1sdk7fPC/t3anpmk0Fm8RyVLPfFwNy7w32mPS8hwPL/SVHzp8KOgWIEEe9ZklZaaYZwUDdq
NynvmMWTH03cd9q1z19jkNYo0G8FWMYnR44LORnZ+nJdQjyY0E54ojlOAhhip3Mf+W2FSnG2/l7q
N2sO/315KPUdkr1sx9tDJycbGUNdgorGlb4PR3i7zxOaIAsQ0Iq5oY6nQJSSwxsR706xRu51iEHs
LqNwYR1bIz35inhosAeUb9xILBYX2pvDGLyALE+6JuL/OON666HctyWtPVRt4MIRURNY9YSX8r19
REfXv8vX7fTly2wTnz44KRIeHXueQQ9SaU4oNTb4dmTd1/zf2nLnDHMK10DJZXnmm1oHUUwdO08Z
8MsBPoUvWFdG8zFvdcMtgduiSWIQFrB/PQR1oR0Unj0tAS6aX9iyCP28aZ/Y32n6+HeKcwaor0qn
Yd5+H9fRlkN7+HrjGgDTWUarkpxjq4p9UYQxc9TF8giGgk9IrxpfMsVkwDk4VEJ7SO6RA9XeW+MK
PYsaT78dXjmWTWBG7DL0PwtecSf67u5Ox5AYwtvUTT7dwmAWu1bisLsbwW4kAtZ5QZJkQ7B5B8wF
CEgFAEHLh0oRAsgXS3+pIlMCPBCo+0gGBQKUA0ltGMkErJPvQp1OJFkD2+VoYPZybhlxzgY0RcJC
TY4ObwTI2duKo9evYzWR7Rzi67Vcw9/OetGmlpaDWwOm6vdT7CJnWHCZZe1WAWxu0GJ7rfJmkdYB
RFoyCGXB8kXvr2pidcg59xlUawSxHSClzRsWkJ0H2h+9zyeNEDeoMWioKGUwwt1V+F9vxJ4YuosH
iu77qkMfZBQBX100nxtPSO9NQv4hMzmOftfL1iWSZ0emF6H97no0HFz7tHlebOUYX6Dg7fmvxiIc
cUruZIunEIZ0hFqu2UOgsb8PHI2TZ8M+Scfi6Yaovl24gwSg0PWzVR/i+aJFR0bQzihEGaVJJEkE
0sXSLSltL5/wa6/d9jVfBK8ZfpUTxLR2vshb/mYnh1Vn10z52+w/xP8So37ayqGGBmBr1uS99F23
g7nYC7u+PzwrqWLULPmJrkdIFn4u7qTIvBpUdRy1g068m3EZpHoTxQhQaXNOFKPBM3EeHleIhxlk
D3o+fm2ScbIyVSRSMT5yWYUuRntM5xPX1LeDQRvTP5t5dV8rGJwyIQ0l9pXWeG8Tm53wIfh1SSBa
+yfhubtC+DkSilTqqyJI0tE4bbNcwe59+xJ6zzB5cH8mZeUa5FkUU5j46mz/QvuriDObZKIVtxux
JZaLY/Is7RuE6DlPwx7qlwlonRhFYKCC61cuCPEfl0QVSgBFUFryRaDt1yHQ2gy39MXCjIO52upP
8ENpVFzL1baVJEKAE83kHQd7P/ZKqtXhQqlMlY+hMzlV7pKO0qKyEyJSvfVJhijDlhFDaYW6ZLiX
4stpQ89p9m1qWwWIm12hUddbr8QvfGOsA1HjJRbwHs4pdY1y1cbUDkX+frrysuvutN6neGh7vggS
qtfgirS8s9vVhp6EgGXa5qm/VkjEhGindWXDercZs9RU8WS2/PQSL316MtSApLgkkWlw3W+eVDVz
x2IWPJjkEpX+HG3cJzCINqYlQmD3cjDji2rTb33qKzxdxs/eY8dB9qsyKaoEgV+bSujTKuejXyKB
px8L9ZijugzFl5LTL8TtY0Pn/aaGlpiN7BzDrpwS/Xzl3EKKN45VXSTOEPAD02X0L04flRBbiaO8
fMM3a89tEaZFEM0cOEme8gA9YoqfFR2v7B4bn+rg949UgKLGZ9eMnZvZdHoNtIj+2Z3w8s1u6y4L
DL1BDU77Ou84GkwGpH5bGMDPF3u80aXuXkqjqLIN9sUVdRJKTztPtlKTrdNhtCLffHJ6B4iR2tVF
ktW5C5NUQR3VFevVOq+sm/7WQor4JJRAwZZMlFwKZe5pNS8+7ZS0T2TpPp1+RJYRX+1fRw3ZEScv
F6fwW8qCKtq30kSyNUTVU30vaAh5i4QXQB4/LAh/0H86MGrw1ukV8KoUyIMN5eRkv8qprQSgbdHc
RKvwcOK3J4Yh4AFS7MRbeppXu4AuxlE5X7A8N/yAW5aW9dkxPaCSVs4hyBmVFpPvklrINj4cCl3y
35B4hxh8FxfbZnPUn1I7m0sm9QpUmaXUAtdu8kYlR58xqNq0bmk3t9QFhkAC5CadMBTtZpEoZVDG
Enk/h33riksKPDZvGWVUAelV2zPY658LEnAQnLoOqPc33ejWN4Luh2n5Yln9q+/CV9d/qthN1s46
cm+qXIG8clzCRq8UI/+YABbqnPfeRQEvcnx6L8CX3sp5icOBYmqz8WtxpEpDWC5uZpGFYDsiPQcy
uoqmyDOnqBCsS/QV4i8M83UI5kYi8MGKRHnb2AqIiqHLya1r0HbApK+74Ht54oj0o2so9H8h7Pen
VskuiVQgjF/xUFc/6SUXn0rObsKvH8zZCg69frvtvL9s0SpAvIRC+486ds6sMSq2XTzPB/HsqWed
j/No+zJ3y87uN5gVNC6lH/n1eCVf2Wd8BNeXA59Usz4E3EHzsosLCWneyQgmzQmqAvvS/7Tkljke
99UGUy2HqMBnEuICRDIEoS5jk1q3CUDnlinmGGuNO6osgyMOhE8Bj1r2Fxst2vLgr6e4zqpyKmxG
nJGtn7nFtY5QvrMtckZjF1YqFmItfBQhfr7mHrndm9eqzuqpFkQXscJr8STJ0+HJXQZ98EGcT3yY
Bk98Snx+k1pZmqvYRovOV6cYdbDcfhWtzbRw4/6u9E9M8LR8t/v5T1zpYw8gMaHKrZE+A1jE10zm
HBBPcnbVbBy+YOm0D3s08NoAVETFOTybHav2oVdeLNE0xqcPoca+ZGEpj/kzlOUN3wO2lsu1kbkG
pWs6TYamHNwHlFrDRJPkRmUbslZWQPx71Ff7D/59ag06TkJs2elaxyVkYa2to1gHNXUbifml4Dc2
hQK+t98FU1Syf7z6uieNmMJ+mHnYZmR1UbvMVW3mt+BSGAieemY/UsOEuNcrJ+xq+V8SHCBzTIsJ
K2rYIrbPc+0mVZQVXE6Bh5BlDAM9jeSS7eXW0Hmpjk/qmAolF4RTStMfbGYnylvfRKNtYRVHzfID
IeYr07yI6L0zaW1MzgXU4r5UKvUXHigCJvMywa9Kx9QFr9JbH1F/zG/KrH2MajeWc6IEuSLX87Jy
GEa0HwiL2ih49dPEgg50GFlZywI4bnM2NFC2xHP3GOxbS6fxDUczYy5BuK8Vmpt1VXjHKLyALkyv
4H1DKy50VzTnBKIcYVpQbRJe7zjRzVXQqMKIXzSmCSYOe4+/+yFf7GfYY8LeOEozFmtMS4u70kJX
GFifV5tRBM24VMT9YkkRG3++2O/QpAFCocDBEuj4XZdvybNU+FYXaMAZstAL5gqHAWUtkiEBsMIv
6x7Wo4bUgB56NnJ6YUYAXszBhqdXrp6DGpjbWUcwPWmch5+VsaQDCK9R8Wv0og1kiujZKWqTEJLc
pMuoU9os+d3B7tTAWkK39TNMqPdcvy0jqhx8/pG9BfK9SpSbg5uUKO2nLxWFjImV66F8c9wYbXmN
r/0hxctaomhgvUCvPBq5QofqzG3UzSTwfPrX3CFa+AW3PXPSuJiC+TaxvKFIdhiFqcnkAje9m+vH
VyLA+PvDzT1/IzjVSUr0h9mBbVOC83/wvdS5hteGDcA3Ij+CU1QkF1RMoKxerj5BzgKF8st3U33N
8zws5wJK4Pgmef4RgM+DzkL/gvyFd8ydpaByw7oNvwbRumTfOQhX+ekyvO+ml846s7xbR9BNZNnU
GGTXZ8J6gXVXRXJ7WONTHvSiUQjIYvtX6Ryu4R90bpkVa21CsQXUwwC5FRlka8dYxQ9QYJJYW/5z
ZuC/P1QF3fvtjXfm0XuQQxyFpch3m/BMKhyBIQdnS9ZU7yGr0fB7dyYUqgDl9Ijg/HeH
`protect end_protected
