`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
SVYe9dgEEQx1meAfjZzarciuksM53aOg1ksiD7a1IwqRo9sSs602Z5FaMhDJSFIwq883otsHt3im
IDsKKiu02bp91cR4MsC29CbjYitqiHYTrdf0gFEaq7xMxdnZVvF4chhNvuEwua+Gon/t/7I+m8Hs
ut9KaCxCMhm2YqYCCkQPhQ+OV0aUxINtnrRI6qC03h0W42DAn5YgjeDO1dczSpZoVZrFqAFQ+OO4
XjdQSV0RwNgjNrtk3TSIOG/ZsHkCe10kQQtDSVNUSIwUKDNYx4DcMlY4Cg6mhG11TVRUzY/iuMla
WOFNN/7G2oZ//LUrLT5vbk9YFkGu4ryRMA3vzKULT5A75i3JaNYj2WdrwePmXldeK64Fdu9ZzyrC
fMbhPx0Yf+VDrCpJ+PiWbkX4JYmlgAOZ8YpUTfOkR0Mui4EEtiZUb2Mnv7F51pnGmhcOIDEMnlo5
SApeAczs8xKDG0ezcpscT5+EpCCWnMocgAja6vEhpycvOeYu8+yp81AWekHYG9daZ0S7yG1ZMMtG
Vw3ds8jZvCtjhDoz2xL9k6P3GU1J4Occzf2bpX1GajvBwX7pwU75NS45SuBpl8JBrSoWyNiSsltv
DI8oCWKjovTxLEBbVN2IWZuZvf5t5n0iJ2nlfEOG5+Dac76GLJ+nhL+FziOlAwJPbd2PfF/meIdu
K9fPgmjS7/DzFiNjmFK+I5WPQh2Cs+IADOLU/syrxPFuqnzXK25iXr1KPbu6nV37UtqWz2qeNKL2
sB02aY2wEFYyB50VfPUkqs/VvOb38x96ja79G+IA7ZTpjyaNroX8LpFI+3pLIrtbzvVKvS++FDeo
MalNmaw8tejZqWv9kiUkLii6MAS/RWgsMvBA7oG9owWZnP7Cy9TJvueJSr4OQnKOzz6ONHbrHUyi
1F4Q/J6Pi5bkAlJ8Z022erShsB2kobRsokRK/e7cnT1kSzVa2S4VNwrklMWtAxEEFzhJo/g9xpAX
e0/igxtP1WWrV4qUj7nX5k5YhpYNTEsGjpEuBBMlQLXZ3Sd0U+QELmxMWXmcdmh/P6GNT6+1GWEC
z9Pej0TzHsJ3RYE8fbzf4ufcvzYE2CRSlmyl1JWOMd/di7mtUXlpfIkkTUTen1pbqoPlK8ELNK2g
/kBl4rMIu4I/ma7gGJ5zUYQ9ftTLf3Xg5iP66m6RJrZafgg9ajrtEqOUS19qImvRxNnDnSNCitUk
ahpbtadeOKkH6AvFgmYiu2vB1yoAQKf1cPMSYn5buRovvKU9EnF4K5mxo5N0vPHwKK5YdpN4ttzD
0MF7hLY5SAoTiaCm1nnASkPOOczDO8RjEm+q5q1i0kTg1ouv83aiiiB5kQT9TaJfvQhBEUYztgYd
JMq7j8TxpGyEl3jnPiNykirq9NKcJpP8DXb9i1eeU1X7rgkPukY8z2YemNqmWwoBvw0ns5rG9DE0
Cqv552h7b3dfAhYiHtsJxWAfXjWMM2VDj8HM315xJgwOoUHuutCp/rEsyZ9E8Tt4Gdfdgl8frq28
29RDrTZD0748DFYhjil43DI2qBpUQtVBYcyJW1TnE7Us4jYRKTNXgtnDoT/duZcnvYR9P3/2SZAy
MFI3YRpmhf54cIfjTAjJUo1KDXdc0P9u9voIvCzgGXXPYRiCS1kI6nMCjaKHXr70LseFYO7SU0yV
SZwRGY8jiNh9ZM7qTaksy7hnz0hIL4hLI8Cf0LV7liWRXOy9p3CO3LEPg+FjQftz+ANDqbQz2UBe
tk9+11HFFRvXgujv6XC1ANnFR93NmaNlJcGFmjTxmh2FfoHxViFiBlAhSKsDbf3c6FgE7uQFWDSN
kCa42rjv1gYI+sCtWBogwmwW1bRvxNIGOj/guKx2MMZ5jXptA8JIH6IAXrXfWrb0hc4m87hm6QaE
C25huYF/VtjgdWQV3lT5sAtwQYZ282wye0m9uso4gp8jo3f+DDP5KnaydNer+ScKiNGVe9d2wx8Y
71ksRUWYRt7USAEZOFPfUBaaIvq9Y7m7uJGhq4PE8Vqjo5n/htC2czXdG9GZmKz3rO7h34p8Q4V3
S1ajt87WKy0k9rxeolYZ0xt8HEpPoK+4o3x+3HJtWJeUaV3cSYfp8bszJsTuIawJfvFqGjKpIMLJ
az/S3xgx068eIr4VcP9L+OUw/PQnc+0qSoanoHnAsyLjukgpF6Ub+DQ9I68aPAOKTnMSpLqK6+Ps
oeyRay1zoIg0FLbA1V304Gmufmh6RrgtnW3nKAkvg+wKQGTMFrwjheHAmf/Q5NqB5mNZ+ZQniDsA
7NxsZtSXOBiPdkfoex/YGqunFTPpP4Ory4O/DVQSxUE+UXaLPYrwt2Ro7qfbn+8TwxTYCKMO0uQq
pGYVIEgV/oSasTPdimr5pHLCZyxXD1llPzlb8f8s1V1PWPAf30HPCQzzsyDkMqrKM7tHekOihZ9S
j42xYViV5Z5qbEC0RWcJ7wM4t6IDI6Ytzt7VxlWv7b9L1mme6g8Y6HhIGryweeD+9gYsnXFHnyNc
DeU+ee/bEcNC02AKFFhWBv22Tij4BirQQimooJUNBDHO0IoYPzDnzpSXCiZnvvEcOTxWaG8F0K05
iyMNyl9nTSL1O0yAOMu1VU7Lrzx61/jlOHLF57dUvJpqv+WgJbwuBdQnxT6PTuvuW6h0LfKPH21v
0uW3theCjwfbRjR+0VBoW4UGjIcCiGvW9DyVA1GTa/1lX8+jXpWaU6UvkhFlpE0wgAB4fdYI+IhK
NtYi4eB0JJpV8bU7PcXpekHawxNJDFLsvbr+ZfJ+GKMAjSupAOjevpU4NIDIBkZW9HRsl/kuSY2T
kGDhinwav2kegJjjPdLXZuNA4H2PXMXscZxcHmPST3th9XhbVn5nt1iKJdo2HmapiV9vTaREMEeU
qjERLKWt9LVRGZfIpjIMVyqXddDvMcilAlAuWpeSeRRsptci2K0OME+vs8CNvKraumf4WSe5yj1w
RZns+n5KR1LaE4ehP4Xj2hXqnNOdeq1eKCjBKQDbzuke3NXYiFdBj9Hbuuw6g1t5SsZAObtlKDMd
8kdkgXMjEVy+luVsEY5gVYQfrNv102i2pLBxPO2vXjqkk4PtvUyqJZs711GZk41oUTmBxDx2fS1a
/xGlp3EmMO28UcbKIWIdetza+5ef/vmoXXl4dnA65c2d9swIJ8V4IVPv05GuYjIkB+dU53AU32Yl
KN4TT6FwZBjPalmc8vavzKNc8IWoRHF7Ua8P7Thjm2nTBu0jsUwJz3VccKEiowylIAnYitoBJy/M
PCWBuvNdOb89zwIO480kdvDyCiKQEuqty152fMK6iv0bPqm2OgJgjBvlfY5tc5Wogmw74h1M6WFC
ULvEWadQrE7tpfnS6Uef+5aNApiM6u+qBMyeQwlqxoSUmf2o/Yj7X6GGAoc//JWo7SfFSU/s4fEK
GnU5w/LQs7NIQmLIfG5f5SQNCthyEQW48I7Az7ynn/C3HbLmybEl7AbG74jQjUwQ97gZAGqCTjcV
oPfBEhAu/TV+7zd4ANsY94rXpP1rDwAFpKbt0nOGk4lD4bbQ9eG8Kl3BjAEZ4ubCLR64F1CAIm0d
MouDA4/fsCY+Gk6Ki+4Id19si11lAfjw0znEVhSHXp7FR5W2xIXKzRr3tp27HrkDLZ0d98S0k0uQ
hJc1z9nExPVvzoBRTPKzooQehPBQZ/rjqxYiTFuzsn+mrt1rqojn2eqPf/0xJwCmTv4dOpcUiGRu
rFa1MFiEGRJ31T6xY/ayuv2G87zBsvyT9XGMdu1twPZx0CYsLV+vxHijkg2MEisvWCuq/Y1aD2aU
KTB89IPvZy4ltGxlDK6TH0bX7nyNLCFuOJX3daL7HdVy4ptJ/xnMGU+qxGgHAi6KgdnnTOnbtVpX
fAf58qUI+tZu80TZweU/7jWxiH6fGwrvbkIiXyaqvXaG+KEs38uRerX9LPdxRVf6cRYj2gUSxsh5
4vl58PQAXt9NGkno5UkpKJAnUaW0h33fWOZUq85gpcyFyJjAia/8NZf0EKMU+oXz5WPKN7fUx2Uz
7y08Q7O1GO/kImLpQodDdEhHCBdcYWyEj95LS7I9NbaFlGDaZO3PvwRo8O0/nBmJfSlNy4cskoEI
AsQA7a7oQzmr7RxD/wE/XECjw3stCCY2V79896jAasArtMCG4kNSsSOFFi/TDQFXxzShx8PKThpq
tpZbqT3O2nHzAEfEa5U5WUgwVL/sQI/2JfmerZKv0buNM/HPHeSSVn8qLPVwOJVfmGVFFwM95eCB
f7k1OQLJcd76OFcET0EcNrLpY3P6/UhzLrZ5MEdzHiPUrQaToG5Q4c0UUzH3//No+ZtzYYmf7G7U
gmIkjViqgHl+EMpF4Ybwvjp3CEIoyO94ZgB+NCK0Gwa0Y3LahKOYtXmBtFD6aNmZ/K8TMcoxFAFQ
MfLSUauPjIIr1f26jtCwh6qWx3Ce8BlvO6zaX9hS1KleRHeiaDOCGsgvp8KyUC3FVjA/a4uY7gg3
nt8yot85d/fuzGeCbEuiia+vjiGJnvtky1licOHIchF3tx9MckOXDiJ/aMhH0Y8KofzNsvwkDpKV
obEMnlk666UN0oJ10l/QFklnQP6llCQq9teNmbQ7nvBLbd0S4pbMZGQxEFpxrrMwyxNvBraGPBxL
CjK7MUZ90K9w0hGWPu+4tKILiX332X/7j7jKrvc4nXotmlkRiZlm3OFhUf9q7MIaLIbTwW6JGvhj
kIX7OEHlNjEYHrU1o14pSIrc4LOXyq4owZYlcK1ZTIlPUf/M/PTPEgP4g8tIXmhUauLbVrBfCIZH
NmbTliq4jKvFjnk5GMxbBbt0lN972HipmVGDVPzm1IGEtBcM9bGVBrC1Cr1OmpBKLz2u3jsgO2fc
25Y9arqS/fxtXrkv/xGttA==
`protect end_protected
