XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	���^�)ZyMU�|PA�~�����*�;=���۠l
���7�K�UF��:	�v�+_Q_Uyyԥ����GCO
����γN߽���$g(�{���	�#,�U��G�V�n��py�R�Y�W�����z�,���o 5:��x�������A�F�1�:+��t?��6>1����{�I�E�Y�q���y"��j�v��m:��2��y��ͼ߿���N���ߙ�����:�Yz���V��&V���`�Up�)����{2��~��BCG���z�CC�<�]��}q��I}���Dn��OP��_���2�d6�Qܨ̫.�^e5f�'��ܻ��݂�ދ�b�U]������=�P�d���"�I�->lr3���-�be�$3��C+�3��X[s��i��H^)D�쥨\�v� H�R�%F�SÜ�A;�~V�N������R祷�/H��i�����-?���?-�+��xaDz�,��i�R���:^7X�L��X7F�j�\�uw���:`��ߝ�� `0@1��f�v?U�I�ԝ�a���S��Gzӌ'˺A��x1��E����^���k���|��M��Q��@�w8g�l��k��2�[c��q�2E�m�Ľs����H�9ɶ�ڜ{�KU������t	W�?��2��rL��ҽk�G��)N_�ӥ���z_!DԐQ:�w�$�w�MP���:���f^(�C������|q$8��ۃ���2�}f8p��"���������XlxVHYEB     400     1a0`�'Y�������_;f�+䝡�3#��8��wvO�I	F�����y���Ome���/
�φ���q:[�h/r���Aq$� �G@����q洁������ُ��r�!��>P�~�.��UT)�ga�p6Е�Y��&��	)L��0Si����W��j}G�ć�x�e�n��{�ܮ�L�h�˔���?zX�0����?����J�u�!�Lj��Q>�4���@�<�v�`��(�Vj�=���A���L��Yk��1phu��������X�FHbᤸD�s��>��U�S�+�E 熺�{j��7�O �Dg�)̭̖i88=�l�iO�d�CN����K�RA���߳�G}��60���ybP3}��v�fd&�s'T,���P�2��K�X*Pך�DGg��B��XlxVHYEB     400     150Xis�h껪14i�\�]g ����N/T1;���z@H/�K��/��F��Pz@����i�؟�����q���ﭨ��_�;��\�M�]���o#�m��N��r��Z������Ll�_؂�@�nC�H[��
z.ר2��黣��,G6�	�(�(�Xاm���6�;M3�V�(�,���͞:$��m=�oAA,k:ؚ-R��w�f}b��}*�zg�2���PM�W9�i"m��8P��X�Fq;F{���چ���Q�d�p�q1����2T�{��w,���{n+�/**^�Z��~9���t%����x[��=��`�@4��әXlxVHYEB     400     190S��r۝
H� "��"��S�r��<���H�Q��`�\܀���)����q=��x�J(������%�qP�c'�F���x;�PQl����؁I ��9��a���Ə�DQq$4c�'6B�u��Q�#��.4čK�z�-<,�o�g�o��5R��-�SQ�9vB��M�Y �8�V��.��������ʥ��K�}���З����ڼN�3>�'�����OG�`"i���(`���*�>��})D�3M)�)�Ht��d�^���S?,�̟z�m0d@e}�a�t0�f�G���^����4�%a�B1͜I�#�!�V�����(98!u��6�-\~��kaI.�׀���cA̠;l7(��>�nݹM�)�ի���CHndd�XlxVHYEB     400      f0��c���Ɛ#<1ɮ"�[N��۰OA��DC�=�U$�O���L j�����Vb$��g�[�=f��֍ KXr�^�H;�S�2:�wZ��Õ�hHʭ�v�<�o�&8���@����2��F���b�&�L����t�P���E����q�~�2S� �D[�hnEx��Կ|��daB��@��ҵR�����6J(�}���7�/�m;�uB��n5Ď�K7�oRP�[��'�Ό�΋XXlxVHYEB     400     120� (�J+2F��:���n/�fK83jZ���^Ǭ>.5M3f*��y����Jq���u��gAK�4�����Oި�:I�9z{B��*�"�ҋu�+�J����vktF$2�Y8��p����D_m��[**y��G�-#�u#�8��C[���1z�5X��kd|�	Zs��tS »�b~n&fz z�κi�fn�Lv�����o]!s�l*v.��N3����5��]K�S��Gi5��B'�����V����.�C澿S�9���0Py�F�S��a�XlxVHYEB     400     150xc��E�B�����%���R�4FM��0^^!���:���[DKCj����tGt{�lD냆� ��C��K�uk�R���`�� +�-W��l�!|�Z:��R�Δ��"�h�����`���L	/�/
����H"7eY4��V������
�($Ё�a���F�N�[������-|��l]Ο4���Gƴ&�.ypF�a�MQ��y��Ҍ�<��7�{}	*���RѝC�	>�u1c����� o-N�n�0�E�]Ų�z�c}o�5p����rg�c��|�K�Oqoj��y�Va��7v��>+��*�쪙��т��Ĭ�Y�U�>�XlxVHYEB      ee      70D�����}6�w ڂ�h�	ŷ}Q��N p��x���)������uq�oӕ}Lw@�t��d)}������K`h0@�L��K�e��,���^&��8��t���~0�.�