`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
+gBWueQtcbqr5TRi/RbnvQC7oI+jU+iQe5Q1bgJkhIePbcVKfqVjVetwGuz0knq9My9ahD85yQkM
blwTfWhn2qw36H24AX0Mb1yqMKfDFfHCEkNeyMo/w3OO3COCq0iR/tkLGPA7BaFuPGnAFz/cRA8+
Av7q+1BNL2gNdLrznpyOt5pyrf9vpBr04IuiCE/eqozuI6M8kyncOZKXYytt8LNfpRz+kYAE+acv
71VC0vYfkfJxaYTkZVlLEgSOoM/hvsTSkQ0UOAvNG6NmMWNtt0782Q3SyXdy+hfFrTer0/UUrvy7
71imBwNNUvkhnmbL8eE8ZgDbm1QrBqmM6rlSrWxgJ1NK89qPtsK69j73XPWNdbEadpUldztRAyRn
TorLNMC4NjS6YPKn5QxaW//Dgv9xRKjECuHx6TqXcm0GXisQfo8X8i+fgF9oRO7ukXcw49CQ/ReA
9PcrLH2qZcPIvq/hkOU7XFViTPCJQJrQk+12wz6jtpB6et0C/52tfOe6c1Dy/N/YRcY1pULtTQeT
jXDMXOUiBKTUKAoIV97JYJs+eS89DQocuGSMnEvx8C+CxsNV+ndqj6pJSLfHkoEZVyZg+Q8FOVhF
v9IXiQGfWKpBeYoYGlzBs5otMfde1UmuiKFRvDZpm/PyM3WbdZ+AV6VD+uaOwS5vKZwz2QyhPOlv
T/i4Wnk5uLpXGa1Q9687gN3Jd54DPTEMZ/toPG9bN84v8mDaF6CVgOtIAeTcSa7WL7V4tr3pBRo/
XsRhRySgHoDdNYfZaC0o4DUmaXhdyIiV58yj33hr3/FZsfWNpbCYYgADSbDJDt1XbABqsdn6O0n+
IuTDWgHf7JBDbamQMf6zOoA33h4SYnY/XUNAFy6+l580V5Nz/NxMyRlRFe2owH5pOkbf4jP47oYK
8kzYBVLz+UBaIA1wutPAQKUW0rMVcP0hqtZ3ZuZqoIPyqM8w2KM6kQBzGlMngKWYYsi52QPHtG6g
czFtJEj1oF5G4eu9R971nqW9Ls0AIiY9oUIDHkI1qtf02YCNYcePfAWOb703JnxCYs+3O5fWbn3E
eGxO0dy93mmz/N4txyWPIqsLvVBueiBrd/TdhHrjoOw4LokXqj989lU/SFYaaBsfuRwbYagVDhdw
eqmVbBF9HnwNmX/knQ2eMQe4LU94WSqjVUug6vwM6ob1RvBsP86ULxMEHzO1lwIC6V9gNpqMgpsJ
oWV2vSyeGDkwVUMQmxV8ExO+FZ9UxMowRrb98et8mqZl3iE+PGsNxQttQSJNnA7FR1WqQnx4Azhi
QN822jCBJMQ7AW0xAll0W5kcXumeEmoGGHRNq9E3N/kSi7TAclFz3XcyYv9VsCgCURw7UsLhoLYG
GbKudhJvUV8dJlo69mK8qaDDb4GUJRfXUFmHWnUXBWuKa3dkwBbm0xSIIp9L5CkB7wMm1MoKodgx
MRlVmJTIfXIHEBRL6Ufolz75LPtaAunv7qxUdNd5cx7barMFeM4J3Qdhs7NKC+Bgzn0RpUYyJBhE
dO7KQsc/m1hB/ikVxyAk19Uvoxl8IHALL/ZhhE19dkKHXdNVJ3b2UPvKRygxPIFrlTVdKSu4IgPr
70G2zS5rZRassgJkb+/KGZbxSrv3VQhoRW2rpge8v+ikEYJqVNzSJTs3X22izOLVl7uKoCdBtcvg
/V7LUBZ85z1d+eadX9MxaEgRs4L41aWEJonPn4TfCtgGv2+6djX8YsyZYNyTnqJiX8Glj4B78+n5
sBGEyYm3CNCHo8q0qKoYfePsoSYxmH7FBAEwEC4HwwROcj5BoNrAGnKCgQOL4cqaHEuX3U71y5Zc
J2GO13FIQqaNSDTh7gpXgfKQ7pBLjZx6Ew6zG/ktal0iZvixunlqZgNiNSTegRDlVG82wcgOb0vs
N512s8fzVGSNix/ssbdysyXrRIiemvGDlwN76akfeY5Q6wbVXpTCUK5lv9Y8RCaAgS7DOkNvf2m5
TPpCPsznpOuu9bu4YREuGVFBDmP17NewZnNycCB5fhDtYbhgtGkvQosYgYMcc2iQuttfnnftdBYV
do7ooG2V3GwZgoPnjmO90a+kvXPbQhLtut5p9SnThmv0mfzVovj8RE4dzB9WZ4uWv5w8JDon/fxh
shMB9DNM1CjT5lD6Qixr2JNHE6wimWYqhaNVe7pPgjYKVmeNbRwiEYmbQr/Ir+alFz0/IlnsGrjr
W/b1Z48sCax8+kLNOUiBKeObMMXABMGHsAdCSehnGxaf1Ruvu9Wncmqhp4aPuP86AKMxpusOjfUO
F2ebgNH6/gpvAnCRDgTUedwi7Kd2xLsm+dyZTyzm11+jEre+7ICEZVecJlwEB6CUhjXmK/rE2UtO
vcEY69hmUKRjh9l5NfJdA53K7l2lzSZsK6PQweyZwYMNu7v5RKdT3Z9bmL3S1Df13vZulegDqMbQ
tHqz+7+Fxr0tndDP7pdkp1cknLJaAfjN9NS+m3a7OBn4ScKaV/iVtdT4guYaEVsGmMsj1fV1yl7k
4HFQX0GhGkUoKK/TN+NTNZep4mb6wHi3zXxTpaLwo2chD5dvNhC/VMG0LV3GZQzJEEXgtrRxG88W
smdx4cdYBX2ZNbpQHmq7FEb7BSQawyK5CHpVaBWGVj5ZD9Z9x58gBcg+yR37Dv3Mb1RD92T1wif7
wjmtCXAkTlw6fjE8cgrIVFdJ87eHx9xY48viDeMFOUwX6HeBro0Q2BOhq2nh+BVHEMv5jUSLVo4j
h7N64fyXa2VIZ/olsEIEEFM3yj3ccLoHPQKfzb1RLJRpAZoVlRcmC7t8Yv0C9ua11XBzhUKbMCTL
sqKOuPsKKG9+ZzeKoLzN0QY/usJPOW3j2FAQ/q+h2Y2zk5Mos/ztTxll2+cNxBa7byf1zrKcKR/D
ABJt9Sr3AAhiNAGjKNgbghwGqA+5xRYyK8Pm0pxHwEwwV7C9HBuq0kOQ8rg2VEVBjflGYPF4RVHL
hxVcU2m4ovzeYFxJdtE+NPShophndzZj0611IkUD0SakdWmoN6VCkLv2K2ut9k89Ze4GMghlcGRF
2eFguRR60fzn6G7xwax4LHm6YmQNu221uPvhbuBN/XBgZ4rdGXtqzIsqd1WxApD8rtOFLWOIU0zX
phU1pqOVfjyhfbKbLOhGbY8eYHMzzHgakjxcTu8+6gS6yS5Tc9NpLmL4yGuxb1lF9KIe1HIscNPS
0VNzZw5Nl/k4JLECCyHjrta6vdmOvb6fuiyg/EDQNVWMgCqEJYfanIQNAwRk66SiyIA+7eVnp9QD
amMr2NI3P/S9xYqVRgCsQ99PoVDGUEU1CABbdZxAYJ7H3x990sPOYAQeanbDU3loUmL88/AZ5mLm
eCbD26mcuqEUVuy4xdVknJeHUbV0xrCL8orJrIQYgaC3Y2w7VeW4IBowmn7QxCq2ahZpl8Tbt9Z7
6WhJhRMIlUIwm3eEIQccKLFWJd16bdhxMzByJINZJ/p+Dl0YVjgCuQznVPJ1T2+I/R5BlImBoj/G
92cHYoLD+7DsOwGjX0E15EibzRbCzvNOqC7wdebnGDhhbBg/62q0wf/h9OgxRRedXczSJWzV6Mm+
noSkgDlyfLssakCCUOhyAAuFvAzo+/3+sxp9F6DOCmNSNBbJ31FbHI5fB1PcCJ2e4sCtEuAqAUIZ
EDSr8IjvA74rARpkzMoUm2I1MzO7ohO7RhY+ARgx68HGxbK2P8rGpp6SjX4b1IP9lwumR/cj2sSu
IW1uXnTTQL90fdRExb5tNDzMtlMP0tLL1ZGVRszBgQag+/PbFAB0KYH1V8msZIxsXcq3j4/x+mjR
Qx7fy/CZ6KadmsF0JHg31bkYYxbzXexiwz5yE2jeJ+B62OdQVMn/87JVMvefAmyyQ34euJC83NQC
hcGX9hLZxf5lWp3Z0LTn7bf//VWq21cZA36BCQHsDjVYB1HzS7QlD2y7liUbwAlZuC3f9eVI6+dg
yEBtru7mANIKHyHjAxXbdBHIJRC1fbZgIbtoO1TtxZQ3B3JAtYL0sf0jnvnSlbF2ECgX/SsTZnRe
viv5/euLzXCtVzCdhS+Ufws124u0HRURewmF50y1i8TW6FCEiTqUILIwpg2bMq6pDC2l+vB0e5NS
7PGO4wvlmtLgurww1rozLGlnwWMRATjfB0LYiD69HOycJhCVAzaL1GFLShLFpOWVZ4QQmmJV4A/E
X0DqK1u0J/YTdETNETKriZzbJDPli5oJtFwUoVIPIUg5
`protect end_protected
