XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���b��{Om�gf<_����g����s�>w$�K�M�%jC��(IѴg;+��ٯ+�\ݜ��k����3��aD�o�dQF|�vl)uꕫoA3YS�N�#B�z��s��y*�d��yjU`ڍ�T
+eа��}R��K�K�]���&9�K���;#������5<V;$�͞���roB�'J���y�����k�n���B�}�������&Z�y�]�SIB/~V}�,י��Y��W��57�������}R��=x�V���)���� 3v�2���,�d�n����ᨹ�Y�4����/�X�	��GGU/OY�J���7�6ԡEf�hٸ�h8=��j�S�f�������a��|,�~RE�hf&�^�(ޅ����+F�\����p�`[��}6=DmmlڏX���bP��}���~�$�������h��#l<��F�dO{[��P}wC����N�7���1��3�%>�7ȤkCA�,�z�<��t��-V�w� 
�^�K��h��ʮ��/��E|�B)�����3�]��Y��v%U�<^�F�(,_RP!����/W��n�����V�
��4Lv훅���a{۵Ӄ ^��@���d��k���2.+������?�s����ʁ���Ⱀ-B��k�OX qڏJٚͥ8L}4?��=�_���V�W� � ���l�s��a��ˬ<*Ǚc-Ƅ] �J�`|g�E�ٓ�'�m4]�"��gJA��;a7��-KR���~t*XlxVHYEB     400     1f0��T;�(��e���E�^~�}�������a1h׷���Wa���|K$jG��G�_�0�|�16��?YP	yO�������'��}��h���.��3.Ա椹�ƣ$fⅾm� �ѕ�@bД�֞(=$DT�(��.� !�"Iq��F�y�@"�E^�P~Ҵ#����οWov��<�Ӷ�J�.]����a�^R��Dz�=� PR��
B�#�K��H%r?�9a��
:���Yy`�^����V"�Fz1w����[�\�
��|��
����X�9����=l��J�!9�L��A�6��=�ep�ԓ'Qe���Z4�5�
�8�#d��ȕ��W3t����?t��k(є�p�SWT��)��t�@��ay��v��1G3ROL�Ս_�7EΎ����$���_����]N0�����Wv���sȜ����\̧�N7@����X�c>��V�5r'�;DB��3����-���Cě)[�XlxVHYEB     400     130���lɡ����u܈�J���Ɯ(q�,�)^��`�H&Q?7�ƃ�!�uxTgr|'��@�k�?MTa��H	���*�w�{�F(H���(�P�[��m��Dџ��C��q�d�{;� � ��2B/�W���8��ɫ�CeY$�O��:�>�\].�*5��G�*��"�q!�M�������_b�7��|�AU絍J˓����&�{�c�7Ag5/�����w �5Z�;$��~��xy㵱�S�;[#'�{(���wn_7�	"�6��:ב�{zo�}lT�Ny(��.�k��$\0�����`ZXlxVHYEB     400     120i@���_�lc�HM`l{��R�v6��]w�4�׌��4P���e���Ř�P��z}//t�a�N��-�QV��øD��L�bZROuz�f:!_����~�x���e�S25�����)�U� �Sw�,6��W�xd.|��$\?����I��&�u�̛M4=�]"��OΏ�"��T�E|�\���̔�/u��
���l�l�XK�W]�00PU!��/��x���KA��"��/����jb&*��0L �[iڂ��(Bk\��0��v��EXlxVHYEB     400     130W�>y���f'��U��z�pi�Y��YyG�8P���@nK��R��6�DX��ۿu$#�G{���iø�:������"�
<7��(T�Z�DX]�9�#��$c�O�P��z|�kvp��Z��*��G�����C��U�ܠO���y�[�v鄿K�o�c���NA{��ň�3Fn��<�`u��n^p
��Ȯ���6G_Rt��;\���z��:ɇ)��p�5X��\���މ2Q����Q9���P����~#�b��S����q�L`�<���_�Ud�1�(�f'3����G؅�X���*XlxVHYEB     400     140<!T2e�+h[�BJ��ϗ����3dl��X�oY��Q�M����CԱ@�8�r��*d�i_�"
�5������u�è���\����b蹼����R^�Un�s����}
�]�	q�!����Z�$��"
N_�
B�,A0��8���q���1����
���(��|�?a�'r~&��xxV*`S��q�/Ӄʌ�1�n�X�@T���)�uL�D�ɉ��;qeA���Y.���&�+s���)^��z�M�_��U%�3T[����m�s��~w�zEF ;������K?̦הD�o0O^�k�T�
T�G��	�XlxVHYEB     400     1809X�7���d]:�}�n��0͹��/P��S��ß�L�1�!�Xh���V@�S��b��
]epu�#�@�vt��2ҤǅMu�
�W��Fw�Z���H�����1�j��C[8��_��GH;��y9��=ўmja"B%��gW�w��Ϡ�ȑ5?�d��ID�,܃�w=� 5�iԂ69�p��\���P
$؈����D�A^�'�ɭn=P�l;3��sb�m��2y��QVGG+}ݤP�sQ��3��J(�T�.�P0q�7��0~�H�b��F���|�z}>��G��}�N�8?6����0nf!�(	@N�q�Zi�Q��bF�=e�p��vl�_`��Xx
��p3�]���3`���q���p�@:�c�I�E���R��XlxVHYEB     400      f0����h@�s�]�hE��䟐H�5m��'��=��뻰�P�Y�\F�rͫ��:���dQ�&��0�h�\����se�c�3�h�]	�5ro[9��fȟ��(�5�^�I�j[2Wܾ�@2r�ݸ�����B�Bg�A�z��0��t̘���l�\�	�rNx/��"Ξ��tN�1�1p>%����1W��֚NI��(�_ר0c�q(�L)v�D���f��"�b=M7�<�XlxVHYEB     400     150i)C�:����0��)[�C���T�H��VB��'��:�5	��j0Nf��Ƀ?'�z��p�m�|��Iة΄�'��Oy��B��}~�[��?��D�NS�z���:�o���=����`副1�',��x��l:�9{i�(�k0���[�J�W�I�+4�eӍ�a49I_{�54���i��
 �����#Z�3`��v��+C��#�!��<L�@��3LO���)PK���ڭd��j/����}d�&��d69B0��K�+N$.B��[�+��+�����{��w�am��,*z���]Z��{�x)j9�Lw�#��~��)��]r!XlxVHYEB      b5      70��������h�L�\��wn�?�
9��g��U�c2?�d���)8���./��%��K�P(F{\y����v���G!�*�>✊[?;��+�0��`s��i�����%�