��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ь��-p�l9qe�p}����y��L�Xݳ�,du~{�/�mt't��UUe
�"WJ�>��.���as��^�o�r�?�>��{�z0�2|K:��lL��+�4gejCx3V�+*��$���$>n�e�*t��I����5y���/���ͤ0�&_�[�ڀ%'=E�JZ���^��Y#״i��\Ce��噤�7�&Я%�
�r��ESƿI	��!�"�XN*���8��X?�(�������=�z��Hl1NE|���qכX�ʦ5�C6��7������.��ۥv��6É?�%� �.ۯ��<�b��r��`�x�����Q>�T]E��������1�S�J;h�nR���D>1�B��`��K�$K$[�*U�1Vu\�A5w&���䂫v`r�_M�0�#a��ck��B*���9�r��ã8��$�UҎ������ 3H³ʾ�o6ߔ�p�$$�E98��C,��Ԣ�ϲ��,#w���A��"��6׭VYG���i�D�-���|�P�*42�Kz��c{�+ظ:h�w����Rxƨn=}�D�J5��"#W�K������8����o��qѱH����2fi�@��U�X�`���(��_y�������O��y�ųeޘ]�G���aw���SI 1W=�>��B�+��t�!Ϊ0y4�"+��_Y�D@S��>k���B��d�?:K.����`D��(����O�%59��r�����6��sZN\\�=�N'"��;7�F��ȉ]?C"B!}VC� ��Ñٸ����l[�!Y����6j�1����m�LA �#��	��j4Ti(�� ������I�ԝ��U,G���"W0V��{|[y�Z�}݂��P_��Pr]��ۄ=cL�	������wB�ł�1�2$����^�l-�f��A^7ބ+�\1����_0zë5�v��^��]Q>�7�ӓ��`4O3˭� }xF�kI� XL���� Y?���W�/u&���M,�{�FF�|�/U�Y\�����A�nq*:Q1��CǗ�%���X��Z��+$G��!�7��Ztf�}c�Թ��a�v�S��%E㌾��%�V��y�jԇ��.�-$�z(<�X��f�E�LF:5B�������9�՗�bP����r��9+#z�˩O�	c��ˑVvp]�����4Mk��(-~�eטI/�l%)�j>�*4VJW<��`��M�h%\��W��xg���)ǥƙ��$���8ڨk�����D���wL�Y�Q� /�ڦN��S��%�e�7���z3�$�=���*wЦ^�6,�c�hY�t�Rf��I�!(KPn�
�5���H��%�p7��=c�"�K�3����1�*�d� �r;�a�o��_ S�)�����@� k�/�ޯ]|� �h��0C�<*)bc4�-tҟݼh0��af�'��RV$��T�V5���L�iF!C޴IZ��_1)A{�X&�F_Lxn4�v��^9�=é�&����Wl�F�.�`7�!|�6����Z-^ �`��&�a��v�/4'H�%����!��`�u�o���wt���h�mah#U%xm�ۃ��s����#0��X-D��(��ſ]QfG<^7�)[]^%6"-XZG3�
�$�`���LV� ���!a1���(��O���^�hr�r�[/��I���}xZ��Q���g(��c�pB���0�ЃӚx�SdxN[�����Άl�A��w���A�6�X����5���A4�ѡ��;+4O��0Ե#�&ւpGG�/K�K���N'���~�N�8N[�&wu��9��gr�����1)���,���UdN~-�+�̲��@#:�#�B�.!=(<1�L���DX:�[lE��L��}����oJ��Rڞ>-�d	g3�a �5:_�#R7��J�EXѨڣ�C���lA�xM�֯C��;w:�E!�dH�P�s�;����cRQ%�{����x���P����ku9O�\�6�Ź����&<+_��U��}�w�a�.Za HA��]=�2[q����bA��SG+ߚ��N,�2���� qJ��᳆���V_�+yJ2��)�_2D�+]A�m1@�b��_V��2��x����-�	��m�*���'G?�|�ҁ����G�*������X���N4?�t/+���-�"£��,C�B���"਋��	b?4�M߼�DC �W�V�-���S۫�o�r��G��%7�k\�I�J(�A}�}u+�����0%�p��0ݹ��y�u��F�Ul_��5��Pj�~7��
,�%�՟4Dǩj�;o������xWu�\zQ�7K�z@�h��\�y;]	HŶD?�Q�fߞ�{f�-�Knǅ�d�ms���NN>�D�z���:M����`Vع~�F�Ѫ��#�33��t�؎*-_�`[R�k�h��~���J��Pzv���׎pN*ui�:A^�=��b�0�saY::���J�?����Ð��⊮W�nt�]GG4j���٪Xk|�q̂��@�ܘ�5�B��Ϻ���o�� N4�x�]�^���z�OY��<'��q9�r�}7];/���J9���key�V3j�Y�&R��j��t�%���=��gA�ȯ8'`���B��1�$pL����L�B����,��D#oh�!	(o����9�����e��6�F�]�j�ȟ��%ǉ��g�i$�g5��$������8�imG��(�wTX�P�H�ʒ ��ukR$`�g+aR'��u���fȞΩ$)@:y�`0(��犽�{�LR�%��I��&�L��i�B
�;,�-+n�wX�e��ȫ����+���wĜ)��Op��-�*d3�)�3��[wl\I�Jf�J�L�:��m���s����C-k;��RԠ�<f31MGa.RTk��]w���c��S��Y��]X�2H�i��c��[�4��:�U���}��\�y	4���]qC2A3s�8�nePopG��_�{H�s���s�)y�==�����`��n��S����
r|�����ZE6䯸"Z�"��X���S�o�uֽ����;�Jc��#��x��M	�(I[���w�J�ҩOk�圵8�(���h� ۮ������wO�<�wɧ[���mPm�& в\wT��_a�Fq��*;w�9ޔsB��߃C�l�b�Ӗ�^�*����Pd�g�I-��g
+�x�	��f��to!2,yP���o�%����}�ܰ�E��x_k��7k�WX�h�bQ�����F�х�&�������v)�6�(���p� (��'b�X�5��&���^��*�n�1�qMȒ-t�˷gp�J�GQAn�u�!t,]�oָ��`?�#��9n�`Bj��x�&8�*G1�C��{k��"9���. p������ ���3@f���Ly[+�Cr ��2	�˅���Dn�1���\��ߠ\	##!rZ�&�.v��4ַ*$��(nŮL�X��-�k�h�K��ٶ��θ �5��A2��h��h_�V�qh[����f��*�@�`	�R���~	Q/�(7��z��n�HN�С���#�� �'��G���.�
V���a��$�t�d�&Ǿ'f��i�V��+����6%��ѣ�:[���'NE�Íyq�b�-Z�>�'=���v�:hB�ۼ���y��۵Bxl�V����������昺B�GF�m$�.v��:��2�7�􇪋��3�S���'H��|\�d�|��t�ʅ���}���^�D��6�ƞf����h��kA+���T��0:���׉ꠓ���u��ʰ�vo��qd9�4l��"z�.�q�m�G��*�����Ҿߤ�*��Ǡ��4��*����r�(zmL���4C���.���_'�"L�4%�\���G�F�mۃt����_�֗`wi��*팉=]�P�ؿ+��ezk[����t.��{����3k7�o��VbH�K���rWGY�M�[�^(���ɚ�GХoY�+�B8� F���C=�X���#�ƈ�l�3�7��-��!�w{~�n�^b�&���ȣ`HTw�����o�Sh �8��醰��_.���J{T��ԅ������i�TP��̣Mv�A�tq��U(<'�^\z��?�>h�������?�0^(6��ge���_�MPH����*T"`����w~O�r�0�>$�>C��H��i�U\�m�,6$�t�5��cV�+H)ܲ.-�ݮ�z����R��Զ�R��)�.$�Y|�P�����R����ʆ��U�|M��R��J���TF<�0���n�'�B;�R�c����Շ�m����b���d��b7ǥ7B�p�@�������Ι|�s�o�����o�u&kZ|QNj��	H��Fl��<��y��}�Hڪ!
r��=F���5.����ذ���d8W%��L�vՂ�G�<��9h��Q�ÖTf�a��t�`)gDP��3�]�,hB[��_�1�@!\H<,x)�Ɯar9���v�0��
�5�*�\v*�!;rF�`W|�H��Y�R�P�����-�Ecx�h�e|���W(��$���_dY4��dc�����6�3��ئs�F��8�i�L�<ᛧ>%p�Y��\�I�BO~����V�7��Vk\N�o'�Q,�G���U9����A{)���Օ�A�I�>�G��T���e��k	���u���o��ݨTH �t���e�?v��࣍��+A�r~�A�7Qm��� |�E`�CLyۡ���
�'#��G�W���
�_,_�o�cS�H�����F(�����)�_+'�Ӌ�3,t8ǣ��8�<����y�T��4�.( �=Ӥe���/���8oU�W������H�&x/Z|�F0f� 恁Y���h��Uҙ����'�n�:�8�I�<�C��a��)Y\�Zy�~�x���f4B�^R��L&�:M��?��vY��i�����!���B$Xgd{�Qak�H���%S��� <�w*���Ql��x�~���W��|���<�����cs�ƥZ�:d�t���t��nC���������"'m�=Q]�̋,/���5��xz����yYd���&�3�q��э��5u�_$�w9ˤP���4t�g�,|��E�O��'#G��QYA_��=:�GO������ l-*�~dm�dm�	�h��������$��\���?;�8�8gH� %��ú��
�/�2��݁�)d��1$�>^;�E��5�M�������0���L���5�1Bo�{�,����/���Ù��a�BΏ���)C��׀h����l���"[�B��f{|��ue����t�ΚA{d�gVe!�d��H�:�����Ho��Kj�V%����$O>a(�Gۊzim��\���?����DC޿,�Ji����@x)����}L���q���҂D��^g�⵩��TҎ���v�FN��������$�t֧?�?\��ܽ�p;��h4��l�2���r��K�DH���]�n�QA) ��,�?m� ��oo����%;HI�mM���OI�ȗo��a���BvѴ6İ��MФ�t�;�sZNl�Ȇ�����,�̗'�%_�߹:1������M$)�5m�UTgT4��a��C=� I^�iB�s�����2��u���,V��d�;�z�$�d�hS&�i��N_��"O�+�j2��}�
����CYk����zoP�Q�S����������D���'��*���ڔ?:I����?	>�O8������s�ǎQғj��h����7n����#���x��U�0w��5�n)��{4��l�8���1.��k�@GC)3w>4�1��g����Y���ܯ@�"{P�ML����$C���kY�<.�Y��I��"�uj��j�3^,�/6tn_Z��ːT�,�c��H<߯z77�<l&�Tw$�_J�	~rdo� �*�$��Ad��d��ۃ�D����l�(��#¢���O�+;{ka���qC����O��O:�����gc8�� ~�J��m�*��V��g��'�b�4���Nh��#�bD&��){-7 ����B�Yh�%�(����T�$m�n=�)bő�kPs�K��L��)�@��-�����b����dC��0e���J�4�Wp�uN�~�����ɪsd�u�ƹL.�ko�x\v�|YH$��N�����PeS���#a��TE��gP� ,C��_�L6��#㵾Ie疥�Š�\|�^ѭ?"�0JĆ`���=��Z���O���5+¢�����F(|���2��f^�A�ݦ�&1p���5�d��v�1ݱ���N��8�ؙO2���H�As��ה_��,@󤍕���g~#-D̲�s�7|J��'�hq��~��������0Gl��h��?,��@�"����`��UA��Ӝ������WEwz�@h�^=S�T�p矧��HJBjw�_sO����tCb��_~��p�e��Fm�>7�N*Q�B)mfZ�c���],L$ԩ*��z��4���+3�]ƘI�%p�˨��s^p�NG���Z����b��^Ӿ���
}�3A��\òX�$R����|��D��DL���9�#A��WN���=�iC�3��H���7�X�+���HP�vkuɻL �}�9�f_A16��<~�S���[K��=!�íuK�]	����л�ƃ�<˪2_�=k/����[L5����*"��޾���^^�}�ﯴO�}�A��<@3�[i,��S�ƝQM�mhܐNOr��V��V�����A�����;�I�?�0�=^Q��͒g���Z�AÖ���{��Ï��}�D�L�Rc�ų�@��Ə�f��"2AC3�+Ix~��kC�OG��(a@��_$�'��\�{A\��"��������O�Z!Z$�E�ncI1 "ȷ����#)=G���J|�k�`�BptZ�N��N�V��z?��'�N�]@<����XI�3���{�5�t��#�B�go�u--�O��j�گ�內��#N����hY78[I}o3�B�S�5�K.�	��>���ٿ^e>������ρ�yS��%oV9�"��-q<�#o�U"Aȷ�n6�qU��
�7�\u����N�'cw���Qّ}#n%�V#��<m!��*I�ѽuo�3���ì
}��v�+�t�`��0�z��}��"'J��	�$N%K��\��w��;o�����5��C*�����V��kd��3��o��p��=@iv��K��|F@�<j�	�/[��I��A�P<ǍTG�C �E��r*VJ�U�S
�Z/��Kp�r)�
_�8�6~[ߛB�bkX� q�հ��?3	^�\-��-H�S<N:�)'X���<��1��"�bC@+a�Q��������'/&;ZܑX����иC~V�=�nen^z���/i���3A�u�����͚��;z�/��X�VwB���{�E(^�����{�!�+3�N�����C�J��������;�6��PWMy��;�r�\#S{3�W�=6��� A03�;�K�O6v]Rf'y��r�H���ci��@����<x|_X�����b,�YpD�Fc1Yz���ut�!���w��4��#��z���N`tK��BS��IE�	~��n��l�G(������o�I�s�5,�����b �댟�2@���@�&� ��&oy�鹇�H"��5vqW�FU�F�I�8
Q2:����c��t5�<�R�Ҭ&��ɽ�ϸ��"��~/9C?�2�i{UP��ݓ�LF� �I6��Zи����:ZY؞�����ם��܎q�������3�l����� 2���X�{qj8�|ܴ��b�[�
�/�^��V���nD�1o䢈������;r�>8^���tn^zQ�h䙃�?�t&r�(��U�#�>�`��h1c�$�
AN�Dk��RƏ6��|"��e9)(.��)I��0���]��j�ً��u���B�}uQn�T_��a����e�������|d
��9��[���Ê�^���^��mj��͟H��c�a�9����<gl�Bȇ͛/R��y�^�i*}\}���J��jU���4�KG;!���F�������ȿ�/� z&�ո�&m�w�^��q�iZ��[i�t�?�$���oc��&<O��bĪ���V��i���E"�����Gm3o{Y�#�Xڄ�ο�˓�iK����~w���9���˗5��i��5�����x�!����͓ ��8��s�c��<��(�0)�:�ZZ��Y���ի��πp�˪y���;9���a$ȷ^�zj�B/��%���B�)ȗ��q�vJ��N�����^���	RB�<F�� j�'��I���J�Dq�h��%m�Hl*�VO��64#0U���}e@gjD[��/�.&xxŶ`�mI�kzN��o���F��\s ���)�}Y����F��߈__ע]�9���PnM .xu؏���&��'����x)��F�e��+�w]
P�P�թ�m�*lC��l�gEH���T����#}H�.���XD��*�X�����6��:P)�g�D��dq������u�l`�ȑ��X޿��W;��Ͱ���}N�C��<��Y��m�(����,O}����U��������"�	O���}��=�4���j���uJ�^AJ'�U�/�_�"�6r����2�	��M�Ǭ�ͯ}O��i��n�/�z��3���ϵ)qK�PiV?,�N�2n���c���lrA�>�M=;��d��#}�7�B���N�HKA9���`�6m���-��wj�}�խ��ۚϑ����)��s���拿�}=�ũ�t4O��z/�SJ	Ҷ`ͯ> �N�'����2}��90�
`	]e��6�c
c�4tb�x�yT����3��A�uSZyKd0�rF<���|h�w�����TL/��C�:��-����M�;=�2��	c@~ ���E��
��/�?�|��۝5���0�MDr������v�~���۶$uj�&&$��tW@A�܃������#g�j_�&��Jn�����&��-=��t-C�������@X���`�{->�9�ކ�w�N�}���4�-�V��=�j�~���J;Zz�Yd�2������}�Kx2a�-ݙ��i�nOL^�����;��#�VD��7�ǌ��d3�x)O�D��&�|߆������]�)���!"�qp���r�6�YA���l����� ɴ~�r�R��vl�%�h��U�r�,�L�VQ��U�O�4�+V��"�	Uh��$������.d"��B*�BYP�|Wf��������]hԢ�@��ct`y5���m�៑���B"�a���jIX���iߤ���H����8������kF~���ˢب����<�w�Ŏ-�D�.{��7&C�O"�2O�;j� zeB~��5���Fd�V>�=h�:�Bp�)��%�����l����?~Q���+�a��x	��F��,'Y�k�h��|V�2��S򪵮ev�Ғ鰆�RS�.�.R;X-�2�'��k :I+m��I �y�Pc�Z`�h-�����kݶIkS�لU��oh�0�W�ț�:�k�V
�L:J~n^�
`�X����YVs��x"A�4�&K�C�@���6a�ď�~\���d<�����qi���jH�2e��U�`̭���ǁ��z$�99�R#o�9��E��COHd�j��w��K|�����z�"���#��+�|�ot,��C��Q�Y�
���KP�Jy}�
��s���^1�k/�֦ϭ���`�U5,ĘUB���ؕ�����F�,�q���(��9@��)��8�u� >NQW�T�j�S�܉��ɉ�Rk��w��,�Q�E��po�-A���F���tA���D������sl'�t��gW��S|Gh�$���A�,/�� IA����RG�pnj"��ͨ��b��MG]P�	g���q���6�E�i�.�yo;jd�����<anA$�. c��Ɠ��V�&V���r��T��sD#����N��al�]�
�p^�!��WC,>��W�p��}4`	��DP0���x�<�߹ �����:w��j|�䏤!7N_�N�.��SÇ[c5ulF�̏խbxj������YD{iU�C3�+R�ZV��ڒ�񑎈q�F�=x��%�x�5����CU�z)M�nwlYf�=��p�#�o�n�����M��Ja�%����yʢ�	�qi^���kj���*�*�$�"W��|e(v*jeJ�h�]^�VN4�岂�l�����7N��V[�"���慊bP��++Ȃ�����#��4 CM�RN�.����Y��'�^�I��w�Ϛ��0qw��F ��R-��4�(+Qk�2�~V��n;�359m�ӫRaapen4i��䀺�:��[+��C��,w�0ڕ1���-v�+�-�+]���
�����cf�+ɂV��S;�Y�ԙpܷ�d2&��c[�?�Pe�B�^&��M_��-�Egggt¤c�1�Fb˶20�#�ڤ�L�V$X�Q} v]�j(�[fjAa���l�en��;�DBn��Ɨ=}J�V������3�&(�,�qni58���f�@������"��>��J�/��ߝ�#���tr�����L��W��Zp�T}"��G�T����s�ӗ�&�(.�u�K|�o�wt��p����e��8@{�"�j�����_�Y�	�a�bnW'gM�,�/v ��/zS����� �0�\��p��X�^�1F��y�JYL���'4�B�ڹB/�jˣ�L+���FѾc�H:?n�
F���j�����e�$-��H���x�9��%�0
�x�$��4�g]�I�Nʿd��yM�u�����c��R�jܗ�P ���V��,�� ?c���?���.*��x�f\��`m:[�2��~>T�%%bqG�[	�IKF_U��:yy�Fq���ڎ?�ؒ��"�l)�A��Q2L�W(k�S&�6o-�coE�:X�f���m�#�a��L�1���g���z��F�b��z�C�5)��o����'"F�L��/ְh��V6G��	��B��&ܔQj���0����w 9�"��e�cS8p�Q���r�P�qIY���<�CH.�;b+`�
���V$_�����8���Agai�tN�l)9�� ������C7���PٯT��-�/��3���h�~�����:̊�h����m���vD��kZJU�z	�Ay֛��u'�!�i���tE�;���@�T~v�=�S����PAQ2����<ƷϾ�ס.}>���X���Ք��ol��j����x��sMMav�e�&���&@C5���j���������С�l�d�SY|l����e��z-��q;�vw����)ٺ+	KK��_�_
Ā����2�@�V*{���|�D
SpA2�f���>5T ���v�Ci�o/hZt��j*�X��#�sL,G-����T���%q,���$�4iR绐-�d
Ѐ�5Z�:��%1��߲q2�d�J~�J�z8i�I#�G@c���	��0�nx�W3�[�f��S���	�X�SK��A��X�3Ď�]<�!�������ҽ	f-� lgR��T&��UTd#'�A��{�ST����������A����ZOT14D��N�[�?pN��q�
<��>�]����?O��	�cK�)�S2z�8��v0��R��D;��dN�5c2��K��x4�wu�˂�xd���i� V��!F�vn"q�7$Arn"�?�,�<���*�:�Q��x*����TU��O����_?Y�%I�A���tU�w�iTv�9�8����s�[p�mP���Ʉ>��$����	�1Yi=l��f��A��r��?�8Cf��iܿ	��8��wo�H+Ո���	 �)���)��H
����o>FH���Zn�Z���bpL-a�AKA?C�p&<+�ʿ��	'H+� ���p)��c�p���3o�I Ҏ�e���݋:��Q��u9;g�Fѵ�͝����@��* оd���b%	�;��I��c �4�����L��ɓ�\�g�\]\��'�_��&X'�]���VOT~��۵�w1�o	� 3m��^E}�·�c�ƨ�pP��1���i�Gc]�(ξ|�zb]}�/�����kX�[���.A|*Y���CDN��Q�~4�Q�W�q(�����>�����W�.ϙ`�ltNet�yw/�+Y�D~��B�a��V
&��ɂ뀈�LR��;��H���$�T�w��\��#h4�K�g$���k���S+���Wr:�K󒽿�1�g�\c�2��a!����L��#����������hwR
QB��F���ȉ��9�!��I����������?MW�+��\�*G��]���Tv_�)@�g{�M�Qg��ǣ�AZ͗V#ڧ�\"�ٹ���	yH��䂣��%�Tf�I���#}X�N��ତ�T2���� v 		R���	��ԭ���ws��O\!�¸�b�t��9�%�2�t���j���0�/�E�!���4c���f�C�.��J�u�C*!g��%�����~Q=�FQX�'ݫ5#�U��mYF�sJ��hA��.-5��ھzT��7��qu����+	<��R��X��W]fFH����wc8=*IEA�������N$Y(|�$���w�D�FǉVI;A�F]��:�"�pᣗk�_<V�W�t�����K�K#(	?�B05#��o�ƹQ�-[�pY�o^�����C�`#��3��떕>~�:���*D�y���.�q�)�h,���7�����O̦�TN�p��}qAԛ �@;��Կ�f�U�h�1n����p����\1%9;}{��w�cW^�����)�o;Q!�r��:Չ?�!����beW�+.�D�f{�ֵ.�[^����
i(La�?���d몹�YD�yT}CH��,d�{7\d{��&U���&��f�n�
��Λm�X���
n �W�W���챋��� )/Ŝ �~�f�ÃP7��9��Xpصș������&V�T��AD�)�}P�������nw�Br�����6�!|(��K>@z�8���Y	�1�QmɎ%�|d�"C���"�s(b�4��=�.�j�c��G?;��v����RGM�K8�v�#/��� r������YQ�*=����uHy�N�A��F=n�Tp�P~�1Y�K͢�b6��EՎC`��Z
�L�6K��.��HDπJ�����{Yך*��ӑxd^N��N���c&i�NL���̈g߼7v։8�0�=��Aϧr͹��OQ� ��4�'�[�(@d�-T]�3>ڶ��I%Ť3�cn���&2����)0��>[�1Z亾����ɳ#) 26k�5���"���5,�����6A���й���m�RT�'M��h�4�0���$�b>�5�r����Qa�$��c�~�J�N0x"�_���;�"��"Ԙ�lәӈ؋����ȋ�}�&��ĸ������9�K���],b	��}�6OJw+�^�ZI�</��(-�	���N+���n�
2tMi��SE���:��St����
"��Nm��n� �7�i���E��n�ђ
��nB�Ց|� k��u{$
V����� a�(b�o5ːI����]���zc�U�C@XHDaRg�Ѡ{�FU��-��������NdMu��%��뇻�}.)#��'���������
V��E�n"��'��=Dh�L�"?x�E��ֲݣ�uh�r���
-���Kl��X�/_FvF5�L֗%\�!#ǟ������|���%�u�BؿA�o�,Ww��&�SC4���_QW:��JP���*�W��`y�{ec� q/�QK�M��r@f�
���P�>�D�8��Ǒ�P���;S�@(�$Z�z�'b^��֢��(���;)�y0*��$q6���:��͉~����(��9%��@�P¹:M�,"�!�9����7[��+X�f��N·��!F�!y�X�"�Uˊ.u
��ޮ��I���Vω�:�r������Q�8�1D�Co7_l��+|i㎲if�U��mQg����Ǽ�@PI�����Y�ʰ?P4���n��Cf�O�d!\� ��A�(#Z6�[���NT���tIZ���QL�����S�+6P�v3��*�ė;�ط��0]جB�o���5Ұ�h����Sj/򈴗�Ȃ�P�����ls�o^�`�S�h8C��Uk���9�hPɬP������^�;d{���$p%'��5$T?>I�g������c�><��J:���J���`� �����kέ�)!u�	 ��<XTT��,z�C)��媝�)�	��� 7�O\DUY�$W\˙�ޞC��x��B )�����0	m��%��I�F�^o��*�����W_t�h8"�S	6[ċg~]w���f��"��Yc������L5[��f�^�����y�%4�5����Ϫ�kc�4�җX�a�Л!q!cbE��]`��*>9��ght�g�PJ ��ͬ�ᔯ���I�!�ޘ�N�m���K4,���(>��<�L������������+" }$G=��a}�4c����g+.�V����dM{{ny1y� :w�k;#��vv�D9���Mjv\9�&��KJ�ZrU��/4���4˱}�����O�uOR}�[|O�9sgǈJ{f���u�`�l�tYگ��|"���N�ʽܢ�8[H*�k*Z��j7��Ho)i�	ĸ����'v�mxVG�#�j�|���뾈��S�a�D��>��yT��[�� J]+���q�:,��DYAL��>�B�I��`U��_�&��HK-� 6�h2y�R|R#��_���0�#�(Y���¦��$R���V�{l}yP��;�/��G�]��q�tu �5 Y{���M��>��q���qo9mJ��)�5$����D�T�H��Ĵ�z��a+DE��w?}9���zaҶ��tv��5�㢨���p@?�����Q� �6}����r[�uQ��:�>�HX������ۅ5��Rs��� ����)�'k��2qJu
���Ч57�:f(�����x�B�D��C�]D+�|şv�K��-��'BI�x#� �vA�1S>@8�%F؀A�-�k��l�Qr��%���M\0+oO<l-I�����2Kl���-�w�qn-mh<�&妆(R��;$��\caQ����e� �N��L�{��h.�m����$	�׶�����co?bӳf�=|��r��B#��PO��H�3PM1N� <� cd�By�E\�fzH�@!Gا������*
���Or7_-�dy�zc�^f5�����(A��X�y ���n�
�K����W����bUG~���І��?S 7<Ӵ4�RH� �(�7RZ��k��֗�4��]P���I��k߶���Q�n�T�o�3!io��s9 �/o/{L��B^����$�c	�pw}���g<�uG�!�wG��\�y#X����߄�[�q��sn.����3�J�'����!�ƒ�QT�?��̔��(t��Td�P�'�X�A�ggX���������+[����Ŗ}�CR��@G�t�Jns�ԁ�m5^�0^�� 
��%F)m�͂��}�m��g��4r@_^��c$E��sQ�\1�z^o��s�\u�0����/�!�����6���"T� 3��n��a�SXP+?]D_�K�5���a��L�Ƶ�ML� -�-h$�u��x5II^�%�PYC�?z�n�j8� ���7k7�;=�='������'�-;s�;g�0��f�KI�s<� ��ڝ\:�5�84�{���}�V��Cd��J]�L���ѣ^���nC�Fs��6���!��d�rw���h,H�|�W��җ2�IM2NA���n�Ȇ�'?��F�,�y{��~ʪv�J��������ܐ,K���9�����t�U0��_�~������P5�E%c;�(��0	��-��R����8ty�1�v��?��/�>W@Tc[1&˾����@��*i�ۇYxB���c�q�<�|���'�jQ�EA�ة�'�P���v�'(f��a�����		p�����]Ӿ���Vu���"�[�1�tPZ ���A���'o�󪕟�	���s��]�8�����k�8���z�N���M�+��Z��b�_q��A&���s:�S��a�I!���ܯ܎���  �z��.ZM�����f�[!�*y�:5�Ƌ��_o���P�̀�?���жc�e3�p�c�oQ��G�M��rՙ^;bBR���r3I��z~�#���M�B���0��
����R�RA(�m�3O;�.�����F���멝Rdm���k�N���BB�?�xh2��I�� 	��I[_���鶦n�?H�|�H���Rߛ��n�y^v}Ƚm�t��A����H�5%����Y����q������?�['i�,}ިuV7��a����!O[X�w�_���⟈��\|C8D���K��Ú�~$��I�n��`d��ڴ���)XA�h�"Œ }9�c�D�*c>-��+�T�J��)�B�y�;��^-x4޾m����W�W�����]��E3"<��X�e�t�3�<��l��(�����=9�J��u*XGD8u���|ќWЈ�T%����SwEk�\@m��n���.4�l�ÿ�z��M�� &a�Q�����뻉��§j�Dvҳ�q�H�ه��"��'Шo�;��#ِ1"+�g����O_���?�M�!�-9W�\�m�����%�fsUuPC�S�0^��wr����|�f.7��=t(xIM��Ph�&6�@-��>4�T�"�����G~�|��r5���˹�<mֺ&�IÒǎ48�Ro��׭x���,ɟR��.��@˗L�'�hAc��g��K��O���`bV�`���U@T �����������������pe������Ǟ�D��8\�*�1%��Ci3&[��7u��v�	¡�;IP��Q;�I�����2۾?<
\�0���b8j���ܿ}������������q�A���Y=�hM�G��< ��;��[�u��laD8
C`O�C+���F'H^D9\u2�?+&µ��O<�1}D.D�8����Rνs��>!�e��J��7�a�c�0#���뫃_t^2]!7��>��$I6XC��@?�`_#	oqLpC��k����vGmzĲ>.���w����,�/�Q����ծ
�C� e�7c�^gI����Ab�]/�O6û6�sǤ��v>��L�촹y�s�E��=1�͎��
�G��#�!u�c���N�ePh
�i�,���W]�M.w��@��8>�~*�{��0?���n���~��/��i<��W	�Ƙ���=j�S�E�C�������ueq�U¬��
�d����$0��d��l� �u��t�wǗ�Z����%ʠ�m
0�B�Q��}ȗLP���q����f��B���
�$���>� �7���c'il��6�}��-��(��$���X� *H4�.�s&�t"{�:%�
h�%d��5�aj�F���C���J��ٲE��7�:�������4��3��d����3&�a[���:���x�T{Sי#.�;��tP�\�
�˟)��,���+2i���g�