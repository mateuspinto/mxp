XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:nV���6��k��g] 0|,c�"�X���>i��m#�e��
삾�#16cH�@�(x�>���?�"��Z� 
�>9Z��)�0����b s�T�;&M��������ORM��I�SU�0��Y��T�ų>ְ
0�
Ui�����s�L5�H����DC2��؟�
�Ž�y�\�%����m�`�ͺ�r�+�~˅�ԇ��:"�����~�f�3&��}��m[;�A�(�Bv��g���rS�?U�VJ4-�2gz_P;�V�a�0��9������sQ!Ĩ3�H5z997������1�>0��N���x�F��A�z/G���C'���Ͻi�v�[��y�J�CfG"cߡ���u��H��k2Z5��B��d���~��c��[���H�/��,[����.�*GX>@�<hl<=�E�y�戴]!���ܱ�E�'�b%�ґaY0�;Ig���Ȅ�J��a��3
u?ո�\t4T��O�	O��n����Ks���yV9Ҟ�խ#}	U�D����U0���q�$�8����r��X��Z�~�b��]�����rE�c���������C�K�l`V�R�bHt1.��[�2��	�VP���I�糭�OS�\�u�Mx�5 Vc���,qVj���A�[�v��!��_�<�8��7�!�R�a��u�^���1�m������Ǹ�f$���۞��������z������и�יJ��3_��.�;/AZ�
�u�-�P�E�a��Ra4�%(3����XlxVHYEB     400     190�W5���;0�M���&��;f��D�Pѩ8���_v+b��I<*C����D_�\VTr�(+�L��+�"X���J��g�ef�� @ɻdt�ʔR� ��3�C:�"\T{ 
<OE���̄��A
�������򛘃.��J�� ��;���L�ǭ���{9�칠`�_�b�.�!'5�c�SQ��G(u�� ?�~g���:� ��/�$���1s��u�L67�z"^������n-)�H�(��I*z���FJ|������[��.�r�S��c��FT�5e�
�5��һ�2$��w -�w��|/�[�uy=Xق��r\�٬� �7o�b�Z��Y�>���,K��jmO'67���M����%�z쮭g[R��0�_����5 s,1�>�XlxVHYEB     400     150����k�S����s���]�/N��W�-<"�����9
�ç���"�,FE�� o���kV�db5K�/e5��2��c���i��$`Rw��=��R�zJ����T���)c	"G��Oਡ�"�9���S�_�t
�����&�\���_��.���029��*��E��g$�_��hgp��+w�믳0�% �-v��ԩ��G����9��sSΎ������k��8����(�egBN����#ך��6W���7���٩~$h
Y�b]�?80ޣ2ŀA�T�|��=����c�Z.nEI=;��Д�$/����Q^!��N�_�M걡X��Rk;XlxVHYEB     400     140����^�TJoW
�Y��n!Qt_�!���*�(�+�Ɩ[�p U���=�V�`[���Dp\H��������Y����`29[U��ܚ���߄2�w%�GZ$�d��K	�Πx�aU,��~�����#U��H�s�����W�*֠p=�=P^����r� ���AV@��LE�������������t������T�om��|�ʭ���þ�H!5�uc��~�u^����J<��s�z/mT+�T.X��~��$6��J�l��2^dAe�D� �XJ��palI��o4)���~;�*��N5�40XlxVHYEB     400     180�8�3��q ����)U��P)�@����̫q��������@4��Ԛ*�r_���϶b|�f�Ν_{�����u0�>�<Zn����&�K��s�^�a�)0�/�E��ʃ�äɍ���Q8^֥�L�dt%o]��=6R�Qr���7����"���~�%�Z?9c�:�&O<^s�mq�|��>(T��0MdE�CV<f�������_BP�7���M�4N�� �U+��/����x	H�v`*XV�����	�ܥ����P�,����G"��&4�V���_��/��7��4i����[G$��dG����}7�bN0酨HI���]I���k�H���O�?6 Y��1Fd�\OC��Gh���@���њ���2�XlxVHYEB     400      f0i>�ef$�S4������B�$Ƨ%1����^#�%@>��
���ͥ�ыBJi��}��}͕�~O���]�<ҟ�-K��v`	y$w�v��+�OV_{��N0�&��V�E� �`����	�ꋩ����l\��2����A;���F= [}��ZF%.P'�����/U�e[��J���-�wKB���T���ny���J����p� jV�m��ˇU&3P&��mKe�!3�c߅�U	�c�XlxVHYEB     400     150���"�˯.��NYA6��'������L�M��`O�� ���{��6���Vܤiɺqϵ����M�է6� �I��X�T�P���gF�8/�g ~1)�Tf:w��TTd�z��[X�5��OթE�i6j|:��g�CY�)]�ʟ��ˀV%!��*��� ��uo*^�{�t������C�X<�w�/7gN<��ʏ�<8��I9򸔤��#���
��P�ÓF6�D���-���ϓ��'�g7����߇��[JUBK�u��$�	+�1`���V��wl�0��'L�!l�k�)l_��|]�ya���n�w�8���G���XlxVHYEB     400     150�I\�K���6��:5\��s��2B�@,΍q��	�6��RBnHѧǊ��`b��✀�ͻ�#�
u����W��8��;:Ɖ��b"�E�\1�I��u��I7�XI��1 ������;���y''���o���C�O�˧́���I�^�+��I,@qt�[͞H��0_'��7�T�Z ń��t�!́5�NK��iN@�҉������Iޣ���C!r��}Lz�����
�������:���GaLNPlt��mEo�fZe�G"��Gm:�2*'w�𳉔���?��ra��j'�5��m� ��lR�� ��ۨ_�mDʬ�6m����XlxVHYEB     400      e0I'1�M����Z7�lTS-�5��§�AO0��LB���r�H5cѫw� �w�;f_�&�veOR(�����A�, ���q%uRٜ%ӄ�����P���ܩ����ת��poj�g���(��d��q�,�,��6$x��{Yѱ/����UA�L���cZ�'�2���
�7�K��3��:�	Xk�i�9�B$J(���o u��p����vL��XlxVHYEB     400     180E���[Q�0Ah�!���i���gM�RT�v[H%�Jm#\փ���S�_��9i�hd�=�8H��|�����o�=��+����h.�&��VŤ�L@Xi�.<+ع��$V@s��~v���}l���0ҝD��Y�=��f��=�B9����/�r��u��d6��'�n,�f����/{C#~�3�	�<�����IE���+A|�Ӆ�z.�L�߽�[�5�p��{�,_�f�W)s������I
�	�d��p��Ϲ�;�˭��A'�*˜ۃ�r6�����=J%�ƙu �àU��������r�8p�?v&?)�N<ɔ���Ұ��C���t@�0~�ͼ���n��w5�e�n��!�l6�XlxVHYEB     2f4     100� �$������$au�)n�8���s|���; "m M�z��O�y�q7�"��ͽX
����%xLZ���RlN�JB�,�b�)$w ���W����������}�~����G��#�9�y
!]��}�1��㯫��ښT���5���&[y�W�N���ӈ��$7�˒���׌��\�G'�+N]���QDRHsAkBt$7\o(Cv��S-q����ӻ��~�
C�����P��ԡ҂t4��Oq���<