`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
opahaZhnIlfeHjAnKA2ADCcCYFpGnJms4JREvDjbJFDUoelqF0s+Xn6W+bfziph8ZnEalo4MoENb
ypivZoQTdJmpSgTqVyiC0zpBcZ7LqIRrzYGm8l5fXk0SHav3DY2+V8Uj+WwJRFxLvRqIW4m//xQj
1AFgQSZJw7kMGptErspb3hl5IClCpRdx5ZAVXycqOzKxtVTw1WxmjCbi8sY7HSuFd0w7KcY8NcVb
leJZNvb3E1Jjvi+fZmKhmDZiJi/19IKol9QY5K7WBtV+8Q2ECuOPBoLHsLTTNAQdQ1aLCJw4jgNu
xI9JktBP6nhxh8zfQII1VfJoKdmejm/npsFW+g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="6oshvH9cnndMbGdfk+JdXGj3Ye2bDV7/1m/Bm9xQBVE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
XLFnnzyf+ohWGbd71T0KTozKz+I4M34Imj+CVVNVj7QhbzRCIz4fAeFLAWrVmb4xMinEVeVJ/CXg
n/ttOAZkzu7S6TobvBeaAF0g8T1iTZlLB2t29/+K53Dr8MtD9tWQ7V9nEVmxUW3+pl7qQ1mvJnvw
JuWP4i9uXdrTBaGlu3FctUToCdZTShRswYVPEZE7fSlcj4CA8MDupLubhxM1XPGTOGKoGbyRvj5F
11fDsWdhM15e2UogAN8X1P6ZLKG/ZmXOhpkCfA4UWgyMeDwofmL//D7iMO/3zFNQdA5kxeldY+zc
KpKd7NhbK+i2DPRNJOCE8ObiQkjgquzosc3c0+WFmzyvQO58jKFCnXrHhrrQOGEZbvcdx0pPayg9
sj7tp+aonn5LmKynRYItn4WwMVyCxfHK9eO1rYbdErCxFCppftz8FdeSq+Y+Jc/0pUqcTKkJcwCJ
vWRQPho4uide0uANcsOUdhIm4RyqXTXDKOQUYE9tlvf9FBPc6yaqYNkbBIAljg9OUUAdXMkEUrzd
kcFz7JxItgezrq3YrPi4g1E6w/t6K/7NpcSMZfsZjVWUfit64t0/h6Cn4ikrfyqV4cEbphdGbREq
k8m99+FA2cJ6ZfTynpf4snLl2nSQJByQs75sOfF5goijdUyca+apSDnWvL/+cS4igKmtdfmR8jSB
XQJpfSTLzRSFul13h72LMiWjfpspf4gm/u0SA0mQARcJTSSa+TpXQ+JbnyjHJYvbxZuUMd+bCZTh
L9vJ/JQ0JWhpUOTD//tU4hp03kARttwtNhV9eJgRNHXmATDPdSZkKfykEjt/je5L3PsYi3E5kYgs
iQnp3tnoHowYaBb23D62N4Ga8jRIREY6c41iwWiGAbayXjlXiC6SYvfhVVyvjj7S2BaaZcGPUiXd
ulpeUMgj7w1PmkrpfoQ1UaWaHU0YUqZpBvXHsNCN0HwtLlCLhMYOem6svzDYZ2nXA2VX0W4s/nrP
q1bnhybRTMraQ9KQVpuhugLYRU0aU6vuWptmgl8bn0JGh2ARZVqD451icmm8WHX1nn9azCUByP9W
mRccIlMgrZeC/jka0HdH7M4mgyS5GN2FRXKp4aMkQvboFLcR3jbwaPqAAOiJCnHhJEcYxF+hS7lN
1zwVo32cXwlMZ92EcCdTnRKt81znwlk3oHuY0uJhuTw5ZDCMbEEJngPh1kMventw2TrBR9IBKqrQ
Sp863NGw0XuszbONoZSKoweL8SY5bZZ+n6MvT1pQ4VO6+MXkIAxWkZuJF36HT2JkTnw/i3F95wxl
e5mrAQRzbok/FJlGLMqGNxtZ9hldx8RUGL30V7q4uxbTbeL12cRkv9lPf0Ncyrbz7oP62Q0opXmi
iOXNEjDyiRPT1D5b3E7grkJlU4EYZY4lkzFM77bm32AwKWZmaCC2psdJiUbZ5vjTLuEL6dYpQAy+
HA4dCs0eFSV4iMkqOoCqu4/zt98oMaKwY4J8bn6nuT6BgTo/LUzVyg5bnu3JO3tnJwlczYzkyExS
AmmRPNO9faK22cBF6KR1AX5GaZ8NzwikSa/kXdZzUBtzB7+8MXiYc7hwcrNuOiYLIDoZZkSoi9/i
FWbiNZim26oXLj/o9tnssaj+blayb2FT9okNW5PHDfVHevDlU5tFoQdUUWVJ6j3SgRFTVfOSOolW
mFLGIJwRB4WkkNlKsUB90VGZ+G/s4cnD+QEGKvIgSCbQMY1+bS9cD29IoiadEpp5beMQ7cO0dSFl
Swe9wbCSoHLUeOuw+9R19qksTFChE+ib4zd1+G9i7PwAhgnXl9eeYW/lioF7dYkBckAXJAR/M7Ze
79tUaT4yDmpbhX2eDMGqTZIYy8OnialCjavFvH7OuSXMa8+3naB6ixg9FmVWdH8M9kNkvvcQFZJc
JvQKChab1OkuzOj0FesOSoP2E8FMDasMgamRfoWNJTgCAFS77sqvbSp3mmT9d/yaXncY0HnVYI6L
YoTgjUFCE+Vf2YjKIK4e5e8ZJZPcmVGReENnIFbaXCC+LcufARO331IxebFOvNvkLZ6NaKQ8jd26
ZKLzQhC0/YT2b9cvI36TqkYfZNMOnbyk3SXG5qkEAgnErwoMbOCAgq5AyaWmj7Gm6YBMobwA6ViJ
gqibNLH+lyyJVtzwJPeMR7xSzQwhollc8p2t0PfYOamWt2RDTyYLdbBOypWA+3HPlQFIufB3sb6V
A4Zabv46G009Z6J5T41fRjYzZ3IHIeT9vjkdIxpoPNka3tqOKYbzlPqxlBkq3FEqSwMKIxw1UxJL
Q3dZbr2478w3zxZ/KMqqM9mFa0WadJ8CB4/wokhL40yDeNqi9qrqgwiNnXdxkfuf0jAScDFoKmqc
2aWBlu2jp9T2SxyuBF/xIlzjym/ju8K4U2ZMgudu6ZpJjFCUZ0RCMPmljIcW0xHN13BkiHFmkU9b
3PMOcHEKhj5YG4MR3eg8eP+GA1Ljl/sqRFmK4og9OkVxWhqk2SQfqxatsrYp3V0tdYU5N46HIqE+
ZnrlRnYH9E4+fn6LSx0mHNjtzed8mBSlKL+qY2y4N3ngVFiZXWHNOKpCjGRm9yg88ixRrd/Eoibs
uCIthHnXG8/sorj42iJxlUGauRSlMFp82+j/OBY5BQOrsRIr39LCUfF5m/vX3NRBKUIQD4uAIa9x
wKLJWjMU6EzrFf0+6JyorQCElPE0Ta3qrl8aHZAAYoITPDkoRZKosl0x/DvlkMvNHYSOJ8vtar8K
b+JxHLCAjxc00OW96E4Fw5UgfAdNEw2vIxUWZZQf7BOfl2HB5FIqPCWlC4cuDDVX8OE2YB2oOhek
kIoPkz+58CdoV70maVqqQT0IRBXu8N+msoRV9Vux9V7BmSR1uCLzLyf8Dz1GVH/hjwufAFciYar8
kIzdDPsV2ABBLVKag6G1eERS1DsYh4Xsyo2kwTwR0EBDEFLm/+O9kfEfwGWa/bcPCTzERSQF9baH
2ZvvL/zLa6+TSDIBfNis+owFEGOAxJA5Ju09bMEtKFPpRlTOdLD/rKoYeLPRCsPvO30CSXZuwmSm
ss/qQtkW7hvuQDikRxILV7d0u67qHLaXln+SSuBGIN3t9V30VlBMfByR9fK46wAhw5Cs0QVc7uUL
/xle8lPbjb94jMECWnb6Tjfk+0iygWD06g3I9SsWkuatfwOBXVeTc7SCj58UQbiCieERHHfG21jA
+fi8DsC9DM11qW5KCTyAPrUg6Azkpw9iS70EFB5V5PrANH9XNqhwA51AaDgLClzU7FgwHZ/VUgIq
mnI0oqudQT7phPPOSVsMBnYaGwvc+msYgUAUFdHejvHfjqAkazxdtZxfJ1iGPrljSB9QBoQ5wvxq
7gvy+j9Tr/k3+JxAldHhC2g8OC/0nkUQKiKgNiurVLwKr5MpvmYyyGOeCie9+Z++SaORvsObImyX
lYNo7W6sJnjJQotMeXqMTTYNAeonGcrnN3fOzPSkzhE/BOz9qBaYo6/Dr+539fZkXlFy5mO8mguO
1blw+nRPX1GC1F8QjQ108emEj1iJAjCX0An0uHL2WTlIXLekPz8FfDnV/e7iDyntVidE3fqXdj1L
cMDUI8klKyDIhKJOkW7b2yvtzb6lwO9wWGPxST9UeHa7CF6pqMgNxjggn+w/R/W8T9l/Flue/vZM
a6dQHJV46klC9kJV/HCgDSrD+vCgir8CkspKRSxrv2SbQFmLyiHhD6gmKfh0PrAliRq7Y60J9KjE
Ck5vdiMRwukq3qLKyXFTiW5/xj1Gu4wLyE4doKIxCIxPwHKH9yQ2j7czKEwWOvm6fsHFGjCVYXEi
pNSg2NmpQmjsLHztcmyO+csZCQlAyY+TbEnkWWrDcUTXTulMZBnQ6NVqGOFF3X8a5rp4SPbFdhrL
Z5LZ2t+pk8ZA1jAf1/ht01SJ22hnE5ta934hZFegu8VopeCcaMVIc0SgcwqK7g4b39dTZPTDS2wj
NkpxEXPeQyZfqXj+BQ4IjzoR2mRX7DcoiGWIDm7B+2b7SUkpHfq/fOl3onQO04nn+y7yfKAI6tse
M8OLueeSxWkJO/zjk7P4qRWnL0XCpABnGFCD0/kcjuTOe/wXHutcGCTJZNg8LFHp/wkLZeP8FS7N
ciBIAIExuMFiT+2/Opuggdhl1xP8VlLna+z5cpswUQGA1k0Yq5ZZRAHaWPbOCKrrAiRz4/ka92WQ
aWZWPsTBv31lkETJyRr/KnOB/b2lh6DHdVz5Hg8b52yzz4bnQpfUVMjnkfyk4hS1/mpavUl8ZGoi
5BjYdbNnSMnfVeKSW5fSqFhfczdBnXav7PSl5I5L/GH5lp7vxhcm9SN0y2jrUIdejOePUcofJ0UU
vdJdtHEoqXgK4YA/L29gLe/cBUodAEis02gKcJ2SPTit5dEwIlQuJr0HxWMHVfR0Qj/t8R/q4Aj9
ceEOXXSoa6XmoBoTjo3zGk+Nb1AOuYsfUKnvUDE2Y7mGZdXQwUZcQPSTh7D3EkulPh+vs9ediNG1
AenfPklNjpoNhx6KhmFS0WyPUdu8/CrFVOvRw1lw49+BxXQGoB7Ogpb5oBQe/UFi6IaGw+3JKPl+
cgbk5Q4CmuIceif+2elcMMp1Y1o+l+Cd7mVOe2HvwLVXh0OnINKhxkEGRxAs81mYjgcHgrilk+Q/
a/9C4lFpwJwmlTrNkyr1GuZn+bypDvlPnpK24KjfG+2yDrA+mywNWSDhBieRF6Ml5SdbXCpBdpOu
+jISHq/Lil2c0bJs0PXnMpXa4fchIw0yEFvvK5QxpqOoDD1fqWfiKeHYmf1qyJkJlYmN4yCuEhFj
JwSnHG1Jlcjw2tSFHZcaZCn9VwimVLVLX/3vb1sfGtpJU+BshZxrrA1U2tAhWJT8Srbq8HqDX0Wy
BHCvOtfhyRi8yp24LkrXwlP6L2h52Hpv2/6C5pDoyzbclVSt5y9f8/Obb74ZFIjPn/BB++k21D7o
X5RLJUgJwVaNLAgkae+Qb1trF+bs1VIcgrHlEvhe36IvPax1rtMAPbx6cCH3wN5K9K4+FkuD2eqU
W1/CyCWdAFstwmebUJV3QY1Pg4YXfbhzMQ76GqEW9ekVWjvfAly7Zl6ScinlZ9c9VqJkPKPeotIi
c6cO049bZKgtAlC3/HLwy8C/HM0T+D8r3oGYXIqppkl2edbGA6fNpM+CpgI7NCFmYKoVMHpNnIrU
LAnXDSIEa5UO7/PD73J3ah4iMxUbngu9iHjC8RbnijKPEcY2S55Ol1GpacyAdOQGCaXqDiPKyXGE
DO7Jptts69VO7KJSkJ/rAUwyEZ3HLDp6qRp3xTQxyTinPwn/roSlPCF55w+qCendKa/h+IJvY+XS
Bttnub/m7B1vYUcXqXqJ7FSCSa4l0yV1dLLCt8LLvkzpjUrJfG9P+ji7u5f0nwkG88GqRvdCtoaQ
wFpqY62zGRuu02AC3mIQEnmiAvZw7kcITeT5xPohUWsnYuM1XwAk4YGYkEjbAv2yWNqvzSeNYQEv
fMjRITow5meSmlrB+ms3n7UFZhRwCH/Tt+DIcvAsJQ4ZEVMDrVQNiLPkBfvL9lcr/r86IuKedLGO
O/llorP5UOwTaaNeqBxISqMNsD9v74aMyhV7jA0DJMB5YEzjSCqiHwI7nfEgE0r2VLYRMdOWodja
k5BtI+os9MxeQc6xSPWb/3uOYF9Rq36ene9Fp2s6Ct5xuM8O6I/V/MGZw4epC+wgaLdQU9wkzaVR
cby704ee9o/BsPEysoxOySjl32rIznFv6oa+sCoeizDzTeFCg6INdifXwzJSGF4QlZWJxD/KDL5G
HrQJ9AAlySXptcaAW0QO3hvc4XBfJLj4o/UUnFwz5g+cE8X4cuc5xEl4kZVTtVz+06os+jxgQW3v
8LX0Pe9/xlt4/sb2xrfX53+OZMtS/wx3nViYmj/u8h+7Ph5X2JhWYbHgyxi/jP0dk1FNWiB3Rw9U
EvHTy+yl6b6lD/scK8AvA3j8dA+RZbvtIWLd2HYUmGfmRmYMnuSBPmTJ9rYnpVfcj8HFGAdh18Fh
gmbjmqmtFQ0GVuwGYVCvZVOwPnXrfCiDXuprU02YXC2rm3+v1TU7/bIX+kWRhA3ASuzSYBh/Cozb
XTJZHVGrlhG4v/xNXSA5B2JBeh32kR3MGH8Tqoo0sI4E2cRZBvqUlj2A2qzGroSC3PqIreWlhilj
f/BOSkOrWcN6JltLJOlx6ZlY2nWIKxnihegndsedN986cLxmUbtooLLXZxvE+T+SqcK+4+7rlLbb
sbywg7O/HFDx7ya2Kn1ouet/nq5K81IvVu5gdbOE6ERNSFFC+cUP9dUstLs9QLklx30Z2Pwwvors
3VlJdcb/vUJ4iLH4Ro1e+Uvp5/9IpYvDGFmXck0p6eW2lUcu5IpgmNNUV/uY34AlB98nM51NxQsu
YdeVjeKBJ0HRV+wzCoF4aamUh41csWrhPLAglIHu3zKXi393HOP965B37+vBG2Q6RLUhUjNsUPiN
tZxmMbSdPqRmYjI3HpOl28zO8ehJt3zOqaMj2w9qF57k6Z65tLIGR9FOJ/jLhUKO7B3CDokdtOfY
luiEh/Ovxv4IyX79H9Ab4jYAtL/ThbDFUKClkzR6uKrBVtoF+33/eQhOUs5oh6tlTRAyLlsvskXg
eFBqvkIYPSYVnAYpJu0S2ZQrVPtMSr2AhqB4//TGJWtEgBja3A/AXaY605jZygGEVtSekTIzyxfP
l66RED5NnhZ/GumLHSb4zIIA2ujUq5L1fHkFdn5QoM/iD2ApPPmqaFnMJwZAXEFwsDkgnA/zSEbG
OUeRhAm9oNTgbfZ+YXSFY6c0H2UzLsFL/AqSH/Up0To3d8GoA1LNbmaBLVXGMKl0V9+ipsPQkrmh
4XuEK9vAAUJ1zFzRj2g+aS3hYFa2ameDT1QM7l70+NHH2fsXwp2HIkGwQZ3UAeQoK5W+rPWpWxOJ
TYM4s72RsWWMKGuhQBm70G1NeRGPouLsWxnja9A6JJ+BC/ClKaSjpn8uxhtZQQvk1VHx/bM3BmWU
smndYoyFIaZi/E4U/eBJftV/uxCYnksXSn8r0dwVAnL04bg0SP7mwzfTF73aUA+cNZ4gjkIxZs4J
PIeWQoyevTFTB0VkLd5o4Xqi62tNgzahAa86erEBYX/l9ZLm+UD/dMX8jJKQheAdg3JI5zHhkhGt
hPaHDvAQyp4KDPBxwrK+unIvVGC9NIdobQH6A65vsqAQJiHXVI7hCbPd2RFje8klF3M5U79B4tV0
rgxc7KOsHCN/vwAph9GGbaMQPoJQh73DaD93596n58mvdW0Gu0tvxEfEGAwPAVzVcIiORNILh6rF
ifqXJogkZAxgV4zpDGJQsbLiU9eQHW3XmIEdK9O+PtoyG8i0NTKvwlIMiBHaJUTjJQi1CKdiWfQ/
Tioh36DvltZUerNZEXH6ns623qnnDHFJ7OLWx9Do6b1k/vXSS9J3YWAjwLOzfkO9MrYAeFl71kib
/KQ13M9xye0pnQNb4qSS03nZLgKDO8ubEsHE21VBMTe9KK0WvvgTE31U4Ta1Du2SzK6iFOYIuYtM
SOazkZ0rC7brJpz3Vk+mncvXpiFilMZt0GqynRN/sgroPDpm2KGCKrbl4lAvTi51uK5JQspPCGad
Q0mUXHoP//kR4oBY4qbqVjoR4YEDOW5uxg1iZcfn/jJtqnlatMA206Sy1zDMapuOturGa+xbmh2r
H1F0sbu1YbckKQuca5M9P/4adVoYW+RLsYIoqKv0Sj404L5lZonc82HvTJU3hkz8qzjFnZfjFfW4
j5qJdnjk79rEVA3eHoMi1yI3onncBg2Cfl8B5J5/8JzEy0HVaxcsEeObXjbqiNoEU5TGrlYbr9tZ
iaFx2uu0p+LYV+5EIGkzzkfEwrsE+QcsQCT/ylNhYOg8eLmZtpLhuiCEb6Rbrt4xGRZPVdo5ALOG
H0+BGXJrD5lA0j/8IdnBqkwqZrY4VpBkY8H6wZxYP76mmz7hO9jL57RAua0+olygCNZmdW/jkUST
0J+tReEN7xZOvIsuYQr9sWDDpTpHpKLo8EBAd3iLIUwqHc610UVIpJpLPKNCdyNhIGrKIoEG5iwY
LmXeY/r6WM8uystRc53/p15TCLv35TLdiohZZIqPKsqz6CKAH1dP26PZjHv7mhdobwzuNRAY8G/6
vX+9McWNN+5zW3wcm++qvX1PwK+zwaa4tjBUDk6tyj2n5P5EgVfzF226NVAU6HiHrPQKAAXv8Am3
8vmsiAhQvuOSszh5JLfnO4K1P063u21U4JG5qVozoYmU3HM7uD+iMNSDI2kA1O0r9XovhoC1mDVP
oa8aq0hHNgy110Gq9YSKD0FC1qU6KZsN3iXl4mNS4IwbDCVP8Ou8DQkqM/cxT3absQDZjdEbxH+A
6U2K+twdecNPvEgmmF0yB1h93up1SlSguvhJwOZoBsxxISBjlg5aIBWikQlWKKeOUcp1xg0BMTGh
jSWCNrspQ3+8x3lHiCR8j5SGSHHRhnr8VKwNH4cgFHxs5WV4VzlMe3LDU4Co7nrYBfnU6UuI/fK3
Ks82u7XnDHX4JaQmmDldV1w89PcVRogKofvRMEmkaIRlMW696lJjFDEtEFMAdr51OJYqJRIaJwg/
+dl+J9jvRsBkyfc2sTcL5juRSt4ZuP0m6BnxQOaDtok0Laz1Kiji53ZKeEU6JmMRkbl+LwMDSZ3X
e45rbHVQ5VAk8xoSmymlF7bFGR8RrQGhLDLMl8yCuRXlKuIPuyBCT+Y7RG93ejRqZA9v7EFwimIi
GjO7tAmwOQ1L0D04TN7ma+/M6HQhaSMnOqAZZJwhUev0jDd8dhXg288E5nmIBSTA/fDoaUYy/5Y/
VRHhXVilEgSmTEVhGMrD+lY0RTbP+ACpAao/a0BrspEDEJfEaGPtDlNz7+vuLq3EjJMnhj3VoSjn
u31AaHfN5j4/EfWZYgjWDaD6k5QifP9+W2Nv30xLbi7wjgXamFSE8ZkcvYL+gYfABbNt3VG+quTe
RUyuTRPpZ2nf6er3wYQ3J3THdZZcfZ0hGUycbV81zyRftd1JFG6OXUvlZQmciaLh0Y2AjpYsOgv8
/GPItr4JxXMd/GfvC+8IldQBbAX/6cQywokT0XEeTROitUqKdpYqKRsvIAwjT2c3efXis4uYtYfY
xX0/x8rqlys675QVwXuoRf2MQInngw9OfdnDIGPjeZf5IMveM0l2HeevQ1aZnKRE5cTSGoqzR/hg
W/16uA4Ipbiqqup/AD4hAjd63NhvHR7UkhXvOrctcovuSQCgMXU0TEwznsXfyD7y4ftXQLOwYjjc
rnzZ+RNEose+2RxqmrQfn05+nP2mzFUX7f+Re11/WyTLk3Nvdx8BlAp8AjDgzPdTMpr0GHyV+7e/
bmmiE/r4rP++LsrB/8VGIpwaf4q5b2IKf+SaYOHFiijKmei41Z8D+eE5GOOsBPnvsl13BYWXUuCI
qefXmRjzFH8PSECM55kFzfehjHNyduFtjz8L3ZEbCcINRt3w4Sb6SAzswxYJbJupXrSKH36+uPUJ
y/AwqXjgLaoK9ifSfIPaeIT+pt8HPC/YHXqDoizmCNfJbwA17RDiriCGii+0IlB9kSro6eL2jDjc
wirVGBhWmnkFjGrXbjYXubJCw8/VmUH5umInehgVJPPLZLdvxQyl7hk4IKtJZbXzr9Kvtrgb/Uxv
+DQmWbVVAnmBixzhOjx7TeJq86d1mYk3slJMgwKmTfaB4W/cnnzgkMG5oFHGM4E88uafKyae15Pb
aFIGOSd+rT7DU6t8Nc225yOJArGR0aZGK/v2S+9V+4ybaFDWP1q79vdL1TX1tIjGO7M0liUcEeOX
lSS3clhCkdtCPbQVJkJ5GXj1Dk6gIrUQZGMzffeqP9N8Jpf1v5aIQT8fk5T6VZ2guXIZQdtXJItM
cZY5rn+GqkYyx5S2xKM1Nd8p+snYg8ZhaPNVhAHh4Djo3y8z/GDxcASjcKoMb/GhdyYJw0eRH/Iq
amViw0aJ82XGhnoge8+X3VIxFzmSYzo+U+EyvGIjhuj/FTzlouYHSQhl83BzqiYKc/D66Wt8zB0Q
iJqO4ETzLtbNLAJcIlZB9ddr3YYwEqk63ruDnMTNt01vN+kMfj+0lPXeX9ZWAXnnxvQfTXYFpLAT
MqyoTGUygX/Be4Xb5xYdhrWNNPtYPW5g6Wyy/E4/C3S132M2yId6wXu/pDUr2+0pERHFwMRatUq7
fEQdiaQRXwN4eWUFkWuAP/wpt4/PaA12ESPWp2lfBVnqoJNBHUeCw4W4bjKH3ZUuyUAIOjeQdRUt
7HoctegsAQo5l54NGBKFVfbA9ft9SP/oEpsaNpx01I1P39YizCScOt1Ggf4P0oHnimJfeFkShmPY
Raz2GB07gAodffipbOqFXZ7RW6/0UPPs4e1WfWGP6fVnn/uCsV/BUaSvP99Kugp1RHa7RfikLeFl
b2SbR8o5Cw8UhuKyYNxdQXlyNww7xo32tPXR2xzcfhD2vesZG2xzkBH/kPKIG1xHW8Wq8J1JjbyG
I1zEWHYoebn/GP1H06pDXd6q2YkUG44OcUt+PML5xwkFu0LjB6v6jTe3XmHVEE1tUFXWV+s/tG0R
299jAfWELng/JRMOeakIt0Zja1X3OiW5Kt2Mq66Zh4MRoKzBNuudoL32WRdQL2ZpOWsT7WqTS4+w
Y6QtqeNbl52IuE/4QIhwG+vFcy6WVBfTr4HLyjV77AKTKy7FfjFEC648yofvCOXMKz+Y3QCBjd5w
XQkAFh8NAbINOLYSYOdB1mcejOp90zpA41jeh9tcYoliNELUd22V6at8hslLci11FA6OfKYf6DM3
euH5Lfy592RKkbjZSr1kpHE3jbilvxgrKy38ctnBfll7YLZ25QNyu2uiruhg1QphGDx1OUPusawd
DDN5Xl4rwNYwcVKubGqKB9t8DY+Pj3t2UyvtUW4W5vAN+07PKy5gUu28f+9UmPnbJ9HWi/X3t0cY
S57sr6JFcMwg1BCArOCYBMjbc84Wq8N0i7nDDWexiCZVONeAKfJfZvgu0syBwRd/t/9WQ3FY8Nf9
X2j7cKzmQTsjVc80JU+Z4GqX0wOvkHHLVgIs/xQGQbXLVKiqLM+vpRKseK9VCnWvaBlOxL+kPC20
vTp8sT0QofFhEir8c9cFeLrrLs/DHHd0/UiWF2kknjJsqsz02f4olBxqEzV4/VWkR7MOPWePnj/1
8963MSpQefgNgv0L8skntG3q5H+/g+JfuHPcwmx1mvSiWQA3gc0ptupWhRwwTUneRaLfkTl5cHWF
ve0+XtUuZtOolAWwZPtRfZ64GYDXpXqd+Td9QUeGHMPuLbOHhDUVgmLkdFHt8P0ecb46NRv1mx9K
pZMb22Ohvxu6Zlg/4WjbscFqq8yDcCsFEGVftorxvTtLJOgSG6S9IZYDujG9UMVbRc22jG+mQ74o
QNgYOn3NxM3cmyCuQodw3XWzL5kFDVt292BtWSKLaXVU5C2Bp0jJMb8JCYumso0GurbBLiZUat0B
KraUpe/etWLP5ty3dbf564vRibaU8q5G1uGk3ZA5h+Bo9K3Wf3bM5BCwcdEPfRwqciCRbsL3nGn7
j/BhedFFqXff2K3cdft6hgsTzia0iq2staFZP8chGdA9QZbMD+vOFL67A5nPBSizC2Aro/3D0d7J
bY4UKhS70cjYi4TYaciQWakpu8624QqaKnQfUj/f8zdKZVR8KLMGtAhsnfl88SBUw5NLRmtL0UnU
5mq2BF7iGggnw+O2q645FjcqvNodcdsvSrdkqy9rYbVi/6AO+ws/W5WS3TuSMxdl/3XWO4ZDDDOB
JA1G/1gRJz2KaL0c+4NOZqPg83XgRUFRODdhbg1iV/yopyj98sdnTJnlaCTo3cNMwfyfGEq7IaR+
B+gJ77KnkPWOOfUatMWbZHeSMA4Os07K1wNcejaqGO52Hny3r3nf/LR0wqVbbG22M6L0CXwhejFW
P/bW24S/1N+eGu6r44Ofcgwj1V/Y9sbFHS/HQgjcThn/ekHXwylzCOnxKIaRXjX+5ylJnHSWy90n
AWhQPb8hjiS5QSt+gd3e57NB/+6amz4DIEf9xVmRcpxBF6tuup+LW8Jpl02Qg21ipc652KtrsL4V
nV7DG9WqWpb90a0rxgXf1bkjPARXswx0qFaKA2JcqXBrubvDLmwf4jYzP4DcA1WqIX05IF1Z+c0f
VcNjsLInHFk2zq5OqIIfTf7YiuqxGhURhm1Ro/JbZtM+pBNw0jEREgQ33LUWbXge4jVsden5u0aa
auGiViOS4okqw+Y5GEscNxhmZWmKYGmz9VuMoPtlNgTTu+ID1JTb5tzSwqr2Mm7we9ehagJNUecp
GyayvE5nP+/dm8+NGPRbdmfF7NxKkNQgWL412BsPxSrO+ZuI2qr2Lz5zvgS6GFTts35Tnqlfwcch
FbqUFXFgZL3efVGGDVSGYG67yTqIjfMziV1CiJ9jIPBuVczyg2t58NJ7XUsH38l2RFhdrhjZq/JT
DzDacwIRAlkLZfnp6s8wFOvtnQuQCwJq2dMt/gmHN3O442nGA396U5VYXG3km6Gyo5dW1Kjh2YKn
niwCAQd6rTtoiNLv0nXMlIlUZRzCOu1klqC1BbP2ZhZRK+m0PkhnPGsaSTalyl1BD0vvgS5I89Ny
uYmanPt6JNuYuHBVoBZ1zDdlb2o2EChFrNqW8BZH4JC9fKpkcn05r/Cvc+YHEmWBFIrvEi+N9te1
iYxcsAlONxKtwOhjRqg1TN7HMQTunbjKDZv7SZeO5wBeJZgmGZVTw1pzZyw6o1apEzhHQuNUloXm
xk/b37pPXZ++vVX8A735SILQk4tiwwLeCEUdzV9K8knTGFr4C4foD45c2PBjiZEKdwEs/kD8jdmj
lusN6QuOE2gd8RmZPUqjJaRDLRyWw/W7Ve8Qpg/FMqMh65QI1lTKhHy8amFN9NdeQL+ymkNsDLhd
cZoSz+hgBxjd4hrIeUgJHymjwh7Lnv1Vh50QGVjg1xvImwrfgjoC3uDTc60Kr3AHEmIvq3MV2Ai2
ocMFURw6j//GDuLS+y1TkiIcNJSwwiIpP3JAf1IFzTIPgqapI5EbBs0Eg0YSKjaLnaWfdtyyFhld
9sCdlaCN8xOyVnQriY8b+HhSrQGsA4T5Z3ipcC62+qEKTxyI7isnad5wJVTUrwLS0PQJWeFwwvNe
fNBA8c5oBNwl7Jz6nqOz3w0tQLfB5K0qJg564IOqIA+mXW1rSRkwFQzWO1bO4lCMrcyMEqpiKddV
vDi+hR/6x7KfDIQ0L2FpEw90HdDBpheLXri5yoYpCnxqIS5J3k78Y5LYOLtpT2EJwdYyJwLOx1Tw
DWaq05Dcu8ZStCnDMvVFHvDg0czYB+THqg==
`protect end_protected
