`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
yxh2jgKD0bFlrBYPRiiUBDARMfUMo8Zkxc5QhvFPh94D67/do+QhHC4el3ovDl2Vr7dEmynYz/Tm
T54VKnmTjJzDzumQtQ2/NDdA3sPAh3TY+Ij/AzTXZPhL2/l60bnzU8T1Cjb9ZrF3ziv/Yc1XZl0Y
0m6i7bwBh/X/WuQVZx5Ji6vPO2v0q6qA3V/HHGjHv1tQZhzLIWpr60s02NBKIOaLKK1Nx91WZBxs
qu5rS8lf1qe9T/S+YGKTgapxDXFqLJ12YHCGpjIs5tEqixYDcnoCewulmn0GLWn29/UjkqFUEcH0
TKLw6ppSpml/D4aQWmDyqfU4WatUEYLb5+/v6MwnPSgr3IzL588iV0NLDJU0FxsUpZPYw1V5rGHE
nI3Ma2tJsVBuL2MHY5YIusuk7AJD1N0EMyoSAoR2LZ39r2VQPvguTB3OO2aVx7Jxml7cJD+JQWIQ
MHHFhbk2lMSzsTmiFQA75eLIEjuGZqxT7eaMTzivqVLD0vbHQJdJ4lmUsEW11PdgkiOqrcAXxrWj
+6JoaP9DVPjUUzCikuH+WAk9QvVmOa2U5Smh/qKGsfuVjRO98sCQowviMnQe+FuSfQWTME2eq4Xx
96W57z6Dg0tuTQL80QYDE4By/ExYlcfGaUC9+El7Ti6qFOBbHydicafHKs/xkT+6ae67BdHXvrN8
rZx/Q/W33xE8nW10gHUqt2d04kNktOF8z3gkcM/exSV+Ji9PKXh3m+DYqX+X9D6Hkh06GmK5loq7
f4Zo3mqMTGD8SJDUWRrFK2uDUqyIe5geIVUjmTw9yEMTpwy+pSgkVHWTSNKiuyftH6s3cLOm5OzU
SwWeVR9g6CMXxnrVpPZ8Lqa93wuUozDrZz93bnAkQaLFDi5cQNWhEeE5/8taXu7eS1IOu1fIFIKa
aPcG93lL8aqwRuUXCeXAIrPxnEmD696xT9Rra9Uc1nHNLxRG6LQBBhxQ2TOgwIDTRiobD+zlRotH
v8L5YcjiO/14wAwkkoz0875jA0HqLmjI63kvoWBx2QBR/+L7Hr9oFPCOG8U+Pi8y5hfPCRk6or0x
VW2CHEET4oM4Dj8FPmN8Qi8Q6ss1wSUeJpPWpC6E46ttXVwNsYgDyMBEeLNRdWqi/UDU9RH8kvhi
T17v63gdAuA+brSIujLYVSgviO/F/Jkyag/MrCpJqX7hf0wRCVR11XLhE4JZh3ND6B4HeiVypTH4
kZGQvxEIJizGTnjn+kwxEw==
`protect end_protected
