`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
0USWSUGxovGsyBJteYpEodNM9bw1h1uV/JAessUd2LzJQtEMuZMDt+QZVvkQ13dUeTRMH93MJK6c
ABvdtuiJwrSejL5cMHFtVxf7sQ2+SXg+Sl/pHV9GUXI0/xUN+NBFIv+sHVG/47G5iDCoVve1HTXc
Nm79iAjVcbP2VM+87cOpoCTaikCdOEfNoLwKcRJC1uFjXwAwJaT0gminRgbgBh5Ka+43yAJBPzjY
MeX4DBNHJZyUGIbRw36Q0I58Ks7gYjahB+vV+/PJbQXK20jP4pfOhBa5wZjZrdRsx6d2QffKwdxB
2B5b/ICwNLCGEh0Fxzngz5KZ7NEbAfKve/AWmE+wjTcGARiX1AECDkR13yRPwNoKU9W8VXP+LOhH
u6L52d8+qPn501PirBkMKvFll2SbnJqs7R6ScfhZeYTRgvjei1phpFFLsFLYlv3I0muKcr+ECumx
lQdEvhMUBhhVG6dHJns1DMuRhEbkdHG4i3nbwlezJ2DNUEpXhnU3VH+GD/p3hyxKWMMEQVuDutf+
etnyepIoD7shOe3ZsCIkcWqgeHDkMdzyPfCSvNXTdx/nhGT4nDLSzUbeU/odnZxWtYx/1ar5hCli
SV0Z5Uw5aQW0cKEMx5m4MAVDEofPuxm4EupJtnKyfffsbFQ9/yf5GbzWY3P16h84ij/vLj9WeWsP
du4q7hARZPHl9KYWH63CRKnvfJWY4aUdBpw7K7KKesngkSyEK1G02EAmSarKYMtl+8IMgH/IvRcG
CGT7Qt/NTynDq4vDyHBWGJQ9NbJ+kfaeSngGmhUkJpCXiXqbHVA8EXNiPlOhUdQDmoTpyGq+M0Pg
6yx5zo834gNCsXxnE1SE34l9HDppgbM/X1Xm07sIHC2cYC3toKrxHS62srJlhm+0tyE8Dlw7pe+H
6iWJyMCR4pPcx0nGZGjdMHnq+B3lE8JM0gNEb7yr6zRDmjoFwjVvTsWJ+Yc+v/brzn1gmZwNeeOg
1OO4WFdcbMOOeH6lob+T8IvNE9AsZ3PphScem2ZjXIi27Wva6h5FjQmJuM+LalRZhnzluCx1xBFW
iiXk5zo7wjYDD5yMNcxZe3R1B5u260VMdVRwS2piHqTFYogPx9I4ZwUiLRmWNW+vY0QbXIA11xMs
b5m/KNrPEt5EBl52sZyYrAFTK+N69jNLNBf4a0qkJYXZe77MHdlzrrSeqD/SuWnf7SRl2sm8mKt+
ePqds92PLXUEBOjO7J5XLHIFojIUl9fnh/3XH3dqEYQBAfZ4kqIgW0Lul1PnaEwJ9IDIsQ+QhD5i
O2CL7rljj/kACODjj1VNWFIVyDIi/AA0l14uIQ2kX9e116pBpVavrhDWYyI+YgCBPj7D4XsCo/IO
NfLR08yXvJfeYeUkaC9vwXV4T6jIEbDQblOhvp654RyAk1LrGDRs919JUx4pyLKZv0/8k0XBSeTl
c6VfwBNuC02Gj9wN0TZkDoM2N/qjxWs4FZUXjoaQtPwQSLlx3ppShenm/whiWFCN48F7mttJe+QD
4in0rXgAx67jsvsnWtqIEsf5svt1rUR2MuFwT4lx8DrqZ2CGuhssZcHL5yxuJKwP/VbwclqW54vp
9gGGf3bW70041UWzVdxZxIvoAZwjFsMhBGgoR4zcdh6qsJMkZFiYb/v8FOn72G8j33aeXQsprVPK
vx7Fflh/trc4Y4uip2LDIFSU7/s/pLhnPr0QEbZmSVTjYvz1bjQ6+FgxatzOwUuywhKsxNPVOghc
qZCtKLzAAsuB3k/wFEgLKEjCJkNLVf4D7johlqTCKvoqC5bPeDzxIVyNt4lNdel4YvryRN2Ds3Kr
0BoobD0jkdMHvoaF6uWwLRMVq0Z0TFukHVTFAZnpQEEjTz49CmM/WuxHRVSx1C/BscReNH4GFR7d
ZdZS8feUBMHYY1PUAuCjgUKjUoPxuJmJ9WrJ12usZuMWwqaqnZYmPS2227+ZiZQ7cyEr0DPjHQVE
dxx8Y+PwE0g3cac3O42MQ9fJQUoiXHbZtVB+Y+z7DjlEIuwIj5zuftLRuOW/TZTkUzZ0Vhq3lMYz
urCO3r8dwkLKSTStvuJjyN+c71AA5KGcXsi+//yYbXZHStZJENh+DNFOIWmSIbdDZzkT8uqnJBEz
D4Y7UOxTJctSZdj/sPjc9B+KwN9EsAvyzis7y5z3MMWsGC1VaqaPAK9fx72LuOjnu3iPuJc5Dw8x
PTUwmTHpLQ8t0+ckCOSb/JGipA5Dc4hgsOFvyCUbl88f0TWzqG2tBjAoj4/VozhEDI4MQalFW9q+
qa7CR6hXpYLgFhQgBLNVydHNEuKdHqgAaRRO043+QVg9TmYH3NrSt5zrAoxtrISyr3Ddj3dz3bjy
8eG7xUyb4KyECITKhqTzOq9VmtC9LrgJOgQV7dE5Iw00Ys/vpngKxv9m+pH2P0or32YmQU0pXq49
CsUsr1LJzglKL/dBJLqIPA7gk2reqzw9lR6K67UkjaKvIXKrJkPflGVv2Y+RoxyaYx9cZqPkhsDV
FEI512is+o6+WEeYIPcc4IeJubSrgzPxDVQGuAtNSBkH/nJ8TlMkXbfAiE/tt8Xn1puJ2GGvyRVC
8rArNFG6cDbRhnt5G1u6LdWdkkh0d469waWxKeo7inBqtjzpKsJ04MJiz+UZ+lsWds90B7sbLgRr
AsqocxlwfLKFGT1+ZnJSwCjSg0xzDJa73AyhrSRo7ECPBqccQVxtSi90qg49Sv5gF7ZXUgQ+rjNq
BjxUfYgycPL0WM9ozIUCDZjY2p1/X3FA5gsjgZdzaQizHdsK+SdO/q/dAretDSJ56rA5aYEOmZN8
GZbZlPy5BQUvsgOpz1gNFaWMe91FkCIMsJn/+jA2TOB24XLtsXtNRFhDXEtGE6gTsnxbYxGEs8D/
CuF/IhWloCRLG/Wi/jSUVdROX7MIOddhQnc/4iOVnMXwy5KsOgK89tYSXjOaNhHL2XHD3T/81ZJY
NBSa2m1ATKxh0IO/9hALCiuOcPi+ze01YmrRTUDui+WKgSBNn5XMzk4FPEb8W/DIs3yrso60IrC0
AAuY+XuTgnL3Kb8WPbALshNnEuF7/zqmZt18jfCbFBcjGT83gonom9jZPXC9lWQI+hUe/LVArsRp
5t30OjJ37vLetIitdBzbnWaiXzapLoLXGUG2FjL8t8qXUg5NhhK9hbJ2N+ne/Ga1WSUuazS18YeZ
C2DpYo5ZvCjHoomrSNENPoqDLsF24er5v8Q3clREfBUOBxFNQZjEBNoexAoOD9GcMZV4MaOjpyem
Iia6622L0x2+vEipXC+g0WAWRkzWJsZEPOH+Fyavqp9vkcaF0FrHg3/H5kGGcE96hab9tcuNWwaQ
YAw1HqN3POTyTXduK9Ijtcrk6DEVkpqYl25bpAXP7o5kZRHtNq5MrPEQXegaYNsRBb5BzPDUOaez
bd/SWc47AQtTLLcbHSX36p/kae2FmJVTnYIoeaMQow+9Bqv6hZVAz+Gh5UFWC3o9u5SXNoTtcnIr
7ns4KCQRz+SE8LfC0IL3Mi+8t+NyNgCmmPSYUipqmD7lOEigT1sHPLCpR0cWmdARC6B6m7fMnI8X
7+nz/F4qUUi/aR6kHKGV1ntRas83rBU2rlde26UhLiKMUd8wNqPOzOwGLD7kl0vX+Yia+mzUzScc
yhoAzphRypej70V7kugj+JZe4RK+3hOD7IzL+z7roU+RBfUo5MbNRVy2KvizoZJVmwtmbsdZWMmh
NnZr8XibDUYnu5K2Eum5d/OrsBpER3qoaP18XF0qoL1IR9OnOeu0vtZbIebPZ2cG5Fosd1KtOg6Z
LUiBqPnptGQsQBBT1URlqekHJerHr72dIolqzvei3+CYc7hUQoac75S/p4KrONOQvvUVkHffE9No
SEOa29urDCn1PwN9GhKfFHY+36B2o7PLiUlALS46nABwNpiw1qQ8z7xpBQx89oe5wy9X8hzYQmmW
BKRR9Zor0LXAMQs9zLNApjQyFjdZ5imYsftExcCjgsMZ4H+FeAPaBlpPgXEr1JHTCxVyjo21vQXn
Ei9OWz5l2C6BV/naY3Bwc+lA9AvlWAua7bMRgoINp+wT/66A0gq+UKcXVNp7/RcULetOhX0/OTVC
QIuZoervrneMbLB6QvxDmFNKsGMY6yiakw0iuVyV2dsick5WNDW/tFHTY2izKvwEn5q0ZNeBBaC/
SnMHM8WnfSn4qDB6pwt+YG8bOPv2BiF2w5rItvYSipNkUYpDM8O0FzqLIBA7zCCmJ/2kRyF922Lt
F0nySuuWVlS1U5ZrAETs+24aLMFhzX9KJ90WJouxHlL7YqBRXxeOVLISrcBzN0u3U9VXv+2je2fW
XdIgCZbbfGmPblGXritcNvydmgyFUDD35D2f2fnuxJybqjHD7rioTBsHiTBhZQt3PShwwK+QhsQ1
GBoRZ8lZvESUI0Uy/C01wc0E7neqtG56tTxP6z7e6elciMeHd2tid63auEH0NQC2pxMLpyTp+ZOl
cnp3Hk0f06O4dPGwnfqlwKZE2tyNznoF35EuxJ9JBMA5ckm9sxnn9gFqDiHeZl9x9u9N8+2Z8hWv
JaemPkAW8w6nCPb6cAEmeVHraZjitjDA0bsPVoKcBw/nIvyjucwSHVGNe0kkG1Tqt0LnZfjFhzsB
Q7ZYyvatI1dLTM0aU1z1GTazprHw79hLWLzjTxkJnSbRoSXcO2CY+mzQbIm89CXYubydRasXFEyk
ppFmseP5MI7re8dzMbwtIUHqUSIXAC30ogi8REuCdeIqkopt3Urd7xzP54SevI7forYDc5H980T1
dawAVwP9pBV4He4WMy7h+aiegB2s/4hzgws8zdF5+C4nHV/sWlQltkUJ8EFqZHuPVcfxauUTUqLV
eeXnii3NEFlyyCv1c5HqA8fx03GpNLAmCQTn8xv3zSYTAx+gCd5t2f6AUEVqjDMloCU4/a5S5Vup
wPK89cG9BBpEYuE5d79DiQCMWt6IAMYmiFkqvtzTRnbgXWNvqRn5IE0xi4Tdml6hiEl+IyA5sOmk
Um99u5XhGijb1OFENJfThxuiJRP3P69O4AChxdicz2JUePOSK04b9RJ8l5Q8yxLKgkh2HLmxsrVY
FGlBPD3HAaj/ObN5X4sRccVRl9JchE8xwNcX0D+Yghpo/BVzzkxF4mNIATsbkyJHPoxkrtQ+xQzB
r5S6L4WQAtr5u7VMY26tuymwzewCW7wiDv+HFa1ReWK9IskZX+O9L9cfE3jC6jNpX9TGFSJvAsZv
kfej3NP80uNAUUwj4zRJgXFvZUCrtx3FpZXdDsyb8nNbIH7DDeOyUQZX/gYb5byXZE/WHEn6Swxn
nlTB7KnTakOLXcob73HGNmupW0Kpw81g1TX0ka4u3e+TNNDy6eN4v/RcKXhbEGgqyCaxRdEkhphI
Ob62kB/miiIf1LNf0yhoUfJw/VBCRrm2RzsZeUE9zsbFqVaXYLnmM69n8t8SBLfv3JsUleEW2HKp
zSJx7vviiiSvq5ArYa78aFCMzGg4d393Id1tEpNOv/uk4URBPOR08rDmm9FOFfNjVJjGGOnK//Eu
LWhI5Ou5FT6XumbyYuspRLzRHbcGIvIudKy08DhTb8fmUIBOEbZWe+rdBr5AbeWvHtKzrppnZVjC
FYsaolJpaBWdTXPrM30VcU1BjcpqLUtopZMeSghVcefxkbHiO3IvSlEPoRE03TsXur+3kPkLr5K1
UsHWwwNS1RrbzcLZwxbKCglRsYgmSyN5jPCp8UTxVAJ85YKriPv2H2fMSdNmJirZ0nfbbcDArDHf
KCpoqtbYZFZDIa9fj7Bd2opO62diQD+JyQVpqttY9Om+tgTNDgneSMPxRCurXWgoxu2URg3ZSO/D
0/ZoyaR5/iUmsxVf0bdLXZCFrMuj1SN0IinF3juF3SMCdg5B/EGcJQtccWqT3lcxBBjIB8PtUt4y
sJb/uEIbYDaKMoOVCAK4A7b/LKa07B7Kv3nZVDolWCbA22rraqrTKp7qqsZUDtfTpJx8ukQRldQ9
cBrfy095bSfUOvfzBhgb8KMx+kdExHjv50UW59CUeOs5hwB4DPMgW+X5lOVdQAagaokSDDfjpNvc
8UUjOQ1I4C4WtxiUT3jEqdmBJOtFAgypz2kTIsv0yIJigRztdb4OMcc5j6VFiRw7uxDv3lsscjgD
ashV1M7WGF2+6J+pxTrFgaIsReKbqV4ktqUKBsMYPjOcIMvPssoYIZubSBk+66I8gm33/pv48SHj
/IOvB6BqNk9At8gKs0AVdj0k2nABf6cs0lXnItXaPxzemf1X2maDHSk8EjZIyCvRwK+msQ89vurd
UGQC5OvXtG9X2oe/3cB2hs8EMG2c0iRaGp7bkoD4sKsjwXaCNUqYJULOfOiXvbISE0WatvzhZVKD
OOTGBf7bPHmIgQoUFLEP7NR9PugofBMjRrA5gQRUxEbhCwaVo4hKPcaCw5CDk7m3YeJv3w7LwK6i
mpDbm1Zp4VX/a/cxcqwiAlBe3eO7a+Xqfdk9Dpd0LUrpzA4riYp5LmVIBy0L2xn2nei/lyh4yfJz
dHawJqW59tE9IijSGVBKRUYMfx7HJ4SeQOx96CPP0xyMRtfVNwwn0b1q94huMspxOEKt6Bm0vhTC
At0bPrWsHcZ4lhX3kdm8meA8Ep3KYlRrIb+eupJrTlfRb4ORcf4qEXDsxz4Fu2tyHCJMvLXw9bI1
GIRtC0yHxFshlGXvrSdUzFfLEsam2/QTSX81uoyqwkCX4LN03nNxCa7iGZrllX/4FF++QFuKyR90
DhdHZBJct4gdPiJLj4PKdYq8KAdYkL/1/ntTxrvxAk9sGng7GUTGCqkraILslhIAzfSsewQoJ9U+
1zraW91lmvr91RLnAMW6lCr+fjl6IF3i4ss0kScM58eTV75Uhhhqit8z+pv4jUv6JBo0RGrreZd9
lqXKYGNXEYqPOqjGNQbjRfZhXWv9fB5GrMH2YVqhrvgDOzn3qpkRj67Y1XZficVXOjeDjbNlBZZV
RLRN4KiBKXxL5fFvcOSRmD9pS0T0WNdFyLrXhdwiYWDLiov4b+3ED6AlHzi7RHG9J3YyJ1y12iaJ
AAB63PZvyHJF21C2fJna5iha/KB71uMYXJ6opKa6Xta/NitvC1Qo1af4ltGhFZ//aGSlYAvVmdKw
2kgj2eXcI7ILcD5ZveE32FYTsirXXcbnW9Z/xgA4lQgZsn33oFY9j6vqpGhoHpyIyX11LuUWDkWS
dEXGbsMyilERNSdWfWwegtrksfq7zb4+B+As+rkg2p9BhTq0FNYYbFkDfJqmfmMlBPwzP9J86l17
0eVA4ZFqxvmmBhFOF6acJmq1mH4+ouRgcRIE8J+6rNZngdn4OZbFwVMHLrkPo7L/ZiZY2d/P9vRB
nW8oV55vwptS4CvJH2v8ZhDHSIpYTBuIdTPbK7Zb5RM3kxTwdiErwTsD2TFqViv5QpGlmReTJgui
gSpz8O5sRZJVSMh79+tDvHW11XCEZRY3zKeaiOSA1H0CabqkFnqIFysSsbfiNnj9VLvP+m0Ykbae
f1TISswkaMzXMko0cccl1YGFb15knaS7qzgc1GLCQTolGnD0E5dj7Ijia4FiTLPkTnB5a4dh03TI
k63AWkbN61Vdv582hLSF4FkiM9ax6MuFnrI5yTwLTS5bnqGjQLb1pJiGy8kx/JGIFm7DfcoLdLos
RxodWGIoxu7ZyhF9xYN2LIZUExfdC6XpB4MDhkaRPsjK97xPHrTYEaL1mUxQPWXq2TpLycVSKGS8
Fk4/bN7/NbIx79yaApvJXXtZOt90LHGMFh7sAzbArFuN1dmbPa0M9atmYjAqfy/169LAcUzrsVXJ
+Xfz87b9nT9J3iTvqQO+Z90Y3EfdPaAMPiia445lnLwkYKVR8zq6EraaKwnvXxrqX/fvlxJJiGpp
OvrxW2ReNN00eHsb0HFxsOWRzLVsBwxwHkWusbcm86RcQo/ILp3/RLc08hFw/9Tp5Tz7+A3+RObQ
0WoVYGKx6MX4aFYeTHKowrkUeLtb1JTZIDzLUzGlRQrq3cBAW7IiF1zSNfBiX+bHCTVpnKOuKP8f
3fswC87bP1Anr4XDqlzLswTXtgeQTwo+IAYaxz6smWleoL70ms7reQexx1aHhnjyYCpUIoZ220+8
H7QpY2h4Uacy0kVVoWkKulj+hN6XuAc0MFoRPQ49jvOFy0UvUW2dGqiXU0rBaAzdgS5ilGkFLyK9
6hGpAsuNxqxZDe1Xa876z67z5lwDvWuCGq/vpJU1rkIkn3bAo2NCKm4Z0bYjnyjwhvRp6vTQ7LtS
67oq+1UsnBTlWwad7pEXfTraSwiAgLdspU5MIjPIdTqejm+s4qGIP9HJRaEOnHDVJmi0FPZGUx8V
+ZNG+Y8arr5zGgGo4iuICdFcvyRUMoeHAbWQygmEYkdCZUjF+u+pQY3wHgGoN8GdOODkDUKiY/Vf
xUU/ORwAreRo26DE6nmIc9FdoyfqSm+OLoqIInKw1b64G1/QKXDgeskED1qdXYLCzsSzIsO8QF6H
BzsDP1ayjEudzPEKB7T4cOOP8Dx/eC2bbtxmYXI27hPk0EhU4VHvjN1UBi7pqyvBd0URLB2ZD8UR
iIZfVWcVdHopwi1/LvEHj7Gb6px0yeKqx+M6+KvGMusLwMFt+UJCQgUgOGfebCIraVaxiLMEZ5kp
LO/P3maHpo9ZLcq+KnqooczyJlQEecPN8ylaP3RHROe4rXyvj9u9mGPKz5z8NbcDveG6El3CYMLO
Bm+sN2EgKoMXckEj4gdKYXQ3wg0NoNjZPUZbG75k1ky/rFiUEiHMoMfLTYe7Crhbn6/gdieL0UiM
cQmYtkPf/DeBQXTG3mRzDsFhql84N4DbM9McCpBVoCBkilm0VOPD7WDb47+QkzN0bOvikvig6LRy
OAOJ6SDGS3snuRzK3HvStUOm6P5MJcSAcb10aRzdhMwef60EhhG5hDebq2KTJSje81eF+lisvOIA
m+HIxf4I9bK0Z6+whyPUP0ki0GiKaVbOnY3VCLLRztyXokiRUgmohw0PeORDPabgHSyKQAHdeCy5
pE+AKQrSe0kpXs5v+ieU1trtqKfgJ65sXkXG03EBYZ/WgDkoZBBp6wbX5VPO+ZGfiXbQxt+01HwX
wmYBG9wTlsO416Lfo17Le6OVZCfrHxHpFKZTAX5QHcD6/1+30mvnOUmWECdg3UWLeZBC3DqRHEGN
OH11RBrXTUDkjIzO2ZQD1UxkSTO+B0KWyy9UJBCY8zLw8+132/MWnvcYlF+o7GSa7XrgnW1st3bm
pV4ZdQPLDkLZRk3Mmh8TyqJtoqEdBeUFOlKqE41Z46AT0nuDZ2KfOkpMYlAthLYhNwmrYuNRiH7l
qQdDe8XgGYDRPLPg7sddUL/mFZXWl3acqHcSWvpTEAmkTfKtvgfxPIOcmvgkdgjaHNCTNtqOnYdm
NFt3lDUDw0AyiYLB+3jMgUFaZW02bKOeubtanmeyNQbexyaM05dvwpPm/9zqRZUDSZ9+yu9iI42c
mtJRqZjHD0mzvfJvy3+BknnfNAkcMbKtnkcH9i8MURSW+ySTBvZUkk31sfBUwXAh0jt5dGZBs6fj
6n4bGdfUFindjnt/ctiGVaKbmdcSd7EsBNjR4dGX8Lb4jdjN816QQLVdgi0HK//0Ywziv0igOV3a
Q+PGk0ogECWtZRHb81U8qIeeTuU3qO2wnyFWC+a+MzaXa7fL1YK5JoEG3iIplDLiD5fKjx0pT9rn
BP4E6/ucpEDsPA/4Kn+jdQVhFhR/LDt2G/OuF2Ur8evt/93COE6/Qzc/5OM7Ri3OFsmV75A61r7J
6nd6pSCIASdzg4zmjcXSTegHM9tU3WW0dn24lqxGJudjB2Recw6P3YBufp1gyNB0p+heO/qvQV/d
QwiVDB64i6ne0QiveWVUYUqSWgsV9dLIFBdTVMoz5sUseecDXwsRFjJJ7IiRmldJsGRX+1Bsaoza
HkbFhvrNvrDb+gv5LwfmaYO8FbuNBnmOaeMUtRaPpWhVPrPGmVTAIgenBzf0ubK1VGSKGNsHbkyN
SdSw/57wkZIRgT1yJYHLmMBo/nnNvIOcR+Ab/kqdYslOoKKl5VY1plrVpz90doQO2NEwVHTi1Oow
SGViFkIznhJKrpvV7iMTQA50JNfHoCKOWEZpX2vrQNnepxRlSDFbcTV4Gro9BvuwzLhJ6ZCKPOEX
8wVu7xOtsd9MX5YvzLoNmqXqCFDeBY2dT9jyaNpIMygaSEVYJBjILBubeINBc+9xGg/Nk0WTilEd
/tHHvwt6R8IJ/7WiZbl2LtPYs5eFLXCZ53ItB+ESFHNEq9ZZQp2D3o3eWPGzS1OmWVKfH4z2lbsD
oi0Ep/rTV2M/5zDosByp9rRKQwLzVucuGNyoq/cnsVm0bA8egyzyMPcVcZzFz0u8P4Uj6vnPyD+j
JhHnUVbTYAajjrNqbtdq4ar6qr7j6T1sQs4Pz2dnItr5ZFAVRmJ+EtHpvJKP7oMQP+gmRz8dYDqP
yc9qH35EVCwJtsc5IhAvzQjJLJWMViECj4rZrsftVhR6+uu6MVHFdvNpHYcNapSHrfSKnu9Ucvkg
A6gDbe/BnzChwIUG+grjuqFQ7lOyiOm+R4Wg1VRaSYULt3vTmx6PckIc62rSFr3gJa6cCuLfjZ7y
2nY8pa/d1s2bo6eVuokvEqSKwmYIeLsUhS+fRNFjPW+byArzxUqCdGqNIfXwKR0GlKYSVgzGJg1+
Y1mXEmCEa68q+funJzxmrVzD0tLqMd0JjsSV/OgOawb32sGxajdUobJ/G0qtpyyMRbpiJzh/JCq0
RSFFZsRU6opTOfxOkbDXPPXPPiail4iyO7eZweLQWGLoZx53WjAxGg/cns9b1PplEwWRBqiqfiX7
T6EXjs3l1ywu8ERFXESv5bdN5czqMfRFNl4J3qQRRba9nq+XQWzhCuP5jiArm9Ze1cWyVQ5nWYf9
NdJP6A1f8klfGliL9gf5sWGQzFGjKzTkxPlLMpYFAtzkn4pAuOShyLadp2UDsU0llwCMNVMS41Cy
KJMV0S3Iu3ZC4fWT8f+dwMSwsKlQYNn+bQZv1r2pvHAPuWnRLX7DshfKzS0pmkZecjUhhbfTuJjb
QNj/fEWY2L1XxaMG5DccFT2wDc0akZj0Cs5CVK5MCmXIQM/NWCCmC0twFiKDWXT9Sb5BaCumoqu/
Q7Z9+0qG/ydzVG/Elj3kHRoj6tJMdtVzN4VZbcUM4QLuUvzNnOKx5ttVIQ20Mn36HUFd8K/OZpa6
5C1so4Fv+QwYqyFioPBiWajZlHJibt2HkrEX31mkUHmVDwcWztcuqu2z2FfCY+N2avioAOcPvoBO
ez960AFPEL34dtvz6YMIipP/VQpHVpUm4lTVmc8eBurUs+0I7KDRPyuClLr9ew0hLStnAnmgIdRZ
TV6ymPo//TivuGGkwQAO62L6XWHN1LN1830N0/Q3GbaLJLq5RknVkWGA81yttzIbcFxw4vAC1HcL
8MLVFmwc4LF4kc4bjXKSlRSKIArWfV1I2O7nfePJfy/FJ3gowYscG2C5WwG5zkKeKGYZPPhEpgU5
zY4ceyZyN+1dJK4eStlQn9B9/YD3RD6HbVRlJquoaGYILsneRux+aP6mBJ2WrRVXyuJGEIe0sMYI
ERQTRP+cgTQhaC46lvjgIvqCOoDWgejY5sOj57+UJVgen8dOyX/8gaXhrqbgyHpjgTngZEWveS28
BnGNzhWRnbKq+1ACYbPkE6kLuVvxBEjws24eaVOEpIWsRh2CnfCJZWyqsc1pmwGZr4NbxAdKKQQA
MBRph8dAhl2JCfMAAjlEYhLSCsSyrsKMczUn4tC40dwU173Snk3hJDgxUm2kanGmOO+hgMI7+Spw
HOsxO7ooydyggPNQRX17kwod8P6QQen4HPegHv+VqFGgUgjFwJEYW7XUulkCu12PWczClnHeGfqF
cdSxwI08M6CINTdQ+LbaiAFvXUpM3oumJhKnRZZRUgpE4suZ1ANSFwHxvSDxXXMhWa88bNz4XlYf
HjZt0YMt1w5xScGuVlk4g95hNwOpSHnCqLn9w91mLS4e4f9CKxNJsr9sX6iObRm6wd3DLXcRUueN
jWgQtB0peJ9YL8OuxDLrWAq4MjtTtdLiMqhG5oUalxLh5QkYjfiVFm/ZjL+oBDpYSfiwF7rWhQx+
AFeQZAd9WU9Gw0zBx8dGue9+eaMIOlrAesWOYYgUijO1ujKCKmSfmL4Uf81pE5ksoq02yMHJcjqh
z0kyULO2afcZ2WwabNPWkY1iSvXJZKkceG3q04s+rxpZJqKD0Y2hSfMIF5OPYQ7qTt5vpX/J3g8/
WREik3DqQKA/Uxaw8hABZJpKRi0cHx3wcKM8aM4+9DwK2bQtwVtP17qfqa7TLgTp9VFug1Wa2btk
flWwyl+3FLxpFuxG+1ZOpuJousoflr0bW5F/t2ysX1xZcL2JaBLaamqprG4yEYxBEkgVf5SfcRnh
ULZVMarqAu7q49T0sQ9vafTu25vO2m8VmRgOrLZ8ba/rSlV8HVJVGCd+S2/3DtrUIoK/rCkThq6E
N13KeFUTizjyn1j6EEdk1rJs8y1o0HaHGde+zxaC2Kc76xul23VtOMNdD1nJxEtiqq4756Qsv/eB
c9VqX0jLezyh40T1o+QcoXHOVbp9Ke9pA/OobOF26fp72alXlrGO7EQVM56PAWfzv7iZ7spswzt8
JcywTgi4G9P78MZdhqoZslF0HqXRW24aOPU4owJ5eF0uBqMfpTaWESaOCNee0WSUej6DLFMjhG1K
llBOrhRVh6zdNEPym7wGkc+QfAo5Ff+F7aAB32kRvOFXw/qncbK9uPKoyOtcp8MGZkjHasdyfsE3
l69L97d/MvNzFmtd9PJyJtqHVMeK+D/WVvlKZhrJatP1QSvguYOCEw5pHBa7BjMHrWhvX2a/avLX
9htUHe2Yspsb+a9Zt80pHW/ECIkbcJtMm3ukbw5axgFX7XG1GHMchP/gGo3sshaRy2UNah8ElaNL
mQfb9IOvea6F79x5r4DgtMKJPLxWQE4vXmRCaWuZdOcJbipfhv73gXKev59dVW5DAhYvKIobLs+c
qUv6Fbn80iz06DAEgp5MZh7wpAs0yJwM6fQJBNc54lHisrY3X31/xJx3pKuX8b9Pgejc72LKU3nd
x9UiPRgwRn7oMkAJO0yuImte/e/XMEz4fxRHZcDxGl/LVqDy1Xi26HpIbp1v6T+n22EeJNx1O9bP
9N9GDyS89sITfGBO7bFyQGV2mJ64IwzaQlGWBWxcaL/BMKf3FT+y4YF53KPid133szhc3hNO1Fdt
2d21mvSQuA9ZhHeeIuOInBh7mVeJRtflYJc3xaJUS6Mkzi0upI3gv7MziaBLGIT/zAYoHbL5RT5i
fzGYiyXGnA0HwTNA9JIKwCuwBbk7cb+zW9MsaOGPoFsANwuhQdo7Hto1duyoct4j6dW/qnKg6Sd8
x8qpgLTY4Va0Pe9iE55PuQ0OzjMcTVqH7zF2jlPIW+5d7qaPvTDZXHAG6e5vltfyt96z12GCYVAU
lH7X43p61UL33mYrXr85qU2vr2o1iHz43yr4ZHNeOPAi0l2fb+E6Qw/t3b7pcCJX6bCUUMU74uJj
Q6whYf5T31BpGIBjsMjpA9CJCSZDilfxXim2qq0yBua55YWe4PnEKlpwb+BHMhRE3zCFglm2HrZF
e3uCFTJe8CWGphNbzLe0J2DJFALMXtx9DnfK8/HhIdeCxDc2xJTPSx82epD/Hh+BrcfZQFo/RjGL
c4JHw+0ZSuxMDik+eP58MAGdxUeWcSJkFtgqPGXFQHV7exeUCSptC9YNltLfDgpiImZfmCC8ql6d
M1KyepAPoBz/X/dNKQYl+0EvRqmaQOwhyNWKD/7Vrs+ZpjINqGfsgnqILszUa7I15VqkG1NUgJdm
m4ZbTUY2Zl/r0IPlO/MvvZx5QrBuHGaV6WgvhPbGTNzxFKiZ6rQOAwgJgZGWyDK0YqUTs4AVAMLX
BLEOJrfDdwbzc3+E0Fh8fWmTS4zLkhBVv/7bkXd5Hd2Jj15KvwG5O/KNh18t9GWmcJmdBJuTnAtf
/swxXWQ60ywCB9InQDr96AqXfOJIZLMDYBunZhmcwx5GWkWqtXo88//KkAqpd1XHDj8pCXEupUfg
T8HP7a7B8PfNXnQRUxYMU3ZX7myLPfpmPIMmkm1LzwuDRafc4n/RbLG5sKf2WBpytxWbfm306aNJ
8+vcRSZb7eZAa6uoqDZ1nqeKLrurqHODjkvMsK+TcPyXNDPgP9Scp8irEOcMKl7FkeHRC59eXfuY
bXKzjGoB6t44ezV0AOtGCcCox6BFw6bpSIMz2F456YA5HfghTCWm9QFmk8vMjW+h1mKVaRK9LZOd
8gVGTn8yXAUlxzxutYxF+MVRpy9JHAspZBrtSSgzYJ7Ogrd/S4v/M9Zm/rhN/JTG3m6JpM+dNYpk
r9dKT/4H/KcHuLHhPYQ9WONLb1lHf9L6l1HZTmRu60pZ5s+RsfHFtRst/tvdYGvDo74fIhCrzbJv
VeFwWlHcj+tSFlYj9T35NX6GGmJzPVLy4dHj8CWIEGJ9E27uTDYVfyvAt4ybQYoyKDAA4DHAiWOY
rNP16a/cl5k/sYq4R58d64V/Go6UJJh+b4iaQV6OFeAzTY4KhCkcCmER/TfABHDa6YnDE0aFNDye
qbAVM0TlqoevvcjS8CU8Csl8ALnQ7bQNWwIN3gpPJGdcTsNHnq2safQ+2zbtV0m73aYZWrCemjd5
Tft4WtltPC8XHIWZy/DiTraQ1EXl15naoMIE/XcvEjCwxt+wo9pakdZ+Jl6zjIniHZPCrqVA41Nn
MuvsCsff7GDYaidruJ4eDPBX1KPDApQFLrBiBr5u67mBemFtcJ+ZDBSr8PeeTqQQ1i/+eVUHSsUe
aAExXCsFKPuXOneHLZZmZRpAWDOBMiDu/XYBHYAR7kcjDNbY+E0flJA8r5I1cNppvr8f6nf7A0jP
nEWblNSb9fyAcS6WpEAcuY38rQUFRRBy1yX+u8nhfHHDUtmmi0F6EKBUmeOOZU1qWjNDV2G1/3oI
kiKSsfqFaB6RqpYk2Y34K854TcdLvX/Rug2lHMi3HeiUofjs4/GSRVc1KdNmxD3u6Sf+IIcem6nP
lJeclNo7duTo9nOU4eBH0LWAm22fB586VZPUy92J9eZI8OptNatbpM/WlIxUJVpV6Oot8DkDPud0
tFeD1yFxFq6xkASz5xD8kk7GG5PvsaA2aDLi4lf7I58ctFTrub1chZbQEqTosAsk067r+AwIbPKX
NYPPnjmSn7B0BVDgh3wJxH4BWBOBXeqWTzMheaGmOrTvBfiOXLwJumIBoMxljZPIplWaW4sDylMd
5Jd3kLA33jADAMWhKWvaw6Xi5eU0Q9LjD/s9GxRUUIPsPwUU61WMppQ2hJlD18v/dGtfOeXxJ+kW
4TK1tUfLnx/IBmQ0NssbeFtyww/ENm4UhpCywnCxh2Huci5kCg3iDIuepaU2WiE69OeZ3e19vsVY
fiKScU5p9hWDbfSFzidtFL/MMtGZPLj2o6V+TDXwadj7OSZUY38SINRbDj8Mri2gzSzwoAtoR62U
CRYyyA6slHE8+tSyv3K044CP3vMtp+gh6aVZpSWB3G7CvFb49lDnVF8Yc3Hvl+tDgLV39D9ee9pE
Zl+Fo7TwqAbvtWeMF9/rPdrJgFexbVVZk5EwX7Ofw76lUUKx92wJepRPgV715njTaqgisQNDYr38
yOiHNGDi4Xht3IcmdzLcMK41ppy/TEJ09IWq4tluTKnkR1tfWzOpAusDiKt46ymdbODWfVp3xxQT
wrsGVmJIXYS4HIao8hzEwPUSd6Gybc/T9/V8jBLYAqRULRwINSuo9/ZhcxPM6tNOWKcBmXjfDRnZ
Xopv8StcbutHxzLKe2UOUD7+sAkTUdYG8JWMNYI2ro4Wt725L49pISLzwbL5VCrFYnSUi/bDaBjM
s+kRbEY9IouzRXH7xVDk689ITjrtlJuCY+7NrzdTgRHUy8Y1OCaqN6ebF4kDBR/Ykz2Sh6eKeeZ2
2H3f94uAAtwwrtbDU1IHv04PBgxz1xgFoc3EDomgTHm9LVMo2d49CGizhMoZCiENmxD48O/cajND
oJNcq/7ng3Y+fcr/tAgstAo9Tl7p4diLBHIz7MjYA9ij/3Lv3P3AzRUAj+16Uo95747nyWkn1jVX
ZWOa1IF/0bRTTUPL8wVSwKpknenURQJAwZoeQmoUdAoWTMC8tBiPgFcvLLUvrZy1SZYy
`protect end_protected
