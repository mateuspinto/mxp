��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���S3�3��E7�LY�JC�ԌtMK�U�m$#�����ֹ�*�|��Q3Wb��4��t��%�r\��'��/a�pPX�B
����VUTzuD�
B�}��Ön��?�)w4��Yc
2F���9�8�Ф.zB/�j�4K�Ѝ�a�ME�Я$�T�_�Ră};�J��.�!W��Q�A�HA���M�6��W�%!���kZ�z�*��`�J�Ra(�7C;�d�O b��z$��%��PI�J��S��=�l�д,!yx_�(��a�[Gz�`_���hq�	��pg�#'�7ɉ±l���P �c�� (r}\�d�fa	I�e����(��,�^l��=ڵ]�3_؀]I�\��dt��ʚ��#��3t��H�3��2�{�6>�Px(���X^X�x��^2��o&4�`�:�g?t�DЧ9�(G�z%�*L�E�y���Y'��ȼ�����V �43�X�%J���'�:�i����a�ۏ�8:��r�����缾$�ozR�sn�7N�I-����.4y�R,��M'#pd3g�;��I��W�ꖑ>�G�N{y�w�S���h9C���Wx\.י}�>%�&����?��A�6��ž�ԠӞ��K�=9��p��r���i,�٪���6�]:w�k,IAa̓Y4Z��BnTX*�v��,*p�T�g@��p��2�A!/�rSg��C��`�	���=�Ԣ���7�,�%��|S�	A��~_�Uv?�X���-�^��6|,�\�N?��v�ߞ�(}j�3]�A����Ҍ�N�L�.~�v$�I���>�Y`ϧ�Ѯ�	a0�U>�6�m�"=�t��cEsu�ū�u,�a�[V6�����h��Jd�c�����L� �hί��X\�qk�K[&൐l��eK�~�D��ɯg�R�>��=�/9���[�{�����E��2=�R�4��KaV��ϝ�AzGc�@��%Gz��S��������ٸ�*S�$jxXr�w\�4��e]=��S5��>�n����V�P�Nr^�b���[Z��)r�����I����wV���TǬ�l�cj��1@��OM�V�f�E�`�n�'d�y�zc� �s��9^f!�i��91|7����dag��p���N�U��!�\��5�ȥ�g��	������~F�
�����*����rp�Q���5c�`�O{����m���:⺜X�I_u�U���Q ��}�D��ZM���Cp(���i7oZl�Q��;
�l_�Wr�i!0X�n<�_3ʲ�q�����F
���3l2[�kns
#�k�nb ���&�+�9��c����r-V�6�_���å9����;����LVQ��72� Թ{��^���[�G�L$	����-TA%_x����d��!��VtZI�V�o����/�^A�U_*�LOl<���|��=��_�n�ȿ�-׈���āfaɠ�%����1��_kp������o°���2v�>H�0J<�Ǩ_�zg~7�ͦ* .�B(DѬ�&��/�Fں����~Jn�^��lؠ���[��S���=E��&�����v�&�kD�A���Ρ��5(� r��	�4�J���+���EV������D>��Nw.R=k`���!E�>x�� =^��}�!g( �����;�5��P�����Ȁ`V?@]OeJ!.��q������K�ʵ4%6/f�c��D��9���;�B�� _ �S!���s�!���&n�,���~��I�dO%�K�5A/;#��V~Dv�Ѱb��]�q�fs�	��Z���o0�0sFC���&5�m��S����x�Ê�ǫ,(���vV�G��	��J67��Vde�Z^�=&�ȟ1�ݹ<�j['�i\���G�J�RM�T�����g�o��ߢhf�a��Xv���2d�ϧ�Ř��cR��>M�����zx�C�"3愕!Qz��n�L�q�e�"�R���f�۵۽u��M\�}Ձ��ݑ��X��o���E�&�P/�XT�������^]%xGU�����;�Q�͗��E�
�R�T�����ɐ�+rG�Q��0�Ʌ�~��*z�>��/�$��s����`?��!�%�?�f��W���N�%�(I�ӆ��B/���k=`6?h(�}!
�֖c��ʞٔ�/��������H�e����ӛS�/�-6 �L�!��v{J�aś�� ؍�li���e���x�AĄ]�5��JQѼ�L��6Gd�e��!�@��as�+e��̶	F�!i��>��J�<���C��gIE��tm�2��U���a�o��Y���hf|�=Q��Nq$�:�0f�Oxg��3��jp�4���2�h���gg4���)rv��.�J_��NI�vYT�x-@�>hK�b�5H>�M�,��w����%��#ju��p����+�b�O�Ƹ^���_�yj
��#X������=Dб5ad�['sG/�=L7�ſ�u�8�I�(�� 4,�p���?����hx�hPK����1��GϏ�%���Ǹ�ȱ��ͱAMX�Mev8Tg3�%gL/ۄ,��h~�H���A�$���Ն���a�
C��YQ����%/�a��+�D�E�90�����~~t�o���~�۬i�fF ���*�ii��6���˛{YM؄A}�^�{T1��`	]��v���~c&]�/эl?�Kf֘I�QC��O�[���?���1Wd?'�m�7��k�U���d����0���Ofjo�J��1�_�!�|�=�i���<nSU4�(�2��=k97by����)��"�<��䂱���CP���X���7���"}a��r��Z�d�k����I�nw%���	-av����rM�[mV�B6a�4��~<�"��J��xj�>.O�\�߈���r晙
Ow�#)O��{0�轏]#�иD��*L�����iI��6��.{+���C����
�2£�{���d@��@�ҪǓ���ח~�'�����5ْ��y��I��<[��T)�����m�:�����1:7���0L�"��Az��n���{Aw��!sx2܏-@�5N�{$�Bd��x�t Uk)̭�`�l��Η�W�%o���W�;,-�VKjt=��Z:�*PT�����w��vJW��Ӗ��Us\�s2w���ٷK�ct�b,�^Nu�`k�vT��
}f�/�dL��(��~�'���9Q͎6\�Z��RLr裆T��BM��|baVw%��3�A�qG�+��]��f�E��	��ǖ��ο#�β 1��u���#c��8
ᜂ�Z�XU�a����<ϑ�k+.��
R��<j���*<��F���4�tvQ�bz��f#7�^b@3���[^�.7�{�/���/	i�j��+5!,Zb�l��H�
N�3��{��Q������2�7p���������L2�E"Ԫ�م���j��p���fAˑ�����T�X_����x��x~J�8c�V��αC�ˮ���@R'P�W՛����<l7n(��1�LGCN �T��Z��8΃�1'nx�s��Ck��J��%�5�f*��1+E���;�ǯ��&���|�hB1-ZUH<��c�?+��`Pc��
Mb�$�:B��%Nj&����0�ԹQ�wW��"ӉLr�'*����}��e��q��{�K{Y���e���v#SM��t��e���-p��>&��D�����*$
*���Ol�s���Pǔe�7"8��:���^�{����IE���&�������_4���y��"�����?�ʏ+- u�	�82c��3Kg�蜠��ؐb%R3� [�0hɴ�"&��HO��N�ÿ�g�ݪ[���p�B��e�!-�����۶4G=j���$�N�C@��|���~��.P��ˠp�pr�#b��V�6����Ă��(�']pNL��0�r��><	֡P�����?�כ���O��(�U̏��-hu������hH�wD� >�J�wAPYb�q��D'I���#6^C�O����泅Օ���0!M��U��*�~J�E�<��8{�if�0�Q�![�jH�o�h�}����ݪLV�a�9��������a�"��`~�~b�w�!%̶��us�d��~��Vv���!X8�$w���nr�"J��oS?P��'��,TΨ(ߩ�LN�\�ūe�����m�1Y*�̰˹�G�����ӑ��>�Y����얟����X'�*#��i.ߵ�k�놅��@�A��R�� ��C6���f��3m�S�D5;��9C��>#1CҦZpg���ĔX[W��$ҋ��<�5'�^���gV��ַ�YQ{�37�Yc��h���l6����YL�Qŉ(�t������]� �c�xS,\�"y���C"y��۠R����L�=($�$@OwO��lz����;���L�d�J�m�)��v�w���QMdR�*&Q�����s����2#�3 �E�����id?��L��8���5a7ژ�� >�[��k�u(z�EV�>��$����"�励N��i�w ���rW<Λ����Z�4�̰��=�*N*���tL*+w����J%� � �G�\��q����v���|޵]+��iX"�q����w-M���ևA�{��`!�.�o��L�1ۙkL�s��|x&��my�N	y�,�i�����l��(�Q,	�3��B΋W�F1���_X�f6p���c���u�Sc	�2�1���w
����U>��6RG��a�"��"���Q��J(m�O0x>)�Ju&>��
a3��ѵ5� �%-0gOj�5oX"�f;��9�h$����΄������b��B[^��Y��n4�9�����,3�6[�������ot˂��J��a�X�����O,��B]5tB�i��(����e�}�� ��oTZ�7)�LIq�� 5n�)��UEŜ��N�O� /�o ]����K��J+{��^�a˓�-�H��w���ab ��^s�B��J�ش{��T��{ꄀu'}8bUѡ���K��&���M�K�N ֣ܟ����婨T�\ܲ�me�4L*�h�	x�)g�c�q-�]H)��$�����(x@)���f�f@{����"�-��}��� f��-N���r�>;U%!-�>������K�~�'���C"��{73Sxz��5���x�a���YF
���C�B%���_��q�^�=��<~���31�eZ��O�lE)_�ڳ-���v�����ټ'm�e{+�,w��籰�p� ���w&����ٻL��?��Ml�'Ǝ�3�8���d̬��� ��MC� ١2�O�?�wj�M93q�ƈ��S;#m�M��GЧq����[��7D��ekJ�5����Fa�n�c�½�&��d3�X�nP��qc�����J$0(Ɍ������E,�B3�*H���$Ks�d��]X�
g� }��Tm
I��l�ӗx������'ݷ���M��o���Y�F��R~�A�4��I�Q�����W̚ߤO�������ӻ<�w�j�������֝��_W�F({�!��l2��]xN�8S�,ઔS�VV
��G|4�3���XQ+�K]��E�W� (�����NJ����y�n2T3�jfE�'U�w3�m��`끛���E�<m妃�'sMR9��+�݃����	�{tjKI�I�()�\�2ku��8�?߆�x��$Dp�h����yn�4�<lx
3�Y�y-���G�ˉf�uwD�}$i���pٙn�f@�f�6�s�����P)Xw��g�
9�nYLf.�a��КX��v�m��MH)�����h�uap9^a����E߳,:�YԪ��&\����+�8rU�܊ҸW�o �M۟� `A��ʁ;-��� �P�_,���	�c��YW����AnH�5�T�ߪ�ɷ�cb#|Ȯ���#� !�>�!�ܮ���Nntؚ�px$N	K.?�c|�x�#f=�D]ll��g��)˪�tA܍ց�{�ӌBQJE�>��/k#P�K��M؉b���S; 2ɣe�f��n=���&�P��z�gZ$��(H͂ax/��]ߺfC��6_����ngC���P%ǒ����5�0�*Y]�S��*ǱQ�A�D�G��?��A�o��^`̒�b݆&.!yLFi�����/^��E�)Q(݋��eIX�h�����-�)!n�k��v�$t��4O���l��)�ZL(m��^��#Oi�Ҽ��L���k�������?/jC��;
�� @'�zCwp��(ʕOY��q:�g���r����O