XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\�椶Io=�������h���þ�d/���:�6�Q@�`z�O�8�����6��aֻK�w�B��\�"9f��ѫ�������4+*ƒ(al���)V�X]Z�%J�.Ðӻ��3ՅIKa\��<̔uټFc�\���	�zK�?�ԭ���:�VϘ�� b�;���xX�����}�夒���v��d���Qw�ēG?�1^���/�v.}�E;H,  ,���(����S�G�c�.z�jp��[.����l�ը�*�V�?4m�.:����=���J��+S�"Q�z;��(�]�2���Ը����l �Q>�?e���g;1�D�z����.�on�Ke��aX��ч� ��N��3�dkH�V��e]oо�yZ�e��t��V4����6X����kT���Ub@z�,L��A��B�P��2�f����|o�h�:�F�հ/��Ϋ�/���_A�>���֑����L�j��p��9�؈�j�tO�?� �ϸᖴ��<
�m�)��.��u���}����{/�:�T�Z��t�ky�� ̬Ǥ��A�;�N���)��R���!�KX�f�lgY̵Y/���HҜU�w������tuv����b�=�B�Qss�ϼ��o��o���\]}h�*gcgt���MĮۃ�b�GB�ꚾ���w�}��4yRg_����Od�=����~���Q�¼����z��:U��S���?�e�&2�X���%�g��f��x��+�uv!T����%��n*�XlxVHYEB     400     1a0�:�;{9�e%/z�Ċ�b�~������eS�����s��wB�*����\Z�a�[j���H]&!��v��fd�\��a݇��G?&փ���mB�P�GW�(��C���D-{*��ݥ`1���DP���6<�f	5�?������S����u��q*����\hgU-�s,�����Q��ob�&	V]p��}^LܛS�(0�˱�5��˩�$ˉ^�z���О�c�lL0nނk4��7)/�AuT�K-��}~8�g* &�0[j������}7]�2��z��}�v�󇠙�-#v�6�Hժ[Ϡ �|Ɇ�R��o���6�|e�DǠ��Ć��d+G�=<	Y��+�<,{\��@�߼Q��)�?w�)���q�;?	�� ��b�O��t㳐3Ҫ�XlxVHYEB     400      f0"��$E���+��{zR��S��ɩ��,���9�F�?(s�9BZv�\7B���`&	�����^+-��9ۼI3t ���3S��j�W�~��h��T��A�#�]�2~�{'��0���G�C�/�{8���Ĥ|(]@�_�0�����(�c�|}y�t~��2��mH�a���⁖�nϕ<*T��D�f���x_<���Q�t�e����o� 3��M�TH�	բa����kXlxVHYEB     400     180��n-p��N�%��H�S㛡ɭ�]d�*�՝�D�бdq�e����^�g��'�\M�u&�a��9��ĸf~�$Nw���J�D�ȩG�xV�T��B�?S~�����.��Wԁ	#��EQ����v�JtZ�F��Ek`
߸�h�sJH�
�|O�W��v�,��Lr��Z��\�������ug��N���B����OE:4�z�%�A�K�2M<��3��?��
�E������_ӟ�B��1Xn��k�l��xl)ᨿi@L�V(B�E�7��lpa"e*�����<%�5���H%���մ��`����ť۩\9){�h��~�YPC߾�TQ��:��/�N�(�X�ۘ0����yC孼юi5yJ�g+XlxVHYEB     400     230�Uw��ǳ��5��,�`7 �g>(,L@���;Ԅ�-D�� �AY0`D����_g->1�)�q�Q{Ǐ{�h�m�,p�����	U.���a�S��/���E�E}d�?��^�^V�[��?ѣQ%\ܨ���I��c����i,���79�l�����xmj@nH��C��*�X���e:i0+�*�S ;Jc��k����G��:�g���y�o�	�C�{��p���}Aj�k`7���1ʅ�un25t.2�[y�m���)h�%� �j��[0�����=�ꄥ����m�� s��»�����M��.�c�d(]/5��c!y��0a}�L�E����Y�ȉWu�^��-���3 x��lb��7[G\<��?�{TV5N�N����&乀h���m����xN��/�wjMpr������x�9��l�F�;���Z�$8�v�΄\�B���!�������q΅�\
��Φxv�M( a��Ϙ-y.�[����(+<"�
�x�c���d嚸5�OO�|��w
�m:���]�.�,u�0�Q"f��*�-����h�_4@�l�XlxVHYEB     400     1c0H��h�C,R�Q|9ż��a�p:yG&HEz#g���Yz�0���l]̂���g���$�_����J����;�̘��J��s=ٗ���,m8���	����Ԥ�?��kQ#�Q>MթU��0�Kk�C��<��t��g_RBⴉ�]����	Vq$����O]�?q�*�(sA�|��D�rWF�� 2�B<8ȶۙ���\liH�X��T�%��kS������M������t���&3L����ڮ�o͌z�G��PL�2V���P�v%��S� ���H�mM5�|͏O�Mk��)�*�O�{:�H�)Seƛ�8�?Z�2x���<\j��0|��4���F��O�>�dq�W[���'�:��9��5�ǂ�ڪ+$�v��uE{��-���#U�:E�����N���.� ��B�w��$/ ��
��u��ɳ �_�t��qXlxVHYEB     400     1a0��:N��8ѲH��K���)Za56�r+�}����pgi����@��
�dZ	�9CA�}nw������45 m�x��W�� l�M1��T5 H+Bh, pn׉��z�������_�ݞ�VZ����%C@��Eb�$��q���I�,ٽ���;�uD�3����Y��k'c@RK֌[L��̽`ـ�^���_�f�%���aR�(�4&&foe��M��Zn���-�#��'V�&� ���}o?�o��sRL�wl�����*�΃��<�/�&8{�NG��i���h�ė�?�Ք�ۮgĬa6�'��)�' �Y/0����q��AYB�F�?�@�o�B_����}���mI�ˣ�n�&��Y�/:�؈7�_��R�%@U>��WVS��{f6�B�D/���XlxVHYEB     400     1a0!��C>�`����"��B��=�J'U'���c4�Nt������X�+S��A���Y�F��n�����聙ں}j©� � T��0��q��¢�U+�!a�U��������k�"�l	?X���P!��_��m��%,ӛ��m�̦ѕ?7K@;�)�FK1��'m(�I�	�%�֊������6���u��� �A?;Qd�[:�p��B���߷�N�J���LPh�H|�ǮA�ĥ+���ձ�G8��o�'�i,�!������N_RpW~^p.d�e��m`l�m���ǻf�������,��7���i�GA�4+�����2V��[��[�����f�7��l�T��'(y]j����FYC�Z���mn���0#�y5�^��{��cW�?ϲfh�X�{(4`N�2�c�XlxVHYEB     400     1b0�*����tj��z��|=��+�TH*�.�d�� �s|42���e��9���cD���{��h9�4���jn�D�(أ���W�Q˺~��1"1O�G%hGIBH�B���W�h8����D@a��T�۰ľW�7v�V�<�!Zxۣ�U�����M\��	�I��lnrH�g�ﻔ���b�"�%�XB��1��:�0��mđa/��hW���r�:Ѭ5}������*��2��<�&W�Q��b��+b�wp\��x�}����i�?�8��w��$JC7mˤ1��xH�������|�9.LY�>4��>�-�u�nI���ѻ�u�8��_��1@���eQӂy���z)��5��tQDoش�ъ�1M��vY�mf�2a���2]8Y���p��(��lSM��3د��XlxVHYEB     400     1e0X�-K��x���%����s< E~y��n�M%�[�z]f�+V�Ղ5�)���J��>7F����/s	����6J��	�%	�W����9v1��o8si$����>)C��2�՟��O�'{�ǳ=J�Jm��^T����0�F<����!BLk��0�R�Fmb��xG���s3����PH��%�`<��Pʜ%z�w�0��N����Q�����]�H���bR�I6�DZ�K<qu�}�e۷��FJ�s�%�c��e�	��ihl�\HB��0�}��a�8>e
H=	��!�i��n��| ��{��,2����"����G��^�c��&D�>���({�Ú~��P!��f"і��I�^p�i��Ϥ=�_8C���Ԍ`�����L���j���&X<��͜"����G�o>*!���w�N ��|;���V���	�z��.���K�?�傢۝Џ��hFh�LpXlxVHYEB     400     170�o�?�F\J,�����E.ڟr���s���:������?�۠u���¼�\#ϟq.���!����� ��j��x=�o�;���s��sOuy�����F���2�L�r���TU�fr�^\%���:������4d�]e�V����.BV�t�,�*q���w҄7w�v��n�a}Q5��ѽ������9���6��:OcA|�����w�����y�۴n��89APyyw�7v����8l>���$_/:�~�i�U1�1y�\g�ծ��?�nl���]�z��F��� 2mc�ԁ¿���J㰎q9���>�&�l�U�	pua7C��
"�"�΍<j�|���jL�K�A*�N�~�a��(k[�XlxVHYEB     400     140��\��4a�j�����x**ұ7ʼ���9�o�Ǉ���@��4�*��KU��^0��CuAW����Vz
�,�!4 > 
ͪ�1�g����<d�)�f�(�7&���M�;��Kӆ_[��x�0�6�?-�#�ta9���f�;�Dd̹)�k'���L,�\�a�/�7G+�y]�����If�f�cm�Q=���-R��	�)�����S�����c�^0��-���?�:U��&��V���t0�G�_�¥�*�oQ��nA��涭f��~��@�r;���)sA^�v�&�w�!!&����?�xr��͵�`�1�͠�XlxVHYEB     400     1405���^b?14������Ɍ�3O��oj�\<��Ҵ��L{3��ˆ�,�hN �)Vg�PDU�1.��k3@��v\���i�`�QN�QN4)I��_��%�_��n&J��!{��@dt�<��� �(���-���޺Ԟ�אI�1���ȠM>D�ә��4ͳ�t8eHc�iq�1���S�h�e}���,g�f}�ʃ7=m{+;ɏa�<�r
����H�*�|���1�nu�t�C��D�:2_i���������'L.��{{���������H�eAGO�	I�~����\��T������XlxVHYEB     400     180��CA8�\8^�51U"%�C-�7t�'���noE��P��wj���>��X0ȳ^�M �~AF�#m�AcU{>���6+qK��ى����}��������~�	H��s�xRxJH��r0zE��<8p�g�J�3ܛ��}3�s�}-�z^C��z�o��Qa�F1g#+�9_�E�O~��6joߌi ���$��ee�:4� ��HY>���"�.ndB<�=�9�.��[Q���-��]�پ�ω`���Z�8l���:��sn,>?����_M5��AD��[��ZkP��ʁl�Ҩ@jR)�_������l=E�{����.D��ʐ)��Z�Q���U�%
���:q�em��À�Y.����l�u낱���;��
(�XlxVHYEB     400     180���P�*t�Bn��3���L�٢̥Bj%u>F�a$`��k��;I���=8�\�!�o֯y��C&q�	�-������.��.�IQ�ڼy%V�"a
������s���sd���+dv��Y�����<��J��QN�����죌�ޟA��<s���.�y�UZ$��D�W��)�}'�Q����c2C6�Ӈ�I~'���
��w��lJC���5�̌{�#X��F��5�������x2�,�W�1e�}ޘ@�~%�k�Jĺ h�i�l}ry��~�O��K���K��8�C,���W�[v}Ky4U�
|!�L�4�P,�|-�����!����Gb�Q8S���<ɼ;'d��+��;1�.5K<� ��[XlxVHYEB     400     180B���vx޶[�)� ���#���l�t�H���a�-KZK�ݝe�a��ah%�N������E�'�{�����Z �T6cל@L���)�������G����6�͏Ǯ37%�;h���v[��z"�Dc�}U��{0B.�A����o��X���y����(���w�(�Iz���![�
�/Q�z,��k$CL^�����r��I���'��>�$`�-}����S���l�1�����2O5I:*2�B���yj��(_��o�e��9�S*rJ��Y���`D��{e��yGZ��w�.��BYu��5����>�����2���M2s�㬈�*;AS#f����nSw��E�~7�`O��j�bЁ����XlxVHYEB     400     1a0���a$ �w����~r�Զ�B�h\p���h��0<��<.��6fy$���m�0�]ӧ\�����Y�sp���禴l{����IC%�����$�<�����	"3���/E��.���s���j�L$S�:r�t�	)���d=��7d�>�$����Ig����M&J/B5	:��ƠKr�Q��:��[T�hR����Z\@���3`���Cڵ�e�Q��tܺ�E�e���]�jI��:���h:6I�%���J�$转������l�@��TJ�VZx �O�$��g����/"��	5�~���,�rI�J�����9���!����H��Ghz�����M)ݹ.���2��r6¾�|��@��5�����w�>��e8Ll�9Ԋ� M��1�j���lk�yb���F�gXlxVHYEB     400     1a0���h:���ұ�]���WPe�]��Y��&��ff9�_al���~��N~i��h�®Y���S�5�'�|�,3���.4n�-�V&K�܃(�:>B�Z#�����<��Ck5a�/�0a���H��v�$3�S�>�B��)����U_� �3��EBd��2{�����u�}Ņ���T{Bi��]F�����1`ʈ���B)�t$��ϠQ���vٷ�#x��_*�e�0���g'�%	�&[G��τ[^C��¬dd�"���ZI[����ѐ���i�o��������`d�^��_뱶a�J3Z+ۜ8��R� Dˇ��4:��/�w�����t�
|�.,���d,��q��E,@�(��Zi���	Jj���:��ʵ������X^n���+Ξ��l�_n�XlxVHYEB     22d     110�F�VI���խ��8�%'RٻU�� ����%B�M�p�b`;UQ�\���w�9�^��Yp�4���ro�[���~RX��
 W�,��9�쎻��W7�d���KWϭ8��L��3A9:���u�@wل�ye�_~(�xGb��bf���A��Ē{�s>����Q3�j���1�Ɨ9�� ��r�p�9�����m�&AlҡQ�i�0ٌk���,���rb���"��{��kR�J;l�����@P�!�wfGh�g�Ց��