XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ue���~z�w:}�OH���p;������o(�o��tbH�(���掴Nퟝ��þq�ը�{j�~{#�����U����١%�ޥ!��mJ($=/�}91�2,kǙ��%:��*�=E��J��h�T<!����� �Jg�"W�[i�T"�-B*ΝFPK49~����i�yv~�0��k	�͒7��_��8�n&Uuw�
��x��0U]�ɓ�*� ���F4vy6��Q������}���r��?�l���5�ς=ό�c~jݼ� a7���6QMWAʍ��˕�PM�M�͝ �rU���u�Mlp���Qg�S.�i�*�|��ǯm �Β�	�'v��s��s��9������Y����Q����ʝ�FC��Ύ��B��n�?�]9�H�IZլ���#�M�JP�@�� Ca�?=������M;Á�\�NS���u����t�2{�~�Z��R3��RG���N3_͵�ȷ�QE���`Šy��{���	]{.f���21���3��U�PTlww��Y_;��$�@�+/���O�|��+Ve���mj~�y��B�-!�5���<m�W/����~��ޛ�lE�]@.gV3�:?~��Xcijy���OHߞW���Ă�N�1�WS>�^��%����?�x�ȏ��z���o�Y��"v�V7���0����%}�p/\�Cؗ2X-���sO�k����QT���j���y �W�{ь�d.N�԰��mm �k5��p����)ֻ B�XlxVHYEB     400     1b0	��ƶ`�9�_;k�n�9�����,��=����ņ8�IeWT��S�UѶ��6�z��[���Կ_ɜ��s����x:�c��#:#./GQQ*)+��ԅ���@�̾���O09'Z� b�����aC�2�B�_`9u� I�\�aW��f�}x�D=T���!��=+b�8��غ,�
�O���e(e{<��y�q�9?�8��?mim¡�yD�d���/������78�g��/Ǳ}TivXlNM�Am��9��������:�vr�_F^2��}��{����K�a	��^I��'�}��qC���W� �m���o�5��;P-8d�F�W�"t��XOZ���C�ʮ��.��
Ul�jfC���s�ˊmJ���Þ�����WT��z��Q���b�;����)���j�W�dn��'�+�16�2��<XlxVHYEB     400     160T��k���d�,X���ݶ��~1,Gl��<=�A�{;��L8n��e��:=�~hVP���H�n�B ������$fq»�����a�iY�_���x�4�{ѓU^Yu�zX��_�H�T� B+��Y��b1nO�P�雒-�L=����^5��K��!C\�`]8��{L{ e���p�����\N��w��
{���Ż�*�i5фt�W2qB�}�����e�&��S%���H;�1S3�m�HDE?H4 �b��JmQ�l�p�'z|}���T �[΀5�t�:���m��P¾�����Y\d�*���V�%��G�Ҧ��7a�L����*�Í���2���;��G�#k7l���XlxVHYEB     400     110�Ԩ?N�[�̓�zݩ�38oKp��c�E�?��.^�K���o���4v^Tu��0�����8;Ƭ����P��4t�Sni;`x�94Q_��>�X`�����I�AK|���fM3�g���w��<��f{�x�d���h7/�����	�eFTgC��ԫ�"�Ia���~o����q_�����U^�X�H��lg��ٺIi�U�Z�@5�B�-�{A�<A�WK�&���,˅6]VZM� `j~u�{�U�o\z�I�	����*�XlxVHYEB      42      50�m���J7������_\!r�ү�<�g�D�{�--�z*��3f1���V��wい%s�,��4a���5�,��