`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
s+Lcv4HmUN9xg/Gxdbrotdnozt7LdNeA6NQmqttLNE7YxRnlKRFzkO96xNRfWjH6zaMihU3KPvr0
qzOlCjkH2Rs3hPEs8xXfVcuGOuYtHh2w+RVWrLRbC4zi3PE7cfnHGRSN5k47Jf5tPSXrvIAuZDyg
v6iRxSTS0mXzFM9baDnF3/zolsuCTbwb/wDWSSGVV5jtiyV8yELx1tHUgT0SeEdNNP3ituxbcMYT
6J4wNCYoEzVLucJURZhfnsEl3TP8kY8h4KXrz2XIS+EfVYWHNXN0pGz5QFjL6TvTQp3+9+l2S8Xg
8kL/yR34uTso3gBTpFYmLT1wTYOmeST+ys+zplPSux5iqrmYuGNVHCYlmT0g2Ov1sJ/dmo4LVgf5
BPkKcuOjysrkucTIWrzLUPW2pFaedVP/UYk83Bo1cpCRDxMMSKmqHv+50scz5pK+ah0hZ4bp496l
iDeE4OJPelcpIVTSEHBMJKNUHThsVrsNMvxTCDms+YGZtjWFALZ8NV66rBNTNqoaOopBImKVo8uL
x6MCSce29c1FpLcOHIOUAQrnzRzv+ROHohrAq8tBtQusA8TX6TM6UmfYNi52acv5qt1mZd1xf7LO
SasOCiwpQVN0kSCLDyw1CVTKjVyZQeVUbtKl41Cl+4eCCzYh/RxoVlU4p7nHHLVnIX6ztk9dCNvI
dEtYJO2kDMOVldP80z97aS/4h/XliIxrb0WxQU/NBromEM+Twmt9cRnf4MxYK4qDeABhPJcwdTsO
p44yN1ZEVA6cOSM2p/ZRZR6EkYeUeicBQqhvHlGqhyg36MJbIDLi9YhOx2ShzSyTltGU2YK9vkEP
xV15OMvsZWikLVoXJjLPwm8LSOjM1j0s2CgT6o0JqhdaXAG/n/8cgLZEVIEfyDzBwgBlVSPhWdwM
o+wBzFaE9aAeaY0mH20rQj0AdJH8eJyfXNjE04iCG5yxxcc3btae8b0ne6+5cF/mXvNLkMdJbQDr
hOz+7dKJGTRYAoAkblF6LXlhWcZJfio+7n/30sXUfTBwwfrRImaCOkSEh6KWHPl4bnwxi64PkWzj
BAupaOdtiitXvgR3mlgKMDqyMqmuc1tAiwex5Hd+lR81LxnLKtW1RK82PG/W6CnwHtRrXKtdxG3S
t6p3M8Hc+rX+gToGKmMXKA4d4wexmAQQ0TC6lm4OL+m/CZ6w2U0dCFwhtUeLdNOKO0X9l+CRVT+5
oSIYYfZx8v0qzYfyOPVlxpQS+EFLocP0BsGfEWV2YgiYKcSK7FUcJUt31kzdjoRb8HP3yBk2bZxN
EpnCCc2qF3AY+23+Guv0yWQgQtDTyTFpGgpx7NUBzSVSc1/XOFCGTLkdnuuNSOkIYV4uomgcdeHb
GM8b7IVliI1/vhBz4zFy1fOJIjUcF1BuHHX83hvmUjMbvf4WPMYNdqu3IVAkciaL6LlJGqddGLXd
DvKNFazCnhLfvvsl3jagj0vq2w3IOACxsqf4GpZGyiwserBIzu8s4wqnvll8P78hUb7hgXOQlNEU
JS970ZkyaLxLmWdF4BrrwQJnR9gqub1dTRhAR++hgSWUx0d36aOjBFK/LgaJUnm+5hshJ2GvPWU/
n+fyQTxjDl4+p5xF2DtvNOe43dVDlxzC2SZKzAaD+Uf+iqPOZrE1x3PzZm38CQzEgIs5QkzvX9Kh
8KoeXzMJTT//XmFVGxRbXAsR4HpY4QKPkdnJwZv9U12AqVuzRH1whpDz+E1kViR2QO9oC1nHDTqP
YDDcQr16f8V/KNYMwaNs5r/NUsOObX4G7G4VbfQz3iR0YNY7qxE2rJiTI7UlwgQZFspsGR4Hw+GO
nLG+dWS37YdTc/Aq+xneQd2skEzav5pWx+QTDk0bUpAXLy6YirXbMplInpncCeZ41VJr73sMPw9Q
vTm93GvhFYaqw2RhEgpCm51lOiuyg4MEpCzpAHR5yF9AwlUySGd+Q9dtx/fs9TaX6idTGgY+K7g2
uloH04i9fby3lfDJ1ZGI6+CRzkJGVCBTzTR4ludWzy2pRBOSHXCdTx3w5JhUG25zgzD1fy/te+An
1uCQbLqavu2CX44fmWQhcVac1qqA4J9loBntcmhX3QfFt+6m0yshULMlUN67s0/8kwJY2Jrkpmvh
T68wPaAyjmtI8pOexKG2RFOMklK+Iky5s9EJxVBCwlOfwejUTQgL3nplMPIjfHYGO4WI4Idi8zVZ
wQUeOYM1yK2+n95kG72Rz7osAK+UjppN2GHrrn687P4m095J8e/Adge+0vie4je+Uens8ABotykV
pq4+oAo7XCr1TtBVjjtfnf17ZlHBrzXkF4OIhD8LI/HxHl9FtiRMWV9xohakGYCQwUvIdrwakmdy
2pHOvvLR3Q+VrqiMFstAkw42mvm0zdQ2VLlb6NhFsc+yHcvwjLVe7jk3qJJ6arKk544Jfs9MObMb
rDwJa6DpsiwclmE26jY8/UGdzz7hX0Y0IJtl/u6QscxwW4BQXp5cQHJ047dMfG7pGCNIKyVb6xCS
sWrSQOrT74DMi24IMycSZx/r1RbILduwcvKEHZj0DAPsNyvd8AGJDEN34Dfay3XJVR04GUrkeGth
VCwio1ukxICsW6R/ywFFbnEh2o+R6cCQkYVKfpaTVCCzjAFLwXyQfUOAI3uL4HaMQfIt+UWkUZZc
BQKeijuJI6I3gq3TcP+WXnWDdpFMXjfjnwEat2UVwrm45PGa3tdolLQWe0xpB+NL43b9X8rzchrP
CVCUBEz6PakCv7QTKe/8x4iPEt/sAw6bylreetWBESQiv4+v/jIRkj+WKTXQr2PXzCwcgdldPPxt
TXTlcHC5MdmvkTEGsn0PAwz7bRq1gErg9UNiQnxd+Xre1uF4rn697pXehjKGYm6pZ80trLboZVA3
I6raa6HNO9F3aHDUPMiiCp5Cp77Ch4LzC2fnQ+4Tk06x55zOxbPiGk11j1AeFzw5Ikg+Hg0PEyGP
mCW/PVYgd02N0XPUrdyX/fgTdGuXaGn1SmjqfZTTQa0JNIXt3VDtz+nPgqcT1MzeNWeRQUA9eJA5
kMMztG76Ti8s3oMxfyvpYgeW+UPXPXWEp+Egk77asOUXy0QS3rC5ywLf0seqoTVpf0w1oNcwA67X
1RUMIeSpUDPi+PT+VX/d8FmLow/Y0TwrTAkRZUo/1tp5Yymk9z/SlNwZZ9H/fQnWhmwvsQeM693M
GtFMTJ3WVM98JbV55BM+7AYIXwJOG6+fLEK9X1gZueT6kp5eynAnfXtkEPUzq51ajpQnQzVDBapJ
Zi356UGqj0Voo3SKKakipvAN5n2Y+FZXgjTAFRRAaoPIex3rX7pCgLoBnBtWCfVxSI6fGXXxSq/Q
FskxOUHEfsWVX+Hgxv1VIJAN9wUar8g0L8R/rsnlAPNAWNDE2wpE9QHBs7sl+djcFiZVtyl6o1Ay
Nkx2V88lzjPcxNlk8HReodcSeIfD+xD2ALSFkZoIUPStix2UjdM4JaM2tiCJB3Dy9l0k+x0guHD6
1lvS2dDK+vZn6HEQPYcnzIom3zTTT/ekyCn8yw+GN2F4bLcN3kCy3xUXyTJmajdL0xlgQMPEsIaJ
0NBJ1zFiQnlSqp5oazdt0pyhLdL3/VCHjbcmc5mrTYoDXI2bqlrdz7apuiDx8b+lNsnK5AIakxbw
NMkhOAAuDKe1GvrnBbnz835EiAhwvcR8hA6JHuluMDi+BrOkyUx0Y716dyWTbcon1bDsKTYOIUw+
/r3xoMlU/7t94h2+NgSCQlsGIBidRciDJmYl1x2CvOCh/vO+zq5GinETA8xxMYO+vt4o/AG3CXNh
lNSPrOIskPJM11nnaRML7NapB9UIcJvlpYP3oM4ZO2qJdwbfAiuIyR9Pn5yffWFCMIexFplbV0gJ
x3TCx8das7YfhI730yaPlAmff1VGk+p7qM4reXe927HOS0wh8zsMe4r1usY1fpD1fkVez8+C/zmW
iM/nomPH7pFnq7jtnPTlUMBu3uPRRiiklyHvGM7TET8wI7viHvA+GUL/Bz6F++sZJDiJRthymDf6
TWYRZHGIUe+XAhB5ZnrE5VPcXk/RCn5H1Iq17Pk27YlSDiRuUuUUSEIlLUI+d5wUQYOUkYdBmcBJ
8v1/EKF6BOQLK5xOhQ8E3hFMXUDHue2Xmrnyx4Xl29j9MWCgv5Oa6HyaHlEdLELa8nY6euksW1h/
WsZVN8Q3UKAbc0bvSe+SxCnn35wCkduWaCkotpcGoKLPAhv1WqrZXpsbaU786wKXxFYp+3TgpH98
qK1I6SzVPjqQF+HpsNTMucl2ewhdnAO6jt01JhXT8fQVeDZJ98EoyFtNMfbkKuzNtwF9QU5RIeVs
da6RZqRwRP0LiBX2OR0RgqVzpJ+CccWFypJH4T3PSAZNlOxkeK8dqNGAy1sKu7qt6SVV5AnI7HfK
UB2c2L/RxICIhrpKOzVinvcrTLBNe2gk8z2y1I1UHvaE16gPWQHlTLWW4h+RzeAi9QODvlK0nc/F
SNDXt8bc5a96VCnTn04QjjZA808bOonD2N4ZwFezIWPq1rCSPWU+cNBQqGQoSezdMYoINAnW6kPj
YaxeLr28wfAB7J6XzLLiArOOCvhNVr0946VurheKtiVFvmj09RzU0ngj1ktz3BHaVIampVyj1dT8
gxCwLjbSzx20RfAUWHlH746kzrEaXgz1p9MMrqbylr0EeyEWW59SYpmG/hr6RuRfoAhsSDOzUf+n
TRXCYOPVsqgKGRAexlsd8LwmDrBdgFH1sMPEONH4R3ItrqBVFk12B+PyHIu8MOe+eu/1WO55EUG1
BQSWtA9Nj0W7Fl8gc893Jb8dqwlkQsQqnmh5VsQ9XrPfwAOpKyV1A2nQZeJww6gIaTfFjGDS/fiK
g1eaUuyP1km0eclNqYjs+g7vAr5vPFKvfkDKnQzOqcr51/cqYGnKmK2qviZ0ayVTJndxJz2egEtE
VPWPf2FEaskCEEpCFLjxPINocTtwXr3v5zpACmYcopHEtwfCltM84T0MuIJ3NYNNgpQdGX2waJaO
SZkwyprbR1X9AVkcCNjkUvxZJHI+4cZnRG99ZG2RF5VdoL22+aOPgVL0ffQgFTwMrmUCiEzKQHei
OjDIqOpexTmW70gyD6U5zlllIUEjqf4HB95cLCsWN75FBTAHAgTevcztNwda75C5AJJP6Pt7yPSJ
WhE7RFLR74wfPl9T1MmZW2xb/NbCJ6SYQ/xCMcE9ODO4z/EP9vB4tX31mtNXXPmqXV/SUNxoTwuY
cOi6+lQS4eT8BKqlquYKVr/dr3E596qnAB4NkACkbmW9NUgsFodxjDaeS2FWTaN8th45mi2mQL8A
pPEM0hufFAMD4BAWhLYgjr8Ebp5qRMmNLk/jiVHiNjC5mK8yGz5oe7z8Eo5NF7WWd+foQGJOoWr8
ATzH275wnBLzEtLEGzpMXQYs774tHxT0IcU+t7UHSs8jnLOG9qauWzs/sOdTXy/ug1c0nxFDu9Kz
EUZcbvb61G+TaXeDtHaClYvi+P5auJuIcd4m/TjEvjBjFJhYAvI0mwj52Ze4DHmbxZ8w879orrsH
Ldl5tkyQlZ8jh3Ft8of3tnVHjd/VU/9SHcuKLH7GLg/HXUflW51JPB6uiURR6tirF0VXw/zvDGgy
n51SI9xYa7k/EBtKZfHVJfPwZO9ZyTGBBNksOxCgPJBb2rvWm9vd71XU1Xq90O80APh094jcp6ZK
bQLln19EsHVhcs/xMLSypyCwz5zsaZ6RVOmX5mP/3OcikZyCgo65mjgz2nvbRBs0k0ehdXHZZiHX
P3cAbHVAxo6ED1nnvF07tBUA7ztrCA8MIb9yFNra9GlK7TYHuOIhW2BKL8mH7Dw0EKYQhBXAOPxl
Z8QtByuunRZeMHD/jbOaBkjPrZdiixnPdBl+XexR778mBWRGDt/paEoxNuW8VWgqDz11FrILhT0c
57z3lqImwvn6x7dI5iKcmoI9DyDNVFPY581G0x1I/YHliHpQI0A6ohy/G/uKVlX3StL0Uem33uVK
1gvEwBqSFw1u/V8B7FyINmpDbi8GGYuU0dZBvgRiUEc/a75M4Ec5Q/2+pvdzC4W4MZwBJT0eQ48f
sJBOzrQEmo/WmlK5PVC6jGQGx0NujkvtFAPNRR7FzZ+84AvTkNtYPVOJ0MTGx1DkdQHx2WV+QEP9
ew543LSuHJz3VnOA7JS/hiPJnYfyaMb0BhLVG+B04EH11rI+39eNfSdCynoyLTcVyHg1uxBXlqev
lca+fCI7SLyjd/vd1kgI/PXTQ8gkX1ntfVSe/DJE2wIjGBlEmRn31Vf2bM4xWTILsIHi/m9zQ/1G
hJi7Cb946W+cOGpIKlsRP6dNRBbGke/zrsL9uUyPplTXMhqzbbnjfPpxO7I5XqCGEcOyCQVl7iBn
iPU7c83sQLMNlEVlhj7V2koVuX2Ea8p2uQAriz1u2kUCbzo80Sr0stUG4Flr7Gno5j+NazyJd4vl
9Hfd0td4oq7FYCcN0KRHiMnHqFMHJX3Qk3MFxPY9kPVFsLX4udvpbg8OyQxfgIAdaBTURm6Xkh6S
15PLGb14vWxNckX5sZVrUR0m53jI1Rlsacw/Vlfj/2w3jXSoVP8h8kvnudxY48a6UWhucIK/p77h
VflFvb/c2xHdfU09x0xu+7QnnAwcg7MXyr2iLgTlQi/E9Fk90PV4M2uNSllIOgj9e+HJatOzn4qL
NjrvYeb3pTi23GMK8BYYobp+EAzh8aw/c7cFycqdsk3qUWiKK57a1f4n8CaHIGy4PdjPEVg5PeRG
QeIt0ZeaaiT2rBUN2VeOYDa3XhBBvAxtfm5Q/qs1FpNvHiwOGEsWPMhUdu/j08JsSKsvvNWeScaX
WMXVVn4YWBAp1EHQ9D3EDG8zzNVejCLxKMVcUTe7hd53jI6Csahksdg9Wb5GJYj23aS1CktTcS/E
xynVxbDHuPQKOPTud/bFqRihYg+Xl9P8+SluXkyYjfqr6IQQDlRtqetUE1W7x5SCWVqzm7fnxciZ
BCcnv4P+Lqy5NuE7sOSfAyKvV044IqcJVG2ALdo/vc+1H1Ku41DMlmGSyV45ACFuCCQRvD+1VlKN
WZltuqd9opHDm8z/emd889YwGDMulJl1ynXlqcHTwPEnf9W3v0FadsgKLcaka5O9ulOJ7KeWB0bZ
1uxRaJLKNC8OVih0pqMzzsemtghuo4JvUkgcTQxZgp3bOkxYR8gX7V9ft6RYDlrulfdmYoc/IwdC
XhElQbW0RJZNjAK/FRiKaobWA8beWwrJ5jHNrlX9DuREt6fOTnFi0h6bp2PPi9VHuciO4Ng6RkaL
J7bKn7PLfjeK7GWCjOYLP0ydMxdOasKZbNAk0cJ/eW25PnhX+HpN+S20SzoM9ogFVNABQN6mHaiy
tCsQDpU2rMoQL169erczJ3OzrEB5zWKdL1K4MbfnPtsaTsgBr0x/NB9vGQG1UXEgNNs4pTq2vElg
TFMT6ypIx1rX2rN1VSfTdKHxSutraZ41XOBi2QBi6aWk5elaMWh4UgI2JiAwbex7Bj7EyCTSGU7T
/Sb0dyb7uw8D5FbEUXhmv/MEIRntbzGfd0HHQRDL/G6I3+lUoUc1NJ3e1qZTof6goTJaLxJQ+7o6
yQNeIXWGzz3IfLpC+A5GIR6SzZeksOPmu4smscKqXlFKuqV9eKBDnpq1tRGhkW00eeU0f+3ogS+e
TyKGkG+bpaufjZb3rd8kpeKWL4z806fona6mfcdwrjkFj7ktkD5QzHF134bQFMpQVJWvopLvjwMk
F7cvq0dnsklIWSuZid1SoqW7OW6m36cP4u8CgqdYtXpw7MI2/Ojpugf6hvra8fACc4N/L9Z+O5M3
AMPFtZP3CYC5P7xk7Gxm4wm+KN0Za1ksd/0LWtDX/+OTC/96/+MgqBXzLaaJT4G2hGM+B9WnZ87N
SVJ8fmbprInrT/CCxkVML6Yh/Ty17fWguYncZUPESP/bptRo4RyOz8EypvEcD7hsVdrU5naGq1kN
/cO3OrYmYSjDTrKYDZ0paTLeQ+xEjoIPKRQ8F1+DsJ318V6aGqS4WrBcMCrDVn8leCS7bnPhDIqT
A4BNEgM3ysXgM28dG+mS9nP3vCwxHmSay0LvTBp4GInrYkxp2TuECeIci2gt/O1c0SjWq4PYInSo
oFatUSlrCmr9TnEJS7ckIF8HFy8RriTOciKzIml2PNzKXeQuCGdtkpLys7gKoZpqsiRWl2lz8bsM
0CJAwqVVYtw+pt14mMRnjUDmH6nIfuKJh2wDWi0mRYaLaw01xRFYxlmiu9bEl39U+Cj51xJGmESd
IBtC1F32h5y/F9TaxOIxnSunGu/gdz8q1wi3/tIzVle0sjjmABS+XCtj/f4yipy5fnl8tqjnrA/W
1vi7gPhagGKSJVyCJmfj3qx0joQWlEWc20u6oyL0euNiSNxoieX4ni3rL2PGPJGXCYm17ssGxIIE
N7jBDf8DH7x2ID8EpCDpJ9V9vBQvbdlo0NhheUX/mlFsgL6KiCPcrzWMpRB6bRpHg5s6lckAntQp
IN5y/qpP5s/dj70XXeArvVXMETq15veqvU8yi3/UIqWxwjRlFBAfuMYcpjRgCr7uYMQjBZMVeTJb
hfKN8BABhCCaSZlA54OOHNnnH/H/VLsrwTYbsJVXziCxA2qXrDZxpZ/8CQTYNVeKu0W1Wo2Ggnbb
7V4Lc0qeBgtsm9rsmXZx2iCe8zlTss0a2x8RQ4YYP9IjvBVdwTB7fFrYsO2CWFgrsK1TdBhbyuGE
OxxsnXF2VQyxYwjQx0YIVENRvCed9ovOkoPX9WH+KJs8WgQf8lvKcH6HvLpnJjfU6oZ70I7HTUIq
itKPTznPZKn4rmJWBmIdjTvfTt+5vDsvaFr2Mfk8oTAX8OBrAbWozbRKqoDo7anJPbpFXXyOtLtC
r4jdzLQbHF0mAgbf4aT9GkS0Fkt23UCMzsJobCfdqQt3fGpD4eqOiYuXeu0S5cjwqviFMBvFXgMg
DwlbKrZaumtD7lmJWooOnbER4Dz6D8jhbiYDTDs79/mgbc8i6XTac0k9J2M6b6+Soo8zMvWGyudY
F2iag9QwEKCJ5QjPuRa12y0+9Z8QqgAK6pO6MgsHvddLmDf88FU7eMOAnBGTY6Otf8kG8YMTb7zb
QjGgtYNGV0S0rPBTDUI1U9X9f3+E919FjKebmHSgbOQTk7VMzqINnzczwYDjXyKtuNal4v1bwqnc
Gv0T1NNvkJoJIQJFVNidbYFXAJT+BDFvXP43WN+tN8h4lZKMzpuJF1CuCh/y1Bk893jkMsmxmWGH
fhbzX59egBQTuxh2fwFby0P17+CNmM0D2rFZ6L0zNvRBNVaVHqF6+Eq6K7btdHIrIaqu+8d+I7Dj
fJC+iixl/Daw/YRCrwB5AFF+5QfIUUJONQBH2Pxbj7OSq3k9mykIxhaUnjX6kYVHbigf5g0rPMBZ
aMlvBKxBVrq58wdxr1hdVRtiuR6kctNzwl2mAB81XDrWqwzNcUgFfBbqx67ZTSowoBZJKGkBU5+B
rONGUYqlAkYqQ82Ry3Uw173MGIhPKdIJNen12xnZEPE4JTgtWUzsGZvJwjxDs0y9yZCfoRLDIiH8
SdbWRiyyFdUo8n/kuEugNSG4xUXVbWwEZUU/KDLepaww2t8UkXFRAjS9TX79YjIkqCiCop2MmJrk
IUUXLHueKO5MBG4kp2gubgacJX3dewrnc+FvIIKrF2EXWCi6Iyt2j6FQrl9dKpGLL6OT9X3fryo9
6XE/Rf2fOOClr1s8SFhPobak9h1LAFrDZZpTvbZExEDr2vqxDCeJQV3nc++gE4XcUQS0AEXKyZsh
SOSQ0sAXiMV37qlZX+4c6qA+C6IEENy918hg2hVL6oGI9dHVeL+3BXzbdBtLVxEhpD0JQORSfL1I
bu9gt6b8RF65XHFDlD/a/UAIxyANUcS9OaJI7+Jb2LJwDO5HleJPcQQBM15ydQ0vM2z3zCbq8MeS
lie4rQe3EwP8iIBSCaRBphjw+5jOJWYT59f/Mnk0QGGYcBB9C0cbA/ld8T2HYi3v/WvdJRDIVGvj
eYc8nsGVlMzCoJ6TY9WHPwCNK3KyrMA1SipRkCyw7edQeDNWIPcB0wieigbwMCdbHyiHNbo1fbnP
5aXyGKKgm+fw8J8mRNCpe1vtRAUECB/hIAHxTWmZnPVGy2xfehFasIAaSd5Acy3W3r4oxeL3WwQF
mqr0Q8yb94q+GDCPIDtXfI7H55fRIJ7wBuQJYAwxxFNuURiLs5ZKCHFCoUqLtHg2mUqUo1SeITon
+SJXsPC/uRu+K/Iud4a/xKpp6yv7kyTKhVbON0Glk8tbAlYeUy0cZp0K8vayfRMOY3jXKtUIKkOG
h/fG+Mxh2uy13ok2nzD6UMLXv59phGl16lSDNf1cvK3MaicLRLPKi8jHEwDFWM/buMegc9F9K6eG
0dHDI/5DLSsS0H650Mb2xgZP0RwHVf5vd3FegPgIUbHfD8n9RzdBovP8jNQWYvf1Hg4k/ffU9BAz
2/2bRY8dfKsq+6dbadUwVnyAiCLlVIxc+jpQVYUUALu+3LkWIb/SyY4K2YUlS1giYkPTaBN1dzh/
KnAAZcMY4wqNsXEIy3WRhcNZgL8P6ANs9K3UDHjyTCpJb5CqmUeuUaUXHViq0jWipeGuLDrGCRdQ
FDmqL8bibNOJBwjdXQkMhaZAzw8tQ1lhlu1+4yD5buTmqNy7sEW2wTus8c+skUx/ivRp3FZQsY5t
FRHYrAWRHMuiE4tr9ZOxejcH/DyAsvsI2Nps4YDzK1oqcTX+u03J326KlSmhaUZbjSrm5d7BW81w
BOJpQgkxY8Y9cCbPxQuHIljedrGnGL2aaO38/HyjvGQF09YSZqs0XBrXMtXmwCd1OY10bnEyTtSE
ugn8B7bbAqW/j1vLGhPKx5dv1Fai6706buo1f+skrl1CnsTeln/3gjuGufiMKjhgzh6Hg4mnLGmG
Q8PkzWXpt7+HIFIIedd+maJl4S4Bo6d+eCUksvZ6YA7RQA0ZliFOELIhETR6w+cVBp3bllG5THK7
fuaj9jXkq+6k1wcAGznQKm+Nuo0FmrN+v9po2TXDMC1Q7H7n/RWrAAdB8TW1g8mZVwo8CAw0SE6x
3pnqXKGJ1iL/hAIXi+kst64AjGPuqu4Hkwip4r9Z4ZUp72/bCODpNa1J3Ybrq6Xr1xre23tYSwd+
UFMcxvq5NdXP3s1MNLdP7iOTQTTfn4kUEc6SE9o29QxwUG3m9cE3G18uTUKe7tl2IJGvbam9uuge
7p5FJL1FQlSMW29c/2EGoli71FAyMSr1I5Y1cjJ6zfgev+zOGVMV+nfwGTTo/bBfxMsofPMM4HMV
2gCzoxRUydoVYqyLhCmA4C8DGsN3sz9PdglMXMqk9Bn9y3RVCBXlaXS1BTeoAJo6J7pajeXjil6D
hQaxQ/DxVTw9DsY9zXfhc6pC4U6nCLjNU9wEPhCbLkajiK/yuy04g2bsuD3JtG7Lj5iF/UWk3jTG
1zfAI08rGxMLI8rdIVu4f9V6LM8SRrFUO/fzE0kdMx1omW/ficHx6FuACGfXrnQ0i8tYt/ZyV1fk
XssEfeELgdSS+bTV/gzpDtdz/37Dn/66mQyxRueRSAPYg+rXPTdZRrwpiM6d+gqCEbPVypdnOOZt
xo74py6629TpA6gHnCtz8SodQlZv6wo15OTRfSm8nzkxi3YQvTl2+lATtXUr6WkwKqw6/EDaBanW
s7bd7iXUMgtUhrSEiKqMmN9ttjE5BPerrbEJlVrMhS5OjtmSEQTmuAKd4zmEkwScCKOyFgzaEFZ3
Aeh+cZwmS4iD6onzAlSERmDW/Jv9/b77YbcJ829CUGC1IT7bNb221QWvdmBwtUrh9mClNPrZyGuj
2GSo045/Q0ZUjNnowJbaOMOwG3YM7Hh3SIt7YlUECV51GVKZsT3eQA4XR0y+07Kq0p14ephImcYo
rQHkYT5bRk1irxovvk1zD8ekZ27NhWhEzPkBVilCnf+hPjKs3oaHYuUqZ1hMpr5nOzkUr0Ipqk7K
01/9IyBRLN9EQGgCJWlZVuFkENQkTcQwN33rNxivxhBmaKW95t6ytXjOJVWu44AyUwB9gV5pmqoA
6zU4jxboigojmUdORtgOshQBbQOa9N7+QGuwLwJkjBFyde4zSs8szFxQDoWuuCyQpx/cPf/fuz/0
yxz48WayaoWn7vPD1a3X38NKG6RxviAJ2gdbr+IpOTE=
`protect end_protected
