��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���_$L�s���u��e������7MR
����w��6����T�w�X��sbI%$O$h�s�P$%�bh��g�"�w.�/�xZ��̛��=e�bJ/.ۤV}6R#���0�9m�$F���§�}<�Ԡ^.�!�����a2ٞ�j]�8u����`�M�C��J�����[��>�^��R~Q��4�t���D�=���V�
')���N�:P�ԓ4��L��,۔�U~����מ6]�mPjRL�⦢!����˼k�R�H�`��+l�3 {��΋1�H�g���T�W&��RZ���Q�]٦!�rē_�!��]uJ>�P����	�J��`_�h���c���H��<��@�i�'�P��2�\�h �����R�k���c�/G�N�
K� ��-M,N���ySn��W���<�[t�����R����_k��S�jH���~��������r��2�y���ި�8��h�-@B�� �&�~�[��ժD��L���D
~h��K�cy��-��q��؊~/}��E ?M�ߌ�0�&����+��+c����43���"�\�~��//�'�#[sH:�@��_��u�~%��^����O���=�����u���8����h�00�[���?f���:�5�ޅ\0�ք���ɹ�?��kÝd�L�E�*�P���x�Yu��v��G��Qh�L����QB�|���u���W�c���~��
�>}����}��9�%��4@=F�^oJV	J�a7Ծ��y�	Zc}�K/C��tp��)à?�"���J� �uh��=r+#Ƨ|��-P����q�X�:�P�G�#w-��7�E��O�(��ußE�Q������zk�+��Z1nc�1^M��WG�����b��a�B��^�	B�[
K�6�>}�� �#�L}�;����"���r�SW�;���&��P��sl���DXD�=����\�f}���`�(>��gU�q��gx=�����,��Yy;��MH��&��<�1[dG*`?�JBq��eE�K�#��V8��Ǚ����W{kx����j�����Q�U:��J�Nˡ��kmDR��k&c�V��������bM���"��YԠjC�KH�/0"֓��ٴ�z0S��4�A*�>G��}���Cku��V��yDmA�$�Db-u%%9�\ފ��]�K��hE��6z`��<�Ub�DP�*��N�Z� !���G�,�5�Z�EL!����_ܙlI��*
"�;�.��RW��HV� �22%8S"1hso�d��:O��H�AQ xS�����*@Ag	���>�.���g�J����}�GHL����m�D~G(L4 g|��#˞�Dk�W����\�E���·�p.		Av��^�	W��ցf�VV��y�f��i1����؎g�hb�z�or�[���n�.����z�c�`ANG��
J���M���+��҃�2 �l�#�ט��OP���ɱv%�R�KuA�;M�1W?�i&5E�Q��U�Z��L�[Y��1H�}�=~g�FI��ƙzAS�*��#~hG�&��=���ܖeY�����:�@5s%i�I �����%�I��򷯳>k�T��5��z�/�PtZꇏ�N.� K�ܼB�1$;ش�U�E[XefJ��o�y@^�i��
������ EC.�L�+�!f��ojV�-ǒ�(�����Z�}-���6�Ѹ��f#E6kB�\6 g?��'~�SHɅqG�޲ޝ��������;�ӈ��͙�>(���Z�.�����2]���%R���VЪ0,��U��Ժ4sG�Td��8��b��{�SC�N��kN�N(Yrѝ�}d����q�9���q4��>	�]�<�Y��	�'i� ��J���t���_�VŃ�{9y�'A�җ�kg�r��8��m- B�_?��ʕx=8*�_�xo��6�_����y�5T�,b�xi.��^�tм���f��u�� �c�������,�~w�d������e�֨��rw��T���Kl��N���p0a|(|��+�|�u�̠�VV0v�Q���}�"�yR&0����q�f5��<#�r*S��Q�Y���v�}�eX5�x�j�zv�)�(8���FIG����pBZ�2�ѿD�7p'?xM�h�������\��Ҕ:׵8x�J�� ���[h��fC���?����.L��_�l'��8%�Nċ_��c��\�L=_"B����/\Y��2j�ӰB�"[�"�YH�g��v�A}D�Rƺ��q�j�,�ZVF��c�W�����M��*�+�o�0���ZA����rq�W%������x��o�rN�6$���T��K��y�`O�e[�:G&O&v�v�h����r��]�����W�V�˘��-w�l3U՜��;�Kah����mz�7sC�?�=�����-�G��d�Fi7ۄƸ�]����H7[���j��
޻g�G܄�(z��oF��=�(�>�|'[�B��y Ε��A౯��>�T�aK��bB��
���J��6#�F�N@4)&y�Փ�x*�E��r���� ݜ5�ۀ8��f���	�GG?z����E�Su�v0�\�G�(X�akRQ��4�Z���\��A�Q����_䛀��K��!�`A	��+����WJ�t&�����A�<����9��
r��:AniA��7�����Xv�d`���v��tD=Ao�s2����(Z�'�}��q��9�m!�6����҈��ܑ��YW8��M�SS	���l�`ۮ"�r��o�#r��\��JK_�f5/��v� �ض�M�5�@	?	��8,Ȑ�������E����c�,W
���!�S�F�#g����p�N,���g���'�D��tM�D���_���>mY'jl ��lMR�b�����{�4F�N43vnO-�=�����l?�>��?�0�݁���(
&������@/0���`�\*y��S��k$����)��0�A�c�k�a��vt��^�K�����#��o���C���]�50ٱɖ'��E����"�3�'��Y#��j�}�Û����ؠ{!k5�^�4�����EmSS�j�!Y���}{�C�o�7�s�}��&PJ4^$ Y�
X7�OX��7/�}�t������!��PH;�#z%�N�!��5���~,+k[@�LKrs�(/v_������b���e�\��S�/^Fp{�g��[*���p#?cg�]�,ۃ�#�
��ѕ�|&z�Gu
�`��Y����f~���;��R	�D!mIR~�Z����ˇ6����~MTF\q��Do8<��|��C�e5�pɋ�`�+W|��a����Ȅ�.;d�z�|�L���wH.ȷ�"�Bŭ*B�2$� ˻�*wc#+�.o���������zw��C��±�E?��L���F;���- Xz����l�l��]��c[ � <]N�II���)J��P][ۧ�M�7�V�5�T2>mt��B��xּ9ܭ#~Z���t2ZL[z�00A��4r��ɮ֐0�,�`��̈́���N�ƌ��N�=�7.B��Y�i���>%��\l�{ʺ�jN��H!���n�ݽO��f��7b�=�L��a�c�:����%ŏ�Xo�I���
�"̲a(��/����1~/��t� ,��7���`�`:�U*��Р��!�A[W��iG���h@��Fu=A��Ҷ�\�Y;��8����lZ�y�cP�Ѧz%y�V)�u���2}AM�j<����䀴��%`�W��\48"�#�G{� ̑T@�^�)�9r��j�D�%M���Hb��-��A�C��{ޯ�ۿ�P�d��G�"��OH��8��<���xӮ��ߑ�}�u2��%��}bq'����>��a)tq��A�{[&S�l��O��r2Y��X_8q$��=�&� ��������TI,��YqW���0���r�&�Zkei�J���4WEHF��a(#q���V�����*5\�H�P��E�%�9�v�k|ȧqJ�,��	>�ri�B�Âo���z�{���y&હ����R5��P�=:�-��POD9��x�pX����9@Z[ ���`hy՞�&����[��l�"#Z%r�R��*�I��o$z�n~;z\��y�G�<��Uqj��#���3,�Vumq�E��Si���0v�Nc���������[]�cWE@^��Ki��ب��{��8��h�<̆���<����(�(��ɠ� ���t�h����5,X۴X�?�s�cP�#�Nl"�F M�[����mqs$�s|������ˋ��F��=\C��,	���ਧ�,�Q,�^c�}�w[?D�G�	�i��͆�&~�ڭ.�dM'*�����b2�!������ʱ}�E��1VV`/ɬ�],p�A�Ë��h�_�9U"��mK=������K�Ԋ1��A:�K��*��g&U)d�[{C�10�St�hi���e��@�7���{ ��5��]�X��v��?��$�	,���AP�����I�"h�$Ѽ���q'4�(�����l���߹v6�	�XW���&V�́�o?pB��B���S?�M}(���SZ/(牚s�G�uh�n+�gf�t�ߺ��]�|9���"�1k��q�F���+�5��3��{��N���Ub��ji�M+Cx��B�/�[ƴ���?�9��<�b�qUAO^	A��I�(AQ@}�L(�i����GEt �tZ t}��1d4�=��@����)F:����W�k4����8jz�E�O��53Rz����EAh��<H���R��cJ^�{n4i�A"�^����%����N�=�m�a����s/��7���B��aj�����s_����!F�M�Q���g��2:*���k��C��{��GL?WS�_à^�Q����\�K�1ߒ�U�4�xU��q��W�b+[&n~�����j�l]"�1���ڍ��̪��;)��� ߢ�I�B�Ӂ�)�s#���
=W�բ&=���'/������(a����}�Zt4�M���8ce�+/eA5�4�5z��>:1��q�����	$O܇�$�����P|u{��/i\v$�V��swoaf2�Ŵ}����1U�\k�R�Y�y���q�F�)D�C�k�i[���e��H�*IA�oY��ְ5ߜ����p<'��c�%Q@NQ6˳+��R��X�V�$��05�,@᳢K"+���"�ۍ�eGם�����z�bwwb�V�Jf�>� ��+W;�;�2�q�Mό���T�a���K`�YGU��a�ը�cn�l��ο��O`�(�G��B������ чDo�I�W�����	��ޕ�0����@�#��D�H�'xZ��z�gT�I�����K_Z��z�),�O���:�"C�)]@&��l",�A�ۧ�(5b����Yq`�7%C�`Tr$F�5��o=y�*�v��(�|�#��p咑���!���[���wB����Sf3A>�ZL��С�%42X�������.E�j�C��P�Gb&�����'�DR����ĭ2�U4z�re�*��ܛ�ܜ��!h0/|�M�=k��O)�Ī�C��ϛqbN!=�i���M���}�e��iI1r���zӴhU�����D�*�ԯ���c��wqy���9�uA#��B�`gncd��2��N���2�(�5�#����֎�������J�LJe������
��=Z�oN�ڳ,����9�;�sn�����:��y��y!��O�.�.�����h�2I�8��]T2t2E��6�_��jH�N����XL6ǖ{1E�|R� 1��F�䰨n���%_O����'do3�Y��~�I���y���)�o�%�^�+]{a"M����TPb�[c�Å��]���*�O���h̿O(����y�h��~Wh�̊{A����,\�]��^'����1Û�&ض)�TN������pZ?1pS�C�a�粈�UMkN����>��`�q�Ɂ�?�W�iaOj��*7�6G6�]��:��VU��L�F�um'%�ʽ1��}�K�k���2:�
2r��S=[��}Y�s��q�`����k�&�o �4��.��2���h*����T���"��x�.�i���˿6l���(:��W�S��AY`�&�Оn��;�bi<�W���
��9<��d�>���I�\cG�PQk���j��FQ����K�i&Z����xXH�Ou%�r_)<O����b���C����-���9Y׻�H <���Î�zU��􁕸�"d��ֈQCdL��-�[+:�p�0Z6����*����d���Y�#�y���ц���+~�|q6�D���E~����S7�:�7��D�n���;� ^�'�I��z�D6f��*�&beo=(�uG�gc{Hj�ڷtKDUj[�^I�mkq�q�Zv��}3�XLZ�\�b �X��t�{�"��e����y*�Xl~��ĝM�aO2'(�s~O��t��V����Zz@]�!n��=[���e����S��L����H�y�ｷ$l4<���@D,��#K7��M�Ϳ�!����-鏻$�8���@ω�����k/�,�a��S��f�%�:�����v�����+{�m�Ok�qH��l�����ңm��ꛝ��Q2���q�$m�T�w��5�/��Y�P� i��(ٟ�+T������L�<��3������������9쁂�ʞ�����>�.��ʠ���ҙ���{mY*K�rL�oqc3�U�_;
�������1!�Q�w��ؽz������r
�~'Q̻΍3�����-�f��Fg��G��ٞ��m���}$��z�+j~��{i�΋#��aC��me3�4�4�>��N-�ӥ�P��o�����Ռ&>i��p���3������w��v�<�-�C��e��	��a
1J"�$͛Y6.���_�㟶r=��q�+�{CPO�~��1�#��v�:�:��~�'��`� �o+m�6n��c�|Ժ�Go�	�	�B�xd�)|�/�G2��L@)�S�Ќ�p�ܞz����{ms��[�5��2��vz���Ce�}�	��Ea^����h��hF�ɜ]��8��"ӆz��S����hc�����|W%�2640��
k�J� ��vՈ�vc��mDOU�4���7E��/�T��(�p��/����+T~�� �E��6�,�/: �D��j~+<�HT�;���鎗��ì��O���6�5�[B�,BO�ѓ �-�q���'_�>�5�lh�KJ.�z=;F�.�X1.�]����R��L���Z꣰}Ґ�`	��������@�	�Ff�0����aWX�b1�^.�F�Zٝn���C3��kT��!o�j�
������2x��bE�g (w�*[�4��~�M��� �z�)q��1�D��|W��T=����f%��b��Z��
v4�LVS���`GP3,��Q0�vkV��-G�P�3+�ey���\E�����M�z���Ȇ@U�+�n��jPH��M;ҁ��v��lP��q�R��:W��c�ޗ����;��v�7���פ��1H3qԬj�X�ά��P��"��)yyމ�\��ڋ	�j�Fg�Z�1G�]��`&,jol���o�Ad��<�O��w0#LNh���\���M
Ŗ�ma0�����BL������d�V�Cq�=�j5�y@��6R����.}�QE�^�	;R>3�H��cw�;��S�������7o<�<�6a�{*"vH�����Nh'�1Fz݁ƅI�\��C�<����WmP���VI�y��@ͤY7��z;ԗ�
6���!�40.=N4����!������)X|&m��2�~�JF���H�	?��K6��X�(_;}qP�5;��\��M.�!��a�;��G��EB*@}�Q�c�|�峲]��Y�����1�Y���������Ң^:P�4��鹚1I�5�$e��V���&����8Τ��@��?.X�z�ϐ�nH�>"�U�VqG�BWT8ب}c
W�����te�|�Ҳ1�Q<��r{ÃWx���d}�L$p��F�
�a�)��g%�(w�b��@Mʩ���kQ\��uLj��!+\y/�8��&�	�MtF�Qy|Aq����3�K�@G�0��z�~�eD/׬M(�Ն�O�?e�?���?0�m�� �?��?�_�k'�Q$���\Gˆ��C��+\|�0��oB��}�D��hv�}�)�� V�]:���ZE	J�	�'T���i�&}�"!*�(U2˪����Gș�s��.�oS�|�/�n���zya&�yq���$�|Hn$�OɁ}��)!V�>g�Z��/����\��������Hq��_gp����g4�|��/y��y���C·����( ]�pv�/%g�kwT�B<��M��A��6�&��ƩD�JY;P ѭ�Q?�����5��7�	��O`���6.)i�k���Rw�����Z���GPc�y�.���ᑌ�#C��֬w����m��	�gWs��-Q�謨�&�t��*^�	��p��8@Lf�7J�QS�A�h��_��;Fy>k}���-7�� x��ǅd4q
fՀ}-��z��5�{�u��cy�Ȯ�Z%�yu��,��\� UU�l�z�'�K�����S����(K���ٸ��a�3�����k�ᱫH�S�^����_���~�r�X�h�4�:�![۾�g�P�;6FE�P�Wu�d����3�`�b?@<ե>)òa�
�p�3P�Q2���/.�9x������\@I��o��>̟��"��࿸�"n��G�,�c1cT�0z��[�y�-��4��{	?��?��C 4�DV4\&�p��r;2���r��Y�U3n�F�0�~�� yU�H�2�8!_�F&]�X�
�$���8��:$�4c�)��hs��ڐC�]Re�9.��7�&QY0�PL|t+�Z��L٭�L�/�����$�y+��K}򻄱m�h���!6m�?R[��Gۨ����,�/Fբ�)S��"䘃6̗}�QV�a񽱛D���
�rh���fz��}��GZ���YìL�L.u%��ڵ|\����`ӑA@r�z����qͫ�޻�=�y����`L�:v�v��wi�b��g-5m{/�����G|i���ʐ��t��AןѸP'z�}R�E�0g��TK�I��5��m+tZu ��Fx����#>כ''�ܴwy�9v�(<yy����N�pj�g���tvO�J\ϔ�l�QahPĔ������)����kx��%/0�H���rW�
 B�������;�IFa�/�x���g��>�x%ٸ��m@��|�7����@":��MF�i	�ފ�q�����x���1��lWL�O��-�>�w\��]`��4�ywx�|�eտ�/sw;�D���mE(�����j�k�.��g}"Y���$� j3Q7{ʕ _��
��O�ط���>(J��b/_:dj4(8U����u�Ѐ��ܒ�.o�e��(90����*aE�����3�bz�(�r�TS�o��N>�P�dƭ��u�zP���{+õ2+�]�p�������d]��*	-ҍ�ļg�?�i�X����1�fGj{_!3e�fq�V����3�_��-S��\�'�M5��7�|�"�(�Ou��z)�����e��T$O�C����^R9�.e�ؐ�|�������a~ ����Q�D��D��������
�HX�N=d��nҫ�3�����0E�H��
po��=?��+��%\"��y�cE�����Lsۻ�l��3eZ�#
���9
�Y��閳�쏃�	��R�E�x1�7OL7ۭ��x>�m�_?��!l����xA��m�3�%.n�
�Q��!��7��?�$Nn��1�ܰmFC�x�x\)l��)���j-6���@~jL(k��s4O͌X��*!f�$ة�
*f=��b��xo��;U����Q�
�qS�Ȁ�l��&e�N��q��1"!���tܑ��.0����ie��־�_ rZj#U�I�TN_��_�7�_��Ev�"v�<�6<������*u�ڔ�ב�N$l�H��ܨ]ʖ�X6���u!�}�Ɵ ��Av*�6phѷ��{#�����F���ECi9�m��E��(ŕc����)+K����#��2Cy��RQ/��yşv66�g�؈�]S}xw��`�h��vl4��ց��ݬG�;�t��< )>��ۋ����:>����>;��v�>I]IȡG'�c�.m��h����0�䷐U���{��W	v�Y&*��[��6Bʂh�m4sRIB��G�6Kn?^���������1R�&>~NS���
�����6�[�j?t|�i�1����QRtn~��fz�<I1���͇ix��b�m�ĸӓ�)�F�ʜ�%&d�}C�V������	e�ߔ��0��W�c�ɑ9���>��f	cC�kDzb��F=
@D��)ֆ�L=�'����|	B�s�5Aۦsŷe�a�g~%�FAyk�_~�FvgXI&><�W�S��a~����Q���ςN�{
T�H^_-�N�ص%�,�8�2�Us��9�]�`�N{���r��m"���P��B2�,���=s���!o[�u�F|�|���*ָ�@����淲I�\��Blm��WP��N�������6��F�9r������2o��.��"5���J�J֛��� ï����[�*�W]VJ�B(���5w�޽JC�1��?r�����^�Q(6��:"BQ���:����4�_1�OڴYt��������&��u<C9�D��)v��i�7�S��z*))y�0߰40#������vE�2��W��wF�6��'L!C0N�5v�M�s��y�w*���y@N��a��;;�.�ˢy��^x�MN��ec�2��*�����W!��n�v�` �vOa�r���v1Ŵ.Hl̙�֍����!��P<J�����3/	������(��	��\�=�|��jC̓�"�d���2|�_z%M�܏p��!�C���<yk��p��Π��Nt�A¤�h�Ⱦx1�l.o�B�F/P�/�l,��*�-�k~� �Az��t�I�5+���� N&J��H���c\�0��^�/��?l�-=��|�
ŏ����I�m���sE+@>e�(d^>��V���_�+T���y�w�[F�m��(���[7;�����Kn���N�a��'�F�晵�:�W���6w�-T��9=����dv��#2�mR�����S+��BW���ё�
�u?��ɡ�U�1�PO��&]�]���QQ���6Q'G����v:��G�3���<��=�K��w61Y�+�WVL՞�ۢ����tg�2{�j�#Pi��{�T�0)X�̑(�@b���ɋB��Gs�����������\��Q �C�{ah_ڜ����[ ��(~���PL��t���'��XB�e��"�l�'�h)�e�5�'-���φ�j���fs�; ���Ї1�2T��]�iK�#�N*�����H��dx��ݭpĄ��X��1U�oT��O��;�+L/w����RvF�]�h�Ym�h�?�κ���1l��0LZǅ�4��\�z�,���[�t�$h�ќe�W�?(W��b��ns=8ϒ��Ӏ�{�[a�W~��R$��	(�AӉ����@�xzt�	W��`Dq���H7իʋ��_���a־B7��ldy%7K��kD�-e)�l2hI&�N՗u7��ơٚ1�t�s�C�Un2V�9fgH�D7H���Q�G\Zw��`�� q�%����G�!qo�^tD���ڢ�w^��,Y��y����vj�$:-�9�4���(W���ɱEz�E	������%v�I���l�|�\ɀ���h#�N=g�����zPv�Y���z��\����2��>�|@GД��<��Gzq D;f����(��rq�_���,�_��Ġ�\Î~�:0��E�)8�i�C�������A�}�)�6.v�
~���t���\F�l��@��|(E�`�C}�&J�qw"�@vݷ��j�*��\�2����
�ʖ2a�����,<�Cق%..��JW�2�w�ܬ�A�-\�R�
5:Θ����#�Ԁ��uw-@�Tm�q��|C�/6�׶õW/��[rQ��;ˮѤ�G��w��L�'q�����D)��b(��44�߭n�|�[tn��w�r�@XWr1M�>�z��xr8o�.Gc��3S������b?��!�[���9X�A��?
���_W����hłe5ѐ�@oY�<��׹k	��_�B���i�Y_�ђT���.��K�6�6p�X*��T�Skͱ�wZ�jy��l����)��a=��`�>g��8AE}�`<�[T��&!璗ֹa�\Tܴ���sHG�[�$"M�zk��B�6ȧ�ֺ��h�A��7��/�MES8��sXKf��(4�w�Jb�"D�v�M�؎I�O7Z�3r�3m���5A0��Ʒ����"�7ޝz�IP-�qH�X�m��fz�QQ0G���ۏ�,ص��-av����]�ڶ�:02#�[;(«��$�ۑ&���u��<q��W#JPP�TjT�.3���}j �M`�P.lcT�2��9��`�z���WE�O$�ܭ�d�6Pc�6 ���{T��4�	��
�+2�l%,iB��(k��;(� ��SX�_.a����	�D/ ��O�����K������`H��#�/���~��K
�pHC�塷C{E/�b�&�Z1<E����G�L^2���a��/As ����+vWI��%� f��H��Kz�L�I���M�q��[�|�T��^�RS��(��Ӊ.M�b=�CV��࢘��L�~,���<�֚ �~��
b(���e9����^ά=�G[�B3myr&ͧ���V����+� ��4kpG&�Lx��Ǐ�.9��'�5������(��b	�4����m�#�V���|�PN���k l���S�=<���ךy��Sѡ��^0��l���Qx��C�Ҵ#�sO�	_23n���d����)��MW�.��$�2 �?�U7ɒD�[p�_L�3��~D;�ly�	���r�6�awǓ˼�H.�p\C�fh>���q�
�7p�q�ڍ�|"��*r��F��BV��f�d�G0�u�{j{\Zw�]�oM�v>��}#0Sh���N���Vt'�P��>em��H	��-$W���򦱓���*%�O�`�o?k��0�B�Ҡ��AI�ޡ7wLh�|�\�6�6P	14T@����D��FX�p5��P�Խ4}[^��i�n&~�d{]��j��F0Q�~H�o�~�6�{���8}�)����K������¿@9�\Y���N��?ٴԤñ���������=�YlȘS^|�ȹ:W{*IO��8��W�!Ǩ'N'Eb��o���]� �*��R����;�9�W��Z�~u�NT�ʔʤJM(����-"������B�Ŕ����PX�U�O��kR�bN�e��w_�7�s2|QT�Pǖ�F�������|��5]=�qjBf�<�;^y�D�e1ll�v6zS�{�//v�[W_���ZF=#jq@=����}�3'؉ӠE����&k���8�?]����=�~�[�iX��h��
�,���h_�Z�\{�ށ��P�?��8��h�z9�)�����Z�@ ;㓹���Q[��l����t92	S�@y��W�%��eH�c7E�uo�CU�A��{����_������(I����SO�-�|�R��̸�|k�<��'4�5�Ф�GlC ����oz��'+yH,�o�Ba�QSڮ蒸5I�(�~(L��	!���{��.je^aR�|y&�F��>I���C�����'�9�m$;4z��Ǟ��h�G��n� ��=$�3cF�N׾8j���I�q��(��.�-�gS�=�c盦Y��_�]84�"�j7�D�tܨr��\�݉F�ƿ���L������W���eI����]`�ҙn�)t�~����m8ޑq~䳡hܵR55cD�!���*Y���G'ߣ�Ʉ��c�d��!'��<�T5�+#KK�&\.m��)a1��v=[͕��M�:h�F��7�'���u�B36=�d�v���WN�佟�S�H���Ai�i��κm�����R!�qP����M�� F��e��}Ģ-����4ή-<L��B�i$��}�'������Lޟ,�$-"@H�r��;n'��f�z������8s���u��,�yO7����:b�U��NXalF�~Ƞpd�{�u5�~��Ȑ��f�ʋ,�3LL�W��7��-���p�v�N��5MȰ]^2*O�ke�eA�;��12i8O />�n(g�u�`)��zE�^�.�;sUlWРQ���HG!f�<�-��&I��`]�d��	�}���⺤^���*co��a��G��=!�<:q$�l}�7|m Q���
E_1��'Q:&�Gx�(b�������Y3G��.P`Z`[��b�}3���)���;�)�����Zh�:k��Oqe\��v���=~p}=m,n��Kh�=ɟ��y4ˁU���
W��;`LM3cXN��a����d����O�26L ��Ѯ�b%�YTb�/��O�Mg�<����`!y�%�kx$���k� �ze�?49���=t�t�o�i��/���M�|a��h@���3Nw�5a���Q���jw�k�o�� �򏚤�xP�mkm@'�P-����S5h>!�E3j胢�z�#�1l�Z�f-f�]�>\�
�T뇫�nc�1(P�\�&���
x|<gtqb����HVƶ�^�ok�P�!�Z�h	�d�k�CGx+^�E��)��W�9L6lJ�h#4{5vv'7�4�6(��*�>��1�����h9�����Y���'�����K>{<ڴ�Uu\�y�!&ϵ��S��h�+=l)�*F.]ǆ��l@U+s\%���$�cX��9p��0��,��O��΋�D?�?E�&��*XYɹ�h�M�(��=Ƥ��Q|!U�ѰP9�A_l�x�q�E'�z��|���:���$8��tiɴ₩d����K��)���5�w�k=��z�'�I
dl�� %x� �Q^����^�de�����Խ�s�-���L���;��+���w.B�3Wv�M�m�lС1���Y�/rr�m�G2��ս�&lL���i�r�Wx�s��:/�a��tF�ŧ_������!�6TW�/��%�K�b�I$�`D��ߒڈ����J�}�bP��'X�f�W_�y��q�V) �\��MغƣҴc���M��Cq�w��B�zE�ZW��teH_�	�E�xS��	��.%&?M�[ƈ��2���R�B�J�S�v���>��v?�O|�i��	��N��:�No��ɯ�1�|<:vQW�c�#E}ݩ�ʲ�������X�%v������C�nEvb~$�;׆ē�K��89̲A�N��O���Ħ�b]}��<3F�l����v��U<񞿓�(2�^bl�A�������'U9 �?j10�9A��Bw�F62xU�LN�I�_�J*��VSA@������/,�(_��Ao[2�b�Es�՜�D\V5� ��Gزz��;�|sl���,�*����*@א^�QB��f�sf,!�S�*"�[DW�{����nT�Whk���:���Q`�drg�aᲇPH��
;�Ap��ʛ	���#��ˌgl�Lu��V�3V ��F}���Q�ϲ��D As�L�Ӳ�n�Qk�8�ኄ��{��Y��L�S'ov�0qb8�G ���L�>�V[���3̹w[2���VR��8�T�2�7�O�i�^�Ii 4�Lh��'6��`��>`�0$�񣓪���_[g�T}:�;�1k�����Z��,��ۄ�#�Ƞ� N��@b=&�r�U�Q�ni'����2�� �m�*:�-~Xd���k|a'��^ۗ�,�'d��|�hb�#�x����5�?h�W�*�)
��d*�a�f�5�`�I�h�FϏ��k�B�!2\X������J���5o��hм�����j8xI{b*U���6��c�l(����Ȑ�\&�^�ƜFô'�@�#xKS"��0����a�_���}	��"Κ`:lsc�VݓG��nk/�NM�p�e؛t\+�Yb����b���z�<���|{�%7@mE�i�9���!x�וi��Q �~A¨����@^�_����ϲc�ʯ��a,O��kIՖ�?Z
���.��!���ċڧF{)��%��M�|!�ߺ}��=c��[4�l�Vh8, =��[�������U���n(��x�0 [
��:���vE
1�L�&d���䓥F��~\�&$��*m�&�,e�<L�H2
f4RUv�ZSd?*��q'Ԥg���%}(�"��{	H�ȭ����?}k6��,���g�����m~�r��ෛ�QU!�.׍ᨏ����+�t8�}�g1{��
^=�T~�6N�`����F�!F�O�B�eZ��^��l�F��A���א�a��Q������	-�0C�	�������>�Yt�w[���dr�K���֣��kI�?�i�R��?`�%w���cq
��vb�_�w�����uF'�Q��.���͖M&�O2asp# p� 2s�U�u�����E���yg�0-(~�A|$K�q�����.՚ �C�-����5�u#:$��)j�qk�"�WuY�%������rM�Qx-�[չ�~��?c�OtI���P%]����Zi��П��E�Œ��k�w�sA�m�n�W�f�e�m�%3��r�,���ɔ��<"&�Bk
��.@3�b2BԢ�D�u���A�H��	huT-�AeI�X6َ��/mf����	"��/Ⱥ��{
-�'��1Poi�c|�l&���)�����IKǇ{��[:Lu�s��K1�I���ɤtb���� ��P$�Sa+B��R�GB��`P�xC����ǤȌ��?�g��G7e���h�}-JV[����4T@�Qٷ�1��^��!k#!��2�uOH���d|g��;�T�X`#)����L4��[�E���%p�5�:��I�aR���bg|���$�,\c��q7�<�7�i5H��UwKq�~Nx��үm�^�Ӛ2[vC�tE����%H���w��/ ��"Gk���s�ݲh��<���9յ�	���p��L���"(�ɬ�;.VK��HЅ�y,��1�|�sm�ع�׿��4wчc��l�2�13 �t� g��g�MW�{<m�^�kR����|�-+����nZ�&�<^��=z�<�J��)��@�] ���ɟR2���a�	�4�}��{�k�总wD�{ĩ�M3I�L?�m`^q��&414{T�Xr�c�⑊������gq�_7�0���L��Q�wjʞ�Y$�U8M����l#4O��X���u��բ�� aJ�	ҧ}�qZ4$j31{/i�'F���-�T�����Bmy`"���%I��Y��I�2�'o��6{�K����#纩d� ��?�ƣ�SB4�����v g8ʅ���?�����d��8�6�b��H���[r�D#h�,����85����k �HF��U);+YCy���*6���O�1��	��2�L������AH<; i�8�e�������o�F/��Å�&8�O���P=I���{$�4Y�:��y�����{�'�e�	%���P(����{;���YQ���"�z��Ib�E��� O���1}�T�+U�IQ/����On�����@����אqr`�.�h��s}��N��7�� ����Vg��.���Z�V���4[\��\
,���!hܨ�N�R�|��V���`n)L��"�3��~%!�%3�`���|����z���H�����)'��	����C������w �=��<��	��yb��ǒ	�"e�����	Ԗ����F�Vdm�7��	�_��J���(�b=�q����Qy{:E�p�_?�����q
�!�&��G����r~���/|e\'�6��6(�{��7D�@1	3�<慻F;�3D��4w����gm�Ri�l��s+�(:�y���/%�V��O�-���"�[�t�� %77���h��Y�o4������m�>����M�VGh)��Pȣ��L5nHSh `^+�rֻ��&|
P�j���d�->x��p��NU*��[N�
�͕�<���ͪQ�gEź�����-?�&�h���ئ2]�0��� �m���{V
Kc���;w=S�D ��go��g���d���*�F��p��r��;��V�p԰E&�e��*P�ޯmk�?H�8M�tmd ��]��1"G�����T����!�a�C���^�+V%M�/���Z[��B�h)v~75,O��l([�?�;ٿ4FɁ���A�9�B�[:���e+t�ݴr�LZ���iK�榺�X�A	7R&�Fo��N F����{��|�J�)��o��8$IC!y吺��'��|1;�����?�9��&�[T��{�5�؎�?R�m�N QZ�:B�Irs�X��a}ob��|�(�?��M�P�	
����1ֳw����d��E@돍�O!�_��Bg��=�i�+�E��$�?-�-O�ވщ�\ees���"�N�/V�|'� ��+�Eԑ�i�F�{�J�GY;���3���~}qK� ��}Yw#�����B�� 3�� ����.���W
�!�GlaI��M���̷$	��P-nos�b'�%�;m��5$[�,���N�!$��)ƭ/�1�~��V�=	�Ll=�ΠiԇS6��'�� Q�erVG�����΋�aB���8�d��B�rYj�	☰��&Wo>q�wn����(��1�2틲�(@���	z��lc'�-Q�|���7l�@�rl/z��b�.��a�Z<��ܧ�2u<&�1\�
Hs�k�`�g�9��Π�������?�����*N�Y�(RW��l��u������@����n�+�&7א���N|8�Z+\Luo�f~-�H@��[aj�X�"�4��5��R蜶��6���ʈ	�瞵Ąq��
�TM�d^�ϟ	�>^��q��4��n1X���!����iI�#��H,�F�[�9i*,jV\a�K��A5O��+Gm�F6�w�%GԕB�\sʹ�k��%j�0-��A��A�D���v����#<~=n�	�6p��rZ��������O�.�Ҫq� ���f�pٴj��1���U6�010�{w��?�1BB�X<n֊���@/&�j2E-F��(|�J�A囟�@�~�3����g,��4�7Z�uKhoyη�H?��4�"2�3\��)��zP��C �dJU���z�s���Ԕ��Pl�X�lӔ�||���*�2���Ŋ񠏮�B�L�T	s0������x^����J�u���y��:����>Q�s�p�2�{�|��L�(sl�&,��W��,������[�x��L8��w��r�+{=�i�6J)g���#[�c-m�^�G��;�*����ka�Z ���qq�� ��Q�U�.M�Ot�`�l��Jle�������#h��9y�oj���ߩ6���QF2�́�1A��{8�o�5F���� +��+��ڦޘ� �+lu�V��{"����S��pD<&��?�!��Y�9,b*�٥�$��g�ju�÷�J4�s�5l�}�R�7E�I�|sR�~R��3�dx��;-�܁V��2RL\��v���z�4*��l���r�m�~�d����+!_�I�=Ѽ��]���*j��o�����Ey�~4��i�>K��4@�e�5��d����ƛ�2Z2�����
�-�:'ڞ�o�ߝ�%X)>�Q*�M�(��kQ)���6٨���
�_Ȼ�!��F����q�F��1،W�A�7h#�p�v��X�l6��D%Ҥ���_���j�>�M>T��chu~����c䗌,�O��	Z{�v}[�YqN�^���q Y;W'|�a�O]pliǾ!6�_��e����n8 �<S��8'�œ�"-~�T:�O���y���ƹ5�~J�_#��=�<�S"����$U�3Q���.q畆0�S��1��;P�;��g3bWD7vǫ��K��ᄃW���Y-����g���q�)�x0���s�> � �m/t��%��z�����L��d�9l�^Zʑ������9�3&
�����1��)Hc9O,��	ъ���Ї'�Iy�x����L�+�M]f��'�4:��<�4�	TN�r`�A�4�жI%7MuZ�鮦�iEW�G`�$8��9��QJt� ���xS���4�!��K]h|M�?�=>�އ�:�h�%�,�;�ș�fϐ��=l� 0��4�[
�Z�a+]*�d0��kU`��-�H]���31(m���I��HK]?�ĎJ���ZN�24�8�-o�z�m�j��*�a���y c�����7�����N ��5`�$O,���T#	"X�Z��s(�b�lE�m	�-�a�j�`��F[�o>p�PmXH��>���	��9ܧpBǏv��V��X�{�Ǘ��C�n<Q�"��ܫƯ��H�� >M9���'��Tc�b����{�Wt1�܌�QHO�T��|�ٟq!l/o�g�G�{Z����_|�+}g:�m�f��e��^��U@�����P�S�����Yb�)�I:��B�jm�a�	B�爡X��sV�,�G�<�q�D�0�3R;���D�>\`��ɞ��$�bV�6f�����L�u���)n��v�8����'��V;��`��h�\�w���~nY�b7� m��_���1���[;���Vq\��S�l��?4�ǁ��Ŋ� �����농w�N[�
K��C�MSJs��I�	��y���Q�<���R���+�:qi�Y��ѳ���j��4�mKպ�Z])�����E\���2:�D��D$�qPbN�#[�͔#�(_�X�MB��ߵ�e�+N$����m������d$��FV$��W�=��z.����h]��4p���i�����h7�:����� �3I����^�+< 7-B����&=*�`m�O\�fj�Q��̚���|%�g�|�x����� �V�u�Wy�����qBF(P�0t*��,�i~T��4��/���xq�x�U4դ��H
�̝.(W�i>U7������0c�X���x�C�J����e�핿}�f^�Կ��?�o��Pg\q��y-'���L>�KA���(-��=SIC>�����ᓨ|y���}�g�cΩz�j@�#�'mnt�5.:���C-L$��uEHQ��K��G���f���+�!
""B~9��-;z��H�z��F��c�?K߿�W��� �zI��^���J�k)�C��7{_Nq���@�a�d8���%!�o�3�3��!#Ƌ�&v�����@��D"������C���S�����de?����DH���!��{*(f�rO�5�,�hIW�D+���Iș����	�;}���##K`?C�������>]�SD|����k 4������I�����B�H��6�<�<�7L�[����o:�p��)�+)GB��ǣ�%y�6�X m��!��X[@`Z�-�$�WQ\Z������dF(��4qS���I2���E_F�6�d(��z��vc\����?��
�&|O�c���4�g�Fk����Ǉ��]
KG��؞ש��^���@�JbDN���<N�p}�@���4�\"��+[>�1U"�t0�s)+��y�p)˞��� /	4�]���
r�J���p�RC�`����dt	�+���#P�ss����/慸�e��.��rZ�\��9�܉D��sT�L����Gi�]���T�!;�>�u �{c�����"w1(`H�=�d°��a[���Z�,I�9XB�F4�1�@��&��%�+|ɞFRw>�e��ر��I]淌6��k<R�| y
-����+!<��=(�]�%4v^�Ou�q�=7���*�Z��Ya��8|<�3���pE�8b��+��Bd�lέ�"�}�$K���!����5޸(E���
6���kFڛjD�^C���o��`��U1���i�40� ��/Z62���~4k�V�Leu;�ͬ�i���,"�34�l�iۍ5Q�E�0���)Q����:X����u�m���)�1��G;��4�����T���R+(��&a�?�W�D�k�u�;�G�$P���0.�Ҵ��W���i�!��Vjg�s7$��7��ޠe�lF'Ŧ�����F~?E��b�8A��@'p6^pP��yG�<��8��~jv4��P���_km��EeK��+�:�"��8�ŬF"��������8��J� �Dq9�w�DAc1���;�B4V���1�+� DS��<(�K�&*��M��wC�E�c���@]�Tq�7��EhK�ѽ��6��H�Z��z�x�`�^�{i��`��˗۩���w���{3F��������T��ǈu7���#'k���qdY1e�DĽ4#Ņ`�ɏ��3�/iP��O �J�?8��PjwJ�֦XI�-�w!�� G ������o$�tmv3/��A���n�=u�1���B*����h��+���dY4���߼���[g@�c��/ےš�b�;,��a:ۤ߼��'�����GF��xG�VUQg]�װ`���b��-��a~F�����Л������	�AG1A�D�R�o�'2�^���v��e���`p����X'�cٶajnb)���G�0j��W WP{�bHv)����v����50�O�aZ.S��������/��X�iYﮏ�Aoy����*]$�Q��=h�l�M9��;]V�6}�m���Ϭ�.�d��9�y��w�����j3-���8�̻�@`F:Of&�Q���~_}}���>�`fSˋ�_*bo�a���	��w<�w�d��R�ڤ�yI��5�GX�]��K�^<5��S@���І	��J�r�D�S��<��%�{i=�FS;я��p=Ͱn��&u�9\�����O�mc��*YD��rQ4DC?�@S�
����K��N@q��߹��h2?�N�i�zw���E��ɺU	R�I4� �h��
U�Ak��|'O�j,�����$���QK#<�}�*?"Y���Y�Pf�jY�"�P�f�9%������k�	v��q[�kΓ�Ͼ`=��l:4����S�~K�̾:G�5+%S�=�f��Ց>���J��$4�=(A,��g�;
��RG�	*:t�l_�k�E��m��^
{�Y�����q6���$�@ZF����lĺ����Yu)�9��WƵ�
p�_�7w�5S����'��D�|��Q�VڹZ>�i6�4jx���>]�=!��\�.!A^�+}z����k�;��
���o�O���j^m�9�!"�|��쏔T��T���p]��t���a��tKa`b��z�'#���*p�N�c�Ą�)}Uw`r+����f�Yb�W����qU���]��C���Ls@q���d��JpG���S-�f�
?����a�U �1,GT�m�ls��f���0�$tJ(��!�+��gt��p+�a�r���8���I�u?4�>jb��;K��8%����~`9�Q	w�5y���Q6���,5���������䣕|��<�!��p�W��"�OD��{^�ΡL��.���t06���e�`0�`�+��!vX��9jIڇ���&���V<��U�-B�s�F��ȩ�˜#�K�/qJ��OoGoki�qC���H �� ���w~;���6���2��N��,��(Qͺly���7�]�y�Y���Z�C����f�\��5���&�"XT?�_b�	;;��UEC���g��G�
��e)�	[�N�ϡޗ�H�a08��<L��WS�<�}�@��q�ni�s
�]��<Cn�.��9��0�p}|t1;��J�:�h�6d^�C*��Kh��w�������������g�E9(�)>Vǿ�������9l⍬m�5I�R�-#|t�� Lg�鼓|����{� }���F'鍓�sT�<H�r��N9�nF�c�3uz���O�5��h#���D���"h%��7�%�na��d>�=��W	�=��|}�il��a�L=�:!�^}n\]�q��y&W)�uEK���a���D|� ��J���2#ےR�eN������e޼�ь�-zph �s�$ 'ʹ4p�Z�?� l�*EI�氳t�]ӱ�Sj�@9\��'u��J�����WP�'Q}����@�K�us�{_��������W����q��*t�s�0��q��Ƶ<����rϲyR[�%�+�<��v�!�ǶTNA��U����Y�"�P�y|9d�s�畊�abP}I�zed�e�k��7�A vyUy��'�6�W��Ut�`�>ڱRˡ����,���+9���wܜ�{0w�R�Jߘ���-e�Sok_׋o/�z�Ւ���
&����*�3ڀ�謐/E���HL����X��o}Z�D�iS��$�FI)�F;�n�H�΄�c=��=���Qﲁ��ּ@,���5��
�dnƉ��˫���V��/^��4_������/f��G�����a�����I]�s��aP?�Y�FB� N�Sܔ���#��� ���B��<X�&���]��� F� � ��H����ҡ�I��[�$����L��HA�3=��g�d&��z��}���"m��KRh��@����M�8-��j��T>o�
����	q�O���-s6���&�8�)�@%�Q:�P0��M�������@)�6E���w!����	��6{�eϐ�F|� oK�v��Ӻ-����@�IME��gj�����q���.�Wp�a��T	 4�r���u^��$�`�t���Y�,��e�TpS��r�4@~�ȿ����NK�#v)�h2n�;.Um�������q���4�0_
�E��?�N����ω�G��>���ڲț�B�DkNЗu�u��i���C¿�v�yٵ��\��e%���2�~.2F��̂���T���pK�9}����(�-[�a�P�)I��^���:�8^-�B$�e���M�5�*c��Of`م��s�[���Ρ���~�=��TD�v��@{�5����6l�=����ײNu����	?'����I�OHԜ��Ⱕ�Gs�3��7-�.����UQ�����Xa�mK���ͽ;-�ѷq��MzC�����&�#�בf�u�z��g(�ۨ��%����SE�}�l` 	��"g������L,/Pu��'v`/�ui���"Ot��{��n�9Ǘ�����A,}�����R�H-��n�4�����;G�7W�|	�N�=�jha�|��P,�a�K�I��x��X|��� .��j{�`��ob�<�v:��E5�>ŃM��R��� �6��t��iaf�7h���l�� k��uSC�{�q��yA
��b����Kw_�i"���%�s�악�M�<��zB�jx��ҍ���R6ֺ���x(�Z��~��N��e!x���X/����y�h�]�.�)W��w��R��\�q{#c�?c'��0�]ZQQ3��YJ�{�kq��rc~����b�\n��Q�+�d�2pI>���D�J���=-����d-�w��IE��-��f
�ݑ�aC�7g� ���j�Tfc��W<��A`yw]	Q�(���i�M���L�D舏��ipb��%K[��G�~Ic��0=-��H���Wxl(� d~B������������D^�y)n��I����B࡝�0���Њ�?!}O�����?���0y�`�(0�Ѹ���[q�����>��)lD�[�=�2]R��gǵ�`�#d�L?n�UK�,hx�G,y���s����y��m�f�	�hjX>�O�'�y�������*��KQYcRnP�@���pU2m��6&����˦+ ����$pT"79A��ԕ؆M�Dݱ��R(���:�t/ڭ��!�A�����;6k�?&̋D�*v6;Ň�+�Ɠ�=q���W�Q�/U�q{���b\��}mt�f�+��HD�&�G5Un-�c�~\���E���yO|L��>�"~�`��Q����m�sI��m��r���������~�u�s
�?{]�}7��4�5=M���SN�	'���M����6EK��OV�qA��Nb#w�$�6__Ѭ{���u��D�'�Ql�a�������I(�3���O\�/��3� ��,m���� m�U7�$��E�[��cD��&��q~��J���t����j�[)��"^w�6����v"cۼ �au����� �4{�g̋��Wn��7��&B�~��Ud�4��O�q��w��G�¤)g��\���R$�����Ѭ6mɲ�|5g��q����e�'�՞~��)�$z:m\��F��pw���� NsO.�'b� ��Ki!6�z�N��E��۶~њ����I2e|�#+K��C�/B���oI%d�̘��4���di�q]!��=����Y�מ�aH���A|{����8s� ���[�{*ӂ!Ɩ���\�����L����Dr�H`Z�e��_���zr�b��<[�r����aʸA�!��w�!��_�r����@/]޿�8Z�sy��#�0P�_|ə|��������Oıs��Lq|L8�a�*y�W�#�W�1{u�}�,i��.�m�YO���