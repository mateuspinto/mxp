��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Z]�� �+��+6�8�)�2�<��?:���#�obxt$]A`s��m�uJ	.���{�fd��_u���W������U"|e`�h߯q�|)S�X��q.��A��c��ߍ2}t+��i�k��˜��7%2)x��w=�o��6�U���`����m��� �G����]T�?�1
H����Y��р5��!cmǛ�];��uk���ȇ�6�r�y
Zwu�ͮ��$��X�_\���|�#�)r����iȖ^~[��	��yxp�ch��˙���o�oƞ�RYk�D�?�=v��,�Cr��awuT{�R�s�������z�9�c��UHP4.�E���ԓE+;x�/�)Ztd�,�؀�}�RQB�r-N���f�q�Ib@QU<TB�K�v���@�����ó����p$9�'ߋ�?�ؗ� ����J�g��3�f�.�E���`$x_+�Ѕ�yFU�A���0�����81]����x����Һ�Т��I��,s=�����
�A0$�GP9$R����N*��P	j{B&#3�Q��3��HC%]���7*��	���  4��ş���\�	Ia�p.��eH�(C��|���u{h�-�:7X!L�H�� �`S��L�Ґ{Œ�p��c2_,��d8�Z��ܷ4r�c�+o&��v|�������ޕQ�d!�FR�b����4�R���rF�o��|���n	k���?����Q�Of:����耇��G��TA�Zu��q,�z��/��r>p$�X� D�f��qI�S1��-ꁳ���\�ԍ2~�S$�ѹ���G'�T?MD�]	vnxh�����|'`�0}�����kd#�C.�����һ�N�P���P&���h�m�����| ���@��`:c+�Z~yMzA��P8�.(�c�kNk;�v���ۣW&��1Y������D���4f�Sv�1�KAp��-Xfȅ,`�7kmN$�,U�W8��϶ǟiR����s���|gbūQ��͜ldA~w3ͻ�K1p��]Mk��}N�h!x�H��rn�w38��؉ג�4QDH��*�i�����>#�i���V����L��9�\2
:N�@o�RQ=�n�L	c�xʉr3\�^/����Qa܀;�fMi]5����;X�G�/��Z�P�n��K��kBJ)�t��)�-�4xԌŚ:�>����w�S�}+j)����y��{���Q(�W�h!���s5�@ NDY%UZ��q�˂ln��s�{�er{y����[�Z�o��r��Jr�����
����%�����3��5X@���F!��<L��#�z�?���[K�!Hw;��� �`^��B�(�\��"聋��}e�,҆��X��e37������i��d���-��u�\y����Y8����2���_Y���K�9!���qm�g
$��`ƞ�1�'������L&���d�<��_?��5`�$I�T{�/��m^��!Ş�n�&���P:�.r$T���I.�D0�ݸ��k9Pq�@{�����+�ï�	��bZEtB��ߛ�'t�X�N��x�;��*����?�@a�0{�DtK��������F� <a�Z�+u^�O�Ɏ����]��~�Z�-��-k� �4�S�>?��I%кev3 `���]��&�о�ݲ���(1tʺ����O�*��񑚗�|�Z�P��\���?R'�C���ic��נZw�w�4ל�e(Qy�(X��7��~Pw{(u�I\̆�G ׌�d�}�A(]�fhC��';���� jˁ������۝��]���r-���B�"�T%�bY�������\<wCV9������Z��|���cg��ײ��~zj<���#�k�6>��5�]��Q��\���}2�>�����g_Ohm������O�wʶx���	,�`k ��.j���1Ƥ_�۪	lΩ��/z���j
N�CV�V�R�\9�3���뉊�޳��b�����m?��E�؀iĠR7�9::N��i%�g��o�ᘙoǷ<�).%�1b�]l<$Q�����?G�D�6A��%\!+k���z������_H>xÔҋ���&�$x=Óo6GLXB���Dk����`M=����_�jdrKɶ�J�TGA���PL������a��.=��9��t�i��������sdhHݓ^3/GV�\1���&R��2~ԅX�e�2͢�F\b�Sd�椰u���,*H��0[f�~�qӸ�X������Un���R����.��?�׻�8?ا�ϫ҄����C:�ǱP��)��<X���;9C\�iA�.�����x�(���g\�3��$������.�;�E��+���+�GBY�M����-<*���zcP,���|����V�������:��M��gU��dA%���T���7 �R���Y�Կ�[� ���%��R ���������+F5Pࣔ⚜mZ��g��b^���[���woK���H��~?J�3��s���T��<%��L�!Z�m�1��%�����dU�r~�Q�'�h7�H
�w��[!�$�߲�!��J������M�_/��~E��a�d&9`��m�x�Fo�+�НvD��t� �����p�H�zY����-B����;�������[�uQ����/�_���E���W5��|��+Ԋ����\����՜��N�`e4�b�
.�K�PㆁM#S��䫍��h�RM?�a]���� ��*��N*��LM�\R�QA��. �V�n �癜��޶R*�xH���G�r�v�	6�5��{����$��L��[�
e�n��U�ߢѤ����yPN|�r_b�|�f�zZ�4h��{1'
�]�
 �^۪͐�����,cLPU�'�SU죀���3�|�Jj���%ǚBU�B9S�g1b�;_��R*.q�-��E��`X=�	Ò����[ѩ�F�6��#�R��S�c;c`�v�);���E/��-^�#Pm�S=˭dF�E�L_��A����0�W`��^[��F1zϴW!���z"�S�8�v������Qդ�<�&�, `-j>z&Ot���ڲ�J��z��B0�uBp2P_�&7�9�������K4��H���T��г����s�u��e�-��v�昉5Y)	�[�L~�o#�X�Y=)��ۙ*��^��<��� �˞+���-�"W�9k2�,�Q�oQ�6����P�3E�A^�����ǽ�ZR�(�'{?��$eL�[0����{Kj�w�T��}��͇�:*�9B�W�F�F��R��܏iOQ/��)H�Z�l�Py����E,&?�tz�����?�a���ѹ|v�a4M��W�=��Ө�n9DE��ʄ�=��4@���\��A�a�q+��9�������1��	4�Ti˞�PbF�k�Ϲ�|�д�sG����U_���?k�f�^�[�#�(p�Ġ[�R�dN��*�ɨ��ٟ^��x�;�u-?�1���v�)N�~�J��0i~m�3��ʳ����jU|i��5dY:�}[�0䓝w�r_jn�	v�/a���|�R��]]�<�t����K��� V��,��5�ǌ�9�Td�ܪ�C�51��}%��o��>��}S�@�}�`-ʫ0�+�O���X��
=1C��X����N)�:��F����W|�uj�QR��.��)4X$�m�A�et�^�J��� ��� �"Λm�Lo߾���^�o��:X:(�!�?j��s�ȃ?��V��GI.ۇ�w���3����}]<܌�3���K�B�:Xt���N(�T8���Վ�_��E��s�������d��=����rg�������{Qa�k,T'J���zU�S��X��Jb�`K㧗��n�͂˲M_���������<��,Ǽ)���F�M��*5�Z�����'~����P:�bư�C�ʩ��I%���������6���=�v ��ׯ�鰂�&s:K���5<��Q�*��m9��f�_�^����|"uan+& #̀n<(�A��Ŧ����$�%�NR����f<d��uiHi��ϰбU�( f���[��'�&��WVm`zVj"v����zQ`u�Sa@ml��>�vގ�8��7���߬���X�)�����nz���}�#w=ڂ�Q�hSW�˨W>.5�m�NP��d��w��]�g������|z�{Gz������ʸ�����vPa�j��s;1^CF��&j�͞L��0��C"/�O�Yo����-t��J�����O�8hTC�fĉ��ܾ[]RA���\ ��CLS��3�#�:�X����x���ċ�)�(�Q��������|n��$
j�Q��igCMX���I��PO��܃�[lvX�5O��5��`8��b;��$-��5�����؛�+ɍ�0]di�M�*�!�M*�!p�����m�H1Ǝ؟u<���?�z�yd��љZ��v��a���q�TT(��!�_��������tǴgqM^����� ���h,��fL2�NrҜ�y�H�u��P/&#z(�d��KAv��=7mB���ɅF��`���Y9����aA�������E.ͬ{�Ll��D����X��{�U1�4�����jh���`��
Q��<�`,�3ď�2��߾XxU�PO�L�6�F�� �d��ls����^&�Xˇ�$�Z)�C�C��]��>���ٟ^��p�*�+�ZwD{��GA�#�_���eژ�xs�A^����G���۳�;-.��O��P_9j^J�_u�XDy���U��(MS9�P���OB|M���໤��<"tbn9o~�ȸ�������y�����0���^�V�;j1I��FO�����uɑ�KA�2���J��π܃P�DL�
�9@���Ue�k�����x}�H=�>��}B��c���I&v@�`��	S�s{��������M]�Il�����f��y�����1yU"�Jg��g*4�kNb�{��|�\�(�)`�j����<r�| {,�n7��  7;�P���Vnڙ�!�Cs9��!ʒL�;����]%�RS�MI���8��e%�M�����"�CԼM��o���_V���f�&(���i6�F���`E藺J�K��'~(��_uE��"qtɧ�;�u���?��S9��5Ld�e�}��*@C��s�p�1Y(/�m��@0?�4����B}�=/�I�P���������N�2T��ڽ';��Ǡ���B��4��d�����1�}� �iIC�$!<��I2�+K@��7���3��N�ޒ�}3M�	C~;�B��)E�OE��bg��W�:ч�'�P!����z��q̓�T�7Ub�g��p�Uy���P��%��&�i�5��+?����%[�{�EM��S�����dD��7�èR.��W"��q��N�wfB��D�o��>n�,5���>]�k��fH]f�}��lI��ͷ�@RT�#$y�<_�G]�"\�F���w+$�H��:���zҀPc_ �(�i6�;��J���jj��u�ȧ�fP,[��mi�6�D{�y��2D���|�r�8�ptp��5���i��*�X7�-bo�z��Ǽ.��m�����ϗ��Q�5߽�5`��=�F!ms�b)+��x ���*hx�2����֦��X�Ϸ�b�LyE��gÔsݰ5Q~|赩�;�;�u�f��	�L>��µ/�]��h�>:ݐ��i"��l��~K�Pvڪ-J�Y}Z�yO�m ����!���=:=N9g����L��/Q�+���|��[�U�=����4����O=tW����0�c��p�$饖�5+s�h&��H'��O��֕x:x�������,FU�*�q[��0dLJXv�[�>b�g���;�I^�pF�9���5�U`���@�Q,���A]�3��(���Az'Մϡ3(5�H~W�q�,���Ŵߋ��5�[qׅ���)�=)�K���L�/�6�:k�
�э��0ŲPa��,��A]�5��1y'�+K��9�K�(���塀3S ���1k�Ӣ�^�O�>u7Z��+K"�Ȓ������/���#i+.>�9��(��A�qî̺sdu���b�
��?J�,��oK�qڲ0z o��Ǩde_r:�L��ponm�ᖨ6RI)����DD!��ȏagO����0tǷ[��X	 U�D��Npy�����y�D����<Uܞ����i���o�oD3�C3�H=@�س���M���"��#cT�wR(`'g���`.c�?Ď��;��-�Ю�����.�W(B�jZp��(g[v�^X4��1���'��;�#Z�?|^�X���؀3�-����Rr���]��U���NÎ�����l�:m.&3@v�B`WhL}g���P�$'E}A_@:x�W ib���^|M�&$]Y�MQ���9��9zISd<n<;����tgi�����W��_ =������)3��Cӹy��E-~�N�!FW