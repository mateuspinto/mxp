XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W��d?���)>�GF?�&C2ω�'~Dnt���`+�|��P$�5�^{�%P����f/(`��Ҍ�dE�!���0��5Z�5҇Xm\�!o��F�e� ��gx��攩N&��J��/���#��ɗ�G�s�1+Nb�J�����c�Hr"�]3����G/y��[,���Y������ƨ��@)���, �����I�����!&;����V&���͊"=7	\X;�f���T��r�7��7�����]O���"Y�.nFOt/��c�v
���ɧ���eCnY�:͡�E4�Y�0:^=,∑^�CV��F"P�~G
�^ڑd�B̧�]E�2�rj ��&��O�*B�;��=یk�G��6�(�
�Q�����M�S2t@�b/^6(�y�ĎVK6�t@�:��K��3���S�Ƙ�p�r#���=1��=#���1��TH0{�Z��7߳I���jk�6�g&Al@��f�vy��c;�חC��+
U�7_߉G���q"�����c:�	��)����eG`c�24k��ه0�8��<O��0�[��x�
�l�K�?�?\�]π����lԚ����;�[��y��m������▥�1��t��Y�yӘ�F��֟�M��ȧ*�S 6��{�۵��кm����)P&�Eӛ�nxФ�"�'�u��e��#�>�5ʐwn��I�F-�k���9���$��#�~-���,lf�s���N?r�i��8Y8o��M��D�����^��XlxVHYEB     400     1805b���v�(�A��5^�-����P����z��M��]���6rw��G�����2��}F�"W���,�ǋ%�:��K�'#J�5l�;�Zݖ�JgX���X����dŉ����]*�R�	��h�ר��B������2-�3	|<�X�d��;*���'�V≏
-�B�ԣ���`�� �ܚo;���KC�ˀ��4������C�
<cs��o����c]���8':��;q��;�!)��FR�W`��:`#-�<V�]=`―3��&��9;��^Bm2�#y$O���QG�As�,��ݓh��Ǥ��B��S���r�Q2�}��(��
�E��ɓ�熣�{��s���W�B`ŕe�gx���wARXlxVHYEB     400     160&\���uŕ	�9=�%�c�@�%"� 춶���\֬F�oM��,�r�<���5��2H��=S#���S����^B�)����\w g�0�>���	D���w�|ڿ�����Ɂx�*��:�I%?w6(�/0f�~?�sJ�»uJ2��qS3��'ڮ����Jj��^_]ڊ��s��?A��٪�B��_x@zz��c�~�&�t�[ư|5Gc����d���{���� ���cQ~����ɨ��nӴ�e�2���r�H+E:�ɲ.:��Y)]��+�{� x�rL����=C�b�	�R(��
0%��͝6ڹ�Ї��?Lu-���'rw���󙶑�XlxVHYEB     400      a0F@�9�l!�J�6��G���;𽞍�A���M���F�71K\�=� ��p_*���t:�w;��nvPo�>��IŻJ����@�!���1LHE�� ��~��4����5&�7�xŅ�7�~�ap3�)ϳ�,��Y�~8�xÕ��ϓgʃt���XlxVHYEB     400     140��bG�E�alk���Śy&C��>ɫq@�'��*,e���[����E�*L�`GR=��,{����n�;���)�����3?erj�vw�����3�����;�v?@6��N�@\G⋍�m3!#O���t�KB�E���B�s��y�b����I!��X��O�iX�+P�; �\����Ƶ�@���ޑ;��&���-�dl��r�B��˙9ӵ��}r�b���ڮ	���*L�Λ�Y��pIYαbU���o`!�jx)*ˣJZ"2�x�YP�/*ݟ
����+�8���k%���o���L�y�:��J�fSyi��XlxVHYEB     400     100<#M��l~��q{�g�_���,�e0c7M7h��<��h�������������,��1�zTd���J9
�r��r)�hk |q�}���B���V50%���y~���I# ;��gLmm�tmw��=�&L����(����_'�N׻9+�`��sū�ɪJ�68 �S \���E��[�.��� � ����b&M0��]��Oc @O۞YF��]�E��:h��c�z�=��iCX)t�6m�oύXlxVHYEB     400     130�P`�?�@?�����8���)���CnK�.�c�^1J��C�9W��a���6��E�Wx)rʞmw�yBZ�	�F\�З*�e�R����CL3�W�� q��'DO�F�E��6�E���Q5�V0
x��_no�+�8'�ܪ��)�Iz֗��-S恜ZB{#C7��, ���/.F%��VT�,t*���7ঃK2�Ll���XT-�R )���i&:��]����N�?���EA�	ڈ�@/b��g���L��[�a���na���ȇa�1��%�zh���<�$]���bL��0[��XlxVHYEB     400     140��n�w/Oo��	4�]�Q˴�2�"5�{j6�S��n����g��g>/�C��F~�-p��\��8�N��{�ȇF�T_����bp�P&P�[��(��:k4Z�0(�}�1׺�;��h �����;/�a=��]�&��*p��2��ʜ�^��������
�p ����En\9N�ix�'!�mq��e��0J{�<6� ��|�rõ#`�@v�Hy�?PZY��S�2�����mJ>�g��ɚFt�a�
�]޳��TOh���1��j���f�1?2&v�[nE;��K�j���X%0��O�;:�е�&3�9vp����XlxVHYEB     400     120'JX�
+n�9F�L��e腉��{e�^ ���V-܏�u�y��-N�1�M�G���#�����#F�\/���A�Z��@@��=A��T܎}����~Z���׆/��S�ۆ-�ϵ���2��A����&���<>a�օ���8�T`ЋF�[q.����c�M�{�{��\�⎚�$l��'ʈ1rn�Hc�8�e�؍���@�z�! �<d��jp=�lYƆS[ĭy�q�$p���I�+m�9��=w�lZUL�_�L��+AO|~��B�x�lWO�	��XlxVHYEB     400     190�ɽPaBZ���|.3��_3~�b�b�3TB*�rv3����K�H����G�w��d����&�;@V���z��H�[+g̲��ބڶ�Ā�X�[�K+`�UT�|:�Ou�Q�9�Yw�������s��{NbP1ݕ�����lJ�fb?ڥ0�'����Ӑ�S����N�i@@[�Y����4e����X�4�W�$�@Ծ�<�i�N�#�qE�5\)����ě�z�i�g�v��u]�U.��Q=��Z$VW�ᶾ�%-��rm���/���L)u��&a %���@,���� ��J�[jE������h��T����ƫ�y|�I��|6��y�8e���� ΐ,���2j�����FiX� ��;�om]y��l�v�v�� �|��$�|\��$XlxVHYEB      d3      90m�� ?�� �bJ"(����7A�ùw��"��.��)����
T�mɑ�����q(�#>9n� ��Z��$h��G� !n*`[ ը��ez��v��g�����*+))yG�$C��ۮ���~1�G��!�!u5Y]�k�\��0��*