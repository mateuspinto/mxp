XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �Q'i��L>U_�ߟ�S84i��n����W�k�z�&�Ϳ�16�=��{����?�s�N�4d��&�.̗Mv����	&Ia�� =*нR�N'��N�rt�}��$����6{�����"TR���Kf�� 9��B��豃����_�GU|JNV������"�O<�o�e�R�u����!Y����Y�ÞE̮�䒳9#������o��+v�4n���\��(���"��W�d+~ƹb,me��8C#.�!�-�v���qD�6��k$��C �_�.��'j󄰺0C�^6��D'D��4Ņ� dr�{׀_�kgJ4G�r�4K�7���?V�D^X�Θ�]���\��-����;�#�I�ڕ.� Ƚ�p����� �<�'�U�]G�^z?&�{TOB��u��~>�p=1%x[@�g.�l�H���(��d���,z�mG�x�����0iR�5= T�F5>�d���Ɵ�	��M����&,��R3��Sx�*щ��tK� ��~��K��4��FL):���0N�F7�4D�H�?.���2-"�X��M�bE���3o�2���:O4pU�Y����/׭r�T0��V�9"t�?nM�B��Be"F� �ɫ�F8�����#x�;g=�����@k��]�6ق��7�0�Hc�Q������f�%j���|��e���W�_'�������	ziR��Y��N6�����xEdNqg`γ��ٰ��i���_�-|�^8�AY=XlxVHYEB     400     1a0&m�('ͳr��Y�%���iy��i��p�β���ef�
�7h�Jt�-!0]I�o*G�N���{͑�+�j}U���T�o����\���\�J%Bt_������끐~Cl��(�`Uޖ�ޜ�����3����?�"� QNa
<p_�<"�>4����6{^#��P�]��j0�r��]�[�q_#�q
S��@Kь�Uo �AGk��Z�]v"i�K�+���:D��KC`ĺ��E�xX��p���CZȇ���)���S�"Kn֥���R[���\>>�]�$��cAU�7�+�|��1��W��£�������ͭj�T�����J�����nE!9���F�[���]��G��5}�
�M`ު�N��C���XlxVHYEB     400     150���"Y��H{�ױ/�"̖�)�Ѝ�����&�3���,8��Aؚ�*0�.�PՓ�>��X�#E'1�����⼓����G8b>ڞ��T5А	�*�q�0ë$�n[T�s!���'g�Χ�{�Qxe�u��%�I�D|>��/�o�q�P�A�}�ǵ��^'�w�n���HB!1��X
��d��
�׆�W��w��pk[�7^u:%*P�x�:A��\4�Am�ڝ!�p�߬��o�T�~�N[Nd�Р�%&��`^�5�#��*�s�`�r(\>���x��>�Zt���pb��BhN�1P������4���%�vXlxVHYEB     400     190q>��TkVw�#dNpv�\�y�M�0\��y��
e���Ć� �e7��GW����s�gH���c�h�	�o����r�E�� �rj��"T^i�U�=#�}2�f�r�c�`�G5�����D�֫Z�GK���4Y���V-+�`�p�[�5�,�^����i9��+<�b�0�	�F4&�Fmu���/��W��}g᫽���K,�g:t�ٽ�q��_���\��x�d��`!O�����E�c ��Uĺ,9C�}��o��<!��'�c�������H኿�a)baƬE��<���Lw��أ�%�{$�3:_��=�X��N6�*7�;�#�/��<:�I�CƏ�τ�e���٘WB1��fґ�=�9L���\�[xXCſ��z���wXlxVHYEB     400      f05	I�����Pr�����Au��PpŊKޗTpѕ7ެ�Q2z�C���~pA'�F4/.W��v"��kO��OOPo`.�.)��>N�F�O�4�U����ĤQ�l����ߋ��?A��&��
���Q_�ր,Da �N�\'(���վ������k�()�X��X;�yo���:A��t��c��ڱ�����
�ច�L��O�q��%$'�s��:��h�ԓ�R��M�����nXlxVHYEB     400     120Fa�
ũ�m�h�Z��G4� iW�O�"|��m����������"9����ɲY��6�?�k$]�+��
�A�nY?�7��2��*m�{�!���9M丸
H$���R}���V�~ ��������|���S������i;Y�Ƞ~���D/׌��5�����o{/�Z~xImk	Xk�}���~��|)�<�l�%��F��n*|��(��sȬ��x|n�F�;/L�|��[d�e�B"%�����5�<n팻�4Se0��[��LԇO��g��P	J�XlxVHYEB     400     150W7��2{�ntII�d�+�{ط���X�B��꿏���/�u�H�n�w�P��wd��E qI f�*�4�Z���/yՉ�`GO��:G)�:U��[k�RvI{��_"*%��.�]^�+7�$Ҁq�-a4wi��}���$d�b��$k�<<Z]���g;j����;HJ�4l��)�B����"v�ת-�A����p���%ܡ�[�������V��SQ׸�{��A��`��r+7���;q�'7tq$�UC'j�]�Ca��6�Fu����.zx�ω/l��^km.�tH�M�@(�A�68�!FV3��ݧNdibqP9��(��XlxVHYEB      ee      70�%��2�\HId&e�ЪD�x����F��\��_���_W��%�^�_�jYA�Y皆Y�E >HY\0���(#�O8c/��.X*c�p��w�Ip�v#�h��ko�.5$q�