`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
j4Sah0l8p21Z4ZJXU8YCAL3Vf6ZsYRp8pYDA0O1yA1sNoRulEzjzWOeuR1eG/9x0MI4UNa6hCY3a
3jYzJLaDG1PcQPTqw3RA7We1L09QVsMVHcG7xZyfQBmUkc8gysadOXmVhbOoQSBgy0nqL6mqHUkX
pyZbJ7zOmBi7CzcT+iJ8m3FjNyQhzByQUqYbEFoR4ihGv5bPWoZmXVtrOkpz6lAeqsoSdz4ThNP/
cPEIbfsf4rQdPyl9ymp2KHdsc0A0WgfqOZHsMk1/YVXrA+/8XtoKkn4VyqUcx1YHcq+HTVJ0SLMH
E5LlvtHhP3AzDsv35ujgHUXeZwEkLzpFwiLSeg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="PPvPUqIpPzJUzy1FIRVM9+cIk3X955VRkcct83iQk+s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26208)
`protect data_block
SK5rV4y3qujshWQazH5SObcPmdAUQjwXSv3urUYN1UN+hjVCn/FxlZhoqM7JLOQv4o3IUMyn93TC
8A3by5djX31dp+/a48RbTiA1T1RNH2Q25oanWRkREqkfax84RVuwOsz7LIJLXuX26w6Lzl36qpna
g3MMqo0drWUPlIbh0yvlmXuVg1UcMUX+yd2gpWu+BVZ4XCcFx7ocyx3evCMtVD9F1ZsqVLC8OHGj
pVSmTsQyy0N5kYu1pmk75XQ8VVzR5X1koPHMNiO4zACB3n+iKivu7xwbi4+C+FdUis1PsMBstTj2
bV938uxZqL9B6f3s9ZS2OKlb7SwuKA5gNbmRF2bILCNG0zwn3VK0hsLxSwe4+Cqn0x2r6qMNvy0A
nbg/a1vwpvAfTvBT6haFyVXvan7vZxpNJyyMsYhcY1rgswuLnBEts7YYIMaXTy+lWegC1UQk4NMj
1LW2nUb9j8AWkSwxMZkShefpq1zbuc+CNpf2/DBcqf+ysmOQFJkSJk1GYP/JXmGQpqvPEnxSeXYn
8QZDoqMTL9AGbmtjoBnm9ZLcB45huxR/VwyEG3nMgDQJa+SZf687zSI9nXD1xYet9whAO86frz1g
ZyzKzSx6KKwvhYgJuw9o6CCjaWvckoPP5ybCnnGgF6AIicAvslg5zWakYLXVLgtoZ8stdtTPhz0L
+8feH4/npgSv/DE7rrRfUl60AU2czcazgX4KpsBU2iEu2H7ZLyrx+QzvbIyjDGIWgpgbn8qY5mrz
c8BInRPvZWdXjVHjUY7PdiLOUEA/2r22t0pDM2V7J6LNH3AGaIDehzxHSoPzaNPyf0X7h+jS/xCP
J/j+4RQx0W+IZV1a4cr3Sprz40SGkMfpe81AQyKRgaFoJHoNzIp8jfli3wF8wqRJEMvBHSPY91Sd
OZxBeuaNxVgG/tSfYYgmKOth7jCRvc5Z0zMeuk/M6Jn2JBwX5gmztVCAwxzIntf2FR+5TXQhOZVA
A+7gJC8IdnRCqagoFEqJ10/vKmyqulUVEHk5KJ8nTQi17D587VOmhzVIErPoTiBoZ5qOItkhorzk
2jc32UW1wWuqEJIxfPioL3oVhbIraHX0sOpBVXa0QldBwL+SLt8ADqfue0WP9J8t/l6712RS8n/G
a2kxxo6nfEgx57t0TLhia4E3jm2E5flfpF5nOZ4qm3UBnN48oZTXFPqJOrLAAtSnwSwTXbKeuXtd
0OjTGKQrWj34ILocVjRGC9LBjV8ZkpvRKkJPkwxT5WBNsb1Q74KM741CWwaSXvjwFvH3s1M4MaR7
N8uNQxURhB2Yvj8iyWi+QsjEwu2lC44JJzeY39IQOTud61SNhKgxdwvwaDUO3o1Je2ptMhowPHN7
qa/f1qTPU2IxkpHyiAp7xZ+Nzy3FD+JpL1VWH+oODmVDvn7qLMxtGDhvOt7YrjWpG0Ucqf0sd07H
caTnvBl2tnTU29kjqkJv5n+27PE9yKcvMlycGM8AAAoBeXu65nX1+99x+SY9kmQ5pV3Di/4Xz6Ii
CNHi6bKxqKifbKaGGCydqzytqiw0JURd1LuQemVtV4EPan/4yfj4ONwhsZI9j0ZfW/AhdXoehs6b
WO0qC8P2d87Br/YPPhkWI25eMSEX7dxR8eGJJNi55LRa6PjMiFnRPzVPY2z4+hjA+NHCgDgmWqUZ
gsacNGYPJ2tgiTSntqspfgmdIASvrjifh92WhijFteYdASNjDmcCSABy3/xiUbfPydiQ9t7kNlJ4
rlqZ7U/wPCzQU7/n1gExy1KbRUbv7NrP3cMEp3VxXl5Z2a+AtvnfbY36Si4x3lDu3WRDuKs3S0lr
jFbp9LCfIXvC59NxtKUtY9pw0cG2wBwD7avP/kY5e153I9abWHl2Av2TUy6rEXlVE7b6el6FRjLT
Bri84kZ4eUwY+YBO5f7a+D97VbzjFb9Qnekc+SfZ/1vB2t37E6vA3kts2/y2xlH9lWNCQ0HWH83m
R0+sR7m8dvpvmNMJsZTzNR+x9kgn5qUanYsf+TKzrS/1Aqu7amU/2125HAwk45PooKLQfhg6QIfp
yWyY24f/yE7hCc9IA6n335a9iQxGuaKWAETHJ0c8DswgUKV9KfeTJipGf1VCcOe8Bi22uJQIMS8j
P/fAPjL/E/qBNwt745m2ntyHtf8c/8HBTaYfmiB2iPG3cjRaJj41tdH9IFyNrLBssuAV4OP0iFHr
/0V1b7lKx8EiTn4yLOFXGFTlTY9Cx3xq7vFVGpn9tJOvZbYXqrN71Lalif98KBNDt4eyutiplDOk
M6QUwE2Oxx0RfqrSKregrhy22wA6gzn7IsZvCN/Lxe3mVpqfydyy57qdDdsZUdCoa4XJn5sUAB95
OcwQqsmUYFNhRrwmXIcRmDXGD92Jb6jlgkwyE+Wt5RmP6HhCT1pt/bms6CX/7286f18KL+Wi4kEc
JjmSQ4YjNgCGYUi00mR2TginmM4HPEwmRkhicI7SeC/fPnZVa/thXivMMKZpAOqSJV8639Y3bxFl
TvatnjgTwL7SwdiTMRblMqTlnWlSMCzRcbGeALRAxTxQTPTTtDgatLpqCXsGEgeJzrcXDh2UD+MD
By2Ch2CSy2oTdd8dfx4VnexzE8mbcqN/PSzNnMHZpLhOHx+P37w4oKaecljBtT71hKrytulamhSq
1B4BMB/BQOH4glVTZopZhbalH0gp8IaBjY3xjFyorKBOPIO4j6aBjZrwboaasZ+w3JkerSgiYIzT
x3iC7zIYdXLqT5739WAWrgi7xPU8UXjSyl8Kth1eI2yejqmAVUI48GTsTDEDU7RDPNeeqQ0TjN8n
ibPONqI5VNmevcDWkqF1e9P53MFCjDIH3ESW+6s9XrWuvdvQmJyDTA9coUvu0uaQmzV/K76Z7J3B
t8aBJTzNULyvELCplQhaWcNL3A1JPqFyJVhiyXDERt/OwzXqishZrHvmgwKI2sv9e64A9nvf7l8f
+nRcyThja7/IDx1LQuGkxEKWdmt2RKZ4jKT0P6QeigaTGULtTVv+TAq42tJPRX6fT8eB/mg27DLc
PR+Qz12uoaT9L8vrd0IGtxCu+ZUe7rgZ3/7cg/37LX1/B78MI6gUfl56mzS3U+1uHSqj7d7KZ0IA
t8u3TKWYQBXLGuXK/5XqJaAjoV+VjUHyMnvbWY/JBlYHEaY/JGDi9wg3oio1owmyvSQ9Jmkm4gOQ
xLL7dmm/rJ2ufyTV+8A+VnqfYl/De5iAHXUcshO6DidzcEUtLFbPHWyacyeE/TJvQQ935i7udCKu
b6tE/rTRuM1ZYDDKWl+XPWxYmjAoqpv4Lx+9P7n/c8PGl7mjvhzes1H1I+Y12vokY5iLbRxuvykr
BTDDQCTDmMbJUTB4SKxDjcGvl4YaonVm+bP85CP3+HQBOfiuODADbonCS0P1NV/xOOVLy8hIiWFk
Zr1+xBwsTpJlW1lVd8j3McPeqNm4zTCeBeOEZa980gJPz2dEvE2IKiox0hGLNyxZmekky0AAC9Bj
nqV41b9290Wjb32BmOs4PI10vUHKckjx4uoElzAcOMj4kl19S/zlZ5JNup7iZtAL+1jt4nbKMnZU
bNuY0JuEiprghr73Oqmb82RRwpY6api3RSUbWpYhmbLvusEDviVvz/CmsiX2ZU1lJcXUv/bV01nx
Yp7fvf7DI+XpP/GAcxGgj8cdGnars+91nEmk0OiBX7sxG6REB/s69lX38giK+Zrnd3FM07xWC8kJ
z33ZiinjNXgmf7uYamqRQLzAO3jvIf/fq9ikP8uNw6coN+h6bZeNwgFhtd3Qos9Gvf+RH5r5GBlo
/DJlo7ZQXGK38SCZGXr3E+gFqwjFRieZUpqWS9Xqpms9U2ARtt0HxqXMnqIt29uKq6uBTEeJSZ3L
enqjEZbPYO2IVR6DmkyOvPKcJQm1S0lxVRogWbIQbqZieR/1px4sxDslaot3HwWyn1eCOImvC1OF
yF88aobTUee5hyFOuakyIiUjuLUauXD+dlhG6X6pIpfNRmEiEebNgOUI/WyizT8gJxtHuc8mSmzs
Gl6gMQetYNy9XQ2XVvqJU+1PzjgIkL41uZOW6nwvZgmvI5cUx6QJsVRM20kmgdOtfyMNod4+YgaI
5JrUhpVPDlKWTlx1oxOAt2x+M6rM3iP50k1+y8mcm8wWDqMNU0D+wKGdqv1X3WvtrzTsYOe0ebzb
dyvkwwaxYzIH/MF/0ApugaYYSp3Dj4cu7jgjGA4mZXCOt8a5EIzloa9eXxpmmzSVKajdHeGOZ85M
wx+X0lgbJFwClUUctbVkWMegUbVD4vpESEfbAo1BgYNzjUnz+p0GZ+pBlco8O6m4TDhaELOeZ3g5
Y+2r+thFSh4XTwB0idePzZPC18ljw8+LoE7kpl7RKhTBbC4uzwEpPYMc3zRpI5bwXy+QSqhtepaJ
xm/WDA14ymn09AU7BREqclSZ9/DQ2K7tJmfZXJiencf4hMkAMoz5kDsL+ZcRrzN03nH3oy4CisOH
ynTCVujiUPUq/Z2IoHcZuY55y7CoWL08bkliZAGaALv3QO9jBKDTROXt9reRSU9mYl/7hF5gemzQ
YLq13f+yI8l1XBxM0x83SU05dIQd6Gi7EU5roTIqz2+tqsp6FN99/VZQJXSbg/rlTzMR0apTQCXR
QbXqnP/1SUI97dqzg0eoaRA45Mq40ikdE+9AN+8tmJ4f9XmthYTsJnebM9YKGmR2KUceVVUXg5o2
pUbBN+RjKHldcW3tKGlJ1SJ3Z4WBsoFeD4E7POd3kEBkEZczY/mP39XzgzbR9D4yH/c6CX30Kbh/
s9lV+6W+G6jYIw0ccpBpmw6dUoAOTnYkH+NODelaWoFSGFWyDv5eeEjAuXXAOoNP9qBWQ9CsF1rJ
zYFDcc0Ak+dE5IC5Bp8QDo4xwnCGkCnVkhG3X/7hn5X4+Zcbb8hSJ2zTjNd9wDoGtY+Fh90U+it+
mKxGI2VvpOwJgOcgYlPxVTLRmNzqYASna+vm7JlvdnRZYfPHxtkoAYMGW8p48LU9RtIFGCraqz7n
KcWbGBs02n3oKGjr9f4piDUPJkc8Gy47Xd99rqgIZvc+WIDIyPfvUlIzMVuEAbxom8hJNDz8aAds
P+pPvwWSkjGjhSOxQMiIvrF8p574R66VGp7iNOJXdWoxxqjP1suBeBVKvYYgUDIsSicQO5Z4ExIL
MoroBw0clsOg00c9OS+6n1s9157Mnnk1ZRkje5Us0jCcPXmcTU9clHhGkVX3a2+PjooyTaxeHy32
5+2pVO6tfxtvM6KavftQWFhF4r8CbnEq4fz8bGyG4vBEhINgzGAEXGdkeUgBfgIMvgJjQSp6Jmth
T751p7uqUpoTtB2ECKUogMQE3cY6PO3+0w3cz08oqlPd60TEbc4GbdFK9YxXaYQtTYJDuA+KVISQ
gh3cLmaWWyUM1ZwLD7ZHvgrCQuul+ByVM4dWUDP/El28YJ1y6t7MeGgy3E+0znkpoAxBMF8POVOl
8kS/yM9AIsWNa/0j8jMBS13RP9bsvNgSU3OCqAiDE/WI2LghRVJCkZCYPDXEQwwhyKDa1kNfGJ9d
t35o5vfIm4ULfLeVlv6qiJi5hKmh1paKsHJhbqlJHO+fkDOZUySHAp09+rVhL3erX1ZK+6Pojwn9
aBTiMfARW8lngVHO6qL896dzrfPnN3bfzRU9+P2RJ4QPG/bM6uvISibJPJHKFD0nOj1bRWeTzqc8
bxrrt4MGdqBJCBYdbczFxLUgcBykqw9qY1Yxt/zspVZyX1rDXAtp7HSVbrVzu38AtJeTo6OCUGm6
O9SnJy8nevUw0ndDjGw4d8WklKpshXE9wouo012D40NCoeJNowEWG4BnsZW8dnas+g2RmgaYcmMc
AC4TxUkN1xtGrEh996e7I/lx6ClxtqbmUemdDsPOoTvszuDV6qhzYv4V6PrVNRiEoQF9T/YvtkYy
Z2CQy998SBu7+o6y4ZG1o3xFuCTeHvi+6eOOFKO6A4wCOJ0EG/nyiJ0H/tK3EienDAaNIrTOC5rw
uu5HakS5nDvC3rPDC2oFSPKC0j1yIyvf3sVQ2CdHrLuvmHytIsScBGG80uUCGDN2Vi5b1fKc8oHd
AbhP8pkMB46MHQmfHkq7/no0jopeGCaAinUYFMKZkI/xdWffftjkXkxTFyTtE6vo1GYpayIvullG
tJPkJMsToK8eZeWyg95Nw8oz9tfVx1oYDau6yeHuGfEdg9EXnP6GXYIRc6pnx1ADb+/0ciNPH+O4
Ht5LCqJecianaYluHL+Y3IRuq1aIdisapM6eojhLIrOUbokFsVGTI6q934RJaVWY4XphnZJ0kOgh
vNPMX4IO+yfXZ/jKuH3V0RyihraWDeJ2SsJ6WR5m7SnhOCaCWwQGinqEyOLB0vMdQoUUZX8Xa/4J
hlnVm2lzOfOrI/5wGFCZo9ZOtyEHIe3dD5te7naPC3JChXHlAEelKDved2L0g+cS3mwe2kFj0rpQ
BFb08MvJXY6RQbqaaSNU9cZ/80y2UfJRbtYo7QlwJvbqI/HaQDI95KoX5i1ihILmzwq1s83noVrx
7KFv/2672QVnbIGpjl7sqT1gz4qnhx8UugU0Vu1XfzAJPqcRlvI8YFJYMz5590lgQqlFVgLuVTj5
yYd/BcnIf5vdPHsxdyn0hhtRn4uszuZLFX0uWEFJp91LSXkSrVO3mjxWNdZscXn2lV4sESo9jouG
ZLr03GLbhSQXQ3H1C5L4yHQEBvSj0svq/DBd/80UxVtyVJzndvR0NCi9JaHtkh9b9gdvXFqgthP1
aoWVYPAB6IO60w1E8nH68XncPRKRTfR1KiYQbs7lqYZvySnEKeq+VombC5QpEtMLx7v3pmDEnn9G
qQVCVFULup52nURrCbCxp8gTzsrGGSjzfiAsX1sGx4b9bxfJTzeYIsLkpxy/Lj3wp2a9J6XFyI81
KtdDC1qwBLEnL1sKm5BWmI6u3RfNYKXMwSzF95fw+BWyWizz18wcCr9bGlJLnGkOvY9w76qNLecs
hDzxK7Ilf1PbniRo24QmiW8Wq6oBexYUfuw/MZdxEMYwRQURhe9f//kCM8zDeoup/QVdbcri7S74
gAjD+UhCo/+pU1BHVGLvxeUnhVGwyeuwgSf2lJCNxP3T90BRafHrQuqeLfPzmwDtF2vR3VZfsv3r
ISGVEcqPB15OkiAKi4xxEExWPH6n2ICLhf03bRlJojn+2FnnayWpnrY7UThiijLvk0kjArqRr26V
dACcQXyAIEgPt/pMOEG59zHMBsieBk575MNFZr+N2T5k3ZD4Dccl2Hun4oMktKfnySM2DwbHzycT
2t3eHLvBCKUaKhpNlYJs5fRCqrbKixwPxJRs/30bvSL0kumpWyr2D9cVLJ5OzPhXHXAcHs06ujDK
GdW7qDQ3EWkp0xOaVJrM2PxJgGQXfpRxmWJVVB45t7BEDqUBGTq2GjgZRFH+gfe5Jy6Pfii/1KeG
VhxyV6i44LJebkbPQFMe+/LXXz/RHc1XzyG1+6kub41GCjIOkrYmHgT81AGDsIu3XvYMhdwrVv74
dXzE600bFQ7/TGZJNThftlolR51rRGom7pKIHiGPDQ0k9bOkBCXyGfdIN7UhXqvi/Q9CCycUW56o
/UWdWZ8OoCYLTiLn2DJ+qUwc3XDYhbHeuf002dfL6OLmYaG6IKzQSIBIUedcq54wKIRobAvrULaR
Z+/bgsHtHmDUzf8Bx9hufxOTR0kM4NoR6vz87kEG+uSy5q9VMvSI+mxZ/qBTVxjnG57bZNpVoH37
qiQSfSUYqbQ7/q2S9mXczGI60ZZZhUDVewKVpBVAlH9Otn7m3PZkn2XtiPJ+UQjcBNVnMcjpm+i3
g6E8wBbP6peX9XIUZ9RqkRN8CVom232hVXApypaDDRB3Oy5hYxBgpCKhaePMn1RYMOyl4gN6L9cT
dfa2Jp1pR+fwSElWrxWJTogRVfRbW798y9JN/oTRZyapmTwjNCjk9S57DudBkywHTTt0+qSlGf3V
IqSQFg6bUgVF8K989T45OHWZ2HCTV5w232LO1N9HgqiooRyyQGsavNkc0QI22o4dBpe6g8NSkIpF
8d83e6/eJKc9B/5bvwLBs2v0wClfihjXpYyy8QkssvG0qN5OQniVmuWVprjX5o8CY6EXDI5BSGEH
asDItFWnCgMFqcm1hih5pRZQNqZ2GaHvRiXO6ArgFSPQ9areCu43ftuM5ncUoSQWkTnE9UXovQkm
mSAVhAEkfSPdek8QCtOpBptG9ubKYVq51UEeV6dUI2ur6fg9brJTYzakzTo3kIi8ClVfTfUMJNJl
Dt6PfASBP8ju0+HHYg3oa75ThfuGdO0gHeR5goKFevm3dLLSNb1+1/WHcU/H0/WFzH49eYVrf/qH
vRZrsI4I+gLY0fRGBDSSto/JjewYDlionzqmM8ZDPZXqHw36JjmPyMdTXhLtmO0hdMWpV2vDC5ej
GIM2t2d7k6j0wa9FmpyekbeFOuSkTzqqaqlPFNmM8aHbuFY0/tTxKtgfPhqzHBdj0bGICGLsMNmU
Aa5/7uu0JMGlElnLjL0p6ewzkmq5rKJ5QmOb7SWqJTRiueQvpFcMY4L1gLw7irXuzLTEZTqdNeXS
pmEbk5TZAyNQ93PzGZ+F9iW54aSWIUiZBBCBBLnelvZvqJFaRDesxqsc01MYu2aP1NPifT4p45lE
qnyPLv3PI39oPu0d0Sfl2a5Q9nR+t+Yyi/PyZUkEmEYm+DdxDNXyzZKFor0u+GK3vBjoQn341Epy
v2Y63R1gDglFO+bzRsvq8aObM0qNYDs8ja9Z9EeruSrrOzobDb4Q9fV12atjRdSh7q1X0AMwyu55
Iv4CBW6Zm+1GHpxiE+PdC59LUyqvLvN6BQDLLMeu4bZGDprbTCM9HxKI3KGXV3Q3djQ1TeG6vH4F
kPFIwPKQRWwQa8SIseOuXhn74fzmnCXlaEfb5u5RtI6is/2rRu5rEoeiyY0lBZHUImBQiMvIlyWI
Jtq9UGjpPvqLKQCYcydTDV4ueFUQ7ICJeJ+getbE9RKJlo4TWJZdg1BCyf9olHGIY2oRTFUWIdk2
uyOalkge26Ci41TfDNACn3sG4B0+ARgPx8weAss4qaJ7raeY2wksNvf4NDuwVO639RMaVxOGIcuQ
Ej3qEcc8TFKzmZ/9HqNCydxbLB9h++Rid5qt9yC3905OwqtBY1HqgkG8Mh0cq3/mW+C37/XW1inf
uHjJp60P8joIM0MMfx/qG9a9vYM5M1EKnvTRt/oym/O4n83GGFivNnasjtP0SAxqHBumwVYg0xC2
MpdKj0bd3HZJUAOXpKRfrEnNGmAn/MEkDZNbsK0DF3rZi8BHm3klVn854Ni5lgT8U7Nw2YCjalUQ
msbmR4rURKPlux3wHDHfY1T3d/0v2m6QM2TGukP247/WXSDrp7DKUN76JX8Dtn3WHMOWxTA/fgOd
XhJ4cFi6pr6GHRgy0pp4YKKAPlrFqX5q3wneKwOoIWCG+HJVKBHG9jsFHl+BYctICwZR7aMofJzZ
oVkNVNv52FN+H1jtt+aHtplErUbe28ezTNXJIkh72DgyW6kk6M/OAUARkDmGCzMQWgQF3oWANlGD
TQFAJam8E9x1jzFEhvibgkWX21doYuwnjjIj/HPKD4LaO/m60r9k72CabnwFa77MP4LQToPM+Dpg
90zTdHMSYFFK65bZl7ieklyu38IGpIcXg9nwXKtwWznrMx9n3r2SF6OgE9IVnrCTAIARTpGsL0O/
7C3L4NJewYgFJx89hy/a2KvEwgCRtvIFsKyWUpN/NorzNogJCyIUlQ2lR/YCxiXJQnnxiujc8WAa
K7ZexZlbMY0fh7W16dGlaKuicMYUJhjmViK0UiPEIKRy2JE3aEJHn8+bcthy9WSbK2h8zt8/YShF
+NxlDdatqLFPN08MDcA1Fb6g8IWPxJWhBD4megIE/hiP6m9OThPzWdjENSleI/jg8GIlqoupXlQj
n+2Pz42gEGPhEvmqRsE03GRH7uLYvt11T1LU3zl4rfKwyARDAzccndWftby3oSdWA2i+jh7vvIZ3
pUH1WCc1v3xXXF3AXVk2EiO6D3VJdlbXz2jN0wYiIYvYdaoK69EE91sClcSnDrKTsQCEsM+i3NNU
8rjl/wIyA1vBaBTkeU1SvMf4n7JbYyzNAsDgMQI6JGSY/GFC+nmOGlc6KPZf0KV3BdW2coKstKXw
L9Sip5mELqkM3Kv7HVNipSjDvPVnxHTmGXFayONNYdPzwCJ236CduTnm2iI+MVptQOMQI+FpJzf3
tbo3S/haJNFAvU1HrM2uJY1w9kzl+aNVE7KXR2dF7/vWSZ7rSsxGMufOL2UTZAVKoD7Gfk1ennNM
M8DLXJrAMhjsFi7aVApfSkKsz6yfY4viN1WxRTP5XC2cO68I068kCq/3JJGshUbfy+dxi4ZJSR2j
ZyHC45QNdohdCtfIWXXjuEGK8mMSf5Pe/BJqBpFL/HqZyX0HjTBX4Q77WMLBYLcYDV6IgCOhT9Qk
JJK0QT2lxa/IRpAxyrbuACHq1BnKtcRXajbwjxGalr2dlXoPKhuxYFPQU0nlGo033Q93ubbWLR5B
OCznKXOt1Z7oJOEVeZ7CJsjoAGJdsT3DewAlhwmgJhk5rV9JmU7H3z0RrZtVCYRl/HX8sxJ+cNXo
U9sh1QMbiXwiBRRnklLu0UJ9IqQoM+RsFXimAWomFed0D8TuTdISQBJlijKp7+QEf50yZNHUxuYr
Ft2wmb4CwnGf8Fcna/L+qy+B7oPcMzCzY+ZkZXk8nq2FFLkOEb5YlOH6Qx6+rZNL4g9Dq0r6ntti
kMsPtPX7bHU6CJ+ARALRWnfa1OC5w+TiP4CPfbzaD1XEAQvEJeqlqPQjBCmpBBlXdnzFLgg02MF/
PH4HsFv8st8KantUbUxOaF15DqmfigGsZfnNJppauIgwW1QEFi+u5CYLJnYIFRlhYyc9uZQnuxWh
/5Ywyi1CIVab9Oz09gqC8hPpA0mpqRUhZ0F//Acf0zprqf+I5lY/s2pSXCK2Lwg5a2UQHcA26dLW
oxbIMuO6+Tha6kbbZ8MccpzntYDBlYbyQfGZAkfC9itoAdsnrZ/Ovkl/lSuRKjAfAUgZgZ2odH7m
WLieWtKyRuEqkdYirMWgzyQ2gKgYJOAU403utW6uNwzFeVkWFAYT/LPAzc1mgoGgv44RAyA2hhD0
6rwmnR71RuIqqMzAJg28JtDDrr9A6bDCc4hj87zQH9Kg5YkE3XETcpQeZSrNunQ12JB+6oFMXlt8
Qcy0gKRyy87TDI/ki04u9X+qDgjD9D+6bt/9+oAzX1kx5AYszaKMVajVd7a/92HYYm4PMlsYxzq4
v4u0Hmn3NAZDzU1jt0LIsmb6x9fERRIZtVVHKWMJxck5RuL79pG+d8mK9g+fEP/kCRzTjbfYoaBd
Pi9fDzCj9K1TtrSQITIrxmG+eqOOXjQd4FY02hCpDPHlLaxzH8HT0ND09Ytki+bp5ffUCQLUZMSR
xEjIu6LKVbHtJ2QWLU2On6/beyNEe0TX8VChknK2sI9BqIiLAEsp9HTQHYkTozAcUvYvC3jWwmYK
NMZpk1rwgoOAUsDxzqtCoTOIpA7i37OeuUap/VBvWVoKve84gR5f3OaNvDBrI2ANzG+cde5PO/Qa
Xge80BMifLPA05A4HSTIIRTuuJa7u+krHTfjlKs1LdELolt0aHxPUsox/AZEuSz/dURNdwphYjSz
20bTyPz2ueYaniDiVSB6dGa8/+rB+i0IxX2faE9wHmJIbC+sPMKTg3h8MN88wZWkAKIrxB+08Jdh
ah1hcOmSJ76rRyRSktH+3Ue3xbunV9DlzEaORxwjYDKwWKMat17hX6yEEi6ELVmvAO2emMmil0U6
7lH68qCGQeQxiZK0PgIxl7kWuSKpDq9wxcGWOlP/hnADuJBeG84keyHyvQW2Y6kK1GYKkYiVXgRT
ELYJl4wrSiuGb6g1eqej8z1TaqheTLjfSJ2ZAdjVnIkxp6/fC2ZLJLVK8ky+EPaesae1fpdmyQIO
gAUEdljJ5cQPBKy4zHxpoGNoMPNLVGLLgDK24kOrsWZkjHd8mA5v4ozz/plOt9KJjRoYc8Ua7W7Y
fqEmOErtrnNNIGyi0RMZiyDBtWRXwdy3vMPSx1Q9mJjLdT0n+mQs8zGrSdZqF11hR/x0py1UzjqO
jweQB+6T3283CkpJckTMoxSn4qRqoTFOcfbLejWFW19cwtavP84gTO0Tai9XHf1xKZ8Ns3g9hlDW
epWyqENNNB3SLqI50CZ7xWftmegjEm5jfQMur/rjMdMBHmDSlL5xaQBLcxe+1fzpWdJ97JZJguFN
YGZSKQnCnDocHZ8oXQi751afFJ3Sc/pG8bY0cwAOfjB5NX5b4RYvG9EKhRPhBxjQyTiTChdB91il
mzVHL8EWKfX/O1vNhUMbIGxdDmG3i/ymbXgdMjr2lHnw4X/uXl8/FpRR3QsK2Fmm5QfRip8AFCyW
gBctpcd4opUnh4AXdIvjjS5MV0mfSTbdg5dmqQ5ax51YjVUvg2AHhXqVMSx8z5w1rT2qx7N1Qqf5
cquTfQoJlpXcDfRMs4Frf7b2Z99MAOQzJ89TTQap+GuazvolyWAemdybJmoEOmIUBn0NnGen26bk
ROckE3BU5itXnaGrrXkj0MCmlTUmQPxPh0kTPOLhyd2CSCukDLKLeNBgz3YaQ8QpyJjYq0Wz/C/f
vLfNcMRKBS83l0HjN4tBnLCgl4LxmE2vkClgdL65zd5yUG/3kqg7UNQXjSxr155d37rJngoZDnz+
0xt+UUCmFOr+0AjllYJJ9F0+RrA1FJ/1BMLX1F7G6bsOSGi+KVwKpS+boLd0ziKi84S3RPINQkn0
SDInzlh73ZmzwCzVoi40GKVVF7Osj0kS6sV0YPzxO/B047d5KWaf/cXxkLK8XoBNs7jcl0ncnQE0
jviYwvBUWqHAspgbjNseC9sifeMdAI8BKs2Shs7r5jpQhNQ4Yes7Hugh/17ZvllFmM9l4KjU+36M
urGSZMxpgxURg12vEwCYDMrOFw5OJS/VA3EjoOR9DC0+1On478H73o5P/zDJQzIabResdhf0ooLu
OV7pB28YKcwKUKYewHg5jBu8ee6MIpDgpX08PkpeDDCshkVLw/DvdFgZsy6HlzD8oMF3aK5Md4uq
XoP5b61SazDsEzgr+sSIVnvTAWFz8Hs8E32UriLTXDC6hRxKlM0u5eFLizLshuLXpPX2PW5RFHZc
mB9sZ+nJTDb/BPCT+siYpVI6uKLbNl0baYcPpok2Ax9PDJa+Y9pDdkblsBe6GJ7yu3O+vpW8GH0R
t4sBoQIikG7dGfdB20HP1EtlHF61NREzwt4K7qCiuki2W20PDJE0AvtDALqczgYSR2Oe7G4LCILp
d6XZKHRlR/goInPtT62BVyxqQwhFMbfbc7tuBcSUwEmrwIVjmCRMYRp2BaSfG2Fjr9slRJ9n74QR
ANKpTfOJtx7WmWV0ykvAQkTkkIFeRw/zZa2DiPjtq757yLIaYnSs8335peBEuE9ujzQ2ILB9s/+q
WK2Sg7LjpYRj8MunnpWYuGMCktE7vEhWFG78lzTkiE4mHcoc5HCdKC+Bt7CMviqAu2MPWsa8sG0z
8jGTkMMRc/kxl8ERxAgJ5Akd0T6zgGRmjHydcDA7AkwHt2AyGESGo7FACWvieMHFboTSeFl/5VgW
PLMJB4NQo7oNU6zwq+6gQvFNYHJRrK6UcNYmv7sj9K5UvGOPfUdbCl7VzPrMYLjKUJUw6hopU2r7
rxaSleVkLcgt5ZJyWEmsx2yx3QqTnjJpu7ngHZUc8s6f9uhzZkRAOlQvG8maY8RhkmAKT1sZ0KD0
b3QaDs4+FXvtHjQLC/wUPAlpKX8JiNEEkkHlZdHzxgV6qnQXSALEYDGG7lqeU51LMuEMZql48FtD
UbCTikyHQX75kpuWmgKDWeYqAWADKoLVeWNBX+fi/VtIw2qKFfbOgcIVeKYbY24yoRleGrHgG10/
6rEy4e7TsLzaCK4dMgJebfJ+G78fISFSL4r5ccGJRv5tNWE9fBx20t4CKOf9J7js8PmgxURWelbi
ya1AEGKBo1cDePKl1x3cR/pgBcwyiD0cxqPxeCeIkMJHE3A//tGo5sjM6g/s/YJyXNwAGQ5s1AP2
/Uwnilj9ls5jiZWiv6EMDm3AdkOzvnj0FR0TkhHIV4ZPZD6SxYvRag05WrkzhEA0x1p0VVdkHYVK
qfhCicq3447iZ2OUoke4kqfp/33fS+8lEQvsCb6bc/BuHO72ZkRm1HJNq1L2ikwZ53KXeKyq0H8C
happGgoACA0n3XnopwWPKQVmy+zYQnI32zXRxi9hME8sJZJfP0HlDuxw5ECn8MtYmo3TXs00jq7F
AypSlhwlmo90cH7zdfofEtjwyMqr12pX8ARcszO5dqhk8zciOvGscWiYntLvQ+HtcmOW+ZSjag2X
MMrYKlTB1amaj16t0gCZPPd/f9HSR1uk9ZgSmCCEm9CBaNh9/4I8UHR1J/zESqpC4cH1GAyMOQAj
mFVrVqXNAhT7lYN79K/OvUPExpPCw2F//dcReuEkkwPXLRaapH0pPA5qk3yx/Vx5Tsz2bH5POZ98
B3f71H1BWw1P+UF64yctqIoDjJ56H7pwQ+ggBTPYpXkDJs+7wySQ6sfQS7MEn+AzBwO3QnvVvKCS
AP+QvOvWhBKsCNOdRLuVvB7v+1Xf2o60YxEpQxVLxf1DXnStAMyfeVwe0s3StilwyIazQt3o8tF6
u2htS85Gel35UUKlyg31S6QTAcPs7mNkDEjR+2PKzmB2rlTJbISVpqL2o5Us4RdCazPghApTKpvb
kQEq5q91I0DI9r9I4yEhUS5SCpWlwVMXdfKjbkhETPgUp+w0pMtstdX1EJRqjJQ5QVJMWGuunL/v
humiHRF8SHdoE65+admLc754JPibEpyumd8DYb/dD2y777eEhwOKPEYvFJgHQF3Clo2u+w+B8icC
4qOHWAVaq3apLoIHEj7aeBUQjw7wHhdVrv8hgoHUDo47Xxe9QLrt/lFXzhLLtOHQ+05+nXbYXCg6
nRsmh9Vt7YG2nPaYHcVNf26TEP0JfE3XLr39FgZsNTVZFMeIV0MXvocnL/fnUfDt6anfUAnW1JX0
u3J99udRPzsn8Lh+Wuz0X2N5VHfdXvy69y/xHcEZ5YTHfcGlcHgMCj6GgKKYjtcRk6enaNHIWOg7
oHaiOudhZE4N+JityyHYgZDBuU8QRwU3VxLWLSga48YvbmVoEqDHWmM5CE7N1v2UsMZMD6DteIFf
TXUqlJGFtSjIxZtV/EexDMhMvaapEj76uHDl+R0O0OtOHATumH5JxYrxVyjLDkOteYVopt7nHvvd
U1gUyteCt0ZuSlPGltThtU3KJps4x3DZuY8sin2FAEO0rxFZ7p6i7nbgvSiDuseh3svqJlvmhG3l
dL/5JmH25vqy6RyBmCmBI55ZWRNchAei0uknPJ3NV48lbyDYfQDn5VxEKGLtv18905vi0Nw+qbO4
rRYtIUpA2WGySeiHqJMtfwxToD0vNq0h9XVKAd8KymPE8VAgjY1Y2DmpFlk9PnEWCyFAdd7zmQW9
luCi2ZHPBJeQcq+0pSRg6BS5feX9GuGMwCPFHmCEOhZGfIc2x37YNr3+6ER5pnOPqWsfaPyp8MG+
hgMlUKEC9xJH+PqmUKCHf+lAGDNno11ZeR9gwl5mqTL5Sg/5Xjmk+KkdT1ar1FjcmJ1fsUvthjSc
qgtzQw4GmGpipt8aKkZ1vEbIiQY9xDw01mNLvMauWy8/odNt7/vPKDHr2gH08k2krfwDXVNX/Ag2
c1XHtYnSls0zlyWNVWNdQxeNZqNNQBdDprZbPuRK70vF10z3eT8WB0hPEt0v4mw7KDDXDuJZVUWM
WoPxE5mCnQ+5gZh+ui1pfidtz4L9VMZrR1gje+uvMSzH4hXRghVFG7LQFgoCPIqerqlnDiheFXYn
cxf2CrvrkNmfprNH+VpRJ/CoJUDb+trES4vsbXvlO7scYAcjn7r82RPNAIdO0n92TTryi01967OB
l9Ja0a0q9sl9ntHiNgwAN2ntn9pvAbTeWh2aYq4C/UoHPtQj6mS/5fIRXUdS6jg7/g+xOz84atyQ
mIFNbqxn0VbkamcTfGD5B/UcSNUYASkuTe16mIl4KMNUZfmYTDgCO32mnw5VX3YxK99zo1T4C71/
8BEQDVyqfjM6BREu51Pc8/GDmCJnxbRMOIUwMrsGfKEO0sAm/j48RzlzDoMGa2lfQ+CMFWD4Fk7U
RFWcILH82XTdn5buDd9TsNYXFHwFAoquKyB4j3Lbnag7fa7LHn5bJ6X+fCIV2cZ2EGx0TjFlaubG
cUqHUBkZsjfSRYVZB/63e1IdekjwrEIYvxQr9jHIaS9vYXPRN1I8tTfzCbSKGfx/4sUtSj2gOiAh
8MJRQhA8eureVf+pdDtxnCRkEEK4O7fBBHEdQsqHE26OvEILq4ogN3b1UQibz4OZpw4c35BWsf9T
72a4b0MLm1lVlvE7nzPZm2Kq5p2QB7u31vzEN/7zenYLlSShcC/s0C3mb7n84343Uj4Yw3hQCdZU
SPX0ptqw5bGVpGu2cpN4x3wyTBpoX5j6uxSibiQm72EMvcEegVSOTxTcmtz3FEbsYwk5ws1Df+pB
T8yQWVz+nM4MSVbvmDH/fF06BBDLOTGsVcCS3N/Ix+ZVbkFobSqKwoD1sfJw5ucRKHZqBWt7fUCR
AXERRJzVje1F/DsV0b+XbQ3iAbkWbD4VXfROoL18BZrOtm7HkBQG3jfwrCfdYxh4LlgdiwbZkNt0
7QOhe4V0RyYXPsTchfxaI4O9g/mZvOsSl4czXv5QPk35HZ3GpBQyAkuUA+M/0BQ7tAxW7p7UroCa
hazU0LVJa+Il7e+6GmOo96hc5soa+Cq0l+Z1FJTa55qpwr1WcnR1U04DYD2ufycwzu/Tw/tkmtje
a2z/IkcAwEoh49uQHmZbSd1meJFG3BCYwfodWE++4wYIyVZxglqSuo+qxzEdY6WaFhu9Zn/ZFOUO
R7L3HCuIr3J2gV1HocvGNLZdSDl323kT6EoIpyB9fU5wrHvR+fDnxaauXIFlDFK4/Un4XZKgP68a
qL33ukDkRFTpBqTas+MKV2tWqCsGQmyipC1Ak9C+pyS1bOWMcZZGGT6TEodUX8eRhFBuhOquCVY5
+I8rjuCxAFzNgL60BLQuMD+NqC2jSggf9AinUTOfXIisX1Hy7eIPUBgC2pwdleUEfEe16bgkD0fi
soQnU5UZ1lThZXdnXMJMTRijmnOgMiTYmZ5RUXGGyFtvFPJnZiZV6mcLH63JIRY0qQqypw+swwvt
FPj3cP0JFOkSMGaE+WaNBUq3nkbRSeSDFHOzKwkZufRLsg5QHDnxWjOsd6hMXFZ5eUPnFH1NsG72
O88usWwH/D/5rpq9fZ/7eGhP9bkYTp4Y2miSS7z0hR8hVPM5iSLf3dbHEoZL374k4B6l/jvE4DUX
esE93pgGmYV3Gx6Qxa3UgcWjdZ60jf3QACgBGkl4Kjo/uWnIO/eFLbEciP273b7zmtJ89sUNveq+
JXgN7dteORMRBrVlqh8rQRwyGTHTqHRrP+RRqvHbOjilA0aXgWl83FXJzceabR3e10fJi/H0Z1gJ
Dl4pxFuUwH0Gn9BvVBtOCaFkBdk32CfVNFnl658N7Ign90O4bls6JANiEPNVluscPxyHaVBf+o88
D5oVNEFXDcSI/Z/n5k6nXxVBZ/JIbpT7CU3NGJLAOHer/EvSW16MyvgA30sInMDSCh2ScrAwC3WT
MGc1TdPtoZLGNACIUhsH0bBdyvXWUe4NQij35RqSU33lP3OibFYX/oDas9x4IqKJXTWp9bhO//5g
+DwyKWSkyMHyaqD80IxiPh/GTXzbRgs1OeiBYqjk7SxgHZ0qh96si8w4Zdwf9B3VI1tVX8fwP6gs
fT6FDLwVgwZi7uzUuLhUDEfZUGFY+SGDgjvo8gBalzqLvZoGsL6pMXsgU9vCgt527xgHC3vj6Q7G
dhJJhTqIu9gRLJaEQo7Z4Hdgwzcw38vHmCwZ4zr3RTMxlPMyTq02z2INj1opYhQrwGKT2EXBEs9g
0WbLMbIkxXcxiK/ng/kbCzf3aqg7IHx24dIOA1bzGr7UqC2XigKcuLPaEuDDTE1b0TXi/zdS+v+x
0YSfPgOmgvbNVMN3htoOIUfJlMk8WEiQ/gaQBBgL9z/HxXRqmgqbio95yOp61r4q2qAnRoX6QsHF
YH5sb7IzJw/lDnMu0q0D00VFe661Ju7hIWzXKgRVqnpCGZB47vowMeqei3DujODbJqWZ1cynwOoB
95AnrUeRduc5hgqw6jYd7usfMv1WGm9dvA1Pz0J+uicKddrMXYUjsnZjjBc4MvqXqy2We1pi0Vtv
QLD44GSIaK0L1pNyzUzjpBpliseyt3+PBnXAcLTE9CwuE+oTfi5JeZnB1wMXtUETps07mjknUIEj
eDIWnKCgkEBagLkk1F0zvDs+d2FWk4p9l3bpDHq0ipUwODhbqC53R/UoWgot6KBramF/FlkrH4Ml
7F0rsp2qoyWeYBrBxoc64JKX/pStLKhg2ALnjHMzEWAHSaYDyFblNZF43oFlzRyPlLQS9SYwvdJ5
ARu1lqUqNezB3xfToAsA58z4Go0mM7VzpuzG4Oq3xjxQ6sMoDiBxsHavRjTT3X+pJzc+RZaaDcmt
Go2dMY6yHmr0RsIa8AB33Zs/FeCwhJMFM4ZUBvrw/j9x4ZXPC5eYR/ot9VTmuymy0sqIgwXjikyS
icGHvECR4d5nuNJ1TBWrCkywmh6DLJaEX8gS4mfnVNmvm5QPJ3B0vPIisQ4fWQDteDESgqVw8D9A
vfXwRLQaZciHllg0S4x2ytSbhz8E1osP9mSdJGSBSxVLQLuthNm1Zesnva76P6GcRc+t/1bcSYt7
pW1Z0DXXXpQGrwXobWv1fBX9u493r3ihQRS92R+B1nc/ZJC0navV9KH/gamAYkuGhMuO+KUgm9tO
rX2GaKo9iHEVT2IJF8g98IG86ai/WB8ToBCFLaAgGlJhNb8kYs+ytObkWUaqTkgbHMyjZKXVkLiN
rhp7vdsKaiEnfgzQHGJ8G2ZL0LBPrc635RWwla/3dEkF9G1qugdNXZ6Y+2GAFH6HJxGmA4PlgGSY
3Yld7ml589/alc+mGC4RePwvEHHPf/ryFxI36G9h4VQZl8UMy2GM1Q2clCcv7P3/3DzooF3nEYys
Lmicf7IzLVy9CF4PDXPk1R8cjn1yD32zin+fjOtihxG+38PrAI8W/PWFB7TxlpNPQevdQs7hpSrh
KrnE/bfCEyOb8bB8G3E8W9lNf8wee4LW2d6azygbBzbXI6njyHV1ntuQqrz5zRMRm1xKOKYP22fa
2tAtGMimHVjma8KFSqKg8+Nmkam/045CGplKyOsDsaLMgRNXN6Uno0QgtZZm43UXYdjyFR1UOxVT
vA+MhUjvJef1AUxQa8F9Ji/UesphJuCsn68vG/WgfkQQJIIXX+aIjcSRaxqK+Z9cS6I4EiVYsaua
sVCcwaBqbX3toDqpMWe86yH/v7mNgi74690hBVU35v4+288pvJ40w9SQX9ttL7nmnvEFkN95szsj
t0x/KIQJFeCEK9Gn3Wc7ON1X4k2teYPqWoCdO5jBjyFs9sK9KwPP2ZpkRnkTrDb0Np6+7AI7NcMR
hauHh65HEN1W9kfbid6e65NxRShR1EDeR82pkbsbe2Z3U1Xjl5co2K17Ps5H2aeGYkGTE3bIGUFK
OS4LWRVp54H4vJB2IuEhVtN10qQ16JlT39XJH+msxnGZ+uxvPmqLGof7rqv+aanAlMeWUEwfoERh
s3EU0PQtduFpQU4/TjN9Cz7FzJpnl6NCvwrrKtxzfroDXXSvueIrdH2hswUFjXCcK9+6lMd+UJn1
jqWTBZtflLBMo9bMZr5cALBXcdmb2gruni7y6lY99zTVznlsStwq9CdHbFJGdnwxLyqFwRWBiO7b
Cj8Ga+ruCGP9cKSeFgVSr/SMU8QkSGTSwNhVV4P0Byd1e5I+IX59S6W+0FM3YJXYYIq2oGu58jzC
9xHsgUGN5nLKTbwKLvhVo0cGatxqo+9iZI3bMoSt2Z7+ZilFgTh7Jp0o4ysvda7qe3m8bJQE63eX
AlvBkzhRBDQm4RT6L9d3jwa4NtfIiTFZZoNJCf+WTTK8sfvQzB/WRHaEIZ1Ul2gS0SnK75ocxquN
1txEMsLBdh+nu6fkc+/WbDimwnBuLZpJuUm0E1PKKPGv/QVZPWmXobNut3mvScDQgaFapsxPo++M
1LSu2U+eickQ8mL+hGXDuzrE4pvQ1kIizwoZHiwGJuAv+kxSQ1STAOGLrCbjZiU7btN3JZM52cgq
1ERB0pJv01XdyyMcO9QFoTUkN0kH+an4xWXVwXoWekIHQa7sG1n9RsCbyPuIOT49r+hjQKx1RxUG
JQ9fjKqmu3QGWFhGWyA/MpUwlSwLlFSFLA3MLe8bfJQymAO8VyiZ0WpREttfm5wOh4At9Pi4EvVl
SlNs0m4oHc4zlkv//cBRSK+9x1frjFh9tnQkM7xoFb5WAAUVORHX2hqs//ZJ+vEv9Etgf//i572Z
sBfh6q3igBQeep02iK5HYJK7xoYmbYHDxBY+beil547PTmuPZh7j4CnkQw7YWL2fSTgJPAZ1if5y
/4m0tVLsBW7RW8L87ewGCZCiAqq76tb4repWinv/P8CfUmLQPSof1xUYWVgizoyKF3VAtL2AKVLT
9wm0eSt/nvlodIppfEb8QY/2A1X2/IOXZcI51tu7wgBZ0vDxGI6G0+3QLo8zZOfpHemUFhaEL50b
RZp4pnLx9wXVTuKKlJ0BeWsu+n3+oM7S7x2nm1jlOqBLOzvfMXju0o1YJm/UvwMQOSd9FR5Z3Y9z
3s3Xu7kx7BTMF6vV1JHP8E8fkn4ot5v03nJjpeblor162tJYn72MLo1jLJQmB9uS2Cdt4OH5lxfs
UGTGjrGRM6gyGbtFe2GB/T1jlWVPAZubKgu1vLpt4GGiqXoq3ciHz+r47rF7r2bRYBVRTea93WcN
B9F3+6MFyeYclU0zVuaM51PFlaN72mLNvxwo73XUAhQgG6+KxRNvpGAnReZGPpfFJ4VSHJAULQao
kaKa7c0ovNa7mKDyZhr2BCijVO6SLBj0Ri7bvZ8UDlemKGxTwZ+xxJvd6qtij4MeB/tToNAc5cA1
/xnBbKziyESUtUDUKnFJ4E69wIQ6M0f7y1AJT23SCOtfWOjkLgivAQtoVfMDZ8Wtf97As/2pv2tm
yjooUGfH8YRE2AUO+b36g/uMlO8wtJeHkf4g3P5a2boCyq07NLLAMzPvUpHiFqSQBOG5ibV1uFxU
rF5gvGT/IZH9pNIu0aDi/xEWxj/HDPzmGql1cMaDdnKIYSrcnugtpgr7sg5Fuqyo3SkqXYj1ptrw
gxZVunQtoHYtVQZDH4mhJfb0w3eNIIlxy4ePtznvny72+Be9X+UYjkUSrKUjHqSOPbnZv3IFaBJO
fpoGMG9Hx9PV4e+oJNk/5whde9BPZDNsI+aLqyOxJzycsRwYQzfN0QBx1t8WW8H/q+moYuUj4X5h
yYPZ72VuYPpVZIAdq5NVFRUb3KTpuStXfKovCTRKK00fNbbPf3oN4zIep7gt1IdeTBERgFXAUkri
pngcFPRM+NGDpnXffT+jAc8jDCIn1X7/tr5pX74hfEPjBBpOF4bZ1d0zQ1AK/6yfOr3OaDh4h9dk
0pE9Axhq0Cl2kPYOEIoPqmVP2h2HEEwnfhyHcYRzrC2RTwIqE/pcdzV7ref2/TpLclyl79LcxH7W
3xVwZNZFP+ptTy/aI225G+2U2AJWLblUIC97OtoErVuQS5flj11wnrOO7XhMqD2nna6mQlSmT/As
ShRi1ZcUB9ir5HInyyju9ITzewx2YZfpDTbwOdy6sYdhe7prjPTMRMAvyAjA6dQ0vxwR+rgLVCta
NEmb4KNCiWIyv8C6mrviWV/W+OwH4hd92T7bvMNOJf1IuxILOnVPIOSRcmBXJ9mE2bweAtZPM5KJ
0daTEJARbo2vAmuy3ohATWkp7dLn6vPnE62XdbktTbIMpp6WXY4cq9am8igzw5C5fzVbiFLuYbJ+
52aXEFjvXP9G16u4ym4e3FG6asA+1H0NbEGM98JsDaKGX7nw+gKUukR7o68cvEAhff0bjLW8Ccht
t3h7zLf/nOP0ymohSNuYAy5Mcnv1hX4gvjlkHGyPAjfaepsTWEK7sOyDtOkegcmGETQskoblbzsz
DxscuYHlkzY1qaVuBa/eZAWF/oTg/ImGOJHzhOZxjBF6MXPbxc7L+ZJZLfY8eOYBF6e8F4MMPbXV
LLsdhQL1nFtIhYNjlGT0GoNnCMS0yEwM4Ir/lfSA0WLnRiPv/iv5hpyiEh9+OtRMpfmYd3Ez1Job
yDqNkqFEkbj4AnkfrOMx50ogL8yq/eZCuuUh3CjWC+OI34TaN81mHDxaLlpv1hCEolzMwKRBqpxl
cddRXvaKHy1VTwpJARKvNvA71atocJH9yPSawUubaBD3BZZOl/OIG+Cy/x3J/AXzHWEo/AXqsxhy
Ct2WAA/f78m1AEWC6GaCihjY8mr0AfmN7YUW6vhsq5fx8yiDcA5kozhBhkW6O7HJbOI/9HAXtpWe
//4iROSrV22BZP7/F//ASHHKr6Lm2womoVdLHoayYR0SCRBsIfLsNSdQooi+ro9MB5d31xWwZqCy
Zcizx1MHCmOAzEqTQHQKLvmESekyRsVYrx/8vDZJ2KQUUppZiezm5XG5B5ntzM3hdmh29XOZKutN
EAkZ2W/w60tqLSholpVNlx7GH9HXtAAKsnmOS+7jopUnUHBYj+GEXFRaqMqJpiEXUw45KgiE1PW2
byzHdkWVy4i3Hl5w82UKDwKUiT3VmN6oqTXBS1VWQhrgRwyyXo47zBsYEliljkvWCwDl7oPe/lXY
7m2TdXSys7Alng1VlmYSHkfsSmf/ZXJmLC9+g+NBi+e/VzyF6G8Ql8db/Ojn3QdSfifuEdRK/tVt
LZ5R7+MF8+gHjK5CpCpfKSyXPKZJJ6WSFVZ4uNOU9/ldhv5gv9RlokHFtWIcr+sXwdKGdNSoiHJf
xy165TP1UWlmkvzbxm+3p1rD+p64687bHABZyTqA9cK/qNwih3PpeYXGKKv0e//ir1yHX8sioZEb
Tmue/vAvOZtHmYYRj4G5/jC0XsAXVFwvClVTl3WIGUkAf+xQNx7K2wF/S7phoyd1J/1ekJxG2+gl
0BFz41PK9vP5fCLnTgKRAfRdUARv4rsXzIYiMyyLpKJKZH/IwautuMAQmF2PniB8UplZC6LOZjcG
TOYnXypp/ClRJCjUJZXIVWJv5gunlsHX2eWZpGHaNo29yL820iEPrune6gn6Hnm84hHZUgZQr6ze
Is1xI+/5ULmCXUcmXG/gYp39dr3/ZI8V8BrIuNQqYW62hRHf6wEtx6gg+j2UYnPUe4dp7In1Y8o2
Qg1jjGNt3ElBCvqkCwX/9qqaEpRGrbDliuPPgH0sFm4UhqwBeudAT2zBitdT98ea08P4BiU6Saur
XIwRlzzaeYaTtYNh+rQ6vIktB8nRebk37ZlNCLEPDwj9G7/c/BrDZMKto3OAmkyxtUOGfGjvRtIN
Qm6R5LVfUw9NxuY7QriiAeU7pjkGJiQRAGV6xQA6xMmk5vHFfh+alQgMSPcH1pXKIliTdtsQ745P
dOBjAMkpnleGsyUWYKhN320KSrTfO0dw5BWoCfGc81+5tHgptKpP0r6PGhHJSzB+3Vow0CLnKTrS
vZfVaBDaYSmJa7yfHF6Kiwhvs2NjvU/jvXNMdWzE2xbZtjSAQkMszjAHSa60GFgDZEgCfwAFjgPi
WvYm7WjdslgkDg/yx4j52927zt8OcFkR5YSS9LZWbqN1icUlnZBOIhCfOHCs1UNd3fNjUkIvBrLi
1qfNQ3AFp33T/8V0Xpns+ITT9Zxe6gsR6Pt5rzPlqKWWjHMF4dBtkSKdErAr1R/PjWlr2LouAYS/
19bPcAFbO8V9A1qAKPOFpD2pGY11bIKpVx7rPFtKOiTkr5mrTgJVGPoJLx9KXh6Kw2Papf67ajGu
XVLNadCkGpGbQnLZGfYbjtiOQ51sl8rxtmOwqD53p2f4R9WXu7Z3tyqeOv/YjabrjoxamOVcIeor
1n4LAt98oWVOfDON7Yos6IpZam2cOx+ocwb89gBHpPMQoCpi6Fbpv9rVZS1T/W+gsFstxriXcG54
lnqM6mslDf52v5OXfRdLRnkvagzhqJaDbue6tfFWGwOCmAO7IXcQOAjGck5CJWHCQjJkJyO2FOWt
w4ejVoMXvuAcT7TlCWQ38cRCl7d+paGzqhluLIz2J5ThSC77rdTXIpHReSyX6MdJn+iePWB7Yy0F
T78XNkx8Z+e24jbPSpvA9heBbqznzKV/L1zJnM82UTGLGG5zg8a701N3w7iTqm1PTNtS8uosMtW9
WTkFhCwb/ezUehaoT303HY+c6Q7DLyJ+iZ4n8Emei+feZalbwb/bVbKCYGSQj2nvMQEn/qESc/pk
RkBQjedFmMVkyiwjKWpeUY30408F0GDGUFWz8sXVVj/fZEG8cHsNkA1rwFOATKelBwLVcA0QitoS
qerm+GIyosAmRgACh4ybxSKsCs9dfFM4kNOqzWezZTn5YrzhVKmXYomU/wbR9sBL3LsDekclvqzj
W21R4zTTCXm8X1UBRs0dJodN0BC+4jX2VnaAopvWCEjZmpDnpeM4uQX2tqFrk0FnE+jYd873oNjb
tW0kFKzKC027vWQtI2vsSwxWObBc27UBG89VlHFKh0mRKmyYPYJ3aTbtiwFmEPt1tzwkkGjQFnOu
8tEXwGB/61Jqz8CVzPwXs7redKbd7PbpGO/86e8HjZMCxChfdBmCL3ofgKEV0tLPXUAD9w8dGKmt
ql7sgVmR9urV9aI+gTJ59MFfeil3BBoIiSCuWoryQAQcfPBsbSEBzy1BsPYirC22jP1g9cwDHJ5V
IZx5h0TZg0hV1z+KONj91SH6P0wAxAkJBQoK7FjokVVqVAcUUbf81vb/qsmOBxYndlSjotMBwzFv
c9PPvi2NdR7cZZ3fXDHsMLoRVc34hmpjsexGnYjU0EXNjteDqZGIcNqVCSim2dkMsP7vn+zbQWCd
Ji+reCnJ9RS6d9xXMr/cDzOoXmCCbZ1e8/8LW/y6cOzX60C1cntUNObHXPDMDCe/7PJOp0uxT+Lv
HNvoVVv3cqrwa+ngXHo8cUVdX2qPMOV/mbKexVzgcDQ5bfWmYfYrfXJbSFzxZjihN1fotOj4EaU3
Ti3/7Jsg4Ij9xVQv1CVPJewK1y/6aZYUGlgwusorXl8hnrevuRaySeDuWjtX8uJU7PdTBRdvI3gv
AdCREQzzGQ1ZZHQqvN4ylSD/BQrZ465Xrekiw05C+v/GynP+KG7nxNyi13MXZr3tc/gTtnp+fqgK
qVMWGtTLBC9RfpRUeBmE5TLexwcEk07fvLb81l44o/E3nO/Y2ccQ+rCXUhlp3IQQBg3LYgkDUlPw
GF5PmxkxaVrujHkak+ZiogQUqw9gG8EDOLEOl64LDKU6UV9JPPl4l4uVSy4Vko+RTT57Rs5hXaqz
LIs0cstQlJBHaVZrbF4sjG0pMNsCbA10gGsLHwgK4H3X25KKq/Kt1worz34r9Ynj+ByXxAYMVcC7
tFGmElShZRuevNkWM1NkZBuzUjnpl1yy+z3Ac9AC26mIAOC9zMbV+ke+bbFrKofzcHx+8dn36JeT
CY4OJ90Kz/zmEBhSBS3wxgJR8figO4j4vXC1XnGj3p80jYON38pYpdGbTLpTP+Pdxs8Nb+3CmCKP
l/pgcns9BDlb8fyWqTF0Wulqde5viwfo1g2NB4Uas3StsirD0Oj2kbvMgIrXoAz17DUkmOfD/HEy
gJ+MB1gzyye5r0zcjNZ707ChHxgt1rR7A93HXJtVtuQwtDxKht/fK+DKl2NcJqo3YyH7ovOz9MoQ
xBtuh2jw4lDtrdcF8hb9gksNts6hfutGspNXAvLLKoL5TSgwI8BzNGeBsDJ0xJfckyGXFDIJ6s5x
B/PdVMZuy2XMdKkciNiDj1XWWWU6Q37R3zSZlLrrqReDPfIvCr/ySEo9Ixk2CvOVWO+snH+MglL5
Or+Yhqs8Kd3d4UzTOSw64L0qVcX50OWqRxjY9iHC9YwsHUUUxlXM8+0NHax83+FATjIcee4CEIk6
ygToVSfD0KSivVjz1nPNdfaP0ps89c7Vig0uSwEQdF//8ws0csgwlw8jg55c1kVAYWyVAtLoBGZ2
p2R6fZ3HkF0pGwufuG7kHPu0lhvbDAjECrd62i2XMYO19po589naC6A/trije+ar3l/KmuqhINVp
Kh7Rkttvc3mpVWjySkloyT/T4M4RbNkDnHN3JHxbKi9/JHh0+jhTxFT1zhFdlAKCbDcAGWIhVYyk
9KzJKR8j2Rkf8sKH797bWSjzRTcVYhupNd6NNKWDbo8vZkX9laRJxAH2qyEDFbZXYVR4zwLChPZx
Gj/pkWt30zNxMUlVuT/OFZsPn6HHvXBLpZT00XQMTz8esRaRqcRjam474NK3ffP35cBYSOSpdlFf
Te4/lmvkxZhZkgH9fIFaBwXhPPumjd65kpg3xz/WFcxlfsMTn+1FIjsu5Gz6Oy1m60kbfMB1fyC5
PZlGL6dts1OLwXPxKys9R/pipIdZ1fNk4KE3x+uTLmqmcJGHeDat9DWL5+ZfjqGYSrz+RrbX4kfC
YmaCiEu6wRpUZ7aezpoP24KLLNryjbV3+Mo6/8HMZnw/wyJhwl/jc3ZkcQWJzVk3dQvGZQi+vwxY
7Nq3S2gM/8veECJ/J0inaiQNrtubfwlck+CdTeGb3sZNdWBaSDbZfH8mJFyDiByvVQDzsmiBoe87
hzUXz2KuIRgaw06UTyyH11aJwgleSI2Fi57Z5G7AksyNnPmZpOQH3fqaNsAMrX/x5rRPQUpSg2Z4
gfzzrbH7xa1TJMrh2sTs7L1pT43Oued8hM9oAGGyhjBdaILnEq3d7yE7n1d+d3JeA6ign+SdiIJj
gsmqgQsF9+chRhNOyqFQ29jQnnOe7fiMNgP1qdP65dEAIt593tUVYzgLg+1So+JNgMDwZeLyjGRj
5fbpq9A99qu8YcQkMRzoro04IN861oyyz2nZQgE9ymVEWDSxkZLyoIShMksA7UXxvdcAVhY7j8lh
Ejgk+qQY/BvsPWZLbMSPrfoiGw6cZC+fV+UxUoa3u5gkegzVA1zweOtyt9c5Gne/YHnvG7kBCDRe
gFmag7Xc+clqqLtlLazCyDIY+zJ9qkCivW7SfKPrTdL11vo37QM96NyVy4bnSRUXy6rCwo9v64NK
HnQw92MBNj4lTwy4fB9sdW5FqlA4DyPMSJdXCMafhLGxyq/2k5fNUXRb0W0GzHHm53z1gXjhCU8s
pgiN2Gw29p1YtQUO6i9Qu4DDLOfvsIcmnH0wpvDm/LVDgHiGOUjntJpUn1HwcX7nR4K2hCK2x6yN
TUO7v84KAFjao0J3+IwRkevImcgiMZS15AdIAoHc5PLXxEYaaWRBhro3Ug2z2x5Gu+Kyy/1AiiL8
5Qk52Sxrra6fIbUe+Sd0O+9GMXunJGZ1ohZsDnWw0lyeDrhLdgeV/6EwH9txgmjZY1GrONWDm/WJ
JyySN08pr/ubGQBInHcC24V1skxLoqEKHucPsy+M+yi25sNzB2QrHuq1iLMZ/2Yt8fV8UvWdFcnL
XFtoQh8/0mX3rL7IKGXqkD9bhBfHeQvGqMU6BuXQfKNQAMKyHAM1Zv+6bT8PPhCgn+1zxKYPsZcG
FUXQNWvLO4xzo546cnnH9oZ+QzqzAt5F8cLsUbLNdDwtizkuqrUxEE8KPdTCM6kuo++pQPzb6EuQ
2foFutm25uPiEGxavDI6Z1Im0giw5PBkmPX0FjZvxJ+MU/9vyaXEqDd1Kr88g8loB4omoQNP4753
vDri7oQZNFah1SH7GnEQMDBGX/7XV+a0RXO1X6xnQS7ZDOyXGplzsWOoA9GSvzpGeCgPeQeducd3
lqMHb5zwI0+TLP30KK4IkamNzGDEjQiPNQ7nVSi4K9bVj0sLOvMCzuRAUmWNSlnc+YxOwoPNX+JF
azG7Cc2eLR91dMLZqK6QACFSJljPV9NJljIdt0S6MveY/vfNC2IfLzvX2culmHuOewYRI13VIV7r
pIm4lRUIbAgrSK4KDN7V2XsM0X5xKAWfbnPx58j6v358mPMtOSDVXbvQAa/zT9roKE1se42dlxAN
byDh/iKPLoF5Fr5kbHmKqAkWs9PaWnB5F8F3Z64zOwcxbx3bJDLSJyb98CwvjDtyZ+fPQHpGKUK3
mtl9OsaOi7I6N14YrCZ59oPK4gRHG4o2N84HbIBnUzeAmjE1KXoDngGE5uetCnIkOvRrSlxhLBRb
ajC8U2NTaVVVaCdspzoEamncAYnDYCP9y+haN5z4szuFF9cZ2yKwUaJre1nag2M9XVbEtJk0/OUm
2Df7Yjg3t8eQ7DCtHx03oFMD9UP3idLBKaAu4kmPny57xX2ej7+Hw15Ja4ciqH3Dgw4JRCN98ZEB
DkIXtSgNbNFxxAq4OWynzWbLQtQsjfipjI4+5HIm/jqXQO9Pke40gK5RMfJAT5Bno4KqM2Rz5pJf
xqKMs+WjbZvztDowN9c2A61SiClm2s5mFCHfn759MALmp/vNXFwO1mJ4HIdY2vrXm/ErtARvrgSp
PU6NICK+g4CtOdcZr21Rkh6fVVBu0wSPXBUWPw1xS5aC4QtPgFVwUs1d6z41E5nQkp7lt9/x3tQg
g0092W0DPf1qdXJ/6+OHtQWI27N9NaXDWrAJYpGENIK9Si4TlSdyd+V8JedsxS0TUN3F60p7G42t
SP93NRJ+ZPD30AcoOdYLfC04WVl01u3U3ZKMDYbLL6yDZv6Gautt2vUDQASv2wzwGD6QkFtbNC8F
XUakcA2/U90mTpGtJt0emgdGEZMPjrMuSnPhvA6Ipx2YScUW8FfHpbfJBUGU9QllkNtmV31S/AZM
ZN6Veffh6LJcdGnRT0bPbRruXYJhAOWRyfXFmr1NHClv3kF6CcbMvauPMXGe4mLaNmICsniQoUOJ
JAC4UBRS0HY20+ToZD7ZXP8dmjb4/cj1DWSjtPaa11oupVsK4wHtL+rdnStv/EKoZFj4Pu5skwH9
a8cOJys3ghucpBows0pYNprZ6Ru6FvaYqQ/4YyHWmXB09ouft4sR5VOpISHXkDkrvhLaI344ZP8Y
E0mM2yWO5AQS6kZANGhg1UwIKYayYFbkSFwDylSBa8A+xulub3zc5GASj7cqvKA8/W07uB+61xRx
4tNZYVg4pT49zj0OC2KnB+tO8mocmQ5FP6ZwqKurMlLtBgrJPAzN8iYybsY6TJJsViiT5SqJsVE9
PlQ1uesFQUubFS/k7N03PAwdCrRHp8DgQ5E82gax2ozFxeWtKU29lij72CWfjMJye0lm1REqwj9b
9hn6inX09zQxYLbv/gi0R4KTrdfznvNEXBHBWVZyghIftF7Xud8wlpsDtnD1aiIv6l+UHiBuTKLF
wPNe87oGQSvo46O5GsH/njSongOmduMSv7AAgcKWmdOPDQqN0nl78aJEIuSzRJ0uJ4sDeAutAT6z
pnAfNmLkRiB1rmb7V3uBKXmZ1FYWRa+cR1Wt6BOQW9nA91o+UHHfmzS9QFgGFIWI1FZ8iahg+Pq7
MEaF84V1susZqaKYvaaVsqmVukDlYB5NFpvmwh6FHd0kZ4eAx1NgMKIH357yhbvX4xTzMw3ZkKEo
Uy6PXeD5wZuBUcyZoutOhyt/XnP6nwSmEUtZRz98p8x4bNn5UlHaceGpaOaSC9fnDuxMeHokNMQT
LCOcKzH7qztJ9DLZtVYmwG3h8qrFYnFeZm3h1jbS82huQf6oZzVrbLjc4aeAcFgQ43K2fZpxySHT
S39mZgLQAXsStaSDP9iYPGG0ta02NBuh7bYErJeRq7Dn7eDkpH+aXKfFhqPTX2C/G9pFSgqfWfXM
DsieX/i9XT0tt7D1YO6KHvhjHbuZQ9uAj05fcfXpY+2xS43w+A8+qzOcJcZY4uALylp6chEJhDA4
7PpE271Q7fTWYSXKvrDh2cIg0I4OjO56l0ty9E2ITIVX0cX5IfzhbEheNUVkj3f//Ztf/uA79GoR
ierYeeU5Ls59ircOtIg6cKfan84qC0DHYo9QEC+4hqCa1REgwjSyL2m0kwb6Rv90EpIxCZY7nacH
tooc+yGJ3/PfEvCmDQcxIIHCBCyxmjr1k8GAPH8JrxeG0yRLu3L26BEHGVyfxN7m6oMOwWdKGKwe
nk/ZOBP36tZTwCbQ4vG8MN1iaVyBoPewH4spIsOWcB45FQazpzJ08HiyQe8gU42q4Hmu3n/Mg5uI
i7idTA4Mpr3k1tAUzqngGHL74LY9sxYdY7dvvLToVGMwFg0p5KZL8KKftcdlEKhjB+apm03Xz8hq
2BysEtLgDY7gilnGT/e38o/dem85gMBZ2IJ0cvsGl9OQdqnTbMv2rTJSD0u0g8mTMEHCe3wHv9ak
oYm86cpb6M1bf+4FLEb6BmGHcAuQo5srkvLqiwwqRnT2kNa1Dqmnrb9DIa5EC1mhGXp9Y7OleTHN
w0qB5iM26m0ESBB5eEmeWOwktDBjPv6J2V2WQ2mfMqZVMgfkQRftrIXMpeszfYR4Ab9luO5L2jvY
tByHc5oqr8mxils3rL+IhH60gP1dOIXkPT1Gj37PfIXFFAq7XYDRTBp70pP5FHyKMznV/oA4gFTT
6AnX6aG0KaXZa1Q/GsrltKOyDkZaQtV7qA1tQs//aHWSUHWPVabj1TXuLtyhlKYFfd9EEgm1AfXz
wtt2iG4VC3FONq0j55jovJ1jUzcojWet+e85FS9kvEpAZgCj8l92xPbB8/AdEqsl2XcORiaZJlIk
RMnAntfWQPtDpcL3Z/hvII4nYbv5+0gl0HlOLiQs1tzJVzfsRIRu2KqcF+1tq7h2xcFglFgqJ3mh
7/MPz3KMLnR4IggeKgCLMoA4dNoUhjFudBNFGZxBx+p1FDPMVHpm8KBcf0ke7jboGi0DJOW30ZFu
HOGS7V96qa2lMhEQceWUjLFRwC+mQs5IQa61UFjXaXk6EPkO92m1OZBU76OKZz8x8xyjhrI8mpPy
aJfp4i7m7dgLGt+LsVN6oPguDIcCWeA/Cm0H0/i9dOaY4HnHMSlKxwuKLfyYjZYbjXTuF4DBzPb9
7ROLh6IHiGPZKprdxLaWd/3kSghM2QFYS2g2l98MdrMLYZE88fbrGyYPrtOKpN2jxmlWJNmAVbns
7LJ1oR3BNGPQOkVBiql1p60aDmfQjVpoDAyZMcumNL923JdR6Fbd42VPb9rGjCm9fmAZ5IYmSobH
bpzbX8729ftxABs4g98WahM0D8NJ+oECsweWn/fAI/3ACipTkNtjWkaI+2txIE5Mr1Umf7x7Y1rO
lSqIOcKPzPxg2Sg9pAxAy/EJ9xMEqc+Vd78XH3lZg7uQ9hIJhcltgEfwOHxpqmcKSv9OqMuxtGBX
iXN6gwPaGknhOLDMxPDkbDf7yJad+HcyZAaPmhPBdnvu1Bjqe5dRrZGhiFTTVsXZAge011TcH/ng
qDWbPMPEunga3/hqpmQM0OaLQtDzBSHojnH3DuH2bU3ZDKLCbVwespw2NG5BeHwfSfQbxLI0KkY+
C5Ab1TDaK6zEioz9hmgwfN/Fg5VJ1tk7QZ/r9bEwkgy+91gM2NKBSqE7FEUqq1wVaygLVw5vvEob
YmY/r8rHD/92hf6L0PmZrYolhUBpyifb7qGLH7F/8pzISDXcNMFKDjmIQWRLvD5W/b8FyTy2vOGS
tXykqIQh/7okuHgjUGWJlSmIR+AA6ceGUnzp0BEkUX0kqTMz/8mhCV3gX9tiuyC4GfX5UXtJxqyS
13ba4U2dmZVlo8aEvwIVAmOEUbl4ZQCiX6tE0RayEqVRDrVBJHP6lbG4VBgds0eHSm9qSq1BEfUz
iRS3qzfo+67x8l4+FP17ypj36pVpKKFry0fB0JEpT/U0yNHiJ9La74US+GK8wxJpCMdGSjFLTfl0
lBsYptOyea0xK8SH9nv23/H3DkkwAef2XI2JOUC6mSPFhJ7yeUOj7VyOxPG8fZxLJh5UotcsflMi
bvb0QnwHEJR2mTNx1Q9yZAoGauGIkFlziFtsHgUilA/DRRSvqBie00KeWanW9ixgk2Nuiwk2vIfD
T12fa+wRf4ISW4fQFNsV/69prSxNpjcv7q4O/RbjVdjtu3X1v44dghcBvasMQjD2Z+Rj900cXa5B
XoafwdD8t0bxVqKwFJnoIhgqtJEsyDmWg6hsNxciLZXNTlzIwppuukQc17IbT2qhD9NqmPf1lILL
6uZMGXhUvrrsUTa1XtxydFA4/oWNUxTpjTXSfUyHj3lWm8ZLzAeXZwoUwzRInDmYiNKBByugrUNy
z2VaKOiTJIW66xT6SBmhWdfuCXY4KvuIuFT/LcDmxPjKbx/KXg1UxsrpBMyeW3C0NvFWlMbP2wZQ
j+bpwQ4Kuoz0wI186HtJ0TRoHd5NaFe5bx7JmduRXNU8kDpnkx14h3ZoIXBvO5xKeo1JRTHHA1rI
Te7Mq7XSdWP1WpaWKhv/O6zqQM3NhTEPeU3vmZjJl3eP9AOp6PQ6YCjdhAjlFIOr1sp/p7zojQWe
fqLD7bwH7MJPCKHYjPJKfiXfgo8oTRZReYZRs8IZp0cTxVhrAg6GSLOTgr0czpw0QX0c/eHC3Rfc
fe+86pGsHTw2XOn5kRY//Pr8pjXSqWliTZcRAmoTG+Axl7P1NdFMJ9GawpZYhJaPRV2zTtyQ9dRa
LWOvmafcMO+reMMnV0r7Hy2rpjXOj2Ibr0Xgwke21Dd3lHd9fB7ynB4KnXnBfQ+OHCTbFMOTgBjq
WP9wmAfmrFU/VrBTBAIjvflQCfy5Y7j1xutvKk8ysPob0/1s13eiza3GiWK3QFPXZanYWi4zkKjs
vfMnwkuQkySHIR7L2cTXmCu5hYitZs7ORnCMpuy+VEFiuqPEAD4hGy4osMyHcENscxCverL3yVen
KDDu3IgEg7ILbN8SaU9Xnsr/oyMLQ/dcq/M3wrN+/FkYvhYTEkyFgToEB3gsuOgesN8qb6iBYzBD
G6fLgm6PVacqOP/amdlhrH2iPo+GfD2RUiuMaTXsyv3jAGakc4BbVcF7W8U/r/dKDa1gVbshZ9xO
NMq29QBgOKKtvVR6oBuQDSaZfwCDHw1y3I7AxxF+kUDXMTyz7nUo5Hmhy4viBxcHi0Kr6Hhfbl6W
yYal+Fq33FSx9YiisIgxaWF+aX5c146nyfBrAri8scE6qknPkrGQrdIzMi14n5G2wRDvUovkiMOR
20GpjLFUgNsqczfGGB+dKRBPyi0YV6N7nN9Ccbm9myOjC3vlIhvQjuj/FpzCdAt5mXXn7DOQijTY
Iu3kTBL2DuG1FFek/IuSfwwAKIwp7p7qgOiZ2S3NKcNLbLJTOw2wM5YOgY2R7JCfmG8tYIeXA2HG
AvIUZ5bpf52oIYBnhNNHF+1Vs/fSbdqC0HHuJ9GX2j7miVWRz+77+ciwTyQV1mFO/a1WGJHu/4b+
tbwRunKo8avYdJ787mfOjuRBG34KUlFtz9UlpA3fkejgqhMFQ8ROXag/78fme9oRkKimGEQOYhuX
jVOviD/V02ntPha9Bsnbqj0TjjfvIAJFng75TIGflMQaRWTfql5Z4huEyltefTxgsccaFXttGuoP
aBbXJ/pTjeeWhYxOmyQkDFS91IJQLZZDHFqH0SkwHNJjV6p0+IuydT5bZnl42eVMoDs0DLvg1Fxr
BkNgwwCYuGARPjH6DUt3zKcTgrxHfulJ9NJXvJUj8FZGpIh7qv3z0jdvpWm7JjYNsAFV00XCWhXG
v+lIJaI/Zea/a60Fi1rBlKX7Ddk5RxJqwfx1RyucOD/kKqW3o4Zm1oRB0hk7yeUoqWtf97Cfm2ov
vWaNma0oSCLb2268q3USOF4Mn2IW5+Ob/gbAkuvqb0bHcB1CBMc7vqNwu9dSdHYniYCS908EtBcI
52wRs65V85GD6EBVls2uaZwNTyIlOIb12FmnNl0AIJHpvdJzU8U8FSQYUBl5gFahi1DrHiitbaAN
gKPxiVbwiAXH0Wxz9p9863uzJw+i4zXKX6SLEnff2wPx8u8zwvecc77ZlGgKM6bto7PUlwWqwFlC
dnBhqz+ZAkiqrpBx+/ds2ELIJLNUe1YImVq3AhIVQwQToNdNbBWQuEceYv5TTjbgRFvyMUOTVEGr
+/PnpDWI3klQqWKWHlurFlfZxdOPuT2lpNU2LzZlz2d91y1LDWDEDsGvzincN6bTlBo3seda+MZg
GIEhxnhXavuol1t6Iw3BMszsRiXj1t5Iwk3+COfCDIaQzHJ6wJjcUxzSq+tUzXDyo2CBqGLXzjrr
MEd8hGnuT+UaOkeBnDDgfUepw1PiA7JX4go0QoajpNAOp5YY185NaE+TV7vuGa0oKR+JtiZ4O0o/
hzGlysHHvWMdf1EyVMOA14oYQSceKyKs+nfhtIxYBn9rPSP56VFQEPDP+F2jHeIhy2k6D44Aqz8y
hXclD4k5bBLyMOWORwnuu4ikloxoHzbfWQIBDmXgM+VZwH9xG09lXqGKVFhXA9GYKHWXzxchYt00
+iQCUNhav4244Sm7pts+H1D9yIMh1dhRWjR46Jw7nVyd7SJyRj4++O3TzNrBqSZYmwd9hsaSwLJf
QDM1kxyqApMkgg5dadqdCQY8iVtS9YJrNXAoHkGHZDncEhHYX5Cffde8/whhUd+l8MnrB92MUywR
APLo3G1708HSSsBZbkAW1sKz53WScjI2fsOu/mA+6Sym/Z+u8+O7I6IBfZ9WaTsUMeSzKOYE3Jzd
WbS8tLObtO5fbwXgZ5unRjcj0lBe4kmfkVBnyQXKyes97vW6Y1mg7LSGBNuD
`protect end_protected
