��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���_$L�s���u��e������7MR
����w��6�]��p���0�_���D支��
/�֍�}��Whf1������H۫ǖ^IY�
<�E�W���wFh�ۧ�0�D/G���b�95�WnB5	����_�������'ׯ�]NF렯��3\ں		uQ�Wqʥ�<� �n�ۭ3�q[�����x��1T�&�o!���Ca�pY�]t�sjH	^m�����T��q�3�+ȋ��g���ۚ`]���)X��d�����P�n�i�O*��l?��*�g	�Ĝ7c�L��|u#d��_����Wb ���j����$w��	�!/ ]h9`�Ox�CG���M����3���Y@�<k'�D��i��XV��q�����8��n���'�85&C��ɣD��?�ֻ�Dg"|iP������I�g���$2��#���p�+�+��_u���Lo�a�IWYqgYs�����+�����Iͥ�ˇB�`5J��?s��a�: z%}�11�A�;�__ ����Z\���ob�pU��w����
;�F~�(~5=��d���5*������nq����e�^����!a�����3��{d�.�X���+@��˘�

G�~ւ�SC��D�h�6�a�O�1��uQ�-�v.��+��t�k/�R�uu�J�d�����1D�gd�s�Z?�����VP*NӥC @������G1S��y��c)bj��&��(߷D��j��@��h���:�Chw�&�x�M\�]�R�Ú����������c_ѹD�1S6���Z��X�������4
�t5rk�.�� ���$-7�Ki��bu���p����Qt_e:/�S�~���б�*��1�|V������fm�י	�X�&-k���F��Ǝ�z`�܆�26�*�ϴn�C�r�������i�W���+9x�v]����,�j^Z��������Foq)��V:rs��n>BM�<�^�,�[����t������|&��Y��Y[EA���8�i��k����<\:P��џ<�%����)U��jn{�07=1�=�x�;�f�Ke[��K�$�1#)�N����}����%���a�vP%SP�J��K�`���u��]�3�3���5.j	�	��"���`\��W���U>!��@��h�%�ɉ٩޾�$��ݍuF����h�l�k��&�N=.�oH�ή`b�en���5�����z2L�Fb���Y��: �e�A�ͺ���p���䦣��or�>���M!o�Yd��B'��W���hgq�g�Cg]$�}i�n$�/a��FoB�_�BS7���Hҿ�UKJ��p�kK,=d��^�>;,e��m��*g��sK����s���_}�^W�x�
����
��c)G!.;M./6�Ex9]�$����\d�sg
��� ^I�W���B�;}F���]񔽘��xJ-wp3�3�V�s�;!����n�K�]�������۴~�yщw������ۡ�t�1�D.���%*ow]�4��wL�e���~́�����v"����eC�>��=*������8�Sa{��!�s WR
�����������G�z�U�օa��[�^%K}2?��&�i�� ҹ��z�.oa*8�2kh� �����愔d��3lM��A�`�[������Q���	D��r�����%h���鮰���S���OIDa5�S�f�4���S|�Ϻ٨B��+����g��C�s�����c�i@\���U��#�Ҥro�א��R�65��HZ����l�M�K��ڕq�7�&L5�J�2����B�W�<\W�]��'�ZVX���GT�
��,��6�'r��_m�{�O˗�ďl�xȒ�|ԑ,��|�;�!�ŝ��#�y�g�:O%nůed�본?�g;ڬ�g�!��Sos�Z�_&����%a���t��.���拓��Dм-�Yڢ�\���B��Rٶ��I��p#s�H!�n6�p�����z�}X��H��	�b�:-����0o��ř<�������:�'����[)�M�(_[��C<�d�;����B\?�ۣvZD?Au,8
0\tC�b�#�l��?�}#�1�fKkXu���H�lA;"GY�;Z��"&�b/�ݤ׷�/�fINv�rE��߅�_YZ��_oc[�ܗ�t�E-~�� �z#�0އre�y��k\�<VHOK,�cg�u�p�T���K8��W��`�%�\�JO�?�<} |�ʋU�_��y4Ǻ�*~7[��wS�Nf!s�:^bv��E���Χ�~�j8jyn���k� �y���C�Y-��Nr����c��J�(Fu!��f`J�,P݄�� ��TƯzp��I'��.]��
��6�Z�:��]|6�.�jI�$���
��I���$6 eB�U-�z�dڨ2g��:X�v[|��!�j Ö�J��$�?c)Ȍe
��j�)�� �_l2���4����M%�y!b~��8���ˌs���[	�F�H�cf���	�+�/�}�`�����b(�"�g��҇oyar'Q&ӹ(>%����N���g�q/�8��	�Sk:�U(���Z�ϱ9��x�A&2zn^d���eH�'��'���h�y�$0v�V8��ca�8�,�, x���ǵ�xh�Cd��a���K}4�|~���>�l=�μ��9�XzGk�aJy�q�%��e�cX1-�b�n�&�<¾�-��D�|#�>̟�|c���>$�(���6���N��a�KNL�61V|�^��_�]�b��A�)��AlG�����˙�1V��P0�"��Hs�`C;/�PR�F�ׯ�F�xpl���m׿�p����,ٟ�R��)̡��LB��#N��4R�*C��l9�N:ӮSξO�gtQk�1��/�o	Cn7o��z��ʢb)M�Cy�e�e��0�U��5�/�/I�߾�a÷[[����� �-�ك�:�-��n����-�~8�yی�.|a�7�� c�V�Uz�����y��T��u.nM�ϊ���|ط��K��g�;¬ȇ��y�բefh�;#$�)���L�xu�n@^�*�l�Ա��Z]�ɪ{��������Y�fD�?M�S3)�oihr!�"juwMͻ;.^�4�Ĉ(�'�ҹ�֖=gV$fĮ'��g�!�ڏ�RW���"�����/[����N^�����T��
��x�Xw�{���L�a�l��)&u���6�u���'H��;�o9�	�9h��r��r��<�|o�
�ď�(8�!n�\M��G3Y_����++
,l��|${��?��r������73/����|@]Y<���5�>�����s��Q��c�����Ct.�|GXG���^O�@��/:Ll���P��0�c�D�~�Hs���K����`z��:;4��"��1��M���6� �~�8{����f�$X(b?.d��Q��=�Sn~[�2�ͪ{w>B��=��4X�@Mx*�����+e�1���`�){�YX�o���ֲ*�O>������^+�x_�!�;��@`�f�)h��IB����ߟ�Q�)醊	y��D¨?��G ��ʤ�\#J�5�Q����e4[D���+�o��D;I@��f�S�6��(�������yH8فu�7�:]ݲ-�CCj�}U����R���˘˝���9�G7g���^0�����_��U�r�]T��
-�:��eb/�WjT1%�q�[�$�-;�k�W;�)��-�1�\"�X{�)ߪ�V�ث�n93Z`ԉ�)���翶t�������u�:����`T��E��%v_�������iE��mpp���| ��GSP���c�D. \�ܑs��b2�nc�#�ڶ���z!"���b	���%�&1t?�eZ�Z��F<�~�}�r���4��)�T�sȌ�)R,���5����·=�OK�I��r���%c�*��� 4"�!�I1(吀�+�_C&�`�����:���mJ�C�e��ƨ�����,��N?�����)����j��i&���K&!e+"�o�̸��u���0��Ҷ��l��Y�����д��^�ӫ)�7C��;eY>��W'W�F%��|+3s��s��ݼK�@4&V�OZ�"��ed�6o�c�D��1C�tѨ���U���eU���ˆ�C��-=�P#C��-����R��!4�it��C�L�% ��6�����^c[�`Z)k���0A+r�rr:�?L�IR�����?�ݯ\�I<���α����]"��d`��EoH?���`��j>lm�.&{~0��%�@�e|Jf���{;4�J:�f�e:��1[|n=y#l���\��55�"�q��f�߲^5Gv�`|�1"�a��=�g[��@J��(����[1$.��g[��A��\<;�H�x�	:p�����
��P&�X%w��UT �J �Ye锈6^���I�U�$�<+#b!l-�2:��������Q��"p��Ei�w��B_�O�uW�0ā�	oH�gI����I�_T�W�L��C����blp%�ש��$�E:�KY��ǧu��Y�,q�6�w����)8msM���.��O���d�ٞ>����eeS 0�S�R�UaT��
kϛy:���a�Bf�Z�ޡ�>�՘�Uu��N��3�Z�Gf&9�Yw?z��'�^�A4I[N���w�a��4�~B]MM�����R�h�-�j�=���DZv�dQ+[��� l�O^M�w�e)a�H���<&[�'�]	N��B�H�Ⱥ�J�J��19���4�LNM���@[J���4F4�T�y�n�JC�
P5���XzU�j������# �%P# m<�٤m�z_���T�Cf,$Q��y�&���6�L�LdpP�Y�!�@mκ�!���[��j>������b �0�m�c���s|���+���^�.z@�uu����{��w�{y����QX��a+��^���O/;��[�ӈX ���?�/�_����+�.�^
�60+Iݰ���p"s��6��.
ƈ���� �*�S����KG�/�.�)�r F2;K �ųZ\'�9�f��
*S�����PF�~��g��B�W
�8�'(�t��E�`��ݔU��PNJ�߈�a�6�y����J^�>%"�4-E�D���ܡV1�@_��S�$�t�'�[���/�b���`�R�iv�2ef��\��R�Y�hP��<�Df]ٗ��(>0�ȄF����6^��Y�l�R	i��%��Η�to?��/�@f
�*c��YK�H�A&z�Ԏ:��(�L�̈޲��u.�$��6\�x�+UG� �Gh��(3���(��w������H��8Rf+p#l�{��{��`kM�{��+f�*V��7�B����_�U�:���p��� ���$�!����]f�����;h8xƞ�im�����e`��[��#$�u9WFF���h��:ӵ��/<���r��fP�6j%�;A���>1.��]���L�J�3k��Z���`hc�8�œ%�Q_|8�20�t�NY�P�zl>�F_��^@i�X��Iϫ-�d�J�t�8����8�Ps�Z)���z�^{����� �֩(	�Ha���M��dR�0b������+�e�hpJN'���vʒ�
�/<�3jg���WJB��)ӰW/&��<�~\E'��|��nU���Fo�O���6�򣟃�*�����' �BSY|��Н�&�|,�/?i�
�!�_-P�O�!��<sY��$[:��V�&���`��ΉTi�R�$4:<���z��T�L�dW�}�+����P�a5qk�%�?f4ي=b��\����}�-�G&�W���n��kMx��=ow}y�<gGVjc`\&r�$�+�#��SL�3cc�@��c6�}���!(%����j�E�v�*�H��bX���y���q�r0x�vU�Y��?𿚗X��z�#	�i����|WD��a'���K�3�!�S�a�j͑/�;�-��e��3t-5��s��&�ھ*$�{�1��h��'�J�Rx����dy��*���z6��c�>U�����o���q�3Ʒx��N�G��AV�{���|B����3@�AB&5j����i����]�<�Ĵ��ȴ�NZ��Pѽ�H��]y�.P9�R���׻�A�9L?������
+�lE��!P�(��5�+f =�_�i�b�_=H���w'�nG��n-LE|)J%�S��i:Z�0���	��0E�Q,iz}#a��2ySݗ>��"��Y\.�sgtci�h@?͓砠S1�E��L�g$��'̗��9FC������jՌ�nä��ħ:z�S����1j�x'���?<]�����#DEF�رɒ�2�7'�=�VޗWCĈ����}v�$��iz�����ݕ��X��{ѯ�A]#$n�%2s��>M�z����iu��o�A7�����~;����]t��'\xY¥)��\
І�há"�&��Ɏ���1����VW=�����;��:ȷ��YRC�<@j[l�t�U�м�Q�O���G4|��Q����F��ӏ�.�IP4=��z����V�����ġk��b�I?��?M�R#�E|(%8a���Ν�1���}5�2z�yRE�
?�hy��ZM�uM���xX X��#3���nF˒Q�e�e9l�V���w�n�KV���ߤv�9�%߿�Ô�xGK9M�(K��w����3���37@$�%�}wo��sx/�n�V%ۅ��Df�ZuR��a}zY��I�ozgR$�.E�L0�D)!5䘿�!�7[���)^4b����$;���c��T��~�0�{�3?�5X��/[���BȘ�]\�'�}�Hdvg_�<�WO�֊��99+��%���F��T������?!�$��\v�_�`E�~��~F�op+�[�pQ�}�b&D�4Z��3"^���b�>����E�~L�xޮ�|��� Vp>J�(1�4�#�U���N�ĞԲ�Ȫ�׺$$��og1��U�js���k�e�]�Q`$scPA�f"� =��Q�  b.�K������"��c1�J���<�X"�XZɪd�R���kh)��\A���xa�`��D��S�L��fCkJH�ڥ㦩jm�v�L^�W������г�� �X��4�e�/���($����4&���T�d�q�.b�8����o�4�����K�1&7f�v�W,��$�X����8�*=w%��ك��X����KR�����Q�AQ,���CW2��%�����J��:��&~�讀�������ӟ�B�Sē�~ݽw��ԯ��e��:?�ԑ~���PJ{̮��\�6H��+��îa
Y�!�"��R'�`�Q�vOR�ҭ�Ps��D\Jڵ��^�E�A=���S����ƥz�#V��D��P]x�&��Z!l���R����|w=>Ԙ���T��$�?\���PߥP��\���E��eR���_֐7�Ęy�P����~����ɺP����w4jGлda�̰�7�mG��Y���糗�׫����9�Q�W�>���C��������bG.���ݨ�\7�����io��R���OV.�{e�ʤ�L�'w�g>T���7�UjW�-M5=Ì���^l���V������� �U������zD�ˏ�#�'M���׸gB�L�ώ��l���|;h��
S�+:��R������.��s��X���mq�)7B���i�����֙`��7AI{<�#�X�J�-*�Z��Us��{�~d��Cm�fH�+8�;Dn�wv���«0⽽�5�/�HZp��������x�P�G�uF�B#���\��� ֱAB$�T�Q%�Іk�{���*txb1{�m'J C�J?�笰=��P��#tWJQJ���΍�n��pǏH�o%��<Bߺ���T|PF��ּ����xjemVd��x�8�3��*W�sp�v=�hl�/��줦����2-e�cuX��ZΏ��rG��|Ek��d���wZr�h����[b_��dk����/�_��~��3���+�X>L��+�Y���ZU9QB�$���(�� ��u3�K�y���m�T�Ցx&KP�����s���ً�"�}wQ�R���D���(w��萠>�	��`��\f`�Z�2�$�H�%�j��[�z}��ϢA��"�0V~��7�P�ct<�Wy�qs[�Ɉ��Uq�)(ٰ{�Z��8�4�OB������; ���v�c�m�����=Z�.����
���LBZ����	�x��rd&E��ܓ)���8
D�����ed@
O��Àu6ׄ�FT4�?V�����c���$l��2�'m�އ�f~���di�C�j+��{�B6�h��dW<�z����[O����"���Ђ{�����YV@��	:����T�dmO��	i�-��5���fA�T���.�Mi�~������h����K%��w�;6������po�Ԝ�i\�W������C%"]e�KP4c�6������fS�$�J�;��9LFV���"���{UB�_�;z�0}}�Z4��!'8�����a�
S��eD���Eū�exq��<�Y�ZG4'p���Vj�D�v�e`"p�=ղ��k��./�;�����+x�Se:�`Z���\�?B����@��l�������5�M�c%� �/�i}���^���z�8�N��g�p�-�%Z��T1�X%z�\*��;�������O�0S�XG��K\TSWt�,�%�/����&
��V� �%=H܉�Vw���G��� z��]���CB\l�R�[��c+�e"e����S��.����i���
��
�N�߀���Z��� 4����L\�+iQA+�ђ�"Yt����u`#nВ J�U����/X�`J��I钅��vSװ�-{�l2[�&4�jY�|h�� )jN��Y�����Q�[}�u�K6��`w�<¶ f�zl^�go�9�.: ��ŗ�g\�/��h�U�h����G��ӯӪƶ���k��Z!@z��Cګ8V
�@4Bu���p=3Dx83�� k�O�U��j^f i��X�D��9Uγ�:����\U��$j�43�Z��-��F>��NI��q����\!+�l�V�j�c`�ݶ�ǅrOݞ��O�-���)$X�,��s'��:���W�_%,��3���1C�a��J�6vP�	�@�q��a=	+�
�q�L�ǝ\d�.r�t���BF3�+8�!WYՇ���+�(j��|��m2J����^H�e[J�> �1��@76gn^B�q�q���yt"�e��wM�r�J�1<��䤅��s�P��odʚq8�fl��{xݾÑ81��{����!nY�1Č��2�1�,B�]��uS|�V��ۧy-H�>�O�ћoO������bHk̈��?�A�2��)����R[��vx^W^��_�㵯249Cz(*�I�@.�b-�YO�
 �l[)��F�ony�Hs{�z��ئ��.TЯ�RXm�4B;S�ڄPoJ;͢oR�����m���T�e@L�;����͠1�
��h8旚��Yo�&�ܤ
%W�ެ�e���I�V<3!`��8��oʈ�B�^ފ�q:]�Yҍδ�I��E�W��Fx��o��lXt��Y>:�N�J3x(��$���x���t]G�?�+:�yq(�0gc�辤����k�s�֠��O���#u�Z��t��-D�&�'�_���l�T
w��9���h��@��J��dF-'nHg�i%>�w��oM!7zo�c`�!�#A�=N@�ܐE�!ЀX~?Ɏ�1:]����	s���V��T)������e���B5'�௧��z0�D�)�Յ�J���ښ�,88��D�%�a0E�f�ݕ 57�7 ����x��K��Yذ�\��0��(&����V��,i�����,�����O1A/g�(G8I6�nkG���0U�*��n�%�\~c���h�*'w�����;�UDn����j�be�P��������t�Ý�Jy�Dۃ��sC���*�j��8�^�nިw�N��+��7�K�*�A�� ?u��L8�ݺ���1�Yt.@]��0C;��@} �߲�4�!/=lx�o"��������S��>����n`0_?�'�7��5�L���L�[ý(��������"r[��p�|n�9�%;m`�{��N����U�	���[H�mjk� ��Gq1��e�r�e��ɞ�ޗAx��^
�3ԇI��Yd[f����?w�{h�����!��+�N[��3˧.!�W5�wa�0�|U������I�_�C1��j ��+���f06a,N!��X�ߋ��U��c�6\��o��bh�������^#n�<r�+�����]A���'Z�/���%���BQ��3��a����#�I
&�>�?��R��m��~h#�*��ŝp�ᅯk�����0�Hq��e��nGF�4�����r&���'�֒7��WVÀ�}�"����~��08�b=�o�C��*��=f�d9 �U�^~��F�b�X2;��>������fr�� �k2��9a^�������wWAx�tcCIǱ�s���{�/���5_��-[�m�0��qV���݊�նx����t�����d�$�t��S�V��?U�8(g�#
@�X^�!��īzh���r10e*A��g�D�!
#=��F���a7�$�i���w/�~���0&]{Z����n�n����v�-�s�B�'.�ʭM	TKë��t,	E��nοV�<&q(�������2[������/�d���c粦�c��@e2�5q���֙�Zs��԰ef���L������!p��!ј���4�CӃM��y�B+�0B\ TN.9�'��>v�̷d�-���١�	��29�[E�����py���i&�ho�B���1���	y��T��y�幠^��+Ũow�BU�K(�&Ǿ*M��܀
m=˻�m��y����yt&t�}W*5� �`�G�x4;����a���a�`�	n�ݍ�m|%��: #dQ�l?q���!�
��R��*�d��ܟ��o�&ʤ�s-�L��?i��N��V���rB����n�<k�$� �>P��Y�O���7��m9AN^�i��J{2�{^R��;M*l	��x�.Wh ��50tA��"lc1}'����P�����@e����)��`�%D�ؼry�]�Z1���t$��҃ؗ3,�����MH�qᩃ�����¦�Ǭ%s��GDM�Ä�_�1��:1��A�U��0���	1��Y;J>oa�=�m����c)Y�>��-�������U����
n[,/�a7\(����i�D�b9V3���v7�pJv�1�ǭ��5M
,�SBZ̍k�,U}�M����C���h�rA_2��K}�
Bs�c�sgf�]��a�Dpת���mG�x�� :`	tpŗH�q�S����Xy�����.k^&��1��MiC1�R�
C��?j�nefB+3l	�%��s�$�q�v �4ēn���P�H�$Oq� �4m&�Jz�~���B|+fqĂw١ouM�F�8����2�{{�Bu��Џ����K��Y� �fz{
��xs?�Tn����ƀ���-+�kC��8��p\B:� BU�]
'2���um1]��K(;/�������j�G���R����EP�);͹�>�R_\�{ �dS���l�U��p�Kkl��1a�iX��\VCe`�K�h<$��b#�Yö'��tI���&i��הN�7���ht��N��$���lyk"���%�:��'��ѝ�]2�@Ƣ����+.Ωk5���<��J�wYj~�B�����j��/�����#������b�����(��С;Q���F�1���^z8^.�3��|ʰ��rC��ٻ���q!nv�=[�'�kʪ���"�[���5k�G���G�B6޿��xU6�^5D0�]��� ��{����g+��+�ȈsK��R�M6sq3��	_*����}��4�G�|_)s��?F�)�G+� g�햌1J��m���1տI_K\_����Ng�5�0��j���*�`7}@e�,v���Hg���G=�ɍֽ&K���>������ɸo"��H�׫�Sv�dYP���~�Q�Y��!?���<�T#��3�uI�A�/������L�/i�@�A�j&`�����8C7[�	�'����^j_�-n��.ϼx~��R�(�Z�����|3� �(�u����/��2YV����%�&��'�C�-?ld�[��C%�Le\�u��U[_Ϙ1�0.���M���+`�(3ux�����U��&�NE!�fkn�[�DY�Y�ߓ)Ҙ����>PC���[
���d� ]�Q��&��Co�JL��*��n���G���JJ�N�I�,��0̔y�!<�w$�Ab-QuT�[յa����O[}-��r��&ꪙ��Y��޿��rP�����3�:ά~�Lw ��zۥ��wlۓ?�4��1����A���b<f��2����Ӯ�W�He��0�:<�:Z{��g������CV&�y�,��?*D�=f��+)=��gD�m���K�D�|��X�W	�~����	�u�:��-?M�>`��i��;�E*�j|sz(���lm��@�l�ӺI9%y�=�+���D��*Z��OXr��X>.���;�<;(��?�>M�Zm��qh	����Sm'�ۊ䖶� Ɲ��F��F�*�ڃiT��
kyT#�U��r\��ȉ� FDV�Un<��נ�<�jƧ�t��궙��GD\P6\�;��/��|��� ����vo���~O�"��@� v�2p-q>���=����B�e����3�)-�]>���60�!�x��lیK�	�T_��&�A!B��Z�ۖfC�8r�Q��|�y�N	�й[Jo���4�
?�?(dޘ���`Lu�nS�H��PW�%�>�렩��*Ȯ��U���hL�mf�dD�4�͔����v{@U�+�A�e��(U@N�����h� �\]���,�x��"���G�K�a��G �:��_�����{�Μ�ZX>�:�}�S�%�.0������= ���e-$���"Kʯ���dR�(��'{�P�铰��I_�]I���y�\hzj�����^�7c�?'9L5����0(����o��P�=���t�%��;�Pr��]��0�z��B�ۭ�_+S���L:V ]�:�B�������zM�؞�|��rEI�W��Og��~E�
� �V�\uy�
B���J}þ!��ԴsRp��q��(}��ڭ�u`�i:ڰ� ��G6=-+ƹ4�1iQZ�]�}"ruC��RW@�<�?eR	±��KZ���T�%�S0bZ��4*�|�u�U��-'a"^%3���򀙳����t��S�a��fT@k�1s���*�ioC�̷�C�h�f��Ñy�,(:��@��Le�`4_�+�9fʻr"	�<�$�EC�e��9�b��5�.�J��N�܀_WR���kg�I!��#�Xy�����-�әJ���W���d��X�b��S'Z�����GörAZ)0�c�I��'V��=��҃�������)�u���1�ִ3��3�eh�I�"F�KN~�{�+�`/&��so쪹.�n��d["����m@:�8�H�[��6W0��O�b�)8�R��5��k��EX�W�=J��knV6sf�G��9;]k\y�4`/�J��&�
�"H^=sq%F�����Ex/N�,�i�+̗�1,�E��զG�j�	ߤ<�= �t�ɫ/�G�fL�^���S�]����J�����aBl�&x�f%�Z�Zo
�j�g(����9(�K��}���`�MAЯ�|7>�OB�d�S~lU�0<�jQ�0���=ޮ�Q��Џ�R�U�q$ J]�r�:�$#A9��)0y'H��e��5��O�ʾ���$j䫉�g�Z�y�S���k�s���� L�e7��W>
����'^�^�sE	�.Cj�`i2��hr�r������r�<��K�J�[p,���>Sm��0�G������S���ٮO�?�Oͅx�W%L��hE�?O���yԆnjAI.��5��M�Nw��wXf���|�l2hb��(�A�~)��̝1^���۪��銴�sº�A�W���F}K�g�A�}�իnn�����J@�o����ۙ飲vP~3��P)�(�C2���([סa�l�u/�I���j�f�687��#J���ޙRl�	�:t�g��Bؑy�VBg�g�4'@@��L	��|vz���)e�w݊N�}ܻmf�gwv+�s�4��䠌s�N���,�,��
-�� ��;���U�e?�I.z��5j�u?�+�M��a..����Fky����_Rc��Ĭߡ�3����~�L
i�m.WjH�<vI�C�7)��$X��U~O�uNT	������ư�W��X�>���Ŵ�b͗]����&u �uZɹ`�z9"��9�њ��|{���ݼ���6v��;�2N$M�iiA��-�ҺKy/���+��4WkJ]8�P�ϔ}����堯`	I��m&�KLUdA�,����$�����Akb�'�Ak�q-��は��Hi���V�V��w�q�,�`��`�a���$��35��()2mGm1�-�=��R���l�������c���A�{$U�
N��N�I��������
�����2Y�H�U�rE�`=�C��5^s�+n|����v3�q�fAڲ���<�f�}�{����Cq�-lVu)�(�z>� ��De�څ��@��*�z/�Bt���5�!��$��������aU7+��E}��Vs�^Y�u�F�&1ˌ����}��@d�=�Cv���s,3A��w`Eg0��b��M2q����LQ�b=�^�����V��qG�If�dˬ�v������}�/���d�˒(�Ii�(�Fa]t)��o�f�H �X'��C#��P���i9Ϙ4�Cd�&Ko�leO�G��G��� h�7Ӎ��^u��_*���n�cd����F���\^�$���/�NO����c�&.iz��EH$K���&����ʩ��?U�X�8W�`By�Ѱ�N���`P���YC����l�^� �Z�3��Ӂ�A
m4G� Fj��"�;��Rq#� �~�5���eP|xd�!S��1�i��q/]�T!e�=��.3�Z�I����uvqJz��E\�$!I[��u������Y_6)db��������
�{�"$��tǗ[����W*�ugzX���*ƺ����vD��<�ٰ��7����P'{_�V���ӂ�H
���B��A��V�=���x�q:c1�.��+)���j�/n�������m9���Lʵ�F�O�B����D�� ��s&�K4o�|�MZ�Zݡ�Y�lt��?�gV��dag�$�٥2iD��iO� y� 5��21��-������m�?^毾��ܽ���T�|�[�D��h��*VB�o��9ؾ��{�g�s�����>�#mC��Ѽ?��gP��[�)�8[H�/FU�Bs���)��xRs"�(p|i=�I��},ʩ��t=H���+D�����C(�`� ��{�R���"2���]s�e��G%���D��J�V��a�� ;��+�l"�b'_�\Y����Wf�)���p�.����4rΝ�E�^�!F��g-^"eʠD�x3g3�8a�D��0��Qy(ABj�m��BA����%��m�ܢ1+�̂d-��m!�Ǭ��VN���0�Q����M�UN����{2c�hə� f�;H�0\�J��J|>�����9�?c��k[�b7dO'v']ߑ��
�:FC�l�.TQ���<�^��+��G���D7P1�߉�N�B���αd���ah���q�0�Y_`K�`��U�!��|�"
'jc�"`��ū̈́hi<�\���b,�^�N=�cOcpm?�a)�����CД�sk��(r�>W�O�5�\M-����� x��C��B�Y�q@�q�M��Op�s�JJ�]?NmJ�L�8=�e�\�ZQK�{��}I�����i��N�U��T���Z�rQ*a5O!��Ą��-X�2ǋ�q@^� ����h�����0�'y��aP>rC�(�"��Cr[s_-d�y�ƥ+�~�InA}⨜;�y�5���W�s$�����'��4��x��<ô p g���]��)'/�{AI-�v��*��:�8����a�F��d�WB�g�80�K�Oے0���]��RRES�\|�3KB���%����d[D�x��:��44}�}�1�d\�v��X�M1��D�S�F��6��fR���r8҆�n�]8`آw�����Я�D�)sd�
,��x�x3��m3Q
�ϒC�%3l���Z
��vubZ~�f��޼н�uϼ��v�D��������xo��9����ES�~����n�9���]h��<P� ܹ�Fy���H��h�]�d�l�f�P��<o��f�+GS>�8��8h�RIYi�ƽ)
�[F�lY�[b= ^Xr��%z&�e Elo���!
�tZ��yi�j��U� �V�<��(Dp��7�$�5� �D�S"'��bU���|��vx8�����F���x�M%߽&���;I��]� �d��e����r*�<Ds��ϵv���N�}AnL%����E^�����BqS�Ş��n�U�/9P�Y=����Gkʋ�\�k/���(%��-8�R[& #�Qp����}��Z�<��yU���<U��7̭��]A��&0����%B/u�I�ז���'�f��t������.���D���_�9-���41�\$a�p0�#�͌��nW;���C;��~�]OT��g���+�j&wt��7������`�.�х���'h�^���N1��љ�^m�B���qf��W�#��pmC�E ��|7����^��4��W�q�N��p�GR���
�{IB��L�{�w��_��(|f�SG�+��R���G�`f,� 	��J�����Q��3����8Ji���u�����C�~s���;�J��
��sz������u$v��.ԭz��?��3Jc(��,'̸iۻꞤ�'-�iR<6M$���|!�mm��.��oZ���(���\��� ��/��H���·�˔T�G��N4(�Yb�K�m����9w1|\}5H0z#��WsR��G�����l�L?`!_y��]-ll��l���5�os��fw�(z�%���F �}B�U�A�^��bEW�pAM��8��f�OY�O`{�_��JK�w�ϫ1��������8Fq$�.���0$��pGu5���UR�zB ]I�kV�蔤��.O3�0ތ��49Q:���K4�O�d@��{��]��w��@լe]\"h�Fi�&���l�-�n	~��ޏ��B-�I�:`q�Sa:�rX;�n;;��p�	�t��(��Y�_�9���}���ۙ���f�S��ܛ��̻S�:�T%?���_��3�i�c�rJ4^v�+�gf���Y�p�A���}�I`a��u׆�`b.Z��l ���1p��;�=�Q^d?P'J��M4T�%ã,u���@pG�2����9�����7�����pv�r-r����Z,��)Ǆ��V���;�^R��}v�1�Q���J*X�Y��+]�� �I�������tX{*��؄��1~��U�+��%��Xzui�r_L�g�-�Қ���� �|�#�R�n+yG^�Hh���{RU�� �Ez�L-�֤�o�!�i�-�X�8��Bͻ��zz���3������Z3�a[�5"���s)S}���*��2ˁ�� _ŌK+��I�##{�}S��R�����wB�� �G���E��FB��@�|���=#~���*O��kXH��{4ϗ-�U\���DFZ��Q��:#~��uS2�9���M�ˮ�ly��78*��W�Ő�'л�����ŐJ?���($ӾF	獲=��P�AǛ���^;_;�A�M��Z1��a�=���6��P���V�=���쎃+SO��������c�����E�����Q�=kCz&���9��P9�#p2�̼s �Mqg)��kuz=îS�4+�z� ��.F�j��vb���'�'t�U�Y�߉�i�����9�\bG�N��V����A;�h�W�@C�#HO�z���R��鮒|r�H�|s�����.�e�I�/, ��z�)��n�.H��)�g�08;tU	���g�'i�����"N�L�����Gu֮Y��o��m
�~�}��@�W���;&�Oo=;c�+/�����5JJ�b�ጮwJ~���v-"���V�l�����!_5U��Kp��4��3v������f���5�o��vR�,L�-�HZ~I����U7T��T|h�0*�����%�1�qY��)���ƞN+�e��Դ�h������K���<t|ei��Z��1^O<��d�-^ vD��L�P��$O_zq��� ��rwS��Kk��p̻�ڥ�>V0�0xKM]?R-�f[Xgj%�U���Gx�N�-`�����짉Yu��c���1 �Cd/�ѱwD��l�;�HB>��Nr��c����~�+<���زp���6d�L�U'�'��� ����DP?�����+X>���"撈O��cZ1g�x��GC-�U�pIvk����S��������SO>�Q��6�e��ڶt��6݅���.lUq�Ns!?�����rj+ �^��Df���V�D���۠��+*J	��m=���١{f.�v�V��SGP2���,}Ug�j-RI��P]u#��i���G��Zh1�x���N����O'ȕ�"d���� 92{KnU�Q���,-k~;�28�Bn����-jG���_@M>�i���g�I��b̐��F�K�V���h���(Xg`��T��`�TS]�C`�7�1kWm
�i�㵿��Ln���p+�L}d���Ұ-��w�s���}e�p趢��YQ���pksYG#ǭ��hN���,>��j�	�x�~i;ˠPv�Y�T���c	kp!�%��6�!�Ym����;F���pt\�V=3����A��������WF���!Zsn��/����{���~�z�mJ
�xJD���i���Z�W��T<�q;�����Rq$�������B
��>S�ʮ�8�g�ഠqx&N�Љ�Y�"L������/=�˞�In�,+�c��Q(��uE�r�7f�s>*,�!�Uc��y���bR�3K�D�P���Q2�6Ѡ ́���tL�w��I$���h�ںU�
t�f�%�ߊ1�𿑊e������k�Յ�i��ϔ�ZÂB����-�4��u��ҋ������B*h"��Fہ?0I޶�'m�?E�.�"�����y�D�:���i��ey�ғ0���d�}��eFL88y�V�������X��`�A��/fD�Ʃ, �]^���
x�#���V�Wh��27s5��^٫lAe�6����-�b���9�rwjJãB��S!��W���\(w���e��C��Q7G�/l�*�Niy'a���(��oo|-�G��;Z���|����_��qc<7�.=8�lPL�{(ϣ)Np�?�DY���EI^�Y���j7�&�����N!X����"�v�ܦ�����IJ������������ojJ��Py�RГ���B��(���;4�����)m�c�3X���-���� �8i�	h�a�YWmG�s�A��ϐ
�Ϙ)�A��7e��e���8;`���(��O�����@����]����|=E�B5� �V�l#V�}h�K)u٤b[y������!l�5��V`��#�/�J�瓎�9j �,Ԕ�	T���1Boqn��a4��X��p������ ���կ���Z'��M<T3�������Ԯ=����L۸=5���K������x��7uzB��ٍy��L����e���SRR���7�w�\�ι$�M
����Si�έnb�yk�P�(t��z���U� ���]|��~��J�p���ߤ1qR���oO:r�	c0�^9�u���şa=�=&|��#���΂������I���X~���&�.��A��z��+1��3̓�wg��>C��!���Maes��_ciW}8}tٖ��O�~S��N#����DM6lo�wf��GBh��S���
���-}+�Y���B�����؝��Q+���.
��	�Ju����t��m��>#���:Oǘ錁ջK���B��_�So cZ<7Ř��#�:��'@�8��du
alݮ��۽��;i!Y��^�t.z��`����e� ��6���/�=�ތ�|�k�U݁�����V�+u&���7�Wo��ey���#�2��s�7G�!h
Z�v�wc�N�˼f=��vG�,<f�B��������`�)�YN̥g?.?�'C��	;j�Q�.��5"�B�N�F����:�1f�-�А�)��
i�(�p[',���am?j�#<M�����4��WN��.�C�]a�<5x`v�N�Ě� ����v��>A>�cb����~Ah��9�|�ড়���6ǝE�g����T��Y)��&��Qe��1� ���Zx�����
�(��L(���4����6��>�v"?�1.�=.�t���|��
��=q0���g?�f�'���L���$��������d�?�=q
a6U��h����_+�-9q:�C�D�=���d3�?��X�Rr�������,�!κ,�<���bWJ�DТ��u;�0���~ϥMઉ��eW?��4{���:�+�5��_���hUP�X��{���EtT�$���z�2�F���r:�W\A���S sZym^��h��׸'��n(� <�tJ`���Q*�0�&�T�+��֐�o�}5_6tn2 ��Q)�����w06=d�jHX�	[@�MɉR�~M%D�P��������%{��Ҽd˲�wո�¨�#p�c�>�/-���
]��
̸�� ,���tX�5�2�(��%te�l�n�}̐�ٰg�����N�i}_����Y���p%��.�]!%�1&J��m jb@ B�rC��������xLUm��C=��1����߶�(	�eW��jJU��s�Qk7����+����u1���o�<i�$�G���}ٳsS��K�ޝ���ui3hmWØ��>�H�*`�w�W^:��|�l��0XG�>�b�^Q;����(�v�#7��Xg��X��oh}�d�7��J���y��eyT{�(&�ql8)6�)��%R��V�X����6D*���Mx��Hz�)���^Փb���Ws�?�e�Lx	�2�BV�Ox���3�{���c!���SS/�P#Z��F�(sS/8�o���C��y��%�8���З����o�x��պ+L��^YiV]V%L�펍�x��!C ��ɮD2*��$d�#k���}�<-�C�͜
���i;�W��@�I�Z*��2�W��N���MF��G�̾?�L�M#�N��m��n��3�o6�34ͯh�%����w�������l��
8�4t�V*��B���?�U&��ۧp�*3R�,ГD���:�s��I�o\7nGt+A �)��vҾk"n_��Z���h�iՌ�?!���5ce���)�}�������5t�~��%��0�jM"v�I]/�q�(�-P� ݥ�. I�J�|�LO�Z>cd7��ہ�6\��s~���K���ڑC�
�h�DI|�츌�Z����(�L�����B��A�5ҵ�Ҋ=y��z�NT���	��]I�d���\Orx�g��b���*n��'Eȟ��5IF��X�1�%�~]ZT,�Z]]�ّ�����~7��A�6�9�w�Oa]d{o��D��d�AK��(�8�ob�E��7pW^�}��`iTGSR=�
�����0��s55��K���e�#�SP�2f�DI���N�y��q���Q9����/ͥ���-���?�_��F<�p;Xhd�mi���=;�2��m�J%�B��^%{l���J/(�""im����i��Q��Z��C1�O(������&3�[:����eR�9_�4���9pt�S�B��N�۬0��UU@�j�C�2��]��
ˤ+w_
V����K]�;ؔ4�E��{��!���ꭙ�Pޙ��kSM3Uˣ%S���S����Rd���K���&�]�r%�g���A��K�T%���A��J��Qҏ���]F]u	�h�����w��N�Y�N�Jw"/4*�fGz���hv-��m��Kq~��pl����B��p�0�nPa�������|��i{��;�y0�k?hs��ǹ�4긾hևh�/e�EѸ�>�� o{��I����6�3Tx�!l�l���o�{"����a��H�:��^~��T)n=,z�f÷6���y�w�/�E8�?r�tt�
Z�u|�y�^'�hv�V�'�0�^�3$F��e�J�)Q؄[R���6}�� �=���SM ������m�X�޹č��[�-R��!�h1�SKP��M�*��p�����1o�	f��)���"�T�;��O6 xX[�>��M��h:=Jq���8)N�=r�q��[v���~�q�l�z��=vq4�_����)���E����X��Sj���p��9�����C��+��M�xotc*��k]��8�*f\Oԡ�'a
�%8��G�柖��<�ΐ�*.u�ˤ�����u�~���B`t��I��:M�Y}O;s<:Pi�<"��X�L�R���lu��99i���N�u����0�+�qܵ����5EE����=�B� �k*t����D�O�Ó���,h�[g�d�ֳDa�?c�k�t{�����c�yt/v,�R}�w��y ��ߴ�%��i�9������f\�T�9�[��IV���=FHQ��.`,��rCi��1tI\W!�YW�L�H"���Œ=6aȂ2)���O�����5��u��]�����^�����h��+�u>j�f@��u�Yv�	��i�����	ބ�aJ��2�v�Q�I�(/�vZ]�iE��A�.��Mo<GQ�?DcB�)PH�.LgZ��m�.�p����:q#4��^��a�S�C����+k��ץ�an�:!~��!<���1z��������M���_-�ݵnwb�N��w�H�4���@�v�W�"&=9�F������&_����mկ9������i7<��Q# �<ZϤ��z�N��	R=O�vJp�G�zab��^ئR�(5��h{�tV��j�h����+x�>҅�L�T<���eʑ�>T�PDPuv��p�G^b��#�WC�9�����ϐ��6��|����C篽���k.%9��j0�k�W���F���j�<.7L���w�hMn�7���=�/u��(tC��pZH� A���0]�kU�n��7V���`�t=sW���9�Eb���-����`Y� �3

��A����N��vo]�ɱ����mQ[v���NҖ�%��(�t��y=:ȶĞ`��aq=�����"�����A���w��'�,�㑾�6$`���l3�IWW�v��b��(Y^�o�J��N�_7h�Z�L�V��d���[����W�]U������ږ���7!��ݰ �o���o�`6"�|�_��Xs�T�#w���nK�!�}�(d���L�R;Ƨ@��VO֨�5W�lJ�W�P��'h��)��O�j�g�天����=%����N%�����_-">*���R�U�x���>6�/js$���L�x־����h���"6��g~����8!��l+����9�<�?�KM|�&�jp����Pv��|�3���]��R�仆�@_��sՙi���ow�K�����H����|����+�|#(�~���
b{#��R�Xe�JZ���c��_�p�j���5g6-��c��}%���!>�B �!�5��,:��18�m�b�%&��<D�Ǵ�@��:�Q�o��M�
�X[�>k%��~�� Î�tߤ������4��^�Ж�i=�D�D����qg��f��ę�Q��]|�W��>V՞d�Z(��Iq��f� =M��u/��JD���[_%'�?�y!�#U.I�[g�����C�H����c2�a� W��s�0�gK�\o6QZ�X�p}�%����������}I�������Xݪ��A�c��\Y�1u�ب=o#��d�'��p��J?De:�{�:Cu�~\�����x'$~n�p���r��&��ѐIx<f��]�a���l.g_�f_�@#��������S4�����Ȕ��Η�G�C�1�.!���0��oҚ���I�����vs�2{O�:5� ߐ���8=Fv�D��� �;%! Pgq,�w``���0w{��@8����S/�P�*���[�w'��DB1����{�b�Wt������=j3��ԏYd��$�
�?�*�)4|��E ��7�I;_����ժ��� ��Ϥ	l�����-������%1�����S�q�g��ֲl��}��l ��n=�j#8z�@�K}�	ٴ�M�`a�f5|.����E��ט?���Ĉ%Lj�3���tNԶ��6u��}�:�jY��$^��6w���^d��|�/�f���2� [h�|�4�od(;w	<�2I �}��m����Xt�%��nK�VMsK1�?���O�����]54s���N2�(5�Y[9hΞ���a�aB���ၰ�%�k����k���^�hap~���؏�t�?J%��az4���Pw
�V�*\�0�%�P������f�rhQ��h�M����4���Hg��t{^{IUbN��~�@k�]!C�Qs--P����؉��;�~h
؄�:ÉC�;4�~�_@-�b�ߥ8��0�3̀�{Jd�;��bE�ߝbx	@�~&�d��sO�h�-�@�	l��^�\:F���~����&�P�V��e�s�Eҳ- ��T:]��T'm��頚�t���^�_W�Ң�,(�B��r�uu��5��:i{�b�9��*��5?� 8n�
��VM�����#���Wkv�%oL���Q&���u[dA�\}��55�v�>[�9��)�A,�`����a����?�:x��f)�f\ӽο�F�Fp�;�8���p���qׁ��Y<���vu7��\��%Dl�c��ܲY��;ŗ�I�4��0���/�����.Y$��,�^d0��g(�O�A�gi\EM��٠��HA���Σ�����=�����׾�ϸ:�8k2#p�3*ڎ#mye�y��1M�A����4 D�=�տ0Kش�	.��/���R,�П+� [����L��,w��2v�2D��!����,�9�]��CU����s�DV'��}�4f=��9�Y��^)e����.����a>ǉ�d!���`+l������E냳��������<��9�]���'Ľ"� �e��Z���nڱ\�"�V�U�v���	�.o&S��IrݮP:�<(�2&�n���s�&���u߿��̳��� p� �B{��}�F��h�j�/VI���T�UH0X�� ��]�)�I�v���F141���)j^���ι!��psxGբXk��z< �� g��E)�`�}~)T��lZe�>�}z�LV��%s�n��M4�ߧ,�y!Y���wZ�V?_����<�7��\f5�7����p�$�Y�}z���~|�L^��2��e[��L�|���o��G������ҵ��L�����ja�iO7]T0�Tȗ� /Z*m;
��D�?��nPa��~bq�>�V^U���xqI��@V)��H�ͰX��9�SRQ:r�⽃y�&y�
m�4.5�Yg�I?Mɗ�	RFp{��m���U�� sl��ŘҐ�q�Sg�6��}r@�h��궽���� ��䢫+c���q�T�MI��$�� �W��n�2۫�#��K���M7-TR�.��`>M�=7^|���ZS�xT"BR����,L�6S� �%��W�n�*�'�:�����{3��F��}�?QL��ڄ�$�~�.-~"Pnq�C���^��]�Qf���@`*�%�����r����m"~� 2��$����NX�*ס���J;
Dk"Q�y�gQ�cp��I*������,OB6+sK��?r���ь��2�M�8ղ^,v%�
�����(�Н���oԣTq�J������|MNn?��	k��ix J�d���{����|1��g�ބ�^�u��xr�/��/5��`��"b���uNJ�o�����\�I=�K���T�m	إ�.}��^Si{�Q�͛���^Rx��i#töY�0�� 3K�(��8'�	x��`u���qd��;3��[�DY�@&��ñ+���Lϳ���}Ӹ?K?�g�Us��#KW�.v���u��H����G�J�W�h�qŎ�򬈪��&�ѭ�N;��5�� ���O�Ly.]��;��<��d��=9�&�b,~�S�4�w����#K�b�7nŭ�!�)P�8�Ӧl~Y^@l-��>c�K���(����#��1��z7�"�����c��F$�R	B���q���w!����l�ͯ7ҩW$ۗ�a�HM{4aM�J&v!^�
��]�X�����j�S��Bh�˸�q��*:��eMtn�#-r�9����V���ۊ�i<.r����nՎyz���>}����㶹����;��"���l��,��V���N�-	/�#�Mz"�����xlKG���W�^k\g��_`���1g�/�מ)��Q82x��)���:�" �.j�橖���P ��r{e�`��o��K�ה��