XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����PQ2�}�+<W��~�?�(2:v;��ĥ��u�T�$����o�E3�o�
����r��D��4��_eq�/!r��Q�.߼=���hw�Bɮ��W�>�N���n�����fppu ��*2)���vW�]�9�dGE���9 ����̾^T��*�Ál� ����#U=� x�<{���<��\������Q��7��Մa~Y&��6J�ϊ�dЙlV�����7��~6ekO_7�����<��YF�\?3j�@V��|v)�4��k�om�w�k37�9*�I������`FG�oԽ$Ǻlǯ��m�(���D�}f t~#�x��r�.��:���qO��j#�2��Ms���걱�f*�?� �KwM���a�%Y��H����;!���v&И����!e��RVlS�H`P��)>q5)�1�pw���.4&8f���v�{d��]SG1�yó� �$: ��Z�y§v��ꨓ�vԖp%�h(X�(�6WVx��2F��q%c�Wq��E�.���Y�RE��(�X�i��Ċ�y�Sj���$�N���`�lQc����}�+g�a�C�nr@�v��`�K�|���>U��C��D�t�J�=�r����ZZ����B�M}�~%�]E8[͟����4焴�XR/y��9��[!i�߉X��kJ�q�������{���g��㦃_z`FbS��?�q"]x�;+�9��D:�E|-��2�����F[��{���힊騺q�Q$�XlxVHYEB     400     180�]G��u���#Ϟ/:��%Ϸ�zZ�|n�U����w���!.,����0Z�� 4>��^H�`Ox4ܲ�n3�_
��""g��c��٪�I�+�@��v�~�3?��l�u�媰hs��dT��:|����/��y5�|�eN�o�x����ϒ�Uq}VF����px�<n#4�"*^�U_1���cІ�T��ނ���0�ܼ_��Lu�m�����^1�����n��cо6�Iu曚 ۥT>�Cd͓k-5`�����,	?�;��̖����ww�EN��*�� 7�炟c+�1�i�N��u4��.h
�G�j�2�[�_�������0p}���!C�]�%o�Z�h�:�<8SS��P�%$�o���?K1�k>�XlxVHYEB     400     160��b��iC� #:`?�HCD7�����ˢ@oG_'j�������;�K7��}��*�q(q���I��2��6G��ۤ�~5�]6�I\�������挢��yC�I6w"�/�eŅU�����@��*Xo��.���R/'<dBYZyJ>M<CX���`s D�3\�h�vӰ���� �Rw�1��7	ř��u2%{���Mhp�Ӟ����@f V�����䧎��4��&)x������g��(��[�:�G`��Ϝ�����%Au��?�r(ى��R������oU���F�B༳+������zC<cLM,'��I=�$!�����œSZ�#?XlxVHYEB     400      a0!`�	}�E�Y�\+�4(J�M����߀�Y�g��o���,�������͊^J�Fb�\g<���E�ǅ�I�����\���8�{P��� ��������(�\����Яb�z
 �#�AG?t���\f�D����9�h/朦��y�w��é�{<�XlxVHYEB     400     120�I��(�b�祎"W��KM��0*�N�(��#�/�2���;���3G0�����DPH�y��+M���w��$ܵe&���If��p�F��x�ߚp�����$,h���)��hT�w�̩�F�@}1X³xǙ�`�mbU` 	wzu������a����}u�;�D
*R���KgmHS��_R�v%��s�Y�rG�0M4���ާ�@%N=�
a>��>c��!�m�Gj��OY��qN�&�h�E�5r��b����Ջe��$�p	�b$��XlxVHYEB     400     110����MK�>����65⾂�5!º@|^� �(.Tpu ��T�c�BK1�9�#A�)y��zcid������<�����_L$�ch6b3����[U*SD��9������KL��;�s�=cBQ}�"��H�ن��c�@e�(xM�y>.L�MQ����s���j���̩<]k�766�>N�~��WT���p�hA�k?�7o���8��em; �n1+�̇��w���h�nEm��Wk�L�Cӡ�@������c�6�z�XlxVHYEB     400     130cl��n�*� ���.�Bl�#��tr�Zp�|�զ��2gk���pc��T6��J֝�����7�?q����q��v)��V�D�� �Hl������3��S�!�0�1�Nc�U���zd��W�����y���R���	�\^' �>5^D]�Tl
;YV���u�,"�R�`�$C�C22%#� MC "�!��~0��M~TT&��8G�_I�8R�X��\E��t�ԢR�_�?cB�vP�j�İ�#6���A<�h�e������JO]�x{��-^ x�~s���u�]��,sS��W^ � �c�X�XlxVHYEB     400     130�n7O�[<g9��n���<��I$4�x(C;�<���ԛ��Fq����i��S�1�x�7[IZ�X�HWa䄪�qV�J�
���7���n�ժ.�i�Ӊ�U���,2�=-I��ڶn��%L�_r}aaE�m�p���=C��M� k�>�7`�4N�$$�~r{JD���F��Tt�oJ�+��>�ZƱ.�O�����U��a7,>)D�(=J��l�B�'���ӝ���X���ޣw�{�����U[���������~%��g�-��'lV�:�#3ۚn4��5�2M�����d�S�XlxVHYEB     400     120	
M�:�i��vk����5�!p�|E��.�x�1�}�����E��:7����(x�:(�s�bv�z�nD7%b��705=O�����}v :H��0�+u�����4A:�<m�\C�d?�� �1�_�zAQ,,^���@^�C���	�m�й9�l|���P�*��boowc�,�c�\3��x�IG�p����"*�q�VW��a.C=�c�O�M	�D;i;�4��1���]IVz�D[ v4%Z��w�#x+��D��㠃`���b�樠�+XlxVHYEB     3a6     180��o�g�0�V �|c�M��̳��P����>�0
I�ןs���\d��EU��i9
�ʇ��D�Q��D8X7�T�r#=U:#]_�l�Y�C���75Ү�wP��� ����R_�����H��)J_��QPI�S\E=�i�MKx�ـ�e�/�"��"�׸i�}˳�i\SjV�(|�i���y����;E\om�S.2Cn�zF�H{����O_O�KHP�&|fz�����Ny)癌�V�<��ؐJ�Յc��l	/9%��о=���8��IolC��+E�֦����ӛ�X���k�qߋ��;y�>��2#ְ[Z��8Nh�P��UB�kLL]#ڭV�-�t����9;QV�s
�_o��e�