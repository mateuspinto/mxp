`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
LRmaskcxiNv2Te+yXg+macnYjh85wZ83GaLhYyAcSAGq6pwMC4vl0b4XNv9bkx9MmXhcfdAilYNz
RyPphtM218tcvzNYKNRxVjVu+V1c3rDlIdIhjN4sEI/ueYjI2LGQquh6kmVYMUfmTrrfx8v9G7vN
fhgAhtLJMKxGhhiinYT8VTrO4dB6sEzaYECbT8ubtVOKKNuxt1Z9g8tYbPPzf0SNdVQdTgI0nWx1
B7IhtBFTyucR8RJjmHdc8m6Ydfh/ba1rDzrOzr31soMdDuG+z0IKzDN+Me606bhdqy18B65InH2S
TiM/Expdghpbmhtqbz21ySRPzRGiZ+WO0OtodA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="NQiS6ZV3DJ1yS1n1pVIJxex5DXWq1dagwWc93eIAxGY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14528)
`protect data_block
cbYfIl9FGG9zc/2HcgkImDrJPzY13OFNiajwL4s7frfoxeVTFLWtVreSWL5kvSYE4X1K1smknm8x
lMBHDeiIwJ9CULK0jemRUwUyx0JadtzwSMsv2+prrSVpSv8CeIQLct7oiUNICAwzfGGfYjP1DOTF
hTwaTJvaTbNSTq2UOG3WWeAYvlohVUnfBucV7w7ZB5v+ocQF00DZWhOp3JtHgMhhgkKHxm4KCrqY
CllD58TQrumdfdBwneTGGhp160umBKHiLxV1ocW6qjO5GVL4ShsV/QGLR/ZnJVkN4ayaFrfOC4Qs
rLOHQU0ZaqwphJKBjlGoCcYRkis2acPWwlloWnVbJLasAWnPc5aD6HaPaRnctZMW5QL91tQ1RDh6
/nqcWQ4/dD9feAsfjtZIN/eMvo7J+a8h/OwlTXEn00vm0cf+T0ZArXpKxd6WnaMcSupP06V+JDTq
vX+x1n0BnafdzgBXXk48xyJBkKzIBODmyrYmMSLQbg4XYR7HQhaYpRCbH5wDCSHEqGofTFlLhkCp
bFif5Zcgn+QVovn5FMP32gdF8YjN0sUCBbiT1UNm6EZIl16e11QY3/ln3MiZU3zOrF3uspo7oZhi
bw/mKJ0sb6s27ukpsBlUOW/oFFGuO1FAodVvVCY/GNk/3xPGjt15xDzjaJke7+Gfl3WmRZ3b9lDV
RSa03ARnW97e3Q5FO0+JT7FYE6ygHBXyAee48u0iXlisYwc5WHVFpk0nywN2SrzQ+pLqXUhKFSDf
lGK0uP2kpXi7QMaAjiUkE0YlrOxJvVncgxaqnCVTg/VGeCUhlFkhzg45OCC/q3GOnh0jnyDe5+t2
HYQYRvsEsI5bj/djPdmJcTfk2RYhWBhE854PdOouJc6xu2oKcAEjpoKt/W3sPuwXl9RrEg9ie+At
RQGcvj4zsa8tEaSn8CDKGhVGn0bz7UA6V9V2bYnpitwl7b6Pz0VozHbzYbs3dmThun/n4elxg/jL
X4/m3E5gQk2U1frJf+IklAxlSIFG2vHi37JtLBy9QWqKpR52mw0U+a6qNaDfFTxEFWtb4/hhiv/5
fu/ruNMksyCf22DmEBBk2PWoLbenr167Z3nOgJ6mzFSX2I8bHQiq77mDG73U8PGsPHcMQNa4xsL9
t9uWrmcG43/GyNg/pavuj19hBg7nuYhb4MArLDxntMwdN21o7mLJGRrOzMACAFpcoPI0ir+X/mSf
Q/Po0krzm8L0vimABUNPCJ+rj2BGiHndrn1jbFSM8xa+2dXs2QaIJq1X1yeAQm6UCtmkkteavVVt
fhigyn4caL6ePYpn9ukMl6lMBo+1MM5TuFCQvSB+AR7mDYmco62ui1t2kFawOtSKUwzBjA2189mz
/MVPLaym29Gy6sfUp+dov9uw4DxbdgDaz+t6zoVkN79TNZEjSi2XqhAyI8BEjo9ohGXFx1JhcXyY
xxY4OyXT1ZqxJ3PjS8BIyKcdo2HfKvJ5B3L7u09Dz096ErI+KTVIPss1IXtxw2GLaN2NHZPk09Jx
idHQazGVZpVPuxPIHpyE4kQnxM3QnCBK0GbrEd1Y5BY0SIjNanvbk+DeVPK3DtvbpM5V6VLqvFju
7Wqh5sfxE85G6OZ941CMk9VNoyMGwEHAOHeKrShmODFwpKnQBNLmD2WxlQjIPl6talB+Jk9jqaP0
sI2gyRdiuDhc0CBQOmFUP+A/Iziku1d+0W3E5VmW61/UBn3xtuWdfoj4v+pJnbR+iuZgQH+1YRX1
12qxKvD6EZznS/7o6QNDV04KQxbI1HutFpD988+Nfjxyz+o/y00ju16abAEbxBiV6qtyNBYMuWV4
Y0i6YVxdCZAhujiH/HtshQ2vzf9cthcm+frpHNv/GF8Ws9yoSiCK1gKZi6FqP+AqxtpZWJIRE58K
a3PmCjdxU9jNwgiKL7H8utLaMKRWYyu94ebJqmciW6bXefbHnNk7wjF0kHGXbb4FGgVjZ56NEjeI
5G9gFA+BBUMkInog3itfssZGUhdcXBjRxJJ2nsQFMwk8WYj9kYTFd6xzVf+kPsTj/mm0AjcGq5wg
3tRi45ZcYX+KWgFBdXrdwaNUa4RfJ/wP5NnTByamPWsyddg89sRGWzNwIMVI/AEIG+ObF4TTWhuF
SL0nBDZiBMFyM9lwtQJp7/QDiiwLGovC5AHnwLHN5cXcAB2Lr9KZx3XwWvq14pr02RvMJQildExZ
GFAupLPLRbw2RMMg2dpox/CiUhhZ1G+mvOgzVRQvNv74EWnNS3Rl5tPY7Sm1CAfNvldTfA1oNDCo
hRgS+AAw+Nzd85jeBUu9NCZ7BxsoYh1quooS60MmYvwtvprJy07TlFIrtR1CH0xOjKqkVvxbi+f4
hvUT/syzwCeKQzoyZ/XQcSb6EWPuw4ym3pXroLBEqLuXpSp4k9tQVNvkJTnef9uGwnK/ZE5OH7hy
sJCs98GKubaukbld4sBhMycpH3L5ZTorEWPgvj/UXYrpdKPzffS+YRij0Ef2aV/AMaIgJRrMzlLo
QOTBk1XfN64bglQI+OymH5vmS4C7kiNbuQ/rQAd4SC8fn9cMXi4778Qi2IVleOPq5njajFrEdOOy
g1QjKmfb5QfO6rv1fWCrFGuu/PG6Sc4adBlllrsTEKhdkJZMXTLpuX+RotkgPMmFPUeMYXhKYCWt
VbdGlEIgAt0D4WKYzFmfxTm4LM0qp0NUjWhU1sp+u/o1gz7UQHLN3sJrvnXDGdf5CvIk7JfOcJZ/
z/AcuFeQiurW+Gp7x9LrL+Ko0IqiX6IL2Pjrsi74+AxNA9K06loX44Remww1GmHJIBw79j6BPrQw
DgUA3gyH/50oJUlTl6QBMRfNmseShd3iJSUn22FbUDbRPd4T+7c+Vfy74ECKm6j7UyL7p6guBXKf
As0I+oh4J3HEYvDbl8iLZ1KoDywYFpR0330b1ROpSsA1qUlt6GbMV29YO3lEYOlu+C56KwJhQVhx
qdRsLabhSS2pLinFSbOxDGAKTF7z2RxxjjCnXBIiOzVVBNH/wGiNm3FCPxJWbSXgUHbl4Str+mrk
1r4aJd7KB2QdbUGwx97iRykptfdPUNCWa8dAKXEk/v+ohZQHDF6zfEU6n+dwHvFCBQv3TH3OwNRg
Kny3yKsZHKP81Y2KTR+CasZnKldLdZGA0ynQEuELBpAsGRKIJJJfZC7jLYKRdgsoNzhiZaewN85p
C+S9a+WaKpSX2kLS6K3dwqMlhzWPZ60CJiqc9LJtM0/WQ77LQNGhsgDj6xL1BK0vuzt33iL+A8L9
DDISrMfYgxnJQvPpCIQzMUE//v+LM60kttCV5GIbFtN87wV9o4KCgyHW8UPBiiJJMaKUq/FHcdKq
rIJubdIOjVqZcBPb9+cPcPc1l28zIY3vMkdfofExYu4/rnofdYOyZg772pukvxkg9dehm4LzGuF3
9YPkDjX0Aw6pPUha1yXqcg8CEFsCT+zeJyG+bT9wvQVa4P9MGnmjHqMy4s3bYnhqZ3qdJ4OeZzVc
flBElM9DCuYO82/kvhtl2CV29gzmgzPuHVW4P5uy7+dJugm9s4THL1B7Us8O1UhpzwrpYhJyKodw
1HpKZTUruypSfcB23GIj5hsojmDWy4ohTV7p/71MJ4QZvwk8r4S0yCpHhPMiJYYji2rQmwp9cVf7
6UN2e6dNPn9++jZCuGpJl/Kt727EXUZxMQ/YUO2/iqkcg/BDB2cenINkXh1Z8T8tbLJenpnawnjP
Gx476yNOWEgfgDlQ5wzO3IDbkQkDZssSpqyDPTh9DhgVTBh4jO/op86T/3oh/lbHLyRpA4iSr7qZ
pGpih1Wl87Pp4bWu7HXUHISg3ES/Ka7fjY58mhVwMSKdAWWtlIN/6O1pbHchrQ0Hr3EdfFORKi6L
75mTdrCwgWsWll5qV9/5/vI+OlFtK0Nv5ztp5mgs53RMAik36Mc0UHP34pCgjAgjjEr1468HEYq7
oQ1rcSVjUthp5fFlbtvB0wewmZExerl3tfrJ3d5974yLDJ9o85w+T+7lf8Tu7tbsHVjve11c0wIc
HK8yE1Iku7StxegQq9EWczPxq0KJLEDyQFfPo+/3xWeUcHdouyTVL67eC9L3knE6DU1OPO5Li2uA
Ix48KvDpP7jJk3ywBefobXu2yc1xHnPVwafJJ9f5pwNb0NisgfL2jqa+dSOR6GfigdnoKpAmJbWS
ihYMVFvy3cQ59DQIeOFNSBStj0Hk0ZQkPwhMQmjE6v/KnS82WOcX1Lqn4iCf3aOrXxNlKvjDhq2w
R8LX6tHs+ij1tqsJU6DJ7DVe1kSvPBP2wD1wbhWTVi7+DPuyJyiJ8J9ES13hcK6yUu862Ju4JAOZ
Rv/I6qSuc9yINwY42mtULsgaE9KP/jYZ0HhUIw5ptmo8Wl0VrRg1fWdysmH+nKzYXjkrJI7N8grU
aDphKTbRlMx4WyiYT8m6JeELVcLyb3D1azTvjAXITEgIyJHVpMDzp+hyoWg49hDX4EwKCcnI5xQz
p0wQL/i8hzk36+Kzs/VcNZgkQ3+ZyUckx1Bsumy7FUEKh/pR3aWgE1+M1vVSjr3yedIGgvqfNfAH
UM36q5LltMmMDmYAwSGtGiRM956wmIKplOLGECv6bRUDJw8zBY789FXeonVDatox2rA/Eqry6sBe
sNIwXaKrjxWmE0r/3ize5ivgyow5jEX/8nut/a5Bbyk1qMmtlP1z13dJciF0kvDNJqYv+42+TtBx
1JK+jF3F7l0upv+B7evfd7Khx+q/Vz4pw9VeuCOsrPfpulrhZushuDmLYw8ieDoZ5sxs6fnhP+RS
vVWa9aH2FpqWn5igDin0Tcho+u0SJofP0zx2WP3Azt3zay592cAx4rPFtqFf4o0RIfJnduazoWaO
yFhJ/1b481BpuRuH3gr3oOFcANO9qOa5mJI0zMwpnx2+FQJnqfoS+Ir5a4zaJoB4vyPJdA3NrIyi
Z/S9EJgXH0Z1+D3Unheh5SZMrVkxBv+1U+09JqTQArkml55VaHgxxvN0BN1xJKOOoizty7KwQtbs
+6hz5+AjIbywgA4zPpW18c53dDmYB7R3QUK9Z5NHE0TH6VAVqpw0VdCJ9LN/SbsZpaulHGfMCpyT
EIdyRci7uQ126V0NlwF/v4DJIshoQmSmg6mDV9WEm8O0MNSG85IomlGHEZYoqSbT3wvIN3Sxl/XA
Cz9w65kl4FQ7we9JC2ig8/LPFDn7uDMo4zxnG5OxnxOekR8PdNJ+NR/Ag9eXxnpOhLRXK94Vvt3Z
z1IgECFyfr2SUgTOl3FV0FUctSYDX2fttqFJUSzXhmhujnoh0sjL7obzxNIkuEsW38ECcxR8j6Re
q17kUWDkGjtccbFke0frIjF7FMEB7h8MBAre2NAwdQJfc+VciQ4lXk/YXnKgNckiZ9v1ik8plsQ1
dso+N32CpCgv4Vknm1cC2E2zE62voxTjLlwOnHID99j71O4SUi6heFHOmayGrwoZRqL/Ktqp9v31
eQPpGQbTfLNDAkzlFXtfkpTZPzHOW5BuzauNIUniI2XsqfdBJ83ibOtAp7bObBOH7TEBGazKkKkB
pWyM63BX7UDO5eIuVN09N23TtYylFB6hAchyO2847vpQi2/3nM/ILjrigbsYhQv2wCflsP75Acd9
Lo28uh6JMoulFE6FoJzE3SeZLaAkTkuKOXZ6MDF2kT2LgnBBPqrcupL7UCWi0tGhMvPqnZlM3eUn
oY0zoY1hPxyW9RVS36wREpcsZTr7wYLdSaFwg0DoXd4oV2iYCOHKYOlzDcmQs7yqX66gkU8vilD+
UINkggHfhEwEwSRwVNx7AjwvtN5qszL566KavsFDvDdTU2plhDBVZT/IKkv1YrHyNS18PfpWpIIP
CeGukA3tO1tvSStRUb2QqlfWTEwd+oDJumoDORoQJizQSgbuebip5gl7xn6iPB7ov/ywDVQKcdoe
tiNGakKfY1mRi0T+KGIO63hwzMou79zLcVzLVmAWIgfXUPAB4bE7loExyaKHjq5Lk0/2ynIzjaYD
x5t/c61f2nad/arYLIniNLqfedy1IxNb1i7Vm3qIxmwFIz9sqUyJyZk4epVodXbItXUuC6oLpe0G
5OqPm6Ag5K9XXrh4Epk7Z2Ejlsuzm9QDcrt3phHp/BXDWp+y7UiwuHsxmJYGUwNl41F5rB+q/wxW
/NLwZoorMzi/ZKNuf8zEjlgbn/+vWnpl9Z9Zp9oJL78HPQ2wLWc2XriidXAmu4xKAtoWCJgBiRyJ
kotSFuLHTCvToL7PB5HzvDxdeWQo1sCmgacH9K9aQpvzEg4olFgu+jF9zmLgHtkTz4hwuRv4+UB8
5wkGvNL2yqBn355nKwBXHXltjMGbcsR5UnSocL5H13wTsLVUrStV20O+lBxRUEDaOb989kMZt01N
dX6NYDnr5GTXEIDKxHNmcfVuqw53PowioZlXyGUSdByhvLiY4wpKc7gLjdBHStZRqDkDrq/0Wc5M
JIrJInOy7PeTDaF9K7J1liFqNwQkeR9zg5p1x5+9bOQvsj6MaQRojUK7OkythOz97dTwG+UoUKLX
i2cuiXsXjM1g+6bWLMDrddLmotgtONNDv/p1qLLXFCDMjR+H162VEVL86/4NpXGdP+7CEK9FTVlI
fWEJho8LCxqKnFR9Ov0k7Ds0TdFHkvtxm9Ietr82mG4bRyilL0EpMlYAnumwJs6X9sJF0shzEeji
T/B4i0cXSuMqHDcz3MHrXa/afoEyr6/ZQkYZiAKEcB1CyRCdNdkKLzNGh+VReAGVTqpcIspiJXeo
nmu1TEkEX0BenA9gyT0eXXGiD2jlzQzs0I4xCMgAADVXKbxwNbYn9hMgZfz3+AjTt0OU8epJVXYz
ZNVbvr3KumfOFMsj3KEqIqRzAqLEzbmbw2piiACb+tJiyfwLoLrV8MEg8L3Md7cNPCL4Z4o3bV5H
c9D5X8ljY6iOCnamLFyip5mpc5Zw/HYb6DLJMFiaJYE6O8hUEkKN5UuqL6z/IVz20mxZjBfiQuhH
wdEVLnzWrDgFHaHO3Etn/qwwniYu7Xdew9zIIWIn7mzyXCkuPmxQF1W0Mp8ca2/PMwaNZn3S+S/a
oS6mcOok24WJ13cmKAkjqFWKR/DVGBi6QEdU7M7LTM2jiFBRmZ/DaSyO43Uj4hAM2IA45mydWWh5
BFGvBEbW7VgNxg1KtsSFCE+IR0G/ZA4COwjF2OznBizRIXdnmNPIcL9Ec90Dclc3caZ3ET01RNuL
080ywecF+QMb918om4r4lmTNtlCgvO+YZd4G9hpxml3jINS/SXJAMYIt+Vuf4KunWfrrgs30jkng
S0QMDL0dOIuZUeAbp/8wxhjazyMhYjIAATqjirGIAWkNPoRRP5XOepBxyfLgk4wbFo+k5fQQEUHM
fqEB/QNZ5IhER6jx6TrXSm8wQJiisNJQKsZiDCCHL3sTHllDaYrXljCCPhqd+L7Fk6/GQgJB7ebx
HWTg2oJeT1LIfoSAw+6uIQGV0XBwUPhOdEaZ+3vSbNN/iwa5l9h+Ur70iTV3C9oF0AvoCezIiW/x
tY99yv9a2B8x35kas+GjCPWpZqeyul4D2DixMMTMxHmmRInVfVGeLKZ62MO5jrd1kP/HDIDqLjfS
pBKanuLygT8dp8H5yaYlX6UePLDs320Sdf9hTjCVqo8SpCWfAkqLLPZFH5UhTWdZYT34GMAUAs0O
dX3ljlHddigPOkXkMwzJOmN4cKF1Orp+romewqgegYgeT+Goo1e+jex/3LtJECIq++CZOm5kiY1R
in+DC8ZsDCzUOwU8qJOUHLr1W2Johy4Ly+fmpWZKCe8b7uk47SobZd5fY/V/mz7jxaEXHlmnkVJz
aMHAerIKGpAWkgrMisxEj8Hh7CC1+SEOoUBfT3IeLz+OYj01vfUNFADVJvAKUMpP02faiU6XBUUp
BPAtIDGlSy4SRF7Qhh59FSI5o+R6CSvj1sOyrYF7aExPtaG51y56BwcZJ6h+MVpusPiPgliqPlZt
n13a4eUrVSKU+TbiYUtptMqWHfu1fs152OaQjIvljh47IGOyZjV9QRUwldXAGnfA2r0N6L9hiHDi
wcYMxyUYeWfFgWZdse9plCvgUrdjScVMYfh1+qc1Lz+8ZjY0z0aHToXHXiPtqGCj++x6hq0/LQzG
WNoXJz9VYJdTLi3wjAHEEzkJPNtw0bjdQ50C4dnzTn7Qu9tTZgxO2BbvcQ5zW+QxHtye1dNv4Kd+
mFAuo9fHnir0fcQvdf3HFQDFAzqcfI+rRcYGNSi93eD9ACatPLhTYHb0kYKCEpHAZ3Bbr6sitTFU
n1HxoDKIFgBKqQfPyoY2cv1OfqxYfdTV274nYyxmVUdu4p8rvbxoqXl4wsbPq+TzgucQRg5XYyIG
O9eZHwqYDpDjRQBq0hf54E03gs4Skk2xq7ff6s/8hWk8BKj5kVWuzeEMAQ76Cz7La1ArnpiKu1Ii
3kAr3evbmTypHiho9S22lOcLoGeP1i1Lg9UDOPAo89mIRTrKJSHquwkZMXA0M0aHPaVE9MwosVq/
0ZIh1cJZi9BE0jhgDSHFJ39SBcmjAcnlC59JM+naoqGf9RvCD8N206whjomB7v6U0Cfhzx1ozL0R
ovhIR+QFZ6mJn7VvHH7pIo36ncwe6Yr8U6I5YV3g+NWjPoIXaOwhCO6CqWkTbUC5XtxeX+SGoLOi
n4z96HEf4aUrsUumXO6bUVUALhJH2Zf+MqxHCdJ5rGH9n19vYSXoHv9rwQ1i4ELwjwcJ3Q72kwli
bZBIwKSlUqUgat6M3yk5qc69yVr5Husd1E5uyrvdxw6Fw3RbRYcU+dHW1KlTQGlD1Qu4dMXDRiDm
mxgKgj3zBJ2oTG4ZmC5R/QjzBqcrfO0ctgrtxA6iKNbOhfdDxUhFJ+itpLR7QA4UB5xTvAXqWYDJ
5s0X/YY9hL/XzH1YVeYM7trdvnxCbzYPdYOrI/cOrvQlzZ71gCTXgtshUhkoxkM6G8/lOaowxX0V
nnQAdnuuhhpOWL7BTzTwhylRvzuMGF52apqlTroAB7eruliDUeLmWDG4VZLGXCPIv1j/LGOpjPDY
zQ9orz5NFoLKKoHU3xRT5NTGviQTxDY4BJjU7TSIOncbeWvYlX3qTom+qu/C0sjKlFmMUPVOAS4h
ejCireabaFxhGdIaGVdz2oyZNPmOoIPf0WInStBiK4IP6FkC/UFI70N4lcitbtY64r+4Fqqv6wOZ
R+6IUyLw+uvApylvBf1UKv0nnumfK4V+uCpe51P7ea0k722ukrb20/W5Z8rVD+6PFfPyelQUij8r
Jujd+CmyP8Ec0dBUftSFJhPXAufm4DpHd6VeAQTayNB3gvnSq+9cPlOF0sJ7B1m2nGjwMCm1TZCi
oRUK4phRvYg/QYtrhVBW3w4Vd3bIj0vZJ1ngcNysNVa9Zv6hAfh8Ke1i5UEWJOsq0HruPVJ9HoIb
kboF+8u7Pi2iMd6hdd8QlMQ2Rj14bLWTc9PRp979SAkGPaxAYNiqKSKkUP1vPgCZqqLghNim6uud
t3zuUigxylMf4haGtmPn2Bnjv2W9rr7MuVitfFricoDcCUWPXC6PXbTfrML2Cpw6vhhCid75ayGH
HvEpJvDziYRfITBhEM8KadMZ176evc/2D5EHUd1DfZAHiwfFIaRHIgGgK4kTtkTSHuzzf6l8p06H
Q7WJ0FaAkx3O08PZA4S4VSP1qZz9NZibMndupUlrF/CSnel6/R1nO04qjzX+2LoGIJRhLGPY84OC
FYOWW30JxvS+EiiqcqtawBP6CBOyo6mC11AbkPmVJVxez8Q8AwbvF8Ch2W9D8DKDlqXsqn4mQEHW
D8fPYgM3B7BQrK9Yex3iRjc0480atIM9TvhlkdvXNlYWYWdFsJDSiaNV0YJ09oI9twAYG+n7608m
UALhQILspsm5c6bWtN/MrEM8XdwJ40kpg6yroDL/LS0vRn699IfPYdC1kacHDXFvLHw/1B4a9C/T
DkvNjKBhnmn9B/be/acaNPi5XxUqw4tP3LS93PFJqEqnm3c6rpd0Y3kwFtwc6ZIx+u156AMEhV26
VO0nJtMpYQwNo2r0EMfyBNKnhly5e5M8or9L+3Rnfdkv4AyHuHMzi6Hg4qdkoYCdYJqDuYan9gqg
glBqMyXOMRTbqnjG8oSSAH5xqQys3Bu1qHaPsI5Vntf5cMtdK8zMNtddKGhxuvcbhp46xvDv0hTI
MDN0dUnmILHEeDHhCh/1VB+eijFWLdiQvgh5I0kuksJ7a5SPEjV1J3NFeGn22Xd2xAXa4i5PZOMv
BflPe7xO9RC+CBSWZ2+4QpvVYyQM5IbVgziQ17TWeyKyHe11wOOxqRjFkz1LbyDaFSecWJk37O6x
OF8rYOrCdq4nbRVwa+PuWAkz26f3Pb6THwZh5NMe7M2ws7B/MQG9l3D1YWAYpMt1EF0va1WwDj2a
d/QvPLAqsvjOzWSWs8M4S3x8jMByNfAxPkm60d7Nk/icGhHKUe1NDvDPtMGTUBuXiesX1SNBwfBZ
A8iPDJ6+m+jM40K9ON2CVVFhxwpCt6Y6bVq9MMs7N5qie3S5K4V5hNihrEoCEBQ8r7EI6z6S7L2m
trGNfBXWtRd72CIr8174Om6sHu7x0bVJxq+xKbW60wca2LakcDMcf+uD8mrWnNeO61Qhb7kI8qeA
fr9+4KldXUjGnc88dFvAxROIqdp/b592LARVtscKs6A+sAxbJSHGHd84RU277pW2T1J3qI0wjitc
Ez7d5g62LdP6+ZQfHXQTnLiBjM5EkWy2EJiPMfZ9gZsoOIUmVRSVoHLuiVdcAL137klH+zoKPmDd
ZXZocvZ1GO5lYOZJnvZlxrdmal1Q4GsZOkKL5kV6i7cGENnXrcZxb9qoEN2G7tMLE0jKdGymPnPs
UXgsIlBRcXFVlp/SyQzRI94XvfQYDbQ3necqht5rpVuGbd39ESTJHY0k9qR4/+CQUmwgPYXqSZhs
jNgcuWt7hIIeAiViqqWM8ZoaSN0jacOmcYaPpo85APOIucZYPJo4koOgui3ST9DFKuQRGQwIc625
ruzsfwRBYq65jmGG38srBVnNnlHOpWefxB/9o24tIoC1TYb+71vWlbcG5/FzJMW6blWhmV5JvHhP
G4t+3EPbFyLz3TOq+VKDfL2Nhf6VyXs4v6wgG3xrp8LaX6+Ay2lVG65Ll2gOLmoWaSOQC+h/HAnO
hjNWACuXA79pajjZ8s//P7/ANjRhlmH5Tx7EUGmrgxgi7rWX3wC7hiD4j+jAIxnQgp6XFSVuX6y3
LNuLLfKIl4mtskk0jsK98MO3uXRDhZ7ift/k2PCYTt0nC/wkWSehe+N/gw50OQpwho0UTHnwLZyt
99Ir1EMiFDoHcM6/ITYEOBmezLDJEhEy6Rlkg3udilVII5XeYEnQnUX4m2l+tVDs/OI3ybb07GIn
yVP/RG0ZmY+rm4NpvHG5DnMsOOUaF6Sfe3erBI7ZAsg7pwZeFALJi4jc1AN/ipalS+uzHWQClRCM
j5oe68vo3QVJHig+ahm/7lY3mJ1WgLyEVbKN2WWaQZHiMX1lD/h8/CCbh+yyJHYT0RPomFFav7uP
C6u64iKpFSGUdWfdZzDue5RgIFeyLSmNE/O3tR/KD3GkkSXtw+71e10KLM0j7Fmw7Q7+gBMF24sV
TMmUhHfGu18qJtL8ca9DnU3WqBgf84+cw1csAGAf2CdE+AIZYXmkdytcShdB/hFM5rMIxVhBXoMU
kkqS8EoPYXBUTgCjWZs+1ObEQREsW+YmBYYO+6U4jlAGEmjtCr6fGkFTl703TedJLK6uPk3QWFEo
MnP7vcdBByjBwGtfk/+Yfo5L5gvjRRkjogS2n0I1NolZ7DA1NNPPMdzlQUL3NMBe2sV0AnJN3rNy
C/BSOVxxryqt7lWoA2eAqvI/bCxzyCumMxr7JjtLsCI7Cvoj4OZ+Ao+FpDTNJ3RTx8rQnGbNyu3J
1ITw5gFCUs8N4DDOGYhUEHDtLpti6K0hRiLw2pT4/FEgYNVW0JCPdFjg1VaqrUD8/kbyTgDtWfHf
qw7WuSK9WlpBRR6RwkygY0YIcsY8Lhbqak4RF9M7X5iPsm2kXdBufBU2zC7NolcdAPqZDm84lvHL
dM8tMcoKon08zqbIrGfd+v+Da5qWCMcH4LHyQukr8Egyq9nDTo7CX5XA4capXhifClruXqeDiUzD
0BYwgGsQeQNM/W1AhR5C0uSO57m8UmI2V7XEgN0j6tyq7WrH3n8WomPtRSkb5DC36XdGMDkOddl2
K89yJRjZQoEh19zqnliwPVdCYXsiRdXJ167pGZZaQ/vxvxfFPGgWhgDFlZW7tUiN1TdIC5UFEyXq
ZKDg1enkhYNe4OX2Cf+LhLKsBlnc37NyNEP9wDSfk6adSvT7BQ1rcUtAUDHvnkF1YuCmpdBV4zsx
OSC+RWH6qXSlP3IaO2bAiaVx8H+XIbX8Udbc2Yij69axHmq+ajuMJPlwngtHsWNSViVASqzMYK7u
xNf9C700EGKxzq0Iy0UPjAaUa0S4s5gvLvbCqTo5SF5MhRlTiobhIXljrx+WAmvRF/7FQ+TSLfTK
AhWH3NCp6JWDfuRybXBVbH53fPKz9PwlTtPXGb7fR1sgehV3yyTR9szgP5QnZrq8hluuJFKhRCvM
O5dSGAre/WmYa0LalVHIXgbELAVYhSnq47dg1tRhc7tnI2sUfOqjZtr95zuLhe6G/WYL5B8egxZN
duzErrBpiYTOBlfHSELE9D3zsE5A7B4CFJEf5bvsI52yByYuvDXxC3/Omv9sOb6hgzLgd71xVPw4
3faMk6DTCM/RH1vER+w2h1gI8BvAEiJsXGtEayzuiLGeqLlpj1Oc3HonaRM3v6jTs/xzUTngrlXc
+szl+xHjVJ/ij0zldsPg6X7glxd20JbHxWrMwyL938IMbzPynhpQl6nSFcdjl/ZLyhLN/lbG5C7N
EL/nl7xXb4wRew7DqEnePITcJ4rJv0sNTNRQZmPu5TCaMiltjdp5LBU5lVSvhLNXf+HJkqnyLBNw
uYcNQSaAplADJnOWaOv3vJ1sGSUYvIv0faDzaEsyZL1r6wL+2f6YtyczqV2dYOgn+JlTOlflNjk/
FAgSdJlzwO1lFxyfU7UWE6SJjsKE3fpnTQ00tSLjv5qL4/mOtNctyv9ypbx/tl7nUh0A59d7HtaE
NAQRJwVSDfeA182p1elcuC+rTJ6tAbrJz2vb75xr/eLXVDT6RA0HB8/+NlUAG5CGha5So49Q4Y5A
RZ8vvdYwNcocCY4FTnf6jeNzUJueWq+QkPZAwCdhT/9eIjH8WdZ5Yex/VhEXLTXE8p2L7IeGU45K
1ANGwVDXJBKrMM23nhhYACxwFrz3SRc8pamXSKVY6RJA43xvqT3RuMPUuZkfCevddk0lXNMJv3ci
X1jew88mFliBZaH9RVbepv5070L5dAfk5+PQG1718rOCHTZrxfxqsHoswewPcoDECfbiMWAkTcn5
uePkZlkkzmT5gjUzRTg9sM86rh5TPOkskeYR8PkMZ4FPjC66+JtnWwMAyEQUNpuAdDWkPIWF/WNy
0uVu4yQms2+1GZpsRrT4lBtL22X6T0yfxMg248KlFsMnidTVfKc4oVpy7MdLyMWAxuZvMeL2R/7J
ZxGWMBkUgqsOEmaFTEx35isuewzt0yvSfZPY5CDRa64GV5S6Hng/OZJo9IsylChXlxmz7lNYCl3a
GAHLKj0PqwXAjtrqviIoi3w7a083YCggAh3Nikb2oDtSgbH2Y3ERONknP8cQRqf9U2hPYOgW5N8t
o21feF1vRgw7r2eWJqbQKtdF3VIkwoiE3HEYywzQdq95uvakNml5D6qV+NO9mQ3XDhyrAPnUxM/4
k7Me9R0e/LP8mLg9f064Iu8PoMWlGxWXR8dQg5nMjLe3E0Lx5i4Gi4IwItAkglT75uFmX50/U5De
QUFp7CNHw37PIBjdl7HmQhkgHy+t86gw1jlngSlEF67WHoHLgJw5ArQdeBCtmkulMGhCDFvOFpMC
Ps9o/FyckICfuiJc5Vw6O4Hg6lg9l1Bjj30Gq3nIxAAfaiRcWJ4QhZNFE5pQuwBJ2r4HCYjSuZYU
YjD8jS6D+PAg1yZQsBZRn0NwytJVPpc2U4BS9SqS7OdR/2nulDB0I4rzicoNJSIw4mPMcjs+w7PF
QdhBjb2fe1H/4n1PGJ+YFTcKs8E89Q+40pjJtKvJdXbWGmi9TBW+0uezqf4M3RuuD2RiTz6hWq03
s480uK+o1q/4bTXWJvba3diyxXIgmucEY5KrqMT+O+zp6YCHt3+oG46AfkGjipU4xKxs3/VGnIG8
EwSwF4ig6c2gpSSsEAu1tqcK6hxZMKBN12FxxsIt2jgo7iHANkrhbT54YsnFxhIrLOIklNcf7iEd
uJrXzBawCxKl5HAQcHf05Q5rTodDjEHYmza4RLNdeIS6k7GW6B7C2Em/YWe0HgBSxCd8Je3lCciV
jPTiSpPTcE1eiPmX8maMWlAbXtVck12wMABYOyHJy++MFRfpAkeFQuGXJByxPlC8EuX9S9VtVGG5
1F8M9lxltqx1n+nzohxTxM1leVCgBEV5JTZplWTd/hHdZ3b/fId8aLsFZ427dH4DpUBlb0CexvsT
Rm0FghgOOhHgN0dSJmFFjR/vf4mvBSuhwIB3rPaSk/KhDXIsf9vJvpJO3squDviH4CVDpxNTX+ET
GtsVsf7X2PtevOGVCWJOIsyl8rZWKD+jmjL0Wvj5T9VkLBWxXnudccjX5MHR83pSQoPi3EsqRv0s
ym2WyYDD4QJ2ZHEm7Gn5wm6umgUKvirfVyKG3zhF2UMg2oqXliXVfLXXpcbhHd1Zxy3BevRMQuJW
09DCSVV/u9PxsLtBOlO6YtPnQQKiyCdY2qwf9K021zlmFklXECW31zuU/7fU4FeYKhedOeY6LlKa
yoKWQYCLxZKZ9L1DYpXK7YLIoXvFdFyuL9yt62HZ0Pcxc1gVbiHbbC9A32MSvxakqpkV0T0OZUh5
qc8a8ON+SlUdsEuMlRKG/coX4VTPNHKxOcCPtNKa3n9ur7Xo3ZvpQiu+nObDTHfPd5ufzGUgDTDq
7t+hbN6fZK4zj8vJN5Dt1qnruIrFQAfLRkSE684T38lsDIh3shX1U/e+BNTwII3qP1okKEnxLKBD
Oqb9BySlOekn+7il20U46i5el6rZxTdOOeW5T05K5wc7zmQPMxQZpXHI5bQBqGGu6KtW96weqwFD
6f2XRqlE/K5h6+OOGuL3MPZEbzZDkN24sv9AgBf7fIpRWLER2B+Icxc/eWGMQ0KpfFLD+8yl+0re
eLl6uLAa+AKbacFxCIjuaIR1x7qz9t614zknCBnG//AuIxIgaw55ZLeK721oRUTbHZK4dZEphGME
DGmyAde2A6C4a0dWxS2G85a6+cc/s64IGNbBSer6XKucVhryBMyUupOh7TyTSgJdCSXdJRCGFDvl
ZN24/S/Mp3r42d3EUiAKsaqGdBjGrdwqFbiTx9C5/JSij6fo8cw9FmJ3pZcbEldQATYJaIl+pPrS
TLxRuDCfsm2WdlHfQxTmXrdYaz2FfMxP/KQbkASMCZQZVadIopGj53cMrrP4h/jPh+y354yR/aso
DRVB+L6FfmWv1oeJsSpqRMBDETYkPDXlWJOx4MW2biDVAU6SZsBXAqYl6nVk8tT6ffO7HN2TSyTX
LBPxCHIZeGmmquafOe486MTyBWqj/IOaPKp/xJItHzy242BOyqUwG9a4kVt8rdYP0QjtGo42WuPd
1VfV9tZ5pehfVoqYvwggvG6ykMIF/2knA6/yzSgGFnUgPANcccVXl6OLxcCmH5I/fNu08NAgA38I
XLD3tV7kO1b0YJlp3w76MbYl/URg3OBaC/J7esSiry3nin9Ck/o6ZrYbIqt750HdDGe/zfl4nCUA
ibnZx9HN0OZxZP2yauURTspHJIuiKdWwm6M5cItM6j+5QuSkmdlzHopq4rSgqVWGD47ve7u0jqLt
1eGRfjuZ9X3pv1y87s/K/REaByYGWok8v7ZsaIwJrGaZ5lgzPQNSi29aFCDuDx0hxVFpc5nqP4H9
9AnGU9nqE3LKIT5OQQ9FTPQ2d3gw+1t9t392QLKcaKa5uALKcJvUPWw5tofDzzzK/xkUEJPoElDq
aMwl2i+xYTzyQldJAYwxEYrPWmYsURkBbRcao4oRPbk/xWX5AhYmrn8xnaoSjl8/AZN2lENZwn/z
ZQfHQy/sXAqN59l6fQpYe/zdj6po6sceLqi7XcaZMxYOIDOLJatnmWd7whlVjyA33qm97ieRqStN
NnQgz+HhCQWddq9PQc6YA6nWxfgATWR/HY1KQqkuYPevEVLl9ESRp9Zm5e/rRLsmt9ikTrqxhcaM
hKMQnsRvnSkoIYbK6S9wWSt7rEANzdhuYESPk6Iub5QxlIhi1afFxFNRz/onny2H2cPhvQTgRule
TfQjkKYhw+GM/QFF5H+uF3d9DW12gnrosWOIxFJZOsyOchpx8WoElkT9TlVWrSGvHi2V4MuKHWfO
WJyOdABkQkSgYpjj+/cuX3vo+oMGYFYgufMziio+PfXsGmskKiHYqWgo8uDG37ob2i4WC3xhEZYK
oECUC8FjX9X4HVv2kfJIsKhntU5XDilv/GaNmDnxdl57YpUHYmq4aY3UCIvLc9z5qsKsTMGyVmxh
YYbV7ue4SbglhGiK6rsksm1vUUm63nz2ZRhPG7Cc3L2ic68KRkq2RNH0ClYoZuxD14jAkbOgPLro
JcblQ5ku48KMBGmnaazhr6MZnBHvoqHrv4BwEhm6b2Tn/Fu6od9sH27eKaObNnor/iiJ421HiWUR
jxUm1FSaaarXCk2DtpsFoU9w8SnKz96ay8dgFey3dbIM6kEj/oGJEtpYfZqdChOZbHVXuk7FyNM4
GKmi0ai/GEoMmTDx+zRVJYsFhIfpNKRHJd+dmzW6PWltxbqpylhPbp3eKfqah4jFJ15mfNy9qJVF
fs1LmRdEMY+rQoUelTP1raG8r4odBZEMQnoZM4yTqJWa9aNzpz0K1sQaH6iiAMjHKjSTQXY07aOe
OTuAYjFJmD+AHdY1FczGHk+HnTkBPS8z16CCu7624TSGw3fP1/uuH9887LK0iFE5V4fY9RQyHQSR
JNNCScJunV/oWDCk0Ni/nHvxBgv+laUaxiJ6t1oamz4fUB7K47ShQUAunCXdOHNqK2w51OP/Xjfm
k0qgeE+IORyKNFdWZtYuoSZ2t4lAtRCSaKPaU/NHpaCbk7q8Z4Sq+5yCRkxK2PNu8Q/bXbaVEHZ2
xxFU8NxbrNesMchIgS4aVRxSAvNPYselgV6yNn8c6OqLeO5EWhLwDThBzgZPqJdOYU9oZIsZD8pI
v8zg/uPrXfV8j+G/LBgf9GjnN4V5d9xn1nlpW1J2lTfoNvCQysZpJo3n9iyc6qPIVN+VGj/yc9J0
xAxbu0ekM2vZS71v1j4ZewuzN4YI/oycYQBdODEI2ikTq4AghSUBwPOr/aA+JsmYKdOUeAgtWvZU
XYBNweJ3aIqD48tt4pxKXJlUZlgB0VKVZrDeZT4GFjCL2s6eXJ6cbhWoKOfbVF5JZRBNFfXBlAyo
DzHQNyaAo7KC9QnDXolai3m2f8qemKafNE7nPMJUf34sRoiLCO2EmohAnxzoocu6mYNXjVgFXsL8
grseZ7QvJx4GRyD6BMvsXBuWqMiONbYgpZ1IF6GkmKoGqmLjxTemhee9qKTv18keIsX7traDGfHw
UBhQ07U4n7y7yEfG6dQXBuRBjyD/SBe49Z/wYUCUkhXF2r/VNbGB/k0rBpXWP2STMozMv6s5VWF5
B1VgA0Pv/mszL7YOBMWGgD9VZWhvx8tLdg4bnYsx7VvGNrV/qhlUEmxtHvg1ErgxiYwZ2wIH/rcq
TAEJN0HxU2MOwyEkitt+t07sf5ttcdUy3SXAYbfwz4u3qEXbkcJ2H+Cn2s3Nf3P2/IBMzRgpLEQB
SX4MIjlfyLuuCIX2SDYL5797tp1haGIBp/aeeMmrc6pOcTCNnFg75BDQrMqWkM8PE04LiTmloTu5
eMNrTIYujGLcO1DPh06SvD8XzXzj879kZ+ZtxIhs2+GH4gwo5r2voNNOjMzVD1vmnzPtC4xLCAVM
CSIi7ZnsVhHnucZgfkFvaisukmQFAiKHEJaB3Nj+lg7yofwWacDrxd4mZnFskwWQsfq4yvlEp0PR
zJaNJ0ihbx6Np5Mu4X7GsmxMqINNovgGwsprn7oxyZmXjyK6Wc+3+lewb0e9bqyZ3itStdafj6yJ
x9EJXkWPFbS5VScZ/AyBQrOZLmiL2KvVIXSKhFJhSlvD7bVECDYD8vrNklY1tQM3MEJ0ub2DSoYN
q1BZospDLlEW03J1Kdi8/YLVFrBNC0vD5ESGMr/8/EduFPoVaglnEmwI1tyAJZmvBQL4pEjyNm6A
VPypDKsi8zWWAtgX0cNSV+VQbyXWydRNjjyDn4HRCPy9N5Sw27pFbPINtCIF7ZQ2BWae0VseF+1K
TkTZgI2Y+beUa6JnyyA93bJSrZkO3cu+WpWoIq/aWX1zudUrS6MktjpNA/Oj8nxiCnXRu35r++JX
pYrjwBac9T5D4u+6zf8JuGmn9N6gNaEZbJ2oLFmxsLSeZTPlMCb0vPD5y4b85RIcUT0Eb6NYYC1O
E4dJwTmygIbajRRfbiu0B3bAdoZqyeO2jKiR8Pa+szVMcS4IiCJGjAxf3aPXKVeI0fxwYjB3sw69
14n6XRVbIIrBn5npzQw/YRKnbTCQAEKonhRxxKPMuaskBJY4MrTeZ+BWSSuNeSs491zn3PEr4nT6
tgZgqL2lWFgY80yYUU6GzOQx305+ilMNOAW+kxkvIwTG0TFMG5reGsJlV9xwR0X7QKXUg2cj+zYq
dxSp1m/7OG0VkP6YhI8WU5oVF2GSzzNgoou4jOmmfJeLTtXXtxtq6CvFV02F2P701PDnlz250zxE
IlPyAuH8lSc5rRrco+kDotmRr5Lt0WpTv+7MxUteWXao3L5djrUopViHbDNLQZXsVxJEqI61cJ1S
Q/W/PNL6BFJh5gTp3rOGsL0CZU4BNV/HhjkxlQJzeijzXe6UxqV1M5tLu62RhkPGefvicD46SyMI
1NiH5vsQkdiASB4MtfaJiLw7HYtaxlIVAn2vFFFm7gJ8THEv17Mg2Cx1+nVfAlcLIYGyyPiV2Xdi
IsXh8O1R8UsxlEMnODo/nVsYePIXxJeokc0VNjLowkdA3foehl8s4i1MvdHnjW2ZDHervvEg/JMP
OtmwkK9gEay3hm21+6wxQlSQB/hpwK41//ls9ud9zgW+QS2f16iHEAO19jB6y2eZmGnrglydzXnK
AyZflLr7CsmnSJrlE7LKjs6M5A8Jwr7MkjwXinsRp0ei2ckK8b57WUoUqAmj9VLO9Hc=
`protect end_protected
