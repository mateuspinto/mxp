`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
Im3YJdlsXYmCT6EuGcyrzpC39RjTbm3HTYMpjmW49rILQ617rM57FWP8i+BHVNU8BZdp50VWH0+Y
H8FL+kpL8HtMc98GeqBCdiRrOyBugR7wstXpRHTr24ISOCWRGrBw1G0/dKhMg/FJZSiknOcgrAtR
fQ7xCi6cTJi2aOo3VVMi6wx7LyEESuqv7kuNEYHDL7/DgYcjjGsun8xfv/LKHAtgpR/YKW+Ci4wB
nt+BTUWqNEO2TNUsml88Qzz5cAXhoiw2lcPZwRyMe4MonfefxokXXLyhOsFcS2EMlapov1KnzhoG
iofjH/JoqsxJp/qUUycaABgI9/YvzjUS6o5cuNCIBC72YGY+SsI0DvPAMD6zsltYQfVjJ07vl0Kl
R+NKrYkxjVBqZsgUoFWwMPllnEh339/qSY+2mbVm9OsCDSSc9jbCNDWQfw7rerHPMUQNV8wuOKRG
TBVVC+QP5c3kWG3jLdVLl94tMTpMmak6/tnWnshNtR0sjSPFjNNJFJgr8ZzqN4Cxxws73gyexgo3
VNIiaT+96qmvuTMkHGjox9d57ZaE3YfczoV4FrsNOJKlxqHAJpemNyjTTWwwH6kZIPekbZ8SxC0y
IX4BHbc3fqR2Sus1qKcWmbWMQFjGAw5oZbEXxTejqb3VmERns/fq+c1lhAnR5/MlOZ0WxO+F9s32
yy6icut6zSFY0pc0oN7s33GrONEgmia68j/34nKWPO1sfOnIdmrSUPyQUSNa42AeynmYetCF9KnE
ZHJ1TvKHaRoISqa5pzvR15cmLaES6xmN1hJOLH4STN7oLf8Itt0qd+A6msAUVLR2b8jdVD7OX0+Y
/AGHylDBFc0KtUIIDRc6XRnv4Qa++fMiY9nnpsCoq76cLsZLufEDxP4otSOdzYtQqD2GupCeC46y
6/0HEtlylpbFZaTNOHssi2bnfrxSPT+z9gmkswemnJYzyduiz6t20Q1DkZ+dwCu7byEAzplk5005
/YWFwDbEZDq90LdXy2vgGBNJLxM6JHgPBdmHR0EEZ0GlmURxkGCn1zkgjoLzjSnb6TmhYWxhR84+
0evIBPv4og05QpbID71CL5pcCRRasVN5o5n1A4+vlApC/Uy01GDpx0MZcPYJUOb82MtTSItqGSvO
hZD6wG+SC4xE0Y9+bySgq1xYKCwNV0qNDSfdG0eA9Nc+Qyf/g6MGB/Ve9Zv8RDBX3jyR49/ihoPn
5HL1IyHWlUvB3ay0mxJy93k6B97D4EXJRpOrAatWiMKLWtWF5TRkP0Wp1sM/vBqOiDfZXI/BSsti
D9YyOq1ss+8y8v7C+5sX1/fPv2dEuQp+k8BVJO9JZu0tdba/3S74hWYyik60a6Vi2yQOSo8/6XSg
W7+btz/OqkhqtqJ0Ho2AIkrj8AUcg0b3f0ovoYkvoGXGb+uIhfb8ehyH4i59AvleN3Tn3uF4hdM7
3/vmu/3Gd96hE/2ZtuuxaBCegTJ/RUb++qqOe8aBeulJk39co6b3mCUPPZAB8blhoQnqMrx09pr2
xdQ7DbQIzaNw2YI9CbMAhr3/luGSLokUMgDA3Tk4ZZGZouMZS7oIaf7jpAIRXAdgBc6sdw9N3tDY
m2CAi85o59ORg4zTiSTgvVnwkdqLtJL9OUeIvyyIqlB7nEzp92FOPj8FlUt2dM7x/Uib+2BIzE27
aZBZfe28qeLLBe1u+YBVYLdlEsrcdySC/iMOUxfa8ID7ainDuSSEaUDzI4t+q2Gbt2A4XIPQuH+g
d9IV5SOzHdx14S/r51D2IySHY0E7cdtHIy3fnnbdnByiGfcZMTVHkBfWoWChFQfxrZdwnMrnhufZ
BEllXZI/gxWyyz2KMaVhAGUc1oXZe+X3fLX1CURkz/LldKFoL5gijmY1Gz+bzNCdm5/02fMsCPJ2
NAd0DrnKlwaa3oUlBelO7A1dD2my0E+IgdWdlmhihr3c26C231l6s6CicMML/KqH8IPXyM3qzFKG
10qxgz9bDuFLYKDnifAgkDv9tO7548TyELRksmzljIKpTnnmwQtDoe5Mf9p/34Du0l1lsmcWSPRy
PbvALzhhInCW6gXc8lGP5Q/liSOm6wI0/PcmT6gGQeFo5XD94UnX2exHsVpU7qrNEbSUk7Kjno/g
+fokCo9/tKEBcbFBJ5FxQeJmfu+5x/soLW+CpHhT/ASYoTWAsFqAhs8QlqML+QKgOGplmpbT1aAW
JrKSp68Bmo+D2lZNtBmkWpNC4/wxhTLAwmHGNs6pcfHLJiedMTWrB8T2P7PMyMXKiaYJxnmHhcbw
p6NTcwzzitA7ee56hqypWXwKrLlnfF5fYsYb9oJTTFn4dwNY88syM2nl3BoSC2sjyn00Zr1kzmZB
JbnVGLFsMCydTtbBsT5+PDfNnsgwWUnE6uOlfYm1tq+DVqwYL21eohBO8k5vmturXXQ3a4nLzF8f
Zi1ScMlHj34Y3cS3cRyIVEulnq+qf13q6/wv/RxWv3WGEqqtC8i/d19tn73aWlQZKyIb1Q4kZVmE
QJxs4rvywjL5WXehcOeIVHzZPJ0D9FiWZPr5eu5lP4t0uQHLBOryMS9gp6Pst+R2B3u3TAw/pIyQ
f9tYA2ykEEZDpgor8f+Oq2+vWqMLp+MJ6hCGuk+Mjume30wu11V8X45uqCdAPPtMkwd5oLeE+GUT
3wDQX7TVIwlW6Xh6F4FONM4iCnPog3fTUCq2Qfs+s8EBH6RLC89ieaxt0s3vmaOdvMFt0rXimjGP
8BQt26AMBgv5ibM+sF3hoqfn3smd7Q/9t0o5MwrtV+RrkH2yrPvIn1x61HvJ6pfAaNZV/ikAb2vB
7putBNbg25AFGv1e3MCpdTy7ePtmlfpOSL6279UxLa6Ku9huI33kCRW56TTG7rlCQj42BBgFZPDL
arUfnZ1hy7+qYdWtT8/sSl7ke1Lh+CvHOk4mNCyot97J96iQC478upJ7vlmLX3gUVN8RFAqiyhHr
pT7eTSw11yrYuTfA/+Yaz1nyMKV44wbnxvYQOrPWNWbqElkBBP9ND6J2+PNwLlf888fQuH9YpATa
FweF/9x6/Y2Q+FEIeQK0lptz2OYCeLZE0sEm/VwvLCYbQ9kS3Oj+AgF80t6JNtrmjqBmBBihM1W0
aVI/uv84Fa4BdQW75SQ18fFSj96bFLA7AET3600am6ZuIjQEhsMHjulu4UJ1G+4lRRk4vwxz3gDf
71Lv7oZ3TOobxG/gx+sxBcb3bti7eXb5I3W6+oDrGqy1bBBNVglYal5rmX25gCWfgVp7DqEv6Aww
raDwJ/dFu0ncCStJ+cp0bBbwnUS0rEwkrYWD4cfw0u1okEeRluVD+G5nHtGE/cYTPekBVSp4Qhu3
G8MaUtN54yJciH50ZxM9igTvksrxuupXHcSyng6DwivzjpcXw1SeNyr7UGPzRQmj9rIwZYJ8lzWz
xC83X32PkC/xxYOFpnuYKYbDZgPUW+0aQJ1CI0pz5F99DsM2XyJf5ZgBSciUem34ImiLNXR8Mf4u
Jv0Hm+UGskR6XkWiHlJ9rFnM4Z9MIc3v2+5EEtx9mU/X5Cl/tq3ad6IxPL4o870b/ix429Mh63+7
fBel8tPIr52H2R9sdu0ZIzQJ/WcN2WIKkMBjKyD8mYSGNv3waqnNYDRLIfsnDHA0RWyxxT3ScCcO
6/UiT2CU5StHDzN9yz3Czaoro6pzpn0ykVNz+pw8J8Kw68+96qtQiBUClkUXireIKiG35GHlzgp9
ayNJnEkMyQPTBpFojoUmp/8gAh8eofVTSM+Ts7IF7vC6RGQEht+roywFkZaf2g5VsZ6peXvFPU+q
GfsQy1d32aEE/NCH+cMEPzrKXR+cTtV+IhWkqsXSmC4/PYNnBcHGbm1SwT0orF1A6cX8nVMXPBYk
fdl9nLJoYxGxlcdY9Kz7tfu31jDSrsdlG+Fwzyg/ok+43B75//3+ORHztKLxTakVDuYD4atbTgwu
qtoOqINUpXPyCRlwYYangSBEo35SJ/laKIXGqqzCIV3KzcVFjU9rGhyjemt9Ab2qUFuNw94ASVpO
+SxLIGjr2Ws3qvWIK6OmavUPoD7F5uys9JEn3JKvKxu3xmofeuL3jnYiCDH2Y376r6k4P0zBy5QR
fZnxMsIiPDXkLAdkKcF/wgYebGNwcDScbRy+gGPfhR6M0CEtWueL+RMlUlb8Pt6AVDFsw+L4W48D
NPaRNBitCHBL043gJmcgWGxzmkh1pzeTlAojWbyN1q+//GqfaelirrhTBUB53CDvZj+wa8LL8/aq
pspukSKBOf9d6py30vdxzbhFZyWv1M9zfC1eAVPQAnPGSHMJ7iHDdF/iCLvHp2XCqoyL6eSyotXb
HSY7txEsYXpeFCtOe/3i1Zkoc/9QBc+BK5ZWmxd87MqUSmcjjkjDL+jLtIz6Ec+ShseW+9t6/diC
7KR5+zkXxsqpA9quWSb/F7lxvm3gGpaGEORiFS5oAlzT3XMUzuIEgucNXvHgg2lIo+gmVE4cwQD8
nmsDAJFqwDRt2EwP7nkQF0wPxAvJOWAGLkz66H0ZyQxnH2ckAWJ12z9yiScCs7ZACsiOzML80b4Y
kD4wkHc7MamEm0tG2mY8WpxPw6dPp0kRiY/ePDOVvZzwLxfl6K8g6sh5PxYW9qZuvoGlnt3xu1lA
wzBEQ4wS5vzn6dW0oUkCWDEybEMRiK+tcf92JzCqCOWIfxkN+XNxQh9LNTd6w/MBUOoRt3ezlDJv
6Rc0oyhyaz9TclIJU3RQ4EUwwaMN8K53hEl7/huuNK47A0KdQGC6UV1cY9m8LJA6MypDro7odxWY
bXpH6aAloh0YAH3pVx1mcY8vCu1NqEZUPSLVIZeI9Q+7O0+MGNAXUtjkxQ/s/LXDN/R4zgSwtZra
buBRv05C3J98x00W1RSr84TxQu/Fn3bfuUyMBjWZQEiDuw0QYIqYs867bCkx+shXv64SDMgweWVv
q1IEqrhsn/UlWCoejlaJ42+8yTskF8IKV5WL8YoifdNYOY46ld7p2I47C6O8C+qUiFOK70iWQ1Wf
ohLpWWWRVUZgacFXn3fSX1EcKHEJYw1DJJhzc0OS2BbArLG7y4x+LIIFOmKoiRtfc+ViOsJQ91VX
ER4bgqjrRRFGAGgBV0m+FVJVwLtxoeT/gUa2kMIc85k/Ae9rrFgis8PBpzD6m4SPnHg8FHw/FOnL
ydBgOqb78ZDl/0b6Z9pxRM9i1fK/okEEWi0oPSo3Zg3KeL1v1bJCFMZSZ8vrX/EXxv3vgY5y5lUC
iV6p43vmZhl3j+aQe2VShsmMK03n+QS1HPdXy+Rzqv8xwfFm1LWHJzBx/f11szgNFtzItenqJ21f
uB4acSaylcgUYZEjEQKR0Kpui5KY26rqfai2CsSrCNta4tn3fMAqmqeE4vnWR86+/D4+LxGlYYwC
YzoY1kEtXq5nHwkgVD7Db53kguia3rsZz/NVXWYizfaFghvMSdtWPA2wO012hk5kKhdwtPDjkrDd
EcznIROch1cjRFH+ZhHwI5Se175UjmBpY93/3pAbZmzYk4ZWyDF9FMsppc6bmvnUwZIgprqtozVV
JGNiuM/ySGP8R9m4GfZk7iV0EvVgWwDgZZ8lCWGYeKrJo+1BA/CPPGasg1gdR/8nLpSt9NF9HzVl
GpuMPf6dkgGZPs0gO/zyK8VkaH6K8sv6XHvaZ01MgZhsVoGK9E/zTrwR61/xnvw+FxvNe5Ri7IKB
XfY5cK8Vuf3zHC6bUlwp2GuPBeO7CoT0exV1MzNJIgvXDW1jDWvbpH1zA7uPJMV83v9PSPXuyVk9
Mr5Z6c/VdbiZzqfswojJnwp8UueB+d3K2YxQSaV44Ee94eIIT5U0uj9H/1VU6dfOIH0pTy6Aehxz
IOSqD9v6PQYag6ijol5Tjjt4g8UmzJVr8k+Qm7GAEYxbWt0WYNND+kBO7FpsyvjoOOQsmVnXuLtj
nLVMa2mXFbOuVf/BXQRjq/6GtLISd108neTIXbJiP1R5eQMngTJznRMDyOqyHZliBDKcukNd2pjy
bb2mbSgy0fLozGHoxv8zJzn5ASyudBgdF4ZrDac20dUEF50dVoQ42Z+USDua5jcnlHiaRkeJncb6
kuXKTeECacbyzH1pmwzWC4Ok++BGBBdmWDWB1XcVMNCzhQ5+C7kYj3Garu+We5KxU6+fEwQjBtzZ
bnl0po9CjLPWhTcb7+gJ4nPRrn+j5EIbt/GcE2tQvRlsI2W+JXpAIbLPkNiyODCk13t+lfoXakaS
rprRnT5Ln2LnO5UFgWqOHdjxmtLu7qmCcTQT0adLeI6WEecoZkn4Vb6StbGswVpFL+mHUf91Lhcx
lPEs8ZaUpogt3p3knoRArZmsSGgWzLLBO05CqYJd4LkfZV9+u6EHayJxkUjwZSp7E8Tt6JcnIGMm
RV6Z1C5IklZBbH4KTwnN89a8U7udih4ywEEX2ieJ2uLioPDswQKOBU//mRghTAOrFCGTR6S+qPi3
a1DoW0KapMAtg3iecS5wiMo0qf1EADcXrHI3MOpJOUbuZamLSNrna0N+pH+VQT7udcWIzQo9n0Mg
vIz46TiyGPjeypK10HBB65L9UreLGhPmAPgzefMhiT3pGNWOMXixPntbX7QXhLLZLOYFq2uq7fDg
MBX4G18nrlDrz76GfcJh621ZWoO0Gv3yzxQp582Zmkd2O3ClqTqetuc9ohAXg/Zvc9YOgFzVMqjM
3K3fpbgL5Em7DNgCveomdCv4VnArona1z15lEzU+w1A/qNSLcNK1a6EqmJTKjajZ4Qo5yPwOzKfM
2ePQoCaX1EPXGoqYD5F4eFNy0YiN5n7WMAkqAPTYLQAArSUq8bwk4z6zi3LtWkMPw4Sf+VG+Tl1w
3AddELKbJpiIede35Y8FxEDLSnG8H7GhfiKEodR8Qo89pkCD+n8+eXZw9e2EOrz/tqHhXNX/mzv9
y/HSVuEp1t0QhtVG3U62QwJ5Di7SC9vIe/Ki9gHoyXWbQbDTnpT3FLQlNAkxxWG/VMiTjqnp5Inz
EDyf1mGsYIhvd0m1qKkbWEhZ7uYs8vkyMo8XjLMQUjYBPmPfnMfST8K3WtbZ1nuGmOTwI/+R20q7
IxTB/9Fh0rAcTjR9FwjGE66T/qS8h/KmzAcxqmejfJza3MzhajQnKftXjV8tEIotEqzM1PSXYTPk
Fc4otTfDI9+OULPoTDXqRM8oevBy6yzSHDZXr2TNVxRu9BJeqRGoWSIfZG/M6dDsDHG/nTm19y7i
bULjjxx0WgO8EcLL+fk87CVtP5qIwy85VPYuHmuEzNSZooqxn8PSqxiiklgFzjbnOLGHHcWWv17A
obOL7wz9lFoYT+w/AFKBi0/i881S6LjjkcMQesU435w571fc3LKmQ7Fwn8yPa3LbpnsvDODdftL2
jL7czr+vVVeeaLPrWXk0qykoPwMGakOP5wOGjdQVY5MdL6aWdHJFKa9FaT7h8Bg6dor5zNbV7Lhl
dWjC5m5tgIeqdG1+oaZ7cQwJnTfV6fS1t2ag1nMeR+1lipRjhZAxQjkmaDsm2c55f4uJ0gtRXxh9
tgHVS3WoiXM41C+AY9zBZtu3r50XkTYAyci2xcv5UOFa8Dc9VQ3SW1WA8rteRm+MD1a7292Ru1zS
5ggJ3827Qox9DIpk8h03iKz0n42IuCq/pM3x9ycUKtAaIogE+Kz0GbhLN2WMmR807L2XgP34Ocfo
QLZYB5Nxsba6UyIA3GZcuA6HnEBnT+bJkdgeQmwmG+maI1KCum0j7vybUpvFDibHwSqdTXSb484C
2WvwJHIW/FwZA2YfnJ+bd6td+HK7FaEZ+hWUm+kfnYbmXhDgk79SRLiZvI7vs8OtGWEnBvIH73yN
xjJDqwbT9d9FAIzfUarq8TkVmfnBvKcXD9aoMB9CGAiAwrjBriVCuxAnjxf6JjsCz7lOKIS3lCKI
2TX6vTXGoIDC3o+EUAnMIRQ6LVUhJJndk8QnRyPstEmGZEgSQ9jDchkYfFGtwplWmUOiD96ygi6F
hlZYJLyLzCXktEbKyRmzKluoR5lQA5aKvNPv+nyCHslkDMzuH6r6ByHPyeaX63rs26nh2Hnpj1Ly
yV9kJxLfRZf4S2RcTs3LXJyiGF93GMwydXiuMV3e7rx6UvQTUCAXxu1uwAdNR+Q2x37LinOatbcw
UQtISuA4Jz/ERgRJAyuXiVA6hcb2fnV5XEdOhVYkZb+BJuKFJkXT9xWNOOiKgAnuUQIEoxnHEehV
PYAXiGRHsFI22fqIMTKidZJFx4WQ58JVxFHVWjKLDXwk4rOwE6vVSz+hsBf0tOftWhoIJ/AISybn
87AXXsaoZv4pK7xKnn6uX/df0PChl1D5ZcWG/pK6YVgs4EFH4TLOweMhfqS6ztdvzDGJ23o1mAPQ
noDE3FFGa14tIFL+bPbFoqkj891iww0fFkepXW5cuaipIZGLMn5LSyJ5bWDR10ttUkv3VxKH/0O5
wmD3RONLvdo+jgJ0eyC699BCJfFxx81vavrNIdSVOyaMknf8XfmmJs5jmunD41XGTkRJN/FAKf3J
kT2DrUsx52/117s0uAkxPlCtB8H4YVicfhkugFd0GAIvXtnCDOWd12PDQqZdnRQuhl8pnwou9TXI
vZEemds/D/aDGYL2VG1jM37I5pm24ofeN3WIfwoxTEOuS3GkF+UKpdakRecwjI2kn+g4ryblt1FL
9Gj6/6YYJlRQHf5z4aK+owjJC/Fqbjqx/ZBFCJPQj2r1/yBkUNXAdWdxNIFzeopoBqzA2H8GvwVM
4f1b74qaULSNQy9kCYwlTc+ZvSw4RsS6IWe2VHpCPxm9WN6gu72GRiV2NvywT8Zd9bRBqsM4jWVw
Tr//PnF5EvB3hPld5dVeShOcAAYk1wrU0NCleDuBnoNhd6qX2FfWfwtFmQVcRm1SOa9LhfayOMbi
sRK4XIEERPQr3cS+4jxWYi9qLeAycjptTkUhVOTWZP+moDnJ/YlSxPxtPFatJGNoMvaLoD6KdoCp
4FF59d8EqifeF4WsR+3OwzH9OxfxQIehCBqN0xYgCLXI8kJPmpSDwDjTJZAcONuNCBwCysgSByw8
i0RKdfu+s3vHGKlkQIwKHyu0lPc4VwGP8jWZAufnsusgMvfwyo25B84FsmRfqXHLbIygaWKe7O7g
Dp3XJ8npJQApCFaHojiXbJkzmRaZbCr6JPo+NLKhsEf5Yv366On6GL7MlhDOz6eAYRopoSpK+AR6
glKQ6DckQkqOiDOC19W/9EpTL/wLf0lCmOjZLTTxPb/oihpMyPk3qQtttwKM5mRFGPSPbPmmK0rK
a6+mX5nEJI7dH/oloCevp45rLmbwQsdIsh8KFPEdXbo26lQMppM2I/JMJng7fS9iMr6+2xpaXMZ5
WXP4BB+fUD81qVYhVNDno90gy+Gn2NlhqL424u5ztfrgL22WlAtNRcPptYMX7mgDzSP0Fa4HVosA
2Xy5P5r7AEZT0jk2eCx/epLXbH3MOpyo7HgPNFFck9+PH8HF3H3+NwfNHZL1b0vx+BSielbE41FC
BxRnPjIbBLBGCI1GvUcf004cGhqrmLJlQ0XNaps8YKC1Pf78XbKwSIaUtzsd/lb43Jr1DAfjXs0u
7xAlIvmpcIUjPtWyo+8G9rue3blk3GW2llnjWh0FnYRXitgQdsYQBbeJmrRvlEHnxEDih21pncNG
QqmZSjvL388XID7XgMOBe0rWq3ysGLiw2kwXVAppxG8tlCOQ2Dqq0JPY1jNP07UcjQtWMTHI40hm
gS5iIS1fMzrcgZDpf7vpR0t66zGcg+ZGnW7jnb87HhSc/IZtFmvw83UHtojS+ayIZAugPevvESB0
2x5ccvqrVSXjGomUEwY9DOW03OYrUsLB3OWfzXZs72vjtja1Frkx7dt1pXW315kWj9EsGMA/XzEV
QUROwo1Ue69YxomWJJ2OfOHxirY6JypnKP+Yt/dKPVxIdPeb3FnawO++gDjUAwfygEqCxVn49ikP
fVRonE8dWOZJDdnEz7DgA+k37zSqIoEUtgqcMJE0TxhRSHA7JqcGhbNadOR3vPVd4AdMx3cZjdk4
5wBJRrtrbz+9aM/UycgthMfpfYLp+IPtlPmXfM+vdZWHGWPulH+KlyeLKEU2fqdHImCVEkT6if0g
pmu9mwTM5eAsak9TjGgCwSO5WceQIRMZzMrTSsa3rHKgeUzC0hAtdWXffsFqhKMOcQMy+K5SfRQ6
AdNrtgKI3grkK6yTNOdsw89sgpAPi/T2MIrtqFefdit2b0G2J8WjKr7JV19gQAQ6W3+KZFSc+/pM
BTHD/+7ziEUlxdDtYARQdu4LB3p72QP6/mtprrUnEG8PBF4aE7oKX+88qbinUg6+qDEWIH3D53vg
LQ1UQ9tJCvgxEduIR9Zls/OEkPXVIitnzmMTljeHR2RgP1HRwbuXDURa3v0zoQ6D2ZT7t8pE2XR7
Lz+cpLRnV3cz34RqQJkX4KfiLNwHs2+Cpyf5UUErdbGylRtMQ2F2ADYo0qRTkI/BPIXtSKt53V4X
ZqBhzMwmUwT5y4qL+1VuiWyF4TBImuC9OafMoGYnqS2zrb8sQYE6D5lMX7q5EpQPDk3Qr1ai84Ma
Bupx9ikGppdd5BldKZE4TnaG0mtHuZJbgfJpc4n59Tulco480crNxZ6p5QG8le/2QJ47zS1u4JvE
W9iSQfmop0FefONF2lUAokEa+egEpB0zPyvgeHQlNaKqFM9AFMm8qa3Qm6sHcnScYWzLpbvPL7aN
FzrBt4W5WSZIb4jkE8p2CSpTgTAGoCQ3WA004jjigHlz7B5O8Uo3KSSXucnDvfRMLiIl0jDB9t0O
xIIkSeWSA9jc7lOsD1AkAnuOzV+0QGdUEu5hDIaaTQb6oLl0bdiX7iq3hDYDxAkIeNVxdUwYi6Lk
bHtln3SJVzpqEfOfKn1hn1BIYcYWc7aC3D7vijeOfyRlIxlMvH8yzjD6XaL9fW+9bpPpPfCb04fu
DzZ4u2wRlWHLRKntMDNdV0rQLvpeo0Og88njy8Up1zg8z4qZMjzyQ1Ra87sfzLjmHUYPkVyYHKnr
48hZYW8Nqv7Aw97oyTMW+lEcjQSzA5Sl8NIP/CRhRNMAuLRSDrIifS4aroitUPxaTrKBqxYQ631c
5CLZRPb/pic8NvZ6AukHsNLn5ITrvGfPqYOg6TxTyPs74D6a4USbESsqHSibx+RWet1baX7cA/bU
yYwuizeyDIxw8EGePGe7Edzql0SB7evUXEisXHMILR7UELKhZojqbxLQ8xvvDTWlG9FXPO71Vsyw
mARKxgLFp77BT9Wku5LPsuyG3eX2F8craWxJSVKJxPmmq/rxGdo/4yNDZJQcs835pxIIgmOVtPNn
pSZGMt5KaohmiYGjqo2xy1cXrtiOygY9XPG/UpZASk+nHE/YWim2kpGkVKp5ylm6cF7K/Auijrsf
XvYFuIEnEOyZ4cDNKd57T0RssSIRCyYMkPLjTHxlNnRmVMkRZjVWVbStcrozJfsdWWYUEO4djaxT
uEdm+g30OozqRZrywaVWCAWkbe1kfwccLCaowHAeofWC3NqzBJIcKX7XWLWRV0oz6Q7vk69gRcRC
9gi/VOgjOQW2UuVzwM9E4PZBo6w16q8VU9CtO7vSGFjlOode8Lq43gn0ohrDTMiAC+kVzIcXCP0V
/bwTgnHWE9Eo1fgUkAotiH7loBy/oj0Um3VmqEyTiKxOFFRh0JVCmhl5xf0bCsnNBUPkaZKoOELK
FGEAlW2woyyi9xAGfEFYFNY1GfsBFb+8pBlYVNZJv5jJiFntGr50k58wtN6TWlwWqRjXx4B1hAJZ
tMxxGFP3ku3KNoz6MRanYEqguqj6HA4MpE+KPrFzykxSp01k/WQP2c5IaY7onfIqp9M7oVGLUjOQ
Y4dgfJgrHmC93kmfSp02VzNlaYXL35VLwVBc7grNRf4bafRlAWF1ikU6tGbTksO3UO5825LVOcpA
vpdMZbScToEEuOpf2/mlvsX9YhqqexkBzOiNjuFf87hBXpYRIYFSedEYdWqTwmXq+0XDcHBo7cM+
fGKJZqsUfplJC9CiArxbGRqwMADZokS7ltCT7lCgetmsZ7//HbpuHl5CaXOuexlfcdNrFeryDynk
TXgDh4jHqCITsah8RZHmKlY+DSY3JxhMIKCBMjiEra6sabkyAM2OHz1TefcpbHHQuhtaDYhJn+ro
oPvH9ULkyHFz34VzJd1SMDBb0QlZjy0D+9b0pJgY3CoZCmPXX3iFB+3oA2X8uCHUYVQ5Pq8qm9LT
UIBFxiVfPZJbO/VP2KSGPpL9Qi/Cop2JHGEwjgKsQ3+UhnLIpTL/uKAF0x1bmf+ECeB9DibMd2uS
JopKRBMjevmf+sApckf1Auwf/XjaUytsiCfRgA2xL8fguNtoBUuTiMFN2Y7Q3BUEW3PsnmlXSvey
66frX/9hKnUneMhtXgBFSSUBheQXr7xFK2Al4PVpfoidIRg/4kQARpemsk2PUNJ3GYfNXga4IevR
1rzWv2U18zeZScVm4rsnmTQ9g1Uve+2Vr36K/D2Y+YBvc4BbBOfeEo5wAEVGuw7r6XCTScdEJ8f3
qyAxBvieiEAgDBh8gb1Uj754dzgAfPt45RSQJ/oavQPiWdh16Hgwypm8ecGcEuWOv6oTm44xTwYg
cKL03wBOBO0rmVyrho1Mpe3lYkEyJE2gAa3umHDYF65oAHSP/Jt0T05sn9ljaqHf7GYk4eA9VZrF
VisByLhJt64i12UIXpnHiyDsGY3CE0FAOJveqjO1wVxMrsXHf/37Kd+SLqTkHN0PBHVXbzcYemIF
bqq7zCvFTAv4YbKaw36TIlSpJ6z+wl/JrNoW/1EwDp1ICScWolGY95hKOHjMyefKaxrZ625lddfs
XZHGsRXJf+pPy/1dKqbKxmZWXU7OiWhWkBfH7AZbRlQFF12f1Z6NLYDYE5yk62o0wt1XeeAhXZuN
wl8+GN9DEeeqe2vA4GJ51Aug6LIMykFBIpnacmwiPbBGpOdWFXNhxctmF9pLb4EnfvBzB5adVKmo
NNHFkZME8XmisMiqcDSSybf1U8BefTHkmR2KXTbRUYIlxhRpy6fk6HX3uIvzNeI2M6y1tHD/y97U
8ZBhOMWiFAiDpOhld1BuoVa23x+kT/92eYS4DgV0ljLwAvann/8ViDqA+iDC6j9NZWXYwP1Tf1RI
PRadDiDTToFhHC4PHdxtuw1B8vWO61W+8cQs46AzUltXcAKQvzl4i/pCCbDzEgpY++7OLt5Fxv65
BOCY4nZUUVXo0Qa+gvx4/zbcBwvw65FAan3DbRO0gpKtieTiow+V+BgrqSB/QP5bYtP5yjGc9Xf2
pBmwKl6aS3MIFL9ec0JEo33pjgydGsNlpi2+WifbmET1Hob9BHlp1FH3lHk1xYdjFiiQt2FfaE+R
cdwWrPwnfOkW6eU1Vvctp9KWFOy5iE7VNeNE7eELogZSAfX2M+lUoOgggzOgIgfyxYMn037cfy/w
ySd61GoNlFm9F104ikYKPLiwsoJQBL6KiJPMU/iXIINEaqBzXYmJQxQmrgKPrcunD6ozzyEZq1YI
JY5CCRYGmDbasTbSRqQYWwbnGeRrFu56MzyWx4WfasVeyLS1708c31hlDd97UDOze0wKTHrDF7DF
m5xjhnnrynb5GYjPyEz/zkmMt6lB1tsOvZ5NKqbWFdbOUBNXGNm7aZoOYNSIgVt/J930gMABI8MO
lz5+6pMq4FVz2g9uLtuax3HCI5GsrJnCB7PY7QTWrnRIq0Ld+L1iYHPupFyNVCLzjIPucjiVjyCS
vUvVfz+isVbV599qUshw9NHQaodEqPzogBO8DUmPUjzpQX/k/AJdoUbpBjJkirT/f457JmZIGUU5
76Eyyo5FkgtyF6Mt+KkZsFyVyuzHfJecSObFlqETjwo2oMwi5yPtK09UGaRHwqJlPQyA2QYh3qpu
WaZZQYGjpXASm674tHW/453bIxIoO+/Zq5xdIxN9fmnVoHK8p54VSvH3ZApoKiOZmPbwE6jQkZop
ki4FF9h7rSlMAMkD0XjYLKe0h5nGBYrCOz5XRL2gI6DNRjJ1et4FjffivFZG63zP2WCVkYwrAuKY
/W6Kz96Dhya7Q3RsFoVGF/imXmItks7Zj+5/vvSVBQLOK+6UgJbciujgRthHxcvdfN0jjRp/LHcU
WDHk1MPi+VjSzUCSEdJ98NoyL/5Sj/EVzs2b9Pi9exZ90u/VkkX+0eIJ4PFiP9AG2kFx1dgDXEJT
KLglATbcbBnh+WOT/i4uHHi4MePieY+DR/zSbDULiLo0jJr4RsaWzhli2yBJNV1/UCXhTlPTTYuK
aE8NvxfPX7er4dbZYMunhOcu0awK2UwLvel8GEcZ3y+WxDMLMkB+hH8ygpNm4HH+u6ZVjscHISgQ
WxNeOmk81xyp9EC4edw0mbhxqHXKZDjtVi2OhYZn21/x/2Bgp7uSH25a3naW/5uQTS1n5eNzaNQB
mmAWsSEhx6oMa40i2yYpnwuV5kNPRV7YkREhizGllLzV5MqLL3XR5Hk3vPes7eAd3RwAwqXLE16x
v+Utfn0pXGZGRoRLV6BPWT53O8hnsXwIIpcmb1dMnYTweJZxJ9+eLIj3GGHC0Yug6yVGcopF7Npb
WRLMEb3m3gCOt8f/QUJ2Q5OyXMkn6QdyX6GQFO734+DHkoJoiSB+Xm4aCg92DWIFYx8BZ5WGB7Y9
pY0XbdlBFQil/R256ygUGywrJhnZTesUkYRgGSIHTwgxlQQoh/TRgljmPAYdRI+BGSXc4p34tdB8
HT86mAXxrJNdOJ0HcKrK7cEQ52+koNkqe//tGtfC0Xku04Dd8ZTb2u/wzyl1x2hInw7ODsXNeZ2i
b61Mq10dnqXeUqU6Ncv1Ijcq+hsX
`protect end_protected
