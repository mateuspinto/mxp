��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���g�"u��L�k��	R�&N�Gc�݈�
f��U���i�<����Q�j�eb�ttt���y�lo�?V�-U�W��(h+����z���=h�*i�g�CS�bXpc�M�Y�x�Q-��{|�u�� &����5��wHmaU!�%SP>��YA��tZ�wQ���>-�Z^*?���*�;��^/ÅA�`��98��ܪ�Y�K#���/�y��y-o>��A�~��j�d��ΦT-�"(=�U�?{���)'���kP�5rI�6�,�y6�H���`�='ٜN�&j�B���a}jQ!K��|8>�Z�]���0p/�ąiB*���^5&RHG��mj\�o3|��k�'��,��4�[d�2z��+j�M���=-
�m���D�	���������J.��'P�i�-���=�z﷊�i��!4�A1��k�-�AU �I��`1�y}�+H`0.3 A!dH���b	R�����GI���?W$n�3ͥF���� ^��=^Y�_��m��a�ɤ�73h�[>8�������h/��wFJ#���W؅ݯ6rbRR	��CߐK*�-1=T#����v��3g�yC��������B��<G��9G&A��\;��mE�ʖ>~�y�PFZ�i�f�~
�iL�52���+�,>~�^iX�j���G�%s�b,�˟���Lk��=z�g�/�Tv�,z�l���ߎ������v�;,>?GtF�v� �9o�S�����d��n0nv�G;�{O~XH�6�&oh��1�i 0��|#f���#��	�E��_�l_�'4�]��a�C����E��T[�x\�h��f�֠Z:1�] e�8�.�zV�!�&3[�����H��i ������vp&�L�󷞫�Z��I{���1v�K�+�x���wTos�K�{��D������$p���[�O�������������ut�<Vs�N��9�6�D0�e n����*L�d;�����6��kBaT�o�3�L����Χ�Xx<>��{6`j�y9s=�`�v�|Ck�[���t�����O�|�4��:����O/]��I� 'ʁ��s�4���s�Ŕ�!!�9j=�ѥ0=�j+ ��P����:�OHb�}�l��ִ���4�A��l�	�+|�P��;5��6�.��P�K��V����CD��"DqW��rF��MN%Q��W�t�N��k�LC������f׎����5�{����^d��6��v`�"�wt��g�e�Ƹ<]}BCr����>��ɿo[�o��D�0q��/��7��b����Z����xm�ivmv"E��<V7�?��ۓ�D����'�>Q�`|˳9� � l�Cw��u� ��.	T���/T�,I��Q��(a�<ȩ�.�@P=p�Y���:(u�����BlA�T�_f#�^�0مRV�ԛ��6Kw9*VTle�c�7�*�h��7�����?���"�Ϩ�ˏJ�����P��a㈳���E���9��ά_r�`7�����o�cxHBqmr�����g��E���n8�!5�;�T��[WS���^c��m�3�>���Z ����oN��n���T];�����4s�(�BEQ!��aN0R	^c�Ŕ�d3e�d��yӔ�+8���ŒH�,9D�Į��?��E�}����|�B�.F͌zr����[��$������<���s����a���(��gg���_tW���v�8S8ޅh����D�o��	uJ���C����kf=_�������)WU;tp*J��t2�?�� �-�A�~ِ�R�q��ΖΉfq[�Es�z0Fu�F9�/a�h-�����Z��߳�h�?�`�i�l�������v6���"���Gw��D��Q��س��d�;%I#6B���E���2d�7��V�N�J�Z�	[4�B�m��L��-��a@mo�H������vn��2��#5lT��1��_g�?�'*��S<2xs�l�[󻒽���G:�B���7��g�Bx<���j��AܰMy��L,Г"�/�b6P��y����+�?����t�sZ��|��G<��\ֿ����g֣���E=zE-d�*�_�'�k-�ߐ,�EX���d*���B!��.������5����8��x=����i�o#�(ţ���Q>�ꊣ�R�Q;/�*�X�,����ς/�_����*�ts�0F9����a�a�� �K20�ɠ82�.����i��yw0a8�&��(�K��AC�P^RK@I�̔���V8N�}!J�	�	�YҢ�c�"�ĲQ/K�H�0]�i���|D���	�;o�'���@�i��û�`Mq��3
����"@���j��ZP�.���绮0@3?ؤ��)�P�vˎB�lL��l�<Z�� f�Pط�l�������ʏх�Cx[��2��£8�k��)��PDX�-�C�"�*G<,�9v���N��ߡNy��3bu�� ���cVd���y*��IFtϒx�}�:o���_�EH�OC��tl��uA�
A�L�D���6p3r�I�Y� �<�^�����a;yz�Rw	����A���1���(��+���n/!*����*�T+m,���)I��3�߈2��
xm^��rU�j�]#:��Gx4�"�O���ZEo�r�9�,��qI���t���x��||#ƃ� KF�+��J����p�0�Al���|°t $�:�0y#���xe�����*��5�>�+Ŕ`��z�R?ʋ0����o�=8�G�*S��zټ?�eh�H�c��"2:fU��sp��l�A�k�ݩ�5prEP�EVg�6���
���;'�7���qg��Z�.��P�EZ]��������qG���饳�#�fU���v��K�%���@$��ڬ2{-A��{1�A��X_�X1)��2vAl	�I�+�R['��{��9�_�W����쁘�v�1�,x=�o��`PxHI���_�ѱ�M��^����x\�&f;=�|<U��:b�b9���'�t�m��ظ�w�R��Tӏ#ĄN�RB���$�v1S��R���~z3��Q��wj��Lnj�����W�.c��*M����ca]sG"`����	��ea��U�Uf�	K�}I�g�����G��S=�z��ӓ(`��s#��lr�R����}#���Y���E��ѥ�>���+�;�r��U v�~�Mщ��@���	±��_�[����	�[5��� �L�˝/����)K�]�l)K �"�#��U�C7����:_�(dN̝���W|�EUD]���2v(!L�4n�G#�d�\3dj�xRq(}�x�� ��rz�������EX��J��3&��>��\5� �XQf}*���m4�w2ڧ�i���W�oڊ��VO��?��T�ë	<?��YZ{<9����		4��R�73ն{�R�$|�KC�An$&Q�Y0K+RzLz�ܠ�Ww����@S�D6��=���_3	��j��x4x�孢
�y��O�K;���j�D��"�����n�_nvRr N�R
ȇj'��1�pa�Їi8���ݑIvv��<�q�򵉸�� ��l��Db�a��)]�l�_䎽�M/����z�Y��k��.8��$��W�i��V\C	j5�(b���̝��ն �u�v̀��pG���1m78��!���ʵy�u�tB��7oK��2"?-?n+����`�T�r3=�OoB+��:l�MO�w�b?DSۿo�fc�p3�Qn9�-ڂNK�t�mO@M+ߦȒ���\�F�ű��4K8QC����^Z��8�Ul�*���gE��y͌���B�vAm[����2C̚���(ݛFZ�o=�GS�C.�M�і�����1��Be�����<���]$��~o�I��;x�6̑�z��Z�/����mKe�$x��-jn)��Q�J\$����rz\׹�hw;�yUG�)��Ƚp�:�m���j�w(Y����bi�J��r�z�ʈ�Z�j����	Ҝ���	;��y��+Ӡ���=T*M<���|64ړ����GW �2^ ~'/%
�w��P��������B��gWczu����Ԝ�n13ۮ��A#?��E�4���PV�<��c���(�6�zq�\�]�y�C[����K�ro�@��p�Yo�ϲN<���&���̈�>	Z��q]=OH�&��Tm_���P�'tW�?Z-K��>�{&��*�\��B.�.h�^8'�&%w�c�ǨrI	C<1�[^ oLDN	6�wl� ~�۳�j����*��<��hyY����C�/:	4E:�)a��(:[��:����Y�����jO��&�֨��2� �ږL�X�4k+)#v�B\䍊�A&k���7����A�Df.�Տ�� �Eo(8�=R��P&ڹ޿�"wi�k�"41�H�S�轱j���9�_%D����� �ʪ9{&X�����ĺ�*,:��FiU�-D�l2�c���q7��W�[�>���!�{��߲�4�F3��=dh.�v��� ��rL�k��o�I����i�[@����e���S�R�!+٦�
$O���u�ϑ�=T��~'����{S�jsFQ�3pvp�\��7���W��@�p�ɇ�E3�%�"�k��LFU�N����RR¾{Ȓ��|��:���-Ơ|���jT��hPJqh�Ȍ6��������?����v�r��
�j��%~h�����nɚQ7���#���V�A����rfL�����-�>��O"�ٗ��쁢�v/�sK��Y���٩�Q�> 3�w:"����8����J������T#3�-w8�Y<80�흺�pBA�K"g���t�k ٫�M!�B�Eg���uܱ��1�_M����9(�9بH����Ϧz�o�\�K t
yn�Y؈#��a����ɢ�*Maz�7�\�%K�u.Q�2 	ay�Ψq�`�U�	���[�L�,*� �t��O>��	�*�`��n��+�N�l���]���.\K����;��ľ��@��/��k�~`R��$C��f��V���6�0C�Yg�,
p��A���11���S{x��"��n]i���OCX+�d�����l���&����\���N���+G
ؽo�Ls�Ԇ���ʈ|��4r��1�ۇ�x�ԓg�٧{�����i��k��k�����b0��A4�b��N5��x�25 ��f���g&�%�|��O��f�+U��h�Y�*^��q�v-�.av�'g:{>x�[�^�����0
F��M7�tb��_��0B�ZH���qgCџ�\%`�_�;����{F>���I �	����J��
x�(��`M������я�ޞz��1�|Â?5��ߩ��>1u�Z�iq��zW[IH�w4Qq��/�~����Wr�i�1k�CT���O�ma�]I�M���~,�=��a���gO��Xq�r�r�S�6c6N�:�>�-�,=z�0i�)D�Xs�vʆR�kk"��E���ҁ�v�*o��"U�����վ�A��a��Z�P��5!�w�Z��Ej�M���ZEW_��H�e*�lKl*\�\$�ggeKJ��_��%�dl�'SP*��Y�|X9����w�J*�8�J湧��8zJ~;*�WZ^�YǱ�!B��?�PU��ӹI+�U��,5�0v�ӌ����b�0���\��ѻ���A�Wżf;!�2.:/|���z[�p��&b�?Բ`
� ]��P����~9�	��Ѯ-��ir|�rS��avcg0z�l#9���xx�zаA��J�1�_����enH�� �U\�a'�JkL鼷���+�nT�S[�R
�����t^,����?���^M��}+l�6r�M�8��.�Ӂ��$�#\���a���ɗRn�zM�v�������$�m�Ot����*/Ӂ�z�#�,@=˖O0[E�o�:k��ط�4���zZ�Y�>pZ!����0�
X�E��1�,^�<P�D�<(���r�vr/��G�pz�1*S���Z���[vR7���i�PmN+!��G2dcAk�Ӌy�TC�M����!8`�q'��אk���ȿa��z,!d��E�5U��/������k��H:e�Ґ��8����_�<��i<�oZ�o+�����[�8�'kx�o��>,N�UJr)��B����̐n�gg�������s�SG�@_�.@S�h�-���⹰f��x�bv�p���k4��n�IJ����/�,�i{淖���u�ѩk�b3�����<��$�,%s�ݙ�Ma�͉�8t!��\�'5	t�q�=Ś�	ΓFN�ܵ��M[K��""����:����ɗ��vI9�̛�+ٜ0@�KӪ�H�`�S=H�'J�"J�8�[�V�&9Uj�r�9XX!6{�Lc���҅^���<Z��'ݤ�����d���ƞ��nd���/���l�ӑ�u������	����\p�?�8�����%�V�F���v�-�v$ʻ�����@����I;4a�"�v�&��+b6�c��M�)���,��#�.��7c�/�D55������v�l���S_x���e�P��y�~19��_���%U�U�g;��$��=)�F��EDzɍ�����(��JwT���}ӑ)4��ə��z=�p�`fZ�h̿�j@{^ڄ�b�[(�mOU�=#0�`�1$'�>4h1yRK��9�� B�Cᢳ|��F�81��pL�rAhc�tN�'�qcGC�T���=�(���br�2��*~?/������CÔ
c��qd�pˌi�X��:��� {��7/�B�\�oEEe�J(��D��Q��S��	�%�W�4x��ι��9mRթ�&:�X]�OW�G!�{��'�G��6�߼�{n�%�G$�X.W���ߍ�_��_�8��X���!��e"��ђX�U�5��ṳ���v^j�$��ma.n![]�n�;���]y�s���X/貌��-Ɏ%�)����`s<�:�;D;��)ݎq��K&�p�D���P�i/�Dz�]�/��!~���{�=�/�3T��f�x1z���h9���Y��r>l�Gc?����=;h��V[��=��r�Y����Wh?/.�$�a`nP���_?:�(|dF��{'�q�ո!�2���;�*��TǑǩ9�W���F.�q����x�?%J@�/m��xT8�q�ϣ�3�r�m��82v1E�h!��G�s轫�L=�^E�e��{����2�J@�����ذб|����@�,0Z���^� ؼ��<�Rz�rԋ�]Ȓ(�6Ԁ[\>Y�I�aoX7�	��]x���1԰����l���"��H�r�cz%#�s"���]rv:K�?F;><Y��.���D(_���}9�c79��`�!���,��}Rn`��·l��]�B�ʬlױ�Jq{�$e*��5�r�Ck���`K�9۩�!���5��'�ԧ �l]�j��a)�i��	�Y������`��)4���x�������U9�nf�� n��icjMX�f\�����#�,t����Z��[.'��o:5G�Cm���պk\!p��^g�%�o�܆|����qP��v��׋o�ı�2_�\d4�cI
 cw�`'C�p�C��]�>s=I���������Y3���a����� �~�����Zt+�r2��u,÷A�Z䱘v�A��p���H}�[��4o����M�?q��گ�]YF/����إ��\Y�L�D����;�_�1А��YqPs������6A�᛺�̉S�T͹Sm@�<�e����+R�\(����G�f�rB���m����m$�Wk~�B,��	o�.�`�d����F��2"J����Oha����N�#��y�ֳ��/����U�}�9��D����#��g�D�|E��O��}j�����0��$��\\�m����	WY<�1�s��x��y��*�r���ϭ�oK+��t�''��Ȏnl�b�0���%@XC�ɴ�)�4x�A��h"��?�3«a���c�T�i/U�$��T��o��Ai,�n��l��d�"W�?&~����)�`���&�*���c)�#�.��Fqh��9���D#�~����tʢ��KK�s���|��7	�F��sk��kc�7+��نT��i��Qg�;��7bS͏9�6��Ӛ�\�G��+T�i↜q<Xw�r��r�B��4q5��w=��ܻ7\?7�FD��Q����qS����G7wμ�btg˞Lo3��������kh2f�^�vuOФ����d�M��Y� �G�4ͥ�.a�O�}X�R�iB�C���:u���atá����r�?k3���a�6h^h��(k��M��s��mO���=��ƐK"o��#4ܶ��/���ȵd�.)-ŋ]�i�}e�5�Z����i/�l����o+����ݦ��s��PP��jsD����n8E��#bK,�m�]Q����=���Yr�諃�j�p�ȥF��NKkG�#���,oǃa6j�;�'��;۲���Q9��$ۥ�P[��D�S�{d�.�!�F�����vjS�fp�r>D�%LC#�I����`T�9:��^s��|����	��@,�#X<�s\�ӯI�1��P;���?�hW��X�e)׉����fO�Dy�
���v��8G;QXg?.xs�J$�rdY�
3`�'$˖gT&q`�9�7
�:4�ÓKnN)�o+���|� -N&�r�Mx�����>���6x5U�Tfັ�:	Z�Y��e�-�r����x�kY�S�����	�7.�E~�[_�1$D���/C�l2�˽ʃ��8���'j8W� ��@G��r�o���z;�\��PE~$��)�f��[X]���|�Z�+ ��J���Y�n��_2�T<�f?(�hF�O ^ >h��aҎ1'�*�������[o�u���I��4[��L M����቗�TL-8�+�w1�����M4B]�R�yI���W��i�y��%�� 9$��/�sMG��{4�o�x��s �v���r�ń��o������n��4/P��6v�*�r�Ӫ�u�4��1��\����i���ד�#���A�'��]?�Nl���5����=���9�բ�QZ����D^����p-������fgm*�c`�íV��]|�8�1�C����ң�"WH�,��i�B֗;�2�~�1�:���E8�fj�b�����*:�ޗ��T��|�� �o7�-� \��:w��J�^M�u��o��]��:��W,.ݎX'f3m��<.��Ch���$�)��a<�2����AW:\�L���c��/�[�O�XlGD�K,�/=��
�����$Nb�^�l�pM:�����V)0u��
 'rnq���yRUqj�M�~(olr��692�E��[Q M�#�V7�u�_����&M��Nז��yռlW���RZ^�4�����+F�]J�n��W�?o��������yK��M�)��s��lUM�=��*�0�k�.@h�H#�=��g���l��d��z\�g,ҳ  ��@�>�J�$i)U��_c�ހ"EH�|��e��t;r_֙��cV�˸�Nݺ�g/��]���ʉ=��˵�=/4��.�v[����s$�X�Դ��Ð+�mw�x?\n��+����;�"����w+���A��1-���;��g�X��Q��A�]�//ņ4��~6��:�"xZC�I=��	�e<��w G���9cY�\�z��+�k2�r�ڭi�ѳ�/V����ZݠϤ���J�h��?)��-�:�C0�ufOJ'�٤�1�+M�gw M8�"�h0�.I��_�@�Jl+\�쨠=`ْ���`U���C�.oΫ�������q>Q4eX�zJ���q�(�"��a-*����:�8Q�������A}�k�x���I�^daȯJtҳ���YjLL�=�;�P������Ӽ¥��3nKѶ"���?�`"���k��aE���%~�8�gS�ִ�v�ѠH�܌�@%�� 0��"s��,�_��U����-L�<빞��J6옩�e1��&�A���۫*��Y�wM���y���jXx�	y�,a����tra2�[|�׏�GT��w�61$
�Z_J�,�WO�7:��'�,��b0��`�^�}�J1j���'h9��s���lP�q���^�jS��K�@�]��?<��Y���?�y�o�����c0>z�r�!�ݷj��s���!� !Ռ���ρƫP�o�Q;��VmC��V0�f!4uq�no���p�#�㒻* v D�j�3�C��4L{�[�o�G��|��߸\*
�2k���K{�������N�Db�ח����h3�ű��b�@_0����C��>�P ���;��#�f��hk�@��s�lD�[Y]!u"����]c,�0��8/�jC��U�*R��H������~:����l�2��٦�'����0Vqx�b���D�۱���6�K]ă��b���3�Ov6�4��p-%{�%���kbZ�d Ǭ-Ѹt!�B�17'���6�M')��e�<F�E�9�4�f���n�Ɓ��ll�[:^�u_f�S���Q m8����	�3����u�5�sR�e��x��QR�:L�\>�s���v��2t�n�8^�R��]���z�UnW����%��8�_]�����F%���">�+�0�R�(�it<h��d�Gt��e�ZNT�� ����+��TQTX){ōk����~���):����e�M>h��\˲� |́@דk
j�a��G�@ٸQ�85�;�M���yYw=+��Ҩ�?2Q-&*�ĸS=.��E/^���,A��o0��Q��	��;_x�#�0�}�̊���i�f7|)�#<7��ȼ-iU������|����ȹn��-M���̹B�*���}tN:(�����䨓�?tS�2T˶edǅ����U��ﲏ��M]��#��%da��xb�Hh�me����\�6�?�iy��\�ԫEE �����4�̰o7�ڎˉ��f5���Ģ58n:nW��5�� KqA�n�kXG�k��� �X1M�1��,�����k�.��.^��'����O��tnmv&�Z�Gash����	j���괇�����k8u�����
K�u�7���Sbs��H0���0�M?<U �oed���f�rxr �m�<���q?q��p�cgH-��(5�'�J�D��j����&E��m��j�*4I
Ts[����H�C��,=����ݠ
�c���O*��CՉ&����8+H2��b%I�
N��O �~A1��x��!��έ�m��;�$����"��3�ӟ0R���\Pj6��0��f$AB[��*���;��㍜i�Wt��W���<!�f�:���M�.E�p�J��Sߛ]�G ����� ��r�o�ȡ�U,,f����*���s	pcK�-epfȾ��!"5�n|-y������5�i�k!ƥb�I�,�9��� <���aί��+���\�i%��Ξ*6�Ź4���0��'��Jy+��Tč����i�Ѥ^>ˏ���
Y�E���-��j���Q���s���` ���'�Hq'�F{t�^]-���c�I�Ȅ8�����ɯ��5ȀZ�K�Q��1�q���:����E�����ܐ9�{�c�F�F���C]���ˤ�:8�y6����X@C�_056�jE�/*�.�1���
�iv����,�kOY`ީ�ug�VM���"�)KZ� �ib:���|��ߓ�ڃ��=hV�[F��y���u|b(u���R�D�h���`ᗂh�G���>S	W��C)F���ˇ�H#D~
���#��� ���(�$3"��;03Hy�Tl&u�h��Ou�2���\���}O��y��Q��ZW��s�T�얫klh��Wk��UNe�'��*z�kR��H(�*�P0/�%��tJߥQk��,ѱ�)�w�.��w�d �D��Ub�е����`E_\%$!��~ހ�OZ&��q>���v�?i5����V;$zv�-�V
�u[ћ/���	O[�cw��R�ā�V�t3�<�ef2�x�\������!�V�;�[�����@J\�)+�D���G�̶\����Ok�`i�U5Vz>�W�t>��$,m(��*��2������J���X/�Ճ;��C�   �U$�n�ںS[\i��ڣ�!`As+W������qK3*�'��e�G����v����Y�����i�B ��PF<�ly���I	TG�G��k#�XS�c����p�jo�6�~�#�v�1n�;�paX����ʒ�UQ��>���pb/A���9���T�e#fO��&�(��è�@�aMF� �B���:����s��C�L7�"E�K�|w0~��~_+=OgQ��V�U����b�E1�m��s�&J�'�;$�W�������ƻC���v�}q+��.@#t�����T>�x/��S��ڗh�c^M����8I��Uuo- PP5���)��\�w��6�R��]ʳ�k����x���r�="�,��I1�@گtո9�����"&M[s�_�/�@�kT�'/�[�<1��އZ�/��Y:t��>�&F��tL ����E��W��{�j�<X�)C��wyH��l�2<�u��s�;;<���e1ga��O�%��n�c�=��i��:d�z�K:��!�u�����&u�j��4F/$���c����Kϓ�O��!y�mPڧ�$���6�Z3���:V�a��nʲq��-�BBΝk��bAt�C,�
Ν��i�{��,���1q�f�4,D�P�*�f��R�+���M�G�u�V\
�I:�5�qa{���3q�e8*��or��.A�F�4�4Ԝ�7��8 �����7Ҝer)��)�� MI�E���~)�;P9��p?��td�|��6�����D��G�n`�>O�]��Z����i����)cyB�d��{�ն� �}���v���Z�Й�R��Ohԡ�o̮y0v��1k���z	QqFA�d=�����wn��Xl���1��zїiP5�k��A)x���dOf��3�)i�p�09<���&��N���J����E�hdײ�t۞���E��q����`Rt]�W=�3���^i���i��Z<&*$�U��аA��}u�'�X|��W�Ԫ{�g��k5�8�]w���v���F�=�*����
*�կzqeit�"߽� t]����͖���ȳ�(��Zz�Zgڕ��(�B�����yS�ɲ��*O$P~��l�-����$�nھ^�0�љ�;gR���C`�(�d�C-6���&�j-�˧�t8�i�� �iv�픋`.K<b�y���|ξ�H��8-�.jIe���0ϐx��r�ox?�ꈛ�'gNaL�+�;�����.��r��~9����E�oۡ^��3hea�ߵ���mel��s�P4[��̂�5�����*��e�~"�֖-�Wﺺ|��<q/��3�,,/��S��[�t�lz����Z�ʾd�7 �y�B"=���L��H�'���	��_�����o%3��P�ďms.+�;�}Sv{^��R)f��Á�M����{������b{��ۅ���7���\��:ɝɑj�ց��<�;+&�ĳ^�̬y9,���t���E�F��A^	i���*K��u��F��'��L��++�z	�A�?��p~��M$�p,X&�r�ٟ��IL/-|Y�c���ZG����1L�P��ӼM۪�$�A*a���@t>� ��nd�� �cv 9~Z��G�^�����m�e�e$� �eZ���O)܋����H�����OW��u�sO���̸G�ێ@W|q1��՝�|(�2�i�C�=P��:�Їq�:8j���G�[���+�	7ı$���FM�P��Ҳ��"�	���,�:��]��N��2��h�)�O���=�L����x��M�up��i���2=��O�:�Ѵ���H��n�=�_̏6ĀT�.��������"�MIf�q�4����j�Tnp��>�T��Rsh��q�
p0%�D��	�Y,0D��\'������:D��B�7@3	����)՞�����=v�:���i܃�T�z�T��r1b�g*5��ŗ��رz�X�\��Z�<"�r����K��x�W�,$5�I����	8ǐYQ)����88�(�-ġ���w4�A�ͳg7���eiN��gN����:(r\#�B�g!L�k_=���`��W]/��^B�z���j=�JU� "@7��r���7c�*TR�l)�[
�|��.�t'����bd�d����I!�Rc{�L�Q���j��X���?&��,�ǋrT	� ,�
(��H��Z�n���2�"��]
򻟮u+�њl��(C<�����U+���X1�X}�~�� �����f������xO��C�rQ(H�{�4�ǎ�D�]��{��]���o��@���Y��z�e-�Q����F�3 �=��b%�O�$�e��ǵ�C~�a��h�tT�CO��ڷ�@�-(�jf5���R��q;�c�PM�ԅ���e���`�ï:�:�������ƌ'AΫֱ���귱��S\oW�l�`��֐d�h!��m�*��4i�ض�3W|�Q��Gf�s2|�>�)n0�T��c�k��M��6�@^V����a�2��4��M|Z
��E"x]�j�$�o�|M�Լ��2�KQ��"N�)��^u*�)��Ÿ�?m1�[K߆��1�&�	����Q������'XV��t���L���w+e��$g6���g�s��+�D��2�bV�;[֡��pq�4O�����0L���-3���U��1v�{��H��we�n��XԔFP([Mf%D���b�,��D���jz����XiuR��	X��Vi{�v����9M�(.��Ge����ٝ��lM��"�x�o��TW[A��zCT�g����B{�p����X��0��L���TH�n�Ņ�.�k����-+k#H�^B&V��h>�����Bu�/-lbF�}nS����rq���S�\6?I�!&Kk��Lzد�JQ����|oɗO�]SM���8�L�Н�Xˇ�\#�O�И���<@2�~S�㕀��Z�L��UQ@8�p��9�"����
HD�G�C�2GU�]͠�� 5�J}�{�Q1�^2k���ԈP�� �a6�#���|�΁����Vc(
,ŐD���P�ǜ=�,�L�&�u�	�Y'���|�-F��ɕ�QnEt05�z'�ed�޽���qq~�D�o����+("٠�p�`��|\<G�������g���yq� �p"h%�� ����G�ѸLH	[����z^ƀ���~I/��יP�8�H{v�Ι�^$���r'�U���\�� Ex��5)� /7�nj����l��:���׹�B5�#�qA���У��}簌#��X[R�����w���e8ͤ��Ҵ5��R{DB�A.�i�35Q������R�eߠBs�p�x�2!��3o�i@+�&�7���s9�Ҩ��P��ۏX1��V�Eg���lqR�M��
ȁ�`�72���C�{�\j�+���vf���m�r.�T��������Ĳ��}�<.���
L_{�-���|	�W�6�z1����w.���Dw�Ys^��+:޿ҹ}�؇�����ǣp������L �)c�e������ް��s���r�C�d��)���.I���3�GrBKJ|��"ԾYx��V~�P	f��N߇�1po%Ne�����H^"u����H� 2������U�ei~�7�x�ڍ�Sz,*u�5��.S7�G^������#P�Mw��0wwr�LЎ�RPf��LZ�����j�ۛ*�1�Nk8�fP�� 
$����~̤?�`t���"-Ϯ�4N����J�=�݀  �"Z�a���Y�T�mؙ/k+ �U~�������t�i�g���zz3�5���r�A�*�6��Oo�K��e�q��sQU��K���[\	.rT��x���=dփr�*o�s
��%*X�$&�m���!��h��2��+�3���!���:7����:�Tb���!4�͢CƠ��\q`�P��:fF����+_g��� i��a.�<�O� g@���!�60Kz ��px}D��@w����\�J�T����Z�t%C$��7�wߡ`��0��~�"e1憗��,@�M����cm;�[��f򿉧b=co�}�mDJ��(���I���>�$W�-MΒ��*潼?�#Գ2ה���I�D�T���9� h�u��`\tt�e�H���0�}	Y/��?�l�ƹI5�������,n=v�3Zw@�o�4�aLVڲ��'oNߠb��Z���Z[ffұ�X^=xi�cd� 3���	 �����Z��zr
�oh�.�H��!s15�5�Z��'(�V��A���H��ۏ���_`�?���iZ=|ïi.�� #3G(	/��!���ň�-�ڹW�'� ��J�*�0�>��G����F>�t܁�,)���tWn�X��ԃ��~��5���n�5�g2 堨J�ᇳ!;\�DF�Z�H�ܐ�ޅ�ԆL�9ӫ�5ɬ�n�������(F�P�*g��gƱ�b2y��3X91b����zz|7�S'��
ݜ��Cb�Fq�W��2�0��u�猨�{�T�x4�b�r��ey�d֩t晝����Ӻ�_��F7LMi�H����TK
dk:�E����/��$]O�h��!��*�:��sG1պ��+T�~3o`~�3���Mi�Y��/��fzxl	�u)mcL���#��5���o5�5��,�CW=c*:0���x��WDL&/:-�����^VC�����t}nOt��B.�Y̎#-������<���$X��,"G�n ��RSc�y�V{�7^���\.�{�.��IOn���t�Ei������Wڻ�H��:N�+�P֕V�啣�UFu�O+q�H���A�w�����"���l�Q#�xD��f�R�k�%& bΤ�Ig�30J��RDD�4�Tx�bi�
�ըy�XTO�ph5������ȕ��S��\�r����l�zG���,�UP���/���d]{�R�#��n���Ep�~�c�P�{��G�j]1��FfԪ+t�I�=P`���}4�&�NI�����0.�Ƹy�~�8ٌ����âȤ�����׆�@��x֑�+\[k��F��<nձWrx�p��m��Kc��wt�@��_τ�����P�bO^����XI#g??O)����T5Q����
aS�kp�2y���7x�� |�u�T��j�Оl' �n9o�1�KR�+�v��]���?�i@�(��X�o�q8Bz#�k`Ls��Y4�Y�.���Җ��<��q��uگa��8�PKNu!{���' *[���B��#`��ұ�,n.�F�N%_�R�'o��JO�O]>SQS��q�˾��'p2�����j��8{s�vB}��V+i�X�����ڊ?��ɰJB�:<c����GI��	�%��:����e���dV��c.j�w˚�se�4d��9��mX��Քz��>Qy�x��x��S|qd��)�u�/�^�~�bA0�������I�վh/��U`[�@005��`p��*�q(a?���P���v�$Dj�ښ����JTV0��]d�R��4���f^���%�f(ǐ��*�����h�� �뢝�hllŒp��`ȞG<���;+�/)>�_ur����_Q~0��}��'4��4|���
�d:!&M(E��҈%�����1OY���-�wh�*aK(1RV�z�Z�4�qP]|���R�F���<����4��#o�v�E���Ch+0.��@�X���(@�L-Y����YWPU�Lz�j�b9��K��� '�qix^�Wi�c��S�1J鳢N,�CO�����d |
hԏF�l"T��oH�Yfh�Fk�\@� 3���g.�sؚ�,�WZ�0g��
�}���d�ӟ �iצ�)_e2�}7���s��׎7��
��&n�1����=Qc�x���HB���Y��4����#׺ۏ�⬸r�F��=��{�[I�|@rbg��������/�X��@HH"۸���_I鱚��^�ޗkY��e�����[k{тi�s+
�;��2��G��$R�T����	m���<�S�ZSן��h�}m\]���q���[p�u�\��)!)ZF�H�逆x��T��r���������_��|�Zŕw%����k����Áã"�2tB���8(��������j	�:h���b�t\�vi�����e�����i��4�����b�l�d�	�*��d	 2q���~���fv���E�^A�;����j�X�K�K�{�	?�]�%1��_Ʃ��`�c�d�c��$���ʲ
ˮ����J�޲����N`Iʨ��-��o����2�s��DO�SX	��Px*�����Q����-;�ŮH� A.�f5>�����EZ3�F��������$wd�t���Xti!��R�����	V��I����6�L��?��G+z���DBEޒ��[:]�ɡn�P9�)�̮|��^��ukّ���o�/v�LQC��ud���[� �P��oE�1�z�Y�py݂wx����3�%U�n��2}�߂+�Z���H��������Я�w��������}�������ƭ-�M���S�'�̰?,�B��p�5�6,g
�wT4,�R?��9�-8���3<�Cy����Y�jA�ä+��d�/�`��� x��7iֶpZ͔gBd2���B��L1�;��v�W4m���-pv\[(�û-�M~t��d�m�[�-b�YY�.����׳!�To�d�4�%�]�q��2�ڼ�U�����~��V;�lW���'�K������a�^9�t��.ö����ͽ�#�����n�֝������C_T�J ^�6Z!v�,�X���߻���6ˆ4��䲅.����ɷBו;�&���ɱ��
�jS+���B�)��sa��1OBD�	��G�Ԇ�,�N�!�y��|�u2S����;�@x����o[�T�x�l�p������{���xz��wC����ߗMD�[�:8�+�_,��Ō�ѿ=+�A�y��MZ`�W�Q�+/{―�Mʆh�������C�v44-�*�=��GQ).��df��B�D�r�)�DE��_*C��d�{�=qD�p��ϖc�r9��L� U�kuQ�T�im��R
\!C�EF�I��c�S�~�c;d�L	� jP9���������U�t�� �j���ϴ*/��������q��;ɴ��n�'$�c^���	�G+˭�إ������WI�v˕�QXS�B>���K�?�CiQ�-�QOZ��q�y٠i��J&�����WAmK�5h@�j�W�0w,W�r����m���s�;?��$4�!����I�Pt�;��o��b�L�<��FqM�O�>��\c�Vg��kp�����f��Q3=��0�3�}�u��tm�II��9��(���mN��"��]ڰ�#�����l\���t����}x�MP�b�̈́dV��1��-����7~�X3��~)q�*�����{�m{}����$�u䈵�z���D��Z�'j�GzԡN>-��O��|��I���c|����B�f4�H&S�}z�m�D��qg�=:N�ޑ�,P��Fu`W<��sƮt�H�_��b��\�f�8�	�@�B!�&�r�w���PR���w�>.���k+í����+�$:ad9ᎅNO�ۭ��u�k4����Z������֍Ȉ��s@i�������Z��f�B��������^�<s��T�E�iDj�==�]p�O��k��~� �>Y�0��v]sE�Y���q�Uk��9�o���A��Q�]6�!t�%�jO���8}�ɢ?�$�[N����:ܽɾ�[�|\��>l�F�Ý�F�r��丣�	��itcN�J"r!�~��t�=]/#����Vxl�@ 1JG�
�)w���<8߲#�HcQ@'<5ǚ���� p|���>g�,�Z��Kd�D�Sr��~���`V��J�u\HQ�`�P�������Q������2��5�	����II�q}���v����1��S�	5�2J[������:ɺ�u��fJpYb�%����&�O=������������q{��L���7����\��(��z��}1N����P<�L��C�
\���S��(&�������kܰ� 

�����i(�g�ox�8|x->��_ ���,	�eׂ����'���GrBd��+��T/�.kt�>����M_DU'���KH���moj��R����V�Ǒj�;7y�R¢r��	�m��}�6�;�Jb�����b ���ʭvA�N��Q�<��jH�}�DUO�5�<���'B^�$]Ѳw&L�<���՟9���ك�+�˯���1��FuK�55��XY�8������{:k��bZ��іeW�d-�,��xW���i�Hv�kjƋ�����1B�ཾ�	>�H��y�$v�ZDJp�t�������3�|p'���)4WK��{8��{�qu�A���&Q��|���f��/��7�����'l={��و�|��`��1tT��I�J5|?տ�740�O�A�ʲ��^?<��!��$d�S����)7k1���n�]�=��;�6!h�u���N�?��yqfD�)���g'�db1)���J���$��ʞ��<|�+�y>O�4K��ˈi�^"aB��&��3�������<y֐[�����N�g8�<�wsp;0[7�t�5{�w� .����6�*B~~�7����#a:�z�:����xl%<�мz�H.�]1���)�D�`�l+O�t[�ds�*v��|�+	��["t􄕩�����J���]�|]�]�C��n�4Q�qT����6���Ǻۻ���B;a�4������ٕ\��hͿ���62��}����XQ���{݇��E~V�d�!���0������{����[���0�����1Eܫ��lo�e��F��& �e�P�p{΄���0��Fk�v?��U]7�]�n�`�E����^D��&�n���ߌ'�6��"���;��P )�ޜa	N��T��$��\�N&���%G�10�u���# �s��kRq.�\a��6V�#^�M	Ds�zj�w�3t`G`/\r��h.�8ܔ���ҭ2M>	�`�����} �{�K�D[ͺ��C�[�� �vd�2(��f`�L���Bl�g��_����i�^]"4�c�6w��P
�Xd'I������<r�1cޏ&��h1:v�}�JSQ^���J��c����}5��a]77Ԓ�B����� ������L�K��R������Y3]�:��4ߌ2��/V73��UjFo��|��X���u�v�9���R]*�l�	k��~�-�2�x�Hn�ַz�M�87upO��c�_����,�M����V���d��U��J6�9;��A�aM����!n�ɚ,�b!KhO����y�+���f05DZ��E�}��Tp]����z5rK��s��fծ��yy�����-=)������n�I��\�ˢ_J�/�\��5C])^�l1MLTo��.�s�!�=�#�K����J2�����f�����IK��+~�l�a!��79Dv֓u}��xő�[g���N�o#quD��j�>�筩5p2̂�%95r�q�E���.~�vgZ��%h����[Mj�c/��%5���ŀ�No�t�o5єʝqW�+�}�Y�H�ۑ冻���W��
@S�,#�#�S��æ�w�'#�}B�
�����j�t-
��;����f�[�*����7r�^�]F��hۥ�U�Lv�	+�5p��:)�����ӽ~0���B��ޅ�t���l�%��T��{CX�gf�ۃ���Xlc<��ֶ�)fٮQY(�b���	4�D��\�#*]��V�tg�{�	�g������EHtR�>��:Gd�s{�EoA�� l��?�� �y��S���� �'�\�+F�����I�X����BS�C��S�r\R���K� ;�p�!|��y�b��bl������@
�#�NDN�@JQ�C�˸$�&�i�z�q�,7ϊ^�������@ᾀ�������A�5s���*�DX�� �X%�oHS�����,�fzYZm�O�=s1%��2�v/R�̰lJ�߄%�Up6\V�͊,����>`��D����lV�Kyy�=����qG��d��C�������ik�(,�|�
��E��QbmSR�x��Tįף��<����5G7X}�f����0�o��>чH��m�}K�h��Q��q�}��/=�*�#Sh��`�w�	��⾻��ǧ�"��]�'sXQ@��@�Yȑc��|��:,3�8�n��N0i��	I��~.Yf�j�T��tk���z� ���'YE"t�0�`[;d��o/e
8k􇀎ATJ���0��TX�2sby�������?��l@mT^�@<�p����c�<=ӹ�����j�+����c���EV��w��p�"a�baK���x|����[D��)!/�]��ِaE���☤�+	��>}�ώ!�r���X�L�~ba�!'"\�����~//��:���$�|78�;��F��ѳ��_�C�_0U�}BqA �\��LKjG�����_��T��5.��	z���!��b�^2q�T����d�>]�?�O��w�6��S�PF)��Z䪾v���.�7a�U��ҡ�G�im^�'�����XZٌW�c28�S,c5Y{R�H�x��I�6-��<��D�i��1
}H�R�q,��%f�J�`��;�"AF�`j.,��Jm��F�qԆ��!�\^zNMe��j��;�w�0�أ#���]���Q��?��,})=b�^)��QSg���i�h��H/�'U{f�4�K���v0NEm�`�e,N�2c��ءČAΓ��D���u�#������4�!�y�_���� vQ�^��v|�
�K�e:��a���dt0��{ϼn���VP��!#H7�i&L	��'l2�X����I1U�&%�i��<(���"E+�#�p!aX9#��߈���v�El������B�ӑN	�MN =6u�0u=k�
Y�U��^.�T��~�xSW��F́�P�_S�O�onD����W���x���]o��Ȩ��Z=�5��v���W7��9��6M���K���j�0��7ji΂�"�g�D�l�M���h�_RYXq=b���D�<�����@3���Ņ�<OM鿮
��I�=S�1^E�#�*oҰ~�����w�W����L
��O����c�m~�(
,��>�m�3��˷DmX˒5Z-��Qe��b2+�&_��φ�C�6)M����r�^���4a�*kB�Xk��I�Q~Ig("���|��R���<؋�(�P/�e\�o����tj�5l�I�#� �;@ۗH���-��?Q��R��ǩ	Q�`R��%�CjCڊ+=z5*��G�>�y�~�[g�����Z�Խ�v�%��v$ {&�*�Ui���w���#�w���d����Ox`)ES�ka���!�D�_���R�l�ә/����V�>�~��3y�&�M��r��K)�$kK�I�B��ҷM�bȟ���c�?3�yF��0.X�8���<�zʝ�lk�5�m�J �7f�[�e�O�f֎&�[fPV��o�RW�smb��q��p��ӟA4�f�b��I�QyH[i�aKq�"	0�B����7p1l"�0���?�d.l%��\c���f�?(u՗Ɏ�B��ze��8�8�\�f������7cn3W���� ���m��u����~x�c��o�i,���R���t�A��:5������17�g;}�'�!K�L���)�A�8{�H���m��O�O�`0�ƍb����MjKBp-�rD�Q��{{���h3�H��K��u�?ל�}���+��,�<��Z�1�
1~:���ǫ	�Ĝ����cP�_�9��|8�޽l����_6帩�ߺ�kv�λ��o������\�ԝI�d�Sjx5��Z���s����7�����o�s�~��6�Ǒ���|�u[_�+�г�hJj�0^����g�=4"�N)S��r����ne��i�.]U�ڊ�x��:E����{�o~Ax�y4����狅�_�@^�?mLs�(�@:�k�E����m��5_�M�rXiM���PFW	ݓ�`؋ ��K*�8�+�*�<�7��H���!Mv��F��Ҝ�?
:`�}����a���L���^��H>�� 2V!+��PL6�3� 4��8�E�>�� ,�c̛n�-7�¡���̻�Vr<T�<9�$�ks��f��K;>�阏����a$�BuP4 X�' ����"h�x�.uh��R�z~�5
s�bE:^O�x,��R���X&:w�\G&���0��Zz�k��!M � �լ��#\P���ք� \�'����4��f��G�����P�s�;~���Z��]��iN�é�yB4���+�ꤜ�ħ�Ġٔ�O�]_˙��!�]��v��y�S�p�a���x�e�ĵq�@�b����p�ܔ�����n�Z����Cᙒ�}a|s֙��J��%Q��_NqC<4w^�qN�nt~���K�`e� �_�`AF*���^]@���cW��~G�9�3�P��$�;Ҷ���c����(�j�H5�SbJ��PÒ�@G��`�x�eW�Cp΅�㷻l��)k[�iP�򠫣��
�o�x�	i���y��{��n����(z�k�f�E@�'x��XУq�?+lI7!��F��F�t�����R61טؘ̣�R�[�J�J�Fs�hЬ(_��e`,<) M��X���z���\�}}�)B2f 9)��yH�hk�k�\��.���W9��&t�(�a����猇�LϠj��AS=�ӵ�U�KP�
�V n+��㒚W�&'v�i�{��}k��&&�`�)�NG���e2M�*!g��À�ښ5cVFl=ܖ��s���¨�C��Y���&%�|����Rq҅���P۲.����I3��4s�6��G�ܜEWq�&��K �,�����B���f��ﻩi���h:o!+N(���F:�B���h1�:�A��%Rۚ���}z���TuJu6sed��m4��!�kZ$s��m���͗E֐#��n�b47�Բ>W>Uv �� ��Z?қL��ʌ?�fq2����/���5�N�c��N�f��~��q5<D��RU֬L��L��f���aTu�m�S	�'�f싥҉aR�(��XKu�X���(,s3C3I]M"����]j!���O��4�M/y�����TH�~�W�<M_���R��s�b�bB`,*��L^�9��홂m,�n)Yը�՘Y�����I���q�b�#�y�f��z0����y�2�0;LN6A�Fn��#�z��1���j
7����'�cti�7��qV��o������ϳ��MF;.���cC8�Y��{��d�� )Nł2� ��xk���>V��Z����,_��"�61[�IT�W�������` ��W5`&nE��h�ĭK�Ͽ�b���)�g�l�C�W�v9.Ҍ�G��{�oQ[9*3�o��^���gPњ4�<���!�"h����=���%ŵ\Xyq�	7�E�ʥ^�מ.D�%��� [y���Gb�W��F��w�Q���+�\A|;������ ��mF����8,hd®(U������}w�"~v��1��&R�#E�X����>uB���^C�{W/S?ٹC麧�pʕ��^�^y7��[�Л4͊i��2����!*A��w*,��S�(��ښHț��}3��������Ő�5����,�!�����"��K7�'=5Q�x���'�O0~Sڒ��aX��o����=�k�l�h�@50 ���K��^rx���v�~� @	�F�Q��>�1|����lI�Nhx�t���A��ީ�� *o�bG
�S�����I�l�hB�Ĩ0��ߜ�[�zRO�i�Wc��/!�X�N�%<���0�(aI�og���K��N4�0a�����5k�-��@��Fe��Q�ڮ��3��m�� /G����6�{���K94��qq+�*R{���-��c��� DgDMRr�j�kqL�֟��(�Xsv|�����I���V #��le�Y�&}����R��4��Yz�|��w ��'H3u[��<j.�u..2�%��pBwG�����/�e����[&���t?M��P��aA^��r�J�<fQ2�.>,��(fzst�R:�`�n�,�,�1���t���;)�khX�7����NƮ���>φ�B�0W���5a��5r�ѱſ\gC�#���BV�䔄����U
I��Iց��G���=$%h'y����+�Z�G�	L�? ��Jz=��x�m!Ŷ9����C'�Y�VB�&S�2�i����c�
%�tp��3�۽����
9��*�p���c���|M����}q�ɏ�|R��Paz����;�ӑ��� ����{RK��Y�����&���	�C��v�{�F}��-�3	�e�y���:/�[����J+H?�	�(HD���Ю�z��%�M�a��Z��ޥ�9WFmJ��,�%�go��^�MS�L����?�R�j��C�I��=�	uozW �����|���UVyTE��6�   �B(ge�Q�q�F��a�w�w'"��u�p����~{?d��̜�{�8�&K&��hMD�R���N���>�TW���� 3�2������RTR�����yV5�Qo��f�U������GQ��|�w�R!��CW�؂՝��U}��6��o�l�'�	�bq�7�����cM-���y����A��o��cv��D��Ȧ�܀����J�A5�*`����2�|�-��F�p �������,�l��EG͇U��b�i�BK�CG%!^N�gb�j�	��_/��i�V��ą�����P�Yёf(T�/��J���i�p���"��`�ཿ��Ly�$���ߚ	C	y1��\��c�l�
]���s�c?�Ul�Sz=;��r��c�̘�!H�p���I��6B.]��䘀�Э��A�q�(y�g�d�|a� ����R8�-qP�#�A�1��ҳo�f۫,�.�o��4ƪ�
9�3q�Bg�L	^�,I0ˢ���wX�g�4�$ivq���dQ���<<g`��W�t��]�����zgi\�r.z��l��D����й��þH
�c�9�+Ǳ	o��[J��=2v��c�i'�o�Hw���]�o��k�1'��c�������c/zI t��/��km���d���%N��9�湹���vJY�GF ��-��	B��"xP��"���y�r��8ԏ����.Fy������h���h]�m��_��J&�~*χ���.a&���������8�`�G��f�5�Mi��]O-󟕡�z6�]j�!䋓
��KB���BB]�G��f_�P��ʶ�X'	�@�:"�R��iv2^��cQ����k�Mi8[�+���1(�`�~�H�zwՠc7=gu�s���Z��R�f�F.�Q�8���5�������-v��	,K��}�������Q��������qΈ`>CTL��������z� F&���A�p}1�^���51uf��gmr�Czb�Dݷ����U����"�|��o�a�)ZY=�@cK�.��U�9^�2�أ�N!�]h8���I�褸��W����ĪAO<&@3�x^��"���4��W KzD��0{:f��$������=�+�~�� �]vk�5��ۦ��ÈG��������ˌ|�Pw� I�4 8>9_K�b�D�M�.��R{�r���Ic�;+�k��n0^gaʩe�F�}�2�&0f^c�_�:���ğ��L:f�+Ӝ��ȧ�G�yq�Wd�a������TS�$pC��2����+po�F]��%�.�q�Z��q��ު\Ir/ё/X`1�7�(3s2<�Z�4t˶ ҷ�;'��Jo_���'�/�E�1���u�����_�|�#D�H��W����?�XQ�$�?�`��ĸ�|���Z�����l�g�������xa���ot�)	p�P����N!�����oW�sF�Y4��+�~�����r��j���]��؀����&�@u�U�+������$�%��Z���r�"��M��o=~�=%M��b::Y�*cz��4��a�d��
'�!X�ѱ/���4x����[���<R�3��r#ydm�L�W��CÆ,5�Á'�*��e{aJ�FC���[����ȅj��g���͠'�j�7T1y��!4���l$,�XƮ!����M�:��B@��; ��;�<�� }���n_�f����xV{�4������jm��č���6=[n�����\�����zք���h�N	�9�����ɱ�S�"���N!�F{� $W���?u��{�i�=��<ʄ5��m��W��9Ng�INh>���#k�Ɩ���a��<�������^P�({jO]D�X̱���Ӟ���&�01��f)�sæ���-��`8�ǟWl�;����̭]��f�E����="�%0ۀ�H�nZ��<����m�y©���g¦��g��N݇ѳ,�^}��ǃs6��� j�72��sD�J�q���L�|�����`�����ȟ�����e�V�3l�M�_���m3�Ȭ��0���Ӧ�G8�2�>��;N�UTO���hz�'��EZܪ�F7�����[�u��w����{�{5���饥��o?�U�Inx�{t0/F�6D4��z����b�O�}h&΄��V�Ń�����]�^o,w An��0q�N�X��0zG���Ќ��l��֪��$����s[�i�?K:;1�X'L7<=G6ʽ���a��i'2�>%��]9i1��{��l�Z����mRlNC�|�8e��D(G��G�Iy�b6�����b�������?�'GQX�#3mU2.fQ�� ���Ņ��������� ^6&S�n�	�	d��;��|9F�2>C���^+�Q*:\\C�*�PT�<���[�A�ӥH�g�gʸw�(�L&A0�d\0�OiK> ll�!���ʿ��,P��*�!��:-1�*C���<�\���'�L5�e���aw�B�<Q�5|a���>����k����+P�/Ӆ~p�1/6@a�4���>�?��]���!��l�o�]	M��U�VC�_�.��s�H�M�y��D��
M� H3;��� T���NQ>z\R����zb�A^K<t�n��a��&8�`K�jQ�ń]"��jqF�
��,b��5@��[�p|���.�fll��H�U�/���?�+fH�:�G�@���+z���Xy�G^�rx�~Z�5>,?�����T�ծ�\�`4���� 8os;�h��%"cp��� �I�P�x�v��w�"��Ť`� ���&��7�F�9�ᨨMڭ%�i���i3��p�+8z��e�(�j���3�(� _��E���4�3F��M�)��t℀���� p��z#�n�����E�='J�\�#B�s2G���r ��Le$[�ק�O��E�Wۑ᪀4�%�8?�Ro�C�,W�Y砉��ǋ���D~�������)��j+SY�^9�a�Nu�%�6pVQAύY@������)E�Fr���҃4]LZ��z�%�,@�jJt�D��/�<�Л٢ob����kz%��R��~-h��W!�ü�.�#o�k٪�|��L�K�9W��6Rh9S�`���J��B��,��":f��oڬ��E�X���w;w��--.�s�����=�p޼NHX/tb9�V'�wk������\��/������V{�.5%m�`���5Jp,>�m�	C̬�k衱��*3��f!�E`V�ɯ��|��\��mT�5<rO���QP-k_��v���xj�{�%�Xq�*!/�]���bd��s��ԩy��O����L�=��!($�ĀW*^���1wCv���~���z�KB����?eT�&���?K����5<!����5�3�x��fTY�0�|&�'p 1��\u��u��$�'����G���h����Xכ���� ���y�^�QP\��/M�A(-N����zB�Q��C�-��\{҅���q|��A8���@��.�ڹC�E33oxja���y6M>�LHܔX>^gW3��w�3��M�%-7��#h؅R�҆������p���' [뢷�U ��@�0 c�؊�``=x��1p;Jv7s��@�L��맴��L�����_���U��E�L���;�vRT)�]�#U
�m��mC�d��� �կ����l��!��W���ͱ��v�gJY�_T�υS	V�z�Nq��-���r����p�7�B ���>��<�ybOU�ۤ$(��h�����q���x�v`v�x��@�y;�`�J'�k����û|���!w���O�x1<#��`w>�im�����2�w� �����+	Q�iR=#�5r	yS"� ����Z`^������$�aO�
�ր�]��.P�0�.���?�c~{�7{�	fmA����N����������A����ß�1��/��n��<.�
��A��EW!Y�)�^�~���ަR��$Tb��fI��f�mg\�JP�U�)�}�C:�O�E&<�L9�*m;5&.ɬ����\�a	F��/�Y�gd&}6��(�I��c�,wS������D�/>�rt����9D���>�|
Z�U��@�LC�(G��UKJ�
>�zѼD?4k	�2oz�)��-��H@��)��xp4)a��ӽ�^9��Hm�J%��p#���Ύ�xV�__>d�}Pk���d�s�2����Eif��Y��hmON��s�����pE��x�Bq>8iW��FD/��H�����ݴ}����|����C�؟7��@~���^���}��A���~�-hb�MIGqp��_&L�	� \1bˢH������t��#X�4��25��z`�P�<������j�jH��L�f�ׄ�
�ՠ��qM���:�kP�)���z�F�N�q�"8�g�k�;�nU����Ǫs�z��Qb�����Q�X|8��-^���x-eU/��[yU���n�.��')�@���/����7U�$Q��j��Ij}���dy�쩋W�O*P���~c���P����P+a%��y�w��8�`�c;��(��S�B�%t����?d띠�?C�E��Mj�|�u���)1	R��ȍȸ9;F�DN,l�+W�	�+�$��j�R돑��`��ժZ}�,f����G��o��g��� )�P-U����Gp�Ț:��+e�G�_I��^��d�j;��X������Q��!� �S��L���1�ŋ׮�{�"	�zL©�~+Z`}�?�#ч��}�u��@�ai���Vm��6��9�6������X��ذ�T�:���3J7���;�_� ?�xc��K��(?*�?����k_O�@og�K{w}���+��&��Z����s�/��G4�o�fcg�1�a��:�/�Ȑr��m5�V���p �m��m��a�;unH�qX4!50�"0����c̶Zh�v��HQ�JW��l(�J^� � ��J��~�U�#������l9(ړlU���Q��[o[7t%/��z����!HԀA[���?��<�"���MV��m=7�rrd��8����[�E���m@��Ћ���3n�n�
�[��3X|h�w��x�RsWq��]�m��5:	��9�%���T@Mb`���c�4����誃��ܡ���`�z��k�/W[ ��w=n@~�y��	����X��c.[e��9�T��-����5I�n �>��x�2���@cW���f_S�W�Q�l���<Ua�}Ҫk�-9,�}VO7�����e� ��=�[ST(�S+X�k��ln���Cv�G���r�y��*��G��M�LT<�|!��|2��f��d�&�p`��v���������j�T��N$Z��$0���]��t��M�
����Cci���%<*��=ҵ�@��Ш!#΃!;p��0
!�����#ݯ��.�N�k�⢂
=��@���d<ł*���r��w�9A�ʟО@�ҢmAc���B'���~|����V���S:��S�s�ǘZ�4�.pc�`D-K���RZ�7���>�T٫�AC �b~Y3J��@*�t֯OG�W�)v��0v���rB9�S4Olo�k}k�V-f1�g������%�H��k�>&���J�|<Ta��nݥ\	��SN��$�("�"������
EB�x߻T���=@�*:���x�K��_�y�a{V�{���������!vᘬy�,��z�]/(wl
�lS�S�����g��Ɇ�Y�K�/T�B_�er7�O)��,:���P�L��ͺJpY.�봸��h��l���A��������ߢL��}���M�$&YuW�0/�Y��.�0�m������a�P��:�;�����_z^�4����+����Ǒ�rj׏�1��~K��	"��Ϻ�q��L
�Cy�.F���U�?��z�^��y��.<�-u��F�0��,�"\Dn�U��7gq0:�.�i��Ƴ��:��Wl�8�<��(�X�q���YINRj�I��̃ۯ�����p4��ev��W��FW�0E�������{u������z.+y���	8x�l��r�`���;O�_r��C'Ӗ=�|�}���5+�6���d�Cwè�����+�:��%5yr�v���O�e��d�Y8�Ӏ%�{���D�p�A�'�熎��:=U�=(�6l���_)`�|(M�q�n�X6��Q֒���pLMa�4)�d~���Z ]B���W�<�Yy��o�$R����q����Ѩ�Iƶ��z��O��ms�i-M�ъ�u�g;�:@0G����Y�P7�-�#��d���yv�wUgY_�Ѡ#Ĕw�{��Z@wj�t�7��V/�:ޓ���i���ٮ���ä��a֓���5��u�u5T�v�U��#Ɍie��^G,����j{��#!A=|�M�P��쀪,����4b���,���]aM؊�s��*n !<>7>���Jy}�5�b�KO#K{���3Oa����A/���ViZ1�� #d�R�����q�x=+'��@v���؛��'l8q@����䖍����
4��ɑ��Fy��OY��e��L���1<�q��)dԄ������ƙW3R�C�N���qB��q��f�eKΡ�NGVwMr���1��Q67�
(G0rn4��̍F�m���k�+���.����5'����g��?�_�t��cs_0,j�1^+0�i�m�,�M��~�[��v폗�E8���B����`��H6�-a����+��.�#��~V}��$T��4���c���2ڭ���~Ƞ�k~�[���1�����۰G?ۛ���_o8�=d8:
f����>]�/����X��i	���&�t��o���!��=2������"\��Z�p����L���Wt��T����0F���M1<kx����ci�[o�dcf�n�X4����@Wc=J(<]|��䏫Z���X�q
� ��[/c2DDH�U��X�!�tS�	Ba<lr~����9��D̭�".�QXO��4�;B�O�����KUw�G��i��rNC6%���kz5�
53/5t���3P�����]���m�|��o(oe݇&Μ���~%�U\Kf����ݐ:$�/cuIQ����.���$�@�O�G��0	�&�d?k�A"3���������T1��`��h4D�>A���I���<K�5R�k��ы��u�+��]��b6���J.�
�M� �<�HF!��ܘ��8^$j��P��L���=�G�zU��a��d�������<	x�"���G�<��D��'I�0a����:��|Y/��g�oEsfta��H^�\@�B��b1���0�����i�K:T-@;>M�>�yG��O���u&�
,0R��ƌ�#-��K[oE\�{l馱�K�
F5(�ٜ ��i�5j�U7,i��N>��080T����r0(*�Jt���"xz�A�mv��k{E����%����.l��O4`cJ��� FK5\�"�����N�]�C�ie��D��+�T�nG��m�*���ǞRnN6/3l���@����]�X�B�#
V�r�׻��.�/6Pl��H#i4KeZ��9{#QF�"m6<��18Tji�;� ��0Ө��r!\|\�ZB���Hn��;���k[��7*#��8F�,Ϲ�T�
�V�i���ߟ��l�+.
��H��M�(��H�Q́��Z�	�º��HD0N4��;�Kr�T�#@f�1�W4��O���4v�Q"O��v�hP�G���dq�$HxLR�$
� y�&tfJ~�.�� �rĎje��'0���]!�Q�5�s�3�H�Q�xtփ(j|���<����0YvQ�=��15Ȅ��@�&��y�*�>��Y�Z��T�iL`�P��"�s6�'�H����ϝ�_Gz��C���hxحG�z����Xzs�y��Y
ѩ�f�^�?�Xb¨�����?�wH4U��XHb��KO6���͔4�y����z���j5P5�(V	�@�� 4�>Y�5<��}��[]%�|�ya�:�U&�+~^��8qZQ���FC��ADU�EO�|��m�us�Z&Ŭer��ع���R_9��~PH��|5������y�Ow���'��I��w�Z1GU����6��Yd�˳����o	�7R3��b�D���iG�i52�pVގ{��2U���H��pM��\�Cg��|r\�`?�$׉����hҾ_�6�eS���ЌN�⶜��d��`$.�Y��mymp"]��vx�~�;���|�f��QQ��A���"��=�0��(t�`Ԍ��c�^�- 5ƵڦGo���MI��1����`d�mgZY�o�F�!Y������;(�
t�i���'�=���őل_�,c9کVǬ/��̅��,��uE�\sOղ70���^ɚ)�Z����b%�u	���WzVO��W�y�m�����:�K�5 ` �BͿ� ƑR��l�L"0H@�C�� ��7�;�����Èȣ���{�s��%���)��sqÍO���{��$ć��N_T4��$S����;���1=V7�<�>Cb�tn�H5rW�֎�Bkf^����#w��w/(�xC�+�3�Pu>�f�G��ٖ��5��c��i���1�^'�usl��wnih�8�b�9n����/�Y>B��������-c�������b�>��/;:ӕ4�0N-����Nhj����:'E?��rLe�zJ\�JZ���e�P��(<=���{NAJ%	��X
�F��%��=�g����z����@������I/=���"�*�m�^c�	3�)���Ҹ �YTbE.�� �(A.���xP�ۙu�n�i�A.���o0����$���V?���y��Rɹ{�N=�����b�f5��	�0y#x>��7�.(������S��I?U���7?9��ؤ��B�2Yܝܸa��!�(֯��	d�h �.!�qd�9<^p�C:�tҞ3��>�qy�72����䞵 Hp�lF������;g�U�)�����F�kH���wq	��f*[�<�X�k�U�xވkㆉ����,1{z���� ��8�9�/���� ���DO��O쯌�3u*;=��$�	}��]���Ybm�C+Njt3ȃ����O�hOn�ɘ�W�Ƌ��S�}����л����)2Mj�M�~�!�~���G�6���I��v+�����K%�kN�A��"��$< �������KW�P,
=_�o��-
�d���m��=����D�7.�H?5���Ŧ�l��rxZ{���jY�ܓh?����c��!O�
���1�O�����c��T��n�����K|���K���s�nV�^E��|9̃?7���RO����so�p��y�L|�����D[����E;�	�y��PH-[�F�ƅ"is*5��78x�,��m2� �B��r.bӿڏ^�L�:}�}��mQۅ���C�۪ׄB��_��Hw����t�@*���dss^a�+��Z�=Sh�IH�rJ���.�J� [�*%��Fd��*U:����I���>w�n�S\v�MY:u����H	�7����U��@�� �/�@�Vb;��o2��)��G̅��۱8Y
@Y�����I���v���r�(軺R,��7h���xTc�$7`C=B1�ɉ��ӫ�PERD����k,X���*��(@�Eo�p+285��b8^��x4+���z>���Y忥����n��"��e��UJ��F�2s��hѰ�fz���6V��PGj��CLa�p�ҠJF#8�8��ly2ȫ�3&�ݾ�]�+t�f��0��C�م���b�]�8r��%:I���D��:�5�u�oD.�'r�[7:�a�#̉��R��,�����#���֤y�:���.�͟���"�%9���w`X�����>�hjU�E���#`�~��)�3tp��g8>��*�Rm�$+S���W��3����[��G�C�jKM
�,�8�AH���x��&	BE�`gv����Vm��3NXy&��!@Vu�nK��&��q6���-�`Hʊ�S�S\q�0>��3k
z�W�a�d(�q�¼1��-�?�%�u]<JL�m���{�U՜��%�ىh�e�׊ŋ�y�_�-�@�>�
g"��J��P��I:��ف�C�=���b
`]g�7&nת��a���v������`��>��xp�wo�7�vsU���'a&W��P'�t�i�QӚ^��]�xg�H}�ot	� ���q%y���,�$��;;_���G'+�X�3���j�"������(
a�=�H!E��uz�Mt��ۈ��ezP���%��W9#IOU�:ǚ�%6����ºS�ϦT���g��ɛ�q��=ެ����$���t���U��zHdZc����V���gn���dR�PA��2v��j	F�텕��]�4�;
��Ng�]���{�;6
���"C��uX�U�H����C��+�Oԛ��e_Y􏇭;�{��H�B�Oyϛ�.2ʀYG��Yfz1�WЇ�玍��?��3x��эO�YW��S��$E������{�6��O��������hqE�V�����|�*g��}vYf�|�7����j{N�zOz��?H��E�e~���W ��z�G��8��rת�L^��IOw?�x[#?���O6�䁘=�d�v'u&z-�ZҌ�d:��D]~��ѩ$į��}ˠ�'}�*m��+�v$ق���;��A�Y�H"H�B�E+&ks��K�`�$����4yI��؀()�o�P%=^�y��:�gљ��<$�n���;E�sj�	��+�r1s���	�5�i8� ��\W���i׵_ݜ�9S:�@�)�fX����}^5��s��C�R4xL{dfh��F��
�B���좜r�QMl�}=��)"�b�S��6��<ǟW��
���'�J���ٟE��!��c�.X�)d��ve��E��ШZ��uD%�"I7�����E:�� +hd��
Jƚl�fH}j9������Hzp��}�J�	}m�@O�|2��f��3 ���"�����ܱ�s��w�Z�3V�tKޖ���@���_�1R�(k��Au&1vpCS=��ܣ�(��`����� c?CS}���],G����Z&�\�,$v�=	���S��[��ʖ�lGN�qbM.�%�[m���9���Ж�\�� E�2�#����إ
:�:G�|���>���g����f����$8��'�v:��ʝ=������q�:�%�U�,���o�2�g2K�V�*��ɵ�1���@$l{��R9D��_������%�ZQ���F��h�$n�:$�����'=�3��Dq��(�&q�p��\ ��A��vl]}�6ɕ�RF�6~T��4��4�O�� <���۹8b8���ų>g�}F 8u&*����0͊�Nz�OJ�t�>n�������t JId	WF�-��/� �3�a�&S0������Z$��;ȜBh�C4���8��'Y$߮�����6ƨ�Y�H�h��%f4���l�U��(5����^.{:�l�+�#�����_�M�EȔ�q'nG9�Qfќ>I�١%���s ��8���=�|%�HDߊ��//ZF4�	�]�����U��.�t=d8�-�V�v�Cm�K�����o%η��S- J��"��4/�[��Wi���v9�G4�}?v�o0.֖�K��ҳ���Z�M���	��k���U伂�k��cY��^�Ty�0�v�g��D :G�9�-�[�c�R�)��w��{0R�v{�N
7c���Y�#�*�:;�@�W�,�� ,�t�\Uo}�0#��_qP��0Ƿ��աإ��E%���z��%l�*�M�(3��L�V�ǹ �4Z!s���ܣ*�~,��]�ָ�u���U�"������g}26������u�F6!2TU6�
��s1ᥡ� [�9� Ү�=�R�:Ԩ�U������30�ڇ�BD��;��6�K�9�ӣ����#�M���V�n��
�-N��<Vu�$�q�H.����A�+0�2����d>�![�9:p/��1�.�q��_ �����2��{��E4P]2�ʳ����7��R^tݦ��j-0�rs�+�!|�/�*T������3w�Gj]�[*	�xrY;jŨu+VP��g���)<a��h�>�z�z��4��2~pp�f^`�A����:�a���WA���}P�eU7����=6F�c��:o��R;�^���VSU�Ƥ��PS�[nf�q�?�C7NV��ܐE���~/S�kEpM�k�}cS�}�;Ƹ0��J%a�1��;�"aXl������i%$��3���!H�{�5F�[؍����'���xsh����חVܡ��˲?^�[�l߭G�'�;���}���V5�>�lgP�w�N|C�a��=�a\�m� �/�<(/U[D�L�#ϓ�� �~yU�Y1*#�_��0�l�q���ժ�P��Y
֥	�$B�X�d)��!��"�m�Z�dkV�oV��^ -��U� ��iv�i�.*$�2�Bڴ�]KOrK���U��d�g /S�V�˦f�D(c��+Oy��#���>	�yc}f��_�H�HS�ϋ,���C�L\��5E7J��<S�BY}/N��&�`A����y�WV����L�PRRUSX�}�^�ֱ����]������U ���vW�y�J�&�,J��S
�$VƼj�`�/�>����;%�9�lj��@���i�[L����&���VpZ��h�ۊjR~�؂������J��_�A�i���xk�4#P]A���?(�����Y��s��p�h];�݁�ً�J%M;:\]�YcZ����ؚ�u��V����v�P4R��-!(Z��eD�%�I֘O��>]��I�h����-�����v��܉���9Uz��P�~�9Xw8�7��ӈC�HQ<�*2D'�]F���.��`@yB������^���������o�_�Xs�3�N��0��w��-b)^��ϲzȴG>���Dd�,�4�)'�8��`$��G��A�9 �o%VڮT��`���N�w=�=\�����;�@�	p����OL��l@0��+)��I��Ы�-j!.i�X��1��:�#6����Z�����%#�0���֪����f�.��Oc����-OpJ�)�*<O����H.~wo� �ҟG�︗��@g3a��Zڍ���s�bp�d���Q���w�|�C%)�I��Hw�*A'��ʔe�Q���j���� �h,3L������uZ�%g��l�^��&�*��%l�XIp�ĝ��ɋ9\s��!�K�6W6^�Y�'X������My�?&&�C���<���t�e����U�TG�k�/ƞuN�6�p�3��Ȇ+gb�@�l��4�>����[-#m	a��Q�`��#^�32@(����E��}�+nf�&�����5K�RJ�C���,,�7f�>�@��^?+�p�C!�N��Eg�H��Q����M�,\�6�sc�.�Z�3��`p�3��%�(w.X�%TH��JP�wg�M$+�/�r����}p�g��s�0L��Z��/T�/H�v��4���M&�Q�g]3��lҐ�H��bX=��uk�X��̣�@�:g�d3Q3��$��k7p��m��/.u�j�;h�*Xﳙ��l�8�i%
_��cY���Ǡ2���G��1*hͳ���}d�P��[(_�Q쒷oU��z��d��ȼ��>���J%էi��k1z������xGoD��9�Z��dE)ʑub8�Md\�@�f�iy{����� �+�	��h�d���f�����w��{��^3ac@�Y�H�����j.��%�Ѹe��7V=$�:	�� ��:[�0����n0�M�I��(<p��]�> �R����؁�8~&��MS尭-�-_����)��w�m�,K'd+m3��X�n��|����g��A�V4���w O�^���J�M0�r������v<�� ���E� 6C*��[���r�	?�Qa�#g���f�4r�+�y�'�5�W�i�"�T>|V�,lt1;�x&�}�{nvs#��d��	|`�<�6�����>��+�����(�рO�Du�`���s��������r�HA�낹H8�:�!�s!_��E/�����%@Ul��%�d�;12����"������uz��d�C|��&]��.��q��2��2Ȏ�U�L�}[�,gl�6�}b��u����޾2��8-qT�>�u[���|	m��|����d�b6���9M&�A2��'x�,����.�=B�RoU����}�{:���
@RT� ��*�(R!$+Ũ|�l��?�C�*w���6����R�--���)��KHpu��/wۏЩ��U��
��?0j��P�/F�y�Х����M�������Q�
I2���Uz �$}�2[�q���̎��^v��At�:W��m��k�֚��uA��C���Ih���ke�,�<\��ߧ�v����:]�R�J����Y09+u�=~{D.0� ��Da�k�Y����R����%��S$XD�u��B��IX0�]�'��f~�m>^�9sz=P,��ЄJu�0�L SM���i��?�5��P�p�Z\�W�>¼��7����
"y���q�iw�5�����~I����=JS^����)�bS4�X�)ݰ�?���Y9��Y�^�9�|�'t+� _İyQ��U9��>���^;%9O.�p����Ys��u����Y��DH{�h��@� �,��F��~n�������zTϖг��S��(���U��LRǛ_Fӷ�$�B� �p������D�E鷋����O�)���I�=���\t�q"B�R�֋$��s���_�ջ'Θ�Q������5��s��)�Q. �n��b�cc�����ۦΐ�T(�	��n��V�hN`�t�q���v%@y��?ԧ��C�n��&QT���QQ��v�f�(n(�H���R�c���^�[��]��Y�vL���s�6��Eg0���9u��P(��+��Ҁ�v��e<ك�,�1~��zހ8_je���J��9����Y�T�9�)y������Č����Pv[?�{
����������z�Ɖ0�!Rb���`F���F���ɿ��=��4�!�C8g�z�҆=�������`s�C+j\QT)�������b/���#�ZA�	~ o)sYx�:��ώ���&b>A��_�$,|W����$�~��S�sn���� d�ۖO�Ĥc�P$��c��l�޶��!҃����i�O|Y��S0!�g��~��"��ex/UQ��u���:���e���E�&�������&��d`����3�V���zc����'m���1"�}7]���q�mS�g�0]��O��'x0?�����S��*�o�[أVDj�a������\ǭy��	����m�@������N��"��9T_�-�?��<�K�����5�I��)Ǝ���f���s��;Y
a��\2)�q��|a�5Z������5Wm������\m��!��2�>�n�F�{k����^@�9�J��	>�e�)�a՝'��:G� >.4x��&�A��f���X�{����v�^�=��"hz�+%��wǠ6����g,�&���R�>�e�{l��,���T��^ow�ps�%����\<-��9\��x�����Z�PR� ��νˮ{�ڍ�u�1���Y��\[}A�
Ing.�a�!y�O2%�2�X3'|f-2�MPe#I�V���i�߄	0nq_T,M�WiJ6p��'G��Go[6�X�R��1y�C�/��Dr�]������si�:��(p�zX5�+R��B������!�|)$���o`��	�%�k�><��9[O9;!:�<S$�O���b҃��F�n�^�#����L���U5���S<d�>�ґc?o�-��w��:,	�~{c0�1#4C��#˂vfWn<��8�)u��Ņ���XX�}s��[�B��vx}��wŸ)��a�J-pXy��'=D���F�S��#�t�jӯrmol��٪�o�Ij�2��&;�����LWP`����k�d��l��@ n���C5�T�����"	`��Y6 Iq*�E�����z���_�5D5Ln�d$�ނ��J"ſv��}|*�Ѡ$`ygks�T�;خy��P�ۿ_���o6��
5v�4Nr�G� v.�, �UPo��';�������t>���TQl�3�\�z A����ʵw�y�e�;<-'�飉͢�TTʉ�|Qp�I�*�n�O(���9�4t��C��E1�x$�����+#��Z�\n�!� ]��&�
��T���1��:-��K�¥�)k�\���u�c�)��9�$`z��Y��T,��
�u�NzJ��e��>:�K�~�%����e6k"d��ω��̰M�Hxڥ�R�l�T��i��h��5Lg�~�������ܣ�����.&�	i-�l�0�����D[dDU`�";��?�~����##J����"�eXTE0<����4��5��n ��GBC�΁ug�{��g��`��������lX��H���`�KzcJux;mϼ,��B�6%�J�����.���LK�oܫ/�fD\E���.ӓ�({I=�ٛ����*X{�/Û������t�(_&q<��8�	cp�i=���1��\y׮�>�:=�@�=����K!�t���2r��'�걒ie�}o�MO1iO����Z���0ֱ���������.���a0�R�*�Bϗ������B���_��̈́۬�Y�R�C��ظO����R)�9�,�Hk�ŁD��Ć��3HLF���Q�<:+ť7>T&,������}���R��ޝ˭��o9b���A�*zl�hs�`q�'��I���9�5ʖ�Q,��c�񕩩��a��I;f��axaM�Z��� 
�#2qq�}�'>��:��&>l�$���P��=��굽ތ��H��a����=�U[U���Q���⊰� l}�U��ʠ�hE
��2r6I�S�`��l}�p�Ц�OZ�-'!�)�qGUgZ����t�1����U��X��N+l,��_�v�ۨ�&�5��C��_��8���-���43n��O�o������R9TF%~+�Y'�NSD��-&Z�����.!���FqIE�0��l'ƗY�6�e� ���W��+�s9-_���l�R�<f{�}�n��`tĔ��NB�9*?��Ð�x��-1��)8��@��:�*[T�%}'��{ȫ�sTD��;m;�w���]I��fKNN�	~ �S�`�)cC__�U�a+��7�L��Ws��Y����H���eI!��Z g�up�VH1������"��+��(�'8� �D�ؙ�MC�� ���P���Vn�/`�!����t�/��j�g~�>憍�h���r�(Ե��N���$�Ԯ)���?��$j�3����*�]-�6{9B�lG���%J��側,��9򓈒᠙��Vt���dSզ��mJ�a�.0�D�<����X��}�m�>M��!RB�T9L���M0O|�ET~"b�?���G�BVK��Fk���%j2�d�790��k���������<W�W7t�H&�ݤo�%�e�������k%[NYb�D����jk�C@v����G�l�7�$���
����~ �m�V��E����Vm�0n���1�<�G�H�ҎpebS3%=���B�H�</�_��~G�o��<�?�"��Oz���6�h�6:m��P�b6�:H�\�jC�U��Ϙ�<zJ�[�:�2��׬�l1��1.pB������)r}Bq��\v�90�����J�ȳ�c_�ڡ�u�]����i�؅�������Y�S�j���Om�؇��t�"�.t���9`�Jh��`9ӎ�&9�C���`W��轊o-���Q-�auii��cJ�9�^M�N474*@��l���g�F�Q ~�W&��n��dZ�"dR����EA�~�9{�����!Î�v�Y��a��5�窥o�*�ll�����,�!q�RZ����\�i�W��/�
�X��A����?O�U��?��l/p�a���Cf
M��!�	��Zx��rJ�fHP���F�~�`�qd#G�S�e�7�"���U�t$�v��/a���Y|x��᧻��_y^_d�B��r�)t@);}�T���[���T�L������n�f�6>Z�I�1+�	�c.!�����xV��ƕ�t�(�ձ��5����W	�� ��2���۬�������Yw�R�G�V�(Y~�挵�-x&�v�$�t
��\(\2@��,�fs�f�,���H�p��OTd1�Zt�C��X�1Sˮ@���E�/Q_�ۼ~mJ�8��I%�E��D�Ro8�ҖT��.#�ئ;���t��<���id�4�?�d�;f��x!�?��h��ӄ��a�V!O�Ih
t�Y��ܦ�7�6ן���n���&P�L޽Kv%��c��B���rA�қD	퍴ó�������	��No���P�������2
':��e��a�ňs8��.�ߟ`g��q��|Hٌ.}��Ϩ���H�һ�/�^��J���� ���|��X�_�?�pUoO��܈8���J���>�f?�|����P=q���V_�&ȓuS��7�!�K���Ӯ��'O8D�pA��H��S���#`6�,Q�&P�w�w9�8�����W8զ�m"����cw<�i�P�n���0o�0X�j�I��_�Q�@��|���p��w�,��T鱣v���+ǹ��Īɥ��9i�5���n�"O��浨����K�`ѻ�s�]< bz��į�l������J���H8e\ �&�yV� F|^s����-����%T���o�Ϳk~�M�Z #h���%/?O�>ڵ�d�#}�����`��](�!G�l(����M!�ll@���b��|���Q��&Rnȥߗw>�5H���G���/�W�蜳�h��?�N�Bש����+�ϯ4ڈ+�H�
��ɢ^S����L���mh�4�Xޔ~�����x�>I5��+D�-u=	
jj���d�Ͷ���Q�K��
���>G̺�l?*{��ům���u;�ZgܮEH��i��'�+�A�Fdˡ����	�����s�^�1,���1�M�	�����	j�!8�!P5�C�Y(DD���WT����v5cw��+���w�;8�U8;��~�	)�KO�g�xmr%�Oc�=1k�8ڮ葌��V��Y�h�����"̀m���]�������햮K,���_��M�E�Я�r�E���.$Ѫ��H�Y�6wE���e)��Ef��@N�=��6�B��q\=&�G�E�w�.��r���5�VD(9�?@^UzK���5��cH��'�Q�{W@_d�W�jJw��E��`�W1H7T撍$�/��؃��G@��G)
TN�ڭ�
�,�[���;oў�'A�.���ĵ"Xyqf�tT長���ù�� ��$X�$An����ћ��LתFa\��\�{r�_���+���Q�(�� ��"��'�-A���$��m%�eۖ�a�:v��"�s�2~���S��x܌C���-��Y���W�;ӟԶk���z! ۃ^�Փ��PE�)��� ����uR�ǥ5��D�0�7����`߷~���?�ׁ��>6��!z����f��_��V,3�Meb��������/+}e��Aw��8�W�c���Ps���0W��C@��H"���Dǯ�T����L9�&�{��}�ߵ�`��-(�;�Sdҁ�C���t�E��+8`�/>�z�yig�G9�Q�-ȅW΃u�T&�4�'����'Z���To���}̭p*���V}��L�N�d�'���Q�Y:�3��#��J�Gks�OI�~QjjuxO�;����sKd�T� ­	}P*sW��o~.����Q��ű9B���q�Q0��0�Ȕ��7b�A��;�q�ޕ�c���E�K�F(N�1h�a~&�����@���ǌ�h��!H�y��l��v�8k�t8���$�ߙ�`������ A��S3G�:>��≆R�	�%׋��,;Y��*oW��I>%���W~YOX�⣗���}��q|18@�@�^�U[�����l'���|�J��SHO����D�F�i U��7��Ì�*��/��_�6�ӎV��O�Y=�1��3i������J�H�ʔ��}?q�l��p��=���F�����6ʍ/M���vm�����i1k����#8�ü0��=�Оn��oPTA���
�j��o�f� �?�C�Y����j>F�/�\Pc��݄$ߙ�1  Ǳ�g��D�Da���x�m�;	��i�(�n���xj
�?!�;~�>�$7��Q�ۊ��v=������+����m��!j�C��+�`����T��-���NL'��L*�t?Z���j��̯8 i���M��+s	���z�T�����bC��p.�FHTQ��H_yv8�����g�4$�P._�@����χbh�1޻� O7�	D>��lL��|�!E��Kt��W��ld�Ȑ�Cƥc:�o u_qFq��Y�� |x-m��]�"�:�:��%�%~��#�+�U��hS�}��ϗgX������"���l�s�FR��������{˞^0�M��\��e�u��ҁ9F�9����O�������!�]C�vv��n֢L��ɞU7�Gw�v,)ܯ�x�V�G��^��|�?B�n�aȕS�ͧ.��dԚA�N��_��צ9}�>�f�
�Xe�w6�ə�� IR4/�,-9�Z-�z�+=o�'VA��5�� �n�3��VQ��G��7	n���v��[Qt&�I���C�&��|�󫻂�9f'vm)�A�F��,~ ����!�_a���_��`v��r��[,<�T򍙱к�U��	��c��S*+�sZ
�O��bh��yH6�/������R��<�X|H�B�|��c��Y(`F^�]
�8bA��h���/b80M]�w͓1yVZ��k������V2�MJ`7yδnأZ޺����E��5�y���Ѱڮr�~tA���*r�٪b^��I���iL�-�pϬd1��&
`L�w����!�,����p*q��ӚZ��9^BAc�AZ�P̗~x��h�.G�������+�;���Gj���m ��@!��i�7�Q�� ��ۄ�o�%2����	N��%7K�4��k�.'���V��բnXh�x}c׎?�INM)9R'yW�ā���0귁�V���Q9�V;�=��@�Τ�E_�P@��׼���s��Qq��Kr/�5 +a��W�Q.���[t
F���v�dߤj!�`^��M�L�|~H�����Y!���5�e?-X]8f�9oV�cj��\���td��f�F�B�A5���R�qu�Q4�tj�GKH�o<X(�-��q5�HZ���O�	��2�8��a8��DF��#6"��5u�%��E%�ͩ{٫BOe�H?/C*�Pw��3e3�l/	_��G��˦k:��	ʢ����ǔ�aA���Q-����
�h��(ƢܛJp',N��i�B��X��B��0��I٭.��-�s����J�D�!e�àz�X�M{�S�-�!U��v��D��	���V
]�˗Ǽ�7ȑ�o�
�9旙ߦ�d���I�u��hUO%�oo�N�r�%#��J��GS����a��	�Fd<������@�o\4�>�D`�jA��K��v'`�J5�:y!�?)[���:�ے5l 1sa�����
yJ�z��l�'�µR?iZ��]�8ׄ56a�}�G���ӏ�
*j�'�� b�7��v0qش����X	�\ x@����ę��4�0����s/.����88'Hyx�p��{��O�j߶� d�/�X���?�fYĤ��y$i�_��Q)�甴�vmX��[��
b�|@0�њ�L����	�4�O(��k�&�A�u����z�{��nG�C�tR��.�8%�~.n8�B_�li�?ŗ%�� 8�{_��U;�hl7: ��R(�_�0D)�ί��>4R�IV�������1V���.J��5|!��ߕ�0�H�'PlJ�<��ǩ)�\�Xw,�� &�sK��c[�7��[���cZ�!5r�Ќ�}+:����	ܦ��V�\��c��q���K���pn��FR�TXvx��~�cS$��ǿ$ua;Y��;{����`܂E�r.�h�ӝd4Y2p[���p���m����H�f�$�ޒI��X͂ ������QI`����>%_:t�tF�>�=?g���m���D�trS2�{�@�����W��s�UT��D�����G*�c�*ND,�^+�z��u�~��ğ�2@�v����:�z�귕��	�W>��4��Rc�%g��%�Idq�a36�.�ÿ-�	�.m��1�ҵu�p=k�<�eoH��+�lD[M3��қ�@��T$6��[��X'���7�B΁]���&7*x�/����"�A��/rT�X��[tG�>�*������V��4�:�B=;/֖�6*��6i�B�0(�I�**�0�tuu+�勎=��$��~Z�9�=��,�D%�n�݋�
tn������3�D���\ mD�al<$�=��ܿ������*i:���x��9��=�Av�b���H���i�o^�m�d��1�*�hZ1,	.wC�F6��z����u%X�����W�w�IE�OC �s����_���^1��'�+]����?�V���ou�rY��f��* c��