`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
JmU0tzxS2HnvMUHn1aYwqjwkoldqWbkwPaKpaDVtaXZmX4Q9izenTxU2D+Kyal4Ye29lC/CBV0+X
Pl9B4b8d1hQiqm/+q7fcmSPnczQALy5bOsf1tC90sUlUOB5aY9tMSjqcTMdY4D3hdYbB/BLbk/1T
sntioqw/5CR6dOJik7BOwAzf57iep2b5qoPFt7bMKqbSRGztHPQ/+fErVOw0Un6kKg2BPdXIPc3P
ZlIvhr7vnMV3jmkHjJmiznWpVUE+RaurTMR+iRdwZ9AX2+ZgDzrRO8Ifw7EkWqLXTZSVeK+EGuDi
RhzcemcuySaZKjcf5UlVl0W7bFHdPWIvrIHstUd+rrMxc0YHx0ID7HzI4+aTcWH714VcSuOO6RJL
j9x+je/POZK948LlEdXjXQEn/xKTiLeyHebM0fm+unfDb7A4fkPQ490JOurwRCqlwcxpHBEtbO/B
g8rEXWVX1S10SWSPIMEOX0iggx/pnN+L+QI5O1YsZYq1FH+Is4w3BmUioRjNPJckFpsECkt9ghOJ
6ng+MAqJ8t+KIMBvyws3hsNpVNfOawQwrJL0vuOYlTGX09aEqj06i3Fffba4w811yfA0qFWEqK8U
4+c47s/x23CWpQjSblWq7+bcP1wAPcGxpuhUwWbfK9d9S6WUNcdwIGjkrtV4tDCTZtSM7b23YWht
ICs8xpg40MrCUEQNFbwlDuLI5btZtE6bzwcmxvES10URS4kI+cui88xm+DSlS3RmvZEuAS4OREYd
7ANr7erC51BGjAUSkHk+RPXAdHI84Hn7DsE4oeCREJ+aEU/dEtUNTbyfhIs9crlD9eIvYe7n1UPj
baBwUdeeZS71iSx42+rB8oysvJp8r1ODnfBwqwtLCcgRryxJJ9/wCRyDqoP2808efwSrX30Sqs1g
dgYb3JtxRTCf+Ptt2OqjWSDbslj+wRBZnC/LBe6iWyKN/9H5omcFVv3fVd+UP9ii44bqF4iQJNv0
/Bt57ZvohND33LAPTkufe5wHbGo/ySRadIZnPVQ/L8hlCsOJhliDk/aZHyqymVHKNgi/Nzur6Ve5
EYmfh5jMDMCW97L09mhP3+BymuVme/ekUpxUQpkuYSp8LQ+aaMpYTJXhV8icfgZdWn2/Dj54Xrbb
TVbvHELD+j2xF1/hgJpUvwFUbIFdlXHLkSeEN5nNsp7QXZMr7VBLm42AbKtfTyk6e9pvCZH9n7Wv
beOgkL5AbVfxvImrkO8WlaP/nwEg48NTuN6t4C6Ha94POZtBDNNP5iUi2q3puV5vV818qBFzD6Be
WFGTzh9tyud+S+V+MW043LBthtBEcMcy6dp4P/NdRUyHx1Xvxh+Yy87HLROf1KBZ+KLlDgEPInT7
qFEqeFtHXnkUzlotgb01Tc/oEnAcLMrV4DynOL+hpmXrWV531GG2AWoAutBEjzbFaIskX1B6bUPx
WMFRdYDAiSDPhdh9pRwhoBQp4hU4bwxlk8d0l12132tjF0LqkmvyWRNuJJZUqCcO2g00Uv8iM736
2vr5VKFe62XJ2D5hHyRac3hXdUzZ2Ykz09FrI75NZmJzKq0jiA9hZveok3RanRtUL3DtR7ZLJ6A1
8kewoI9gTlUpOMgxgos5e4JDmh5v0crWO6EikYJ1fxMdcIY23R4DLUj7P9RU9b+5o29h88EGrjpc
EuAj7tFdWlMURCTy2jR26mRoPHsIEzNrPC6qOOQuL17yY0CYO5lltX3RZopVU3RQ3KDQHs2TSe1U
+AV/0j6agsiL+sYE3lpgD9EolnIW7d2nUcRsvsXCqRzdOFru/ewGY1NUKP3V2o1pxOORNcwZSGhe
n8a3IxqWIPkIx5pqSOz+Xz+rq7encfxzCcVBf+RQmleXxLAosKhFFTwEvrwTmiihrCIjo1nu1ver
6rQfR1Jvx5xpO2tTd4BZAHpP5Rf6ImQ9uPQGuWIGOc72gEQZ1Di5qtaINhjoomdUXHrqhVkJzGw/
B1yl5xnQHHKM34PV5mLEdR835P6FgrK0JUukTDcyzi9ny0fV2QdFnEMsKfLcDuC5DUKkNYfVAfl2
h3YjgAj16yxqIW9NTHgH5RyDrlX85mJAofelZXsB2aZVVFHx+v2j0AQ+7BkFFOXS9iFVWjcbFZC+
+YgVpiCPb7TSe8MSpBNpaBK0sO2A5JnYFLncLJxpQemXDRGC4bGUWJBu7Bg+S89aTDuCKgCaWnUj
43+QObukAbhmj/iGa80tqgi3ehZJmNGdNYie/V7d3mof8ZltnFleU8Ey5UfSzktWWf5QCp9S2GAz
K4wCfYfz2Dv+DAn0Se8e9rNwKkX7VrNgXKiLaj1pFvXyrxcP5QwK40qzoQH4Y2FEXX1aeaKHYskJ
g5XGsnAAwHwIw4agWlW1u416cdWmzrqIzX4za8egwoGyP7lhn1uooPK6JhgLgSrM5SbFPNxRavtp
c2mkdHbcv6p7o8q08IGaJepX/lLHIbf2KSNWRlqzf3N+KE4H3LFFsJxvgqIqxYWBaqTK9lo7ue7w
9i3Lv4zrsfDSwJx4NDeZKzOqg94oBeYZg+5wvrjNdYtWj8YTs1DLapMdPbDyPv5dphDpgiLLgCx7
FRp1kSIAvPcgxBOLESaq+qZUvgAheawbTw03Nt7O7kOZ2pJDDajHIrAilpoy8ENNsa8XsACLCnVd
49s7hHA7weBr2x6/rEnuWEdZtFg0ltQEzdCblbjj5It5JYeiaF01geu32X3Q6Wb2wZyvHfaQzYDk
8NcScqd3GptFXhrYurgQWuCj7VM9TjxUX7TJyydOKVjGMCluBNchOrVFbGs3Adp+IvbHTMRHEq33
HHgxWtPpnsdYFmofq313UOTEqNJ2/afRjAVJqrKBfmHprBj9ln+hlukqQ9WKewtiyzR4LzuFkGG/
sf5QB9R0q+bxWQR4IY2EJOyKxFgaDU/7q9A7705xxYLqSwUUKpgVsCFSMzGxO1Ug8b1QOwJr5oda
O2w1I8CJ1fWPZ9/N0Lg83MIHB0vxYrGV5OFXMZlIfIV1BAutP5HcGKcG94kL5nUD+vjmlhy44dBR
JjFfF0RVdllmszvjDz0M2DW5HiPUT9+dclmZRoBIPRtfEFugGFo+yyvG7TSIuEZCDVANgozZji58
RdiCcZy6SoNiOMUZislnvb0wyBhTes/SLeZhsI8MVuVXWslkhMe+hYe4b+MBtLIm0Fd1JQSWGWN0
EFk5qTsytUCu14b2axJFtapxcT4prSQ0oJDsLVbA/4MEfe8suTY7d5XUUsEgXVhPCOIywhxQ78xO
FsXZCG/rfSjntlLJMGdmBBoXkIG+nfhpC1NnQMtWdCkGRH0FZvv7eqolEe+uRNiTVdiDIWAhW8VF
D0Gs7px+hBGsf7udC+kuMEfkfJMEmNd3AsQzvLYoSVW5/ystuqmMAIXO7STP93bkMLgvlMYREJOe
9x24SbPID2NmELvnKe9JVrmZ2Xs3it4suKTfpObhuEAMFqSAIOUWLRmLVxg1YV93aVEsKGzXLd+q
Yw3vBvBU08UcgwaJlprvKN+UNBNz1S0lYypeeUQAOkyg2o5u3AAqUZhcvN0z0nTdKX+FrLA+EbfJ
hYt4KZIgnkitdljkB+tluFTfjfEZbSncFZgpTPuCI9HUKd7ykVytAj1wzGlNkRWQaSQOv8E+2dtL
lsLCpcgO4SMZNBElYQ+pD+pimRozBHGjEZElf/kD13GPc7XErZdKly6ZrOCfyHkMq8PNAtdkYncv
cMxGUycJv/plsTuwG416r4ZRzUirPS7GoNvWNCLZUh8fVLuxiCIhrgCxOIWlvhV+N1KSX8zozmdj
GDVyQ8YVRTlSVOAavtZiM6Z1A8woNM524Gbu87UMBFuPcP+/5DSrF1v0i2tzFBTs4QmXyxEL6wxc
whj2XnPIUBHdHsLeny+8Vmf429FNnZyAvRHLjNcbca35wM9+qXCN+O5yBR6MhhId0Sxj7GC8Kxkw
xd0r1NM88SVuokTm+hO4/Wo7qJPfSEpBTGKwghbHn1ieTtAZz1pS7Vbo8V0+evRJzNNe1M1CLgqS
Vdt3DV20kE5r3lEU63mG9WgdcgT8Rb+sZg1grNFeraanG+R9fmzrRYSAhsr4C2jUa8iAkWqDFDPq
/qxf0tTg43tnZwq2FPfetSzO3ps1ck3wGCL9jl8T17U/QNPkCUVHbYPLTnBHPzJRO8OJoedsC0uK
BH4In5eqFZfA1mstlcLEGWtUA5qS2iI4kNEctB1Ry6r8z1KZY8bRe6D86hrpVUNoLtcLWSqu9iT0
IU2RkZA0qGfKP2EbsFBAtB9x+LG9XzWnY2fw9UihAl1Iw1CCGv5I/v2YLg/JZET3FBr5NGFMoy0R
XQZGPeGzk3lyoz9K+v1LY651LqHzegZsJDhs29+eTIqC/sPb2+AsD4ltpnOhlwnAGkOfHENJdowI
7qGLcgHlMRZTeIrJzKZoh5N+sU/hFLKUZypXQM/Llq505liywUCRHejqfcWFRrVrD1LA5Vo1ggmf
GPO1TT34dT9t1gw48ngiWJLpzBpbnUSDQjpMAOy4+btcydP7DzM1s/xeK5vbCVg4pPPwPCaCDtZj
Qzy2GTA8pNdXr59mZLR7ykZtFPfC7COUl1zqDOcSnIIxXe+4pL61CYg+PYTeUJ8E7oy52lqrH3t0
p+wFyn2lyQCmx/hMcqBjlpCWrIMC7eTQdCmYh/jIdktDuYs5sRHlKGp1olYtbCa/bxz15ZpdJ1+T
RIxFI+F4tGoXWoesU+6SmG7Xecv4TBIwJC3ay5tD1hCg6DjE7jpK2YHPZndJ9eyUMWmKOCsM8Ojh
jIR/MtCszze4bgjQ/mKAKtazT/EqBBwj7rVzMFFgnwkVUVU5xhY8i1ift9DPFrarKrbinftumqmY
kknUCx6797AZ9g8wETYOha+e7Dz6cFUifmWc89SsCWXxsFYpd4mkwzmT5SCBXdvPWo9Ymy7Y2Lwy
yZ5q3Lcj+Rrz62d1Dzy7gxST7eI2ZwBqu3RiY/XVYSlOuhL0PQNdrY57d4GcFZvojOYHNqm/0SsJ
jvhergaemg7Vy6GHBzByMZumuMhDnTK3o+6S/Bg9afSig3g7enGJwnLDEii0h0LLuoM7SWpJAfbU
1ybBfgRLmT7y4OFdV+LpQwuvy+Zk5T7HqzD1PWXNua6UodOm0rtOfkuc4VvfRMNb5e0oMM75Fosg
8Vq5thbOgr68I9xt/BW2qbnZD56Hhd8QLEb5OgA0EWYNiaW3b9fZrvBxpWRdD/fY51Ki69wLCCCt
0Yz+jHEI1FveEMP07IP/Y2nnZHoanpvkbkNNGzix3c8qoCjV1Gtt58OiCerkuBb54Y7wDaiKEJRJ
Iva2Ymbb2AZq8/Uq38bl2LlffgSHzY6jLvi+XJXwRFfGhVU5cZU9l8tEKlJBJLfoVnNNstPe0LX3
yb8pGhPLjB0QqB5NhkXhqm7qPqyLq1UcaYiBFyVe/eNJ0KAcuKEsQ96UuAqwFDEjq9n8nn8Aq+C7
FdXXsSs6mbD+ittQK/3/biNK8SfLSjtcb2Cw++iL3tGcCxousyBd0X5LrLClg6ejJM/uFLjk1kuy
84IkznWKp577JWDOrxUXL8ShTegh1Fo3WqnYxro23mOWIJAMuGlEJWSZU6CzVZ4hUVPhJDmiB1Lh
AcFG7Hpl+ibEtYqv25YsMIM3/5NCfK9JhQqj+OXQYOj4WEP1IIp7q5YTUavASFvl/ER8OPmresyY
ZjazhMBRwPheKfzeWqKQbcKbftt6ePQQ9wAS+JVvG+nvt6tSvt0q1bNbWIXLp2gVEiNBlSq1zZZt
QTXxruQUhVuYW2zWAvG3WjTxms6bmTtVWNV2k7F2yOUsKUy66M4F8NuVOvalFwicvXqQwTV0CXEr
f0PdmJ8cVk6AWyJlv+f3bm7VK5pi984LGd9PStLtrt7p6A3f1rB0oADXHe6BaczHBuuwSSs+W9yu
b8X0OalEjOEK4LWDTnSDRLrCXKBrfLdABwEp8ZhaSua8+iyQOhHbMQBZrkHSphexXmBjN6eBwxYO
Ht3AEV6YMuYAv2zFYzP+f4M0nCMahNOSAjEBZ1hPBTZkAR9l8cQQXsc4bMHN+qbchiswPMdl0o0X
tJTWCTPsivzVLaK+D3JlQ2kI3IGBYrKUfKa8JZUkjHYgSfZmB1LKkNjugK1BDwBv0TH/3HB7K5gG
LIv66RRP61RSETMBMUKlPRI+DM+iJlmabUTo/2xGAjffeCaBJt8vpfrhgX7gnqtpzp69cnz6wyXw
7V07nRGXC+OH4fulGffXnqHIuq60MnUub672+UWNpZPqgb/g5AWthFDZ1G9il9FC2b7reDNP4tT9
rNXZ/5SWPnuO1G0eTK8ONxy1Pf+aV6JIMlxD/WqC4vO293ojHAsXtOZnQ6eo+EfAOXjBYIPMt4i4
TVBTd0ViHRhvJHr+uzixWgPXAXd/uT0oTgHDjr8v7gM3osPpOsZ8sOlyyFU4gEl3jBLVitYAaJ5a
gSVJ45psWItoFzK0rpanhVhdlTOtvfqndcJRfpdohMbn3ilDv2M405RYFAS4ddADv/K0s3CNxUmS
KjQTovKHNmTw6RoQ7tjZMXt0CfcMHf1BRpxYMGYik0WhBjrLYlCYOCk/4Ntvd8P/uJLxOk4LyTPb
GPaASPOILHyd+ffQUt2IRpt/LHd/irhLiXDXcWzsaZ7EHUHOiVNpN+j248avWuAKgXEyAOGlSzLB
dlwyU9yctxtQiK5sR3Gbro05PPaZsDdo3Pm+FppsflrM/4kFdpUr0r0vmKEPKXXP+Usng2YSmk2V
iuBB4gEGVpySJhwsgqw2hpsTHoCwL2wZCwzEKWQ9Fgdj6O9KIGcyjPyYUgzRBWwjqZBh80NsTHQ2
KQviRwm79jzRVqn3GtwdvgUCWj7uIIVcniNCFQXxiP7RZ8CVKNPCZ7hfnrI5+GCb+oY3vav9keJ7
9lsXDgixGr0y+ez8Xs0uWqV1zdFlGsC3nbCQIw2MEj9kW5STay4CIpBzTC96NWXHVmmikEWUTf9h
7jqFiouGutfFR4FMAvjRv5d4zkeCeIkHT0GufZTrFIBRrqWbInN0W1pOk5tNEUmYG4/3UwMrUNUR
rtcDqkdd2nKx5x5zZdImLY5LL+bpnlDQD3IvPzja8Jv49bVrjhgy8dORn/7QgXgmHsza1LHla+4B
4uZtFB9ku+Gy+nA64Iya8WtmSyTfjDe0F+BXMQGLm4U7rz2OBAtNXVgEDC7rXOZ/nHHDvyLtZ57G
FER/MingTsCW8hcDPWIJZbb9nksftgMXZjOyr+mdN7q8Ow8p8kqu/vBbnSiPpy6eLdLd/1fW3rwZ
rU8363ymYbrKHT/a5aJzcTp7ldGlkxDAGQKPw5i94DtyoFSWCnT1xbJm4FpsKJBMHbC23ayGpQM9
JEgMQMVhbAHayBgRuRAygBnAWiVchsmd3ovgrWbeR+TODG9yFuDsIUvne8YZVD0jimH0aGsbUUxY
VxYP5AGvPlF6mnF0RSYK51WmTI0eQGCIe6OZmYhU2GLPK7l7nDvBSOu6gvDV9EvMtftc+6qOKvNK
zxvs9hvIxxI78IdiT5TeZoM12iKnJtoln1ZVlYwYRR0jrZ8f3+un1H+6ZDPTQJBH7m8K8uGrGoSv
qOUEo/CDNpY8gvhIeSrKuVs3OTQOvwVVylycQa6tpnN1CdyImhpyXeaiVJLUsbb4chw6p6fI5n6J
vzNLHOUIN0SVwWOIbd5CDpnOIOR8QoaO+C4i7EB2A1H5cs9uQblj/ShizbhOhw2wCjbRXoboknBF
gTmjt2F8fYuP/i0187Zvki7pMxj0slNBTdcuqkaYnlFqb+Xol27oDnqRPbF9441cV4kczXYTi5wJ
JO/6WpOaQnGIe/A/0KKByxHjh0BIi+m+EDWQSR+w92SJKLdGa0o9t5vyF18fhwk4FQZJJ64J8qiI
/lbrWTXCegq1bBzK0pRPOInNuvYXLDciMkPJ+AREji8hmeZbnvCxE1BPCgb6H3hHYAPpSfe4x/wZ
13ATnYJmNadgN5XAOY4+JQRHzibep1yPly29Y2K672nEDMJsSHoAhlLZZjrW9rmLtJLov3lA8SOU
aPHnU+p93o6aC0y4n3QxvGrhB9O3Tsm0F5eXGqSI0zKOg0DuP1mFLMaO/bPgkqu0JIz3q9mBU3q/
zdJQ0yoTz7dtnhn989aJtPIP6PVN9foVqt1ITJE1iCLNYhV5yb0q6VuNS8YZH49jYR1DuVPjvvQi
4s221gCLUyk3fl2z2GGohyTpzSChSi/LwXQIuZ+Nhy5lfZYf48Nop5Mm4H6PIbwoUlHTryroVhUn
qez9qVJo6/cv7Uxy2cHFYzZ3QzQBFrGHFx/cObeO8ZULhpQjB66rdL5tDfZhG1mMsI+kush0CQCa
630CqPI//FBPEcIXopGJuDR4OZZvL52F75QzfCfcrUb9nVdzoGS8sY6gJUpqguheMbvCjxrMfUCw
Br5qxoFw8OI8xpTbAPrRUMPhPnQcLDGCSHDj24HKg2S0LGAJf3xXdD4k/786po2DhktJ2G/RKmK5
Jw2TYQbRr7J2RpG2at7VaPGRuDl24wTLYv8SyMgrUgfZH6kgXyPbeH2n33KD4v7jkWu473jKs61Z
S9iaju4uEuc1C2l7n7/Gu5Ve6cAjhSxySWsltCCg5tgc+h5QN6BF/GdhBa9nFQHYmcU3NDcNII5q
1B769axCTGLeLwxEznwp1KDjou5A0fCI+crtKiCgK9BsVlWFxqnrB6keaWCHzsC7QJ67bKvhTSqQ
DgPC6pWovsk8kumm9d12xMiwKwHhBBM988atgLvM+gXY9W+jYSaA0oCR60D/dRmcWZrBERhHt7Et
+8ddNdm/9hqZLrUP2LEhHBHZTBtT+wPhIeUK6VbLSKY7xNygeeEHnjFvtc0HjaVIuyHJDydsEb+1
3ZcguSk/T/MR1pSzItzIk993Kk3rnjI1/DvBXHfO4y9nx4TzNQKkwaxNwWb7V7Lk8tEhhyZgvpKw
1oS+trqacrO0KfgDdiHmyZQytiFRMBomLKP7wO2tdDTjYuZ2Bx6eICjnhxsy/LCC9HrEWEsVhGeQ
byEVIExCwJsIwFn5S14qi3bmVIulDk+m74RZU7C5NgeG5zqA4WZLkVLlfvPPQPt6ES1FCOYXJ48a
lZZYmqORLPeEl3hZG4QkfUVWcdR+baBerhmQ+jzIDVlKOvEa7qMJNT5tubxdNPPAmq0vDPKYHLSR
XfvcMRb4qo68GCUwUXvBtRmma6AkNlx233AM59SFimijWJeZ6f9aG4D1OJmM57xQ65AZXImIfrvI
VUEqU1TeWgmCB8lALAdQ4bFjRlNzVsNi4lGcgtTmUR9NJLVX8hx7Q8bsVfSQ58KIHlgR5coEDCIM
+K4cignV1FphRq1jubLwu6N9D+68TzLc2JiXsjDbecHzEHSChmRQXT6OH80YvBMfUkqzj8oHF6Iw
XC8VebT0bR4NKgatdONmoYYRdWebeqNjXhvnqhqmMZZ7gpUEbQweIwdT1R4gRq10RpGfV5MRYRE6
KGGvV1O/iU/HNHAMiVt4FC8+eJfcliAuigc2q8TUBt2iWMhqiIyxQdeBHN3EmkuXNu1xKAhFn/Zi
qPtU9a76I3G3KhOvcH/s1PNMY6zyyP1z1pncrer/sKWKJ8WpoZ+DyMA/991rYkntYMqkQ4a1ozCt
O+6aBCO+YgyeHmCG6NGjonLY0q9KupNDnDHBoHNbOqR3eEtOW6GeQQq6f7VK38BAa1iVbgs2Opcc
jhNzQMnqSfYTDQP+2h/0ZhaW949uGsyu23hGHigWVC+tQXDPSKSLaA4kX6ZMW0VuKyn+SPAR2Odi
YEyfYc2MnD+SDYHAyeHTWqvT2IqDJ1ClOzOhyY38MVyD4Elgf91TIJGiv8jdgO2BOIRzxFM4ks/m
lxKNE8jPHy4/afylMWZm9Sp/ny0fvptmj8w4iLtxtMDbY9LNtLi4x2IW/tu1v/Hi7Zsja9t8imJf
IPY9FZop0M2A/gwp+3DcK9NEJlljJIDGhX0tZRT2NF6SHo+Qq8yX5s5bWrb6ZrYwKli7CcJJyUr+
fnGfPJbFg6jT7ajKEqeOHaQeW0ThLXrL2jykH8NN1yk1Gy1gvYXWHDNgPxPcDJPm+ti4BweBZTG1
sdtOwney+O9WYHRK//pctdOqvyvNJabQPbmUz93mC6asdO1UPi9ClH6bErOp1898mpLyYj4NRc34
w4UdVwGxhs19EZuAfguuf4ZER9s9DFiCm9waCs1egvfBbdgefRaF2P9dqPJJm1Xq7ibejHulNyh2
ktgL6XtIRe1+s4Mlt/J3WdKHCIvBC6hPu3EB+dF907abrS/UcLQqqcbVISvi1kI1PRUPZlnJ6g3Y
NgFGCP6fiuYjTG1Olb5NyIW58SL2z9saOqYP1U/1XFQLOud5OhSLXYpQ84zVDmZi0x7tz4oRk0TO
dqDc3eSbggCLvw6ep9jp+Rp5re/FlPeysGDjR1MQUz+dC6KJeR6C2de303jd1LocJVpRaebnBUjS
pR7262rZobIfHQ1m8EyPc9wIZGSipB86UfToEH5WvIYo35+8qAOS7NJD0oNAvtpajukBzUUNKVVZ
kYZ15sIH96sg9N6vyO1pU3hwrSez/yjPIXmWRb0pvRMCbExGVy8ZF9ezKN8EYUdcZv5O/tQkvbRs
LIXApf/7724k1Zk71WabQtVCVa8JRNXk7WwFMubum8LlEYBsiwrjukYBMQI/5hIZRyIHmZPdvM3Y
LRAyX9qEHFQdnNDkSe2a+NBREDEJJSyCZlWy3aR+PpLeKdAdUoMVZyUBEe7FZmgdlXApeYFYlWIB
l3X4YzUz4Pt9QNt39anJ8AAWE7hH2y2HmrA4FUV1L1vb0BDGY2uyK6A90EOWYMTiEe2NgemUCtkc
7XIZkooVuuN+3UBn7K8ZXe9YIv4wkkyWPLB2yqQmRmF8FwnwVqkERpqvE7H/1YYFmVzIP33k0Vwl
cbR1i2QLyfwHcDEBg36aK2rBufH9uZ/rqAL7J8VfLsY2XQ1E25BP4+TgHRtZchrmB4ZWwzcxR5cf
T37V9+l1FbDHLntjMMB8/qcnyVxCKt+U+2JmmPhhsLgt4/N90IWLI+x42t9KxmiRRiJB/F6PeODv
lXjellwxxUsuFKAEp0bVXcCcaAQagaMADPleWaX2n/geOqek7rf0viwCNw0RwYuc6UlyGm8DVsCs
tC7jqISYHyGJL4+RfIHwhVc/kQ3PIwHBs5UoX8ZLgG1EalQiWsc0I5YwEMowyoH97lt8FXn9v2P6
HEOF3yvuqwjZ2qREMCIaK58gxKyPK7oUfc++AY4hKtDEqzHhF2VzGcnlYZrInYhEOBwgn7DyxtQq
m6SlBjDr55fFKv/YH4kr4Iwod470PQ6HzyAU/oDpZTJ3j7MhHLBZ9KubnpdwFS1otFL/cp537X1r
c0dm6k8fyLDCZgm8FMOnXoXB7txeIV4TqinLGnpgTF5GokZd5Xt4kJS4JWzNG/4XO30Nu3f//jyh
vIWggOZLftn4gSsHMjLPfndDXWAEdjVwtJzhYj6aWDTAbsyBAZRIpUisu1ZtG3m0jumt9OMa5t0r
YKp8tif/ryF1oQBiKR5bHCSRKGGnKQCl6WKx24EOSF7Nw3zPuNVik8MK9ZBl3X4CUPfJ7LZ4+sKz
FRAdvyxerVNzVYAXBSDUFbMYS5rGcl0Hzum7fwzv0c7CzEiiNt7BkAQhVJjHJmUDjgLfUBtJdXtV
nT4Qvt9g3mjALSxkExwulJ2l9wj68XeXzEcr7cU/ZWf8wEN1aHuzOflJYLHwV7vOssvRt+c5+mor
ecG37c70AdMUY1IbmkY+3B/qAw49UcIja/JcHETXFNxyH2WfrYmIIFt/s1v8b9cOHynLqqtDjwyW
osnjUXp5xGM24OXrLA83H2wlzCUm3Axq1TJJJV9HV3SOQW4KQoTToFOkiuf12bE6XTiWeSEr858J
Me6vdZ8iLVQO9G7qussHhaLiIIGPpAjB4iTbuXQnFcYWUHBoItX6p9AdgUQv6gU+/QPDrEQorHkU
dlqMUvs51QoCCsDAyqtJfcVUY0gsi42NBZYotqMKFU41ssjxl+Hl8SfNCau1HA+utdwJiOMPO+vz
L37IHfPLgW/9amDi+5z20pLvN2V8oa1+euK/rJr57YgoWcTBH7bR6ZfReBrVyzI3lLko+3es+w70
oDdi5BlP2RNKQOk2GcLvv8vSHYUo9rM3TKVvU/y37A8GGlAErMK4TaRiWEQP9YS/Qdp4bnvnXp0T
AaaXFTZefITGJBPJnKOYjdkpvmgv7FPcMys2eMfrcM167/ha2m9dtq09+lpohG0bXtKV/IVjZsf9
lXUb0bGWR6q8gxXivfjcdn7IehpSimVem49Xo46DxMemQ9yubJKM5dcfVaPy4PJPre+QzVXuPV3d
035qDFqXThCILRCKQaDQnFC9u6EKC3dD3ySel9naphxq5RhStBuv7fT8WtIhGRjMC3beb7hOCoJ1
fbCEWIX1tr1iemPnyVvyWjupHPJV1wAHnBS+8b3laTGurtTRsvHbFtVmDGRLMGGmLr4NsfOykXUa
dZATD4an3pFTiiq/J56yXBTM/X03gycryFahoL2gQGwedas2KHuk2z/GuDm9LGhjPm388AN4W9xw
58M11/j9s6WvKVn/N7EJ7pWlQRjIlHwbGQaR5RksCzFP0VpmEHe/x5FHURMnqbBDI8+gylKs35eG
GR2+9C96ymMGoNxxMM/0tugWSBGxYrQYFbL7Vvdx0fXkGjGJTmgNJYHCNptqVTiH/oIplMS7v8NI
S2IxdXyqG79ZpcY0Gf127D+G7htgA/oaxH1fB6YRSIPlkX75m2dTjf1rQVNWMekJev3+Z3Y/7e05
sDX9ieosTysFvqKWlpjuSrnmf+gK8boEaP2zFKvLutRSUcAJ2knKlQqhP3X7XO8onPMzHsUhqtvw
lhdnWJByZQ86BV4moQO/jf82YUpD+Lia5YgMl8k2j2YgURCeNNdlkp1lGKTHYSKWk5UilVglxfv8
O8Br1D6p/9lhkg3uUfedGSZUC0aCc+BHv0Mhy2ZwxnPhV1I1witfUDNv6wybj3AQtxK3dMS9oV2g
8ISEYruFITd3Yyog3XCi5pWKsyNlktPpYwn8sZMlkjHeiMPiFtpFcXQN3v6nfqIb+AEzLZWv9FqP
hjjWo1GL71/9RILJzk/N02rMRqKX3tBAJesxCfCGCW4jg7Rlo0ekmfxhf/J+WI4FTI9z3v1m0Qp0
FXkd2B+DAk6/tkREnoFLTs5bQFGArYsvoGsCE7C26+wS1IId996G93/NXfGLexnVYcbtDdYP5/ki
ntXDMGl6uZnCKzQ5F8t2lJqUFOsTTGKKcGkNdkYDZKvEkNcdu52VuiCwLY9DdxLnI9z3Ms2DZwg7
NlxKILNyiSYClb6LOQSt5D4eBhXFeXIh6YXQczL2c41rLng/IypnY2oMtxoTu8Se6SEBUrrmHS2x
UyhkO+shbwSvXAQyPfffEeWvq2ZyKedzTJWDsDxzoc4tBOuivJiqtaXZgg2MfueXXjdfCo1ajkxF
dUCQNmGL0prfllwNXw35vhmWh2ZEnuFtxUtBZE4noPIunfr/3l9wNTL24WRt0lecd07iBG2yjxG3
oHacF9/BCqLEoQiUWfnGlc0dyG47a9hs8I0qIIKRyY1HpAGEkneltij/vSI2mQFsvQFXaK8wHWVX
rOEyfJYk1d1YimYPdXk4LB4wthEup+/RsH+A6Lbo5u/NrpR+4VY/j7ha05lLBZku8dnmcKM+2dvj
rCXxv9w1fDXUfThe5/4k40XekLgK8kdrh2RmYQlMjDZV8h/aD8P4G+3zhkdMBk6d0HqUTQYHFkNa
mKNYetdITKG7emdZ530/6TGZBsYM8EprecYTdZzVgdMWDc0eXXFbJ3LKbqhCTuNikJPFH6VJlM5t
ROcbXT+Y5GCsbCQ3/kT2Yi3HiQPP5pgf1RlWbb/xS5g8O1S3CMrwLdEu+bAeLB4K5emuSNq8WCt/
CFOLuKwBzXre+UalS3nQ+pdHD5uNXPWswS+OoN/hLaCEBGpbWvCEAvflvpV6SRNLH6xpbL6Ss+eZ
hzkkb5QJcOl1GUCLqN4auiIooLKN0zrnGxRJJVGEeqHJ550s3z4QgQU5PGKdBsbn5XKanJ/L+ugB
3tG+UrLi1sLsNTNKgbzVN9wKsswRzLtkXYbUBUyq9d2s5JNYRm6eStRwxCByQy+80C0FKDdL7E6Y
FSURUQkMA4g9msLzb10j44VjNQzz/FznE1AvqSVNDi/XOurm9ngmO4D5p/ArCfQ2DRuFJXkgvhx4
3mBNiFiRKCmyOLPu8RW/xIkwiIGPhiYmJ28CBKhRWywMcJu0vP11p/7jkjaTcCQRH6x8XAmq9d2P
EzfkzkQWAmD+/b5dpYc0PRFPtEYBYsu1PrJgUPwK3wlUiFf9vy7MbIIHh5bcZbAObQI3MvWRvjzo
DFrtWJldVrWz5L8Qgxfhj127XVeMEEpDhbQfVRqVK3JV6ZPp8pT2XlxSCUXhHIPLE/vlOQUds/5i
E4bzkWBiyo3oypxDX54nNLkiomhJK+Kd7faII7GEl2g4a8B6fm3R4VzwHjvHwo8wMDK2wIY+9ip7
kXYeqzKvXYr5YtAndmxpYFsL9vzJRu2+5FG7DvKOE/pJ8dRBZsqEs19pC7f+ZIBAcvmQ/fiZPkfs
XvMPXDUc8mUr+ntAfjIPxHh5VSmfEZnbUmeLYtoBcAoFADpKeciccZiJ2zWgWSmwo5nJzBo1iIaf
6zxKMHWaqb7ImJYQewmW0Yb81gI4cs9pgApgObjsrWE5gmErrGB4D5DvT4QQTg6BdJYhh1xgtuMg
eJYOAKJOg/KKjYz9VsHrHYf3w375+pKiN7LjMbbNIW13H+6lvCJN7ZskYd1B2q34+Jm0W5VUt3Jf
TsGBUz+sYRhkYhcAJLaGDfEJoLNw6ZvhUu+lNRiH/C9yYT6vFsoVTkfXBVxWX5vofbDFOxcSsxNX
nBrt73KP4VuMhnYOSjiFoAXdNs8RXLNZKZO4U1vyeCT6zbhl0Q137H+8+XSroWPZXqZJuGFC5bps
2YGpxLfE0tktCMWi+iNelCntGxunlMA0SBweZBteYIWk3+S4cKqj9RR2Pbc9Yxiy0vy/E4bTwzuZ
KWMa6gMac/qyzPyLfJUn4o4BlviUwcO/HB4n8aiG4oaIzoFysdY2olrHw6I0UbRydKwvlNLpXw0E
oy4nMRYCOkLVAejLh607QC5lNmtG6zxh2L2NulnBZqFfFo8lyrBxSQQ+4aAyUo5cFl8A5N31WSV1
+Bf3yZrtm2Cw+p64EkaFnNKFIJHg3qr1jREp5lL1Br7NHmJLbJOz49y3QPw1wuzYCzqECCmBc280
I0Q31Ip1nCiOoWYV7NbcHgidC1zTuojU1mNvUFL5nECafLINqGHV+8cQYiwCNgouSUbNmqWN9QP9
syY0h0MWIP5U3bboUSWJOcfE8MVPDt6y0fHRhvN2CRXS2RhJicod4E0uUjMjFanRj6/wuVTpbe2Z
iTEiuiLNwhRu6DrjMNBqh+6Wdbq0k4zBdnX8UHcP4xfI2tssMyChGEEAOcXwMq/HwghdHV7S6D9R
cnlX8abq06UNihdbBl2UGNFmiHEWPUAYfnJfls/u+aTe9JMSDC6u/qm1/cCzBpi+hUuxYJ82KAOc
uBBuIkt4RluArLvgPxfaDNwLImuZo3xUE8UKcPGzBxl9eeppzemImDa98DzU6MHVlGOhg/Lc50OD
DzaogAo3REhfTku0eBWTzR6symufdufxHQkNuldv/5j7mFwo1Ezm+xL966egVkTf2Tjd+O6t4sNO
OFJY8a0cDPVn0pd3WEkICNe7PrZZulsADlKLw+Sl/o0575lXVXAOROs7oThILwENhIJTHMDJj+Cm
DsUCsXDR5LjspdRmlUd0YzOHRItwD48+lpmeiMBYvoJXn7xzKPYaWN4a6OghS4vLuzvbUj/wZQGb
9syI2wXq5e+8Oxo+Y5BjFhhdZgHmuF0P+xmXSVchh/iaa8j0IQFIgDEOJv+RlU+EfRQCEXQonQ2L
dOyc5KhvWNHWXzesbnMg0C2hyKxSfStSRfht4oKGoIGjXwrFWhpoWjjSuKyuOpTqXWAQmfvhhINf
eefRXXcRl2gB4HWQJ/QgPm4DBCfez0hGIhMKU8d7xpXo0PXmOdP2Sj3a3SLA5UlNVKghR+fetbJf
y41Lt8oF7e/hJSn7gXuUYZzesUc8QWx0QXhGSszxlGRoyUKSyx9BFj1zejxBM1qtpE/GS/47Q8MM
MbuU2vt2CF+2Jrh393eyBbrZNPjuHzcOnTBNAWo8prwGiZnO0KmsCklJ6nSiWCAs4Av+BpXLybOS
21/v3u4FLPiwdFJUC2+sNuY041FxguOOFK8BEn2iKyodU1+Ix6RYoHy6pUkxtzpWbGKogr5XeVpO
Ql2k3DbYbN27YWvw7iQigqelfP1z6jwsA/zlZB2+Yyddw3UhzwT6XH/ifjVzNRA8cRFkNrpakygM
IXlDgthjvmlzCUAMp46XQ2jq7PQlVu3CcOzSDfrzReQYMVzP5Ug+QYgoCcDAQn3luSfL2u5LzxO5
/I5i5ldD5UAZNivQWJb+IBIem8INS7UtBIlR2i6HlHO6fRdJJ2TVEp3i0SCvheLTxS75snyE3vlo
h6a+G5zcnb1rUIcGez6yLpAdLlhZQdKxowv5wjUcUo+hfnUiqOqdBrfFZnjzs2/2GwGKBW4We+GL
kea0wDVdCcWK8xRAPnK4BmFBeYcbVdtONiSja2PYez1N0YCU5wG6kP4JoCFkRUtIw3sY/igDEd4g
FHKyEdhrHqbVoqwpuSb4yqiWkkZo8DnlLDG0HaF3/WngA98sgmFcggNAIMskzPQ3odA3LD+lboG0
ZLSB84wxafwcZE/dVC7X89Uc6iMgd4vyI2sE1HgOzfc+oTFYgDrfWR786eVU7Gy0BYgUKEPdJB2l
hbOV76gKVEhVMOi8BTp444VTqPjZHMiBajhC4NIrrqC3R+Y+P5jIBdeLvkmU9zMNxkD6UbN11cWm
KG1aDkmwpfzoDd1FJo3Dij6XcuWSESTTEM7kYm3KsBeWYv6YxxEjr3j1MFoOmQOCKqy64o13fQAx
5Qc7lQfq8GIrJhCTHK/4ePHGThrJtMbazg88AuoGSla4u2aCYrWcOp/uIUjTL2928giz+ub0KMHX
Yj4PZ8MbI82Hcyrvjl6LIo4OyGHH+bEm5Lm5+HhlcfaEw26zcx87BrdKyycbMzfi+sQbd5pgDxVJ
GnOSiyw+gI+MyQ7yL1MsegRmtEesBVvvOHQmkcBhpEdYc1I4CnFzQ3vMXiGeR9vLNpWNZ5S4QM0X
dXPXgBviX6BDqv5QGlxYp7uHN1UsLuWPF4HFEr1Ag+rlFvGtD5G3nJ6r6YzpFHJGDivYB2B7Um4G
98Sqn/qsvVsU0nivKeYbcQqajUgik05gcWXVmbHHTfK/KaNvZouaWpsgSDWt2S430eXMqv+RsezX
ssZCvR6o4xlKj41jvD7oDB1h5XyJXSjwvgYqRLMb2r/7HUJEwXojTf2QRS6o9SBUnpbldh6hNkre
gYQH+9jzez42U2Qtj7eTqED5qnLKWHmpkESN2NCg4EoDmmMZPfbsOTCxT2wxeoEwB8NQvln2iRDA
sIychj6hDLUC1zqBUY7ye47IzrIM1hOmVzD9SIUbttOTCNS7Y/KfhtBTy/2uL4QCwqOo77bFIaoj
ec4ntzmPwJ25dgRoj5UPeli8qeC3wkjYHK2dMva4VvHnkp5csVPrjd92AFWpAeKIyRgDBkQw6YbU
GRvhi1f/P6rMYhXYHR7yCfwd5t78DVXz2fdCR5T0he8hp7TxTCoOyDYjehmThss5SV1dyxv0YKqW
jVjhIkNKjh5U0ju0kqxkCQKAuZQMVRmYBX8R7bjnrJFLRceyF256dFPKK+fiAIVpbpPCxMhKgiMd
cuvtjNttjGkBKC4VvszhfQDHRO86WncmADZ5NylRoYbDj0mFr2aZ8ABfbIPImqNFcrwDdCGGtx4p
JYgmp3/GO7621oZKF2CyVJbsjqIVnqtzbdzJmSpTLZnfyAnIfiZ6c2VmckymvbN6fQq1ragdW15x
OCspnUHDeMPj4uOwDYbdfwA2YCbeKsL7z8MTbYov9rlN1iwSqsTuLVIzHRbKP7JwbQ+vFHAgmVOi
KMaKHhfdvwz3ZQeYL0vpUNqTDC1P5ITFEsGQZvhCNwZtCjaQ8U450ND3KHIU9I3RUbrgBVQSUa54
HVgH/co6YQCBMPJqzrKMQGt7j+6l7R4cT/xL3WQtx0XF2NJ7xtEyyKXDa8wpCn/tOpR7YNmkW34S
5IB/9n3tqNDbira7HGTqgWRk0ekxZB72kMQWB1FHsnjhY+vAeyNoQogBBpFjFMEA+sZrVZX8IYKI
o1LXYiQ1YofEQPQVxcloKXoOqeOlfjHDf0wn1gUTtM2fu7z3TcnU3lEcB63mMl9jtkhn1sJ8oix1
bzPWOFmuNP72D8wd7EtnX1e/BPzns0/7ZlQkR176+i1+RfmPp35+xggBTU2umGogVahZd5rlnrWp
4UxC555bYG93cJti
`protect end_protected
