XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�9�=�t�]���T���G,@�M���R�hAd1�`�GZ�<	Ǫ�ƪ,N���7��v�2������}���lSI�N��w��nBYi� ��r��@χ\a����%�:K3/O�]\�|�ݪ�����F_�2ͧ���e�@��X���2AQ�ϒp9�]�#]��7��oV����Y���G�bA�1t�N��Ia[�\��
j
��w����8��t]�m��v{㷆{2����ף�L+L��@�fL�tX �$M.�`���5�k��(��`���F~ﶃ�լ ��M�v���Z��l�7��`[�e�b����a���$�LjQva�/��5�xA�mb]E(�4�����nۜH>�Z�1Nj���U9��}�����q�� e��/�to�a��[*�����?�8jCr��aԥQ��<�|�`&�V�'��p��R�Y�����Ǫ���q�&Y��;�˙q
WQ�� '�[&b�(�f���1���*s�A�ӻU֒Ж?$�{��x�s��÷��������1�V��S�ʙ�k����7%đ���&��Q	nP+���2*G��	�����me�m-+��מ�MI�\�<䧡�#��
�~� 9��}���t)/��ԥA#���*�Q��)��R�0Rf*<�wbOխ�[^��ݜ���쒡Ց)XЄ>������2-L<�+���`�>{%�9kbX�O�p5��?��7����(t����"��l:9���&�����(���U����R����XlxVHYEB     400     1e0�\���SU��g�K�֭�d�G��/N���\��˾8]��l�PTV��5,>��if�"��!��챩�}����+�ǲ]V��2�n�I6˽�T@����
s(QG�4�󀑪s,oŗ V���<� ��K�~�ىr�%�|H$���%)�YP�zL�֥�Xf�~a�vA2>�9嬩!�p�5���69�h�>������ѫ���DEQ�!wtO���\B�!m�Z����8ԇO@R@�O�r��\Ex4�wД�DDz�2�=�a��G���3�ӍԪ�{<Ҩz㗿��Vf`��Fb���hd�,��O��߫��8�J�rF]ԛ3��[�NpﱃEO{t-i��Q����6v/�ґ���M�>��:Hx/o'�[�r-����9Zc��\U�Ȑ�~�~�3�(m�����gXw5���	�%�������{����n>��މ�9�=�O�pmɌ��-�J��ׅ�!���i��ɱ�XlxVHYEB     213      b0N�� ��	~31��P�cc���i�6[�J�����FRǛ,*>��U�N\8G����go�3��7�x��� +A�����̝^ �c>Y5!\s�p���D@>χ}r�h�h�Q\j�gk�j�t�p��.4`�p�8Y٥1`�����hj�S�_ϸ;���G�N�