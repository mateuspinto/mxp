XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g���'s	~��A$Qh���ep���왭,gC�X�ɀ>�*�Z�~�cwԙ�y����O	�˲Ŧ�#�D�e���I�U[ ���=���5Ӎ[�!���ۧ1?�-���Ż֞PՁr������N[��/&�j�)_��H���2˰���3]��o�G*�"��)�+J��ZX,�<�KZ�,M �2��6������M/~X�f�� ����?=�]��M&���������'��$P�F�H�	7�7n`7�[���&�ǇD�� �'���`OM�z2�IF�V�6��4h*����v�b��^:��(ݜ
eP��R)-F`̨��Yx��Z�*r ϸ�)��R����C�Fጕ�(�=������i�t����/�yyc<�~����Z��:h�����'�;��� �,��Π����ہ�e7=4_����,�*�3}6���u����v�̕j��h�ܑ�G�l��d �^j��:c�� �cc�o4,�PWwRTF_>F{���	���Ō�`y~�@��=��"�GȾ4O���˂�<�E7/|[�)G������(�ı���O��u�^����+�����Fl�'�+gqL^��*��c�~ �xB���G.��\�{W7��8�L�ڱN�2���Gԅ]ynx����|m{C-�[����ݷ٧��i���a�8����ط.[����K���G�E��QQ�L:�e�Ѕ��]�4��jڕB�q���:0��s�!��^��@-���ZͥK���=�U�'���XlxVHYEB     400     1b0�6v���b'i���VE ��Y
��W���wv�6�L)���4��&&��!c�[�F��!>�s��S ^�h����Yte9�#�� �z��H#����E�TE@z���.zS��oP"^�(,�����8l ����-�d���<����%��eJrP�wF>�b�v/M�3P3
����ͼwЇ�b�_N[W|m�f�#��`�z�o�u*���Q�`/������X�B�_Ĉ����o���h��i�p4i{)�6�s���ߐF��UC��ī	���m�a� k��C�۫�J��2��//C�N�lԶFm�$)��%���
*���r�-/��_�g�)�;��q���E.!ύ��1�5}�Hz����H�;�-��Ӯ�D�ΞU�o^UR��m���;י�m��w����H�j�XlxVHYEB     400     160](�
Z���ə�H�e��jJn�E5�+y6薡�J	ڲ�[1�x3��徲�5�ʴ)��qz{����J�ש���g�;R̦�tሻ&b��bb��Җ�([R]C7�Om�B���tg:�^o��Jbu><��tu�D������8�-�
�����;��}��]�N4�����{!t�"�ي�F���5&��"���9,��~���|!�T��\&��ݪ�/�*\m��x&���V�H��nC����ڈ,T.&j׍5�a���.�=�"���Ջ�K��~�	��->��Ǧ��=��v��"��?{�i�j^6���*p��۹U�����`P�ꫜ�@���},1XlxVHYEB     400     110�V�K�
�t�������s�<Y����e���ƻ;��~Bz8�A�8�S �N�'^��]�I"WV�h����TO�.���w]l�ε�\P���Js�g��|�6���֏lI�Z��*W��Tc���#�(��&J��\[ubO��#��=@x	��l�S�-��(~棄�߱��-�hA=�:��.�@?�a�;��p�E�$�~��a��_�v��LW��?���[�c�ý50L �t� ���?�w��动@Y��9�o�#�q��b`�2�XlxVHYEB      42      50S�g�j�ug�&_	?�9�,���k� s]gI�1�D��k��O���n�wL�Ҟ���7���8��7��� �|�KB�