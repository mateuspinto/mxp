XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����H�����Օ�Ź-��,q�E�D�@<�N�ۄz·TE�_
;�߬�����Y0`��LՌ�c��tb<[��$y���1y�2��_c�68�J��&NΫ�$��K˘�Z��{����2� 8��v�-���*n�i��`�z�@�8��?g��Hk�����+>}��&���F��Q����J%��}x7^�)���\��J��]�@�u��P��i��F:���*H�����4ʹ4bN�nJvB��]<��f����y�]��(��Б'v�$�Hv��2�D�#	h�몂���P�:;�ms�e�G�%��Bk���R�����lb�|C��e`��^d�/^UeS������K��A��R 9�22PVJd���8^���5[*�c���L`�܀T�P�����a�:c�ל�ڈ\vU��e�Gv.3aCAUĹ�z�/~ ��w��G\-��H��ÿ,A���D��}v�T��R���;l��O�2gbx<�uQ�������e�2㍡~Vl!ʃ���C�XȆ���|���W����t��+&�b�]n4v��ve^_u�W�-���e�|�C��{�3 `JGyP_�Դ��j��8���Mw�lc�/�u���>�oO�����4GAx�ѫ u�"������,511�(h�ƘIY y{~?�-���z|�[�����s��W������u���zi�U�C/��%��Wۏե����y��O��FWwC�n[V���`d��L��]K#�F숤��3���ʽf��K�XlxVHYEB     389     180�Mцj9w">V1��Ki�AM�lL�9���gZ���eBh7�k�z�����'���5r���:N�^�)?e1�/J���Z{��]���vT>�!����aAz� �A
�G�g����"6]� x��Dp3Q�y�	��s���4\�]�+w?�������M�ZdYdr�H��1�F�1��2��Q�*�S��_��
�3���~�����_�аX菖-V�9��3;שB}�\9;��z�$K�q�ݒ�7�����aC�S����#OzLo���p��0Y_�>��1��k�~^���_jƽ��&�Y��1F�po'��3G���dy��(��{䗿�@����g�>xg�k�+�1�>y*�2�$6����I��c�oo�