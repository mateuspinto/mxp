`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
faokpuRlrtMfmOoETVnbvvI8ee6RARnWb9xYQQP56GHeezmuVdh9e06VPJn1sy6NhV5DKdjJCk8S
SSA4bZqQ4XF7lssXSX/AIEzxLjxOrW7GbGKX6MWk76TyYRvFpmqn0tct2TnYJF+g/kRDL+Dpo8bb
oKcnM9Oxqkv2vq0zIK2UF9vM8qtTPtTJVQq11J1yyXv+IUhvB2fiZ+cZUf7NiFhyvxH3R/AzxJGb
Zja9OC5zhAeY7aYrqogyft1lNdm5jS8CnZLt8Hy7S9W+LRDLRD5liYD+NIEQAmORGzhhR4r/Ci1O
a1x5ewIJK3BkBx6Il49ljgvEFnFI9kakhqTzYA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="mpFJq+FrFtrKFNQcYELUttKMnTZcD3UbvURYe1HN6R4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
nAzNh0UlVd19Hg/Dq3SnIZrGwNpcrFg+EFVs0dQ7+jzsKZdQ7xJ+JXWk9+cjc+AWjeJKaBHueSaZ
RrQOGrEKuLFsEyJAuDKG8IyITg+xBZN0aJIa7cpSzLMNdw2nGWXOAYibUAJvWK0ACm8MpUGEn4a8
K2ajifnkWmejoOFgDsiBFoMhC5+8sWf3ISF54/NpmDOo4nbOkgX9zPCpkooWpZmRoE0YAOkdydn6
leF1D5H//NPzsX6nxFtoYxbl50k/JGeexL+YSPRWJrcPk/eEIMbGhh4TWS0iNt9/MOJtj2w0dKck
kNveqlTqagnqU30DqGLsqPIpbIq1USGLhPwuSdLB2f8n/kXD4KV5AE2tEEUzA36StNOo+OwxVTNB
kj6YpAChV+7WsW666/0xE1IFAcqGQoJ9fghHuVoTHYzImSWhrHgnqKxSFOEImU4SMbcrLIzSi24r
yKzrnNu8V34NF4ouPcnFkLLiMWx6yX20s0sXq61c/D4/hjlzzOIhL2TJhoUlnhajiSBxG0UigZaO
dDFY0pe1ID/QspFR0blngDRaL6OjUo4qC7lbbfJJOa0Jql+E2Da54IFqKV4fHCmcyMliAd0EdtvJ
3T5L4bzxDOddwnFuPwbjkwLjnMlDvy9lYd379pGGGWrQn4spo4/sgCsIJUK/496B0LKSndlbiE8b
pt0UqUcfXFayl1f8BSRydglhsp0M842SoGTQEuOCmVzT30bqWOENKA34yslHIo+2KjWRTWY88cRZ
NAxIrnKg5vnnX19v3wrkfx8b2LCZvZPs0yTo6MbHuxznwwRwMmNjolhRaSzzgKne1eGWqECnvn9Y
FzoRH7Wl0CuvmibCoj9Q08QO5Hxlj1O920PUuY5YnxUU+KpB5Qo+JQOw1BOo2RhcHHFeGHbpPAKc
zwEqz4z/py934WAh+bkY+1KCBdSa3fO7q5Al6WnBHNb79EbAlWsIcoBQJDnNQjyTyros3ZHT2TqH
9e5FFfHYqZ4fn4LBOn1kvUokR0bLBkfiiYZqQ8x8bTw5Rq83JxzrNDCnoBKRJsRuv7WJxD16p2xn
GE6YBgz3gOJpHu9hSE5KTFGjc/EPY5Q7FAoEsV63rfYjAj52SeAnsGQSCdNaUgZV/n+TVQlQBSws
gIGQbT97WXZvBUseA+8Ktls98vyTCKkumfJ0wXNb4MLcwleZy/OaqHa/67pzqnLU2GDPOujb0lUH
+YJ19shtaWA6ZV1akVWW1X5UfyAKRUYMSjiixZ00GFgp6wtfaiDVH/OXXOmw+6PtdQXbJiy8usy8
Lo046z7uFPOIZ4NRPsgSmtMlLd39vdnTeKIeKlrJQh+vwkCS+R0IO4VzNV3UepS4/LaJGOLM+9ju
dMe3IfjQdaX8kkTX6Yh9jd/BZrkzsHYltBjPtR48rQZZPpwtKCtKwi1zw7nFrwSBDo9JLcNHF2uY
7SecDekDYN2lQmiLaPY2SJyuf9FoK/WSpST+7Kc3KvMI3JxwkvwSR1+axc4DtrjqoaAJCUNGBA6m
F6nPt5UATS3kXENxPO9DjnWvjdkfKEvtjmw3Q6O+RSNaV07U47WCHoFnZS5H1KrBa3ddp3EeKnlL
lyuq3dposHPiK61lUQQiKt3wvEq0O2uROCnds1ZTxWQxOtalZJMC4jvtwhqDFriPfGB6BnmvbV2f
4K9/S2cQaaSHD4MusqWojE74iqKW85xXlh+UPV3X4bm9C57MbF5QIgfCNUXhp81RNd8pY2qSQTUy
dS8LdBhGu93baWT9Tweg9XKnnJDeprNpXmH70waHtFzf0gu/4OSxV/Ju0Zw7VUiyTlQw42sCjI9n
gsCmLUUuuP7WQp6mTvO8+BChV6Fjqn9D7XMsFkgiiu6cXK52ca9V64btexMRwL46oRTQW/Kmv0/+
N8JEDgy3YND8Q9MLv2j7C7DZC+sfrSgyN40FP8fDbLdWf5+bPuZwJ4NiLIkOxHiR/1dhO0Zw1/lC
dEVqZ43HmAF/OCbLFgn7eIOUDt3FwYwCq1+Sn8xnP2RpDGeOo4w1aSVY3DRPsDZ5NVNJ9jHzT8Mj
3MH7x3kfA2ZXZ6shwTxjD7XnbVc+neggbAfxE3zpE/FzYnKSaSr99+qQf4q5eioXjLjEEF6aPhyU
gg68aSD0MhrCCUgwIb1nmlOJ7Jh6RQTV884TG6v32ZH4rm7XtAGViT4bpyuy92hcWP5RJrYJhi7m
7rrJovZszdSbxTcV65lkvCtVFGxfedB/6Km2/wB3joXWBS+LGYUZi/HUuhQCep5S+qNW1qCSyfam
FM5L6EUGifFDfBd75c7KxkSkVeETPdb2Hk+9OsJv0o96Xtfmtcin+vQelI0cOaEsZbCfn6PqXNp0
k26xW4dq+5tf1OeOmmPJh9bCZIHC+DdTCxidteWId8UeTF5QVBQeJsOj1CtwcWRi7vwmmKFOqO6C
Sr2UCbmtyMQLle4Xsf4FPJIjMiNBEEyqpoL3erzs8WSXt6n8dfgNTLzi93ldldL03XLOVW7YlikG
vTVg1gRWa0+02hXPA7IvZqiNmSUjoWii7ehh1zHPmf6o553hWoDK/a2dJ9mTHzGHnhlr2dIfbH8A
Jp6evOpcRYLy3FSZrhhHoeJBl0PZ3//UI3f5GR4D6+apakznzpM9ceYBsSTOR+0cHZ9Kr/8KXSEx
cAUWO+YYHZsAte074/0i2+80kwzSEAD3no8nFxSzMZrHrfHMie4P5dUce1PZn7vwWmTKd3oeMZqn
Fuyyug/BDSYaFG2yLodtjB/vASxLG2dWv1XhoToWyWHxzFjbvAKHpoRPzGjwQh64a1FRV7Oet5be
ypGc8KyLxTPiPeDWupd4J/ZVZuYEQIzM80QwCdqWvv+jisBGLI6Uwl4bwQq4sIBDCtnE
`protect end_protected
