��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���UIn� ��V.��T�B0\�|��K��Sv:���g	�y}-���9�����'��qp˹�*h�a �C�(��p.j-��P<
��e�ن���݁����,�>*���D��NQ?<��y7�RD6dk�I�
��N���lz�n����-��gi%]y'!{�i��:uݧ�|*�q����k�9�h��'S�U ���b¯��QT��<��D���	�c�6��@��:b.GƧ�ja`����u�W�)Jt4t�Ey_n~KnA�.�q2��s�G�A6�ec�-�7<�YQs�Y�Qȕ���'��, �ik����,D.Lo�5c#��7�du���"�ݺ���kj�V�������$��_�TZI�LC_�"�: �6��W��*���(�i4�vD��=�,�+� �}����}4�k�I���"����e2o��d1�a��Z�bV��2��l��n��ː0@V�[D���S�'0Yi��_�֍c����O�bݳz,c�J?ާC��g8f$M 8xf袧� �.��x���}�)v����0��K���ߝ���h��
����׀�sznG_g���&��	$x��� �2���@����5�L���br�ʴ�f�O�/ډ���ř�>ù&�"�Ͱ�Rh���fL���� ���;E��EQ�?��z�W�s^Z���,8Z�n&p�F��c�Z�m�`�� �DĿSBzE2S�o"�R�x�^�'��}4;`��K�C�R��d���<C�%H0r�4v������u���:̴+�����n[⢽�M.E�]y!��Z/iJN�c�o��=x�ޟoaU0�bB�����W�����rj�=w��<����$�һ����0��*!�d�*��C�'�I���\��6����5��fK����%ķ��5�y�ey�Q��yG�e.�o%a�ϱ?3�n\m�0%.6�v�*��Uh[F��%���N9S�:'����!Ua��b��+¿V�4g��:Zm�+ Re��br=J5���w���$����>"��vs�ot��R��)?Q��L���$����p���ܟ{)�L܆"p�������3(��}v� ���Y.�+�O��C����]{6�����5�k~
��EX�(�\��((V�	����x��e��������N������������%P4j\a�F[Y�p镵�_���KT�^AM�.	I�,Q[Lh��	@��7k��V6Z ��x��T��)w��Y*�F��g����5�K��s�����O_m+���(-����X�8ϗ$��AT���-/^߂�&�ȃ���h=7�;��e^�گIa�uh%�;��+�E�"c�
 QB�.o4���7ח!$`σ+���]@�	dS~�8
��I����X�F+�{^��yC?�K����`�~��������9�9�`D������4؏L3T)�`N�6�K���8���a[���d���r_�%o@��7��x[�sb7����y�C����\ߖ���/�`uxȟO Z��n��zZ�-�ٶ��|�j��^���
�j�����;��ǋH�{ʩtu�����'
����u��"ө��c�A��:VQ� 3S��&�W!х�sŸ���������ιC3&�����M���˙�fr�*A��K�V�%�{���_�'2f�W>XFBO��쒾��C��ş�/���9�J�O��S���Iv*�Ч��ցQl�'�Eg���k���F
�󍐄�k��5��bH���<��Ef\ߔ
��ėAd�u���%�yV�����+1��22\�D&��)B�2b��?�����&�@@w��W��a���h# �OX�uM�nP��L��4�B�����e�X?
�X"����`m��l09D�q���3�X���bmүT�������f3h��,���kd�GA��C��]�7MG��b�Z�n2v��4�')�dc�ԓ�q]cp堦�CeJX����`����UP[E�S����0-�o<y�V@�:��������X���$�=�6܃aP����L���?���]���)FՒJ~*9��ّ�߭�C�i�DRf��D?1�v��KG�4�ȋ�/Ʃ�~[G�2�5��8�i��M�#������+��|d�$����w�s9Q���epO 禄�B��5X�Z������\hg�;�/�WB��	&�)�`Ȟ�J>�%ù��Db�ŏ�e#��Q���Q�`��I�Uq��jf���IN����p�D�)�=R�j'}w�ev�v���N��V�XP<�ve&̕�.8��<�vp��E~3?���I�����r�,���e����Ku��[���� k�<����/G�	��A~xn��ۡ������}1�5u������T�䂁!�Y��6�������m�;QҚ  ����}��R�6nYV1����%P�6�On�6,&a	'yK��<�+�_7l��Z~�?A}��������H�B �Ȋ�<)l�TYFL��e���K_5 �[�P�c�.��cti|������yα�\4�w���5b�AU��̙�s���q؀՛nc���i^����F������7����AŨa�'aG*je��~��5�m�8�c�Ƶ�z�1�˯09�Yy��wz�(?�����b�xPg�F��U�p:$2ӥ(�H�Ďb�!���,�yj�K9�j���*99l\ �*��Q�R{�ms�6 Jҷ-�+�7I�\��T�5O�?b���+M�� e�����ص����&L'�ԓ|C�<*Z�.8���>�Ė3x�F���5(U����� zS2��~��b�_c@���H�?�QB��~x���{)�q&>β"'����
Օ���%eڸ������E�)RN��ét���k�I�O�*�@U�o�E>���0H�+*�ei�֍i^�Ts�L��z�_���;�z�'JA������]�t��ìU�ع���_����#R S�o��|��	^܏�-^ �Uhlv�H枊ŠS8�	I@��.�[����i�8ȥ�q%M�9\,���$$���w��
qc��Y'^�a�VS����ZY|���C�	��#��9F݈'�~�[v�?"�2J�������xˬ�C��Wҳv�uK�K&�Lr?�Շ6�l����2�*�-O,oSWv�"H�roӚ��������!i��1�걻��r��H*�E��"�D��{@j�Ys̲Ozܮ�xһ^�!hQ@���b�4��A>��	��Q����S�ν�?������Oȧ�-�es(N�}*��n�P� �����>��P�r�/�N���+-䉝0n�^Ч5���5:TPC@�w!��β��z^�ɗ�y�z���m���y̗l���+j�w`bp���C�ʑ��s��}
���F�iĝlcm�GP�-qSm|��U�^������?.N,A�i,ū���-*o�SK4+|�L��1=�<�pӡ��E��aj/3�I�#yd
+��BS����� G�������RȻ���ș���*����ɨI��I���	�>���˷7�7G��ZL�rby��������L�=���E!��Y��:�-{��0��x��m�v�&�&�5���W@q���O����?�~� (s�h��>f�0z���ө��עQ�5,�G�>m0��M �^�$�oNBλv�i�
��0��䯚~`�Q����q�炔�^krɧF�*tG$W��ٓ�wͰ兕����c�7^�.s��"�SX�z�@-�%gidX>���o{�{����pҽ���[�c��'6I��;&�M�"�kF�s}����fi������2U,�s)��t.� 
95?�g@S�T���NY~J�M�x���-6o�yZ�޷�
����*���h�8U*3�0�L?����E�`}!R�-C�/!-dwe0���g�T�FѢ������ֹ���mC�am|GK� �����v�'���P�ƣ�_��Q���<p�T5�J�4�T~�?��v �CD����І���M��`�i�;!Vd�`h5);��ʏi��-g։ƨ!e�;�@��=+q���`�W�/z��D�<<�cS��ՠ�滼R����y��L�R�^Ȭ#�Ş�U�(�r:�����9Ddf&u\�.Q񂚝�x���ڮV!�٫���p+���np
;t�k��&Ou.��M��:m��>�"�p�p�V�e�4:9%_ܼ�g�8%�)���A�{A���]̪�,��׮'��2ߚ�v�Aͧ�*��Gn�j+a�o��MZ�קL�զ͙2�r�אo���R3|����w����`d3Xox{g?�n�H.������$l����k��C�?r��#��!51��z��d��R�P�#M+��(!��i_>�a������Y�9���m|�Қ�1F��`�E�qVB��Q��H_13�G����q�e% my�a>�X�3���W쪳��mX�~�r)�;$�qU���cd߸�������'�nڬ�KȂ��T�)�u��߈2{��y���͠Χ�*�V�#��QMT���cI�e���Lѡ1��vB�JQM�kJ��4d��ݒ^_-�p��RDM#z�
���/�XUS�Kb�Ƅ����=ۗ�5�����fD���C��߿��'H�Z�0�@,c�+5��o�_ñ�G˩$(��@�Hp�V��~/b7���=�Q��BX�_
V�Q5f�v2n���^�vEY�d�h,N�4-r$<��p��Xz�a�6������?fEJ$'ܰ%�MQ����4O~�%�GW���e; �)_��w���|�O<�a�/���#�v�\��P��a��������r���{��B�kS�"��"�R��Dw��6�H`�?Xz!��Q�F���>�(r1m�ͷՃ�t����2Zp]�ROwO�"?|!���XK�� ���X��9�S�ޛ��3�H^�Q���N�p��M��	K�>�<�6?��
	����L|zk\�I�+�����۰)X&2�����u�KŚ���^��!���eD�S��o#v߭�E�j�&*C�y��s4���4|�g��i�V�G�UW�:�ޣ��~`���~R�q�t�4��9M5.Q��pLT�!Z��4�8$�)I:רŉ�>��&��\$��T݀�y�^(�Fxۤy�y�:�f�~��u�2#6GN�D ���I�"��_.���)�@.��F@y�\H� �g+d�����_�0r�r�GzXc�q)�+�Ɯ ���,7�	��Ip��e�������jc������S[�����hZ��נ] 4稹q@0�����O���oٖf�S~�T�*��D�ސ�"(&���V�7�s�%s����eL�!���(a�r��\�Y"�}�f�0�r�X�W���@6����J��S5���Śl������R\SQ��fG�]
�q���GG���_�Z�� ��T;B�N�R�ٛzG,i�_����=�.v��3+����Pݵ ESx��$>�ͦ}֮*��H�^!'��πK~�)	�:` S�"ֻ�F�K�d-�)mo��I�b~� ]r�1*�#�=i��*$���@�0� )�	@jR��z���n��0��ƙ�e���H��/�<ia����;y#��熔
��Q������T�)��~C`�+6� ��� �UL/�>͆ca�Z��~�ŧ=���I6���]���m#��?���s��۴��T��:q�'9wA=�}�'$�l+.Tm�X��N-���ٙ�]�Ns��[c��5�#{Q�6=��2�x�h>�/rd�\kB]<��
ތ�mU�S�#Q�^>7������/�!h��P���ze'B@�0<���u�36�. ���� ��s���*Zf��D@�����&+ exxD����~R��~������F���kl���ɿ�`��i#�]=߻d���f`���7����8�^�=,.�'��l��������J7���T��`���0�7f\�,c`4D��#�4���#�AG�aЃПБI��2&^��
+S&�*���}eP���'���B]1%I�;�w���8�=�>韼0w�I(nv�뾦�0�B��6�C��AFy��~׉0n#�����������J�|�"Õ��N�bLu���ݟl̀5����8ԍmw�ѣN>���g��X`R��Û�'��=)�ڀ�T3{�)���dǹ��V��?��s�5��A���]Ľ��g���S�J�Cu����u։�f��Ȅ��ƭ�p���\�o����)�0.G�`i�Ks����-�;T9{�WU��>Yz�1[-#p8��i�#��TS��;�����;��fڟ�)�v�Ⱥ��9��1�ͽ4��{ .�r	D�=#{fӢ9$�-�Ǳ%T�Qq�҈�F�r��� �"+�=v�ܤ/��d\���X��u�%�x:�Q#6�[,`�fA�Z��$6v
9*u���_^$$�Q4t�ۏ���ޗt=Q�S �1A�(�����p���z,��qO��2���������%@�N��t:rS�q�YmՂJ�I��7����0���޺Q�J�o��	9H���2`�c�ʹY��r�b�a��S��b0�=;mAwx�o�;�LDL�#'qGvjeiP����]jAU�����$�O��V1���rcC���S�Z<���<e-�[k^�� ��QP�I�����Jk�Țj��ç�9��n�P�
">P���gv"43z)�[=��d��-�)���p&��
�Pϒ��,�
�P�B���_��Ci��c��_o����l|���M!��j�>'��.���>�fTM�����q����P0	�Ѣ��&gs�z��.���8B�Y��	�2���gAD���f���y����;m����T-E�~z� �7)�k$J������?Y�hCl:����U4�}S�ѷ ��\*'��~�"Ui m�� ��.PP�r�X�#��~���Fؓ��(���~T���@���� ��hB�r��Y��{�,_h�CB�q���妭7.=�/�`e��1�-Ж+[��cl�{��^��o�����٢Hɴ>�ub��Yw��Ug��x}��Ң��@*�3k��A�U���.G� ��JN3*WoLs�w��.�x�ㄙl�a&��՗�|�ȥv��#!c+x�s�:��))z���	 \�"vr34?��<��4h���pl�h�ʧ�
���G�q$��_�M?Vrc���dx�ɸL�&�f�`�2�q����-J��2,N�R�*��@#�VsjeA��K C���ڕ8G��O���]9r�.�$>|B��Ycv�֚��S���0����+N��;v���-*��"��	��!B�������&~��1��a����{��X��%�������Ǐ=�]�i�?�$z8Vb !�U�A���k]/������r��=�b����C��~\)ou"��||��DؔK���J�U�K*PD)T���?P(/nmem�x�0�䠚�h^�,;I��?T�M*�����2�V+D9�겿Y)��5^�0��,��ƫ%�.��ޒ��̽*���$ՖU:�s��ft#�FF�=���̎�R�L���K��h[y��[����4���[���j^M�J�4�� CV	���&�"�MO�n9v�6����o`����/kB_ЂS��-�8�w+�q���D�g�b��ʱ���dV#�B��T̒��5�&���s�h�)��R��� e�y�"���mw��+����=Q��!w������uW)~��K�~�S���H1 '�kk"����]���I��#����@����"�A�ShG��!����=���9��?Q#�����A�Lx3k�]���*��h'x�jv-��=��/Ƨok�����!�09�	��.K�_�,�ٳ�?���V�ߜ6=�3D�`K��5�~�n|�g�c�����Krڧs�v�U��/eh�ir�ٮ����Ho��p�+��2�X?��G�J�X|gZ ^n��m|>�w�����"�� �;`��4]���]��7�Wv�%o���'�%���d���J�o��a�6�dֺ_yR�}�H{�����`�p)���3"�a�UCNRLF�������|��(�xU��V_7�ф}j{b� ���O���w�GU;��s.S�m	mW[D�L\ʅ�4}�h�>��A�؛������D����&;8�Ōdc����5%_�L����) �:�[��a�0���sg�9�����۔ǰG�t�C�t�]��>�يq'J��a�I�K�f�f�X^lw/WK���3Cd�ץ ٺ$�5C�({����;@���Z������Ê��-h���<�'�K���r�o3�J.N�id��K��?����ߘ5��PiOՍ{�����5:~��	Q&�ʏ����d\�E��1b����
�CVR7��!TM��맘	�	>3�>�����oM�m��2��VG"L��ZOد�y�Z��qFd���$�1�^pÖ;R�fGI��.c��o!f�d�H2h Yct��o�$�
��C̗��z\��=��t�DY[����g������p3캝IFg}E*�Ҧ�����͏�K?XԾQ!nu��ZV�B�ԯ�>V �$VOuY|�����=�z�D�5&�+�RۀB��2��Z�lu�B�O��x`GOb(Ȑ��j�j��z\V�l��m2���Y)p,���`��;E��	�r|Eط�M6�z OSTc�|�$����j>�c惀��}�h8�V-�E�ϣ#m�}�j �6�T�c�1�O�@״l�������G��V��'+R�q-$1�I���Z��Ph!�:��X��0{of${���0"i�̞����+g�n~�4NZ	�������d��'��̊�3w�	� U��co�����b��L�ѹjOV������.8V��/~��
9��@�n#~�N�b���ō�jdn���lm�=߿�o�Y^�*�H�aGQn����[;q(�����׀�Jgh�W�Dgj>�:nh;��
�.��[b�ᏼ�6�8��I]rA��`����|[��LGP��}�d��\�F�?�]$Ud���h;���c�q�(œo����"i��l���q9��rXG�se�jg5��������WB=�n�%׏��u�r��=��я�k1�A�T�8X~��F��6S��� ��dK��tɸ7�Rx����=�E���>���\��i�'4�T=��g�`2T��#�ڨ���C,Q�+�&�M�I�T
 �<P|A�1�9'��lqY�~��+`�4���1e�v�e�[�8��L�W�_�^j�$�)�t��ŪK�O�R�4N`�U��z�oC��'H89uL]�En��vC}�:�`B0���J؅K���1�A dG��K� �Y)R�o���?�{��J�?u���Rތ��r�d�^���x�d���kcʽ��/�M����D?�'DHbP�(!�cS}$����b'��٢�>��e9u����i��y�O��d�J�Ԓ�ъ����,��)��׫�;�B�[��Ƙ�QP�-t[^���U���B4z�dT��8|Y��˟^�3�?T��᡽�+�f��	���
�+��Ƒ�`��tP����z�GN#M5�����ʇL�r��?;&�]~�Q����D�fY;�PU͒߷Ө����.�e��>��x�rA���e�i	�R�@�~x/�8�J��BW\U��q�6�/�������'�u�ƬT�騣��*j,j<�U~�b)�1F�J��㯎�ͮ�a&�l��W��w�1Ԇit'?wh��d;F��-m;�=��� ��Y�(�_��+$��/�7�LQ�_)zq���y��~Pt_�l��x�甿$5��o�dS'��/����]�w���������5`;XPf�3G7�`H	SN� <�C7��t��/��gٻ/|@C���לoMc�aH�0[��ݝ���6��gr�>�>�`E��+u���2��a1X����� �c�Ym` 2���f�2�\�xS��<E���П��>��84�G��:�y���9��Z���w�t��<�a���%�0�`̡�oA�t��� n�E��%ޢ�U$�������k#�6<�Pʮ���ث�1��s&�Jb��J�@Ѝ���+}��5L1�����Sm��R�nWr��dϠ��\h>���#�˓O_�Ɏ���_ֱ^K��$Qy[��&�P�ݦ7ρw��#�(b���d�y��}��rTf�tM��4�۬�7Wm�K��W�,���	������,��[��x7��ܹ�r�
�N��1dL�i�0`��K���j�'T�+�$B��i�^���g�b���I���EAWo
kit����K�8�����5����c@�&KN��!q	���w������=՜�05��X6����q���5�j`O�l6�@g���")W�mn��	�w��J����\>��� �2ZO�-F�Xi���b�p�?�lWZv�4�o-�XQ�����C?)�c|$�G�qk�'��ݪ��|�H���,����"΍�������kƝ[���I}6�m�>:z�%�\S�T���:"pMQ.j?V�>�*��]E�}e���d�ʉ�0ӝ�j�2<5���1�mhI�`Ѩ]��F1�>��	��Rj1����{��BT�ct
h��z�qڡ�?��ub�,f�ttl��u$��8��:#�Rŷ��;Lm�p�6d	@!�o=����s�"`A��[ţ���u���K���oQM���6���{�n��E�Ǭ��ZDl�O�g��<o��]��2����6��&_�,�0���o�� ����t ������;�͜��T��f.�)�)�D�>�$��s�5^�٘ǀ/���-dq���p���֏�@�H1���e� @����ѸZ�\�&��t�V����ݧ�ʰ�\L�?��+<�T�6���G[���&$�8���o���\ѭ(P� ���51�{s�ǡ������M� `El�@�ԥ�Q���A,g�<b�k�ڿw���B����T5S[���о,��9!���܇���.h�ǆ�b�p\����R�S)�^ �
[��d|��.h��,O���LA�1|����Y�q�ڸߐ.��F�_�~�؇U��z����t���e������9��^�!-7@���n���<�itw+����k�-9�;���3��c��~��Y�[6Hs�ެĖ���D��K�(N��Î����#��K��w�8����)��{MA(I���mt�v���x���5��3��s�X��(� _"�W��\�\����� �Ⲽ�W>�����8�H�����=}R�/�A~䆊F�gQ&�U��F&O��䮩��ės;�;|��֐�-PwKB�����3w�䶥5XL�D9�k��?p"A���X��P���yi�֦� �)������v�4�v0�^�13d_��o��x�r�̧�������Uᦐ�i]T[�u�K��!����L��uF�r{��������Q'��a�Op�(@GUQ{W�zC��[/م� Z�I��*$�����4�"��2�~�9���SG�ь�y�m^�FxuB~�w�?E��
�=��C��ںi��Nf���+��2�?���H8�e�v����y�pc �He���_�g*^r�"��+�Wso��FE5��/v�W�c�x���{i%\�$R~H�%Y�	=6
����ޫ�-e�C�z�B�D�%s�$L���+�IK���p��R����t&�Ѭ|zZ��j,��fD.��8�A��J˕�/�88�ߞ��8��ڳ��������A����[˷8��i}W��(��C���I[9���n����su�(�o����E�ژ�2ďb�$j�7	[2��={�C���(9
k�AM$Ᏽ`�CX܈T��P	?$�޾���d�-���n��)��ɀ���-��{̄���e�B�4F�~?F�U:eS��������6X��%��I���[h$���#�MwH�?P�%�h1|��O�Ԋ4J��ٻ��{B��2:4��,�aj�[��A�?;�	Ws*#Y�`\���� ���kN-����ya�*	 ��4P)�2��VRR7�D��֢����4�H7���5�j]�|�9v�g�^5ȯ��y�$PtW��{3o�
��7�v!Ђ�U����;8��1QGLrA����gw���>g�BpS+�Ɇl�+��R��M���eM�P���D���o�����V ���49z�kX%6�=;������t��,��ޮ����^P�rhI!]N��E��4F�ߵUc�c3%x��X���V<�2��5�=����)��Ϛ�����8ȠzG�+�7a`���C-�����e�����2���W�;s��-��/Ycé
�!�Qm���� ����k��1�c� /ޱBt7���z��oϖIhz��z����>��kK�E]�8��oh�~�r.�����_��#8������C���I��[��O�]���&��l�����ԅ�Q���P��� ��`,�
lKc9BV/��6\�CEg�p:���
w�h'��`>su�B_G8ɈM_��Ӊ^���Y@�3-������Px�Tx�i��ƍQB_���%xɑ;�+D��q��_�E0+HՖYCk��	�O�1kM-�i?5��1������lE��Q�p�pdsE�L^5�^3[pQ�2�պ4	[��T�:8x����#��*J|����~$y�6B��C�1����j�T��I��t�a��	Bt�]�4 +I��c�((��b���=l�ԸE?�\:-F_3H�ZȺ�(
鸼 |�ˤш�H_pi\�g�(� ���W��,��,�k��Lq�p��?��
j2��U �>��J��I$&�)�Ԑ=f1A���y9�^ȕ;t<��~|�t�%��`1x�ޑ�_��������S��,�N������*< �@�2�PCJ�ty6������K�E���yg��������؍�G%`IΖ$ʾPf��of�j�-�kq���a��w�-�"�x8/��zI��/K�7V��-�����ٕ[#V�,[W�`�Bg �6�-c��P���w������5��)�X�ɠ���c�����Թ$���T��#V͙I�.X '6�[�}Cؠ� ���!��6�OU��n0��D/Ax��-����xh
��s�&U<[r��8�J3����&.����-����
c����]m^qApy��%�i�ϵ&R^U�m��@�����fo�a�'m�
�Q+���y���,'g���
�����֪f�;2��/����a��
����t*�}6��\�+ߗ'� 6����g��^�z���pQ��0wA11���Duuh�>R�Ą/e���{L��D����pv��@g�⑮�j%����z��4��]
|�+�\U)e��s3ӕ�[�C-�v�밄���L�R�Ku+(ٶ��N�I���2�c�j���7�`O�5�9�a����}�5><x���t��'e���u$����K���4�ǒ,7����?g��MR2Gu	�[w��;�J9������<�:���j�/\��v�dfp^�M]怩��'��^��A��ۛ�k�@�2����{�کSi�I��*r�N��~�����mFm�s ��?��#�i<H���T��:Q�s���v,ww�-R�r��ؑ��b����]�O���(����%E|i��e�PC��=�F���&�K�����@�qE�����(����^&Ekz�F���/�$��!���g�F�(U��}0Q�sH�|�|�~^���mL����*�{;4?n��'��\YFL��D1m���f�n��4�t=sb�0s��H`�or��N�^�4c����A���x/>�+s{�!(�k10TD���|SK8t��!vT�2���Hr�m�H���p]1���x��3�0�/��r(��B h��W`.�;�l�H�ٔ#�x�sw :�#���Q�Ď[��;���o.H�I�o�ʙ�`��e)b�w�������]�	�|I R%*�;���B�$B]��k �w23�[C[]��5�
��U�k1O��@��L�<��^�Ϡ��*C;��3S4$����U)�֌���!�iE���X9����~�A���c��n��f�dŪG&
Q�qA'�1�ˎJt���|�N��j�ю��v��P.�۝��G�>�,����$�$$�h� n")�\�RT�`��uq*&n̰L�㋼��}Un�p9\Y�\/s=xT*��y���ڧ���X���SPbO3�`J����G�I��a��|�݌��A�#�t6���������4�j�X���x��٭d0e"�1(5Y���6W�v㗃���7l|Y��v+�4PYI!����s��w��K�:̏�#�Q�j/A��ڵ/�	i��@){Q����G����Xy��%N`8��u���X�]�}"UY���ڭQ#a~%������;"To���P� �HF*/7y�`�C<�״g��&"�x��|@п��j��0M�\�	�8���lgw��c�Dc�'���oa��r�	��=e�.TQ��Ì4��ʆr�?��b�q��a���%��+��p-ϝ�8�G��[��A�^q!G�� ��d��*��?
 �1f�0�l'��u��1��ya����-ġ�kc#E��!D.�B� |m	we�E��y��s���w|��'8�
O�|��}�yˀ'��-��*��+.�6���'�70��#0M�(��jU�U{*z۸�n3��+�`�������C�cw��q ֓B�[Y��g`���W��3��Q��[�1��n%���= kec��<L��� X&kL0��/��.��2 �U0ZR��R+�'5���i�&A(�^�,�ob�t�7y8a��D�C�l�z�tw|�eC�j�T��-gԃ��;��E[�v6��|��f��6��b��!�QK�%��p2	|����u�ʢ��>>:]���)`C�qF0�47WV�x�!�#���,������)��n�O��u��5og��t�´~��Fɋ�.�m
��kH������N[q���* ����㹗=;xZ�\`����p����35�cYKm��);Z�)؃ԗ�4��!P�m��k��x_b[���r��Q5t�y
ui/���c�_x}�x{��c�� Qy�
r��-U�§���Q��>�֭c��o�[��Dz�ت%I�6������r�+Pj���6}7G�_g�["z��M=��N�im�������&ǺÜ.Y��h*�{Ǝ�u\�5�HȘsv�=w|@�W� '�8����r��O�MVj���>����©��	�{�1��?��J��&)���*Q�q��O�]�iM�9,۴��N�x����KVJ���r׃�Pr�u��.n�Hf-��9�Jk���m|?G1!|%��G؋s %���ĝ�I�QO뎺Q�+���3g����>�k�'���ߓ�I�,�5h�� d�s�h�v�u�b��\���yMD�#�`"IȂ+��F �u�V�dE�W�4ޏJ�E�:b-�Ň���������J-U�<\�����/դtӘX�O�O�̲��f���Y�Jd�Lg�mኴ/)�"�L�� ���8��p[0��� �� _h ��۫�����kX���A��5iPR�z\(XOCK0q���y���Z���dC��S*� �Pc��`��Vvv2'+�ো��*����0�eD~�0�����ƋcBh'�9���Toio��w�p86c}����]6R��e �i0Ii���G�D�RS8-����:KA���Ƿ�c�ޅ'���Dr"˶�R2���N��R��E����:�i��Wxf��7�%:���r��h��H� t���ؿZٟ&tj~���>���Q��
���������'g��Rw�Qۤ{�H�����D���f}�Q?���%���M�T+�'s
������֝buz򛅀�ӁHh���R5)H�7*�?:�n9	�Jz�w���(�x��E6ߐ	<�fU4Sk2��p^?�~����h���g�t�$��-�O�Y�E�7~�2�8A�gi�$ֵ���a"�W�{��zӘ9����ʛ+%����N�RE6�T����g�\����'xRՙ""�`1���x%?;w��=]2\���Y8��?;_~�Y��w��=!�c�}�S�ͣ�l���AІ��B|=7�n:�gV��^G(�"O&D/���+��kF�m*����17*���/�	G(��mi)���p��N�a�[|�w�����nvs"m�)թ�F��AR��ThV6�DZ�<�:�Ş�~�۩���f���m�U$��I��drS옸���d���B@JK�ӝԵČ�(U7��ѹ=n���%�+���oo��$����g�S��%�ۮ�?�仿ډE�enY5ͳ�=����4Q�#>.u����7ʠ-�֫��h(Qh��c�V�T�#-T���2"�Գ�ʫ}��Z��,|;{	���rѿP-��u����<�m7�v@�D��]����h!B�#mCo^��k��G�����/h�*k���5�xf��Kt���?�
��[�9�!�?m�w4�B(��>�m��n�5B�� �\V���B��p���<B��AC��ź�k�q݄���\RL��m�9���ED��"%�Z��>�!��W߰D��G�%�����d�/�l�W���эڇt��������
�C��Ч�� �nme !��+d+}%UI�3�T�� �5c�y���2���L��	T��ż\c�y��<F��n�H�X�d��ڞ�|����W��J~�!]�j`:k�^����G�����E�Jӗ�|+A�8��D)�FV׆��5ӵ4Ԩ��&�A���Qu�P��g\���i^{�㰖��m�p6C���c�k^�	ʾ ig���<3_�Hf��[��
�E����C��:�JwF�^�ѧ����@��wd���hR�JMK��[
��-&GM`���h%D�Y���7��D�M��5=�!d˩�@��^�>�Z�0���LK��ȃ�=f%�~>�B��>�/�vc�����ￌ���q�\������oh���j�q�PD�%eK�]!�s�q���:��#?B�"��e'm�u�C��|:F)�I���,�7�Y/��D�9ꮽq��l��!�ee�����l��9�pmY
��r��q�_(�� ��������c��	���
�mS���q���p�o�����3��ӏ��QUw�8tE��]!��Fru���һ	
���3�%�($��m��enj��V.���֒��ݗ5I�m���n��B��Mx�N^j�����cЙB�ik��W�ql�F���1�"%p�ҩ!SВ�RJ��JM��e��K(��b��h��ȿ�p�����=�q���a�0x��I�Q!��%
�< �x8�j�-�U��:�vԮsP>��R&����8�������ZR�	N��.wO�"|�@R0��K[̒p$<�}s�6>�h�ו;$3-��yd*�N��d�P*�Xo��V�S���Sп���N�h��� 8�3I'G�&uM���T��B2e���&�>�ԵvD��
�2�Zl��&��yS���`):(!H�C�����E✂SVi���+�C�2&�S�N�b)ݶp�}M�g~_�Yu{�:�M4D�இ3A��sCkv
�?���mTIC�9�geX?O���Ẏ��s� 5�It��s����"��X��e�k�+c���ȗY�,k_����]�k�r�Tu�yY^�@���mפ�#�NI��fY%iIb�C޼�!�P���"_�9��xb�y0��L�w����qWX��
�j�2��͍��a1����-»
Xr�c�]�=�ε}�(a��x�Y>Vd��`Yͧyvn�W�*z���W&V�@���F(��.�{Շdf��ͬ��$��0��̈́0��	ɺ�+��� ���j�VC�z��6�O'Z�W�X>�I%��'9)~��p�4��+�c�:�ؿb����nɂ��'�"�~aƝ�3ݠ�q�EF+�:Q����CՈE�~�YH��	zk#�cB���w�1��#}��cY�3�"�8s�nC�D��u��rS��z+Z̻*/�	���iR�C[!O�cĠ6��	�5lc�{�NR��cڠ:2�������L�c���I(��P? i���Tp0y���@�G��I8��ϾV��'D]h_��o>�
ÒO�����q���iWN�|����!ģ$fja�L��������Qe1	�
;�Adϲcl�T��a�dH�ڵ
�aT�� I����(��x��	V�@$;
fd>�Yq>���7o�z����<ss�]�f�b:?94/+<0��o��W��M�:S�̳U^j�nn�΅>̩˾��4�=3�v�q�SS��(d����v�:n2�O&���0$��=���;Y$c���8�!2���ޝ\_G�x�n��(����-���y;����5K�.�f��|���q^Պ=r$�����Wż_8g�b����C�T�A��߮���y���8�Bc��w3�D���8 ��'�+�JI���LN�#"�� ��b�q/��uq��%��ѐ��~��u$��v�5Gpʹ���9��B]����"�9���q�� d4���[��{��ONS���c�Mg�X��nˊ��
�'�U�+�p���|��}<[����_/��ߣd���ޟBA�C�\�m5�SBx��K	Q�������,��y�yI��6"�N���w5t�Ҭ�\Hylmф.�܇f ~k9;R�E9	���8��,��b��U��8�_7RV@��g���4]�Q[���1sRV\���2ͽy���q@��C濥*�ޢ!^����$�ιB�� 2�uy]�����K��Y
<r�˛r����\h��Laݴ�;�����OU�ּ�&#k�
	k�&7��b��&b��y�<�O��0\/�9B�S)��C{\�๔n��=WO,J�?.�����Ʈ����	a��AEwk����7K�c��� z�u�n���Աv�i�Q z�T?}
;,*+��-���¿ᆝ�-��V~���o�f��U�آ�mX8�d�V�o���1l|B��@E�H�B���Ҙ�_o7a�ǝ0���3Y|Ȧ%%�t�<PG�4N���D8j-��&��G�\x���M��-M�
��\z�g'�I�4ʆ����;P��Y*o(�e�Q�{�S:�P(>!�.���)��K�40"k�al�g����/�JUW�6CL��z&�)����ƭkP��V��>�\��H�C���k4k�P�".vV��*"��6�,�QƼ[1�e���đ���'f�[dvK��B�s�����l�����{#� �N�����\��ׁ;�����%DU�2N��Jk�(��Z�9�r/-�l�A��~0�!��-��9ݧ��P� ��L���=��I���Wilb~�H���#1����D!g��)ǂ-�.���A���À�~��c�\US;Ţ���q'f����d��6�T:t�Ix�.7�z�Fu�r7Zg�E_��n�_��P� iP?�*����2��?��I���E�@"����
��c���L8�_�Y��:�u�'_�����,W�u��ع���˱Y���d4��m��Ӫ���~���������@%��ҋ�֜D�|y���� K��>��}��b��ԸQ��'Q{2Y��c�a��.��"iX��^���Kq	���bQ���\�}��V��}-|gm�	�]�`�eĭ__=��d
�ƣՉG����4d�� Zתۃ��v
�UI[� L�|��uOP.I���l�7*�]��E�m�	~r�8vW<N4v�r�-�)�rrR��A�l�l���`z4�cܦE���Uʥe��a]V�=�O���L�u���z����R���N��3E|[L�c�WMp&ѽ�u�(a�$KJ�@G��|�7��P�2~�xq%���Ai�B7o��F�nv�Y�j��/�&y����sb�D}�K����?t@Ɂ�Y.NN�ѝBTO��WO�C`'��n���E�ߠ�ȴ��e�A\k
������n ]ښ�F�Q��u5�]v΍h�D8GOA��h����j�(&�_[�1U�R6K�ϯ����c�b�R�8���Z���?4�g	c���/JC_���3�%j�p�㙐�F��B.7�Y���B:S�2ؿ'#�ϛ�o�� k��os`g~��C*��^�2lY�|u�p`�o:mv����c]l�u���d.�]Y�R����L���6�@��F�5$*n<&�ư�囮ZD���4�,�܀����R��Y�4�ލ=U�zͽ�\m�T��lWN���%(��f^��j�D�l�����u��`��s�:���졈�h�eQ-�H\& Co��W�Q���i,�B�0��"i���Ԧ=2��(SM������d������X�R���T"	S܏���ɵV�h#���,�|�9�/�q�C��&т��d��R�T�DmR��vӘB��5���������lsu/K��80�׶N�$���p�a�#G	ny
"Hɝ���T���K�^���GhN�{�KU\_H�]��A�l���m�&�]�C��A~ ��oYa�|5KT�R���̓S~����Bk��8�iW��j�����@��@�ȵ'@t���^t)y�����rE��k�P-'�?��)~���!���� (*9� �����͊f��.J.���V�u`�w��K��=����y`�
�+H�1辳A��X���rm/�լ���B�m���u/E��^u���2F�mI��]7��.�������Jh2Wc��;��&��������;�:-Z�e[���rG.Ls-�`��L(+�Z���e{XH^*��d�˱�쿖��͓�'��E�*�zԯ4Dq�$�%��]�k�=@ 5P�P�
_ڧ�:�e����'&��Th>�)cAC�y�Hkʜ��!��JM�����UNp/�f�a�
u�Dݞ�O%'g�]j��p����B��58�j�:p>پB�~S�t{�u L��c�T�|j�L'��h*�0�;z�rM��x�!5ధk�*h�Q�zu�S���P$����+z\0���Y).a�7"�9�Ѣ�_������T^�����gUd�'����N{��%����P�_jh���cbWVʱ\m�?���d�1�/�%O��"}����y�9����g����(�d�Ȼ��K`J��|��s��fF94DO%ɜ��a�;�˫�}�>��`�KP�&��(ڱY�C�"F`X�����.d6]�8������H�������Pp�1M�����;C0Ըy��42��Z���ْ�l��x��+�ś=�A�	�	�1�"�0�%T��dk�#�'��@9��uw��b���d�A+�u�g�^O�s�1�MDL�\꒣���0�m���aou7z�B'��.�[
R�oIƝ��+P�����ʺ�a��3!��A��e)0��Z�F�z�>K���b�X���=Γbkͭ��W�Ų�I����=��k�y΄��ٲ�C�]qy�;Q^fb�2m���Z{�@�u�5��̃�*�|H�i�]����Y�ڔ�D��F��#c䩱9�hƤ���h&�����W!P�����v��-E�3�Ͷ�#~�����鶌=���ְ�.�'�����L+�:S<��4��B�Ϸ�����m��x�,�T�H*�4�I�M���~�y�Ȱנ�A�W��+C4f�P����,R�5��(r1��+]D������jo\�Ot���D�x�H�=�H�9���+�����%u<��<�~&��qc����/	,�։�)�#��f�H{�9�'��ÿ�m�V�e�K���Lt���L��!@tG�&.��	/F��p�~TΌ�%�?���i�)*n�=�1&Q�Pk]l�tR���EI�^l㓐eWy���8^�Q^8��y�ʅ��+랁��(�-6.$��O6<1yK14s�h�b�K"/�󲽼A	 ��/�����THBT��g��Z�Q�y��,&��0I�l@���]ٻ.>)�`W����V uS?��o�C�k����6ޯ�֌��.���v��`�",��4���l�������D{C���Fu��K���S�i����b���B��ֶ$p��ke�)ߦ+;���������r%pۤ�+�7��V��ˊ_�)Nb�'��s��E`=�-�N��P��H}��<'�����]|�=B������ݱr�ZL�Tws�ƅ*�,�������L[��l��@}�{*Ŀ��Q�T'o̢sa�R0;���l���S��gZǘhT��R���˕�10����w��Ɔ%�1���1"�n�T^��n<
�³�@�N�^��U�����Z�Z�r��/�M?ki�_{�[b��	�`:�	��W�����[@�"�û��4��e����r��y8*���V��R�ˬ6�Gw�/��/�V��ϵ�O��<�
�j��~���3�W<�g!��"��*i�.�Ӝ�s�+/�C����E$UkL�jD���X��乪A���� �`��Y�g���ze�'�5ʆ�m_}���MlE
��{2�G�A)8�
���H��c�>�9[�]�m�s0�G�૥��9�9BM�q���9�U��*��+�iI�8M��}����=Vc�)��w��rT��:o�@�S�4!\�;����*�A���0Tѿh�آ�OB�>�� �cAj�ab�B:j*��v(������r��XU:["&h$a��&L�10g�"��q����+]m+ ��?f�=�i�YW���a�ӰI^ϱ�[�+����f�[�N�R�K�[,�!	�||X�6�K8����s`$�{\[��c�
ZD<�;K�G�};�>��d=�V�8/R
o{$����f�MR��p�%�Q��V���7�C��)%��"X!��|}��,��xB�����|@Y�_]��U"���7�K���~�1u�3F�L|����b�x��#ʎ�JzH�0�T���bV�-b�_�\��ݗG�� ���L̢{�gh������n=��ظÇi�H*�lܢ0Y�`�a��X&��qnD����NM��"=�@ ��=�+����t�m6e���f	�R�N�%�V\��-�h�l�$
�����,�����m`���@���q�r5���%�����ܷ�g�L{'�|���Z����&WadІ f8\����5�n$�w@��D:A�D%���������6����X�YO1�E�(��i��z���x��N����<�[:eI�c� �V�8m-W8z�mƞ��!R�m���J��j6_�Q+۹keY��g�ݝ�N�F����FB���I������#3��B��*���e�RdNB�	����M�U�q�g�ST�[	@K<�4���j�2d
�Yw�HK��z�tXK&B�l�̏�+b�C���Vt&�Xt8E�G]��\3��=@ z��S ,�VFF�];������۲������D��j��-){83=��I��u������WB"��}�[y���tjb�;�7�6�l�32�%eD���_)�c.a5e�Mܢ�Q�$B{-���\8�����V�yO"���b��E��"� `�$�J���­�/�62uT0�F�0��>p�܀�9���A悏��É��|lhbi��*a�iy�1)���m���l��ؙ[�~)�ӊU³Щ��Myu��D��%�YK���"} c�`V=8y	Zy�g�ߖ/s��`N#����^cIP�G^�p�Q��.1�M����#����B#2x�7T�t1�s!@� ���y~������H�5�#=�,D��{���0�Λ��]bX��N��c���7������z�FT~6�I4�b(f_�l�MJ���zy����#��QTZ�9�j`W)���.;Nq����/��\L	,Էd`|I�8��+1�vn��y�ȑ����z��f]�F�qZu���>4"Y@���*���GBKٻ_��U�)�Q�G<�i�j��t��L�1�&;G,mfGq��b��s<Rě��5uA��=�\I3�� ��?ΔEY�;� %Qz��Oѐ>uu��d~Jyr&Fѓ�H� �9�����U�:,~$\.ݫ=,���I3�\)K��5����`�q.%���&s�U6��FW�7!�xzW��l{�-�Jv��
cR[�s�
	r�i)�0�GvD�;�!��M��1�kB)S}�A����y5�I;U��!-N�x�� ���)��J3�|�+�U2W��$ �Lv�l*�T�(Qa���	�����Dv8�b�o��.��'����U<�.�y(�<i�8�ZIh��ܲ��=m�7܊2M�I�$* +X_3����05��Xod��W��w�`��$�v����Vr���R��o�k�Es ����.��By��3;�GUBy6�7u6~3i�����Mp���S	�jm�}�<�d�V��fh2�N��N�c���M��5��͖���k��`�6��5h����腷�jq�:E���6��?ئ|o�˞��[����������@�j
V�+��p"��E��?�4�N��Ia�t��	xr ��rR �r$�Q���ނefǢ��S0ϓޢ���0��e�?�a2��H3,� d:��U�$<��o�~��|�gC��3R1�_�/���w]%�|���s��a� �A�"��C�)I�ҋ��Z� �Ż\���Aĩ���;��l��=���
�?�y�����r�f�[rϓ4u��?��}��F�Tw�G55��qq��.d��~�B���a'����8=|'	���7�8������R�\2^� ��I;tT�qk������ʛ'dOH���2�.����������	`��2sC�yUAGap�x"'����u�G�/��Ƒ����\E	�t�	��=j>���|�
�{f�/�8�k2S�d�;9�@%�0H�ê�Tk�<5���By�镆q�l@�ezcgHIoU�B�:�i_G�ÝϩrN�a��$�7O\y�k|��>�1�Y<�+٦�ov;Hj	d�����R&wI���VE3o�f��Wg]�[�}cQ�T�m�wi��d��Po� ���ڳa��ZL<#�TQ�L�H�*��@�JU��=q�0��QC7�8m��"�^�IAD>����8j	�k��>%��+0�A���~L:���������j�_��y%YV�|A���xd�tM����Q"d"�yؑ����V#F���)�0k I���j���M����P��_PC�ʞ��8����t!���d�-P��]�����*D��^Z��"����'Y3s�Q���w�>>�
�:��p(J��|J9܁�MzDa.�$�zߞZ�s�Ⱥ�d���.��$�n]����u$R�;0?��W�d!��o�Wiz&�̙R�1q�_���Ƭ�'���:'�'>3�GM�_m.�Ǿ!J�A��=�rؤ�����\��e�hxB�����)+�/���j���������a�j�q����Z���/�A��[���^��`�E��1��e��3aD�Һ&�I��@�T�A�q���8����{�H~R�Y��J��5�|u�_=0���&+�a�-r����s��*K�YwLhA�Tv�g5�Y3=�r���#��F��?n�sD-�ާ��XO%��[�"AC�ʔS�VW���"/#��e�Q�%>?�0;���TjG�>���=?�"�ޓ%��kw�]z#�<|�ʄ�ۓVV���D��2����sّx��^�&�m����1$:�1��Y�Iz�M��p�
#K��`I�#�{J��G��J;4����ї�'�'����g,�V'���8Ip5�H������s}��cJRF0���K�	���7��I�����r^yS�8��Ɣ��ٱW�J�l������'^���.&�1�j�����D�	�6oпd�+d��P�FD�	$Xf6�!��Y5��Gfj�V���E��k�N�J��Ct8�M�ܸ�ɮ7��^�&�{���"L�&Q�!f����1��;n)�k�Y�櫯ÄJ���)���)����*��E=]��]#�Qn��3G����Y+9������AT(d� �Ck�f�ɑ]�O]zqk���
�����3��M�W�M���]�U"�א�3�����Vc� fv�2��h4��[�)���xU�*�8��A?��T���~E�
�%��g�/<����G@F�d�I����Zp��d�����O���v6� ;3 2 W-��i��/hɷN#�`�t�
>�gS�m���%|u=߆k��dʠ���S�3J�/�B�ɖ��T�dBRS��i�Ѹ,��q��a���^�Ym�H��pAh*�j������@�1�b̈́�D�B�x��U���|����HA��Tʟ�t/@�H;,f��Sƚ���<e{BΏ�ʴ ���jKv����Q��u��.�����#�6�R0�ga'�\����W=0]��Nb��O���'���+T$�������
�9Y��
��iI
����W.Ϸ{���.�4�c�;H��Ȓlc�1UJi�a�}����e���Y$n��ͪ��4�]k7Q7�O|�xq��y�T�2�X0��n7p�k4�qSs��U!���k�#1�����w�ڿ����x�V:�^cu�^r q��KWSN�Ze/���,�����b���&k�1p����vm�)ip�+oc�D�A�r�Y3jl5���k8��.�^Ǘ[�E��߈U�x�F��o�D�,�n�@���u&U���5	ӝ!r4�atޠ��:�t�Gx>L�ԩAmc�6�'R�;��VӼ֢��ZQ)���g����8];&�H���tCBD �եbi>c+�T5����u�z0�E�����'5�.���#�ҬnG��

�
��椾`b�����=�x�Y.O��h��4<+�2y����.B�!XZ�6���Kj2��.�!�*��^)�<���1�3�pPƅn�ɯ����&�j>}�M�L,?�����~���gT@���Nmv1Ch�i���]���x�0�׸�����z#l��.�+V��w�VQ,��?��s��-�RiO������0�$����T�sg���q�[�>�M����FP7g�-rڛ�� E�:=��%!���%���o��J�E�L��ԍ��g��f�p�(��ǜp*������]
ө�D�$.�Xд������>���Zf�Ԗ�h���*�]b���?絗�[`�{�u�g��t����C��;Xm�%aW�pW�ZR�d7xTmq����e�?dq��4�T�ў����X��1;*�'^Eq�O�5���O*#th�F����0D��~Q�������b(V���P ЊG}���eGV��
��|J9��1�?X_L$��JY�4��l^:W.% ��7�'e�UZR/�$����,eŹ�1�X�0C�_����'[�l�`�6����F&8QЬ����h���h�	�����cz P��>�: ��t|]��?����-bh�?�i������i�ʿ,������"D�z�&"���K�fP?�]�p*�~�+�����\-'l��O���E�S)��S�ͥn����a�ko#Q��&��g�4�o�W"��N�Pr����-w���ո6�;2�J��M&��B^��67��Xڶ2e�F������ڃp�z�kq����.�5�E��0&/��:Fb�1�*��J2P��<��FC���0��.�7�q�7#M= ����Ҽ[c����:0��o/]�z�e�^c���f���MB1zr�P�+m�q?7k�Q��Td�ъ�e|'����ށ��얄�mټ�)�U�
�t�\?Vb5�&@�5���}��0:���5)+��v��k;�s��sܱ%>��C�n�|�/�OM�$z�d�/�ȍ���-9PB^�x��l��z���''�2f�l�	��i*�*T�O9�S᠘���&���Mn�K�.%���.�z���ƿ��2m�C%� ��h|�6�;V��8ĚB��tש���|��ԗ��Kf��ނ��wlZϙN�pn��b%¹u>�W��^
�x�E��(��*��O^�;����o��#���v l���{��Du�u��o<�*�ی��r3@O�h�;Ӏ}��8��s�/��n(�\el���X6����Bn> ���hw!d
�y�is_&�Ά���P���b�f.�]����aG��U^wK�� /4e��7�ڶ�:�_(5��D���v��]�K!��ը��CRVz�v�<`�"(�Xi��
��m9��LY6����£ȉ�.���@5"C�ىlU�d��lBR���ǚ����<�)�7��W�O�S�Hc��y�Q�.�F���?�} �E��E�C���?~�]�-�W�穣"��7Z��U[]�#<^?��?ɴ	gHZ����� �x��@���*,�ɨ�!�'{+t�XG�M`wHd��o e����\e���N�{�[̎��2��]�8�m6<-} �k|��%g�qJ�\`U�����1 �[���t�UX�>���>�*�tR]K�t��)k���֮N>挲��S�<[޵D ҧ�h�������2a��$����g���qԛ��帔z\R^�6�<X�K�f����)��֛v|��j]A�H�T�'�(�<pY��7�<��X�����Āt�o(���iNJ��>u��Iq�)S��2���d���S�&c���f�Q=%�}��.���9�D�@�5��Sɹ&�
9����9�=�������)	�b5	��z"��ή��8����>�jUn����:h�����Ut�'�i��9U��䠆���wcv
����	�30;	���ѓAQb�i/�YI_��h�����A�[��2�x�;^tqw�����vr�%0i&��0d^W4���^�~ph\��Jl�y%gbѻm��q��B���1���+?`�J���7nt(ݽ�y�鬼u�Ϗ�P���i���a����6i@R���qX�
���1�$�e�>q ��eAF�>��"�
��?]����ǈ\�̑C��kΤQ�/��2��D�pv�\�nH�<zL�.��3vǏ���=;���r��K��s�0��iX3�|��sE�Q���JY�z,�j�ﻳN)��4��k<}��ܴ�,�wls=�;�s�W�zn�⩿Q�e��eL�v�9x���C�'��҇�C�+���1=/�n�5����ª�X�*k��ѿ�(Ny�n�d�B͐�T�]���_JX����� hk�@�� � 1,����`5rIU0��57��F:�|9�f���l��I�F��|��Wu�C����rO�*�_�|���3t (���M��ߔh{�3Nng
H�r�"Z�tq�e6�BD��ڈ��Hg#�3���1��蠁�V�xʟ�[�ֲ��nƎ
Nl�S��,Қh�{��M2'�!��^��N%��8���# !�m���?���y�߰�Go��X�l>*��E@�v%�}�ܶ	6�M6�*3>3�{G�~g%��̊����Ж<D�d��)���@6*�6az(0��\��t�Er.$P�M'^����W;�� ?.3��}�x�-��~�8j�k���#(ޝH�΢��?^%t�
��}� ��ˀ�r��'2�a��>,��6p�qS�=�� �d�K��,R�K�������v=d|�4�O0��l�9�mę&�,Q>>,�/�N\,���h��{�$�iNv�.�Hv	3�a5��p������4���^Q�[d
��Y��`Wn���W���CD�u*"2�q�K�"~x���Y[�ˆ��p��j�����Ƭ���8K���� ��
�P9��+�];Ns�D�FDp�w2%eu*p�>W�͋ZK<�3��� T�fΟ6o���*�j��
�5Ŭ.�Z�%ۣ��_�іm��n�z�p���-'\��I7ֶ��څ���>�C)� ����Ga�v���
7TP�{��������gT�ݣHA�s���1��F��MB��A���=�d�����m�y��pE+f��t�ѳ������>��g�E:ڋ�Y��T	J�R�L�����65 r �Ql�ߛ�S*��o��yi�n��[����<��d���1���PKE��C��4(�ک�fe4-��nfjy*
iר� �����\�5x�]f��2δ��)��%>�M���es��jR.;��c=I"j��vK��Qԫ!�,V� ���������0@1��p���2W����� ߋ�b�WRAq$i�g#�|�ڡ���쬌]|��K�T�sC܂�`>��P��}=͑S�&��	��i�)u��R3a{�`���nV�9�| �t�<I�O��i��E���O�Ě�Pf�H8N��DY�����5߳�{����#`M��뫯-Z���$�0΃�嗙^1�O�	��@�V�EC�nǩ+�snP�����ᐜ�����߬,؂@�t�Z*�ėA�ch��������=YZB"����b��{�uZ����AWɎU:�3:���S�CP�?(jV�r���c�y��?	?��?����}항�M�ɲ�(����|YB(�]^%%� �y�̡��0�[���<?��g����9�|��vq�XQBԁ%mB�����9��e��0x�ںHe�ʡ���` 3����t�Mbܘ+���<���au[h� ����&�)E͝���p��Ǽ^ﳡ��X��Ӵ�4k�`^;޶�1B����dzu�����R���YQ;����B�fv��W��0cS�t1�	��-�9�82%g�h�_�>	��0Q�3rV,Fa�GW�EZ�'���Zye���;9�������#6ϡ8�3����ݓ������)՗_m
���P.�*�����jJ��Xu�;��3��v�F��r�Ğ��΋ό� ��m~���v���st���r8�
%��Ѭ�<]�"6d}{<ĝ��vi�v4G0(D=���,s���w�c2V�ny�C�x��#�S��&��s�-���IE����- �p@�u+~�.��'��r��
heX�y�xoT���L9�~�=��[K�hk:s2bUfIb�ܦ�~�P�y�o<%\�+������e��UV:Ҏ��[�>��םT�Q1�c���Aʿɠ	�Kz�kI��1����L��W�ҙ���� ��EVm���P*d����2er��aYh��� cր��KA��	�}� X���!�]mt��5/җ���R��^6�I��j�;�x�ډԬ���?ٷc�Wy�J� q�t�jy1���l'*�qI=�����?��T�SA����!��(` A���%h`@�� �~����.����k9�
�3i���td'[�(����i[�$8����C/�?�G-
'Ã,�#Xk�\Le߾�c���o'��b!�`6$+�;f4����A��Y,�L�f	�F�P���9P8�*��w�D���$.�6��$Y}��2o�}胙%U�,�����g���I��7Z6��49u'�n�_hC�$V�FDZ�RW�,g-?��1%ҹdl��v�5s̳A�#�n����_n�P���J�:V?f������*h��_�`���D�Q�׈S��F����~J�]�9p ��!�\ycfQ(��r[����xU6Mk*l��K����d�5sE������9g�m���£��L��!����/#M�Y˔�&~V��A�69�Edc��L��C�W0���n�ְt�)�۹# V/_�N��ύ���LFS��`e�n�󞡗��'HS��h�S���~oRBa���fQm~	c+�N\��-����>��nP�K��;�wI��,����}%�Vy�I��W�O�[���(`St�v��2M�e$ �@XB�S���pq�N�7�z)0��������ƨ�~�A�m�mq�N��7�ȇ�Y݀ p �8<�{�l;�����j�/����7��?��SY2/�}�Y�(*8�������\�h������t�!��K��+>��38qЙv���Ѩw�s¹�U�� ��l �/�\�	�a~�/y�-ٞr'�M��O���3lx���@�m���*R,�O��ʰվ�o	��0߂�f�ε� �|��. n���F]uf�����Dߗ�\n�.�\����3U�92�;�'�cX���$�cG�s/Pi�3���+�;'�j���]tdN�_���"�5�∀<�����Z�L2
��$2�c���/���G��� q�]�/�}]_E��2uP��6(�/���bn�9�%E^?�+ϴ����c��-4f���R�����D���qfnW+����H�b�Y\-�:��?��@����<��c9�gF�����'��8$\�b����#ͼx99����Pi�R8�-��1�/�%��ҍ2�,���#l��A�(Oyw�l�G�v{��=ج����R�.B�T����
��iÕ��<��#
�oln�v�Q����@oZ��ۋO����]�&<+S��g�q�M`G K灘��%��F�vF1Y2���-��@Yُ\�m�%L��<1��K*��N,�vT( �VQ#B{�E�]�����ۚ���oj�)����n�%6+}4@�������m�����A	k�4t��z�a�+���/��S:�є%��b��ap ?�fS�lIcU�
:i�f�
�T�h����Cq��]4l��O'CA��5q2��_�/eljn�J�tR�q׀��^�;�_�KGΔK��w��k�➨D�N�WeS�J���$}�9��f3����Fo�ix�OK~Gy��a�^�	V�xA�K�s��x�U��W|ۚ�L����#��"�I��M^�|�-,�3�Uqlf/-C �J���!�@6o_�s+��@i�����������m��|Ȇ@:��,*/ֲ�?��%bsk��.t���zR�ȆC�:�P��(i8�\�f�	(��zN�b��)�hj,l�se�jR�aK�9�:U�g�,�\�����ơHhzJ
!Ӥ��'T&�gm���*��]�-8?];�4��A'I��F�b�x�֌������a�yE���
Z�Ř�~I q0��ðwl�P��-�� �T�)ö����aiw�z���?g����X�Q����}�E����@�X6D�wCz!nV����K�>���}�iVh�������_(�-s���T�2c
��i����h��8^T��
�ū����]>^ť�����۱�ƚ���՗��V�ox�8j����5�����De�rt�S�,���;N��5dV��$F
�%1t�X��R��i=��#T�[4�K�d�Ūj��I�5 �RшqzMaIya��"=Fe=���� �
���}7���}�n�)�U�/�2i	c6�4��߆f4��
/ßoMj���&�)?�L�����o�=��@#�4��_��&	'�A_��|����}���C����������g���	�Y_{f���KFV��������#���V��7�A	�gm����Bk?�>�oW�ȧ���U�g��9�|�A�[ì�����56sԴ�ʻs���"�ٻb��KU�lJ�����,�v�-�f��=�0�Ca����5� ���j�7����Чr:�Ї9�Weth��ޝ�����G��Wє���ۢ������ZX�3����t�a'w�����^ݟ�c�#�� �1�FC�P�7J0.�n0�M��>u�?�<?�Os[F���(y��Ȑ�%H������ ��[ �A/�͒�1DB���[��;��B� Lp0�@�m����9����C��m��<�fA��I�TJ�g�4O�ƨ��x��#XP|�^��V�ŢY妄
=�F��5��	�q�[}��@>�e��^���	�l��6E��Sޛ9���iRE�*��u��B�P�զ�b8��M.H`4�=~����%�XѮ%OQrKVv�/6��i���lO��(���$�~���|;��K�sꡍzEv
��0ӉǞ�/9ݣs��zU݌��Pߩ��y�0jA��*���$.[�sA��4B8-�d�bV��Y��,/vL�H�8����Ň6��&�C�/{��nE�/˛/k�����1Z���&�x`,gp;��7�� :��X�?��QN[� oL<���su��Q�&�hñ����:���֝^�|���SD����u�T$� ��_[��b!��ezi��f������_��y.�)Ҟ_]'�t�EQ���Ju�:�P-ϼn�ȱf�CL�6�	�x �0�;����¨�h�x�X!O͔]h/Ǹj�f��6`��ͨ��j�7�%y8og#i?�B�'���J���?k2x�W;�����n����~�:�+�g��y�[�h��/��h�s}���':2n����۞�1@zC���n|��y�<T��#_�ܖ����YH$�������Vz��o��#[&!-S�a+�b����pD O�sq�K"ƍ��R�Ԇ`��ϡK�[8i�I5�I��K)���[��{��$��V�F��&����Oq+e��Nm����}�"��by�
���0'�xP��MJ��r���J�F4��63ﰋ<����\ �c����[�'Gp���gp�4�j�x=^ѧ<?{ctS5͢r�e��=EŮ/����o�>*��|ǳkq��{�����@c"MaC\VyMk.����R�}��]%PʌS�}�kr���Ֆ�KG�q���������EN۷�H�r������PA]`�=[����v�~y�*�>+|��mk&�U��E7_5z��|Eċ���FA��!Vke!x��� [�*��3wrFb�|��ԉ��:C��L�pJ��#Q����� s����\�ͩ��}���'́.���(�@�3U�Km>��|/2�X�&�{CZ2�j+{��dʝ "}xc �O�6LDx1L�#D��?��u�$�e�'�
?�7���m�st��keNl�����ؓ!���I}͍������e�?qa
���L|�R<,�.3;R�v�Ҏ�5�ᤖ�C�Qf�Դ�c+������a�p����]��� ~�Eo%�Pb����ڳ0�p�[M9p3�~/���qq�q�M�x�/{�I@AW�s!����Ӽ�-�H��3�x{c����@[
t���b��M6�+¼"T��_9RDI��]���{֧�v�aۜ��JS�1xP��P��g�� ����>6�v�)̫�I�b��$.
����܋)�P[eH�7��Bz�e����v١�xw4x-�|7�Մ��k��N� �������LB���r��|�q�-�J��kj�a��w�e@��Fkz8��Tw��o�=�K:"�R}��`Z��qq��LSNl�S�$.F�we�-�~�ƍ3�_:v����>,�l㎙
�I
��dj>ĖvF!���T_��
o��9[���$�oCX:�+ǉҐ5攞%;�T5ZT�Z�l����7^��&�؁�D�c�V�.¡]rז<��}����p2���d�����+���u�	�kܢ��q��'=��Po���\��[����R�Hb�81��y~o���k���*���Kd9A��4�(�֧�6�#*R�׈���wɠ�He�h�b�\k�jõKXC�̮T����F�Q�Ĩ����S�������$���U�<Ҍ4F�X	�\��f��-*�qBhS":6���oS]�nS�&����oW��7�c,��jg�Y��_���� �U�i�O��o<ul�]:�g��Z�R1ef��̏n� �2&.>�n�
#Da���)m�����M��sV pn�]o�py���8A]>$��C�^�����\�閃��w�z�1V]��=��� �Ib3�)ֲ���g}���D�_<}�I��)����F� '7���oXB�DHDT�#�b�����Nh̑z�&�V��J��j�
 ��ؓ������ަ��xb���C5~�O�^��oh��e	O��K�+�ITtK_Ly��I;r�]�r�+B���m	�5�Fݘ�5��*2r۾������?�+�
���hr{���n����1�g/�2��߄&y�ݓ����Go�up*�q����8�gR�s�	��#(R���F����B�֥�*jR����qAR>��~V4v?��I�MP� ����r+�`t%m���g3�������O�׬�e����:�v�o!���G��y�G�]�G��<;����Lt�TT��~Nu���#K|��**MX��'��n#�&���F˧D��������HZ���f0ƍLU�-ػ���P�ԍ6rBb>���*��E�)6��L�i���mC��bS �h��q�#8s��ʠڔ+�ێ�!XS�"M��٪2s��U�oM�B��#z���w���h�{v_�)��J�p)%6��T?�Fb ���륀����f�w�;c<b���!=�J5���i�� ��E��t�V���Ʌ��b+�/v�u��v*��!*���R� ���KQ�C�t�l 3�sl+-v���W�j���t�}3�ƽSɥ����y�}�~T�YC�ъ˱�$����ļ;,&<�N�ހjJ�mFx�}��i|?K����"Xl�ر�ysS��E�(D�*��}=�o��k��1u2/
���N�jM�Ɔӭ�#ݟ����U7�$�5<Q�X.8�≯�P�j��m ��J�eb�%�K*`\FS�C���)#nE*!�t��(�+���Y �P#��G����@|3�Q�-Up�`��$}�9}t��|���B��7�@����C�9�Z�|[M�Vq���,���9��Ч�Y����q���ⵃ���ǃ�Z)RM�^q\9�#�P�Q��YF��K�խf6Wg�r��_%�$A��N���ðP���I5�8T���Ռ�(��\���ȵZ�ZB��7p�c��Ã��O�x�`�9��!�h틯�2�R!�BQPx �h�t�p��F�������px�n��Kc��#v[� �� >�1D�z�.�D�^j_�=e�:�"���!=���=!7��5��X���P����h�/�J/�U��ڑ8n��TI�Z5N�u�	�P����D�MPx�5�M߁��+��̞�t��N�t�|�~d|�F2W�}xTG�;|�Y.�F�ĸU�]�5)��av�>lB�z7mڼ�Л��n|�i�=�k"v"o��B籯��0��W[���qt$����xn��_�"���m�-Q��NhR�D;8X�����<�n'�r�Ģ��49OpHT�5���gm	�X�_=@��Y��u�4��<ב�z`f��"::�3?�onf�aЛ���c�!��j�e8�+n�XdV�ZN.׫e�x�Hu�YS�����S\6~����	P ������vg�zt��B��O�4?��q��:�˞�1�+�d���a���4z%�)y��'b������M�21�uqM���[�ڗ�l�_��ȭ ۹�h�*ɫ�s�/��W��A.���`��}C�DDe%g�)0��F�����@/<r4���:�c�)��<#_͚��u}�Ǝ�;!uV"z�!<��S+��e�K(ޑ�ʮ L�0c7����Y�[QA���q#P�g�D\���y���nR�$�
����s(�����\�Q���I����YÏ�����R�~(oq��J�7�e���D����T�)��7�ц���ӥa�\V�3��V&�9�K@�W�2��Mk��с�`L�C"%��#�G� ����\����S��wK�mu���tMy�_3[e�[�6�V��X�%|2_�-r�C�������qK�M�0�o�H2Y�X+��,�ѝ�������㒝��g����j��D���O����<������+��B3�W��*t�e�>���
�"n�>�>wr�����w�\#��H�*�����fO�u֏�?��i�Yޣ:5!�9�V��#
9E��T)y��D�Һx���/��}T���'�SȆ�ryAC ��USx��v<��~�`�@$���!sKtTG�`Cr/A�L�� ��rG�e�ՃJ��W�n2�d#�+���&��$;�����XJ��ys^J���پ�"UKTf!�#�JK�cy2�鹾$�]�[L��d�������-��ț�5pp�c��rm���$X�R�6�Y�8Y\ѦG���w<��̇�GB��ݒps�wGρQ�h��WLt�7�:9��vBU�_r�2� �ߦ�륢��"G���� �	[�7�o�
�Ybe�����?[�d�������DW�ة�h���mDW,ݘ�p���eYL.-5����lT��O��"7��'0ٕ��u��%aW������#!�OB�W*چP�y�3�2����&L�X�
��?_���۞ȵ&��J�]'E��ER+J�_@��dZ��,)x9��%uLc��_�Ѽ3E�
�a&X5��	�� �"8^��[�{�*"c�W���f>Hm�	ئ�J��o݄h��x���.4����;�l���88�R�:^���{�z����YҰ$c�t�����Gp�W}$;�\<��8�h�X�J� ����O]g*W�um)д��(ֶ�~c!�L0�+1��R�E�����~����W
���N�uJ����pi�6�B���k���;XG�{(�:U	^B%��b4וm�M0�������6qO�fL<%8qJ* �M� �\�j�yx�;&$�n)N\�	/=��qlF&�أ��3��R47K�5���Zߋ[}�Ș���Ԅ �����xc8��L2���0�ɭ��<��g�yQ{C��U���YK�6�L���}��:h.��)��j\�k3�dۋ&��j�|��袲+Z-��/����_]��)��A�C1l���������,Qд�5#-̏C�?]�u%ߤ�I5�� E9�.� NE�	�bkv�����k�Ȅj{�p����.�\/��V�k�+-6 24g��Ͼ��#;[v��� f��� <:>6�x�E����ʅ���c.��늁B<�����F�1���UmŔ��Fz3��o�ʏ�0R�]F�����>KB�e�z�pP�߆rq|I�m�#��|h[Z��HBr�����}>�i�2r\�nY�Fd���U�w�>bZu�'��a �#��G��0_�}��fX��{Y[?B�a~V�s��~�gu��=`��c2��5mޞ���G��em3Z�eL��7}��h�t|�(�%�܈��k6���
�_ߪ��8p��qz#����(��ղ6�3�@���6���5[���X|�Hr3z�0`���8���E��_��%����f1�HIw�-��7��I��?��"�5zC�:���R����ۻZ+j��j�.5��	�������(.)��5��>���3L�p�4 )u'�rL=S�c@I�TB�U�$��<}r|䕇�LH���'����=�α82�>){K�O��!���:��_�C�j�I�Ð�5�@υ���.-�Չwޞ�4�-Q;?���M&ь�AJ3(vh�%C�IH,tcC�)qn�@$�v+�#�J��W}]*��cJ\��s��W"��嘛Qo(��l�!���/l/^g�[�=����3o8���?A�������.�R��'��5��>�l��X���5��vm0�>��XjEf��=>���?w[U�r��U��sg�2�:�ι�^�'��f�s��f��_�cy�u�$Xt�6&S�>����C"j++�X|x4dR:?����#w
�[�(=���*(�.QR��E}A��8�	��!&���v��X;4ggy������=I��q� �X�L�W���gm��S�E���a�$C^�J�t�F.��e�?rӱMIA3���l>6���Έ��~������ϖj���ԙ��x�Q���񦠷OF��Ҟ^}7e����Yi���ߌB?\^�1O{4��ː�VX������\e�@�B��f��Q��ڗ�30��Ԕ|�4Ձ��o��X���/3u&W2��:f<J/ �d�fF�z�:F(ށ������g4��*}����y@'��ˣL0:�I�͠pSE:;?,�[�=�p:���v���A�޽^|��d����ۦ�]�̈DN���b��ܢz�2�D�k%�`�iMs�e�؃���L���!����9��'���9�F�^0V6Kp�.=Q�h>'�MS��S>�?�Y�0�XRk�[�K0���b'U�>{_'&[��>]��h��?�����?#�Xz3+C>#�e����U�_��]ے��A���6�Sz��M0�Q�xO���]ft��&�N4�������[���q���C�ګ��
��^�+��S�w��K�N�0��%��`f���8c�!c���v�y��-��E"��;W�؞�
J��[�u��5��\>��}	��l� N��ŧ�	��~$D�l��[qE�6�-U��Ġ�]kb��Lk���{*��і@:Ew�/���
ۛ���/{�,��MS�)=ֹ��v��ů�c"��x��+��v�48��H��P�AR���b@��{�R2��׺�P�1�����F�o�.��T��Ñ{�x��U�i�nwż�6�ç�ħj�� ��3���O�1�9���tg��		�("�b[ƭ�ɬ577Ѡ���HתJr����C�k:l�*�_R�!��h��l؁��8�}�������:O&3؂Y�sm!c�\@�mr�P�����n֠�3x���U�8���I�e�J����pCY�W���0�Z��}���9�)�	n�We����q�T1omK���݃��{i�q�c�&˺G�t���w�bm����Ԯ^t���%��e�i-_� +��%�h�Ҫ��칖"ci����V3��'�c,kr���.?�PUo�H�8!S�G(�<����o/�
l�.��i�Aq��m��Y����q�(Jq����+U� d��%�z�\�G�8"����M�˞k��Q;¨��u���m�nՠ���%�|x�K�رV�3゜���"�Rm 4�����d`��9}����G`�#�x�F�h�ԗ&B�k����B��c��e����VP^�-z6J����n6,���[�=���rtZ�%�K^��L~�\��J��!M�V�Sk�`�v+$����*mR&� ��c�Ɓ�v8f8=0z䘟b1)�������t9�/�sД�0�M}/mJ8�b��!D��}>�CfQ@�g��?yJ9��дNq�O^�uw,[������R$�P�: 󕥴@"�[���dفu��_Q�G!MU���[ɻF����՗i(ԕ~�kA�B�1��(UGQ��sA�)��2W��d�(����xwɬ�FƁ��_=�wH��]L����dȉ,w�y���H}H�j����)��t4춌4�ٶ�l��ܜU���VE�?�xA�tx����Q����R�4�ōV
�Z�4\{�6>��c�.��&S`�L�C�����b��J�x�lBDo���E�n�.�r���ը�/>��!M�>f��ߦu[^��F�w�I�Xպ�ʢ2��>��#o��5EUv��]}=C@�+�ֵ.�m$ao�����r��w�v[�G�����!nC!o,3<�ș]�,�dt� �	�E��:¥�e��<���6����V����w3/C۫h���:U7��,��с������/m!Y����xj��I�h'}�+�M�5e�O���>w�ݲ�@�/+�/���ZZ��|P0	 ����z�p;�OZ�3��m"�y<��ȢG����e��"�2�Z�vZU�(�,����J]-eM�,������	XϷ@E���~�lw��w�M�2�d�������C�4�W@�Lͅ+f79�j��Ԩ��y��)�+�6�֕�&<�<ZW�dCLek���`���p��/��E߸�ʀ7N����䓺�5��	)��ȃ>cԝ6�:��$��.��� B�V����ўg"��=�[���zH\
��A*�w�p.�w/�8EM��� �����0��ȃ�w�Z�|��-!SRNy'h�GԪ#Y��ݛ��㖌MZ}��L3$̇��$"����Q�t��yIO�T�I �t�x�� M��N!��z�\�9*:���|�5�.��H#=2���cqLm| �r�~4:�����b���0��ڡG�"��D�9��ЊBR�~�ڍ`����@��|@V�e��t6]<�K�_���?5[��HO���-��{�]�Jy�9v]u8&�<�P��ӴT��j���B+bAq�d������&��28W�mF�)���i�w�,$�)(I3����f��&�[�}�p<�s.���EGȤD?�j��%����#�F�՛���OZ������)�;�w;r�M$(�>�\K��aJ15X78-0e�$��2�q`N�X�=���x��\��T��SZ�5��Ne�OSܠ�C��H�LΌy5W>-�i�7ۆ�p���vЕ5ԇ<Z���;�YmR%��.���� ���"�x�=d�o�	�@M������Q�*I�U^U�IE_Ϸ�.&Ҭ
.�M)w��[_��2]U;��o�6ލ����E�XV.ԏ�G�o�ߪ�]C��g+ԏ1�W0���!$Ƿ�@�ۄ�XB�{MK�"��`����g�og��!�q�vD�&ZY�ei����R;�w�v<�DA"]�.�^f!�=����g����U��?Y��[[��A�����������7�馠I�j���%t#�~N2��":��f\^�Uխ�Q�m�8�z'Q�U��Smrr����R�ˢ��I'�]H�@�5�F� 7w�;"�8�?\��?9��u�:F�'zFó�����.��V���)�AP���d���
_��CUo��̱��$Hj�[�؂����`�'ړ,7]����K��ț���=���W-r(R��p����1Ҡh�2����^+�?���>+Q�f�:�KMbiw������Zz~�dɴ��}>�x�S)${(4[�ݤ�XXN�^*u��W���p/��SD���~�!r��v���V�^<��D�� �a��uA��l���*d=�`��䐦S�奲���T�Ƈ�҇�W�䜅�\�4�P�d�l-���gn�6<,U�;�q 8����)w�*o�H�M園�uX����~G�f�+�mdJe�oL��Y�����q��O�p����Aѹ���T]���<����4N�Қ�[*R��B�j�7�2Tҋjq�����	��c�Ҋ���T%k=�q4�H��	���Twtd�;����!��� ��V߀Z��_�Z1[Q��A����>h�L�I�;�r4�o��	�Dܑ%�!�� ̬-��Ќ��l�0�~bw��< �l~d����L�x�k���ɅNA��Cp��Ա�	���X1/<�UT,�!�%/���֑�L+"v����Fi���\��=��Uiņ�e��H
;ۥ?��dQդ��Q��x9 [x�� =��wL���L�B�"�S�0`���ȴ��.t��Me�/xr�)Ӗo�sy��_�b2�o�O���G�H�������������uyD
f��w6��G[S�P�2��i�����n����H��~�(�l
3�q��I-��Ѻ�{
'm<aTTֹT���vh_5�M���%)֚�_�Duj��U���q��@��	���]9u�n��x���}�'~X�TpV}�=+�/օÖ0�ԇ��������V��À��j\�*�b�Z����rV�w����uZh�����iܗ�$�&�b3�_d�����\���]�`h�9a�c-�]���t��V��G��2"�^�5�+��?�5#���֖R宠���wZa��Z|�Q��������P�'!����~`��Zn��}AC:�s,�����K��С��u@ �e;Hۊ�<$�0~�>y!>�7l �A�]�ʊ�!�$\�Y���SB�W�(G?�j0e/�Q1���xX+Hlaz�O�ì/���4�C���I�+k������w��Dv*P=�ƵA_�D@ci�W��orV�7�M���8�}�D������ڴ�|�UN�}�����,_����/|��#��Y���(y��9�g��.o�Ih^	#�\�e:�;��.�E�J�/���̹������4Ԍ��b)�y!'v2�dQ�̕��WH��fE?���b|�ߠw&Y�Z�搬Nh|�0��H�3��=2Լw9�gu[�f�5��h�`���kz��1(�tw����B�X.�F�~�@D��%x�L�zS��#�M�ǧ�C���L���(E��!*��e�8�`�?t�Α���V$�_5��1�"ޱ�Њkߵ_��G���ɮOK���3��e�����jY�G����dP�T-t�خ,�&����YF�P�hl�~�"�� �i`�	u&�i=۰�ǕT7��$� RI_��ߪ����׽�1��9"%�PCF�ck������i�瞂 Xf�0�<�l<<�ҩ�54�͈$���%W,������O"ύ�o��=k*9A���&��*EawmѠ5.Rvי6��gg53v�
��<���e�M�QiiLhM����-lf���F���� k/���J�j��:$�N�V����,��N� ���OH5�O����?F�"9
�&"��;�J���]w��#�.��T�,��
��.IW��'g��e�_�_�iӰ�>B�^��֏�1�@�mtޫխRe�/ ��\��ЂY#�f�����L	��vf�RL@ˍc -���?�W8�;8�@�|6��TʹW6��h!v�L`=b����po^�y�<�M�><�n��K�bǲ5˻-��D��^Py����m��@��� y�i��t�`��v��H��	�w�ˉ��������-t|�v����<*��Գ|߬�6�2ҝ�KV��S���%Z��|]dAj3�K��*L�鱹`���&l�C�^�!�Y�_��c[�Ԉ�rjgٻ�}��M�#���&�z�0S�^���ޝ"�<���>����`L��eÖǇ�x��>*,�3Ip��O�����XO����mc/���(��{��)K}�=T�rA+�õk~CW"q|��'Q؋н��������=��d��e�a�#If׭��Q`P�GmbaP6Z�#.R<=�%���l�Gv�g�9�@*�W;M!ܣ䄵amrk���?:�>jE������3�����Ӌ�g�
@}Nq�cLc>38`����p����#B��Tek2+j{~'���8��˶�f�Vw����y]w�]]v4&$��E��DʊR�;�=l`�s���եhA�J�T�XD��M�.�
��s�I��h���A��+�$���<m�k������� >u}�{��!��?�
�ڥ��k��5LǛ8�g��Ù�~e���@P���e�fK�9 �X���V�yx0�=.���f���x���^�B��l<���Ř��Rbar>DO~#R)}��P�<�b�ý�rb��=zZ)9U?6�@����w|�u��N=��rY�rcIӳZ $"�/i�yW��G��k��D%5V�[�Z�r%,\�z2�Pڿ�njz�ݏ���;yU�U��M��X��nF�P�Biv�h	lzSI�^$��
�� �Z�E�������y���ܑ��<�.BCƯ�ǯ^��i�Z��6�<�c7���"��Ԗ�颳���a���|m�y�������+}·�Vu �� �(�	�oK�4�jz�q;�O[dج1���i�bO�g.�mGcj�M��Yg��KF�0M	.��T'Ǡ���a�{�K4C��9�	���ޥ�O�"�����Ly��?��7${��(�~hs{`㚤����n��,,�hM��]���>UE|�>%I�i�{b��`jJcLh��i�w���)3�}�3��r���OI-�|��`L`	��"˃T���L�z�r�p�+ 7i(��&҇-�̞��j���a���T�����q�&!ظ��	oj�]��؎J� ��%D���H�eȮ�x.+$0���7a�XO�X6��#�KX�(B��{䝍�T	��c�q4�M��cLp�9˾V.F ZX���b]#�,}C��oc�w�V&�
�d�1?��Vow��գ��u��a�B$�l��T��P�M�q���D�"n��;0T��O{�M|����Z�������Gv�8Xe�3������G�isEc!^������I�B�����ֆY���tU:-�$'L=n������g�s��b��T�(g��Lt���Z��l��H��gc�6��i_ޑ�͸F��/�gJp�wN�@�n2]y�q��!}�\�h��"�[���.~c��0I/�A�ˆIDc���~���ｲ�.��d�^_J�x�&Յ���p���Ќ�{E���*e�yP���}��fe+����38}Q�ib��t2���Ee�d�.lL7�B��+����Α���H�M���[��n�
�!�s��U@�Gog�.֏_#ϕ�TS �'c� @�c}w;�A��{�m�T�kMB���up��4�}*�p�����3i��k7^'�,a��&2Y�K�P�1 �J��K}�G��Ε��d�����pX#x^!X��OH�������m�����Qnr��n�lVQ�,XJ 	�@	/?�rѰ��:��:�
])3x��
0邆��?�NNG �dH�8aǷ�(���m����+I4��r��0 ��2��F��ԯ����L�֏ɑ��}����Ύ�����{�'B���Z>��� ���ǳf��k�qQ��.���jR������*q��՝�Ou�8kToK��]��<���G�1��C�Dr�+89��V�>751��J��H$�D^]y���w:jK��P�<�ᘼ�����6�}2LJ����~{2BV7�8�k;'����s�UN����Q̝X�,�+|�Vp��${{�ȯ�d��-����z��In�c�����g��4��,�q�r3��6k�q:P�����-��?�6�e�\%o*�1Λj�&~����Q75x�����g�Z�,~�v7���P�ղ��3���Ɓ��Uqn�DD/;8�tZv����#xq���v��|�ѣ=�_;э��T���x�zo*���GL]ԥ�Y8������1���Þ�X��;y�v��%�ˊE�5�6<�Nom^�W�KZ2:S0�yϺ��sI�K�H8,���#���!� �6 �yi�u���i�ip�>ë�������Dh
��I������5��h9P��D��!s�mN\�F�1S�i<(G��[�=�)8s���S��,��90��|��؟l�d�z���L�ި4$�-���Tɉ�s�j���ٞ�h}DD�k���-,��)��?B O~/�kנ��'��}��
E�^kU�o5�a�~�W�vh����5r�����7�����gi�D`��j�ŃhwsxK�L��z���Hς���e�r(C&�ú|�s$�r��'qXb�m�����,`��cp���.Ϊ'��ZT�O�W֧��<���m�����a�r8�%-�����tΐE����i$���_fL;����F��Բ�}���3|���_��{g�i�X:;�i��`uNOS��R��>��1�a�˙��ֻ$N�9+�Okv`)ʭ�Haʱw��w����(�B�4
��	��B���y�.�*�@�i19�S�������ʋꆿV��>i6��]-#w�3���枍SSzց,����QkL^�-&��L��p�@$��:�[�P1jER)Wzߺʪ�[�kuy)R�Ɣ5�r���\����=9��5Y���abI�R�����Ѩ]i\�>p��5�G�:�8�>�W�h~KH�M�2:0��ރ��.2V��
�5�ԹՇ��9��3M1�*V�����+�'m��t5ff����@�$�Ź�|���) Y�����y�F ��M�F��nD���3�#�����R�{�yݔoXB9^/���D)~�6w�޴o\�*<��B9�(9�/_��s��#���0/���h��8�	�\|���A��g|!����X�o�ɩ�H����1�-*�L�5�PQ������6)����Ldd�=��͞.8p���~Cz)�3zW�c^>� �����\iy]s���!+\K���Ғ�2fX�8g�����~Pw!Mʸpht�Gm�1ϴר;C�������T)̆tm�����;�E2/��8sO�m���9��;#N������jO�b�3�l��{��#�P�$O���X�,!4� w���5ԡ!���vhg�*w�+n_?m���G9l�/d��-Y=j�N*t��Y��;�s|� Mp������t`o��|�ybH�_����ۃ�$��2G�#E!q�r�#�(��ɟ�����E�9�T�[�M���3�#�9�t�bЍ�o#�����ӫ��n��H��rkC����%�$��I'�U��!�6�`�C��[�m�<�4�zO�MS|�l�Z^4�.#礃;)��l͸`��Z$�P�D�z�f۾H@xs��tԖ]>Z�~/ĒJ�5�~���E�H���W�ڲ̜KM�;Yq�C��ލ����k�Nowʙ7"�ƊP��Caޚyk���{>���8q���1�C�;����@L�q��X�;�r8�o�R)�=��A��H�a��M�Gw��=y�`ܐ\,�1B�/a�%���XС\���_�4d����2�L�~�<ȭv2�,���TY�d�����[&���t�f��1Zh���r�UI����s�R��g��=�i�L�s�l	�S���Em���Q�n"@d�7�ƶc���%B��h��� X:l����(���pZ�t1I�Ҋ6�Cj�1)�`n�'۱^��^� Uj�é��\P=RX7�m�8,t�[��:��z��K*���l�'-��hů��㻷 �"De��T.c�=} =�DTg3��0���?��{=.4xr�K������-�Wv�>���!�>�UZm�`�q�� �7BJ��N�B���_tB�8��(�<���d���_��?�
�����9��I��RO�Ҁ$�ɴ9  �s;ב��̢��O+�1�_��L���:4�_�<��n?J�{�4������IQ��u� �8N�2��̻�]�z+�bI�NQ�������r�%C �G�!Z:?�8���ZIOxx�t4����7���X`Uڛ�0��W[�/ki�n�������#�hɋ�a�X��;����s��0K�Hܸ���4B��F+��1�`����d�D{^�b�q?��@����t>Q����d����")�]u��¥x�����Dkcs�������g������/>�~6�oW���ؔ��=Mjo���Վ(��=+K��L���P��}/ȁ�>ޒ��%ѪQ�۩dZ��A���`C�����K�L��&P�#5!��#�ԸF��4I.m��f�.���{�&W��=$eث���2}�x�Kf8%��}�Ĳ��� �O��������L�cC&�[�Ʈ��h��zQ����qe\Ͻ+�����ƻ�tn*�B|r>W��j����ZΪ�U�B��Zj�9YsN�@������ز4�w����l� p�'��;���]�o�' �=/��=D�i{��D��)�7�,t\���P5�z�M��?�.1<7��wNF!�P�������A��ä:��%�"��-���ɻ�}\���~@[QCߠR@3;o�M����4J�:�k���#��+*���� Z̒�s������T�gѬ�R���s�8U���YͰ�?��b�?R�|̸@N*�qڼ(��y����)(��K����m��UZ?���lw����"���v�+�"��0W�3�5�a �5#��Ҝ��2��������Cjc_WT;�Q>�Aҡ_�M����Hi�G�Wo4�_J@� ����l ��8�_�Y�Ł@q_��3� (���H̚�v���!L}�?�ezUY�1JXz^\Ն�ﵟ���FAv��v��US����
+��Q���+3��U����n���܉�%8��++eA�ۋ|H�@��և%ɹ{�؃�%�C# _|�� ����D:2�t��KyMMW}���I�>�mȍd�F�5�������^�>��Hl��u;�KDU���:���<�xIva���D KC��u*��\՘��,�BSS�����,v E�LBr�VR�f\����M"�vBT��;��Ĕ/�G�9in�����9N�ٟ�g� Kj7l+���^U�kAjz6���I���W���i��7,��w=Kb<��	�K!�T�]#���N��� >Y�X��"+�A=_Ο��� �u�q/���l:=$X����|]`�|���c8��m�r�m1��e�3ϫPY-��ZK��W�
��Ư<�(D� � S�WORd��iD��eإ/)�U�Q�i�(�xc������N�vĥ���3F�_F������vb���
��$��x��*s�ޯ����$qU$��){n^��`��V?�5�0��Ք��X�gP<K�jʉ_x�Tߪ� >1&�TB����=G��5!׺��DW��j�����Ƞe|'�Jg8�>�\���u@��N���-tA��q�[�4�;�a��rmE���1����`!i�bF�w��fئ�V3Ǖl�j��ޢ�}�+�	}<��Sj��<���s�j�kɦƟ��n��O�}l��$�E��;N�q�$�k���r�`�0!/�X~�`i�}>"0v1�m&?��ŊzIN������[�����Ni��Br�/ ՚�HO �$_�+z�1=Jp�C�y���\�~�)B'?�u�r�����%%���!�ʊZ��32����Հ�U��I���*�@|v�1�ed����;����jO��@�	<��@���"�&ܓ��sw/)s�ɉ#�ŵ�ל|X�(r0��Š����K�Qz:�H����,&2��E!�O�p"L�7�V4�ꢱmh�˫-v)k9me�J���C����
����\���:�X�W\NMa�������A�A#v��j{�(�1�� ̆C��L�(������y�����)7��
%�H$�OQ(x'��i�a̼����UFbU�S���֟m���覯�w @�q��+�wY���Fn	�l2D���/���{��~��S����W��A��>�+�9�i�9���������7�_۶��>��Nb+�-2!�����Z@�~��~D���S(4���Q�`��Q_}�k(��{`*���x�n����o?�}�����oP�B�0��~2���3�f��ʐ�����i�x�e���*X�B��[0.����Ź|C�K��w�伃piI��������"��Q�_�v�o
��c�E��O%�����1�,k�VFw\��dK�Aڕ�
(ܑ��N��=�� ��7�uY�y_-�6������k��=���xk*L-&�wq�-6U�h������V�~ό;�7R�(~|Z��"x��z<����Ïu�2�&�Sck#j0��E���\�^O���1D�f�/�gVi�P��=�oJ*��!z���7�7[�Z����=	�*H߅:�_Ƿ�ş�2)wp^)s�܏�i
�a�^v����1"�~i�p�p�GIS8�O��)�'�m;�2���1�)@�2	Ѣx��F�?�P_o�����>��dZ�m����4TƤŚ�>�_x��~T�X]�;��ߨ�R`w]�l��9�ஂ��7�ղZ�u�̀�d�|>R��������8�%t��g8��a��^?�Y�Hʠ�J��1K����w�i�k	��nd�����WʜV&��}�m�;�Q-U'�4�ko�&��W4٢*Gu �}Qy��E��$���b��uGs�=m�ͫ��|�z�NU���+SW��<6Q�j��ۻF�~d��=� �p�	�"F���]f�ژ�s� ����"�QLu�c]�b�Q��J�(ޥ;���������?�۰|��fį�n�c����Hgr��+J�3�����| \Hmq���R����8����6C��ݦ#6��������-�z>	ݘ.�qnďbi�l�ͺ0A�V��3n���q�ө����Ȩ���k|Y��|i�KA���b�( �L��Xq+{�������3;xِ�:��il2\ P��K�k�F�����`�6�%��dR��ös�O���/!^)���ݜ�R��4G����������55f�����t�[[ �pS�we6�YJ����/���J_F\�+������Ӽ�V-�&����ʱ;���A��uHȘ8F�X_�G@?���(�r[�8�/��g�a��%_��9ӽv��m��Z��D�g�I�|��w�'�eC�@���_�rVQ�|)ts� ��4���$�Jo�{ܙ��?xh��s�D;nA�����u@�IY+��������#y^
����;�#���N�eYh�[����IM)s`�u���'��C ���6�j�Y���&^F^���a,����r��Ý�s�����@���.]�5���W�{=z��')�>)��.�\i����f���h�H�w�+�,���s� �{0�봤s*]F��*l�\����T��
�3X�a��O�r�@��✈���G��*!�M�ͤ�pv&�{�=�c �0a����J�YB�Q�c�G1��45~��sx����`��鯩�Y�A�j��.}Xؾ\��$l�;z�t�ߊ���*�mx����,��i��#
�~l'U�Ͽ���PE��P/~��G�ν&���)�KQ��a�^��J��0����mT���q����\���"��0(��R&H��U����(|[�f���Yu�p޽�D����:!6y��E�^K��p�W�}Ffd'g���ڟ�$#��
��Y��A�:���[T�����v?WїI�_��̘(����.��ZY~���)�a��u�L1f]-b��:}�ݾ䤝���:]��L��t�%������W��)��JLA.�ښ>5�V�_@���G�y�^aD���&��T���-���j$��a{�~}�K{��w#�M�0Y�6��\FZ}Z&G���E�E���S:%��~�FB��8�L��\�������''˦?��;�����k�;޿��S��̞2פ���L���w����y-ӿ9Ys������}b$L��2��7�WH��GPz����A�(P�-ɮo�����ط�(j���>v��Nv,�l&�>9>�P�dB�1��Y!�0�E�����Wa���+
�1�'sRI�ьA�kKycY����|R�U�[���<���!�]a��h1U���Э�?���>g��r�2�(I��b���{X8���ȥ�N��r�}SiQ�����p[��7:��H����_�����!�&���4���Bz~5���6\one~�$�fkpǭ�2L��8[�@7���f�ZDU���>�� �뭧��A>�Aj�]U��xkh�r��+���Sq�����㗎���m�Ⱥ�y�*��?���m[Za B,�~���r�g�ەuHBA�+����Q��ؤ��������v|˙�X���:>��9r��Rj�Ju�+ȠR�aY]#x��o�}+;�N�)ܛ�k|:^U]c�Q��С��9���ֺR�G:��3.�K��%ӆ;���~��9N
�/,���T~��&[C�j�6���u�MT�u�No���u@=�Ocŝ�y��U{�W�3���|�QjY���ȡ�H%��f�fLH}�ȣ���pg�d��p:�esd��5r�#�O�c�D���~�(�v��V�L����8PN�J���A�YM�9o�+5XQpk}�vK3�;�O�4���Ϧ��t'cMg�(��;��������YK��amKz�	ǡ�����r.���$/t����J�l&V��6R�ܦc�����$�]�u��[�{��~����k�C����"�'�)�Ѹ��U�3z�˝�8��B*$S��pJ����N��2)��Ll�^�;�`��"O4��皬 ���p���.Z��ec�*��ʦ�y���i���}9��4�#z��]j��0�9�LeF2uu���wP�GO��l%����9�KO#��]ɛ��!˟���b���U�q2���Ү�h�$���z�s�be��ظ�"�Z�w��ђˈT������ս{?��i�)3i/������l����1f��$9upx=t��ݶN����qc)�Fm��TY�F� �Y,}�(���3
Gp���yʤ�8��.�Bh �I�m^�ֿ{�����Ǌ_�����뭿�=���t�T����e�ڲ��s椏�H@�N i�	p:�4yKQ��Z�a���z_3�̶�,+,��]��w+��G��PƑ@�3�&�ǞG̒1���!��2��_[�(}�9�7�z?Xl�,~{G���
�{<s����e�t�^ƿL�,(�v'���ktX�TeH�}�a��^熋h��s$b�^͛�������5��(T�0X����_��I����;M|ݴ��q�r-U�;�D.�� l~�Z������:��m�H���(�hy�o�M$�����:����w�0-
�`�A��ch�#)��d�������m<�H��=�)�7���ʥNR�~IvaTOA������2+��g�ٿ�c�*�ݵ�ʶ4��GzT��$D*JY!i]��
���
/#��M>�>5�0t�l��ɛ�x����52�=� �H*��M��ۑiN, �`T�x�'B�^	���V^!x�r#�)mϤ�H6&�v�Cti+�N<�=�I�\��"�7���ϲ�{�2�F��+�kK���4`{�(����Ȫ�{�Y!k�t���E��h!�`�(.I�!����YArǰ�@ܘh�o�__5�3]��U���UKY�(�^uƬ'�2l�=F��.e�΋!��hT�f�M���JC��UԮ�*I���q��;n=�W�H�
�����J9�k<�Z��Y���ˑP3H?�]A;r��J���h���\ i���!ȌUEk ����iP�8��%�	�0�ᄇ���.��l��u�{b��6�����CR:�ݠ��,�/�$�eu�Y<~�U=3�)�5CסuADn�;O�	���H�V( �hY�K��Ca�����:�)��l~���#���s�`��)�K�D�-މ1��+�b!H��z�f1���嗱2��rӿf��S\�݇����٧�ex@"�8����\���X��(I���0s|���[��|:"LS��Lz�}�&d"�v���,]�������~�~����n�W��ŧ({������GhQ�S����̽�������	��ʲ��|~���e���dh+�|���d�Q2x��.��n��1�@^&�`aS�=��	jK�ք?�<��U#���.R1�x~m�`�=� +h�7ب3fr���B÷r�����O5ͼq��j ��TL��s7��AZ�~�c��3�&�VZ�ř{G;��U{r���s�����b���Ƒѱ� �H"�mff�K�����Vd�?�����1$���S�
��a�"/�y�vG�'\^��[�%v�T���b������O�%%"����Q��f��k�ξ���_ְ������?83FңO̘���g��3��#L\3�\i�s�̗t�_\1`�s⚟̷7gQN�-��=��>���M�[��/3�ز���)8
�"̪mo�8"`�ٛqH�z���T����M�)�VƩ�a�X/�����} q4Q�!X&�ײ�8�/����tKH;^,
������`�:tq��{,?j�:�����w������Z��4Z!��P�����6���d�߃	5]����}�_I$�k��al�3���N4�6��_�����&��Z���⁾�v��0��T�w��W���C��T��ˉ"\�T�fC��\��fv
J�?0�&<��J='�� .� ����<G</�g�
|��w�6&y-�t����*L�X�B�a�E���/N�f��.O�ek����ފ���?z/lڵ,\�7HH�^��zJ�hJ!��	Lv��i)YgBy�MN���j�3��rtp׏��gt��c �s�xE
�������K�WÔ��� ҷ� �"���_$���y��`��yn6���s�|CQ!����kX5Y�!�~s���,T��+=���k^�����K��c�3�fD]%x]Ӊ�̫C0!�����c����u���1>
]�˺�k(6]k�S�W� �,4��B��1p���R|�}*T��a��O@E�O��ܰv�3v�n�3ޯ�0D��כ�,���;��,7�6o���d�~|�8My��D���=޽���#T۞dC�)B^>�ǼM-*x�;"������?��޳�ו=��]n�@~��gA����@.��
=�~� ��N ?)����ҍs�Md�޺$�����%��2����u���k���@���-ꫳW`�J�}M�����G�}�a�
邍�u�����K��hA}�8�l����/@�m�����4�vumv�Mr^q�������=R
M����î��֛��Hh%��v�0��ѐ����?��U1#�}M�EAr5�|����!��턌[��X��"c����6����J~%�g�ò��[�X�o Si���P>Ya
$�1��W��/3��e ����p;-bd�_��J��#O��$A�޴)�ԯ���WhJ<1KTzDݽ�haYd��߼b�q6##S�ֳ��\oD��ȏ�=ίo*A��X"c�m���h'�D����$qn5����nQ��d]���d"rO������kI�1�o����9�>�����uUt*z�UΪ;Nȧ�nd�{%XP	w��n�G|��,�MF���b���O,�`R���<���}�g�� ���[�V�Z��9q�<8I���*,� �$LO�zZ�D��K�1xj�s-��<��^I>#�!g�t��{ �&ŭ>�(�I��Ms�d��Z�)���<�Iq�֩��W�{l�z�3�hL�ʩ��-���9�v3�'�3���v�>P�(ˈY#���Z��a�i�z��3C�V��
|4���(,@�	�-&�Z,6���g�o^t|B����
t��~Z>RC5�-p���q猛��� ?���/�'t����
_��r�k�8܍�.���o�F��h	;�6��_�vF�ր"?x�mo�%�!r���v�,��������b|@�6�}L"�2.#����Y���u�_�����Z�S^*T��q A��d�"+nS~�o��T ��f�{^F����ړ��A��CpC66�v���s��e۸_2�D0�:���s�ETw�1�-b	��tX���#U�8�%�y�=���$������Kq���� @�<!_��%�����^eO�K>��[�$�����X��S�}�-g����! QQy]��є��0�0aݡ`���aN�U<n]� �)���9���7.�&'�v���!�CØk_�h �z��t�k�Y�x~A��HG�=0}�\=4��V�p��ؑ��_@>�~V�ʶy�<4����z"A��ߥ��R@n����?&�������@�RD�7��9nJ�`��h3����2����Z�wif�?�'�v�[xhg-�T��q�>���T���/g�|`����4��U���LȂ/�Ea+J�G������ǀ^�F��<`rq��Ē�D�X�����;o��v�Iu�'�^�1�M)��� �c�gCR�lR*�F��P#/���1��<�U��Z�]Wvf��D�aM�j�n�@ �5�Xy�$^���&Pူt^�Xq��ӂ;뭤�>=�ͮ!_砀��^�P��;����h��e�+�0p�t�w�M����l)"�Ica��}� �ڐ�]ɤU��v/*���|������@�/�
�b�e&HV	'Qo��FK�w-���M��HvJ^�ӌ��3A����,��ZF����hӽ�>�\���rq~߇�5)�X��Ҩ5���a�=^���k[�&�e�Î-n~��D�ц��EY��^�ʧ"'A��
r�t�\d���.���s���ȟ�"maX�;�[��Z���/f_P{�u\卦DzB2��.%P�|ҫ�2Z=�C�e z�|cw��m{��sR��)l��؈b��/�<K&X���+hH���A������!]�j]���1����;�n�;�Vqk���Ց�����G!�ŵL7��$�\H���m����}��ꕬ<?d&w�e�OG��*����=L3��X�W�UlڟO���oA�(��^#2B��M�[� %B�J���a#�]�=���y}������Z#��������+��l�*�g���5dş{��.����Z���:@���Cݕ:H�;w��v���^\���.__i�F�IS�j�ͱ�%\k^WNr귤'�av�AEk{�Y���x��3����j�0�g���b�~�����6�n��]2)}c.W��؏����*��s�za�eQ6L�z5�J#��B���4�"��oʹ��[���T��O��p��}��s��2Ni*9��jc`��#��Nq�J�֔p��2����JA��H���CP:w[�q-e�M�s�Ԓ(T�{�$P�W�c�>����S�>u���d��#�t���z���<3ⴆ
�{q��h�ϊ��0Cu��G,X�o$���[�o�5�S��#�|ԯZ~��Y�X�;�������.D�B'���z��s��SG�����N�`�d}�:[�{e߾g��)��Ds���5�D��wп���*��aP�dV$O��Ւ8Q���40a�˼����� rk'#�Z�<�b5�*�<uJ���ђ�����9�����X�礋�b���@�-"�N���d�0:�\?�ʋb��>`&F���X����N_B%U��3�*�!�h�g�l�Q|0M�I�*�<���aki�t��[Q5�� ������T"�%�uz��w���G#uw���
���N���p�Y�4����a�����%[`ȶ�g�n�|K��7�}dKRΨiNF� m߬�T]��?���5Yf�B�#�&D6�0%����s*in9��x.��,����Θ�X[�Y��,Q��)ɤx���*T3�C/�֋�*��C�ͩ!�ްǯ�a�d{3I��x�}�bu�[�/���HI�p����w��FrJ�B��?L�JT(����>E�-�^i���Gꂚ)��ة���7&Eڥ�4��V��N\q�W�ޘ�,O���Gb	�z�e5�q�$����V=�s��g���dHR���v�3�L���e��]Yx;��ay�����b����+@	=��R*�����;����X��\6�B���� ��3�jw�)ƪ�ք�v��A^�Fk�$� y�0��_cNgw9Y��
���hâ����.���gY$r4���S��Z0iu�~/3�
�5��e0O�9�ɤO�9TU�(�Ԯ�I�ˆ�d���l�F��v�R�#d��3j����=tj�����(��|���yn���1ǖ���A�7�����o�ܯ�X��Q�L&�hcv�x!ZIJ�.H Bhid]�-�#U~لYn�������@`m�vZ�+S	�1o�SQYVRz�G�c��]�����1���#iD֑�yw��xW�c�m֮��0�I�&7�!���yGu�JJ^0fa�&&	eHO�����&�<�r����nz8��\i�g�O��%M�bq�Po�J���X���]������p�swd�4kHB7�	����h���tP���qۅ�ם��>��sY(�Ӝ������i,�-~)�C_%�F�|�I���,Z�"�ȿ<#/n�x�jN�C#�{�x��A�/ޠ��ZB"�+�������_[#��nNNm�:����
Z�Z+�߯�a~���aB�����'\(��f�]�5;�6^O��&rQ&�����l(6(��z��k�}]H'������:�0���-|���F�X�m�?^�����[.�V�8H63�'�膋����RA���<>���}a�g�lfAv"�9��N���/z]U�v+#+�ƽ4Ql�Kę��2 �U� ���.f�yu.v`�tp��j|�i��H$�'%�̩����pY�e����.7hF���j%��ݚn��I�V6�ר官f�",�a��:wդ�p�q�	��Xf�v����6?��Q��_?�k�l^��G��;wV�A��X*E�C��Oq��td僌���fE%@�j
g��$��O��pY���sv�5x��hֽb���OzIo�嚀�� �4�A�������	�����.����(�k�&}��j�i����g{I����C�믃����|Ȳ�����5y��쩧�a\��k|~�r,!��3�:�&gל~Ӝ's}�B�z7-BV��2�J�=���4��n���.O���m�W��]k�+�uZF���L�gQ�P$|Cɡ\1�*�C�Ǜv�Ǵd�\D���)�7�ԤJJ���!sŇG��s10�å؈C�yk9S!��}�8-*�5����Oꃾ ��SK�XJ�P#�R[ٶ���RQS�cW�,_�$3�i��lU񳒓�,2��-EЏ����/C���!����Ń�&I��Zҏ��;�iI���m/����u���؝��G�	p���z�t��~7���Y����(s�쪥ܿ��t�Q+����6W�[��C�Lk;�&�u�`�[��m�'&r|c:�M奨�J��ָU1��y�}5�sԸ���٩e"T]�ŝ���}h��T[�����S�~+��an95:�1��U��a�k����W10���軬���Vx4S�"Q��<7����j$��o�)0m���ޙ���3ݑqQ���g@h2����Ze��A:x������)g�ԓV�9׆��<����▽�ע���|�0�jm��pY�w������KS8M�K�w�%-B�Xni*&T��M�Jv	��Ay6�Jw}6�m���NWb6F �!	S�A~%�F�<��t��?�v$�I_��(c>?
h@��{$%Ä���<���*�+���/�|$�Mkc0jS� �a�������T�jz����7S^�3�d�)��0B���醙� �P��#�g�I&�ϲ��?c(suF��Aq�Qa	�fҦ/�����bR��|R�{��Ë�"��
��"Q~�+�ө�#�����#?�/a��4�ݚ�O�m�I��/=���$� �4`gU��%^�����[|��'3��` �����ʦL!�$���Ĭ�26�_�O�C��B|��o �rL�J>�}w|@s'P�,s����?(~x����"��`�$��z�"F",̦���NX5� �V�v[Թ��t���S��l��JW�Ȕ'*�&�4�ו�>xv]���
e�=��.��w�ՊX��t�[C^�t*[9O�h��t�
"����)�Ǡp�� ��+m7�����V��In���[W�f��>X�h1��5�*��e��C�dÜ��2�MuRH��˳.�۹�QʹN��MŨ|�����|W�a�/bYq=;�7�yhw���9���c���Kc�c$Eɏh^o~1q��9	�؉��k]�&�j�5�V��*�;o�EN����1�/���\'���pq������|�Nx���#�Cέ�۽��Ɂ�/h��F6\q��㐏�Wt�hG;'ε�Y���B�
HP o�������9�Sxh��6��1�l�h;%\�(���lf�$�eƩc�}�h��m�p�[*vɦ���פ�J%�8�4�o9�gf��"O�&��N2o#�!���r��'<Y�7+�Řy&���Ͳ��+.�'�1��Yz�_X�c��hM��"�z�z�9�Z7�i,����v��40���i>��?�j�R2<x��}�c���0�~E�����MbGi��+s�$|��G��\�$��PW;��o���^a�b���������!<��Е8�8�{{�/�9l��AU.i7�<3��$�C3}?�C��{�=4�o�&����\�*�0�E����4�j�4lџ��ʄ�o���R�� ܚߌC�A��}H������^�شT9������<R��ꧦK�� �?�ՠ��ĵ���F���+�C�h*�I��:��6;���ɨ�����\Y�r@������;S|����$I�_6)���n�TP�d�=R����"��uB��T��^D�*
���
��$�9 ߂�JOpv�A���m"�Q
?{b��e�nօ5Ys^�a�g<���c�bI����H�V�1>���ZϢ#G���յ��/-[=�9�C�Y9d�j�ג���ez	zGDX��&����<�)�<��w�p�?Y��W�Hnj�©>�I�3?�q%;)oك���{�bC��#jB�+���� ��$a$�.X1w��tSbÑpR��o�z����!�6Z�O�<�)��6荸�E���[K�7wV�q��w��CNM��=zסg�q�#�:u��Ƶh��O�^�H���gN�aV����b;GcI���H�F_a�Z�KI�5����������:��ʟ^CwJ���
�M�L����~�0��y�;X���n��:7�E]�JȨs��8�1��5[K!���!I^�fw��:ՋPR,Ȗ��A�.4C_�䡮FN`+<8��;�jT[Y�Q���r��%p��	�.Hq^a0�~:�DԎV*�Q�S8d'#]��E�~��Q"�׃���<K;�c"�G�`]�mU>5��
�`�
$Y$7Au��Mlf�����s@ ���G�S�	U*\��5�yݩ���	;�i,�)C�vuC�������ݴ�1ǟ�C�Q>�PJ�.%ad5��Y��$X4��6b3��ų�,2d���X=sgwC��Ѡ1ZM�6�#s��9�h�r��|9�F���I�{�����MIe��I~~L����7�� 1�Ӄ�>�dv*���L�$��r9⊢�f���t�|��?�ӉZ9�v�:�#�^�P�`�}���뺗 5�N>�P	� W��=�!�C���u���v��Ҋ�fa���$���uo�v��=����S��ً�j��z6�'Z�����~�=&�׏�QJ#{bPm���	��]�S\���.��BSinp���VKǦk���9I\���������
������~�qy���[Mb��X0;����j0߆�M�:5����AǊ��ģ�*%���*omq�����m'��oXG1�򾯧[���g1���_vN\\Եf���58��>���oD���<>�����8�)�X��֎=�K�ʶ�<�u���.&[��n��&��X��/d���H���
Cpo��x�((`z<v����!SRc����X 7i%��P��<`F5���|=I�� �i�_1�&a錄�;Q�q�,b s���
|�8[)�*�9ue7��U}Ulw{]8�x��'hs���oo��k:�,�|�Pkh����ujL��12
,"&p�o��"�G���)*������T��`�Q��ÈV%�L)�1I����y,��f_,ȃϳ�q�+4)vok[�F�\H@�����6�4� �})������mm;��;dI;fHH�����lm"�;э��Ĥ��@�j���G!=�#�y��,�N�a�+Z	ݑ��SX����ن�t��So$�7�l=2��S2�w�A �gGv�+���}�e�h�ك%�������(8{�P�J��貞M	�< ���ݏ�S.f���9D	�s; �r���T..0?���ڗ~��Ss4�}�<����� ���K0�����F8�Ś+��Qf���S<�c�����~�w�����X�Xy�occ������·��_9��e�긦�������}t]���7Y":\�8���:a՜�G/����x��I;���|���Cຳ���������k�H�zW%+��J��i��Ĳ+���bw�ߣχ@�I�9&��y�M�l��BШ���q3�5�ЁX=�N���j-���z������� �O��a[�ާO8O��������ծ<)?��pK>M�ٯU��\	����I���1��D%�౛D�`p��-qΛR5�*��ʱ/�7�/h�{b��-��: TU���H�s�/j]h�}{�v��E�SR���	��(�#S."��� �1'H�EK�ՠ }FV,�Wnч�?L���R��a���ο��i�"��mˌ���D����FÁח��O����RQ)� R���ȻėJ�s�%<���MV�sC�_�]��@�ߴs�i	ҧ²'�-��E��J��A>�0�Ai�pv">Ў�Q���3�{�H��,���k�w�x]�֝�7:,¶�����N�4�KȂW�4�<��j�	�X-[j�&��CP�����i|���O����O��3�y\w%)Ǜ��
�a��A��)�RO^����M�ގ2���!�73�O^��~���h���v<����={�����#/�m'Ӈ�,{�3�=�:K�H��}����֎lM�����Y>k*o�m}�L�μ��D�_��6b1[z�B� �
�y�",}��� 0l����}П��/��J3��ֈѢsK��BmH��$M�nl�A��ǡ�$ط�-Y�;�^�'�m%��Έ�P� G���o��+���yG�7�6���k#������.�� 923�3��d�Z)����L�t�IEܹ[�~�c�'��ۿy?.�agO)V��@�{tTS�7�%w���	N�'z-�B�����(�ݩ�Y��ɶvJkq-7�i��&���Q����I[4�����?h�>�;�H}������;����` �Ņ]b��O@��Кk����N���9��<xU�w� ���ESdV-���A'+��~X�L=�u��X�6y���~?J=?^	
�bД�M �m�ǣ:Y�
��gkq�sW< A����j"͍�T(Z�}Xfz-(��1����+h�����3�#7�6xa��ʉ\�2�;wB2����c}R��p��=?׷��:��-�T�!�<Af��f9g�O��"���PU�Mdv�@)����?J�����@]��M���9 ���Au�q���z������C�|���]�"��;ת�K��EPf��,
�����u�nVq��r�ft�-�ڷ�?=K.G�����.|<7�^~��t(v:DN�1��ef j��Ϊ�c��^}Q5&�?9�[��Ϙ�0����|@�\�}"I�%<%�u���p��H<�h��\#�¥j
�g�F�Zң��kѐa}OEK�~��YS]�a�L�/�_��j�fL�<iFyЀW	�iZ験��UF��f��{5�0���B2��/q���G�H���eXeb!���ni��j'a��*�����	�#}���*O�dY0:A�&�U���V[!�$$�j�6M%-ە�-9���wf��Z��wٗ`�UU,yp���<��x�ZƓ)TwW�h�d������71F<v(T--͚�x�g�Z��
0�h8�Y�M�D �Dg�-9a$n��	�,���p�$�4��w�a��Y�W�x!��!/\[�7�k^��R�%Q�5�vQ�aC`���?}B��.n�ҝ���E�ÕN�5YNE=Yd�w�N���fK�:�5�3���Ӫ���Q��;˵n�y�B�a����͗u�L�OA����9�E�W�|�O�U=���隣z�L��dWO�E��a�c����5M�Ӗo�{�qi�0���T4�}���@�r�����l�|U�˩�e�ձO�9������#z���I�yz`����{& �Kj�&|"-(�� ���ޭ��~ vm�[Į�ڡ�{.��?nQc�1�
���tU v}����D�����喨Y:�PwG�*5���ay��ڝ�{�EO��*o�6�.	���>m�~#�5�]3��G�$����mFkr2*@��������2u���:B�4JvwvrQ���#�\7���O�,8��a��M�5m=�	z,���ƙtw҄�& �R��`�����Zf�al$4ϗ@Cn6Ԧߑ�
���)������� ��9~�����g����Q�=my'ʏ�Ik�ǉ��$у���5�IJ�w�%��&�SG'�֌{p�p�n_4�g�v�����5�aȤ���O��&���@���7�6d^��C�l�3�i��M����'��	��ƿo�V�A!��u\��O���	i>t��S-����zjڀ��Ճ~1Tf"T���o���Q�Z�[n��X ��p5����϶}�`GN��2Rds2˳��/.3�:<���F���Rԁ��F�-R��I�y^�s�T�t����Gާ���ڭ춪T9���r��V^�c�`0W�>yI|UE8�����.#���j.q6�G�����ɉ=��X�gg�!hLQ6�G*d�}8,[���Q���O[Dl=�r�Hv����؝G���
���u�q�\?�/��F��+�/�h�+'�&<�n���!�g���F��>��5��S�Tf0^�|1e���%`@n0TH]���s��u��[�]���Oc���BR���(택��ڏ��V�m�N���\�B}�}�i�.��h����+��Bܪ�V��������Z׈��ب���������w�2��v���_"��@�1R&Y}d��,,ECuX��%�	H��)���2��Oغ�̀������8�����T�II�mB�[��`*X���,�yv �?��fW��ɿ���H���SR���嚠C�e>�����0���͠ 6�����I\a�qԇ�r$3m�vDnn�-m�W#�6�BE����pdb�>�֨&|�Y~�.��R��i�����䃽�_� ��LyN�HO�es+��/֫f�� D���$��3�����	���0{�������Կ�����8;;҈��eN/�:���2Y~��¡�' 4`�6�-��ƲH��Eƣv���^��.*T�q�h(������`MY*.&�1�I�jPAI�+���n¨S��@�	 ��}gu���������I��>`+ɝ$��mŖ�T良w᧾�O��r��j�
us_'wJ賳ㅊ�ߚ:�,�N�K0�\�:�Y49ԶN?,����T٦�ɔb~��-�p����S�2}w�`]�D��u��}�	W�F��dǸ���bң�
�����Q�?�S��]e�.�Mq�I|����ĳQ��vfO5�k��f$�� 4����ٯ�a[�vyO��5Y�B+�H�>�q��lW�]H�iv�#0��� M�r �U���5ҧ��CS_az�?��ï��E͢���A��7��c�Ѝ��_�ys���[�P8o��IS�S���J�b�M�o*_���0{i-j)\̝PkP�k��v���