XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!FPO8J��-f^�.##Np���e�;c��M����<IoX/dcn9ZXh�n(T�S��M߈^/��P9�Ǯ�]��Ӧ�0������ ����h&=��7���Ta/̴�Rö�K>t�)�P��7�S��6�`�vC�O�]����P�M�9B7;�,�Y���%��@�/�!�I
9�i���1$�5ʂ�`~�b"��i��~g�C�Nm�@��kC�\I��c[	|�麷�(���݊?A1����f0��������-qՑ����pò^s�[P���	���r,7mdu���b���"��ZK�6%��-�,�l��V�g�NS�`�0�x�@����� �a�|a��4ie �>�.�:�gK���fz-T����YM���v:��l���y��( f�2��̶�༴P�>�Q,v����p�+�4�SKaG� 
�A��c��p��e�C�đ�4/A�*��p��ۨ��#,y��)�.���;��H6.�8��f�=(?(�m�d�ns/�t_�Z|K1)K��,5�wcA'B�MH����(��������{���e�w��l,�}��:��9%���fΎ\V�r��Q\�P�F&�B��4K!��u�Ӏ�iI����N3�T��[�έ��nN�"��?H�N�J�9��4�ʕi��7��^,������ ���>��g�	{�A��Yr���Y���6����T�Z�ǟ�U��5�=Hlh�J���e�	O�)x��-�XlxVHYEB     400     1e0��	����B��B��*9j��xܙ/�)���"��b�h}2�Ȗ�"LՒ�jT�#�_ Ѵ�T�P)m��icA�;�@��0�PTv��5X&�Oݲ6��LYU+4)�[�Kٓ��Z��.+[���R��Ql�"�I୅�=-�[ ?$��h`��]l���D�O��|[��D��5{^���Z�"��R�Q}dQ�d(lm�}����8t�-F����I>�48B��"]�G	$
Jx�����ő�D���.#]� Q:sZ ���6��6�X��lF0}��7o�e̠[<�묟�Y�\��o��G��������r����+?XUH��>\�FP�|�U`�? �ZLDwˉ���<�̽&���E�*�B%G���MvĐ�n��gD"���ڱ���mV�o&�txݫs�u��a��k����!��Dy�:,%���d.�8����B�E]��PP㌴a4ȅ&�p�3�A����s������2N�aTXlxVHYEB     400     160(<1��|�����m/M넢�.n��$�J`�"���UA%9�ՄD�������0ӭ��o�zm��҄8[�ԥ�-.�8�F��&���1�AK�h��!8��Wvk6��e�;@�hV�I^�R@~���z�"wY�����+N�q@cч\8Di�9i��渽�ĮOu+�,ƽԚ*��H�=�ҍ0�Z���~^[.�@S��j���"��'-o�!@H�ma;#��Yؐ�pū��J�������-(lP���(�hF�D����t�	�Vfv/%b̷���#�*$�4/��єd>��|��N�0c�}�1�5�2��1�OPx3t�"7a'ES/�k�Θ�߆�4��E��I�XlxVHYEB      50      50ac<��i6Uj Lw#��SI��@�I�-t%��#y�և�Tk�I��@�U�����CF᫆����G�WK!Dth�V�