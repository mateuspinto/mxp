XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����'va0��#��ѥg�WrD��[ꕽ����Z(�>��f>b����#A6ߢ��-�f����tc>�~D��W�^/v�>�f����d@���YKI%�С� 0T���a'KK���~jrS9k! ��ʣ�����0��H�*P���weNKT�agjT´g�y:��������f��)���c���R�+��$]:������(e7v	o�?��tS��T+�ܥ=����N��+���@��
-��C8E6�q;�]\`���F">�$���u��{2���o�Za"_8nw�oJuJY����%7ź��7CJN�<�ך�Ʈ�Il�K�MG�M�L�y�E{��DO~5�ǜ��;����m_Qr��RN�7<�M+�k�1�y���f���ں+�aO���-b�xD�� �����@4����b��<�OE5/)��m}��x��0���dq��nu���a�I�ܴ����W��,<�מҡ|�g�T�ؗ15�Y�����sEy�a�$�y���H��G?����^���j����0}�K�~����%$��������=�h�:��vWLk��#y(R߭j`>��+�c0��V����~i��I3
frwcP��p?4���bM�r�������(�&��=��i���x��%h�\�TAp�aV�*d���V���7N������lK�+��q</a��RѰ�Q�����K:���! �.��r6�I
'����;�W�0��8�Р��KoX&K)&KIT���5�OXlxVHYEB     400     190�n�[G+6��D�]ӺN<��4������$c���}^�n���9��i��eznS��.�=3Ś�`γ�T��VT��8({��)i���u'W�0���B�^�u�dNxG<�7��Od"�����D�jWw�6�l��UH�'.1�Bd_�ք��������@'ɘ*��R22����τPz.tP�h�O���{�'��@��/�N���jכ�) `��w$TU�x52C���r�ߞ����!��*�H�{)���o����1��t�I���\���v�T:a�&�H־�����=�Y���8+��w4����У�R1i�6r������[��ˊm��d1��~@/�k���A�@��l�����I- zj����>\E�XlxVHYEB     400     170��Ou����`�X����F1̏�� \ ,٤�Qv����)��adc.�ָݝ��q�8�x���V$�c7��lJagn՜��U�����j���B���P~6���F7�9��=���4�Z�J���iB�E���U�pH�$[�d!L�h���3q%�I�y�B�������J.5�@2J�b����d��V�ե�+���(��Uoa>+~��Gd���(`H�^��A�&"8��υRG_e�k�!���l�?CƊO|yVp���]�w��m�g�=�B�����2�:=פ��+}�W�M�\�1.�73jvOԞ��(��g�l���;1&���0?��3*`!W��b[�R���Ӆ�?�țXlxVHYEB     400     180�:O��o{fޔ|ʟbx�Jգ�e����S��5��~%��o��R�O�s���+�>3�?>X��f8|	�o��yS�ʡ_x�+��ɬ��"SI/P��JN矍l�"�׸ ���P����ȭn�aܣ��K�C�x�>�i]�0�͠�� )��Lh���#�a�C�� Q63$��wL�N�`밬Gb�p*���X�ňҧ�K�Bho�7g�p�,�W�3q#t��G"�6�K�������'V0��ؘ�6��8 �v��܈���/�|��"7��yY�&;D%����'���8e*��щŧ(F�ů���^'>��u
�Aee��*�L�[`T�6̌ڢ�����#�Ò��gb�e\��7��,��3�9'��|Ǉ�XlxVHYEB     400     150m����l��+VŴ|#c���p�f�u
��'L^�Z����*��
�����#���)O��6��N���B"�so� 6PE1�c��Xr0���p�p����ωyNm�nH�3Y��[+Ր$��~�3NW���������͞R�����n-���N���.a�H=��h���c����mos�)Z�̿6�m���E֫���>O����P�/�#�i`�8�N�M,>Vqf0��:�.kTP;�>u'QMҷ*����m��ݞ>���6k��\�>��xW����AR�*�t�0ێ�ŋ�Q9J�i���n:�z`��"��M�wiS%:��(>���XlxVHYEB     400     1700�(M4!oi,�.��C�[�Xy�^CFѼs�g$�o��7�!ev�C.M4��>�����I��I X!Ż�s���wL|\���Ã��%!�~�y�m����hj����SXl��"}=�]��-�IW��N�����紵���G���
Q���Qg��N���2l��tC�#7r�³;�.Q3��˫Ƶ�o� w��r 	G`h۵w�y7������omy���"aj�sH_#�"x��C�w~�6�_ʍu�8ӹ�I��F150m =7��'"��a��
Lg�,�VH6q{�$lF���dѴ ,��T��/�ȫ�r ���M�[Р�	c:����������H�=����N\� �Q�jx��\d#�A��8XlxVHYEB     400     1b0Q٥���bR#Y� �P����E�!b�C�2� ��;�>���jɻvJ���+�c�$�,�I
�h}�7��B>��7d�BỪ.1K׻����� t0_Ѻ�V�O���h�8c���=8|�q�����T�!��K��'��Z��IKq��R�_�ֿZ�Ф��1����r��rC�yo`��ר+
�Ѩ4�����$[L'�������k9��#�v����M�M��R��<y6 �!��K�)
n�]Љ脅S7��T��:k�O��./b[nr�%�<�P��������7�-��t<q�b�.d��%��XD%�r6�($=�9�� �TP4��}�L]d�f��ʤO�&~d-j>��������h��*�x�a�/u�O�
#�L��yB�b���C`e��$��w�Ktr���B
��~�j��D2���s<�/XlxVHYEB      e0      a0������dPh�Y��.�FLC ��ݖ��#���� [2`�������y�&4��뙼e��uR'�$����=������������&L�ʞ�9c�MKS�@ǘV�5-��EX�1��XйZ�q�����̦���>BGQ�)=�ZG�f���U�V}�����