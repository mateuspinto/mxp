��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����<VF��B�k��o�*D������b
/�G�d�}fW:GW�h6��$6^W���z�`W��Y0d#�G'8�y����	��{~�W�C�������^��z����O�:*4�$3��vƧ9=���Vù���n����atu���V,Mr���Ͼ���ӡ�[ȁ.d�0�JV}$�����MS���I4��9w1� ��U��ՌMԤ�Z�F��øǼ�bЬ� ~J񮅴�ў��v�z�o����G����)W�SOw��\���,u��W���'w�+i`��:�)������|<��cZ�=<{b��N� !��~@��]?�R!��Y��l9���.|-�6Ng��`е_����.o@�axA46Ӧ�Ҏy,�um:�>�m<e�h��ʎ���g����Toy\!J����f�."	8�
��`a�	�^���{���F	*��Z#$n���?���-��p	���GLYЪya�=J?N?�aE���([H'��~L;G-�.?���&Hk���C}�n�'�w;+�&�O"G*��vM���&]�_�Әe���ك0�7��1m�$*o�	P�{�B���3����������C9 o�$9cG(��ƈ�q6M����B<b�U�0�7�����9�?�=�Pi���0�%�%���`dI+�����1#u�� �gڿ�`�P�8犤o	�^_���<��H�s;���1	H��1��6��W\l��&�]�������#Ay�����aBoy��e��gn�`�ep�.�=�<EX�����{K�և�Á�����S��eoa��}�����_���W�g��g�S���ý%�چ�Mb��g�}��/�h�F�Š1!6�t�0`�귾m��qs�6���t5P��=����C�}�<�jh>�^�-���2NwF��g�;g޺���V��=��]:�$(��O�[F7�ٯ��7բk,�4��o=��4�pbCm)xK2徍��^iV�q���mN���X�o=�Ҏr�.\O���SMlZ"�dϢ���..�n$�J��^ăI���UY���<=l�2�aBh� +�� `p�K+�Fd���S5�<V�+h�ʫ�g�$Tnz)�!g�A�E8(i�H ��)�b�?�w�p�#�eyJƑ�ۊ��zO�s��-�~ǭ�qNN�R\��f� ��@��F�G�2��eE�#�H�$[ff<�2[�	�"ej�j�r�|}H���3�u��Χe�3�x�R�%~�Y9��Dz��Or�!λ5+��A�\��=���k� �"����b�bc��_Wx�N N�4͕������R��c@�n ^��PA,�r4Q�D�1\n���yeB�����g��i���H~N��k)/;Άlw	9o ��-п��D��8F��F�S)�F%ΩǄ��=(���;����n%��<���o/Xɀ�y�K6�+��hY �${Y7�x ��8���!g�G�������U��k�s��/>+Ge�!?��+C@���sj��+y��M~#Ih{
�~��iT'�9��V���� �~�'�.z�y�W��&F�>�4��5E��\��í-�=҄n#�o�ڶZ�N��E�G��8$,�rY�屯;+/r�3��ŗ�8����\7b�<4k��C��2���s��DȈ�j�)7�G�$R��"���5^��,�}GUaBO8�xaAj)-�$�hܞp��O/©Y�񝄧k!���]\+]+���6y7`�m�9���r-֤��"�O��G7<�u�����^����Ft�޻XCX�^��x;�&˟&���N[~�	�&�B��/�!�_,�q?�%3!���e���{�����q2@�
Q��ظI�ݹq��s�+2
r���6t�_p���+�C���m�P��t�
���~?fT�7�x�_����d��ѯ��*6_Ir^�9�sv�a�
��n�ƕ���(Ul��n8������Dȣ�o�+��"/��׮-��*A�>����s���qHDe�;����?��U�4�12�scX�:� ��93�$ �"g]!n��0�1��Z7E�L�+���~��+��KU/z-ӈ{)P���=������@)R�ɰq�L��R�k���|��
j4HPlL�O�����94�ρ	����?��Da�+]��S?����ν?p�9��Guu��n���I����.�{��4�~D�1�<o�S�5���,�d��У�Bˣy�AE�F��_��rU����V�o����N���ɨˤ�[KZv�W/A"�LP��Dv9�d�4�L<\Il���JZ� �w7���,��ˎ�m��M�̉�)�8�Zf���g�KbI���	!WUt��o�W`1�ltx��v�ԺQf����>�dT@��!Su�u�qZksb+�	��!D�����&�j��w�N95����-�u��( 6�f���,[i���%�c[_�x�)���x��
VKT���w^Tt|��d�*!2�0#"�>��W���f���kv;2YB���^��
}�Z ��M+������Q�4�.��T��y�8�,^=��	2Ҫ���y�R�8w����t��$����"H	C����ņSR��e�l��3(�I<oc,���y���i4b�%��؆�����D<⼙v��v.pD�=r-
! �$� ��3N�!����%�b���yS���N�i�zx[�D���`�ޟ���!�?{Z����@ه��}��T��?geʎ���`��z��&d�T��פ�o:πS����P�GU���M�R�p�q����a�� �C��Y��zq�����c.0�~
��"�z���A�7�����f.���m����C��S��.wϤ�?P�R�x���0�3�9Y�����ke6ˉ�$O����/�U��"��5������2>��
�b<^�� Ah��ƼP��Q�������8�*1 6�ӟ���,���`*�"�o$c����c���x�1'�ę9_:��r��?�Q�ZG��AE/�z��{�3HXRq8�B.������b�5��-&z{K׆R�����v�	�g�tz�} �V�F�|�;�T����)iKkU��t�z8K|��I��e}�\?T��隳V����}�X�c�"R���:Pӹz����m��ۙ��J<O�o���pm��=ܪ�����wR]������TrF@mע���/$o�����p�bI����&ѽ����g��w�k}��d���&¶Y�#�D�2�6_v!�P�I@1:������k�$�J�#)�jM�4v�q��w�w-����m���N����(�~+Q~�V�*��TW���4�Ή�z:""�W����`��p��p>:�h���gp���x�8�c�r1�s�Sq�a�,)�:���UV����׷_y��W�E�8�K�j����KM�p��'��=Ӭ���+�R���|�@��gB��>sbs���7;P���Ϗ��M��I�l�=�u#���A�3 �*1F�y�'�/�o�Q<R��Q��g�>��3��D�l�J_o� k�dlU�����p��Ș����r�M�y��$�K���}x���$-Ģ"������&��R�e��*�����Y:{	o�N#���04��B����"�΅��R� "����xӶ8���8Vl	�������e�	��}����l�k�@hvp�z�%�7l�,�.�?���z=̕΃�d:_��}�_��¤�4���)�����0�����2I��z���d ���(^Ċ�K��.~i'�/��ޏ�vyo_툟U����7�r��޿(��n����]4~ǻЊ2��+��r<XG	��/�sE9�p�=1��<-E�,��>�<���nC�)Y_	�ʪ���^J�y�ץ�F��44'�yֽy������EW��B:m�ї�d}��Y'''��^�$�?
?6W ;H�[�Vc�l'��4x±~�H&yoo��S �̕Ç�n�MM%Y/���a��)-42�6����/З.Ž?�h,'YB �x^X����+��6�zo	�}ֹ���r6��?D�ff'\���>�g6GQ(��*�i�L�?#�X��4�#n�11v��W�"4�_Uw����e
'�y��Г%�]�-Ѩ>�:��If"�.40�ڭx֪��k:�N�Ҫ��{�n�\�,��W�2���f�3�gPln(��so'I$H��"���`QK�{�|6�#hB	i�WA��+����CjxDzc+��p�cȷ�	y�m�I[�i��Uk��oN}�)ĕ�+���?ALt':�z}�O�'��[����*�R�K�7�l
B)�N�.�����M|F��������_�\��C��n��%Q�l�՜OR�x�l�+}�y���d���9JMi���� ��i��y6F���������5w�*��-���'�c��K�f��%</��8��>��/����Xz&,�2���18A.���դs�$ ~3۾�ǜ3���r��L�;=£�傎
%�+�$6>� u�ɾ�z�;?oK4��7��4��]W���HfLW���J�[/�#�8	v�������`fp)p�Ax�$���TƖq�Q��,��n_������� z���r��>R��(�]�S�[FY�
�򖠾�9��0��I=�"��Q'���8�-���������4HS�_��y_@�[_�Y�)-��Ӓ���>�O�̃������q���"��=���@Z!�Йt�]W�I���'#EV��}`[�� ��$FoY�8�"�����f��F�'�Ǵ�*Er�Iu�;�j3��.��b4綽%�����E���U���S8V��h��ay�b�l�������������߁eɬ��K�D��,���M����sJ�6��RuBٲ* ��r�e��:���dpKR'�Y�[���(��l�����S,x���ϯK��Pu?��itP�z<�^Rf�i4+̟�Q&<o�݌jr�uo2ĭ�T��s��bd�5e�}@�7���'�
P��|����<7�@~!�O]]�{�okY�
��d(�Gu��"�Վ?Kv~��Pk -��b�ZR-D׬�����S�C��n,E(��~^�]"~�S����OfFU4M{�pn�o_ׂ+��NI��������3V#u���,�rK/��G�ם?E���_e���?�I�q(�n�����׼EY��3F��P�~?�\;5'������+��~��h�N�L�M�<=�C
#g arK�)]�Z����U$`)]'

�3	,�qHbҋ�ћ��N�g��F:5�4Lz�O��Fؑ�Ά��V�>�M\X�P��P|�S���dYJ��T���a�w}3����C�j��y;�֎T�����o~{8����ܫ�r{_mJ}sj-y��e��~W9C��Tgca5�r�uHq&i�>�Oƫ}B����/��:��^u�,�i��{?�:�
�� `�#�����e�g{��J�n�(�_1P�}^�f ����O�K��p��wu����H����מ��Org5����Y�e��ɟ;�
�k� 7���k !`e]d�Dm�/�ːh��%��'|���0O��PhK���r�?��v�E�e�	�x�����1d7��b�� D�`)0����8a��^���G˺���g�E���]d���r���{�[n"�` >n7h-#�q�ʣ6��+���J5����d���}��Y�Du~�M�Ī��70�y5n�"�7
Zy�*c��T��AT�3���.MF����Y�-U�`4N��W�r�I2��n�$>��3�h��<��Lk�_r�f@OjH�v��6��B�<gXkQ�/�6H�W�H�"�ػ����i�>��'=�k����=n��K�?D�6���pCE��m|���CKe���1��]]�����w\�,�c��ړ9�QӚ?[�0s��"G��]/�-�����kq
���rO�-+�U�b�*]���
6$��$�8�H�䎔���C��݂@en':R�>��+Od2�~Ax�<���A����V�7P��1�3����7����������z�%V��ŕ�{�D�u=���%N��O�����&�ȑ��77]�nr �����&�󾯹ż9�mu4�F9���p[�́?�$��'-�G�q�=��)���U:˶mN����Dz�le%1�����`�)8/-'�#�Tޮ�0hv'����
.��#�;��lj�uܮ�
K������YߎMg,$�j5
�@0�}�'ΚP���Vk�����c���5��z�ŐD��1�t�z0��^]�MF�ɍ�V��`8ƪ_x:�͟\Y�ƕ�3��Np9�&]&p)�'BP[r���~?�R��ڧ֌�RO�����	V\�
�+�么�]{���'�R���O�n%E|Ҥ������f����1�,�z^�z��T�:&�� [�9v�aݛ��<~!�N琂>�iT	�wZ�"�p�ז{�ZdS�a{H�I����*������N@� 8�=j��r�H�օ�g'�@�����@�m6�/��h~��^��t�?krB}�c�0��l������Ý��G�5v�͔�[�G�L �hW���Q>�%����x�����5*b�Y�q{ԃ��5���H�WNۣnAm����[�-��S��L.>l�.TU�������3�sJͫ�2rd՘������u0TY���Iz���$�����.�����N�z�.�K�u_�3��@��çQ1�/F����紀\e 6��X�;��ϵ�;˓q45��?ڏ�qz��}^м���yi�|���-B3��M�:�0?��|ܐ�۝�¢��-�#�C�r<��X�
�GF�>un�t�-j1d�$VF��X�C�P���3aDRuܢ����1<ՌQ�S��l�f��ԀZ�T�+�O��*�%%K��X/	5��9�i!C`�i�w��"&9�U�*������%�ƩmrH;�V��q��F���T��>_C��03E`<K=��=��.'��پ���!�#�X��\��j3��~�&�� ��s�������/����;�<#��J�+�S9ĂX��<ŧ	�w��y�G�R�i���ua�T[���L�DE�����7� /�i4�'��#>����<�e������w��r��ҧ�pX��R�tT��YC�!w��S�/��}�P�.���*���n!��i�6O��t���ЮS�Z'�"�˩��@͢�ǈ��Su����D�`>��oF����#���)�-��E�v��рrZ�en�g~� ZڵN�tl�S�J��)PL^��]m{ [�f�F@K�p��1b�D:��R�yqJ)�y�ea^3�"��5�����j̫S����0��a����I�݃�3<�4�ё5��p��G���x?��G��l]H��Whl�M�k�T*3ō���=Dv��[��K�^���/ގ��pBJƇ�Ł^��ٝ2a�9$�R�ct��yY*�����:�
�-c=BC�5�T�V@E ��H��~Y(���-���{����_-i1aQ��64��dã���TZc�C��� �dJ6���զ� �5�N��Ȣ��+����.s�X������~�hrYs��R7?�����c��L=�ɩ�B��Z�p��F�=�apy���ԏU� ʓ��p|���#gJN�I����AҠ�4���gB�\���ZI��Kq�?��^�=���!YK[�F����q���F��,��*R��.��T��d8�SJ�,t$]����cV�G���1hٚd�LRzN+�ǽ+n���ZNbD L>#��fT�2הT�;��eշ ���b`�	;"0;�� J�����b���C��o��!�G�1�
X̆>���FnO�|#���m	�Y6�w+���ҋє(�9�y���y��w�w��~M�0��sE�U�U�T]��|���46�|�^�Hk�Mܞ,�D�NOx��Es2��C�9{r�"搻�C*�Z�g�NJ�?N�\~("-�D�lp5�d���>;���iH���� v���`�ɋ��5��"( 2U(�3 ��BB�RX���m�}�jy�D���� 6��/\{']�༇x�b�P=�!=�_���c�kp�ڎLz�X��&�y�뿀�%�L]�Qa(T�����}�����_���������{���ƣ]l��z���>�T.Tې�ޖ�����/?�5٬�����7EK�Z� ��������:��o���|�8�6b/����ck·�XD;��m��
	46��_�HF��8�����}4[b��9_��n���v�lI�d��H��U����=�<|E�j��7D�E�{�����h �"$IUC�-�̙�2�<���������s�4 ��`�#<>�3�g�ii5� �D#��1�}�����|�8ZL��?���#�l#-�:�E��#��O���<���ȁ�t3�?ٕI�dm�="�%b����ϖ��e�**�P������� Z���{[+���4(�2���v+G���_������:A���
�?#�'�'m�ğ��g�ɯ��� ��;��>=�߈}&TP<�'.���`�ֈ��f��Z�a�S�>fTK���S�9��<7�r�nA����B�9啊OzX^EX��zIQ`g�id�tT�]��l����ro��ň����#v�Z�wNё\�9�>l��F +)�� .?
�m����n%�O2�Y�/�����3zK�F�?��(��	�]2v�}F#ʕ	kY;7i5�����=�ȕ����-�����E�15�Sjq}7B+���!c�{�����aH�K�n���QW)���|�o_����3� B�1)������' x1��g��zg��o�]�����D{�hU�"p:ghd]�[�M��xG���Қ������w�`��'��+M�X��/旨�&�@;]Y�R�,�zZHī��-$a��kL��.U,gW�
��z�)�Y����Z����5X[�w�n+q��w_�ȑ`�3�RЪ+�޿�HZ�<B-�����yē�ݶ
�O"��]؟r�ơ�Y؎�\��qû�u
ֱ���l��W�W}v�̐W����kQ��7��i��h��!��S=�7��i�{�&����'�R"B��<�g/���/Ɇ�\��U}ʭ��2�5���Ӹl`V@cM��̫��iG-��<�����(�� ���r.�.�>8g�f�����eE�H�u"��S�|D*�8�{���/<Exjz�@��5ʫ�>��e�бD�`�u��S"�*W����һ�����%��0~��h�Kf\I}'JR�ڨ������.���Q�z-�ް��k��Ξ�>��h.��pEr�xAD�k��Qh�=����7Y�LY]�R��e�:QvB4��q>?��FyN�����S��"8�A�������R��λ�F>�َ����e��m�s�|�73Jo��qD��;�tb��KG*Kv��<�)����@���x6�ْ�ZpL�FР5ad#�4�hP�Y�ߏ`�d3�;�A��Ⱦ�H���];�[lQb��=_-��8�R��C�	��=��J4�7)L�F���A�X��Hr�jaD���"� �H�s��\�C�ژ��X]��/�@��9�9}l� ɫɳf�*�����zT��p������	���������ݧe�pZ�*50I�"���A#�����%�%�G�(��x���B(���+Fb(��$um�6rt̓����	˵ɦ�:T��˴��{�>��)�Y����T#�����C��P �U��U�L�;�x�
��?���^���>n��9��tYҍ�6Z�W'����Δ:��r�^�W�h�����S���W��)lЛ�,~�I��3��$�7�^��D@��o'���{#�)� B��3���As<���Q��Nl���$�%���z�Z�IzY�����}K��yy��*��+���}�(��hߙ)%Aon�1Fqh-g���@׳ ��Z���4�,d�>0W�cV벨��-�:dA6�(����i�(NP�*�w�2�fD����{-��:�(1Z�"��z���M�~g'��}"��!��N���6���-gN��|�R������H⇮[h��֤�O�ݹ!8
r�W�L4�uͮ"l�Ѿ'��\�2֯NƵ��r�z�)��Aq�.��*&���^46�j|59�zP��>|���8�/'��!$�!q_���}���k?M�"1��U��_h�[�?D`]`��N�.�a�]��(�0⌭F��K�+�d/���m�Ò�6�-�t��:Ģ��ϣ�X[%��`F��~�NgƷbA�KN*h H�d���y�𓥸�8 �)���B��"�nm��%��(W�4/ZaV7�>�p"��� LGG:����%�zN
IC�?�����t�g���ru��Q�eu�,�r�A%2��u��)Z�����|�{o�Y�hس37�B����%�ӭz�{w�����ۅ(%x̯���J�F��� s&��M�z����u�E�Р���Z�������Mr/�4P��,�M�L��<�������i2?�Ϧ��L��~�b�����|���Y$TN�=Ί�gE�.�����6���h�Тym��/?ơ2�'9\���6���!���v�ܫ�?ã��J��bZ^;N���o7 x��H��<;���C��yxheں4�Ϲ��p?q��+����M��wR�_�@@E�UͰ���=��������-{6*��	t�OL��� G�s�B��֎�d�������j���2D�vI>�/o���4�~*���@f���=��h�CU��bLC�/>%��
�Ax<����$Yr$Q�2إ��8[~��NŅV����cإ�����/�*��{:L�dks��W�Uf���i��4'��������Z!�j��ndJ�ˉ$��
$�!׋;|�.��Ή?�%�y�z�^�ʕ-�D� ���H�e��g2i0z䓿�Jl4��O{�J�9���n��4�eX��k:'<}�f-7���w��Ι]�_ך�o���ǟ��D�RT�J��k��{F)�ޝ�������ˉ���eG��j^N�w6�%5]
�9���Ce@0���p�򂭱��e���Er�P�o�1�B��<�kG:hU���ǜ�S3�Beő�(��Q�2N��=�\w�W�viX`T$��ߑ��3�9�wg�
N&xi> xM1���և�t\yϼ�4�3a�BKV+�c��~L���ɮ���a����T�1���d'�	�Nt��@v}���D��E-w� 䡣?,���1�
v)�T��%����tx(���$�Y���`�Wt��9�w1���b���C�a�u�,6l%�O�wZTTk�'�,�RW�B�-���Ҟ�G�:��5uKq�^��n����p���lwǯ�%͉��(���)��=��#�>�p��*���O�_��g�%C�
����ޤ$�+���
u�f:H\P�I)3k�z6I�s%s���w]`]B�&��^�+�F"�����v��'߹ �M�,��z)���g���GZe���si3PN�WGZL���,P<k>���N�$�mk�)�G%��Me��sJ��W�dόZ'��xT�˪��9-N$��g������oy�<K͌a�B����wi�3���~
��S'*��17��H�a�6-�@!�����Ov���WA8hI�Mv�X{~D���{����C��6��ހ�"��yG��qm)Yw�M4��1��B�\ ̺*�*
�'��mr��y�2qk��x�_�\���>�#����הӤh�ihg2t��-�U��p�8Z � 2�ɢ�E��=ˈ?6s��l����ڣbn�Eaf�@�L����ye��x�a�֮{͋l n�@akK'�����y�n��Z�.&��<%)����I!��X;L&�-�n�W���!p����A���O�D�nNq�|����Ѿm��{�����gQ�)P�n����QfG��Mm]��M��s��]�w��|���G�Vk �G�;ӟ�`����Ͷ�uڥ�)��6���:�W�2�}w��u��Υ�\�m4�Ѫ�i�5�Ɓ���z#�����r_�k���4����T[�F.�uRzl���>�;���3��VO���Z�����f���RIM%����%/����@�C�� �I΅�\M�L}:�3I��⠜pҠ���9̱���"
U�����bB�㡽�;�C��>��������	�j�}��sB91/����.7`?��<���9�S��(5�H�p�ݫ������3���h�\�2�K4�x>�C���\����;{��a�3�	�A����s, q,ϸ�=p�Ҫ���`u���Πo�_!GC'ⶵg�n���݂��:��`I:i�~�VM����t��KY���t�������crJ�)�ܩm�0���f��������]��<��1�J=&s�Zy�D-�>w/DOv��3p`�g�'�L�~����˄��3�kfn�?��;����"N�~%�XH1��5IOO��OJZϮ����3j?f��ҭ�0E|'j�%"4P�K�L+)9gk�ݮ�leBGi��'�h��)��9N�)���;�Y �<�[j2[�ˈg+���:��I#?х|d��8��h7g�I\�<;zuI�Enq�3��5�%5��z�Zz����Q����ـ,�M��f��*D��|,fcQ������Y�l�\���6X��[aƳ�]��S�'G�V:���/��S�����r���V��U:X���r�M����u�a�FbMܘQ��@�f�l���"Hk�cgV�:~�5�^K��Ԉ�byp����/�aS��::�i$Y�g,�N��^Z���޻��|�Q���d5T��.�G1�Z�\����?%�@�+�&u���U+� �/o5�;�冄D���i|�� kD���&bA]��x��T���"���c�>�+��PX�=Ǎ�+�`��$	4pg��ik?΂�l�f뉞�_�X$�E�+�{�|s�Gfo��'��Z~�=��2��z��pVx���pϞ�T�sAʸ��M��S�3Ae44�S�e���l�)�'H�s��l�ޓ~m��9idi����(�Sd�zC���W�ߘ����ql�T�C[%��	?��;"�(D�\h�ԓ��&�s��[l\� ��I��?,^�6��g��VFq I4?� �=��\ _�d#��q��]$�ܛs,J"}�^��FI���W��Aa��t�h�gH���T���sqȳҴر�1�>�<��=������>�H�<s�^�S��A��(&�ٷ���M1�̭d4�Jv����s~����7*Wr����|8��X����>C"?����W߭`D��Y�x�k�҂+A̒��Wb�Z�p���E")@m��~��­t5!O˃˘8����3�\��ͅ0T���?G��`���y�C��\~	�E��R*���㳍��;�
����Ե{}�dݑN���(p-{1Lh��E��~zw�� mR�mc0��->� ~gM���L'�l󑖢���*�t[㻸*��i.�#�g��lS�L��i�ߘ���i��?����'��u��\{�w�j�����h��?��2/�k���{�M�X�����< 嵊�}4�ܺ�?���?qd7]1�,��R\6���c��i'�ۂ�o�;b�_��E^@�W4�@j�צ]�9�C���tx�D/5�i�f
�6��ء#8_т��m,xL1F�z�`����Ef*U�3�FJHB�c7k���乔���B�?�6sL���$j=����_e����j�"?&�C��p�[�8g#���my+Xq�����}��ő�oYgK�\AϷzBΰ&w �x�*�&�eH=cz�./�F�xv"�T>W����"�>���:��
*M�Q�G���#<���=teZj��}�Mܚ����8�%����|��,l���[^fd(��Ukt�T00O��|l��Z�6�!��\��
�/�ȻP�6��������_��vsӃ��o� ���1�r]'6��J2��O	�i�L�I�-�	ŝ���x?T%� lj
�/��UN�r�R���{2F���H���|-\Q������t
f)��8���g]Y��6���忻hW.P'�f@��5ԅG��Ń��gxS� r/��H@��N��~gx��<��O�0@2��)�$��Ǻ�s�d��X�)�l���"��Ik%B���d�2���^.�\���`׿�Ăy���ssçVʠ�6sQ�7�mT�9��G�#Z�Ǵ������ni��^��W��O����b.׉�[�k�R\A	���M��Ò���>8_,��a�ܙ�$������P�W��Ț�'�������<�1��#��/�P�h�B�j��Z�iYe�!��9~�$��5�9r��v<h��f�Yt���A5W`�G�lS�ȝ��}I��ؠ"��{$�7W9�v�zҮܼ��ۏ�#�]U�]���)J����[�ͷ�|�����/��գϭ�uM�wAse=����p�K���Dʱ$l�F����B�ԁQ���g��6�����,n$�+kΓ	��(B�u���Jb���Ｘ��J=/�.b�G�o i{��o���G�!�C]�8q}ZW�i�l#�?��D�i�ϋL'@�җu�8��m�������Ӽ�
�B]�ԇ�rd�Fe|3!�K;���0��n���Q�ܨ�'�Q1�s��?���ʎ#������$̏���j��[p���I�D &ݡ�����S�޼2)*}���sJ���Ŧ�\`H��?�"�
����T��.����a��>^^��E��I��Np`�6����Y��e�Ǫ�"�� ��sǁ���,2�}��[�>���m��ԋ��nW����5cF�����\G�IZ*�ze'�q��u8B�Rn	�3V .�LR����e_���u�]�|"��Z� �&Վ�������)��.��^��%`���dC��R�֮�`ɓz�`pV�'�7s����ѣX����=E�x��2���I��c���{�ȑ0qy *-<�Uz����Å� ѬOe�j_��2�����Ȏ#B%�稈��I���n]x��<�nY��&}���u�	����ǉ�����'*�w���b4=��8�C�b��J�dcjD���7�Pm;�vi�� ��4�r�1����)��� �6�a���[��R0�ä�А)��C眞6�tw�1(�	�5�X�@��>B�Ҫ�啖��t�:~lR�Rw� �]b0��n�}�5�/&u,n%�� E�ü�σB���w4�T���i�T���ݖMՂ�ۨpw�˻osy�7�f	٥\�?�揪�p���y9j?�Te��ԸKi/�A�n�ۆ������e� W)U��@�ˤ�fw�y�������-�\)4L�DD>��������EU�@�9?�T�J,?&� �#Dh:!vj��G�TFIҖE\���J��b�'�=O������|��tTX��*�H��z�y�~͍puO���V@!��l~Q0z���\m�>� �D!���[���ʶ�C4S�Tp����؋k[�S���Q�Q�?�4���N�{9�Ofݦq	�NEb���>݌J^[�h��M��p�n
����'�|bi���|<n��3�B����5�h�Nŝ-�e��Dw�Q� k+��b�T��ߨ�(B�"�Y��XW��^�2��}0Z>N�.�f���z�	��
ae �|����Q5�(�OH��˩<f#�a�	WF�0I��Q��T���+_�S��@cw��@�xa/~ka;+\�
#��B"A�"G���o��D}�r��ҖT���E /�A@& tx���,kMu�ҺG�U�0����?���Z1�Og����:V���*Z�o�ͯ������R�~j�F�=g�*�0��J��\c1����
�C��>.FV��SG�C�����3R*�nFDCI��b�U�Tƿ	��P|�pS/�ז�=�	��1AQ��!¸`|���(�o����^I���O��R�D ]�#�<�wUMO �4�#ȩ��C�p:Օ���Y{F|�嫊��9���҅���ق6p�=��wv��ѵ��^G��L��S��xL�$�{ȅ��/D�7�1~#A�!�E�2B/\o�����5R������ί^�4�_^�6�3�@1P�o�t���⪔6�6.n��#~�D�  [z�d�=�+�y �t5����77����7lIZ�w��A!� 툲R��%�-�T����h� �қ��\!3�tA��
u��}�t�<��U68���
��ӈrɮV�*�PL}�ͨ���+�2TyL6;�t{�Or�:�$��dǼ��%���O�ŪcSUL�wq,�L�(G�1�`�݅����6�n�������D�pHv���4�P��x�+�",��Ƌ�ځ�e��yQ����������h-җ�Y�J5M���@���w�4�Mso��He�a.X��`=�h�o��X}�)_@�>eOb��~fa�4Q��ҍ5�q\�c�p�)فˁ�'�m�� �]���B��MM��cGl�3�Ag��AEh8�>C�^e�:���P�(��m:�A�@�ӿ�LJpu-��$�y�_ѥ�(o�����/Pj�(�vv)q�<���-V≡u0����p�|�Z^��nƅ+���	���düm�T
��/�b�(��%a�]}ƌ��"޳R��i:"�.U��4� %��։���ů˫��^P��P�:�C 8�c��fZ�Jw�2`/Q�U�a"�$��N� �,l;9͝�+e�I�j	�u�vOe��1��$���iX<5ߦE��Ƥ�.� �p�����Y}v �+�4p�m���t��_��eE�bƍ�<���,8�r���{���͉�K��L��_�����k�<oq�-��c����I�a����IusҒ���)
kOqT�o�;N��)t��c6`k/�B��ۚza�Z�P"�ޯx�7G�P�Z<��!A�p�"w���ϋ�UG2�o�G֙��Lp�)�c�0U� ��
І-�8X� �q�+��(5a�%4�ή=�/���h�ȉQ,��AfXޙ2!a��:����`n1�n�qKm{��Z.b���w��QQ�J�,<
wO�V����LƵ��Ց�g�$. �)pb�x��LI�O�=_:E��J;�y�;�*��}����3`�B F>�@9��ZcU�(�s����rj�������HFO� �u�ĴC���bc��Zz�w���Y�H���j�I��.��F0�j\�>�bH{��z���ۯ>L�W�W�t�;��(�p��W���0�k��Q[�_����E�|�k��|#�}�l���O��~�B1�\��_�O�4	� `��p�;��^�{w�Q�|�#��.�\��s���1�/��?O�m����N�ȩ��giM4=p�w��`?���N����i��<~�eu����!n��e�m�P}<�߂<`!C����#PܮR������esx��9�mj��2��.�,V�(��~s�r]߸��͵�T�g�E�?���i)9=U�ki���H����q-����������A�qj�Y�9��`��yRQD�ѵ������a��$�h�s�]3�6Q7���6��G���K:�m;Og�r��*fV�Y�$? }f���0�7���ܯ��M��ܸ,��cM��jř���q{�Z�w�/?�����0C��&�3 t�l�[5XaƂ~݈x�DD�����R-���w_��ش��(`���e� �`@;m� 2;o���r�o�X �,��~*|7�m��>��{ܐ	�#-'t��Z�4�����an�BfS���>w�dL�X�Ļ��Շ�]zϵ�EG$3��i��Iv�$�49Q��d�\�O%�ъ[o�]�iT$��A�H0�|)�MV	�:#��y�^w��ϔ�/s�u�Rס$/��Wa�!N���In�@0`�CQ��P���D�����Z," r"r@_�%ңI�U�*؟�����):9�R�f�9����<:0����(��db�0玥 ;n4�\B�@�Ln ^��u�q�,n��C��"F����~nL��)��*�O��ɖ��]�;3}�i�y���=�'��/p��@�ϕ-�T���ִ˭Ct��_!�ƭ�İ|Vq\I .�'�kV��j��R򰮴��nC
�hq�J��Q��C��Jc��v{��
��M�����7�7[���(����5un��c�Z{9��JU�Z��,B����Z4ceQYX8:TI��:��o$l�vQ�VyE3�����l>M����>�����#N��>w׃�D��N���e��AjQ(�±��%�LEVה����ʨ��tcJ����4�5�.�Q~q��z���5���o_b�G��G=��u�V4A��[��4~,y<�e���#O޲x�W=��׃,��DE��uXU��<��~���Nf�em�?���ѓ����+�RC���������/�ob:)����[CƓɝt����'��`�����)�V���P���N� �9������R��z;I[��_Ӻ���-�7��TF��Kd'��D�Ly�͞���rY�(��͢��B~P�k<�r�X{��$��4*zG/��3�I�ON�rw�|�k�GJ��M����f"O d��q��)���vj0�;�-�g6}���ڍ{�	}_�i�8Rl�ď����]GB���n@w7X*tw�P�b)A�W�R���!+Z����K1�^��F���E�x/+�O��w�v�]j�Pq�(�⥉�?�Oovhy���ʕ�Hz;�L��dtK`�]:�8������ҽ�<x�O�*� ֙ ��� �by���sv��tt���I����R-��4�wy�u䓅�b�k݃|W��K��0v�A0A̖T鐩��-��d,9��>_�l,
�6�!��q(�0Lg\ 2}Z �|p�����I5��`�\�4���%����~/<���ա�G7���b �MK|���5�Ȼ����0#G랁�$n3M������ő�t�����d�E�P�j3q��� aԵ�Q�C���d�o��h�n*�����F��o�o���Ȋ`�|���U���I��tϷ@�-�Y�g3��@ҜCY弲��lJ�Jq �V���=L�}F/��Dط$:��/�#q�p�ԧZ��*!�0�o,,Gq�<%.Pp���Q~ê�E�с�BpI0|��� 	��`�p�$������m�<��A+�o+��͠-�㽝,�ݝL���>מ���u��dV6X	
0g����/xG�9�_�6�g�䳤���c��I�y�e��=9��s��!�n#����:Tx���܏����8W+
�P��I���h;�XaM�^�H�==Y�:"��,�;��	�SVC�pKƮ��>�:>q�_dZ��Uw4�h��u;?��w�wW�Nh���%���<�:���O�I�<>iD|�S��eci���zF���ʝ�V8�uG���0��?���L[��
��L�h���!WJ�<w�y�d�v�'������*�i�O�.��o��yp���f+e�ScЮI"�}����'������cj"���Q(���lTڇ<���x�3]2�ѥ�2���
�NU���j��KB�)z'���h4�M2{�r*��+��M�M�]�j���q'9���>��rn���1��b�C���?O)(m����n퀧�`Q�	��d��ݛ��ٜ�a��l_]R�V�c.T�x�U���|e����l��'9~������+�"�#�@�hU;�hB�y��)�sd˨U�Y_&%h��X�SZ������Mŧ+��}b ��nrf�������d��ڴ�+[�~@ee��9V��1��w2��K#g�X�m"V!A+�-M:#C����QF�+��-#�΢��.HH�u�tacze��Sɱ��,?ۦ HN��@�}�L�&D�ꥨ����t�G�Ou]o�\.7k� �� �߀Au�\&RgWj4G8D��9�?�敄.�xP���E��"�OQ��������p0o��1v���d��\�T�çk8�k����n�4�7q�]�+i�)4�Q>��y.i�y�u��B�~����`�ˁf�xB'�ȕ��gG�p@�^o4i��L�N�_p�wb�`ϔ���z� h��$�E�&E��FT1N�1 ��P�n�@Z�3?�Gy��t�Iai�nQ��D&]�%z(��1���M�3Ɩ�2�j��
�����Q����M�"Y�)k8q��� �!�4��"�b|�؉N�.p<;ɽ�	�v���/E�ה�Y�Ԙ]�G�^;N����C����_^�^E�_h`�K9[�4�&˗e)9�m{a���D�&�A��z���o��չx`h�MN�W�I`�%������N�x�/��`�gSH�Mj���#QV	�q��%P���t7�{`"�����uC��l,Ο���'��5j҇kH��\E�
�����>bS���J�	��{��v#UY���kAX�X��+dF܍GSL�Ib(5�I�4CÿM��j0ü��w��	-w��p�VS���i�抻@�.��uz�
�}w�M)ZH������\N~޼F�{W�	lYD`���J-ޤA���)zn3U�D�lJ�am��MV��~��,͢]��V4l��M���H_vN�ѱꀾ�-��s�?���C��p�oW3F�?Uep�	��ޭ$������`- ���~h�"�h~���1�^��g�f���6~_�4>wUh�UW^��4����[�B�� [CJ�^ڦVD�s�p��o�Ϣ��d���DH*#�>~L�Q|��q��*d�w�m��^eЀ�5✧��VO?��Õ4N|ѡ@���� �4գ����ӡ-7�ޛ�$ɚR$��"}>�~�di��>�d�@�G�1����鷫��9�}|�f���d�`���LIq�qw�Q���HO�0$;:9�vzb6�_�已��xI�N�
��|�������`���� 7�7�C/d; ��%�����Wc�d��P���fS�k��ÁP7}SE��SCĭ��LB�ƒ���@����y���`x� ��i���<\tҋ�ۃ�;+��%�eGɤ���-�6"� �W�13���_��Q&��-�{|��lX���Dl5=�>L������c��� 6_1�e����R�yKޤK�<��Fݱ7ч�Snѵ�Z�̡6�׼ض�[Jp��'*R���J`�d2j�Q$�{��X��`�3��1)�ü��k��<��!������w����8�)}oA	���W�V��sK���1K<ƛd��'�X���^�M�O��@�@o;���w�H�L�`�ȹ���MS��D��K��[��؃�L���f�\W�[�%i�}��W9h�B�5�p]u���z�¼l�vt;��_�:��N��2l}��xi��̤:(�>}2;(MKK�`\�h���K+{��.>vɦ����]}
;<0��<��g�#�6X�ʐQ�˨?Eq��-h?D�ÍT�۵�y��P��iֹ���0wZ�/@�X7r'ޕH��j�N�ĝJ
�|��W=���$O�yG�ݩ_�R\�4n�Y! �a� Z�K4�37z��"\�xU�dEq櫯�wvt�ȼ�r�{��A��ϬB�8�˥Z��296����fi�J	���rT'�g8�|A�'f��H��S�N�:���u{�}4l�4u��+�.��K��@��U۳��W�2Ns�׫�o�@�vFcH�n�G���e���, ����P�|�סk�N���׌�L\���6�Ϯ;+��?_�1_Q�	;�\dNַkR�dt�E�g�9kME�8���&�h�F�����x�r��qJ��Y��2�A'��ko�56d8�zG^	H/�N7	�N'���°��8)`��b;v��O`ߵ+��|�w�ڭ��ʳw�a����|`��o��#��)��E����HʚE��:),^��8�;� �D�����-C��}5����%]{�q���i��*���;A$��ڞ��#X��Y�(�4Ź�ܚfl3�0+�86�ƅ�ԭ���T��N-�Y��S�I�����Qf��y1��},V?e��n�r�Ņ�7���_�N\�o+_t�@�e=N�LzW�O���^���S)WR)�6jX	���B���:���4�uZ�;v�[Ą���eZ.������/}Z��<r��K��p��
�+Q�kx�Q{j%>��@g�KGAT-}m��K���9w��o&���e����'��
K�<�$�AR���G���FQ�[(�_"	���tre�=����=��t���;�ۏ;y=O�� \yQ�ek�����%�c崎9�]noES�_�̝�+�����h�\��h����	���6d#��E��=���	�����)9Ļ�GK���=��N�!t��-����}��%��9�p�RX�sЧ�N�yсv��*y`�#W��Nh$z��v����"ۄ�r�&O� 3�<��Iď���\��X���*���ns��*u��=����U$qk���������$JZT~� fD��H1��o�Y��g��~�7��^��5E�~ Oo5��+�QC��]��0���M�w^�3Q���O�q�S�p��T)B);1�<�(���	�.��9T��i;g^D�C3�A'������Sf��ܧn�˳�bi��s��J�
��QDլ��l�)�{N܇���@7�~�ٖ,��_WFK��Z��F˼և���d�� ��[��u{�u��Ey�dk\�����LZe%��C�xHI�ڟ�q9eU�8�t��4hn��k����l���*9���҂�����cƨ�"���"����1��83�H8'��c����qE��b;�V-Q[�01�tEa4P"��mY۠;�gP�l����i@v��4���$�x��1P�������L?��&<�@�4�s�C.�$�-���Q\�G2�~@���lR~*H&p�۸��g�q '���1T72j�\%.i��RW��`�]&�f0)"!���gX;���A7������_l`�Rز����»�Un�#���A�Hk)���Z#z�\D��e�n�`���&��SoV����<�M��f@�u�,�B�8��2M��F�����u��`��Ǖ��wԪ$#�Թ����&�t���eb���Y"���x�֯�IP��������Y/
w�pa�*��� ��sA���������ى��{�4_���E�>�K��&s�wll����D���LI�4rV���9���g�;#���VD�6���Ք�R8��Ù�-+����^pܐ�$��g@ĳ��;i�Б?ٺY�f�,��O�)e�� �:A%
g��� 6h!���$'�+����[tÝCL�c��N��U�����{�W>�0��d��pxO/K h��mk{�<)ĸ�8��@$c;��D���c�V��ګ0=W��P�$��i�b㚩�)����z@b#7��6�FR7�Z���ik�h�]�͍^@y|��:d>W�Y��kʘ��o	v��f�����B?�)�0E{)�;��c	2�y�'!�P�*�!���R\q�id=#��d�V�boiՀ%6�P�B]9~TP���v/w+� H`|�Zz�� C	�~�Ӛ�*���9���P�/'e- ��+��+0�gJ&V
^t�C�Q�\���6�B�0T�c=�%n����ojDQU�cz윛5e��z)&|�SЅr`.~wQ$|6�c���$�b#�Vʝ#@+���9� ����'}7�I����0�Je�A�ȼ� ��������v��0�3|�jN/�65PͬK��g�y��w\�*p�!<o���i��-�]���9o�7O��s~b�;���0���\��"'�t��V�q�~n�i�_D/�������-��E禾�w3�g;-����hQeZ������k�r���d����O����:lZ�V���<!%�h�f�X�F�bQ�v�]��EVx�"鮷��TJ$'��ۙFht<�f��C�%�PW`Û�޿�<s:��?l��&\���S��`��27�sZ7T\��l�Fd^xZ}��LR�r�G����Ĩ�Ŧ����v<,�+}�ũ��|A/PS�4 4���>�=��B�Q��z|E=�����OTԮW�*�O��Υ"�@��ˈ�Ol��C�̿��!�k��ة;�/�̯:\Sru�Š�0��R|��+���Y���l��*��ʐh@l~??��C�Ut�k(z੮�`��ħ��g�w�3�c�n��9j����hoހ����������xm�uP�r�C�3]`�f][$ml�I�".����3׉/�k��H�Y��4S9@���D�~��ޣ峌�D�^tb�^��$�܅!�;�?��ǼZyzU��xi�����QK_q��컯IT)��W��1�F�WZ�>��f~� ��&�]�~�[J�h[ɇ�ceE�Zxޑ�':O��s4$�pޓ#�4�F�rT�jbPfGY��]=s}ľ��b<��%�B7R�t��0�{�����6��YE��ċ=eW�B.Ol �4D4ԙ7T��6��h^c��"�<	PB%�К�'��4B����`D�!���n���P�RAYX�X����Q8Ke�������7���\"�-}���r��cO�@�y��>ݗ�j%'�Cr�ͮ{y�Ҝ��_���)c���IzB6��~z]O����;�}YC��w�Жs� A>CR6��oL������|�8���(�y�3��&�}�PZ�\��˲�xP�Y&Oth�}�N��)�sp�"s�M}Z.{��uR����iecq���՜F@#9�듍ɒډp�v��+iA0�1���R�`TL��ZuG� �~q1Y���n�1��u&�ť���}�zZ\��KYD
�;����?��;eNQ���j!�Zŗ��Z �>��2� 4Iš�2Y?f��_	�2��j�r��㎄�)M=CH �Q���q�zg��%I 8.�,	F\a�B殿p1I9��.qo,��gh�0�cR����a���`ʝ̜�E�s�-����b����I��R
�j�4�d�T��D?����j����#(����g��b��}\�*��p�����3W|{�72މw	f�fsH����M�-V�Ge<�@�j�3IlNg�=~�	�;�ⷽ¨�O}�o�e*+�?.�ifj|�q-?�X�)9���
L�<̿�t�BX2��ҋf����un>� �� `�x�7[��9�ݽ����IAȏYY�( �:H��pf��i�K�p����jI/Ʊ�=Qbj���p��h���X�u4,��3� ����8(o�Z���Qg�LVgټ_�6�>Yܷn𙆜u���m���tE��C;�j��V�!��U6��t�����+��CO�;�8ڼu��g�|t({(�g���ڊ�s0��<�y�dZ��գ��*�������É�R�����_���p;:)��߹|�k��&0vz�Oa	��ȥوwUN+0�{�XO�8]vY�w���.�g���%鐻���~�	��#�r��<n����z�B>v�MP�GXW���Ԩx3�(��djeЏp���Q���̰����G���}�-���Y��4)��r"I(�υ�UcAST� �K��*����w�%.��]�_�A:����t���'��Ɂ%�S�Ba���~�v�`�xh> �uNmJ�w�u[6Ư�6~-�I�b�>����(��67���f2z�4:�̆���u4�'Lz�C!�y�ɽQ`���r8�>Mb�����v8ɓ���إm�2�o�L,}A����ϳ��e�_>Í�A?�o�ç溂MZ��5&��N��0��#L��|�o�����p���"q+Rl��4�&u��Tru�w�Xv�R5��Q����A�
g��I&�ҶRL���~�g5(���?��
� A��W�V�XEܻ���RB�}*� 3˨�"��#������bMFs@�X�Q,� �n*\!���-��-3pn=c۲ba�>{*&���
��X�X3�4��XSPh�����bUNY�p/��^ݲ�c7�(���5���ze�0�����UԤ�ފ���_�t����2R��ڟ��bN+�W�����NӺ>�����Ȟ���A��2(�PʗK��y@чq�Ӷ!c�M�K��/wM����r�!��ⷜbH;ݼ��Xo����܋y�%�G�˘~~�/5�p�j�Npg�<y@՞�P��`��7j4h��t4�(�Q��Gjt"�JO��7����ѫb0^��2��];,}"ASw@<��0���R�M1�Gn}�����A_���p�y����)�M�(W��i��6'��e]���7��뙠���8�&SX�G˖�7'c�a>�D���̴!YE�`���9�9Z�(�R�5�]�4��x��W[CyB,����ю�'D�Ӭ�ao)�V&�NQ�?����b�/��k�|16��85O�e�Iq���n���j6H�i$���~RG��]K�vB��Ű����S
i<��J�"{1j����k���p�xI�2�9�K9����u�r�q���l{/�_3�~�u��F��#�M��.r�l�����izϻ�{�+���Oܗ�M���@q�Z�^}�y�F��V�R�k^�"��p,�]�G0p�:��j)?#�8�q��H�璬^����)jYM�OjR�`�L̺���A�ٟqk��ߔs�����ŕX�@��psb];}����:c�I�Z�mV�aSd�Ǘ�~���S3�͌������ګ8���p3@L�8ί�^,k��h�����t�`��~�K�XYa��8����g:T��Z�4}��y<��"9��F�8�ƹP��߫c�V7��'��>F�o��<�§�^x[�T�d�%7�#�P�'�u�]��#X?�o,ٕ�٤Xn�N߳U��W�����b~hr�0�l��=xj��-lF��;7�/�1�����y��d�gd�P�eA���OJΔb�8|�3�b�ć5�O�s*�C@g�7(�ܦ�B��X�5�u�@��a X�0:��e`'n:#s���k�;Ѱ�����	�,%8�ba��C5>/;|���Ƀ����v
�Ɩl�%JY6\Z�D��C�{���<sJЈ$F2�����At�!��?����rڂd-J,�T��?d�]�ބ'i�{[@kF� IYZ}�Y��>UW��G������(���{�7�ҜT������p��LOXs+5��2�s��U�f��Yʄk�@ �����K�;8��ZY��b�cĚ���c~����O���k��Јy���n��D���ʷN[!՞�i5U��E3�=+� TW� 3f����� �U��N4�}����Â��~��,��A�:��t,R?�ƄV�L`>�������p����%�u��R�˥�ERz�QI'��-�> ��Tϖ��gBі�kT�� �M%�i��\���/�1�,��~�����iky�R�4<�Ps�A�6���X"�K�	��-ƒ?dy\�������v����0Pt�z.�N���wG�9�ϣ�8�H��o<�( �v�Ӭ�^̹ʎ�iUe��P�x&�ܧ��+�ǰ���pf�]�E
L-����E�''��P0���u{�8 0���L��1?������SФቔ=ʔk�,Q���Uԇ�L�$Wϭ�h�%֍w��<2-5����:N�]j�-ui\������D9���"�7����O��T�h��Q����;�1Uܝ1v��AΗ�U.V(OX����*M���Qbp�Z��Lr�>�SXb�!�7.��Z���D�����,�3��% �ڊRr�l_/_���*����W{�T���<W�=�r�t��O�pb�A~�J��c(T]��Z�r�d̨��D��A�4a~ _����SxG��D[]OtQ�ʷ���R^i��х�I�i(��vH�F�n]����S��=�{��O7:D�c����٩*�u_۔~aԁ�ވC��{������ ������6��B����n��4�!,00��u>�>�/](+r~K��˖%X�j�)�h���)� ��Wg���L�a{��.���r��h�f�{��M�X@?e�R���G��U1s�;�.����*2��9�_��!'%��
�b �_�����/�U 7F�H��N�8��ɸ ���BҾ@#�<8�7k�S�-�i*l������~��_�k�v`��c�x�R�"c�K!�I^�2��e�e~^囄���K'ڹ����<6r�d@�iܑ<*K����Fg������sA�L�'4.��k˨�*뫔_�5�m8FĖC�?�T��*���&�8�Yb�b�P2ϪөM�3g��~�H��^�bx��ǣ��s\
�S:�4D�w8p��J�IH��|�M,k!r%2{J��Z���m>O�7��o�z�>T�q�-p3楏�f���;�ae�>P��ƀ��Z�C���]x>r��_�0zO�1��!-~��� �)��վ\5Ya�','�����f1��.�5��f�$gDC�;�y��!���̞����o>s$�����VFw���1�	*[S�����~�.������`��}hQkH�6�^��"�}���E��8蒸@Q���O`��8P6�INW����=��7|$�w�(c�<��	��e~i7�����<5�T����\#�b�L�K�͛:C�CwnUP��o��롐#���yc�I�0�S���s^iLL4͹ i0���yCb�y
�]��l���+f��X�igk�K����\>g|��4`���$;���������;�6���0��7��X������Uwgc�B*k��[\Q"T�dcvG�i_
̶���8?��	M�"?Q�I��nB�;</�?D��a`X�a����PK?����Ղ;T�C������=���T�����C��KGk�'/����!�CR'�<`?ç�.�R@W̯F�-:�Y���:V	榃��]��Dz�v^8'���́і�Z��F8��F�qЧ���j�@��]{A9ЦL��"���*=֬�~�����~v��S�+'�����l���X�:��H_YY+�d+�� q�D�5f[@aU-���6R!~VQ	R��t�7��?��͹�SGR�����Z��w=ڃ�Z��!�ǂ��ƍrX�*�He[[��xS������x�y{0v�,��J�b���t��&��Y	:����&~�ȊzNxu�p1�}���zNL����q��v�������*	ICH7��`�yHR�f��� ���LhD�S(B=
�d��������C+=��@�<:�@O��>VC��Ex���u�M��M����ђL��p�⯽l�������@|g|2-[hI��O*� �ߥ�IN�M�{�.^I�y�h�Y�Ɩ7hW���":cCMK�Ilb�n�eңC�H�*/��V��籥��:��m�%t�֏�����Q���D��.3C��K��������iL� ���<H3�jYoNo�˽�C�GO��F9# C|�k�z��T/��2�hB^�
{Ѯƹ�+�߱��7��S�6'k(�8G�C�i4S�u�d�Êe��|HVǇ�����E!�3V`ُ$n�Ω-�:ɗ���KQU$rd��4�n;��A�\��jp���!�p�����l$49炽�g�1.������ΓwF ?�)
Q!f'��V�v���)!���� ���
�����׺�����M���r<^���Chۤ%��+��|n=Ԇ��] ���su���@2�罟y� �˕S}�N��eR��9�&�ˣ�L?���,ڎ�ڀ������O�2W�a�%��R9`�\"#(���6��O�������'�;"-�+k�B9\tDR�n�P[��r!��pE%>c�~��ㇹh�l!�v՜^�pT��؎I_���e�ES��=�`���GF��[hBv�Et���~}h��xL���v
�
�;��Q]�H�S�+Ő���q8�r����Bn����(��
�h�'l���L1����ue:�t`���}N����uy #��֭��;���m,�ֽA��:eF��ܿ,�"%�=nI���e�;�;�BB��##^�}b�[�'�w9��Ɏͱ�H��ə]�5t$��S��UbP-k���$��{{q� � ���p%	dp���'�߰s�%)0�{�M�wovW%�h �����&}է�N�"�	��ӷ�ŉY<�N����9+��`�93��6~��j4&��Jl�6ꤞ�K�\�^8����&���G�Ҡ�"�B'���	g���փ�@
 ӊ&�c� �8���lE�6�q:��>!w����\ �j�Q��v-���(��~ |8;L�-���9�|U��\����ˮ{�q$e�CYĵK9�z�_����e=�,(���k�	��Qr_yo9�j���^�_N2�J3/w֗1P���Mb�k��#K��G�� x���ٖ�̣Di�jz�_��*���!.�I�s�?�t$�ˤ>d��[{S�qk��i��4�Î68�u���r�|��28�v��L3?�uؘ��$��|r��bR�y����l/ge|leId���uP��(��7�@4�
��y�v�7[���}`|�! �� ��m��\Sq��A�O�/��ߤ�+q�� H )<qa�FMV��S�#� =�K+�?^�����6�"
�3QK�d�2�S�+:� 6���G=��⥉���O*z,�)y��޾�ǈ\0���\�Ӌc�A#�@{mњd���ߴ{ =�z��B����0;��)}	��!ޚGv]���<�3�S�ҟvm@�Ƕ
S\gqJ�v0և��g�,�a��s��U�[@�,����b�)��]�}�]�1C���ۣ>�����ul�mt�3s&w��q�� /�a����X�F]�"�r��J��!�?cեNu��� �euk�H1�L�9�k�T��j厕�/l?��v`ESc�5ץ�@�l>]ðw|~S���w��~/�X��p�\I���3RSܻ��$3�H�_q�o|��W}w0�5:VOr�ު	����3E"CL�"A�fo�48��4b�B��-sJ2k�&��hb�#�'���S�Nwj<��9�`��X��,���g2,�qA�-�R���xIn?�Wg}'�h�c=���~	���@3u��/��]�`o��2���́D�Q7���V����w�O��1������s
s�eߋK��b׸��&DG7��-?m�����y��58��_h�2f�(�l�N)�o텉_['��/ ��������jo;Wؘ��N�
"��vT1Du�B��/�6�fs�&�pl�>�A�"���{}yi��R\-A��h����~�6��Ԅ�V��b��T"�������)¡�śC�]ԅ��n��Н�d�ɽ��-��/�b%�2�����ם�?�9���Y�>n�<���ƠwEOk�1}A��P% }����\ລ&�%�_�i4�̧�����.�,��b�,K��J�$��A,��o`���DЅ�}WO(�����Y>,;���H�"�-���zh(F�r����������&�,�|�ķB^QW�ۻt�@�pIZ֖f��s�J(��v&���q��h9X�K��l'g�^����"T��80�wz�;Ujj�V2�@�n��'̪c�;Uꎽ�m��v^`�bV/T��=F� �%!�y�!�?H0�ռ�tؖ��m3�f�?�N5��aUފB���ɳ��)\���� p��N��_׫��s����X]��`�g�f�&*ah�:��[�2鎧�����k�����Nh5��o=��'�bk��i��-�t�0"Sٷ^M���zcO:�H��;5!� ��u?<�O�T`v��h��@����7er�I�`9����<1\��{���Ὑĵ�m�_��yk3p��8��+<=�r��/f�(,��щ�yu�n��nT����J:��#�Al�a�����
RW,ۙ�wkW�)j6��u�ƌ��4���Ra�F
J��ߗ��ɜ�~�Q�_�@R�M�B�ժ.�N�r���^Sa�3�%N���4�������c�`����䊌����^$e�\�*��$A��] �`��y���W�/CH`�*Q�$d��z�~!��)�Mx��؆�Gc��ǩ��7�}��4�"�%�:9@�=G���'��?pd�0�%�Td�)['���� 6|<[IǙ�
pd����z�w/��x΃��;Չ����Ƃ��㿚dl
����.��Pz�`bzFFZ���I�������4��[6�R	P.2pa���u�pꀅL��V�材'�d���p���I	�� q�[]�������LR����W����3M��w�G�T�a��61m.�������ݐz�'�N����@�V�AG&�3��H���(�U�9tiG$�EU �<��B��)�R2Qy�C����3�mY�e�If3��L&�0�0�.���0n��Vfu�G��{]f��[����}3��C�|)�(�-~�'-s�_#S+dM�ǴY��D���,_.���&-�e�v�gB�*,���O�9��e�K�Nt;@�3t�H�"��dآM�g����ꮿ���Lk�o��	�A��l*{5v\=Y`��ʻ��M�~P�:XN��2���u� �(� ���/瞋E+alWBd��g���vE}L"%+����o�#Kp�J����]ʤ�0��ƅ�{w%x����������%���`UQAcE�]�g��kb��W+i�	[�QJʏ�4�����1J�b�3{I�^Jz1?%�K{�+�[@fN�=�o&���"�YE��5��7��S&�|�5sob�����!�ўi�Ӿq2���2!�0P��p��M�H�KC�V\MM-�J���C��rHl����|#�Ip%������u�H^8�#۲��M�'2N��O�G�B���kE�:1��MN��:t@�����7d���\�2�(/���E]_q�E��8��v�?�^R�[骵JWSYl��(�Grw�B?T�P�ѧX�
�%0���;B�]�v��F!�'Ȭn�8���3��Py/����1�F�@�9[�3�D�Te/�!"�Cm�nЧz=�#ĘƦ���e�j ��y/mӿ�IL�v����Z�����;d�!��9.��SL�� |]*3-�H�����	�3��:w�e��ҟ�À5FXTJ��9�;CRb'I��z����`�}��������:��k�F��<0|��C`�Z��!ʼȬ[�*04����f�i�M�"�̼��pd��-�J����h�qVd��n!��T�<,�H��-�. ����s�H�c�L1����cE�{pC��E��n�C=}��	�r���z��z\����i�w�2#�a�Xs���#z�}�U-�%�����E�7���Z�˺�J�g��୙]�t�l�.v��B]��H�`��/;�(�i�':K��[��>`/v�Y�J�}WS�G��}��>��9E��ͿsXu���dU崶;e0H�4) �&]�'r���=���4d�W�2Q��d{�Km���Vx�*��:�ʽ0ӑPj*��z������W�/P;�-�k�,$������m��W�1����8>�Cg��e:G���f��B�%�ܒ��렀4�/(�w�l[[-��}E�p��&d����POպqm�#��z6V.�7i۪�rn�K����x4�ꢗ68�|R.�c������4J36�V+i�ݑK*ұ�U���Ȳ1��H��0�����_� ղ:Pj��Q��ފh?��v�_�c�"��6[x�W�U\Q���,uP<R*�na�p��u�P����C}p�$B����l������$p�"J��q[,ѵ��Sl���S�q��� $��d#3�89V��kݵ���0q�X�_2�;�r�t�6⏧��C���Tk�~���V��s�z�^�f��Mp~QR��(nf�#��n5��͡6?��~�� 8�)?��eN�O���(*Z�Ii��0,��Hnah��S�̥���>\��]�?x�m8�_�͆���I��[̒�ȧ�E"�����ҚJH_Z��6/����J��� ��r����� u��w���bIN$�u׍��e��u^����[���#�5���n�`Eڌ�=�v�F��we�]����ې�Ѓ�X��->ʜy��B��]��g)Q��C�U|4�s��U�'js����ej����6oƶKH�Ax\������)���,�9�<�6dl��� ȹku����'�����	�6fj�8��Q����7�����>��W*T+%��7K�8�רe���e��T0�4�:v��9i@���]!-�B(�x� ږsTk�O�V�,l�Y���7_�K��w6�*��r@RA(�����3�8.SC�T�Bo���:���r�#�E�h���h�^P��y ��0���gGG�ē��	���!q?����pU��c�ܯB*�*W��6�E�6�ߎ��u� W��4+�L.�N���kXC��f�k5��m~N����<H�/[�A_$qo�F>���w�:`σ�Oa]R��TC�g�N��.i�s�R�:�b����ր�6���8�څI�Б���c��B��c7=����zt���R�j;21��ƃJ�Ƿ�D1���@!�[ '�p����!�'�3M�B�5W�jU��:�fݗ�;�X mf�.�^T�P�ܵ���N]���o$����|�LD�L��V>و9|v�ǁ0�&픦�b"lƦ��	�Y:�5M����9���41��f)Q�[y5�g"
�k�'\
�T�yD�IAlT�ܕ%�焢�"|�}mC&+Nm��m�u�}�F��_�Y�wf@�\<�DZ&޶�*J�I�.�a�Iq�|[Ht��щ�8���@�Mʹ:����\?��a��$��u;d�;����(��w���0K Ӳ��!��b.���/�A�w%�t�	�ez�7��O��b����/�&N�$�h���/6�I��n�VZu��t�[�a�(��4�}����`���W_�w'5�l���й���e1���@D���O�kn��Xx��^2�7;-���E{�H08>�h?p~�^�[L���h
@W��N�oT�=�S�/�CӦ��ے�*G��Wx���ݪo����=����:~J
t��T�2����c6�j�X#ڢٔ_w%D	�o;���Pw�@��p:s�^Q�Duћǚ���[.�f4�O�e�fD��S9�N�'� �Pᴌbӹ�ߧ=�N���zI_�1A� ��W�g�"�v�>G��0U��*_c�z�٬����9d3�[x	8f���|�䠾�~C%��PޟEqn]�"�����Od[۞����IS��a͞�?�����D �ƾ�V��YS�-�gQkg1����h���2�9�A��& �k^�ΪS�ziD;-g�
\�Ll�8��Cwd��-B�ΟgM���u�U5m�I5��屐%��]w�l7z:h�P�x�x~��n�R��x18�1Ƈ>�F`��+��_l���/i(#X"^/��肌�~���c̚]6x�q�,��5|u� �Q<P��p�F��dG��&��y$l�ⲡ�vyDKÔ�l�"��^1�:E^�p;��	���x�}������� �<ƺ7�h�[O'յO������{���G;�O]��pp-��[<�YT�
;�`�A�+����*�򕭍`�O��l����/�ft��r�"j������y�<�6/�-?�\_����_r��noݠ��r�������K�j���.I1���da�}���m��[h���&`�M�a��G��r&s�w��p�e�+������#���m4<���eA�m;T�?o�#��tt4�������zT�+��b���&3����"-[�����܁B��@���wZ��4x;���hZ�x#qZ�RA&�*�H���bf���"4�P_�j����p'��3��Q|h۹�CͳC�������.���?�����C�^�v�Te���z�d� �_�G�#rs��0<����`��3��0r쁮k'�vShG�[�J(���o�A�zr�&�D����N�P�Oը�$3#�� '�<Ϗ�Z/��=IW�)2�U\�邮�:��]�$�,�`ad����*�ˋ6�
8T���׮�B���Ia�#�D(|�ӹA�5$�����!L��uyŇN�ى�R9/���g�����¸�?�|K�ۂ/�D�hK�J�FN�����]JQ��B�v2�_�� 5h��7 ��-�ˤd�bI����\�H��2��*:hͯ[$�W�D"�L�{���^;%2hK �x 
���e�[����h���Ea"1�2%�c�gP���)rB1����:A5�P1�5�>�ؒ��*�͢zE`�˼G��`�����X;H\ʙ�����4d�%(KHA =!�s(�/�H;�%��a��JM4`�.�?Ԗ|}ظ��b<gyX>��eIX�0�1����Jd����H�w�g7F�_��t/���7
*_�(��3]����q��o�ѽ����lnB�b�)2z_��$��*�<�N�Wg�䓯5v���[��Ƕ�?tsL*��؄}�ds��:u��-i�҅����1�`���"��^E:�*�V}^��t���~�촋b>���ǯྈz�۟�w�%Ȗ%K҃z��cj�`s�0i���܎,/S:�"��F���M�U�Z�x���L�R��\.4^V��h��Kf/�悛��y� a<HN�dnm�8'*���k5�Ω����n�	�c{��v0u��xH:��,Ƃ��] �_'Y�I��<��ɾ�!i�0����j2�C�����y�����us�*h?�C��y��0%�"�޶O����'�?|�m�*�3C��G�?�������'b|���Pa���ϳ@]�,��X��j:�1�B�^)�&y��4�2�fi�H��xJ��s��b:��iw)��
�\E������M�j��Eu��p�u���>�ʓ5��yyM�5|X:���F�j���V�8�M��4NF��Q��aH���v�jA��p2T���9+G�GUQ� H�Κ;�u�9�h���z�r�p}��Z=�[��P�gil��Z沓�z�X�K�;d����U�Vv����d9�u�f����?����r�����M�7�������kߊ��|�2�,��˺��T��D���'T��g�����͖n(�%{�O�:�A�@�@��H����7�7��T=�(�Y���}�Q�[��*�M{���Q8�Q��'E�E�(
a�U2�Zc�������F�+��"��T�Ay��9�|�ߪ�r�e]>qJT�!�7
%�?��:��� �.މl����ΕV��Տ�M� ��>��L���G5��(�d'�}��H����,�5+q�7�m�/�8�5�ysX������5�rm^�Sm���O9��s7}�"�tK��~B�!����w� �����9)g��5oL4�
�.�?�f~��m��6n�[�wDI�q�$'���uZPN���ëb�kh�c�v������I^��ZM��D��*�)��1狿���M�jzT�mN{;ͣ��_�㑮����e�s��{��2kL����"�|�-.��F�+���Of�f�C	>SY`��nvesa����ē}/��3e%)��a��Sg&�O����_����QdZY�@�P�y�?���(��]��KH��ҋ)���D�(�Nm�ǲf ����~������Y�	���c���m1����P��Ԗ�{�^e�<cQ��a�����#�*.7dZ�_ݻ(R�P*�4�k�b���	/���dW��z�9R�vU%�s�\�z~b�~.���"Ҙ�D���r��D���0��o��~z���������7�Α�Nx�|��!
���Y�-AYh����{���]L�Dףf�B��c�]#�9�ou�\��W��I ��K7/9�(8�Yd=����r��9�m�S21�!(>g}~U��ɶs��!~(�ޖ,������ѩ��7�5��M�O��3������
Hd�uF`�Jy�pֽ�Q���@-0�ȵM~���l��_��U�"�p�J�/�C�He%Q-J+�e����n�?�8"�� g&�p��
�ǿ�v���I����,�8�<&8l�,�;�Ϗن�T6߉�޵��\6���wn� 7�(��Uw�W��>{j�*�\�󑡡Mo4��D"8'�����jJ�o��%K[���_�9�K6y�g��2��9���������D���*�ӓt��hG:qe��a��O���ə�$X�&u���G[��hӾq��؎��6���pKh�4]خ�\~�K_W��q6�1^���l����+�"��I92�;�;C��F~�ϵJi�m�igD|�]��ģu�t*��]�|��k���I��A�b��&���	�(�x"�v��Ƈ�4L�g4�j��]T��b��� 	�H�=�����ͺ������6L����q�x{�̉YJ�[,������_����lzNشK\I&���!,�0۞��MI@ l�h8�9�D��'�9�%��w��}w��%��cF��+)^=5�3\���˨@h��#В��0�<��/������R�)h�9�����NJ�_���B:�̴��E��r=;rP���̒�'?8b�4�i�zR��@O���<۾���M6�P"��'�ܭ����k�9�j�
U9�^�^Ͼ�^�6��V���������|i�>74�ɤ9fd�玽���h =s	E��Om������UTڬI�*G�iR�t��y
d���NFX��J%J���3BtcjT�_O�"� �|mj@,��k�ÆZ$|�	�V������r���=�h��[w�6�����V*n�ed]��� ��f��E����,%��1�
�f��ɰԐ��ֽy棿�t4�#�%�W�褟�����n��Ӝ�:>�<k̖9�B����.[3��m�=K�ڃ�)���mg��������~؊�_�@�B��m�x�<�["h$���.:�GE��w��� Z����.[w?�'4q��KM�/d���H]�BV��Qx������ad��ut� �r����c�\8�� *����s�}_ԦN;W��it�ބr�q�?^�������݅��V��Q���dղ�U��G��~ᴠߢ@c�j��6]�]ǹY�;@ʕG�6��TVj�9ѽ������S�� +�����=̢�N������GhhS�=z��k�S���&`@� N��q �[Q�T��Q~�f��\G߹���\�:�:Ҵq㮈����V�㣱*5O��i+%��o�"���P�_XV�3�ݣ�E�8_\m��s}
uc�R����C��B��B(,�g�v�*�|�cS ���H�|e�HF̎�Xȭ1�:=�������N�w��`�>i#:H$#�+zɑ�[�{��y��=��{-������B��R�\
� � <�K�)5_n�+��MM�G�V��'e�}{�恚� =���H�\�㯾\R��lEE?���+�Ίc[����N�+�_=c���T��H�[���}+ރ+�uN��nȃ�����G�+k_&�(h����ܡ��o��#��Er�{�d��{�����˷s��|����a�$X~���a�|兾��Q�IcgӃ��,����3���������1b-��E����8<� 48�y�������8�m,�f��:各�m���a�׌K�pT�b�L��n+m#�4�_0`1��z�j�N����hAЏ��Lc)5g��7�-y��4�n���� �L%{�a��P{o����@�.3���/�4�>����XX$��ʍ�:����u����㯿���ZF�Ɲ(�PU���salx=�(��7pw�F:>����=��U��t32S��#��˵G�bX�0�3�kաKWYz��ѧ�@��%�X�y��8VX%��%4M��	R0-n8�2ұ�x�!|������:V4ʱm��1[��1����ɤ!ҳE:w����ϸ�1��V�C��*kn����O�����8-b���\[�B�TZ\@�HO���\)��r�ծ=F��J��+�07[g�T�L���� H�8�J�1�⁗7]� ו	%# vx|�q�J�+ܨ!/f<���T�2{x^�TZ�dA[����,_�NG=��0nͶn�`�M�iߵ��ȋ<�$F'T!x�8����3N(k���ȅ"��Ǫi�"����N7��)4W�����/�*���o���D�����(�F.U��G����0���O���K8!
ϕ�2��^GJ��u�4���)Y�L>�l���VnЎ�nG�o��=�}��0󇖒��i�/�g��U�O�&��^�3-��J[S��l����V7�H֌T6�a 0�z��m�^#SI仈rǥ�Ka1��w����ye-Hu� ��Rsa7$n���̲`jI������dw�벸�$]`H�/�X�ĈC�nJKf���{�B ��j�7�j���2Jt7>��̚=L��	�4���jۚ�4W��1�L,��{B4g��t#bB�`)��@�ݸ	�Q�tA��ڙ���l�|JKO�Ɵ��^g�A�n���vџ�Xv�?�K���S�-ic�֮�v S��J1қ�����x�?ΈQ��Z�.��ɤ�m�C0-&3�J��Mf&�����D��KH��6� ���ϳ��mK\�\K/s�a�a,/��ö��ç$9�LE63�d�O�$6l��uPV�kl{�e ��}g���h�� М/��a��ؓ��1;شi-��9�}���F�M|IYh܄�[���b�l�5�P��
/޳���h�1�n�R*�,lb�#,��5 ��ySa�]"��Z�=�?�*m$5�̔���BM`M��&>����ч��!��1�V��͝j���M���UI�}<�1���6Re���w�E�o��k�����9�Hq֎~�]io����2Ts���Qd���s��Lb�q�o�($dIe�+�g�"�{��X�K 1{�a��g��lZ[����iȫe�j��c�"�Zy5!%3��a��?O��z���nN���4�x6;Ͱ��!�g.I׻�(���9�?Pɺk?��%t�_9A�c�y�2\._C�e��6�uXX���뎦&�n�sUu:�iW��?g��c�j5��C���;V���|s���	u'B���UJ&���"�����_<�#Ld_� ��aKѾ35K���O��c,��0`�7@����7Qs�uc��U��B�7S�b;ix�E`��e���/9��ض�ȩR����Aط�ٵGbk]5�@S��c�e�,痞sAI�
�D4�4L[qQ�*)��J�[��e��BP�]%��m�%��*�x��TMţ8��!�����bH�.m��Y��J� \���YA��#�;�@F�M߻�?��p�7���m+3Y������/04XR�H[`48���q�4I��M^�������&�W?�$"yI�GE�q���	�z�R�tl#&�b���������6�����A"Aė�v�"���_9���շ��m�����U������
�����������β���$��Q���:䯊��q����31b����r������ΑMw�3a��D�_�Z�ߤ=۲v�`�G�r:m~�Xr�,�|�Tڡ#�S� �e��ǁ@-[�WSx3G,�@j{��621%�2S���Бq��l@��D_buI�#�)
^�ð�H��^9�/6��x����J���%�pC�2ν�e�R�0�+�Eȥ�K�0������i�.tf���u���l~I��p�ulY#�қO��]���Lj��������r��Ա>�E�ߐnI�K��"��4D6\��P�v+�˗��򳃹�F7�]���+�Cꉆ�a�X���
b�T��֬�i���I�_�x�Omd�ṓJ��?ox<���n��?�6p��$U�d}����o~�Z0��H%ѯ]��,�PR>�)~��,�Ē�[��:Q	�z��΃��/�~��W|�+�ǚ�(᳍�t�:�v���}b��2�"���e���:;��;������*������d��i�<$
ǭ��(^P��i�('�٤��qIt܂�KK�օ��x,�#��"�t��X���.ߨOZ�`�$a�z�0�/�/%�lPn�wx|��x���:�ֲ6b;�'Eh�Z�ld�'r��2��/� ~��ug�EtQ��J�9kgy5B����9;޲��&�����W	��n���I��e1H$Cj2����ШAʟ�(��Ɏ�hc��4Hn�H���5��Mm��X-�|H��!1���!�s����C�x�~y�v�µH9�:��2���c��0w>Դ�).׆��DSC9���`8��l����p� �;���<��V�8&iX�;"��E9����Ch����Sγ��~�Y�]�Y����-�vO����v��QA\:����Lڿ�p4sX�t�ҡts�2����5d B��5FD bu��;��.�q���'�QRH����Z����)�������m̙����LK�KS���� `���s��V�	t�N;F�z.���0g̛df�t���
�=*d �!@��M�I���bٱ�<)y�Ut�-
*Lڒ���������
J����n������~�	o���C�k�y��8P� v�w�Zu�"+��TtO�}m(yo91���V1~�e�D�E�j��0���}��U��!�fNsϡ�s�1���'�ʞ�����y��h��Ru�XSg�x��q+�	SWXZ�z/�oi��
������5�'�=�����c/?o��U���3��uj�F!��F���˹���qAy���t�&�X��~�Ǔ�M8ٿ��V�D��`���������~�Pc-{�L���DxSI�QUԋi4o�֡^$2�����@�3�A~��.�m2SjB������C�(ۋP0���/PV�`X���)Yi&�,�Y�R�}`����7tm@Z� G]]}�캨�lsP%�>�;�Z"�D�U�ό������o�ņ{��x`�ܒ���q����L��=`
�&iVy_<9���I�*y���I���Ox?���gD�jܳ�W��Ǵ��]].D;��^��	�JW�-��L]Mª^X�ݣz�i�����u��z4�Ӗ4��PrΚ.3l��Εv��v2(߃Y��L�'u��:���KSTUTG���(�.��e������xq��u):jP�d5�9�XxՀ
�N�k4WA{T4k�����A�C�b���f4ɉc�۾�G�����S�#��VO�p��Y<�o��yy���ٱ5v��Ku�������NZ��=��Nӿ�x��������+��V�'�\���I�L��m[�0"#����B�GB�g���E��2��&<X��dn�Fg�i.N��L�� ���'�}1�Uf���*�����ܻ�m���ɮc��H������T�>[�[�{�5'܅�X�MB�f�rB'S��дH�����f?����bo�@,x��vp?M�	���Gܜ��Kh���p�)��AWnv�}��!��ԽI� \%?�*{#$��
T4���N�5��ຐ?co�h$$�sԭ����0��3�2C��\��p��+r����f�%i���URD_���zoO�tA���G�x#��=�H3b{�睚�� �����Rs�=�֝�p�C����� ��E�u���oWi�V4�U���3��*3�ɖ���F��d�O�����J�-S�a���^`��-��:�\�f�����w��h������.9�!e�% ��U���|�����9���FA�SY� ����M��ߪ��ׯa����&���R���2Mwp'���1n�TA{	�:`�rw7�[6��N��J^Ɏ����-�rB�i�$�9��G�/#��2���LLx�^�����q�?��A�[��XK��C�����+��_��?$�F��n7��'̞��>	gJ8q��q��#�l�ˣ��Ԛ�{�Gd��mq	}7��y�3q�D�
i��z|���\:' yE�����FjlK�x,t�ꛃE�<D����/{�E�ep1��1�IB���%��u<�"��l)��@��.1�$���p���ё�l��G[?��g���<IT�#��]i8B�9Өr�E�n���*IF>�~&�PnX~�7Vc"?��1A�囫�tʧ�k�����5���ս�yp��]}���_r�*�X���2�c~�O��l��4_7&��k[����V�F��M�ۣ*��ns�:����>L�^VF�Ƨ�*td�#+"�߹����R �3.Ը��Yد@�u���P1���Z�92���9��a�I��g�X�Ь��9��x(�`��s����>h�J�B�оc���}�{#�y�A�T����f�0�ޢz�8F��
E��J%�:|��+u\���ؒr�3LL��r�����;$<n�<�wa���.� ]��g��?ӛ&��@�q�?�?/���P-�T�t�hJ�L�8��RE�v��Ćrؒ?M����W��� �Tzkf0wyF���*R�/��dB*�5�7����s]^�6����
æ���c��Fiҍ�n���BxV�Oy�ejm�����Ł��	9w�+@��E��Jz�� Dç|�Ų��C���EN\c#��
�fwޑ/w��@{@	
&]� $:~�KO=h��D��k0���G:�`�Nf����m>�۴�K,��gP��>:�,��>��\l����B����N5$>�q%�H
RM�C~�d5%�*,�f
��(-�l�7��}hH7�e���#/���s��%� �0���B��  ��W�����%\�7�Y�����$���]$�X�+d��Z��*���neb�2׆v2�>wy�t�,�d���d�Jy������sv��5�@M��F�=�F7ׁ.Ȉ9���KE�`L�P�w�Z�d�e{� u�lcr�b�=��_�-2F�<�Ё,���P���N%�X0�ԭ+!�����pR���M`�
�]�[c1b
�@���eQQ���\���d�[VK���ݡ�B��H���+g�	���%5�l�v���3��ig������ۥX����[e�)��y]�`
�<�����K)o�6�N}�&���`��������G3ϯ�O�R"ZhV�w��/�
ޓ�2S[.��/��D(z쎸7�JH�~�)g 
�/j��Ic�����u�r-��Է�6<(�1!\@3�졲��o�q��?��2N�����(!���f�v�3�Q<�{�ǟ3���5�-�{D`X���m�<r��TWGH�Zn��Ea�}ЉH`}�yۘk�H�2��`���`|����!�Wl�Z�v.�kt:�	�.{����R
��2����%/��91�M7����}7Ͳ�׏�Ǚ�% ��q|m))�.����w#vޫ��UJw��Q/^���K�D7t+��Z+��淐
�l{~-DA)ЙuR_������D�>"�=+ר!��^0�P�VF����o��HOE>���kJ�r+-ǂ`'�B�k�DFf _�YKڗb�|=���Ɣy]�a�����/aK�K��� ރS�*=eG��}�_E�E_�Y&��Vө���<-��[B��Qr�k^;�6kg֚��/K�� 5Kb>�����->�V�7}v�9���滰�X���]!`�%� -�#�ج��ub�q.�Ӹg6rE?v�$v���b��+�I��ǌ�'�aY�D#Aeu�xA>�2��Lq�/d��4�#����X.S��zm�;�H5�ܡ��8wu���<@���/�7�Z�^�2WKIO%��ψ\2��5_D�O=&6D9]G�E�V:ѝ��(���o
|��8��^=���?�-��P�W����}����D��Glx_��'h#�ux�*Vz��%j�aK�}��f����c)o?A ��x1����� �Z6�d����c>�	65x�ٖ�w.2>!r�m'b�a��֚J��6�9wI]���lY�B�&b#"�o����X�ᐍ�@�\���r�#-�9�]#��i���9M���9���AZ����: <����}d͐��^��h�܋uℴ�ȟ�t�a��w����&�C��c݈s�H��&B�gv�M-q�Q�n�)���iCp��Z�C�+�oCs���6�H`K�Ĵ-�u�ܹ�\)qS��.���<�[���su�G9p�Q%�,�!N�du��	����d����{���j��x*W��	\d&f�Vp'��c՝�KU�߈� ���
�%@����}.���n�$� E�N}c�a�~���E�M�,Bݜh�m�-�Ȇ��V|���^'_+�W����Y�lڥte;��G���X��f�s��)��U��n����S��xz�w���+]��%�ckGn�W\6�J�neh`D���v�_����Fe�(����O�d>�ht�tTk2��J���P�	�x����p�5��嵽��|ω�� �#K��ͅ� '�ly���>�����4�5���O�w�Ф�{(����d� �ch���8�zԎ.9{_�����gkiZ������[�<dy��㱀�X�@vl�fL�������_�I��ŗ�G�5�OP@�L(�;���тB�%�݌7_�������?�#@S��W�2��l&��el�a�G�Z�y0�Z��z����"�O�HXyѫ�h�zǬ�j�^'S��O�j\�� v�e�CQֿM���F��x"%Kx���L���z1�czGt���Q��B�$8<!]��*�I�-�՛t�yلz��5�	��%j1eZs�|��F��3m,���ښ�ࡏ� {��/�&']PBPב@�pp�ۻu��v�%��X���~Z�Ǐ���nr��^�F���0���%�$���V�J�Ȟ=%p=�s��Q>i�G�y�*����o��%J+�-+/���?z�];�p	)z�@�$�o�,J�=�Tx���'�?�J1矱�r<FB��(Q�M?��'��3o���|�Z(��.7����)eT��i�Đ��)�Α��������<��W�-گ�%=տL�鑣m=�!�s�o�=��Ck��QT���քBmt.�a���w�8J4���p�.7�e�I<�*1�y1)qH�#-JF�D�aH�Vib�Gu*��j��܀��7 �� ���i���md�/�g߼�o�[I����@�+O�Q���5������'�q9S�)�T�0��u��:Z�.�bDN�o
E�?q����4�Q.��:�в���a,"s��.������}
��GKS���C���a	��?�Xɍ?�J?���m-��Hq�빗�c7�q��+X �K"�m�f�=a�����1����.`�Jq0�ěR�������т{���#E8N���Ƶ��˘]U��#�Tj����i��_O4m��Mb:!�2��=��V3���ծ��e��>t�@J��a`���R����QL\���B M�X^ȼCp�4�*sӤ�O�������|r"{�Fv�Y��k����>�Z�!Y$�3 �����k��D�s��r� .��Bʉ��Z>s�Kĥ8NS�ͺ� ����0��=i�z�DE��o�P�|�F�nX��H��]r�y$`��XYA6{�ŴP�bF�䳔�x��.�tu�Ag֔���϶����\�R�5�����x�#�ǽߍ��q��%7��������_ɹ(�W]a��GY�������rS���Xx��Qw =m��^�_>h�b�&�KP�֨jo�g��lӲ�����)|�?��xw݋Y,�гРc�[�Cp�5��9�ݐ�:XXG^!/���ZHăרmo�7ݝW:8�i�t�v �>囨�5 2���3ꝡϘ�Z���ZD���!�	0:B|{LSoM�KD�f�"O�Q�̈́�^E�?���4$#���뽍��J���-�C�N66���2�a�y�$��Q�ֲ�Z�Q4-WD9L(UE�4�bN��$z/�8�%~G��]�i�"�XҪ^��/t��>7�n0�Fa���p�M��`�7|CуUw"�yA��K'���$�בlƀ�"�G������(=>
��>$Q�%b�j*x7��Z�5%�&��ɮ����R}K�B{R�u9Fm>�<qA4:#L��P,BxH�b���P�O�C�a����]R�c''�;�.���Ŝ�I+��`6�"=�VE�|�7�%���]�;���������}Sį�ç�s��4����S�|���T]�b����P֢T@�6�xW��g���:�s�l��|��|��O�8�(uJd{ږ�k�@�P��YZM>�U�<"�����lJ�mA%;p)=�҂gR]T�3'8.���l$��C�3,V�@�0�p-�"��ao�o~h�C���� %����ԟ�k��W��T-�k�\*�d�Fz�p�w����%�*w�P���c��|��H5�]^�:`3ql�Ⱥ��H���)>E�N:����*Je�(J:�����_n�
s��;g,v���=r�P��.q��Փ|]��a3	��r��G-��TK�Zލ�+Z�Z�t�����ylZ`,�%T��Й�*�9��H���k.��!�)�3�������\���	A-��ȑ��:!g����TH-wÚ�+���?�r�B~�(�\:�/6Og�@��m��1��zW�x@:�� �DfB67��"�@�P
�X��k�ʽ�-��	X�.rOf*��:���M!U&.����iJo?�����Ȟ��~��BЗd��tztu���&&�H�WƚW�ՀqV��pN�Sͷ <�8��Q�<� ��Y�%굃��v��^�/R���<X\�A"���G($����w�5(����к�?��|��H�u�<"x�=���٠���M�r���l�ϊ2����P�W� S�k33Z1L�W�n
e0'�� �,kp�����7����@H$�_�k)�(qX)6��S���1��O����{�Y��t�v���U��]��\,��mUT$_Dk�����E�D�<�.��Vެh[��L�R�b�i��܅��B�*j|kÎ$Y�2�cX�&��%�{f=>�s��WN�Nb,���3�f5:���j~�;�Ѓ���2 My.JX���h}��վ���ct��F5�[��p�������a�/�K�䱏�f��e�Sp�Z:���Y�sp;��VN�ݷ9�,�XA6��v�{��!�zS����8�c�V��4W�%��1��"ӷJD�������O�if��=����ܤ|�\��}y1�2XF$C������N�$�2���H�"e���Λ��w'Hc��qM2T�e0Wr�����͖����<.��L����ni[��K;�Pn=��FD����.Ň]��Σ`���yf?����lfI���Z��Z�ڿ^��Y@-�0G��Vp��U���m��X�������P���k�/���M!��:�:NfL��N�i��,b�v]�E��<����F���J�F4���Na3��d�~����vJ�[G�2��H��
t�Yb����H8M?��t�Mk���Y$�~lG�O��5[ëP7R�p���7���e}zLWep�I-�����&�5]����]&�Ҋ�0��:�����~)vgVW���ZI��V���i\);�HO:�PX{�g���qU+v�i�������;����(�%4�sh���J�U����S�P��{R��h4����B���6%�&���Żs�K:[f�b�O�Y���[ٳ,IF��{���ڜ"�$gX�Ԉ<��Ѕ2�j$u���9�ct �C���h����=���<��Q��gqO��Sx��D���+��FgtW�'l�	=�Xݖ�ͧS���wB�rf��ݎ~�k
�	����"cD\z�I�"���ǌ\�鱕	����3��l����L8������C����F���*,8DJ��r�j�N>�DX����u�\��1��=�R��4\ƼW
�
3����Dl�+"<��/(G��cv�C-a�M�%���N����[/Y������Io �돃ݞ�n�u��X�F�Abn%��R�=�FW4�V��2�%����R�����ϚC�R�����]��U�.��%5�RJ���� �w��I�e�f�o����0:��+#����ȁW!&�^K���MG2�+X�@(B����しSV��i+�&Jk�`<�IC�tt���$&ك�%���Jɚ�(09e��k K�5�|x�
�l}�����G�Ak�Ֆ��U��<�|��NW��HƇ���k���JK��ө���Z�9�`˽U��f�w`���q�-
 �^�}0;s:"eW��T�L������~:xD5S
�X�#]��CP3bU5�k�(����绔^}����w�Ϻ��ɠ��$��T��>?[Hk�d�����������W�#��Fn��X�?e�7� (�)=��)X"��W\l$�cH�fϬ���\���տ��,U:�T^A�7A_+���K�'c�F�Y-�9�����/X%;����(S��,+֭m�A�Ǔ�����47��� >��擬X���M05������v����I��[�ۡ��X�����Q��_�M�܀]h��ϯZ�6Qb�z'��G?a�������'*
7�)��a����[�`H�|j��u��\�[���a�:&�.𓚗��v�Օ>�Q�,w{�֒����s�i�ͣ�]�Dd�g���T��I<8l+�\1�}�9V�v��'~g�" 5�_��]BYi�@pD.P�;�"QV�,�����o��Hi�+br7"U�
��^���g5g=�FbpO?9ԖCX����/�#�Ӡ�o��?�4�y=�B%N3�ׂ�_�"�F���/ͬ0���oN��>��Nx	k<�X��pH-P~�ꢖ����r�!��1�3�2M���	������4dǸ��/SOȽC�R�l`M<	ǕN�f�9 ���)qp��Awg�J���1¾�����R�4E�+\/SW�U'K�عP�y�P�C�,���ہ*�aX�Dİ�Ь���&3�E��>�S-�͎���sa4K����GY�ϧ�u�x���zꭳ�HKu,���z�Zwz}��r���RA9�p�`+2�C >K�f\;i��N�1�d�3��&l�m�U���6=#�3�s���j��>�W���>�F��D	^_��E��w������ϝ�T;��d�,NՑF�>��w�~����9�S�J���E���<"�a>���yB\&_3\$:�mc�訚_/y:��֎��tԪ2K��K�Յ��Ğ�N��v�,�b�	�̭}��`Ը	�V�Zr���B~l�q��W�s�T�Tr��諗r P�#)b8�ǆ��}-we����\8T+V"��k�0��_���5n<��Z�^�J�S/&0�zTE���C�M�pm[���5�#���>�tR�3x�^��]ud�2k�@�g{���K�g	f�XQ�<�)X�Q�R�_��2�zS
[�͟�����7>���	��of��AV,�����60��{��"�,WOi^�.�x�����-���sf��RAJ�[L�s����@��O%���k c�Ae.5|9��Y�e��u2��{�@�ɯ�
o��E�k��:I�^6(RoX\� �y�O.;��ǫ�����+/�kF���0$2�z�,�CU��iP`=����?0��&)��N�u�osz��|��E�Bx�:�n$X�3�Δ@9.�B��ê�{G{��A<S<�T�ܤ1��BN��>h��X��z��|�9�h�0�70xC�8ްs�T�� [��x������u%G�Ad#3{Z��}�?��ki�0�� ��!�qT����W��`,����G_����Tg�b�J׃S�O?��~��_Q�:x�O������A`�VH�����\�gB�q 8�pL��J<]�3@��i��0��H/��1Do3��9���X ��"Sl$��g9\ �^m���8/��|aع3�3o���$�\��x4\9V�������PU$����M֥��^��u׼���1Y��_�T�,���EcY#�kЎFS�654Z�;�����,�5�$��I e7�Q�e�bO����!j�{����2*���e;���҆���$�.'X<�#����")w+�x�!@�IH8|�)&$�_����,�|�t��x�)�Y-=$A�+d������Gs�am[��HQ��0;���o��y�d-���}����l����A��{�
�Lr,Σ�u��:i���M�'\%�&���kT�]��;ތ�hl|]B���#ﶌy�t(IdT�?����9�����͝�i�^Z��}:T��R�7`�2��E�_}k�c	�Oz�п|�մ�<�Vo���k��og���8`�OP�Y�C&���Od�ZE:P�_����>>�u�S�q�YJbz�2�
T���N��o�*G,ȶ�h��fI�M�G<Ň����A3΅R�t=��Xz7�U���eG���C )4zw��yy�0d-�F���}0#�!Jq�\�P�_Q-h��Zx�c��ojHu�\�5G��e9����� NBt��B�����3=���[�_���}�7���_U���D�L���o�$I��P����f���[�E��3h��߬��S�q���3*��d��⻶�5�4�!^�T-+ڤ�-��{�J���y�tbH"c�׋�[��8<RA-ˡ�X|��h��{;U����V���zk�Ț]D7�u�X����Bg4G�]�����L�i�.�}�Sɹ�Ou�����-1���Յۻ�u"�t�ú�x`�y�����E�5�k���º�hݦ��k�Up����@�F�<�G��H�����tԗL��-:���D�=ĵ07�y�H\D�$���$H�r��y�đr�o����(2X��UTX,����(�q(�M⑾�c1N���&�l��#`G^�uf԰�y�h15�C�N��o�:=�D]�����K"h�&�k����E���\���tǵ��Cz��\���2c��z@A��~�3R<+zi*�8�?�a�ּ��HT��.q��0οh9N��m���sXAb�o� ���;��"�=L��'� ��̴RD�M[)J�����Lh��Ċͻ��P�⤕S&���@9����y%�	��ЮC7�����3~� TZ+��1�%2��[�O��l��syw�׹4C�fQ�k�&�.vu@�����~�	d3�|b*�Z}��Z�JqU�N+� y���̷BV�-���d�"5���L����J�OĨܘ�23�/q�����6G����fE${�KFP2�ki�9b�-Yu��*K�d���I�|�F��xsa0w�у�f�sE�S�X��J�9	~mc	����O���.�B�2�,��|tx��WQ�c�PX0��X���P=k�C�xoJ�u����,�y�o#<�8�=�w�R6����ԓ$��� (���G��ջף�*��qI�$==��[?�y��GQ�:'@s�R�j?(|��Y�'Y٭� �{�XU�*ċ��w)��հtg�@x���S	������	|����L�wK@�BSz���QbQ�NY�����M�o?w�SDGs���?�OG��Q�q�Ȫ1�zJ���9�zO��2LY�������ܖ����3�ubL���z�����{N����	��5�C���Zb�u�߶`���y����'`�4���Y��sw�:i:��[k\	]��e��/
�5
�cj>^V�?�h�HW����ʄb�n.�*�Z�}�� ��F�}i�e�jBITw{�V<Kh&�D'��Ț ���٫[�F8��l1��Sl��Ι�R*���J��� Vo���8���nAGnc'⭁��Z�A5���y)��+�]ҡ�������K����f�ls���� S	r�CRt(��>~�$�a �F{.�VE�^���o�"�j��[r,�����U*�[A�`��'K�9���@��,��0w�@�:�F���G�fc��2��v��'b���5.��XZTCId//o�ǣ^bTn�pQ����y����ȅ��Aw��LF>��ơz�G&g시�7bWS��|=��(�W��B�&e�'0��f�F�U̐��dc�YI*�	L�:V��@�K�k\w��T�`x�yG����UϽ9�g��|�?n�b��
�qsw?�d���;օ�jU=l�u�j<e_R����A��#a�K��a��찊љ _��c�EM'�>-1xc t=�wn��V<v�k�FD �^�-�F�����N����Ԇ���M��}z�~�N�i_p:ܯ����0<�n�!e�}���Lt!\\��1���s�X��c����!"D?-�����]�#�9!3���t�B?AC�k����ջ��7>��� ƕ�E��LѢ����p/��o����O/�B�%Ղ� e�l��?�=���xַ���]�@�IL"�>�w�k&{^�fc2���o���qlv�G��k�f��|��Y�I����]����Ð�W3���P��	�ӭ�Ϣ��`ɗ���������ƾɦ2�&�u�&M�jxoi�T����+?� (�\G�}����v��6\�b��b�G�Ֆ��Zrw��9�y�M�����N��cA=�ۿE?��l�i�da�m/���𡥒]2Y�o�? xf,7.�{Z �4(=0��e�%	�_��-��v��ʬ"� 9*�������'��͜�JN���p'�p�e��QM�|�#Bf��dA��zv�P��=�;,� jxYH��r�R����S��! ���u�Ԝ���~r>þ�s'�
M�ձ�(�)q-�<����|).��� qy��{��
4-��	՞�������gh��愓N~b��G�Œpڀ�s�������5���%~�/ܪ����qZ�����:F1�����(:��$8%�B��N�w�;��O���;�3�wO�R��:���7D��Y��=�6G��e�׎���X�IE)��P��`�{���7��Kq����]��(D`�����lr�,���@\��|��	�:c�z�qV`]�|�@\��/��aݿ/h��S�ʝy� Za�	z:5?���7���Xu��MtW��k��Q�:���uRer6޾�ҺK����탞Kd4j��z5�J���*��Oa���~�	���2"�Q�p�������(�j%}�Kl�h�~�b�d��p%�É�l`pY���z��w2��Q2��.9����F���w�g�Wq}�L��$�y.��]+�z�Z�A
�xu��h�����[vA/�zS��z(`��ܰ��D{CP�A肓$p8���*Y�������UU圽��/v�9�_^D�j���as	,��.�{i�mJ���/����t�Zku�l��	kCnCG5�#�k�g7���V3-�;�4cE�/���6xFS�bZ=�ހ�	�وB$=�+y5%�Ѝ����y��$U?�H
o��g�w�Q��֧3@��.p{��[)o�QT���[E�^���r�ƒ�Mi��șa�+�6�qQO���@J/��*�Y���R<� �ߠ�]�R��dk/�i�%DՇƦ�4e1��u���]B�&E�ۺD���^�ǽ!iZ��t�T��K�$[��	%���-��t ⧥�w&���xg�Ѽ�v溴�������V���|�u�B�u��%��/B�]�O[{�����F�]����$
[E��X]*���/|��{�۽.�-܎�y�X,���n�t�;���(��"�}�Q?�Z�T���CY҆'l{B���XqiF��(��.	�s��>Qc�JH���	�c�����@�ٞ��Cr'���lΗ\���/�Bnº&�u#�Q��yF��#$�x�0�=w��y[��0������޽�k7-:eW���u���[�j��?A�}z����fwO�G���4ި�s��X92%�ֺ�kj4�@��ji�����E��黉��%���8��Xk�H���	E��C��#��x��"����i�eT��,����4P3���0<< �v</�üH���"�ؑ�,�`���6�q�!x6� &R)>qh=�7�%�mdS�!�#Uq�� ,��թ�Y�s���AU�V3�
�U���#Y?�h� c=�q�Ln�q�����^���� ��^,h%��c=��Hًo���],Z@�_u� 4k݌����^�_�:ޡ���n�'���F����C5���4.��-(o=��|z����s���x�H��cN�������,�Y���.<2�S�]�OI�Id�!�3������5���7c6�H�[Զ�~@�Z)Qp����u�`�ӿ��x�}�';��&��$m4z[�&��D������у�e@���6+��`�:1:i�/\�JN��kr� �G�����3/��[!Q�~�#�\ws�)Ó�F^$��;�z/���Y=��5Qݹ]��$��ɯ�҇k�e����|.����֋ﴻG��i�ef�Q�V�����p�Q�g�� �#�N	��%�#��<�:C2;!����Q*;XVf����A��g$�f.�6�S�R��XW�y���L�
 �r����r	���!��1��������跐�)4:�`�l��"vP�O�#�EZĈ����Ⱦ�tik����c�Y�]��8Y~��=wdu�����i3k�-7��-���=7RE�̢]$u�������'�=<�G}��Gd+�TR�,H���?�2��%�䙩����Tҋ[*`���dSv�R�H��_O|��[��� �r�]Gu_
W�!<��.�>0[�8���+�F���ڥ�-�(#�s��͇=����@I�c*��l�����L��I~��ӏ���G��d��H�]gld�l�� ��Ī��?��Һ���)���lx�(��\����1�J<���3��r+�ؠ��˔4��v���C�m�	�V�=*���	X�����ǲPí{6�Z8�L�zlQ/x	*lXv$.�E�p�p,�uJh����p��qְ��j	:��[E��q5�3]+�Pt��"1��@�3� J~�M���Jk�:�b��5m��_��e���B�0U�e���~L[��=7
���l}���f:Y�Gw�X�D��*����m?���ߡU�9��BS���7D�˅MI��N�~ q��8�<��U�Y�~g�~���}��� �Q��yM'��syo�=o��@������W��y#,�����`�zȷ�Y�\�`�4���M���r�S:�5�˰�D�=s��6�L]��3�_�Α]]IG*����s�9� ]��WM���w�����J��S`���MH`CMB֪�Pi�6b��&���.�����'ϒ�d�����6�Ǐg�
��pc�-\� 8U�p�<�sg�>�R!��r��F��<�ӦC�[�\p�v��=6��֍@)R���d�]�m-8G��9K�#�����/������ۈ�U���A��ђ��y"W�_�]��x��g�(��S����cb��]�J�dR��`g��+�%�u�g�I`l}z⮲Ѹ�d��!=O@�w��]��ds4�~���9%���M�b�Jb��cf��=g�{a�{*�A�Ga���z@!�k~�Q׉������_��oGo8��t�%_.�����ǽG���Px��t�r��+�*6����,�o-���D	�b)=T�\ֵ��s!=�����ȒR6Y�m�W��K	��7�X��qfV��C���M�(=���[�1�b��4)ݚ�W�W��>k��~6jJ�'rc,�ꅰ�J.=A��<�N~��<�a��9�a��e��K=���.	�i[�� �	�pQS���Uɐ�/�������GM�c�q%	���t}�
6:x�Gr/�P0T�^S�r�՘D��R\k5;@FF&�T��H[�H��B����Gp�Ai�^��Nz钦 c�N�l��iQ%�1���B�v�not.��[_���1����+�t4���1]biG�f�;3+_��^S_J�ɨw��Z��=üI����3�r��*�.bo1�t�y܅�8���L�� �r���S���X�lC9��� |�sDi�R\P�>�cqY��5A��Y�������y��׍���,�ob��3������`�hp�_fk0�Z]#�@��G8P�� ��O]�9);l���b�J/�C�lK_&���#�g��V����&ʆGI�T��xI�N͡`�|Bٕ�qK�a���1p�$�	�{]��M_�?ꉪ����K��	���N@c�t����(�h,�ڀ��۟$�Q�mp�'I8lZ��'��#u��9�"�J)'@"��V������D9�3N�z8/J&�����δ�E��.�
=aɿ<���<��u"�ߥ�KQ�ŭ�<�DD�m� Nǧ}/jKZ�J_�t͝�{���<Z��&�+ot������F[@0$���7/%�EBN'`���ŷ���ED�H�8��DA�~w�ʫ�?O�A���{�	&^Y=~`d'#{7���n��'�6@O��=b͟�TY�,�c���|�����]D(�\�^d��Kbh~E�iHf�$N��oֹ �����d\�)�ӰbD&���fp��f&2٨�їP�=�aJ�pN���'����[�V�vc_�P�K�E`�@�B�.nr��L^r�W�X<�}�-�J�W�n�tܢg�ѽx�[���O�D����g!OZ�ĎLZqA����S�58�r["{��>ۙ�C|wN?7�3�m�����G�<��>J�,%�z��?�O��+)>��i���bzW�Á�
�DМ��q�D�X������>���z_�Ea|��U�����ZY>��y@y#�0b�n`����`G������ӳm��Q�^3X*d	��c�P���"/�<[�V��R�b �9%O*q��(��Hv�����A��;�A��V�ːړ����% ��{�a�<;���^���K�ת�qޢ5�� ��9�Q��Q����z(��_x�>�g��}���Ħ5T̷�b%�P�
�S36[�}#-�N���+�,�HqzXʧ�ԫ��gφ�˶c�b]�?��M�.sؚdx���X{��%
�_�f�$����Rp��ץ_H6���mO&��{V���Qay&s������ ך���n[V$wM��s
���,u�
����!����0�l�'��K��EZ]a�)dV���%#�r|��o��������d ݄e�F?�m�����T�k��A�ݓ^��{>1QU�Ȏ*�E������h��w�oR%6�A�u�nۤ;2%��^
Z�ˏ�J��]F��,��Y^l���9�y#����Y�eF�9`���'�r�i�R	��}ڍf�4阐�P�n�.��AZb��}��|#ђc������i��2��k��g��Dփ&�9߇T�䌅��{xOˁ���3��Ū�p�_���di.�ADd9�P=k6��y��h�k��Q�E]��X�8�r�G��B�iu�u��$ș]��e*��Y�p^X�S՗���by<����c7$�0,ut5����t�(h���'T�U��(�9zOw�iTa�%��x���$H�qe����r�5�4�{���?(�Y���y79@9c��F�P�=4&f�G�=|=1����픘�ڤ�)��¼T�p�Z���x,9 ��T��ΜP[�F3Ŷ���}ds(�J1�K[?m�Fd��u�^��G�Jj��:���
�U���ݎb���<���d,������l� ~*�鞡H����i��)��r�4��^�lx+�+���.����X�bREҏBʁ(ؑ�z,�Sз�:r;�5����>���
�B��Ypm㛅�ɼf�g��$H��	;��*̦�������d��5ˢy
����fn�>������]�~�Tg�h�
�U`A��3Lښ�pb���&����h��� �-�f/$�����πd�G�?3^[�?q%Ұ�����V���"�'$�@>�.�W��(2�$�b����h ��f�7{�{��Z����/,d��k�5���ǰ��o�����'�p=Ī��xZ�< v3��zJ�,�e�?�'�њ&w��.��Qz��J���R������Ȍ��m/�]�w�]� �t�"(H��:��
9�	ZiD� ��WFǹ�o����<�>���@2�`�nF�:��-�=�WL�k�=s�����J�,Π|�)�z�[	���3���$�ţZ�h����������Nj��]'knS�i9���x�5#�Q"�=+mK��ۆJFt��EM2�o�)�D�E���AKR_�-�L�u|��v3��9Q�k鳣�����t/ᖑy��OB#��~�5
z����N�vgw�ĺ�h��>y����^oEHu����"]��)�\����Ħ�0j����/Hg�C�[hC�+���i�ts����cz����l#=SzG"Zn�1#��+f)�����:���{,�6�
x�$�̸1��OR��N|%����$ ��>�w�܆ҡ�z�ￍ�'՚7�f8\����PӇ׃.����e�$И���U�o\i�ɥ��?�����@�6�(��)6����@r�����^�[��0Ѕ&I�W|D��Enݷ���ŝ����`�3P�/��Z%[7PX����E{@���b��_�?�]����"���z���,��� 1>��8�XD\�����%}�Ğ�3G~�F���e-���\�΍����Hli���J���49���]gy���o�`�����
Sv2U�1�ܨH�c�\�2m�i���	7?%V�����̦.3�0���%�T���mN���㙵L���Z<aۯ/ı����Զb5n���N������\�*�w-�pL'<��p�$�'���HL����]�����0��������¦7�.�N��+�]c��0s�����}�23�T{<�͝*^b\,�����c�1����N��,٠�t=Z�<7p��q8�X�˒�:�d��6Ζ$Q�WQp�ф潘������H��j����"�����vDIҵO3j�x�`�]�4E�@0"��lw��h24^멎�So�	�7����/�-k��­�E>e�4j���L���lĺ@�2��&Z�&�'����8\�S�^Đ�v�lkqI�B�pm�g�g]v�Ḅϣ�HQ�?���'��,��:^+ǜ�I��

h�z,�g�J�;P�M[t��=�ю��ȷNa����BB:�	×�K&�tZ���2d�6�CXr~��)~M��t���{�X(�&B�_�ľګ���e�:���mC����F�c�;.�GcB�]H���f�e$��26s��=t�ޯҝ"g:������~�� �=�:�?(`M�&��hɲ5p�M���J\�eZZ9�2~��#��N�W�H�b�Lc�V����y_��.&�')@�����#�u��ƈХ�@�4P�@�4��fU�t
��IZ�1�K�'�wm���u��anc�
���}�!M�w[E�?�̊�*"��eW�~#(��x�\&���0�QW�&�E�Z����iR��������g�j�ЃD���1ҼG�Z���v[%-��.u+����I����4������	;����?W�8
7A�T���H�6>�C�;��Z����x����'Q����;���a��T��m����)�H#�����V�ƍ��'�Dg�o�?V��z�#ȫ˴��H^Vto�ܘ�tr�X~U\;m\�U=�u��<��vYN���P�薀h��`%7��!6��%l���[����3m��[`�֩.��_���G+�D��σO_��]te_[�p?���D$�U�Mg\�S[��.��ֶ*�+8P�e���?qb�U�o4�/�@��'�$|P�_3݁��H�K1�W.�6+���Y�EQ���ٮi+$�$�ZL����4�\���7V���aXz` ( Y���GI��'jq}dY�v^OR�4p��(��{F�՗/�"W뺓�hɼ��B��2@�W�Y��{&t��l�ۛ�ː��r�z��j��.vZ�%�f��M��$~�4�6�(�(�(b�+��n�
zP��L����c�9�Lځ
l����m��E*���Y1bl��~�K�1��]��!��U
h������K'G6���G�j��v��2̬�ӃT鞚DYsU��|��UR(�'!0ԅ�K���+9������3Yx1 4�B��J�s��I��8�\��΅����ߠ猞�&&�'�}d�GVP7[r���d#Yt��x�����G��l�A���[|`�$ �8 ag��j�a�&ů�-�vաW�s3	-d����=-�N�OJ̍N_u���ȺG1O�Ad����}&	�h��N�M�K�-�5�l��˕�.���	�2Eu%&��։r�y�
���z�]z$�g[�����ų�(�A�evO~ �?׫A!��wa� ��_�0�% ��'וr���V���@V)tY'�uHV� �k6��]�`�����'��Ӟ���<�@�>�E��U��c�x�A�C	s��f�1{[�!�A��iL����[L%͕���������������y�+��|Žq�y��
a?n�Z�B�1)*{m��� ��#�E(��(��� ��
���_Wb�F2P�G����[ɉ`4&#)�w��Ň�}!fR����:m�c�
s��B���X���>��Z�����rO=SO�l^�l�Zv+Aږ�������o
��f�L���i�"�+3�.fT�Tw!_{vp�&�nR�X�kVɕ��q�x O�t�k(�?E8�#�;:]�<��1+b*���Կ9�W|��xx{�k�5�&k�n�Ԯ�C~��@/T�4�2d+�1�I�/q�tCC ����☜r�>�SÒ}*�jq(����� ̼�Wg��6�{^b�'nt9ׁ�nB��d��^e�ʫ���!y�d���4t��j�H�����������N�Ұ���� ��r���� K��b:T������V/�{��
UuV��D�Z�)d����5tQΉ���;Ā�M)��r���@�]"~c�"(�B�-�k�@���|�<�n��"����?$o�'��z	c��k�A�Q[G�P3w:�J��{�]�]ͮ�o�p��E#����M��g�����i���/UC$��?�����ЯKǈ�7C6ڶ0:�⌞�Xy��O7�V��S��!��M��430h�1[���d'��T��1��e�kI(%�)�:��iMo��H�{���U#BZM+�� �}�x\���<O���eq������������T���[/E@�'���w8ىJHd��,��U�}Q"����4���p�l��rb77ؗ��Z9BZ SRL�f�SΑ[�3��002�����}5�fc�	���`C(�Q���n*�9���R�GT���?u#c<���("]RA��+u)����*&e��m��xǺ �h!�͞�d��r��?�H��C����ڒ[�����q��uC����K�F�I�<̶�PC	55�tЄJ�����l��sɤ8�o���s��T$�(��WvR��+8���&�AL[i�1���l��Fm�s�A�Ҽ45����3���(� 0�A|��y�k'QLF?�r��D����8�ˇ�hް�`�z�,ٝ��K'�He��֨�����҇-�`�r�#E�����8��-|@� �Nq��~��X��?��0d�uPZq+c���$�0et�@׻�Ԗ,�L�R�kP����&�������.��8�3�E��j��qi.Sn�����u(�����rˌ��{t��� ��r�O�1֍Y.��������{+��&q�ه?�}h`tQ%U�j3NL��h�R%���)���Wr`�ƙ�2Jx��b�>��i�û�UA�ü��)d�eCd�ϰ���Vw�T)�@|m�T���e&��Ɨ�j$�D��4T�w�y�DɄ�]1�Y����YO�}ճ9ͣҗ-���MC�<)o�����h߉�T'�l�뛠��� {IЂG:��X���|S)�Dgl���CߥК���/���-%�F#��6�X���,��_�4Y�>K�	j��A�]��M�X�����đ�U&cyho.i�����K��X�	���*�| �+1��J��]��[�!y��0,CA��v�}�����N�,iQP��	aDlT�7Z�o���r��ޘ�������
6ET7����_���_򫾔[�2.��͖��
�k��i�{�~�BpR���7W��X*s��L�X�0�zt�a��4���;��KTҶ%+�5_3,g�5l�)X[�m)q/8V�AR,y��������$Å���v\h)FH�>���L��������n�Y˞�9F���;��X(v220Z��}�A.�d I��(t.d��|�{�����B�.�s�n���kL�C��=����ny#?�\��ɷ���[Y���s%4��q��Gܔ��2������A{�̤j�镒�G �χ��Y�z������G����1�y&d�Z@J�*m�SE�6�^ͦ��m�S�_�qz��-��<u)m~���q[m�3�e��x6㖉���~���lB�/��n
�L𒄘�3d;�������vc>F����A�=;0�䥶<g��ӏ���#4�d���̆KP�:�=V2$��qXND�D��+n�
��8��x�HՌ���P�5�W���s�M��q���D� 4"��sx�d�V�/�JO���w}12l�!R#�ם�s;U΍���&�|��KDc0u&X�m"��D�i�kU ��'���"����H1�
슟=�@D����\Ec�r`Y5�C�V�X'.�89»f!�8
xt�?�L�7�{��+
N��s�o*@<ْV��x�x��Nc�lǥ�9�=]>3�x��njWqX{�("��q2`%��j�.1g��A9��#ǂw�Nh��L���0�O;�}�	�\S��@#ב%N�%�7Co�h�R�!,����=��.�YQ�HH�1�
B�̿���������X�]	���fz��\���+gK���{,�̫^���[澷��ɬ+����������%��M�Cd�J8>�`Cn��H�m�츩��~�Y�]z����e!�^����^l���ÿq�_|m�ަ)\^9
�{�_�-TD;w��{x�rl�(�Y�Rk�K���s�f��� +˜��\�=�$��6KU��F��N$^c�~��ܰZ!
�8�w���o��Q:�ck���e��%f
<3�rN4���x�F��F[<�M|�7��!�=�̓3_�3��c���5)�v����d�?*�J1�{z��s���F
7���GPڡ���Ct
�;��U�ؑQ��H^4'YY�+|9#�$�ހކRm#�V��B���[���*�f��-<�9�(��+���Ȗ�9O=D+�j߁96��ku��3j��{�