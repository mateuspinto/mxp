��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����������q򊒆�
�X49>OC)�GM��N;s$ZT~�ȑ �f��t�yx��MC�6E@)�߻�$�w��ռd��NR�[ݶ:��= #i�s�W��b�rb���Sи�T@��7"�:Tn�!5�'�;~���A�7���e*,�8�GwB���7ӭ�j��b��ª����0�0�jV@��)F���)4����݁Ӣ�+8�}��T�E~e����\Eނk����
V��A���p�Z�$ �T�0HPyQ*�mz޳����̏r��L��y�9]N�v���-�hXx��	(z�-,�d�	D�Q�h�\��Cn�&ˮ	7�1�����Wm1�5���u�ӎ �j.� No��=+�>W�KΈ���I��g�x�E
��M�b�w}8j�iJT��!��:���W����YV���VZ�%��ӝ�2����l�ӄ9�$0�q���o���j���{�gq�*JP���>����\��lF�7���#�qm�5i!�_䃌e?/�#;��MqCx���F�ծ��ܪEW�Dw6��^�K�CUg��C���%a�?�������b|�Fd[��R0bӠl��N��� Ldb�)�D��jyX�QIk�P���\H����&2|<8�5�9b�y}j~�MeބW���hH[�W�{킩���e����6���#��J�����=��1�[ g���P���ՐZ���]�]?�=¶��ȩ����N)>�ʎ�����Wb�DDf�n����4թ�m� �%Ov���WN^�4�K���W:`ʥ���I��0�%�S������A��PdH{���B��J�� :Oҡ�z")f_J�.�،{�=����-Z�~��e�?���J,v���< ��V��e�f&G1����I�3	�jϣd�l���Xçl�*�~hL��*P߽sr��U�%�\��9l��1(RX��ӊ���������,"t%���̴�L���$!>у�}�0�A|sM�0]�l�$O��{\�+��cB�7�"8����3��JP��9o 8��g��$��[�)S�ۻ��n�����:�T�>�z���z�a,h�rW��?��*�i�(�}12��ӣ����$�[]}O�$.;hEA�c_^�ּ6wʿ��,+C���U,��w�S�	mFi�S����c:�l�]���VA^Q����?G�������UC��q�^0lf�c>�F��:j6+dj��Z6��)$�x�z�ݼ�J�BNF:޾Lǻ2��
�eqb��U�EֲR��<2����+(W<Q�ܔm�H�EZ0$c|>�R#?�s�S*�5G�m�7�v2�&��.�ls7��V�F�F�?��R}0�	�C�U������?N�"Vh������:��)�N[.?��S�M^��p=θ.�1��E�����$��W�{�0۲Ã�Ic�榱M[�i\e��� i��q�ʅ��e�fF�*d���D�j�A>(x�6���^J�c���q	��'ZSS�/����*|�c{�ӷ��J'�U�Ct�հ1!�V��ma�_��e5'Y������pZ}"�l�%8ڃ��{A�:�y8��������Z�kT�B5�Q� [�f�q{\g/��Y�#MD�s��,�[���g���G�.Ø{�1�f?0�4z��9"�I�dؽ*�V����w� N��L��q�ݞ�SD%|�ZS�Q"k}��Zw|�%���Y��8�0԰��2/s��o"�� ���0 ���)��S��)�:d�
���N12U\mY�s�0��-�A�����w��IS	oLs�h�d1l-^B9� %�Qa�1����%Տۏ�6j�0ո!���#M":��JZR����'�5/���:q�l�I�������a�?$Ŭ# ��{�+5�d�xb_���>���;� 98>��E��m�>m'���aW��N��Ґӈsm��� 5�����2\�Ke����y��^-WFp��,����5�"��h�z�
F���dlҌq��P ʊ5J��R�i��M�Or� ��+.Xn�r5���@0i�)W�N�7`��4&b��՜L���{L�����>6-��jJ��=H
�Rh�G88$��Q�xQ�Gf���T�xЕ��R4�Mo�LY"E�����;t ��k��L�Y�h��s��c�&r���ܮƓ � u�!lǸ�Q����%_og˂�"1��]��s-��*�[�e�Xx�(���N)Ǌ"�h�p�(o�H��uѪ�������R��d�����GT�j��*�=�S��q ?��2ڣ�H���N�#�&��ᥠf�P��2 �	���V'�8/�
��a@U[�8]��2z"�_�oiN��f���˂���#׮j-_%���:k����MFi�'���?e9�ec�D/�~ٞ;&z��|�K���V��zN��ȵ�u҃sh��b'�ȑ*����$�Nn��-W0���5j��1v�;�&5Q�M˂\����z���G�nAc�2槩�@n�Q�u���ɴSLOn�ۜ���=���s�/	���\�7m��nW��|�z&�h�rW��;ͦc�����դ�W��>��0q.��s�%y����f���׆��H���KE裖�� �V#�oE�3w�"*��t�!������ǜ�5�+�:��Fv�ߛ��3�4<�6��l�c�{����$����nx$�����8�X�b�>}u�, ��os�_�W�� �
�1�LPn�I��D��֡��-�� �~� @�A���X�x�2 r��$��b�ï��/�;�����D�����Y��|��x�����$:m�b��	�� Y�_#��C�B1��;����}J%}��5-�o18����<�l̝`hz�{ޮ�S������]�`m2�^������E�a˞�^���F��8o�̻m�������;bLs�R�xm���@�;-�n�Kq�҈fC��͢�	cb�;�/��=�̩�8C�S���������Wg���	������E�L�[l	5�#j\�6���e��C~z�����ikof��s��ޛm�q����XGh�6��!`���:�dݞi5��k,r��犠�29����!~��-�����1)^]7�9� �g?���Km�߼��a�H ,ڿPn�����|F0$�nο@���D��6�(:�������N?�5�6����z���Q�&Wn��<D��Ӱ���5����K*�͔�^�'<3P���C�\���xS6 ��:(��8p�k��@-�;�����e��" r3����du���d�'[��Ŝ*��q#3�
p-{V�/7#��)d����s&�_�3�sp�êl�j�+)��.���ˢ2į�޻v��&kr���v������ƻ#�̦� ��L��X��ջ����5ې���$�u�c.�-�xk�� ��p�w�Y�����!$�e�J�qX ��}�ϜsҰ�eB��ۻp�@���a4�O҆|Aߨ�W��-�o9ݡP]������h�����r�[Gn��d������@	�Z�i��3	�N Q	xۖ�5e� G�;`���>� � ��]��eT2��T��f�)4c�����W�,�H"�N�vf�U)�M�}(�8J�=����]g�ޫ�0\�O���s����c��Lײh����N���ƩBt(����Ӟ���P�)��[}%�ԫ��eU�D>����Q�d
�~k@E�'��~�*�쉪=Y�5�E#�/���������m��������q1X8�	>�'�{�~����W��W�~RZ������B2Mɨu�g�h!^!-G���941O�mHٝgH�� #�(����ϬϽ��aa#�����9i�ph��](�F���� >2�,T尦S��O{g168V*���'0B�y2{�5�� )sA!f,��W�Ь��,�ŴM��n��#��y�&��<-rLTN�H�������#:�jg����P��/D����X��ǐ܌��X<�t��4^x�|��?FhJ�匋�	BSn!:>%�5���;�b�02+O�M���𢡊�3�'�-%�(�X�*�G��8�����v$+sS�nm\K%d�q0�C���,p�^�j��dV.��c}�kb�Jr�?��5oxc����/lZb;��Gn6kK�'�3;��Qs��p���ZA�����>)T�o`�M���
�W�޶�p�zq�<�gQ�4ve+�WQ�D�sb������7	��u4�����{oB>k;A���,�7��=!���(&Kӵ�nx�Z���[R������+�+T�Jv=�h��