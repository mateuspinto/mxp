`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
bDnVbTb5kE4PZFSxFXVXNS4tyE/Ss1hLweLjh65AoSz5VhjluAB5UmLlkbmmeRxOMO2Lqf/qzJJ4
krXDDqrOsafNpYZ4MpAqasbjaCaYPi/eCOH+SKnsuDLi0oIzP4LtBoA3Ox/18GOMuWmdz/Vxzk8/
bCq/4ktHdvnSFZHf6Jcik1l0CLEE0yaLo93MajbBIbgb5Po3ihrurxGs9KBGxBvkiyozCUEXsZ3I
IlX/a63dL5I/TIWIddl+1Ujdq5YRc7RqwD10ONvE3YpsSjD7XgZdlIPxKIeQPdvjGgwVQKNrqlnW
M7VQ1DkvhOJfKpB8hrw9bvawyd3+MGB5sWoC9gBC2qAD00T+GMdnFJgErrc6HOLHT9ogOjkXxd5b
8aU4yFCqKgp8WvQ+sfsaZ2XwLynMXRRTuMwS++2rZkFaq9REyfsZbsJxEDl07CQVfUpQne3fkw47
tppabWvnENadVtC/Z/JIexMB5cDYcxHnC5nAaHfmEjdp/yhN1NpQ6A+BDq2D+Hi2n51fpm0Yhnk1
SQsnl4+0LJJAnbqdJyQZVKT1U+EskTY1CkznATmsMSCEM9PWoxsIBKA4asQLdbWpH/1JB4HrQsfh
SjgaN8xpeReFFlTI1myuBls9qRiFIioZ+ByrgS2bgd4o6a19ZAC0pkpb4BVq3IHpqsKi96hLGxvb
ZW/B+MiEnI9XEHIjwgUAtcOblH5TTS9rB7am+KFap0cdNWiH2ilvJ8g7dVYGg8j0jy7xFsqTjnr0
fyjjWiMU0uM26uAcsyp66OdzWSPLlTqgwk4ugWd3TH2UEZ+dAkR/MxFZkaXXIpi/Gwbc3RF6Kmsl
oCQfGaH1xmccvIGGkg/lI+cwJEQB+33TXD+fI4hcY/0peCBvB5o0BuJNV8UGky7emOH/+DZ8A2EO
2DXSmlMoLm3UQuEcqLcwhemgr0qpjtID25JsAIvgIM4FOE43S9jTb16GKswNTy59yZ/LtIuGskrf
HADqSYjz5zo4yc/HVccXmze2fDJ+vkHa1RlzwyGXqgvxY0cCPqWgkk3Er5pBhBTzRBXJc6pH0TrH
3zMdzZXC2kcYjxANd+OapTzxFUtlDw8+wUDMzzuwouMOiSK7F5KVdk6U5I6RZnCL3dPdJGkBT5bh
m3IeWWnDCwKF0DkxFRUw6noo5Vrrp8Ok9syCVpwnzu5ombIqxDDV6FaVVdZXUPiBWN5I6+KIiLBS
ukqiZE+sQzAMTDNvZI/CtylQLWsn0cgHQqAUXQ1Ax9L82dX1KCogy9+rkXere1/n4HUwzVPHfLuC
94+POZ1Xi6sRqyTb9LZpXRfIVjSCa2OLBgTdTR6cF5E9hpo3szHUyLKm/gXE7ml8hiuWTRgARSUJ
55onXt7sdTl2Tfviw/ERgDkDaeS8D/kkfy+0Rl+IZvor9lfz4mJXgNdj/KlOXIlRHws+bwKUMxCJ
QWlLXzB228hgdE6iCdUik2x6Bzk5/Stu+c05w8r964tdf8XQIA==
`protect end_protected
