XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����P-(�h����Y�*��hı��.�2̳��?b�p��N�*`�Y{����C�6�Kw>='�	ay�`si@<þPteH�6$�h��5(�hK��RD���y�V��|�$C>8���Ww�|[��vi�p��`3�))���m'EA� �U\�����Y/��ZH&�n��,�c`U�w2���c�|���ލx0	`ƕP��-Z�1�����1��q�2����H���;�)��o7nW[�v̹tIeRw��^/
�]Z���/�]�^}<�)�'�m4T�_��r���W'�CpR/Y�|GIV���3n��0H䷖�mF�Z{�����N�?Sj��w%��C�E(�)9vej�o�(ՐfX*�*���qRD��q�My��S&�����c(0��t�7^��!w��L�BS����ɀ��D�2�ʬ��zzv�z1��j�s��	-j��"�4t;b��T�d[U=���J��_���'�"W�M�k�xD�o�N��7��0��E�^��
��j*6�
&�N��WBL�Q�Yx���z1��#x�}��3���Wk4�*T��F��D=�+y���a1��|z�10�%u��)"���;3�����t�|.\�@F$Z����4��c�=�5A�]����U�zP3��]��<:C�U��k��ϻn"�{��J@�6AuU#��=�yE^V8"5	&��gh/Z~0����\B�⛷	�G�¾�R��c7}�������[�XlxVHYEB     400     240(8��[Ͳ�	�>���-){�E�QV���2�Jd��R�^O����Ab�Z�x�	��i;��ϑ������+N��������v�F9��."^j+:w�^�4�rϹ����	��SE��8��J�]���;�c�h��Mm)�|�y.w���/����W�z����f�d��������O�d���%��00�V�N��K�ݹ>��3^�C����,O5��$(-	������Ƙ�Y�A��}��ޏ���/f�Lt�?���׵�۟���'��h'J���G�R����C�M�Z�M����AL0!\ tsx����Ҟ⠟�qe*��,������J�����U�p����P��e�O[�,����.:�̶��E���<�#Sw�`�&Quh-�7dU��`~VY�G��u��*�
�J��� .�0�}�)$\%�D!ǧ^�E2�R�5#���|�]����*��+��23Ah����������������8�`�LF��ǀќSdE�(ϸ<}X��]}�����+5$tL'k�+zkB��㛖cBV�m!WrM�5,
���P�d�CXlxVHYEB     400     210�>	�U����~=�Q�(�ޱ�U�zz�2Q�J�����Bb_(�hu�16��}bY0>R�D�͹Y�ɲr�	Ѝ�'�����?�⽐��'h)�xs_�c�2q����H���>#��2 ��*�'X��j��R$%H��:��V�$]~�9[�_ޭV_�K��ءl,���7�*���󇦬�ڤ����b���k�V�R�^6�	�~IU�H���9K���Y��,������}c�D��Ih����r���Q�ޛKV�ި�Z5�^:���Ϥ����O̦��?�ͅ�W�<o:�I=.�H0X�F��ԴhSY���.�:�J5Y������K��/c�}P,���=��3�Fyu��q0���W>0	�j(+�ԭ������3 �öǆ��o�z�Y�[����I��I6

�G�F�qq�h�N8ne(��؁칺Z�R�;d�,_�|�+�yȶy?�0�� I�<��Gk�Gt)�^ ��?�Sz��6p9��{�1�� ��r�f������T��:��JzXlxVHYEB     400     1f0�S���ٙ��b^T����T^�^������?��@\�\]�Cg�0\Ss��*�;���E��Vf^�[����G#�K��U"�� ¦�{�mHIl��P7��Y�{b�Ѱ�\�7&E�_���S-k$� �?P"2���R�U�a �?8b�8���������K�\�#/�3~#/���ndV�,]xQTg�I�ʇ%K� +J��L���y�ة��o,27\�X���6��D{Iа��<����?� �ý���1��.oog�� [�S�=R�i��1T�@O4������@��9�;�m���b������̘��Z������<��9(�	�K�������CP�H�$B�v�W�$�߆-?q�O���5��l� P9qI�ث!lz��y�7��1��.��	�Ͳ^
Ѫ\��ia	��šo�
-	U?��m����t�9���fo?���L�f�4R�ȹ��.�T�;@�p���%�-#�&c��?���q*�nXlxVHYEB     400     1c0�����6��<�����Up3vl�0I�=��S�����"	��l�t۔�{?�ݖ:+�H�l�w�+U��B����8�Bi �28�,n�/wD� =�tJ�[�ӫ=���Wo>-���U��8��u�4Z�����uբ��U��[��q���@�5��0��Z�e��#ɔ'k�� ��	.�(�o��{�r�$���Gף9���L���d�k?�۹w���EE/nu(��N�K���藡�����~���C�L�(�'W 3(��i�Ҫ��c4B�u��` ��?Z[�����L\��O_l$Zp����B��u��UI7�fr)�ͪI̼X��,'�#	[sf��ہ A�gs�7�찕��BS��ƒ$V�$�WZ�\�V�
Y(�(�w��x:�C�$Լ�$�+#��(<e_�Oc.�#>8J)O��c�l�)���f�<XlxVHYEB     400     200�=�S��<���3��0ɥ���|�ϲT�7+�W�n=���Ny���w ϻ��pP,���ˀіM���!*"��y?ut �#)�Gc���q��5��V�W�o��{��]�'�������v�(<
 ވ�?�����g����ge�k:�L�|��i���Ga<Q#s��ǈ��A9 �+F�<6I9�k�1j1P=P��ɺM�Zz����~���e�%�#o3�,��i���|A�\�MY��
��.xl�P� �d`�Ґ)�����ւ��i:��� (�|�&搐}&yX��%�(|�ْ�5��3����V0�U�'�j��թ&���i�Ln͒ߑ6>�%��rPu^���x��N��S:1p��h�(�薎7q�D:"_�z���l��"ߡ좹c(il�i��i����\�m,����m����-:\,�i8�D2S*J'���J�c�!�`s��/���2*A(Z�^��DM����d�<������[?R�c���ת����� XlxVHYEB     400     120�D��5�Ƶ/S��h�p��f%��:�ρ?_e��a/?
��m?��7�奟�3�gR����U�v�p`o��N�W���U%A1��f��(!`�:N]P*�U �n��4��Y�{/�A�G�n��h7��\�������!�Z���_����;��h�~%Y��!O����!��l��\���[�) M���9�&�p�/\f�b�K`��q���Q�p3�^'|e�d(�Ny�c������d�����\ä��]H2."��"n,����v�JH�h4��QgJ�����XlxVHYEB     400     1a0F? M.��dN�P��h;-5K��{��J���5A9�G7��`X�Ѝ�Y�����pU�J� ���b#�b3g��$s
X��~I.U�`��Xx��'��W�zW��F�Vڥ/�x�>Kmm��R���'y�����I�O�� ������̔�U�c�hf�����*B�b굗6o�?,cׄX��:���V��a8 ��������6�L9���;>�2W��m�W�B˔XQ�x�_�����k�ͺ�8������%�yP�fH%��1�ؙ�	��x�Soܭl9���*Y2��e�/{ǌY�l�m7�I��=:�m��N&"?f�O�'�>��F\hW�'����Sd��yB�Sl�I�M5I� �1P��
)�"��о���n!��)hH�|�b�L�ʙћ7�X3n	x.OS:��f�XlxVHYEB     400     110��3���}��^��ŜC��C���S7�T5�G�s�^.QvŊ'/Ǧ/���x������	�z,>(�U�� ����f��;�Q��s�G��y]�q��2��]
O�xI�S2ˤ�]��`�〘�z����I�L��$�iQy�I�{�-Kt���AcX^[�'����Q�/��wͩ��*KKN���Q����W%�<���G?C�x��To�Sw��r�鎡�bؿ��\�7�ﺰI�����j�+�T�?��
5zZi:H&m����s�ВXlxVHYEB     400      f0��_��ԽM
� }K���{�ӓ[���ۯ��u����ٺf���%��&e-��Ė���W@�h������t>�51���v���M� C�.�Oo*Wњ���������m(�p�p���᜴������V*h�IF����Z��!W��W�d��M���g������L[�;�v%�!��籂���ھ�UX/0�_��'�#���fsjf?���m��h��z�~A�-HXlxVHYEB     400     130�.�[�"{}L S��<J�,���7�|������Atb�rIY} ��D��+#,�\�$sz1�YQ�~�KV�F^�BE��c��9����9��A�a|ݩ{&�vt$?,�gE���U��_���`#��iK���Zb�r�a�!鵒W�ƾ]�ɑ�b�1^��UY����0�<En/�M��!���'��|=����?o_��"X�ష�$�?>
�g�6��g/W����Q�y�FP0j�4� ���NIV'dE�������d��&O�HRTr+ǡ/�/2�R�䒰`��XlxVHYEB     400     130w�T�I�O�7w#+���e�hȰ{�Í�":����Ʒhn���+��c�ۖ�A��2{zY�1� ٢�rRfj�o���7�7eV9P02;�Y_$P�~qrSI2�g��K����{�Hظ�p�?E\
��z�%3TƮo����C������j p����$q\���z�]ŭN"���8�T-��Z��I�wTz��8��k�o�4F16[5�Mc��52Ѹ߼'�/OO��Ek�q��ݸ.�A��A�s5�Q]3�S�'X�Qr( �]]�p���lI{B�޷�o��y~U�7�����(�XlxVHYEB     400     130걦r�#Z+�d�CD����[G �uɼ�[�0�]���ǤS�פ�Sʋ�dM<6�ʝ�f� ��>̳��CLV1���{�k{�W��P�a��la&f���=�TÇ�;��_���55�%���8���fQ�$ ��	�I�;J��95��h�+ߵ�\�
$@���q�w�����vZ^%:Ҙw������:� XDeY6'��D2�N"��
�!�3�3�VٝW!�}Z9�.%�&目8>۰L�D����_��?�EH����B��F�� O֫$*-�[�m����KSzGs#�N��,��e����ǨL�XlxVHYEB     400     190�Y�c����_�����R�����c�n#�be\�]\�~���?�yBW�_`��ï�+�l�8���UXD��7�IQt����_�w���wO�+: �s1�̏�9�Ź��U}-�vl���"�k>�����yQ%3�hd���ǲ�N��}-vv�\�:jD�� �>m֣�����.���3�QzXC�i�(��7�׻���
^�D����%E��%��eN���4�xN|a@a�^7�_����We���X�;.�-�k��A�1`���0�'1G�ڠ�,�>�Z �릨�)U[R������3Бm~��7N��Z<OeN�0�X�($z� �,��5܊e�Y?�=6F���b�6���V?�!�"43X��n"�|�
��}�����rb��XlxVHYEB     400     110���q�N��o��^"���o���u�����Y�1�Rs���v��߫���k��_�{� ��ۊ���q.��Xfv8Ӂ93��Rٱw���[��v�u���Ӂ�q{S�� LY:�!kMj�
��.Ar>l�Q�4]+n�e��YQٲ������ ��F������d�$H��zp����Q��j\�r7d�� m�]���DK�� 
G��r��B�H�,u4���Q����p�7XA��yUG����<[��%�"��A�9���7��v�XlxVHYEB     400     1b0v���H�uxDk`d���c�WDQK��m��S%� �C7i� ��8�h�x٧�y�������v��[��-apӧ
���?��B���
sB�d
��\�p��/m@M���Όk�|䫚��Ht㪞qӚ�l��-��Q#�`tr�v�C�~�)�.���|A\�Od����:��lO��}0���LR�����T�w�_�o�]6�(/��<�X��*�6��Z]�O����J �*O��X�iГ�����+�VQ�?Lϸ�S�@��x�_>�/u$��X~p�	(�"dW��y���4g�c����FqP�GnyhH"Q�g�+� k��h`���]N�[C�*a�:��+��܅;��`"�I�1��q+�sVR$�o����W��r�ّ|�����"��?@�lQ�F���_�/o.������������F'�XlxVHYEB     400     190��8N0�S�w�T��ք�����č�_�E��JQMe�l{C��.�#bV�}������t�W/�G�VQ��԰	�m�G�l>B탲`��<]�Ӗ��?����y��.�1�a
�.G���Vy�C��MR��'�f��j��'��Ն��֋�p!ܑ�e���8�1:Uy�v�;�݌��i������|ۦ�e�FJ�m����(�ORx����8��E�z�쀙rը�`|��ohj_�	a���5���i���!��ޕ���͌*�E�fD?�t,H�K�b��7ck���p)*�>Eg��b�'f˟�X��4z�IU�##�D�r>@ox�2�4G1y��Z�kj�'���4�\>S�$HE3e���g�LF���i�8�G]OXlxVHYEB     400     120d?縏����[��D�8��B��<+NZڂ�"U^D,�k0WzuNJ�+��ޅ5�^E�;N������Sݹ��F������ H�i��Y��\�3��A��z䀓�r�� \��`��) �*�z�LW
�1�,�Z���:w�zG-û	����^JM c]��)�(��D;�hl?vU:u��|�+�gQ?�����	H����Zs�sqE��g}ȋ��U=�����LR; ��.��"��}���
b��"�!i	>�	
���\@]`����ġă{ɻF}�-�4��XlxVHYEB     400     120�^B{+[�����0$��.���?�Vש�.�'ŏDy�>������lA���|��X.�pt�n������>��	O�S�{	u�)Oqd��������Ӷ�&S�JV)�2m����7�B�ʨ�0xk�ZT���m�6�0��bc�|����x��N�{soh��n�-r�Q=�{��W��H}�s:#"�����8�K�H"������,s�F
)q�V���yS��������������(?�/t��+ݜ KD�y�<�w� N���+����%(��ڍ"2�3T¬XlxVHYEB     400     160�ԑX�k��bZ�:zկ0Nw{�1��#�nkL�\�:�G����I��~(�&����B�4H�d���֏�t��{Y,$�r�B�ũ�-5�{������\&Uwغ���Oii�#0�E��zˍ��&�`����G��Ae�J���9��W��NɎ����"�g��8ٷ�uXQ��
��%İ���/|ԇ�?�Wv�H���2:;���9ѝ-�G��Tͅ���h����ץiE2��ʁ#i��a�iz�����y$�(b�Y>ء^p���h+'���kr���r�C�PHA������l���Y��:"x����υ�□��1���:�8�|m4���)��-� XlxVHYEB     400     150��/��=D<M<� \�E�1�fO>��� ��>]�\�r��I�P�
D��H���Nf`K 4Fp~�b�jJ�t�]E�	�_�H�=�tq��p4��g�J��wH�(�q�C:�����~=��o� ���8 j����`r� ]JZ�WO����9�V���@XS��P����4uw�a�O�g�X�O3�\a� GUV<i�]��'w�A��N[&x �Y��/�g_(-]��u��,i�ڿ�����"A�>�R�f�jMO>wЏ7Fkw.�;�ŀ�%gH��:��o�
	p*��z�!o�|�B�p-a���)<9L�6h^�9�e����n���>LXlxVHYEB     400      e0�喴{ǝ-OA|�dlP>/���(wq��7�w0�����ڻ�g�Vs�������9$�-t� |.��#�ő�׀/�vR��`7	�z��ߎ�crqGץ��������CLCP�菠�yx"$3�u��oqc��?�)i,z*���w#O��I�F���p�3ڣ�ǵ*"pFxNO(}�,c���cj�W�op�zaP�#uޔ�q�U�g�/ c�>�<��ԃ�R��XlxVHYEB     400     130s�t�MM�p�&��/<����S���,��������w��y�7�Du࿟4��	��K�!u��烠
uG��ʣ��R?���2j��.�ֺ%u���߶���l��e��l{Ы�����M�
cĀåf��[Ŵ�$%�W���IQn��T'i�O��G�3��Ҟ<���>�|J�U��Xz�4�w�W���K��҈f�C����6j��T�Ok�m=CX�7{����R��mgӁ�b���,n��"���:o���'�g��NM�>����3�d�mi���Y��Y�
�^�Ѫ,T�p7�Q��P��hhr��߲XlxVHYEB     400     140�i�3]�D%-�k��JL��``�IR�Π7&���%�xH��X���Ar �;�Ņ@�7��l�����[�y��ʚ̝��Ri�z�)nXH�����3d�FI[��Q��략V��X;gh�:'e�Л6�/CH�c
"��n����e�	f����;�y�$�����n�_��r�&��P��κ������5v�E�E��j���R�#Ng�ɓUk-5�J�i9�A�2Y��<$��&�K8&1�)�NY���-T6��Pi�5߲���������8᯿��0�d�A���K�d}����0��XlxVHYEB     400     150��<㗐jY�2�R�/��-��q�T�j�e�/_�N5Ώz��y	֥��4c��28�e׮����-�f��1=�ZD}y%8��]P5��qJ�De���
"��+� �X_\����?�H�朳`|�y %� t��SS�NE]<'��k"ydh��E7�q��=�OƗz��W�'取����-��S����>�ØCt$��7�e��}�[����]��#Z�/Mɫn�i�pݿc����}�}(WR�Z���#hfy$ܳ����'YwUT���8��ޥ�&ut���mK�#��қ.Wʠ��3 0 ���.!n<3J�}��N�u��XlxVHYEB     400     150]��nv�?᭵Q!�L&�㄄���L��J��~q���k�H���WZ��#�N�Ы��5��:	x`�����:E�ӳ���5�g�1�����D�+!�B07�˖ij[g�����¹$.����Dy.��/� �j;�l���˗)n��sgW�\���`�c���+�ˀ�*�̅��^�B�Jh��p�2{O�@��OM]pmT���HX��OO6�Q�l*M�m^r�p'F7��G�����P�$}}�]���)S�Jz&�s�6r
w=����;�|:�����h}�ֆMz�v� 'f�����`5�����ڙ!4�=�����<M�juW��_�XlxVHYEB     400     120ʬ�SV�a�V?��f�_:$���߆c,��0�l��'+4��z���Q}fA���8}s�������g&���h"�V#��IGǓ1y�q�|'�J&_{�u�1]�5�d28�W�K���\Fby����D���n���FVOu�S�p8
��}�Dx+Y�(��j9���a�s;��P�Px�:	�G]�b�J�f9�3���7�[vL�*�<z�I�:�r��|_����C��s��+����K������_[��\=�Z���A2)�V��4=A�O��LXlxVHYEB     400     130�t^5Xߙ�ʰA?/~�4G.�������������Tbb�Y��;H�����mo�6F�gM���L6����5�Q}���|@�r�����)��t{���O;�~o���I�o�O�#Sܪ�J����A��r�tt��BCc����BzL�B�D�46I�=?�@g����RP�;��Ԧܤ��l�U��$@����i�����w��:O��e׶��%���h�t{UEL���b졈3���y��۷{�K0���`v6@�4?�5���P�<,Wr�l�Z`&?Z`�%V�i|{/G�(��+�n�XlxVHYEB     400     140�+�r�QsNm�1�g�=��p�G�Oy�c-�ze|��n��b��m�W���1؋���fyϦ[ņy�n���� ^t[tV�/�޵6�~a-�4R�S�+�]�˲ET�D��)�EŇi����,��Kƴ �ol���Ԁb �m�	���	Lr���H~�M"9E]�~�!kJ���$@r��\Ŭ�o�zܶ�C&��^��<�e�tw�O�ݰ$�Oc<Q
滎jp��
U�՗�z�$'��ϙ�^��:� ��0$ĭ��_G�R%j��%ᘥ`V螈��<4X�������P�T�>���p��Ӫ�{��XlxVHYEB     400     120g��,=r�[`JHM��^'�L��4*�9�e��'���`_w�7U�;D!��u����*n��]N̤'Y�l��!�w$�:	:�c`���/F���za�o�ܒ5w�C�K`,��u���7��4?4�`>�T6������ZH���l�0����G.�k�i�4~V3���7i4��*?<��ǐ���0��6�N��PI�t���F6z���Xۙ��a.^E�[�t��\�� �sUМ	ȴ�n���}Km��ߴa��h8cnv�
�\} �ݽvXlxVHYEB     400     150���ߏ��/T~��݌�}t�vR�� �\�]5�N�V���}lrL�I�Y�ȳ�49��w�&:����G*c
D���Vp�x�,[����0iG��N�'O
���#�h�ɥ�'�,U�����1���nht���yΉ�}w%Qm�x����յ^tn-�X�k=�m�$�}w�W������z�A�]�}x<ę���-9�>�����}K�~,����
d%<ai�ie>�WCh� ]��Q=\T�V��Q���*���c��w�YòN����S[	��2p�������o;^���q� =8� ���N{jM(�ƀ�p�GCy��O
l�	ИXlxVHYEB     400     150i���y
Y�Ȫh^!:q!U��я��H�e�Y|��$����/r�[�`��Q�c5�Ji[��B�yM.�i��˷�ڴ ������f� ��h���!|/��%��+0�_Kw�T�7�bE�k1U:S�3�10���o��P�C��z�ܥ��0�&�/*qN�D��i��䱐�"�5ɣɏ�K�zl�D���O���A��hh`*�A|�#��f�_HF�o�5��E�:!����*�M�HS�G���QBW<����f��D�-��l	I�so>�9��z��s��|�o��3����wޝ58�	�sk.�\T���Oٓh2����ݾ�rX$8XlxVHYEB     400      c0�*Ѷ.c��_�!�`��Z�/!%dk���\17���O&[���k����+���K40��{�g���U�M� Ã�FA�w�$�bGCY#0�wd���QD*m�N���$�k�x�A*L4��hj�!�p����/O�T��V@+`�F���"�A�h�
��WZe�"�,NA�J� �
9y�Pk�.�XlxVHYEB     400      c0`���dox��(�vu��K�w1���"B��Q����31���w���I�s�t�m�Lρa"�

��������R��[�a��##iU�ڒCC�p]�ՆЇ�N�2�=�Fn;��ԆDcV]������L�2m�l�iu�'f�c����]��w$|�Uj��-����Ĭ����/�_�3�XlxVHYEB     400     130�C�P	�]"���}��Z�UxƲ� �|mZ�s�ރ���ށu✾Y6��DN�6얁�v���,��v�t�N�GJz�s�).u'1�wJ��4�Y�]�h�L������4�H,[� nYd�'���?>�4�SS�m�� ��r` 0�ʙ3�\r}^Ҙ��������M�a�Fwa�ǷE��GE�ֲ�)֗���d#�����<�l�m��eg+!+ETX�>u;[�R�e��*'5e@�<r��}:��R"/"��V��E����$bFv�a(4�̧wl�3LC��:B��T�̡��/�F�DQXlxVHYEB     400     120f���W��i��\���yF2���G���6�5�H�x˾ʸ3��e�ZP&�E����� ���-�|�c�&�A/d�=X�W��d��S��B�9�k�%8��a�\���@�,6!���[}�=�����J36��M7������r�qC�Z=0��� ���K&����t�h[-Ԟ�13s��R�%�
i�Ir�!�N�*�KS���ـ{h�H}�-�ī�(�%���E��XW�=z�=!�ʻ�5N�÷W�~� �=>�h5m��Q-���8�F L�bz{v�i��$XlxVHYEB     400     100�:%���/LVp?ީ�왨���DZ��U���-�?
ia�-ٍ��i�l�0���I`>�׽*�8F ��{��Y�iS6���(��@6� �ƝK5jg�H��?!3�j�)�c����S7ZV��=\H7�^J~Jڱ-ƢMw���f:��mI�����[�x9��~�xsѐ�9��Zp:?�b���l`��3ȥ�3��b�k�(�P2��������Y���*h�8��w��y� e�9�ҩ��UZ�Qџ����u�XlxVHYEB     400     160��դ/jn��^<H��٭o)*x�C<�˶:t�^��<b�����]0��WYNCQBH����g&T\Ic=t!5�'�('XL�&,��B��\`�SMT��/½v9n�z�g�B�=O�f\�-bn�T��f�3ߋ��~��@v
/�igT�W�����C!-R��q�����[����u�Sl����ே���rƑ��J�\��}�gf.�uK�}�jBm�!��l��UAD@��zO���K����ZS��G �PPMaMe����vIɂ%!K=�YBu��2K�x@)�E˱,���צY��c�"E#C�S">ۼ�r�� �M*k�G��?k�uKDV��XlxVHYEB     400     1c0��H�}�صy͠K�?!���]oZ���ҁ��( :�-m=��܌ٹ�h2w}�f�m��u����0����2����x�c:�i�q���W,�����(�2�?cA�� �"��B-��</��'�eL��l���M�S��FA(Q
\V~9y�Z"s}W=,���`�n���]L^�ZЍ?.�r����	;������Xܕ�M�f��_p�P(�*z� ;N�d�H�[���-J�.� ��CQ<3�����zԙ�fݥϝ��@R�4�Tq;�O[�&.��iܿ�8h��_��5��hے�a?��y#չ�*!�q}w�y����_PC�Mc����>la�x�}���r�m��4����ln���7L�
����tjn�#C�di���OP�5�cUPz�?�������x�>�>3��;_(
���Q� ����^Z9T�����1�XlxVHYEB     400     1d0����Lw:H�1NoeJj~&Y&&����g
�~���+T��|���m V@���J��+��;��,�-Gi��I��J�͡���ZjN\�����܍Bѣ<Z'���ǒ��=�3d��04ū�H�h�Y�0�4�)/�Ԇ�սu�m�����'���W��7�����n�]i�O�<!�k�o��N��h���z�X[��(1N^�f��䳻�WO��J�^ʄ��QiK��b�Gv��p�iQ���)fC�ѿ� �w%'T)*���Tv36�LI�'��C��3�0����ҽϷ��t'G{'��g�P9�5�n��=QQ��g���3u�'�8�x(���+;�,�0�z��+q&d�YQ���Eol|��9�{��s=:�bq���
Ӷ�Eg	�[��)�s�E����(�=��͙2��u�dL���t��T,�N��<�R讪J.�s�Z�yx�OXlxVHYEB     400     1b0�t!���n�%�&TȓX+M�,�3:�"�x[n2�d3��V^��U�T��(�X��CZ��2��GBȋ-W3uR
NI���:��g_�8&��욼gt�z�y�S��U{��T�X��o.@c����i|o2q[�=	W���ԏ$�P�5���og}��9�p�챿�t��C<8a���>�ҍ����I���1�K�^���
m�\�u��zs��g7'��LG�k)-�pV �7�K�X[M1=���ZRONN�.S➘%|��R;C��H4��`�yΆ^��b]!ݻ,�"�Ot�+x.sn�	V�o��~`'rv*�|g�����8�	�h�e�N��Њ}9���Cѧ�/VG�fPǻ
��֝Cr^�VF����y��B"�<mб��Sҗ��ZTH��4z�����9�f�w���{�0�-�f2�o�V�XlxVHYEB     400     1a0P�0ޮfø=���I-b$�u*H��$2�����0�fy�B��`�sg<W�+�d)�I����Du�^��j��e�2���8��i����
S���{Zw �݂��r��ݜ����ڶ������^�y���O"��.`d�u�򶛛�˘|k��S|�f�T��cَ�I������~�W�(��,2	9�Du��� ��K��<����eD(E�7�͟e�\V����5H).>�;*]~�A�r^�N"�>[��g{::E|!�(�98�g?�l�
�b�YX\�V�3
��6$�@��9��TO5��F�2��y�#`�����̈�H�[Ϊ���Vk��m.X� M��o��{v�����_�]/�T�T�`����`Mf�4FM�X�J<k8)��S��XlxVHYEB     400     160�'�ms�BǸ��2<ZtyC�a� �>K2$��8�,�:3�\�Ӊi��`T8�S��J)U�K?�N��z�)q��)����&���c¸�o�뽹4q1�"��{�m��>,ѫI����`�$ν2�����	��c;z�}�`vm\<�;<~x���qw����,�Ԏ��Z��"kr��Ua�����$�Z�i;�x����b���O"�CtG�v�Fp�#>Y�9����������VM���a��_�
r{�YA�|rt�Ǵ�K<' �_^��/ڛy�G	39[x��Kf��1ڠ��BcΞ���-j&Zr�Đ�ف��$|&����c��c�#V�O�լIXlxVHYEB     400     160��Z����ꯄo�8W��\^���l*�Aؐ9�\/q@A���ϼm��8�7eAXx���$�?�>AiG\ ��n��i���6ڽ�Y1�G���4Ǻ���Գ]C�=A�
N�ć�ĕW��F�ԉ�:�v�Cu�&k�]��;w^���9����ǣ��_U��}A�h��"9@{������H鴏
j�)-�>O*�
g��y�n�6+��Ds<1h�WO�{�x��g��Wx�U����=2���'TG��5F%~������;X���%c�S(-�2|,;Y���
��$5�3cߜ����zY��E�Ĳ�x4~�\y/};䟠�1�[�J6�J��+qE9�&�W�\,K"�^�����6�XlxVHYEB     400     180P�>ٿ	��>Bb"��d{PbVa�|&FuY���ؓ� 
 ���K�N�f��T��tnt.��=.�\�r9+"Q���8��0�Z�����g5?�)ꩴ3��w�W�ȠQ뒋�� �ל��{�+"4@�zV\!��U��.fs����G���w�L���2+��^�,�}����ٳfl$���2{8�kV \��h��*%�H�_B2��vJO7��"��C�i]$�£��k�p����b��)V6���^��͎1���x����0���S�9���7�R2��,έ��3���/�?����!9͉�6I����{�J��c�*G>��dv�Z�#���:����>d<���᜕CQ���Q�D0����ҥ8We��XlxVHYEB     2ed     130d�̃���["��n��F�)�Ӷ���O���"��$��j�9CЉä�{>;���ً<QMb�t49�1�����f�5�#�Y<��Lٹ�;��S���;���Y �0Rb���Z@&�\H�3}ڶ3I؃<j�E��m�;W��Sb��E�宯���u8B wr���~l�t�+^_ܟ�=���r�����)rnZ��N}�~�w}�?X�L}�qCE �'[�3y��n��X��CUFOq����_#wM�~|R��X0M6��4tؓ������r�1΋~-�j�D>���o�Fx��S