XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�a�2���}{��\�9���0�>\ۿ�wj�h3!a�%I�f�
� �[,"'�\�������J_!����V�uC��PR� rPN��o�3�|��w%Q,��K-�;�^�W��Z����?MUġ �YcqO3�M3D���w*%B��j&�#�k���w�l>� �=��>�T�j ����d�m��ǒJwz�;�䄁u�"u_3���ѷF烶!#2��p�(Wȧ�Ѿ9�ٱ�6��Lܟ��9֡c&��IuA��V���0c�2ʏ:�Y�X���x����9�-%�-��I��-�����gZ�K�����#������d�o�:���u�9(�i�Ճ�k4O�H���$�R��e���ms�0���!�)��Z���0����\����4M������v�~�Y�Q��"���:ۧ%����k,I�ߙ{�H�E�w�~u��n2UV��5�\U�.uІ��SK8ܶ<���o�8y��f�F��l�C�Q���� 9�W�N� ��
��9��.C�F�2��RHVF?�2�)��Q|�jqXVH��R�7c"5V TZ�AXN�����|l ��q>���\Me�E2m�X��s�4SRד���7*v�C������`�!+6v1r��/\I���ޠs�q}�H�a_8k�*Bbi��6�-�jywÀ�;|�9��hX
>�˳�n��s�M�6�A�j�o�8!��p�(����Vߤ�̓�`G��ܧ����.ˌ�u������H#;5ih�XlxVHYEB     400     190��v��t���d�#�}/�����L#�0�����{���#�>U��v�4]�w�t,������`����&"���B��r%��n�ܰ���3��X!6�^� '��<O�B��
W #��Rӷ�/���w����!��
�g�׊�3���<�#�&٧�{(���6SB腩�����|K��1Y1b�=���K���/B�ي�|�MA�a��J��|�C�U�S�]�R�:�m�he�3�%��`�v�ԇ� ��I8�����7	֮>�\�4�*,�w�&�W�ٹp��}Z#�kK%?�p�K�`h15w($%.�f��ȷLyͲ}$"wB��;�U���y�i�mp����,P��Ҽi����Ʒ6K�p_�O�]���{� ��I")A����H��ؓ��XlxVHYEB      3f      50�m����b�Jx�+&j�t(@�SaCQ~=N�&��λ���$n}�R���ţ|�A�SF@@�=�'��h��ߤ���:�