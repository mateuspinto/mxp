��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����Ol��v^w ���Ʃ֔;i)0��D��J�{���uw����}M'�gB�7W�ꀨ���vǻ�RGL5�Ƒw~��O�_�Ɇ��gPq��7R�Znv�.��8H��� ���K]���W�^_�j��0�v�	Dg28+/[�u]o�M����.�b!�Vey^[��!A���c����+�p��%�=W��xF	��޲���|yOa"^?�ioy��:V|�b��IG���B�E�jb\���RH	�v#
)nPU]�ܕ�=`����5q/�NM�y`N�UB��HJ�O�G7 L}1�#���[�׽|��8d~�A�9��՛Un$п�$ C����j8�.�Q\�"�}�:Q;^
*Gd�e)�;������Ue�T����=��u���D�w�i��Yg~�Ph1�� B6��-����Yf�F�k?
&)�S[�wX+��N��oI�����&���ǰu�����|Q��"i���i�bع�2�z3e5�E�]���=o�a�0����h�3��MQ�`�S%S:t�|� �|�x��ܕ�n�i�X�hnq�g#�B*a���Z�f=�g�`cw/z�>�U�����*����ف��nh$+���>��G���s���W�D�j{�^؛C-�SǪ�<�J�P����P�su�k�5�f\dI�F}��������SK�)2a� ��x������Tz����=Cuo�賝��d�V�ϷD�=Kfɗmg@�I��\W(�{�p�k��\����J���PGG��}� ΃,[po �wsh��l�[bt,91�Y%���O�O�G�Q��^��)�����f�+=�6z�w�A�W�V�8�2k�]��H�+OtQ�O���%��)ȶe��'%Y�,��P�VY�LA
o��~�mW�'�6�6��5�ŏP�����F�lz��O-`�5��\�^&	�>�%�0`��iEX���5���Բ�G�1�v�k҅�ޙ��Frɲ��5�'�`6�,[]�rD�{�J
��^d���Бn���X1�����˘�D^��!������X�C'��P�	]�ɫ�ˀ�)�B@�(����)=5��6E��.��{�(yȹ�)R�F7�!�� �����bī0�Tԕ�B��DM鏈��LN���>1ؤ��l'�����^�L��
��+a������]"T�6��܋�e9�;�v|����'���6�9m�A)�m�m\J}g+��P:��Q0X�}�4��)A	��2�~̽7�Kc�`�Bt3"q v���S�9X��7>m��z�Ŋ�V�E2&Z��s4Z����G�������0�h	����<Ryo�����0k_�s3NҶ�Fiƺ	̡�C-7_�����w� v�`";����o�L�]k�`����9�
�A�K�l�`Dx)>Y���@?��D�ڟ��"/OߙCA$��㠣�/D	Ƣ�7ȁw[��G�H�$��ݲ'��0��r��
�G��Ο�m�/��k�q��>�� ?��`�@R�xMd%������B��;�q�SÎ�Iw'�	��4��6~wx9�4��l��>p�.���tv�})�B�rg�o�֯����X�R{͕�j��W���d�Ɋ�:�>a�k�է&�"��S8-< �#~s��~ �*�E���C]���D�=��� ���R���v9��������u���?%I��s����a�z޻�2o�,8?l�@[+J�;�B}K�z�28��+�2�F�2A�����x�,qF��RjD>?7{���-~EU_��<fu�|�n��"��G�׳ٽ�Zo�3�� u�33|�-��:�\~�sB������+|H��;r�KWR5v\ �+�D`{Ζ��D]i��F�3�.�z _&�|������Օ�bWʺ�csu��#����o�3M���*��2�dWG�����6\�o��kZ�'K���+���/�&}��U	���!�������[��V'��3������Ә /ô�~Qy���A�/|f/�:y����RR����d%����dL�q>�=V�0�ղ����y;#'�����'cg|Ǔ^G��_JA�q��>��r�ta�Z�HOi���d���rg��=#\���?�+������CS�E~"�����!�漠�m����>�6���B���qL�k�z�8�]�H�߅��e��DB"� �_\�f�Z-�Y�`��QJ�LN��S�G��-ڐ�<������=2��%h��ܫT��2C39��L��in��������{K3t�o�59�B�������H�W<
�|��M��y��O���c�'��&ź���l�rY�O�T�'�I���f�先er���g�X+2#��E�f-k[���̍W�!�Z�ñl�W8�P�(���;����G�� )�����H#taR���O�%(�C�z��MK��	W�N������ĬԤ�&1B�&tJ�b$'�,R�W� ?�mݟ���߰o�R�=�W��r�v_�����	[9j���}H� ���y��rs�&���=����.R�@��Cq��G�Ǧ0ޥ�Yl�pX���&=s/B�g�
!�����\��tR�C`����"�>����N����n����<%6�[481'�M$��֛�����	��#��E���ߌi[��D�y�
��5s�0�X����`��A��k���DV��� (����<.C������97P�O,�3AR�+Fp4�z�MI@��t՜��j�m�����(�4�L�QIB^bJ��fDUB�|:�BJU�:%W�>ψ7ub��vǫm��=^�N�y��0m;�����1taјă��K-GA���d�&�C�����7y�����yҨ�x�Ú��=�)W�u5�f�{� l`̻�@��5��Jћ�d��:N �v7�VG�b}�29t���e�I�Ep���r��77�i��g2��VE�-(��iڳ��I`/�8���
�/JN2�ܝ�:�fb���m[�-�����)@QQ�f&;O��Ker��Y�ZV4���Ǧ��&�[��/{�^����.9<���nF�l�NB��!%�mXĴ���3l�Vɞx��.
sd��|��\.�p� 3�w~ l(��[=�~/�~���6� �=q�b?�5�����2��RU�Y�x[��d����>�֗xw��cC�Y�h]��;�
!ny�E��G�9�YA�Gℂp�VrT��d����]OX-	�H�p�EW�[�g|�:_EN�+��*��	��_��팲Y�)Ѽ��ԩ��ߞ2��{�0N*�уb�s9��.Z�vŬ#+��� E�ɶ�x���ձ�Ě���d\�@�[)k'���n-<���}���-�����+R�ʯ�YD�	��wC�v!LN�]q��D5e��m�#�?=�=G/./Dt5����y��/�}6#���K��m��~B��Wע��iX��ǶUv,FC�3����?���܋*����(r~�1ƌ�	��P�b00<QK3^	PuΔ�1�`Ֆ�i� Z`8��k�چ	礟.�S�C�W�v��Y	���-/�T�'�9AP2�\�̬���ڀ*��1e�8��@�;	���\@ER�X�c��Ag�Mm.3�ഛ�Q�������(}�b�u.~g7f���K^!Q 
��ю$��5�����IO���lKtL�'�B7/��h�%���ɕ��מ[���u��H�8Ɨ���)���K������Uo)��jI��獿o��Ǉ ��,� ���~�A�⓴��W�W�b#�ƛo�(�3�A����f�4��2\�!��1�@I]�:��k�i��bGXg����ֶt�qD2���4�L���O��0k9)��6|rM�7L9E]���4�A焦�Yk�\4�c m��w���yW����b����|�=w(Ҡ�t��V�)E�*�
����!�8!�X R�&�A��ư������
T�&�7�lV'����:�w����`K�;�$,H����%�d��q�Ň؃���,~��0_��)"�S�bPO�rO/�pdl���U�{Ϸd�Oҍo�P�N%��K�r�6�ɻ������e�-��r��+�o'�籠���!� bc)NrwTb�nV�����Sq�+B�4�c��=�3'≐"���kG�NY�w���V��B��$�i����E@iX�����JTM�C�^���&�Ě|$<o�k��sL6�E�	l5�ۤÇ%E�[��:J���N%g}J�#A��MJ�{
�se���h�u"(��`ƴ޾�p-�y���;�1���������l����ty�aS|�~'�>��sv]�տ��o5�������,2�<ty�����_�=VHL��gy�t�S���f�u>Y�#m�*�i�ے3Ŭ:V�}=�WT�;g*��_lIϳ�앚�Q
�]����ft�4+c\#�@Ό7�et����i��bSI��I�p�nlm�[��S�pZ��"]]yq֢
�+�����+ߧt�����ݯ%�1+浄���[	�uKy�练J?CȒ;sJ�)���X�f�,���d�����9�2ǧ��#����4���k��]f�������t=\�G���#�z�x�$Nb����ff`F ΄����q�g.ǩxR\�d�լ�2�����Yx҂��1~sa���VoE�ETY�7����_yQqL��Ir1��aǂh8g�P�_�~��3��mhKP�7(��]�`� 8��31���c�����u�F7&M`��Kz��L�N��vU�X�ik�wك��$+�D���,:DFOa2zȬ���0��S�jF %�{��Fs��&�ec ^a�ڒ+�����ܷg��oc����S�S�K�5�@��[��O�=tم��#��s�j�9>��(���a�g-A�މ@�n�-�O(����mk.��L�?��l�&�$wW�|�r��n�W��ly�Q���Zڮv��? ��<{HLp��%�	��XAT]��<� ��o ��㤖�{S��J{l��F̟�O�~�>�z���~��	K[����z"=�A�z�F��$�9l#��Zg�-	�O>P&�8��L�
Ͷ�A��^��^3:��I�+)+@��P7o�/8�K蝘��{����x-F~�[��Zɿڱ�%O��ۖf�t��-�[�H	_Y����$�9C���������b�W��'�5P}&�����|���L>�m�D��6ǖ�w�LƗh�3�.��T�d�I��n����h{z|Q���%�;t�!|�>1�����+V�}l����Ƶ�d+T.Q�.+����q�
�h?���6v}xM���7zD��QI�|k�B<�7���[JAsi�����
�n0��Yzb���L�v��P��!�7\�c�7Q�z�qDJXᆘ6^H�<B����#Qew+�g��m�b���NJ�(�X�U�kv�8|�u��65����BmE�ڹ�r��g���c,n����xL#���,D��'�S�"�T�Rm��z8���B���,�Koj�&X�i�$E����p0/���:��|��Ɯ�Q8l�;�`Э附��L��$tD����
�%�wx����'9 ��C'I�@TJ�+:���t�F~���*ډs<�Z'��@7:��~���ȝ9�z�N�v�xpҼ�({�B�5�.���3a�ܱ�[���"8�@��txbE��%�V���b@�a�G����8b(p��96�Uz�������$��>C����+4�g��Nέ�	2�s��Xo����'Uc��� �d_=(�QX��W�����L_��M�kS�$e�D�F�t���<��%����=j�8�29���k1�3���N��.�����������t���!B)y���fğ���Y�4����	~���x-�X���{sFTT�t��Fzz��(c�6�F��c6��!���ĮD�T`:�k�,�ܸ��Ћ���Co�AG�S�[�t�$����-����;�?� ��
3w�Cو�£���L��ROt�T~��Z���G���n��N��,�-R�%�����4=�ƭ-Y�:�9�xv	
q�$k����`ܙ�xYFf��$��W��xtFn�4��ʧ��Z�n���=+��rtH�[��Pټ�iY桍/�f�v���z����ޙ�C��������{��K�?/�� ���
M�S�WR z�s�<�2����z߇�@�.���XJ[f�J�q��A�c�8z�Ζ~�ڵcx��_U���B:�b�F,�%�C�V0B��4��K���*�y�}_t�O��q�&��T����"X��pTúJ$|�]s�k���'�d<�Hs���% �6���IN!��تAo�q�S�zX`�����ήF�"���'�Ya��6l��CM�T3�KoO`�⥻�"�j�