XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�NZ�\�Z ��Yc�>�pL(��|�:���@�3��?Ɂ��~�󈷥�]��ܶŏ�����n�������\�G���_:.�v�^Y�ֈJ��v�C��ra.��)ꗅ�����b����Ey;���4�-��Q��l������øa�	`t~�W�]2�z�����y��"
D1G�q5_�%k�hϪ ��7S vR�Ƃ�A���26i�aޫv����4�U9U��.RD�vUJ�@���su*rhKU���ͧ7��?r\
�pdsᯚ+�.�;�wP���9ހP��:����V[�`�(Q� y�x��� ��\�F┽X�U^�'�����`�����¦�8�}\%-?�o������bm=�K����?*p̍_|���T%{�F��� �@1N��$�),;Yza��y���>�o��9�r��9Ox�����шb ��u�S�( ���ۡ�n���ݩ�T�R�����jRu�P����P,e�^�N'�R��1d���A{z�����5�e��YA&ֆ���4B~Dx@9)������+fvT���eF����r'�@�*?�&X�H� �h�`����/`�74��Ŀ������I�x�e�ӳ�a�Xd}��R���(6��z�pI����2�_�>������40Q�E�}��R�[/&3�����z��ln�<I�Do@��T0��Ŏ�;��0��N��'�f-m"����)�^Qd�p_��3�&;͋s|A�=��� 0��(�.u:揭���cXlxVHYEB     400     1d0��M���B]�^	I��O`���k�<~�&��2�觿�L�α��c[{�nL���qI�~��Le��a'94��Ċn����W�J�}���8�uqķ�n33�wE�%V����M��0���g&��g��~7���EL(��"��{�/�2GIR��*bs
6?���ai@�5R��4V��6DNJP�?3� 
����T����M��V��t��ȱnQ۴R��=�谭��<b^\5SZ!�*(�Hf�����b���=��Zw)N�⫀V����vg-
W�n�b��'a� Qf������/���K� ���)����׸�r�}�oE��NЩq����rZ�'����ët�W���٫���K��q� �����q�;���~$%��M���e�K���`�{��O�&��� iu8���,gv���/���N�ѓ�-���j��Uw#&�\�ͺ��XlxVHYEB     400     130�je*ޣ�u�����A�P�/�z=,$�EW(�t:i�IY��Ս�bg��}���e<g�赦Y�k%�i`��4
��Q]F�5��qa���D�a����D���iC}Dh`�)N<�&�{�[x����齌��
�Y�_�슄�\�l������3{���K�yU]�g��������=û���\�.����?,�LO��L�SP����P*uu���D�>��lE���C�*�S��l��TU!� 8�d�C	�s�:�0��q�'�^]IWN&��j���5�4�>6�p���d���?�����YH.XlxVHYEB     121      90� �$Á�"��H%d��e>z4�_Jl�.�ɬ6Y�[d�wXyL6���sǎ���j��C���B@RB��:���L4���{I�<�2Es���jW�>g[1� �ftd����QϪ|��N>L^S?`;��d���=