XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ǒ(���K�4�w����a&���]����?�9�oA�cY9�pJ�Ô1�"1H�*�{2~Lg��R���$��F1��'iJ,`�Eb���Ѯ�W��ѥ$:�d���'�4�#4�^_|%~ y�.����hN�S�J�hHB���u���2�@0����{SN��Ax(�eY~��ґ���Gb�K6��^5��T�^> ����x������V�:��e�{��w*7��r+������Ih�[b���ڜ�A�
ƣK�{:S��X-a=XuJ�qB�m$rPb��
A��Q��� tI�����o�X���@��2���[f}N�>h���$�;����`57��>��M��N��<�������>���$�W��C�;i�;wնFl������1[@��[S��Jeܞj�J%;PV��ѕ�^�YL���V[�<8E�˄h�o��?��+F��C�:LgIPlY���'���k=t����V�d����){�KՂ�Vp{ !7�}[$�
y4���lDӠ<u҉�Rų#���3m��(^�iCz��jn
�G�1�����i&)3n�|I����/Pӫ�NCW�!�Rb8��4T��H|)��.�1��Sp���#s��?�~D���U�5~����J�b�`$������>�.F�A4���i<�˵��H�c�������bG1�7��an@
�9�#�vIbAqh�G��-:Y3ћȹ��pa�#�>����9+�z���AX%��|��>(�G�"����XlxVHYEB     400     1d0e*���9�A!G��Bg�`�_m ���eӳ�-��X�.�m_	�mIF�����tňAb\3/4t���SI<6,$���w�k؇­6h���᜜PΊqO �����Mu����M��f]P�z_�.G}�=ܚ���\�ɰ�
�RS:Kpw���k �C���ԍt��������tf�f��tlw�C ��_��~%z��LT���Ge�YkgTW��l��h�z�F.��4���"ܚ���<�8_hx*�P�̚��aU-l9Y0�I����@$F]���دi5�VPܔ NSŖ0\�X�\����X�q;�?q?�yR���[�L��j$�vV��q2P�s�gP�Wߪ�3Ќ'y���N���{�*{`��Xr�E(l03P����z�>��q�-�\�}�x՝=Xz5kG�q�77iFCvX�E	\�n����H�А_�U��b�z���@����)�>
VXlxVHYEB     400     170�w�߆��R^`�O{�v��"; �$��`Q��9�F��ܛ�!�K�� \>�ot�|��;*E�TA8��*�ˬ9�Z�Po���t�y^��K���@��W��Ϋ��
"ܖ�� ������k4�s�������,e���5�w��L��m��gCX��mWa#�d��J�F��,��6f�o6���}M�o�l�,Ŵ�/��%��ڔ��c�N��N��s)>p�2���ѡe���'ۘL �\5�@0��Y����CFK����Sy��&MMhDS���d�m�7���-��((�Qca��t������:��BD�C��`#�ĭ��+
�6��?���x�
�n@dZe]@�a�+��!XlxVHYEB     400     120��H�
Ƭ�5
s!4Ǽ�A���ZXo������x`�I���˝}�K@fqGN�^�$���G�����l���i��e���Р+M�'o��V��V^ �{�Y�|�ڳHЉ��XR��۝��pʰ�p��FcF�;wU�p}0|*�X�� ���&�W	Ũ��&Z�	L�=�&��~� q�`�)�Կ�Q�roi��("�f�ANf�i?���l�v!a��/��F�O����#l�R�j��JF��}�_L
A[�_,���h�]��34Ƈ��A���XS�r�(XlxVHYEB     400     17045�*����P\�����eH�/��%�4A�U��{F.�0����d@)��4��Q�I3F��l������*���poߚ��'y�鵌�{Nz�ة��X��������:���D���Ƒ�Z%Z�
���P:�ǣ�����yH�R3Gy{�f��6�q���_��س��@X��c�Vm�Q��DN�|���ɲrgnȵ���h�R�c^���hy����w�{7|�l[�"��}{g�sֿ���\������-�%��"�H�<�u˻�;C>k�	|ʳ�1W_uԜ�BE^�"L}��ҽM���A0�׾�=��s��g"`ɕ&��H�5�W�.%�� ~����� �����)�!XlxVHYEB     400     170<<Y���`[�"%nn�*B��<��	.o��~�~L�)��^@ �I4��N�jQd�j�<3U]�@<Mn�ՇC6k���^$B	�Ğ١=�s@=�=�G�.'&Ef�"�6x�s��H�9�j��F{|����ɫ�:�n��niB�+H2�#��">ߠ	O2��
4}\R��"�eP#��B�v��1t`5�x#>T?���2
������m��ߐ�]�v߬�1ͱ�SDit�Ө��.�y���dI�ei�H����o�����U(�!f�^�}���&��X�qLf@����S��xt�A\�-�J�\�jy�E�G���;�'�yS������E�m�E!�j�v���b(�FG!\NrT��@5�4�OXlxVHYEB     400     140l���$J�<Ǟp?��<�I�,��s ��6px����x"X������=ܦ~��D8	��%q¤�G��ףH̞@���u�s���a��N� �Sx��D��J��zf���o��_�RZ�^8åxs-)h�����!��� �N׍_▾�[��/'�ŗ�Z?�])/��Ś�����,:�\��'eb#e�7�{s�MX��4����uͩ.��z�h�I���%݊h�S��x�]�E�:���)g�!~ė��~����3�Y�
��F:��c>������B���k�ʺN�F���~Uʽ��9<�It	����ڿձXlxVHYEB     400     100���ݩ�jRJ�W���Rrk�۠O1����u>8����bFWo�����RHI"y	$���z>�SV �������r$�!dz�����'���w��I��e��!�88hS�R/�;�.���>�����8��>���f�Q��m:�I:b� �;vEX�\�{i��F1鹝�TVz��O�j���V�V*�d�����c!Y��ث�zl��Bu�{̯��,�O�Lu�z��1덎���P��U�b��8Yh�ݩ�tz}XlxVHYEB     400     170_4p�bX2@q+�!g�'��-�Cf�+�:����&ZF�2�:�����Q>���2c#?���^}��?4���$}# �D5��ݎ"Ϳ��#r߉����k�su��'K�����Ӧ�R�S(l�\����z�#����2$��
�A|�G��ǉ�;��x��0ޫ�؎�>�82���
V�P�T�o�E��ڃ-:A�cU����q�m�%Jq�g�(�h�v9�(g)hYa2��{:Vj�������
����	�YKV���B�����O	��s�����-Wf�;���%c�Ú�u��`����R�F�%���M�n8`r�`U������2��o�����y��G�O�aq��>��	������%�XlxVHYEB     400     1b04���{�^OIQ}Pw�,��SF��X$�r���jM�������f��e�7�t""���	{��}}��e�*�����,t�1�/4
��P�W��}*�K[��M�Gz?ԭ`��υ���y����X�c� d�<ȩ� �$�S���d!@���/Ҡ�R���G� /A�9{�BR�d|�e�@s��!���5�>м�xD<�U��-2�L�%g��x�u]�UIT��#@��n��� v��s%'v����0���%���9�8֘g	��t�O'�6ѹ�	p��+&u��1ef֎�Z�ہr�7y��49�E�
#�R��ker���y�|%�P��z�,i�t��S����).7�KD�,j��@.m�n)U9;2=��:��c�-�X@B��BI�J�:��wt����XlxVHYEB     400     160�h���ˡ%�h�V �Y#nj���v�H���~��F��_57Z�Ŏ����Iq:�iM���ߒ�z�P+��Z;�͈He���[����]:}9'#�$긷H�.��桂��MtK�j���>\��c�a2��
��+,��*t���WRhF96���G���3N��w���M�s#e=�������yR���|H?���x��֏�ʪ=����])Nd�󵿝��*F#�TB��)E����tk9H�b�#,itui��x2 *WDN&�/�,��("E�:=m�bZ�o��M���7䖲�<�e�1�OF�+����{�z��z����I	7��;?���0���wjT��S�MXlxVHYEB     400     1d0鄍�9°SB|%�KWb���Q���3-�( Y��/�����n�Le,�e�x�YX��lv���u��e$*"V�֧+ w{�dd8}�L�{��� �� �T�t��V�:�KeJF�&����b���>t��"�RʛȗW���N&Q����0�� B_
��dú82E?oq�".W<�Ѐy$���o��P��N[lt���<�x-�FL^�mk�]s�A/�oM��V����>R~��%��~���(B]_��T�i���Yס��2�V-4�)QM��t̋�
g	���ȵ��{� ~��j�ƍ-��" 3}i��^#g>��x]wT��+�Kd^3����~/0�)"͖��c@Fs�VέsVT���EƉ��������B�$G|:�pt:bS�bɜ^�|�(��s�Ma��[6�D	�� �'�N-���ɜf��[́֗����Q`����s]��5�XlxVHYEB     400     170Xnϸ)˹��b����.���*����Й��$�4�~�R�����%�w7Ir\��k�	��؟���'�@-�FL�v��Q�*��
X���M~\ܵ�؄� �����o��+�=����\&r��ܪM��������c�l�0�H�w�����RĢ3	�����܍{V���ܧad6���!U�����)�;�r�5g��]�J|�D;��Cq��E	��8����W�-�q�p�-��6n�*�����D)G��ۼQ�^5���*$���8��]t+ �ʌ�VC�5�[��s����8L����K����l�|/1�Prnُ�����Z��;������d���CO��FV��j��-�/��XlxVHYEB     400     160u��ޏ(R�0�n�YB߿5>��'����ii�����]�L�	�E7��l�����"������̎[�zO%��+�#�7�J���Di��������c������g
���x,/�7�[CN|*]�Rv̥o�淌3cZ���c�"��>��JÅK�FY�~�$Mur!�o�j���$h��1v�y�f�#R����I�.��,G�20N���V��}��aT��)}r~@�c��L�0m�;���,|(���ܦ`���2��]^��u�=�ijeq���4�۹���ե�MiIZ>�!�I����O����2-Z�&p�5-��l|k�/À�Î=�
XlxVHYEB     400     180�àA�<��pP2xMD�$}����4l��"�P]�%�U��a:2��P�H�T�-7x�MI���]* /˦@���V��~;�r���x6� �썗:�l �5,,.MzK¢��BP����:��y���~��)�dlOk���}F�����ݾ*9�k|�gj>O�M�I�-N\n1��a�P�hL����j&I�)�37���j�G~n�s���5��C�$N��y�J�_	���l�a�pg6����7L���&$��,5��Oj�@;�+�_��yF��;���4�; �Eі�q>t�t��3q��^1:�;.���-e�ɼTm���xU0n8���*HC,7QL��� zt��Ԝ���`��]�k Lll�y@����XlxVHYEB     400     130s�M�s�9<����o}�Y��0��^mOᑖ�����'���$���2i���Ī3���F8ؔ�3�VH ��뮖���u�G,'���%�@��B</�FL��Dt����4�C��ؠBH���
;)�MO�g&��rj�9�a����DC����k�{���(ͅ-&P�Z-�@�R|O0�F�3bȞ���l>'`	�LZ�J-+�4b��-P!�� ��ub�V&c`֮�����4q؄��9E	��'��Ok@^��b���H�Z7�!����5hsC��gE�:��@D��,��9��pzXlxVHYEB     400     160�~�ڪ�����۞y��������7���E,d��\jO��g]�`�R��?nn� ��>X3}�:1��j�@Za�x����  �}@ �Z7]��i��.(C"B��!���V�cX�1\���\�΁+_G�2�=Xi@d��\�lK���{7��"�.��/ğ�Q ��W񫩄iH;v(��XՅ���Vm���ǋ۞ш��D��d)E񲟞N�a6eP�S16�
i�/�̾��|�2�r\�hop1�q{Y�,q��P���1���>��4+�$��Zߋ��)��$4��cP�R��\�LV2"a<��FƦ��MY�����!ho'f����H���}��g�;&5XlxVHYEB     287     130�6ԩ�'���C����)��~3���xb���c�j1�B�L8��ہ��$=?�z�*�IR���e��a�X#�̪������rn߰��H��Ԗq'�����
 Ǆ\%�xX�q$��Fo�V!V�azV/�q��f-L@�Ѣ!k��}|B���u�� '~q>6ʄ'����f��+�B����'��]L�{�k
���2D���Lcd��C����a�[�(�W�)bd��}t �#%���Q���In}��g�\`�Q����O&寙h\B:?�KJ��`s/BUm-���P�EVE