`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
SsTks+RVFdcRUmDEZhjAs03cVB18XmCDm8yDg93y4jgjXurgXbfDOztYZ2rt03pTkeEFiY4X9PD4
crAeR77sFct3yMdXWgI60cRWdM6C9eq9wR1d2NWvRpW3/3ezT9r4n+1Dh6w5x40WI/4sE8PPWv3g
yWQsNBLyb8Qhk2t2Huuqos+pQCdSJV5O+uIefCkAX8c5plPdB1Hw6AZ53IgkFquIx7w0MCa+dERk
aHgC/VamCYS+SU1fMoVxh/OMX8K+xnt/kfy9RW5d7/Qco0jM/Se2VsfO+AFXTXKs1ADNbw963YZV
qK0AOPmFmKBLacjyNBCT1F8HAXSZVMCcVNhUdoFtXqt2+BaokLy6S1hTVW68lp5LIjhg0WdZyDXu
x4iSe9zYNKVaPWKMz2YoGeubIG8XZsUMegU5n5Nwx8c5twrmh4Xa/abVGObij9D4k1Vz4C6K1ofJ
GVID3350IEJ8J9bWsYCjeCpStHWpjcZrPBCpf+EEtvNp5dXwB0Hq4WfqJnLNpt6W/klxIjX76CRK
gofp6aZ+DaChmOPBADH9o/O+gBVO6rl8ovWIJHgl+zq06+dxvez/ZCfjzgoisC7pYUMkJx6/7qSR
z7GCdtQXKSZTboV+62KMt7irNKnu6f/tZUXjiZQdhYHfThq5dxoxk9JrmbGzKsKqsdnOhcQggT8S
B6U9H+V/PGrXxg1PIWM1R98YaxooRqaB9vj8K2oEWD7bVnkGp71XuyfPOH09XXbvpXbfx1g019yH
YgW6wNVCbRtC5Fc1mGnOoD9zLMf+8WMRr9fKPGbDZfh/xezKy9BVkScoLMP8zwYFj7bbpgLDNrZx
uE4bMUbBJU6vJJAL3g3JC+owlupaQ3Ul4YjxGMJru+APeJ3qHCSx2nyr/nA9r7DUBBFo0jrAUItH
ja+uf5SsFXOkZg2guLrkaVm3FeHXJPsGzfoY3SvmxAkoAq4BG2mYPjXh1Tv4vRmurHeWSTi0ZPb2
uDk+xy79pO7MNOV1WDVXt1TN5Fs+oX902v37MTMYClLUht/vvRRp6vr7g2xtb1EJ1QiENcm/tRh8
zUeg9CxtP3kYHS97h1yRjeXyeg6F3cfEY9fJ+w3YObyTqwFCVdbdml8xUvU95qkQBa2igiTTtam9
m3kP3Ofc8WIuK8O6g5taK9v2aX5Cuyc86aNfEohhAWNKJgrY532Nlgxy3W8TYUr6F2PsJp0mR1Fk
WK1WZeUse0Wyco8TiyMEoiwmS5FcLNr78/GwRFcedhBwXKcQLpkoW5c/sZ5gW2lCOtBS6Ohgyiii
y6cdlFgMCVMMr6tv8XQ3CCvvaqIMI+6TCDzYZu5ERTIBWxu/de37ql95Kqy9xlmSk506paPuVY/w
3l3QoQVJb7qOrchPala8ue2BD9iiYkZaZIy3vZmYV6D1+b3XjLNm02+P4Y0KtgBhHqAy/tG38t6q
UPBic+Bhd5nYSoR5lxkew3tda+XxDXrHDPOFR59kfOHJibZu2QU6ox4kOqLFwc+yJZTMcTzDQkwx
6JgmvBXHSc3Y32ay6TjsY6rceOdFDEIniW2cKFtCeqQf5OoyuSENbWyB5lFf5SNyfApwl2D7tG4b
04VwkUu2iZ0c844VICqgIv2cAbfDjXWvajQKag/U3veOA4AVlpCLE+BhqbFbScC0uKqT3eL9LA5/
c9LbI9WpogCBElo9G8N9MYm9pB/phSFgyJs+BAXZzPGv7xhnJuPAPgLyhh8WJu3s+lsaI/xx7osR
M8e95XH1ndrR+CEgUNIlr2TSXKnXgWCBWFuVa+ChAtA5LWqq8xHU9TGOKfkVDPkqdxfqYMlb+59i
TrCw+Ubb+Sn4ZJDWGBm1X/vmxarLXKRuiHWsoU+t9fB8ApfjqYD9nIJnUbASmFO+f2ZKX2p3bsTI
RUoNQGOGNuB/xwghcJu/Qzt/W2kiqQIgDJPxUeSGnz4yDd07Wy6togDgvBRfOHQRVE1sW/3mVZ+A
M+o5jeXbVPG0QmwfY2AGBjHC7i9+0DZ0cP01SqEgqdotaNqFVqSD7/gQ9rbeGkhQCJESlUaGDQ7/
5xxGVH19J9xtgD1weLBgrQ5qhNhxynil9NrZELhxmUOqlf+W6ycES/5z8h2EZYdILzGUlMv83hmL
+3Gi97cdjtVhr6JDyJzKubr63xFZcqlzNsHfUp6OU9zjP414I54+lqnx/g2fzXXcaTx9+jRPD/S6
0iHHWeqlGIX292d5dVDFBQFmm7UbyZxbKKvNh6M3E4xV7SDNqmJMkgpMPXLVhBXOJ8ph+zAd3JAk
zE+VUau9aFCLh8juzk0XQ8TQbAic7AwJvlzT7KqzHR86Xyz24fYJ3aWAra1vpnjiCYe36ZcEPvM8
Y0pgancKgsWwOD4B76/86n5eyg9Dm893g0ieLsGLmtPUEcatmiZfDX6g17eB0Q4CJD4adGNqZjxt
VQaVWDBzLyoSjQCxGnRfWwnnPmheqNx43tQ0R8NtwLmHuQcogHBFaN8uYYrNaLJLYj6isU7s71Ff
LXu02PaKRYKlqqyP13B+pr4hrUoCDW6bBcBxKsZThVq1YGa7EyxiPW/VHARmwqXK6tilYs9550Gh
3r01SJ9lLeG/rOmcINBi6hAfu0NXNIM53kmT3xN0A9OjEVu0EVyAJ0YPWFTZVAaXrk1el+iPklPd
Plh8u5BGdIfhSbV+mnsqyfmnY4Normy5AhNQkCaeV1L8+T//ztRDB9Bd8w922L6zvsTWFnfSCqe7
apiZper19nxHIDiWBGX7vNlbwowF42ZYpuQCDrxzt/PCI5Mujs/E6BQNtcJkV6WUVhmkO7KvJjWr
mvQRyh9ysa8TFIuQ5GjuiYB6VpBJ7w6QHM+CjKZWHfUfZHaRHON/WHMNIPIBz+WqWNP0BT5oZiVf
PiN9ZFJLug8uz5UMlN5N+AvIrnCcg3u+SVXz2H0eIPYLuxM/iFl5Gbwl12ijzn6Q5ANNxwVGkVIF
aciVcMKHqEV+Re8WZ2KyiyTqa1d/z1okj3fpl71Juyfn7f3B/0Bp5Ny0R7TrCkgCwxFbfJycJXLV
OTnCeNBTqFr1J8V1kxeMuNAEYMcR9G9ieR3P6Nj1LjjgRSPb+MeMtXZegDOyi1hUOT2wZIENC6bS
YfA/Axq8kHc/yYgzGkI46yEN8mPby9iEpBrsW69v8qalvAC5nqJrRkREaJFTAnZJq7Y/Avh1TDBc
S8relUptIJPPgehx/Nm7m8+1XlEFIlUPaomyxrLZ3rLxzrEydk4QDmu5N2MTnjAZq3RcQXNQVw1K
NOYceGR4OQPb1Ywqy6f7svZgdrI0PlWRL0Uq3yApJLnAblSPSW1LblZlHfAdmm0b/OVAejlxnLXT
4YaYScYMQz/5f/dw8phfXOcvw10zor36ZGhqQT44TNW5rZW3EHL+fdxU3j9vt7m1v8iFmL8pQIaw
TOv2RLkT/A9w2ItpMesUsFRyXzcfQGpS+Ecz/UcTlsmDa8Usn1D3t2RHfDsGq7MZ6QYo3mTHgyWN
QWrIcYqgf/fKTZ4IP/4B387H4RIANb2NMSWfrWeG8ojMyEtszyzVTLq57bX0mRqQnKgQ4rn3YO1i
HXoZWjURex07FLIJXHCTBZ+J/20QVMFj7w5xhtO8xNBrfUk3VF7SG0toLuxVPfnRFxONrI1INj2h
FFCBQ/fwERlq/echtC52txc+42jskP3/IX+EAfit6ZQ8KMI4J0O6ahKc0wDpKtN6B0UJmGK1/4VU
8lb+qWDEy4rGZzaqO0TvPfPdbn5zS2UpHNvtG0ur1ausRkUlFef3W9SuXFbmiQSBD7GYx/oJUuDE
iuofa/fqKxTlFaLubq702Ph3l3EZI0l/FvKQrm313zN+c0LLNAvh/nOJkGjwDPeAe9MW+iwzaKt/
urncZ/yER+UWiFqnixe9t5KpQfzmim6kXHzShvN+rAm2n3jGi+J74t/oVTRlgFqK1hzF5Geg0mX/
wElCBGP8+ynW9AditM40XsEC8uwcBcTuJxH47kRgzw1ZWbCmJGjl2zeSlE2zjpyK9r6WiPL+n3ED
FkHPlwcdu/pQ2RbOeyPUS90qGKFUcVzb93Hgawp0WXeM9WTZcn1GaBnycCOjlqfrmeAYi5wJAkOW
3Ae/RN5mHT6ExflC91ExJzqqIMtjUA+fCFGhjunDO2Ab8j0cmFgAq5G8KQEliAeq82tHQziKes01
xt/p7oa5LvPRU5f/i8xj9GYviJ5gCjjqxNFKeCqM8ZEpnGT2zUUZEZcbEYqhlwEZJJ3S+3ocXQiF
bBfsjqbi1Avus0oLeYKlLKbReH5HNOjFRuubUgbtb1hq3NoOd6gnbjOAv6HemwPOAHF/fTMBxV6w
Op9vPJ7wGGmlewXYIyxyBTe8NqeU6Di+hxWFpqI2VnHmCRD+S7blNMjRkMmJ9ETLYD663gJj9/8b
Hu2aIvnT5UU90JppZZEQWnyCxlH1ccV9r61R96LpYY+nO3lJtfXllcFD9hqU69/o7i5o1wGBKUNS
XbfcVC2mQB/WbAFiyiu3WzzJTCF7j75jy+c/eYwijeZ4/oKS6j+0mLxgl+1QF4cmtlf77vBKxpu5
tUWVHbb9zr9O6+52SY3LS9vUyOj2hcnHs8Sa12S7Zquxo2YZgqX/wCpMoZjrJ3DRZHVdEu5UmJOB
BFV89nN/HxkwrOG474Hitairx4ucqGH8x3Q9Tpoc+rF2BdyGxU7fpy4AX7w9NGts9OcNQyAklFrO
tkmyEeTuW70hrfusyE6FncNgBhH4pjA3fM2wDTr2YYUeX5XY0ZNRi+i+9ncQl+i+e7cXICsRTl65
/9XbcXirryW9IuQj7gsScMjXiBpnM46lBGhXWuwERQ7eWYtfcs0BA+EQNWYaW4sm8ArkKg1rAcF7
dHVwXtjIxDK6iTV7eiXm4Q==
`protect end_protected
