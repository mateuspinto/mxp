XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�M��q���C�geQ`����@�ˢm)�n�{'����'��Λ�R�A#�j4�! ��Dщ+j������,S���[�;�]"-4E�p�F����z�-�B���6@o�"�ئ@:������}�܈�Tz�)`j�_��sp�|�-ּ9�p(�w���E��>��2M#�2w9:Zt��RK�K�α�
ҞbD0�����M��s]��Y��O��	nJ�5D4U�����HC�� �39���Ha���²�+�*�3!�]�~���=�/��h�W�4>ֿ� "�X^�B�d�޶P][�K���Ǟ܃��㊍�и�0�'�v��9Hx[(�[���g�(��쓒&Lll��2F�� 
������U�jZ�C4�j���x�ٵ P�$�M���\�kV�� pa'i��O�e[���j+)r�Y�vNl[QPNߺ��X�(� ����%'"Q�/��	��>�K:�y�4ӥ����Y���,C�C�j7�哊�t|C�a������]���bU�2�����%/>�r)U��Ю�P	�#8���e�s! �+�rΆ&pF<���>�k�ѫ`^u�O���9)��2x H�;4֙��%r�%�e�ժZ��6�v��J���J��=�0�Y���dL�����P�W~D��nH����c�[��j#�/�WVI[1�����q.�>��6�(b�P��z��[xk ������m�u��M�K^�X�m�˙�}��!�2���t�����XlxVHYEB     400     1d0�	�WG!�a�2��72�6۷�n�H�����lL5�o(VV[�"]_4��D�# ^�q�eBb��Tf���o&�W�Tp��Q%�|E9;д��+�!Τ����J�L��.t�R�H��[��A���U�$���$Y�j]�]��Q0Z@6�Ԝ��w��K{#m��E�R��6(J�%0��x��Xїڐ+��3�K�P���̖�^dߎ�n�_��Q{ �
�]3��b�wzXAdqTE�돁X�rv K�1Ļ�ډ�Zj6?��R.���jkd�~��R#�:�j�}�>�H-.+F�e��5��B�bE��`�ֻ��@X^&0�W�J�Vr�-i�p�1B�8��YXҡ,c>�k�����;O�&�Oa���y������|��Ս��И	�����*�9�n�WV��`+D��h	#�l��~p��A��* ���u�xZ��#n���7�cs�U��XlxVHYEB     400     180	���A�]���9	I��q�&�x��s��m��](Dq�"��n3^�.	:��ƾ|��Fp���T�jEL�]]	�kAf�-�zb�:���A�����-t�T?ajl��Iы���m��X>]�Q���
���S�0��#f�s�s ��E$$���Bo��og �#�ԍϫb4�5��]�*쓶=��4^u4�jـ.��弻U��]k��s��1�F���-�b���PY:�e�d�ň@�C ͅi٦	E�>I�"*�bg)��gY�����#����g���uΥ:^x��!?�l���A�%�BÑW�Lp�����˓����%�/L���T�g ����a��T�#�Ζ���Q��l�2��X��M����^�~XlxVHYEB     400     140A2r�@>ƙ���~ u��;�,Ha�����F!�wg��>�Bݼ�&F�r&m��P���wQ�?.e3���zL����)��@*	��n|=� �Xz5�p�^�k�p?����Jy���� �/>�P<�j�ɳ�C�xCLn���m�	��"�k0q��$ĸ~X�,F��YH�cBɛ(��İ�6����t��[���J��+:Q���!�榎��M�ma22�U}��}�=o�S��n�W1�9 �#08����dFC�V���g%C�D�z�~��-����[�<*Gu�r$w�g��gG�8���e��XlxVHYEB     400     110���c,Y[��T�B�g�W�/�=�z�����ht��c�`z�&���F '�\�N���Q��h��U%U4�"�$��Z�d$��6D)�]��	�Q������$�n���5D.ݏn�	G	:�I߰�~f񗣦F�FS4�<p�|$���\�Ç���6B��L	��PQ ��K;b�O�8 ��p͊�l>�Ľ��#����w�V >��8�J�8����Zly�9X�9%�4ý����N�O.@މ��8�)@�Ӥ����5[XlxVHYEB     400     130z�=�����9iA����.S��P{t�:�$Z{�����6�J^�@|��:1���*)۬O�<P׏L����'�Tܧ߳Z���H��[;�n���d�ܩ�'YV�k��m�mF�2ᄸ<S6k6Pjgd�ԑ��ގ��F���WQ������#�e�<���^�\�����IN9*��ߗ�Sl���D������oK\*����V� �A=�֏��O��F�BP������M��I�g)����׽l;���|wL&����c.���
�&�ܝ��E�H�5�p��Ci��(Oh�3;{��nXlxVHYEB     400     150��W,F.�����TϏD'��5�z���Z����|�	���K�m B����u�
��q�<�K���8͗�)�J����҄��i.ɗ%EK~"2�8�(7)�[��^hIFz��*�s�y���l�]�$��%�C'ɑ����&q��yA[?��v"����EB�l��m���^�]ZG�Q�ve���� ]�u�X���,�s?ˌ�fl�x��u��7(�#^�,n|ȶ���(XE�E�r{�K��1P+�y����F�&ѩ�8�zDs[�WQ������>�%8z��;���ۊtT���K�4�{��������!O�-�-XlxVHYEB     400     110&�O��<����a�z�D:����zX�J�Tf��y��)���d�p���s�M4%^�)?}VHq���c��d�1�,/"Exv E�U��W�-��QI���ּ�۲�X(,�B�����7��{�rɉa۬l,����+g�,+xۍ��m�l6ۧ�9��iOz�{.���j���&�4��}/��I�.V���=|��2V���ׇ7�E����Wd��L�|7i<��� �B  ��)g8�Fm�DJ�I5o/᝗�mv�d�h�5�H w	m�mPSr�XlxVHYEB     400     1c0���O�b�5+bPS���Z��v��L=�(��r�v�����.B�t����K|O��~�S��m�_Y~:2x*m9?�1pvan�Ũ
=������2�~���|���G�c�TO�W���Z�EoO����ѸðH�V+��!H�8�S���c*i��| E ��yF��,��$�-�|�C��ț).t��s�̑u��;��foqC]����IsT�b];a�j����è/a�aб��8����e~��ܾɕE:�Vg����泄�g��Zq۫y�v�����].��_8�B�W6#+�����f�l1ID#����5��	���s/����xù��ڜP?r�4N����~<j'	�-L�nPF)��J/I+Fzܠ�����b�)z7�<��y�Bfb|��*���v`��,"N�Y��K����,\d�Ċkt|�P=Ol7]�5׼�XlxVHYEB     400     150U.{C�g��ׇ՝��t"��^�i�@���8�m�<�Ǐ�q��O��q�qjpPL���ԑ���dBS�>nM����j.-�e�}������4@��3<� ���TN̕�O�_clw�D��lOO�Q�HC�G^@`������8��*kC�+��/�+�KeӰ�����s� �p?^��\����i-b��F�p��~&�U���&���O�s!� ��2mU��hW�.���ʈ��a���qk L��._|�'r���&Ѳ1X�dm�1;Vk�H�f�v�G9�!���ԝ���c,J]�+?~��OtkQ���bp<>�����
��A�z��1�X�|DXlxVHYEB     400     170�����Y�K�Py��a�Ck����1��n�[yi�У�i�����S���I�xh~Ie��/$�E�ʕ)�9��)n�Dp���������Y� ��wbđ�֖W�%��J:G^�_�&����{�i?��L��t�8�X!{��䕉�H�t�3R4��p�@�E��=���y@/y=�Ow^�],#�X��6���~F2�O2�?��r�	?Q�M��D����۟㌗���<��00���u��ؗ��.���=���u��Wb�4�p������Va��js�sG,�w����ɦ�z�o/D��IP�i�(�b�����b����cI�J,G�1�	��5�d�� �/cGC`{⑤b��XlxVHYEB     400     170Y�.Ζ�2%����2[��*O������C'6�$�F��p�T�O|~ ���?i�����{�;n25����b2z���`&$����Y�hE�a���Q	�����&U�aL+�l��7+�$>'��~d�R~/E��1�"�z�Z&��&oY��
�n�L����9���eD��,��.����;q� �%Q����BG๑h�������S������J�+�4ńʥ8��эl��o�ѥIT���`uhH�	}�J��
���młuE�jW^�5���8*���|�º(t�\���!b
S��y��hi�O^�P)����T#TV��x��vD��~m4������#.��c�Q�
~�kUHw�B|!��XlxVHYEB     400     1f0��W��f��nN���m�Ҟ������Bj��&���X��̫�Xa�fi3�~K�x�W���
F� ��DX���t�;����p��כ>�w�z?<]/yy0dtD�4�ϋ�O�7�J�-�/����`�� �!��"#J�h�MCMs,	�8F�8<a�����K0Շu%����ba���㟓��:ܓ�P�SWlP���>��9�w���Vxth9�v�n�@��K_͛�[%���f�ap�����?hI#O�=�Y>Y�1y�a�X�1�s�;pD��=�	��Oj�'9�a.h��j˶!4�8e ��x+�v����B�؎e��5/�N��c3ʭN�Y�{�y��1Z�TEx6����+A|��g��|.VQ���bg��EZ��Z^�2v����DE:"2�&u��UΛ�ݧ�	I�FE�+\V����2�x*��X�K�VVY�iW�Bl%�h���R	{�w�j�7�n)]h�� g^
}���k���z�XlxVHYEB     400     170��f�+�;{������(�}n����Sw1�c>f��\��^�Ǉ-��'DZ�[��v�O33�����T(&�)�	~'��?i����ߘ�b�mӒ�meu0��	2l�ʝ�����,����(t��L$�V��L1 �퉉�j�Z}о�=F�^����4:M�[�Q�Eȸ�A�F 
&��Ho;�����Q��yds�J\_@�� u�ٞ���K�rL LrX�M����jL-?�^���O\��� �1�4X����c�;�l�@��_�r���2�$��y*�n�bsPK�yᗰ��w�qbU��6;���Q׽�lt��ۃ`s��R�y�s)���y��� �8��Ҧ��bw� �sXlxVHYEB     400     190�4G� ����p��E�����9O{�Ա�ؚG�'j´���04kj��"�jظ�h�s��$�M��.�w����0�a[%��Ռ�Ns�C��4��d�<�xZV��n�T�>P�[k�{�2�{��՘~w]*X�/>oԮF�o�����9�n!�wx;k�1��б���Ma��j�!%R��f���k���r�C�ir�:Ai��a�d ��3��>��'t���2I�y��x���Z�%�N����)��C�}��2�9���h]R���?h�D^��1�B���㉺4���j��ؾ���P��W10l�7'؅|�KKވ�)D�R�Կ�+JJ��u��?�lt+Dhv�"|D�%�'��˟��h��5��X�U���Vpww���_XlxVHYEB     21f      e0���%�|�~.��R��C�IVJ RЇ���D? ��b�S��y�8�v�ْEzD����!�?��φ�L���D�{|�nJ&K~%N��'��C��L9�U{�������E�����fz���� ���H��>����p�﫾�{`��i�P��e��`�l�`�x����z	X����w���#��ם\�V9�ƾ:M�K��ۙ�.��J��v��\�f]2?�;