XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�X�KKX<'�����^s1��ܚ�Z+4M���3�X������� ����)�:4���9�-N�Sѿ�W��G��&}�gX��:O��5�]�������e���%N�]�ּO��ы��;T���`�F"��Ǟ>>�&8���f�I�f� u��<�HM����E�H�s���h�PGG��"!�|I����U�峨���=�a�'Kz�Ŏ_�0Ζ{������׸��M���}�뛉�t���ta~���Q�t�ێ�;�%5�ڝ����Ԭ&h�3OHn���l(n��9��E	a��Nc���x�@0,uq�e�<�~��
�D�ՎD:��E��A�[�I��X}����-�n�^�)ݩE�s��@(�XD���5X���!4:�^F/^h.�ΠN��y���&,<�D�j�\�7��sQ2�U���Wo�wY����%o��Guޔ��Sb�L��m�wP�lLI��e�K<�•� �\�X[.�	%�qm��^V�q�g�|���[�\/�Q��Ms˦�oN��8��h�����ذû�)2-����o�3�eC���K�����X"]�|s7}_D,���0��d&&������n?'o�8�r�Q���ɑA�'�O�4�o��X�4<ݎk
;KqW�؅���U�D�pu���W����G=,�2x	S���o3���_����6n�o������MR������!E�B�s�S�2��9`4\�i��?h�$\m�Y�* E�ezٍ?s�o6,�XlxVHYEB     400     1b0��޸��K�߼�(�7�T�4�=7u7i��
�<����ѦSwM��\ͣ����z�U�����v;�B8	�a/x���}jw�t�J ��ix���W�*�N����81{��ģjMZZ�'ȃ��g����i����]r46��M$e��V1r��HF �L�?��aLO,�8"�ȐE�	�ڶd���{6S��.�J����$wo�����Y��s�f=MH���Po:�����f�=/�+�:��"=��袾���p����
�PkӤ��8��s�������i���X��y�ߺ��i��k������/<�=��L�G���$T��
$�����P���#L)�N�Z�����^��������,��9���%'�{|]�� �C�o1	Gf�h��1�YICI�~��x:]!�w���i�tC)��l�XlxVHYEB     400     1b0El^)^��TED�6&񠰖KX���ho�ƹ������W!";�}�������C
#��?��$w�8>w���˙Bv/�k7��E�r� U�|Ŭ��6��ȝ�&�&g"�J��R�������9�6�t��#HZ�"¨�CZ_'���a��J������Kx���W(�lU:��v�Ei�|����A*fg���,���{��K?�:b9<�|h����B���L߾�H�O-��6����o�*��\�	;�6%�3��b�����$'�4�|��m��4�����&(�غ�Z�Ax � �3��tii��؟In�VM�D<�p�40����.Q'F�,��8t���S�Ɗ�9׊��$�����jѦ	���� Y3q0�� �reՈ*n���x[�������׉X#r�s'VŐ�XlxVHYEB     400     130"	m�뉷�'�����:J<�I�C%Q��zx*T�6��ч�D���}ҷIZ�L�X(�f�{�
� �L4n�������u�xH�)��:�n���� gT�~;�b���Rv�a��t%�F�S|*o�l�Y��dƞ	#�.č�4�w尜���,�y��
���T:�s2Y/�L_aQ?�!.�l4/wx9��"����}���L�R<�a�|�90k�4�W	G�/4�0,W4��YwKB�#Y>R���@pq��l���5��p����C��A~µη��AY$,i����y6�]4�T�r�dyt�	�x�XlxVHYEB     400     190.&�r+ݏ��C�!�}$��Z���\��ј��=������0O��C���MO���iZ5�.x�N{�/�����?�ǒ�k����2��7�k���
��1Ex�"2���9ʃv1��"�TL�?��1AP�=�.���uȳo�q;�9�CY\���K�=�e�������%�;�	x��di�a��=}2/���n����Z���k��&F��{���=.��(wv���+~�LX����C�W���5��gA��D�v���rl�GC�`ت�z�qZ���2TxL��UV��c��^��C�{���ȏ�n���%�(��r�A�D	�ۛT���.��e�� �I��B��ל�.�ҹ�"�
�����rX�P�.}܉�ޟi�$f����5(R�;���66��&XlxVHYEB     400     160��̒_B��(-�d����E�,p��Z=D��H�jpZ���;�NG�t��	s3i��m�d��1�M����	o6R� :RՁ�U���z��R�1�<<j�2����u}}x[�#<[��i�,���	6��>S���<�|[�F�D�I��	p�*�˘|����ȄX�Yu��G���0�qS�鼳��1������z��m�K][�7[��3��'��L-���h�E�D�V��aY��<��).�>c�8>̷2�!P��j���MY1�T��
Z�W��H>�k�c!�A�Y�H>���Sm.�t�%X|�o/7��a�����\ؖ|=�q�h|R{���A�E�`ϒ�;h�%���XlxVHYEB     400     1b0���\Z���6���ψ����r�E�*�g��\����uV�^Ϝ_�v:&�ђ����;����f���J4�$e0��"4$1P+�V|jL�6DVq:��`r���J�~8Q����%1�ǀ?�j��%�߃�=C2@�ŋ�1f�V}H����^�����V��_��eu���=�L�.*�O���˹��ߗ�m'c0�~�eT�0�䍭�V��T\�����{�g8�eDNV�j`�N�|�h��ET�,Ifs&�['8vq5�}�r1����ώ�����G{6��-D+4������)�x��bmf^'
�Y>{����W��Z��2Ԡ����{+t3=7�OmsW�6��Lگp�.g9��U�����&��t���qD�[�H�|\4xP���A����}��n�5��5S=]�Ҥm���7�}XlxVHYEB     400     1609�ףs�z�H��l�2pv<�� /2ogQ��وeO�H(B�+d 9,h����j���$�O5�슮�@K����}�P�"��'	�BFt��u���_ ~��ڒl�p!�>���<�@��$�#=ˏm�P����ڄ�Zo	g������Ђ�zB8ȶsy#�9����S�2�Ϊ7�p�R�X3Y�.�~��%d�	?#e}G����V�/q��A�Xbϸ��&�%�kA�rh(�;�Y�(�8�HϪ ���E5�k���=q�0���LAU��`-:ˍew��dOE�]_g�j�t=�x��������|n�j�b�!��d���TlܧκP�����qo�,gXlxVHYEB     400     120���CF��x�]>��%�6�?���^c�����>G�n<�����pU��� ��_�_��`�x� {��H�}�3��y]E�a�@�}F�/�"#6$�A�I�r�y�`\��(�S)��)�A�q^����ͦA���J�V�F���d��dJ�0��G��#�vIޒ�����{���{-��Qiiҭᣔ�SA��)�i�����\�66j+WQ�)d��B���ũ�¿V��`�����/5D�r��?f^Fxã7�&!����*`D��eS���W���Nc��)�XlxVHYEB     400     190���ɠ�ϲ;<����$���\��7T�ؖ3XDN���3>�[z-�B��5�'�:B2�0Q�Å w����:l��]�/�BJ�9���f�R0�|	�7PBxM@�9\Vg�� P�t������7γ�[�����q�9�^P%���������O}�>��^�;p�����%&�u���bK4��7ӟ�\�&���^���U��%OT�+¯ʼ��n�[2&�UimU0�gwC1����8T��iAq*��HL��k�0S3碜�s �$��T�U�BW�]��d��������R�P�������}r\�s�rȹ��7��h祊�+Ѩ������+��!�g.@��E�΃f����'!ץ�x��"�-���^�e>�ۼ�
-�g��rXlxVHYEB     400     140|SM�����ƕ:-��J��)'�H�ư�E ^�V����~�g���T��t�0�"�k�Q'J&��h��u�b��R;�1�?h@`�7s�8\z,ؤ=w@��S9�<�Q&��E�g�̃>��E���q���~ېx8�j�@D�.��р;���\��2υ�g߾E��4X᯻�3�}9�"���]\_��`�T���S��c�t0g�H�
�A3��{�/)&�或���_�U�R�>�_�Ȇ`����2� �%N'��/�����P�.���X>�B(�4���@ĆÛ?|�G�<8�ǔ�i#ʾX�.�� y�m�XlxVHYEB     400     160�4�=~����}�R+���!���2���������K�OH,��RУ���r;��x�>eÝ�3e�}$3N�����e/a��Z�����*��W1����H�J��־l���{#�c�fp�ϵg��4�3n��
I�?[In�g>��f�U�K!�5��[��f)N�i�5ʖ�DTU��Uxg̋���|�Mm�JzR���p�fv:P)��Be�?�?~)�}��Õ>(�TDY�_�R�k?�A�K�][p���hx�1Q�!'V�R���VlE��Ր;�2��Y�½"_=�h9;0�����.�2d�R�D��jA�-�M<�zη�H�`�ҟ�����t���1����Z=&���XlxVHYEB     21a     100��+�G�0	L�Ü�4�"����x��XA(��T�jݳn��p�B�D(2��z&V��5p�:Y��-|�Y|��$�6���od�_I+\9�(̣���ڍ�*�alD)�yԶ	
.qX�en�h_g@�3֒���� �F�tw����=G�s-:�~��
��UK}MOf9����ށ�I��U�Ա�z芒�9��V�R�ǵ��o��Q�����w�Hs��,�%�a��.���h��eFmF(ZI�]ggu��i�