`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
JszaybEyzrykmhV/bFdd+S5hSLtuDf+6BsKYE8d0YJPMzrQqQwMAjb+THY/f6RL8+05TeJqybhSs
BQ3/zFDh8ye++nGSUHZpkHEs6IpbVdaBE2USj9KgBkDsCmdh7SK/5tkKCRez727ml83HSPCRUmds
sXMDYBpPQnJJeFQG62jWYYwhG7KMmg45Ku2wBN5xbXgnqxlxKMEi99ML0GIjIOIW+ithqlM9ol/R
X5CRJJafJpyE3iAB5KElUCvT/L+Qi/ajoDm6kX2yr+8WQQP81Oa/M7OGURbcGGK98loytPfXkMhA
on1M8mWK+NibqO/AOKnHwkdrk+wW0RD40TyF0T7576vEjlF+2yfFwQVqlMarIbNA8r/zql7B2VUk
nP95Bj8byjnX6suneYjcD7zpY1BB8elwQQELZEhlvuQqEpKXA+WWuwiP0s5Xsr82pu3oSV/sr5NF
20RnPlx5Pz0vC7ZMkRWWGOucs5vV61aR6LUD77yuhdjFeG0VQLYJvqXqSqPYbGqHMF04UgWy/NLg
PwPyHLbSQ7Ivp+W0PbMp1LAYbikQFPmnH1WeItDeLdtHANpYuISw+758wt2nFa0j1incRR+mOKyW
yfLnJCgQap57GUcK069Jka509dzuugX/WpEg4umwTb5+H6oYBuQuPHTcYOLiacaaIRHCNJSYdIlu
HCJ4PG7GDfppBiFHV+GLFh82H9nbPyKfVvAVSrmBMWEjkL54XZlWWYQaCKnJaaLHiigbzRyATddk
Uf+Um9zdthEZNLu1Ds7NabOp7+moGsrqi6r4WI5tVTBq6WjcMZHx+161uuW1QSNE+1bfhMyHaIxM
YWZnLHEBlFiObaD7OwKu7fZ+ZyAexip5G3z7ECIt4mvo15PwK42scZAKEnjbwBkNXNL9yjJXK8dm
+fnTI0+yhBVh9cwe9pjEDERW1BMWMzqCp7CjnUroug5OJpR2PmqhZ6Baa5oRJ7woXeGFkK2dtwPR
RslJECFANAPxp7jTvpvkvHDheWTvyI6SVMvj8W2QIpQvmQLT+P/rN/TrLPEYAJkYNYiVG+hoM/z8
GLSSnCzH1trc7F62ASVjKealHVzBwL8264r3UUbxs6xp/Sia+na+LVCr5gcL1T83U7R+Povf191d
W/y+Bs6Hix8+uWjoyc3MTG91lV/hgvK6vZuqcE+oGV3U1y2QbDXMfFaoZZHCkJlaW65WXFSJtAyx
2/Z96td2/upT//FyRdAL4xvs0Rcll5QlF4US0B6VMUXSENb7eMOfEVjbqkfHbocvekFZOUDFzsXX
G9DxaZMgQtzHlt7ls5HNPpDZx3YAj3xURirM1ycYHabL9CqCEbFzT+LV7NtEG8qTfE0xXgXKkb+R
Vj8k2avRMfSH/6yRWwVH/gRR2Ok79o+gVuBtPdAwvbFaSuL8G9vhrCHLnxS6wZiYieAIvGsq5xgU
5k8wXFMehX7KAusZ9VlByu72D19CXVd5rJsKjbbwZnQmqwQTtgdbjCugD0AAfKJoQoB2NuRD88U7
DEHPUJfo4eW0ExecUn30uFGoS+zBg8eNH0g811+lhrQ+HJPyRhpmUXlG97x0D5Em56gJpisRAaf8
dnb21x+Xophn3tYXoYSAeGvCuZlPc610UhBPVt2J3dXYob8x/MgogNzb1Yrt197dDqmML64fPWBg
LzZegEl/Q8WrrB1gOw9xcuKAJoKJIgsvNQQ+T9XGXxml++obFMYGaOCea6YzywYlLyMeVAdeGFu1
axMyLo09mwCbbWuQjNh6vJ2OSxYzK2Wujp3AASHF+yEXVnX/Eym0f2uMN3Uw2sPttbEEe/1+PQJy
PA0XjQ9JirxdAR1hsCuTVX5tenuWAo2ALyYAdE2zLdSpw0rcHpfJ0/cAzacwvOYc8075lW6NigS+
I2DXIdYsJQoyQjPXY7hMlI8k7K7eYSDREhaamTMOIJzBhnd2llFnN9hiaTt3hz8pSoftjAE4wF8W
NbltX2nvbhMg8H3iPjedhF4CNI4qzVGKyk3DryjBTxgGwIkJZ8LLIPrjchWjqauiitOeu/T5l5fs
2x4gwfeShS/MLJCNuzKJ5uzHDDxQnFuICbhEXogufG2p9rwjweS7sNUbdRmwleJ1MdlodkwdD4nZ
9NhY6uUa5+pSwZlVa/WW9ijkfDTkXyyi+KHGM4SKhHnMcf32Epa3qi3eLfXnanLgO+L7DLWivz+F
+fsm4Df8F6ZfGh9HKBkL6I51og9IBcYB5+a9r5TOeewQpnUaB3mAD4neEC3NfyyDcJ2VBQgUU1ba
8707Xr/SiQ7W+AsUouoYmtrNhUXQyZcLVOD9+EiehcZKarwsgNuDXXiu1DNcHe/0txgxebDbFJ/u
AeRT0CDmMZtk/d9aEzFtwqgk4VjZs/mFAxLBubi4u2g43G0kceXIqhkLVhB1FmRxWEbECW9acY8b
JJIiEWHprLfNDCp2Zsf31ARtluxo0WH+LDpp3G4FXNwdhfMICM6WRlJvZml29Hg0LtDb2RGixDf+
+uSkk+MXCSYeqRjRzMKdHMKSGGxpmOr+4dK3eY/vPeYkxzkJSdOUrMTfdZg/yJm09wtdMfjFH/i+
MZ0sSlhwoCAl+6JluRv+0xoXN/O9OKmjF1tt0h5km/4pXrMhubIgqgZDvI9pce9xBDEEIxakdtmf
jipwBX9AvZ8juOtLqJ8woe/dL0AtWx7xAOGcbisu/04PNok1PYwriU+1ZgTqP6aM3oPiVHVR8HTX
FWZUDlZbWwOE64VZ5CvX2eX69op/0vQOcLHMQ/1mZ1SHbJ0OqbcFJ7QFTGmmC7QxEqXnCnS64JTp
HYlpdwmRkLWMjdWkNmgMpbbop3e47bcytTXXCJiuwO0bReOZBnzZFr0jFZEQ/2IZO0I76TcfyrLt
1kin21pU6aoUNG9fTc2HnVTG+lhdLa7QjBvRe5g5Bvu1jbN9vJdabnGfgr9baBBhb2MzwYOe3hDY
Or6Eb7AFmsS2uyFMX1DNKUGe4Do4RZdCaxxIEflvoQNtmC1t47VkiUerO1Pt70bk0UIGpg8MmGc+
gEU0wmGDUCsGFAy06fEGxtxes7qZqJj52mrs/zqDNVdSLAOZg4qeGT+5sb+yzWo7nNMX3R0ppy2p
aU4uYQkQ2w1KFRiAuooD7tPI0097Wez8cMp7CamRU4Ad1N3CzNhwVbwheK+IHFhLJ7A8UrognbXU
77rPsseNdXJeTxVXQOM9E9ZsqTAIB8x1zWjf33vKuKT0XqqZLjjV5ec5JYtwttjWSKKCr+USZLI9
mYzW7q5Ec3+Y5sg1GEtwQ8b3v/pQ8wx1yZJtwPjc6AgdQAJnmJhhUtrcDFlGTwhWmTbupZIa4X7k
GGLsCXV9DK6EpuPGJccZs2YJ1CwY/cgykEh9pknHH+DmG3IH3BiV5dw5OheIpGLsBFHb6XcWOQkj
lpb3Iet5L8yQsag2Ce/KV9+XTGL30Oed5b6U9ienDbTBtOpGr2cQKTajuoHfW7rJ2LNP1DryF7EL
zcxLMv7jOf3uM/kBqm0LJbXh8TJYa8eBcXfIaZZ+0/piQDRXWVv/LR41b6di/tzRu2KD00gjRYSV
6dpoT1+v89DVt3m8HnNu/CCHy1L63a4DJ4b0JqBNroczGZ6MRhc6ZSmXFEWlNc2NldmYSqiriG7+
4yzbdyqN7e8nQikGK5i6+jH4ZvQhncMlO2BZ6tYLRk8Oof9wwkBLPq46W2qN/Nm9rq3x47lUfTXN
N5IBgy51x8aASR42giIbna4Yt5k2F+swZecmhoasA3f0dqP6RcEv0VLjYJR7Ymv1ae/x5O1ns8Jl
Jy8m+CFT1ttG1tHy9QNk23eECtG8aohCetkxzDP90U/l/1V62u0CrnRUMd25EcWyi/WwwjNOroJ5
O89iGdTWvvDxglVgguJ9IQ04/KuzwRVWvzsTfOQw6bOqzDwucSkrlYStu5wBT+10bI5QTqhX7Tzw
p8evrrhgHn3QcAlnCUw2DLGs9J5zYEC/NZFOJDOm4Zvsx2k30z6q1EZ6eLYrNbl9b93ZkA5vt49n
REkHwgNyq+4yod42tG5xS9Pqyj9Gup2ySk2O7CIRTzskajfvt9ug2xWRXjoqWLiC/fHvH6kIEe/m
vuIv9t/1KhrKgu4gCSrl+4aAnrtlt7WeE7IjZKDpnzkMx6BT74ldpD4blrpGJhnoDg6ebL+WGKTz
gG3hH63gKLW6BxE6JHnuE7eStpCwe27eMR+N9AanWznvQ3CqVhomugmPaGgJe/h7GG1Yzgb1UfhI
ifqHXaWh7+P/RmX2/nkDC8oTt32/PF7FPN1aAk7hmpvkRAOxnISegmJRRebro5DtGp4EmvZKsSl4
QC2UEAM7q+HDOzsShPX4ALr4Ut5h1ifRHrlcqF+uxIoWHYX5qSo3oNNA/OOnGjsz1M8zi79DE0Cf
yJYAixR8HynUkWWyW6tAnLv/MfTeOSTVZ0zc+aYcT7jdRATbd8F0MtHjWp9PEYlyap0HtFPN4Mp6
DxVrZoxawsMJe3jyo30oXW8JJr/fGDcoh528utRpQw6AmYQOHRHZHHUv37Wxg5FnONKgy8R2nXBr
0z6Ctu1eg1T3HJ+Jjxpp5iZUX7yhLWmsPQVAVQQNMxnNQDEqTQwgAgPavZr0AqaiZ6f3pMmMjTnX
VWfXEQWuCV8/UrsCNZ77POiWX796Mxkb0J16YkR4J6/VcTJGyZW2NU68YpoTO+aSfpOj+ARcFtSM
rqdLLA11VKHu4glLfnWctmGm3dv+uDkZle1KlVfTu5eEcOlxrO2W71c/CRjP6pVM5QYUK5e8Hkyr
TPdmKhNUpVVSVAbUvj3CxO4sr1+59Zt76RO3K8LIXCI485si/mBuahFtITixMn5A9ZKNoyeuqb+k
L+0ZM9q7sU+K0AuM5E4Gx6F+V9/53i2kTz5DEJ4DkWJyoaisg9+XA9YYtnUcbcaSImnkEzTwJdsI
1S5eyacixAyUtXReQlHUDgRi7m2UOaEXhKjljIfhUprFxbIdfSqZY3mkSqpoolTFZACQeobyTYlg
bwIEgMURyGm/7qRutuOLHvqbaH5GFjFVMW/19QnZCDp4Udnh8dqPEDHoE1nZJtbwtQ4J9qaJHf/C
kCXaZnHzPQZZRl4TvBFaCnHm3ZVV1MQl7GV0ObazfUE0R0ZFObpGd7rM1YuJW1gQFrenJ2qdLFKO
1v6otfSCAa23I2mZEQFnOtygAzDRuGRvX5QwHSjIGyoiGs51rwelA0lrzHxK/yFDlc2IKyB+AqXi
GHrbu+PpfcvX4rAZhl4Uxe9wKm8NY45rO7xMlKlmo+AuN1mPQ5OutsNQin2GUXajZXed4NtG6QXI
iP3H1eK+NyIXa42hmi/2PVzMHr2DOfr1yklDiBVH1JSuzHmcnmlEa8pIHMIvCprBw0gZgHmULcbq
C7x67/7lb8w95L6ozJI8XPUWNZtKxlPJAkXfTFgBnOS5DipC6Cp/VoWKuwteVQIR2c1h3Xnk05CZ
h3eEAu9C84QsaMrOwn/b/7KNanfDMlXYFZu8sEy9Zu1SR8nH0RmDeyKipN7sznThWHGMzoOTmA19
bs1ytZ3Al7lz/jyZNNAlPQNteCBwoUSMpo6xXsm8yrXdr7XHNusB57USbTs9BZ1fiuVbxUJCcYOr
zSCE/5y3FZAlvncalZcNecD3kUHm6ZwxiSEPTtgdeK2n5pRAAuHMwC9jgsIgHFlVj8NAUWttvk5s
aU8uzeAj/LO01Fd5i3n0WL1yjaE/W5nbUamGIc7eN78zCaEnv7JsCCkH3dggRKy8Mm+Wabhjh4yq
2vtiDJQ85E7riDZHfA1JRNJhxEC6B0x3n5xUeaFyu4++K9NlZdKN9ghPDtcr8uTyI8TFcfEyld7i
V7/wt7OB/Eux2kOepFfPYT3D3gOYF8j7febvyS56PsqFgpBq4iOIz70isecmPAMPXVPu1YDzo7aO
xo3ZCW58zerD7aN/Bb4Lk8w3e8ZuXtNHxr63VzDnr0oQXUnC3tzvPeQDAmeDHqG9THx2S4n80kxN
Wd19XVGFUaQ5kbwTYGh+zHJARK7t26WGfcWwaR+myd5t5PzoV7B2C1OYwJQQjNZr4gjgxe48bqhW
xiljkmv9xwOdFhArkALzpZUB5mgpjPpLVKCFieZaQm4OG1xLDVYYaahmlOJlhTbrkN1/wRrosFKz
saAyPiyqbIWUMtX9bHkK8zlMeYEfLA2wy/uMraIhbne5dMcmAgmV8AChLyWV0ZmFjkrS/xgSOUTG
JCSHRvYllPQmv4Er1vYtxOzT1cflCcHqvAu5EDqgZhoWpDC/i+Y9pkYWm72MasGpTDhiH1jdsn7i
sEDmN2rZFih3PxX6TmvOAr2NQsrRRh6O/eSxuzhMpGQmhGf+pzae7RKFCWltoc8Qu8PRioy5kGCh
Opcxe1dHWhz9RjMfx909+2MVQcDkDzIuPjKgq5j+ACJ8SxJpuis+386mO2q/6go57JzRgVt/KTCN
MPDtkBiGnMQqkJSQ28c3vYf2Vc7+fVcgoveoTUT4ogoWhPxz/2u6X0CioDdrYu1S63xcUjhgXsKl
q7XR2rL5FYEQ/YdGt3DkgviAbkxur+iblrJpRbfe2x5U/v5byrNr/U1V+EzfdwI1cxuvLGVeY4b8
V7T6JWYONxgSnFTXai6ANGqhazas0Drl/kF47PAFLryX9uELkA8uiJV87o60VyofdaRuCiIAGDBS
qCobLs/fi5TFjntby1N/bRzueGGHxICVEawWE4J8qlNcjzWuS7z8j6P1o/pz/kTIuhUC+0FRwqiq
BHFpnrh/BPxb3TzdTd1QPvSAJNnPXKu51ng0DK+NG3FYKkll09CGAel6R0glK/wCHXPvaRPm6QQ4
htoUP6ARBQDVNgiB7rxeKrfDjdBgEkC/vbjrLd7YuJ65zBpDbRUi3Mca58HmpVFHxbcTqsQCmF7d
GaZTyre9YvLQPUiGjYJJZlZc/fjLY8rD8AJtAhotohj8FpfYz6E8Npv00ZWY7TkGPRVsAkspvG5c
eQgHEKcE15EHS9jN80wkEiOxrSzbe+z9NlqHGKLGGPFS3hFZF4IDjUd4BqpOm80qp+1gfTB3rVk+
EyG/LjXNwj+hl0q4uNXKUX2u/voRLvWLhIYDJ5svuBOFfk1mG2z1czsgl0ZqB2GCZve9tSPz6EOV
DkBJ6FAi8zeDdXQA/aPerpviv1ZEp/343ry9ciCGqzgKLVTpVM9dHOEp3xWnNwulwyBkVCpiKatt
qFMfNcL22xiy5n04JkEok6LrMNrQeMRCCuyclEjKQDdljZVK9AZJ05BbfD3mCeZFu7ElRuhZOVjU
ZE1/ogwWfoti1Pf4jFs3aLraQyENuqwe3FNc/qhgPHg3GJ861B4XY8avosABUhyZJtnuNBrEZSu+
CQCK+UY9kI8sn9GSfU0KWhi2fKXqDjDG9tU7P++VQYPTJxUfjD9T9zxbR40nkBCoSxmTV/vsZn6k
Z6esg+F9gb0aDeVxie9w6idbfi5ND4llqGfNZkFY+cxyTBBs8mEpLeXWLeqII1bzhtBO0gpFp0Ra
ciQradI7wnmIbVt1KYKKoUOm0ASB9miWTJw3tSN+UUzYUnHXsRNOaMBrLExc+pEohmz3k2r//fDf
tJDWCT5w5G3B1+oggpf1Uc4bRs+zlCL8wHFX7z9nI9ZhLweaMcjAmOFSUgzeJh8JOFC479IgXNpY
1+qLv1YrgnpSoNloO1SAlZtN0AvqcHeB16JI84NvsO9ElwsBxksfY5jJHmQJduHJhz3BEKTfjlVB
XHwDzEcFgx2/kkNAbgSxBj4BJOxIwT0bDLwL6VWD9KtInbE8beXHgJDe6yG1Vg17r1rXq+nsfAOf
E9cJfhg7KTqRcMypH9RXpg0L31xsdO1s4LsGBiszp98i3UTd9SmyfKg6gl6yMmfHHg3Mlj2DofGT
0nIt/+z2a0ryWKsgYWq8zU2LJNKkCUpE3ehUZfTQXRbxkXR7qB6Iw2NQag2A+7mX60p6sHGIIfSh
mkX3p7+MMV5x0JIDNSb4wcaisEp4nPi5JCdqGx35PVRPnFzQHEUGvABoL6LVR33ELHhoDXzNcOxU
C4JPEoFmpqfqY1/X2zGkoCMdverIdc4jwylyhAMLKeAgp/gKUdJ+6l6jHJ6zdjE1Ae4YYuMvtlxL
QzF3FKU7tYVuruAPRgUzikGbJMtONyyGSsGvpXGspRunNAHqGOzGPrydmwXLYtcV5Ms+yo8Fw4ZH
ONJC/SlsApy3V6/zajHXErOmWOswqdLFfV5AW3oZltDP4gwC9S1hW2H8Y0OquPdd0pBQWkN76VIi
tpdZ+KiH2ur9UyHwBePO/pamHaFm8rRoK+sqNo95GgG/810NdGi/496dOfxAGvdiff/e2lGlqG6V
wy1z9XYE/PhAfbTf1dL21T5Y5lUFVBqb7gB1m0bsK7Wh35+VEcV+obUmtRnv1oCibdlqZwpYyZKP
aFtSgDenSk++5PerQsAjxLIPED0SgEFTpBqsjRgWyRlg3uuirCbCXwih5sG62GLL2mOiWV0iX1wZ
xLc8pAaxuESbh08r0QtZMwVKPVvlooKBNbEccXhBumP9nRuZ4GXU6im+pTLpXNIr1Up2BAc+slzO
maduIQZ3foxuFWe4uI7MvPyLKc0wqdLekPBvB+ZhEBxrOkS0CKrAOVs99w8AxMP9w99dehs0bYEo
Z4aMUJKtACGF3aGh9worvpBpPTarKrdXdFJo1esk7ExNKFwbcz1CEDgRGUTYcI28GnM6P9N3EabP
cl5Y1RJ7DdNk2nh2h6V4EvgcoKgTErdd3hBvLDWmMX9URTnkg7QhUnDnyGaTJfrfYR7FLgze9MjE
Ocu8Kg/jG27WV3m/krEQBEdLj0luhJRok75JiysVJeOKecMBWSpjUJbYaYxXqbtjBarAV7DHjWWD
VKORkn12Hj+ByAIKdxYKs6PBC13QiPbbFQivR8JxCdNb27/ghIWrkFOS+cyyBhoSUfwir4KeLzO1
rtZMycguxRl78OGaZSQgtcE30nRSLymMh/IGh9xCXIxPlqxXlaSjHIS/wn/CPvXArYWFtwX2aNUd
W/SDUkz8SucmmEOqIPpNiO+zzgrTpL/0ChqoIJCLNjNarknCVyDxw0WxCHJpo4PfHb138x0o8zU/
hCih+yg6WgPKbKG49Xj1Rr6lpqQvrebx0UHUYMumU80GK98Yny69Ihgmnh4UXq+3OV3BriOmHYIS
0UzKaqqVc6+qYo2jqWF/cvx78Rq6hRWKt3YA/NeB3MRQrVeNLQqbtK6btijRUB+xreciNimx7cWz
iSJKaA1ZRPyW7YWX4RfcKnZmC5+qBkw7IUqg1ddmKQ47iN2MkZMk2EVjZgFqP6nA5xtOYZOBXaXl
oapta30KnP8t3SXA3wnnvZSMAwE1bPQi9p0APKsiVRlExt/JJgfw9L4g4i2BwlQ8kkNh63vcFGPh
OXQeg5CD8QKNs4siK1CY9XqQlK+C09Mmngifye4pracBV2wxqXeYopYiXjRE/9k34yHhAdYXBnPz
39H0FmDlFu8ugP8nf/N9Dz8xfBBOW8EsQkM3UquJtAV+Ydr1i0OGFNkCQnbPVeDuQRkzJQ/kSbOI
mnSDOGYe84hOX/pjRtstyJdcgc6I7aS8qpbWUHuX98QKvnoqEMYFUnU+Bx+fsN1YuNGdT01WjhEs
tknU+gviaN8T5LEfHGzVC1LYNN/ASJkLiE2KWAMsjUTtIs3FRjLKGmh+OG4qwrOttTJpB68FfY7J
vRUdO7Lq66f2RikDUe8y++LW/uxNOsVQS+sM3gyGASWF03OEWHLxPHQfYXr6wnCSMphorVZURDx+
q3noYtE925nkOsSmpQApeIlk15emcVNRlR16Xbqt+4AiBiJ7XawZqXUk7L9H59nxxYryb9BD2O2J
7o7k85lLHH9sb1On+AFLb4uXZMD+g95znq6j7zkiK2yqpLzmxzBBghCBPFeoiWfXWw1V8XrVTWgc
+N01Qyqt++jW1chlxwHG74OIMxNPQ4O6Bkxut3OOi9wP8Bhv1H6Y74Sju5Hq6QH9Q4wYZdNCvncX
Ar3PNsyZVZhiFWQg51zBvNu1ELifKvH6L2qta4/8WJhTV9IvGSDLwR0E39FM0kxj3e5g6/Q1OPoA
T7ellt4inLB4D37GrU80OfrAU7YWcbKI/z8xyoanW+hAPS0Z6z/MWoXTKcCkXm/PkucfCh0py48Q
qNfSXH1ISZePOGaybIhsCE/UMZ495Ng3/YqrPDELpChg3yxYAYy91EnSTnH22aWo/F9MnZ/bj/B7
q7ObY/7dnCgxyxKEettbbtHYoRfwIg9qYkuhgRsQ1PGzyfQ3ajmgDLjD6Bj6Oos/CoP/X9F9yEbD
sgE/zuGtz7khTVZCdSkoLdVUFF4ciRoG+uR1GXYVrEyNmXHb95n2o+Ijl9UA4cLpb/ueNUU15Lre
CnN99PHD2GMb/aXDXXGdS3m8I/UaPVTCM2XtPhPjT4rYYgUpc4KwlbNaHp1AzuqdRGVOATDkGqyD
7Rrr6onJydYQ/K5T0jCExUfd04wSHEvLM/BG9/9LlHvzanTPkHCaQzh9A4eU6oypIUu2EaDFMI2J
JqsYDLIRfQeKfwT4668bBBR0Ov03Nof3rc2TAVw0MMpTBtqD7u+Ta1cpE6dHPqOWmfHbhDRrzdcZ
dT/2b/jAKZdIo5wh7f2Z4r6GbAw3wXSSnyHC8EivV+iZw1uHwCp7ZJDqzCZbLHnN1LfH96B4udae
SKXdS0hJCdjOig28vUSX8FPxGGLDLhk/yMrPxgOxhqO1luIpOurLp0FreoyzhJFg36Tkjon6NvRW
EwMZoDqh5PKXNRBO7nHjoDv8n6HHSo3xlQJ+aW71gGULHfz083UoEtyiM4TZwCFsotwGweVwYp4j
0LZwhQUfRnEdnw08JDKKAS7NHySt/W2uNs2OwUZG0I9099ZS3TM1tqlTkysTmSP3jJ7JBui7UKgz
oFKrsW3MBd/ZzoRKbJQACUKWG4Sk0HX7RhaJFpdQw86rlwv9tvgHYlkdmp+1ra9u7JKCkfuT90sY
K/nsR1AurjxZgilUec79tGIX0fqHenu/tc4Upqz1wSHh5v/5VzmQ4J5lCUAC5BVM4CJ0XxcgtLEx
IDl/Hzdf/fNiacxmlZmLUSutolL+e99OSMKAMNxtNF9Hw10zW7u/84jb5OHiXNGAhqUQPd8ZdQbA
Sj8VUljpjyfA/aZqX6GgbrC2TCK6MTVB3hWdi3SdAH8ZHgxzaWFT1tr+ol7sPZMHbioHw/rf90G3
+ZE/nwRsn69Ly833NkemA0JyE480vF1xhsF1oxzRBQfXOVhofcZqVO7RcfCpBi+e35X7LNhkHQYf
T3o/7S8l2dSjoyhu4XEhOHcCnl7mQVJkjDi8ueNp+uuQfT5PM+GObjZomDloT7IlMmcKEm2BmQ7U
TpeHwPXmCiEkxgq3ZkuF4Cmbp/AyhhpbGft0rcdMNDadHfvaUDJvRMDoO2efuealYJgK4XMPTWw/
057VWA+Ht4qOIwxSnZMg82nEIO6p4dtuk/Hqr04gmhtYvqhB8ZfOm7d/L0M+QmxGePQDK7stW058
llCXk7HpNHcKnajmUEpaWW2S+NPV4HmKJTq/njdaOva4+8SptZ5k9hWfK4BsbzyX2wXblgZygP3T
d9f3mnDO8X+HRMn2RcosNdnC7C7EgDJEbPRPDhCdXjTuRQ32UYi5BvSJu1haiW69Of2MnMmXVhGR
2GHKB+kSQjfHQpGLpqcUjnlZaDOtUUrf9SmZeOjq/Ajb5j/sTF8sPRyZnmPnrsqlxrzQWm9FYEvF
fs5uaR1vteIkRDZk+ofvmcc90Q0LLggR0MqsEuOoEY2JDx7oepSV9JgIXJ/FhXPVBklnshP0J4S1
PD3vDVkzZFuFWaags0uA8GFt8hc7jYYkWGh1tLF5H0iVIQl7+MiPK/iwbxuwB0EfWyDpfLNpbCI3
9bx0vAn3wSKvEREPAB3pKcey7p7kWmu0eFFQG+vG1iAxkorDfsPjjSfjrRW+IgSs3tgb0H94uLjS
nUxNTXbusS2d+GxfhAfnCRNrcQL0MQ8BW4uO7+Eo3tQTVb9M9hztp1iq0LqJmP6tYCemrYeSAa7V
7rB0iME2RhOeL/1nqJppj2oRK/IM99p33DMB5c8vLaI8nEeggdIe1fiaM10J9p0fsR2Mo3v50pLZ
uUJiLoRwsv9FbM/aKvcJSOb+IUjq0QG8firaVv733yv2EcwDSZroMP+Tp9yVRg1lxIryHE3a515T
sS84T9Rem6UFzd56KElCGCw1rVB2qualKAOOORpDAQc1XE/riGRcIj8g/aRx7j8wYvT/eqPy8Enk
TiRHDI52Or4d6IFfPtsCviJRM1h9tRXMIbwk2rzgMNccYOwCPWIecXuY5P/bsAvdTdWwPZaJpY7s
pAiF3+rTaS0jhUEMD8MpPvzH9t7qb/wd2wO9v3+KnrCPMaSNRMRTzCCPgMzotMXxcqo55/lry5c7
aueu8ahHW7vsDCvjjYbmRc/SGR7dFLrbQUsGz2McnnN3WtKfAuRADqKhW4D72JLlDZiR7rHkyNwv
necZTToki2xiw7nvIDm39chwbFBC7ZY2r9SF3el15Syf0KCSv5s1e/cTcJY6v5xuQNSMEB/Cw6Pb
nadeoUedJIGRMXc2fjohYiKnjPjOrE2sdCBKLURrQgg+cMuiBq/ykRMwwPZXon8htTZCc6MN4pRU
vFp+gSsbGB2dTZti8GoWaWHdvXaq6Ikc44f+IsFRgLjAe6ifdydiAmGz/2sNrsHmJDbFTwWezjAb
g8jdVbc/0jRsx/9dLCfk+RMncEE6XA4E33vJVBao7tdj5Ly9wDwypqBUMSQz8trBl9JNAoVqFIdB
5BdAPSMtWEW4KoVR8SEs29B6IKX33BP8D9j2DrrCJKHKTU3xNaaYW8K/XcXtwNTgAFlkH/yfelgK
XopCAlu+xY25sisumMximDYSZaUiEnLQHt2plXjkdL7bQHx+w19cwB/jNV4IZHTZY5eU8Zpd61tf
N8zUuuuX7+FoA79+LsiiT24ZXIB4T9PpYcYXAEHF2i7nRWoS4nyg+qYiLAPGfN18i9kFr74E4xZk
L8vZfTpHOPvTamAIyffWBKN3CDeAj7AoD/0R6dpReP895Auc9ZbeYg48/H32zZxmzvdTunKsx93+
oQ0GnRhqRwC5sHZpcLivnoVw980E3GXuyvKRNx5V5sj+7m5IIp3L9LW7EpXAxf6ps2GObJL7v1XT
qxxRP3VrrKp/y9goD98+sRcTN5tKJ4vI5GqavJ0FNWUtVsDZ42QHVBOwIQYGUrB/P8wAtUr0Ngc2
pJihbTjAXVxTBgbBYRLPCBhoHe3A4CS8dLRyXiVJAUJVa/b/QYn/jEeEJ8Js3Y9sslxcXnw+iRAV
bBY6EpQBP41RNURki2bpgRAZ7qkG0Ps7uyNlR+mYvjLzE+z9eDdlUWYDDENx2IbD2+bhZTZ3/+BE
rNslHYPK73DrZKGlqaStGIexfRSnA/MzPZ2NsZT7J2Jfi5pYvCiSs0pU3DQWSfJp0owJV4H+CjYL
ZAfRoDiyo4MWE75IHje8lmvSTUCuI1yy5Gwo9iz5SyRp3Zwm9yPQqh/3Ka7G350FASS1tL645k6/
/jTmmwR3CkunW/IS/i5jASpOtJ6Eqza0qK2qwogASCMyyDmAtvSuxrzQjo4h394U94XOxl3O8JpR
hnnMwr46c4g9l+I5/bw2w8MT0+TpC/dBhlHdja8cAsvs92I0yGBMXjaQ9/UDJFtwM2NmgUE5ioRl
PANmEzuEvovOpQCzt6RXC6g28rFPisNOCkRla2V6I8vWXLIUF9EyuXMnZ+753YDcDnbay0+nbxLo
MYiktzw265NYjcFmm5y5TZksJGp7PSH/kCGS/UYjrYhlIoYjjs8XMa+dZeBEB1GriwesW9WrQ3Gw
e/4gbEGpif4rPk635lpGCn6VFAXT5Z/A9tGtlrn6Z8g2IgAZ/Azz7xQAN4jQf6NtwDQKPTzGHUGJ
U2XY+bdTe5xno/sp/wu1B8QVShpCI1tqtyQI5hu2+QWFcWTtwyVZoKWFn/LPwaLqGLxZS08YmAhh
L0zoQMNrAijm2KzLF4qx6ebJwZ5iLcV7uLBcSPenq5Qclx+9ZxBzNjPsSofpFAc7W6mQhIWm5pj6
FerFmR+lOHXcHNyMMhfShTwVgOA+4s9IK8EQXzWtCtC8nyLFrVpAi914KiBPM+dyPNZgdYDlpBi/
Icq53IlUke9Zz9On29v0fvFvfRSkRQbZnAW4lp515wsDoS3z289enjwwgR+bgvDq0H68eNuxodu5
HVYggRpJCH2RvcmpjeMdtoB+Tmtz/CLmYGh8+hvMgVLdJ5lmPXDoKNiT6sM/nfWSiV0zP/yukrEM
ti7gOTLfkwm+/QHy07j5H7r9OUoRhnaBZ4yV+doY06DCydh+QqXMDn0ZaCfsYuV2k5GzWgj8Gk/G
n/AM3gUWwtjRdSoC140u3mAYVVhNaLrsuynCzu2PFgOSohlVG0yKnL6YdncBKIhgCAw0DoFh+mhH
SUfeynZJQArE2bTF0SvN2NNNWCMlZeOeAE5PKGOKxwUln0jvqe+nH4vol9f8AnHhfWFPkfgv8WGZ
44PnzgiuhZi1+WeQV68xAG+uj1Gu1iU6fdb9eAw8L5ONFUggoAYvfHu6CdEvlDuIk09+/f1HXA4J
Al00GzQv27AbOCDcA5t4Vjattfxrq9CspLnCpaZcACnJj6pvgK+8gad/4JOAYqRtkPXDIIsStfNc
2HEg++uICfhFKJuFLRTGfo4iZkSluzyAUTHOurYU7U4mbTXY3w8U/mlGzq/a1d7q+z/exKu0qI9V
E8e+/rRwyvmi10Iu5RiNTPtXKaVNtupYpTdtMfwIJdbMjZxkxc0p7o09G67erTdpJn0mffRMQuJN
1T1tqErg23uErbP+onLInC5efLb7PlKD0Gzn3e5kLifWE3jwXRisGtBBiFA+wNkkZ5guf3aAsmvg
+JtdADTq6S/uCRIX4AwBKMDGrazXyEZ/W+nXJvmIZEnBY2/25aNNYRw31SFf0rPEjEDCK+7zaTT/
Ojf3ENRS82AOE4rG6rguchI0jIMsA3CuM83TzCS6qoeDqZ6LpIKPja8IXtEqOeO73W7ztU6u0wx+
odqBrrle1VmPj70r+hD5ZFrDznCzhFuYk6sckyOsOU13iOphNG9n4eFblr3zfP2tpacfIndNSZNK
7fKH7IzQ+7U8l2z8fYiiHhDsNa1yWZTntwDkE5OoC+Hv1+bRxSkTMrGYFMs9v9XYuioAP1SIGddO
7H0Ty9cLcU0WD4nEfeqheDI6yc5zbUZQY2TBX/pon9jJX0blFNaGq4fnUn4vDEbNHzlKUWrk571L
VTB9TTC0P+3d6vsuX6UrmZYPWj+RzFce7YVta20cLJSqvHspNlp356MTGkeWXnqBJv04LtYSNIUU
2uw8eMLdNrIxFatBqOdpKvFPidjZYocR+NL48ePxxWYFW8nRyDGszZizqYUOVo/bwkVc9XDOaBYV
U7MXHmDJ9O/kaMD5GeWNkTUPCaUxH9qb/MND6Pz0ntPN+OvMvLoUaKrEDY6ZrO7mcz7/iNFNqWMY
Er2GNYVRka5dvO2TvQTy5keVEddN/OL/vJtwFuxXS8IQ+QAlt+0jKxpCZesbG9REb3mOJqDrFCEf
A7y1HlKD7zsMWUNrLUyIojK5E4ERtdW9NfAZ/KWW1RHb2Id8+4Z6K37q3jHmXMUi/2xOjRnMFQzP
+Gl5QYnQqtFHIUJVYASb7nHF/2XVl7VjkGa/PSA+VQ6GxxiHU+ItEuTljistUFYQPW5JFFAIpj1J
92mqRfHpD37ljGvsqLsHF7OB0Tululaibfrx0AkXh9HRab5jpCk8XlDd/lrFNguj5vwiCAes6RnV
q6Qh7VItQInfKuPUSZFv+6nh76ajtAP2yU26dQeOuuQ3ckYl98JPUzT/D0DF67sZCXCuFBb8nZMv
CAu8nvga97YjoLqh50VNdhowBxePKaBOk4FURVcx17gG2irHD8KzNn4A2OJaULxOlbuiCpUmm4Z4
7S05UX6VDcyNDCc5B7AK66EzxqmB3MggNP6YIOuh7yg9ExCt2oi0xnstaYcPr96wEVO58bcjagwh
84mPTha89SSRXIgtWx6qxvDiM5dVgMz5180S24LOQ3ZXF2+L0tgqkm5XlHw230B3qAHf5Oc+KqsR
A8S80i19n2Dxoj6fDTvIbaRInDh9wCQ4cnKdRdE1bYXnTEwinfkDU2DEj6tppPiuxouekfsZfsW1
N1nukhhbIqOV+WJGzct1mHEfH6S6xPbplxmttaW4snZ83Ce/mrRkpJtv0HcvLqqIxxfbVs1UxeoS
NLo1Rh2uf8Q9RD518RTNEoITIR3AbTcpJSn3KyiEQhgyDuLGr8AIc/RBnlYqP92uO741J2SuY9ZO
MpoQTxTQk9UKgIEX8dkOroRuYXav2YHFmN5XUKLb9i3h71vYFwzom48zFfuXn04XpGojZH1Fi3LG
yH5LNvJI9wEUTA353hmVyuw6D4Y4JRr+GOYE+lvPPVnzN1xT9f7EjJZmeI6RxiDxSpGGW5d3/PX+
BKWvU/tasB6GxtwBsWg80rNwcf9penxie3kBQn+nIYY+X+IuNdXPNKVPEHxRUAjWxO8I64HjvbEI
k3WPyS8mRtKEDrdXC3od+0JXsX46SaCjm1uaSHvYj+aDMn1rQpkbZXiI4xl6hKqWw6wP7rYt1koM
dMQRkxAFNpLIUHiOAo7n2mR5D0BIpZX10EZXeyb6DUAZsVyt5Ag8c8UkAGnnGt8a7QCZ+9h8otSQ
heEjIHXaGu+Lhy7yZxFPEBmhSzR833XO+INs2DrwxQNWFAibfr1js6ATcFyXFgcI5pF0UYu/ilA+
/xg1HY/DnTi1DWqSYR96DZDr+2H6snNdfAKgNKDXH+SW8YsQ+MujTHA/jLorpFXl8vjgb7o52ppi
sIJUx5bgqgyJ+o27iUJtO/eAKUOJ9WJBSelvrgthU2jzx65uE1ZBfKJ7VKaYzOJzleCZ07vInuMb
mogzBHUsUCy9Ok9BZ5AUZYXdmOeGNMsDHzrUrw5yt8gAbK+BQlfFd+3wS5/BPFhcWJDUiz/ZH6xW
fm4gyJjKRebniCNF+W1eN5KM/MvHUQy8G8g2ZfG6RtxmqaaFkVNDk+wqpbGPo9zDt3N+sxmGASoV
FB6ROMwcMmxlkVdVKCjK/fXyHQo+myyhNIQu7IKHxbqQ4QRbODJVhnORgVJuzQeFeElvj2M6eBn2
uNXQMhQCSnwt9kigfDSe4mdN++f8u1AVPhPQuhW+jh1pH6h646JqM9MyZap8cUpqXUUjbhaD87eN
izCS9BQYhBe6TbZgwW846zyHWmMOc48Lq98CCBSThPZcNQAD9rED11nJ6eWwNlRhrcSfcYy/EEE2
mMARynM8rekgr+iBrMP3v5hn2hsxJm4PNOrjou+4auS+w0e0xFAqkjv3Qkxss3oy2UP1DX9CR5VZ
f5kkF/yqlnAaDM1GDw4aAAnhYSv98YSRXocLYvjx/5o1YT2XulXh8/dLE8PtwcmlGDiXlPsTXwKG
Mf7UKVJMMPBEEBvrdEq84s+lmF6TKYIScHbuBMRfFMDixa7GegIrUevi+jPO57AqNAkBkrIkkK/v
XF9Qh7WRWXrAA9KE8RVSNf/ZzODdVQscpivcnsHT9l2hRElfK9+i/bzmqjiIDra+9lfVgkOZyZY6
PwuH7wnb4APlPBYx48Kc64dwHpMsTVaYHicss9QUZ9LBAX05e50HsS9qZ+XYIwbat3+L40kUvhLo
1Px5P1pp7UpJvLudKIng89CJIuRXjt7Bj0UWVvIdSPSzj6YhtutRis0+NH7cs2INQ8Xw7m6VmepB
Sq/zVwvZqlaDeoNRdk3izz4C6vaKnuYWrkrOr5GCXDHMvjdtOy2OMHaNXxhGodAUEdcHWlQ0IqiN
dv0fEUkZSLfUxilh/1B2l37e/h/V8TVtDL0ZeS2cG08JEEf4ZOIjPfPcFbPqo1ZvuGO4fLZgpT0n
uzhliQss5E7+cbonhFG87wF0uWGqxdryaizHivpQnk4vzbevnN8ddfQP3ZDqEhHDFgRxSrKCRHNf
XLu8NWMttOFXcbtFvhalN/BOd8uq4KmX4U68cdGl48RL3oBFNs3ukxWpWpnJQ70M8LXQwYA+yAUk
lGsejGofmLLFqyHHllLBaOtgwNcI5tjmxKFuVwOgXhgrtTHd+WhPWxopvAxWRM2vfRaQ/Iz7A9KN
9ERoiyb95cKFOncyPKhcX7e7LKpOafrr9o5LWOIsexj8CBO9OumTm4KKXtYAFl3tKABxeuLE/Q1q
Wyr4WbG3AljefNdVQx2Rju1kLCB3GwMk2Abv4TeKfxOzW3Ju++BwAyJNCZsV86ocs0i/rkLoHAnP
Iag0ZBLHbBNkVroJZ2uE+gYD3RFHn6pokgFRMggh1IrTgmPFPzFRn7vEj5aVBnYYb2jj7FfFQh82
AyeNiWJ+r6EstBRzaANT0XMxmnWB76T5lGhefbxqSYES6GeQR9oyc6t9Ng9y97NNqH38mAlzFXYj
dZXLhjc2ttQcbtv3R2yHB6vsn3XKmaR2Fz2rVtx6Ld7Tf5F8IAaO9s/rnizdmTlsMEtjKP+ji089
lcKSbKkwRYBoc3wnkQJMdMs8RUaP5tkljlDP8aDUcjYVBbnlRvw+tuhr6vFQPN7iMLGDgo6w/ZEH
z7OAPbecg9cOZKnzB2n9tUgRfT/Fd492wldJK7dYRVNtz1L1iMQYvrSkv7XbegufkmDoswgtnRAS
EAD3VeH9E4t3VkyeeoI346SdaFWz0IqPbDgVnJz31S/mJgv+8/xsKb8nrGbhg5N3S65ldRavFQUw
WXmzLEdbLVojRJa3SQJ1dABm2kCwR8ADKdhNSfRkMvrEQugGAKNDY1dxy809fUpodR4BH+DCv1Uw
OVgAu7/o4kYHsS774HKiYeJFiTsL20ELnma2bpNDljAoNZ+ibrpClK/t81RYMcq08WbnCb7GEtWA
GwiMiOUFd+5TeXEQX3UlCuXM8NPmCDA8UlT8D6aS6zb2NJRWxgLvsvF5tyYy+SwXfxbqL+X7ImrD
fl5x63ohHXWMsFIPD46t+a+JpGh3gXkJ17pmCBfDwk19yJuHMeyvkLZnfrAFCgKO9310WIeUmCwG
11JkCL9kynxXULKNI9pM0mWdboHVOsntqhF8BiH/WcUrZF3UUtqGfYI/cH4OR6Jqd/KK3kVJNTAF
duma0Wxy65THKYI9vn++rLfup/FkW5M6yrTP++jOCldEv3APR1AYsrwZzjdJf5aRPuiBUc/rqcnK
4FuOiQdfi0zRLw1XOcGXnVcmygJrrlgbhindBxVZ3LZO9y7XJkhtftdeluiBufCrDvag6VN//f80
wW2Z4A5WoP4FhlHgdHY82rYFgaKikajR2oryiD+W4Bw2EzUXTE7WFuBr6DKirmiuqEfpBwg6B7u1
9GvWdfde0/ebC0t29ckkWeX3JqHfMb+N/q1crhLLaWGJigRR6hTMrwU4AMyPimuoouXkimYTWLmL
Ou9Z/op4YzCprNHyPF/ikJ+iif3cmC/FtK9SgX6if6hoI6YKMLESBqgTTQw6+xNh6FW+B7xblRyS
ir20sMWUrgnkn/CmclUfFrIOHNXOzQzu6dCTmHZNLHF5dbnWhpNG9PUs3KLKscWFqYKc5MK3YsYh
mp+oUVEuoOIGikvaS2744QUzS/qRId95xaxk6NLs9tX9j30MRsutSL+nK3662pRiPsbz/gDcOr3e
Ht+I4iYTfb5RrlRFf30NEk6vsXiW3aK4ytTS7wrqWQyMuFvC5b6Vqpq2X9UtIZbF5x7TWWmFqu8d
ILEM+pbjDQSCxWOArkYBJJGT1mAhpYOgpjQcCcxVpDhkTw8Sp0HxeHRcpCYQisv9k2TMXYEKVm4w
Nkz87WjNtINtoukUMGfcxlMcTds03pDT+VRWhOgX8hUY9qmwhywmm+6ojWjQSFeRYG4fdX5k+6SZ
VC04rs1MXMvw0EEyxdIzB/kbWtr+5MZ3f1lp0Zd4Q6tAIpej5vLrVmw75LhoDvAOEVxaW5gcOYGu
lGBWZvpg5++4GRMgckS2UBOktx6XmlWUgnv9y477CudfaBi61Rsd2Pg2mPXR9okBlRlJrE2rTM3c
9g6seLJG07h3kQaqN9N56ssvEXMCqc5NKU3rKXbXTZCxWfiJTdtpNkpG2cLTvqGcihmnRLpo20en
pkcnfODL9mWJ/4x8JtVBj1cS8AVSHPOWGTTen0Le8fKZkMkfO2ZyXkHsfezpM5FExd73RBdtI5+m
adswIqEbZSU/FWdcas/NbgFzJbB/Aj2yRlnnuWQGVdSU8sELJXxOj+QgoKS3F9gtgtkQdxLxCtSm
+GUl7drvzJU4+CHqmewSbABl6tpcKtVABXJ0YCNFSW76xlM21YXhmSI7DCkkneJLpMG1KqB+ht3i
LTxPLNWSOssS6Un+1Z0jygPnGlsW1lFI34rXUP1ddkdCRcHWBh0Ozjtkpz69Dy4uO0vErv1xhVM2
H74V6EHjrer2AoQDsq06mRrM9Fcy09LqWeLfh5TpDPSyKUWoYADo1o1fNv1Ab6I0V2BioQoDT78z
qWDfoRUNDKsv4TipzEqBkDb8AxHqEEtAf3m+PIvkNZg9KhjV8TQ2w/uBt8ckUMuWLw9VXmrm3eSz
x7OGa7XkUPwm3cFdFsL5mjDIuu5VrcJY3jrk6HfkEAy11ko7jmdKgeTdmxDbh00lDG99rN5I8gPm
uO6w4HBPvp9ZVot7fMBNboFGPiEs/vEvg7kCuQPTyf4CkBiyMXtNpPYjCgJTsMp/QfeE4icTV+Yd
CQmmL2vjkmE0r7M5aaZt3qAHYdZTuhZPIVgsfZu2wp/0KFZ5Orb+aywreeOx/wfdx7AgH84J22Vl
5HeQYt6qyQbGfz4FyootRs7YYBYTDAFaYOAhWHYYDv9wRG4LMbQrGpfmsf+yRMA/YMviNlmOBTTo
f6E6IpOL1xufJTh1vcn2BSUQr7+1UXQZ4/oiGUHIOjHS7G3Nrwb/GVdM9EaPIF8w1Wb10vcTBSxi
a6nqO7Tj4I1dvD3BEa/JejhtJLBEl9B1sKdTJk7+FQHqqc3LVeSSXaarts6G+Bm1gpE+R1YOR+Xe
S3ayVCkylDCq5SM6N9oL1Qv2Mu/LSGO7ANi/GY9Y9zXRCo9xT8t8J7jeRqQrijDpGeHtAkLoDlta
IWvmxMF3+oKSCD3uRQjtfvNB2RAUnh7YOuUtXtTU74Nf+dBOcw82SZ8okLfoa+EwgLqG4mXlYnUT
z1M72ybEswI3cO1MWKc6MEneaurrk+9UTWIJnwTNhAldMsJ4Z7OFnaIg+OfTGwdvHnLDm3XLVXu1
3q6kfPqEQhIk27ipP4lwPkEana3yAJbLwZTXZo/kT27iJklX1oALhoKBQILtzHAbnAXAh1atNoac
7tRPGHS9BbLR+Cpc1dGKNdgf98Fbpr2I1EJPkjFUC5yhMTYevEivgVccCGMFMD4FjfwkazoqShbL
RJFMLSWrMf93ibg/yhVGeQLnUh4NC0YmFS0MVQsfsSlaYQDc6XOnjzoUZuxy9pMGB974wEE7OISC
XqSpRVhVVe4vRIcJB0wcV+jaMif99L791FUn0uTdMRR7mVVSSge4RaF5a2fb5eQGVeM1lhB5+rOR
SR1xHUTB0HvUkBEp9gx6Qd3vS3Q/mgTOXbdPoElQMQs5CBckk2APqtoUhyh1tIq72cPvj7LDYdBB
Yx+3t9uE6tIWvArvJTryGfxbsdRaZju2Ibo+noLjRKlUJg3QHBAl5yuj+yElfKzjFnUBIwwstBjT
wU2Zoa+DdgdQOmMV8fc8RujCiE+/K9kKVSHpbxT8FRlJd2QWMfZvu8NATikaNAW7oI+r1xXGgJwX
wLizgjiqtBWaSOVyfP+srjsjl7bGOvLqJNZ2Q3x214IVhaN1FuSpGP1pnvTWNfWL2oXHeackmjp+
9kkmX4H+0nPRc4292DBfhVrkiOrj3lAAqNX7uD+B5xNE1i8Ray8AzPS8ibSD3xpp2OuR1PZL/W/S
wVTD612ACNtugdz73CI8hjWWR5ppSlKvsjC6XimaDRaKWeM9gDDfpfa+nJGXT8sO2mqnMWjUoeuQ
VwkGlojsZYns8KN2ahgAjA/rRc8Pdsg2wTbHlHYlF2UMrZw8D4U1dNAAz36dJ+sDDxwL3TJLXQTU
LBJlQLsnurMnrCwdeR9tBG68sE4S9X4hCjVFWzrs3FeOvPi0U9FSEDNGmtliqLTjkXQF6trQjFgc
r27KxEoGJggEwSWOCSyKonfKqgPaECZRzrsCYlUDsZAT1Id4gwEX9SGJ6OWU6oT8mq/bAD5M43iz
bhfP1UN7tcSM7qaLlaSkG1QVveebbfjPL+sMOsdbEePIdSphs0eySLGw8Z7yk+ifmmI8gr0icrky
iKMOBzb6qzuaX6jZGaaathQjXBzph2kOVPKsd9oTgw/s5Yoaz5svB4uLc1NmC1goxtiT+wF5PgIe
8cOazZuVeSfr1r8f2KiqdSjVTwlb4sNZLLQSYHMdBzISDGgvOtAO+kgnVBVhlWhjGp6AadCdE3iN
us8Gk5Ue2ETldJlf11wpcM1OSjFRTTBbkfoKKELhpfzkdnn7qcb6DV2vxrZ8vyN66nrW/D2FfLrQ
VN284Rp+s8QzrlIxsnI/Cp7VIWE0b0zW6AvT6WFuORefX+t1lAEYHXOuxAaAiY8B5ULBToDmplMA
Lh0n8MsFN/FKwDgT60DgPpIN+w3CaHBN3SUGWDRxMBsimvFQSOQtqS1469NqMaU/pvJBNeqy4y0C
aPvOG2GLwfQZ2pVg+/UCYSVMEeYORh/ckyKaJ5uHJF9yF41NafAsfBgEJ74nuVb+CW9wZCOxnK7I
3DM9TsuoLYjsmQ1oZwmj04+cpaBZWy9JITUyL+OZpA7ucw5kqr0X61CA/u//nd7zy7wg8I0uMf+m
EPW61druLF1GDTYA0Z9saTrhRmE3QIFd4MkrSt7sU9z/XZcTiXDSHWn+wapc1EHPQiM6grLeLTV8
+9BIQgZ6+2enA0Vpd2wvv0HwOxj2XEbneWsRBoTRV1N2GuITwdTR4Zi5WndECDY9Bnh0fidTQAw7
PHBzoJ3rBW0JFNtho9VEqRmUbEtX89f1f4wQEsMjR/IcWOsfzIdcMnw5kDRwb5uTpCxTPNCXy35e
gj0WE9x3UefFtggLIJgqe7ymzAHFl15Ec6MCmHBldv2OTP6dtRlOLQllhh2z03nN1jDyaHEhZ9Mo
sWbjQgWh7ss2p2KgYxOMstPKbklxhZySpfGtRbzZSnVxkt6EcNNx1V7pwpx8bFGntJVL1d3cVGw8
keoYzTvCl060SDHMYp2fiBfmegysuLRsmVntHljuqIq6i1Vj4v6MGz3WupNOmEDGFOTI2dR09ef5
8mH8SZ+Mr1lF/NuZGeHHUKH+6jnx8Hu/rK1MEcUWADEFzkmWWLAB7U/0LiqkIjutUdr3emrom4EI
Ec94LjvF08RgTSDh9pWAGlQNjHJ6mCYCKB/Ashy8RVUYwIFxsI5WrMstbzujlJ6pwmY6kCQ7W7+X
56Hyf+ZsEVxKtBCVTM8t82oqVlHeCgyjtECM96fLWrxeQytgpjkybv1FGXmZiWyl2qydw8xD0ptd
zH2hJZNVMzvT84H7X3YnAldU91cXLpShAKTtAFt5RvrTeZH8p/wDHI2XQOJmAoCQt8avyet0Sru2
OkBiQyHK61GKPQkaJa4y28K9AUS8hYeOfYJ9Z6FXSAqa+J8cpfgKnkYDbzUZ8IPQA0yxHADPOe1+
dwwz8B+cBfaLcqFPQOQ6K6fTVq6J0Wv9hE6bTr8spnlnP29s0RfOZepLOvsFMKb7F0M9Oxh2Zfoa
oEstv8Qlry6Z9238wXMMS+deJM9TgkV/4nyxo7g4IK3FnwnMgtVsA0LPjG4TPTBeGXUXBozy8LTU
eBfxu0g0FMXmMgCnsyA6uX64GjW8WGisX8h3G36bThs/NOwx3QCVylQfUMdak/i3GeNbrfBTRHSA
iwOfVTzsLdrsHDXsDrJie2DNOPfuNCWPs8l4m6mGA+XDu0PnDmFSYiYnKcXR40EAVRSoxJxVlcoQ
aewywMlK232KoWK1kPoePOH7fgdLfjr4Y6mj9vwkB56/em2rvaz7GMidL6i1med6RDDeMNKp6E44
Jaj5xZtxEV01mkF0s7B3RE0iNLD1ajxKcWG5BvqcD+cii5Hwzg1m+EILSoLRRRLYfj8IEnP3Yl6w
/P0y//FdYeUNjqrNX3LTzmP74JxFHPaJPeHy/mdF6HAWTz1l9KyDbpTPtwn7B2e9WjIsMEYgY6+0
8gr5RcR+jqjfY0P0v6V/jFU94g3d9L3vwNWug5fXUGRuj/WMIjnFVaH2zy788q2mS1JkupG6afkq
V1mn/Ygo3yucCIL2Wji41tobZ00ZM7U3SnzuUXHYpykUnEvKIonJuCeWiKcpValU4IJi01f5b0hp
RsQJB30knXd4QxQiQ9lQJZ5brFQhIIBiO1yjmEjJx4wmLQ0jc12/Qb9sdGRIXQ0n6figg1pjd2WE
RDfXSdWr7k84uMnxoV7n8TUb18TNmdBqnjj+0OS0QGNk55gpJ9p/pirQWB39ogFO8UB04HRdK9w7
+Mgn1Cye7p4JykioDinJePB6VyizaDARsAe4wGVYcrOnZqSBMbIxKjegXwjhpoXz2uqKK01zlVip
ClIznNh2W+hmsMkvLkmrdnIs5aZmUuzD4dvTkyzRPtZKldODOIhHdNhDBRHNeiW2ZpRgLFM9tWbe
zbGKL4ibzpJg6KgWmNyP+3pQiaH8LpSOYXRENJ6YE3o2NsLKLAzCpjIYPTO8/nzIrHfbvdSBfMbl
/jgud1abCmhQDqVl3czQ1RSNL8Nw16PBGDhyg0S8ihiG82+/6P7/rB7ANT6sBL5JNpj1fYfK/2Z1
oH3qcyhZvOZSmwGiiYP8PSRqWFNlyiN3FBjS8giAxCJHsLZrTvcss4eLors3FGzBVp7xMz6lNUEU
Bc69zEf/ZZnrtJwzJOS+j5bNUFmx4o31N1EsAfqTIIDnz20SFRhhbEFBW9WXCUR21KR7vOn8nN0X
IyKFIiC1mm/nKe+0wRctJKfqrbbay+YR5OpgtsDTK+FRb7gzcbmhqoCMiudSYvflsZLBt5WORFR5
TWKvoKuLWHEYSUkHHZi0r+rN86u0oa52AoLN5fFYw3aburTKjQLM9rIgcMA4FAeSF66UBoDu8cXw
xid3nX5EpuPet3K4KbCEZsEXJD2PjTJ6JbMDTzUhobMUx1VreDYEyPjyj3j45s7LaWkSkJp38kk8
K2eqlU6rOtX6OHpJpTH7aSLorqsoADhLfwE9G7L/4aEAgTSHrsLMIqO40BDZt7P75VT56a0ffKt+
8DBeG32MOdXCmGlsu2zJm3iyTM+6mfnz+gwf3ISPUMpWMZpWkFE74c3+fWUW4eQ0p726xxz82N/n
DRv1HquLMLIOeBX8HdolsvPANXjhwQzpoGAGmFp14FupIw9Bgr1aExu6yAsBQm0aGzRkx1Wuligw
iblq5WGeuTIKJXAfpNHr4Chozn5yQJjQ/2L3mpjJpGu5DkrJa50P3CS8mqv5paRyzNeCWOTR+l/I
x4lCgX5JuMXkitV4MajNctLowvTlmAxxICWhgKqqIWerH0621CT4fKg4cjkY5xnwcIxeyItEweoT
9xR3+hY51WrVbbD8p2CNIAH6dbntSPRV0YzeIcythBkC171QYG+Sut/qqHsqv6gbymqlrljPq/ve
MKdQyiAMX3t4QfMpK2YsQkJciKHztJurNWHcNWeCNjTt4G5xDCRpiBSqj28SG3qDpax2fTJKsL10
VDrZncatt7pwZu4lGWE1HfV0tzq2rIckKYeCBRI7tPNt8ATlCFe2Tr2nvkvBI5byMBlC4Em/bSSs
MbZNNVoB+a28t0WnseNw5EY1C0tdSmHNZ1+F3FZ9eDDxcanRBdNiQPUhBwtlp9cL4cxIkbjeUgk/
prfpac9KasxQo3njgJxfisDHdVFrz/RQDZJwIH+0MUEfJwYCEMJuTZ7oaLpPmxyrvICbywgbq/J1
QSgDbBLSPc+IWl3YdGzdjp1un4NWoa/De7OPiYlbzkoDgg/dPW4W0uv2yzNF/KQt2YgIL86sk8+s
p+0w4EsrPtd4xGaTwJLi/k3MuJXVQi2fjz9Bf2Eudu4AzNgaQbpa7ihi/lonlYd1h5hqaXv8A3ok
Zlag+5s48yc3mtmcGioNhVEWhxeUxOtuZnMUaOtYSmfJ8CBNUqd7AAlubmQeg7TTHoqVWrQkHz1q
PUOJVeWPLYXyD98gmTGzNebGdmQ0sTAZqE0UkinJDc1ZrOZh9kndu0u15L6E6pzkLGfj3BiWed3T
MteF3AUCl74cjAGPORr/buuHoFb9VAxjo6o7yyzq/AEQndenoybKvqUDJDWR3N4PzOuChKPxJlVL
KG8zDyQu5ndKtSlgEXNSy2RReqX1fIa3RY8am3K9Ry/HI6sCMcItjtdpRnNuuW8RlgwTz1zPpExz
s6S8Zjbq2lxnfsYyto4DIyUhtTqQ0qww0cSKasrCsVOOogifjCavSROdi1uZ2Q7MzBOcKfIeBa3K
q+iusojgAaPDNkLLrxKaNuFvmZ6YJf686CKsW7WZ1b1JjVr0NR7rbP/WIyAdt7TcenRJyT+rlOm2
qyE56Eci4ra1a/6jrOM1tPEySa1AqQGxvHC5TdqEaGT2D+ywsKMMkPPX6Hmw7dpdPDDMUkarAcoi
CVVoUUmyOvz9kE+lfePwOM5Npv0zWmxxWfYPCqHG1aWMojQbFOsitd7wU9i66kbFGlROBhXEFXXY
evjVdsY0bOESAQEt2N7VHOpgDLN3Sgrj4ZDZW0xVGEUallB3J1u7mUwzePzRGOo5P2c+MTiQ2Xui
NpLhwpRYooLZEd1icy4BJTh14FeIvGKSkHnQi7i+r8HOhxhLvhGoptKF1K8Fd++yOGExMOBJlmee
yu3RWiEgLe2c0NsN/5Ow3mg2yLD2zbGCLb5safP70l7MAFPsPJL7xVnbG/gCeW0xlpACboWcOOAW
xqSV7N0o7HmbYKJ6YNZFWrQUt6FMrs5bVcnwOZtXj1D0o3gYduUmuVYul0ND/SgFqTI99RJvU6YG
KCdoLJezmBJxGQgml4ftoay7lv3KwE6TMhqbcOZr5aGKD5A6Zow58RSB4ZKpnblcsbS2SxOu3M47
3Z5s118Xypwx9udZJ8iBVtnoBHjNFWwCC6oV9DRWy5Az41C0V0YZqm2ioPGRoXwKw1iT/Tv0OIez
j69+3FEUL2j89bDboHnjtKfyWNKQBTn6kEN3OyikyqIWUr5Boa55hVya+cef1IEIveJd6UWW1c8Y
v80AtthKDfBcV1hP8xAArHMIlbgKaiWUNL99IVIABksXfvkns+h8ET/1XpLHfbnn9yO5NYPeYGqj
RpF+nWiTKHYdgzpYoP+jE1LxvjQWBFRzjgzNwDeC4OA4vqzQgSdqhUF5pBmzvBj6caDASXTqK4/c
I2T/caIHVg0GQqbpc8K12A55FPfx5EX52fSSOtJk+6xUL9n+JVISORvuzMuQJoCCw0jcIWvoRzPc
U/Q9ATBjU0IJKAAl0MuSYIkyeejqnbsMQDNIwPu1fwP43Pc/aZr3rSnVA1zSpq4fKY0W1be7jcOU
K1FhJkCltXlsDAMF2zNP6Ynn3iXUBA/KlYimfhEHxc05JQIhff3KTpTntJof2OmzHq0TXdYT/1dQ
AIzloefv4zCCiK+HKMCe863vGwb+a0cG2bdkDL+37XEawbcE8V3drF4FLWNTdxx5jb5azvDC/ogB
8IlaJ42qmdDlVfJCNwCBEDUMMuNK1O99AGeBqyVDPSvWow7/H1C/+i0ZUh6oZUaWfqjr2FK2hBj8
jsIS5IT9M8OWbXq8j+iZyzrDOhwaqjmnApnOM2hqziijtu592Kd6NJ0aP01eLkBrhXy7VF3vYDXv
usl4zncksWd20XxZbJw6HHJKY6+bJHcgx1V9lIXkNrklyauuqI4zBEiCfWZwfLIrDs00SdIp+65m
0NdWCTjaTRcXKoup79aM+CqAnUwv6Y6vsBf1E7/HX5wRt8MnLaijAbvPFwD/UNxPue+KpCBLo+0H
aw+4s14ujipT0zy9J7YfswMou0hGZleTDQkEYM9/DECOSWpLuL8buHAdyujY8IV8XyWP74DHFJ+O
uvii+ILksBHSNzQc6nNWuBgdBYj8pgtk9pO4jXcO808wUXlL4/iDqwzIXf9nYTrKKhwsRkXRqRZw
Hw/AS93emckD4xBxeLFm8EnMMPVCCvM6APN+DV+tA/2Pt2PUidh7B97ZhQ70wfDNqFnS5zOsXY9P
6DlUwtxCVUDE+u5LJvzQwpRUCmLxhoaND37HjEXkn4FWrT9kJORyh3in5hb+4xamnvCFiBei1MYH
u7xO25YV/Ei4lH6ym/Q2xUvscOq3vANMSEj+BcCHa5tA98CNtszkaZ0wpnpReElynrjhFtI1KCdY
MSs+l1j+ksv4eArwRLBm08sNPG0u8cwsGpUbtO0Gk7E1cJdxuwUlt6L5UpECh4jw5iP3YkjQ6hQI
aZdPmET+d/zK0b17yp3/F0/iovsJTyx0vTaP99fRQGhh2210bSaGs5b9WtaPdHhp3WAgNyLW2jN6
57iDolfPk7Z8gG5o45RmnIEzmfxd/uTRycSO23OkJPKcw9bd5+OEiyBnGKTfrdmtCTECcSOyesXN
m4R7ECiBY8WQvo+TBSh/eRpEipPp9KtLWZXxS0ar698Y6JyToyg/FwHXoEuoQbUok1/brUqgeXJg
PQq6MNtvkUhLzkE1ju0v0LV9c887zsQwEvfoMSlF+kIOKAZxioZFh71UnCpKoYUq5vjYqp/gjfMz
SRhELZqBnPpKYR4Z0X8NMAnyh6Mj03C+/HXfsE2vPtCMxMs8lLi2CmwGMsUSSKu1KYEax0JjiBLL
ONKZXIKHshHtn+ht/cnV5bQW1axJn22TwgWJ/MU5t6QW78JMSRncDDoDxs7Q2Qmwh34eRPzhRoi1
0iOP2XVrqaivFyaRFsY9xA5dH+cKawMTEwYcInjjz7yUtpauaNZ1dEL6WzoqU9xzGBNwUcniqPDG
w0cta6HvCGifkeDXHJPmlEw1jH0RlQ6jky4lVko2W1hBhUv9cpGM3shFhhWSzD6peS6cnZb1ecUF
gEcDFe0vRYGf8tyPxbJd5P+XIyBs+Sv8RjcDScrmiKiobSiyXjShd0RHGsGBiPa+qY15O6pyYI0c
ZSmcvPpM3ZNO2uBVZPQI+97AzfOry/Wtovq0Eb5EQP8nKrPoDrE3OqLGFAZzcu7EmZn/ldNe+8eD
IcZF8dntq+Ak86y+8alxlcTdjXl+Ytkv+bH2DFfZXp4GBtJjnhZDFKqum5vGstMGBu1WXXxWL++8
z5dsBHIQ8CqKd7AXQJDAE6E3goqh85KzW+rLMjKh/967TDdJQz6Spn/oqXmo/P7Kk8pQaAUxQzVz
D8emqXGOx9ZGk3rebX7siKMW1nAj9YYTVJN59i06cwXJASf/8d7XbmTONFZjJWtcxwBdh1z2EMYX
OP9eU3HOFEDd45trxmoVCuE+ZC7jLkmo2INmtVVYUnh7nOsrQ3LLHgAA9jRqShmFGsBaz3dxt03R
7K7eVyx9aZ1iRD62lwIo3KN1c904EEKm5GDlXytdDjAGybCV5NP/L2lX1IJApUF5rco7Dej/IOtd
+UBxaBW4RTq40IDRhmNabVOl3LSdDRQlZsfoX27jYe9zmFQ2dP1YeZ7N9Dm9540xyEtipuGtPYqO
b00vX4JE7JW0HVXg/Y0JX/s6A4juIFsd9FLUsHZRXkKV4lwXXTzG/PMzjvUbepag2IbXEmFDHONf
aWHFTN7DrxumnufAM81e+SABIx7nXi4xKPXUDx6DfUG/4oWIdQkjzlXHGzm6GkmB/gY2mEMaTj9W
SRLQRmrSpjCKtS3B64nIwNgb+8GJ9mWNuLUy5g3D2yiORynF3TLcqkU9j92et4t4yx0MvjJVvD6M
kIuXlQXEEzHMazwgQBhw8OYf0V5YiYkvW8tSwXoGy4xYxhrKsIjDPtI8VyPfr8xl4xmfctGgGMJH
YuEfAH9vGuVAHn9Xzi4SzDd7QKHmIyDUxSSau2L+ZvXKTSVVoYVMptx9/w3k7KcstC/0TGTn3Fk+
tI5wWiq0+AxmXp+ZqDvmCXzhNY+5QYUqcYvsyBlV6026DTMElP4vRd/pXcKECHszu/5U+/p/BwMK
qCsASaq3i+zMHviN8chAZYb1ruOgJHQzoLsQ8X0CjIaCrOut9RMiQKGmAVuXEshfTpoOVGK7o3M3
53FSS5RZv5W3RX1Ef3rMc2jHhf52qCehZa8yOutleL46Au7EdsxgjVyRkepW7+QSTzRTKfGDNYxz
ND5v6gAQMatqYsX2dZZ3G4tLqiBNsq+S7EKEkstFKVHyS4XfXLDI1DoS6TZ8B6fyl58jXj46myZc
NdHnkZQ9SahHN1z85JsSMkoSiZd6rwDC4wwH4R6GruM5SF8b7T/Qw+aa6Phc0JUGo+i2aD1bSoBS
gYx9VazMN6lUHKfnOqzanGV/vOtX/yNxxhGeredzPZkq2C3CcVb03IWjqMrVHPI03iLE8mh31B9j
V59dmuRkwTXWRBiy6oqPB8RxpnvP97TkGQM+vMwAk2F8v58FSRM8ai2qufk6cKia1zOKXN5hZVqh
e6w3QafcuEeqU/t07MFJU1co1mCCuxdJDWW7B0b7CgVQ3HVf7id90oIa5DZpc3Y3eL4+Fs8l/KS1
XvuVI9Oe03OOp4o6zPekDWfJSl53/jMO7JeplMi3ETyTwyaT1tbxUn3bigCpJMaXv+cWKAliyZzQ
+ICXQ+dsORza9GjOm9XxKwj7oxnUUVfFzcMJOwnXe/gEOgw1+9DUj8bO216RddKFon50GHMOVFIF
RuXj6AM6kUiMtu9t+9HqwrYnvF5jQ9BIrAo2MNNIEjN6pUxJqrpkBgo1PqJnENKc5O4BxgUiI566
awaLULudd9YV7Je9FLR3bsDtVcSneUaKiHrK4pRRx0ZtokXANfxd+WXDMwkw3LLCimVz8YLsXGLO
ZSxgLpRWVdMdyJ1H1T06QXG0H+1iBwut744G+jxI3nDl0iloBNfkGRrNk99SJsJkR+FrC2Qwe/Qv
DosYmKhdqRzbaadPaQI5o3aD1cwjLxtL156W8zM837fRBg8PecP8TL1IfRQyQ50VbQzk6nnQvoGm
yLYLf+WMtdG4LUlWGtuKdYPdaxECurB4UG5j9Za+gv2yr0N4ADW7GXYKbuy3XPEayTKSa4wGd5sL
6vrpa9SGvxknXVF94bFjhSpf8fZxQQOg+2ra4ngaX7NF/BObJ+/Em+8BU8WjJeenu3W7im/AxYTq
79rbvJVU0UFKZZNcILCup9POXBuKZVOPubyNM95C7RbpJGOzd1/W05OcAUaMUK3QlcrWqoyMPn3o
QsGy7z+pMUARrqhXc4E3T9EkBQGIxwzZVvZBMwrndZ7Kig1ZoSuzTH1lVN3QgIu4D/cUHpPBFZLL
xE8Momru5hMQk1ZqBGw+Lp5pva0uz9LISpEq7uzf2NnQq+61QLHHXPMDBEXuG5JsNUAOpHTGD8el
WXLRQUEQ9sgRqoyd/Y2aqVBQnJfcFii5r6TX9AklFIVxprcIVTrWPFcn2J0sgG2euvd407Xl7yzy
kL9S1dp/Ye6Fn5ExPaFhZ+PvUIROgsvgEJOSKBm+dIBjfFdUaYXWu2//MqLsafkTan9z1Fmqmlxs
RVBOjfCVbtmr/rfVVYY0hKTmBDKRRx80o31ecG8Ow9HURJPdlsSORdHAma1d/r2HLvfwJp0BrWK0
yD8NmBT+Wqxm///4h7jIZFjzjvVv/115bf1ivoWnY1CaCMqzP1oVOQPNLQKeXB94RX6ORKTRI28h
y/vdESYFu8K+A0LcPOZ0QyjyGtrkKBHsFbchtwmMOzRY6GA1nIiM/uh7sHI8TXjWmT9Y16IUuntV
ekbeKzwqY93GgYqHV0cfKKWCrj3J86qmCIE/MaOCHJwQcJ5DjVRr3LpIwlE02Yubqn/Ft5zwoKj8
q9dRhEEuY90M8oTpVYLuTpfxPIkkm4m4/abBIe9xeyS+nNoygsNoyXNnGNvjJbKqB0lZU0Y6ZkQ6
vksUBncSlFCKORotFtw6iKzLMZNEX55mxIYzAiiq2s231elE4IIrIQR8o53ruyMbSFqsfBa0VKRJ
CG++q/OXB/+10ZSPfI5+OnpqWKYMdL9HpRZwWsAJVLc3zJ1FVDL30TC7GHQGT6e4+IZ7WdNkr+6x
y/LR7cO1m9VCXcaK+LEJqNAbblwSA2qwTd4vXb8ypVJwUonHWbWx0Zorp5Mukb7nm83rHs1Ruehz
0ZQIvUX/uIb3Jb4epSiSH0XOJkDingzt3YVKGNR9z/nnxcERewYdl0igzpTyreSpfyP6Rkh+anbu
p1e643gfXr5ZtjSkyPxskM35RGF2AbJlutHybdopG3Hibr8qx/MTfkKw4AyeBMaRHae0DqACJlMI
ift2Z0flY6GRT47WVPy3/81X8ohbh3lbBJ1QYM4HCfaGEpZ4k5lbhiHMdUKUu6gtVpB1Ey8LlSty
9AZMyMN3TwbyN76ViAxURVAuXVfGiChiEwbcbDMwAX/DBYksCNsCRpko9Bt/GCvEevnBzE+yx+VS
+BLdnn/+r8HkMPrK3NwQNRDgGANeaKW5j486t4TIFI6vVn7w1tLb17HxIY1D3X7BCCO5rLjTJEw3
ft53vjarJ+B6yCPzQS9cBoIh1tgLRNVmf/12u9S/zqEdwFwnRFVYYOJQEOReXXQbCMHtjYeQuAUf
vcOscZRtyb68g88RqDxcB4gcZnSG4vL9vKrljy95v8vxLQsUPIXd6nhtVjmhtpGWGUkauOCZkoaK
Kh38IldGr3NfqYrRR/WVVq/mMphNnsnBiKcwxTPfdLe0c+nMUBlLmtlUMO+snsS5SI9NFEmt4UZ0
m7dAA7Z6FUXWt3B1JQgJiTUaOrCbXOGVZz4fTPZJUBwtGpw3gAGtaCuO3zrATaApwlHzGaZ1SYlg
aZ2LkvmUmLj9G6Sugnf9rCSt4rsfQtczl7y41lc/niVWcM4vPxplcnC9l6xgHkPc7QqO+2yEf+oR
0CTMVF9eCeKBN+p619WbI/2pseR57QTNkIW6twg/yqhJzDQfTBCcVurzNli6XXxhTVE+fn28nCE9
Bmnegj0pEtwiXe8a1iiO549qppsw5Yz7jtfFlj/977pMDiY3so3ykBUTKTO/y40mTPCDQtbypR99
KUMiYG/O9eMqx+9mOQKMNwx40jHy67rFX86mqmCewYSloqpVNYbmIC1hGqgTqXNnJj9H6nZB9y3I
djqcixrxOIg165z+tUFuH8LbOlO40aeYEE8hEpam9RHlrtSdyslanO4B5vA7ULLr180nZkTqc76v
v/1Cdlio9rCRu/LkGRkTnKGqzFebPw4SKnbgo7KLfJLj9qAt7VYv+IFC8V2EALRj8nl6tcYQws66
4tQltPb+tUqt8yuzozDuz7pEZJKWOFCbA6vxX5JxSmx8M24+05vyANsUXcvM4aOZKSChsgcnUo39
a9dGtrQ/vdgpUGY5R1xLy0cC0UEcH0wj/367CVDFsV9U59p7GZ/5IzH1CMg2LXwsCLfEDNoY0JA9
ZLTdS9Ypi4n89rj93Ep960EPzdnDGUZoE21yaHpP+CxEpBCPZ5bVkqxi6cRBDiKrllEqymC+w/6v
1BzgLVcgFEpYuZRasWv8vgAGik5NehcP/44sPAKl1LXTGyeM9qlVSD9hgk1jasCCG3iJmwDXTNCC
ZiDK1csmGMF83ZSIUki86IF45h/oO7b5JGGjW0sPD5He0ha4sI4q9/NL4BXoTtWqLe82+0ABnU80
cOa0llMMymaiahM2k6ME93f6X2VntIXuCnlSajVSIcNpr9WZErq/FvLSYl3+qjJdacXxw8d5Dsr2
niZj7YI2Io8RsTP0xURShwA+crOE6XjAFYYWGqgspK7vZTintCJHb1xK3SPcCa5JqRl8v/APemBe
LSgTl8gomTxb6l4sCNQV6hta2Q/1xwHrVNr5ZJ9Shs7FnMCbx3vKXdFAh0otp++ZoQHswxOUOpOK
Cl1CTd5x6ix5RjwDsl7CT1JgI2BD7XWiKVl9ShXLXTImtEBIukWaKHIWXidpJvuEqWnjQNUAWJEl
Diy5JJcPymTvjSmGOCs82T1YCirMPA/f2moTqEN7mKBndGpqssetjn0VM4SAvm5QMyGEEiBIsHMh
4Ybl0Urn2Eqpdjb9I/HoxUxcKKZeOjW3c7JJdyBgGvO8ZaQ8wi/bOs99R/i6M0/WL2Rlg5hI5Tfa
69odZ4h6ahPEdql9atiVHvm5qG4xJzV/ia+u2n/N/hJEOiRADV7sDPeMhlZQPf4JGM2d17QYl7br
TZzOawF16sfTI2AWsWPqo737MwDiAh5Yw8O0hClWtyx6kBrSU5CwTSIf2/1C/HhtTuL353ugo7KV
xKOSPpvR1HhxcTM4EhTwHONMyRI6lA6e+5ekO1o1H7ibEhYEUhpSC3FqxFoOY0ZGxdE58oTtsm3V
QKQlgdvecu+eJ45BX8pOSTpTg49t6WIs5cGiWsppTeCv3FTzqnOfQ2J2cGCOktO8kskznUP9xeEK
mol+Ta4BsK+fYv/HXr4+fR8ucG/0hA9zhw15QLNfzGtswhh7Y0J8pSwLBQzb1pIod6ExZEPaJrgE
kYxLBDNh4PQJYNk+m0OgACXcxBVI3wqRtGg+YX6LgRbg1jDHseCxRjeU9cko2KHFUX9JQlNmwhX9
Yp3FcgPsMStWqjl//UaPTKLjXHgAVQq8aTdl5L5kF+V2Ij0iatvwNmbhq47pHAKQyj8l1e9LXCEM
/IE/amfLHeTRS8Xq8PcSdraB+1VDLwSeumlR5btaDRCOFHjFlDQwmXfEUDYj+vW6o8ZNMwa3YJiN
tMRBom/7qXujNGhjTypgeG6wP27W3cfZOsArJxpaKEU/rg3xVoOOtVhlubypGa+WqO6IccLZaqsL
eZqr3ZB4i9g+cJeZnGNk05jHHSXto0eg5lBXgnkFeIMkxtJt7WFBDFNHKqCnSu+A1nK/SR3ktPJZ
6eNHbdjWfCejeIuB1+ibAbw5ZV7DlwITbMAB1jnpBqZBzIv5mZDykhP5LdjS8/4uIIVgGDGiWPQb
QsMPCqArP3l2JSlUF01EE1OxrsASqJXuZCLL4UKKGIXy4t0Pon7S5Ctk0GE3geTOPEDao+URQfan
E3buIdbt1S1eTpMOkt5x+nG/hxB/TfW9syWmT8qbDi6fCa4LvJKC99NSOM9VP9CGFuMwiHkW3yDH
vZHyztYN1KJZiikO5jfC7X7vMO7B0UnSKmmhL2MpY3xDEAUWdxeEjyqph+EcndTB1WPA6IguwJlo
LcPo9v/lO80RKOSW//0FObZEHrPQSYSE0UX5R/nvMf9RZROngfwn/3Fg+32vG4Z4bQPT7vLyRIMq
E90dap27DmL0rb9J3T9Im9UtbdoojbOEkO8EAFmNylMMK+gtmeccWTZA4yq6HNLmvqqBlxlclJaj
xNDXEjr96xHQojlFc1zvLpI3b6+O1yrF8SBYvCpI6ElKaPaSo9CtTWHrJFMkjEKapfw2iDgOnIo9
3bcU7ie6GKo+jJOTmx5du4VZsrO7oCvNmKoTRoIb5w+0mXUkuj3++Lyoz4y7K43RuLDJtB2bdr+r
La3a5yOFz19+RVH6N1Joqj1tO1eiYEjI7KZRVqINTlo0A8YzrrvsFWpxbIlnrIv8BfdP5Bn4fnYQ
sQ7hbRkaWl6IowmpOSQ+mu2fRCOiL9UfzhHQLEZTbS96D6haP8pUL7qkLe8WfnvMrUAIcMsE+G1V
M6HCf1BTsdHBJHy7qxJ6mfxoFofVCQheOKQbSABNr6xXr2Pulpj0SWOFTNdPD7mTEzEAFu4mBSgx
Iqn7OQJhYln+EfCL/BvKUBhfPWHz3/pYdrrvGtMLl/bbtcKhjve6wDuPLLYwI2pdDvPLUnSKMWwE
6rAb+QYqFkki06lS0BpwBOmP1sqiUD/lKRkKNeXep2+JwYF4c5Fw17/LdgXIPwTWCtO/CnpD4fqz
7pyJI6Z+XjnO5rE+WfntScrDmSOfwaBk3FUrW9/1nn+/LP0opcpCpFdCfqPOvUzKar2vz2qSp/+J
yqGEcOhox87ItARP5ipiEdC1tkuZhdrJJI2Kr+k+1Vx5zA3qSTG6qLW/z6lgyA6f6ylLiSBZK/9Q
PFdkdckxrjP3HpnHme1NyPX84F5Tn+W3x90t49ejHQVLW2wbsiqn/b9FS3AmRqcdtP/FdvtFgKmM
2tw7t3EZcEmVrbzmv5eBlpXW+Fb2l+8yzeJopNzJkvVG07adBBvcWvBd/Kkdk8VrCflwc1n806q2
MWPtmN9+4eG2iJyuamJfeQfXIpByrq6/4pGff/0pw4ujS4C3j6k+wfA63oB6SSArvJ3TBc9Ykylr
gFZsVPFk5aHjlZHB+2h+54E2b3ci9zYR2TjhUfFnsgIexOnIOErc+/QuPLQRp/Px0GmEz/dnsnGJ
I8x6hNH65SWDfEyanEu+wO+J/Y0Evmf+m47seKbbYe6xouKPzaKShUOHikYM4gxhPvLrjnCC7KXU
pe2ZQ52s6foeoUB2XfqaalQ9z5VcrXdVKMc2KaM1rttE+Ld6VO3Fd4/+KEPIu05pw7Tfc42CUIHu
DteOAFCZOKZijZbmcKY7JhWwqr1eKxqBC7sovb7uwZVDY8eTwlCuKYf/54bzU5uc2iHT4OxGjJGP
jwSHW2a934vBwdnF1XxgLAYmPhSzaCVLB7Cb0s06yypXik+sIKBYLQg33qA4QfJ4drnupOCQ+RfV
u8fjZiNNkrNK5QayaosEZrfe9OnEBQkEI1fPQXVGwZsiLg8gQZ4/bM6jpFbe9s4AMzJKbuIt1ZF2
TQvKMiJVutV/un5o9oda6IWOJq8fWzR2eOdQALG9d9qVZq15NxCZRYrasMjOuJJ5ybjYzWF55GBG
J4asXLTX9Lt0Ap7OZcT1rQ9/GRbrvWlpnYlA+gNbRSsFn1dGahBseMky1/6olpl7R5MIYOsVSYwL
02NnkaX8wpljTyn3RoubV2MoXPMRXb077cx5Hk7ABQI+GzmXnRPFOqgZI8k8PvrK+fF7k4R08fIA
+5lIBPaMkGND93gVWsMi2u7ixh8mcQjdcH0vDmjQ77LKeyCPasylQ5ZHhnzdmTRAzg0XoCGUNjfn
rqpNqZbRNUsB+YLZeoSh+h4flqN2RAHHapN/kdUIACq7u10VzIusmtRMJXY4aH7XIV56R0liTW96
GDCH07qfZipF7C7KOCHQkLioAkodPxcZ6inmrlYiJ0ntCl6NKk87toDtF7JGKlX2NGkWDL4itmiP
jKFFT56XU4lS+qDssXmasNkxlc8Rabt8nuAdIIuYCkY1bsWmUMGNRmgvrI5pgcO/AxZgTj6Fot7q
I/vnzSULQtaX5mUi73k7Q1LSqSsxjc/9KKM+mP/yrWVrB7ygv9Y8h1JULRYDR72qzYbFjRd3vh/N
2Zsp67yeha01FT+q/PnCdCVc1VzdaYbOO3htG6hm+VHJVgj5bopoTOTHUTtgNdMhan08121Fdifn
BwSS6a8bIY/MiqZR2QGxDzcOpGgtrLliOBF18Ymv30sr/8j6tewwMnFiOXicrT+Fd0RBn0ZmZFda
xaMrJLoHMvPvDpT7iCgCt1e/yjwQYONzT+PawAmLKz7/CcHFW2Vo3SNpW6aUy/FSiROLJe8WfWyL
bqRri63tMvC6NHNZ0+RMeD7d11S5dwbxmOYvJpuzn/O1NIbT7C0PiYv+9xrKMUsJUzwkYTJ9Owrw
LKURduDdAKBZedYqxuaCqmOHGZ676cXIgO9lrErjHDlexAS1ZE99tSo6sQ27JdtmyUgqs30gUyRU
32zV/J1/xI3Pn6noZuUvbARgMbVhCEnwC5YUi5o4rRoG7kxjeDQihvTfl0jRoRuYtl28/sej8BBk
WFd2zLH2obfY5x8iKx7El7W3RAZaH4/oyL2Hsc2wJkSz6YU8Cy9oeq1efZzvG7ukk2fly/HGHwsg
HADV5+F0gQtdfGGUJtO0HCDxufV1TStXo0iCaakUkGKAH9X9kUWeaGCArGiEfBu8APNambjWV+v5
5xr87VUYItYQVg3uL/81kM+gptJnf6izmgMF85D2U0794bLWrr6wcds7RnElST4nvMYohWAZ+FEp
l+kgoprISw6ZJn0Ffyc3Jp3rx9wr+AzWTEpOstNJZWgL+S0TjR+kgTkcr6oFenaiqX1gyzQgkaQ9
54/sgZWx1Zmt2jjHowvSlg8WbSIiT576sfEjmSmYpQw67dT/3EbSawhaEONO1XboHS2kRqybCGA5
a2y0mVAcqo41D/NCmCcZZndXQ3vcQIANg+Cz7G+u/t+cxZEGj3Hy0s74g1JFtGqeU4priblqlgVt
/rvJjNWYk/US5us4fyHLsKhuE+eKoT+VaeF8xWHuBChpXZLI6R6M+mgC3F2OSbIOaKuMjROuymX4
VWPgbQ/Kfs/VA/f7EFieBAbVtqZuFjXKliEE43WchkV0+NJ778WRjaifYFqAe9uzpN4Yx5nuHGhA
uUkr8outKH2APvW1MqHT89+n06WEjMjEve80MO/IBZlOsqNqqBKcsd4iR+gUDM/vUAMDynfpnNIH
30azBulzgSUukkceClWKbfy91SGqqE+alFFk/vnLC2QseMNCh6fgrZNSJlvLXNaqfmk8PM8hhEPy
7Y2u24NTumSVj+OW9jRSyej3VVKnzJGKShoClifZSaokHF+XrF+fHK6FKnCeRM11j4amddndmB8c
v+0s7FZIrcDjsrn/APfzHNkG9Nmq+9egmNizCgmWbvHNKSW+nzNl2oa+Fum7o+5tw+a0XVS1Hu0p
+ZTHUf/d97BwSCBgPBrdTAkKWIBsVSk33h4ZGr3dbVufGOQIR9kWb7Qr3dQxj4wGGr8hp0lmtZYm
EhXiYS6oXhrkcvTwyb/9Oq7TdskUtqejSEXM2uIYDLGlDkb+Uk6ks+Ga7tEO6U4YmoA7T/WBbsBx
2YY05fPNHQhmdj55VErH+nHmpgrKiAAoN0uobB7jec1oAOncfFBqyZqInJeWXcBqb2Cbc/uwc/5K
Qg4sadeaeXcOwkOQq6YhcFsH9FnfopvfFj1JyJp9BTYE3VZcvhF4WPmivASOl3+hAAciEHSRSLRc
6odfJ65mNEs4PBq12au6dVB3AmtFQN/8oUA5ohogkQSVjJa1lUcSOlnhfaKdkSLfkKs0W9M8pnjg
hBCvQwKGDZp6kh6jqRh3w7SO/M2L9GpG7G0Is1XjFVAPI5quKHP7LkrslkY5DIsBpX8LzhA4Dgwg
Q2LMjb/4e/zFAQH0OY4LztYNUBwHrC0VkFeHDZryxPOGEL32KPZIZNerYEW57pV0pdUlfRCaJWUh
KMIvYBqCT/CjM8eDucGWDJKsHS7ddVq941o/oTwOZEUzAjS9SJQCMmt8sMQNoGtsVg4HwKl1WMjg
RR9R/U0a6yo15jFE09OpNtNNeByJJtOMxo7aTOXlW9B+Uffz1pK77ncEv7La7j1IXwAOzN2pOKPQ
SpWddC7GYDeMeHUdXV4jaIYKXAOFWSWfe6cqLpUCAbrMxixqvlrKBvUWXGW7OFiYbPqqYhIbs8Qy
WDTlJ9yMwHoYRxLsPD64Fymtb7/esGSScnSh9thz9wOiWPAkRpEtnYCd89bRtYVKbpRJKzEefxpP
YZBnnFXXy3odOFwgmro9zlEtXhd7EMUdjmjY9PqkgNeZ8zx3k6WcXPrxhH8WcJo513tXGT6f+NK4
L5baXOf0aCvm7Gbm2grp4ZqHDKQ3NZm0/kmLzcCneW8BpYBcFFukXIA7+Stn83OT1INvqMtjm9i0
ztFv41MlcluPiwoTvHWEeCclslhWd86HkctmnQ2tETo91gSjiu6xlkIk9TxwtAwkz0qNuEHeFr0f
lkFsU5RjTsha9nIvIBIxCkiYzfmt6UEco7et4PsFUPF4vmzMF2iOby+y9s0THiTw/SpNCUj+hgTp
xlK+oTKmDgE6gf9mk6POSjNnws/IFijWvA3AH4dozv7oPXd+qfHxca69gihYR0TyQ1IqcYrndcPu
6gVginp+OJGz/xMx+8t4M/Twn8LHdkVqK7gwOjfMdqpi4n6Ve8fQ6Bwz6Bmo3uwLY+LR4h8m2mtE
/7nCqRU034u0lnRv7MLgmklpfpxNd0B8wCs4FzsLQPDrGeWUmlCnt7M3RtmgOSwYTw1NgQDgQakr
aQoRVLbn3ZRMIkLKpxdlTXcny9AMZkmtVk+JwL05wyEj18c+rifFydtJMpWvKD4RfvJetYXt51yo
9K2eUad7hL6VarAYGGCBCQaMWISnMO5EkzzshiB5ss8phrFesrratdGi7lmWPtEzbTe1E9eLS+2W
23cXvoxd5cKbIPwS2tKLqQr7E6wJrzKF2aiTbJyLkEQuUISISwQx3ZojM4AigdCsOWfUu6e7tCZv
gRSvq1FrEwLkzP0Wh3Jt51rWA8E8A6AnLoSoCpiSKcxoesOMe6aVxrlBzcByX+aP1eWyOGjDHgil
5cawlb7JRWZNOan2alnGOkdK6CiJJCmqBupvt5ihq0fz2Yu2qUTwF4DcFQZnpzvHcSToJtV4fBvy
ev1xu+9GFB4gJ8Z+vlFE/AaLeBI4c7dCUvhoeqIebrdsEm3wEB5Ysgd1PK1pb10kddQpenGHrdiH
mrwTH6L5CvmfsLY/ELSwMOtvbaOJtyIwMu241zPx9pCBBAwXp4HeBNqnJ9+vuAJJ4TT9YMDdaxpd
biUHbBdvzPgv3Rcmg/lqR8T299iiYNpafNWh9F9cAyNlsEzgD4RbIdY03vQYMqe+u+Vu4qlnI28q
ne8Rp4hoqX84inPRzZZ3oW2VqVo0YCxWPjTyi2pRWTJ40xO7Rrqykvvb713FWaRBXGAl7ut5JkuX
oAXj0DDZuDVuYqlft+7/XVEv5OfWwJUwsFsvHTRvbLxpLtKhi9AkSmcPze9WqGM2ex0FZFdNy4BX
cjCt/0j5gqsSXV4dcHLi8/88VnhqvrP0Ulc1BCvVKDfyVeRxCDupgs8YwY1GIVpLBX8o3aLyMQTE
bq+9nm5etdLSK1KknHKovnuf3BIUjCdRpC0C2wBwoy6U1+ThBICtvdP69b3+baM8ug4AYv6DJnXq
xtCWcDV0DI39BrzZEoD8VMVx8OnQqE1k+uLqrUWRXeo0vg37+bByfwPtTpwDcSmHlA8PzKPHrlX9
WEOQncQqpTkVZ+Tfe0P4waP+av+9UoqAdg0Ao9/O1h9S7CTV7bTxjtf2+up3ba/yEZZ4GLQYHC1a
Z2xl/um9D5YBxeIQGAQjD4cSCSjB/OrtACilyYC5Wjl/7IYIhp2JQDkvXuQTd9Sq4SLrC9GnaliJ
hw3v8OK824vMhtfLT3Dx6hTCNblhyGSOF1oudr9HNKECc0y0yE57DwRX/z5j11V4MJ6JnfVg/7oD
BA+uQ6ImRaf8sVAYLmY4Oc0hSkpKmte/BoVXXer6mBYGYtZlOG4SbmIClXgMtrCPjWXAcobw/NaL
avTVy8nbZxl0lzFkUowfmCEcZYnqODfnEyh97GsIFq6Uq/bEsvc8witnsKo+8O5eL2eeSl6B24UM
ZtxOCaOo8MW9y43PIefPwXoN5nxRE0FVjKin32EVBcBBIFALaq0syG0kHCshgfaZuLlxx7ATzn/K
XPJgRwd7y3oGrMEyc+OO1ew0KTYuLMx/DMPmh9buTzHBzVzUPpf5xI0/4q/Up3W0/ZUoet95yrq8
hzZREKhlw/ncFPC4dDj+8ne00fjNEU0rDcXWvD9KB7IMuCHMrMRlmie2TvDpg6EFtIwhMy0btIR9
hMJdlRwxYrMV+UnZrnmi9QPCsFR//ouC58+5c17jIPakQpZgiGnVrMQ7jBm0gueaDidaSTUC0SeF
+crUangiBx25JNgUHmRvnE4iFQfEPwS2spRrRKU6K5UH3q5inhzDTW/++Am621zjDtX9KRlUr9h+
D+E7XyzSCpw4PlDuL6RnaouIApn3eRHpSkVTODWnlnsXEhAIsK5JjTurhavYTiZBXAsjiu8eYBlJ
Yh0aeU6l0TyBuohAfdbXs0EWJ9NLMYHvxTsJ1tpcDv15GNwEtlfp3+0tgTfRuWHhndywEw6dNV+T
xeSYM2lvVk6DqdUzmeLNH/Qx+pLMr1e2CBdauC6hXhnb3yTBi8D0zkE50SuJfUaEh3vVYYgdg9SE
nWeET7sSzGtagbhqL+jv2QqOTwWVhtk+RA+8cfDqwR80+gA6wY8BgcoS7LqFiytsK+SK3eiLnpbr
1tHLNWROu5cm6fsN3hZohNQRFW0gjm5CKj3BV7CFnx54jpUIWDenP4vi5JeFgYG4jjtenIcAMfNf
PtJtkpLCGZ91E8guBXEXzYnhAI28OnhAvz/ay47lHiYKLtLH2j3+oqfzAeek0dMvPm/nG5WQQ0Tz
PCk1RfaNpACUBMUKfhYkI9hRPthCPYzN4umPyoI9bdVFZLdxJFHH+FK74ZIm/77SLpGk82JW5yvs
UHcMYUDIPDt2p4S4165UAr+LPtlEpdV2PiSrYMPJbmYJbAGPi17fSjI6l7G4b2qJwh81CpnmUdAe
+qqWkD1vs/NaiwX+1FQOZeNlc0kOht6jm1UGcV0K0rF8QedC2rriB0AuKUeJsk7o592wAhiIGwXy
/Tm5Xu3ay9zu19ag8qNCqoWjA+C8XwyLAb8SZWHRPmM9IQ4fqe6Bgx6F7FnaighnZBOl4+90saSk
z+2o1FR0+oZzmRtF6kcpUMDk2mmJ/vTOVe6yC5wgUYXT3bsH3q3rbJiWL2f8MMIP6qibEh64irTS
QoQwrj3zmsj14cjZFs50sMwQTafhDJ1n4QPB0mvBhHAji50srpoXV+Mp+F2vQuwoosSEuN1KaPQe
ZMPoqiiglbyP8Z+gVKpq27LYhSk1MsYzsLOZ6LOUD2hE8PMH8rB/an+nb8Abw8I6S0ARZAOvCT6T
WzhjIvKlYThxqEIegePgkRnntj8Ii/eMoMKbS+KwfgntP8SBQMyDmwTLC/aA+7JTk30B5BKeLCgn
5Wbvx07YNfdIuNrBGZoQDEC9FgyuWw0/Is11B1Op54Y7krEWMLeIXK/1wX1JJzCHejPkOZ73pG8c
FNvJgPY2oejIiPD+C9vBh5V83KDmNXoRO7bbKaiPU2twmIVepc2XaRA4UtIe+3bsQzOE+1QLkPx9
QVibFOz3833AdBtgVY5AcfUVGTPnjjItpwRbLJgJNtrRm+41orRBZ1D4aE59kmbROI7bFwRq9EaO
3wLFbI08yRovOasNm0mYoThSRArPLAXE1LySo0i8YK+WpWrvWuW3rWnI0BxN/Uji9qAR6U25J7/Y
Y4pn+iGVKrKRJ8RnjhWwuOgYcPthOaYsN+DAzOyRK+fkwmehBkes+y6w5GOgD8kqB2m7HTLVbc01
GUnSXIkmNl0HECfS3QR/AVl8/cLT8mUcYziEiVKK87P4SDw9gzlFi2yQI0EZzbBMVc3AvpkY9doQ
AxnVyoQ4ehB3chQEn6D7Db1n+Uvn1rtltbWZYxGF3N0bWMgDPNw34YF+sd9oWEus3ZuVC84/+CEM
gsAHTGJZAAxNMUYYOkau8jdsfFKWfyyjuCHWMmSHcdHJn32mppkTHVuHKMWhbuG35/qe5uVrMCUg
z5YuV5gSRMJSpwEnTc8PDmj1aTMOohpNzH2bkCRWtip6ajbuW5sgv+ufURt5M+3vnyhIsaFpYf3e
ZDpYEF1iSsQa4fw1fTrFDzOHDikGdMMLdTP7c2UkwxeI0uFAgpNliZFHO/YeCYuYY960Vz8lVr5x
LnA0RZ+wXbfvkNvOOpVu8naV0zJXubNkJo2aHLoytgz4lzR1EbIi45xR4yVNUxXXswmZd4xyt1ZN
XCHQ20tT4dkPtGANUGEqvrYJP4SqABQzyHERsEF1I+RnRSURMLLK3FBJM9c39kkijo5rLKwMhSM7
q5fChYVdnm8R5kX++Sp0Qa5pGh6yU+ZBix1SecoPgMCAzuLJARB77KcmbtQbiapAxmvh3kut/zaT
amCQNYRFdHoiFl0lNse06fojCO7ToInTL2AUiaGQsZyMFS0+KbAJ9ZdO7LUKQxfwk6WM42RZM9vr
fRhVaN15ZkZl9JxSmFGn+E2p/DXygDguGI6JL2zTwmMIVWF1XMC23FcPBnwl1ArKfABCyYS4P3NS
FLbm+3HdgY62URT9EBgIWpllvVn8K7Hde2FHR+DZkjJCi+Rb9ZgYUmpHmDUkjg85QfkNAkTLAIpP
sbdBTBKPZjnmiN8zCuWQQa+ssxoWfQtZgNS0dk8R9xzKGnET1y5euteScFl62zke48qaBrLM1J5+
C/UkM1btg6PU79cTaXapx/9zQbqAd81pAat73RMIEgYHx8JT+GSEzjIU4+qgiBGpG9Xu/CpMetes
SyE4McHbHkJT/AVbEQcxhcpRWfPbn+dikkvhGLtSyekIN9BtRmm7DR+5xeYrBfpuQvrh0eHB7gA9
bYYx/Blj0mQIoY7ZVWH0fbM047TsQnO82f+ymecqRJ9aT2Y2YqPH0iKUw15vL4E6lT5g2fF0EJpd
j3nc/+lC+0zHbBPm2sTuenOTK7n9/15o0ie+InidvdYo1h+e3uZ3SWR4ygWhIWwkIvjvUhVzFotv
B5AAzWJh8vFWlfjZ/ZkeBvphAg/N7u9Q3ecbM2uyPRKBD0rmHt/z4VFmo5Sm7gYF0Ci+VVZGSIFS
YxKZTHlyLpJQsyoJ4CqOGghCRuoYemGespdH67rFCjd4ccJhR9L6pEObdGmir2yflj60YqqRckaa
QAjMoh0m4Ca4vVZYbbzxcnYyHSSQ365qzcxiKQIVDqe6aCP7fSVE9ifmdLpSOf3XrRyKr819rzXR
xEB5KsXeQtDc5zbnOtzG4aRLwU7w28fMldmxGLQJmGpc1to9oNdlhGmzuWuTXfO34niYq2hSLgou
1fmEXdo57dN7TUMy8KqpjdlWbN8uNntG3R8mLSqcpnPjuFL8bINZN2LaXPR9t5+2Ox2KWX+czwT0
vQC9yVwDKS75M4yASm/PfdFMyJ+9Y3wi1Y8ra+EaZYzyxB5LuPwUuVUZGRc7JuBEZmipIlWBMP2D
rpyqtBVrANELgZt/i/udTZU8X8F6NY9vhBNXXzljGr+CgngrF2wGb8XrruwRc3vb/+CYKV+c5Fl/
CY82LvwS0UCzNGTkJknxZkRfLBhGnrCCMdpqKRAkdBE3Pnjmpr8uSKjSZqjLYJCzVrDDwP5IyYWA
25ipzLFuWKgcSeZ2Tsjwc0S9UTTTIp8meZKNMLn/paPZvbJJz/V7IylNvh/TQHyM8O/QqUtd5UpJ
6pDIKN4APKNhN+QUf3t07mlHJZePuZlBPXzGpOCLtrV1E94ovoPDZPnXcpgXHyd8IlyLEQoYE4bh
39bJ2efJh3SgdJbzMKut6TAMxTGm9yU/mpX1lgxEE8ebmnNlTBgyfBvdDGUxgrBb3cBvncV85sED
rUf1Zs/5uqgiK19ZY4/HRmsn3K0CLFiEJgM+B8FSMcB7vx8A/nscO5aclsJ4FfnuQHZKWT51ocj/
GCzykFpdbI3BuvoeGG1MaSup2yGgJMDDVv3pXfFLxoaJoxuVIl9rv+Qd661XxCkRQGIgehXtv9UN
1JtHr8UFK0HFeOjgiXniTgkF7jmC8TG0VWwywcd4IwcWzqEPXwQkg3fg5ogYX5KdFxqtkeyWxLpM
9+3BXAQtSorI6jU+iTtnfcf99tr0C7G4VPW0Un4UA1syMLQZgIEU1Y8zhRc5k99aLyi7cXpiCu+3
vGhGrDUl4U/2JuAFetPaLrMIpnFD1dKgiUrAIRZuknZ/biIPuewMO+t6fCMQku3YlexDnAbUW3QY
89dx1s5U/wg7fs6x4JG2OE58m0pmUIYdW8yTEL3GDCG4k7IZZJOUL6Hw9Iz7aipVFIOiE9bUmCrQ
4z4tMbvX8+QpXaaJU59X3o/no/PipA0gbQxrOCR9fdKR9y17KtIfevg2qSeMPsASRbZpGfVW6BzN
H0ZOlwWFGk/aX3vsDWEWwGr2+P9Gzkfa8PReS1fl9HTBpTXwGk/s5mP1C/YKQRasYqE6KHypH1mf
rmmC87YcHvin2Ms9KbV6H9kzx3ahIsAsspel37E8CjHZpQsj1SlTOfAmmt64j/4Ta6tmK7T23Q7X
3khJVLyX5+EqALgEzmw5HfozxqS+USJn4xQTq2iHawTu7f5eeSXIM4fJ+o/7euIIJtMh7CaUWrEQ
+PzPs1nJUhG+jbAkkwzoP1AUqEA7dl7Vk5LWFiO4KrVTgf0gA7JnkyQ0ARpksgyST6jUmfHkQD+o
SCtHAiOEpFVIvGprp7BrIkl58zy5ChdzgzwLMTwP1B75WqbLKX8MNZ2NeD9m8BvuHVTuQaikgKB8
7o9V7bwUHfXtTIWJDgaXfbjsTlPQbVo/QhRXgRM+8PNTnHQ4bZmAyn2iZtZJKSOPSNp5Sh5B6/Uf
EzrMzK6KpjMFzON4Vw2o/Vz08cTSIHXlNGt4YsJk4TGQq6sWuvdc/nYDxU8gOuk+VJ2HQBMssg1e
Oe1nbJgS08HChqFZNhjns33sZ226amqMpC2Fa9AJkB/+syatt4ae+EglF9vuyaygRbEkZJ5kJgUX
5QyS2+ayhid2V3EBu+c0PvUMs1Q73Tfwzgea6HetSVns788asBZI8rl78xCf0+Y+we8i6oPhMw9Y
VRbGdsPCG0/9+Z+I1NF0VuTSspQM9MaBDMxGzLctHefef5pDSRrxnhfm5SmwyVI68x1GZ4GS9J9J
fgIVNLtAt4peJfa6E1PGqfIsBoPAudjQh8GzrDfkkZdRWVXjzUOfBrcbo/L2OZTn/Gdd2FYfRB/X
8C+GKCbG940rsYTo+8gHnQvr8SXrbuxqGwCz5UjG1Fly5ZwaplYdiIlNxLyqYg/AGRT3p3JZNI8h
/86lV2oJ0CmskI36VexmSo8tyfLZLz7VRPwyJuTIapqMd0Ytunk4lEZ5js+u4XvCHCs9maPtZiTw
Y5+Va24VC+GGBPoNjRxgkKyWZipdb8I2N1KqhQjcFtX6C3jNlp+qJfV35O33tp7PQCFyvPr17G4n
mPoC3dd40GqeVXbNbNeuf5hn6xVA23pnNMKWva02HK/S3xdZIGgErBiBInLNLuDKwU19LdG+2+AI
bq/S/b8J3lZ1xOmaHiHO3Q9RHMvILTC8gkO9yo0kSOJAKNnLuQMfqNH5AxXVioNyzgCO1Iu6U8U4
+0Z5Qwql36FzhA2zeIOD0qaKiCcOtLdQQwuNjc7fSvr+KqWm4AQ9hQKCSO0mnivKGQroFaNa4H4F
LYDxS9Bw136Gb2PGLN5iIFfSi48NhDeqwfhE/Cii6CDuqIe/cX8zyf+ICUjEejqwTWKb0iuuRJmc
FDOfbOpTEz5gWijsgE6SyF6PYXFysXfUrOFwVNRVvD9QAeKs4+cS1t4rMjamoNUBSqkHIy/+nspf
8kjR96oDkVTNY7Vs+ad1qO/hftokd6gcVSYHkhgApLmQGAkULoELTcf9XSZ2KwrnQPMthhbkPKjm
8/Lr6Nku3ziUTYBmhxyFUgk73SnRw90KOZVF2TIfWQaYm7Zx7KALusvtbg6riYC22CoreQ/PDVup
3Q6HeiCjXfSAaguXxbESEZbwvJneGrQl8rS47HymEUlldU+b/7uegq5P15PXIrV3aPyqFkiqvGr6
ixTNQFe5MF2LhV8V1JmcbJHVK3uqYKO+j96IrtpxY5zmAAiEN+fLX1zUSLqtZnPXj0mXeXZe1K89
8uQRdljaqtDHTjXMzl04cv6bhDOzVgnXP/QyXsglCiYWtzaiv01/bFsVrQSc7McUwV1aKCeJn8dU
FZlcaXN1jh190hLBhc4I3UADfbQiy0EHg8pwE4qyCRXLonc1G1CZojCUyRUnwRzjZ1yw1zvw+U/4
QTZG3+WdMy73lkJj3uvxcxri+UAAf0/3n3/OIAYta1zy+zVCyQY04mbdjjpVPxm1DV5QZFIoVKRI
yGLjfXrk5NxAgKf1Qg+VZLyUZD0qxLbaniFuw6CsubKQvGvLLUI0h1ogd4Ml5AMWxo+jTeTfJAY4
+iyeP3At7xf98/7Fm39pDEfJgUvhZyp9HOsnNdbJV+IKQjXBKah4FG13ajNGDHrUz6Y+WyfXRjCq
uSDz76RV2IoGqwnJEmY/a8TxoWeOECDbJGwqauC8xB+iWh4/2u2CEGVBY/CFMwNvLSRgtfey/qBq
GPUHb+KCMntDpSfN1OawPujGQZ90d6QKLJ+6ENl9bbqMhDdfIrzV3bEkKRg+rhEBEB0x4KKmJ2K9
89tKuwpctrJAoNivWlJwdPisrUMojtim+JHt+BlXFpvdQJ2ylnO+pgVXSaW5Up/nGya0xNIQCEl5
5C9Yq3EA3/5IDZrCMTxgajzapGa5T2PoYFYCt0pfH7ME5qmeBptxLojnnLJfinkr4eyjHfECF3CE
PDOl/B7a3pVYlVUkq2QQOSCNsHAjOxF0sfo5zmoZiBqpaO/Ke7vlNqkIiE9wao7Td4lckCMTOSgJ
B+sZ840L8cfwWzwx6dVV2AMlPjlZuqJoNLaHc+hz0UgGNm6cw3KWgLjkUZYBOUi04Er1D417tnoi
VBcgbxKIyqv35LE4PPcAQPji3j797Nvk1dM6ZGmSzcq7wcIGUDtE6a2Dv9gqxoE7yFkyng3D1a2F
Onj9uCFBd/4hixHqgUiJ1x9hsVLJShdZfJQOx7q1NUvijfid67Clmz2MZkfQU4J6KH80tlfm+XNT
jDwe4BaAZ4N8uriCXhmAf8w4eAzSU2PVcIXFE2GZnkS3NO6DxhUWPRCnVtDqRu90kIu2xCRdRrE2
pZvnlh3GoMSoP5St3BxBsrO5jri594cNoF6xyxkFG9ywLhMdxCGASWuk4MiIA1BHS7CHjUae7z1z
8zPdYbeIB4Mwh8sS1dEnvK9yo3JwI8oAcEKqug6QGby0LROmQ/mwBCgEh5fxAXd5xBzOBFZMZAKu
WLGLOApFHGFpIDrDs7ZIU4w+wgYdBzzLRjiL8NxWnLco7d8UwlZOtx8yULmcUxlwTn4yu1nNl0vC
mmdnaOQcB1CdVkSnR2IwYZgLQSJRglTYZcilG0ybAmxvjWZkUD4eAJwd6oYScQpYRswFb/orSTgi
ZPoXokIVSxz26RLDB6lRXaeoTKk3hxsqNcqNkAiaJ/cZvedc8eOg4Tb1qCbq6phiB03xBK3V6mlj
rKoTQW/5KbpMn4RGXFdnXWQUtTnOmN8trRgMGdjIN8tSLuPZ0Y1DQdSe9MZkX8fZ5MpNCDQozDDA
r8K7Y6UQrer+xObZEy68uby33Ichu+Eyx73QZW6cchKvpIpW/IU0REzYVnPHNgfb8e/D+Ygg/moK
j/ubN6ojCwogGkQkaRxFoDecLHNjtysdUIytwd4KGRbuSQ0Ow1iPqqR6fiyYFNW8ZQCDVzXAT97L
gX1uF4iQ88vou4mm3f5itI1hPodqeL3Dw4SxZXqtoLElsmtxXEOqsxKbZFvVCJzm9v8exx6P9l78
96XceQjW4is8s9eB7wfFf1zfju/9kom6roe+0x8dUAx5c2zN3BmSRdvvfEl2hPPY44E58w8kmgPk
tdL1wY/cGm3emt+BQsgGr1zdwLwWrx8D0JjHTxCY2EUnk0bjWcr9RA7ub3oqbWQZ1OTK1LdpYNRE
KCT63vP5XCFai+GaiXPf6JGxMjdgfUkD0WwtcCYV6rFCXhE6WfDS2NV/eOKUKHuwpIiwU+iph5Ke
Tl24lnnhfwujtIXSzH7rePxvyT1Hi6ngzbp0t13h5jzcfHmq+LFs8IyNcZEjIew3WJqN+h3T9uvi
/6Aqbm9uhkDZBUfKm1huEJkym46TzQjmythcSc2yeyT4y+nsy0wWaoGf9gg7sCN+IcFCRyPMixfW
QUOEbCXgPXzPLkp4L02LVlAxhBYtvGCAHxGAhMZemBujlAdtu8bnOuUz7m8WTG0T+7YuRT54vVZ7
qUeHStjy0WqT3UiPkyikdKaoH1QFVg4xeiVTtW7yyZQXxUymVNm3ITjuFKvkUfLYcw19UZY28pUu
3hpJhIWgMaZP0ooEoedHGx4DXHFya4gVlQN+okbXR7kLtewodho3rIzuHmhxX3XWsXW2KoSui4zz
4TBLFtf211XvEJvr/cTEyMJBWkWl81O8OmIjzcm8r1jVeQcOU9nlx5aDzErorVsoOgJZWYUI1dlH
PbAeJMssx/emoZrwnoZ8t87AHrRHced0lgY1MwI8/ZDQyve3nI7JnrKSL695B6ZPwp/EKZ98wxEt
RaWYZBYk0FRqRhF6TELWeGk/QVEH/eAmJD2V33P0DGzPC0t5ZCBrT9f3E7UtNTRVdTlLlPXDu1DB
rpqU4Eo14h35KAdEDd++ieNxelza/J4rW03bz6JRyefwtM8QcloZcXGt/cv2975SJw9gYtGL1t59
tiMfP7D09oygkWn4gUnJ6qExvooM2o5ueAa4bMaaOiqvhAMMfuQaK9pqkp6dZrEnBl5sUrjlp94Y
W3l26o4VeHUTq9Xaj7mEQd9hVHaRv7CZwMk+3Fo8KnHriuOMVUI4yiSW5YiFK8BCy0bom+hqxp6M
Y8AGMPRc+n2EDak5le/ocnAffFbZhIvoUMETPj2NTs4cxN3pj94PRtampS7QuLpUTDdLh4yaPSBC
rWQyFjSEB1N8QDDYuoc0PVa3Q5p/hJxyPWFq++d5NgxYWuzl/5BeLEFFG5I1iIxJv6Wo+/GYn9qL
5+Vr2pOpVYXsZrRnYCB7ekPO9GyzOmTynDioeIjaN4+FRd/pZwu9c6GYTVBBOW8s7op1jK35hikJ
1rAa0LJqsqk1vidI12qY3vOfL3/rZpBqY/3zVODMtrXb0L8NrYdpZgu/BfLLlzE9eYJpdt4TPfcW
0prWNqfJ4Xs3LtLdr5Si/l4fNuYVcaYXQkLdTJxbI3HOMnxLzbmt7A0NHYmtS7Buux+ScrNww/Pz
GLcIvZ6Wxx+ofZHzJVoVWD3i2VlCmyVVZwOxUgs80CtMPWh0A54ldnTsXY+hsHSgCz2cwEPwRupy
1eQzVklDgc0hoqHl/5Iv3IFCaKeiVqmtFb2+aS1s9P3DGyj/64JEuh3KHlGW4MLbuzk15O3cztci
95/boWP2UhGX3Ir+9NSOSKkBaoO3NPy/E3XXXidSjAYq0z7dGfrQy+r1eSdkYAlzV80pOmMK+u/H
A9vVbq6trfje0p4+KlorXLhkBaW1Fwz8BLa2702X0HWpf6EitX2qZckMsq65PNh6POLrNfYYaE2b
GYbHCpWKnmkJ+7MQTeCn9wux0ATC1YoDZMo7nP6GUPdQ8c/tveOpI65TiKAUI9CrS6VHl9fmWwIL
R5qZsU7PYdm8gaGloee+zXWKUOskGAb08d6Zk7y6WJS7jqworqyQuT/CHIqQeUbGiTk26NhktHKZ
bQU0EPtAB1JMF7hW1C+6RZQY7Z/wiTsaAZZlxqd2COz04D7ZsrBi9389L1vwZ+2JZa3ntG34cWIZ
gqA7iiKFobK90g2Ce4tXJKeCs9GritWwuMFsZzLIZblQYjfRdE2LEoAXz53hs6Uzel8nsf4jhEHh
PhXva/oPVYAZeTa+/l5QeWVzLLdM90eCPL7QxLJvMqwgB65/xy+GnbBxBoURpYY/EcfgIxs61XFh
eeNPBcNNAqRHAXSG1UjmMal5VsNawxehfB855heR14XIEUHcAiUA/Btq+dG1s2AM7XstHEjYf4Yr
pSZkKpm9etWrl1WZactgwYwiy/b/W+2kgLZ4LgE1NaS8fACjp0L5s16cFqx+BeOEUsP7LDc5t34J
8crLn7woK+xLGjYfwYiVJmgoeH7mW8Z0lNefAy/U95W+gn3wLDfpz01X1ig73CF9eEqevzToQE6A
PFc6xZM5LAXS6EbduOqbmDHkt1aZR6R6xExdy0itckk9Dm1a6/B6dcXU8LDjkjJTrAnZ+gkXLBDw
EW2b8skicO4OveH/f0nRlDdHRHu4LWzjOWSovinHsI5IiC7tVVHJbcsT7bxSkAvZgO50iabsmBCT
KCyqY1S24eYtomRBeGvwk9+GDo/JLn61gYPGSASau8M65sSbbzpgBtXZbS1r6LTLV4fnPTKRTCFW
lbTW7ghL7z6EQG1GAopFiR4KyaTPBLo2Hk7w9al1qImafcBv0abOSBudhg/RU+lkUFr0z6ln8hnt
rr8YnxxU1y6t6y1YAXqmRJJ6b9Vip8nSl7tWo7x1FQ3MmBAEmhXOOBUDZdAXMwYxAzswd9MjyPGH
WtMFL19ulgX/gc45yL+7lqk1qaHcTR0gYPJmW8PXMS9lnXaIeFZpuvqdsIU1Myr43k/9gLXDrV9+
Wx/nQTwap4NzTzYLKUcZnQcy7cHFUezA0R5LM/hp1kQcqDTFrCaNQwlk0TEagkGa55znj+vD7a6Z
mrhVdKdDIasChLhfhdOZzinIT7C6/8fDOsGYDpCbC1mZXQDrAYFUWhH0/z6zO54gyvY9spYT8p2i
bLlLYqVokFAnP3y6KZKefmzi256kzTEG7SSjH42pZpeGwPNDLD79fsE7qz4n48pk+Cyhc++4VCSR
6w93MVZH1olI30UqUKJTX/vItgSQ0Q1eAD904VZshY8yXO94uP27wdcd66u9zr8+8WNkQbYJl/1T
n7YJMZHry2YFqwoZneyCOwAEzKdfZ6It6bxftFOfe5nzySICATKqn3hN6kICwqsJVjXpzs1pfFAU
p5Z/bAFaIx0NcinwiwRbws/kvHvWM79cEj+w7VVuBVKr6mxVJO0yrv6k6N/79IaJCsjX8bYPX+oB
7RnmAMPC1N91PopojSKoUErIiVPKEWv+IzDgg2PFSb2lhSSUCaQprHJhpA6nyJJUum9D2NFFyK80
147n9yDi4trzQxuw7U6Ao1L1yyhOP9wBQs1lJTqc1muV28K/NPCQW5m56no9oMNuuDv9lW8a+yRY
0JgYjNWN1n8F2NM+wIPVuAA5SQCwpPvjFa48ssDsRHvBdmnskPJMxU4jEdFkpJida+jiIgAv+fc9
w4p8ZSWNVUplI/5Ryvom9JfkE5PJa9y0Y/jnkWQhjcNGztSALT9gmk4wXKSGNmsCGhlyqJrZyv6T
PprTfY3If1T5Nwid1re1kHEMAA051k4LVcBw2ahpwiUfDs6eHzQQKC9tgV/v6Brb3/uksgEfQCM/
2c60xneU/k86R8lKHtu4Ati4COSPCRvCxmR7Joy9cPohW0gggflMVSAUcn3toEK9yKJcLI4xNm5Z
ZUCEtoMUA4ZWflLx4iYAvjll8qDhGiXhD+zXzpj0qB2cbMqyIfS7yAIHMT5hahypIbkBCo7pOSyL
RqqP9ChzZ3Unk3114u4ll3nebIKjX+YswkKHatFbDQmpMxVgsmIGzWfNNMkrsCJKORtV6BvcXKGY
vdZqwklkSOXgGNeqvfUGb36jmNyuTB5Q6Uq9ssiOeRpNHxrbWG6sv9QxhV/rsC6z6/lhEUQBH0a+
OzlGuN3xkMhYOx+9mc0A/CoJ1JOvWbb309u3HO8CHCGS/+LZh6Jr5NaH+dsesXSBQ0ZYDNPBe873
Y3Yja/wuCQmP8lyJzhBkaSJ90SSZiHqnwmRtOPQS59WhVTApbssMKNaRGiXr+OQ5WzjRxFtloPXK
cxMxIC43qYkHZzMZ4Tvwtu0N/4qsSPZM6rB11EOE5mKp2dCoqnWrbSVqyKbhuiB/HQCpGwyILOgZ
iPjEx6wfWdxiqFLJ3/z6uxMSjL1T+NlUUiPYsDKqa9QmgkwRdHphN4e/tXwxgYrgyVun3CEKsUI0
I7wC+3Cq3aCVDReCQSsgcQeyCzkP4qoKdL3VPqf3B0Sfi7ZAtlG0jjqzkU2xeW2FXVo0ENW5STbS
r50ulgqD9jHb5+KJBQxDe0qey6Wg0OzVYdnjvTrTTlZokrIciVOqMQIjkx9DFX5WdBjaN5vTSOik
hQmf1IRgJkKkJnbORIsGgfrsakd9CmmqfXO00ATV8XYelQ4pelL6xrvqzu66Afrlt7RMmitLc4zj
WqigmY7FkFgmF3MHaijV7iq/i5N3t0FUcf4qOc0Vb4B6TU5QuG4I1JFHH+U/Y5m9m89V/PRApg5r
v1wzt+yyA6MMRTystCBRBq69YhjI6iBvbE+0iaFk9ZKF1AaNWBg+v+Srks2bFI25UHG/MytbpWxx
Ffcc98zPIJyZzGXvmoLy+A5Bu1qWC2AYd/N9Kyxo1qBGjT89G0Fi/B1FCraueB7lTxHR8DNLR/6+
MEIPm5GSpeTjHGDXKlHI1G+NrCj9luF4ahUeJ5jRQkBmh5spXIkETZjsFqLiOYKH4p80VhP+g59C
c/ezlL7PxU0yg8A9eOmeC7SSjesqNQTuDdKtVNWqOmiH9ZLSO7XXzYhgZp4wpaP/P9G1gCVrn5eY
+tjV1EuCdxn1YAEzp8YlzosRgj+n4fzzTqKV6ugcTcQ58mjQ/SY2KG1BE8cns30uiIDuPGnwq/De
4BTdzpODVPw50lrAeoXSq74SMUwM6vaOv4lL2clr19ViL7aTft1bMUziMyU00YEMc4FGTBU3QrZq
Xz9nITn6UHlBy454ta+qj54Q7fSwcXyCNWTJXTn8YyYYm7GKepXiJexgTahWr26eTiBQiGBjfP5X
7m+91qBzhkfilj+uE1H/agm4d02H6U+lH5KNrHuZKS9ZsUadT8fZte0fk1lW6DlVZVWEoaiLwCGU
aJE4ZfXdMXw0Dx6xNIaW3sy7WpJqIpShFqSHIj+PUC/dB4h8IUR3NuIM9Zb+qhfBow3gxaeEEGXt
xY8ekntW3mA3HQmAKsjfgqrnNHkGWYpIv5EPgeUMdZQqysnMptBk/Cd2Cpz40FY/WwZ1vyQQElov
hxWn2W3yRzUWtiL6iDFMyFmClSu6j476Qlf7/4CgpVNvNZTybN89fHJIe870CYGoZRUZx7vB4fwi
hwjl0FJ0Ivgm4knB8nIZ+FsVsv2RMlomcEogAJgsYtsTKyo9dP9NfsP3zrqQwyaTGKs/a9dTHxgQ
V7/Dl8KS7F9NaVz+tjIUWxoKL7W/iQedxu66KhyIMKsiFs4azT1NR8TJ1RwTPCiYS+wY8jRCbJyo
b7x+aE1lBsUVJkyTtJG+8zc3DfoJdtmgHAO8jA8W1oBz45LNZ5pRrTuYOExuL51V4nkMyJOcUPA8
kVKwqlulMPgu1kKUfsYNVuCaVbeVQC7xndTOp218YA+0B7dqBnfEuMFgSVSngt0q6O0vIomJIkHG
hCee/aFLdXd9PsMRaQJv0MoANQF5HCgR76NUv9iHNHLpwMkFGk2w4g77zInYzM8WciXkSFFU2pg0
75Gro+cMZsH+RCMch7mlE4crgtQxZsBIYdGGRIUH80nkSWubc940IQr0kFQqvGLiscyG5pAi7BIa
BtFrrmiDGo4YIpnHyRTmz4l8WNwtn+iws4ffdTGe0Rjf5Uk0VwRqifr+dTp0hxDk4IQz+aALTZfh
GRMjD2d8eZ5VNZ5LZuJyMhRZpLJgUMzvhlZbEohWvw8usp1ALNbrZkuloyGX5Pr7CXtoNriI+V1W
R1NJoNFkNv2P8JUJTue/oe/jD305eKUYLyIsRBQl9mHydo9GJxe7iKomsG2V9x7ZPjqnIxdvmCwn
IhiWgOW3LI0C6XOLXLKI/pGy6rpRzCZ9ZMfDCADY+kRZcBvxtq7aqZF9Zr2yO+bpw/26Zu7P4Kyo
4O3jAG2qaOUHntD9xHFWn5qhd0QTk7qhKVP/pLQ3lCE6t7KNkhu6a2x8dOQGMGvG6oezYvY9IqoZ
/MOE8r4/MqP7Hb8hUZ0CrKbyza5PCt+yrI5p9CV/e/M5l7okANjoWjw4UXqg77uC084CjOA+FFWm
HG8NlvD05PITJAUYxz8OOVDiMScw68BuwlA7/H30qrS7zSEfgaERi/jAY2I1ztxFqOK0pgmZvX5r
puKkkEXUzlz4DSd5Zvt7XA4ODMU8VpbUZn3PyiVsMDJzVplcip9sATSqFH+FJ7bBzOVaai4nNYuo
6qfc/MTFz+cC91LzYJjPAKPGP9iEeLHG/Z1ByJCvYdv+sp30oOt7KwOfi31vZHqwsXHv59naZqmA
rEGyNZmq1cBGf4FPmNQFy/IW8cwv8yRIC9opRU0kEmAlwOp7j8ixvUT94aH2xY3ofD5JqejcqlYC
wclhwG3JpHNOOjAtutXDWYwVk/5fPxD4BC/4E2z2zsAGYyAt+WPrhHRHdrnrKdAvak5MBJ8had5R
PPiuKQkkaQYHYUUA+J9820oa+1/Vg2wI3RIQMdP2t8Ygu4Cak2Sj1Faxd+Towva22v4Ae/j6K3zi
3Xz6z9ba2fzHF+2IQGPTbOKyBvQVt5c36emd5PltE2FWw82PfmHavWG9yhWiuOhzOZjQjlBixxfb
jLxtWfC2FL7iuZ87GspVO04Fe9BwKDKR//6MiKfBUUishSKvrUm1gRGCfdvhMxav3ix+38WRjmqk
v6nNbjgTNaD5TJcTP4qUrGDFr6WhlGRj2IPHXGu+TT1pRRUfY9wPsJwpPCnM6VfxMGEm3IHdXCAI
uD0Pa5xb1xuQnraDL0mpwOY281pYBWsrdILdjNGOdcDCyrNqmppVV/yUffz9cQX4MuUOAdJqLSpF
jEX+20TvMYoCYpxPCtqLKB1xAYjbyflB7GjVWkkyMwrww0F1IYsRpU5fQ9Q6z/yDaxL5ejmRWYBI
JaBTT996JrlcHTHWqqiREFm99F+Ad2wj4pJGUpQjhkjZzHJfEu5NK2pyMorOAXWieDtEIItRqliV
0jL1z+RBDpW4LNNnivf3mGEhB0GPEl1ay2YNiPw8Jh592uv8+cXUEakIAfHKE5AsJetfpf4Y9Dcu
OXSVtmYR+kE6sIl1icluGA5azkY2Gy+tSh5VKQs0LMzD+Q64gAW7QtzvExMSZJcNfOZcZO9zecNZ
w0/tuY2nRWL3NRdLDSngbHSe8B2oAeum7lYIjcT5d/2zt6ltPyeaNS0vFg3ceTuMg6dD5vhs/2S2
sewAycECwkWXkEvcPAylV9u6o5kukSFHZEdiLn3NxSWOqz23gSeCZlLiFdGTTGBo0GCGauZ2sxAk
/WGqy+fFhTBChM/lZJkgQmNr5Zy2kU+dV74yVR2H95k1U8u5Yp+FADuQUFIh+qe82naKfxT3nPvU
C28/V61pVjYbWSlcVobLlzrSr/W8k9mkw/mzcEnQqq5IwKxbyZtXSZ3wqwAhLLk7PwaMVCdkZdeI
ng/Oiy6YsusbRjP5S1KBY1rjVU2UAP/kN36YCNjQ2zrY/6c/bCRSigRC0LaVUast4L+UE5rgo/2M
5wv8qiVEpoCr6npOLc5Y1RSKqR4xdKR5kulu328nayJquNmbWZGbd6sLnbZ0QiLRkZ/tYHH7NZl8
92WqQMKQsnqEHA7rMJU2Dz9uY8qURaLCn4ueNo2cLsLqBhyk2jSPS2iCrVTExvpzSb+G/RTkhB1n
CgW0I9A34ut3f1Z0Nbs4QGH/XEAW+TLdyXt7UdSi/glygdSKQ62Vd6jPC7K2lLEQ9RY+sE961HSM
5u7P+u4MYJ6qUYBrXLSO84gBRNO4rxlilqPcX172DDJd5iRaO7IpMpRjD+jhqINP0qtDd1QDVOOB
qQ6e6nRs3qJ7/lfa43ypvWddj1DzIChDsmq685Ya01M+LtOWNCMJsYCqbnceTNg0si29cS/QB++O
fGF3oRCQTh+/41kwilSdRbTwJwUjtRxmd1isorEU3MeDA46T9gzMZNytM21J8jNfm26ZRTn5JsbA
5MONDKm5cWuQMljGV23DpO2l1E7/PzLfwWaNWatWu9DooH6V1om+X/IXD790J8hOpEpt0qyuFE0i
xgWdA4j2EnJOPZHRS/MRnAbDsyOngs4hXlnGmlDDugSmciM980EfGl+hPIFRCBxYLcG1AXOs3JDt
GEHKPz3o6Zts2FDkmCNhyJOwfUWt7npTHtbCZEzxYiQQoUCrpEt4d31yvgmFQ98Nt2sgW4BU32bb
Rb/RR+cfLLFg51zFCucdv7YU5GuF/s66tNUxsNBA3uqJp2kbQmj0uAj4z9W4E+XED9Vs6eihW+VH
vRKnbdZpMKgVarghOv+R6rtdyPvz8miQowJMcOCSy3f5uSh3Bqkjt4rfSILyESyR1DhVtli/sJpp
YQZZr/1QaQiqVFYi+9vsctmGLIx4kPyol7BNduOGTZ1qBX8ZahJuZQLVyAxTGRQjilhNa0wO3sYw
+YfUQRvF4FjF8VdVm6xBMz8GGW/nXtxjvC+JwHs3UeMbnNItfwVL17h49XNMul0R4Z+g+JLLx5/M
Br6N6Tj1zWFuDBVcvZVpCAxlv6JH4twqZHAzKJzUnaQRjNYiXIhobFfO43fmUUkN29/FBZ8K6u75
63QHEi2hcTIT3QIfTUu3WMjPFYTf2bwWDLpRKOI69IgwBipOymaix+jjuho43DzvsVtEbVCrLnLO
2kMipLsMddu3AnH4i3xbaPHIoT6Kx3EZUw6ivf+1igZ4TwZvwJlqWr4B4GRSkkT6UeRLTT5TRDf8
+hg8uk6BBjSCYVjNxazRRrbyc4bbDpW2x+XUOBx+nQWow2SbWebYHa+DCr8/MI+NMytMA30qZ71r
Xu94xv1H2Isk7aSx9v0sSyC4bltRrXROQdcyXQrD3JFGwS2OKzKMoa1k/FDQnCYceSDJ1GmfNMyw
EUCPBSyvWeI91gHN6jHuI/wHR382yybF/ter68kCYLxV0hxou6EOB685FNITvH2bhs4Kx83g+ANg
3OnDV/+hoDGKMJoDosZltFIMD6T+PTkmmLWB4YwL4XOdJEAHk/NqitV2O3dGkNirqIYs5qVNT7hD
fYvXilrULI9TnXITrl9yP6tPmDW4491IsiyL9QR0uo90OXRaDqOYEhNlBUs+FtadAf15ocGodTQ+
uWhRWOhuWUgxvp4Z3SXB9BqMEZa2ea2ZQzVQnYDVU1gIIKSTT+L7WXeuBqJnG1X96EtxYPN5fwJF
tKoBprMiZXJiZ/cnMH9SJ371hhFaCwIjpeNGoY0tAlxt+wtFVIofFzLpN4PoXyf8mhwY384Em2Kv
SlCow4MN56zKFENJSLBt/1ZWw+a50aZABQ/b62rxlhAMDvvSxuZnSCF3lyYbZenCaY5wT8uxxRwF
9Ay1g0bdGSxSLT/AwaoPeZAK03qWkFr6j3fGXNEethT9Bvqt9hppmYYvsVX4hVjCrfvFylRSnAv7
UKEa6Y7fN8pD9Qh8w+q5Ave1r88QL3qw2iwEsUVgTgqeCzJO5rDhZGFIg7loNob6aYc9DiRUtka6
U7b88KaEMsPwkox/sC+fqj1f7aOeSUHOQwfWzp1rDkdfLU86X+Z5NmYGVdUVDnBFrEkJPgXQ8zDn
A8V6ydTehqi5la3uupdWj1omum7JVTsI4dLPer5qEI+CJjQWmltaa6N9C7qEhyQKWPhnEEC8SWvp
izidcdiX2Px/KqvnnW4d/voo84cKxP1DBt5qnm1sD0q4m+YEjKNxxFsM4NL2aczxxw01flOToite
rT5I/bv9+1PyP02QlsIE4je7PoQ9BtZoTZMv+liK6Hswf5mXj0EZSx89xowOkmu158nnA1tz9NCG
Cr2J2l78KJtDehRDxmWB9Ymp6x0+DcKYNl2PkTsyXO1egUW7fX5uAr99aLHe8bEqW5Ghh6PWcNUS
Iwsqj7nTDCrLUbbQdARoiZAiVKG+VkEuMHtTVq/UUIPgXOYe5YMGiqCgFiU1CVK2gsHp3JwNqnAZ
OP/GIKnw9FEbySkH2Ae02fQFfXDIllUHbhqdFwjhDOeRX+qt4RbE1X93HLLx2By0FlCtp7kiG4H+
C5dtkRql8psXedWsisgSFr2KqkakzFTq15G2dtbf5dcmWxoOKPLwwoVcXTn6Md97tM7K5SiQjIFM
+IDwAaUe03I4/APcXI/1zYpCuA1TmoZfwcagXW80wJW3xXNIe76OQGRWCmRa0jcFwWJrkDeyuh16
+1nmC98AFTdepOTroTF2XwYP74Fn3C9ChVb+625y0ppdcPQ3H8EaDUhmJiMBE+PzBuPr4qXRYNCM
NZ00ctpxqhP08677xutEko/r9cOguG9BrK8kmZmEerFdM9xOYuF1T4KL0UxGex53RDLgCvscv23U
rDlB6bzHT1sFFPZH4pMZTuyE1KhoPVzbCz9iKCRu1Wu1zOGvNSIcFfW5gu8Z6YMubZmvCJXhq/i1
oMwvB52J1H1zetEM2vPIci47twgf8ASPV/BjG1XlwtOj73Z/bMdMkmTS04ygPQIkGXP+h31Qv55e
Vy8BK89AJghlgvCWj9+ai1sBwbjnClJRm/6k33gtzO3YIT68IjyL7B4DQvhOwuaY/XU7iaIlgsMq
+CfT0vFoXNv/I5+CdlbDGB2iGYQNd/Vn0andOnuajXbHpqF7jZtR2yzCeyte+4aIUocWwtSXdAYE
9hH408fuUKbgPE/MOpV4JGCaVbGzUL+eUd1te9+G+a2gIRY8QJTFMcFoPTmqR747604V9uh+WmgL
OZdUHtzI707J1XP76j0oKdumZ4b2XFsYakvwieLz1A3L4lThvLRxD7oUYczQgzFxsI8bFYJS+MNe
wFb/Z+w63rKvBUKHwqFdrG2mk/nKZYjYpExl4BJWnYD1Rpt/1qrSWjtSVMOn2EjoCPnXYgDb60xp
6u9mHtvzDifzSKKzsH4IuJaC5TH/ONwFk34r4DOanpW/oQnwtHGTWSK3RnB3w+AlsckCKFuBeNtW
7Oiqh3zIWhdfKwVWglsByQUUOqtSWiCABnODy9H6/AsU95MTYAAP0BxzJDKH7YRETBVvVJI0DhR4
WjncqES98XACxY0asWNbGH5bZK6vw5PJ54ZbNnUNazIthwoVl7VhKmJRTh6To4g+W6fivSVCYEz9
WXBCZvbvoMf7iLh7prVDtTDVcPyzVm63nNkovH5x5R4OxU3WYGlsm31VaLYwBNcVedEws6GONgPy
w3SlEeZM7x+aUyW7zrSMfQBUEaJJBXW+BcktfF4OdKRxaCu/Tne/I/CCu12p9DBRkDlsIhkxozSy
8WQwKnk3Db1Cs0sFLzwYnbGR099tv7D503+1uAU0TxMEk7dLmR6UYt85X31ODJEC+Dh+hwW5VFtr
K75sauRY0Ip1FMRTeV0HcldHznuLLt03MqU4vdzcB3P7VzmQMEceo6rtRaAA7PJT71bA4Hm2tozi
vIxncsRSI1V88JSK5VGkK91+Nhmo9+B9qCGhS85WdFhGwHbxFg2Jv3jvypVAm9UXXG/fy1EbuUlY
qP4Ja9m2M9llxC84zWMSg1u0PiO7TW3geuCcI5scbsgwW7hfLRSebTCQnCuQrJ7qgINuPv6/9Mv/
eWlLnQ9Gjnr3SbjtXfUrwLw7G1SqeuP7Oq/i7QRPL+Y+tXPbVj3fyY2Y+DZq/B45lpCA3f0m0v5x
kuO8cW3I+Iy3V/Wk7qIJknrZR1YSZsGjrqImEmg9wdMqUc743K+8dYk9OQwXdm41q3JmrbKa/1te
n2mfA1KeR2HSuuAjAc3tjdAUzbfTF5AQArITN/p0XlnqGihwV1AyhSijEFl9xEOszn6dIHYnrzRJ
AaRgE4Aj0DREh6xW1TtfoXYNZqNxUuaowZPpWhSgzQF6aCSxmZVa4Ao4iZMSWxtMEtk3gR9tRH80
aVyD4IXRlQ0qqDB1z/peFJCLqvJ9TQPBFrGI/gP81O2sPsQlRKIEjpqCNi4AGgjY1CBHxs2K84Bv
80kz0mP8+CXwrHyF7UK7YVsM3ElYGQVnhYWvtIq2OfUu7hFE1R5uC1N1c1aU2j4T5kf2TF5fdnwT
Sumk39O8QfDCeBkUfn8powy01z9ApdI7bZJOPv9rBgkLbAEKpKGGAQozmGWn5Su25ohSsh49TeAf
ZV4UiH3LnUIyJHicx8bRoMOyTN8ARxpAOFfoiQ7O7UbKqZPoIwkZqWoeApyUpFiAmXBdEgZOI9Qj
CCjem6S/X5SURSjHDeifx+hNAAwQtiP42bWB79JOaYOsIYFuXFSLDf0vbWr75SR3/nFDZfQJg8r7
u6Vh5SeG3zMnT2IedCQYECiIJcZHeY3Lz3y9lK9GER4TEbn87q1+Hr3upNda7M/QoLxrURe8x1hS
Bus6eGzmXJg11V2yo7zCSlgO1CuO5cJkNMchUzMC1WXeqRRViPcMQ0td128qTBehvA94hWduOOn0
6i40Jp1/+Mqnz9Ijsgy21SdnX/V4C5IQUKrCqQdcjwiPfYVd7T1Jz/40WfQV+AQjN4awUiwCOYID
XwrUhAXHRCSQwc81Y4UqNiiUb+mXvDSOPptxerFiB33Djs46045npAgeoRScbfNbx3PYQ3Y+jofp
00h2U8TK4uV8eGQ+KQNFMnFT4aJL7WjW1AHiLJ47Y/AEsesrk+ZhGnaFocrSdnrH0Flhn5em0ARi
p+RFRcsr7nmrnF6V4jrAV2TAA9t923ldbC9gybp9T7fh0QkdeCmJiB8Qcq9X6Hqh8p3iCeT7/pWX
N2kS5AQsfaJvpnS/KkH0s0wIDTtVGY3VcaHrtPS87YnsBv42hqrzdKuUEmDkQg1XAlfi2WceHx42
Hl3k4yS91eL6QzuJIzBRb1j1Nlnzti7m+SXVJDhh5py4hTLqhkMPDvusTbh4AgzK3SQfRC9yLJo0
7xzCRJ6NDwvJDcomg4HnJ4JdSg4Io/fnWH480ko21TK2nVcE2c3HHWniIw6CS2KQNyuzuBpta7WD
7kmgFyg35q8MwVbKknJAHixAyVL4QHQ5CUCdlR/QGu/H8E+uXnEfRz1XaRwyoVfosORVGuhJ489/
y1mTymuuVRX6wuRXAaOCT/mudx86m6pjN6GWCN9go7+StZPqsyee91BcI8X0tiXdYA3L08SrHZ2L
olDxVeL+bQEo0fzRmqNrjZTnik3ML1u4QdZgbyNBa8ABi6r3e/VIpnJELvL7o7gzPFOOUJxSPGRF
HnmkGQ+ccsf9z0VPDSZ+3b2TqD/2uFRIbwHsvg+xuyBR77NrGXoNz8vkBQMVcN1XG0XbqupZlqI/
+5L8wnnNyyudszYWEXZfck8NF4ZJT7rqWQasMQ/NZrrz1FFUWeuWZmWhNUlXPDqT4IqBUmHU9Iea
Efdfy6aiYKo5dkgzv6hKFb56tmdcBqAtWcD+jC525eIcbIwq9iyrm22LzSsfvBbOmgkHC5XZlRNX
IKy7y5CgymNhYvEKdz6ACc5y0RqsRoZ/pxfOAnLPOFM9BCqd64JI7GyjSgZF3O6XTUcaHdfdHZhs
XtaJSVaYYdEuFsm78Fe+eyOlnPA7C01e8SS+Vu34gdOG5ZLWstJLB8hYFXVskRIRvO8ftjEilono
w4I0at5YXOYCLXVv1zUP7zxByw67R8NDQldFKgreStoi+0dicXaDmbaSt9UmINbpR6VNgFJFnw2K
EpsT0X4GppBL9ExBQcuEEP1fj/7qcO7l6AzaYZ+H92beuTXHQ9V8Tij2ZLO2Uz3oJsBool0iOtB4
5mLaOMQqJR9U+pculFdBfIf5bM7napXOJy2GpmlqRoCwjHY2o32fhAKeF7tX4EPbRvDDyqEh714j
hzv0JtBFgNAm2yjzaxNySoBQxWlPWlDBPP+sag1ZO0aJV0/soI/bOVQZ4P8T0l8uUnyoyMqPSh1n
aHhn3helPBUpi0OJkUh4FZPCQ7dsqyxrsmrIroccJNRUMc0XHE4cUDhg4btXhpRftdMQpko6ecao
OyMlL5KXNwPEq/eTIhdGzHZjFSN4BzCtM2+vWoiT5RCX+aPBFdyO8P3V6J3zclKcL/9w/ljeIK24
6ygVvjB6snHbp3i91UQbLafSCmgs3efLdYXOO3umwdOIICQqm6xqeYrT/7G2tu4N7vgkYBKXS+Ku
k6a9cUJhZD2twZsYT8m5lVT9yBJTgf3H5pr/nh3/XEoh2lUwRaTZAmp98PnTvBBYMx3o3Luo2ozb
5nRFPaUkVYM31eYWiwGxMdNnep30owj2yeooWjH8a/SaxyjZJBoWERgEqVP/D9rHt1zCihEc0Zrr
2/BNFBIwrAPufbcdUUw0U4k87qwfSpXldZ87eO/w8CgichfHTxoZQU8knAWhbc5j2x7mCLHThNz/
lEwUXfRzJZRWiOTjdpjn1rhmEOR+/UFQOkYLtfLXB533rgu0r60Lq8/PEvwUqxWiV3TZyIjfCaLN
/0BCvRvE9e3lJ0MZKq0kFo5U+zrf4PurvdJaQX+rFzvXznJ+tN6br6+ITVc88KJg9Swycae4Z5Wr
+CUpbEmDFNOMkumgSc/P1FcaF4MT9MvEO3+tdCA8p8qZE39SGDzHP+qHxYPWRUPK9Hkf2cS7xgMf
w3k4JFn0/TqfvLCPWAvbYX2PAy0k1LA6JAR0V6xE9uw/8++qXaBfatp8aqZNcQBFxzHjpQ6iS0JG
hNKgeRe7TTMKBpINMMsE2zemMHTJRiHnBCgZEopgIwch2KuOUgdZ5d8ERzYaJ3oX56xQxuFG/Gs/
7KRWWrkuex6MBZ0w+cu83/0zdHHo1+J8Aosysvq1t/AzCwu+H71dWlD6WZIL88mTb+stQUea5gvf
t6s1y4edaZjiWiZxJAvUZ0wZY/5m3wjh1dPvYhLjj/ISYBlg2y20Sc/Il7Yk9l4LFqqIgAwz2WjM
xdOGcRjQ2SItjT8t7eyZu6ofIFgHwSFIRGy0XJ/BYhHhg4YDKoF/r5VSN6prv9Cpg9+9yvLjo/ik
wJa8pLbBUg+Phnl2i5oHvl3Gwh9Xj0wDZky+tUqlXd6EeqxtrdcESJmjWHOwMvf6a6468vvwvkeH
hZDavDx3kWIMenCEM8tC0lcyUv0Nfp8113n0vOpg/VD8Cj9jSruGk2XFX4bkcybCZH569kL+YCsD
I1RVJ0XUnmBg7Nh7WchtAm8I+71uj4W5CtuhNYE+OmzY/0cksJmYebJtBH6vqnE/p52TzAiqNMsD
l2xxQF+kBJfP7fuxFSZiYuOreHGE4Drdx5sO94OsndkmSMknI0Fsl8G6cAcorhmtrzNVUs/nfiGM
igET3IcPGCsw1ZNgGA9WyIhp8D7JsD2hgmIj6JPmKaCeM53vnTjdxyhW/Q/kPLByUGaQW1EZR3hk
iUisgmfDnHPN+GarYyrDmIhHOSaJ5Ucs5JKZw+vPU39uXaDjda0VJEBZJfxXH14RJpHN0oDyknEc
Dk7kdajrVq/zF2O/0Fm90s4Udz7tEmX97sBsSTMbznimYjBRPMIUid1URm9ipVk3gRJjjQDK9duK
2K3ly/XLlwLAdMEP65FdF50lVyv6CtILXqw6P4xM6cX9TAQbUS5lNIYQmIvHPqQBJw3Q8wvkFVu1
vPToeI1YLS1U00rj1yh46tU8WXaZ3DSMbTJ5mceVy8qWjQGjcJGiJmW5FEbf9Btfaun8nr3Ao/uC
G+pqs/0DtfVmsVMi8/ZVMh6vajYJup/sZafcp42MsPf7hEtvBshd9QZ8nE86AEQ85cMaV55y+HG1
oP5S2X+7prXZcof5VEHMdBRiCYFIWUE9CLFahz8mrJLN0mxq5FJI1qcaXX01HDE7e2KLxzz0eOw4
1+qheo200n4m6OWbXcO9q0FxUjzx0BlE84XRGYQ5io0/rmBiJZEMgpdYJWGm5XvF9h+7EE2jG3Kf
c2rj1Fme0bO7w1e6hOeObFSLOil8GZ/OuEZGwJ4cio5V5AV5uzu5X3fzxfRabVaWNV5BBqfdXqnQ
2KHfnB0P2jXpOzX4/TqIz1Zr2oeiblsgfKqcLdYviBT7grNfSKi55sAy/c75m5kQEhrpeEOACMaA
274Uk6hrQyB8n5+q2MybG1wC6vwHOWX4K0az1dgoPouoqnZDOWZ/w/YE/JPbkH2hSttUSwY25CKn
poRb1SRIaZE/CJlmcZSJQM4rGHIED/D4NMfYR+lGgQsNFjfYj0vjGWooLPiWQVnbCfmRFYqmloB9
fdWAOIhuomtsEvQ3rhposQukyOpqCvyeSHhg2UFwcaZ6N3aKydj+nJc3JBQEcC2GCQde+K7wN1mY
PPHBkouiTX2xWUMbfLbN+UZ14ax6G9LTbJFkEWbGxnkaKOpepZ4jsKbUpVZdDjw3RuyM8XzOOaJu
VjnDy1/J8GTET1s/Wk/VvtTnb/LowU+5mvks+vD/dm4HMAEQ2+tWQWKOGt0WDw0e3Tb2NYYk0Ppg
S02aIzMFIk80k7ILZoXYwIlxS4Kl2xhUZ7VOmli6zY2kRKBqJABfaPfnnoPIkkyQSlYOh88lUCjG
WdFUXmuNdOWgHdT+ceaGFu+O2Yh6jl8tBYJtrrfATTsZMzbI+WhfpJvNDMKoNR3rvUB4fT2/rHpF
MpAiQskpNluQn1PvCN1h5GqeVdl2OpuH5spXM6hyT45GRW5C0/V/UlDtX9o8Qnjsu9yS1P+kdeS4
s42RNgwamtbd/Le/GMByAB1aPa7HPQ3koEEstNKLujWo0QbZO2Qd7HDkYn6g70KaWsYnNHDXUHvN
1vASp1ABbAOeDElrvw/VgDCuD+hWujgU8S2eQhkgaNhwhlwrQ9rufv7iEMUAxxjUp/6+39idQgA7
8wKPe3Lfvi8L4hSxj5TiNOBZbm3cYyYbl9Uy+mFo3Pwa+/Uo7ql1Qu7JwE+9IG/q+YP1AcrOxaCY
dRqWhfteJgYazev28JQPjYcV481gTW26rl9qEwSY2gQjr1fwZ5M7Ojv/83scGNZ0tos58M1QjekX
jrQDLqAx/sjGRWumnHqNeEe7div/IgQjf7Ug2ngrxImCpyG3g45u1ZLk+6iTXX2hoE/i20ITupZJ
Asv7h75jK4HCxTdTkbKHHuXNy2d6PDcs+ztN1fNnrx64GDXTfISth/b25VQv7TVbnNwpeJkUSGgv
hITACKINOzn1r+cBcfZHqGVOb8PsM3O3SL8vpSn7NssmFUrw58W+BSN9rPs8H7nb9gGwBpvnw45C
vvSev/C1tm9kNHPHkAPGxV/ZAkoFFlZKFdb1e4tD4y03pg8M6ytQO4oIfWAjPAyYKpHwCADBFQZL
go99Uom7wY7lVZ3FdvoZPIM2VAifHL0mtwscijlKK7OOIPjDy+UeQPCjJdjW4/DuAoJvEWopnWqP
2PzfHUuIx6m3n5nKBtOqhzaVOQIVi1mah+uhZUsY75CKLw4q50Y0T8UNWtxjUb4ogRb3kf6AGB/t
T1XaH9HQPPJISqns2SIy6OT9J088EZcoY7mWH1XIJp6/UWv3X13vCYSHKH5menCbs+BtO6hM17Rn
uDbRDqBMkVWggCbE9X1pDq2K0ooBF/nMG52fIjGkJY6PIeEi6mdT5PViFo8m6/AgEbduhvaeoZMN
8GIJcC7a1Y2THpALLzWgX0dL8iTlLvseKr8mT9FuJ9sMposcI6rgLAXIMMI24Ol07moN6LEw1drk
BlutU3N3euj6FO1+My8yziuuZhXSSWG2ppfKyREaZER5tdsIf/hpKB8B0o6AQ40h4IelBryrNQl7
Gw06Uje2uIWEJBjhFFAqR+j5UZY0cxkyS+1Cahnaexn0c861CK/UJDw+0PrdtmMGEoSSJgTMVgIV
1ck1J6J3PJSquFe4UcHdAHEzesnJyaRGbcHiFeJ4Nqh3YwATSDTzqH0moOcjRSxbRm8yV8J/L2R7
+Ke1MJVfsU9d5GR2c5KFE1katq607ZvCi8M6YJvQdSeTtR6kGljyr8QNxSxjBYw=
`protect end_protected
