`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
hojhJkFO02EwZo1gPjHK7Iq85rW5Wq4h7LffZUYaDlcFvW3fl7zJ644dO3vCni6UyJAsqHG9Nh11
2P5myDOMl9DR8qPtpEnHo3qtpn3nHkzkotlVNkLjKD6dhzYnTjwyyaRUg7p5uiwkIQmvQ8mIegbn
68AvV8bAoih5zyOtXUiHvfjDsF6nfYwvYrEqFx9cM43jTwsLEPhkEXbCnw0NQoJsQ0brrS9lJrZN
rw61rFxwyHAUoTj/W8ga3CVpM2hJuAo05jZ27I9Ht3tGaRrQW0stIopnkPMAmevi32Q96/l8ux2T
QRm04IU5fqDsqF5QFntQnLUXZPoAN5Say1Tpng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="+J3P3Pdw4irMeq8HGi1IFoJKaY4w2aWkHgdX/jxYHUA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77632)
`protect data_block
kLJ1jqimYJSe4fNdZwumysF1thTIyvDn2sY5ukGtpkJArS/mftGrK0P5f4QJtZxcOV0W5diCHXTF
3xE121LqRFPa0e8zhIjKjH3WDLoQZByTMLGSwNYWnQtctsZrNqMOtD4indXeSVN6VoTK0qn3lNwY
cPJB5ZhujyI4/hiPAyLH6bZcMuOEQPyVIbP/Zmj2Q/kFdFnDdaDEMMzy4qbvjz3Ooq057wKdAiz3
KvE3eze4wJ6y3//yrMeuCSd4AjmLGVlE5e0ygw1n/j9lQVAMpe8eLpupLtWW8SgeY+S6LwaeNW5B
2P8/3HF7A06G3pLdE/Y4BbjDueRlhZpaT2Sbbb5hwN/oGFw98wjem6QC8lCadiJoFmNCZ1pVlxeZ
x1O7o9svxvwhjOkdnvD+AIjtu9PD9nzwDARY8BgD2RyaEEOfSIYpz9t0arkFpHPVU7ei/JsH5rT1
cMzjZFzBN0qnW7k26E/NJ3E+UAS6E8jLY2+WiV2Gqt5vXJSlqa6VAJjvMwEMewD2rMx1QqgP5PnT
a2Ecg/SbK4VXgGZDuSZZ+uRuDTItATBf/T1ksWKTj6+hFeY0jaCIFNKVDaKu7kShv7aZQ6FHHKuV
i95WKETrIBEH4szjQx3t6RaQKNmjtgq/AkAF/TATFmlAEF3HHJEYkGxMwzQSPtlc2iEPRqfbjQ/F
6yfcX7rvZnKBapmNFoCqKqihLDfTk6dYi0kiAEy96X1O/Q4Xgrb3Yx1qLWcsYiiTfc7/JhmvGqEO
qt8HZvubdUer+KMD08WguVyn6Uv+z3+23/jBOH++Be5EbG2TceJ4MVy5eqf/yF8Wt28CFHE+6ukG
dBhFmtmn1j8O6EBg4RdE2JoH5rXzJqfDGuG1lwS196jXKzvEy6X29UTUV+0+0JqBoxJP48ENLn3z
O8mhjapFo9s3We41B2wU5YxdvBE2gbVzgWEsP6kVXkRi9iCqBPco9bTYcn+oFXoL514WDhYDtyRi
pEcU1kc1OYFVEQp6Dq9IE6jAn7zICAMa8h/Bqeuh7XRNUuweC2sZTdG7Q+BqG+n+6mNXHn6gKO6m
ZLTRxrTERZB1+AOCQFR67nphur91kHz0bMqrFz0eFz75K0sJhkSTNWrPFU6UGr//pagNv2Q2qgMY
rIpqrakbisNHmzfWVHHQplSW3UVGHn13+tLVdvz/NRo1B7Hr2HMTl+QGgy5l989FyJQa4qauNwFw
3o49irBprOeu2JQ4ZFVpf2EyXHDuOekDkr+zg8nCZNOEDkbnMgsKOMQ9MmYan0cQx+5Gx6Ht3GZu
CxEHhS9wZzUHTr4npIuUBdVzDo6K7npR9Gp3VlhMKBvel+67VBzoefBXP8mpeUmQOqTkHYM8wBa1
g4eSxQSQ03ASjq4pH3Y9h0C2usZ2QtVs23eZsDnovidceAimyQvVOn8tF48VdGjv4r52rZ9CTBqN
8aTTPjF4EWVMEve+NqSKSEMzpNRJ85XBvBWj6poF9Ws4z2XhFtlrrVMJYQu+ErrMAlbX9jEVFYR4
+LXjmM3h7zh0RS3U0e7NenehQJFOWsyDPazp0CG9d8DvLg7WsbL4uUUHksdEXS5+3u3eN/FQLG5E
wzJm1rk6h0Zt5OWnrfS51KrGuDOgUOeTHYwRQymWeNNYHvhhunQBo1penc2Fs+lvg99lHzkSHBjW
nnXQQIZfIANJpm+zhYt3hSIXOMQhU3kefKuiSCgyJ9WPerDA7vC9lSk7n27g2Bu/9FUyv0F088Fg
KmFhzNT9ktOO3k+krTL+ItZZDw9Dx6pjdPgO7M9TIe0VPeM39vpw3o9Q5S6LK1me173XP60TUmwq
UO+7KyMhjiBAc1pc4MF0FMD36ju2K8aby7F9cwCvusNBWxAy7vy+KacwFTuo9c6JbRyzazXhFQcx
T8km1RVEz/n2YW0MB1ua1QPhynxZ4BCw9fUyUKr/ysDwYySY5plhiXxkbSVVz5Qpa9Len0DqbdGN
qq5Q+pxHCi1mml/mMMxfQgDp0Gq/E1XlDN9hXcptvRpqnlB6l1CZzsn4CVcTWMPzjMsX6QoCCOG9
umrEdmSVijC3ExrWI+ir2ii/Oi8ho+Xo8sp762JyYuD3Q9KP+kLFt+46iQIfOmtNCqWUCSptQB43
PYDS+PegAq/H/hU7qX3hX0DcfEklH7lPaKnetgCI0jlzERZZRhmIWToZLvnDEbig11k5lWNWa/7n
G5Bn1kcFvfz4mrb7xzVsylZSaV/YQsKWrUWRtp5ly882o1CFtUUlzIkr0saB2XEgpaxlXsvXrhTt
uMpCeNcTt7b4RVbzYgfnkzxv9tGsYiPha11OkO1d/0lvW+b1+nBQXjM2AgVASytITQKM3VYbLmdz
Gw1fvt8gts+/by/H3ikvv9QN6rybVHPvSR5MLL3k4fHM7ooqvPRgxfHB4xPCwcRqWpk3AbFXzQD4
WPC/Rn61kXUN9M/yhXFfD7a7IhW045mK7FLuxqY2DbcxW79mlSpLwGz/71sfBKhXb0KBfwclUkhr
0cPoCmYpZ5oDOkz6ANydE3qd8epQSIy6OYLI8cwjH5m0WqbT+YYSKbdczt62HPlaPgI3harYmEf3
ZIn8joT4iDnfc34JgDTkIf4ujy3oPTgrcWv6ajlSKl8U08Lh+LTejMNZd/EWwsBO7dg6FZoIYz7o
loUUAXN1sBDvWQrjKDGaT3eJLhLrphLRbNo+TxIwJReOl/9RCtGBTwk1s7uYZHFSwKDL2Bztpqtn
dJkJK7rjDecjWAhBBijDWAp164x1hXu4e1Zksg1tBMF6peoklxS+vea3uISAjz1+seyWq68Ncmy3
k2+5IpaihOHYwoXUn+HmqTmJTv9BNn97VJulzwhKW4oc/Cl2+1j9zZEOjSdz0QG42pehwUtfEbYo
ixNOYYdsxxA85YaV2eEzUlMCMkYKxDofC724QCuME85MkjABok9zSDvprqaRl/SoWRJX5MhAub0/
JfSiO0RWLtoi4wSBv/CAYLY82PyplOr3stQLUv+WqrjiTH3SdyuZpC25XpAfwnEYoYnuaC64C9x7
u0asondvZUpJHZOBo9C9dvJgRVTIekhnliScRdGIxeU/5Sp4tHl3F2o8Jap+JMgR3aBVgn/8pKwu
WcQfRe24MDovVE0aU3EYuSIGddAadV26xZiXMn3lLs+8AZAbVvvqMRL150rWEafLytosOKaLwpL9
d8UpnIcroACQB01A4Gjj37Bul1s3chMo936tLvc0xig+2pdIb9ZAIpECDkZy1KUfmSjDodf4J44a
N9V4bXB7Rx98tIFZ97I+wb4BMKUoEglQGu5VOAe6ZxERax8pSnHcT7934tur0gDUSZeedIJE/jDP
bL50Z/or0wD3n/be3qxBuuNBUY/Q+BXSNXH75WESQgXb5cFI5GrnU2fbcYblJ68xrVi27fEwJdj8
jbuWvY4XFM4JppYNs2kMtcZzHjxgCXUjtOe1080VrjG1QowK1o43/EzBD/tk9KDqWXQ078tW3KGx
sJBXWzKZgbG2YT2rbVPD3lhkTyIkwVRpuXLSDIBbv+IGWMs3Z1+c7OZ0SwdvWjRn3VMzi3v1bR75
2SJrM7LpClQQB1LQ9EcXkLE3ZWgalP4ugBMaIuA9xz/CX5tNu1vOJ/CvilR3OU4omRC55fEAlzJb
X+Lw9MPYSgfPLWEL5ZPSepR5xBs/Ja+gDfoHPeHIX0pyvsYRas3vekdT9s7lJ6pz9WhGr5RayjGH
O6K6He/DyhwTp9Aqgg9YiktTNmF/L7lyPnBUSwdjGdUgtnMf+xMofumW7oNaQvC81A4QH6fp2Iog
fay4RVVtU+HqttSI5+gYwwlsRjB7Eps+Ms2UOMvC29LdUGsnw0Cdd7FdJ3AgcwPYFKFTnYg55SsP
Fs19teM8xwBoRwHhpQIkdM6ZSUI+UXPioTe/f0GeIaufx4gzLHNYCIwxK65i56JApuDzuXhVEeHl
Ak7Aux1EX0JhqdYfgpsVImirAub6rFe+FKgihd/PzMrBsadDBbSO2v0p8Oqc3/C3Tz0e3PtNQgzJ
ePbR5JiEkk6RW43vmdF2YfHxVHcm9cS+B+98Q46dWMSJtOdGqkD2uj8Ux2tdXsiEgL6WG9Q3YQ/D
ksxbDJ8FwtLnvDCqXM6HaYBGiCf0DN+kO5SAe1rFqyH0YN3jTev4Rwk0HNfjb+6dBufjPbSNcmvJ
B7/B9IiFtHCO+pWVzZK87GVPI8zvSV+bxMUvTdKGEVxzv88zszD7x4Ox1xK2B7vWWzz3KiP6IIXz
jX+JfG5RIZ8/8T1gJ6lqggRKn+ksBILh5lFgj33b2j0bX6dsismQgA4IKBXzHm63FQIcmJFYoey5
F8GI4+yqgygXq5enH19FGK20sqAO/T8v740XHL0kIrGB1SB3zkNm/DGqAQ+i7OYn1b2c0uFyyt4K
UWOw8ugOoRQ5zSn84etxVAYTw1ljDuU2dI6f8tnWBHdbpflB2xJgA2lke0nb3+ZquJlTpLp/7jtr
cDNl6RreVlwfGBzBM9chLiEj5+UUK1kLR/SMS3SGZ7WuhrymYXzGWfyLPFkahGXdXn7GRlrSKzeW
3oSIOmFxrC1szz8h+pHOXTNBnGseH4pR/1j50aWwyUfIJmRZZUp5x3hQlgLl1soLn7FshAipDzbi
HxeDa5t8X7vZndQZKCQ1H5gKzWZUp61ltHc3r8VVAxnqibDFBYFVnNHBz5ycWIkKtt6pnDgx40d4
etX/1kfQRVqw5b2InMCtLDPfu09ecYsnL+OavcC4KdXPvv9hQy0tL2iJ8hqctAwgavjsvkWXiKBK
GPrbyIOl08uOf7H9/KaGTvSm9UMsoXhX82yHN4/SnbaozoFrYnzoGv/sVytDpSGKxOlkr9dl7uEp
9MVx88SmasH57GozTITPQZgU7rTrr+ZEWm74F2VXRGZ6iCaIpIz0C/xenXr7MygA9NB5rqRKQWrH
AEYm4n8EuU0vbarkK2HlJs6KuIgclBzKLFjOoAFyof7aIn6nnHebStN267Aku7sjgjDQyi27tQ3k
yaGu0S4S3xGeB+zIIPxllQGJwq2+QeuAQtLx1x95TNAyas/RAatHcSKlln5clrozCInEVA6YoY3e
QpUdGnymEDaGEBwiq10X+IApSG/ZpvzzFr3pMKCExXOqCdmNvENqU4TlYvEO8tyTmuwv98V1o3bB
z5iTKfUa35Y8dfcwGgWqNkwxeQi0LllNhMZBgfNSoTCviHRzz5SSq1A269kR2UNYStGadgXvjFsb
/iF7BbOvjIEya98QdbTYbADoScbuFAAGKthEeC8boeY1t5Z/Lnx8rinclI7ZWHYYG5CzIJKhqe/+
gXM+0mGyXwKmhi5EW8Eulm91Kw/WtqzI29tNwmpCSpxdjrcHM3P4KT+XTa4krghLTUHU3XKGzwbF
niSuUgqyTV8+PN5GOXdlmaYJt9We5/F6naXQb0c2wANWmjeGg/J+MA/OUaX0Cl/mc7IRCuCB5XIR
S/gE+sr4ts9/mV+MnPSe5ZZMMcD/J0uNs1VFakWd6yqUxgZKJmO6fDBnGIdhJJIbaQBYSPsy9iJE
pT5Bk1UfS44RZ6h48sdVi0VAL9G4ucWX8efE6c1l3RlSjGBAUo1EaqEX6wxknVYSJnYGEQxIono7
+WGd8C5I2dGFXV2i+dmnbRAW15HnyVTLSP6nY4DGAn22vAjvJIjlEYyPHSQfzP9X9Mt7q4OgRou8
BIvjjKtAoW/liwkNtqQfI+R3JDyCpI8/04jpSKqxqiE5qcqhj5tzxkEnK6mr/noRs3tc41P2tCVu
MWDRkYBtxjqLchwcFFRCHtkzoSDGVzVeqRb/01x7mJRkPLSDRo2uDGYZUfehNQYLxEBHxV/PGmh9
jqTAk3L1ynMik8xDk6+O+A5ia9FFesAseWZhdT4TH0hJ+RSmt7HJmNNYi8M4QVpn9lIaO6guFkIL
sOmOQ5r4xWONtQS4kQPb5OAX2G4Z1PrRwdW834r1I/8HwMQHSsxu4Eck9E6kJNN1Y/KlrQuCINCV
hst2lVXqf/t+HJU7lUBTwtDyHhtzKcfKWnHZZrongFsqw6APGfQ/np+BvCZIg27GD2L4zhHa5O9U
gKwnkLsv0+133Ex+BRk3yHWcyvA62x0SHDS4y55bqCJmXPh4OXvaVoN41dD5avJGcwcILP5AXoHg
w2WcvCD6q3/ojjpdmHfNtKDoyo1XqcdfPyA597dbeuuZ/tc8/frfEhc6chCBPzvUinok0PcWFOXz
74yOZl6dV0KZINdYD7uP/fKBCLf3OgoU0ESP7tkC8r4Pk/fb3123SPUmReeNQVsYI5iyczBab/9K
eFo+QiDNwn2eK/Kyaqxejtfh/ZxSx1ZHzTW5dWqDswTZJM0axIL/WQxIzm0qPu325Z6iIgHRBU7i
j0SAk9HW3U3hHkOsqj6mfnVf9hctqXJk7fHM/fY8QHGhwXCwqx2b94x5WitW/HxNd0vq8GRpfiHo
LRq1spYc4JHrtLLb+tb84v/B/Yvr3yqENYhOchVNCsE4nR26cxDxoebkSLgE6AIT4xAyzNffXN7X
vDfcdch9dYODWVXZ/NFMVex7mWxVbfMn99JpP6895T2uTfy9Y2RHdcOPoJLLV+dyp9rjrd4m6dxz
vhNGu4LLZV4VDP42VEKBAZl/h+e2ImNOipZsXOaKR6dSm6kRTBGVSLVMiZkCA8ctw3FZ3c3IFG/l
d/hak9tqYKd2ulxcidl+fsZv2m0bk1fJkjnuRsdbw0ajxFLie28Mv/DcZvO35tO+Ln/QcnndPTPO
b7XKaolCiBX8yOL/YMBu6GWDf3H29fWKLDZV/UxYD2LgRyHL9YIh9DHyx6fl4WeQPnnLelEeKqS7
t6KcwH32ENs5owEYym4xjLMXMBDGPAsE5zp3L/gpHfNzNi/uWeI6J08kuTA9JK5pQt78v8059Oew
MbOsLuKvtZ2cq3sPIzqc/IV+n3kAVdAvUPkvOEXanB0CwHP+HnW93P9xq7PYbIxX+e+mqZWB96di
LtBmpBZK6Z62AwJK216hqpXikFNUrNKPitai8M0XOAon34DcWbRJKd+/7fiRTPh5Ub9xSaESsxWZ
MClc7AY6n6guTs2GrhkOuCoj9NBKyZCRa8hz1iXWUBWDuA9RflmVfWBIAgDbeKatIlxWe3lHla0j
jwmbKTx6QTz/SGB98qXLtuOp3dOCITE9wixNUGUKWXU37HPi93zQ4a48ta2og3CqfsBuYMpkRj1U
5O8A6Pmasp8ML3UpZXngXLx6hK/QVCEc+nQW5dsyblxjkx75jAUyBybvqTWSxywNXjJergycSK3V
I55++sopUNczw2R3PHKSyfmuCADgFd/uxBVZejsMfEunSn+P3hytCAOPiFw0S3Pml/T2DperD3R5
chfPg5FvSlHbGxzZ+JOlxyGCpU3ZUQUw1D/gpsT3x5AEbw6IYm1C1qaNaVNjRJQi+kKImuSbf0Zc
nnNwuSjmc9igLmJ2nf21IV6JW4vUvr1hf43+5zPFqHRjVnISS905zJrFmRtAD4elksCY5xlHthOa
8du/c6QS/ZK8x/l0YcW17P21Yw/aWJUlyXXxuf/Yc6LbT+dsgkBnmFpJB+ofGDGPoBg+HRsKdMQg
SS6owHIFP0wrWqXAeWmcQDAgNxt43FQ7SkPVKHfgQG7+fJhrkL+0ppIKSFYkAZan9rPd7Joq9sZ/
HCsEGq53WsnJdDy06xu1cb4V9sAyXzc4hAfFaaVyOsAK+piEoH23J+ocszqbXw6uR7b06gbLYt4r
MvJNyN2DsVdIuOIWbJ7DI5Pp0sGAd2El4fSI0ZhZlK+fQld0OoZKn26A1X+wvWHncX6Uql1lureG
g1rOJdhCYBHQRA9i7urc+fi+69UOx/yCACeJO86LpIKPoEoRvFeslQQz8dR0S2UVT+Jc59BZXYhi
19Lo9Z+d7Bqg3CphaWfFAsNp05N3+bEJ752dWa0MRgd5Pns1Hz64MARZBHhM+EFgHOtuEekixQ7B
mZwEZWsqOcnpmRUOd/ARNHEjoTEBefC/Vmenop+RnceBKJjW1v1Ph72BuEuSSPOajeuGrLcm0kWT
fL3mCM3F9n7zprHpSZP2XUnXvK42LshCvzBdI0ut8H5dhgxGCJwmW1IcGFEGzI6wi+que7ts9wH0
u2wF0AHj4PcwvlXMuG6OXDmKxxeXK8xRGEWve9NY3B/8Je3W601w0WnEa3mRFJjpGiwvtkQ25rU2
DryD+x0P7bFJUm5Il8uaQp3GKDjz7gB2xgNbGg/zBRZga/U+WWJJ7na2L4bzz3jv9bkvu8QAj8QQ
3sUF6tGT4+iriCPyk8K5RtJV54W6mDVzDSYJnTQjFAmKZYxwvccDw5N2JRG9TPfEMHPWOwdVHM+g
K2tjnthegEsorwrQEZnU2EckvOib2YQjzWt8r9eaN7GyEtg6aQuqWwGYMEbtjTX5ii2WionYh4rN
NeHynz1eb9qTWQFtJHNAXW/4qMY8fE6XireR28kBBsPhT3isVVwro51tAaikzhp7Mzp7zamg6WpU
Y48cqkGddOxJOrz9C86ZZRTOkyCrD4Zob12VAp1csFGQKgH7IJySvLYVoSR9+uOpwdFbt+IT9wG5
EioR0ipguJZ/g/YrN9JwBDSHQph7AH/QT4h2D7cPw6IYamhVWo8UvFYxZGXkxnf9oILcTgpbbaLe
B8CyzfUeAZtubAW7klBp5g0+a1B7QIbZ6hAzkJfyfIRhs1O6vakoTqutlhyjkrxZENwmc+JL+rOw
EJbvW/MeEjlJjfyuRTLlzjuvYh8BsJQaXk10YA06Q1NbyKWbMwo/Lcp+DyXhnu310q0deUd8oO0A
/iRL/gjungga4VJtYFfvHcncfm5JLk2+B3lPfc+EhQbRbAw5jtZdG8d5e5cDRBfye+C2xl6fLu8G
H5/m1ru+GR0a/v4x5TgH1uRMD5Do2Oj6idBsJSpIZMcInfDVj9eQjSGvYdaSkq4YaSTQFZLvw7Sp
tkdwVTZlX3P3m+youthajiDisU7UebU9xdAfbJan43StTv+EaLXkbJgOAtBxKaiEOoFzNQ/sO6GN
aBJDRE0dbGhTO6M6U1JcG0JVHG4tIpAPIpsc3ihkZoUM0IQMNWfuChezqKT8Kna5OrtgbAu1zC6H
eDc3ughabZHi0t0fzqIrBpP1qjnSbAJLF97zlIyWabtj6sHr04FnDFIMbcvcgsXvJFipqlHEAd+w
mFw/hsZBeKaFHDUOJcWTUYfT+AW4W9BNIBrfoUblhd7lgs1Zond+1FoBWdHx6cO7pzK/Gw1FCxVs
wMkPMyoNxT57ixcRa+Diqm8skdDQm1V+j0qnP3I0GJcMrgREed9fP4gbgWJX7TqPKIlzWM29mt2a
NiciOvf7GKIgZGSHkukYlQmi0Cw9Acmul/gtXqjV7klRN0tUN5p9/hDNtldi9qjP8MD5RihkAoaC
w15FsJIOUmUyULRNj6PTG5g9Z2zbexdJ/haSqNgJ3yfJdFv4QwPNQYCCJNxYAeHeagZJpcQGP/lx
CY/pkxfu0qq6lOsTBhOiEELzxcXPdxTJPQywFJpdVbWXcMLPEC3j6CZXoYzmrqyIwEyMnMQQSO98
TldIbm+F/ssFKYELxUrmrGP0ueO8CW4MXPjspa4Z2ED1p+RVIDiBZliFRISp5mcYJDHVQDEjhCJm
BlljGDmeT/bT8/KBVHS8gOmloBsrMm4uBf/VtiHYy+fZthI5MmDw0S3E7oOm4UvPt4woZEO4zODP
ylfvx+pgvhpw7ZSqbx3AopGt+9iEpUjTEU8JIv4O6cyh9N5GBlTMs1RehzM7S0Mao3+7YQEInrRI
xMsIh55jAjjAEt7pYJqKmZZOGIJJ6XjHpf6TcH9RATKoogr5F3OF76xJ1q/NDdTGgSr8GdrbjWqj
TnJQWUSjshav37Yc2MsorViFZY692fPcX4H7ItfcxX+8wir14dxr22J1smIOd7HGOESlAYcFISnV
/4GEu+9TWSKUmd5yLLWRlb9RqDNFAuBl0E9ISzs7Fx0LtspzyaLra8POAyS9rcWmP77hXon9iozS
bfaX88zDp5fzeA+kg40LBQ+0ICUiQ6uD0sncHSwETFM8bpvRHxry5SbPOCl0mO3xGul8DYtvNS5K
kl9gh0LSZAm+ttY4yMXNAvFOnHc+1KDQIyIydtXnwyCd0Vh2BtQ4s+LJUeO/e502a3lPsX9ZvKeo
qQBXAm0CEJhsmQ++onVDtgvvUiVga5cseX8ShHHp+Z14DoCz7JUeFcucNmR8H3i1ZdDiALmrS0NI
AV1m0lwi8Q5yeis41RIQxwv3kB6kuWiPkjEdhv8ddivAvrfXtXmNyP3Aw+u3DSDc+vQxzlJeLmtt
NoA+OIQjbEU0LdwzSBT2A/zeyWD8vgQPHOhSLGfhvRh/KLPCcLLvwHbpZJRpBrgqk9GZv2q19j1S
tAITB6KWneVhF53ce5T9BsDuTjmI6JT9rMzjktoXwxx8WoQLBOVBnKtGanp8d1DLpRhIc/8jMW/T
hI2cMeYGoMt5W/mysPBu93ME4JDW7Hl1d5P2OSek8133Or/zI/vIrPVglZmMbNlclmMc42zBJxO/
RuHzcOCuziTYSk9nVC4kl8WtfxV3VBa0SwRlubXPHaqZiQ6C0daJ2wuI9p66lAJViPhem9RsesjT
pZ56ocgQu0YJeP+pCgRSStLFunBVDkxgql9gCRfMqmBO1LtlbtPm7pEcWEEGvanjYdQubi9DsolX
sE55A3EO/JTjbCpHXWdcE7f9mZb5tMET6BugcMJJyt+WnHl0v4Z6DX7nzOhxr6B1svZXNAuVgnAg
1vbUVGydAu3/8TPSOzAHdWbJ41LY35QE/nr8CWHqqCgen+J2FP4/y0PbYHZNNf2/TWI1O+NYffXT
pGT3CwCcvxDAang3WYBFDUGP4lYWNDB2XZ1HDqInWKq120BTYb6dteSMWOxJdSbeIeFpZGNDOgWJ
UEyWkOcqoji++RxPdpxG59yUdE4HxlG6Nz7ditaE+unZv3xvBiV5NB2f8vEZH1j2/crGZSYV/72Z
7JYb89RQRppJMCmCtI/CBvYpWMFcA0u0aM+K60yOkQguMOL95bwOfWXqSrlcwZpaY73N3EhQqqSd
y2uZnvs6xa2NdHh/XfB8ep/xzubceGnQuw7Fy0/p1yY5uG+At1RbK+NTBa901RNDCO2rwW4gYHDE
RUjob3TCiKudegGtB5oZu0UdU4CRk9nxug1hG+IcNn6hyMV5XJtT7SRjaOhaE7nIu93T0qUoEvIx
dqrxjVizR6RLdjQtesB6MaaN9uFKGIUIGQ3h6AkfjlRwPcc+yCvBBjjQ2704UjjsffQ06PY2S2G9
kSPC9Vd5HO00aLbsmwZI+oKtIh5ZmYd322uV2citl1r5jzsYQeWFhVF/SdTOSdgqbeFFmIZFLSMz
OlALYWxclGZrkS/QqpB7xkaI8n0+378+jotKp0oUfd4XArZ74UpQiScGIkLEm+/nqGOVPFUrqOOW
nvzaulRQLnsh5wDJAVjbbFapNW+NOqgerIMbNeXO11XK3KG2LgOYq0aLTSd43s7lm7SJXhYCgaY8
WlJN0jFpEC9TsV5kIwS2HYfGvpaum1lZn9Hh2Z+f6T7/aRRWvV6NKjcw11zeFRSpRp3aVDq2pTnT
gy7hf/r7VUF+tlb/EFML8zlI97gMv5mPBiplireKRXR+g15tJkQEEMH4JAtWTY9bo6CUbuFicdBw
p+77wPnY3yAWARDnkAG3KvQMh5mWgTYqvzuayXlKks62FUpJqaS4WyOk7tlj9fSYGx0yc4Okhm7b
R2feCVQO5t1qkjQAyFJu9ENG7SZ9EVKNKKU6Do5L9uJzwJaS4UQUjRUsxuHX00om3cOgsU3/khr3
YMi2FOEp698OgbdN+rGEA/tBijaClfvtgbmg79M5c04DD4tDnrLWdRYw8pEOuDYGZAQ7O18iZ8zb
a03E4SSZKQnaP0UZ0axWIocF8w6ExHVub9KhVu1ObOYp5/giBzlym1Ee+CK7o4YKNqU4ntlVBWp6
jVEwI3EQvIjl5+LtRisTyLm3xSahKTOWArQr3Vtro0IvF8Z9VlkhOxT2qUWxeOT/50jJoTLrk8Td
jWR6UzPbmRl+m+3WH6TMqKKAaMXqfpeN14Py6prKETqvRd2rEF/BMiLCSmKo38Lnu5cG6YR9/U+n
8AGFG+mzs+/tPi33y0J4gb/c/22izwlkxmY/cFMXry/Nmfz2qXewydP/4hblKxwH4TcBmN9uu0wO
EQvUAhxR+ZRRcIcQ4H0LQZgXXxikp0ALULWObslpLlQA+yjtilSZDDIDVwA8y630Ru2Uk5RDmJTm
eBG3ispYBq4wPKO0RzfL0eolRqwr2/auv8wHtu9OZ/MY+XRzclj/gy7kKSSmuc2NWpQwBYDRVMEp
o7jISuH0NdbUT/gJhjfzTfjzQCseHwc+9GEj/y+cfTKKmCSeEHzIjvA2rfxcNSDsAnvr2AWYdXUs
tjGf1rSx7/dd5Y4mnym+pkj1ZPYHIqirwBxjHXBifrp3btWyLR1YAbdT7PR2lYz7Bv+WQPT6bA3v
G26BW5WEkw0nnKRKkyZcnc/DFIeSkbhdu5w9SDx64j3L0gF/LbsFA7VRIuzY7ye2WGUdM45uUB8L
NPt/pUUnP5Is1DAwRCIxlrm2+ls6F+rtLSYe+eSv29nyFZCeGY2ySnAHXoqsAvUsKOMIgUn5A3ix
lAQMDlmHNkeMuZllpAMfEfj+FsxmPAGzMzHttPZIdajWcysfoLV0378IJAQdUDHSl5u+WeufI5g2
3AzUrdE5KnDIm9d/90R+/oE5xltVqgtj6KVaJ9eX/bfyCrqmTeW5eS2E3wfKeHTLvFY44q5KOhkn
OuqwLsHSou2cqZuD3zG6rrnO8gGDpvUPvBOPHTvfw1JfLnedLWBVGllmAD5tZ4kI2LOnVN2bMv1k
vhGr8aeGl9CaIjRrYnBBs7P0qQGRMu7K/JiqMQsGjlGjYskh3plouYH3o7QK/XfuY/+sb4wAn8B4
63yn+W3MXq6RVNDvD3micGKxHgb45HfRthZsW5nnrzxlJ9bSt98+Td8TB+o8MkJ82J28RuhCTMvP
Is+f9JzSylS8fyuJ4MsSigi0vGJ/5m5SXYT+V1E3+4GKUDXLO2LQc/KdRGqloRivjJr7y7rpnxeu
db/ZKghVMN0i4/zCsHleLkLfvZf8fS1KHTrXUtizSg0BQgqdqCqtUoA0VqtkfF66fkAlUOB7KNbu
/JKxwEo0bCNkzdQTGzn8AuOGpuxXn9RgBVnTP1MFQ/g9H+m6avC56kczEZ+/XHEvV3ekgLx4TjJ0
Nu527o73hAtMtxueF6s97qM5iGd7XaMyEharPWXXJkvAALB40N2Qo6TY14vaZoORV8TBTNEwitPa
pLDVliFV3pznnq4zKhUl+kV1Z8tPoy7IfXe4YsgiE2L5UiIyPonJgC12jTOLimssCCBTVjQ7/7xs
E/UnFp0/UKIsRsJGMYELGL4DOoWmGIjWcvLzu/WY+A/v8y/PxrEem+BI/V9GdXrmothEebvFx0D3
qJLlVPbHx2upZQjeEqSiokPA9axkc/WQr3YfeNFtknWJmbaqUm9gmspMvyDuWA8IJo1FNui/wYMM
V4h1YqAAc0uhiKgBWcd1tOFfGVFgiCYuJoJj+x9ymfZ5ANI15xlLExT+X47WNlqWPdHt8iA/Rnq9
I78oQOokhPpzaWQsbiTATFGNHxBMO5Qe/dReZId7iyCGyP95ckqGP36TVGwDIMfl9ZM+G0Dfc22V
J3SWQgrQSbKr92JNEo6U8seRZyHDPLE3o9wxVHNDjaUmc5TA6H2A5Mzyl6nevcajKuOcjc8VKJhs
BLHlusDTxDSEgJJwliUwdgcqEIUPXBfIJZTVvgeT4HGDkkBnOBVrsMivJz/Qqj/5bYYlxLQ+LJc4
8+aBTBtF4xKQmPe4E+aCJV+ctYE4cQIjT/Wm8KMUYuJB+X5q4kbqBO1W0uRiwFACdo4hXlMNh/tb
FioPW4MM4ln1C/a5kJkXdNPLiqo1B5jOqDHH+tvCH5XpM1l3ncb/TrzF/Gv59L2OWyuK1orGkyPK
1plMlqGi+XiJAQK/TZ1SfBocpBZp2ZiSN8h+Oz9+zaL+pTygj7YskQv4TrtJHYsj1quS+9EkrZxM
9jUTMQawVvYZ89dsBynRVGyEfI8ecNECQSSa8UOqsrz1LXRkbAkUwsucA/dn4BJElQi5AZSUwHAB
64C1FaCQAEOmPaqmFdoElUXJsfam53DpAdR5/YaJ/5tbdrgpNdrAWJXzBT8Bp/KviTASkNuJAQBU
yz2IMldO8ueAeVfewKyu4YGRv1lnTHSJKLkgUZHKot9j0yhvPH4xadjwpy/bbP5ZIeIaLdHraqxN
PWfxeAhXWSNwr2P/PQUinz/t1dOaKe7V8bnDsIS6sft2fXQV1AnH3to46Irqrz2fyvE0TOPftiAJ
GVcyvbMH/7+y9+YqQyZLqfOEMAvIKARr3X4XXKTmSKMWTbspE5FE6J1boQpPYIauFmUngf0MIiGf
RBLRWa9jdVSrFbIPPEfe2noY/nrmFI3hnzrMvrL5Z3Z9Dn/BblqQTZ68oCj0zizv+ynes3o4QUEz
NZFkYDnfvM1Fzd9nyA7zCxeqbZz9/PUAN8g4iZudRsaAbGum+YSItCgf7Ws1rFK9O49RnSeBkQYo
b3Iym7PMVjp45WHgUZ7ADaVjtijT20PMoKQ3p8P5BkshraWl4tdG2UspdGoq/KcMfjwBb9Ci0T1K
4hgNhW8QTNpGLEM3jWXAY0OFSeO86Jk4aghR2aIvrLSJ2pPi/zlZ9Ro9Xl6XydPYuMbNEXd0rDXf
XAGklwEzmRKGgitbT9I8rG4pKDLsr27Uqcm+56niI1/YV2TcAenvkk1J16gwRwlJEu+ILBWbI911
H0n2x7Rb6Hus+mLrHY79KCRkyNfcLTFB7ka2lGi/wvglyrUAyXXTS7azlPxxkQD55eAKItO3/iIi
J8CpN0AMn3t5zv6HJpr99Ugfg3XwUOJKL6/hSnjL8/YUx7xzdSJTdxiBozb0cJ2ro3niYM4UixF7
3HaOdQdYpjXl+mgPoWfd4aFrjORTSuEaFoLAZX8jcM22JJxnaOqBSMFIDm+8BtYNITbP+kTaHR9M
mxsSoj03UlkgeDdcFuLZC3LX6gwbc9SSQ4vq7JcfiKbfZmOO8emGOvaLUb/9TQtFJpZDltfmMegf
EClf8JB7PeYRSBMn96r5fVdGMuhMTTju85LcQjfasrkJX6Y1tNemKDTfkbLyUYj8Gap6ivzIjX/2
OVEDb1HuHvCDN8AWvwdSDblxHDQO/g6RFBiyn1RxhXZtlyUdulWW9moRYsXaoUjWBM9K83mdJNe8
zqn4mVsXyRsKrhpj5ZxSZxfNGKRas0pVgXEEKSadJUbJJfAxU2b3GG5GQ3Ig2OpmSHaMfIZY8ibf
5nObmKobwVyKzDWUAFF76YqgL51OAM5RDLszCji2LvAXCEjtjKhLgtEM7gTMGAdTLcNJj9D/C/Qb
7RqIObkaHWFal+hy/iF3kHPaIBKMdjxOp7KAIGo0SNdgc0ZFT5V3WiFi8kk4ZMQkUTPWg3Ia5mwS
ya2jGQL1yRubK1B7/1DYO0dlfH6puLayBNEAIaaRGxJYfoKaifrsuf1EC+c33hsCm2iA0GAseTSa
T5W8+27GPpfZTIu+MDE5OPiFJmDvbPAfdlOQmqz/IHu4I+GA7gb2U5VsVSOWhGtF0ybGXXhJuNrj
rpOxW9l4S5vDoEfYXs+y5+MweiFjAd7pYmKWjH4uw1yS+yvbtbpJjHLNgvY4TYholcVchcatf77d
ph2y3Z+XyH6r83RFr3Hoq2jZV1IjqYSp8i2MoJYUUj0dmBjkyySyYBfMXWvd1QvXWYFs+t5/TyII
I/gDOkkQUOmUTbWURDJ3m1E/+XwK31w0nd/VEFHAFPENsrL2w6KxMKK9bYla0GL3SAnMc0q9Fdhn
h/MOUCJfEpKl5q1bgtt6UbqmoQe9j54pfszmtdI5fA7hL4sKBZf2ME1EJZ4LMiG+jjt27EGOIqqc
HDvmu839NPY6EUuz4if6ou2TMhpczijFESiLlWAnHUOiq5VTK3VGTcUot5w6o0GljYWZ4Bs9hS1f
mBGk3TdA4hKYJp/SLNquyMY8SXuNnxq4RY/ZmdNjrnrDdYtWCmN8aVnSqWB4FUXJYqWLU2r6YsFc
Bo9HygitMDJfJUVXtkSgtaEJFO+klhK8BAL7YAQUUunwYHGAow5e3SryLRj6Hk5IUKJiDmi9Tgj4
gpaPzMXXxzuIkrcr8L3emYd4LS3bLXfC2qDc/6RPjB5xIyDXxkOZKYxmA3ujXs+yNiGET94O1wTZ
ZFW/zCATszIzPrFx+l5E78Nru3oO0uGhZfJmnNhLEkMyyr79qstx2fJcEFP4ZmaGavUcIUYfry5X
oNp373O+Bv4TaaQzhk9yCu5kiMG2BdUiKXLKfR4enYMjmfESbFZSMRDg0hw/M8pc6xPtHFXfq/pu
U4QHIx3oA74tVby/duu1D/skuunfT50xIJIr6mcbr0stj7buc/8yJGUreN9nAwJs/o7ammIyfRN5
TQSpSoSRSlownBaq5l0wFWJzFLBBtfkknil2Fve5sX16bo+FmKSMIQlJ2qE9PA7k8AgKf2IOyjFN
JDLPgrTqPmDIHwUweCJWoP7x75kKb7rBSCaHctyvw7U1dNmSy2fx7RKE4E5L8W3HvjC2+xN94aI/
ORSx0AIUVbIsg7LqNiLv7/eRSzwykjE1oDVoF3FGUrRyrVhhHD0LVDOPF83OTdID9qQSleFZLoXt
wRwUPqH/cCSvko4UfMw8QdmQvnq/LFzNC6DfNbEEYneZoDGshTTg9R0yWoSzFLCJ/M3j9VHJY454
20uYYfYaG7AmPR1n+xQjeRxVWjUw1DE54DQVeqllM+uvzftX8Q4mrA78LmXeRs9QzU3jTQHCj298
B5d1blf3AxhES+LRn08/nWDLTLtsqtixfcTFgCqemE8fVJuCG8UtLxQDShx+i9B8nz5bfiTE7QG6
Vv47ahC+dW9iuBPs299T20HNFPwbXEDkz/H1D3E6QKU+1iGxG3F9/01h1yEzSpInhxiVcyxKZyaN
/5Gg3AbIG7CvszKJeDwDbNm9TaHHlSw3n7NCBt5YRRAfXEWmqziqKMbX+jlAV1MIPmxPfhGuZd4N
7DCnDDyjWZ7E1ET71+rTJNbGxIgrgAPt90XUldPFTWRGDmgyW6EI24NA4GZaRqKk8bsfmVcdaZAk
HBUsr2sJ0NsBqakNeJSa0gDrRvilKkK8u97eVgusw6+KORwDiWzBX04SCrSSHTJhexaB4C921lf5
9TEVUp8K64z7HpeonAKOrGhl5bm9LQ+XDZnQuKzyNEQBrmnFwnUY3RZjgfb8A5VttMQcz7xR/vvU
WT6xadaThxERANWfbxb/0PkU08BS7gVseoTsEpOif5EFeHGo2+6+35uEzLw6NNbBi16q4ZeeRmOS
rg6vbnfTYGd4GymOJS760eH+mdeNFSv/UEONRoy75weVJha01JeomnyRRotYQVKRXZJ3pRbrf3Kn
guAVMLKi4Dyqw1nYH7QKHy+Cmnxe1qdd2rc5BqgoJD1A+D6Y5L0K8Lfq4Kkn+7LWFPGWYIYaF1eW
bkPpyTRH7Nc9wrZ5GXajgpTPwoIcXtzpT4FUnIVmE6RllX/OofdqlVrY134KWgJwPH8tD+p0zith
93aCtMqKyrx1yX9QjbbLiHGfAnsr0z6W2rAOUY/Jm9h62V4Dhn6EdnBsgT9h5V6hkpTA2iy2Umxg
qfpYAaXcC3Y5Xp+Zwo1ZZPejlAxjhXDkkqYMOD4VlZQy6EQ1DIQpYKCCAMKJGWX0spIp8Tosiv/m
RU57CCSnjq2ikGllMNuNBTwnChJyAUD1Ho/P9xSFBb3zi8xvziwFdhj9BssXImI41pCIRzJnWDVE
hSxQ0bisUlxFekl2N6qf9Ee6L5kXiT2jap8cM29uTJCrOgHsb85YgdkXEiEKWwvG1Lpd+7lm9cQ4
IpZogQQgWPhiMYI6wtVYIjXVvB48TT16g0IgvObfZAbYFuti7nuxWviA/p9NYidgUkGB1gvMZ/Jl
bRdcbwefb5GfRk5aUmUTTx/QarImU6sKWD4TzigWqgAFgkDMrVlzTcalXH9F9S2xUWV1iAv4CJYI
zkAGnZy+BY7m/8rAbEnE/mkjS+9fDAnN0uHyhpu5BGVVan8o6ss4XddQEaLnFmNhNP8l9gWQq5mc
yCIJ9NRMs78oSyvSnVALwSjb/G97dsTmNM62DkmHF6qsBIqTMxY1dltYJ9ZP63PKihhHMgwXSBr+
vcBRoIkPK6RFViwEse0OFRiDlfgY7v/8hOzpaFkQOXJUUH69h2WIGy4NjQTOBp12ihVvQEkpDEGo
lpYVeaSAYJ9od4lMqx4zs28Nkyms9ujHrscTly5mfiK9IT/PHFIFyGZjnqXeDHWzFw+fEVrIGNiC
Ps1MwPbRcrza55jh1PIk2tyJdU7ulJ0sbDKw7puIUC5/LlN5GqVMIHnlwTJvHrXeNp4/KzzRwdZk
RoMFmH6MIWdp69IinftcNmPltxtLxutictL6/ifARjToAGLOslx3OO/NjNZTV41kYoRA/xRySjx+
VCidDrf5GSPgkGdY1+yS+kYGAemFQCG0tIz0DyWaq+brX9l8+f0KRQvGhCClLl9GfDwfaN+HsW0j
XLhRpHbTVNSdDkfuJEWw0xU/Ohe3xpOuI7Le9NLnaXbxg4EyaDFsROGIq8EdM6OsW3NryCVBlp8q
orFVIbE/7mJHyOGgYBcnc9CBzPJJ8Is55nKHNLLe77fnwLiViBXP94ZhS11LQaS5nldJc27O/l3/
aohz15QZbvxUGtkUtEbiH9ANEAVKk2rKtd5aTLqkpa0G4en0aAAOQtm3qTCMy8traoHkJC+IwUV8
WISC2V6dsDi7FAI7OZnTyY4Qf78k7l+4ANDb51jdwqsmiZ3WIJ7gW5WFmkIyP+mVVJSZvM1R5BWe
u0H67QLQRZ26gj+7VWM3Gpf/h0yyNflB4lx7SCnI4S99qxw4edvwaonFVbVAayw5XVmHtQMZtv8h
KhNt2s7S9KGD50P6t/KhXrtsU8rVJdY2nbJLlUo975B4yuESSe5dllMd+G1bXxbXYumF1eukw/uQ
qX74N7vHpf6js8OKS66TykJMvv1rsNNBH0/zJTJQthkTIAHVOb6PZdGTXXcXmw6uKMTpKtY6B7pT
FBla5nzayQxRka3Wn0+gJqVpWljPRrGSfz3puYhdY6WntpgmYo7sB7krsjg1PpIJt6cAeRpUzMsl
YQcDaZfmLyOHP+cPc8j3aOtgadF1NlMBSzRhn5LNabOqzA3Ym4aCQDrHuxt9meaG1HLIi7GSFUVX
Q+enqTuL1HyI1Ng5cJqlqPbgNTfEj/pUBFeH++vzjaRiuQY+mxj978EwzeT3lbkEJHLF6W0y50pT
PjReQIaG1/gjSS4m8hNzDX3grOiQfAKBW1638t5q01C+QZEwj/YyrpRUYIpekk+b3Np4Wl9F6EuQ
9rL31tLx4sk2O4kQvLNRwUw3Wy8Rmgt3GCruRbFHCB/5GqGmgdN1u31N3mwu2BiKRwq+ZUJ7DfHS
XSbkxi1PQ1qtbpsdFSZKo6Su7+WdbzM71UU7JZvUH3XSscwZZojuL3hSSCh/u0o+xS09MbT1vDAZ
adbjvjvtcX5o5pDYNlqQcgPN1YIMotwCZq5DClFmTlRNDCSZgnDjRxCU2YPCl8kXFxm8aa6+lDq8
g/TEaWpRWdJSW7XGiPk5ZpKXMBp1zHgyaHn+8+iHeXlJ3Yn5eGO9e+yBhoYk+reFTFM60DafiSw5
PJwsFIoo+vb7PDjU9F14er/hmC4sKISCgR0n/xduOQRyvJE/HoPTpI9y+xtUeLgrV1J7Yx5q90JN
5KDGrO+EKD4OFsGLq1RD3AgFojGIhJDbKiHzU6lq1XTIUbOibmrfJtaZVRce3+t1EmqmatvkcM5w
t444grCLCwhnayVI+xXBeSrJqsBU+H2kCum8O2lOyMgKfP3n856N+ekCfkaGPHQCRwB3V1QkgBgM
MJ92M/DeD127kdcDnts5IJBzEPynnWR0LTIacDthNJOcWew1MNOkSZsm2ihnxdKffTI3HYvhHJPc
VouZ/d9dAVIrprICoizcJ5n4iA7j993kRo06wBmz9g5N910/ST8cf68l4nyfdkrukEnHCQbt3BWG
crkFdDlpxhS8H4nJ+lT1HSue49NVEYLOZZSSkLy8YcLl1UFaJWDkdsYVlBc055dyDlJ4UXd9DJfb
PGdAM0Tleh4U5IobcLkV8shC57w4tJPi6zg3avWTX2F60DpuulzVTugfVwqeuOYo18y7kuNqbqul
hhahaQoMytmEYgAaB52mMQCdg2WoOQbH4xr1kiikz0Qnr/h7Zd0lOuShdwrKmCgA69AbINkvoibD
sQUrRu6BNhtFkHsuOpBnPTVU/lVt6mEZv4/Y3YONQNDzK+LwMd+3mh3UiZ7JLJiUZv3LhIxNGC9R
zk3Ft+pUZIOl0B89P+WTQUoUrPHGVpKGE9C+rkJ7atWSRrBEbJd8ctWWZIXz/OBg3ypIill7XVFx
+gm2Mp3Va/xXpOayUfBCC/kUgw/yHqJyu/huiM2fHKhtHdrSRQDy2FFpzOeoLrH1kXOh14F4dOWr
VFYzW3W/D/uu9DI7/JVTGSPHBP5e0d2xR7PoHykhWevJnGqIClbr/YSKCtvwsq67AwPdJDmDq/+b
D4Hm3fXhw84wUhXIF2hQKqXPamyz6p71DIeD+hpkjmpWqpTfjBvHvzHbwMlW8JlS6AJCNyPRgqfe
DmtMYTXvfdgonpTFQR08OWyQZn+BQcwhyHBAX//NxiMVR4MUtTaVHJiVeFhh+606w97eUSlTFadN
Lmirrel1QkQnIdemlg10Th1eLVGJyE0rBENmd/KtQ1fEcwkUu/B1ot2H1sVtHMetxHYANs0SmMeu
MQ01+WMAXBj56ypwn3v+O7wd4G4SBKxJWZn85gJvQ1JNgW3FPHkkTyZV03P/PCPKE5s4AprgRyeO
Mc+RMpQaliHgcXyGCWqqaB9/4dx1s+GRYzVcQpQiQplg4V1knjfOFnY9UYg5q9HEX5/Kk1TZfm/G
fItQlXvYQ5V4CE9PURQ5Yp/IXD1aMgjYhzRjRQTVVGl8/iRwekefx455VdrrNxnCzwyqrSW3vuBl
MBKnu6Xl7J1h6dwDJ8euz0UX4a4/fZy6YwigL8apKFvujzpIzp76ju0VOmX7jBd1P8qzO0eYzg2l
XspE0yiz4z9B5gWNeeFfbyi7z8WU7XPgqjIfTc04FUVyYenlD5NqW1ChIjbXuNXq1qQ3oSy6A6Um
uQOYe2h3p2Rg5Paw2N8/CfH9ZGSdpDbkZtzVvr1SrnCNF6rz6NcXXqiIH+ZLtqNowgmapA/eiLme
vk/W1afcn8lx2scKEimcytuo/5SpXnkl9UBP8uUOyvVg84llCkG8mykynaiEm2A2M+338WXqXauw
HYhfD7hxy56hziOozMXFA4wVQFGWYOJ33J7EOLYRblzEgSPirPis9KI2L+hOLwk8M8n4xS8WfJbO
3EMQKo+pf2YJzyDe3S3hq09z7NMWkrkYyK88/O4JxCuWi9w7TK95AultQ89KBYnQAh8fvQ9KyS8i
CH2DqUMwHFMEuGijPaDCW6lZODLvg6K1bQ3PFH7TZQR6bqTzvGhqZbv8NZGeX+b+7LDMspWbS6/v
rTpB+/v2b/iKWy+7oBGJMNKTutenHvcbimWlEnUEFOkf+Hk0hg0uI9lnRhTV3GSkIqdyd17Qf6T5
4hjc/nireFY69rvPy8EBuuBDQcMvv/CWn0hbzrv2DRtC2+IQUQ5gEAAgER/YSJ7q5RbvNMky0fW5
H6IfE5NvSQ5k3LuEqhn1NoD4CvK2KMxgKVCESHL6jw8z7BurcEMNDNEu5xtflzkNjsTdEj7l6fGi
2O5vRkqrNeilMKYGINc1TFlSIktmkA4/8N+8PA2DGWoWiPhsprTuTS2qpoavX3dPPM3i0HkyzlRA
qCSOG3IQQoPHkKZgslmirHv8sO+O8LNoNoOLdmQjOsNPb2jmP5khF9z6vL3/zlM+Ud5WLe91nTET
LTgvXS9hBJ8GDXDfYj3mzErMGkxs2GZ9ofMTc9SV/J3oAGKMgaBbGiVXjuHvRoKMgpGNQRPEKhH/
RMJe8xikZUPzXG65wIOV8aMeE2wmUCwOaaNjiruxEbNhX6zrCMVerUr2390LFGTO2rRdLMVPcxS4
6zl4PCi7WFeooOwtLRIybT/v9jpCF1KTLXt1ilOlg7OUnC6BNv0rXwk+Tsx6B9kHSf8e0E2MvGgZ
k+xiCuWqcj1Sr0oVbfOkO+k/Se1+Bb8kXn1x9ENT/KtnpATNQTSOvX0x2og+zZdP7REjucio1er2
JVXVMoOwCgmmsa857GGRa1CztV8jiDd53XynIR2N91RP+Z6rv5jN77jYJFtUnKpFFLik4lGbBLRp
v1vI6Acvx/tZo6fiRABmSx09MCMbgy3gO+gXjpA/UETv9s77g8vGqFpyARlOFyCFD4+AV8OEnstg
p+TsROwzDa4KPbkVcrRBr/a427DObpZGGAHbrtsywzLL4fc3wvOg96QszHbLkURz9MACw+I7Q1bx
deY1NcCk2CMfzTFxvuJJB67cwKJHXrTbFjDlkVmoC0z3HFP2pKvrUv06sfKeVTv2b+zlQ1zbPZFV
096+MIppO5LqSznIwRlxnnDZR/yMlnjBrp0uurWmBjhsrbu9sBPOk2+4UtwWaxzZcOwg3iZeZKBO
C+gZ5W6AOryYC2JMn2h2EYNmM83+a3REL+QnxebgMhMyTibo4fkT0sGvGUkB41uvGL4pE/mVUC/6
4RSiawMXbt0j4a+dRHL3HHxF0coAQGAeMj6gRkVg6P8QXSoNXsaJx8+/lr7CPfmPiXqmIhmrfb+Y
XF4rQRdSVQuHYUtwIsQZ4xCiHqt+ohzV5842nl6lY/FconTep9LuGf6i5UU5A2IutdpLVHqXT+cj
rrg+fH2+ZTg+sMqPIEzOQoZtNY94CeKKZy6Z9XG2QhnE/NWGlnqal3/z+4+pGWhJ9n+sQzxwJgny
EvQw/h0m5UFSmShcTW0/8x6TAuQHsQnaCV3rV483xsNoY0pHpvIpdyOF3CMzQjNWvYaVdA7BOITa
LVoQmaXRp6rfrKfezFARTQdACvVtMfRlxj9smSI5BRIWJTrXeU1g750X2RwECDAcoxXyrj58g/a9
7C/i8uceSuwfXqQkW4qGKFYrujizpom/y/MGdSVMf13Sh4oXVQarUkOidiVaWSfaVzp9hLgykZA4
EVVZcAWmKPXaEWg699Me9wCCHRKHHO/HxTyUQE4ljfGJxFnsaguCIffdGn3HIgqTSQPdUeaiRTF7
ogGHAYEgIzEgUgRtDpdB2nFxYAsAmy3G+D/GaN8SA/gudNb9aNIm0tvKWWaBXlfZyyckon5EjxR9
inznEARbLr1KKQRz4DW/AkEzn1eW+BgRu7gUTRI5PG/m9GDXdcsJw1XmyoMaDzVP8118HzIWXArB
IEgRtB1OfWc6vlhHB6soVxl4nQTODTk0Dnp87VurukkiK0I4pmYDf+QoAKXz7QoWbpfuRghq3+Ys
EJRiK7aBRsIaQraLcQkQ8KDYlK3X/KPzh1swtVZIpVZae6Udp7SlMDc7QiQzoXdUM67dZ+KYsRaJ
OLCEvFaBXpr5q5JJp14r+ySslydJX2nmkSAU+X/XmPKtXqBFzruf5zAQScUB73S4LRuxyrRslA07
4ls16TV5HY4e0q1oFkXdduw+UZoUeI0xOLU+2XCEW8OhV4Dp+EAVU701pCxomiLc4MlnrYFOqN+M
YWqGLSL3TDzU8+6Mb6L8s5nA00LiqZbgYlffPWMQmjVgGkbSZL1j4TRoQHv1a5As26brmw+xg+HD
0YS2lIt/l1zHNKIYN0bKnzXBMAwEnKDAUb7P6wozwLHifGlYHh+wy8MxQMvZCYV6J8Hk2e8KSuJD
TZEzaj7RmnJdkUz3MWuPJCYoM5tES218/05fQIPCfyKnTCY7jBgsJm1wmRJtmqbC7O0qhKGBN4R3
Pc48OmzEqrK9djoTyTNkR78yHmMa3XnQZxcW9SPKERzoqu4qCg11ZubKZ87kGNoJIicp8+gQHJDn
drMtcP17OGD1pkQal04zNanQzun3IUyTuPMRoe8frU6fooYlb7M9sWkqJ2Zxm84a7d8FRr/Z2zXU
3SeYSL+UlN/C10yKblfadYQBciAuPViVKSX3uB8rZYyKwb3PNh0+A5FPHcZJcdTF4JEGYOUuX7V6
WwJWKtp+9D7yWSkhORlSTDnHF2+d7QWsoWCFziyOqAf3uFpJKDI0/69+mq+TZvLk1rpkndds+gCj
Ldu/Uw8tUEVtAuLj7Fg/dv49ebCxyyTW2fn22WyGBGm+OjxS3l5IB5/tAl0uDT62khyQCq4bljOw
VjtD+9oTKMnF9RCwWZuVdujHKnKx//MT9grwJh/2TVvv+VdHH4723rLuESKQDEZc0E2MzM4Yfq/8
oDN1YiLkF1d7KNRPP+DyYyNKheICjgl2buK24Ht0plQLmzwGBwQ6/Uke0J+q1/pxd6rI4/2LrY+0
z8kFGSrHccLEkkHgu/WBbonGoayssEwCg6VDJsM7pPjRTf6AQdAIjvNWuHNw8qGZjutfG/pYlUUe
JXpPQLZWOrko7KVGco4SsbO9v3wKhVLScnV5VSvL+Aj9tWON7riJBmPY4vjDGb8Cb9CTd187UAOr
F82FccULQGQoQNInwCxFs0UwZ3wN0Qj/nLH8JV9rSdIAZD9Nf/8GtKIV+wYJ+0pP/eEsi9CWqX9O
y6vd/O3yX1EpeEtdmebeMWZWGonYiLhdlLDZ1fYK6uH3vg71btoRE9KU5mJ6zFkZM1Mt9traIznq
Q4SuoQmgKwq/271QrX5pViwp6/NXz3dQSjpSEYuQBYrm555EgYlga0tDvg5Y241YKGzfhYWm+rMn
BsYfPgxC4rQ7hiQCKfPdUuXoWzU3Qj4s1ICyt/ka5Ug9n9EZQCQMxEeO4DJaqw+9kqYxr87i6CKH
SmzUiwoN9qgqe2LAtk3c6hWGjMj+xDWMgANaO/vvLwzz5d4J53wj415nppKKvbmpdUkCZourZCyX
YouBvhbpMwKHoSymCZrffvDugIAYEm4KK178P+s9bA0jB2vtTVnBo1nMXdBSof2qgk8Wst5YedYR
52QEtJHACChrqsO9Ocmmq2BqlEy9WXRxfQ9xZ1IUaOrYTEq+c/6Bg8TgoFrRRn61pLyfQ3CZWNCA
U4G4NqJBC7LE0Grl5e7IRLAGNG3Qp+AiLYFZivvbGHgw7Or/O9usT+EMztSjPZ3PVVqrJz4AP/ni
cBfELDtiBCdKS9AjDggL26/DIpGcTUsSBGLOH7KXapMiFvM6Cl+JHETzLT3aEljuuRvFhZm0jMwX
qhs4Q28B38tzVnFHTug4jdv2+/HhuXKkE18p1sl9nIrMpaYRdiT88gjxZVNobn1egq0SsEKSv0Qt
0XkMMPaXMGZ6JItWKGzfxQIjdztMLmawoQ8kp9+ad39AbK8Qfz4vq8mvZWGUNN1SL3rw4VhErB7m
HVffLRAEtDuslFyqHQ4Szl7fjragUcs82H9jSrBG8e+UFp0Mhuihsrmfdkl+Z4HzHMg68wckbw5M
6jBFbPRze/BNPzaoiOrs5RPiSFfNLTHeCXemNELJXr2Frj8raqvCHfo3CoCf7VFpLCNALFPo3yZc
U/EYhUMZIFBHINsAdK8rhOM+qwLrxmBXrWhwOFKPJNBpCF6a8ExHZSmukkrC4DzrYFDtpkvLBiS6
roGuQg3pZi5MpNQQ8byB66I0+gcDwnt4LYjdO7WG63mcV643pul45ZsD2Er9/mabgJi3VTUfe17E
vkgW2XCNNZuywGf7MqXJB998ThD/SQqTWew+Vh08mZMpWp7ButHdlnBtULpM4k+c1F+KoeaL2my8
S05UGQaU7thHqsDXlr4/A3UNo/23aDsJITqv64TDako0/wdyR6414Py86KJhQsBQystejd1Er9uX
9T6uIKB0znigSPGq62mJ+hEpJh2qYeNVMQz5aogmiL76nzfQEt7XXt+uOFeKA5Fl2FjJ5qMh73Mu
YyXFWiQu3TtSdgRwV9rWIvpilR+HeWhXtFKftK8WLw2ho6itXv4uDjn0VplfNfO6n3GvW3U8P4J1
NQXxdhEdLQmIV0yL64OlFu0bAflJL7bEvIjDWEBpxeIHjF6xH6Kn7uH8bBtvs20O+xE6nJdHsBUv
uiwzUnhnsAug6riwDGIh+h4vleMqlOlmcMwhC+g115pCIDtu0N6bmhrBKYj/fGWCI7Y2AR0YNdPE
7TfyLlj3n7AzpQopp5cryU2ON4/IhruCzyUp7wvvNte5xrw4+5JhbMRH8WyypByPd8ZdQUqBDV5t
L1kWF+yPY0KSMr7nLlbuVP8EH4Pxj3s0hHwabVqQVyYKlGqGXJitFyMqhQpZlMc+ygn9IhYegETg
VttaIpwBqBrq9JUOUanvbJoSRQQNZg8qWj17MY/Zc2Zo9SfHF2UsQrvhwRaN5s4itI21vRGwym75
pVSrxKfiGYcCy2ZpmESDlYh6VD83ARLXjDDTdcqlV1fXu+31EhBFtj92IASxiaH1iA0GzjjAFnIS
AySB0nd7GgzhXFRN0zAm5P5vnrWyqWmGzKyz8Y3oqTDQYbUb69S8rHG29V8iwGqJRI0lt7XssVSs
jCLWEDWzsufHxhOtuAQuaHD0rsroY1rwkYSJN0rC792FShwx9yKsk7tIXgUH4ssD8dOGuK7cQln7
GLfwitMN+UTYjs3Tz2FFbLAOIVPdtWBiIdhwtLGL70eOI2uJKjq+O9EYDKk7sHlzEG0dLagSjZvr
P796DJP2xEjDmEUXxOuMeQ4jmOhCsGKPfqsEYkWsL7d22VMBG3ILWLr2HdNnLGLPf4fd76n7F7sv
mLIFkpfch0kD610SNxnlJ0aKsHnSRxkiDGAiRs99kyvGhKvhN/D1JShW1Gl18WgzFLO537c/zefV
DLlv6ZwIMkefcb8R9jFjbEPw+Sr3PrR8cid8pcpnERlPrePXVuYzxnKGq445JHNBOaQiCGrfWVA5
5LoTL3ppYI0kxsLre2/EPNonHDUobOAhm4618iI9VX2fIGFr3/WNQ+vpinmsBHY3EvZ1x633V4oy
gShwWawm31Zz07MggNR3bConY4rdtuXq6pNbFnFeqint50upfoy6Os7l+OsHXzEQ29owLfjRlsIB
7bOEDaQfLSjwFQzmnRHyxZhMPYPYj8o0NCXI45B+qjpC/stb99pz/1Bh00cf4XWehs1u8A+udJ14
tbr53SlzCBoTayXAYhXEX3aqR3x4x3Bdbe6lxE3RO2cE7VdmvJEshElGW4mWYQph6NyHQnDTXqSW
gBzHKE9DLoizprawIv5kgbiu2RE4m4hCvYGSS49PgHNpF4IwrBG0r/epO7M4DjGOy9z6D3iDxQEu
P6e7DSrVJ+HOD3q4BytP3I/dq+B2C+TwZolBgkiiuJcB3rQFSIG/H10LldIAwzcqNQKobrxHlJXS
eHQb2XAn/9s0E9o8UPuDE9QuPxAErmLTFwiJ7v5QlyGDeR6WZMPp/u27IaxkVApa+wIHl5Vt523V
h6vtMN9E3+Im7Se0jCkwdjuUJWLONGK7mCEGj2eVpneDfQL6xzqVy6TaM7Ojk8SX/Ks18PNvjjgE
aX29RMAln/orfCoKY9jnv+NKRA6kgT6SBqu1iV/VuiXb/7x1U2PiOUGoa5YcA/bF7RAsF+WmKeLq
B7W2CM7rjbj7tGdNVMre5wCqku0dHaP3xDQcfZKWwQnWsEZuXPb0a/qIrHe5KHNxQrHYiELkmFB5
z0HBYm+heZovaiDPTdO+9V8Xdf+bDANw7MeKnTsm0Vnj++5qoyY6df+4/hhTgSbDp4/ltPld6/uM
xey2sthT5ua1yP9saBuyYOGp5EBK3Jjp1zlkxWRzKFgDA9ICR5HdHMT1X0xGqAGWhrMH5cRxgvfe
nYuE531DJGaTBQ7rzXyN41eaCgzwn3D+si30UKrsuePKmo39zHCIfZJnJcYpAl8Vp9ODIN8ITWzT
ZwxG2bFwKzTLcOAz4YlwvJmlcumhttUKmd8U+dBRtdnhYfZ9hS7DyKzJaSCPamFXeai9Pzn+d51Y
zAQKa0ciiU1mkj0A5ZQASXinueCfkOyaFxHiY7MeMgipjXr7LgqkjB4WkVfvM/RwUR5W+oRVsObU
dke+AVivbyc+t2gRsOdnuEy6Tb6Ft39Wh7nHp80JYLMiSsnLBlt/f1sX0uWdlFjmTaGQNNjl+sfr
ARggubyu0G6zvxaFIWbXp8ers31R5+M34djWSUsZQStYTonsupp17H/ygTYFWwlSUPNVqmskMFM9
HrxE9fAbBdlFYOCDxXPoCHkcW151a167Dn9OwvfvrkWUOepvwk5pa9+3w8JxW+WxEy3TePlOV0lY
WWFHr65oSB37qShx6GPRZkY6502pPFmCbGvKEDMMQzmYyipAak6r+oAZ7f2pIp4EGOoYAMrtl6UE
EgHCIseX8mtE2v+lfAYwue+a86nAaUARtVWGTZ3atGUrXuevpGcjN2oYlgu5Kq+KtJuW8BA7A4F2
OugAfQl7bsakGAY7Z84U22b43AFNBbk08J8bpQp0QcgXwWYLblxVNueBQRx5Mdt7ec4Moa3/qOdh
FB0pCi1h4wna6ZclorB2mhN6vlLzp3PLZErW4o97vyejavG3FIa4iP7DNF+a1aFMOI/4qvQLcSgq
BVqYC4bP6vHXb6lO8IltlnYumBgbxt0jf50Tlgg5f1qDRTj15fcLC+Z/M13HR/3cjOYxYxTdqCoa
fhOcm4cHtXiaEusnT18RHeiouWj0fwJu6vpwv87SId/IBFtY+BSGi785TSrwHdlrfSfqD6pVtAb+
emRSiUGC14fkMNXEKRSRa+QlGGNcEQP/g3dS3qj6In4SlGHCT0Jgm7slKO8c+32nN+5rreoWf6MF
IH2ugW+3Gnf5IP5T5BXLuvSAZ04c1km91MdVlfx8X2DE6dPdP/1FG1/D0kbl0oLZnGF894uOKgxo
P+mxlErFJAEFtdyEx3V+IJRrzxXnh9NAshW5dUhXLE471jhvk2bz89sc9QMEuQC9Dno3R+kn33a9
KOgCeAO4Fe54BRctrH08NFk9oJ3mM8ar5FbXC5yw7QiZhQqUewziPPLTknuF0t2kKtLq4HhctYat
j1ToLcrXn9C3OnmImtwbVskHcRLTvyBeXAhHDt/vbatz09SnxwIdeKQ58cSHjK2g/fEiEgc1ydPK
+NZ6wSw4SQrVT2FcgTCIFU9OpdCDrviOZgCDE7FmjQM7El8q3SXQXEtoUJPdXhfB0xMyOJSXCaZ2
+EhVOSRRJ6QJQyCOke8WmMrp0KGyhAeEFaKXKYWYm3mYH/RiuNt5AimG7LFzK6IUJ1fpqgrgzESX
raiLS4JYqg5SsoMkpVn5CQ2KO54wbwYhwvqRYtO1fdMmx8qqpYQ7+rOO1m7F4o0Ta8kDiUm+mJci
JCnWftwbiWc32Adtg3y+1KdlgKE5z4O/Mx61sUQU0OS+0s8TC8LkUxQ/V/rjAxGjH7BPFtsgj0JJ
icLz4AwAKIe9AW9MZICw1mnx2W1c7FrLxK+ql7WCtgXVRFJqrKLAsRNTeucd70XKhskKI5m1Q89w
O4uvKjJwAmv/eGes80Lqtrr+CYA9VPob7NiDCVs4eByLljnqethqmugU0zjp/nnsfWeDqsLWGhUW
FtnEK3EDkHcMutKynM77xaujEqlx3LX3nxhfiocvgEGnUzRDB1XL8AswZGWhxFCwPdpUewN4AqZe
G9oqds4RBM0E7HanVDl5qfITNL8YXZ3JQ3VXVNqYLy4sHgGcJx6LI8uy0UQPvS12mHDuoJl3EzgI
TEVhUB7Yo6a/O+vkb7i70Z/Q56Y/VjIw4AwXSdCnNe76oHdB3YQi8itjkpOU6S5D3/di84wnPfTq
hZUtJ9fIo9eUT+/mfHglPdQLQaYsP9wUUA3Om5nDz60wR+fMXQUpsERjKohg0mULq1XZXNeNDOCU
/sgU7PrKNS/19+vxaiixnfkiKPu/bBzzgetsqOlpiiDWiKQe1l5QijfWMFwa3Esa+I4WyoAfAtbe
2Nn8zBq8933aoLktoHdI34xhFVMgCOpNQIWoG/EwtrKj8CpiewoZVdIicKaAlpN38EG0kfOJ9fCK
FtPRtecHlcslndWburAl3KgRZy89ZyywOuH3Kt/McjI33rVkn00YvALXNWQfrJlwxwdjLrQx9tMX
P8YNMcChAEXMUQVy3avjuGjpemBXdJYUtz4riFFIl3Z8Cq1JhMx/JKBl/St3ka292RARwB4P5O7B
mcXiZ3CdyquvEeih418qB0c5ThChOGWsBPDrYNDGL9rcvvEIHl55nZoInxKVPgZee91tXeFH0URL
oBC0luFQqCtC+Cv5zsISWZNuhWnnPEtRMsh7cZVmdYhbiBFzZt/nPjZSP7QfcYTGNKkxeeucN0OU
NfPzFnxZIYBBuQdpKqYDessE7xH/1A9iJyGOHQAY9/LW25uvTzQ5sgSPta9WvBA9RqfDGjgMFjBa
Q1e8pEnxUr/ycL+ndVMuk+Or0ZU8Vve5ARXo9djbu3Me6f+25kwwLBxijZ5UGWcHmNO7vs15xlfq
84K1FgV2z3RkLSYNawb3GlUxVLFATrevH0VKTMhbMoQMW6VMCYw0bn+Q9GuwWY7ZKX9O9+1c9MJ0
zjPGOL5yQ2DxiNqPktc7sUzMWIM5pHgNyq1BZdwPR6VUAtr+9ZQv/ZlcBxG27L76HJhXrOQVO5sr
/BdGL0hj++aGKA1WmjQKS4KlbmF3roIpMyU4mA0f3bbT9LNqR+Y2rmMi8QWphx/w8g87+QTnOHA7
rzKK2yPKlliSMnqKl6Vf2+1SyPdHkGc3ajqnhkluHzQxegmcTM++/03e/N1Z5s+waV4D//tFxPQ7
5duYmQ0DkQJvBuyBM1qLwrTfMQKymHPHy3GD9BCy5nlPn22vrIHd9DzCQw+OwbcxN1A4s44C/sem
jCFDNRb3zaLlXAg6RUIdpARrqt48fkH1FgRPUF58Eq4SghLypNBmHlR4iOL46eoGDOQvNOP9JtJt
PlO8/vWpkDjA5iy4NB3ssSHdNqp14vdfKH4cIBgKU+vMrKh1VaGjYEo5/dEG5B7HWynTz8NgG+N/
Mndp4RWJ8WuiPE4F84dAr2ZnMfUkp2rqUk1trMwxnn+Xzi2XfHOeXzc9ekumtk0YJ2adGykJz1S1
FtzvyozqIGw+Fmd6uAnt7Gk2i7tlZaC81mMFvqFkVYMMt1VQdg0DQxg1ZTUtWI+vYiHvhhzOBI6r
OQEUR3J/1FG9T9ySERX1ANy6akUydJccHo2GvF1wlhcryz5jIAQsskPj6dvmVO4bLPoCbHQd5ICG
BLhn8z2+knBPZUwBB+LPw6UtsNRrEkickM0wmTWQGwpfwl2dm/6dP4ZAv9zBHFp0MogoRELwpyci
qgQsgBbL07yF8KE3A4gqaeiqYIVd6mqkX06M6CL5hxG8/3heKfejwEHGLwGRgup44IBspdH0tj80
2d3ugKb4fzC+obNo0k7nAKlGBZjMJYh+M4Mom3wM8swlUL3rnUd75sr5ePKimCfZKOLQ55naVnfE
vR8IkUjGNpVm+TZbwFXoGIK81lG8/trnKiRBGnRnLNkms23JD8IgcfZVLqD1CoZHxseTq5/hEnBp
t31TRGjU4cCSI7SHlCEdXmCe73DA5y7P/YdCkinBRc8xRaMT03qhpSCP7bGScarZY/L7k9ZZJtL+
Z2zykHuoxvJ3vnU70BHzwYKJGuDhjX2KNe7uif/kiqb1IN+hl9c5Debo+X2IXb4wgzGDROh64vhq
dtqT1lKCrn1w9A7wsIusttvI7JmuwbTd2rnAcbm9yrDA1mttQkgPK7snC7UvVUcqHDz7NUDy/FQj
57J0wllCtHqw0t5YaxGQ7mfAGHZ1/ToGnGtYr2jpS83wYVNPogsEDsQ3HkeAPlhXr7UrANUyE8vc
4eUIWeiXf3kLFdsKkrhvp2VT5JWR1GYBS7XcOFCSTUdkZazkPuC5fB4oZYtLpAQeNYqjGteBfTNJ
3q5Zg0CdLw7ZUiCA7UaOMHZQQE7+Qq1bGeM2fPrvFBbXCrl1HFrBx2SyFfULquLZjED0Dx9cUwdn
/nJyLenBOwwk+nRb4pHg6emi6NIv6DrfgNzDIb8gepM8yO4ARGpntJGuutOheo3EyJMqikZL9Hcy
OkcovWlnRbQOy6pMjthgzv0fGqov0BsaPt80Q33T0OHCkfS0Lu20JLU7RcKFb8pwk4a2w3mh/U4H
rMco3xZR70bNfwWmk5ZDqmbmN8VY01DWWWMZjnPCl4bXXqleQymCLHI5paKJ3KFmTn/Q+P/r+NVb
8vVxUQ1ovHbQpy1Be2ebTisZkmb0qGL2yYADP0Wry5hk14rkRvDy1N9VPmtdy6y/UjZKrw4Nov4n
yd/UD5RWB16JCFJl7lQsm/rNdPTvmDkD+jGVbfXgs+QEVNupkSIMYHMXJmt6jj/yJxnM7o8ruRsO
trJuxD1MmxAFTo0txOC89nwhfO3sPR+uboGgOn+cDtLaEPpR7q84DXZET2vbcJ2xukN6r0W2xRgA
59CYeGB1rsnAz3QW7hqFxF1oyotaLh24i9QQ29fpZrCNWrxUIMo1BAKopon/J+iCpR1nOLxSSI/q
JUAPco4wlLqahlTl7J0NippdYNZflItzdcz+v5y5DbZnzmtqagA2RWn8m9car8ZfkeNZBYXyWWK9
JeimOtcQ8fZqBqKzhnVUK6t3/arf1yR0mvn0Ov2KlAMz8LwhvWRKpqFyV+3MLQySeQWe0fL2zaLT
R9UV1ShxVNMFSDTPOzQXIqSX1DtsKqG2sBdM+YixkbcPxzVIdoUTA/k3Mali4ZmORtDWI2CgcRuQ
ksMDGFKuSgGRqkJIYaL0BW7ZX/4jX2PwJLe4zU58zeSyBit1MniVfW50MKRTNpFDAlY77wazFjWO
miIJUZsaS0QjvE6RDI61Llx9nnFiozXBq67GlykBJ2yV3L9/XdmFbrB9yRt/4Pb5t4FBF6cnBGg7
7VtuDuEW0grhkAj5/bTEUEuIzzYLxXltV8Um0CxDJ1J6SwRCAX2VJLOj58TiSToJcSIXoGnXaMCN
uh4r1bTkghCdP0aJPLg8OuNYyfkIAWH+b3wp9PcWSVdyXCVyvk91jRmSoMooKzSzUrUZy6M8nuOh
CgH7tzp9RUoEl5cOwDdbxEpDChBp6gP/y3xKumqsVIeEADfaYFYFc5gmlLUoZpvOLgSJGUTHYY9p
opPEGxIo+nbyxqQwcIStNAgP9pvJ/eff+QYf5FtoxR2w0vdG3WAcOPuZu5mG3OrLOrqouN5OK8d7
wi7GQ/G3MtlL/JnK0oyDzGYYzleZhz8MDsVkeRmfyZ98Bv1/DH7oHIjiUPwUi/2sY7Re0VIVNmtx
e4EoojFTUYWjCjpW8j/uFBrjNRRQPmp6qY0HSH88mogCZSTFWE3MaJ2CYw4WYV7s5D7vqaP3O1rd
c/iPN1+fVLRmbnitgoJkKm0fnUwxCLxn19T58QtGtG5z+9IVCeO6t3No0JRwkdVPrKdV3X7SQ8kL
TTUj6WiaOy+FbUCeIwMDou9Q66ihZ8FJRIAtPZ6JWm3NFdlwk7lYHSysMlPlGglkbsW5A3Wn2fha
zDU4GBfl/WM+EpAXYteJcFv1jfbIkTzIoXgqlVzaJ0ioyfTvPBzchU7X+Al9s/LXgfJUoA3krAsf
2vGKEchLeCoy4H84IMrF13EZ7DLCm2NlwnSTm5A1rUigQOQfOARufDfgObJsbEk8ur/QnkZii6Rh
GBqE+vJtBruVGIXZGy/EayiQRBfYftA5d7IrGRboLgdbrCeQheknR9mLSapm4A0sIzS+HJdW9jTM
8olSoZGIiGyXYNw/09GqUyLmVLDNkx0polfr4IeM2G4GUsTuPG09po7dQ1TCy3OupvWjpj9Rmchf
MksGoKsbdY6+plLeqsTgaJs4GNnmvtOY7OupSuZdHAUrRzKHbxEuGYte00FT9VQ3dWqwu0Ow5g2C
pFtvHY1NsJEYYrt9yCiOodjidXkh/cghvD2zKWan8fU7j9D6ZlOJB/n6jGqAP+3Q8nQj+tf4sXUA
9/+gv0REWIlSqoMWbNjs/i8Um4wwv3CLYmQvYXDoOg6pute5deO7D9OzblRBd7B86tqkLznV39Ji
B10wpM02I5lzQhc4X0UTNNUscuDt4DbG2oWh0WThvBrgTW898NZlAmbyMBleyeiROg44RajpzPxR
m/sa1tSmSd6kzEK2eRyf9UV/+PXB9Dvs5TE4HidWGkd5+xavq3wACZ5/iZ6vZkTCWuSsA9WETEWd
5q3NB+cIHoHm2pcUCFZQ2B6hm0kM9FKDPZ5gfifwylSYaiwTOCo4Ix1ge27QBGsBsucHJIJoVeo7
6o8owN2YZgbpwf27NJ8wCncQDMiYUMDHu64b7dv4oWteQCnykfRAP04A8oU+wnhCbNTtZMtGgu2P
LlfcT7H0wAmfP/rsHWb7x7vtC3p8vAGSA3U1D3klvVk/L6mYbtN7iGm+MxsHsmFLxtKn2SvfCd9W
epgl38CVxE929rjAWKdRdyNWwDivdLSpo5qMjfpRjGf50zNQdYb8OMVsHFU+xevBRt9XnQ50PAHJ
I+xxJk4Z99hcOXyTUqYNys++bgjX5V9ucCQLeGEk8EdB26B/+CYzj0PVL4mJY4EDfXVu1BaphRa4
i71oiWoImi5c8T5BzC5kQhMvVNnMCh297Sa3JuuemtuFWN+FctFokqS+PiK+8x2APivpSR1Ez0fa
AHs9AVRTd02oyhA6BszLeRrz6HfNpRVZDSUcSu/W5DHd0fDzAzW5hfSvOBm8fEPwF1HZbydE/qMj
2DNvREYMOvQrQiH26g9XR7ZjF0dAtw97m0ul7YWICMD1snjM25xByrHpoTSTVGV8j3fOol+xFZ3C
XzzVGSpEtiQ3Y7fO+0qNaMmm2P7B4+DHUi6jhc9dwSUnNHt2zEi2ZzsZlkW3iWotYL8ygkQWVg/S
DeW80tHRT7nClKi63w5+wnINgNjA8NbE4Yo25+K/jNSJB0WQiiGi+Ltopt0uTCMv4JHUbLJN0iWl
4LuGSP1FwpcpEnv+uJFNALHnvyqvxJRM6NcJwlczBrFA7XVsuWzTMv7RbEnZ+kMnSwHWLwuZADeI
5/BV9gAmtpJYErszgAkL6NV3BljzPW5j0HQgLr0qPxlmYW3yyycfc5g7AZCXH9akbVS+iRjZ1XYS
Sr4zy3vgaGv9Oyytu13cf5/0KoYOIeii3jFjh9YCUrEOdwdFVv0mrpbVJT0N8rKC48va1Vcr+bv4
SmEzNN3kU/R2Gbtz3ozZjUHqcjB54KDZVMw+/PscSQj+egDkznySkfcVJIFbEN92uxGL1b2WecLN
QKBWXAf4uaxJxpkKFqNQ20CKFY+q0jSyRN7eEwvmHqyDXbnFxyh4OhgI6tv430taVPMm/781PLuy
JqmAITGkdcm1VTUYEiCaGrgG7MDm2UY5m1ooXEZmYhi+jUQIvInCF5euGBAXfsBuUqw2g56Q8VPL
pniKGb7y0DZ6uVyEzO974FKX/vhPAClHddtFPu71POjvD3rXB2wVazmHGX1FoCJjmukZfWcWVHR1
UM6CVIwcBfNzd/BqhA0vcYjMtvhhV1BApRJssnbiqnhKERqJAzmnaEEut7MMqVJfqhUz24mH7Khx
Z4xKxKpheMoCZ1JeWo6QzvPKyl30AwclZKV0kv4p+XqHcHMH1fMRcyGyTHZy3CxqBN2s5UA6zjDp
mbbNbQZ27HNoL/ZZuHuDGrM3zCdsplLWB95QBNPWSK5fMx5C9hU1zVri6V9BKtf0Qu5Z+Il933Ih
mEidrV44FqnTQ2MB0+6fzEwoQ/VZ1VDngHfRE64boMzQxXgaTJJ2+jqRFh3PRQfxtCcRkdQDRLnB
iMJpHAQiz924dXWfS+fs6R7zDNfA5OiPjvD8Bs780bimItOnD3EP9aaCFTOH0XDhHLO6xREbiPnS
QqCS5h4FI2C+kDBHUxhnhURMxmzRkgZryA3HSZxTdEdmki4I9G9+MMDg5AvAhvO7i5xC1wO8bhN6
Aw+oRTyRV3LHCZr+w11MdjEP8OnqeiDKqdT6fnu9K2r3Inv9TDIdhIYvq1BqPapy7G0zgTfiqj1Q
d+ac91QAmrK3OFg2HKgQtkq+qKukfriWr5vWXYY9crzVVEjBLtgEAh9yTffhDtp/tugvXtCz6ojb
RtPeKPCGUDLwVjZpLqPy6sgAir/3pBcBPk8fxr1BekDAn1/9tta1I6xThgQ4sAXzhMwDQxI/sq9d
r3Qhs3Z4s/vZ3c71NucBL+oOQaUyqPkcqXCNLF77IpRVPYBTYKMjqr5P2d7JIUCr14fSj2mUyQ0s
2/yxtAJ6+is0l3LJG2lFre5yjgUgQJJxeIT8rHwLk6qRjljQaRLEgbUjF++VcneAf6u3hxjB6nj9
/4aQuINnzrbCEHBJNxgjnRJ1hVbI+0Y/WoLpA9rOlyPvXYZIhFfisa4EYWNUbyP8d5GFG8XU4fpE
lVXI6r/TAOnwq9+wdWK4qfRMu51mCteXI/w+hpN+JiXpnqfpx+uoftdWVGoV3iSI0mb1Hc4glac0
4o9vr0VYIcC1a8yek0PHHTAP6mxayPcS5j6P215UdnScd29PrOH8WsMSFVdm/GsVX0fxZyV9yu/E
AOt2XkcgLp144m2gETXx+TFlBzdyzXwZK5fBHBZsdbZYfN7UV9KUMpBZG9UHzw34T3mg8Fp3nm/h
CqYCUmewfrLlvKARh3uLIH6VkrHNURLGxh0KCm4h5MWxQymd1Pju3ZnyjSugoUDUoCEYaqnG+eT6
FVkjyJ3bgKm4Wq6PU3Rz2BMm7i/Y3w6KF5ovsBD5oTkWyBQSdAvJuWcae3KJbie8Pq4ykXaUeua9
Rf9XLGmf5v0x18R3SXZVyE00vAErRfkTjpPwmq+f7Pu2vlpq6YgD6JxKNIfNThEJ+8o4cWSNoSt7
uCJDBdHOcoBi+OuB5KpeSshQG3MR9ujN1vVfGpST/vg+tV/aN5T6VHIN5ZYZCxZTc7bxzyri6x1+
vsRm/4yrlYQ/nPq67eMZ8T3nMdZ1ZMk3ZJmFPN8mTW+xmBc5MFRydN/1eCwfe8vZizbJtUNElWST
9iuPA//ZYR9qrAqSCVlbEXzMZV8i8Ea64YoGALl3+MTUd62/Xc+RRLvuDVWhQNfiL3zFSrmu9lwd
FuKL9hFW/eYX0Fx5zpsmWcBUrfvDSJEGcLeYCcOZZP6X+0pZT6FyFBvxjApO+qXhHnFmXURgzyaz
QguOvkcSsd03cwR6zPDKFI/uSC3SSPWBAJ9rFIASe2bqre/JcsRfc3peGtNlziKa9fqnTf2ulCfa
22SlMNQmbSrGFgC3KLsLTfq4Azw1dG56XuyA/zloOU4SsWjTEx2L25QfV9LNyOWw3qbcBKLjRXYu
nFt4YcU8fWKjkaTHOyiG6VAGgxEViHLCBSesLlF6SrolpyFDlMzBKyutEjZPfwZx6/HR7ZxYdRLm
pYVy722ZAKzLuTsPAs50LGbhFuUoGOa/yo6Kqgxe67hw9yog0pxZs2FdnLi2r81LomitP25r2OLu
5RO7c1Y6xFhfKa0+mAMFgYEuMGX2KiG7nmgRicLhHr/lP59C2AcMmQjJahwPDZ0XdSxehgmWpkje
FFLfHUXmdFwN5+uDp0IBKrXZ4682Zvn4IHkdBfmUC9SdnfK4SIz2eOsw1GCB2uynyj/iHHA4C4t7
ONASPgUPs0J6uxtdLgaMJe4TlA+9k1nB8Wo/pYasWY2D+DLIZNioYPWXyK2bgWOb8qv9S9nRzUlJ
WarVRiSW9XBX7/8k728EfaX2S2uq4xyor0ya2gbwFfnj+GmpNQE5ca9pj50HgtEQOxLQ4Gb/RJqj
w2oEMCk1xr+10hDoGKTF2DrMH14jUOo5V0ERyi8ck7vph0Qkp0ljk/zxd3spWmGhQx8U2Gg2s2qM
A4+Bgrkixpt2m2KP14xTJj8KYCFkUc9Rgv7rR85SCS+kiDCFybVBFXqAyaew3MNRECLy3k0JkrIa
9Fc2p1ikL3S9z2pL/QTcD7GXIf+8/Sa6URQsoqAdcjF/0HTObXlsCdcfV1h+GlKyxxJRsRLg73d7
bM9mpte3WFv0aGp3YgHe6KdO0C4ARdvbTH52IasYpmuM87PaqPbM4L3zSE6Z4Yt01h+YOsrzZVQj
ZFAAakHd9TGy8G6NfHd88kkAzZLk0Zn7vM4oZkjL0fVvG2BbPqImqP5NghBxH7w4Gi/9Plyl9Tts
9oMnGp8PfmLQ1IK6Yo8Q9gcTG6mDUoUuER6IWNdgfA6NcAt8BKS/+C1QLBqTvvjDUFoOfh4UqcA4
W2E0dNaaCZEN42b0dzxzjBQXFIdOXkUjFAg4wGh19TOTxNDfORoNki7F0yzN00CtIs7qj8yI1Yi0
4uifg6kdYdZ6nl0S6P1kh3ogCr1IjtD3pdTwiwbf2n74k9HzwzuKTb3vNRfkPuRHNhf5taF08a9m
ntcqKa0472tQpXI8oBUkfg3juNJN1cGA9swX6VVnETUhFjXUkXUd1vNfdvq8V+6ELYuBt0O/yBx6
1pjHV3fwJe3oCTsDKlMELeuQ/Dyn9D5F0spiX7taVgRzYqkqSbTJsgLcrPW9PTWXyjV/gbtzjnMK
Dw5WbriMidqA4Yh8EAgdx17cW0nDfXp8WtVYGXjGkDKONtAxbWZhe+DRfv50V24Qt7Hoh1VacrJG
4lb4a2m5HyfJhQAa6ITBF0esUgQqZP+ECw1wMhtXcHQecagrVNRGfqwwTIgrlw8tir9JUVe6YJ8m
n3jMEy0FONceV0TKf2Ie7lplwVF9HZV1/58/DW+FGa05uTQvwFbW01/hvzqv6YrQtkrhkvVzaGo6
qDCIyvahMN/RJfCyyXKMHy0wFAAFmDyDvI6d9YaAnsHX1rfTFifoB9uBMNvqH0sb+Qxf4Lv1qOSu
A4GWLvo63sF2skv6f5YEIRL/SLvW2d6MT1qaKV3YqEn2OyCrd0Tvue/SeaMYSPU6oNz+jcNZdf8W
IQ0LGT1q0uRQh3WdQ2FLuRBgWww7fe8+tNn8yHxlATu3XH6kAQHepDNVu0ILDZl75qbju8zE1bBn
D2txsASLyvgQZ4nd3VRKwShp7m7WixGHZiJ0IuLdNClKmg7aDZH4OmZmnnUf6nL0zbtPwPBbWo/K
D85Dm+GMTlVquqTKoxiiIB0oeHs30F9G7cYb/MnipRkyjMtztmwGhTHM6/woqSFEdbhEczxMuUnz
d5crGDPsvgXQiWNMHPG+ohR/3mg6JLnMpX7xCG5c92F6++Wz0YNeb9ze+HE5y4o9+SFBbXJrc9mx
jXvMUj8CIdbDMLzcs6bD2hl+3r67YCEdFbep6+ajaUjKMcsVp8KCwqaPD2jqsIZntIQJLctjVe0q
3vK04QjMRCagT/b7Jl2erEmSyrZK5n8S78mCLFJyQ1pbTLOzp0N+8fMtjasO3DmArwoPkqdWIp82
JH4uLemCtirfbHH5Qp7dtUFhzaW9uwYtheHdqBZ7tocKfjUsDEa0PtgWQRliDrLJLoz63cWL7ktl
UhVQ/ZP/agsXgKzg2YaS+IsSaLHVIAOcArhISUXepEN4Xa38alhEY8GnjTfxEBBxLezsQ0NNkrid
KTpJJWezoCEf9Oi8GBr9tR9xMYGjrhVnFGy6vJEW3veZ/xE/B4pySNnIXbqIqkko7AqLMTQgLrUN
OZFc2+0+D5O3iweRGxTaZuTUL4Iwylw8Ope2zOe9L2lW5kZdCb5hf7gJJxUZowIp9jNFbWPOv/2E
LfDx3vM1gLfYxiSFbcfm/fhWusYTgMneWn50YboMa6Cklyme3kIiipxGRodLIVp4Ys80EoBT5M17
s4/M+1GI6U9RjUU8CxyCNLRBUVWElJrbSyKlofebhxIFpse0jANxFkq3h9Gc6c9F/wT4aG3qQmX7
9EHgA+ofawRQJBqTG9dyo4gPsZ14/ymyDga9K8ldttEBakQxdxajs6NydYwHhwnU6etLx8YnwR9h
2sqhQaWXZeL5cCsFiCaw4fHtv5rhZw9lHhnGiU1b90sZWugf8x6rYcuAhTBZltEne+IfLWGGu9tC
TCzwbykNQ791zRUmx2KsrPpWmLghuj6huBw/hdI2GIfsRFHiPqOS8FHXP8cIsVNe3Q/c86I6fsrS
CFA7cq7rSI3XxMH9CFYPF43AJseaKWZ6HPMtFpA3UmxY3x/8KEhslQBv7IZlhgzFe8lYGGkL3wrH
2gzHmBbwRuuuDeBlcuaJiV9zw92XfygNy4ua8L8jEbC426586jXk6lajz23cI+T0OXiAqyNJWo9l
abgTtYCyZGw2BCkckt+KvDw3Tm8UE1cnX4gqfbuqpTZ/+eHOJCD+j1rOB9Km7AEH5mnp/Ngf9mIx
L2sX2vcmcDSgcVpbIqZRKjNZPGKLBx/UfhjMpUGBhrtL1C4+aUo3G5Emg4IAQ3QX5Eb6zGWfpBvn
xKUGfMU3vPk0ouYNMDx9hrmImVSd8ylP1bLxV5e4qIkGUtsVUVWyWPgdAwRGZzjvGhTciMKAxjHC
CuJBmc0/ZcdFcD9YCJaFV4azZq70cxv3NBpZmmP1E4Uzu4VHXX3+TBB/7TEbV0Yq5DM/QdEyDRUC
cRXEZkIX63Wl0PWZn9bHPGfnO6Dfq8xwNFKLd7U6onVTYLKPA0XCzV27LxUiA1x/mikvIWPtYVws
BOrSVV1vK2TbNmRQIgYukXGJNugzZao+ybFzo/bwKzHCkHo4FtIyk1WgHkPDHPUlkHEoDvoLSJy1
gNaM8vNwAPtOI7aXXvDpsGhfW5j6ZiiAeB72SMABy5c0FrKRUTR/Wz6jBOn2ODbfWc772qNLHkEr
IJA9IU0PIEJpZW8ZzUZqYH8EIXTz47isrOGB6Uk5MkmHlWGy7zjZLqeT5JhI7/zboBkWzsVqO00v
pGPMYnMlgD72YlzjA7nFQOh4R9Jf+HsToKB6Foj+Emj4wVqxKWsRJwvaLn0X7lf2EX4vIJ6N4NsT
Ugp44qu671Y0DgeosZUTOhml14JScpAO6cPX5S/YrbaG4ehYNZrZQvgOyAJWfYzEIbjevA7ftmJu
G//LW8KnsflmSHdOjUgxzmVnByF8oYK2zc7ThhVSAeXLYuax6345S1J+onRYHuj5C2+fB3Bhg5Bt
NCwSGqaTZKjsof1mqkoJZ5yBUjaSIklGpM+XEDjDz63EgJdMDxkMhEfDCO2M5BqeD4RKe53pA94R
lK0K63cY+HS4OwRc5wsQP6JpDLEqoTPlVp9QI+AzJE3Qiqr6LVzRYyzSuV3zl0Ktv3rQDmmrXkjW
sMoyQksJA0tRNh07D/LRisAp056M+86W+yAfu/CvqnZz31GJhWZ1oF88/0ngKXmvjVPb/Q/BqhDU
xVUmsicgxuk77hu7YuB8KN/6QPeAuB++V2CBfyCwmwCyoSdae4uL4T/qto7PwvV5YRF+MN8GQahU
cgVdE3gGXksecEOTYRVYv6J7cZ8XOQvy3gmmo64LNVz6WGpJDk+9DBV7FfGXkC8z3aVtSsj+hrKK
UCzu14JLaqs45FNrdXYVG+UZU5v8+v4aC+bhlM1maJy8gXJ8ZlCfdXb7rPHtk8YlJ0GunlX8rMP8
MUYtWjk75w4koFFvvI4sC7mBVDIayOFK0w4cPB54fNDaBnmehmBf1HR1+8a2uIRxRQGSW1AWVMYC
D2WGRiq+RgI5E1h2kwTzVcpnZHoJQxWw2PzeyI59pcyYplc19X8wea67YHkExyaUnl7RM5kSjbDX
F1vJVzALLq6NAtSqL+SqHc9Ix1E9+zF8XQ9jBqJxEWMeMZ9FizNk2WA5kPHxE+TXawYVuTGX2E9f
M0TQozQI6DX6uMSHvZvmLsMH74mA0wOmHvaO6W/Q0fsqJ6lTzrBrRsRNTIU4DrjoLH5IDgNLf9Xi
c4A48hKSdsNPwbKfbpsoSM0MnP7WwmZy2SV50tGHDjyYQRhtipemYzj+gnFuAOFO8qvv9Co2XNtG
UxPvUfXjTdRClKxAbSztOfO5UcOW6GpKDQ8dvPxL2ut4vgx2+CSQ2OFhIeoFmfml6RlnflQFFFiz
XQwOJH1gIUBe/g6Pv3+d3HvMKYTgfQQiYuzbkcNn6Gaz10TUUlSqXYnbgLg8N7nH2XBiGjLR+njF
W5TF7R2CtKK+1M9TUnqUeaQbkyjlixtVo2nE0Hb5XLG6G1il0gm1uNSQ7lrqlKabDbGE6pkUNn5s
+7OWCyVBDt5PQ9BrY6CkIC5LPYpE9fFga9eUMD+tVeI/7qB0QxcEP9K2o1hAHr4Rf78wClBjizDT
fgXf7vCyF8i3qV3Kr03g9AN6KT+G7Qvd7n6DS1COsZFyCM9srHSaxUwvUwpFrT42EDfHMGGkpa0y
A7KehbvH03LJzdw1gvbSte1TOMbhnfSL0aHBoelArn/AbgLhD6dRaEyBjPOeIGQxYvlgpGrMxtpg
0ZBH+sYs9wpz4vVOZj7mzsaiCmlvvKfq+FVizx67YEMSkdM2ViKiZZhd6+2YTGQ4+d7d0MpwirFf
U5635dTEhfvPznxqzuCqqtMSogXI8sAsLccMfScR9CbmzAZCPfPqqIbKxaZBTVGqmTocNLpfMMU8
G+yV3UCVQmj3i0AVBxiCj19YcamDcEZfHXDkqbWkq5g6v4MALYdKY0V+Hz98wDmkxU96Iog4CN9k
B8fdla5BB0PT8Dm03OD6y78YddjSf3M43aphdg3OEswu3YLp5uR4rwDFL4FBKVCRz2eO6eLSVL7q
m7dtP4TKFXkw0QhpTfi3e/FEAhAm7MYiUyqf0JqPlgmyZbDRS0XroB2LFO65q2BgJPX+qljWq6YZ
gGY316zeGAz+XwRRAKlBQKMSgLY4yH+L8A+wKi5Rm9FQIS17VKvbdI66zKXDDwOUQ5kySj0ntPSf
7TWMG0uCyhOSM6wmKX2m8NmU4QGM1FI3j8jakR1M2kF8vTA4JWWc3DL7PzmIf/TOmb2fXiHwJ6PA
nNal1Tp/6T88TqBz2icIsN2Evp6cpTWeC0e3SuPAtCtlt+D1vbEqq4BLFB692V1d6zEXx1X+1bpy
bpWXhkyQS/De9OFeKE+yNH1S+OJvfHGF1Pd5Y+1cQLqnY7W0J5xd1U1pOkJrwxXkSDMRRMANWP6e
L0nei0djOXbeaJTaaQQdVpCCJmvgYXZgkg10tEoQHYMQ+EqWvKG8u4FOVHSwDWofBRYlx2wSHDA+
zPkQrZXtyrk0hEf1plH1plQUEU7g5Ny1XNNS5MUsQHrLRFhoFnPEeuEIE+zkq0EJZGA2wNTDFOyD
Ms1lpRPc1KPNG+XLUq0N+PJEIV1UR7d0oopJ6+WTqYNcUMRa1IXDI9bi0VIv1ms1YvWrjb3dADC8
SMC5ZUuKQbVsSGgg3fxmHWYM115RW3FE3cDgKBVCFGAxb4bTXZW8aALrWkE/KwKMdpxIkNpyKTkE
r2sHd0aUHu7UvpoaKzqviboKus2wdoniz6BsmUq6AFeN3qojsj7LduvrZxcoZc0bsWK5NHm8NzpF
LKGPPGcSvhEBzrw72/NLQGFhuTGFoR5xxmRoATH9w9QvILz0yDBOIz4cdlFdXpNl2Paqm58AX04Y
19/zPud6uZ6qhQyYtTFBZQXVOAbnpqvS47/ocOs1frC+IoxFcf2VoH8d6H+b6e7T6fPnF6e1Nw1V
Ngf0Tor3v/HGE40bHhY5H0Zvt+s45ubtrRVV7gYlcdxfkbUnOaEXs3WOb890P40cBZpCNO0kMhDt
zzlVkBit4ZT4TZxgf5rj2gDKdpZ5vpp4UVRlfIDbg9QEv1iP5rnNhtVgqgfZoCQBY3x7oERSMNI7
JjBzFM+1avk2JiCiI26MSVOL1EV03e4RGRw2bY5C2C0Lv5hGz404JwryBOe0rNad1gQrrYlHXd/2
6IXVqYQpbnSeQxnXUFAnsL/F83e0NInsjNPhqJxLDV16P1bDtorRoN4LHOitiXwUGE29NkwCMAQy
HTCcvTmNyS4bbjPvpiWxTFu2Cnc2Opsd7/z0v4qbFd7Mx6ZCc3oXbzdlUSFJE2Jmp/0gGsTHpfML
1rv6FWjmcQYU/AhrguDkPjhkoY/H6bVvH7BOOb/iYNlUalN/+17icDbXFlL0bRK4pbTAREHlEJL+
dZTZtHzLiv1PCAKZFjgdkXSCTtgmjUthGHuprt29Dr04VWMtFd0j3km8tzTFF+3ibUNJcJYShPep
woBik5j3FUKdkmtNAec0p19h8YWZYzQGhhn3EwAxtnI0JgcMuCW1MusQZdXKEf/ghchO4g6RRIaf
xCaJn94uGbw0/r95sPf+Fp3Yx0ewdZh/aJGQBKH7rxxYXqg5YSFL/tSOyz2I/z/LNitchlgyH8Pu
bVeEYlYlvcKwgWqf8HFNdTBm5a+LlpO80QNxcDwNZDLDOM/fKPoMk1WgOee+W6/XmEUpTpqOmCn5
T7AWsvO5a1fVMetcqPQD4KTP0f7uVL7IOFa+uS/gnZBz7vQmmCbe3PMk1kj2sahAOU1Tm+M4X+QG
QQp38fhWAxyukBCOcdaOwwxSB1qXIhYRmGAx8BR40Kj0w3zYv2b5BAEyM5iR+8XvisvAaFgFoI2E
gce7dWy+F/iiUrUwjiFCcqo4zoysPJ3ZAk7blKC1qqEB7dLsOy/OfQ5H+Zh0yE1gAKfpWwblc8OA
N4ibtphMtFyVxqsLTrxYwAd4xvW9FVf9Ms3KPxpQrhC3/VfQyVeOAf787Kelv3LzZ7CzMV3mVNlv
fB3OWdkeI7QnSKRIk4BWXdBb4X/n5x21tQWEYm5MmCYcH0J4nBMFzWXovN3EgyZk4mCv+In9bhFh
ulxdmdsmSkX1EcmCnOBAsbj17BUefhtqVwocuNOVkKs4Kl1PAlQgknKrYdq7NSqroapoPifQ4Cdi
iLrTDsYKQiDrKppKaDHP1/i6agk2OgCio0pPSNAJsN6vJcq3HkOHv3gbdcDPlmxA8mXlq1XFydwx
cXV+o3aJjjGepRRKNW+J3wP5170NSVFrh8cXTlSVXrPbI5dyh6r30VvzE1HWgddqefyx7VcB+wkp
4usxVSSpstVbeeYHFupD3vOquli2GGjcL7VGkcuYVPTugj2L5NbP79++rvAXTRdmSz/yVnSwy2Y7
IAXLyR5kqKcsQWDjSkQohy2fMoAl1IE2FUigTnoZcch1yZ0/G6/+a1o7ImUtYytcdyWceFG36gpg
R+YJ3W1RpL8cVLA7QqolDYfqT3Kptesq5ESclxTbRfVNi869j8arXVE/v7NHp+WZQMx1uiq1REx+
u9/iCFd8nzMH4sG/XEAVKcxwHZ+5zoyAmKOkqE3tv2h7dIf4locj5SlpbP0fWPRWOn3Ov6XdkNO2
+HDKWkP1xthwB4zFxMvMIOozZ0raxaS2iXRbdJtrVfU8tJUCKfro/BRrhBfn6EccWdrsGmlXIX0M
Xi7SsJOUtBEG6GaoeFoXyFKLBiFAW9poETdBGtaVfBNVCs+I24TtYypQCHLbOyt02dxNVKRl+jE6
+m81hrKCXZqU/btxVSb8L0zdvxedZK/DBj0leLZHN0z1PBWFP2i8/4hd6qNaLjAbCr1MfECsnrFv
GTWdbrj7aaI0YHQXm2pBp+NnTEfC6oCyDFQ5GjYPS2toFnnIbXy2HrtnZGuJeIsdR2ESOl/G2ZJT
GYIvy6I+R0I530CQO7DXe8m1tyVWtE1Lzg5RbxOFdlqxvaOONXW1v9Xf7RNfTZMJkPxFbPP7RVBv
tBQUA4LadYyuDRk6Uga2ia9UgIyrc+5hKaJw1E0lN7TGN8Y7djatsnYS12Hdu908stpegg/fSQQr
rHoCDUC8q9N3QSocRRC+P22SgRyjc9wJk2flcwd6nacS6UtafRdJq5dUWwkBl7G7XQRKq4d2jRNB
4h9QbrW/LikxlSbWYDy/YdVbU+vSHs8Z1N5cI0OTMhgkQreJQ2uI/uEsQTK+pK5F1hP6e1+GzoqC
17+v1dVTS+UAofPtnheQvqwqpbfy3QM0svYD9zAHERPUpdbP3YtQC6JiBoHJRDhopyDxfeMNBDto
cRj08Ihoaz7iuHb93ClokicJK4TwrwaUw9h7eaYxozczOpPLTZLFNFEQOJnDapXyoyECEUgAhr37
uTwJ4jBN8OHqwt7fbxftB2imcWYHxv0+UMh50muehNAdFC2lxr+PMub9NFucRK1Lm2AymLJDgL9c
JRrdVQzWfLkMMM5SM7dYnF5+xI72od8Qj20Hk85pi+wyb5GFpIgUNARdMp023UNEMgaCo+7cz7hC
Uw4OMOzEOulrmeT4ur62h12yuVNSsCS534Aq2DIPQaz5CkXpnSpsnZyywlfdnbiGLlBianb0Xz8L
CosHzupyJMLMcOAtKEPUb3BMOXOg78D0OSXvbj2nJqHM997DRg2mr/S26bogZzT+exRTm+hVEFLq
4HBgCq5gt68IHmMkDTG2XQOHqrt39AZM5V8O3VauFD1E8jf61Mgaywb3F7BuZk1HIvZ+WTaQcVbC
CRKkSRmqdAi6a+8xfbw7CGggM71CQfAUlaIhUg19l5vErJ5cZif2CcYjfS+1z8pgYmwec3G0PLR7
GsGFvoNFY0GrU9sKjHtPggLDcBO33wPn6py73kfo4akCanewPSK5lgowTHVak60RZeeqbPfApDdV
Kxw8xYxNfX1MPbd+okUvI4h28xC0t2lbhE0u6S/YN4PEeX4lENCjAplwtHbzji4RIcAyG+veSBgW
f2O4/aDsmuL8WBeI43eN9dqaRnbrTu2YQWnUnYSwqo2bwZUxeIR2z676UEo3ndDUTdSRWKbItXb1
EC9IKf8In912iLrW062TnUrvqUfOC7AarUA9mbc9Pw2c+ZuLozS7plp/UrPAaQvPNAM/L+9YqbvN
UCRZQG4swRvLMuSYBCChef0OHYH1S7Ea7V0irRcmfNoXo6rCDAAwXa7Cy2Coi4buOxce3wvsTpFl
8nM5HfkLp67hpbiJ0/HZzRxm0Lubr1rvgMdoKzc1L7EmvsVljyM4CXX8SdnIs2K//SbFpH4dvvGi
ON2XDynRUmD0x+/hHaTe0RTj7MZBb4WfLEXlAEtbD30yzAYklKcsVxhOGEKbLE5vwMTBKOTd+Im2
W1P6A2R7PukpVIVNfBuBrU9G0SpCxu5MmRGo7xDZk7xWq6MuAPLD+y6sllV8NR5R5PfclJTshhY0
1ku3696uaD8mq747P9SdhLUuQ9mAW+KncHhXo12u7VtjVR5x9qA5C1k8cODTGUv6EUNZlyKgmJeB
xnKKmNpwX5R6HjSQaXrZfLZT/917yvp4rmdNxt/MJ8q0HrRfAPPzBZpV9hxdruVk2JOXCxTUdxWl
HgsrzvcytW1D4RWBkPt2ZPVaEvLRTW/HOHjnkue+nHSTBs0YtX57+zQLI7fDa+XBKWq9O4Lx4WHB
zXwvQlq0FrZEEz83czFckuDfp9fQc0sF1ZdEt4Mhio4Nryb1PfP5QuISuvQPa8ZoDg9uVw1B+uh0
q9mei7C1DOLfJEhoorxfVILKbu40NkMMbQtwEv6nKooWkVAJ8h/In3fcDiP2tVtFUX8gu3e0jGjq
s8xZ4c0/ExQYfuFhJdhkmNoOENkjNl2wGjngs/MOJskoVu/qcL+5oSTuIFipScK7/NywOSf+CEp8
4kFT0yxVb6wHkR2d1X5zaF3IXGjaiRJwmAfPMyJt+4h2BFc4n1CpBmTAzMbw9DQmXDtbyW93JpqM
7XmAW8SHyAG02SGcWehgqlIolKZ9PNCm+xqOkfrWsS4A/vj+yqA2eLPlZu1gWCymvlz7pw7u7y90
+1t86nE0ri32h4G/PZ45ko4xL1xEC8qkyGoCZbIget6tk7t3alIXwJoivDk6CdmfjmZEvfQdD6dW
0Yykes6RY33ovsmVtsLZyzuPO7oqy7p0jfOtp3UB7/u8/fewyoWGxwPougB77uoQs1NORXREkN83
na+11Go+EDnXkCbkBRMnD5S6kk+m2ILdyOwlASCxa+/exGYMfQ5Ly4knXceNu24l34zBjrsLm582
gmXm4v9byBJBi7spG/g0tex/gx2BTBmbh0mNv34WVJ7ZOTDETi+J4WxvF3RORtnV4+Lk124njE1Q
jMJntFsvfpxMQ0Cx1QcorsDmytHd1uoleTCRjlgCSovPAV1aCbsY7XjBAJtoycN55kwcBvKvGOEO
MZQohuCCYnyBGtxv0inqPY9ajGL0ro3jzFDeVLnAjbNnhA5c4aaxnDSDIxzZUcUabdokFF5qs8h8
D8295UH95UJ3I5Rj563q/ETlPv1rPIbRAdSe7IGuHEtxa7jIkxWRr/yrHZG2iH8MtnirFYhQ8K33
p1ROCt+hRbRs4Y1z3SQlsFYZSfLHywCFQXUFYJyOH1GBMGsWn/wcI3Xw6Pq/prsCsa91bX8RTBn1
CpSsSs0YnoLi11KdWEkhlOL8uDTrpoyDfUaxqQavOTLoLfPMpQAmYZXR9hS0LQGPZ+W1+Ja+63N+
fMtNR2XH56uuWx2WXgfSsv7ycQtjnFbAbQzJucYa08pwZHKy7FohxI15UnhYKfrm4WlJFU34PLmt
ZNd5WAqkpPHgEsyQTb7A6QruZcyzkz00ObZwcpbDE0iALN35H6R1F4ETGCFtQmVPatIg7F0urJJe
BoB/oKATVL5bzFMM2i1Z3l2bc7qP8fl6Edf7uhBICzMSk5fuOxlo4PLff8gd2ZFupQlOgK/e+SrM
JhHTcnA5opH0UqeMBb1WoFgw0g2tQFj0f2mtN2iP5mab5Jy6Yotf7jGXkktQQOxHY84wHoe8Ag1b
ZH7M8Sc83+5Wei87a6N+aYphocYo2aN9uM4XfDvFqfXyERxTGn3C8qF0l6KJLugVS7P2YvgP9pVr
L1l98QAUgMdTDqd6AXP+G5aB118W8YkIbIn+rGUAWDKsBov9mPDfX/HdQXHWPSkUmfchmBs04m00
E77OEdhSerBm9wuiVqEgOSFQErFthjM71GZztsi/bOTr4P9IabBPlXvFmC0TCucd8dKDmXpOmtfn
NzvXRq1/3FVKgufHmcIr1uYy/Z77RJxjhas9fpLUiJV6c5WlM9rGk3zOSF2SSv/VknaRtTUpwmgc
rGf4hRCXQ6Hu9bqD9gnGPUPTUArlhNFYFcfYA0FC13Z6kSClFhDweZRUZFsbPMbNKWEd0ryi5wNi
RDCsTgpufRH0FZlLbaPrxtRH4qZXo+O14sqgA0ccxf5MHvRLjC4XCthlptvEY6K5TZGGrQiJmxaR
UHeUN1ZgB95oCgB/ztbi/KhKwskUVDxpqb3anEmrLO6V//Ow2AcvncfKICx20NKFnOidlcFnuvt/
OU4dT3Om837LuYohi7Lg8dj2tMDkMZINW0HQ7w51ilVWlIuJNISM6rU5dqWEQ0tL4N7wHu+J1LlC
Wu81q5B1WJHPz/xPxpbe9GB31rVqmdC3qIUlj30JqB4o55FDPyOb8OgZiDKYc1EBGgIbZVY/fftW
Y8yakWVHyP33ErnQKt+7s6ts1UiK9gcETyafHG8FXandG6Gx0uWsDCPrRsjMXYFaFJjr+ctAVYm8
J0eH6DQNzqTx/o56C6Y9BDsst9RYjMdhFDR4r7QMAtGOIjkSKuDXjW6q3Bx3kiOwMpQwguUySNTL
rzB3WDDC4byDgO9IxclWRsbzOliyFPHWI3V4aPdJutI39inoh0o9LE1eR+7ewEwsOHKChl7cUZpF
+CXrPFRijd1a7FJjl9G5nt3heoLMlHtfIeyI0BvdW3GW/viZWhrjNkao1o6Me+CuKN1jcX6FKZIf
LNRfAWxYfdDWV5/t3hoR9WJbMo0F6UGy2ZyHD7nkTPeHt3aKNYGhZmwTseTA2FtE5UZ63GOrVFOK
Vdcy0AdP0GwhfYtLCn+JBs0kvpkC3Yvku3PRAnMsjrv6O15kR8+7TMTxEntla6GoACJvn+1sdTve
q7R+Nu0WuKlOTPiuymUuo3bHOl9EFsK04Xk8idSwVxiNXf10ZfVlo8fsdwv+OPJWqNxkMzoP7Q1n
EUUJBer9pV1cL031oCGL5iLoet2C49UpS16YM9V/xNi305Nq33freVxbl4RLA9FgAqJ6kl0VC3T5
/tcAffGXJXHM9S2zKXuy7VIkyr0M1UjnANaI0AvhT5dzB3HnnPRzsOfmWUawrcvtLLI0iwN/MEPN
uL0c/W8YGPRs5Zwm4qwwdeMD9QGO5n5CH11M7bRGBqfxbDwh8zoSEBwnDT4j4HUlsv3EY9XV/bXP
BLvChqmuCmDj3w1iEIAiTwHMvbXHTfHQJewK4jSTU+a7a7z+TITQ5oKfG4Wf/2orlSxDdnxBA9oj
BZeRhW3y7vlJdVnsfnnkPStHRwDEgrixy7Lm9+QcPxDiY6XHvsirA6oNT9W3L0rW+puuQnnrUs+Y
Y9cFdwZ9H3bcaknZeSlgJP45PinkB9vyxKyYRYHQ6aek5yqf5+QEJT4C/FgRqWy0Ysh9AGB0KmV8
i+jtPA4/CLlBtkV1jJvjELK9K1aSoQCNjiLpbJGvIZHgtaOzqRiEaev737176BEXMUB7rMOgw89c
5NG1PuSGkk5ns39aR/rwPvHLAtmYfA6iyWp2G/88bygBqv6rqLcCrs2hiXJvH91OYDWOZ+qjPYII
dtLMl1AMDh0WshQpQA4LBJkOSQJNBRPxNOXWiB6yAF2n5LzGkHUpV0gZr65H8Jbuuxy7DSJv9cDU
/0+GN7H1tojKDq5SQ8eanHqgHFyzUz5iCFGLgMAd2sEkj14K+/kvXZPtBRIaoZvwpwSc5wC6fwDb
lgAsUby9+zKZtsv1EaKDC66h7kR5a8dgHuZBR76Md6IVV/I7VNlMphnSg6WKeelOxIooG30Wbwzv
9J6lO1tXcbH2buWagDVogP1dLrqtTzvgPZ2Y3GJv+LphPR+41qyjVbAuBtRoRDo1L7CfDxn3ieI3
sbsG0MPht4teKCnLxYT/8f+ybGYGr67B7lWYYa14T0rZ3R8Hr34PLU/IyHkwMErZ8Cq7tB+zgqnk
EXsn9/Y/0GWGAdXXVTfXUg95PWd8xtYNHwp32lcu7KIk22y8DKVlgJDiYfwVyYhPiL+NcKlKm659
+KEFLcjsSbKN8bHoddYlvaQJ+pfEiokto8S3dZCBzP94CabFunZAhzRRB+ijOIG4WMmY57yWlwB4
ZEqEI4Sd8QXrf1pBsYnsMvb3OA4zcI2Kb6Xr6EwOSuaAwBm9zarzlUMy0QZAGnKLzBCXzQ813NQE
R2Z/04K5qlPWMM0b9ZLyfxKV/t3H55U6bJ5QjptkcW+nCbxwnkH598aebF4EjBOaYlxi4dylTSCd
fBKcEC+cOzMBVqNCz1tyfHQ8JfkRlEUjUwDqbY029g+K5WM05yYe5XJfEKNOETfijHhWI+n4+dRi
kFGdokeowKiNiI+C536QkBoZdZQMezHADyYK5msC3koPKc5vdyAtRRUpMW3gEbY+4d4wv2vFKxWs
QYoU23x9bIvp8qntKwBazNbAZXjM1nYEk3lXnTNbRdPiaG8sC65jhLmxhe5oP3l7aQGaRAFlntM8
p42juhTPzygTxOLdmwmFcgko6vuzrjrH3icMxc+ly5ljteodYotgCQmHfN4dmpvF9/F8EQJHxiov
WSWyJpLPnlZ3n8Il7cXFLy6NglVFyKPZGOaTWNwGRLtEj638iFKnllaIGq/PLLhHbGkWcyTL4Pvm
SBY8QP7X4GMx2hC6u03NGyqi65rejn5Kb/1qI0nfKgMQrmk+Cg1heocKB+QVkEzx0dS8Xpb4nNiY
DwGmW9TrJhfpexR+udTvYzBkUTsWDBquKiDGWotUfaHRX0dmAESRcVdqDLIYzUGRBucEJDTuWCe9
lcNBfUvXn1rxDmuh6R36P27/+zni6AtT/hbv1/y4VHcwVuFkwfNdaJkvHc3tiM+AxsCfrBlP4y2C
RTJBRHLmgPMX4Hs67/XN5JelAymKfvWeJ6zsewqbzFbbg7zd/95a4obkUJMRvNIu5wjVnlaVWZ20
eu/gQSMSTkFxLcE8jHESBNt4TUDjXEZn7LJ2SxyQX1Q+79taAnMk8fAd7TFOod/bLY4wjtuT9lpt
TKsOQNbnX3BLrYc3FHuPT2tqvHkt5tCiEBTdlc/1aHvcgQvlU3k7fR5ZbuxkgW+wlG6FBqvBgI0b
VF4LP4n7AqGqeV66CQmxOer4dcpvFxBWTxceZDNwE/fl76+dcmeqt6yjl7wRwbQ/06S15PJWZHGl
xssrqLLh79ibJG4IaYOFL8opXbb0T/UAI6PgrRzgXuMIBknHyg45vKMYi4dZ6EA2kX81I4E7LxHT
JC9pTRXcvHR3+TtTfyqfce5OHLmkSli+3B4nGrzZ5RC3b8Og5nbfalpj2iingHtqZl/UbsVQ1INc
ilL+o5jXVN0sz4kiQmS8eCfWFipdLjvKkxtMkosnZDfloh+9qZTjg3ShdmuAVgBzPw+548ywKLT+
Q9Uf++WnPYyU6HDWhYuXkUrHoxAHKAgdq8+VIhPe2AbPiaNpGx8xeQu08ilZqXwNQaGsukkM4pd7
Owe0Nbd271TkrvGdtTmUWJrpWog3yVxC655CcK8Y3Jtp3KZHEOPCm3yTcVVcQDXy/OOeShpaGNfl
cEM+T7hKIEUMEgxqn6a95ZxnBbQ4jPauyVnbQzV3POjxgBeb3npQka+6Jrz33I23b7WcdMtiyC+9
J6USNMk4RzoU3URyZx3ITmg6nQ8WTTing0kfbcVHry4Hq7D3N7X41EUCLavfsWZV52BgewmZc/a8
vnO7Ui2tpKUS8naKqGydVt+dvsQRJza0k1IdSdK+ycj0DivHOhVXxljfF7jsVjhhM3flr5fDvvxW
fatnxjxgvhyFpyxDEx3WizTegaNE4lifvhZvvtvg4006UsyPWSpGbfGS1gbXxmDC286henchbMMj
appCxBHawWCT8R9phLZuT3WrFRIUIVVwii/xqurxtvDqD2+Fj2jsj4tezuTyKGsWUQxy8ISZ4inr
vS0f+jZal+pxpV8C4BrGYVHgHsRR+bVcTXRM+jX3qH6QZyogvkvkd3WXV68tewKLYOsiOpx5oVC0
9NWNypGAgoBFCoDc7snRZT8eXKWsRE6U7yFutanUd9Ry8lg1FqRHvh5+ZsM5XcoeQxApnhdaBH3w
7MJQ9DoMIZec9g4uY8Mymb64FyMan4nmYDjddEzVaOzv5z3mAWX2RA6Nd7UfR4/nzn2K1sx7L7E0
DSG6+M5dMVMydL9eqfZbTR+V0it2YuVG+0RvuYbNkWJ8IZJ/Z6/3BUFXeGenrfTzSHTMBquRXn4z
AZon1Xeaxji1bfGIqaByZP9xp6WqhiJODfjgTyk60ApQXS2kBPcn0AwmpUP5OEZdH3LQhhz38VMr
4lHKO+8Zem+Kpe/YaDDLBy14BvuwoLgutU4GfGc80RWsd4mvN5cXhGmNfnL3zHGKAiJIqKpR3RyI
S2SnbYyFFbCZhsR7/hriup/v9+vIleqVAemhpXKNJ/dpXDoPQI8TSOtPR3hAfgAf9Fno2xZXPscM
CmNHoPyf0oBQ+KSZ8MJ3vB8Dk+mk5LVXbzg1xxEED0Lt0X5xi7hHkLSzNdJ8wFEjItVev0/xIHuW
pfXIAh905Wzh+y5SCm/e4zYh1RRLRTUQCjENad2Mm37cUuGWAaQz1Hn5kZFh4ik6OMbqwYgETfeg
msQYlcZhYEX1lLYrkKtqW0cIQ3ikI4NkaYHPR9iQpy6ON5jjdPww+357jjIti51+g7UlvWwCVw+8
uHmrBzCae9E7nGGZmULhiWZ5fW5njdA93OV+JVTVvg19v2HlaY1W+D5lHm7lL5cCUTbN9QBnXmnw
LfEIMJSTfA1oP6YDexMSGb9i7ChtsuwabuCWOPzrFbg+d4FCD9TRTppCaXd9sGAaPiQPSl+hVYhI
DPI2+ZohlGCvk5DrcYmWXcJKtLZsnr0DFORAhLpLVhbu/Eoc241WHlD0DUP/k24ipdaWaq8VrjD2
+Uyu3OFKYRNg4kSF0X2tOX2K2seMYzucb8hNRLJFJ0lw3iXoIWKESTd4tjbUGeWfOeoY5Xfscd6D
mRrmCf7q4KIim6fwRvzah3at17hrfVZjjdrDWEcMUoZrUUA1AqZnfyBlAxcP0DR8Rx1LicK2g5Og
FnS9JA5fOtpY3s1VwGwv4aAZQahROtZMZQixmyEVsz5+E6Tbzo7WlQrz6xHnVkoVDbehKGVfq8oR
xzca8/EdrDH07WKvKQwyWAYgbyO1PxtFtZJfaDQnpkVHMk7/szzobuDvq+O3sN8zAHk8gXNaexB8
UKo/Hnq4Kb/6Zkt79KwtxolwJZmDHFebmCDRKZFKX+dyu5MfWpGjsHqb2YSGIHpSxojyCEuldYzB
Jh/lHVLEBaS7Dk61GjwyRkTNxLiQfGM2rxCG2bxftgsWj4V1o4/exrZrKzhlzlwXdfVloqAw5Ax/
6BDdwUGreGSiSWKZPPqTCF0fCiZOXBuxv3naDivltqkBGbACjH1d+brH0+UoMkHfXm6ad1u0hkNR
GwLxhAqlQ8qmFrITOTUbKQ+uCchTHXpkhisEiDVUdwuM0bCIrRqaF9LFPYa8TzpWsUVES4PB+CnI
njeu1TUyRfuh3p8GDRtlp0L5hb4CIAnZLfDG+xwdKAn4NEziT+t4CUkmeeW+fzY+KUfSNxUB+mgC
F7FxsvyVi1eZ33BfvLEnvs2bBd7VhoAeImS/Inih5YW2/i5zzzIBvqsmaI9jvApuprqpl+OQDVz/
VwYxbWQL2HIIzkqBMAcpTaMhYnW9CppG8ESJBoJxMy5qohJ+8oFsBKzFJYdboig2qtU2kTSvWYRQ
B2icC4sgKjyGlYsxhFymnIVA8MFGhD7zDwlXRSTzyrYI2rMktxeHwOq1FZ8UNFbyQ0E06ISFFM6M
O8XUaZihRpG/V/j8b7l7O0K6UUVgsXG9QJFBP996GdeGA/XCrFG/Wj7Fx3YQrxVycX7gDp3zb+2F
VhMzmjAjmtW7woaRUj6aTJqMeeUFgD0ip5E63U8IHfkHTH/PJlrxb5LRFTGLe93/fLNkSd/WvKxg
EurfgXw86RWiyfIO/boUC6G24O8XW7izjLZ+Vi85ArMGgqARPVn1A0V24g5UREJc+cs4GcdaO9KF
pUibIrtTPjtdpgy5/Gn0S2SIF2BwX5QveIWcg8/AdObHg9rVXuQFs23DBitSinMStqsIdck0Rqrb
Udz+r/P3SzFu32pTUTMSRnY5/UprEb/GveiFap1DtvIMAbxDU/GzwGFogmAOrQgkyR7M7HnsXlK/
TCkvPC1Q3b3mfjJvTeBT9II/42QZIyhym4q0aXAkozKXeGBQMyn7/vjAfUcNVOSLyP15u7Xz1/No
AKYqrkJ0F/LCaNcFCQOBY0vMfzsQyZqgLaIFN0PjZ3RFtbvOrjf9HynbJsAd/hDsUsOwAPcNHw6w
VsPrPlPcNh0Hz7qVblEhC5ydA3cOkdhsIiF3cJyYz6DgTCV0kaN4ej1y3qM39kP62VIJCnBFRVgb
CU3npFcFDG0lAzE1rf8+miUvpYLIlZe+G88m+ndSKkMiI2jWLbP7bYEsDZbWBa91/gs0rlBpix6Q
dDQLwtdqzI/JGbka4SwrurQg3ClgoTh9PbpZC6t+YD8EFNWqjJDxv0NMkcf2wIY6rlbikRitbpDm
8ZQVqGa/+yrc2wAfSX88UcVoVG8CeBEUrkua8Z5Jpr7pbrhIU4BQX2r+ZGj5m7bNEKCeKnbaNst6
Hz/NR0Q1rz/jfawx160m7APR2+GC2wDiGDTDQaZukcheIYLNQwRQwh43nJW0uN3uLUUK6N+YMMIB
i/XgAdXZgz3NNaGoGlo1ZxcZ8KUYadtk6NF+x44XsB3BYE69huldqB+COArRJvQ0vCVyjk7g6APT
sZn2cMdffYb957ZYAtcKfnu6YBym0sHTyhKuyVReqr3GYmlIFmg4+srBHokMcbeCSR4850o4uayV
VnKu9o3Ya3ue9yGFaAthEhhs2mnar0pKoPYAjaTaaAXgz4r0ODta+BVRBZvvhK7cCyikZNAO+d7u
9GxIT1Tr6c8cLTQbxZ3ZTSsk4nmAFUSoaK5jwcWPlvTvJuTXQzq6R/sZARncyA9TQ0FMc6D9uE/j
yxQkafBPzUWdJ3WqQfvIW5tBvxgF8Iq9VdhI22rbb+F4fyC0KNtVkH0Ge+E19bLmZy+jhfSZFiN3
4t9C9TJXxz4wVwvFhkn/oh4PMFCxvXnYF73tZEoTKHzSFrWJDASOJKd5OnMKN2EVlwUTLBAxFrro
dILRyaEoHBv8g+yS0/Q8ymTgUQUFIPwrQv683WGS7hXNf8cTRlLPKBrR1noHJQTXTLA1EUqtZsiZ
2VvlcZ3nesP9LFy8Ez6W2y6QbNqPVF0KFMS+jpwhC4wwPs/vqDCYPnJg/hzGeOcH80RB2C6eFi7H
KvrCl+NDaBXHwk0+SxhKgeSHyOyoFf+jMWxwdA6NQ9XJ/CYPVBVKV4JBcR2ICnW75dHV7Zl/syhp
NRs2imWbAG83gqNP7pqfKeQEc/MykJFtDA5gw6jGCJ7MsdXuAJGk2rzEd37Ymz5rviEDfpJ6HbNz
imTGvUuVLiMWOWnFQf88GYkCczybG6UllchKalKtvWOMQ0icbKPAfhIViVckKC3voOCbu/gkiqEm
wdTwbzYixAswkxSLMIpI3nExktVuUTMHxjmiXJWCuZK50HF2gXGRF711Xf713sSyXzzzNTtTpP63
jFbNiqd7EHe/Ig5TQhsFEZj8E7OHWh4RPizZbExqQj4tbqD5rccRF7shyg7oeEM/3X+wP4QN7loN
6x2ocAvEgrdGOQ5pzxegtaXwJfrTKTKS+x27K9mp0J2dfwXJp3ikR8/cgN9yll1TkCiCTQ1iFZQu
fvhiNrBvjrCB2Lns+B9VvUsbh1ythfeWWws0SuGEpHm3EMkcWtjkaB6kKpS3iUSM5/ggJ6vj+5zh
zuuwdy9jj29CcFfSdov9nHUWDRo18y3y7pGdrpij3t2ko0NCaOQ8FLnfZjNs4DL1vuK+pi+niq/G
D5IFWhiPBuNGAF7yYdSOHtIuD7CO7KQQt87WknkFEX5kxKSeRj+DRQztVLmQWGWaIW1jPU+tDKlZ
249/IvFld74H+WzcQOUjbFUZ+sw+uif2ObMysnw1pq3qBn+Yf7HgAjbtOGAnwZ4bxesAud8hmt0Q
GxkBnCZAmYY4DQnxppWfW019H/OmYdAmIsJNQRW17pPWCtuTFq9oqCejJZK8cdQ2mBfziscrAZ/r
UL8wUzT07xTKvGxLLHkBABXGLHQHGgolka6OCYu0/ZwGRmYetXDA6OEZp/kdvhkdtqPV60mUug7F
h3L4wFVjfLpi8jmT/sns+57PVlbMxHtJpU7cI8A5hbLmGO9mHqmtbUQe41qlDSiiSix2W0iWpQFR
7O4WOcw4lTTcVfECOWksUTFpZvyiAps6D08xJKZJgaT9vPXT8X5igtffuek0oZB0S+aE+Ox2D+bK
048AXp395cXlBvtFzri+i4hcduZHYsL5SVYMuaxntkDT1+hHuukC+d24wMnDYCDsGnotX7SDMOtB
w+BctmaXTPNF5zOMvUwQWqB5wpc9jgDByluj9aiEn7BaAGZMDma4KfyM/y1QkjKM2ISNtjiDjQEF
igHNos5/DetbgPm+G9v0s40U6iVwLRSZiqt/xiIiV1df+FT/txbmFh0IaWhKE+4xgqPukmksf3eN
wt6KaH5+EJn9sMIsWjchiH/qoOMUv/bit71/dRO3ENTUkqfC/bsVlqCMbACoV9L4QSck1Y704WMJ
vtRp8XLJPBwOfAv70f2Q7XMMLAx+oF8Q6uC+GV1pXRhL6v9aB/bkUKISI3kH1RY+IUanes3evRlC
91huHEjMxdvcwYa/V07z0nmcbj3rqQHL7gaAOF/gYa2BvgGxX74smZC8nmjmOiD/ousPW3tLY3Wy
3u0gWnRjWOVZWW9wlc53IPZExrMeEPpzgpXEvZpN/TrzRJDgEiLy3sEsBk4UMwGTCBhhFEQn6oWP
N2xa1vaF3WaWhGG5mJxv0QMW7nVvfztgoghkf0s/s/shbz9CtzYMnXzfvXc2Bq9y9fDbyGLHvXT3
AUlaFfYjMfQw4SeT2MhBh5rg2GYd+1SMyPTMuT9NCnypMwKrMuGUzdO7be/qQDekuzaLHnVr0tL1
+oo9GRF31Hlt9OM6/rShuuR5j7+jFLRc29o6K+OsVeL11Kuq93pM+5HWUt0MEu/BYrd706S1rqV7
9HIJYjqnZSmYHd2tutYbV7eJxGEKHN7QDflLJGRJKUe5ZDbazEmRXOC8yMK2wixaxadgwkCCikQu
EH+gR3+9IKZ/5jt4+n0ATTOQ00QWZFvrkmROOyVmyiIFLJq+Yr+Lz8rj0yLcEPhoF8e8bwqOT3hT
NoZOIdLVpFj8rKkRiILbGy0W0BhI/w9GNwUi2W4Z6K3qIQ/W20a1+MrMkj5vlABDfizV86dzdDra
9089ffQZEjF27B7kM6SjSq+drCyhJQ3Ts55n2LkItxlRZlZByreYY3e+Mf//TadF2SQqx+BxFspn
ZKc2AkDRC62kLD3zcjwa+cQeAaQ+H9Z4zr5y/PWPOyJfyN3BdAyCz7EU2U6VEeJ6wybVaESbLpQj
k7fteXW+n/z4e0/9H5O72GBJne6A/ARY7dG83vVdOpCHpYaZs7UbDYBmPF9DtrKhNFnod3cM3Itf
osWnT5J75F2NHTfcHdY4/l/DkvleITERw9RaantyiWUoGqu2CXJc0sbBhEUaPt31LIpHqWJqrkFR
s+S5Pq/+WOvQTLcjO/nJqNSv/zSBuHK4du1IPKCP8uYiTzL+6Hew/DsA5xeCkK+Pmx70BKZ7qsNg
hxIa7WYYmweCRgxm4q33s6bFPwzmkP3LUgOY2oavKx1mctWIAd4dQTbtukIlib1pSJZ1dKVdSnsX
XPiCPo4QiKxLZSwZKYwtEcFt/uJF9nodcFImKHkQ+xQTT9yvWb8hrq/LOCQARDD7l15Hn3OlmiEh
bghEEHHtgSckhMofsw4Yvq4UMmSlwMFZvL17/BC0PzHUm/3a8JBaJkMGmzdfjTiBKGiUYtCPz6sO
ElQbq/LWVXbe0RYOy4+Kc/4YSNXpmJ0cZgbdrWk6lZ5MwTKk7TV6DAQUk0bMPo/jS72sOQ70BgMr
2+G75H7eHR41vuTcHqizg/s3JQuy/Sz3jdP1i9qLRL0mBm06KuYZpWW4TWcBHZRJBlXPlPR95ysx
wqogpJ+7LIna/r7wq7yJP8SJSicw8BlgNrvfybWqjk1Ff0Mc8NRNJvRuG2CNpFdYD28VCScpRwOR
P2c/W9r0TLBlllhzV3TjVsXIFzth9B87Y/+16XdQ1wl7UVOyFHil0rQRqiRIMTGorAudMQzXsqRi
52Mrb7TZ8Q+xM64mEPNBWuXeRwWGhyeMwVLXdttT8yUytOB+ttcgWZr8nM64oCcGPs+dsEuUDTxO
p5QQAhMtcQhKwvv+G3KGo3p+p53v4j06IAvFicClK6J4C1NiiByEIj9sBS02aDvnlfKEiFzxGO39
FI4ROFiaooAvgwQsf0cyMDgBGLE5tTn13OsDpiYz3JzQMg50WD/yKkBO2FvW4vNriMhksoWpZN1V
pIHMAHfwHovQ1Q9NfwLnzg4dIUZuftJyC8xcmsI/AyapKFC08CBEku94Rg2VdOKZpCES4zKaZGDB
3b4keA/BYSsXlpm1UfG6e1aLcp3eRAg5LbuZH2NoLB5zDD3qvd7fn1Qj26PNiwXi6JJXFmVWLXie
Np4SaqpkvNxS5aSC4Kg2pe5Ezq1LgKruZYPy839sfhuWwNSXF4oWHk37NwxYAkgb9ifyP7OeoQB/
d9nxE6oN3MDNoyfJSndoa+ariXMLvQSb9Oy/K9UyEXaJ1I1yJC0L+g6FiUTmLwAaIBf70HKDHn/X
JIGklo1OzFyLG5IL5YhFESARoh+voCG/y7EQ+huRp20NPaNXuTT2jacupKqIbuyvgQD/R84qjB+D
u1dLhx/OghxkMxICVroYRpkwMqe1nIa8gUtJZy1s9iyrT1jYkElOLYY0SqaQR7AQHlPCAg4T0BEm
ZSHntp9R0W7M3N0kVKX0PXKXWVQ0nSK4uyZIpNAsAW0CT1LZGDcq60P9ApAlBqqwkKfFf+0vas+U
qt6jZjeCn92fLwMGDDnHvzkejZv36Pk9ELdCxtJNdiqyEUy7KSR0A6rCaPAwEmEMHTuI5v5NcWO+
jJSbf34XISCZTTHAB2fV9yHR9BN2NUo83AcNTj6jHezY8A9ypIDiEseQI/wppTUw3GQo8YLuRzPD
9H2V9V3ejA77PMIrYE2snqZ71v6UlS0VlKCTPpJ/PQOiILC4YamnhQS7uLAGyTTQKMyIzzIyEjCX
Ngrz/FBfwID5k9k43NZKogxst8oK6N8Ds3TveHCAmJzSoUblivBk3Azv7/GjT69FjbmOEDUEhmfq
+WgE6R9Qgvd5wpgskfgluwSeg1oDWiEYONvbm26ZAKA5ABZS58oQmFKEJoUFQiimGQmdB4FcKcqF
VGH2EXIHNP/FK/5XFhW1N9XYT4ab4f6o6kSPQLyZ0dyzTC08XdYZ1ZVRr8kgPK9kZoreUxXu1Hbi
Y7elrQa7h7G8EeqoORcQ3pwAtHgUc/P783IUQ01LZZzfjFRZP8J61QzXUYsL5kctXon6r9F+0CoJ
WWGVI7AEroRWtl4N8g5fHYcSxJBNg+6mbXKHh4snMjIl+JjhDfEbq8q5S25Vo/78nXm9I+s29owR
FXqX9rNYVu0XFoVfyUm3cGGwhSYrwnT7CrLRbuqTKwaE12EHCCqS00Xgc8x3XL2XvVOAgBST0yFi
Lm108eSyGG77QRYQsLqcaBdAYkOQ/t/nMTA5UGCqY07BNhJd2nTEUEt6bcTQ6shpQO8eWXEzSsV5
pl3/s3D4GAcK+nK5Z1ZqWJArjUi8xO/8ZH9zG8DI21E8RZm1NZHNqqEuTVSBD7MBCtziCuRqnGfb
0Xqsuc4E5+4skBPXv2m6Wm1NR3pE81Y6Qagz/8OzYkzgii8xaQ5R5uy9934zcbL4VuteYBIredEZ
cQvsPeXJXdPBlKnu8lBchF2AYBVzvD1aDTJoQwYwOgOoLJ5itieqE97higzTiTNZJHWXh/V/pIzZ
d4uKpJn2FHKhO/y32kuR4fmODBpVSnP5yo0r6wofnxPwDr+PVJim4OnPCl/QnPie+stWrtht18K9
iY53XKPy3E4u/9Gc2swjo86aNrsFFVio/JOQjTyPsF0ByrFC3F1IzswDY/k/ojGKsrY55pCT5VbJ
6ekxuJbNTUJ7UZ3PM0rZrWtehld/LEiDic0SbHnKlXL88daIi4t3zK1u8FrxeVoN/6XNxQLumBmI
tZ/zYopTvUe4ZS1vgs690EsK0twYXbR0EKMkmIxgwzZDmWzP6ZXNhgvB79baLmJdlkNdN2L0g57j
nJyVJk31FDnz72lHg2QnyEU+jFsjtxSe1SecqIzYlQ7PQ2vk5dvdVYnB5kIZlWlyqiHCCPt37BCN
7uflPf0l54D2hdJrJ5nm7AZ3M9/QSP8PNEFjrvLlE7S/EJLLPcozPaQz8YIQ8xF5m3X9wqRmQovn
EHzORVg5wtD8SH3xLnjvE+WxO82zpprvL/aUKM0Eqzwu4iqbGBRLrMWmeTV6K86fCA9snVDEa2pY
7b5BzEQZ3XHdF/xNQSqWDp7KU4j1dZhuK1SFgbd+fGWL1tk7ZOQWdVdx5VVFXxiOfCo9m136C4fk
clQphWZRTEmNQG4JzhSoWZCcaT8r0EdYg5ZpUa6chz5ra5GOqAjWOiTcN73acXeug63EwxddVcrL
y5KvZ21ZkMnlDnQnMWjIFa85wAxNDJMZdl5haFlSBX97W2A0rq6IA+oReQ8T1gi0PKVQ6o2VjcE5
R1KU9r4K7RpwY+g+3ehsperzV0Yh6wXC/HqvwjHVY15WcuvZ54a6+fJ3QJbnymxiBEEK/iBrpleV
U4AAm0krB3yxE1xaCWq6k+BlngVe1T/zen/Oj5r+n1TD6zSKXvwhW6bcCRC0zwoxQXXWEGgLNPix
RcWSBlLQdILIPW7RhoJmN/3CZ7K7KCN2n4kc8ZJQLR3YGQR87elv4pkjykU2+1rl566y1jm0VFZZ
+LvGwfYs1J0T94JA/eIjjWhpTO2X0mlxQpIN7vcfCxcVRLs5AcXH85C70nSFFWJZlAcfB3nUHxzk
RwZUkONxjtlPd3cQyj1Wb4J1DQWYwyvWhMF2quqIPngxZfJ58e5g37QwWPaaSgLUPq7sT1mWfu6w
ViQ4JP4y9QhGEFASneuqaxZHQ+yqQTaAJs2wQufUD0+G62kxcGIJhkIvAxJyUFt2z+1DeDSoEV2c
dwJH9NkbwwjVXGbN9bDHrpFeQNTduzDvFSvwZcq1D1ZUgWYRK1Hsr89bCcL7KzfjccEMJNaHiBeH
LR8T4IM2ZkrccOcP9c67ZMo83Pro2e6WUv21bikV68TM2OQmMS+Szp/xxNM3pSitCkJF8/Q5XOaz
fWF0Hv37VzOvlFs6yExW1mJwLkIzZG8meDgSKqCgoRByfj97KPTxgahRsW6Qe2Uc+kfdqgbDMolr
9U6Tsf5eWOucdA5QGZ1tzXML6l2p7+MiF0KAe9RXWL90JruN+8MeYqAlQkCAjJH5Z6iReWvKIo/Q
XylxApT8oHtwyokVdPCN9uPAUxsnIj4/cUfAaz3XpMpv8gSwF4VLXnonevYxKnLA1DcMGcw/U8/B
/3bsxXg3ER+l9N+VQeWhyriZA4OkU2KKfnP1+j9SPfjo9g0SUW8OSY8ZtmzFLYozus9DUCg/Jmit
c2GNYqxU+YYmqnTlNNo4poBjidbXtC0Hgc9pwEO4TvsoAfSOlSwkoVYHz6/cecBUOGD5Xb4ILQwO
EC6kAkynH6yoB+oh332hx9Z1LO4FQhKBoTKYQqJFGtcFzJB/+DvmC6h5icr6uJFInrddGSBVbGo5
GbO5eEMD2xNxHmrfKdI/1AJ12tBXKNNPg9R/SOdDPI9F42MglbI8QgB1wc8MVpJyoGfkUb2m8Vvx
+jUy2UwWAfIe1I5J21teQFEm6QzRk6dKQMbry8w58ABXaYOOxu/QGH1r8gnvExPikSakWdeEA/jK
1uDPx34849w5j19/BMZHepyPML1bKUkiK4IVksPKyU0S0+QczqYnfl3obBkRk/Mq/RsFjnu2DiEQ
dM79ETirKp43bCvIKvGjXw3v1KirA09E+62iKx8p9Rlk0kEs4tXDnoN47EcUIapbeH5xScA647OL
kpt9lfnTp6kp5eKOJSFxSsESG7S+8gEg5k4NY7aTOnLqAQmZDf+2xLsuE4kgMAWge8X0k49QixpB
7Z4Y8Z8f0BzTrocTbDnlvyHT/WrjPkiPnfgLV9/7/AJ1QKxlM1zNfhPhT6S8r2BCMc/RTcXY8bcf
6DqG0QBEQV9VtQfVHvHBC6BpEaM3awcUQOyKYKVNS14aUT1WNv5iqt/P2KuUcBnF230IP/71HK99
FW4n2bL71EurV7oTSWwjvm9r3H+5DrEWSaPAatZXYpR8NdNp+bP6V/RZ6NBaVmnFHGrHn+HfVGVZ
pxHv/gWzOKeTtjKg79G9zqGJ12evZYh33FRUjcmSJuEirxoR6p9yWCmyfdRqOZn1xEi2eZxbLBMM
KhHzdnOl9XUSuvayvtXBMB43xMu2ElFz9SoiqR9oiiX0u2L7MpSRrs6CbvZiFyqb0LF+DX7UPY8c
IL9vpbyUUoCcLlPf3WVhRfQ35l2nmtCSIv088NyIhpTlST4zZBbzfl7dXVzK4hkGsfptEBjlL0i9
6npU4Ef+b0fEIYjvanHY9mMLjMwvq810HmQlnYbXkOa8PcWHkiyKeKycgD5Sy+hzGrKKcYaQsdbR
AZVsN+f8VKN1tvyCcNq+w2utKP5xD9pqUlO/ZfFD7niiIDDTR5bjVCdfKvmRaJ80OhW7yOes9NG5
9GF+d0UlHX/kSp2oeH65SgTto02Vyk1C2l0I/stlmQhbMPFxla1OqlsgiQWjdRJnkgM331Orrt7F
w3+L0VlpU247KSHXzKfK1VHyrqRxrHZVSwONGTroVeOsh1GQjYEcYx7avayNGYV26D9sS6jIf43M
urSs3wrifbVEaijVJhI9SMZBYxX7hhmemjJujDXotmMmDg+CsM++oNGY0T9QXEfrriq7LRZFh8Z7
1OE6X0JwsDRG6s1Sg392mwETbWb/GmSpWCxiABhFdUwHDvhltWlXc6SB3IfEVban+UQm5KP2Gvdq
jUMHdtZzfVj1pAKT7y1nLIicO4FAooKJCSTmluecyq4I4pyFBrpNWvQqYl+Ur6EsdwbWSekZp/kN
Cv/TTgeNzfNliJqHu3GKby7lJ7YOT22ReyC/uvo/8io/4yzzaqlB6cmmnZOFX9CHmS8q353zKyNl
RA63Pnnjd3ViwIisOwlK7G78FBp+jWj0eVBoKHiB0Pf1vcHMM7UVsma5vvf99il7kWe1B0Lin1DW
oQgF3ysbJ7Chc0UlURgOAGsOc7SJlxWW2irNkKUhLv9o1aFYwPYSNFkaIM+th/2BL9TWzat1X+mj
Nkf738RwMAkJ5qIShAk59YbpMcVFFeqoOEDkjwYa8SiA8CADt5u5iWDyToyBXtSYrIY2pTGbPR/J
qdWejyJzyDwrGZw4bG2sfiAukVrrGt8jRCGBN0FpsXeaihdRb4Sjoik3hdpQfb0CRK5Gqlmzwzdy
eUXcb9f1d2PJMKV7L2LRErmsNPNHKp5RfbPAmpjjl+Bt2sGmnjTQTyFdjRKQ5tpdJ/kxAq01WvZc
ZjO0i4mpz3qfD5badp21f7q1ELX0yh+BadX+iPcyRTa/DRt4bPCLUp0WoFzIRMR0e2pTWCJKfXn9
SQzeoJFnrGxbovPbeIHwreyfOzBj2vKcjPUy8piL3Og6LwnmDiQwsBWOQ5FgwR77Z5uWIDU4hKeW
CaoOIhV6kMjlAOTK7rZZqDJ2033Mhv5GTfq24Tu2lXzBTk+Lvbu4gXGTgTOzo0B8CmH30JxYr4gh
oGRpVq5X3MnoZitRjvXQ8CoR8nK6iWmiS3aPIRnsfUPi7OGPpQ3z7YtYgNnnRvn48cLqa3hb3GXA
YhfyNRvpP565KKH1sf940evnQ/Bx2jZifst9bxSe4jhgjsj62Rp8lX9AE/+3+aXRmzKP8UeVxr3M
G6TmLV9bO75XND7865DJG86sOUbTxG7xhK2k5C5orlwlMiVaZ0vk4D79B3esCgZS5fpUuq6sBqbY
bcMFfJNGHQ62oJ9sAhZCyxFM+A9KC4pJuDTGyRmDqIHXfSt9pD7+xo+FwsCPwAv4CTJvckQ1sNJv
D9Gyj0Bjs6ZjhpMZd3jXFk7oEmhgpzk059nPIP2/hjpCdJqgxjYTHJpbVZheZO5OSTE6f+yqqPII
8/CpS/Pwf3uQiptcaphE5UjWtHmTvTu5ecbDbEP7iiWUXPL3R4O+nKXNwomyXJxHfOLCZWFRTpaI
Ekiep9Zi5f+X/Bvg0d04rTBsVmGcpGNoKyFy6Rx1NsdXe0Gh1YX5oMozLsPYIrT02VOTMxShx47T
P852j6/AE8qUt7/U4s6csREznYyztPEfHCGFdPcQOjc6AyvUb04gVgsp4NX2uYk/3qCOtd9ss9OT
fx05fBBCCURmYm9hPGDvtcJDVYNOHlpzaxZJz3djsd6KChsgXJtEjB2RYP+P+n29ukGAkm+y7sEd
TXJeTPhivloWGLragKYYHswQDT0yM/MldMJxXNepBFmDZ5LcskLczWxRrlwf2TWSKN0yqHGGOHV5
DWkwNoazTtIyhbgs7dnFe8ako0V5FPsTQwHGU+b5NUa0L+Tx8jC7hEEQd8KCQ2vHSY1J3mCt5TGJ
JnlT+bVxckNY0V6fWfnbj6Uo+hdZenmdbHfE5hzqtl9/gYUuH/gPtZqknIJ7mybc7AnLCSsqljOe
BQC/V1IEpPeqPWgFyLMLFcO/DLBxka3YIV4V9S8HbZ6H2sLM02wfRaiGLXinfULtXPahcgTNNCrF
II9mWuknfHm6AE2i7JyVyf6KbTSseyoy0vM5et9VkDbmcb4RRNExwPCCh6co+swvL6gDvJomR6Kh
sRYrQA1RT+/ubYox+blnSJEOI6lw4pT1QHqP3qOY80In8Ye/x4EqH0ST0W7WObBmzRvac4K232KD
bCNF6jKZ6tvmYAKJJckvi35E6EPF3fs5M6fZMeycRqIuk1gXcJXRbhH66Y3xQmECNVXrGttsbLmC
311n0hWDSsxMOZZ5Rvdizyvnz0iip3DG//61FQ0Ni+HJopIUyy7IY4o+Ov8zMGTaZIEM1sRlCkpa
Gavq8LDZ1QNTr+GG63nKj9rDjrcO6Zjyf4VuV0fYWD3HCbX8dK75RBuGBjXk4/xyBkKZAz20/EdO
/GTkMI+9NiVwHzu8mQf334WkNldAh63rYDhTuRivCYphYrKAvY35j7/F3fiaXG+nrTypGM96jN1O
QfxioephdYZv8khFvdUAC8M7SAVlOzLEDQB9eq5gJatA9b7i9ge84E8kFcYs6M56Fgh/eUGkauTm
ZLI1Es+ct7zzCPqjBqwYjjqknwX1E7wFv4KB/whvNRJpYzgcVIl3K1eHy0qXsWdaut/xyQFRemyk
/mUuUinS+r7Xap/4KXNsIgJSxahL5VajcXJVuko2weon69Jzzo8jz6o0jA6oXPJdKa6lvBTAMcz6
GA9//5BXQ86uUc26DiKjTYYobeBoDzCpXbkhZ54N8R3Hg9HoARHzo89oLHup+mXulT2CYcLUKSHN
jH8PeZOGYcRVUpabeGmzn5tIwfhh38H3Nwrbu6zBR8XB9ljlL6l8I4klk7cb4+641SaAZq0gCqB0
MH/nFpPFmr5LDL+7R8bICojq0HwJtiqGawxv3kh7S47YE60WvXlH9dCkAzRgIUtVyg3NW3vOD3Hu
aR0gbjFZtPsBLkXHxwU7sC2NoxXnE8v4GJQuPvw2ze1SxqRbjH0gJp3r844C5RB/vu4vwxosOguI
gziNppCfhiEXSf3gMqoN7urWbaaHJYVzS1qHmp8ql+ObqgS0GPJjTGL4YOZ4rQHEvl9SHKi7r3k4
H9Yuw1oP5PNb29OnoiTjAzQ9VYP8IT6dcWPFDlGbHZ1IkocW7GPWXywjDluLvC/Z8ZBNKwe9+46m
4oPar+cLeUaYyi/0X2Rinsv0wPG0ut4Llvoy8v6PEC/C++lSx3j47zXGTtHLTozlYFztu3aBDSMY
SQcRX8w9aOFriS4VrrHBBODM9sMy5RMvfoU/e8YWjjp7XD+edBs6EgKeAbqsokB7JzzQ0MaYkni4
PUdDMWs9EoeMJMZ0uC0+sCNEFf9olQKHc9JXaZFTiEYhb39YTBOXY/6rbQdARKB2gDK6vdY3p3tS
pVmgGScDq2CkvNbnUarrYuB8nUHHQMbpWk77n7B9ET2XPo+6TcQH9GghFhNqNdBM3sHGGiKbFLYl
gRlDzgmAFKi+n6BBVmM7MLQXSZLwVUyDdbEr2C5M8Ht7arO8NrPXmwyUlX2fj4RUrhBN6pJaor2w
R4DK7vm2ic4sWYX5G15VK+vihFOVy+tMIWRbireHnoyJVrZr9apSp2D6Z59rFukX8BQh6VjsAR7J
ILU4r/WR0DImznVNKW9b/B57Imv/IPE/UTuMl2pFfPwwC7qvauEw9fPxdMtyloZV2tzECp6cJHCd
lDLYcMwQW6Us5N039NQKfV/I38qqSG1JS5W4ulRnlWqoI9HByeybfMDfBJOKU5AF1i+dFbn5FTb7
+asfbvc6nQE6pSNkXPvbnn8a43QRhVHon6rWT37KmGO8BwamSnVaTBrdi0ZeCNDKBsmMtHRfEWyl
OxzGfh4xMZhugQheGqW4qfuO5crQOUN+wVuYrsctJafeJPZtnDDf56esH5RVdgDRsxQ29QKhxxL4
RTxNJqHs29ds7ZNy0w7RcrEMVkpd1Gw1/kvLk3k9fFCJNxHnHzxaMJzUEGGX/+q4C/CWs1Gq6JRO
IIywIdXl+srRLA1yHqkGxgNgCjV5cJCPsek+S9Sk6oIrCJ2zabieigDHJgjO4veuex6/5k5plsYZ
/VE9cF9D5aPP4ZwpOex+sB1gEF99epTj7+o4+k39A+fCAAVxuubwTKdp7kwErvnTaIUVeah25ob3
k9sxbsAAKCgp52wnVnBGQV7StBY2PgWwIPqKI5S/yK2pApEx1mjWPN7yWjBQC5tswMNLeNJashP3
CR/9wsBr+2hhg+Y0lutqvtk/nmhNoAT9DbBoQktK5+s6DEvYGqW51tr8NkNgDPZ7v1wrn1whSkgs
kNTWf2j14liX6uMvUA7NSMbST6NAFOp6QewrD+DaUV7VTM/4RRe7B/0JU1kyyMNP7GuwWqnI47iq
QIGZu0s75QQkASAuTp8/0O5G5DsgrS3Mf0A9V4u201SpCfK5FpI4AU3orTFzdKnILCvda2lOSgAv
NYz/mQoaxfLfPha9Ib7hU0S6lZG7ZOqAxZR3N6jJhDjtR5iUGXsS23d/CX7Et+00KTrpNEqFny2S
IkiufotwAJkBaL9YefA71padBpY88MQ0Nb9yQ7h7TjTnlD7wbzSUXclSNguhff6nOC71AZ9qvClb
6zeTT5LmDxOxhuWsPTxxwJY8ZAOIo1n0rlneR78/IDvf2fTyJWrJfNzTL7KgFAjVKbqsZWsowOLB
3WkQN6+WxChKebZ7whC1Qkr+mVzeZ9hdD9TAIgV9te3Y8f1uBHzXgo++xwdpLVqBFpvjEblmHkHD
sOutoRH7pqcScJoMjBGSrSssmDioZbCdIwp4MWTOjn/H8utsyK68rQIn2kMnvtQ3fBqhCx3+PHA2
m46afxDBOEib+nLUnhV5ivBONBnt6SjLFMciZvNWhMpcNffLF2/7+0uI10Cn5fetxad9ralezoPy
qCBpURxl0qfAsDy8qkvfy1PmiNFC9q7CVJTuZShJIQUKJE4Nqgrxfy21HxmbPUZteX+5nRz2Q6kw
Hqhl8IuBO+HtqAidN+5tKzSXrdZTbP8FWxqk++dKb7fDetjR4KTwmbWqnuRyM8aADyTblCXydI6U
LG1FBlr31l2GmwPC8s+xGYjPtRcFneY27U7N+ESwesxFi9noaYWDf7k6A4fh//l+pMHaDaeEVANn
/Rs94BJxuICosLwju0s/sS9Xmf7UI8/NB02STjRkyzulAsLDaLzrxxRLLCJteQJJ86ecygXGtB2H
iR0d41Eaa8qhqQgAbHsJXIJP5tG/MsDr6CnkZaA6AUN8nRo2P1bs88+QLA0nDKC7MZ+MjcIR03Lv
bsogBi+QSMjJJeycbj0gkswv4aDJQz46dV+BME15we9sAe+pKirsIMsk4xrd81U2hj7og43ebEAL
iHkraFhpdra8HXmLLUne1ZHhgdTtvXvA/Gt/aWwsKbi6zYakP3Cefi+WQ8H21t9h97VqSWKunKxN
MWYwfewoI/YU1h2ThmZKjsx+YGvdPfrWvi888o2/9OIwcR8Ft8Cbq84ObrLW3ooaL2WosC2aDrgR
9UM0AGdZvrjn5uUJCMezLa+S1XZwHJ2x8xNghvlXzn2ZRhIHxgkl99oRYSTy6gNEXJOUlWp0VMQr
tHK5t6R1+kgUCDN5N669L+Ne4ixCVVq6cxVAeWFJ49SYbfjMTKUCljmfnPz5Q2VcaMYVUdCA6RDX
XKLvor2aW65aCfXrCVCr2O8zvzSftsJPeotAGxhC4vFXfc84gSOwgXLrpRhxIZmosBTkVWX7M0oy
oNOKXCSJiaXXp6EO2e5HdLhkmL3OjvHpx8/PpdtEruGuUe4n26Nc1uc4biCzpJk3cghG4Wqe8ILk
27VEBpjpWbOk+t2BUfzfXozqn7lnQGbCiIXa3aMfiERCJgDLwgSg2l8nZvSAnf8NBClhheR2Rowh
MdQc4QN6UBYal/BSujRQnv5fV09w6t2jjZv0rUm20SnsGSa5pVF05d++io5yanqfcrn4LD9J61Zk
eYWa5ndpwI+iMCq/gxuLF1FSC5d/tGfG+hh+8Cy0JYQkQYw6liZJbGDBDL0qalPwJj37YGAqYWL0
IUmj6M456b/0guAb1BxA//9iB8iBvgqErTyyOhcZFu2qQj9jGfS0zg7/s+ECusOOZ2iYAHTTsF9H
zYrEqrbZsJKf+xVHd+yHYLZ3hZ4XUf/Q/yCoJuG2AiR65KBj81g+k5VSVjjIvrxvEceNyxZPUKpe
zYSlmr/2jvY4o2GjFQQSkC+yg+z4J4UVaHvw5shibT2fl1nQ5pjD/oL9KtAppA/Isds9QxljxY/N
fDFxQvFVqS67qxFrnD8DCamKQSD0RtD0RmRR/do3+3bbhMWAtR3JqBQbM1+nRU/b6FsG+xlbNRhp
gZHEtHQfCwf273IcwVDDeezf/7vbHMC0RyyzmkC6uqMU4swadTUj1NZcUBGlCGh3QiYoTFQw/Ra1
Ux2R5pZ+qbUrH9CExZECvdIKgeDsKkTFnFxxyLXxKwQGFMyRQ0E0ssCq3UmzJ02qf9arfi1QX+lC
Xi7j0ylHzN/OPnAkJpMWftDOqdnT4ZIyNhNRtz2yvkxAQuDguVzMyktgh+TZcSZ9/NRaHwtVNDqL
Cm5nouAGnmZJ9ctSsQi0O2Sb1tqTf5aip5ckGV186bUYsmKtAYIoxjI1P00dT4NEiW31S2JBqRbt
9nxjXb62R/xryAdckKPuy2iY8ZVf3mxNm6C+8IrAoYOZHtq8llK9PYlW/cZAEYrzu93xlEPRhCZQ
c+zpgDj9HJmnp7NcO4BrUYNxr8UzDFRGLg5cefyVuLnJ6/bjJx1Pw6RVgLJY1O63EA8dFeqrWL9A
fDMqd0j5p/mLmOQr4yOLHKEQXDSAP9BCRyNud+UhXk57TtiRL2Pv5DXPcM+vjgaN0ypBLANmtyvq
v9fG2RQYpclEdU65Sct1nKObkHMjTVU3mcLVgwLFsvx5zqDXpeihVXH30W0FAlh4XgH+p7Ef7C0b
mzneHmPpZhGNFGsQozlOGMqZPFwsu2FlvZ6Rh0PHKkk+bvtdWKUV0yOYYFiUCAVkZaGtfgUxNRWo
j8zSHofQ23zrDi8k/TQEV/cnmuR/QcFVufL7M+MEU0+GeIOSlt08Z9Gis2XSza9gvRAs39bZeGAU
xYmBBF8qseI9MCKXxW9vx0IBAQL3HxmPadSQ6bH6Pj46J92eg/KI5H2dj3+l4AfSiPSWIb0zT0nZ
qVBQssuvuVOAb8GgQZvB89h87ire7WGmsRo8SIWMEGR5+w6VB1k1os0zLmyKaC2wBVOm9w7jhqqp
oI/rsXFEZAOjQq74ASSul5hKOQVbLZLyMIsgRFtl4Z0VAPmIZ6BDbV44RIZBMacYSnYpR9dTqGeD
fV6rQyz4Vj2UNHKVetj33BF394/G0eXo+2UgkdjPmZY7xbpeWTlpdaGDMYB3R8AzhlN8d9IXUj3d
JRqs6wGUGGk8x29YlXtMXfyQm0glDsS5FWHOqC9Lk/1zUGd7bZ+HC7r9239c8/mak66EhaLBDZA9
CUJz6OWA6P7K+a8XIEgBe56x1Sp8JEuTuOEcIYvclNgeZtgo8VMMniJrUWUfox4zXx8sYHi3Hba+
QKTTeTERQ6QsRM/ZD7pZ3rooSNWgGPvplO9N51OCWgXinCQvkXhEO5DuvF6U8SDneyqjWKFxu65J
GWuyabJ40RNgcp9MYKmvBoJFvt7PxD5aB/7WZbUDIT/AcFXngnEqHKU7vGQhquuSJECbP2SlCHQJ
NWFZChMKoi6CWZ7kS/33jZUx0SgDtGYNBYw1gBHUbHmzhCEUONmEa6vo+REyVP+Zl7+Gd9J7vBwe
vR/Kgtof+TGVqfU8ttAPCnQfOCYYFa7V+qdn4VsGJcH0w90CoZfDIMlx9WyO5rTD64qJyQfoJRhj
gTIJ+PiptD/V2afmcZ5T3NKsUHdvFytMbDxlBXa55QOLX3cBLv7FQy0aDKnDWEets7QniSfMk8lw
O9/xWyEuwfRNv+XNE4hTYGwTnIHSaoKBHgenkIad0eyTbB5uOiygZIrudcRv+l7uIPLTn5PaQs5X
dy1nE31qWvy3PxhCy+lvXUmyNz8J+gwQtrkyv2Awo/zL1w4kplTsLPCY+XNUEMI0BbqCtcT7oJlN
wkf1W2b3Hsr5wpt2wOdbN9jdQgz2imw0B85GckfPbYlU1XlMGTfexR9ZiskMH/3RCqFGGY0fwKnR
rTkYgejBycTM9dCV2IZiAGqVX8zHIsgRLgQu0jnJuwHr8uEDiGIAaeKKpwp1vdROcE+rhr8/UXul
XkEzEaFvQMDGFP9Xs3ulYCVCtymOz1izby+/5XUJEcK2k6JVvryL2sShn5xOx5EUaWQClb6xpKut
ZjD041seFrxY2G13hSWY5XSQfS32Vqa5wb9mlCxLsmAwANIke5FWNhhPBYDh/emhfm3dmM5tdRvk
JhwZI8/XG+Ar0jiYFYblcHslO2x8iwvaeeslTAahyPWFqA++pJffkKzzEfxBirbt7kpZYLzkpm6R
0UG07K5X6MySxZCbnFfa/gfWytnOBP+oc8H37WjI5BbreqxdjUT5kmIj2HcRTazlG9QOa0Bad/Nf
1doM9uFLzgv5k+xYjgl/oT25NIpeSUUPuUjA9LcnCiXlum7JKFRsGF8UlhzCc7Kbl6naRKTbmOWG
t6/nYMkEbYg9osRkWUzyG35/KIeoYI2y92zgVAtB5nhmBuNSb+b+RzaRsKK0S62WVI/0lQvD7Nzm
GiZJsv4yLoqiL/OuxYVd+RlwqIvCY6qWQtY4eOGdO+7IllgTseBBYdnQZUu7XX+R/HMyXKrIgFdU
I6BLBAH5ojuMg9TTHsfGs1LM/pspR3/QW3kD2l2+K773fHbcBLxGzZJBvocJYrHH3UnH6SLhNtNR
urbxL+anwu9DKdfAg1BJcySw/DQGG8X2Ml3s1SC3bg7wOOB1Vc/tXSaz+LXQ/d4F1qH2yKvAULHu
TTQ8CVBEbsMEbz0BR+4Kl00kTN44DSyyh2lf2HKaPkZvmI4z1ZlkQ0w2qNB0vQsynY8CcjHyHAgt
HrtdxOkaZfuES9q19kR+Fldu8f5RujcEnYqonYQapmtMm+HXpvZ53/sqRvAVMGdVjg6OkfjH2h2p
JDhVMnqoXTLC8FrQVfqFblfB5WL0MMoh48EgsXqmPx+OI//hKbKHzBVTfOZi79dBvCyLonLPxVgP
EApLqQH2Ma6UMgFB5s4XbLy3uR0gTUZ3K5Od5PQgdBE/1Ijn4aaep3GQLN8vWYsZHZtv67NSrtud
Njp+j4+4NoEkGMWwo71pOrVH2nGjK+9HIVUvCjpDQhbIzIBw5sm8xWvDCEk+fZZ4iTOT77yLv+1W
DgRrbqWtk8OnSw7DBsssB5wTbmKUOHYkOByRycqXXLG7K5mJ7fWOe1ZZcqvljvtmvSKFSwPhgz4r
8lN5zTOYgKRE6/ViF6RtVFKv+q13Bskrujd4PUICYxykt2HEUmT6WeX9NR/CmP8XWl8bhMYk3q+S
tKQBBaT8vXGuE+DJuaByRszx0gW2BalkNaXsE7Ocu3LbCBuqV3FPRqDSQwFWQ3bRkJA33CDqxkR8
YPRPH7Hw0bfKl3mdWnD24YLidAegJ7XXConvxSJOT5FN+cYClUIQVG+uyROb+RIyaWIyBe+Wy/Aj
y4ntqNr6At64POjGLhiNgNUOnv65YOJPmiVvmd4tXD9pDYh/Gt/3lmBCwy7sRpFmIvhjbeAUh2Lt
+DqfRlb/8FB92ebf8wR8cisAg+epbMn+ciGzuCJZ36T6cRr92nVHuT4rw2QgxO2+1dc0Mp9GNCvm
8c1uBhchHZpvHgGHW3Timd6vajFgMCp18F2PIfuxH9/hAuW2MMYeGWX6pu8z7bb6UcUYbbtlo/6A
PXONIZnkk87xYJCQ+z6jEl7cUY6SqlOc4m8Br4b6fbrfY+FYEXV/uOObSqw3vZ5Qp75aXbADNtns
DVyJMgkeoGuMi7hf7uLetKd4hlguWaePUVgzXBBvu8dTLsHlSPPpVViYJeN6BW0N71L5zYXnr+p8
Vvh1AL6gTOUbpzAUDL+rMflb+DLMEVa7gQwQGwt8fqestYHbpx5N/EfQpzJaMKG56d7JWBFIgQrx
sWaoQWDX9CJycdn4INaHqWhux9DmffxO15qQNsvWwMcaLD4iQhrkxzLdQa/XjL7GVvPbTIoeIqyn
HcgZai9LJ0TehrpvLeZmYovPioBLKYLoJvnBqT4lbU7FAIrQgM6w1d4+KUtC0bcLP7vkI+5/CpoC
vfZxmwgAeEdXZwKBDcFhSILIitpL2X8p8W3SeqJWr3nmCajNN03QHObbA5KI8COc9TkX0zoq8PCx
Javw1KoRi5VSW85QUQy+WS/bkz1JiJlml5UIGhKXcahtmPO7X+LwcIa28O0UcztLfATYI8SAjVR+
askcLoKzngYnW+4fFVKPLHPkpoahtHr0VYaRKVDa2jB9noJ/p0Uchjs9yYCjIRu725MwD0hCWw0g
OyS2f+SUhd9iWk1HCUZjJfhwSrWjQdv94ER/082RCjuBNwmGRDgjj+C9NGt7BLm6BGiD1M9Smw9k
ecGQ3QmaNuIBqHTT4UU+zlyk8AvJqRevurYfh/lm8+4TAhHnz/PCBepfk0ODcYhp9kXY5TwMMUCP
EL4W8McVh/N0NlHGaviRsybPBw+qVhF70Osh7SPIuEPF1unFhhCXtiEGX5k5/70fS8ALrUZsEdPC
ljlGhiE7C7W6U9lUtnAb5VP0W0oHL5AkF86hszGVatACVCR26W/xLif9isR+LwDW21Snh2cgTvaQ
IhUXsCveG8qU8K+eFwR7Ue9ic9epMCV6AC6K6aHNI1yTMqeZIXbBvsAXEahvLhSjGsKPt2K6zvZ2
t6Dwf2qfO+/KJXkhBDlInadZsGaeOUXQlWx0SXd5uRLEoWhFTUnZUUZXZBuJ6sIjVRQoKpEFxR3l
KisgG5qPAPEgIM+22oBxRqOg+LriOXE02oc7/pJ2Re0TW+0Ai0Awh6/rhmi0QYcdF9wQODLrjH3c
9vVfJgK3ayPcT3fCd+MUpTxE5Nx4o+kSe9ZjrnbTCXd8VrwRcg3eau8VSj3Ml0meIJ2R+rscE76G
thOIRbeWtvcDndegii+8Cuu50QXJpagP0XIwGZavU75dXdVcycxOGUw1bNLgzb8hgTxzRZ42ET4/
uixvpHh41mgWf2t8yi6XE2P7uSPfVd0jzttHiOtV6SWUcPplUWK8wC9YMnBl4Q9VKpYf6PqReUV1
uifQtKq+c/l0vkQ2ujDNXuFFmqnjavhdT9Jnyy3zeydli59dVC31E8LRaW4rZ6n5mpLtPflRpipw
gzaPWjaskDX/p16mLeHblggkiJYvSnXMZINftGPDg0c3f13X8MqrSjJ5u6Q74zMOfXJXenH/z9A2
j55Bejc/qEt5cNVfChDpyBCPbdPa0uffomS3V3wnmlXklikvvukPp41Gkj2S59OnK6GxY7VUg7Sv
b5CNTzCYgSQ/wo3uQHaKPzOYK55jzMpWP59zNEpKSx6DKd8vYU1ieo+P+ghvacLQsobobVd5hcBh
iPJATYChc2gZPVdOwlvfepCtjrAFKSpPv2OhXwXh1kFznNNMuZy+JOLoYgsfZ521zB8h/BvQxNPK
sP15IJQWXQl0fkiroU1nSiLfRwQvaeT1fWIum3h6eJ4MRljnoqLJuSiAPbPaVo5/CWelXikLnCVS
A1zzX3tvh+1Pq9IQgHlGv10r/lWQkptusenGWAA94hDjX4C437qjjQuhiShbfx122YuDIAQbudXz
LFGasdYU7+oazhW0C7C+Zgek4Q4FriMtyZ8Vp0Zcse38iK5KWmqnsct6ds8PaxYhVr1Mq2/nrZub
GIghF6ZZzF/5sP6Jmzv4symQa6oDTtNQb1Ku7l0oapauCW3hYG3m+HtPLD0YcQfgGDugEsLYmWqT
GNfqmamVg4YwoxvfbnX7bDjfthOak4/rjyiF7lBxPDRAU8oYA1IVWwzTufAbcKQE/sAEzgqGRPjQ
ZMf/SBKzCLNK3345nupBOx8hJZyCvvGFOhtxyz9OFzNu8djrr2ZeTetXo5RjC0sEn6jK6xqtBFJj
ytiwHV24bwZ20uvZ+uPCgQUnxJl8O9ye8o36lQiZAMID2NpEyk4fx1MeLdsyvDP9LnzLuIkJamCL
FBq3M8XJw9U8oh5y9dVnFhUyiZBeE/7cZqOY7Tcnpi9IeCDWCMZw7LdazlYPjzREi1eQ4pJbUyRk
usi0opqz1o8LHgWj3OUM41jZAcbPoO8gQ5/daAwgrVlmu82W68gjXKRLNjn4FXJr7fMMhD7rm4EM
mg/5gj/BSEVSyk46sTndIpVQ7WCvZE9tZdE5qe4pDLJU9gqGBZYXm7y8tX13aYTQ/QZ8BiyF8jev
i0cPQ2k0wRdY+GmEBkvBVwAmNJeeWwHnDCTX/2IG8MRsnZAMKcVM63H4CmT3joE6vB2W7xgSCupk
1deBfu4HcrYIFje9ojKSDskjn7vrfLUvEvwl5v3TpqU0TCEEIheyyntLb+rCdWwCUbw4Ak8tncbk
o7aeNAY94ZESP9S2Ybdnt7AQxW2wQm8s9ESlx+jLlPt5u5DHr1eiCGFgWjt6NdHYjuKFeH1Jgejt
tK7NUsLqI+8C/NWg9D9PtR8IaHT45UNr6LieaQfeXG0BG8YaYmJ0hiVN1nUzE3oDYsQd7xN754BG
qly1Tml2pg4fi9bdo22EfOisO419alcuIwTj6aWh+f/kH5iGZR2qFmTVhCRlZcT2dWIWBfwtmL4h
a0bLF67SZedlkgHfLFV+eZ4cskm4uxHLZU3MK+wR1+h8pguTEE/jC4/fpurkEdhC8/xnzfqm5c3e
UwI+lU/z06WDZueUiP8tUXUP+kB5ggUlyMd57/hJ+Fiq1FpvXOPG/8UASLVnfC7G9HNNc80AfwmW
JViZBxsL8YNWimAofOZQsAEgOe1bKaIo2pHfleva66VJo+tTlPmjqAI3QEDnupY9Y8+c0izGeHB8
E/12ZKWCpSnrbXjrtJzScWIg/cueR9Yj7DWCtF06LOVtv+mjbPFWXddciadyHO99tBtGlzxM3+t4
dhmBjxOzg5G/yhuQd4pSaXT/C/NhRO/FP7Q0/imQYiK0H7zqHHYUgsL4bC7yquqdGZmZgJCyuftA
GdMJAAfZBzuxgNANMPRK/9PhvalizcHhowmT/EXM7bc3bZ/ZX9lQTXY70AuW9vxcw2jhZL9MevJ9
Od/NwtU6ytfZUSxrnmTsQ2oYZmGyRXOT1ay54euHfE6izM99Qc7hBHAgmhm/NmKFN1vwaAcCTRX7
MnKOl25u4PmJCa3+eqpO9fq89Ukd139kvu6w9DN2uTvW2C6FbIg9x1wzZjw2JmU9/2+BEK+XiEHE
GKhYqT02/mtO9NPtcWrslYYJfndqNl0Bd2q930xK7FnuO2+LZlq7Tm2NuBhCOagk3aLYr77XlIw4
9kYSs0axuNfAWdxbp/1sunB6qqrKFa5R77X//9VlMwqf7On7iX+YBh+GaY/B3shxM8B7sM5rFImK
yXIBeM8OVRKp7/i6qybY5Hai18PvWeS4UUM+BvZqsS9x6oejy2lbPlyciNNn9nRCTYCW1hyrD9GD
9JapLvhjoSP0Z/l5E/GSkG18ZuG4hPy3M8l7h3mjR+Gc1JbxWKzbqurNNeNGd5Y7ce0gvKKngrXg
0Fmo0uYAOkXATYWaVc7qbZHgj2B0ND2AXppj66Zmwc9yLJP+YUMke/5J1+bBj43kU2SmhkAeuO6J
mQrKzYQz9Y2fwDeLvrl/vOIiKTRX15EWxGSVzX8KLnB4zSFE7Tb8B1i21IYErias3ervyTpv5EX9
iiMfQGYX4GdhpT6Rr04BJ/wbxVS8GzQSZWrYw6VybD9EA9hZxTv7G/KJCx59TPCM+FsyqsAnhbXl
DdQZ44p6NcDrfOVfJCRucmLVEaT03JYUbhSSWhm/4Iczd7K+4mdR1+1jE9b2fAffUzvMeHX9D47i
TQ26xF0ZRBPssMmxxzAUqG1mNNvReMaXfVZAHlWqzPN16Dl2v7zTOJP4A+qfxwwrBeEO1TPlDx51
yw7du7QgVoQDALjon/oXfRpqUjLTz22bjqRpHljYFMVSghSuB59F2V5GQqWZZcRvnyhUEeMesdSa
tclW0c1qwM/aA8QCwsQiRs+a8zIRosEM7ZVJNtnMBK+eeoIt3SY+3+DA3txc/45TEhAfcO1kTtMQ
AsczPdAd5yIRllfCkgeYeL6b3DyhQr0rz7UHLwHMA42bhd/+OUXeasGAVoqA7ki2y4iq3N1qFpwP
ymTmd1sO0zsVZgqZxjmSF5B0Tb1fjUovon9dVe7znrX+0H+o4i2buPIp/oRAczXCWEkUsJ8p3+BE
T5AG0As5hzw0dwLNAascZinQ8jY36pccmD2n4efFJhdfHuRjuDuF+CsuqLraZpWIk7k7TRovp0q0
WcPTvtC1mEdp6dFwBV9gZCykU2fp4YmwGifkSiRJEvjvBF2h9vH8YIA/xxtI7UVVQbj3Lqnjx7r/
6OsY3L43Y4qT0VMe9RsfZdZAEvriNuGFtgHs4ckx07mGCLOhgMPSQmEc/1swqJ3Z8esKFTw3h7dR
KGjwbPD9CqBJh9r+lJWs1bus+T4zNX8H/FuSvYGUtHSL1VpWnMeBsbf/P94TzcU6uDjSVSkFQSpc
Q8R/Ya5vbPXdsEqeSwVqsgrs+e2p6oZjITmMbVX9giNz3HYeYerYfl34+QePK4M3J01f+40Yh8u7
+cMKnrEIK2Sk+4X0zHbbVQ2FcB+IqWutEV4evqJxU5DU8UPhqrxSbXGN85ws4CII+G8EcAYaGxPR
1D3ik1NpntLv4oHkt85OycxCQUGtmFgmAhcdjW2QsWNrx48NwgwKr0uOpiM3wC/n0tjd259+Hb/X
UmN2+FUDfbi5vDE+t4uuFHhh4rRKcBQFmixfHa+ZndfKjB6q4kXv0liKIfhLDjyhB9HLtY815+D1
olSrFvzt2X4sRygBYL/oLSW1Y6Szwb+cuPA0V54QkDn4j78XvG/y96hIJnKS3+bQY1xjzgTDIqfS
LhzEDpnI6cHPvCp2pY2YA4AKCzJ2eSY2/E+0RQIGinBQiMEkODPtSvXgQqGgrlR7kMVdrbyZvDwQ
MccI9HLtteNsh8g3PnCSAqoFDno5TGPcERLM1MtjygFeXq9veKaEuSEyKfvtR0RnwYvak1Y9NfEG
q3UcLu+Lq17JcPlnX1zK6syf4NHvp0eo/mmZIs/gs19SMcVbV4amBf441J1CMJatoLtaXsrQC5bN
SMC5O90hhKeMBznLt36ZbBJ8EKexg1MvRm46bejPLK/LUKxFSHDYIe6UayuaoQo+0FCwN9R5v/sd
v9scCGNHTy6d1R8I9daJXEboocfwGYLhzf/5+ivUuIuPWyq4sQ1ueX0SEMdb0QKoVzA0sCuAEJY5
6VppT2Tp8wA4n99hszRuMFYoQrwISeRH1qRYhNk72LP16s2zNKIVGO7d+oTTva3omWIKD3skrrwD
PazdX26XNZ1GFE5tH2d42oMsrz4BuLi7S4wL9LSVDdpfTZ63MRD0dFruRJZ4Ec4F2BpGlo7NZUIa
Fr7bZP/vFHwrippvdpssL1LurwKxgBGTZuacoxHaUEJVass2n2Fi8LOCSMPsVs4JUfZN0Mo4Tlan
Jno2eoGB5yetABPbRDv2j7ofBazvJTONvtmqOjsXYXNYNlAr035uJuKE6Wz0Oe4GNtfWkFXDft7y
izBamG/XpE1lrk2bRcXCik1YWH5rm7xxSfVs3Dv0q2A0d8vxezhG3ZpHlJoCdd99/F6GVJ/b9yTj
zWX7OgrbJhMRlJp1+OWtZmQJuNgVObjdxfdkjj+CnbIfwVqz6B1GFtSvPvz5PwcnNLCYAnKtiLsq
T3i+ltS/Fq+qvbSALoeEjK7t21Q5OB76cfj1q0aheHnwdTI5FUX5cz4Mio4BCEW+SP2vuMXtlm2q
vZSSuRJ18cYXuehSW0iqiEEXW057/jKXN/3n3meANkHzKozqL2im4IIvns/ek8N9eCdW+5ka6xU4
FlPDvrPDoJVcIJrP7cw8QHdLw5wtgxJO3MZ0f0COKCs6KSEmJJvC1xe76DssZuixwDC6ueYUgDww
JtEGzkGvDEf47EjfOMj92aoP+zM7YDcvxiO/8IDUTdnDMqfS23aNfCxZqp+Qsum07fvWL3D7l6JS
V4p3fUr4tcn5wK7UsWsZTFrI2G4ZT1QYRTvQfsoR9TGnMghMRhWBLil9E1nAb5KDZsj5UBtTBT+f
IZ8T07uxAeeNLFQOYEV4sdr0JwdL5B86CDtHgj6mGpST91ap0niVxHnRPaBWnh/8zsxLLrh6vYji
hCZH1x3Ve5u3e30JLt5ErBgbfgyI8oIM/9nsaZPuJrgRhU+AQWnjobZcVNTyzdOVjKUl/QXYG1ns
Ymoc7CcESzoehzfP8sWgPF9d5y+IPWqJEG+x37PNIPnPcoPhOd2gfqXrN3EIVV+PvHyKfEbbjCn7
ud4jsosDmp91R7+/b3gYDJhl6BJyhAIGOt3E2kdcNQZH9y0y9mOLfMi4iKRLSOrcOXW73+RlBlT6
oweCeCXX/WFnk+Sjh3RigI9VC3QnMjKR+pjPZ8MtafQuf2lSsBsNYmbLLbu2bWdwo9blSIxHXLfv
oG4MwbkruHWPZYuldXJ4RHB8tk29a+G8ERpw+h43CX7vKYB/YnpUm6eiW8xY74Qq/qz1sGwf+/Od
iZh0q2nAGcegFi5sMECBJTQ9NGaQFV6rWu/PyipRo5uIl08JtZvYqc3LxhdoFaJJat0+3/G3H8wt
s5JCwmihbf7Q0AcsjULdb69CJoN/jnKFKnBCs0zDn4TX8La3SZ/sIE60AdYlAZ7DQsX0Z4Gn4sya
6SaZzO47Hj1iLjw0a7b7yAKS9wqNRnBAKw9B7XBOnlQoTUeS8Ecwbh6kp5a4UNMkKRc+CTOijgUy
tnIZbrbINujse3QSCPOiUJ0TCPLYhin+6rBTOrEKGeTOTPaSe71bTtuIAT4SM9ERKwHF0N/CELUO
yx/bxZ63IBcU0GxzdbALRIUKULcAzU97KghgP/zraJ3c69FlKvKohO3KktF18fnT8zoTbxZEHoTp
2/9xE6PNXwyknl+tDi1M4UCLK6xGoi1l0aSAon6ufsSvAiBFFmdBaYueH+qwKecMRuLclZ2MpY/+
Drss0Hvkm4eHscGBaJzGYTQvtZpJq8Vl+RycsF2D2tcyH5aR3IB4Hv+HYQgrTVVAUYHqqyylTwuK
ttl2gX6uA1mKXa8VEfSw8vxMx15ln//Z0kXhozRcXWx1eDSS3v9GQfd7dxAlebQIi9yLxuXB5TxP
U3UCGJ1aMS3hcjJbr95KZJQFqLOfwduLM1S+rp7Ei8NL2yWFD2qZE2xFVrWon32wHpJzXSjYxjvU
/SSeH+6Ze+BS6CI4sH2OhwhVYkuWCGsRSGSmdrRHFNRwzzq28lEOms/COFTNHKLq2J+JwAZ+X8VC
Rx/9QslTvbC90mp5hJwxSsZLYowAi5FMAa/BhrjImY0nyWwvO4jtBTK5riIkDA0EpUAlqXL6FzFl
4jpYe0GBwxHBwOjCsk6evCdUsMHVPiq7LD/wjyKo9fZyRes+0oYH1ENNZErDsCVA2RVWpcUisb1h
KIttrlCZcN47b6FcQSrAybrFLcaXjPjW3LAMzFwzrrhqMygS6/0bIm6RB7osHZ/nwj7FAIwogsrM
TpRmtIazNxxggb2MCE4SaPUHMcuxMIg5ZobqbCb3tkwyjJ+vXKKmwq/4N/kTbDWRbp/F2/ljOGvv
nWhpDQFr3ZW7CfyJbeXGWdTI/TuVcdjdVsOOL1YnS5fQYgeg+zPcnKX7FtKLiirhKKQ4YVQVMLGx
Gs09Z0LNtJ5svYkbyMk6es3TQxpk5IcCMaZOYqN/y601dEI/MPp6wAnq2oW/Wp7ZN/eMp/j9pqs3
/mLhynkDKkZgvFypX6G+oi+gHNtQXYZponTTCKLpY3UlwGRr31tE9M8wMK5LICh3uCMLi+CMPPXQ
pRAHHMWIvhAzDpB6QDfE/eoATnSrWXkYjzth7ru/uLW3SkkeMpctwRSjI0tJwVEw2fVwdVurTAi7
leUkhW/qnA3fB6uDAY1a6gSZ7+P3MEramOLx4AcXngbVZE2YG+cSUYjD3P9vHLXJ/3bY1m0EbPNN
mpO+XVTtfHbRN2NtKCs9k9u7QHPx5MvbHvZ77AkwB8LuNo2Bn5Yn3d4H5dwsPsLE16wNRBMk7Y5q
z9CwmqyR1x3tsN8Hf9oqSKn0akJMTOc009m4yEVftE+DIWHXJ93BtQ1PWB7VUJtkKBk04pz215aA
mHL1ewbORbL4eyczp4LoGb5fJHCZbXDyGoUE6whv5KHsgos/Hv7xAD2Bxdz8jH/+cgDdwBZLSqJl
9XFmG97qEcR/dmpOAP2HexE14o7mxREGQd3lsMXEuTPYysGtD6Y61qmZtiEvUkVqU7mn4R8PJX1j
HLJKuLVWHmMnKzNI4+o6awCIxSVXEStrkNMgaFPHxscPWRvBkUxFR2R3XMtFLklHQ4zjLelEmx6A
noK9seJsOrCTsYHL8nYcOjzA0rlzTn/pD9I0idkFoUAnsxSro9ffd4xf+Tun17Xunokx8e29+aEs
JP5YWrnnZC3TuaQIBAZEncc9oDtz/uVwp8zlHrpCLhNYshDft5M/JXUVVAOp9VQgcHWH6Ficilyi
eiTf4xz++SFk/l9Kqn2P0wWO/r0dpRqsD1fqqo+H5Vfc2qu4sfbpZJo11VUi9qCA5EgJ4XyT/TC1
5brnY6WNNyaAzL7lJ39Fku4zUTmG50XQuByu/7pFTY45zYqlTLmihVyGCJukWHLsXDn60/HkDDQH
SqbAgcIzEyb2XzweyNi6UBZH144Qyx61wnHKQKQo6g5XwmubIiAN0Oex87G16s6x476WnorE4HFr
AMT/ZrcAiEMXqOA3YjaONPTKjU4RKSE/rj0JH+r8SYRNwrfOM2u2A4D9waQN6pfoO6XrAX3SdQ9j
tSpijvF48LCyPFZNIVlyUwCk8NmLLWMko8+Vni0fd6GnvTMRqAr+iFAb334e+ULoR5ymw5FgvGR2
AtSIBU+EdojxuepaYX6gx/LbJCr0Zk9YjYWVKCX+gJUpjqyw/4UBcTWcPdOOtfoEvoMh7Wd/Iapv
i7dAB77bHXSYGc1dB4HkSpQioYTP7I699/PFs7gLTbpeU8O6A8IhMGY5XSTpE3wA/TuiEdA4o6TB
ErWAGp4/KCLvvXyQTH0q2zGXDtXJbQOG6lOcU4MoFn1MKQ/YcW/yvZpsiKBTVlvtucaqiGlCnDCs
DdDzTx3iNREoqZU5a0DnVWIcYUyCDURye/8GCFfUDU9ZQM2aksvfae5o5MbFby7anx/z+pN24Nxr
4A9+lcPhbZG95xLm9O50pioYh8lfSHvdO+jcMFYG2rdZclrVCCStBPpuY07AiKfbJx7vPro3F+QC
RW+49iy0oAqxP4PvUwHVNA4oLOBnc/RTM/YvEathemV3alrXAv6kAAn9LNaNXGW5d41C1oTuLUms
JidHb5CGcoZvslrSkhzYrIttwMdtENwDn/40HhDATr514bSODHqBfjSAv6KMXjvDcVpzUaSRUfkV
LPF9IIW+UGav9b1mm8Zzo9TrRH/Gt2Tzgg9m0GdJ7SM2feAf+KaYlCCgm5FAgWUzVNM3bGra0oAf
tYwhuuJ7rJXxvuhEyy8ljsCjvGnF9DFtIBiSsw1m9GULYhqcL94XTHEEAPb6onZfUAIHDOobo1W9
9MNaLqqI7ryiDUZlFD1/GQbVVLlKPxj9KN6exkyGro4iCrjNnQRXdYVsR4tu6z95Fw6TZglrKKH1
lVkKAahesJSrZtn1j+sS6/qKWoQbHacO8fAsmlUGSubWMqz9boTsQG8K+Snh43oY5g6GLT76u0p2
k4tcfLuueqYzeS6pEvAughqiebPjYvebUjxkP7nzCGh/GfQ7M1OCletbtyr2KMmgCZHNhS/WbDgG
cFEKQCurZEbWcvsRRKYRuFgwzpxWI9ftDy0qnm9mUj/l3D0QOfg4NW/jJGq7dOP7PRJNnRckm+6T
OSjzy5Soo2idtOcUVOjk3Sut93gN3+PbL+zHD/OSwS8kEoQ59lG9FQ2nLBG1EWce75YkML0bjPSO
xsUOJZQ9zLwx+96i4j6S2h0QZncMIGvZF3XhfDTylHFYkH4DaFGnnknVqu5Rj8aLYXLJQWYP6V9B
OPvQRkWWH6n9rJnbLWjspiOqph9Uw9BT97W1zZYPlqWfScYNMFVAjuL9f5H9gKYyJdaxn+hcdaG8
Q+jBsJE7FRQ7fISbxy4+BQrdTM1wU9BMUxr4/nboKa48k//T3WffAJbTYyXHgCs9wp9RzxRMD7Pu
tKdtQ0JGboXKU8Kzpp9GRIGx1AnapDM/gR6rmkbytuHg9bYoQGLj6D13p/xH5zQTmg5T0SXer9cv
hHm7rMxToVX3PomtUVWbRzGAB4cwTJprv7iWeZXJD2+fnfZtb5hdGW2wLq144hTOxPSTzA6kj6I2
mx2F2GfFVtsfB49Y/h08oxX5QJnbyvJTB1I7nq83nDLTx3bLJrgmX4qTxNDXXMeAWuz0JE4kvt4o
Q3A0BYAWHq+E1uJB1/sr5XkRPoeSY17NM7p+TS2lL8Gx9AOvJV72/OOB93UJlznY/af/AYkpPHeN
8Y0LQ2krADIbuyTsaWwbQ7V8TqpJL7OmxR3LRGQ2qrP+wBw9QHh0vb91FDG5Ta/39UDrBFuWFFt+
X5nO9pDTkPGgleCS26mSWeSzcVqxKgb8iirinEG7g6Pw7J2lQEJorNphEj31q19+2tRw/01pxbcx
1/xND52urXGXKVrcS/Y2gCKxd16bH+hGQU2RITpn+Pgmsou/4ym1l8JB5EfYyfITRLETnpie3tIq
mjkuIhlfVD/9nh88pWgOuk3od49nqBbo/OVepRcMI3ji0puwSZGsnMnq5cYq1bmPh3MoRR24mr4S
fDJUJo70PWxlGXYj4Y2/E+dDAG4ZaopRC4bwfi8WsbNxZpPgfBrYjoOq9w3KE9Ldb1O9HVwCYz1h
+Wwe79VSuTIJR3ja9djJaGCXQqoHI1QxX6SOqflEx3ZxrSSfhC/otmSaDvHjpmm8ARQZ3FQ+iUNe
TvYmKXyzWT6k9sL9nbaaUlazAXCivZwseZV0yJq8pOpNrjClxMoiWLdoOA1pgVHeDDnjSDsE4k8f
q35pprOB9Bg2BO2KhMAXSyvDUjvL3CyUIF1eLJvto40V7dI15+hODjHO/hNbQ13zE2UL1kMVEASD
7zJ9KjugeF83+sm4oC7y9kowkMVBa3bDdsvpZKeLVZJ2wueCabeAuUbg+5xqX5OiO9Uhxf0HxODa
2z8MhiQrSJq7Z095ek/E0YLZi137IPsj8FEkrzN/6bnsoA/kWBw7iES/W0SQ+nhCbh2cEJlAq/m6
L3emfBinZ0S3JMZkyuXBN44CiB2uQ6aJyoDwlKNMyAT/5Ot0vnRnayejam1rvcJ9J8nh4JzehFdR
ISiewywiSQ+n4gAIrq5sr+rdHLwbvjUIXMnb+fnq0eXeWCdDV5IXiSgPzot5nHtbFNjJzWENoNOG
peiU7Y7PzVXtcJHu/SThu3W4JKY5QCdF4Rx/PEqTtoaT2H7EwPbC6LasHT7QimDeYQlHUuqwEiEy
d+j1IXbkxnhAxJH0NWxMYwNptaB53lsOb/1/IDQSiU59YVlCCmFgd5Ct9YrEg/lYIwdVq3fan2hd
kR/831OhcRubMZ8u1qV6jlJN6sQ3IB0Pmb77cKihqHu/pfost7lmPKXqskS55zzo6Ov3Xf5OawWU
GTRIoyA+NDYzEvEpdunMtdqor9mElxDkcwytQnZfREutNP1MNhDH8JaFpyPXNGGt/IU2T8SUI9Zw
H7wi5V/Ox7+q4MYV/ra8PugJeiBjLHH4pscaKK1SrIJUOVDPKAz+FCEVLtHb+oRm4ZwYK8nSmQCJ
J3UARF9QMY9RZRt8Mm1sW8KHQtLKHboL5qi7W7PgZbOlR2VAn/eMKB+F4qmsjRe+oa7Cbl8Uz9W3
WGlez+B07fb0bM7fIZeV2GH8/lR9iiD6kxagj1bCh2piXIiwdmbyU9GCxrEES4nsH3vonbPXtN0t
Xg8XZ6wpAvBkrZWX4dGkNqN6qsl3f4fOaEobPkaW5ezzFoh5pwBuUuMN/9dO8agU9rmGx2UN2DP+
+fbgHFDmsiNNkmqQhc9sfgat7ATtiJoA7xriMmHq8lT41kvpv7RCi4Uzd86T624yER2WbpQah+we
tyBg0v866MTWJ9tycL5o4oq3ysPSFG6oPTBk5z0ocJhVolQlyCyS21KaaeshYOAub0G8xyJLx5Lp
cfyjLdSULaYqdgYZBnZO3B3cpJ+XX3Q6Bw2G1Dk0Ol9eJpp26PRaaCkx1+BYT2k4mjMTa+93u2lR
k1elI8ECNF8ryrxaTWcixpXtsSSmbPGeYQ1LSQPbmxK4ISSg3VDAxO81UiuYkHJODdfpcbXFoF7q
VYvHH0+LomrflEUXQToA+GlbjLzsCUmRFWmWhQcJBiG3UqmDoCNsGe45Y/P4oFArCarrgBUnf5eq
qbRzaREgVQaKtz6JrJ4lNL1Nfcz7kjIe/CKpmjYjAnB6c31ox588QWo1gbyOm3hU4SYTnlbsNz9/
oPFsCtVSODfbLKicYwn/v6zzjmhVVuwkx2hYnDW3x+2Hf/gpjCCUENFHFwwTykP2RINbtCJHrjoW
dEjUzaAdMBQCnM2p7Nk8NKf6sQWGFqLRog0uHG6zdDNVB259kK/BiJdDrYvqlhXRxI+mGqCSkWEe
eT3eFiWsjTk7VdT0gWlEmvBgwqn+TydqJX7bF9B+wRsFIOtxVhEykn42AqzvYRyU55/CBffwWE3+
MuC4lQF4/gpAWP71CtxSEArRU2qxxSdhl4pkdThImjPzESpiRG+FoFTgvh4d6HrZy17z/LWunqS/
sez2mWB+bPx+2N+LmiF+4CXOajwPGX3jWHCAjUFK2OczLklh5Hq8ty46Qemltn+AtX7J0yVHNtMg
9qO7pv2WvHW8Jj2aYVRdXwbRmyfoOkpweabd8JcH4QNXk09KfjclaKBHudintfNRWtWaKAfXtsQf
n657AdVL1qiLb5/lYmXJ9pSu/ZRmkMawvr9kR/z+7ox7hBBYpQ/O6/yO8eq2dQly4tJVlB1xjNel
rD96aSHa+8hqeRT5iAmlmJ9+WQ2sUquroD/GPQaXFIZleqCCGMqrNMXCJ7vYcMF1DfA5lF8BpGNI
/xky3j8yQEhr4n7DtrKBxsWF44MqooWt/RpSjQxQt0LLR0esI1iRt26+KK/4tXlQZHeOnH2YQxmU
GXAX2krVBhdUUNm7/hYT4ZJ18D8R9FCYOfjz1Xon+hGRbTySJFydX9AY+2iIwwYBZGomBvarwPd3
mULC6iZOoSP3sNgeTDGQQ2fSx/nmLmO9yP2dNbdNeWDvRJz8O7OrLMNM7frUYRivKJ6D3bTGnMIe
pZeZ5Xy2vYQNWoLZAuOployKpTv2tva5pTbEhJyZRmZ65SHQ+sNkJyJtZWy/3AgZ2bFnljzcHpof
Mz7XpgagxSzMK1rgcqnzYN1Y8/I1HSxP1xUd9sDpmaEFyP2CFT4pMmiqkYMHZfeXRD01ebkhSn8l
qwKI6IOjz3tPv9I8EyCxz/M3nsKSTTWTelwiD4eLnw0FRlaiweEnsbUabY77Sm7VRnYYPOzigXyY
IC8WAcV3eKKR1dZhMTsLN7xwLnrkZSIwTAO8XqTpzPxvfmlK6Sb2mAuHtSott5yE2MSHia+xo+XU
HMjTejEZGaeYHTG7y9vlIPmIAMq0EE/dzzqMBnRwQ/Vd+hVgTIxN9/G+YEBQj1aocUUMeARHZVvD
bZSrVRyA9stkdSpypuC5Y1OFfxjM+PWAGVx6On3Fww7VwJ7gEC0Q9NEek7fWAs2Pgile6tSIJ1iU
+COPPi5/jWhgLwdahGTG0pVQMEkV/LmRLOcmyQ7EBAKa8WQL5RAM0AyEM+CNh3uX9IMnsB5NwykT
F7F94T03gtJ++2FtAnr1n+Xs4eXIIJwrxITkglHCrm3mqHnOsnu1Fz9ByVXOu0fc0uAi7zCHBNQh
YL14j+czJKRR+pTs6Zl4B1zml+Mtm84iTeVW1v3kRmL70J/0Jx2TyXNfj8fayTCZ7FJPNq3KCd4y
+gDVhdpE9Jom+ZCzPLELTKnEPFtajOBYHkRbKqeu9FDhVQekJPWS/kIn2gEITx8AgQB5vPxDtkJt
psdyv9iRriflG4QJolgDuIzUsFbIIX6Lcrd0pow3M1p/rUiYT1vhLCBMvQw5Ts/uFNga6Q6Ygssz
p+969eSP8YsTUIF4HNlJ/7+BY0iWdoGyJ0gE4xR822r64BGv496Q+Td1EQ1fg4LeGeztie70RwwZ
cWxr2B4ptV3pdl7p3HNKAELbukQZ6CRA7m7OT7lf8TsxtGKSw8kaBTukz9OfXlRW/cA0CBubs7Jq
f4EHRCzsxdV+Rm26qUVxhPOGcT0Os5VpA48evhlgBAXHyRfAGLyUbYRWbmhd7V4fs4HCIQES5/51
5JDxYQpXbd2V8AsrhHvOdtG8uONVnGqWadj23JEyr5GXK+yS0MQ4rjMyN2a2/YfhNwI+9UezpeBx
fbqZxdW+xjFaQBrsbW0dw/X9l0Y9eY5mSa8dvQm0RfySr6xK0vbYPktbfDUnbIXyPqC5xkfGhuPI
4+58RBOE81CSahtaAo4fZFpGBmXbXpobPM6hSLcmVBFWoOSxe5ErwSLc7/HpQWIUoUsjbaFZyqMP
uW0kuazE8ZiAb5OIiMPptpJKgi0aAplEi2doeB0G7Dmj+pQGlhWynNYYOvC14d4P2w9DLdHvzWcM
eDvBAbYAMOdk7JLFm82Y/4JMp1hjfXodHmTFiOS8m05Pxor+o6OybvYRaFLQ2F9A3xyL6s0XuFYT
VlB+gAJTQx/t7akW+JTIKVEm7VkMKFooRTmWroWDQOs1FIW66uX2FYLWr40CWxzTLR/j0Dz1vbM0
9vYnMKxPBTn8hizeGUGTyw6qGnMHXsZici6Fd1lH/scSYMsgSkeUKwvtsUXiJSOGi8HPY1eN9S4B
HepGRyY6dbSpdo+tBRtVkZJGzKED0+lqP0povsPUzxpK5NqsqwVzFO61JiIfw9u+nW8sZYWMinuw
Q/WhNKm2Z53fG+pYYKiULE4LYhBZdrBhOSBKZ5DfdQS3LmEe6qTL9W5xEIeuKxI5prUCHnYjizPK
qm0bSWpKj+HUloSkfts+0z9g4t+Jw6YafvtW5yajMeeIxMeqdZbgaAoe5KQ7YLQhmTZnA3wvvDXw
C1nESukjAGZ/Z5dEq371OwLsx43fYHRgitAw22MZ+KvX9l0fkRzKDEezXtVvdObCa6DrBDrfSwHA
DWSoj0tjNskQuVLaE0iH80mACq/uIhYNM6LecXKqN1mOb616SNtUSroQYCm8myiLLBlFaVWB7jNl
MWkDvCSi6PvvuhDcFNnI2XoS97s266be+8cNMPCQtauoPRM+yet+ZA/7Vp8J1MJPvyRVDFbETzGY
K5s6FWoY1A/JUTdUUTlQ/shIgKEREv+SML2uzpQTNyG7IRUAIm6y3b+nM2pU3zpW/kX8oiqrGeJv
bNkrMy9hO1nCOjxUCvKlbhaAM88pQujlLiv1Fvk8v9sRXw/excNA2SK3GRZB9PEAt5ykFcW52VAD
ei91e1UcAxSy9RLNxYvE65u7yoYiDs5j100+ehsqQy18FXKLRhaWinnvsc3tdN9FkzDas8WBbcy9
vz+vrT7w1QcGb7Eoe8pcra5EHsSEL2aqcuGj+kxn3dSgWk9OoVcrgI/hP2Inw7PtIVqFajaeBPJx
j0o1ax7DA0pdbjVhkaUWzpG0YJhUX7rnXqjf3uctCvmlWqrsUU4xhAYxtoRICDn3whrT1/cNG/4z
NpdUgvL9CQ4BsbNR6vfMsMsgxg8ZjBzZHS4W2cuyVaRgWl5G7muxfvukhBAo9dIYBCbfGeK1p1H9
yk/QRS/rnD5ncYmRVex1VbfkmuOBBBePTZsMrnWoNy/H0jFC46ce7P6ewhbgphI7ZpIt3+HlLGVa
QDWaTEeJzArBtr1F3ead9fwiIoTKg0IOXZsHdvxmKcB2FMyIDc/Zke0cv3lM8+X64lQStU+1zz/e
v3n//092AGSlCc7i2ZzIwcPlVmT7JZlVphtDL2+dWrpICeoRLXInljMe3MLel5/tD55HVeJFL3Uh
gfGKB/dOpvd9y0a+9fTO5YHjthRDtuV7OMA94BqncpsC6WWJwyXSHMA+Xqx2JhiHFU6LLQA0w8gQ
UsbO4mAh8I0VkRJ7JuuQ6vjGN9kaV0jMYYM9m1yAUYWPeYK4TclhjYsyivj5cGwO1emvgherDXDt
9L88pGB2HejMcGxVdt0FioRd872mxYWmeW0WSqXyyBef5nrnLaVGmBPfH078eqo0ee18Gx8TG/C0
2xIKRtjj21YrFLoySDNJtraxxtScDJgdxONjyPAmhY9LwbeTdhvLtqWje5A6EeYGbW+z+Ld7gYCN
0pp1YYz/GkbjERytgrMCcrKFvVw5T20jXEhVtKyLfor9y/IrPRWjQwlQDIV/E8ShnTd8+s2wvPXp
bLGg+ZxJPz1pnhcuZrVCrOpjxZy6lqF6X6hiKAaOp2ogWxIFbdSyPbQlrt7vtE60tYKS2UosSri8
xm1wBr/uWiikVqcPoe4hgfS0q9UH6CalhMU0/sK+IsEHukE393D41mSykSMCUqv8wItbyCVdfTKa
Q4ZGwQwph+m6GoxC7n+lKDW4KXUxtFHb9sx4TxywlvNyTyZiWZ3v7qnoyGDpvv4S5eaV+s6uLBCD
n4/n+DAAooVMdt9RrKwSXOHNoFYr6mgBLvdT1sMa38Yss56p1xebqjHae99+YeX4Fv398wTPigq9
DclPBe7NecdTwnS8a/wN8ouckFcdyAqbSNyZPmgI5iEzYB6X1Tr+0MX1g/qJ4lzGCvYyBeO0oiL6
cmFEc51eM2WzGEiJgWmKxyoM5tXnWSV5+85Ruknt/r2p5v/1O+cmoNQQdzry7pJtY7FDa4cnpxQP
VsZtxpL2H8k2rQgA0GYkXgsn5OtSRFla9BJXRIDfp2ZFXFSKdxiyvv3MF6fB6+Kzp/ahTZy+aHNZ
RtULEeXVAXquKnTl3xNiCnMYEwfvI7fp05Rfx+sMtFifmoB/jR0U5xAQ71uGV9fNiVsOThem175L
PQI4rorqqAwQ2CG+aqw6EZssdT+yCElvikmt6zctIGKFn7VzTAJgIRVT5Kkh1QwPn9zdbjLVEsLk
WG506h0QOMlhfDFlndbdTZSc+BgU4ax7KGtYmngScVnbgLk1bNueUVQZXqQ5ukDe/+hLV7xPQqQr
vaIctVo5Wa6FR9fhX5XcTRv1Nar5Bu96O+19vKTdwgsA6pnGECDTuldBmYrkOoyAyx6n2JcBez79
6GG7SDRIwc4zDa+CU/WHidoYG0xGF7YNA/7EIY0AfnqzZRM4iuoh1FeX0Gqzrph7QX+cym93IKsu
QJt7btx7ydxcfif2PVl+JfO08cbyiNBdihmoLk1HgEIMZDb2YDBPKAQfCVb1uAdQ9F+1GzpYp4Xp
GzF0If+RBhyWk260kioMzvF/bR4gk0Tyw1EXN8++N4KLvFNl4rpkyNlzIhBCnRZ9qXZfsXw5ESn+
v7T8G88K7XkWIK07ugF6EcXXJ6VSgmR2RnMVwUP5gdm+kflf/F4PB0L2TmFw8PjtIDs9h4x34Mqm
9mozhCgE2huyVExYqIm078QmvaYoUQQSAW98/nMV5tmgQwoKM6IrC5nFmP58BwzekP7rxYCFWE3y
Lp/Fjxc0E2wSJBPHwnxgKbFMbLmiFbATgBEBfMhcQFkD8ehm0tS05UM5NbPTsoHQHjcQ6Tq2fVVo
7+a1zZc8Oj68e8RF4RZGyTF0va9jbb5ZiwJNJFsWdOR6IWv6iZk7T31hmqzxZhZFNRPJy6646Nyf
qA7syhqachd+pXKTP5j6hgVOdS9eFFlGnx58sFn5cgVccsXDHKEdp8w90V0poJMiyKUkGH6KJFlA
/Arl3SEnSPWYl7F9gIsfUCCqamRzuLslyAi0XAusN4ma4PhgwXMg3Lrs0TNmbOlWbzznAALgSaVO
EpNaD1gobbM0KCbCGVsmo7yS32vzL/JmyvFYl/SLbICl8bvkrJ+MuTgow0H7PzRYozthg1XxJ/sJ
5kObkKTE8rgF+fRnFnpgR9wNdh7NFXseJqzabuEb5YBr6QHOa0mko04ekJpx0LCYkmH1qCSd/+8Z
Rwh23yFTlPpyYr3z0zmmpFAYyqUMP8MZf0v6PIvaNL+dNSwwCcMt7cI/iOgjP3d7rApz1v6qe7CD
xhAmEe7+MGiKZ6oEqXVg9+skrTcv7gs+a2+Wgr27TncqKI2U4IOzDFzI6Kk7NJIquRAsvr9XKH7O
8YObPDXf8TajDa9Kkj3dWgPuLAZcjkLODZbkBHmJweVLVxo0lr9vquWTpykZMN46Ws4OMlFYbJjt
2RFGI1y/vmBfXoRTiYYLft057I4u2Ugo9RtCGwLLAXGJgdC+vRYTLjJ6Ik82DlIjOGTWWtF7gF17
8RCUDcNCYbBZ29LpKVqFHOUrCAStqeQ5vaUyBQXIXPHearkQtpXfuFVjOj/ymBxMPX6NNeBk+GW2
Xfg2Z/I/LI6/XNWOD2595F8fUziYI4/G4tMRLYZoWI4IrMJgz5DwldLPFSmO+mGNto9bzqc7/Zeg
EeF7qqfzU/WRpyfsHpn/4AnYmxrO2Lfz8hUOMw5l24CMPUGZoka8R3P9FPFGhKbER5vXJtxnBHcQ
EIPCF5jLVjcEAIudcaZ7WrryBGC1T3rTLRKVsP/i9bPcjwfj0SpiFBVz5IyzEwRF15RhNf5YZr4Y
xOFV2RA6GVG+6HMf+pMCI5YeQ7MNJT4M6DG1RvIGOfA0JGZfuYtoLvq6NcWg75I0O/+1RVfZXmRn
LR9kEVGht6lj6t+U6Fbcb8wLnUhWmiZ/8MBPI+GjrPhkL8/1k8zdKMBwNRlHXrjxRqGDj4z3e//Q
GYgMiuQIXREn6ItTdX/4IZZ8XAQkzjTgmLka1PeKPYfczC/o9y/5hyG4jBRj1EKeuSRpM2RRv9KW
PC5OeXTZ9VLYtzurwwcYMWLsLzGVHyKrePCHCx9uxNEBP0r+TB6AqcAkvhIZQmLbdru8Ym5xVm3Y
O4oh77+puf0flU3H7WOgGISWjN+9oOrX6xZsezFttE7dN6UUSlg88hUiwbL08m8SgPpHHrOQsl2p
kyzxSP8N5gqyFXhobr1Mn7oVZvgydhmnQxR9214KsOCMpmLVC67hDQyS3aHaQxryCN7imonFjCP3
R/+KWUb7N98dxP8RjS/Aux6F3i6sCO6EF5vNMk5XXoZn7Kj6bxqORvtCerOLlJLigtF/+4+IPOCw
N7/4Sm52fNRhtgP7qZUqWOzEaOTWciN3XKlER6QPTBxpDjWY/XJmXAWirzn1mnWvv990nib886l7
0LfOGcsPaEKm6tlVC9ci3eJXy5TM3bQoiLZ/EdaXyitVeD673HRScL3v0HVLtSlEP0/bJir+4k4v
a4vDHVGUnDdHKpV8x9SBj9iMb+NopBQ6FAW8Dy9YpFN7ynRo9k1reem1wxXukgddTUNQD05OlYwi
YuGMwsyXamJQPk6XLwK6vATLiA1ml8wX1Eo+ZBVDPBmzIvuJh76S2rZo6aNe2iGqZvvC3iVBOOjJ
f3hwVr2zvbLGO0aUmOG0ikiOJ4To6tdoeGOfwaUUf4h+vevz7kD9J3pDKurlWV3ZacubzsefvXP/
g2nLT1nyAVgIpNWMwOB55XmAXSuEXbqG+jGqhdaol5mU3DcS1yzE2ftT5UgjEyYvrecLPzsxv5qJ
mUQS0cSvmHNYUbHFF3BSBtO7EVdsnVsPZlTAFN82FswfNvURc10keq0nJntMYmGA6gBWEvQPV9eP
0zTr9GDWCZ92SXywkVrc6qhXRFLaeD93Qt/4np5FmQtptHciQzuPGjbA3yBnp2xL55IqO6UuJaZS
+rDhu3G2gMHP/fwUAxoCE0X5iHuLtxKjdnIHoV7rTjtmgGfsnyM1SGNbxRZnFj9Wx94yTAAbTbDn
3emCCbg5WLSd2NvxuquyqDYaVByBuovjSqIPYNCq3jJnmbr+tj0Sv5MZEIl95+DV0FUzDLaxiZ2N
ITIFxICh6ekoqg0MhQVCXvCdS72q47ZDZ8mo/EVDtZlswc6buPwfiKWzKsnbzyC2W31i8gMPSzZI
umGCz9x6kACgkFdqCpup9xcJ9MwXeyNF9+iX7wP1F9ow7v4JQcN6MSIFTiO7a78V1DzMa+8vlxfP
j5JMwF2xWEerpgjEYsk7b0GPvMRIdCLlBCevMcBGjkiWc+7UgFbBkDJJGhj5eYp1lLCtefRbPH7E
8svGJ4h+3O0mbll5Fi5pKbiN1FVbRJ9Uslgw0P36LqnSaEPsyyE8l/4SwOT7VOzYxTV1vRpa8lkf
qpBKhu5S3yHdh6LAbxYjTQd2KlROJnIoE2vBWjivy5IhKePIrmCL6SffGozKqQHt6k29jV85vwJK
VPuizQNrfwmdylGRfECLPcjXauMYiGPyr6gk+Jas9/S1rgxjv9E7ipDYvEw+WYGWV8832oqhI1E+
5PsImZCqdp4JYYitTRf6UwidTGFVvTXbadu41kk7Yq70C2A6g68jjRhScxegJExt7pc2Wor7QdHj
sK2J4zfdP5JdadbO/GA0csJ4jfJ9vxOSJUwk6yk5VNK9R1IgahX/5xQGL/dXNCTeVzm7ZnWs97qO
LcVnJU0VfrLOnNqXIHSYmm+oInYMGHjhwxH+BziuFRJ+K7ouMrDx/cgynjr3bky7WEz4epoc73EF
TAYKfvUWRELatGX0PySqc9Ek1o47o7z0DioKzpDAgKZTqG6vS7q2R+D2JmcjKe4pasQD8nezoNVH
fsaiKRXQXPhdzdBU78CB9mqLQG0Tan0uxW2ABKL2omxL6vyxJmsPhMVav9C1xeQvj2s/SfMNuoEq
dMQA0NUzNOTFqsNOllKP1rGK2kW3JNRMYs1LEJioh329NGnnQGUeBzD5tzwwJtHwcppjA7Frk280
PUh0rONhZCoB0y1kLrHX7+TyCKMAERL/4AXEuBg7MQXc6gEaQ63g27i0drf9lfBtjYmBjQeD7ofP
BDSHUtvnBVRcSSUklslKS/HdR3CDy0sMPHnmweyf/638EGWuy30jiCyiKALK7xs17s6Np7bXAXGr
c5UWNZR/GOcCGQwN/n4vLAORI9TeaYYRnSNgg5UBlE6MX4X0BAjNcOE7v2ZpjRFsYPFPrsdVftTt
aMMhPaD0+CfcfFlNAPy0oEeKg5PWcS9sNio17aDTdB+HP94JnBNUUR4pwyFTfkto9q9hb8RieKF/
ELLZ8ud7iLrgI6GQl6f6SbvfW5Pd0F/xhZyBrTSSodLEUcPdMhj96sQoW/SqB3W/9SNhYnjCGjTs
32rJ5yTUyThNzYOJzcBlrgIHOXApmvWpvycauyO9p1tICsuufN3cwEdeHt4sUb2clkOwOMqjHcOR
iVTJHpVAPqOfByHwywLupLIEBlrk16t1ZPx/VRYBs5We0q0xLXYgaTl2OsY53+rxcFQmYlJBYuwg
7D8kBzdFKfTnuIoFA0Tp8LRU33c+b0sHUTxzHk0Q2U+gQNuITvoshCvjsBGFLGycxpJjkqcrcA+c
GeRkYYvO2QOkoZsDL5r3GYd5NMrvRQP6DxLJNK4lhOEBVIfNeQnbHxwHGdfqqWiuY/3w+qrjuhrN
oBC6MkAcT76XDkaCE+stVeVTRiNiqS/GNzrmMVCp2YmEUliiZ2kIxNB+QSbBNd9W4A9KnyqCbIHx
sz2oP7La/D7wwIY1KSfrTqJmgZ87742J5WJod4Rz57ajm7mCOW3FL4fhXeC3jveuR/JMvh1bYUVW
tb/hpCfxwxaaA2EqLpFzddTuOuKfaKvUJ7PmaPEkdMG88KndpEBXmadXn22Spco1xmEynRhBLvMI
+DHEvqYuWuatEKpccpKMD6IihMV3V/g3jYvBX4lUXwRSqwYVjbrhwLY6TALMN7s2oHN1WB+llvnZ
lFZtAoulYuWnSBMXIO32xJS9jMM2PZWXLN4i4WcFL/ZYjNYN6RjKgExVgVve6N+hiZBkO8DXBDxO
LBDWPeuCoiEGIhurHdu90MLnjPZErdRs5yTnJZPJtKFqxQt5bgK9ynOdITFRJaoIJVXCd5GLlpmL
738QFoftHH1Z/1KZgSE/ZOLBX6sAYiqtU3AJjz93l4nmbgfEfELZ0UpXSJgDFi6nV2zd1BwI1PJO
OvZDsvXg1tVQIJW6wS4mKDA52+CIGN/02LbFdCxSOFRbMBcMmEZ1N+Mt1utV/WBIEiXMjZE+6zMb
DI+CMibz/HBjwBkB+mB2wP1xl1POuNMuDVOIZ1Ecj2prvf0ewGHHbK0K+Qa5k4LjbQxG8S3xBPXu
1dJ3Z+T1LaG27Oe0hoUI971dnPPFw+j7iTftZh0n4SkHDn0dB6VLnA3matA5MZgU4NBVRoThBUw5
T+5WjBx0EMrCwK54B14k+f9/JkC25JGvHyu7yJY16HcWE1id1r6ryUJShlW4i7JyVX/fnPP0z7de
8KHw9DEz+NS8svey5Bubj5JKc1ZycVJi0S6MQVysN0PddZcTccc3jCg+JNEIG6f19ToMuiB/6vNr
bZ1tILZ1G3k1NbH83z+4F9dpFl1kDcWqkTm01ShXSnw7sfYI8+bjfq/r1abgiUgFMIu0QhBILBEc
BJnmYHkr5k/pu9ebrf06kNiPJgdMFXL2GZ+ODJNv3u6zS8YSG5PV7WttiGgeIXAiR+Z/TvtnF8an
vuCEVbRbkIwOGJbO9ENwvGEwCgmupbOz8Jh3hx9MFpm5bqtJB99fYtTj+8k/Ymsuml4ErJh5gfa8
fYpucNvrh7TyMP475CoZtQUTMylcBwtNRjkYxOwNwuSyhclrQkoCKzLU2jiduKGe/TQ3ad6jjGe9
WaIXT3J1yNA9wn/PvXzGpIBOuCrrBLUjCs/GCcJ2aUMdFhN2ApwgGW4CyBNlx15/l8ub4vcKEPm6
bbfl0C843deNtut3v1gazK4Pp6+Opng3L28JFYnXOxHZh9ojQs+6byQEJhCtmtjau8o0J1Gmyk8C
NZH8c6gDqkW7+IxB1T6kuvG1nZTI/2H8oYKup0tmUcCBdVQukl7V/1ZOYwN8nk7WVbfIkpAdu0+7
sw/SBTQgeEjMr7Ac1/G0B7Zf6eOACYohB3NysEHVl7alu78HryBb5v6ojfwwu0GOCO8E+qfv5Kp3
7DqIdqko/HFyC0TPGHZIYvhGvsUgLDpVgVbdmssjT7Xa38zlJCOsAK1+kjDgocdWumGJF/EfV2Ao
9lxku0Rg5H1xHl0QwQz8I8dN2D41EqMTrwfrkRAxgEp2i953GHd3nOc8Ed/99hYQ8TLbW0i+bOc5
KM4NyhCKPLnFWCtDkmETnPKrbYDYGxX6JqQxoZxmWQX8bJ2PXnVFjXm6mlivQ9urmTv9exludKgq
M2ioU4YicI8XdUutwUybIhZN/2MkmB+PfVO/ipKqoA2SX76ZsTFAjA09qCLtczVURijK9isWZ99U
52oX58yVQehnmm9r8BoLzGnLGOssGfIkm5Y8TA/KgR4qbDUfsrcMuMwQ6se/ofwHZZbZpRUPG859
1ZaNaRX9dVD8EvPPlbnS/POiZODHToef3nRL2tDxgAX5Uo+H7sbLWMZU5aZk7P9Sw5lpGCAw1zBX
bVXTEeINtnapb1tYIAnMR46PmlVZ9GCKSrX0UcNuimPeP5jHSUZjSWXcURVWNwcgSlengC643DUP
2rkSa4u379F3YHSQ+SYTdxUt0Wk6eaI/eOM17otOkZB/5M5s16ZG+AFPygKyP64OWUgd71CzMbEr
Q68Psk4oa9xel6ULahzuJyEck1QsAYEF0063rSJhBfr7noesaC1RVdY5Vs4s633v2Lag4n6Zl1+s
GDnTnsXM0EsmhE0F09DKUBvbyaK9dkPAWlbZJz4N45vKlVUNmKM5k8Ol2RxJ0bdjoI5CpAb+tQoW
pofgtKmy2QM9cnqJrTmvrL57OqUrwRncW0rsLMSYFnWs5L8jCKOHENzJZ3IPmaskV15qkf2+mNMy
Om2EpWknLu7HZcYVbxntwItu3bs9TJmy6F2Okpw+1TyLwbJEy8HqYJz5D8WIqkwAZKT3SrJHQnbS
LGAvn5IsOOYHSL2hJAyV2WbtM9UKrpEEAoSqGmXc+tfgGswdWnjlGa7FdeG4UryeccNGzFDCFtiz
hGyHDoTjVkSAZvHL6wPgvZVWCbv00FgNIE+wY48JsDeD74OXw4CdWuK8pRvseRzLQ+Ys1gYukTd3
V548SGy6AX1EPbMlmbNlJBrJkg7kCQ8VCNJUMLo+7E0Q5CcZMWMeBnL79oagUEkPuwDls+GggONP
ZylU2DRffHMZs6zz/T+AcK5nudR36X1EktPtv9IkDjnr1P9UgE7dVL/lLR5ThN+Uex43INrhG+a/
kva5VztsKuf4LwAy4SaIrJGbrs9Fe65FJhTA/03IReQ2mUAQnxbaWL10Abt7Rhsr031+ffiD7Ygh
PYFSHAhcL0GwZS0tVsBI+887Vinfr/cDgCiKSArssiCXDtReuLy9WhUyx80Ytc9ecixO2sD40u5x
jd1kqh9JyfLkB7LMZZA+aAESzNCi9cJBBbXEMMr8VvQyK6NvDGvOCmOUduAC2EORcsnEt5nv4OZZ
lmCve+Z4ZowBgiupmDGo9+DfE0a9PHo0btFUybyGtrqcONMa+A9ndZn1ZWuXe50LrIbLzmJFCMIo
kzTAOSxq2NH8j5VWLFbv1+vaUR9KH2ClwazqEob14F6GTxZWDFboNHuhNVVPE4ELI+kkAWfPZQPv
g2n58bXCJrGpgyB0nt01d9LWQV++DSZGQWnWTQ0yWCA1l28E3sPFkw5sx7z+JSrXrvbu4Kkh/bSB
d6T2ThFE4KYXRO7WV9tmfHAxFpUleTc913ZE/tEnKlGJCmolTqNn4XyYwiarJknZkC4lnsh3xPWf
+rK6mnfYoDIkNfhrp2byV+XAAVnJFrPT5uSCR7T+jHjvkDg8LIj/771mglKPSwILoID0TGIxLq6m
xcDEY/V52ExPS6pQ3L2vwrXARcO/OK7IMlZcstZHinAEsdqSexE+WsWX6VtgPhpvgYfCUNk0iVLJ
lCDhSd8iEjqKKI8gU0OOcDz7cDAI80cWggra8c6v7YX95U635lMyN//QOh3ePooLAy3u6WC98oas
tITfXjj3kxUo0Cj2hAKfd+aQCqvpsJgNoYiAgfQMfCLhHq/nW2duwWtRJzdwgQQZV69tmczYBPGd
LkcG4qSsU6LOwhO1ZSKS0JZXtaY7REw2xU/ptq7YCEY3mZ4P7yAqB0EdrsEe8dPtn93ErTowNiBP
D/OVBZSWwzzwuzVYWFCTVb91KV+L0DtJXbm+j6TpsduEVfLz4RqvKFKLyfc8WRbfh0bnfxaV7MoO
sdsR7Vye7qAdeOe2ScVK8+8vbpR5fVqTOEKPkdR5BzINkV/O34zoaWP7959AYag4z+Yanlu2GJLq
mLdvumOT4LkYA0jgLclr1UJsquz/LiKtcqrHsOnb5OmZdRjLuUS0j7WzQ7rotO8Byxq/mDZW3wzh
5WtvcQsy/QnxJLeEXAstmG22Ao928xCFC8DYGFhdeQHQfUCWFs8ycGTTmpJoIG06/dFqOTtvPxVv
oVHirRDmvV6AmNwB+4OXy9WLC85mRyLh4UnmHGb0dpe3U23SZEv12QUH0zXOCyfXR//FX36lUboC
ZrGVDsiMt2q3NavsJ84fiXBUlXf067zEG7lSD4wiDbOqGcKj9jA/xYrBHrYh6qNINZ53scuHUotI
C5oAnv12jIUOpj6JyKOeAMqP9r5CSiwYruEWqF8G7hTnwSx2YmBlDwuFkIOnuwHn8PWjZ8SzjutK
TIpOo8sn6cboDWuOVdyFuIl7A7xfqaX+PZ3aBiDngyEDufQL/6uCQCDHgKhkTiyc1qH6RLHzykmx
kHvLJiR93AvtAZLfyVdsgXoq5hDxV9g+t1yK9qPII50TaQaHzkpi4DGvPj1Ucodxm/xHbBr2QURj
p/IYOhupV6HoqtiBgzLGF0Iwcid4nkBkxw+bXSIFdhxp/IqOAOI1K4MDnQskFK7DLoWV/Q3RjRLJ
nCAJRpteeJKZJGGUrAFxY5o/pDDZOnV3yp1V92Jyo9ks8VWuzoRKRMu6B/SuHPfV/6JwP6ZlqR7A
JiTQQrwOxlgFzhNxYEZASYTeYlhLutDkCg6/BGweeJNWhg/ycKCxw66dMgdUZvJqRbDkzTXFp2L3
06EY71BLiCZorV/ga3Sj5BFB6FAjILwKYFjSp3mUr7UMpInqakadS+Pb/fXb/t7tnzNNZgAy11dR
ExUahAhIWRDmjfD0ih+kUylSjIcIdvuD53Ihqt2L9NLL2fkZnYnGH3WeMKvvR0u56OzXUnurEMa4
bZt++GTZVetxzQ8k30z0TeVIH7Jabec9uJS8iUdXtJ3YPv2PLt1oDfYa2y7j2oZza1uiDzbfBKcc
PiYGFpI5LIgIXhwKY8e6bHvyN7EqccgGZQJgZEFeVLTj4DCVzV+GXGBSnS/J7lNJXAUfMylsc1rp
/FgLLivvFm8oh+Q9ZaEVCiMF7gg+sggveSnO0+qEhEa1FxXSxD5YvbHZr5qtOeGkqEjbKrMac/vv
LGz4/Uzw+b6hQgmEqrrB6VHkEk86Vm6wTT+DHo/l45M8anF/bIE2MYM06GghS/BHJ9Zelv88YVhc
UPN+J1oABrtN5GmozDi/MrHyqNvD29o2YuHWSoOiLq+VNzOQEFlNVxFp+TYwAqz8iM/PfmsYhQ7x
Rb9p2izh9YrEfm9vids1MtG6spygwbjl8NQV713G8pczw48xw0QLxQOve2Lo17/n+6U6XewZMAAj
UyJzRNeAo/SVGPlslDIZlF3DIdCyGsRnlCLjZejJXtHrFHghGbBbAjjfV1HN8tqkDIx2NtN/Xx1h
loTc3SQtzpmXadlF0RAPJuR/ZS4XzJDtmqOIB3hYxKEfxE0N5FL64ZVDGNcsuAcl3vACWfGXRMZU
HyBMpUtcETrrFQnOzlYDNFlNPAK64vPK+y4qN99pzO+N7gX4XvgnSa2LKL+vNjim9sY+1Df2xb99
Z5qYA/kM97j1UlcZz55je1X4Z0JIui5utP4JGN2u65BOJxKGMFcrM0IrdUq7LGzqySN7xuF43A5c
pbLioCKVoW02Igi7JNGBUF3gdAiKUgzZofMBqXPeCT2B2hPFjoUkuIGky/uFhd5qRN1YBsQy5HJ5
0M2JqPc+HnMoTemonJRsPy2vjeiyoyKXY7rinXPdPprId8JIBvjYciZkRVVpIMDBCoqxmDmZsTgH
sKhEFnQMsPJXcXW2zQf3bMSXP7QK7695x156N0hsmnvm7MBdTUUAql5mehtLOCjTR5TuWJ+gY0tg
AHRCROv2PYX3BoVz1/CJKzROagSk26w47W6PiV/7LEHmI6hwm1/YabZ4spM7JCFzLCwo8KhBYCK+
UZd3VsvcLVob9SauM+rTa1E6CDzGyvn5BHr/JH9mYD1iBN8VKOufRmw08c2EnyVK7Tc+jkNsK4HX
s9KILrXbbEx+VSb/x1sO6LfDV8Rcmsd1R/K39x3qcnlnvRsIhMkVrJP4OJWdu+Juggp8ojmaFWF6
iWWzqru37PD64zBHpFO+8O19zwSpQXrYkaTgtusHp8iwfvD6dXOtaZc75Q4rYg9EY9j8Eq2Nr3mR
XCC2hwYUv6/uUZ0gII+SdzEE8SHlWq+tWjh/1ku80NhsRhIE/YNOlRWb4gPiabXzR7PapZvebe4n
yai2GptQiYtuuKyWu6eRk4irJFgO89RIIsXINkSTZcczvIGh+5SXPpW0PeIMdxSsYTFqdpbimeKs
ceJDttzOp/jovV8Wh3wY/j3rqHnTAlNm/fNL4TgQZ7z7y1cB9Aw/QCiAYDFJ5CHXvpXleBGosXQL
QVJJOiTo7DNIU7B53F2dCRDtwymlU0l/JSIEt+ixe/Olz9cDTuLOjR/RXjfU9bAmEZFVEOgyFKvm
CbIMumnZrebNydSKYIdU7u4Nuqk0NzE4/RXF13jjSEOUZ7Y/AuqmU7Lt86tQ/LG2Ap44gb3LlINV
O9WPUJtE3ZjPFweV+u1SeuY+KJihScX1qbnnPy9Tt06zaJ0m/qGt6ViySxju283buF5C2hr+KvJv
sqV+NHO/KsVBAkDQM/ny+a1YotICTLN4ehZCdE+BXqXlOi1X3tPlpxqa1smpavEw67pY+ZGU6iUA
xr+S3NsKiDxw0I6rqh7OlOslIdmPHsLslRu9T4LkcA1ZpG4qS/zxozlMmk41pgZ+Kiv8rOdTg6tQ
UZZctFVFxhNyd7vkxz937233nvGSU1nFv1CCcq5NgBLTbCELov+KvASa/7m20jTZ7f8Xe1jRvVEd
G58CB6aOxXCeWHZSm1S/P9EG+xclWUe3s09m3sUVbo4FiApUdJ37xrW8iNae7GxwQo6CYPJRWNWN
xmUc6sLOx/GjX8HTvQdHZvQJep7zpI4+GTivw2Y6qKjGDXiISxgIJZb44t39P/WOqQjDmDoGw9WM
YDxHMSZhSqxxpKi8zpLte15Fhf6jpClc51WPjuK9v16z2eOwHm8zfOMORZ7/XeoyZnFR4gNSQcy+
nIJivD044C2zyh5eFYGCBu7FBt311rN1dsisZz8lPbJQ1sDyIbx5dbOEZdhAHk6Mmnsvnr/EPRUm
yh++hdF8lLMQKd8wvZcachQvFzfk2tNceaqlpxq0FE1bAfYujn5/iuKmRqJ8EZ92u3rkxZDGj8ch
/KyU2Hx/iOTcllIk9RRv6bPDkmIdPad2ZUc4TL7JJlXyBz8+1H5qkQnvJ4auxXK+Lg3TWFVmY9vA
hc/agvj7U8KrMe2S76rA2cF02iUMJBF0qPYR8maC6Ey9967mXU2mTGNpL4l1sQULL4mmAVFJPQCV
gd0JOjqdPcr7SZSZmm7wZm1vOiIVYMFUGC1X6Pu0c4Wb1CkNFokk9TAr7nJxn0mnrKg+wWmVDt8O
/TFZb5+BdQzxw+vbgY8IxhR2ntUGRO19B6sgnmpW+wzPbaA9PkwuP8swDJOB3ytixh9rsyjtRNIY
7L3IGzkwB+KwSpSBddo3KhPKqLEocq31K1O7RcDcXxLzFAkaRvI8PLXNzmGm1+a43FiaQ9ro0Yvt
cz+0kledL/tZY/Amsir4a2iKGATcf0Gj/E6DdmghfjYjxpTfRrIZa8h4e08ysIKfAX8eEC2CpFJP
l0kd/haV1Mmislpd+uh/QyRC7KnCK1VpxSqA/+j6jmOfxd9M1vTp6ZZMEk3vqEzcYf2krAjbVYdQ
8i2FcwDhDtnW5DaGlgWa0SvUl8by+DUggUzZjAlieOBma74JIzu+jlN+guZVqteJyvk9DtJ7QqeV
7RxyUCDGE29giSh+lnqh+31bPkbyKSW9HId0Dxrj10ZsZ92mKVdte2PHZegOsl2gijQkNBF/0w==
`protect end_protected
