`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
NxVqOg0TXtooy9HCUSzTAGmIQBpyqCSPn60n1MxkdCkYVrhsMtjbLEdhYKyzJc4KZLwBsZmLin18
j6M1an8NJGicmjlNoDalr3M4KdIhHECexZls18GGejMEUbS+g4FohaZ2y9fKL8KwV+n7kJAzuGCc
hD28tQwF5j7VO4UiULf9E45vebouTnOgZ83uhOuL1GCNpK6yKXE+o/H2dy5dTemVW0gaaMxxef4b
AscTgqk0noMk5O3AmeJNi7BZrWEiLvu8OIehO/7Y9Ni/36aEtoRdquqre6APwnk+lkEB4s2UWEBX
3dccaBcT18NHaeuWe7TlLv7GdSVt7S+O4pmiKQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="zfoZCm+cSE4+4LYgU3ApIr7D9N0x1FeYw6bYlt8eHvY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3600)
`protect data_block
sPEYf436iBq5azbsjsJnTzbFSe9O/h/qi53I8qBbvjHXjk0rj3SB1SsWfC6B/A7hO0tG+S9WfqQF
k072UpX3f1Q7Lt7qQ7ANoCL9/6ZxMdf181nGQWYcZZ2moJlUbtqtehjIZei4YHgrM1415uChWhUZ
bxT2F1vE7DbFu7fJ4BJNJGeWFj0PW3rtuKY4LcgmLHjQPX01KE2XD1Ys8xQkxgWeRYhTGF5+m1hv
1jWqcN5AyFyTzdNpFgeW9KnsUePZdBc3jn8TBlyrGFMjH9eF0egrXPsJFzty1RGO4hcYoOvbdfVI
Gfgs7ap4S5ehNUAPsPvoAAPHGbioRPCog7dyluVYZeszwRIlfL+dRC16LyLv96JFLGX8ELMu+WNW
1exh/q8U6UM5/T/vAoGGu4p2XJynhEYMeeJ0Hkm6ZbQTYuQGIKkcG6sPp4QKrolIc733zPEHrHVE
2FuZ1XrFh+aK9rU3SsSUuzrGSq5T+s2Qt24hGvGjXn/2YjULtm06dEX/apFantnmpvi/qAhtPFQn
rXh4o3zbOtCGUWiKk+5sKXJXmRbcvGDZzb3xRMNIGfBsgJrX8IC6AwVxSWDr7hkZRiaRhG/2OR0A
/lzyfZslh9sG7P8pRqhLZAIFgEzRig8i7YEng5mj+sU4wu6K2rmMEf38tjYQq2qdyqOnEs1Fk3ec
sndGWR+Sfk3er09ko9X6vyIkbqIoyuPb7y4IfU5Src0Ejr1K0wQwUfHUYq8MwksLZYnT7GEYBjsS
y3r4zq7cFilbXO2P6epe+T1WAOJvgIqQ0Gp1qoZcsQz3JplNMAQxIFCoZ7X5uYvsLOIBFI+OoI2n
jgNguclAO/3YAZgLCDRcZPG6ROU+TWgTUua4H5xGhqvFEk7wK1M3+b+HcVSVXQ0nusq8NxqSzqEp
ZHJT0ZcIWXWAVUqbkC6hacCT7Enfe8hHXrPcEuvFLW+sJN1NJ25zxt6gMIYrC9T90o4DNhBl3KLH
fZ7Fs8HgBXl5BMHqN+dGR/f3K6vuKRL7p3cXy2rgNR3vCfJMmP6HEFFghOKOuA4f0ubNCZvsBq4I
MlbQGl4I6PFx8bj8f3YbMql+j13I8XFo3jFJ5wxoRgDx+ANeaVG0qBvZWCgk1O0HOrXyHd6QeLZk
K1J+56MplBRnDw2BW31NygwNog4/ly/pLdSbCzNykrfIn9snS4ZCFnBJ+pWjsVt1H5PkA6X99cMq
TZMfl/d3cfaV3oIMpdN5OTcdbkOGe0qxkeK3BzWzcC3ptLAVwewOgAZPeCmby7pI0XMd1SfhcbnW
W+CmKLpP/rmjcZGTG9RK/y7OPIzwp6nDszcdtXHuPjPxEzgB4PTo6h6JIqSKFjK0d7qCf3JWIfak
59GOwOfkMJDwutpcf9rBCTnnclmRAQfBD3ZCLHEQzVs0Q8lnqnJq8906q/4j79D0srmFYt4L0Yxz
UUSApDAkx++TVHyktVDLHppLqpTarjIEFQgwHeRvyNOc4R1vfRdDGLPs6TD4kIUZ0e3+XLg5ujdy
yDxXsNf3aFwCMYRG+AnwVqAUawt4RnOGOKfVk6VScqGpAO6q0hb0QgUb4vQIi57uCSktlPr707U7
hakdCNjwy1Syy+eOAc9r5UFGXGZQNrkpCoykaimj9bAd6qGEvKi3iOorZvPc1U0ROl1SHVx1FH6t
7GgMHTsKwKegv6O3vCvgPsNvNLQSb+k0FbXUv8Moj326kKSzHRFyraC7vSLCH9bUYqi4eBu2TXnB
d+yrbnuSalQFypnQwrHeY5k9CEQKSMulyChNYjg0dKynXNIOlBs3peziCXgfemHBs8xzFW4rPdHx
xzODjpj5I3PBH93B03tdzrmW3LJObxbWJzJw/LD+LPp2erqw/JH5/slsb85L4HiGiVwxzfs+EV7H
GMNWzxbOu4ACLug0iA6jocQRloiMZ/r4IzGFoP/0/cq82cDQGLd/ifnGzzb1UBHMKcR7qE0i6Pgk
f2mtNRY2+BD2x8q9ymm/evjmFLaJ2EkG6zJssSOWH5y8yz8waeEndgtkDfTB/g8elW+uVCQmIDfh
91vIBEq0outjRAlXMD8tXnUlnMIq9eGYtBuboC+Uw89LR+MeHHDCOb4EBEsC7PlNKCLHb4Fh+T7h
8Z+QE57hh6PK8UewPKA8NJs7eNxc2Vn+XKhx4Hlpx/v3XNkwuDXnbkqW+mz3diAvgJpDJ0BiI6Y2
BYaPk2wyEpizO2PJm+qw+KTHtVLffkkU5kZjc9NlV1Z1yyNtljg3uQDTOf+ZfGS6Ih84/KlJN7e/
pgy545NuPCLDZJLcjzKCud0nohDfFg3aj4Jr7lCia3Nk1ifunaUQ2Sy5oE83Hmep3lIcrRKTIhwF
2kahtHUOtkeNOyeDTdTYpReYBNwmq58FRuxdEog4Aq9VMU6JNX9HwOx9DP+SFgWL3kX4Q+UDNZlD
euPw+PLCyiedzXGvdXmrq5UN5pNCw1+9aAKwrem4//boZ694i1CtJXfo5MCVL9jrnMURh84MjP3o
nToO/p/zuJCdG+X4y3P+VEEylkygPFkM/neKZy/fqwrWQMks4N1p00Hptw+F/H5iEDSir5Sq3Spp
GciVTlZAElf7Ei1yx+u0XGH9Wovrmqsz09PdpmVqeETGuQfk5OfkWyjRxwcSkwxZD3pWL3bLVmDm
HNaffZh9zfkDwj6xs2sTT0zS8ivYJONpXchEylGcMyTuRSXx0JYXj74ioWco41VJ8GFFwq+soBWp
fkBMEDZOpeSEDoqMFBdYxR5Yf3IQkutVodOU9p++/JnX0KLOmcWTb175Y6RLjqeXk9k7HUzRycs7
khvxJy9LM8KpIy467uocAcpNtxX51bDN+gjS9OIzer87cZpp7CZxo1J00lAD1inAn6hWBmYJ+32P
Lb/IBtsjqUgPE8glD7bwNdXK+9U2nRRcdrMnA3PkwQ/iLqV9QSw0UKXbrCoIoSiaRYvogT52ePO+
OPBb9m5IaVcxMhC8p6tFEG2j+vK+JWqZwjVfXQLcz3DvFuEbHJPkSjE1YCqXmiJNknGWy6wuIuPG
f65Mzgf/gNziYu8kz7mJoQRDLhueMB+64bToSuc4vaScdIl1kqj/Oxl7gQzSaVvdE+PmeRql1NI0
0z9qbHBN5nl2mbuiuNuVLbaLww0s4q4Lprd+Cq+5STna4SsSEHkr78yZyjFe+1l3oBQTcB5QGfmL
yhuyEmrgX88VcJwzMmYw/ObtCcVzKGoZVjMb8GjbvaYNXzz4ShDUN1Z8OOGAm4l2oVoMfJix+f8d
N0Be8JvQEf9MCmKQeh2kfgJJSr6Ign7H6H84sRlEASVVq4WfrCaewsJQfytdYfJEP7BEGURUZ6JR
RLGktrlFqvCegzJUvGvfo/ETR/fTrPpmqSQCkcpz8pGS5khLmZT7lpfAnoCh61G0OBdPCINedCZD
V6PExWKomn+xgVYFh+fha3EKdyHneRMfYE+rnhgCpY35/UpgyI3f0JJ4kY0dIkBovegYZ82xBZFN
w2w2aqkEQDzqqmiY3r+g2oDnEZBIvHUxuWnS8RJo4QRSS9LiDJj4H6DE39WioWNQFCZKOj81VKIH
ucj0yt7XsLbysF1Tl7EUxPOcWfJCHr5unXr1sXknfVlWb4uhW7tvZ5Wvot/3GioMXXCgHmn2fNet
8VU/25v7iU91HHwaOAm5KTkYD6IwGzvzxK8V/2oNrgpNq0jv4mSR0b8fG7zzn0OssNLJpFRsqDZQ
pEZgn1U9XWmQR1RpOePCdTURh6l25NbPNRTqVjrBmd1PqAsjzuIMru2lsK1BbWVOe4BVOdLMH6vY
638DILL4gKiyen8H91c7TNku17vHORdOkOMSIrtzbuBaYrRUTk+1Q6U1IKAvilu9L1zk1YUHT33E
SinnW5ErNS4icRgLekngCAyqxwnBu5yxqyDDMhTxPnsKaqDnenkIa0zH5vwDk/zhOoMWmUiLptqt
KLfxFE2gl83x6SqKdU6RThkY7HghYZanhsh//srCLX7cwDIoURHvC/sQWzKQr6yv71XHmuKIe71O
DIRxZND77Q/gwP6ZyVadJnBinSTkX/gPVgkqg6y5yoDIfFBiLRRXVAO2Z0C70gMJlQtGDoj6Rn0T
ok/dLZT+nHmfEBqus6BiZrwLzW3xP6nYT7KAz97ZxYasSdWEaXBSGm3LJZSJOUh2BCbQx5u1eEyN
1nkdWmThZC4IHaqo5/CKrpy5Xqj3xpY0VlYTnpXYGOYp7Gu86rqWrGRLWAwEWNihRb5SDGKaVlZN
xmJF6yE9sxRb/7ET1fxrd/qvO37S88REJZauyN3bsxnAgEm+JNrLmBdEu66JvwrtVMDPGPMxLOEo
Vr0Pv3q0E7Bbb5s6YvKGqK64+Xu8SllmmoSaVIkmGKkwHnuXxVX3y8Olkx8vvkM5amnnYRNfwYc8
ixJF2fEkzPXkpppfxuGH3jwzTJMF5FQnESIy8gU6+Su+sc5gTFiDynQEOBAT1lxmjbxARpHYEuXv
I3JjPh+tZDKclLlfq/Jn61s01kL/FeOlu/MmFeAgDPXXF7f3ja9zzmgYZvQheJYPTEYXRywzB5KZ
6QBSScKX8zq4DVdJrKKgZHB3IkUzDGBcQ16UYrgHJ2cP+HPjBEujqUAWJapv4qI2ULS/ksxBm6Mu
Vgx3Z0rPWlSZlt+0q741o1D5wnDwVkjGTD50v/AHEJBO4ZCRxzj3lEF+vB5ftOUMj2fpNTXQf5Xx
UsIlLXTbW6gCft9CKW74sh6DeySIa/zz7BNmI9tPu02oZF3X/QL5ObfcpU+Z2WCzx8owu1d55P4a
wiwo6isQkRpm
`protect end_protected
