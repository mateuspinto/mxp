`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ch9l2m9AO6L0RVxtn3vO5SKPg0HzlDCAkRDooKPlGJYQ2rVK4e1I9bgnuYgk/7RA9G9Tl8Qmkat1
5jyD3dFDmJWmsUS8UTBKH/4OERikXdWgz06EXwMvjD5eZiKf9RYm+N0+eHr4h4ki+C57fATmP/zB
R+pXxgwA/PMtecOGhAzALLrGovQlXhgbJsnAeWH8q9Sz4bx2UraXOzYHwUtDOCL651GhpAxzu79w
V1iNkOlrU75JaQK4mhw+feTxwlOQqHdRsRWtS+nk4gYdM5bjdz6g21TCTNUVZ+XH+2R0bdHYyQ4R
6TcSNdU63WlMVHixqmxefZxbd49d7EAyqboXWQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="io2cDZ82BdOFJdrBpmegF6jjDv2sp1wEK13sOFtOXOI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
lJkcL5792pOaEkW/ZmsGypkbPXjyNusyh1coRTOAFCNa9fP8u8pmuPuvOwc6zf2IQZU+tKvsJmga
F/dUQ5fa6LrxN62tJvd03ymki5QHoVIMPHoW1tgS1qVUuTGa2wPhooEJDhmf3zp+imYGlX+Q+Bzg
itOB58iCGRCqnSk0PcdWcjDm7zZE2RiFGUN66aZoH68zPfwtuhuAq0K/CZIYYs0X5YAbwpYG+NUj
9wSHxpaox7GeTu5htiLZsBm3emofoYHojFGNDBSg209vFQCGtWo4wu7psoC5iryriAKUUdXamPaD
QCaKo6OWEIBxUcWcK//jNmD7ixl1fpkLFjgK9yLX+byNmhzlt1rUwEgjQQRBncOoLUcG0vvs56e8
xvRfGef5SEkVitZLBhQT9Mw7OdFOdSVa62HKRfPNKHz4fFIa13AOrPy7jx34rT29Oms+OhlrYeui
PF4Y0DJ5CItpnnCvI1yZtbVdmQnkOTwl2amcP0lhP1pzHTsj5qZg4zNOpYUVxzvXgYqRHo4XtyK1
qveqMK5G7oyiZ/vjANpSe0a4ImdgXIg0r0YD7gpu13A+4PigpjZG7Fwpka7jJTv1KNRMKvjTyiNV
ow+2sIPiEuFZcbeYMcjTtT++KKlUjitjasXIRrU9pnDH0jeqN/3jObkjfFay3+i+eJSJDVwP0NSh
mxEZ1leYw2V+qoVxm2GHXPVvcw7Nw9pnWSgbE0Sk7Upi6/V5UlSgXoR6aI8a8qSgGPaboCURLgO4
SE03O355eLSMWPJGN+SDJ6F+4MSN6IhiJbnRYEkATlmU/gBr0q+ku2xBTwfJX3n6ZOlXfs8MHGk4
jZqwlzagZrxSBDRFPbTWTt+No8AerXkFDaLcb8+ZrTtE64jGMecnpdSDG0AwxBXaHnjsydQPJnrO
vSGV+xDk4GwoZLQORcXqnbqHodlIQ2kpiBE+i0swrrYsXKgm41UcuPX+Dwy8AW/CFP3mdNdRvWlZ
U39LH/GVtR+jU0Rg67pWddsVSGYkn+mslFYs8WdPND8WfTO/TH2Hfhcixsrx4GQynPQEq+53jBQ+
tlzJtstlpsIOxZUQdeYYLNn7NmIt7lmPb5eoef5cyAnO/Getm06+O7yqwmInASXR7Sz7ICkmvRy5
ASBHmioYtI09nCRziIpkO0pgFK4JuLKHeJd3HMtqy6II7pcQ+fa4zbE6dQ/ypi8ojj1XugXY+Txu
zJgEyrl8BHNtMHRZ5t6FA9+U/nA5AmMk/Ulbm8ZSmnD/vd2/ArdqI4php9UdWlku5yAufbBS1tiH
HUmvvZAWNgee0dkcz1PBJisP+lRq/9wT+S8D2dCbn3CHEFHAwepXiOSvkBuoMSJgAsjpPecrBrQf
PUkeeGw1YDyFJkTgTFjKKbwFYAAlmyK6acT3PdV8yJigZ5/uL0dd3FheY9+sxXHfapu5NfwwglrE
o9BeI5ufNMSEGEHEek45H2kIPnMgxog8iuCVmNJ2TAKUyMhUaXbVXmfSJy7yb6I6ErDXMM66v/i8
B/Hyb2cfymO2KMk69swAGHhqTOLM3TKrCYTJLsInHXhQ2y73X06QG9ppmmff+TouPpD7VFIEHRuc
P7NK8bu/d74qOklxLatRv+gfWmX0w2Tq+Fbc3rDmEL3h2qo6AmVqw+gPO3IUPWxJIqkGBT0gjznm
l7PGQ2Ks2Baf7fqiAqlbA9AsJWp5OALTNUN4/NPDZWb1/PZAqvujtTicwandiXLGn7utp59gYVrf
6E9+kNn6KC+ulcRpuefpTnzcLWgr6rl1HYehRNbQXN8DpAseJCw9hxQzavA7J/kUpYPmJncTibgQ
Yp/0hO+rWDkRk2Q8o70dh0SZ7P/JQNvVs0kLleYkFF7SrKsum4kvkYtrMePOb3jZhCFbj57+Lak5
6kUIRMYQUMEL35pB1VIpqrFX8ECu4ephIW+VwI7vk9hbXEre8S/pLCn/BmrlLlCfvfmw5QIgGz1Z
u3bqSjXKca2Ib9nB03d9NwAiD1BnqTHEjfgTNOnS/DqAQjyR4jxf9GiEobvFZYP1y0pW7COfMXxg
1S6C6zltQNUEbwbnkHhh4bKzl3VpccCEnbO3Mth0iXlGhbHmcjMd94iF7s8jehYT9dvWcFE/X0r/
DgS7gKPyTo05iVSv9nBWYFUbzB3siFrHw57L825cWrdimZyQSU4CzVZaESA3pl9LEGaKcngViZql
a67hw4nDkrA0wHzaSKvaeqGgi5Pym0nPFgSv5mXovpzKNFJgcr/6N2nHC8Jra+EtQ94yHV/N189m
e6QvYQ2qqHPdfHtvXW+1MU7W824aMovKTnjG564jr2svxkmDT7LbBHrzepdCW1xqMz+tPKPjSFYW
yGvQG4laPxl1IEf6n/vY6SDkz1riTX9TYZlSi3t2JVANlkru6pZapQZuhIExenGrS6rxFtCSVgNM
OtV+lFOqjNtlgzkFN2DNye7GA/6aEI8vwOBp8OKawwO2xNN472r5vgiecIKLpl8eInRV9HfRirKT
jhxCs87ySYG2LhhkVWvmJm7uUcV/0SePOemCKDb1oNtGlMSMsMAzbcWRk6ytBiVzzjEJnI3jIDoP
XmxdcnzEwy1xWelwr6C1HfI92lVHdIFWbJZVkwy2q0X+wejcADnaekJ1mCnqsotVa16zcL2VDK3p
RQ/MVDrbKbedBIbPPGI3z/V+2pNuLdFgY8VXjMh5bWP/FIfr39sAks9Gb4l26gTur/VIxjItZq0J
Qdj0CBBIsJwpnr0zn7G248fPxV1lsUAh23ui8WqRebiavB2V9z7R8UUSImyCLZX2CE7qEgByoCWP
iFhhBMuZbv0CRVNsS7J88vIlM+ka5LvT7qqBo0kdcITwU58nEm1pAf0Gd1xmFKBqLLdDTZatA/o2
mzY9dBFl4W1U43bcMj+5r3MJ2cyGoZpKHZVNa2J4aIh/PZF1PjBrtBCQtgostlDR/clIEBH1BlH+
EVLgFpQoLtife5/HUb1V2p/copvZCIS0zIPyzsw1+mFZOyYTPfJjt0Xt/9dV64CyW0sZy95WFIk1
yDJcsMq+A1H4/3juv3p6Ej3j/CbHAa303wtPSYeX9iw796e6JWYyj7Na4lLxlfiNfLn389T1jI5J
QmivpHTQvAqafGoSQbQ1pTjO6lDuO0ZWbltmIw2QdJMyvyz0m1MWFsq4owov3ebB2dNywubvfDf9
493A8GzB5D2s3NzA5Ctk/gArYvQZuBvd+ysWEvmQNkMnrYL2xDRlNcw6PanrREhATeDvURszT2p/
v4Ibb1kc9F9tvtLlpP88ZeNxpzMNGEd4oLc5v3g2z4gugIYZG6eRIhHp8D9p8myZu9SO4yOJVWtJ
zs9XE125yzOW8oa0UOVPExi/wA5ZBLXZeYyDAzmRhYKrVbYKzVMM9XVfJeHB5cNKfnUT4XvojwFQ
QeO20v4h3/MrQU/5e6jg+BgKsbir0e+pejeRCYLj3wnnqt236DjUGbb6hTRgJNlgytqAHbSxKmgC
N3iwX7JQroTkKUZVQi1VZYyDalGVlN4mhbcJaZgKlmWci+Pv+rltr63DUv8CV+9hlC6E4mProkz3
oniBNJPa/2zV3VeBzA/9A1sRGdohLOUm7g9f97Ww1M30OxDbYDvxDY4e9g6BZ8tADtFNpngf7obf
9jSv+UyUbTOg3Jva1MSfrWewyz7p+CucVUpxqvaxBi9WsyvhFoGfBrcSFYKkz8mGuHfwnrxnYS46
205z1j34po4qQWo2FHFO/NDg7X64E48RikKBCw8P0MvDvMVHutCHJ8Sn3ROCDn+6Bz46gbx9SdnV
cgTzWYbAJzlj0qoPhy+XDR7BeyDpHSLMnuwFzp7dvfrLfIiForLj588ocPbKSK8+bLFOjUbYorzs
SKfnSERHNq0Zx3GWpzmSpYv+44LrldoIQBffkW1AHPmKmEmf2FPcyT4DbBuejmtxqhJDvlU8ooKj
vdywI1R3DfppwHopiYUWvD4ABUXJyuD8g+KrqC0HAeoic+9TictsA9yDKeYLG9CpansZ2ijZ9Muw
C0w3xPRRCRBrkEyKN0UcXrA7gzFy7r+N6HywG7/b/v3TMIqIxUA1FY9DhtHqqhlEeJSl02arXEsC
pszMF6av0r8jFB/L/5SMsWNrKzl9pZz7b4SxdGQerk1/+H9/UlSiK8LpXb3gke1ROCS+pTJsBlHJ
zpmeuZrG6E7BYEcY5D5VU/gz0cOA41TPAbI+IgWty4Lu1DHh1qhoLiYHNjP0oBRlZwIf6E6Dxpbw
clgp32GDf5AWPkO/zJwWaa4oeMhnmq4FATxFdcMYeRUF7kXZZpExmUqIJb1fyeBd/bZ24wxiZ/0T
wAFS+pw3AiwBBVXwL1HSQSw+RUNDC8Bl9lHFHGQxkA6/O7q+AppiUnxkqLjMcocWVlqLrqsM4/ct
la7ArfAXyy6Nw3K1/8vxlo/cvTgCO58FZrqT6j/ahWFdp/T2XTHz8kVq5Q6B5R16RCnNTcG+7ymC
8WXOKkk4t+uekjQRcc30gA0DGilsPM/dFktP2+eFNBOFDA12/XnLuCHpu4rZFWeOq2KkMkIe1Nqh
WPKyfHouH0+oeZmebI46SL3q3yd0m/qRgZOaxmkU9JvgZqHcuNYPn2xtC45DtReu3wJqSNmGKIhW
oqMzjDd3cC+RXSofTrt/EMRmXXbf+WPaRpb5yK9t1RcrB1wfOI7Z2VbFdMUvbyINqw8ARg6hvnTh
mBUZvVLGDCMnJVkDIrqw0yYgE5JWKxnlAeTa0qH2BQJC9zR4MAr79uAj5wVUSD+vRYEt3OBNUXwJ
VvXxSgr8r+o/IAD84YKtdG8rXrtF3Wmr/gB76K/q3KTtYv6xAF6UxjCMbSYOCDt2kYmUIAglwgLm
HTRsmJVQ/2KTuY8fRRkPY01kAfZlsm6ydaos/IaaogIaCyXa6jtQn39euP50PUyIsE+T731ZF4B4
YmEPF8gqXyICOYsjDjVrZi1ZsC/9z25x3YQZSzwA+2tMBTzIfJVjKYhJItvW7M3cmOoX4XQZQXZW
/eoSRCyxXglx51HXSnym2eX5KBePbwZVp+vcDFLFsstU1eWmxfdENFWIodGPxqwaoY8uwXakA8qJ
nTin+Fmecx9Ai5lJmKp27mUEU4DL3B7D5jUtz8vHMlWx5AKQEuj+tZZ8AXMWjBEY6Kqyr0GA/h8T
Qbc7btdlGmq0iBo0NdEMgz0sqInCWEVdiCPycpMJW0cyBFTaXZ8GODUh8GLZxlMuMJfZKP1qlRM8
oW1pBbmALhKZsKtrERXFV8IECJo9z5Dmbon2wvOdV11TCLl6gdk9CA3BjX/bKbunfB1TMJMQKZYv
aqpFp8J1Sud1nPrCjAzYy5PDaiX6fxuCiWGtkQv2j6jsQHCRwAomXomalDu9cU6Dl2YVW54W2oj8
SfO/zklSYqsb8k+/peK04e+qhP8tUzbEE5m2dsoQbGLfg/y4twAU7ZVsABmuKR1NzCfEn0fw/Ksw
kbS79gzN/nTEebmEcOLtubWUJPMh5Vn4gq8yoMFqLy6/eIjPbGGN9U3jopqN6PhJMVLB4mxb3+5a
XQdPUdhMgCcKpinDUbvzKvCWLDjG2Alb21dxT5wrK4vAw9ZUGB3oxQWQGvXamj6gTz1lz05eT/+c
8w9GcBLEH7QbftxHokZkrMITu1VpeWLSLAuPgwbuQxcdZnteK48D6VosEJg8BMtAGEgokrRAHtgT
GrlHN841Vt42TTniUglbbMNgYNgAHu7+VR044eqiA6/YAsEjTyD1fmksArmx/fPmEsXPZjZhZKt2
q+6w1+0qsyb0+M9e6nx7MOwAXU85K/X3ZwsLiDhn3H/8tZODQbX2X/DVjzwENRJIpC1p5H0yHVNH
d0p0vA6aSug7+zPWwr+WyA3/suisnQDivLWwQW6A+6phCTLjXJUDm8Xre76yciPT2c/bbwbHN8l+
kHZPt1k8Cb7zp/deDki+t1d9Nw87X0+DohzCNpJYhBmfGlI3EegoNrgElF9+dAm4Y/FDOvl54nrP
TVbtwWrXYensv0AS/utxRLDuR64vNQ9XsLI48Jg53qDPHa96BHa7kptg2lw+7DGOxrGXTx/+HLmX
QLBo9KdnNFimJUj5+5J0weOM5+01lv3vU4GNV35ahekJp4d7C5NgXMf3B/tw8knysOERcfVds2VP
q+N06Zl7CGbFANIO3OCC8JJrqF3Z3D8xuEF4rB+bP4n/TAyL8WIKJR1+z4ldzf4PVLCxEZqcJ604
9i4Vb6PGAt6K2RsGgViGExMtDWJcaa8FIWZEd49j5lA9k76w8x36cCnnIFQG/tAC+w0vFRfNAwzc
3a54DzxgBnC3ekILyTkiJqFgaRBNjRLv3PvG7v/26/3y868b/0OIFOHWCllvwhiFb6oZ39RPQEhC
Q/WPtj8etQDx1IiWn91V7Wx0DWKEqSiECqM3SezC/P2TrYfulncuDLIse4xjuZhqCwiBJb2vlnyQ
yY71yEB8FxYRfoexfsAOt4Eku4YkjOfT3ebWSHcIqs2l8Ltl6OniqijG/G6RuMhE/NCd/LBgQCIl
UQkNgFOklscudo0VLk3srbl/lroKlBqDVRIM2Gd5jdo9IrBVpIx7jQH0c5t2JhkbI5k46sw/AUQb
iHAdoi4aDo/cuAjPEsOQ375wAnOZGJfr0DhLRXIjyHEThNclHsmdp6NOJZsv1cMNjs+6AcVtWxWV
sSKC6qWa4xFjq7rsuZAWQM52RtkNIxKuBvxfBSIbFXqeUmsg+NtY7apfslQv5+ZLSXCYLXWy/Qmc
h9/RaI7RZwnXPSSiSe+kleqVqRhF/I+8ddzOEnrN0d+7Wb6hIqVeoUvumbPJVStpZYoH6++fZMY2
3WipP/vz0/f4UvCz6786hDfx3T5eKZiIoe8F4JUM16N6EbTV0IedoB6eUyKejRTOgAmjBLbTL5ZL
xzLlbSJfAcCutjD9mxJj8kh2AJQarC4e6Wf7ScxgRYp/9hShKXCLSDroT+5ZDu38Wj8i/4WOB7Jm
bdkJjdnBiGzfSpLK8VN4Vrr9xcY6Nay3plE8idRnmrrfq7AANYODBadayvLstjPw2rEyVjasjlIO
YPep2h4ZHzRZVXIX5LHfelRpJ50XkJeNF40IEC6nyFPsihYa0T752WQJjw6gFfi4bnEoylXThIPu
A/avvYbhqDhbvQ5Rbe3ljp1pdZ+mQBPuAEAd5iIFsdhp373zRe6RoIg280zW8JdhQqbdIvTCMm6p
wGYVLxD2RU422S+uEHrsWIgdp11G4JIHflaB3zq4Cv83h8ZNTJoFhazCCfxRcCYvl/m49Y8r/Z+k
VTY4IjTsu612R3812rdfnTJcP4B+S2mGRIczu5remKvN6G5q8Xe168HPNwZw7DOCa2BuqKfGkui9
XG/SCmFfaocoW844YooM4B1+O1+uhC9JQYt3xTrapTOqwTgdB8csSrwgZW+BvWvsjTU2P1+odv9j
o5iIgCHD7O5DmEFNOqadaWg4rB6U+eF2HDZloWWu9I7vu1gQW18DsbK4UKG/C3VIvmt9WG6VAxCN
vdo3K8hTpAIa2alwkUz8bamPDHjKm7I5TCus+J3VLIhpziSnxRSPmxTsWhhBB0hYqoGhpRqHZ1HN
4T99Mk54dCUCBwixWUP1iGPJt+k8oEuZdpR0ofJpB9Lj2VS63bY2aKqTSsDhOKYsM8M5bAaxc+O0
2cSrJLWDTr5fgGVTAsWhjLvD1ZnEfrADsbMf8/0e9bL/ohXV8PtaRmj9kSjSo+OtcWnR73rblPmg
QL9KX2wbgFozvZIjVJxVUzK9EZ/6E5P9T6Fqe9p6FXozQxdhnpva1ODSanxAuyrnvB17/2Lq7/wi
IqVOSZW6KRQ+ATLshG0yvebY0W+9t3on0XNXQLtIzEblag0BWvkTuTFkKZqQ+SxvdLKOtoKU1Luz
OYuxdv0h0cR1aywkMQheJ4DBFro3YPbYieHzVEOgBZn1+wpwsJm8dCrf+rXgJCM4v8tlkDanX7+H
LTZPRKdToDqqn+5JHVcfM1U/2ExF3fG7UvClFwUC3fbXz1YH1uykR4USLRcvIfS1pduL2qNrx7nS
2FebVPZExqLylasvCijFTg+G4O95iPrTNJPeKHIlr11zBx6TdujHe3eDmP5BqiX2hwy8vSuNG9bx
5A56/fA1Eb4qfQmWF5j2CZVBX+slu4jED96DaHYgJlRZvdT/K4xL2xxz0+E7Onwb1dxvxjaTA8JC
+UKobaJydTgaP4D5mIt+YgeJD2+ynTOVIlZ6oZ92MXNNusZASuM7AgRanWpBq4mz0y7bZVF7f1pW
3Dr8MJAkNtc0I8OwTQlOXWd7sN/Nbh4nLJpwp9l4QoxKm9ha9BN10yQ7JCJkeQawGYkrtpEyEZMw
+CXiZHu6+6cAxA4bSuaXNQ8pu3xcKsR3hVhJBEF37Yg+CQ453hfNnhrXmRrh0dOa/g6Oy5xSOoH0
9P/KZ2YaqamOCnBNB344Z3neD6gF+KPtSDuHeKTYWZHW5+l7xNx1Bvqtp9MlyrsJc4ZPSfjH9gwH
wBjG5uAVCAE1ZGcVWwzDci1mmVDFCpy/ff9GQggmzSqF0JRg744hIyPztytoB+1r2Fkz6fYf0683
bptX+ZjMjED7sUSh7i6EDL3hVjd37pQwXUjZ4fwQtGqdzWy6/62bH9rupHThybKG3O5t+xdgSn/B
jcfXhqB5fWYPmYhVGxtPTg8DTzAriv+8tkK4Ngzle0yGvKjo5Q2yki+8FvXt9niGTMOtkeaB4bir
0eP1TaRreKQce2gsGddO57XemP5hm8TrTI+s53O2P2SkXTkB23UfRdBF2cZtkKsF97rIWNEsUaB9
+Hp5FHXhzrZ/7FIsDiTKv5augeYp9WkLdoZRp2iiNxClDSTqeXsbcWeTAzDoGjiIZzP3SwvgZ0Qs
QiP2taNM+eB3G2ktxfpcGruEMbz1Wp6VyYnFcTFvVBE76/ZegBoh/8r8NhDoqDf1HZTe0AIuLWgy
JIWRncqXwc1kckKs5IgxM43RooYFa/eyIMSMqdW5psYcZniylWHn88A6F4pxJt9Rh/Mas+WXP2QO
gfGKqaOkw/HZBBkqrvWNhgwdfjCNc/Jqoz5PTkpgEpCPeajFde1aA3h88pwNINbpdHMV+PUfbp1W
STf6TAk+z5Obd0TpOb8MF19XxO6w9qzAiUnu9slDIqMbo9znsiXJ7rYEFo4JKHwe7TxcidVxBg15
h9wNmCtWzJWsDqfp4JUTgvaO4eagLzDGV1cGq/fimKUAqtG3kwIPtR/zB+sMGqbwsOKr4Cqz/ihD
hdJkwOuPLLLsS/zZv0dpaK14iaKuJ/GTVdFDLkFCiiSx4nkZxWi4FCQeg3ZcVDL96hicgb7y/Q+Y
6QEKkwAb6sO4f7qo1xBi2D+MzGPg+SVYssbyk1L6mFjMXSEKTn5njTAgN+7wltffTPTYly7rNtLZ
TDDHrku6nS0P00AGWxzW2rg0M/KdWFrtPRZZ0M9fNckFBKvw1qeHuWyHbJo6quA33l9kbmSRdbQY
XYNCyXk6ac190uOI2Xv9wydK2nsEQ9A22EHrSlVbCyxeQUiKJ1ukBX2rIhHDiWnHezzeRsDDcKSq
ExD/pRK0eL24tAkEcdBwSa4qTm0wLI5w0iUtPwGgl0qqkX/FXS7q4W8xftLlbXwiS7au9s022NTP
HOJpXyCmvGErcScctJXlOBOY6RVy5vBzAUklaeqbcVhgnKYpReDWxwtFcTuWE3BGVeVGahwEGRfq
JcaNoBNmz5mCkYZySYUzSRmeM8w8t1KoUZZIXIFQ0LVCzjp9Z2Pd0IFWpX/V14WLFM2Ay8Co7VVe
oiwzv4s1coW1jumKfdQ5/xvpcV5nepF1Jcfoq8ABI6EfDKPFBBxairvulmQtx9GShupX/UhwoVwA
z+H006wD2XRcvPe3jg14q7L4One42W8jfbJr+pqXj6jtZ92kTmytjYuwQmyWX0O5x4BHxMTazcrG
pMXSH7gwc/OvRMhyGLird7EJBTMxDuHviYPnKq3luHmN0K5GPBS8qAyUobBWBQy91sYC3ZZQwDbN
A9W0MSt9K07WvBvWffY7o5M4D0VvvHFWPdghynoyVJGDvKRlry6+pVJqMMX9d3ywa/l9kJlZPf7K
SLIj10ORaI7WP2FBMWq1Jg+M0TqTEh5DZzdsaV/IT1DZFIu/yR1l9C6PjpgOe8t5dedalEUgBruY
RM2lk5S5uPycmGGr1iU5LG9qgIOnzc1hMSH6ZjwBz70sModeVpd40asdIPvGnXUekT0FiGeBPoC6
48nIa+EaWYyinEfc64mnwUN2zbHCyGBsjtQnh/NHc6fYjO4Wr6S5rK6gLrpTOpbm2+V2Yp0a3iYv
qikDoyNJZHXx0zFigzZNPlhrYN2bOHQBDhltOrikPnZur01v42B1B0DenCuJun5UmiAkV5+AsMEJ
z7xiesI9essZ0r17E5EGOgce2YPNALjCLy13QQ+SX85jf5+P2bNB5m4t4FcZvaSLaqMmg7UFYbfo
l8RrEQfLC6mhZYH5gAuVmx/faGFcrVl3drZkn7X6O7o5lT3HPAHE+e0S3cwn7jhsM0cHmrWre9OQ
QwvfogSMXFaicPhvZvze4OGji7orhaAOCcK3tZCXyZghCaLK7JZ8uaXy/Nr5ZoWWWAP3oLjCYvV+
rTg3+7b9Tx6dXRawEFQ+kHnsEV66qA7giKhkOHzi8PQo3XFu/Vobd+Y0X56PFGTRwzQCWyl52NMr
hmLFSwByN35owbBJiR9BCZKKW0QMDGyqPhhqLpBaGw1ZsY+EDyYiOx7rLN7nEy2cs2b5bj3CnUTc
1EWYcqomVcEkXKj9bMh1OX8c3LUCQHUsYC1nOd8+bTeMEc/dJ6XE4EsMymzLPEdMjX7ZueKZVLR2
IXXN7pCe7NNwcoFRbbJIpSXhtirZqBfhjxIq/emGL57Dna8zwZuC4SGssPV9CJOKcG9CmjaMleQd
7Oi/qodIBHn7pLGe+MiLePxG/KGh7HCmX2W8pmLM7SDIHvYpIeKfdgFSzyjUI6eqOT8LQCUpKAqq
SvkL78qXgFko4u1IGrnrFaJskFaBQQqSzHhg0zWOo2n5PUnCD9AFwFkR8PVd0WpiVwWsAH2LDFZL
u9oY20eKamq8CF5uBrMXk24PGCuawkZbWKpmtFalH8psVwhI3F0cTl57ri2BnuY2BqHTrkZAxsn4
Gptx8MP8JOJ32yVZt9CskI/byd3u8CdlzgWGZMzJdSAyKQKmkuouAkD64my7bOa3bqTvSQQiFfoW
kWuydD+6JokAyiXzY5CFK2oORld32EzhAlDezU6znRkcPWHoThcAV0lUGqp/wovKFBvpOmf0spFP
wjTgBc9HRGC1ZF9g/l2F6XEQQQsHefEqRcw5cLOWxxdsE09nEIs00wgnrpZHhdFJIpZ+h6bi2GQK
3fbULI+g3Hg021Pn81pZSg+7ivd8eowyxPambyn52uyjsAQ25Nl8Ihyz+mPw99Pu7Z8hdDZL5o51
23H4yONmNY2cIQPGBnWALPf2ZmjZ8v3poZ/b3Iw2kp7e+pB5aQjy86n4M4wOWGDPCOm0+QP7TjY9
e4rWxAKWPRDkHDXh1QNsL+vRoWNHBtz2X+mxiSvU3RRPa3BBAWjRwgQItAAXNLPe+UTNu6n04RVw
X+A/1wf4pgvTVsNMPGX0SqP1bFjLeu0af1ljxiJ778OQho2FrXIdSCPH82weZcPpy92qoSO3suh+
hyZUHWauUNpAPy791+TfORvcCEGFkS9SgRTzFoKr07ISdNPY+BMBj84H2MIO6O6lKNAyIXpjkAeD
8sLlL2HKR3TnPrHWOOukpTjHuRy3h0hqaUNXoERu751LyWGxqvx98xAju61kLg+pMUABFaiKHv6G
MYdV7Zd/HGjPEh9/05g8mFa6X8IW5XXdxac6tMCsiz0NnmBJeTlAcp9Ke54EraPBjDlxmqgDNFzi
Zhaw8GP10qJpES4C+sfdgu004aOqwEs+fDTYD6HfPt2o5DyGqqpWpX+xrmUvVXyejWbjso68YGLn
fBY1nfCqbPQVz8SnmMp1a6/MQG1MjXKeCoPP4WzNF4XT71szeqWP1J/7m57MRQB5zxN6gT7E5JGJ
NvH7wCiFE5RuCCLp9n7vMCI3cHAxLY7txP+eKqQMVFbj0bM0KfFdI1fhWuI/Gd2SYrxLaNZ2b30w
XZLlESWlopa1y62RgPbdTzlcljfD5zcdL64yeL4VXk+6BPGiUlGCr2RvO+0+GLtC8CMqp3rIYVXd
QISdpfzeThFdkZitmZJ1vMUHZuoVPnN59U2HDRN3PBPIRN+8NMtHiz8N3Xpmyd9CD0h7/kIjZ2Sh
qww0FJOn8DBBgWXRc4pImvyNoTApshvw+IvV0szAvCX45xoyDc3YAIt3fiFkWcm1kSstIqx2RHuc
dDEsKCaidjQ5OrSXeT7eMsfT9nFgd9eBHOfx76wd8cfKD6Oibp1tOXPkbQLjRqBDzv8w2XbBfrVW
3J44IA0SBESkHMeBE4bsEnxvsttG+i+3eqJIqaTqHXy54oVdaSHL21PpuIpxg3jO6pjzBtxRNiXv
9GhXKDCYbRgCScykaUrGYp8fnF123NA0MtgxDmVHYST70Nk5dZX4f3m9oyLmShgMeqRFHnXJOwII
KzAGKhyPo+cskIpk3Jo8hfVv6TejKVeleaRequr59XgxoLYantCFHhpkLIUXU6LgGvPBQViNbo+9
vCNHoR1Cn2wshTgZmYV3718tWcR8ZuegdkBtzURywEcMCyjduEpM1XdlGdZ/8jq1Kbw4LMh2qhuQ
djRUtKv2Qeam+TOHI7F+Nfca5tO/BzY4kEKZdJCQbPIuPSRFyNpBCrtxHnG644iWMlWPf3mZoCkI
pUg5TpWn171jGm8Esi0TT/mxH9PbErPPgSe45M3dP8NaQqkSn7nJ0+ev3/XU9APMJP4O9wNhw1km
IpCQq+Jr/gVLs7oxq5ci/yR4yRDgn2WIrMIPsMPf93YMadZNL2oDslotAGR42aqjNBaXWMygfbSR
i8j5cwamWSScrw8SP7mPgGSjlOus9i/flFgm6CQhXAmlfxY2DVxyCbeGam8IZgZi8KS/3d6utSzn
NbxJ/qZv33DfjdIhB1JSW0lZHwi1nj3ocCmp590kQJC6Dyo2yz46V/gol4ObKYipgCsUCgFkqIkF
Sr4rYw9uLdOCCHox8JAqrCnRJ6fF3Htp50D46hiCBBUrtPS+t46dk9eq/MQKXhHt01esLetD1MCL
8++TpwyGMs7vC7XxXUqR0QIZtJwxiWyQBr2l48KRR1+E8YxZZhrFSfFMU0RxUxwD5jFkrpipUpbr
x3r/uGOyENVx+TrcT2u5Ezn8d+R7jBvT1VOCfP64jczb/FjreLuzsQXoy6waOHl2z366QltWtSTt
WZurhh0KHj698FjXSOjCE6pcxZ/ljLVaD2KSTRJbMoPB6NQEwl5KxFHEc/eZeys5Pda+yUXsg3Mc
q63mEGtp494nrZbb4eJu63cfvsmEgp9NSiwcMGUTW3s2eDGgKUP4yPHF6FTvS+SjSMGtXBgsKhgK
n7Ni2TrB3/eLYVhvYjySR4a2JsbKt73pZPLC3pl+UnY9ItkJlqK30y9bbhN6cH56Xx3DVVXzCJSw
4YVudFRbxQgPgsdETiu/D2oriMtFVPLcnuDXonsWaV8Twzoh91tOpuPSlroi8D3vYcvHAlbooqLO
an35GrrY7kA8gaBGqEaS1sauDtvDw1f3CdJ/7JVi1m/n55qsQlCOc78CoJMMZuB1N0y+/ZOEF+UJ
/leWEzMn4AOnjgEZKo+0gjG74/ZYOaG3/6SZY/ZIiyNXHgpS2GjDuY8WTpRUetzhhyeUHlmkc8lR
bO9x7Y6rRs4Ndf/+/2kQwaCB6yPphYjMFwPOiXgje1nsD8GNRfURrkXWZsgsxUI/QE8IXrYTDKEB
ftewOkPEU/mtXPWLhK5CVEukD9gla5MR2j22F82rgNiUPmY8bj6wnN7an+cvY2HrxM03XewtQ3XE
cxq2IpxVnm4y2PEPKd85wlY54vVStM5Ze8KkhBHbrfPVpbhumUH0F3exvwiaTg8SxgG4rWatS2gn
A0kCyyMTlQ8rcjBTkbodblrwNcVIojFSwiAB5MiMFMRHZvicKsJ0Gv4bX+Dht0ZT4+muoTyaacYq
on0RkREV6JCftBMw8IvSF8h0DPmNrH3bE4rxZ0qC2lIWgPDn/r0H45FxiEweSKsgZiCiB0tD2dLK
xjXpiNlYHBB8i5h+8nfUdgu/wudldDi0vnlNsGxnD6GMR/6k76dBt35b8+REoh5HSvNjPdYnPcoa
KHcExi2Ca8Ve4gKK3c3QhNjgFI3h/63dEiY8uK0DngkapeGdzhTjFI5197ZjuHefhkBlf4/bNooU
MlF0cHG9n6XCrDeReBt2sdjHzol05azvQ9JcKiTljPoDHtv3SP/3f6xqwvq6GvbFgcpYDMw4vBb5
loicBYZIvHLJwN0qVh7AHkkVtCrsnJllvb2FC8RSz54Rg+vHORl/b6lKN811DJYwZFITYljs3IuV
sr2eKkbMKEMcownyfJuy613QGEbx87yb7W5Lj5wtshPiPCThfPxDIS/Kei/VFGlpXUQtaiEMenh+
7Y9Vpr+21L1ebECV2nA4m6tVbXebWTemlXbcrr/9N+ebCyhZ3uN9tAkPQfW1L1Fu0RW2yzAlcWQQ
ZMdEA/bZxTQkpfMi+jUHJ7Jto1Me5+eH0NNBGDbtccxunGejkAoidUmIJaToAOY3z3nl+KEx5lDj
T1kQC2vU7m6XqsO4ofLpA4ro9KcFqJjk7m8hiwnYMrjQZ8CuoTkWrkdE4lm/hAMgg/r8GMGjGdn6
zKkLek/7lnyfh38H0QLSUGnsZ3ZHmOkUqWD9jiT6Cy/2MFuTiJDcjDZkTwUCfxg1aebf8HA6/hG5
h7/CTrPpXdT7S6SlwYZOJNTjGw1ANEF06CtFKShEHj+i9QNCnm++Dqnc1coN0Zbc33jx2/95IBrS
+4KmZKku9ShhdZyTLM9y0Evg8fjOtDSb5fe61VL9SQR9eVXJcrggjZ7qD9G+pLZIYAMFdfUFdWen
F/DtUkvkSnmE2GkJMUwkHCy++8Qa2vCwah6M8OQvWSdy6YlnaZdqtAGZAkB3h1kSD1ofu7j3wKJ7
kwiF1GOcUCpRii4Yf3hGuHHPNfyKdfxq2nrzVWVNiEStp8PZQ1aoPAfE7OXDjbog7/8FC8z9jCz7
UM6G0/7HhIP9LZCZD7gzA+dzyAobmDUzY9r4nQIJvllEspr4Q0tPWJczi2ByHABAyoAWDhiUz1HY
bcD4jjbEgeHU1TlOZnDtGfsbmlHsksCPP9077d+KN4WzjOkr1gJjxHAWjDlhrnnt00w4Ur6X1SG/
XOIWzzq7jeVi6G8taK1yqishIRGjy66pmYp5X8sJx5jKYq0INvqK0RiVBVTU75gsGmIWz0eYEVDV
YpoKu9j6h1+fwDabjD2PbPD+94iZw68f17PHFo2Ge6orrHnleUOV10UqIKpbSg1ON0GVu0/YcR6f
Y9AyI63Wm07fFqaNnuhj0CjV+fh7G7XNGHCTmftfUrNC6o2M1AByIqxI0KzlykuWYfIJMk33IU7D
7g6p7PPweBd2cjnSCLHF0bLq9SEgvBUNOLN8npLPqWPstMWl2egL2S0Iv/prYPt6XqCPXfti8Jjk
inTaRztTVuHsK+ZFqIycEaLqufXNizGKEZuYtypBB0dN+mp80p8rsBk4aQx8yR9CLl8Xb5b/AuAU
iJldSMK//FOtyp3zdg3HKAfjGptdsl+7EjhQEDcVTEXGIPEV2SCRYmROTLGQ7Yme68qROd8YhESz
9hFHat6l57FQl9P9pcU8j5afreVGd089q7z1PAn/fqF96krVfZvWqssAuhq/uv/azy2wf9xWkP0I
FmuTmWJZI8hBP19LxE7pIjvhJmkXrwyT1fMS2XNzmxgkbzmK/8W5wmQfBsyjPxl2Zv56zh0t/0IF
f70i48B9MXeOcOyeb0yvurulZzMAoByPB4hqPtguFcvaAj0wDWkPToS0CGip9XUEBVl5kBO9oXfq
U9G1zOXu13UGTdKa5Dg+i2ZvMNfe8y7TEojEkzlScreOe5ymz9VvQLX1u11V5TBhJ1J4ySdo9fTb
iEKLmZscczur2s5vwCa2iapMAm2x19xZ2CzMQ8j7rChk2zFcYJ0Bj73KRcgsOTG59CaWbfb3VFFs
0ncu6w4iCMIvxavtygIR69todl4SwEWm/xzP55ckT2tCTJEer3wQ2XJtoEn7eFSfWaRkMwWnAfD2
fGo7ThnWMqsFSsMU6vQoW73xrFcIyguV0DuNxQoIUcAZYvOl6iaWX057JA8qt49MEbc4nMnez8Do
v7tGeH/DxxvkLHolSkNe9jfymVG62Oj7XF1GnwtjXoEHa0YVq3uDE3+8Vxfyr7ubdrwRzYmHkupw
z6oOlvrn8WtTBiZNk70P40r6ypq+UkcCMQ3R5tmy/8eh2besjlHX36zOw4zFwPNSPthEzokeihLB
3zkwp1tvSar9e5HA267fKnZJw+EmvtdMDaSThGHB143Vl/q7PDMCHJPkM+pmEmXQ4PKOt9q4zJmZ
kvxfE+BKELdptwb6KfVuEa8WeQXHekSihxjyMYh0W99r76segechHRAUw6MmfHksoxWeFctR894e
TpmAK+kDOXaasV8DdE5lxLcJ8cC8h62oMnS0g/o9TjXIzURkNM8qDWgw75JySn6gqpxEOmjXXHjF
4S2pGMpQnVzXIXvczQ6j5hihtAA3Mr4puWYmTCPfo1zqMH5NVASR0tZhtBTWTrBxat7rRqK5UUMN
YNX5huKmHtdtcYZAxMYY9spmgRtqNJB2xPerGxel2p5Az0P3HnqwCDKtkfW1oqnmt6D5FtenxXLy
xmB8ynWM5SjZFqnYv9EKoegO+e1GGH0DNbyJvyVfEZ32phZGToYPKjM65/FQG+fFZw5YwYV/CJP9
0vCr2bdZkI4uMcwlDKu6a+cyWe922BXrzFlGgdmh0RSFk3tBB/3Jhq94eVzbPDw5/ZAOEzCj2LJJ
dSG2Hv05ZJ33HAeZvio9d9JtqIYfPeKW82aoErecgggW3qhaYbBraf/DZD05OOodDLs/73fP4v0O
hhoFW03hwLEE9EMPDv1szAnMXj9LUo2WLSOiPuMwF4ZvMKaJ63i1pGGveg9lF1KX4Hp3wrmlToLX
hSaqSu6lkmH2Bu98jz4Szs3xQVECLv0kp8HRevxHtq5CfFQQvTp3thMpfaWDWfT79LfG/wMmLOoB
w3HKHjPNGcpZTrNQmz/6fsiwKQDfg0FHT8o2YAwJNP3mUkznfxxkF/PZo7WU+dhmRpPDJMb8OptT
pxWnOm0+9xup4Rq+wVM7wvxLxGHy/VfXo3XBMDAupKLSWC2kiPBHGvC4S25c+OvP2YtSg4/z2oGS
hXnfUKFAcH2PYI3Qkj5DXIXHAS5jB4kzQ8paJy0AWHhG/jXhxaDGwHz9anFtH18gOns5jSuy55fW
NkNbBKnR8yXiaf9n/2ZhUAm6Q4h+m6j0MmwZ2/VSrCDqRbRADaO3w05swG8bBevLrNw3VuxCbGt7
2cP4yXm8OXVtprKvb9936Edys5OpBY82PYWngLEe517P1uF9IUgJlElUo07ag5oLZ8M4T7+xXVum
Q6Q1BQHBKUENC+cIXjHuUHCXaXT60jY3dSDGVKsHQSkA/ljNpDuOgPMVhuCBmvjn9uPcPeabMfub
eU+vP6WD3GQAPBCJPUQaOPu3GafdiJfRj4B+e/8GrcBlhJD6qWlowCRU74MgQDpwqCrME23YQ5Fw
MjkJjuD423FcFFy/ZlLsZrc7l60c8vHONrzf8N/dpC+ylC2FtXyem3PU7io6mB41/8cy7D/qo1E2
cAN2f7W/0hbAW7TQGIurJfOR2Z4lGzklZpd5WpMTYm0/GkXqy4kOZv6Xgcecz+M7ySPCnJLRUqQJ
beppu4l7SmEoy2AcitfYkd0qb8dtpS6trqCrmCwsWbimhEhpzQYe8/y1Zwb96k6o7eRwzGpvZ3QF
VyRygkqHUBaSKcgR3c2gXKRVfw92cCmpBYQ5ABkZlogybQoRGocVAOFVrmyJZfWZOzaxTGHfJstl
tJFV6hWDPok9G6XpGvGJsv3qqdDYJORCRolLtRBoaoMLV3v6orYwhcGGbwidggQgHsPnhVXZfZkg
Hi9oz8ACVtSbqqoub57tmirrWNVj2wTu7aIdyDqpvbvLvZLKRjDn11AXLjoWJkdVqR2D/Ylx9qLU
Jok70B0K1ruGfeBw7RDfW/Yfw27QLolmO2W9uOai0cVH11nmlWfpGUzIw03kCCXZ0tR7ISmhzNpk
w3a/V0/0wsKk+Axm19QOOFyeAnU6gXf2cRHyWjJrGz1Wtdf8gMM1JsRgkxLjQBojpwLMnLQCC1CI
OYlGtv1yMiWP+AGyvihXzkq7yTQsHXItQG1fS2trWiVSrXSLO4aaiTnx0tg5y3TZRS6KNG8cnDpQ
pbve0aE6VeKFvrMYDiVMOnAWk7bMXGEtJdKT0Io4sUM67VnTR/KvBSFcoFcT24UnkvX35swVxxhK
48kFSIyDjfMHykZtvzGe4g74HqBkC3SxZf5iDamS/DNbJiS6QfCVGO8EwDAcOaVCe40957KpDyBH
jvrpjhjzHBNCUsbZo7Z5okcRevOmKo8T3ztVRLYgz08+qp0FThT0dsp2hlDo3rq6WXUku+BJjw8v
iC/vdOmp1EtRrzbjLqA76+M4uzpAR6TxDdc6ZRKUV8yjcpQJnv4+12DyZ4U0LvtRoSFN1lhVLIIK
GBWkIZuc0Wipzgskyz7hTE+wmO04ZtO8+PeDdfcMXjxEovOjfM7sPHpe6E23oJIQqVdgRn7nAUgm
Jf04BEcOKtNnh+qG1WoAfI18V99b4a6/iTA9fgDpSJIp7H3LM8sRQ2Cxvl/BnXBjDtRpITIqYPTw
Ik+e7ahE0UfucZe43uVNJBXlnT+j1gd0vM9N7McDxV81A2kuEcxQ1ge3BCJ44wUEXYS4rIvJI6gV
MoMabG+DEeMN+okuOv78W5Rvrp4DamyoJTdzoJd0VN747pN391O9FUD+yheo+QHiWY6HiXnxVjFe
hnFMadQzfqOFF0obtl0LM44GZxr1+1z7NqESMvXX0V9yPnVNwa6aRQxyvnESMR17YuKXbtNylKDV
TWcqghie3NooeDM/ZryBOTGWcb1DfpGHW8GG9LOZN7NqavSN5Tg14ye4ReNtvwdQWwtPWG8oOfHg
Cc24Vcnn9gZ00BshwPwGiztxFoQXAGoaOVzCFbtjW4EgwpUQ4TUEaX5cVGAyiTkDw+9fLuoM0n94
YJmdzZsCk+KCGI+HW85Bl+pajLNio0m2DO0gxn2uDuywAOy2AAXVzDyzAK3cnZpLUGMGznC4U5yU
/wDcLcsgzksRZGcC5hC8E3zc3uHi5RtfjwAWRJ8c2qVm5F3qtjA0FHLp6O+wUI8mgXgT9++PWj0x
FGFZ/TnESJDEh3+krES+t0RLqZ3mD8cd2TpRVsVxvHrTBUHYNxzeU2ebNttyAlSgVF24LSBJueXs
YRmkyZu8+x2ac9/xrPmU9xSXJKorxphj3y7p5Rb7U34haj8zauvNHqsGYbs4JBlr+son+iPIorLf
cgm95X7dFl2QxqVYiCBarLQ9RDUrZx5H/efHMZyFFvsSP5NabN7ps6cEXbZ62/X0pu1UGVvhKN0z
oVTvfKfSaCsDtJJHqR36/odoJcY5Drko9fRm8kHgmxBwUMDgQdRq8qPI9NyhZId/wh/OnsMa/X6h
YAwLgyoQ0hbD1fyQSGHr+vSZD/rNIiIQW7Epy+3WGYFGZQFJ/rE0zj5C+AqzLqt0v7r9xjgcoCPn
0SQIPLKME4v6KtRhCpWOSRzNegYAjRLB9il4Fp81jVHHS3VsXnSi2Md+Qg0xK7HBFRUxSevpw3p5
OL+pzF2hfWx3m44+sHsYHLXGe9d+1nqViCj6YPToiDY8V4yiYk8jdwvn2hdFegjVZxZbws1PwJWK
zuAt3FisbqwlW7aiaQhBluIw9h6se9tSDAPUGpm1fOoyMLrsRbMUS3JiTZ0of2q8Gv59rmLP2oeD
4CqMhODKMsS5gik52q5zUpKpiVsm2zRCL/AcsLYn5j1GucqA+/XIBXTvQmIXKhFDedjgY6+gMTeT
akRaXcvTTdCmxXNO5HX1wY/KNiZ8f9AOOEagcFMe/OARbzvs/KcBJ17Xxz/KDmmNiZi85/JcrwOX
zRJ5tKFM4wy9x+nLuKhJ8H0iYH0sflyd3avZor7ZC6XwZKFRV/VWid8k2dzZzcBuqF8RfbAlQNgJ
j9SG9Geo7bmruDhHmXGfGcCVDedY7k1HKZyHtm2SYTix93eM3hSbN9xAa8a/GzVsY9JTiLaBbeVJ
2BB+VYohLJLSMkwED2FzE/nvjpYtnc74/Mi0G7eHBtjn0+bwa0PGzT7YBPyd3HDc2qj+FxdVQQJp
Jhjz9zulc3XR5kztXo3n75CmA4i0DCbYiguqfOAakhk8Vc1ZYeyD3w5tndDuAPH6q5glfC83PB4t
DDnSuFAmy49yVDOdvvUc8iayQhnA+UkY73s1pK6FZHJBg+k3jkW/3Bt0Wa0EJ89K8WOycQY8tK5o
/RrbYxUZX3N1Xlrn2OHSjx2R5NYJlw1QofUlOUhhwVxUzc4kzA+7yYk/5885PoSP96aQkuDky/kt
hW8RGcleUOnI/qamWYsVs0ctU2OpTYCGf5Uv4L73EWDtQPYJQROmGBDQi6d91h2awo/nr5a8mjMK
PVsZ8BcCCjoLxeL9sULD2niKDG9szK+tpnrHYhcdKup+fplCts01L12tO9q9iKJeGZKB0hbxbdZf
hjGhajp8mAOlvWzbnfN5YxfDxVCCHOuCE+kk/3q9HxlZEwFiIZWGU74OUV5M5AEXoiSjQuRl/Qq7
IqCGgnFAR2SJnJW6sa3XnmjxkYEKAhWqFboRTLm4bMStW7mGBXw+821aJrdP8SBjKd+6FbUNcTlV
4xKA8OyFMktsjW4v+nl/7LSU1zicwkkwedq81ZjiO/OO7kT0hSuK7VEojnTA+8aawi1uIGeLikBA
g4HgQQNe+YYH4SSznb2PTRV70oi8qqrm+P7CAbA5FvFLWqck82SYCoCE9UFDqDWkuPNKZKrCFvQh
jJWYsNmkGjfdqY1nmm1gkM+5fbLyWcqMZ25V3uiTldtuNVcFncZwhnR0VdmhVyTzbluv8LzXXzB+
0NZoAH2GTbSVXdQDk2RnLNdAmLsaTl0THkDHiNAwfiY0Fj+PNCQY+p5kpsquzyy/8tz7ODjx5OF7
RbsPi0FhFOPo+7g76JDfZyDWQbmBKW5N9dENIJt4ug946/h90vsNqQU1gpLn2/WaMcOwYx1CSDam
TIla3yUuU5mbD8NcMtfniIqIyyEj7X3I+RjPPvMe2PnTvfA632pn/1eocbn2vNaY4L8d5gqCc9Dx
NNHF97Ns/NN1WejuKV29wn76up7gWGA7YD5kOF4mSMWydHn3bl9OcV60SLUYq5/3ck9B7WXbOyUb
HwTVvBpTNHeRfjnFE7laQjRDtFBtSAbeF4VWxWT1Aw2/8mKAejIuOMtOaO9BTWkxgFa13NTUardL
379VlTjpEYwC4odhZGlSonpT8lOBaztN0vb+0u0pkbjrHiytl4MLrvzc59OvmctoSiBhf54Fbo3A
yVGKcRFm+BccsihuvBTf/+xz53O8Ce8QTNNG4ur8XbdW7AEfuZ170bEv0LFcaWoOculj67KZCav+
Tjv6TWqBzX86tXl2ChJZzii8SUNvLmJvR9JO8AsNC3i+5PQzE2vBJNBo7rlH5wqL0EmXv/EG53Ag
IESXgvpCajIs9FN87JPEIUkH9Ay0u7VOQfuoLVoEfBd53uLc3JXqwz4wdq57KyliJ0mYsXNBrR8p
UdEcxVsiUmMyHwStjNr7ycaoPj0m4HNUzefkyc0JHy80bcJstF8Q/NpVTGI/ck/x
`protect end_protected
