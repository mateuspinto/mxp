XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���e2�M:G�~'�<�KЙ��w��w��h>OU;��1t��y]���j9���0#����g��]n���r�������öѰɑ��u�{�x��H{֦�Q���El8:�_G|��Q��Q��P�z��!�B�/&C¤d !.��*���3i�+�<�v�.�7No!�ak$ݲޤM 'P���Áxe�����HKOگ���=��Li�ΐq�	e��%M�N�mωu�?2d7t	��~
f�|�4@������\�T�Q�(\d,�#�7��8��MF�*�פ�gl�P\D�$��������A
�´�I滶)������W?��'�Y�O��Y_`���_��KB[�2,��|OR��Q�#l�.8GY�f("�':�f>N{��󁦱z�|��xːxGUvC-z�D���N��$���I�I�P8�禽�g�`w��A0=l<�>�Gp!|�	e14�P����T����Q9���y���oU��J�R3�K������
�4�w |蚊:�uG�s�5p��ߢ���P�V�@M��ΰ2����12s���>���H\L��Z��v���Mm��bƶQݎ�?LH���`��&�U�[�F���P�ڨ���,qnv�+�K�E����ؒ:�2]���]["�ѽJ��߆�a��Ȩ��liƶ���ب���/�mqQe�a��Z�4�n�A����l<P|k���M�Dzqy�}=�55�v��qq�-�7�I
B6c,���ٮ\��#fD�ߧXw���XlxVHYEB     400     1c0^1���{��ק���94�t��n!#���W�{��F7������yA@��ev�z㰟��Φ�w@xFO��n��k[�&�c� ���c`m	�������4���i<�zԫ1���aĬ)����ʍBF�-\)�Bٷ���bd�u��/���J�$ G��,:)���v�*����T?T�_��|����BHW
:��^���ȶ>,��� o��%�t.5��Ym�D��v��(���_�ذ��M���n������Ne���0U�R����e��C�,�kF���WL�{^�G�_��f|B��H"�I5�)>�m��+xN�5�⥮ߞ��d���-��>/�q����㎯D�Ao�EIX����|0C=Q�U��	���[��*V	�M�q�=�U,@M�W�&�!��א�HaPJ����p�ۡN�p"$e��d<½N�"w��a�XlxVHYEB     400     160���+Q"�C�dK cvO���uKI�B�phٸ���s>���Z��	��&�c�A��~���OC} Q�&�_[�I�-E�_�t�D�t'�K��Ц� �H:�po���)���� P���Y�����jr�E=����>�^Z{�I�{�	�t���:�K p	ύ)wDXQ��K��`���R&/X���ߘ�N]|@!��i��#����E1c@+�|*>��/.�TO��c=�q�Wo0&R-���#���m����QB=�:��^$��$�	��i�\���=��j��޺�ӥ&����/���)�3��4��:��7���b>�g����F�d�*Z�>Q���u$�ޱ�����8B�0�XlxVHYEB     400     160�G���Q�ܿ�5M�ms:s��N�4����Ora_w��p�x�F���h�w1U��w	f�-�	���q�wo���1�-`p��)ѮpB(�W��h<��X�Z�ڮ�3`bޠ��gWt�sٹ��s���,Y�C.
�vU��k��Ѡ�%z��CK�Mw7�II�@��}q����y��+�u�0����
�m�Lx����?�mB���Ns)� �s���GT&㝕<�(OQ�Đ�i��͘�{R�1|m����c-u����ے��G��r��[�BAG,��lx�R/K3!"�:d0���Ĵ��0a�X7,��}�L�3=��♶��_���?'�n kQJ͇�:�ע @L��XlxVHYEB     400     100�q�+��T�;
(�qk?OÔ�2"�8�*��è���{���XtS��P�Qt�+��1B\2��}wd����)8��5����诛���'�H.�/r�O�;��m������9�N�d�r���'��+i�9�O�Ial]�\�7�B$Wr��h�M�{B�_2��?���W��o��~b�,��E���_3����1xI��
S��Kc�󚔀;%{��1ţE��h���q�=�)A'�zXlxVHYEB     400     1a0Gϫ�ċz���B�Dc���q)��W8�=�D����_�����$�R�[���o$G k�����b>�%�~�� ���T�� }+��<�G�Ra��=D��;A���u��?�h����]�ݠ}]�!ΉJ�����ё��}��Q�n̿��^��'2_����w��j�N�m�	��W
I;�o���.���9��W/��yپ��,T'��L&r=������R�'�S�����v�S=��[���@��i4Q �����X8�ϩ�"�\��b/�V��.��M��Θ�S���)W۝�-"�T:P9[�����`Π��4��"��Z�)�*�f�b�2��J�kwE� ��_� *�W*hw�H�.H6p�1֥tBRs-Y�;���}8���-�� yM,M�������\h���XlxVHYEB     400     140|��G�������2�S�]1ޓ �{F�fV�#�DH6�B���V9�^�'G�I	j^z8x�T8m�k_�Tƪ��|�J_�@�\�����]�KӭZ�7`��Mh�v��4�Ȏ������9�(���yT+?'�!�=!����4�jN8���B�-Z�6��Tab��d��f�ә>��z7MP-�����G����FZ�����%����"�?(�������Ym�5�n��xEʐ����E$�F)|joI��@	��3���<��.���G��,X`����kP��'?(���"[|�#��Ay���@D��p	���F4^��XlxVHYEB     400     120�B�鿾H%�P�s�79ԁ�>?�+��	���h�l�)��Tyug�7ݴp�Ҏ�m)q[��9R�`���z/�	dP� ���+Г���,&'�����%ǫ���)�D>�,Fƚ6;U@�� �⣏�O�ۮ^kx���{aKS[Df�Dl�{}ϸ$�9lf��ȱ�w��%�=��� �OJ:-M���(؎e��,���-�0��Q]�u�QE��MV����y�櫍��M�y]c�M*��W�:��`ra
�;�;#��SF�Fn�3[�DZ�t��I��P�XlxVHYEB     400     130̷!�]���ֻ�8AQe����7��!��&�\ z�[u�����bח�>@=���V����A��B9V���*���~|�~#�t��+�u���ti�����>�]���|�jΦ�n>.�����p1=��\i6�����p,�Q��o~B|����rR�o�ڢğ�b䈞�)��dr���o�i6����i�j!�ů�h5u�jK��O��MɁ�f9��L���C�0O�U7ۇ���	�n\�V ~8�R�<mZ�s,(X�� ��MO��l���e�<ᔒ����H�w�+�#�a�"��6��XlxVHYEB     400     1c0Z�;�J�ki��l�8jaA����t�V-�Ͽ��Y�*	60�:�W�utaq_�7���,A�G^gR	؍��'E���f����8���[ԁ1�S�o�BԬDYз3O=�W�O��H�޷qrJ���j��b>��99C*s=o,��m5�Ϻ�Ak�/���y7alP��*��>����UƵ�v6�Bj.ȗ��V��I�!v�?�������se�!������Fm�Z!#�s>(׋��{
Ʊz,�e�Q�<s*~�?� `z��m���h�[�7�&S/۔��Y��-r��oc��,kV/I��Ѷ����T.S�&ķ ���V�(�Ig&U�j�1W��B�P7$��ϰ�KVRڂ�pw�곇��Gզ�	x���5��7@_r�ܨOSs�X��1Y:�Y��:�p��Oι=��;�����d��`,=P�ڴXlxVHYEB     400     1a0��������PĨ0���p�Ԫ׎+h|I�����s�J��3��y�'���bY�P�T#p��t>t�)/i������&IAk׮p��aꞘ9֭Qi%I���X�*֕�zC��_[lp$�)\ ~���8�++9������!/uP��`��c�������M眄��Y�w�����(Fz\S���5��͠��R�z*Z�N��r&�;SΫ���7)t����~�}.Dx·���%�=e��@���zz������q;0zO���M��D���\`������$��)����������a�ӿ�XT����<0�����p���������#F�j͍~����M��ļ/����Au���MN!lM}S.�CmWM�j��V��W�p�W�r�[���XlxVHYEB     400     1a0"�(��/l�	�l����+��Wv�0��{�guA!���ʾ�8	�aٜ]X3�fέ��ّ�1\3.����]�^��:���|Iߊ˴0b� ���J�N�($P�OQ�����E�v�,V���!v(#l��:�6�|�e���]hv��V�,��?���3��
F`�1�q�*��,ۯ{{݆ų��V��x��oH��8U��t��"`bfR���K��t���qi�9�8̰ �B�>��1+2=+=Z��*�����}�����-R�
}!Z��<��<v���~쓄��r�&	�L�+�G��W�5.V�
e�4Θ����W/!ewl3Z�t�Ϥe��֬^�Jao">-aq�
�;�$��K�d~�ڨ���Sǎ3�x �sa�-*w�Tǲ#f?JY<��:���"XlxVHYEB     2d9      e0 �ñ�u��u=:�1���uqr�͇Y��2�s{��0����t�cW��<��#�f�h���5�{9�а�&�3�C���b.��%B��,�U(d�S��A�kX"kd�?�)��d&�ծ��R�~�XQ�)��;��d��g�À�fR��~����4���G)���@Z��h���">٨�@�g�.B�0͍y	��	�"�|��}�l��K1O�mu���+\�