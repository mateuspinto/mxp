��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���a�`q}�-{7q�s���������H|�?`�G�{s	i�'e�6�r��u�
n�3��`w(��Ђ����fOnOƠ؛���n�<(��������#�G>�#�����_�ԗ��p|�nZ,o�jz�[�1e���w�σ��7��S�3G��id�պ��P�@V 8#E�wk
��]l\}��XA�^�&�%��092�ō�SOC.���UL"	+P@��3o�ȟ䥬`َue�]���CGC?�8��I�a2�%K|h�4/�s8�95s����v��=1�]��Aؿzhe�\��K��/��r��9Z����TE�(�<����g��??�����AsT�J$D�	���0�B۸m}࿄B@�љr8��K��m�XDܖ�_X�F�푖'��]�Ͽ��ùWTB���Ȟ����y�m�w��ٺ��Vt�7qJŇk/��>�3r;9ͮ���JH9`h9(͘�b�Uì�K�`d�z�5N��+������ɰ�?���f��
�mM�a�R��<S(���P����x��Co>�����x�j�k�t��5$/�D���6��c���#���#��Ȑ��U����I�y���{#%O���/���݉Rd��'R�U:�I�}�O�a�p9�|�g�T���K���>` S��l _S�>�[tJE��y;\ܶ)�ܭ��e����lO}�����*!M��xu����N �����@-�N�� ����$��J�`#Rh%��:���]�Qb3m�Fr�����o�=D�=�~�Z��,Y�����
J���N��U�cM5��A�Z��6��g�C9(Ja_de³��BI�~X�ߛ�sscԅ������?8�"��$��̥��y��x�.ߺ�ڪ�P�92_܊�Om)ԇa���E��	���:�e�B�D�#5�cc�~�W�%�� fɺ����4JX������3��MX�I2&@���d�Q�Qsz��ȱ�#[�/迋�KK�un�OE�a�����i�j�������\��'��[�8̠'�ߴY����N����F��~V�9� ���]�8GV���R׀&~�g���BXH:7��U����}�k�~�+��֎�,�7�(�J)�zNːھ�ެ���,c�$^U���+ODsٟ�����t��#Y��G(;���c������Ւ"\�vnŔX�8h�� �J	B�Z�/�(�]G�NY�'�vo���_�,OI�0��$�N��xt;������S�9@�2���2��{���Q�f�6���u	�������;��7���W�m
W���A���L���ߓ|� 2��+H��>�?�Jͯ�~�����gQ�] �M���q݁����!	��3�Z��0�����}��ɞ�)\��kg��i�S�$�dG���& ޭ��W3kiа����؄^@6DK�P��_d
d5g�+g���� ?��q���@U�Wg	WWC��J��	�:��{X"5B���w�j��V����	FU�:�!ja"�3���`2���y�W3�#���4ׇ���F�3h�G��l"������sPN�l����!R51A\����fo��ޚj��zƼ�67�z���7��d w����$��ޕԛ.�=.�L���L��v��y/�Ms�z��?I����_��\�k����!��q���e��yX��LVRjuC]R!e@y�4q/%�k�����B����-����K���&g緀Z7,P,�o����g�5~p���gj3�5k��NS�s� B���h�^�C4(l-���A<]�w�*�*D6Yّ�VA^Vɱ��<8V�;�Q~H~����ic���B����8%<�
#!�C�;L�z�>s�|��_�3���Wy%pB�j'����@+�D�U��RE^��P����Z��/���ҝe�obMH�z������$�����W]��M��Կ���ax!tۉN��,��{F��p��Vh�"��Nӧ�5��U_U�\��z8����u�Q��͂@=ũ���R��P� ��"M���5�r�9�ܙG������m�� �1Gs��%���Q���hd%hq��n_H���>aP���=T��T}>���u�Sa�� ���lTwVE�mיd�\~=�h���<W*��H=�����{9WZ��=(_Az��̓#E�w"���!9c����$@�����_�1�>��8Uo�!'/ը�������lY��5J+�8cl*��%�����=@�g]��֗P�в{,��7���3�%3e7N
بx:/�)j
�@̧���\a��-y^�z��&�9=�� �GG??��a�`,�v���ǲ�I�	��S�.�l�:�B�h�]�=#�v�_%6*6����+Ʀ����M�Ej��/n��b�rҴn��z���R1�`liH��:���;��C����.X�3�N7.�Z �0̼in�+��d��Rk���ض���`�`��Gλx��3-!JD&	��h�'o�J��t��d� @���]IJ�5�l�'z�ؑY�!�ⲁ��M���@��)t���f��� ��t��y�tR?F$�g}$?!���>�5��
�;��������$���X!R-���6�\��AQ�/��]�^����������ˣC���`Lj�58MH�D�'���pT?�6(qO!����UЌ�$`�s�>D #�ΰ�(ab��eRxY"�pҧ�=��Kz�e�5v���ܱ�����Yd�5�%$�͊�5��$�_�~�=9?Hy��w���Pm0_7�Q4h�(���&j�Ԗ����p^M���#|FW�&녈�QY���>S^��n��~�+abЈF_`�����o_��غt�N�5����Zdh�����A�X�#�F��)�h�,�GRM�Ycx@U�2�BZ\x�q�N
������
F>��Y?�M�茫̿��5!��+cs7�lJ��#d$��f����9���W�N�vՇ1��	! lA\��(����"}���G�G-h�F��e4�lhL��	." ��2��$i�G(����NlI�v6+�%���b���iE�|9�R��Z�j '�+�?H��[�1��J惾����1�AE;��ǿ�L��Ou�;k}���.��a�P��3��;0�����;�'��p����&��q��JD�1��C�H�]�p�x���b�N���Th���׉�8Qi���/?f�q�ѯ�&=�|I�i�[�+�A�ױ�ܢ��pd0�`ȶ���ز�{͇W�Q���ļJ��#����|�bSЃ1Gfa�0��J�A�)���� �e�ht �KW�R��J͑�����,;M�)I���E�NJ���g����z���j�˦-��;��K���l�6��ԫV�?\��]T~B.���%N�������db�r�G���Vpއ剘��;�#/:�?&"M�l,cҧ`0d�k}�n%(>��l�?���FԺ.�
8�꓃�`��f��:����H�,��QtSJ�9F�pz�߭�AC�!��~�+��A���x"�}i	K����"�v��6@f��p���N#����y�d����aEjOl���� m(�@�D<�9l0�U��]�ar�F9�$��Qv~k����S_�L�������t�4g����x�O���b�Jz��"�B5��6�v�vP|���bzr�4���e��{�0�k����6��/J��^����SP��I���#{�)����sŶ�ʆ^	Ue4�f#��W������Ԃ�h�jW��A�	��,;>�a�RK�s4
�^�V���P�q��Jf̌3�b:ߙ�l�\	�j>$/S�fɰQ�tZʯJ���VgSaH:"ZLA�t�p~G��6o�ާg��P��Y�s�_�~�j��|YFO�cϯ̫���&#	�?�QF|��<�nP�S{��m�Y�q̩��rl��+֫t����#	u�>�6tx�u⿦Mk~6y!��9}����{��7V4��P�	�hc<�XA��Dۓ ���I��*Z�� ��>��#ޘӴ�;�|[E�M��eT�1̧���Nkٞͪʴ�.:[,�W��Z����/��y���0,���h�?1�&HZ>�������*��è��H$��̆�!4���(s��0,�{o�絊{ŷ�����ێ����,�d���vL*�C}W���vD���i���Nu�w��V���|9���s��O�m�Pq��6��O1\�h�9��h�5:��"��&�|Ԋ߃�든q���
a��f��œ�����1?�v5�������C�	s�K�`nE%�K��dOt9J�r+r=��/"^2�]-P�f�Ϟ@<%OSl����>�������������I�|3+��*W��]+-�E��vw=@S�z�eNB]f�Kb��{�=�QCBxݤ�;�]���S��.�KmվTRR�@ߥm\|M�[e�G|�S2�"����HH?Ç�����L�U��R�l�/��<r'}��<��Ym���o3 �Q�����0M�Eژ�*ν���&e���6�fK8��׽�z����4�^R�OE��B@lS-��E��~~-ֳk���-,n[�U�W�J���TM#�u�ny��LU~�vW�:��P��T{|����;7�"E'T�f�8�g$��C��=j��aΩ;	���y ��[����ɜ��(cR�4�_]!�Gz�4z_�b[��q6����P�U�K��xZ7^jF9pdjb�?r�_��
/v�4���rS��q���m�Im4���?E�a���)�E򛼅@�s7G-p�ޏ��R�,M�Y��ܽN�n��%Qm٦�J���YW�}�ks��V~X(m��U�x������=V����9b���C�H�#q�����y�x�oOY]����]; %ݩ\��?�Dp3�g��qˠ����s�Ҷ
����S8��w��"N˪9��5��W@�<��J䧍7�,�aM���
�r'[ ��e� KH\���Wf�is=.����hw��4M�A�bT���,�O�N�z��1�Z�������I,����r���{��PŐ��}�r����)ҞuA_��׬t�Ϸf]A����rg^*N���׊�%i���e�6@�Q����HO�!|�i˜F^(�?Ē��h!��#�A��0&��J��r'~�\�Z���5U'�k��?kP��"Zz�h ����o�)�.�N��-���3$H3������m'H>o�6Mtz���uQ 1�#�ߏ�6pt�E��y/)��M�§�%D�.�|? �RUr���j�G~��m��W�f��K�AG�[�IoA|[���Y���=F�f��m��5MV�4 (De	D�C���l?Zv3"!�m#N?��6�v�A������D���W#��zq�������ɖ�������(����;�h�����(�(�V�J�ƍ�OK��� U>�E��2� {"�Vp��q��I�h��;�m@x6;��;Q��Z)MT�R��w��F��Ņ5]eb 0*Yg7�R��wPF@��-��͑p43?������j�ƞ��sxi�`�zho����M�F�.^A�,���*����MW�4�]�?i���lu#\!�񩑖��E�\%�.?٪��hR��1'x���(������F[A���[�ԛ�� �5iI8�_?�4��`1h&��K�19c��[�"�Ir,�u����U�b�Z��w�e>���1^���.�u4��<�W��������aTrye!����P"��
J�z>�<�R
埌fe���p�2c�$W�x��}�)���U"t�ٴ[A}S_�˄���/@bgD8Io$� Y_7⺚����G�+DMv�h0C�x���x;lCsW c�E[���2�H� �3��\�O�e�`��µ��_^4�*.�n$jt����F$�	�������\���zւ(t�Vq�h�Cݹ�Ȋ&�I�=�{�v��ȓy��ʋ�#����B�ہJn��{'c>�����+'�'����^訃
��=���zFU w��Q��k޿��Y�x˶ѷ�>�������Z��`$��N�;�x�f�u5tR`���sE/?>�[������	�n�Py��X�M��1i�7�t���j�	_�����^��W]�ARMI|!�@����a$|�����p�6_K���@+��{����h�8ha�"Ə*�7�d'˯�%e.�<�"�A����0�+��<Q���y2Q�*� g�:�I���`}��9���Eh��*k�~��R�Cډ�r#-��c��]�pͫ����xx1s38�Ȫ�n��.1�'���K��V��*^��u�;�3�a���D�J�D����`��D���'y�q���٬޹FIʀM��o�O��I	�Q$���"�T�s�?������ṫj�����g���
��.ؚO�nHni;<L��u]g�+0�p�녓�����i��g������%Z`�^-���M���t5�>',&�ߎ. ��H3�+�p�&��m�W>K��?2	ĉ�{	�k]Mٴ+u�=<�)��_&�Z��"�O k��q�]9�#���u/�߁VQ�a��D
;؞�����HN��+c�22��?����l�}����n2������N�$���~���ϓ�~N�Β��\h[��D����(�H�<qmxX
�Ƅﺦ*����%����C�k�B��:����&����m��	�#�Ѻ�Nz���R�� "��ό�K0;K-w���x���y�,�_�?�v���������2��ۗ�
�H_��Kw���}.�����Lq�UpD]��i�͡���>3	۾��z��)���+���s�����.OΦ*�/ʤ����`%��-.��ؔU�4��tB���l�F�i��l-V(���G*�i���L ����x�O�'�J􍘲lƫ̧�*Y�y�9�R~0dqnM�]v�qu��ƽ I��t�Ƽσ�CB�Sg�}���JfE�g?ݒ^I>�&�������|���r�-3��ߤ|���Q�J�D�.�5s�7�|�\�cg�=.��X��b�rŜr\��A(g[;��#օ�C�G��ц�w�$�T���c�#e.L��#3@�ȗ,�����}��]�~�72_!:�����Կ�_��eN�l��R�,�
j97I��Ԋ�ϸ��`�B,�ԸmHw���(`0D�{'���v�m׼j�k�����=�ᑃ�p������ ��5
rÂwH3O�Nـ�e6�9���ֻ�l�$�S�����M�,��,�>j�	V̳Bw����Բ���-����%��S��d��^�����t����3=P�[;�cZ����������%����́�ŉ5dJ(��.x:�Z��j�����]��y���ݬHaD>��Lh0�F�c�l�t2����FC��J�L� 6�d�K�O�]�#nuK m��m�@UP�j�(K�f&����6"�P[S�PL�������!��P�.�	+�?�)�B������Z�����)����+��aF9��[E�6���l����@��$ښb" �q����1T��M��8�=rI:�������K�8����7��?e�n�>�y:C �-~�+��m}}�ҩD�����Xŗ�R/ɧG���X�&<�$�x�Gn.^�BJ���)G�%���Ջt���]B�X�1,�����<ubrQL,K�_��	�?�Z$2@$���
�[]>���8I~��VB��M�B�V�њ4q��'mf���a���'&�E�8Ɏ�/���B��p�Ɛ�j��o+O�N��H���j����Q� ��4w{Ҽ*g���rG�A�q�Z^Jg�8�s2	���Y\I��L%��$ͬ�ocwP��%���pQ�'c����B��o~���ЫK��
=���$"�Qɝ�V7+B�K��m��!W&���3T4�Ofx�5hd�'�\W+���6"�~+߽z�0�,#i�Iq'Q�����5�c�g�R����u�@��
��]����^g]�P��%���˦u7I12C��8��}� �`��2�v��ZWW��KTz�d�%맺=�QU�� ��s���I��ܦ�'��T$,���GR��y�Ϟכ�փF��f�����ݔ��Tf��O#Bߊ��,�(��C-v�GZ��p\�X/��/X97!��<͒���Q=�Z�(7����z2�kE%]5�b�W�Zw�l�A�D��86g%c��k���O;���sݏգ,q�c���(�6(��V�^��H����I�қ��ŕ?
s)H�n;Hf[��c�[�mD����+?��^H�>�Z�X�T�ަ3Yާ��I�v
��>=-��Q�#:���Dig�-�0�jݒY>�c�e���k�Q���>�L�ԥ��������J��X��,
)$��Sv��lԟ���,�k��+V����׻�͸}O�*b�O{���D��Z����b��-�N�/W��)Lh��qϥ́�� �sĺ�45�����8��Us&���4�� �����+]�t1U-��+�@6���{Me?���5$�KJC��ަw9��6�2h��hJօ*x��q�=a+�Y2>�v��6��=��=ap[q�L��Z�֖�Y}Hk������BU��B����4\hden�~S�y�{nb�t��2/�`鹛�ʹL��l��{{O�''�"ȹ�b� �9�P)�8d�.4��̝�k\�&�n��$:�+����n�~n�T�"=N�N�>sm��r��C��db��v�E~E:��
M��W\9UQz\�?���yx��ɣG�D�(�B��P��,VqO�~�;+���L���&�4~|B��r�҈dA���W�Fq�MTh�Ho��bm�0����E��a�t#5鰺2���q7}���4�	��[CA� ��0n�d0�@��}��-Jpm�Ech��ԑ�/�m*G��Q��r� �_�me{�w���0룠�}F����+bX*����d9Uyz�uXX�k�^� �Iw��J��c&��oMuG�<J}��.+	�K@�D�(R���9���o򧕁+��u�cF�F���:�*���b&4����L! ���"�3�$��<L?��_���p`�r$�����1Z���YϹ���*a�ʘ�����sX3z�$q�6�c���~ep���E"U�Mء������Vl-*=Q�}[���U�۷��jFp�g�Kx"�']����pE�H@Z6[���`F��d�D�r)T�Y��r,����_B7ؼ}�K���r����'$xd�z�B�"N�x����!b��yt��U��L�����:X��������o�ٛ�6����
�X�߫͐T+t��F��gP��ݦ�P�k�*u3�{�9ĖgvL߻V����a��3g��\x��
1z ��#&~�/����y�6��{X�if���>�Ƒ|Rt�t�$��xEy_�/�5��BZ��ީt��>K�WZ�i����S@1ݼ��W̒o>r؟�-2�\���� Ërze�?ͭl Ns��AT���|�rql[�o���B [���D��)��AB�P	E�
�t)��W��ԭo�?��foY���M�46g��V@R��=�#�2Z
J����ç
�PT7E���чr�,t���W�@�f���Xr���8��L���N�広��-��1�T@��,���B��^��欨&AɪT�v�U�bn�£	u��`	��"�m��we�up����Eh���J[5���O<^�&Q��(�z�����k�.���LUuҟ���>ͺ3ѽ:;d�F��91Ҡ!���4�[�-sX,"U�!��A�����#D�*��
�E���<<8���l��R����q�6�8�HC7܊V��T޷6�vF.���|��8Z�λ��H����$�����=�i���z3�f߀��h��?��(I)�_��ՎG	��u�=?��-s���Rx�6u��^�}��1 �ߒ������ ������R�:������ /C,�SR�z^���96��9��0t/lO�N��*jس��N�x���@}���?\��k�CtHAE��ϖ�腋�
x�����H���:�(�P8J=�x��m��:��%<���{Q/i�4��,-���؃��µ�����5(�&���ef�'�4(�X���-�H`�x�R28:KV
�hxf6��RM���69S"Q���^�����,Z�Y���l�]�Q�}���|Q��������3��1�_)_���g�J�������9	���Uߏ/S���KL��6=���Q~�7f1-�63�7�p��`;�aatAF4�f����Ȉ�3{]yY��8����jҧ�[�\��l
�����p�_�;�֎��n����Muొ1^���,���&~CK� "˔s5LBM�(y;6� �@��9zB�[=!��DBa̋�-I ?��O���CG�=-�]))C�n�Q�d��#xp}XMw��wH�SBC�"�3�58�c���2=��Lu��/�W)~C�)�0�Xd�����#O��]���5�;���2��Wbq����:K�Nђ���0��Ӯ��VԤ�_?�c����I�n#z��:
`��Ri��UT��6����w��s	1�����R1�b�!L�{�J��M�&��'�UM*��U���D�����%�̀��*��|(J)x���B�&�%������[�J�<!�D�Q�r5���E�>�Bq�A
��%#)�x��0��c��"�f�T?��/D
�
��юŹ����y)�,��<��q$3�9�HX,�K�S�l�i��}{��Ѝ[cծ�^�t;}<9&�5(U/XKK�+�XA����5u��XB�c�2ʖC4�|ƛom���S�<�Cx���܄|I����vd'2�;e�]1!A*��E%q�r�/�؅=��RҚ|��%� ¼�6ħG�1�	<��n��t�B9@�8���L��63�>D�uЊ�2����y����(�)�u;����Q�1,��+[j�X@a�v>rɕZ#�Z���PA!ql�yf!`�Lp(��(Y��~�Ny������u㘱�������u�4��ž�!��P��\s͆�l/�SB�f��wLm�q�h8	��i~s�Ș.݊�j.��	�j�8aS�rKv9�`�q|W[����\��Cu��"�Aw�y���(tVƁ�PO���c���M��ӆW�*�?��9�u_N6�b���b/�0��6F
�G+����.�Fw+ɗ<����VGu����A^�e����+RR�=��P#�-��Z��F�YUD'ܿ�o�aA���U��k�
�qm) v>�ϭ꽷�M�B�~d���$U�Xw�J��5LҮ�g|U��lO���&b�o-���w����� �&�o}�^2�8}�Ǝ J[���بX�S�<�ّT�����a��~h��V� ܼ���Dp7{q�\Y�E'��אּ.a�Z�R3s �kg^m0�q�G
j�Sҽ��Ml�}~���,Ύ��~����MХ�=v͙��ʋ�A{�L:(�M�M��\��'7LܞC��L��6�s_��/�4�Yz{��Y��+H���"]1��]����qڱL�c��8<�Q)�Z;ikᱟN�,v36һ�X5�Y`�`;������-pi,�&n�S9"C�5>�#��Ļ[w�E��j���k��gͳ�s\������@�y9i��⋿�R-��D�s��&_��%���NS�1��K �D�-9���A�.���,cհߏ�aVڭ�M1��v��;袷T�e���8S��K�[%�=��q�ח\u�9��n�ߟ��q�0-��g��.q9vT������Z�ַp�~�or��<Is�C���N�hS�Y_޾Y�A�U�̍��~�t"�L9��P�⋣�db���zˌI� �❋�[�k�j�e"~zq5��;q�l�M�c�PGU;��g���M1O�j�����H�T�{��o�ŭ�,�v�m{	��ڣ�/���R�ʍ�@8P�*O�Ԧ:�K�������*~��s<�"W�U��7�����㜰u���~j���ʪ�Z#`�w���	)�R���$>˾*r	��m,�t
8�;O��m	>D}n������7.�:�禌ԍ�y���YMj��wn���u��i���M'&q���j>��b~G�C����]_}7�۰�~�tm��p����&	��vb+wH
|�t6�'��t-; F����^��9����w�0{a���8�(s�)+�2��bGQ|�$Ɓ]�(d��$��Z���s�E;r�U��+��.hA2����(�u�1t�L�)���[�����K�wl}7j���h��J|E�RB�����}s��
����ʇ�i�Y�_�Q;�XL�eq����pL>�+~I9��^h�ɳ��Z��!��yc�Ř7@'I�	�3���1�u��%�JV��G�`�/H�7g�yj�$�V $#�bI泥8�ߋ>�+A���U��Bߏ�gE�w���;2zjx(䋙�#XM	��oX����( ?��n��`�nY�op�Θ���Q��Iǎ�T�6�����ɳRa���`
��JR�A&1d��d�Y�# �پ�~oH�[o��j���6��=�8/�n�o�=W����w7.g���o�[!�N8/������_���q,���d*��ę��.Ј&�]Li;q�#���˄�z�ٿK�Nvn�Fҽh�w����t�Z-���*��X�o��Y�t�k?T���t'k��Z�dn=���+SXK0�а�!X���{M���$�4WQ��X�_m�}�)� �B3��JN$����*Ʋz@�W�a���+̷���CV#5���@���ܕ.=��
xOt2���6�!nҥ�M�M����и�TPB-F��M�^|tӐ7B\:B.j%z�s �ɲ�3S��QE��h�+)��GA��$����������2r�nn�,]��d�pQ�µ�#JjJ��'��#�͂��$E��E,%�����+��nQe�`J�	p�z�[�\�q1g�rM5��S���e6ͻMUQ��oV 2���-%���2�F����C����6%|���9{�6&���~-�#0 ����E�m��"&s#��4}o��@�\� �D��+�RKpQl�+bF�H͟2^C@�9��]u�%�������as'G��C٩Q����C��﫠�-�R\������H�?"�T��}֬mR��C�6;p�]���1m�n@::CK�X��zćSmi�΄c{���9�b2Y��ӡ�*�2-��w�Hĥ����0��	ʫ�S�)�V��ү ��pr>������ɼ0JGb>�f�Kȱ`��x��)[y�\w���ע^��	/V���$l��r_�t��¼���W�Zw��B�4<�Z�/�m�ZߛLz{�*�!Oz�Z���<�e�|�� ʹT�5|`� n�HN�ۚٶ�?TJ��IR�|��:�ofWz#XS�Z'�n����B��QR��k5|����H��RRD�m��_BD8%��m1�`�k2�?�qCC�W]��h7�(��,��L���j2�A"��50Ȇ���_=�I�VB�A%k�6xv�w7��N@@#���0�'��/ekf�N������y�!>0���� @��ǒ*��}�KJ	��Ff�e��BH5�(��O�}A0�� �؜�Mn���զ�����H��UV|��W Հ�Xd�cV�z��-�	Ϗ�z_jس	�ByD����=��BE��������^U�~wU3[�G�[>ѿ� ߐ����K�Y���x���'��-h�v⮑�'J��~�%�i���[���tӢ�S����(x:Ζ�3g�]�'��ڵ�I��E�,J_��0�^.�y��f�Ǿ}�&DPhh��v��6��%!ټX��h>{)��lqh��T�^��M0Y�w�`��χ��������(3H	��)A������bGE8L~JDS�(�2��������z��\�g�j��.wEF���`T�����3�gr�qK�`~�V�{��V��эz��1	[d<�Og��M0	�P���h�פ�iH����+�/��wndEQ8#�ԉ�#�%�f(�4���Q�b���;�e��aɑC\,�
p$��98y��)S�`O��|�8�‗�1���E��3���9տHWV�9W�I��4�lMs����:+SƃOoZ�F��-�E�ZE8ꇮJP�Kn�Q�8���#2G�
U:�e�99��A�Ev�=� �Tf�WA^dR��u�4�Ļ�8��{�>�¸��s���n>?$0Z?��g�_��ȮB}��k�����Ɑ/����7a8ap�i�R$��ZE��tY��ڵ�%�F�,Մ��r��,��`�M,[&NN�myq�b�dT�t����,�t�2��������Ղ9#�Ne-��K���-is�1��?�ip�8�A����s|agY�C�s������ߖ�[U}�Śٵ/�S�� ��Fz��A�M/k:���y����g����5�-�!�.���mP,q=�_rn���Yw}u�ղƯ���6�>M���>XM��Q�9+�	i�I8���̒h���[$�VL23�1n�T��Y7ǟ��Tc��
D�s�k�GN�a�!�E4�#:�x���������_�5�i.�ya|h�m-Xf�Sf~��n�Nn�
���{~�\����q�}��*/��3�gi{�8x�Md�'�0[$p)	��\�VT=TS����uP��G�C�"�;�C'&X�/̙\�#���ʖ7����ז��&b��=���ĳ��l�m�b�w� 2">?�Nk���ƽ91��(��� ,�1���L����e�]�b+T:���C�#��#���Lqk����۶����	4�| Y�2�7c3Z#�z]ڲ��/%�f9����wy��O��rx�������`�>���4[�HD��J�&�׌��J(74*Ė �A\h��P�,8n����h-��M�XnS\�'��u��� ~��k";ŹU�)u�0��'�%b��>��E楫�3�>�2��/�n��_�wے����y�����_��n^�9��U�1Sc�1:��Ljl{���96x�^�[���^QX���wx�}VH�Ӛ�y��W��|��{kg&-Z#�u��kg<ɐ�&�QSѐE�&�e�-ϫ�ͺ/W?ᮚd��[��L��&P{����
�M��>c'�;���$�$�;�PO�=G���ǒ��%b��	`���
,��V����u�yW�O����웇.�eI�iͷ�Z}��ʑu���ǝ������,����[�J	�1BD ��>�-;v�U�^r	o�!���!��&�Aq������)W�f��*�fkL���z;�?A`_7���Xf{1�QN�S�	ҏw*w�?���翯���PdqA3�T��7۲�[�Qb�o����sK(U�� ��L^d):k�)����],���MJ���V6G����e\\��\e(󢤔]N�:� L
	6����.��H�t�0�b#y\2)>���,܆�$߉�Y"S�m��DJ��CG�:�<}CT��٘�A�U�Ϧ��Y��B�n�r����y"XK�9l3������9���$d9��пTL]�-��?B'�
�ѓ|��M���m&�~4Cb3y�8�m�f(q���J�����PcS?�`�v%�U�3�U*�a�[	�@Q-1�]�.�s�Au�ܼ���^��-pd�����EH��!��e}7vG�r<�}��8Ϝ���7j�<�M��[=���p�;z�y �jQ����h�u�_�34MF6�i�H��Í���B��dr���[ߠp���st��[u���f�$�'p��L���!�U�{������MG���3Sa䒓��<�d���te%7���i���=�}>�b2.JY<����M����	i�خ� ���=y�8����ɮ�с�sy#�B��թ���&ca�`�hxe�G��Qq�9�Q���3�[4����9���I�Ω���{����F<��~9�s�̈́n���7ib�Sn�#F0!Sa���,ӣ�~]����ixه�,Ug7�_U��5AzR�d4:C�9��}r���h���}��ͱ�B�K�P�:Gsi�AF�h�'a��Z�	7 K}d�R]hB�T���ȤThEɩ/�ŭYs�#���icz�ɱ@�����Q��2NiA��*���a#�c���Nk����:�����Ë��/L�9��f<O�DJ3�f��D��ͻ	:NZ��VSw��5�0�o���R�HѺ�;X=ܽ(�Ͼu�	��%^]����3�kP�D�@�=)�szu�C�����-�il��e���R���
����ͺ�nP��5�6.���EB{xT���+��C�.����>��%y�v��g�F=���ʿ݃�'��e�����W���F$����f����w��6��AKh�G�S�0�!���/z�x>� ���&������vt�!���=O��t��Ҫ�-��*o4a���w~�I X����ú&�!�ky�x#5Оzw@��9�7g�Ľ�˅-�2������I|$|��[��Abو�+����K�ko�20�����.v�KV9XPv{�uS�����4T�Bu�U�R�a��k��$������FP"�ʣ���ڸ7����+=u����,c[�� 줳��R�m��q�8yD�Q��hcDI��	�2���CW�kKP� �O�R�/͝���X��I��tB��={�ъ<��\*�g�9Wy]�cb|\q����s�V��<�#č��L��<��6�\�����=��.�j-�ת5)�h'[������� E(Z_5���X�t�r��6}�:,��ﲙ.qHS���1��*u�gt[+��,CQ���o�L��8�,��l2��J0P�<%*2	�t������������lTk��Nd�.^ݟ�o�
2�:���8�M|�N1FW���?I]K m씂x~D��CB�!0��� ��KL�M���+\$�W/J�^p��R�{�rb�
H*
_�&m�u�?�+=��RW��" 
5��v>��N��E�J�CRJ�CX�i^(f�)^��)ˁ�7�L!�psp5N���x��=����f��V[�L�\�{n����3@餃����S#�xք2v��;��f.�c��@�J7���2)�5N�\��"-Gd�}�
AS@ڋ�Ac���jT�{�c�΅���&9����@^�n_�u�R׻��jot�WQF	��%�������\^����(;$�@
j��5_�-$*��!�G5����W+"��ի��ĥ*��q�X�j_���H��L�מB�Y=�j�Z=�y�]T����
�*�=YT�����Y�	��Q�.!�Gn�)��t����s'����A��܌D��MD�u!� td�����S	I�Sc�{����woX�!�I¾��1r��.���x,��?�Hb��t1���)����i��#k�n{��ͨ�8���(W_��1� j'��.�A����� )'�\���k5wi	2q����6���U����։� ��r�L5�(��җ�7� +~s]��6'��Rcb�+-(��a�j�Ά{�����t�ŝ�G�ob��E���M�����
��;	���I{Th�5�
weh���61jCc�ĸFH�ߪ�R��Z�~�8v#k�c7[��ߠ��X9�nyW�rv��R����Y��>��l��eŨ�fZV�lo/VB����*12�g��};.qSqI��h���S�a���@������iP�R���er�>ٞ�4#I�jK�E�A�*�ﰘ�����<�z����Y���!���\^��d��榳F�V������K�6 I�%�X��0���"ҟB�h�ߚ$6�G��RX�v�ס�َ�z��F#������q�V�L~{���>�|��쇹\o�[<�]�K��>�?8�y�I<��(`A]���^��o�vQ@��� H�������3X���AkZ�5ɚ�����8�滋ܖ��`Q�����>*s���Xڹg:���F��y�@Gd�;��K%gAL�v���a�@qd�YC�b���;tv<9�	��ׁ�kf�y]��/H	�p�����[�~3,�L:�¤b�@�����fTµ� ��D�8��p�\�]����d(06Z5"F�3����_f���`�HH� 9�c�<bP�����L@EY��w�ܿ�{W-O6[��l_�b��x�"%�41�����$�!���'�A���'��Rk�?�c�߱H��+����٭\k�7/�
�0Y�E�������|�a���]K���W��oX ����gD*X�H�_@6�#�cmh���H�������_�5���f��]� ��x?]�{�_.*]{jK��.��������O�[D��Q�!r�Zy�;l����/[;�ޗuƵ�1��P��.p(5��Y(J�B͑�R��$;��ciHq�^[�H/v��]o�$��o��#T���y��
k�u)�i*3N���;�IQE(|���6%��x�Ȅ�K���f����hgM��AE,�𚭝;S�%z9sZ�l�ޚܼ`��q�QX��k]m[��eK�ܖN�bX�d��e�#4�ez�J��f�L�<v����!k>&�cK.O�㞾VN��)~ԃ����p��1(`RG<RH�H��۪^g[D$8�Oy8$�,Բ���ǲ��8�8�@�^N��͐:�.r��I��������J��FcX��Lpo�`����Co�X��GQuV&2��d�;B��m3��!���b�-�fm	;���	�������;�{�����D�43x]?7;_w���CS�2r5J�M�Vg,���\K7����Ǔx�-瓌��ߵ@�Vt*\0�x��SJ��͍;�E�Y���W��P�>K�l��Q���1&��5��`��J����k�V-A_C���"t�h��߿H��t �4��?�t�Vx �2�|��fŬ�/�D�N8���dMy$4�! K�s��F����>b­]e;�J�/gy5N�D��9= -6i����)���Ȟ�?2T�A+ ]��x�m~a�2��9�P�$���69�}Z��t���갈�0�M<���� ��%�	���ծ��Ъ�6���G��M�i�	�ކ�dn�t��{�&����=Ќ�+���5�t�s2�B=���4�r���P&��������qB�ؖ��%�G�� ���/��#��Z��xļ���B�R�'1z�m��H?K�
��{b����c���Ip�����-���禠Kz�]���A���\?D�h�b)�����d/ ����' V�߲�:�y@,eQ=�Md��`taw��6�'2pv���l��qۖ�m�S���I�W[Y�ǤR����l���6���M�~�� �W�	�I�5��
@�����7�O�h���V���d%η�ԏh�a�����vR�ݶE�e��}�W�6�����LО�i ����3���?�s�=�懚ߖK�}J⬡G��v�o&�p���1��ֿ�H�nf�nF�rA�B6���u��]�h�B�[@T��Ձ���$�H�� ����A��l�~?;�,V�􄫧�p:�V�����+���A�����f�#EО�Nno����(�H|y�ջ�
2HX�i��� ��,b�a�u7�1$g���9��)�>�������2��.��;%nxN�)hZ\Gh�j{��6G?�S�Qb:�U�ԇ�����;��s`���w�j�V0y��ᎽI_񘶌%�<=H&ZZ��}ɘq�޺E���\��4M�:�\E�D��(� �j�	7&+}q�����)�<�Ql�2v.��d�usp>9\]�'+c��u7EC�]}�2�F!u�x�<%��"XD�:h�,��M {���[Z�L]fl�α��J�0w>}�FH�q��~��0�'z��6���q����=��DY���1�N�4D�*&�0֬\�����/���;t��O��'K�;�3�`D��H"� ű+t����
���eFHu����6�O�P��HQWԕB;=�e�~������e`�B�]�O"�jēs�_�4��tn����
od����G��������p�6�K�1�����+� �؀ˀG��.�p�W%��?�n�Wu�O%��Ȳ>�f��1�8�ڪ�VW*�aM5\"��ӛ�(Q&!�?׭&�K˥ݧ��槄��8EY/@��G,�gi�!������K�k8���Hc�ͧ�j|=�a�s�u���O>���.�N�/��t�n�Z��K��/U���lM�'ۓx���N$Мr��lx|GNS5�$|w7���3H�tF�J)����=�z	� ~Q�e�ٟ*M�|GE/��k��G����:� J�-;����v�/3G%.���b-�Nu{�U��0Kp��	�'�S�sC�����7s�I�;���/zw������j��A��H�=S/�@�� ��o�E�֐�c��D��4�v�/�=&�?�=,�HxՇ���uG�NxJ����_u�@��:��ۼ4��#*w��&8�fy�q�Un�$s������'�O��`;u��u�~�8P|ky���.��W4=H"�{|���\��2{1����h��d�<�}�A�����8u��*�U� R:;#(��1�NV���I���]�X��J�������	u��&㭪G����9���8��H��p�|l�T&��67{J.H�+�CB������q'���]�uk��I�h�]
���HufOo�v]@����w�P�$z���W�	�*��H�lB�Io�Sݓ�6�s�.�:*�F���~���[S�f���h'�x���oRtO�׽3�����*��+����B9�!8T�ƾ޻��랔��ms�/f8�����@�8��}���K<$��3טV�^�9)���0rQ�8V�A|�Y�hW2�����WǧY= �(�!笜�F&G�l0)Y��m���a��/ԯ��%2"6����b댋E ��{I�O-����D�����w;�VMX՛�,?�T�͏�l;�nb	�y�~Z�Ns���ݟ�)���q1��(%�F?��7k�O����1�K���L��	D���ЈՈm������Ci��y��ӽ�dr(�+̘MЕ_��j�h�yUex�U�O�̰<��Y���A�����~`�W$�y���b�u�J1'ﻀ4���Up9����qRN�I����8��v�M�"���_�/�v�щ8�"1�<9�#*:��ë�. �Hg�ޥ9e��"��ܴU��@1�Ay[���
;�l��E�g[�@�"���8pl<�GP�5��]!�u��̙s�[Gm�ӫI�@\#���}���u �8yD�F/�w��� ��z���U��7c��#��� Q�����S�F [�j��"[�����A��A�FÏw$푾 b+�Ue�c�iս��֝��z�{k�������#j��/�	R+����N�)�*� b��������T���̀���/�aN�c��B��r��?�UW��<7�X���s&�����K�a��y))�KO���O���LC�������a�[�t�;@GV-я�orW(p��i^��?d2u\�H�ЁY�f�}
��r�8d7O?���50 �m�8F����X7E>������B�~5qKQ�-���s��I��J:	XV[��8���G_��W'濮�\q����l�}�! t�V�ؼS�� D�?��a��O�矡���g�{F�+L<�5k���	Cϸ��`�ת:��#y�Ŝ�c��ڑ���6���O�0�T��9��x�K*oL'M;��e�C}F,վ�m�*y��l�\̧lwDG?!bf���D�?{�}	j�)�IT��pY"4kV��7r=q3�@��sL�फ़A
!k��W^�R$�8�3���5f����2Y��� ���=%P�kBS8[��Nk�m�KS�IR�r��j?�
���*Mȅ+%��� o�x���3�wx�~g��	)���ln~����}��o�_OZ+Q	�$A3�qnXU��ȫ��啃�̘�ւ��`�[��>�s)<ܞIh�L🤸pԂ{&1�k |v㟉�y�r�
����t�~P�
�B[�N,8�(V�����o��Ya٩I�_����5'��*v�Y��@YO�E�Y��.Q��",�s�h��fiO�?���X��l�A�'���h!h8���i��h���e7O������5���cI�g��-� �e?�d1����`�e($LB:?TX�j�躴�7�5ѥW^(G�5_�z3�e����SYh�w~��;_� �/�^�G�[o�a�:v!_*��8=�[I,#�Σ4�z1�6Z�J�����paՍl�bQcD�`#�@ �9��e�EK���-Ԁ�� ;�����l��
FgC-��v>_�oϼա���V1����1o$0����G�����ޟ���=L��[��Ae���v�XE���(Y2��!�3}��Yl�S-E��EN��_�χ �L�@*L�S�z�Ha٭�P�@�F=!-I����˺ڛA:'��D����R�3����4����|+�uk���Q��֏�.41%�6I�mKЀLe�ӄ�����$j�Q�����5ij��T�t
2�$ɏ���[��:���:��m&pbRx�>�IG���&�o�N~����q������#sk���M~�K]����=_�Ν��������fMjM�~^\�#���7h-�������.�O�ӽ\Ĩ�euwf���!(*��A��v�80%�A��h����h���j�$~T��q�]k����V3����8�Rg7$�R�Il�s��;�U�|��dBb��8(��~
�����扶��i��4�̬����W��?���J �_ٸ�k��Qw����*W��0|���p�x���1��X���Ժ�KS�!_{٢�p֓���o64�c� �����b�xm������������k�YYH�#�9L�����A�௜�#@�P��gz�l��>�秭	��\�v�
��4�D2A�Ë�Ak�<�C�wւ@����4���֗ ͇�]�Q�a�)�s��K�]p�гм@︕�(yy�z[y�_�dR�I^@��Xr�]	�? 
�M�b����V��+t[v�^��.��<&�?=�v�JW�pGǋ�k�צM�+����k>%���N Kw�a�r� �������0�T!ـYP��[�e~��;z�kF#DvL�-9�h���(�4��HP������<���m5m��O.�o7�Q�	�Ui�deu��r�n���&[ѻ.4����3tr*49�iN�ի�+ofJ��~o��(��獤�r�a�mFŦ��D7��*Ĉm���E���D�3��t��?�3m3I���~�#�a�쏷�{�M�r������vw���b.P�����{Z�1��m�d�n%)m�~<���j�^M3S�̂���#���5��X�K�+f{d`O��[!���b��,Y򮤈���Z��Kz��6�X��2c�����V�@�&�B��jH�ۯ�_ى�SլQ��Ϟ�ी�	��a�T>�Ng0O٘?*l�i)��h*,��$��ɉ��Z��W���KWP�>��� �L�A�bN�����wzlL	㨗d��4��wt��Ta���H��Hp�8I>R�Bs��#w���r�SR�f�ӆ�&�6y�Ĵ����^�m,QxG �0{����%��O�"`?m��m)�G-�>de��=Q�@����s��J`6~�˭M֬z䁟�����Ç�\mn��Lf�?Lr�<AT�G�`�b��JQ!��w���<{�i\�Ļ�8\~���%�|��zh�7`�:Q��ϕ�Yy�[dXc�C �؄�!�R��{���bR�L����w�NP8;���˚H��Mc�o�u�D����I �B^>I��j2���fЮ~�'V%�ʅ
���7�z��*�=�_4�Z)�zb���9@ ��q���ꊳ�z��0P��Ĥ(Q��d�nGl���	8�X�Bോ���"�t'�Wڑ�ه�L�ta/*�-�ٖ�ї��o�g���I�'J���|��>�A*��� ZV�/�Sͬ�T���!�I��K�̚��)�ޝB#y���IWY�����(;3��D�a������H�m�n�>���Q��y����}��v�hL�^��t���!��i�����%�%��%EA��&DJ�� �
Uq�06^�27�~�����흶�x!V�&���� ��z��
��)ȝ�HS�=�`�Q���lQ��P-��4���_�lsÈ�I��Z��������e-ص�T����~�#=�=S���&�@�Ó;r�(]�s��L�SǗ�YmS�apc�=X�Ɣ�ߌ�ȅ{Uʓ<��R�YKoe�]q���^���6v�$�eCHW�J��v
y�i��$�ZK�o�������WHN��S�}���/��l}����5�~�1�2Ј�z��S�-$4�F��!\�?+�Et�/�y���ll: ���|7o�(�c��{��:�@=�4u���]��>�"=��ʢҤ�I��vqf� �B��H����3�N ������4'��g��"BJ���X��|����}(TJʮ8@�6��]RĲ���)u*h����.{����R�UN���]���>��iQ.4�w"/U��F��ELq����߾<�������9��f���JK�V�O�BL慘�KOffR8��:��W܋�4�ۺx����W�9�}�v�����K	�A;6��1Ӯ/��]�1X��ևl)<�<����\���]���S �� K@` �?��r������(,58�ĦM�w�D�<E2��"qv]�AIj��.4u�U\)
Q79�������i�I�,u�k�]��9�]x	-Z�\7Bu�(r����I*ȓM���z�lv���9��?`�>�'IQ�N�XZ��Z?��=?:�MY�e��#�sK���f�$��>[I��W��L�3VNi���S.��#X�v��0N��,��W�ti�]Y��k������&2�ňē!���rՀQ9Ƽ|<x�uwa�m@�D�o�0��2�)1)����T�� ���'Kȩ��ʯS�x7�,#��Y긍�z	�����*�}(��/�q^^��FVN$��q"���=��'��f��^J":�w��Q��";m�j�`!޽� �y$�UVh`�ִ	��׋5�RH��S�#�i��]�C�Y�~K;��3+���h�����^Cs� t�C+�yՃ�N�N�4Q&y���yT�K�K����x�L�H"�ـ��I�A�.���=���/p8�c}E80 �e?�/��J��� ����,oe@H�
 ��Y��̷��<��k& i����ݬ�}1ށ"����x.��t���2wk�G��nUT�5����јݒ�Sg���kq-�_��� d��ɊŇ�_&L�#�艅�H7��a�(R�$V�3t4��Κ6v��v�s�(�/�Ve�������!�p�y��p�G���-�g\�a#S�L��!�c��e��\́/�J���]3���{��#c%z�.#�e����0��{���}�� H�/���(��.�p���6.�_f~��M�D�^Ҡ�ܨ���4�Uv-��a�m2"��Nѫ��Q�8W�3����f}��
�[z*@ĵ<�Z}��*�FM^rY"�/�I"MT��jO��ܰ}�=j��'��sr�lj���p�1�� �J���@���r�w؈�*d�s3ڷi�N��'�x>���C��fGx�����?A�=����]1t%�Y\����z�'��oK;���9B?9�fٱ$`���W���k%����El�=]�ퟲŭ�<�+�Y�e�棺�)�Z`�U�8��/&-I"e6��#���S:����}��� Ѓڎ����P<+p�J�߻��9a�VoV�|�y3W�ʕ^�� ���\1Ek��B���ˑ�}�L��s)�*{q��8�t�J�j Hh�6{8^��#Bċ��d���s{��N~1�׃I�����ɻ�8��ʣ��ʔf��B��['OT8޶Y����$E5F��KO#F�K.T$�,��7�WbG�6ɴ�P��'Q���BAƥg3�A�<It�f�2@c�I�J�g�,P��ʱ�U�yG[F����u�u3Ȱ<T+"�F��w��~������!��qn-/_���^a��Q�v(8gæ�5�of���&�O��?N1�t�)�6N��s�/�B���=v��]~�6M9i���t�ʉy��5^K|���M�՚GO��[�X_���u5z���TW�QoH�
��ϻ������rC/��XG�\�Y��c�zl��E-��)��/EG�r�����r��6dw���JYn��q�e��BlScʨ�3�nщԶ�B%��P)�q�d���{�!��KI�O[��ق>&��k��_��"�B���g�>R����q��\TG�9�^��-��?�	%��j���k��<��ێ�6 ����e�'+r�K��4�Ve�Z �����_f:�C������_�9c}�<�� ��e�PK��/C���VG5^��a�ƕ>
=F��p���7��0~H�cA�OJ:�g�kg���|b��i��Y�(~������o6B���^2�g� ������8SC5���eݸ�I��i�t�+��uqa��}���o��K�j���PG�:K�d_�V�FS����9W������Mҽ	f���E�.��������淢�[��C�2��--�AU�e,����M���ݼ+����M�Y��`�@1�8drzm��I�����v��J-&R���뾂�����A;��7��2����4N��?�Ҫ~�C���0a�%A���{�x����/���c-��T6�����B��Q7�mZ�=WV+��ے]�݉���>�|���������2�ȟ6K豃�I�FIA��s*�Wއ��a��Ԕ��������3�J�aZ�����D�֨x��\1��2�d�r߀ɋ!@�O�tA�c�|���[��5�0���+�2f���#$���*Zd�޹Y���R06-f��ѻ��)<����)���@����N�˵8�7��3���^�R22��=�^ư�,�dwH.�ǩ�K��H(�]s�;00w��3W�|'�`�E	4�WEN�9��)=�p��n��iȢ���tb�4�ҖW�^��'7:�̈́h�~� 
�i?��@�D�>U����5����n��C��Wn/�j�Nf6��5�y ��BM�T�W�x���F���|-2,��]]�&�Z��*�����Leý,H����:j�����?���~���3�bCȞ�$M@�X;V������{ff�k^6�6��U�L�@�'���r�T�����C�Y��̈́Q5X���I�ZI5�;{��n�^����Y �H1�3N�!ܼ^�������*�x��8��/�@4��Y�-!~h�$ڀ�|ac�;瓥3s�5�YDO#Z[�t10�C��r�c�+�8�r@AkW�G��E�I��Ǽ@�U����Z���Xy!��f!j���ξ)�~�a�����NA�����,.`vƽ|(�|5|$�5�x���R����V/���].{J��Fں`��׶�q���o�c�FK~O����͍�_��⿳;s��H��ue�֝��!��Zt;����
��N���c�� �V�q���M��_��6o��t]	lN?&+�I�_�4�4�J ��
�{=�d���gN�.�V�@g���p�j�����{B�!��X ��d6�mw>AZG�[�}Il��-(��Vzg�an�t�J������NYtU�5�S�����f
C�����ý`�&�n!H�Y�V�s�&�@�)�6��s�	Sk�Ēw$��sW�|���ȷmyh�ҼԦ�^�_��K~~]\��	C��cW�#/�h�|��Ѐ��1�%��8ߓ=.�L����Oq���$E=S��`�`�a�鯗��f��f��1�L�
�GQ�j�d�>=K<M,�M<TE+w�3�V�3a��L��Qf��Du��dz�,�J����Ŋ�t@E�r�Q�/��4�:���u n�-ay�&���H}�rA�{�^�;���gA�n�,(P�ۤř���J8����X�M^�� �/�]Vɨ�CFd3�p�M!�)`h�k�-nv�(u���՞����\Lo3�k~�Dd���,'k��$_��q�r�$ȕ�����k��<���R����1&�Z����~d0�J�r�~ֶ'l	h��P`M8h��`�A�w K#%w^�zp��׶m��R��'B�w�SR� gH`��FFˊ�Yr�zC!���w9�>:ηU�&n<��??��QK�����Ê�`�����L
�G(�58!�8��i]�HEă
��:%�u�4(��$��>��˳@\h��d��7]�������]�62@;�3}"���BQ�8�N�<�13�}�*���*A�����&��ϕ�*��O�D�0�NZ'y��m�~d�,RA�*�m��������Լ�}-�o��z�G8��pV���j�� R��حz�͛��`�Y̖V.j�&|��S�V��+s��7
76��O�|t˂���΀�ʝ��/���4�R�f��c��Խ�٨&G� \ݏ��~z�P�~qO0�k� �B~Foꭿ�/��\����ǭm�Ƣ�$z՟q�~Q=oY3�R��tI�9�T��LK�o���Q:�'*C�Fݰ`35��-ŕh�c�J����C}��~���]��"-[�i���)_W�~��w����<&���P��Jg��?����+�M��pb��`��˪_�PƟu�.S���C�����<s�i/��!�:��<oY�O�Z�{�� t_�u��h��K�Z���/>�:Ǟ���� ���'$y7�W�SU��B_\�E=���i�D�3W%��z�_IG[�iR����|r�g%f��ȿ�^e��I���Dyg�?��>c� `|Z��`k@u���8Z��V$CB��ZBݒ`
O�ʙ�g�%#bʒI���"s��=�a���܀E#�0�B�<7,�_�3�>8�n	����1U��t:�r����=��HgG���z.��*$=�M��^�)�`V׳�Q��P�C�kkP��O#�l���*��o��9�jx�=W�`���7���x���NLg5;�v�U6L�����B�u�d�� ���jE� ^!y�����?��<����%���k�����m�>�z7?(&�A�u�D�X����e�����*��х����ׇM�f�c����vu�#��tL�Y,U����u�J�����:��� ���h.�Ey�mL�}�[b�3Q��[��j鍀i�Nx����#�PT`��@�K(���>�1�(X���O�O.����6H��;r��(x�C�Lz���=4��y�M0��.�Wڔ�d��X<l��S���p���&�?"����eh*�_h��y�� ���7�y�z#<��"ϓx^Q���PMg��:���P^2��P���fr#9�\����+,���a�-�ߓ6�Qc�ø�����r4&��@ao_��9\�р��Ǡ���ޢѳmeo;� �yQ/S�\[�'�̽��lӿbn���7-p�F���M���9(|�~4q/����jX�b�����d9�Bχ
ܪ@�uK�X�.��'�WgZ�N|.�k-�弬�G�0�ф/%�'�>�2,~���@���r5�(��/�P��-�{�|���1-qz�a
���M$��������(�^��Ĩ���d�T�rvl�ϼ�R^��d ����#@���#��k���WbR�^�6�&���0",�����ʭ?e$����<��"��&�.��?�k
�f�i�~�MR\=|��o���݄ι_XȚEx�.�La�M�Vu�ÙJ8�阀-�D�%)��u�>$����I	��1��D5�j`'9 x�u���/��V�k��7`R9���;��J����c��]��7� ��>��,��Y�Z�{0��	r��zN�H��5��w�����9�m�x��.5ew�q�"�0����E�P�жm��9���{����t<����AF�'�Ux�;� �R�������Z����J�����2�й�w���(h	�bؑ��,S���5"~�̚�ӅSV���sx1��^y�Ws�q�i��~X:B�J�V�����E���_x�pa8g��no����>#+!Է`�����l�U1#���֟YA|�B�LtЉ	Zq�����?1�����j��W`��H���	t��f�E;ʩ�7��%�;<����!g��s��c"1��W���:r�:��1�� �p�$�`��K�n�dEֳ:����y ߓ�i5��7*[�Y�~�W�G�*x����P�e��FSpO��d$o[��q�\��� ��j����U��:���W��������{�=��Io��!5b���ua� ]�+�^�10�EZf�#��̒>.Y`λB�2�@�����^��?���3p6��|�Yo�]
U�jP˺��2R��>��p�hz�i<�X0����_�L��{T�q�_HX�P���^�z7X���8
�]���[|*��w���]ʆ�	�~&3�D$���4%��*�W�m>���H]�����"������C,	V^��p�к�wz^��ϵB�?tg,���ko������o!�Ze�վ�?X�h�P�8�+��d]y���p�����m�]y�8-@�3�/�~�L�K�U���<�Y*�@�^-�]Q{e$�ޟ�� �Q��7�z���H%B�a�P��d�A>f������!���ˈ[�h�琘j
1E�3k�J#�񡦦~���&�2/�`��iV92�n�|H�l�P�V:�&l���������,-��z���	%�vvj�V�#i�Nw�H���(�?��^ ��k����  ��f��߬�#X{�Q�ɑ��]�JX�@@�"gH���������=�$�h�KXq������
�׆�z�w~SQz9�~:?BoS�5�pu����u�عv�ür�u=�����6�022b���DV5�_�!����l��D�����igW�0:R`�2�5�d��{v���9�Q���`�lA�:n���]׫�y%���"W�zH��	0, PP�T�űU�t���bk2������J�S�t�p�u9���6���V���B�ʙ��9:|���%σ�x������6 �� Q޿���A�Ŏ�[3�Ly�yȵ�P?��YưLH��ۉ��P�3��\�V�����D��=�[���M���P��״�����, ���Q4����j5q��>��0� ]�[��l:�W=�����#�Mΰ��%8KF#p�43�q��赎W�Y�V�(��5�B�%�G��jK���^��C�QU��;O҆�fƝ�SoO1���WPz��&a��b����H}���Yqo��LB�Y[���p	��I�5p1=�A��%���<�C�q��]��ς��^�u^���JA�F��СW������2#��6 �7r���2����T*D�`$�	D�I;g��4�Mګ��fV�Q���a �12iT�فO���7-lm���U��N�4'�{{E�]�Y�ڼ!�'���eâ�����4<#t���!�.+���k����YR{���s���$�2�Vưnf]���`�H�fL1LϨ[윎$x#�x�G������vzX�>x��im�q�� ����wB&h�t�<���XL�"��K���PB]?�D��&�]�m������V%;z�e��l�z5�Ɓf'^aN�v���_�J	#�KX�����E�F�����w�CÇ/{�*��ĉϹ/�6xRl�ϐfY�q���KL�M����y
6<��X4G��9xT��з92��qpw������uC�,��O"�1N�D�3jK ��p@��������%4����LE���l�
�`$u�T�`x���Fo����N�����]ۑ��ªNf��#�ʹ��3m5?�l�ק��.�Tnfn���*	��OpO25*���L��P��V_�`r�ú��F�������!����Jh�}���a͹7��Ty���y�a]k����(iշ�/L��W���Q��_k�(#^��W����}ӟ?v���������
y����9�x���~������D�@g�>Fb�	˞�hF�=k��Um�)?��Pb2ǜ6�As�č��2x����i;Z�5�& �!�R?u6y�^*�I,�qG�#�����&�㖁�H/�e���*i&AѨd���LT�����z�:3^�g�W�ox�%�������䀢ݐ_�h��D^7h���ς/�K�'�T6�s?�0ʀf�^��U	W�&���+>/�s�6�5�^�F~�������&����;���]��������cX8�tt��ѩ����7eT����x�4�K:��ם�&�w��=�uSț�K���L��j+\�J��	.4M7�u1.x�d���|A��aP3Jc�|�wK��EQ�}�N`g���#�&W����qp@"Q�*�6��1�{%8Eَ���&i��)b$�^����s��Rn��4�I͢4e�\����8��_y'��\k+ۜ�L�3[M��b��GL~���=���0��`���Ȯg��Rv�$�ͣ=�x�,a:������hi�Y��)��:+��8XnB+8r�Ah������#P{���;���_�lշR��7�g�y-��Y'P$��DJ���������-�|$��ooe�����:f]�i�㊼�0X��ҩ6"#��y���$����z��̜c���9n�7�į�z�C�!��G�MQ\�$�L���h�5'\��:��'o���~�0<��^ˆ{Qj�2��Q���+�n���5���uK�چ[���J��e�&�cલ���R�do�T�3���Ұ0Y�{z������, ��4���[�"���� �ĊM?<aFp38B����P��\t^���"��_�>kv���Kn�w����Po��u_�S�T�9������J�`��m�}p V�JӺ�~N���ٵ쟞b��;���@`>�L ��9�D	�n���X-��BE81,)s�����*�`����(-?������ N���)���\(�ke$q9v�.6���8m(���%#9��?�~����o�ڤ���W�\8I�8Q�o��G��%�Y�3o��C�75��IC���W�)�@��84�PnA��uja�ZeJ%TS�ڕ�_�8��q)ǅ}`<�C���W�J�G�Ъ
�{��!�9��]\��[�S���.��l�m"�����X��s)
�+�����7� ��Ջ?�܇�S�4YĨ(-�M0G�Ϛ�:D���-��Dm,07�2�1��w�ih$&�U��:a ��9�ɤ�c� ���r�#>�n"Uɾɜ�Y\���.�y�e`������Uѱ�{t�������%<��o;٠z�hI�H뾥ioĤ[u�F��V��1��?�^ K�v����"��zo�,��bb��Ј����SA�3�����.���"HS^�C���ͱ{1����b2^�v�v�Ļ����O��-�Q%��O��ƥ��_ch���r%�	�`����%R��]C���^��'��|�މP���7���{!˳��l��� ��P<�&v����|��V�U�Dp/��,��Ad�?ݗ�pW��b�u��&����ւG�E/v�H��N>�+����aR*�2��_,����A]m��n��}�:���^�'x%����3��F=�8��~V�TX�H$�ڃdt)'�Jn�f^�۳~�yyn�W��D�=�����	Z&*�9d� �����"����pX�G�^�Rh��䇊l0�n��9�v�R|N�?��"Y�/]5������j��`!E����}!�*����`�I�`g��3�l�]�őB�����|`�/{�x3�и2�;r��a��܇�iE�����bk�t�*;_�R"b�{��xb�U��r�V���$��/#w9�;\����.�����cG�f�)���_�'�����gA�������4�!G~�~�U�A���/���W�z\���o.�?�R�͏��m�g���K����3X�ML��h?������#Dh�:��������C��?�V�>~�)K��s@�5;�"��֞ZUY��$�wDS>p�5{��9$V���
S�U9mD�`��tP3[�wg8�9Qw��3�N�ف��j��L�.�ϯςIA�B�C5���0�x��ʒ�Fc�e�	�z�K*4��h����S/�%I�(̜ S���P����q�(��W���T��tsp׸��a� h�W�&]��U"�5�����?-��S<�a��Lq�{yܬ��g<��G
�d�}�E�t	�/B7L�᫮!��曙�|��:'������4�R�H%�Le�I��Lo��4 ��a�T��7�����Ƶ�J7���*/������=�Z������Zk����0�2O��TuM���y8� ��2Ӎ*�l��ëIl1l�6��g�_&���6���N��j4��+��Y��b8 �S���Wqa�����d'!����oZ�~yt�@W̳��W�C��a�4\H�ې����D�R!�
�8L��h��m�����W6"\�XfDɷ�Ӟ�U�%���C��Z��Yó�i�Ζ�Z�M,^�4Q:ub/�;��<;��!:d�=����ע��.��%[�9F�7���\��)QV�Q�z`'�J:�T=J��\ӻ�����8�_�ߚ���Bɚ����S�_��D�"�嵠`c�nu�a��\\Yi�I5� �0���f<Wfj������IVBy����Gm������
�MI��Sze��L�VY�#�Bկ��'�kT�4�l��a���aU�ŷ@jh�*����������|�߹u<k��T>�?��4T˺�\r�g�D��	X
T>u�<�Өz��ћ��ps�{ߕ���V��W2hI�sJ��`��P���ts�>���U�V�?�|PNKda1�(N�[v&�����1���c��҅�.�Δ&WҸ�{+���L�X��x���Oې�����rfL�} 
H%������Z��"�D���,�@�rL������+�)� o��SU�@ u�ژF��w�m�lhF�����5���TW�z"L��`�o�O	H.(2d�n8/�=�	e	���]�T?p{E�ʺ���w�qN��Kvݝp��Q߉2{P�wL{�-o4z���Fغ-�ƻ�
1~�nh
p��m0�N�=��\�qR���e
����N�(�Q�C�}-OLa =�*[x��g�F���֟�yGܯ�?Հ�5��������O�V�մ?�����j�;��I�:���P��H�#,��/�0�
��c��3T���g�kr�PRD��䥜kg�jB�A5�V@|��b�8�5��믶WI���H/hjIV�|m��	|}��:����@X���G<R��X�G�L�F �����f�ˋ�վ%�bg���Զj��&@Ml�十�>3������mʟ������<%P=XU�#$���o��x󡔯	y��/0��'����T���*Ӭ��d�9�Nd���#��$ES��1�����E�!Oܧ|si����4t�{~絻���Y���$���En���G�aL�aӆI(ژ�@՜6�>�$ca��=/|�i%�d��b+���%�u�0U� ڑe6#�A1���]���:I�}x�µ���-��e���ia�`�"r+~A��^~#W�bDo啟����jUGqFUl��|����䛴�)����?E�;\�2c�c8�Kk�5�z��Y{Ϙﺥ�������c���/�}'<+���e�X��r�`I��!,&�����?C�_Q����^P=����y�7 � x �k�&~��y�u�� +��h|��E5��^�s8�g�نO#�W��#(��N�� VM3�}�`�j ߹9��D�y_����P?�k\����M�����wI���G=� �����,�!ØۉE ��,���?@�7���Cw��a���(�L�#��i�uP�kS���Ww�e���,8���!�F �^@٢� ��{�?�����5��뇮<Vϖ+�Y,���|�������cy�m?�V;R��R��8�	�����R�g�s�[��G��[d
��C+A9��f�"��K�2I.��?|�ȹՈ*|r���'W�S�*��3		��)��һP�����H�<���d��>��SS45G� 0���L!7Fl:$]�T;lĖ��]�!y� p���ЍI�u���9q3e���8�&O8�@��R������3e'&��,��r!BJ��auc$�-�V�3雉��0{�eM����J�v�~�1�������40��Y��JYC#{0�����2xb�es��E}$픕Q)Xy�r*�&��5�����?	����v"��0ڤ���b����0)��ޫ����!���P N��#9�:���p�^�WbԉQÅ;�6h9���)�'��x&r7�������$�fK|Ntj�n��*��ީx�{�,'J���}S_�U���˅9���i�-2As켰��(@8�)������(���B�l����]����եr���z*��)��?��ڥ�to��'0�l:���Y�#sm��F�]#�]ȹ͒�t1g@�S._S�%��JdٟGBԕE�|���.ޡ5�����X�XK���n����^Z��B�Ua�	�%��&3vz���d��0�i��� p�[Miq����yv�쩐��(�n
+��E	R�1-�iK�x3z��L��>
�My��l��b��&ix�A��3}g3O)'&n�I��Y�^�cz�yn>�3�		%���,�lVm�!� P0�q�.�11c�`G��\�>�o����k��}%Ay���Sò�ߥN&��S�trA�bCm��>�5ک9�_���-\�����*%&�tS�ib�����y
��],Կ�{c㬝�J�r���o7j�I����.�h���s�2���;�c�$1��%��I����vަ��x|��p����L~�t�����
\����5��<Sꢫ�:ut���a��8ȹ�7#e)���'�_y��<��8�a�T�>�â��(�~#~�l���bX�3Sj�M"�/b�cXi��D��k����
=lǻ>�,�)���RhZ)�^�-\���%�D��@^*��)QSIxf��{�l��s���<'���XV�vz��T�&�ӂ!I��Ҹ�	�X36�F�+�lD,c~�%�W���u���ژ*��ۃ���op	*�ب�
���a�M+�8��x{'W�<A=uiq ����^�6���PK]]�bd�h��b?i�Q�׫3�6/��]�j��G�0`��3�|Ru��:Eb�-GHr��mxv�����q\�@5��G&S£c�����<���c�ߨj���Fi�Y%qJ!6I�}�#��wF�h/�;����̖]�Iho�L��2D��R���e`pH�>�gO�VS�*�ƒ�<R��r���}	;��9���ȯ�Ej�& A��������S�T�u�O��Σ��c8��H��$REg� L�Ƒ<������ģ��y�kl0RHJ>m��AS���з_�1���ˊ.���O��"�Uu%���)��$n��we��b���8��ᬢo?�ړ��ĸ�ns�\FR�D�m~dMeF��rȡo�v䟏�;�1|�����R$՟�ʵWX�%�a����s,��g��v��`<c+d`΋Z� �=����	��g�1���V:�O�ky>�9�=�v�V��c;���-��`���.�P^v����x{�0v����b��{6N�����295!���|��Wv.Q�|������ׯ��<M�z����oDJ/�S��^�QL� �w�e9_=Q��y8?yO'��Y+�:
��%JЪ�FW$�>j޻h�+�~�ءҦ�����7b�wD����p�Ec�]x�Y�9����xz�f�{Ñ���v��"��!1/����)��5�Q>����f
��?��o�t� Jk;�*xLO��Q<�x0���Rd���-E�Vc�g��-B=��Чq+�9bs۝_R���$�p��Ms�(�6������ IaNl$�	�C�'�d3��ִչ�8��p�q?���ș�c�+̘�m[� ��l��P(��z]^��^��h�C�9���W@��/����X����F_����n��X�VN���q_�~E�T����[c��T�뒢���\b�g��@���3�H���Q*.p�say%ì��"��\}�&z�NM$h�.hu�:l�	�s���C��[Y��ɹV$����T����fnv?�C�#���!�
��R�O�e')�(��S4���s��* vG��KFU��nG0YC����J����<k�C�o�f�K$����H4ܡ��.E�\�%T���t�;�V�ua#n"z1��q?�o�k�C��i=�I�t��~�"�V$Ѻ�(�gao�	�����8H$X��a!�&�Պ�i��hT}���7%@�����׫17 ;(w|E��P�O�: �����t�����\��S3���<yNOr�������;#���|R�\w����eR����P��j�/�=:{w���ﵕ(����F~dM��!�?��C�]�5�h��MPf��ѹ����僌$q����;r�!mJ,���=�:�F!��T����Z�P���pPϖX��8�]�#�	}]�&��k��2=���5|
"��;��5��uX}��i���:n�����Jr���$}I�\#A�߻��>*���&��x��;�?O垂�Hz�ܔ9�1�������OBE5�}=QT�9�^mD�R]�?��[v�ai�(/	�T�HK��rd�L8������M>��Z*D:�,-CU|k�� X����]���Cz��PS4BI��<�$CR32��>="�(0��Tn:xF�Z�� ��]�Q�N����%s�m����ZaP�0�g�a�l	N��5��U�=�#j#��=��:�gQ���;"���Gi����<��(�7���B����*��e���P(�j��)�l��,�g=�Y�u������-^���	���s[�����S�$�w��X�e�����y�&�9�Z��^�`M�"餯�ʤ���es������Z�9�G��q{�{�f/��-���8ԃ�h��^?�:
�Ճ^"<LĨ\�]D�0�@�����h_y�$�I�o��;$X1������.)�
�=�n�@�[���ݼwl��Ȝ���!n��Z�9d>��
�H�R��\�%5�b� �6���Ij�7��� ��bמ��цI�B���>�r��e��:� GTab*��=���c�(u�Ӵ�K�]ui�2�]�N\΄����8c��e��Ik�;�\a/������ZZ_���^��8i�w���cx�w8�l57"b�0Ǻt��
~�[1�?����v�VJm����v{W���]�SЖ�e��≿e�8N��t��b]8�Y6|���(����zg�iK�d�y�y</��2��hi�tPeQ�p���T�������| �bKL�iȿ).D����jL���j`��ú��i����`��3����ŷ4j�A�m�G0h��߉��U�0nbnS?�A�%�#��l�Z3�%�i�1/Uc�L?����b�S�s�(��kU�&���뮳ȫW�0r�3�2�cH|�*Q>� tZH�Q��JF� \�}��9�����o����d�(f<
IѸ�%����Z��.� qxq���)�zxD5�1��U��n0,�Ђ��{��V�[�{~����!�R����%^
����o��Sk7L���;���E�%[�G���w3��Kl7�a�B�G�θy���
U6�B'�5�U>��o�f�P&GUCJ��^r�y��3��j�@�v�Z2�w�5�#f�~��l��Q����R,z������!�D�����w�B�U-�p��g�6�O3\��j
-I����::��-�� 	u��g�ԩ�N���Ǐ��ⅅ9K�� ]�g_3�(���t��!^Eu>�%��	E?]߸�;���m0���#����R�dB	���7殓�|�$F�Y�e-�h�F\	��[��c�@�z�HFǤ�)�l76�X j�Ώ#=�1!�����#Y[ƥ-�֜�{�)�}�Kk,���b�����?�g܎�W��d[i�zk�O�O�YZ���aqC�s=έ����8F�/��b��l�s��	{w[V���&E�{8�\̶�`�O�G�1��A������,V��E:�:īEvNX#ɘP�}Va׀�`q�&Lzi�pO�3�h|��h��_�����V����A=Q���I��(�&2�~���i8y�ƫ��;���N�@8��n�36����_ԭ"X���+?�G�ѭ�$�������+~)#ۓ���S�R[+��79��@�Yo��'f�|U��Շ(-��R�.�w��?a*���ޜH��8�~b��?�n9�!�����r��f��:���W`An�oJ�������"_��H<^�q�<�K�Eo�	�u��ޣɷ����o�G�rJ���e�_U��I�67^6��2����" �F�c�s]��+/�a|:�n>�����.��w�{�����`A;�%T��$^��Y�?!��� ʧX�bd���9x�&A)6{�X�@\���-������>�����u�^����n��V��x�Z@	�d��¨��ξ�EIa�҉�fy~dH&�9=5*�B>���T�)v�o>/��k���e�n�$���"�0
�X2U�0F���� ��7�@�i�Q$1�$��"o}���d@�Z|/&`B��@����H��t��~Ȥq�L��(�-���;�����̓W]/�{�+V�žw�`�D8t��g�b*f�>��U��֤^�_�������j�>�������{��X��$���~�D���-ʍ�ޮ	 @B���(�o�D��$�Ta#��4�0+��N�Y�Bg�����j�Y?���{HB�Aa�Ze2��mC�U�4��_�m�)�|�����Q�ֱF���������oe�t4H���O� g?ʏ8�9=u�*OK_�ǣ����y"�V�S�ʙ���i�搨�-"+��^wS
6-j\H ӗ��y;+��6&��d�EK��z�̽X�Az3/�!��]+��K�[C���ug뚗j�����]W&�)�PG'#���_$�j��I��:����b�������㑟>),jHp?�!�=�F�&/ި)���Y�^��b�Y����č�E8���� Z��6�W�	)ؘ]ĊA��88�>���2�]<O�Yԩ��V���Y�ŻUB��P\�ַ��-�}��$߂U��R2�>�a�k��P���'mPs�͓�V�]U�}�:_��D.�������O��]�ճ�����A*y��U�X4��.�Q�wD;�q�v�uj6�P���F��(u2"��&�H�H����h��mY�ol|�L/�k渔�������@l�O�]���ء���V�l����Zq'H�텳�P��*V5�r��+�V�3��ؒ���b+̬���p�����،Yc@pru8Ā������n�̨��6��\Ea./m}EpVQ��cL��t-v.�4![�CÎz얤c�-�Xszg��3	�i�/�i�$Q^^�zEw��J�`�菲#�x�|���ų���X�E��C��F}:�+����8�s<��pIL����?�W���]����<VP��/�������+Qq�|*�Rr���mN9�8ݍ�Q��J_pA]�� ��|���Vʼ"�d~QW����>NnثJ�Y�<]b3����͔ҳ�U�	�_���2�t��rB���Kj.E���Rq�ů��f�Y{m��R�J�b挵�<-���P�3��u���/�%���f�(��(����ϐ��n�H������3h@���A��&�#����e��� �y
�x�S J��_���vk`��a�*�x"�C�־�� �
ˆ|AhKDo�$��W$0�r~;�]邸{y�l���p��Kr��@�)u�6d���9��0KR"�o��Oђ��"��S��.|��� a����#�@��oӈ5dТ5�����[�$���X[����E���(�	��\�MK)$�����;B@�az1�?�t�8�
�ߗ%�v�q2��z�6�Μ���/��D��|�ͺf� ��7y7}H>4���Q�_������ߦ�L:mW �2����0���Ź�}������D���~DK�R(�5,�����N
�;Ee~g�1.̰��?�΅��rrbg��?�g{Θ�)�0)��4j� � �-����h�p�9�G�&X���)�����"�����A�A���6�˅�wAx�b���8���G,�lj�S�����>�OV��x���o���V���Я��#q�t�粪#���kb�������!.���h@��/�}�X��e�k�ЩB�s�.V&
�^YY�Lm����|�j(h5�u��V���N{8����4��'����ȗ9�<m�,��UR@��Gۇ�S�G��ӈrDE6i7�X����΍�6�G�-�Ʋ��)�{��]���7 7ګK��������?�BVZG}� +�Mb��$�}�)v	I��!�o�~����Y��k1LV8a��	��������%���f�B�������C�գ��o�yH�Ȅ;d4�_���E�T�������a�r^�h����c1!��r��S�{Tߌ��������Ý���g��1|�I#	6C>�%�ˠ����+�[���T�7،�:4H	���iX pX�m�A�����שyZ� m{��7
�<��ǖ�s(B[L^D��Xfͬ��]"_yx�s����Bk$?�I2�n�6��W��'����-���p)�l��Īz��"�p�e�(BD@{\��0�^|w	�k��ߟ��|�uU!�~�[���T=�<m�Ֆp��bȞ檩�+!tS)��;����2wxӲ��T��>��:��=��z9{�%<ϲ�3ޔ�C/yu���j[�{s|�ۂ�����(��RB� p����?'�h/���,�}`�x�B L3bP�"�7���AM6"�ˑC׊� �8��r��BzQt�௒�_�\kp��Y�vmc8���y����W��%V����b�ݢɴV��4]�����-Ow ˰;�����+8]cYV�0,$@�mF ��ڐD����ݖKv sR�,![ڶp�?�j[��K�]ʹ6K,��;���]�!_ZAg�ij���M7�-�6���e��)�2k>�܍�|���4y��o�����w����<cGbR�l�&al���o-�n���A�i�v}����2!5��ۧ��vȞ�^rJf�"�}2�Y�l�?����]����|�S
&��tq�W0h��P���o\��{[���*(%DJ@��km���Z��J^�y�I����GsStJ1)�>��8��,\�Y�]˂�f�C�oc�ζ �2~ۈR^♥�L��E��@h=@�;Ýe?(�Ӡg�iaUsY�o0�L�,FKC�_o�-r\��(�?�������u�~V��Dg������<8�;�4>9Q%��A����EA�hY,�қM@����؏���o���o<l#�u�����ґ��鳛w��8�L�����:�����/hy=��5�q�r(?J�{�J�sBY���6���u���8��&M�p��ww�1�%���q�o(�1��k�a-��N��J>��N��Kd�#kAA�"2K�c�D���"iXj�)�����H<��,(E����ʠ��J�C`��X�X�����e�APAa��@�G��E=����/�Bڞ����c�S�<�ء����p��N�b�8 C�iO�A�H̀�����:jQZ|Z����:�ʐ��� zh���zz���wF����1�������4�U"O�����YS���=t�X����oBKb2�a���^Ps#� ���`���nCy�0��gv�K���!I	��[/m�pZ���=��>S\�p�;����dN�+��Oy<Ywt7���z����r�n[��B��, ��gغ� 	�zwԩK�%@��z����b�41��I��u���=L�K^�B)�E Թ�I���~,�б����>��K8�g~��}q������>P��X�Y+��f����bCn��u``N�U�w7m�>a�q�:hDW���,ݼ�e�п�D�L�ZZp�(Qf_�q�KIP!��\���or�ܺߟ�C�(�����v#c�cI�q�࣯Mu5�{�t�ʢ��]n�:�F�eN3M�����E��6G<@����A�:�E�"�@��&#��ҠaK��O|�����U��Nf��b�(r	�у5)}�!o�]`�@�}1�O��C9��r>����+�E�Y��D�?u��<�cɯ֔q��RQaƹ��m�/|o����N�0��I;-\k�d��{
L�E�ʒ_�!�����F���v���V2P��o�J1V-ư���P���\:����y�)Q9�@���E�̨b�ҏK`N�F|D�[C�O��!k���
.6�K�
��4�I���Xm�������jo��٭�l~׷&�|�Ėg��v(���5��l����d����S��a�6�eF���7K$��"�U���G��|O���w2�赁*<1�;�#��Xz̓%q9(��J0~x�Τ䨹#��}Lnв�_�t�F��	s;��Cr�O��M}C��q1�˦���ː1�̐ރN���z���P.�`�#%E�ߜ���lU�$rYP����M"S�lz�S��2 >:������;ז��̜/�E[�;���2%hҞp�7�<v�AK��ꁉ!�0���e5���m�h7�\����]!PX}�.i�پiaK���@��6��{j{�C�����W��@x�~�N�;d�.���)����.�H�/\�X���3|P�렗Wq��i��@�he�<�����&lQ+̇��S�DM��O���	��|�3R�.��ۭ3�?c4�[Z7�Oɀy���� =�����((ru� ��.]6�}���'�M솖���L�x�Ҽ~5�����j�W]��!S�O�r;9 P��\�\o\���À`���L�J���|�fC������\�PZfk$'��9ʠΏD����DH���#Tk�y,m���F\�s�x$��4 �`�`o�%m6y���*�D�����LVpb���$�P`@s}a�O:���Z;r�q���B	M�߬���ܴ4��h��q��Y�X���E[Nƛ������Qy����N:VI>�v��G'�����ΰv�7+!h��J���FF�������t`�>�k��j3�ӱ�Y՜��kPO�xmP]� ����˭1\!�C�r���ߜ����&*v�CO�0&���
RG�\M�c��m�~ �~B�]þ�Z�Ḁ�U dDi��#��Q���:L����=���S���%��}�Չ�L��jʶA7G�1�3Py�
�|�d��wXh�C����Aӥ�����X��MK�;*�������+,�SB��|��i=I�G��d�o��=P{��
�<�ߌ��ￚ7<�#���&-��p-��[��6�U��X�����@dxL�;�,ާ��#ZܚS�i�aVTx0ځ�<jFa�����&>ʴ���N�����Dq�?��qAlµ$��у<h����/�����RX[�V�e~ρR�c�>��=����>@��� ��ѯD�tkײUd��N�-����@+ q*p��GI��xɮ�~�����Qs|�>�l�e�!�ӕ�淤@��{a���~��{FA|��f5o\�9��#���8U8�g�I�p��Vn���q��ƦĈMy��$bO0�Sz�QҎ�0ř�Vj�y
�M�lF��¬$�1����r֢:j��
�j[`�P���i�΄Uχ=rE8O�32aVɿ$F����)Z=�'�}�ɯ�/�)¢`rt^��W�ui&��^-<�7��+�0���6~{����8�~$�b�Q[�Y��l�\��	-1��v����vS��$=�4�PĎ�NK� ���7�/����Օ��6���
,7ia'�3�roo�O���v��H)���!� R��:�0?b�;��z��pbV�*Zfr���g����.�If[�X�-��J|l\h�Z��ѡ�Q�ٚM�� �u�$�	C,�?�~J�#ؕZ�H�/'��z3
s���HK��,���e�s��ǜ�l%�l��o�@����}3�8��o+ZqU�@�^��&)cp"�Q����+Xq
 o��	3�$�9<���O'�쀼�i�9�?��ؤ���cBR.���m:�"����cc�����Q��9���`�����P��	�G�>�d�C�Aۢ$�?����Tavz~dT)`9����ră��f�Ȓwm�f��'')�Ǜ���u4B_u�׍E�6<Ay+�+W�N�l&�]w��O�J�t	6a���rf^������ԛ�~p�	�U�)@�nm��ܬ��kA�}>����m�����JM�ΩV)"�^�8843��F	�D_�|�$�Q�9㥴�� ��F���Vܫ�8�8�h�i3�2��r/!����zͪ^jb�i�L��;���0Mеɚ�~o����،!m_Ȗ�>k9PE��lӽιV�����m����Qle�:j���P7�2��"���k-4���Fp��o�Ӫ<j0ҙ�ڎ���`�D�n�����,�ը�k�\�����	���/�L���� ��ؤ����gb���~�I�����.�k���fy^4�u�Y��х��A��ݺ͔�����'���\�O"7@����8�_������hH���e��/���!��i���@�;�Ym��t"���YQ���x��3��oYgvX>d%4��w,'/�C�`��nT��c�C��2�; ��B�*���wV�>9�8uL�]�!��z���@�`M��7JA�C�*D�g����>΢�{����tid��6~:��r;�H��%椳_J�������$]���m}�<���,F ���I�ooF�@l�0{ryK�D@�h/�D˄A�T�X�"S��".�$3��+�dg攄����S%)��T���=hEM=�k֛2gp���%�\p4���F�OG�h���S�_����4a�S��f>��bб��؏��i�/#��K�B����p��~	����W�����,)<D���T�8�R:�������/�7_L��R�f�b-��C�������ԓ*U�?8[%���b�3w�����{#��o����bD����TT�p eq��W~�@��Wg�^D��2)b�w�Jq-#�!*I�@1��z�.;]��`|'E��al�&L*2�f��0k]I��f��v��7G�G��_q�~�
8�V
O=U�{(���H����P����.�N8�9�k0˻ް�{��k�p��:���`�2�Ց��_鳀�>�ͽ���[��lWV��O�(�4(�HlU0�Y0�,������(-k:�[Dr*,����xw�����B0	�����0l�>�	��_Z@�	��5s��CX��ô׏jp�#�x�{�HNc�s�O��}���gfaۭ�&;�2e��)���^���oO-	B�����A��1�zǭ�tձxN���%](�B���/v�\<i�B}�A9?�^��x��x݅�t��g,�9�m��l�u��1x�'g��8[ݠ4e�+�d@$��r两tOZ�-�@ݢ=��z=�]�9q��Z�҈�oɓ�yV�]�Ԝ+#-!�I�8!Z��-1�i[	[�K����`U�~��c�-�'�7f6̚��(b7�l3�ڍ|�8{H�oo`�Kq�C�,����s/���
`M����O�6�k����9��c���B��>�̒�$�pnM��r鹷��q����F�8���UX���9���KIĀ�4[G
�鷲�G�n�WQ��|���L-�x�N�,5-	n��;W�h ��`NA)�=���^r��^Bˏj�~-p�s�R~3��Y,[ľnn�0ix;�����8k5T�W�;Є�������E��(�Z�r] ��:����N9_3��юw���%��Bfa@I�yѽ"�{;�I�b�����i���d��"m3�Cg�ജc�>�Ũ-���P�|O�����Nv+��,e[�b9�pB�-��+�wd�Jh�a�S��gN�s4�im� z��`BI2����R)S����r&��W��%�CP�F�C^�(����|���O&$Uj��Pe�e�N���?�`{�WǞ�#��07���[��ÄT�f�oZR㥿��B�e��#h�g���>q��J�
`2L;^+��r+}ү��Ո�N��Zy���x�N�T:��E��VP��{�1;��!P2�M?÷��ϐ�K��v���8�kV+��?�F��ZX*$33�қ��y�/��\_֣$�p�h+�N}+k�W�>��ʡ�(����6����/?�4�-�ck�Z�'���ES���b�e�_N��4�\��T��wɭ��O	?-�A�I
3�/D����Vz�@�?��D��U�~E�|��^��
�.g�$u�a]�7Oˇ�7�Ar�yt��5}:q��8n�ݤ����~6���+*��9#H��������:�#�z��P]jb��)����$��7�3.�J��?�U������V�ߩ�Tu+s�`|�L(N���bХ��<h���o'-�}��8�'uuԵ?��q�h���K,�*L���q��V��3_R1+v�4	���;FL%ݬ�o�p�+6ϓ`Q�O�Z��k3U-X�S�M�<v�K�zkƯ��o�"�C�9�B�Y�����]��Fh&>�L��o�H��/�C�<�)'�@/2�ƞ8�|7""��9(:4�S*(z]I|4��~���0{��B��L)ɿU-�^��3�3���}��-4�	�@�Q*C�z��e�ҁ������ob���
\���oZ�'K\2f��� n&��I�y��x�hP���A3c"	:�}{P��~�w��,j�H�s�}J�1n��՝��Rɉ��
�nd爼�x���Z(m0�$���*������\D#�w�;/H��p�u~Gm�Q��8УO-�?�N6L����Y�^���eE��"�n�sL.��������+�D7f%����/�X�>/�ivlB][Ĭ��z�,}]�2y�^uN�F��V#_��1[(�?��P� ��Λ���!��F��CvN���~�k)v�5�����ʟ�ccT��4��I~I)7x��՘�$O5�V%bԕA�ϻ ��O��QVq4G���D�l2���
��'�Ԕ\��I�u�1���:�[v��]����2W�N�����1I�Uً^�R�/�6��ɫLn����w�U��d���[!o6������Z$`����g��N�2���\zǡ1�O���E�/�MؒM����=Y�36�En�H�o�ށݧIR�`��M���ِ �@�I�8�D�@�����gWb�`�BO7��!��p�"u�Ȇ�>A|����>�M:�ٿ�2�Kɹ��J��}ns�d=��Ι>�&�gka�憷 ��WK��&�m�uc1M>��R�ѭ��u&�ڐQ,����4�'�ng�F���W�ی������"���hU'������GH�+0Ox9ݲ�-�bhc�vTG������T;����z��1�Q,�١}b(Ű�g�֡"�h�̬�_m�%�j�C�����[��.�d{)h��
��:E|w��P�h�%��2 p%�t{� �~�)v�M4���LM��vPv��mD�Q{e�ŧ�-:�D��<��1ݰʛ�4��>"�!���$�����o���
�O���	��Z�֯���������H����^��W���T�R�G��:	H w&�TX"迟~!��lڬ��l����) &t�f��d3�:'�%�n�B���>a��{\���ǂ+جw�#ڒ���b����,g�޻?�TP)\]�d��}�	��7��rQr�=^�]s);�hw������0��(H;�J(��{�f��D�����Qh@�F�5���Q�r�A ��2?/���fP�(��/������5��Y�M��`�Pss�jN�U߱�����}����l��B�KaMG�J�0D�~����V�܁�k�{�p�xs���>"	��=�b���ߢlS�s�4ߐ(�?|�l���2�%� ��f��3����^�=K�eι� 0V$��G��B�m%� .e�0��M���r넢�9x�z�����%��L'��W��S�R�z��#{����\�(��*� ���Y��)X�
Q�so{r�<ې���
���y�$����N��2��J�(����<�35�B�jy�AJ���h0VQ�Ђ�MR����2w���Mu�EP�go�A�i���^�=���b��)&�R�i>7zDa�p��
+�̾{Oƅ+N���t���
@�2��n���,)#G��$���؅ � �k��_����|.+c��D=_k:p��j�N<���S��ɋ��r���U^Z������-H��S4���KG�CxX��a%i5Z'�+,�@�A�7� �zH6���uuR�O`�2@5�^)���gAk������
5�(
/�'�R��r��f��{�{sO5ڹ6��E��Φ�����B��q���
��:tKte
;��ڧ��5��V4έ����E�S��n�zlO_�O��>yަ�2�hG/��`<�4M�fF\��I���m�lϱ�B����pz��؝GDs;;��_v�5lf�W8���m�^�2Q�,�hf������[��qد6��C�s4&���"8�d��2>����&��̌�6e~��|.�Ɓ�g�)��˯��U/�7�/��	������C�<�����V�T�P�uC~=
���.tJ�s��'�QIlLS�c ;��w�y5���K�d�"6�#*K6���3ꆼ029�C���L�A)GJ�͘�7�r3�?3��CΓ]��>�9���2�̚E@�	�1zy��MY6��xRɖ��9�^�}u������t+"k�,�(����{�L���+��re��m��}֣3A|CyB�s�\�?���C��ì�����T����&�������x��%�I2��C�O�ٓJ,e�[��W|�����y�O��D"�jB��|[v�ݻ$QR�AI�\�o�C׀�i��*���e"ɁJ���Ȏx��.�<UKĵ
��|��Ps�۝��;-3�T$���9����:ϗŊ���������3���ʨ��K��t'N _�c�lbH��ų�f�p�6����8��:b�����+?ޣlh�p.���ȇ%�C���=7����%&�tvm;�}�Œr�w��Ja���VkH��@����J���8�� ���A��s����>��z�~�0R��}I���1���Pq�C>r�Q�0����>�	�.ڻ���xW��1[�Н��S���~p�m��j�q/		7u!
�@�B��.�]p�4-S[�W�T�^nUXU��C,��o�͎`�H�6{�d����8V@���\0�����`�x�Vn�,y�T����v� �Ը��%N8��M���B	������g�k�����7��=Y���(D���)3��R,Ol��Ĉ[��H�_w^��z���4T��\j������>V�`}+����v���R�!;�vo3�rRTx�����B�r��j�B_�́1M���n��0LkX�0~*������J��鴭"���_�Ɍ��t�;�ͦ��Q�+��Q7���[��&Hb��z�*�B�	��0�$�C�2@<٫E6�ߍ���6�/cZ=���l�g���]tbDz;+.�A�aW�9uY���X�ۀb<��!��h������(t�"y���gȅ|܈.#lm�~/��VY1;���&��l���@�*/��q4$�>fs���ڞ�}�����˭�|Zp=�;[˸�us���S(BÙ]"�W�-��]2Gmo��:�AJ�7�I$���}:�B���c_+϶��ha}j[t��{��:1hσ&P+�i�Q��WP��E㊂�ĳ�T��hU-�à�?MA�q�$�]��g���Ӎ�Q�i�W����u$�7७���	�[3��%��z3sT��qi���W:�u�'�F��8�3ΕB@��~:�4���b)X]�T|:��;�lD������;�
?��n��+8
R���F�uH2 ������ �O��%�CU�Ɵ��O��S4iOHq8�̧pd���e�J���y����f%��f�t�J�N[��z�������fV�Y+s��ZWW��G��-���@��zӡg�}��\Z-�0 ��&�\}�v�Tsj2[�ݷ��p�µX}+iI�mٴ�'�p�Qi��ХҎ Q!�^��+� ��n�����Ϳq����q��(��V�1��U�Ah�ᰁ?E��2+ܯ��T��y%�i����꥿
ڦu(V�/�0�H�����Hp^���30��A��I�ΛWb	�����A�";�:�?{*TS�����J���K���CI�E���7��V�)Ѷ4j�)>q�@7)��)�R/×�J�]���W%��	�.��N��;���1�j�,hC�`����1)��qβ�R]R-��]H��
B��y�z��q����-f�עP�@�'��
ǭ�\�����|�$]��)�������`s���)����=����ڈ����Wo'�
q@HK���W18��}���)h򹥧�U�������VbSf��a��Ǐ��ug���+����شԺRl�M�_��P��m���8���2�P�Ot���Fc*u��|rS�P�����e�1*��>`_5�CR4��QY�]����� ��2�q�,�gA�5X3+8qrJX����u�����ޏ�G�'�~��]���zC�`S�)��ٺ�U�_D��b�� �X����yU�ɰf���yc�u�m��&@۝2:�eO�3�R����_��������t"�Q�ӄHD�Q6��}����t!@�i��o���d.���4���N�{j��_Gn�5B��6���v��:��W2:f����Z�׋c�a;��S�V�;6BP���jb��������B/,Iф}�I}�D��o�V�u��Kw�>�9x!)L=}h�z:�:�u`I㎻�X��'U��8[
bCt����*s��B
�,�2k���(��1�삨ʴ;�UEr���Whd�7��砾��������<������D�iW�|Ӱ���{�ta\��g��Ӡ�:�՚\'���j��D�Ez'Ǆ�K�s�����O�?I�W�ÜQ$/��;m�m;u��a��S������3��L�E��Ϲ�\w��7ǲ.���1u"���a�#�(8�t��d��U��i ���7c�#}�D��L:ďu��a�Z/��-�t_�`�Xtِտ��̺	r�Ð{"F��F��.L=!��1Ȥ��x�v�ؘf8ܞ+r�����B�#�B���ed��ߣ0����Łwގ���5d37,�A�h���V�0�
��3��h�o��x�.f�_������Q�*׵���zv�B��	Ha`�,���jI桮�M ��H`�L<Z�0����J�#�i����X"�̔�89;�$pO�O��pj5
8(-Τd����ug���\ ȏ�h�(�ƃ�������*��eQt���\��ud>b#�m���*�CZ-WK��g]ղ�J�(��
7�s��)�v�f���W?�L�����Ζ��Z(p>��0C�A�ȏ����R:��4��z�F@K�6�yf��Hwޫ|ւ�;�����hc��կ@\<�]aE��%c����\ȼ)�(�_$a���6B͝�wR�a�������x.)M@$���"�ຬ�*�v�-/+���؝Ju�N�n�*Q-��(o���Mkj��pw�7����?�S��ԱE��-N���	C�t��gv7>��dE��\ȢX��~���4�����!�sq��ö�m�J�R��3��!"5���A��yj��n�'���'��e�!������>C�Ax��[r��-��Q�/��yҀZ4Zx�A)��B����V� ����s�q�~��u4���)EVﻵ��J|�oJ����g��᠆/ُ�E���ڳO[3���l�}�8�QT	�D���߀L�	.���շW�ќ?���[8��i�}���W���y�C�{�~�%����ԾI[�oi�t�;v��Y����tWL�:�T���A��m/�&+t��)]u���դs�������`���E���^��ݿ��_�w�ة�U�S�y���:l���n�v�}�V0���(73�"U���e_e/>�&0
ó5��>�������c0��L��aa�L�8I�;'�oOO�/�l�����O�m�Y�j�2�D�i�|��14�'��9Q�z�3�C�3�h��&D�5Kc ��Ժ���&����/��-1��L���o#��@�E�좤|���X�c�K�*Gy}�좢
`��3Mc�[՘�zDdݡ�h�#D=��t\-u����M����������ɗm��R!	ui��T�f�?�>�2�,^"m�GK���}�����dU��~k��O�%�׊��@�Cf�q�j��q��b9�n����l�'���-E�z���>^^��?����:@�X���_ ���P��UMN�y4�|ȩ�4�R�
�nu�m$�{�ӱ��'(�6��,��Z^��{BO��?��b��i�N%��" �ϊ�L8x�E+��tp+'
�ꋈ�;�dgAt5wv��@+�s"���y��H�x;�����(�(rV�Z�Nj��y�u�Rt4��d��s��O�4��&�ǡ�G$f�X�7r�M�+��TO^�V2VkCP����X�+J�����W�ih�;g�ӳ���$2�b���_��3�p,�@i���~c� �98��w��1E�|�/�|s�J��J�7�g�FSD�f���!r��.��\��y	T�-	�p�K#&��ӓ��)Nl���.li������L����f.	�ou��&ߟ0���m��Q���GU*IU7;��:O�ޫM�_�Ux�#�n�̷)\p��6���?����n���aI�$�h�����4�,0'$dʬKdC~�q
J]����V;��꛱��@'j��N�"��]cAdH \e��Š�EM��4����=#c��������k�,�^�HN׫����}�_��ys�)v����Eޱ���!��3x�i���ST�V��,J1�[�@Wԋ"2@ �>���Eǝ�fs#I����\
�(v)%�ߒ�P���ֵ��(���o~�<KL�.�ð�w�B�v�\������z/*��b�i�D�k�C�����e��Y[>�?�:.U��{�r�
���b@pp�4�_���Ԅ��I&�֙/�kf�󤌥�A8;T]	��t%�N��W��V��]��&�B^+��!a��)b�O���� L=��7L!1�'5�c.��OD0����D�{�]�ga7J���-���=�'5��9���=pw�}	Z�\|��0��v�0��g�&��k3"�MsFTӁ~ߢ]܇ԙ�}�{��	�=��jSW�Z��lYww����R^���ńڻ�&��#�0�O������&PX9�)e%k97o݊��8z�,����%I]0���̇���(�$`Z<pS ���v������������C�t��&��1�~Ϳ=+��4�x����о����%`T�����K����P���XǍ{U�h")�9�
�֬���]m�i�}��⥲����Ym#+�g�Lg���{�K&�7� k�$0������Ǳ;:~���L;��D6ҭU�ww+�Q�����h��(�����!r���t� �tf�-�rb�	s
�}�}F�w2��X1G>����������n3/��z���zOoG�iN�^T��<}�o�&��w�L�TY �7��)ke?�u�j���[؄�;��Cv�Z蘵`��; H���gr�N�A3�K��<�@��u�� �2w5|s�?��X�-��QUXH+<#������K��� =	��$^�+whI	hk%�RB�	�����K=Zf����i�;-Jm�S=Q�rG��g�0�y���6�ԒN��D�B����(�$"tZ�x��`j��u��1�H}F���p'|�t��zcR܈�zJ�`�TM�)�f'� ���q\�`|XT�s�2�*������h��ԑn݇v<��ʓݧc�6��I�.L��*Bï�>��^ӟ�Z��9�츏s9(�2%~�}��f��ew��Ee���.s��P��(يV�B�'�rj��u�|Ȧ��y��$ �մ�
�h��a�0���N�D������x��i������z}��Y�q���d��HϾ�;��n�9����[U�WZ�D:�A���l��s�c2N/=� ���p�^��,���J�9EK�NGosH����j��˨�7��vK�\��v�RH.N3��_���</6$�2������(?"�R��T�{�#z��˔�c��")�ȏ�%iSZ�ŝA�R����2���9��	�W��ƕ�v:jzy,��Y��=K�h��+���>#.AH��8���"(�Ԛ�A��007�gS9��-v(ke�޹:�Rj�v�s-�>D��n����wI�����;�y�n9:6W�ܵ\�q�}��@ۜgatr՘ h�P���զA�_��-c�� �N�ƍ��Z�67�5p����شnt�����烀�9�a&*tgNt:ͩ���|�V%�xB]MC���Մ��FN���]��-�L�Ɩ�ʛ������}m��	WԟN�/K��WK�3a��P5�����:V�x�����^��+J�<�S{iU�p�Vs�d��n�ي ����r��_��D�i#σ�� �����~~�/�c|h��JL4�8r= e P��-C�;���X���%K����Ai���ؓ8����Fֵ.�S�L�A��Q5��ݱ}������Y+�T�Lbt���^�(���=@)<�r�]����|w =�� �L-��0�b>���ss�L?�%C0�O������v=gܴ����M���@Y^0~��T*)�je�D�#E��@m��К隷N\x�[�'YC�/��܋ETž�A�5��a��,�ܼ��
cO�yg4yb<�W��b�!=��8�dS��{��[u��Hj��ddtFcpq�&k�Uǜ�4%�T�i=
0��w�f?.�s��iTefi�bfRT4]�*�~,���K��(z�QV*+��3m�}9(���ń0N�[���	R�H+]$,�y��ex_�l5{�6lhQ훋�J�u�����[� �;\��O��o�6�ӂh����T�� q.�4xRXEmI�",,�=,q���MU,P�@�_?h�ئ����'������~-�5����($�E�tLˎ�~�����M߿�U��N��x,Xʁ짜*�y����#�hc�+@�Y\�I'��׹�ٜL.��谰N�l����O��#(�,�e~�<��t[���H�H��>]�T������hU�LhM�Z����w��t4s�>CC�<�VґS l���2�ưv��#�4��0W�T�3�� L�R��^o�;�l�P�}=��q,Qqw�k�*�]����vm&`j��#���P!���Y�(CI
�%Qh���5l+VL�T(M����УX��u�L�m�lo�|CC�2�&Ռ��>� >$5F{�n��-��V��)4ط8�U�f�{w���B\4����ͬ!���1�?9�����&az��n����Z��֠��~�H�$��HJ��~�B�����~l�	kZ�fw|VWV��Qe��xb�!�B��`��4Im.e�W�.�:''���?�1V氉O"S���Ƿ����kY3��O!�F�d������M�C���8mn����
76�6�e8�"��^ӘI�d�L�AR^����->�W$�E��G2��ϼ4m�aFWON����}Hz>�%G�d�eK���l���
������>S��2*����V�F
��$ ����_t�ˢ^p}&E����n�����AV<v��:TW����e*��!\Q��?�î�?�ȵ��\��
��z;�{�vڵ��~�Vъ�n/-�쨫�Mv^�AZ���
�em?3c���5��-��$s�2��(�4,�lp$�@Hij���`����g n�!��1My����6�>V��8O�\�h�Wi.`�#��B�
��cJ���$�{`$qz��_+yOV��	����d�..f�	P�OHe �i����������߸���	���1^z�'<^�ϯ3|x�n�1'X�©<w�od����r(l-��t����@�:������ܜ}��(�e�Hs�?�ӭ��^�+�~��V ��$����9��B��ԔkeL}���~�D��C�?�k ���B�^<]��P�����!N����T�rcSC\J����z�M��|@c��a,��O>d�@W�t�߹�j�ʙ-SG����tl��W?R�:�j���3�=1����]��>�;5 �+r���D���|׸����_"�jt��k�4�/��D�����l~C
H��AQ��� �F8@WvLf��4�N?�ͳ��8n�5
�؎�2G�*Wݜ�^�Ʊ���7��z�j��4b^ڼ�:��K��E���v�A�mWh�ι���[%]'��j|D���S-5�v\]It����V�Q�x���>���7C���-����ϵ!��O-f����}����g����,����ݸ��3��M���
���)���їNI�v��[���S��(�;I��jB�AԿ�7�K�v���1S�"�erw�NV�n,n�9��wx�ŋ���j�v�9�F���Ϯ6�1��n��#M�c�L��0���˭Z|�!�]2e@#�0���#v̑Y$�ȼ+���{[[���%���A|1FesI��V�i֢U���X�k�#�<�
<���Z�)�W��|�}bUz�{�s�K͡b�K� T�Q��«�9YMs�������͉;����.-( '`����p-3�mw��WQ�۾1���=���u!�RF�c���UK��0��W�=���+4�a��L'6 O�UXg��Nㅣ�r�52ީQT�_�]q�j�|#[k�>�,=��"a���Dn��7{�OVd"���o�����
���x���:(�y��
�%�V��y�E�������[y��LOh���@R���]D9�_I�> ����¼C-kSj�h$�\�����R¯�S�2��Y�{*<J�<,�F}u�9V��>���j\���l�]TQ��r���A�Sts"`�T������"D�	�mt`*֍�Q�)�;-���5�i7��$(�.�m��$�q���B6��Ch��>����ش�W�,'m-����vm0����gy*�����.�GoD� �9��p��V(�����"��/��Le����O�F��X�WJ#�,#�IQ9���� �jv��*-	.�+��d)��Nx�ⲗ}��|Σ���k��)�g��P0V���=>{������H*����:���s�Ϭ��k2\����B�sF�<�OA���� ��<�g���PW�	�M�����g�ݔ,� :|B�o��	-�Ȋ����ԇl���A[�6S��`Z]=��ë���~�� ��dǸ� �k��(����<#2�N���}���g:#1H��XF���A�^��WE�y��f�S�m�e	����vj�&�#+��!c��R�B@;M����NM��_m�( `U)9�ĖvcYl N�<���v�(�/�O�p\�#��.�d�����zN���x6+�@�#��tc����<�s�-&�.
���
��,pAX*;;_��W�X���u�H�C���7m�zbF.��(��P��0^2v� 7�ꣅ;���N^Û����}�j��Ʈ�n�(�����.!.M%��~�V���Q��aک%�W��[�� ��S�h�c�QC-r�����U�~�6�*�XWW���C��L_0���˺�.���m��5	�|]Zw7nkz'7#%�nD�^����~8%����Y6L���w��q�_e�2U�nפYaړ�_�疳������w�D��H�ET�����JW���L,�u�m����ߪ�����;v4���:ʆ�O��ڕ��O������E��UxȔ����]!�n��t\��nd���xˆF��ʞh��o2������'�Q�^ؒ|W�sً��S��C̛�.�&Ҟ,Ks��E�����$��x���~6S���U��Z�Y�t^D�ǰ��^���s�&=�l�C>��{m>�#^$h�h�>��6;o�;&��a�&�{��9��fP��n,/��v��'Pԝ&�dff�{��a��b��rb���_z,E��@(��A2�f�-ޫ���`�m��'��Xê�T�4)�&�P9�|SzX��|ҡs4I��2��9H싞�kfC�h)!<�>h�ςq�=M�X;�-��%�pۍ�"�K���32V�$:�=#/������Ѱ�~��3��2F]��������Qwd@�W�%Z��|M�z4���<�I�A>���~��#r%��dV�u���._���S�!C,Cq�I�ޖ�X_�O���瘟.�"Nč��`k�O��l��'�]|�%d����f��ט6?�=͹���J�Λ*C~a���'	��A���~�&��v�0�9���q�(͛�ݾ�C=��4��;T+��UIΣ���A%��'��7�y�׵�.a�l��|�*w"g�P�W`���)�h�<6��ek���B��(֧UM~}{;�*�������.�@jZS���f�jo���^�"��KAg!sJ:dk�s�[֚�D�N���s������� ��P�6'A�����7����ٿ���7Aqi�s��ч�HNn�wSJ��Je�|�(<\���_��o:s�&#�d�u�;?�V��Vq9!^H9��44.�oTa�1���ج`�Rȭ���:kپ�4Ƀ���l	?��R�%������o�,+�N���K�@�e�a�� �4�`�4����F�x���sk� @k�.����6��5�`s��s�0K�j�'������<�/���O2���T���T!z`m�R��I6b�`O�����)5�jAq`��\���0� =Eu�\�[9rj� ��1�����X݇���N�GwϨ�H<O���jܫ��F�R���f�d�˥DcAC�/�� I��c��(a��ϑa;�-4���GR��o�#N[����|k����'�e�Աe�T��*%rPM�X�toQ8�h��" �T��:������*�Mp��r5r��@��,�������h�JK�ˇ�v$S�{�n�����	�ĿQ�k�Z�$���@�Sڝ�S��,����yJ[c�o>h��]R�4�!F|�>ί�P�N֨mzؼT��n#�>�c ����>����Cz��S�U6/yi�
󗄛8���mO���)��G>�k�Xoz���9����bPN���lB/��'Z�1�I��	U�C���!�ٻS��HyҦ���Q�E��~��L��1ɒ[#�9�z�Ft�+ d�,6"Oo��M�$��g���E�����-m���m�w.���A����P�,s������aƍt�q����o+��&�c�"݃yE�3��-�H��|�B^�O�����6�	�����]d6�!AA�v�).x����X{ٌTF>U	�&Z�Q�������� dt<�1��o�9
o��t�p��ޱWIm��#��W^�(cp���#��4�'Z�$���Ԟ�;�T	8�ni�9��O�t��֭R(N�I��?#dE��g�ba����1w���ű(f�~N6մx,/��G�v���+��▀[U��� �7z~��7w��;��"6V�S���L���&�X�[#:C�F���&�ظ=D����4�rOD������������Bw����*��!����	�bw/x��$i)�$���D��2��M����9<�8�Ą������{1�6����'dp�3�껶k����y��������0�x�N�����L�k*��5Qsuoh� �Kz�t��qE�z�6 Pqb[Ω�P}�mS�8��faZ���"O���� ����mN���b?��WD-��j��v��`���;S�}�h�)EIH�e-w_��E�-��9��>����#���V�1g��̴N{�3��� \��(�/1���$'�C�
�¬o�T�N���[+�a��s�����"^y.y��y��������1�|?`y��W~V�D���hU?�fT|D��Y�b�E���Cұ�Z��C	�G(�Lb�T	^+�Ǟ�,���;t��L�.��>�?��;���=�
�	�?��'k{p�$�F#Y��7�D�$�Nm̝T�`��+E;~8�YBze��iQ�r8I��)�lk��|��.ݞ�O��>,�1ґ��b��~������Nv��g�F�^�@π��X�������sc��0 �0���vO�E������V+L,�L�������7&��}��T���L�<�k,<cČ�N)�����z	1>�����l����!w\��eХ�HP_��T��ޯ�֥��"�pBi�U��M�E[:}<-*)>S@�{���Q��ꀲ�9�4aߢe�k�_s�L^r&Z��������[��K	3�[TS���{�.�w\ �aV3��FT; �#d��$�	Vm�q0�E��+���ݓ�<��A��.�.�f�㝂����1�U��tB@�.�{z��pR]�E��角Y]�#+7������r/t$K��0���Rq��B���&�^j��îSc��V���h)
@�ׂ��"ĉI�D�5�w}!�}&	��s��1���ښ�sID�����r|��oE�{����o�_[����'%�7�^�HJ[>��[��c�S ����Wb*����+�5y�JT�zC$~s��>Gn@\�)^Lc�]�u3�"�d���װ���
��iR�o������Ͳ�w6��s��*��0>[�B�7�����h��$��[��4�s+��ۖ�&m��ޓqYO��A+����{�]lL�b$o��n���'�S�i|>{5��*6�+._/��/,��W��ŕX 5�\ff]i ��T����̆Bw><��6rzl���$g{TFݦ�sj�����~�`���C�i���[= �.a��I��G�¼"�b/�%�Aѣx�<�t����?���m�ŵ�����tJݫ�@/��Ծ�
������*�wa?�%y�a9/��'�m�����/��}�����B����͸a$�{}EB�unԻ�� tGw���'i���7d�#.W.���9Ja�*""m��x�{*�a
f8=�L� �Jہu��n��9�� ����S�6QJv֭����M�k�H�2�}jg$s>$�w�u�N�ܠ%����W�m�INm����W�}�3���o�q.qn������'nWJ8Y�������a��C=H�������f􄌻Z�7��#����z�}Q,Lp
�-��:*3����]o����FX���卪��`.��I٧����C��ֆ۪@�t��J;U������8(mL�I�G�I��5�A���<��]^K*�a�z���@m!�e;�Ϣ�����,���������Cje���~��W��^]�����k�,'��x���WM=��T�P�l�Gr�
����8VH��W`"4�/�t�We�`3+�+t��s��M��h�S��������
+2�nxu}��d��8m��yV�zy@�og�e�����-ĕ��w�z=���������b߹&=t۫;_�dx!��I��������/�[��/(ۧx�ਂ��X����E����";F7>�6��,�������m�$y��U�����oTi���h/[t����ڞ3�[��d��R�jB�'��ר1녶T��k�i�R*p�e�%9��Vd0���g����[s�.Z�5�f!��r��x.1OB��e��������UkO�kg�Ey(V������bt?*����8;�÷[/UL�I��B��q�y��!YOb��i1����?=VG�fs�X��n�! ��Cw[k�GP-=���p*����n��M�pfh\�}�,K�[I�@��X��+�T�4��>}��-�a��A[��|�|�Լ�G�eQ��k�w�l��>§X����cq�9E����5�=����������阁�M(�a�c��KE�&��/4h�O�5i:.Ќ�B�LHIE-���[~�ϛ@����Ow�5u�������W�9�Td�#v�;����	��z��Mth���}��&���a>��?���<����C`N`���4����U�]Oj��+U��N��c�D]!T��_đ�&���)��Vr�]
W��s�vl�?F�T�𓫶zN���`�)�6�;N)D"@����θ=�P�y�>3���B�d�X��� O��$]lu�X>̨��k,�.���i��+������"1Bm�����cU��e$1�������j�\X!�מ/�/af��S;#r$G�VL�A�����k��e�T�z��C����j���"H�m��,��3O$��@8�|�����#q���=	uA^�$��T�5Y$���|�VG�u���#ߜ��(��y4>�qQ'��B??zM�*e0���������P��R��U7~�az�)a�����4�/,������)������p�:<=K���Ux2il�f��&���A�����]��{�>���a(��㬤���h�~��,����uyw����a�	��lV9ֱB;��D#�F�^�'�(��;�Uu���i��冘���nV,��7����^&L�[@Te{��J%+��>�0��	9���rÃ�;��˧��U��
n�/<��-�����0,�)4c�q8�]%y2��$^"\��n��OGI�}�o6��������&*A8C1=��3�CɛWEQ+(�[2ж[�<I�C�zZ�����3 _����,}� ?�����3���nF�^|\��Z�ɼ�A̀Y���+�VQx�iz_A��N��K���q;v\$}q�"�+��Ď�j�B�l�gLNӶ�5�L��:8	P_��<L�%dG̺j��}U��|X{=�,mu+O�sbn��c���_q��O7�6š둴��ޯ$�].%�C�NGf)
4��J}����%Y��D�����\? ����i�e��˧`"��@f���"B��g���.�j��5�|9��q�x������G��
�RA��7f�A"o�IY��
ME��>��˓�z�5�]�9����uɓ?��B{�A��>�R���/���Z��/l_�����%@�F9���������OwJ��s���M��~�c�*ԳGη���"�Nm�'ֱ�'��'����^>�� cޫڰ,Z�qՀb4��9e�~����B�\�*�2Vq��R�	�����V?}�/P
��PùR�R��"4Cl�V]K	]�i	�-�^�O����t�{n�`5��I�z0�_�yM�ǁ6$�1O3���׬�z�'���pi<z��p0�Myh
m��_?�!=٘eÝT�ԝg\J��Vk%6&����VO]��di�K�*���UT!QN�
���vr�p+U��b�:�9�)Aӻ~C�}��r���?3H��GDϕ�:��r{�c}����Xy�9#�e?��'M9�*��]_����j�����Q�8�~n\K:/��.�+���.���F"-�����_iج`��+�ז@��x��ǩs4ppc��`���s�x��v+�g,ĕ�8��")����B�ԃu�����Gi�I�]�O{,�B��:@�f쳄+{����W�x*�q��\�_���ړ%Cۓ�Lr�'����#Xo"�?���B��'��j gC�cgͤ�n�ZJ�a�P�ǲ�XH<:�q�� X�@'&��o���b/?x�:�%xx��x^�oF_,�����o7wƘQ(E
�zV����pb���?�Ϙ�T
��ꨎ���������A�Иt��?�tJ����%1�a�=_�	��ag��`	���"���R�BLnEٸ{=+����� |Vu��ũOEx���?��/���UwW�I��+6DWS���a�!3v�����J:��H�Ԡ��'�R���vv|B��K��?#q�ƣ���������C ��u�	H��}���ԩ7��B�Ba�2~
��]W�U1��m��=S�ŗ��i��Y�q��__50p��6��u6+9�]���v�a��9e�"K;�3-h>\M�E#����\� ���� z���K��`7���~G6��E7r6.�g�%,/�������)���U-32 �CQ~`�y�EG�`ٜ�T�e��,g����=+���i��hњ�7�Y���!�JKQ�����8k���}UT��Z>`��s&���4��
�(V9˝Mi��4�p�D�t�fld5�,�ô>����o�� ��j��-|�X��7bi������R���{�&|�6�9��^�Ke�!���ܬC���u�M�vo�!����;���.���m�u.��FR�����67=�roTIgQ=,Un}d0濢Ҵ��֮�����`.�A���_|;"�*]��1t�����(�R���-A��xj(��e1Ju�>K]O�
j<n���;�	�������餮]󽶅bCD3���T� ��*��E_�iy5��
��|"N��	��a���\>to��i�;v�y��O��yAJ����uw��*3��i.}�/�|G��~p��U�;0�~ʏ"�K�첤�G��=��4�H��,NXJ@X������k��l��-���ۙ�[����:�[�)�=�U�O*�t�b�]� .%�@�s5ı�r�ً���##^_5(����rc��B�]����ɿeZL�(_�r�L�[@� Z[n��ϩ�3�K�2�֜��qqz�lՇM���
۞���('�2�{@�E�b`�a�����������M�~�����