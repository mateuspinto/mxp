`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mzZ8k8nL+JaWSnVG/FweCs1o0F6XP35bpturASSZPloCTF2FidulL+6pU0TTHOl2IDCzyr2v5lOd
I83c9nBUsijHHMub5Xql8vvipi2XBa9ZARTHAdsi3DniklGGK5neQL28NY6g094hMVZo7ajQHcl2
SOIx8CRPiKPg1bIeYxq2Akx44+l9LAZ7SjvJtTl7NtHVe3AK8u62zX2eDtlif1/zG/JxyBuGPBGW
7sK6Su7xcEmSonfQPFNZcficiq9Gx8J8Vw9/JmUSMQWJttlS9dUH9HpuJZvf8AEzNEiYcpKbzq2w
Nk3dF+bcC9p9ES6uMMg405mHYwXq4DPWRI7Q1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="IVqAS8f8Tx6ChcGRkm+BNPINxhJwlbsnZy5QhLeOHq4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
snLgdAAK7X5qbgg0cWY1d1AwC0M4s+v3qFP3NoIT+aPxJtiVs9It8T+Yu2y6OW6v3Zqd8y8qw1ch
ALFIQy5ZcJ6jC2dfqiOuu1y9QX0dPcl70B4PYqXwAXTOQ02l5dITvDssBNmAZL07VCnGLAIIjQaR
Z/Z8nNMFqYdeXfhH7toMif/JoMroX3CYIX4fhqk6eSHDTs1lpZzLiAlnoP788LKaqr6YLryRzTKC
EAbKRaWG/kUXisaTB45DqhPqdFV2BKS1RzABvZWfpviMKH/HPib8ibSWQGybNyma1tBrTVLP2cOz
xYP6i9IHEKb/fnVkdhDGQjM/1es1aTMEEITCQRQtSuYE3sgMIkdekAaNw1cFNXy/DH28NuTbh9Ev
tGx7Y5sLPiTkN3Y6sOBwJ1cYR5V3HUdp9G71ZEdiyv4641OiWnaT+hCPKVjkgMl/e1D7uZgWleVh
aDW0n7pK501WPFWQvv9j56K+zWpkxAXaQfAXy4LbYM4sBO7FGGVTs/1oC/8LeKqLj57r9pO7iBZD
LpJ6SNAVsx5Fn3h7ka0xurr1ebODDzeio5ZYTt1fsYb2OcPWylWGSeOR05IYGfkem4L69/C/F/O9
ru2mZ8G+BKa385cbk+aiiQIifR8n/ZAX78TNA17qXkoRp1uyRQ7Ocw3vmnG9Quk8cpHd8ZvSieBy
NZCbnP9Nc+rmK1qiWHGpFrlZUzHPdp6T/eQPCs11m9TxwOiFWOW2lFuDST6VW+JKUDfxy4aVD+Gx
Q00ctB9DBEl8pUb3qWt298KdAli8ZS9UoKH5z4s2j6NL0AAJR4ANLVGm5aEqWI8b3Ooee/ndn+XJ
u1jiqz10G6CR16iueKy7wc2m3R3J/gCS5LiNjRa8H5YpXdjmkO7THO4K1iI5sanJ1EOqkvQkiasd
xDax8X4ntGrDv69E+An+UPMcLbF1KFeVDZGb5nJLVPk6v6nBbIpNPEXmjwpVMaGH72yh4GsL9hFW
wzlm2nnlJDDjp9nPir97OgjK/yVQQ8WkFYS1sMtfBEiMM2WONcnJT2lhXSnbm7UnCGnkL5D5P9fh
u2/+SFbzaek0K/mcnklVki2ae/0DIJOa9PGxvqOyKlMWDFwc15lx1w9srLDhf71TE9OAbcZLv8zI
5sOL/IvxO+xJ2CE7Vfw39FPjXf++LL77HNazFq4kS/yWktoiu3psg1kTNzR3JdM/XS2DIVxqx2UT
rYrdJiDbRVIP/InKw9nUpFm8jigB9Gw3FfM1mKd5H42yTVDQBvmewwE30U5Gg8Dl60RWYS1KyjsU
W7SlJj15MjQWNLY66WVk2oc5AfYzS+WVPMlMC9YnMap0yW5/rC0FfuSZZJzV+bRn/rGlceKWDJXh
c8S5d7+/nBwAtpTaoUZwhN0IOdtcR5x2NOYDGLM2cggYoYlMaj+o+EOBK2Gfgp6tUlUPpKl6+Ss6
bKwAruMnVyIKVeVUeb7QY3S50XgSGnFBXweanIrN9x71K15BqTA+xOR6BJ6q/PL1Bs1qDvjdAB1s
cXx9dYgLqG/foVdApUXREuxQ8XUdw+o29k+siCSkhClvfOif17M9J7W9PoVqKMujADDEKgmVFhCt
fbKYS5Gxibnr/vo21WOR0UuYYo9jm0FQJyahoGEPIru7GnbOtBsM7vJuVhSzRcMssmrxPKIaZYXv
ulnenREYRRx38TVML0ianzsDaBWoIzxTMNn/Y+lyVtJkXfU/uS6kOeTiXQaTQQ1dBYIGp6d6DH/3
INDqvE4E0Ulm8yr9pWxq0bzaPninEFJeoL0c0P2ivy5GI7ILeq9081Tj9xDv158Ugs+9hayRjK/V
TpUOIwgdShsky9B/1GBr0VZ+tNCEmiMomMt84CF/jAUdqw6hdcNTCahyi3sRaX9JEiG2pxNAPxUI
RACZmrR/E21itqoFRwuI8yIz40EckY2Qzjj+PPkNCVcQV0RudKfgHnvxrHzxKfaUSJAEXrDXEBA1
sqHSWzMBVG6W+rHzjMjIcOXZQ/UNtPUEOps/z4Z+8T9ZA1t88xt8bI4nnPgLxqxpqH+zpweSj/5u
+El49vTH6oD+b+KLgoRUQxc+c7ZdW3WZiBjcSGQNTRpH7fI9mAS6c3XlcVlbOHGcdvAGJRlENRLf
z/0pcOBRgO/BVV4h9WmXmhLho/5yZC4ItURB7jOISqMFQ95Mf6hS1th3nXvyDB6497udTXUMidAe
de5cXdpNTvimCPeHuAKh2TkqgPmBlK9Mx/TEm4cCI01fhBjQZyWXqZ8YGEeBwSGXz3ry9pXmN1Zr
OL+sCVxW0JHZ3mMXbwIPZhIYH90LdfJmQXV4I9bNOUEhDwPxnJfwV3KiSi5VPkJKg9IjTLLpNC9i
1jSmw+r70EHmX6V/t1yNh1FafN+OEOZ72Oi9lkSFnPM82sJ4yl4ozRDqyC/xCP/oqox8G4ZL7Mwj
qYBmgZTLP9hPZJg1QElotrTTFh+QlyR6hyqB9E9RBuMvupqWwJ/s9MdFaylLj1uGdPCh8/OhyveZ
hEMBcr/DvoOi7Xgs4u9Jp1kdzh9QCR7SsO3ZTKYBIicu9uWvBKEYZdoWhUJdn5kumdKBbkfhdtap
CXQFTicYE/Q4A6mvEbRj9VWOJz8TVGGz7HTiTyXjXm+/XpvKVQFdvWgCFd9KsfUh9bfdbbWEPjM6
ROq5T4mqdMr1+Wo+giowSmJy1jRh1bLv1jpcKpJqlR0m7xivuaTormJdxEe8VYCoxa3yxydGrAKI
4JRpl5+TXWsFoM9JG0to5klHx+buZNhhQJjkUliUjwWoSMug2tnSx3J/s/KyelHOgjo1QnkT+XKM
bsLXtvt3sRubrYuuZ0e79V+daVNcu9pnpj7A3GFz27xNRdxkflFyBLXlvubFQNFEacJOoAwQ7RR/
R9ytNORXNO/K37xCgOoQS4RqjfLUXAZ8UO2+7DaVF0xlWkEFK52r0M8rq/8VQai3NMTWp6IVMmpK
Ir89rEeGPNpRCr8cPZaO3tSjEe7bb31pMEXEBGsu5KwXOnxAL5qE971YjV/q6FdZLU8fwGONstv8
iTf6eVf6+nBQ/ZYuDtmaNavAL4m1FvyuARETJmGm0Mon04d4sJ/2yB4+t5xI2gSXwf+W2SiUkb3z
ONTCQ6piYAB2LAveLyksffr0b+81KQF3zixBTapq963PrMZyDUy/6CO7dB+wSfyxqgR3h4Zp+WP3
O/lmKIu3lb+MZk4HraXHlU5/8pMKMoHTDP2P0Ql0XZ7vY0Rv6WSxXVhUg7LLT7pPAxz+GCjaScc/
I8/aNzsAZ/ArKy5HbBsFcUSeTqdjRffcBkLrhINTcJvVd67fVEO9gNbLEpw9Qxq/u3t8ATO2wFmW
3/7XJoyHbLTKQ10Ywa8BfyGtexO/pXGAPiHepe7dskF5w6G2GvNK7dj94ouMH07wdvVqpy68HiEs
Svq3hnYCwnTxkZXbvKtSlXHgqQIpQncVfLlEpRB9KM97dxCWs5ryWV2zuUHxwDdwdWo6i9fO4WFK
Vw1TdZ8FM2JnYCyJ/7+m7HncCnmfmmeirxJTs6syL7Q8eFDEpQQ5ybcwl5aUEMawy6p0pCuMaCKr
DtVGY31Ebv9XHmGjppYLGxOPZKKfnuzstsTkw2DYQxniky8MijF6UuB5NhOpjd//5yEjUoHqPQRG
WRTxAqtFVcvjwXKdOj/hz7z0aGMCQIJ/dSHC51Uged1RDkYlmaqjsN46ZE5bw9f0bBHgns6Ysaq2
P6zrW8JeaSJnObuieLJp7EOmRsmUcNJbaF1c5MjxUiX9HjgStegMKchFsI1fp9DApQtc8EtrWV3L
l827p2cCkP3D6TdY1iYe0A5a7oAeh+b/TgMyxgFt2R1A46pt/sHJ1GWJTJvEr01Q5mQIqqHFnkjU
9jlAQx7bCBmOXdPOxz2A+x+Ueb4aYWsUv11nBOQWbNRv+1fBc+N8anYAkgs/mKjxMDcpuaF2dLW4
flKH02Xawh7cU1REY1ZCqKa9/sGnX30xIjGGs/ykrvAr26nJtmh4hSoX+4q+rGW+I/6POXRMW1PL
fbU9tyLPXtERggEFuTn+2zV3a8epr2PUyeVQxw2NwmJi25LKau6b8UouOsLW1FShM4mUUuH9sopv
+mTAoIvEvLPmETWJg0fbFJax7Fv4Rddyr6h1mIkW0tGhS6OATYtLDHLV7ykhKrmKxvzTL6TGwaqQ
991JzhlHckMTVHWWjtP3DJhqXOS63ALVbRR8yTZiiXEm4i2r4epBg5elzhXE+EZfx16yVkRiToss
GQgRM6JBTSFnC3yXrrTcv/6pxK5h6IdK5q2q4DjSNih8GM21aq9+rFYnLSHXcOIrhw3v3SyypfVT
0PGK/Fa11TlAq5zB2a6JRffOiNhV82ZwSbp2Xlshe+OtpwWrvO6E0elk6GNVoXzZ+sg2B6Ij1Bvh
l0exrBP9zBo5OBYVNxS/QVjyaqdN8CgbPKi3rsIiPfn9Vxc9bOb1DFoUX3PylAX42elbiB42Cv6O
9mkwy1nRDxWidpiznvNPT1xkQKBGysJPWw4gL4QBxV4cWH4Rw+6dj3W2kY/zlBu2GhpwjiPxlk7s
IcLF0zdxGPsli3aBHRslMmumFTuc8+eXSHE4YdeGEfCw9UHdxIitLpE43ePTr65k+FEausknZq4V
gSixpb3+RLQcw8knP+lwg6IRHN6IUl4NZ3hO
`protect end_protected
