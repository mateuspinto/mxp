XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���uݧ��f��Z��Y�j�M4�ιBz��(�面�z	���؋�)��A�_M��}�sڠM��kc;�.h�g2d�Z-����$� $�됝�Z�>��v��Uzʎ�XK�\��-�7JQq[Z�<�p������b���,N���(
w�.�����נ�)�1�0�@�ѕQT��+о�'v�TUC��LȤ��T���XؽVrN��4m���P4:%g����߃���nyJp�H�c3,)���aH�O���K}�
��r(�ᦉ\�w�L{eH0���Am�EOۊ��8"	�#�������tc�#]��0������Ro���)S6m�4
�(�߱`�����K{VB�p#�+��M1�?{���봧���2J�p��΀ _���Ƽ��hhYᙲ���|��Ս��~��8!|u�w& ��SB׫7Z��I����~$��$�K!�P���f�����-��)�c��<�z6�4c1�a��K��Rx�l�\d���^��ڑ�2E����7f
5��g�+�9޺�m�f�NZ�vn��)�k���'2a��^�<��C�<䛏�e��6�s�CV�����Ӧ�S�̾�v��0��>�F�^
�f��oAtđ��T,��!�c B2�p����ӫ�Ǌ���6�}�r�ݎV���5fb+.tDAp�������ȍ���RDa��{I�%$[ݶF��}(H�^7���P5���/�df��I?;�c��[�òn�����ŪL��Q���lXlxVHYEB     400     190�"����O]|�L��k�P#d���쫷�ĺ"��
M>$���ʙ��{�H���g���p�'ׇ�SCoCd��N��hh� !�r7C\�!�}��1j�2L���R�\��w��c��^Y)6�l$��h�j��S��j5���s��� n")�}�\VS=�Msh��ފ�Nɵ�l*QV���ڦt2K�:Vvx'H��xqM��N��8^,�G��@�U3�e���Y���fP���<��� ��A�1�vĐ����w�ů$�|1�!�'�x��ݨ���3����X33�W�3��!8�.�TY"15���9�&����HM��*ׁ�s��rX���m�U�8�Tba��i���Q兺A�J<zh��i�|�ۨp%^ɯ��'XlxVHYEB     400     170�� A�pT�R�sR7?.A'�ӗ�~�^���y6���~����'	�ŭ�%?���%�����ə�Ͽ���C!�]�HS.�]����%��w�e��/V{w�豍U�����2���(=;_�����D|,��+q�Ȃi'ٌ��6)�K�yӹ�6�Kt���U�j�\c���J9lV(T��k[J��Ĺ��#�s�B��8�6d�� B;D�� ���<���%z'��x@�~cDCoǳc�_�G[���bz��=���<pX=6q>�s�Q�]�B,�ң yf���8IEM����05]I�&%)K,��5�����S�~�쯄7r��?c^.l��Ԑ�&�e����b�z�bd[]7�Ն�f� XlxVHYEB     400     180�Bn��s$�糝�Vj��/����3M��=��0��hEN[3^<��좤آ���O��[�ip�:&����|bIN�B���i~����\m�8��4m\�����%p���w�آ1Y���m�i�0�{�D
�����up�/I�6b�JۥG߶ɖ�V�|��Fw�1Eu�-ɥ&FoC��-�H�0��f�3;�[�&�ip����:un�>i]��������@�]��F��R`y���ؐYQvJ�+����2�n|ZE����	EΙjkk�u<D_]�Z͕Oe��r�T�"t�`J7������Xыe�襣/�J vl�s�K���F��t�͕a�<��+>Z��JV�����&�5S�Y�i��BT��XlxVHYEB     400     150B�מ�gN�B����5���JM��~�:4"�J�F턃$/|9��~�:�'����1��)|��������DO����%>��4,���O� ��x؂�|���Ɋ��(��"��ǟ�B6z  ���ڤf�Ki4�"��dl��S
��"�lQ[_�����ҟ���~�j�'�ۊ:�.Nl�,u7��4׏���ʁP�kO$W�M~�*��	e�l\ 7=����,|����fIM&�2Q���;�Zs �_g�%U#w�l�5�w�*.���۷����>���שJq��|�q��U��	k��V�=�7��D�l���_�i3<ixfG����j=qXlxVHYEB     400     170+*>�S{i�z�Q��g�����$��YB���Ԯo��<��8fZK:�K 7�µ�J�p������T������H�`�r���r`V�cB��aǸuW.������w>+g����Z�7큦�0�C����_O{YjX:It�cSޞ��#+yj�������vHZi Sm�ө�Do�ޜ2���q5��g�9�-�5�e��o�؍�&��������6fI�/ ����Hg�췥WK��>^����}�mir��	S{��y��Y�2�3�
r��@����-�E?�Y&o����3�Y)�?bIף���`9[Ş C���"����\b���SW�褗^`Uʇs�l-��(-��w3������}�XlxVHYEB     400     1b0]]�O��ߨ튳�uD�{�!��0��!��o(7�F����J���3~T^\0ٛ��>�e�-̳F�	���,<UP/*�����Ez@5��v��/a@ &�9|��[r
]�d�n�!<��^�f�d����|3�� U4��B��il��e,��d�7ܭ�&��[�N���uF�W���v6JCf'J^�IRV�I[3��� 8��H:"��gm�g6x��h�lrG����P΂��T
�A蜮�ۗ]����Kb8S��	 S�^]�ٮ!�q���ٹ����9҆�y;Rmuyo����H �<��b���[r:�Z[�eCO
j�����5����#Z���xh���Ѣz� 0��#9��C��8V!�V��~�e�=�r�y��sR[�] ��������R"9#}�$�L�ȵGy���ٽ�˫���XlxVHYEB      e0      a0��X�7�BZk8C�%��nŪ���)]�����Ϗ`�:	�X�Y�1�s�J�A�@>���3f%|��1D"�ڰ���
:r�O4��Y�X`�-m�ؕ����4i�pܻ�W!��� ����\���m�#Ե�< 8��2tn�P���Yu�$Sd