XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~8��HH��keOȘ�Z�)���Ny��P���" �J������\?�h�)��4���׊����ys��3��8�����5c,� ��C������6K�c����˼(ǔĐ�!|����2�_I�⯻([����1C�_P��������*E��F��R��_D�8}|�ԣ[А������ "�QRx1�j������K���2�<ի�n�#��T5?�EV��o�{=2��ԓ�Os�g�7@�����G���V��[�[8�o��hÉVD���p8��E9�ӓ�������F���.Ǽ)p�>bS�#����o�PL�d���P�ӥ>��տD��bR����9�^��ط6�-L/)8qZ���zs�z+��~�a'��X���^룺�}Ϯ�#oߔ/�eFkSЀ����s>䮞ԕ�Px�	ˆ�=��U��_53�d�j;rH�u�5����O0�4<u٫w,\:��I�j3������	7�����S˕�E�/��U#��
B��j��j�.!��B��H^�&1O
o˽�hF���=_����������u��h9���^����'�2����w�Y\m��IM)�B���ɥaG��{�!0���n�٪��$�� ��o��V��NqÂy�`�m�IϪ���ȯ���a��⎚0��e�Jmj��^�����}U�>��bBӗ����	�<�SZ�2�Ob�C'U֌���XlxVHYEB     400     1a0;�>����Ҽ��	eP)����%P�5[g`c�h�}�H�3�4i��n����ޣe~��I��-_1�:I��#v&Ē��Q�:
c�Nz�pp�a�b�0��?��[�\��9$�u��1���xa�SK����f��I�p�ta��Ay���co�2�G�>}\�g#B@�+;�]Z������[/�LW��[Kb�n ���cm��~![���G��d�cy��8�����.y$��p�W�"�~�'�e ���߭a�?��:����<~�ւw/�Ғ(���T!��cƛ�b�.� ��Cʦ!��B$
�=�ƊN�i����`J؃��y����J>�T��k,�:�$,������7�%�>�3�&�|���);�uN�(�8;S��oJ�&���1h^c�}Hۑ�	�W��4��gQ	XlxVHYEB     400     150�*��u��O�爲��c��/xڸ
uM9�S&��ƒk����
�'Q��1=G�~����vP�ƽإ��j`�ȟ�$a=�EA��)<���,�
����N� h�C����X����jb��|b~ �;��*O"L?�rb��t��U�ǎ������!|�I��N�V�s�� � p�~T�sF@+�ܺ�6n�B6[�z�������|��@�<d����eF���iB�@�$�T�!���
M����5�i-�I�c J#"�Į*�J��\&�ʴ�*��彿2i2�m���*ώ�Og?2j���1������+WW?c�*@�U�XlxVHYEB     400     190���s͎�H��Z[VgR���C��]���)ψ�0 �Mļ
���j���&�A�љH�h�]��h� D��u�wG����
�&��D�) J���L���I
��WZ^&�ۉ=��@3��k�pB���TG��3TH�.j;Uѯ$J�'�z@�b0'ό�Ǵڼi��b�\q[(�&0�vd�PG(��)�|0f"޿I�
���8���O����4 Z���L�g"�����>�G��EJ�ǎA��Z��%����e�C~�7�a�Q*8�i�O;`_ǡ!����K�/��%��^}Ww�O��܉u4+��M���k�C�er=9g��gF���'}x���\�8�Ҙ��\��o�����W���~��\���!5ϰE!=�@}آ�C �5XlxVHYEB     400      f0#߽g�����n���%����|\��\4�b=���"�fG��D������Š:\��9����U����.���/�����n	��Y�A,aA��&�<��@������bS2�,h��)�N���F��%�Ր�(�$\w���<!�Tċũ��A[�����]|HbR�Ƙ\`M�s��>U�E��K� ���<m�����u��Y��+m�u�����G+�Ӹ�]���>�-�9_ȉ�XlxVHYEB     400     120�h��aZa;}~��C� ���%Mr<����;-�w44(%����1J�E����q��A��cJY��W�\~�h�V�W����ǐ����PFq����r�M಄�g*U���`����[�������y<*��f���&s��4Hgd�����+�dX��l0	��:�]'��!��0�s���W{c����.A�P�O����ʜ������O\{������ff<���@���D�=�Ɠ쑓�n�o>��G�!�P�ܰ�:I*M�z?]�nJѝ�C�2�L��=����kXlxVHYEB     400     150 9��'Մ8{��=ۜ��-�"
�F��w��{�Z���9:Zj�O��~�a u
P���� 
�������4�V�q5����U�( Ǣ�?�(E��A���(��ܿmM����A[����/M�f�W'L�����(5����՚K�$fʜ��0��|�����-�J;O̽q�:j�"],�����$L�da�U�A�">�u�{�5d�90b�$4	i��kƅ̓4�v�_|�S��v�R���;+'7w��lyg�R��%��s��g���|=$� �X8I6!���BKWlM�9\`��ǲ�q�h.ax�����˵�K�� �"XlxVHYEB      ee      70�p�
��!�@�EnSԭ�A��0��'��g$օ!�rn��=Ҹ�g2�2QA5���Wh0�1���)#��%O�*�[�*e�FV�l�c$�S��!ɖ}C�yI�QBj���̲�