`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
0USWSUGxovGsyBJteYpEoS1AWp7D8zxzJALrqplD4apCASPCvvkAPhyD5Qr4k+0UdSb9pPVE8Utz
aVps8i2EYIY4gRjDZVkBg2i+GDTl4V1ej9OkAVkuH2XCLUOD5j8uFpzBRP+/lRFM3iCz4BkNhvVO
5ODN4HY4BNxc/3+oMH8rVT7cGCrCoNoJkui/eU8oGq5AwQXXOzj37u37GtVzUEY2f2MqrDhjrrz5
kp8hMD89nC443vRKUSmRpIVuckm0v4ClTxJASI2jv6x/H7XrM78UKorzFQBhCLaCJ/hQ3M2Ic+0U
sKUkiuAJUbrUbH+ieogXCQkCzIFmmSQeECGoon2UzsqfS0jsi3sIkJyBygM3ayzyhr76IMBSXkts
XtVT184e5rPrTBMQgOr6HMLiwYlG55ZTpKp4IhvkKgVs5b3JqAl/+2SWS2Y/olaZrCwoIOmCpVSZ
v9KM1HkF9102aVh2JZLMBd+yjTrWuu9KNDm1q6biLO4la+R9vpwlbSQSIqIwo5kkUz/VXtxdiyqI
ELoxekbgKSZlDRzESZCYvJIhiJEYD6ulX0wEsBYf0z/4sIxnq4m+1ZHca7EotA629HquAeO65ADp
18xdQeDgFCYu0edZqFXES8L6MFd67A01diPwwGF5A6DJo+f/n3BKwcwInQemwCI4kyrbPXai6ZmU
E9637QB0ly/KCJg1iLWmvCTlTLQT4kD6miG20ovHhS5s/snkWVGhsz25OdlqvUzEBHVnDDAdC1gM
J3fZhLXe0etUbz1RcrqDRovhBdxM34kgkuCBwb3kJ7PGaIEcFBc39gStZ2S7cqbJeJR4m+eBU1z4
eyTMUY7Ap4o7PYsJzWiMT3ozPXwA07wFob/sKWjtPvMYP16amfsuS8SLZSZBmPJc8tiqoP5CYR7e
Fo+inDgYFGMoHwoAvxT2RCSUja0u1RvrIafMznafEGHyGRSdpxpn3vl4aUuKk9i+qOx0KyrBgFOk
P1eTSabC8t8z3i+uqc/GuCWcKBErUcx/KyfLTCPjoOSeRCbEMBROQB3fIUftqTlK+PRVn9ifpZeq
S9cLvH2Gi0fu55hycnwEdkuROAZnrRcYUCu978awH0uPVuYY8C78B0BI7KzIujrYo3XM2J3nQ8Ui
/WMlmWJ9PovPAgHdMZQEoBUXF3XO72eIsB469HjTKkkUbDVY8iFDmajrObsuqnRHpiMvCZW+VrTM
hbhvoN6l1EurwXGS9eTaqsPACQB6yPuvLs4K8lwXFw687bwbsPwvNhVg6NNlXJxOJ9mh7cF0tnpO
jhj5mgAXXC3d13jcbp7+dvvjDl84Tay3yaQxlrL8UZNr9RKZjKkhSXtSIPUkQ1+QAnVCN0+AoSXa
zTzxucqNbcfD+mNbosm3M4TWs9Qb7b713hYA9l6+YH4iGIJUhX3kttucCF2m0uyjeeWWA7KfjkfI
2EbmLsjdEJacmcgwtf78Xca7HRqeTNXa9nQzu76MQsO7ZIWpdSefHnz2HXl0zmoEsViOlvFpTofE
l25Kz3A+13tKWrqTKmfY+HNUEkhSJdFMBEonicHp7lz/iQr39/f/ptmel3GQF5B+jYp201sypSYG
dNfzeFIQaYuoF89frdO456jBCfHDcbSIl5fA5kN15PtXo/8zUqAOGHtUczz4Uxf+iCenapC3K6OI
plFYkhRJHFZZ4NR0vQdAXgTSCsQj/wqklCSBzCpYka3i3CBYSEeWZe1NvekWIrDpmJTdGU9iLTOG
grhKEHx5UgfHR74sXn/7qedfWYGOFg8Rv5Gjvkz6zKh77V49tC31DoifXShaIoeqWz9quf0uMIJ+
EEE29GNs3i98NvAWOGqr//fIBsfr+wW2SKV5vbzCxbpFb9H8IOI3sS4cV+fEWjWOiQiGFwkAlz9s
VuOKt2+Ul5oMo7NumFidWKaAx9eS/DaCEMI+yod3wK27Wk3jCWbBH7HMEbZF1+DysZsPmidlZJm1
C4w2NbWwiXAOAnbemPEvJ4ObP2ps3e0wtA0rcQIqtzM5mU/IxAHdVrlIsmO2+dZpWAxyavHETeSa
WO7oY2SGQz7NVgSehNP1udTKsbs4Jlz0ypgjcyE4mif59Vv+yf6mn9vmWMwnA7SC9a12Cmyb5esa
vphs9fhAU06wWlrn+bDCpkomSaptRVNoO9/OSVIJKiua6OOkx4umJOx3TUa31q2WFRYQ3yds/qIB
BPH1GkXnNq+lyDphsxMrZGsBn2MIpViHtkJPjmew5VK1cCmLMX5VpSeAIp9ARRatZRcmGhCwXqs8
L20KE2Q9xDeWfvx7JyLKY3gEr7AbeGtoDRF8/Z8bce4i2WNpogpOmbkYaPlrQqRMjvg05ctdTJhy
EWg30fyw4C/uXJqdKP2H3k9ALeYsXkWbYSGT/LRdfsyPHpwG1Gd/ePXgc16Es/AoJKGxI4buF72K
ij9Ew5DvC9WjbBIR/L5Xg69aRzpzNWYASSm1//guHn2scu6PsZwr44U6avTHe8YU5NkRz9x8RAQK
L01NKDLDBZsG1i18DyPu/dd6dGaI1rI/UsXpW7f7Ps5Jhe61GvRxDD6nLb19FlPeNnUOMbiF3qOp
+Z10ZNIWaaCBHyjIwvzNO5/5WG8/lmRujrxmsq65Dy7jpFgiDZRJySdopG1ujOtM+wyIr5Iv/oAI
5sBGwHFU0ZLpN+qRHTv2WUt56moP2p+YxMUJKbr/RV4oc0MRQ0EWOaXtNlO9yuC3M1e7L3mzIMAO
K61LV48OmM6guiCprnaGH4TYS9kdD1lN2vT9Y1jP2Rzar8QpkDSNN3Nq0iaazGi6rf3LkbN9JX/W
GA/NnZI4z2uATi11aanYl7VfTHo4ePfrnmRhqmvSnDK8X+iAdiWvzSrSRDw5h6qh7AaiwEu87+dm
HQXph42/utG0JxPzS4U1ElglhuAOWhOk7lQYgCnjpVmhlueM5UPKrWmxn/6SkeRLF/ZfIl1sGfiS
DXPWXgO4ouuvyzUs3VcRf+2vfto9+7R3fD11Ba56T4al3hKKSdNZXyDuciBKxe3aWxuCOYmH/D+z
sRC9x4FmWeKqYbLBox852cP3mPG9bDwyEON+LEZMCzMeVZGBnhJ5+fGkrwwaqc3SXstN/4XBqxcw
7/S0WSXEn1Oi1VGvvIF2+7E8oA0+15v13P8Ym9W/wMilXTPgafJIQHM+J7D8KG+hVa35V+OaWO1b
IbfFBfrRGQUBF7g+5GuwIj1BhFoOKfJtaYRnnXVtwJqMAMsVqULTMsv2iXGOAOGpJW92jk1Vx37i
CFKvO5FbwPTHj1LbnmJSWboxzoUoo65jVACGdhtN4WUgc483xcPAcXiYorWe+/0jc6ROx70o657S
qywNT31yKlKYDDWCfeu80IFiemAqW24Na9GMXzWoDimvr0staUMdHI70hN0NGOOvYRHLPqkv75mX
jZlUMzXRl+RsmS1mpuncHaiEStfAl6iOwY2LJoaLT7aESoI1lvIhJAxmJGdazUhDPz47udznxIyS
THTee7fwQdDRfwAxClalZ9+rXpty9t6cQlPNqlZvsWmiZbmIW9CPrA0nueFcbzgU+jjVcl8qWpl1
939tUS2PJAsBYb3kbLuhtY9VI03/GVI9aipFHK+lymu5NQ9z8uPRUD4vw60YWU/p07DK3ls7HFT6
omQA9dLG7nbHA4k/6VSjgqJt3NNL+P5VgUWyht3xRs5Df8Ez4i/9D0/CBL9YIXr/OAfSxuXHoGE7
ANjF3BdTM6WDAeT/6MTn39JfZ2m6agdxLrBIg6YhdtXEjLGmb1ERrh8k6Olc8Zld4CD2PkFENkXp
ulcBkSCwrf/OHOyPIZnW2hVDKa9kMkG7fxF6qsloXQ32x9365C7FR44ztC2p9c+HliTS08xW/0wF
7EYOvpZXq3s2bB12b4qLSo9rzYjcKIaSviQ1qtEsm29wlqNsoRKJLbErVGpFngwpcyVFCIS5F5mt
zHAvLykWPFK+7nbo8ray+yyLiXG2yeZ8/FAmDo8o4UozSzVpIj2Sgw/6l/11uq0YKeBlMPM/mxQs
wb6QxD8qzm2jI+KJfji+6gwqnOiLxA6g9X/b0K46NlGM8dU2kvovV8bBRGhBxetpV6NazEp34WTV
2ZNdp6eii+K1L80j6h+NascnRwK/hz1cNr1YMVRlMZRJwZk8p0V1NsAf0c3n/nueuRMvGyXqQdJT
XOWrv4e7j3+jey0dsx4oVcv1Am4V9F5nhK5azTSs+0e8PcofyWlOu+EjfiZtk9ls9US/vgL9gbnA
aUY19KJWXjIkNoG/fB+18QnVrJmzYJmsnSXoYe+tmKWCbkC0mNgCGkxwQecxMYx9DQWrvyDmhJzQ
UBz3HqNAN5g35HnY+0gh4aH07ot8yM546+Yu06jqy6jomZQlwTRS1k64u7XSMivQCELX2+pkrOjC
ypzle6VzgVY83TB5Z2Gpua6roqDJQq2jM0oYoF7xD9XF3oYGQ6HOJXOG0aCWZ5iq1DKmzTbWCydk
iW4N61FbKTak6SxSxDYjkfunBn5D6ORFggSwEgGmfb01fOimGfXrwxhejBwQb3RztKyBuXp6md2A
TA4VLies7r2dV8vB/p2gDCV73LS9fdmxXfYVw8tQWyUZ5zsWZWLemARxoqKgB2JxVr/oQHtMsEkn
sYIK+iVsJlPlI0HQydM+qQGGDBNFEyUn6lu4ldyirTQLy5/7+W5mDYNbq509MG2rTHEi3DjRec53
3l3Q3rkzleC7SWf08o2b5MBZLE/ZvLcuwC+3oV2M/9dfzrChzTcawmfS90Gv04JiTjmNJsWnvqd6
mQQBjmvK5JXE3Gd7W/9imDcv6B8B1HvVSRnlwhO0REMOfcfugGc6womcz+CjcERm/1BdaY8N9N2g
ZL1K6FHJhGB4r1m2ETGmNmNgi1wIFcuYNG8lqS3yGJyBvxiWgA7SudJgitLDF5LqZxYPctrt0ma+
mgQOYdUfs7CjCUe8RDqM/rw6taIlxW3Z+9cmmT5Jgc7Ow1XD4FVkZHON02e1xBomYogHw0fU0qvE
1CvqHXzGywART+6EDD2FDapME83BEakx79xRQe1dt8Kjy7e8yVzgMJir/ZglPBXE9lRj44Ab675t
FNpn//bDDbSoYvMkp7PIhw4ubIvCEJto7DFiclp2z1ReivWbNmbwumcPkD8WQ2b7FyF7kKfhvA+f
SnZ9NBRexa/qX2Asc6VE1DE0QrRk/zyXpxeHY6PfNKyTBQ89dD+oYbnhlDSY3xVUzSf3ev+swUqT
UtdWMzz7taLTl/GvxU+09aKuYAKtnxPL+R5EFpPnvbZH24A4/yEBOPCMdI6MiCqinMWa+n6gDjcq
mUC1jPHluKYQ1i1fTGYylYVeZnqkRqVt2IP6taKY3o4mkdnCz7EpP0bVEde+Q8WUZddfDpxtF6mw
OYH2+Y/jxS5NOBqPxnxNfreJobWSWEp7BeuHz6dctvrcZoSfqJkQ9iuR2526+lvXYrlKQbl4aJCX
0nVNO/CHH7He3mBz1Fr9P0aid+8ItaK0OUfVRDCldU1hUryaSlSSUHxAreHknASmghmeF3Mia1mT
DdVA/oK6L8dwTQeogPThtLJYIE4QS09rfesS5RJ/9cdqTbGCSJBTuHQ2pOWeBwxwDNe+xkvGLOrV
VQ7Jqnk6zpvm6oLHkXCuByVz4HZ+kMpvbNspcgTD7Yqng/qpOdsI4/yI3zIDnOe0ZM1TtzTcUYz0
BDJ92gGts9OeQuVbpn27/B0O+RJOWnKlQD840Ys8gBkBADSYMfNveiNjTykXo6QagXcgaOwcsn3w
203cQl1lyX86aAW3QMJpqtNzVd0xzpqEmkbOZKsTmXHVKeqDD8sQXN3YzS2FRce/sZbEPx5x1evo
uwF5ToxT4fux5B15mw9VxpEsU4IqBI2D07H4HhcL8ZrvKa+P4RoGdXFfSq7iIxcGm7q2vleJqjM2
YioFuvbMEGv2qj5A2kRJyv1pafBBI3oYGfYwFW9OqaDdIjTP55mZMyBu0wsFW0YhSIWavj1GH+0e
6pzrNcYt8yEX/NlX9letr2LZ/d80LYA/9ilM38oKThzIHJfAcHRs3SQvUUaTDo/uINZ7xs184JWy
VF8Lgk12ysfaOBzsKCKQXAXHLqP8VQhbDh4uKau4QVtqPJxXHImRZPs0O0egZQ2wcY/t5H+PXDuf
JKlOi5ESd3kv8V/gsdfdk4Dy6ePHixiZ6ptf6bBDf7cjEmboxUdPgsq88JOLinJN0MA7mNI/OjTF
n77ptgU2fgF1nCUl+bGHMGJkbbKtd6b6/2rVMAfnR6q9yfLF5+wmh0zAWeUGioTpJ2KG3UTMyD1H
sbu7j3rp8AlykOfxSdOvHSyVo16aPGAqwryGDQczNvsXPKc7ToQ7atF0vphKgSlVuKqao2zqlUMx
YkGUCLS0ZYMq9YxVQdRsv51ASJOuGNUwD9zq1PAp4eF65rZ5wDJMMjrsXpn9+8foP8rbqGypJ0Zb
Of+C9kFUQWglzSofo//CJ9wjvdsG7/cC4Md7X2ISd9EU+RcbFH8UYepQJ5O17PoH8gyV79qWGRpp
0sCyeiKA7Yg6e+afmcK+TFoYD5yAl9tEmr9o9AHO1hwAI+zBMymEGKaFnv8wMysTLoxNzoqTkW/f
xvIMht90A9bdeGfk4xRFFG/febt3Sdtlb5k+GYP35lIaeAIcw/8gIGoAJUWOxeNgKlpaIX4klbgd
A2hQnWRS+Wf7XkFO0QLNF+a2zughu2EwOX+87u+vSG/RWCEGp/oYmrXrimnQh3gCjdL7dkfO3sBD
dYbz3WRX7L4DhNsrHmyr7W5XtEmz6zlgfJumDzgqI+w+1/ClVpdSpjjfYLkJ/qoKAf8ReFmzfF5y
flP8KDv43YksOiVQFwh3SgR6AuHMPdRahfIKV3ra35jzC9a4m9zjG9T5cJJa4xirxh/VX5AXRSCH
6nx+Ppft9LvfGdcSEGOTHx62bhe9J1y9t0WI3k8F8EqspLmd8NNnMuKm3zMcdQmA88Ho2QrGxIC8
8wb1WrL+v5FWxNIXuW/uKhzVGGD1k8wIHWke5pQSCtYvelZK2v1EAlhsSpRqNKuKnSDPytckhJaA
TwY07Ldcp6Vg8JDeiQ/4/XeKXSnOdSn0SNg5THg3fuwWd4sbEshRqvsB2g1LwRS1OuVle5HT3WXg
tEOo/AoFMGUP3KeJw2zGSPrvXcTwUYGfAhtQsqa216SpmX9hWa1NmKTswqb03TbLbx3ue/Eqi4ah
5VA/G9oD9jAWSjDytPAsu/1b8kx6JN5KJNEq3RdUyTVHcje/MyPAnDQyWLSQqt6bNTc4DABhcMBQ
JajVOmtl7XPZSnRpRm5WW4TzbPVAypGGLKXrBw4FkGLzY+nPFlcP05gJiWtmYuioUCXKCRpSbML8
W2dsITTMm9OryGMsNVkJfhhgdOQ/jaEQB7FL+Z4zHFFIrlS7GlANdE/r9EQLbnu9k2HYAoTk49o2
6TQFO00JxNBvExGi7bKasyc+mZMnl7wgoRF/m+Oh7Hb6dz/tqYlg98i5ehfV8PhM/pW9mTnNuaZ6
ZDnAi4kUnhLIv3uGHT3WcdCssDL40Er5TCmZvGWNI694vXkIgIl34aFGnG/aE9iuiahUcBjC8ULi
TS9ZMJbq6rNybjf5p1rCoV28lwhADPhFXFwnXZo8597jH9RYpVRmVvFtNiwyHD2us6pWRRsD7msl
8gfeGmTbwznbvyk6zn6/5Z1ihElx+6OluFiL0wOSPhWG2lbqIcaMPDP/5OwBmyfinAWn4KvQarAx
cgnwcfQ2TNCTdktqyp1ZCsJ1qd07wVLnq5wyM9Fz2Vtl7eY9jlT1AoAI5tYS9CHSqXbQnasW3ml0
N9qNKz+LYfIz903jGuldr6+LXoUoqcddX/UNkv8hV1uby0D2VzIMjJjoU4Oy9+5Km6JHNDH5WJ2e
QHwH5OitwCXgqIzlSJm9g+avt+pF6uR3jZ/YgBjDSs35nzhsP0/HyuiDI5fN2z4B9djHDaVhinal
dXu9DB0RqHESU6mTp9/0zhy9OdexTYwA89jQdRRRABcClObgfuqWgjZYflk3gX5gGqyA/4x8sW4m
svf1aDZuPy0ZPbrJ2cz3wQ8JC+iFZF+mSxnwfTPt7008xgzOU4nspyt7k4cMr+OrvRHeVQLB/C86
g6ja94bAdZhITyzdEvcWJNsHbS+JDdHnXTwjGIB8EyiUJ+eNxdFl3tVD8h9iPUf0JuHiZjo6D186
wbFal5iDddfEHNcqC1Wcy8jtM2aMIZTWcfXhQirB+map/T/zlqJMBop9dooKn8UkXgtfjR105FNX
A/8kTz9Uvz+b+wuk2vUHlAy3FPCb46Xf0gQH+Z1yT1zLKfn+D/nFa/pMJuL8h8k9vwkoE85hwsf7
tWtRNPObDB0l1y/6OMoLX3RGnpvRKAZgvbM1MOWXMB21lNRXEiCqnPfo5B8D2YJDiOi7HTPb2ug9
Y1ADeSnSZPwSvpU++c7jE9jSlZWoPbhCMrJs2A6tvYjjTYkuwe5I/R22wPeY7E8D5/GoZoW0mtMC
quSEvOXxA1y/KbnYRaB5nsdb/06/cfRwYdI1oWTcnF7252i1xGYv7sg67x/uw2XsNe1FfuwiJh24
TLJH4zp/M5BF1brWDX+dCn3Zm2a5tTxW1uWi7IYjSknScilJ9I1ol2V10YkO2giuACvH67MKZR6t
Dv0P0CNv3mmoP/KbBbxLFJxNpo9RSF7yd6PCpTvbxsksTNecKiMOV9FnHNGuCm1TvLvtmXOiZXWJ
byvxpe30Ce1N9lkR+6wLtVCde90JzgxZkDiU47u6+n474TeUAD2tAqL18MyqPofTrfKgIbIZfvZY
4q3RD9NjTaHreW6FVtgl/vP4i/IqERE7jyO9/Q5UXy2Zh538Cvz0YHB7ZeNVcd1+nWv1OnT/d08O
PcVSt2u40PfREXXEG1s3WuucWCU+GTNt+8+XU0mW7HGoGZsiqZzaqk3Y9i3MO7bEESY/oI9sLrsu
t2960+wIcBdDrTKlYeh9KJ3GkNkwQ0+qeUXF7SXuIvyN4AWhXosGYucWWSCmteIKynN5465u1gxM
zAXu5uxLWJcFJiCFxN8SrnkSR/AdUdmvgXhS4gKDPYjQieJSc432xQtpp8jczD/jUJFKMVuehp2R
2+jQ8XUmi85XGTUvJE6n35vabqLspPWImlxr2rJjbRMUXVO6kHXUUspA87WuLqUW5F4q0hf2sBw3
gyRDq8jxxFdIZEnBKVLUnV0GfseiyZYp4inpXlWv+nsRUg6SFdwyv4izzVEvz9dGUQnNVgVKETMe
xfx3tt19eLJIixwVSridXaFv3NKSmujEWjB8qCawS2ITIAhrwuxVnUuDGRDapuU37zNsgIEmUQ6O
kYI2d2r8FGIBUJ7ZHgWzvO8CVGh48SPnVMNTPncUPuSP5sVPEle+erS5BhU9gcllfV+h39ZXj+Tg
nVS+bjSBGgG7zWY/J0lfVsfEmr3LCHM8mrvceiJkXiSYFTYqhEWVL91Y61J3lBmS5N8QAHnlbL90
42EbtRD7HtZviomvPusnuF6/XBPd44z9d0FQz18+vDQartFYbrpcICRuiqY3bakKyB3RMFtrHFF3
ZKUQPSOtBtoS30KK9E88Gn2d3UQewtXN6iYTO/HMXJjHZZfgaV8rDtq7/TlSHQ+fywC55u0XyCT2
VI4JdNCP52GE6TGHXh74m3LRnPtQJrhMeDi4l1IccOYkgiO1GJW4FHui+D6GNs9qrd+utwwe2WCB
NEzzM/zQTXky9Sdg/X8sSnRgCIAULlhZAMW52gKtY7dnhQJJTWxc3lS9qYz47smSrJYt4X9H+HhF
vyHhU6FN8WIz9O7JaXZwpHwDLInF2lObczfT4cHOr4C1OnsnEawh+LzyoPCxzD2N4ijGx46eNGyq
QY9gXKu3ohNA7PdVVGArqOMWrQYtJXRR/LGKgvwg1K4JKtphQvtvi4+Mq5n8IsQ5jI3syPujCzSl
KeXbVnCZDEFtu8Flqa5sZjDUTNyE3Ag3hZyOnOedMOl2U+oWHybtA+rywhYxU17LS/Y0AC/FT5/i
TL4MH7cHibCWNMknrP9v4+B8qHQXJ/j44HVkjOlSjAYaK4dNnRAdvPjHG6TUKKY/b56HlSgA5ucU
ap9jt1TUiWYdzuA+GHe9SqskUGl2S+vPNX+R3dW+LeMPPste5G6AOFB2DSCvHTPj08JquKJzXc8V
BHf1UlPKwJM4BraeDjE/zLt2WIf/dXCHXpurQGK9TtWxClmLDznXvLgvCCOhembbpf4fdMgtq8Gj
W3DVgdpWEVbP30DT6jo8vLBGSct6nmTmNplXUVGU+b7RyobiCFpgn3ufVaL1LyjRhQbm0ci6FDCd
sEz+QGWowyKhAcwLSHHvq/V/TRAxO4jCbYpeAZRus5m54K6rU1sOO84CPJoZ37IYOR7N3lIISvBP
FywMozEGcfhe0OOqiDWjfi9vK+DHtHlfxkjdD6FJj20ZJEwa8jYnx4dAfDVeAGujeCghp6Knchik
jf6sfw4t7aZKbpcIk3Wm4xPPOhwJK4lyegWj6RpfD780TnESf4Tnl/DiFWqyEcvxajtpiHnGmELU
PhBz8gLcKsdI8YVdhKfjBzoQ62mUIbkYDFPOMGAY+7FHV5aTm7Qp9kDPPeCk6Y8lHR6Uw96Czi6v
RyEHqxuAqQHSGQ2ctW1H5AUKfQSQs1ZUqvAogKr5GI1zQiiGNNHxLuR540XBdrbXJ3zOxXJGE8k1
AjEs+0Cy1n2fmvwdw7ASD4/J6PBespmRwPyP7G1nMCJfL6ilfuoFz4EhuPuAPeXbFoJvIihFngjt
HtNyyEZXYZTiqfCVHM/QZNny6poo+KewD7CNmwYA29unSrX8l3eWDLNzGUnxpLq2eb91ah1xGsWa
7906KcevFl8yY8xTvXifMA0ZelGkIvofXx4LHvJEgr+yq25K3DwavHthwAW6J2TaKceJnwCNksBh
BsRbV3JBZXOJtQoC2msSjr0IdmIOW6L20iMUGTGwwv1e9We+bI9aD1P3+o+Jk0bhx8ONepV99cTN
eWGMMyWwNsNgDXvy5Jybp4AA4AKYmDDaXeqDhp+8O8rCBI1nB3G4xgxs7Qu1ZgCftQjkknZmHS9f
X8HNMU5v5IVwICzRFXQ6IsqwTT9mY6bQgCB2aFUrp2wwmBcvUip8jK6fofr95MmHwGzeLLlWp/V9
4yv42suHS9+4roi2P0Mx9GGQCOGBfdyvhWT+0n99yqZYXQiXcuVvPGNN+ukZWOCw3NARu584r1HV
M4jg49NZKnf9RhiO+SfJACLIfO3AjUNrCo6nGNUbHto0eXbBsdech7SZv6p/VlylaO4+cLbfWxUg
I7nQenF63/FqRveNjoUmT19buZ9YJujGWnzsvUtxaKOJ/ATguJRPU5t3A/3EFyyvhFXnOvo3RF3j
DJ8PG34GuCUtB4yMVmb6+eccfzrF7RJSGksXCMA4R9DUV7pNs9jl/36ENHVBZphI+8UQjebBfRDO
ZVASiWawroSlqeq+PVDHBiG0ll6pO66407pgUQI+CnapVysI73bfxz24uxZ1DtZ6w7TXt+7b+Ggs
GFlG1ZYIDRQT9fuYVOk3ZgJZDoamP1HTO1BKLN/BEn1BwCUaLpH+0xhSTAOacZSQujP6TdHDEkCA
VPT2CWap3pK5pdWDXZgMKukR88+xCEGWZ1w2cJBiMhGr49GJuakof7pyS/7Gn9NapnMAIFSDUEZw
JhejVilqYyyWHWWGoeJSIyUe1wWAzY/dB6fkPztM9e+kDEX7jsEIEZ3GBsqAl5uSHlNBbjGuJbly
VCGSS+NZ7Fa3YxAoeGBt9BN8OQguhu6nS+ofLGExZ/V0IFJGoxWxZR98YeFw6y8S00SADFeWAOa9
nKZir1Rnfz4QJDItDNUOvWF0N7vog1tjERiSg9Ujxj0xYAfld9I+4nG1mtmp3fUq1D2yVCCWtsuW
sobGrcOPg4Hu9eXflCgJFe2V7j44q1TIQLehpIfY3AwdrIFwtmhnsvU8bBKFqgk0ClA+8qpXFchN
w0HSgKRO3hZ5p3F6MwBcSkdbSf8vL0vW0/pQ3K7/GK2kD/4DH6c+JUeSbu//QL9Eh9OlmGa1wVTz
dGTsuW27ay5YAePeg2CcMLghMfJZ0Kl880nHhemp0MzM3nTDTLhHSYn4Qzg9gm7iqOcoeIneyGzP
k5Dje8/wWjupuNZ+KJ95wqAR3jm2ScDTgp9lLrAF3ptZghf1I+GPwfWBnMqK1SW1Txs9qIZLjXIT
5hGlTjgNz4Hy9DynJ9oJGrMy6qvfz3vZR2NIWxSNkj+I3ziNi+MXzhYognCepUwBPY4EHBNT1sAh
1j6pm49UE/BQ7bwo0ycGAiU6VDLNEhuEyYfmBTf3g1IZJZ0hSYe2tUANtvdzbcAESrLe3qfXwTAp
cFFNmVvhzm1qJeGlNf5Xp+Uz8glf7g26ZThQklmifUNVNZX9jlEnt18xOHBShGmhAyNOCo2957AW
oU2og9TNH6ENP36kcQUZAevd0Ky7Pe9qSEWE8y+VFmWLz+pk6gFh69jYJAClhVSNUiChPZgOxaem
xngX9cJYbZd3objUdjsADMOv+3yo1a+xxo0H4kPP764PGz/uTtKZAW0szE+OPbgaULUKlXNUdT8G
o6VkwDmtechkjH28Wm3UQdtXtbJHGshDOXQZncy2f1AfntfrhCNhv2ugGluRmkajdsKGygKV4Mvh
lWb4fetvUGB7etJXCIeWomITwtpkBwgnQpr5wr67XWJ1WmR7eS3/k199imNCxHij85oubBGSJAip
tdzfk3LBh5YbNG6bt/XdO4tn4itFIO9F/T3RcJjlAD4XmZ/d2hXaRSjcpud7GIz9GpES3TCxmL1o
11Z4gGU4UEhhJgsjbDGue/hpTWypfO8Z06pVMe+WxdwLS1YmfBzflCT+aMxJdMJxkuylbV5kbEnt
I/6cUoerhGG46uyNfcYztwTqAsLoNRgQn7pPv1RUfk8DvEjwFtc6YgxdPO0NyS3Q4eGJQL24jO67
1SdDTJZjQXuII0vdkEw+FAvfH8R6BrGkxunqyiFiirMXezO1Cw2ttccE6d3wf28DCkRh32WCNrR+
DiewsWUSKp/JvRLQ7RzkOsfEfwKR5LGUabw/+Azwcei6BlDbEO9Z0oQTS3WwkT/+CATfVSAGa8qY
hoY1BlducpONxqyHvRzDMDn4bhwiSNIr3iOO9DlipcCTq/Z2I+Nk0YKMkXi4VsO97OlFS5Dr3N0e
2xUlE+g2HQJ9rZ00iVmLIynhR/I7YQj6LLFvYJWNz1rsk9gPIwrSbFzcugCiVqMhVgLZp9clA7l7
69Mk5agAGFdqmzzkVeU0sqFOIegm6tXa+po6UgNDSbK2gx26//U735eHZSdjIiHBiI2Gdr46FLOK
L9CzFNGvxeNcJX7542CryN7UtKjAscumG5VwgATGp9cgjqzbflAPiOKxcerPl2DRUf8VZGkW+suE
WO8v/v+roCHk8X90UYYNjTId4bdMIoRr4yd9U8Zg6hwiTvwGJ8u3bu49v1WSoOqBCo7BY5xBXWhC
BRWePqLnOmozVs1Ql3xnr1g6Tb/R0fx6F96zDU013GWhlsqey/20xeMaBxQlBfUzqDCUxgZHSp1+
Awvdp6MtBKSuKmeT3TeonCKs2qtGddWpYse5N1DRq9sxJN4UCju2pZbSAIpmlOWTQM3RTbixMrhb
5z0g2VZyKmfryw0oE2itibkHHqF2y3+ZajojZluef2mweENcdVjP1eEBHj47GcEdriySNxRqhvCe
PI+HSQohbFHZzqkedXFwoOUL09muJgFc2Sfi7OBKCXJ9f7vb7fbbSs590B+10MKd83OuTIpr0OBH
wqmScBNe+qVvYtZCxnR/0bKub4LPV/nkD8W1L/JW8O7es6Z4cSioDTcFYMOdm8BRRS9sA7CVBhZ4
albDT1C8bioQSt6e6PDUIVSj7le+Kgr8bmGqGdWWyzZ7BoDwcvZC9FswyX+j2Fu5H0E6GIa6rPTb
TCSoNDrH2MJgTnI3dkOhKcTewSbnHcqA3XXe348tjCKztJY084OnoJBfw/OczXZApwjKbYA0GwKc
+XF/H9qBrNCZQI4/paOeIVKIW1xIhx2IqenK+x5BYDdDOzOwOlafZt2yYKlb4BRag7jLp6kfjiBY
koq0F6GpDjWwfCCmlOkbnVea20PoilBnkv50oLDINuRKWekBV0uMles5vindWYvJtOQ4fox7HQNK
Fyc2DIp9opg6hfl2gJJqSrBuQgf6kUKNdguDf0YHZvJyoh/C+qsu2l7IbZ9d781RqLRZ7ufv9MFT
bBN4J8pk/Pk+eSTw0AhbpvMw4gMG5fujjDQOUZz5EvZDtNfMcgYnif6HsbEyAxneOPwXmGggyrgx
MTTH27XRvnczeL1Eipgm19usAEPzA1zvTwGDT5g3fR8QCpUQ0seOTR5qRiO5B4Y4Mtb5T/WunFnB
iESDd97a9NcMlIYi5Pdz5znxOop3mG/GIN2iWskQtlABV790KXxXF9J7PSXosy93bbqwg8LPYjzc
HAAZnqE9ev2nLcS3It0n1GKVdgUYN8rh5XBPaOSR7Aq4ggo7KoipwOfMnqA7ctCj8Atvd1ifrt17
jCPlmelaLkSI/vBFOnCb6WLor/tCFTTGn7wPCX3VYyQPLFTDWVOOQYxyxe8YKLq2oy+MJLl21wTw
V8augQjO74FbJe6DMjhHJTghSycp3v0pItCYhmsj5TTgTBBPeiQ7egf9GefL8sTEFd+1LXYRYx70
3T3QHSUn8xnjxcGGhJvzk1U+NBtChGToI5CMfWDK3B/KmqxouzCVdwrVw3ysdix3juPMJ/NyQoiW
048F7fMRsQIrf95LzO/fO12XVHA5mvznOG20yk8+rks2n8uESEmVn4FuJW7oD104ytnM7PRzahuH
rBc+CUGNVkiKk+KSmPSGNpyh/KqFWBNJZqfDnwelSCYS6FJzYog3kl9epFvZKN0/kbEI0DQaS+jO
weAq13yu3Rx+XMnoUDQIiEi8Ln3apyGRTZJwR1sML3+2FJihWf8isOboZujgnq6ypICY5zXRw7sf
DctAJZ8iyciH9cLqAFvO6u/U3fCNkUcvpjHNSsioVpnGGYNaZxmgotxQaAbPZVrPQz1NuDqq4qMq
6ja2+Cid4uKz00B2vQw7LtYcL592RHiWRKmpTkVVlIh1OnQWGzg6vhAJCFVdfW5DM+v4a8bao3X7
ZQn3CBRSPG7a3CEIUNQIJnwpQZXMvQGIzfShZmKLlqW3HwMB4gFLivR8b9sRn3FvUCzB5whCPnkQ
i47J/XkkWQAuK+enl14sr3ENYD+QmI0YWjzluBFwSiSnxU1cQFnBCBY/Ay5jPgj09mHeuUXR/TMO
VC48MY7R6nP1HobTHM1IdcLppeahu8O4kdQC+o6Atb3d6DVUNfjx/ocwiolzdpRqSr8OEl7lERfS
Eo8GO2yXjufiyh7dAkivLAcnMzXAucStlZQRmWuTFPDJR6efHs9pCLosFYzdRP28ypByiqFO/O2t
0pY0sWKd/rzuB7g9qk6KMTAC9Z+hxxlEp85hLtoXYWeWbjwGdgyUJm6x1xxrl6QokDU4iKxncyG5
zuxZxq2Bgd/8LW7UhFds6P3QiBjLu1mWzb2Q6VffUK9bOV1VPKCHdaAHDaHEECzi5MVE2cDjURL8
9MZ4cMdozCQLFhc6VXC1v4J9Gb7M/QK9Id/JePD+BknOCK1m6Efew7YBxfan7YefjKtTrBQttS1N
BRrTIHdKFN8TMbDP0nVb0iOHFFrs+6ITA3rXZMYMwZXkeDE0lPdBKnQ4cBbuxTWKsSNiSGRMNxYu
fN6n2UNGaPRXvt94O3zNjyr0Hps0V68qLfdFtLlwab+rBEvhmk67NDF3U9dzI0+EBljTRCU0pJQO
GaFnZq5doIg7K144taTnEoRD2Dmv/iRiRSb4n0l8my+2U495S2wrygm4fg7NS7EVZ8byFL0jjWYV
YSyPdJnkirXQUTga+0J2myk2EJX64TtmoKw2mz6iMb1b6nAizd2hlUCnd1GNaY6oZiZnZOyBjIKx
Z6pIpZxgQkebJRH9Qe0Fb9zL+Fj4nxDdPf2KgCBui0DMPl0OoZHKNNV2UVp5akhskcdpn6jaADjB
ZWQ9Q8HnxI6/506y9VvDCxiOje5OHlOg2uAmOlOr4xAg++wMpshET14FoBjeOik4xoKXYKPlqG93
aLuPXkJksEjrNBjHI35X7S2Sbr1b7BEcWh9LLsX8GWWTvPvBw6TfX72A6ymbq5zsLWDLVy7aQPUH
3atXt5Da0YYX2+UoSiHjmITCv/+fY/4o1fEIfklNniVyP5WOYMCTIWhD4FL02rhWOgfSAcMbwtD8
uSU/1jv8MC8lx4HFuNmkDoraXJTMhluxXXkb6qXs1u5TTritK7I7hBZ1WjhSNdxh4Es7pwdQw1yw
5fyD9IZT2WAneOtKRz4eA73PnYj/ghrrA6pmJJvnUwedkFzFa2IeDueuFFP3J+lzAJV/1IS2nAXe
OwnXAa/cDHxLLqgt7q5fDOuPCn4jekrukXoptsw2aMhXrdPc+xJfFHT3D1ffi2DylwLGKGA1M0CC
a/65vgKHH4JUCvZkrdsEUrGAT4IqoPpxBgza/9Id73Lcbz5iRYFPKMEhtgpiQONBoAYbGft56euY
3EJ2szulyv7to/NAoS49jrGdS+SrVJaAh+73TjwOYkDlJBoWsbo7iXCIB6SM0cyZp6BM+tfGPWdg
N6rtNzbBQPxCK6FDHmMHgpRwL7zoLTJXBHSQG3TmbF3Bm550z4aNHTnR/WXHe3yI07IlXVU/Lo9t
RuGHQDHt+KBlLx+LzzBMm4B99WqFYGCn/sfKZapzQjVRnYFHPiB3FN+b0XxCYQa+tVH14ENSEouP
RYn0+vARW9HS96sw8td/vMDSMs9hVi8YoCxd8BxB4DrFiolLXmLdvMeV7cI4CT5NUHBgV34f1rWW
/083BR90AtOstVd6UKjKIcLY6Ifg7syiIChYGeSghIWHrMx/XSM2LewghQ56XKW1417X5gKYFvD4
enBGJSioQwiu3lugIHansWnu3sTLW5IBK9SJJnoGbEm2nMem7G4me2iJiUnnuXGGWa5W3HnGKooX
EtnWkCx2S2aWMvfYiCbczsTlkLo0y7m9zQQhKsyDAC3Nyxq0/sg07kQE3c8C9+gG11fZ9WEiTY0Z
KFLzZ0kJM37Aa070pCCGQNX7Kq3r9flLX28keO3WoesLwYsIl+RV4ltvBH9iXD/5O/Bkp44fUFs2
vBd3jicMEchjVoqfoyIcgTpGSXuwYfeh26pHs3EnZ+HkHztOq0qQ2uXisPZyvKfST7rYXMdIYSn0
4IuKTrpFkyQuU0X2LMePFX1isnzs3Yf9+QFCtk85vHhgGUJ9ayUbAumT63pa+vRhrr3gnqVaghXv
oMr6PYzV4PewMFsK/Va8sCsE1b9Ji36vGRm6ZrXM6P4zLK4RUniN4FY+lOJyC/tjj1ystnrm6MVP
d7/GMYIbrwpH7b7GsO0H+vxx4bq0hg5sEYmS0dtycLs8yNZRXY3UNezrZrTkio8lAIO/t0NP8F6f
WYq34JZXaezUbfDjTYfrgCxqqhDc/gnwgkZRjss5SRhZIZLtTIQFAW4jxpuS4bkSQinBA7qqlcM/
GIS7SCPlLBCKOwYpb3ozyVHMjLthXxYT9OpmJae/jUfSb+seMr04kQqRwdcYjJkRk9WWVNdTbd3K
0k/KudlGhnwotM1ioB4VKfqja4uLhbr/JrsqA9s9Y/avz20Yo6mbCeIY1BAdvoVAJpHQAW2USV3o
I8QO13fq/GKQgePtCxDn4Xl0llfouiycZw5b2bgO18G7AvQoTPIWWp6hlL9/j7/ADxYIqcd4IUsd
oCYl/5CafaumeHsTt7dEYypHcNUNlb1r5zi/bv6abLDlUGgdJFVQ9CUPO83BVN+vAZyvZmdsbNBU
F61ezxidFbi7Cf4EjrRZoEmglHRS/RWJcAVi/b3AwwYCwOMJ//xgx4V9SFwYa1V8b+261KpQRfdY
KMhaiYprpLOKYJAh8P5pKgyqtbuHnv2Ueonk2PNKIMpRfZzj44r41RAFZmk51nX9VcyuPGH3T1gE
RkPQeYCzNthWRn6d+N6ZQK7Mcs1NEGKjQstB5PTwliapjAJ1AySN0YsiXyJFqpzkZdgXHOLFF8Qy
mqrzvRyUDBEhL2nS+3ryIWX80GZ9A/2Xl8CnoSwfFg4J1LE1NuZCMZLjBlMzVCqOsMOKmI3+b38R
JtZIOLP6KucwwjoIv7BliyW7njVhZJwV1L0/kesZn9qnAPLoiBksXdvM+nJmvDUWWHrBEGgivgYx
9NmlhzOOM5aJIqn2mUULTXIqiNbpQejktTEk3viM9J9QPR5Ek0CK+1vGtazyyGYMnf06XDx/0hu3
QbByfWIPAH+hcM2rv5YZtsGRM8+pGX/fLewMEiDHtR92A6aIL14fLrTt1Wvpefq5Hd5h7+soOOE4
vwA5//IAZU5zXBrBumSGr6gbC9GTzsX2J7lfuAz0ExhcdfhY4PvNcF1jC5UoUHNoexi/WOjfLUmU
+NSNaNyBa8D/O9zj
`protect end_protected
