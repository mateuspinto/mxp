XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Y���'dbf��n�kl�AۇͽX�0B�Dlz�y�KNpZ���?�t�(����Bs�|%���0	�9�"���M�S~A�a%0��SB�b���hY뱝+{��`����-;�B�Z(���<44�/��CsB��g��w%�p��s�Ph��)�^�Ŧ������J+� ��J�8%���1��@.f��J�`����i ��J�=*U��N;����n��c�ɲ�/�A��[g�Ѷk��}��{[��4�c�L�p�F�
(��q��� ��khg'o����P�s���x���8��%�*��U\�k���tG�$�s��0~{g��,FJC�8Iӑ�ܛ�B��S�kҩ���*�L�8"� �R֥d�xfm1�M�GcR��#կoG�eD7�W��>�Oh�dn��Բ5q�m��ߪ�.j"�G���ZR:0��"�K7�O���[�_6�S)0K�^��H�}��dvZ�O��Kp�A=?�om�.�ц�\^�_i[PB�U�g�P���1:��V.ȥ������Z����pyNߥ���}*���|߁Ԯ�<�f0��ʽ�ސ��� ��n�fg$�9���'��AajlJA�#7������o}4���|"X�b�'�]���QA�tdv<�*�tY��!r�c�^ɛ�°�˨U�*���R����a�M��)�r��<�"��%�u;���,Lo[�����!������0��Q�e�u���s���e��<Q!���*XlxVHYEB     400     190��s��ZإS���p���v�/_
]�1O_;���e_�k��~�F%��B{��8��9p�9v�����y��ָf}��##�ë;/��+7���\$�\I� �����:P2�>����o����1⿆W[��^���Ԍ=.�*HZf^����Z�� ���dI�qOi�L���/�}_'��s;,= r��d���0�cj��=�&M�����h�=�8P���\|A���X���\��R�P�vh�y��6h����z�(J�W*sy���L|��H}|�bUٮ|1�²��n����ziO7V�?1��}�x�}�&��b�,�Ѡ=4G�7�'�j��'��`�;�A�ʡ!��^����M]�mF&:!3�<�?�D�ƀo&��^�d�;�{XlxVHYEB     400     180�;�z���ˍR�t�$Ђ/�T���yy���Ju4�#�%�7O8��8Y
��P�w �p�Bq)���}Y<� T���T�ĥ�C�j��G+��ׯ���}7���cT����@��>h����7�ܹ<���X�5G�荍9�2���_ XTι�*8��&�ܷ�8v�������(~<�Bȅ�H$
7������Ҝ�]�kAf��-GF��V�Ԍ�̞ኰ�����(���|�
�=C�n�LoDJ|q����W��|�v�E�t���<�S��<k[����U��ך�Lq��&`����	�������9���i��̈������.6�����f�&�n�pEE��r�y:���	���9U�ب)}�XlxVHYEB     400      b0��.$?��@XlZ��xx �*.6�|�;Mh؃Ԓ1�6{���u/���������Sl�x�@�s;n �ɫW���\��ڂ��V��t��,�aF:  Z%�f����v��9��x����%�a)��}�6%���۬���!\0!j��Sn_q����{�k�c�V{��2x����L�XlxVHYEB     400     1703�d��/tH�j�Z�i�TM ,z���tL�����B�G��m��)$���_�l�0��Oe�b��"�94iB�B��U'�B��L��y�2�4��o#�;��S�j3���-B����RMփ�ƘW
��%��j	�P-�"��D�H�/��,J/6��G��_?9	t¾	tF���r���h�8��<$�)epL@�7�j�X�1������F�4�0F6�����Hz4llRyu��i��4=�Dl��1v��!wqygF2 �2Iu����Z���w�Q���)2��#ڨw��8R�n���7V׺c
@�Z������Z�`6��S��A����B�b���v���m�E����K�F�I�}1�p��<��_=�<XlxVHYEB     400      90D!���]=�7Rv�?+L,�3%:Sd����h(�J����~1���i����X���>�CЦ�v�`���Ď�C|�0��NjaH�
��C�s>5Ao'h;�����yv�b�8����js�6�%*qd^�`����	��4�0��AXlxVHYEB     400      90���4�T�+�y@��5���tba�ڟ�ȡ*�9�='P_:{�w�^R%��{�NWjA�k}[ȑۯn@.W&U�Y�!5G���d�n�ė�&œHJC[+�U�R���f�Eg�EZ۫}LW��*+�8þ�\�`}RZ�Ր<�+�XlxVHYEB     400      90�Wi���11 ��*�O
QV���r�.��;iӱ��V�l!7��@�Fmh�z��yk8BG�bg��w����Q�� 5�K��;�b8�`��=�!�ڃYkDr��=� [A��v��z�aV"�j)`�g��.ˈ�f�XlxVHYEB     11d      506�6ڷ����r0�ޤ�����z�'��������f�����#u�&�V��^�b%��� �qE 1^H�䂎p�m+