XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<���z���%)��l82*Ue7G&a��-{���s�>��C�yնtWw�1e�)�u��Ƒ8��h�ՊS;,f�0';��O���K.B�H��}[�A�m01���ݯ���O�����c~p�W�����0����ʯU��L�q�wl�T(��Kv�K��o@�F[z�|<|�,����P�z���B�R�فE��
��seD��H��r��*��ߊM`z�J�WD=[��)��C'�w�t;�)%ғ-AG��"�Һ�Q��}��p�T?��Ԏ�iE4.�'��T��CK$��]ٵ����~ �3�����c����!�9I�ct;����I��l占@od75�>�q�#��n�K�Ζ�x����	��+61��	�]�0��������]&�%�r&

��M+#]��Ǭ|�:��嵺�xZ��=&+��C���h y.%a��#�}�f���(x�u�K��Ύ�w[�A�8�#.��W�Xm����2y]8U�ܨt>�5J��x�����l�׆��7L[��ǫ91�`��(���bt�ۈ�Ձ������j���oY��o�Om�쐢�����T�{��U�S�W+
v�D��4�T����W�X�}�`����Iv�$����B#	d;ƒ`m��I�'R;ȃ����W�
��:[ _E��rE��3rن9���< �\A5�C�P��52�J���ɢt�ǳ�`�3}�\_���g8F���Ɏ�G�=��t&XlxVHYEB     400     1d0�!� �Clk��Բ^�[��Ng����M�ld	�go9�]Yz'���l�3I&.�>�U�#�uF ��D�;�ӣ�ݘb�O�#��K&GX���bKN�t����8n��E���`8�RP_�&@]�_��U7rS��Eyq 4�!S�C�Dݦm}DD��\wN���O}N'e�#V�A{5�"��^�(5]���𓖖�ٴ
�G_�q/����pB)�g�~��ғ�+ݹM�`���P�d��.��x<Q~-�#69}���w����{�X���P���|��m�b�?-�����gIe��6R�'n�AJ����<2�^��)�5)�N�s�]!�+?�g׌�z�'�+���ٵ�k�lzx}A��jg�Z��`G�R��֏���&F�{_[���X����.Ό-�O���ج7�bp��5�~��x<���W�p~����p���S�C�lԥ�{�q����vTR)XlxVHYEB     400     160;ݺ��,��
4�b��â��s�G�rj܇[S��&���t���zjn����uY�ʶ�Y��*~������W�,�Nc|i�W�ۦ��q�9w�	��spU���K՞��T*j������7�b&�y�9=�_���4�(1�/���	�c�M�����ZI��� `d\�
���-�-eƩ޴�X in��jpF�н��j5�"���U�UQ���5T�tN�i�qʐ"��^��^�V.��y5��e�$���DFO����K����=�M�S:I{9��,��O�}��2�N0��TrtgɈKA���eɪ+i������N��:E\����F�T��7�I�XlxVHYEB     400     110M�\E��,���=���7�O��t�!W\0'�o�&�-�Cj}B1��K߹��j�ȃda��K�}ǘfy�SK��z>��6����D�O�VP��p�����¼淕��q	�N���]V�^��I>[�m�EiYo/����>a%b�JY���E����h�Ԯ3nD�C�8u�hU����>���Ek(6�׳����~���;�L��|?Q�E���!�*O,;�9���^�}mo�J\Q%o"&ec(�¥7�n@����OXlxVHYEB     400     110(���E4�79�	�*183�-/���u�ۊI�{�Q#{t�������X	6HRO��=ӄ�a�?����utGf�bB��s��%g˩.�^�KI���Um��ӾT]������� ��)���j�ޔx�JHR�W*�3���u X�?����͹����iIt������]E����c;w��o��aN�͚������վ��
2C)*�=+�2ͫ�$M�Hd͝��5��|&@�}&_��w�����M|�Zg�S� ڮ�.XlxVHYEB     400     1509'��6ׁ���s�2*��t
r3%���ۨh��|�ns*��Ɗ��G��0���Q]Z�H9������s[s�5�?v���i	��7��\�u�<�Y�q������^�B��s�Ƚ9=�?Ɂ!�vԻ-��a`H�:�a��;���>��-��2���ͻp����ۓ<6ٍ�uQ��2�a�hj�ڥ�r�l`?=���-�h��>��18n
���y�����r�������,{>��ϼҮ���OV.)cn䏲I?I"	��DUG0ҌPv�����HE�����Eªo��O���W���p�D��F��٣����v7��X��XlxVHYEB     400     190��Aoi,�δȖn�׾ɧ�dn��1��p�����H 6,l��M�_��A�Ŧ���߂ZE��T9�?�� ��z��"�g��Ű]�?��E�zfȅ�^�_�z�;�;���n
����t��1C`��8!P]	�QF��X�B<�6����2\�;�M{������L�ͫ-(%m|_,�NTH>G��.�c�KC����o����5?�!��	��@��Վn�y�a)�Ƶ�z0�v
}�ܕ���&�b2���7��zN �9�;��Ƹ`��#�����"���EZXU1�B'��~즣���K�x�3]v$m2m��Y�|� ��JR�n��� �E"1�̅>7������)�)9B��V1M�x�2彦�5��+��C-�o�ۼ/Jp%��!��A'XlxVHYEB     400     150	P<���pJZ8��@����y鼎Ȍ��W�j��M@�Q���CDP����;�HB0-*���7V�T]#�����z�x �N�qs��eL`a��_��gi��w>������'�MN/�g���?V$�L���׮��l�\G-ٞ[�<�W��<bk ��v-�x�����N�<�KG�~���}��~�6��˒�.�v���.�7�X�_����d?������&|��H��߅_u����Y�Vxq �9QDB3�(SC�۔ae"?s&�r�ɵ~�/�r�����E��Z�JCB��t
����oj	�^P팩�g���c�8\��XlxVHYEB     400     160<��"��M>N�Uf�<IC P&&u}��+���X�LD��J��b�쑶j�J��č@�{n��7������ ��$Ly#�$>1�������P�~��D�"��sqZӐ�y�
�O#�t�n�YT�� �o�����P�xW(��e�	���6S��b�B�q�J(��z�-��v�Po˻|�l}�ֶ�0�%/���\�l�G�d�#''IP-��h��p���}��k}e~�ER:���V��i���궼�$�Y*$��Β�K�l���a�(|���7+?{���|ˤfÙ��V4��~���Ѷ�8�Uh}qYj?�P�������D7@�|�?Rbժ�a;XlxVHYEB     400     120i�$��	�'�O:���	����%�M��*���b$(k��&X[��k�m� ����4=�ӝ�1�)5}��Y��9�e�#�������p�D\�H�wi�y���8)Y�{�i�І4"4���4�rUc���t��Z�����G�Ⱥ��1Q�֑�>����ŷ�l5 �F�F�W�XH!W�+%M��ߗ�d���T/u�����QVd�(�fӗ�a���Ȓ��f�"2�9�{l��e:�K��/1�5�`j�>ڞ����8C��_@Cb"%�1��XlxVHYEB     400     1b0��#�k15��\�)>e[���i�ր�0���i�o����s��b��{�В.+�Z�:���5M�%3�(�85�jf ڒ�R�T�W1���޿�}��@+��9���k_Ŋ�a
3xiy�lRq�)��*�dmH�?6&�lY�!L�)Rj�|��	�C�LR�G�Ů��̇i�z�u����H��bI���eY^ҙ%ׁ�H��^Jϼ�R���g�_@o����}�l��	ʜ=��{��ߓwv�����y��z��*cܲ��I�P'�P��J��X�@Q�Y��~���J8vj2�8�4��������
X[g�>^J8q�Xݍ�	3��iGj�����!�O:�/��"z�Co\�Y�$<�ǈ�'}��!�6�pɟ�!�{����f���d�0�#��J�Aoϓc�d�5�[���7�E�)�XlxVHYEB     400     1b0���?��Ϛ�����~��`���� �s�Di��獊��+�[wYU#����v��|RcL۵fF���t�(vޠF�Y!(�nWWDw�����7!�a���u	"`���|\��n��:N��"(Q[�+�,����^�\�>���#��#c�\B�d*qW:n/\O7Rxix7{r��7"}b"I���O�0ǰ��+j�l9i>Jn�@=WRg�u�P-�����Q�Gt?gI]���k��u
V{���WI��6mL�5k�avJC�p�1D����k�*8��M���MΡ	��0�Y�elU�U��iּr�wy7�"��k!u��,�x�����7:�'y4؀Оt��T�3��c�i+
�?~�[��P-J��dy��'�Mo�D�{����G\��XD�t�3�V�N�_}XlxVHYEB     400     1808�oƱ�;tq}VJ@z5R�T�o3�����4�ObI��:7P����f��6�Jh����1������)����.�RN�����9앞��� 0���K�r��J(�UA	���1���7�k�tt �|���x'κ9<"��X`{"0 ��$L���Fv��vY�I�dp����rE�p�4��oj.���w��Q�m3d���qK���q�06�p�4�͡��B?�=|./�<���:qe���<٤c5�g��|B�2- �w������:tg�����&+�Bþ�M��!?.1������`��-�}�&�-�}�wk���K�av��V�-��_z���N� ����:��ts�e�,�JK�1�rn����̶ oXlxVHYEB     400     170z�10\�@�{뉿����8�0�.�WB8��	�z�	�(���4��3ا�~9���6Ӭ�E'z�ɋ�!��>���z^����8�臲��LX�zh%�$Q�/D/ �կ��F0D��Ԙ}-�DX���&���vn�k����w'��[EJ����7�K�����+(���
3B�{��0�b+�r����~w�a)����L�Z��ez�vGO�>K�'��?I�C3��X�Mb��:�B�/�>2��1��+���ڣ,�9X��Dw��A�~唟l��z��ٵW�xKOp�&�����������HO�ި��⇤����$:0�;�2@1_i�6FGI�5<�C�V��P�If���XlxVHYEB     243     100��U�����Cb��+ ��fB0�,�]�~"��"T���E�3:3j�NU*(iO�Lm��\Ȼ���o�a����Z�"��)��`]�t�v��uZ�.�h���A�6�>��H�[iR�*�?��a���7ay�Ҋ�輗��s�|�!����v��7a�w�th|>�	�4<�C~}�k��M�\��C7y�����nX�i��PI�]��/��h`�muC�����E/���Zf/�_����O