XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4-���}�d����:�e�����>����_2~��>/F~m�� \� �����c������|fl�Wh!`�9]a:Ջ�R��H���2������OXiأ�gK�n}�m��w4,��K�xv����ZQ9��-�[�N�<��g$�M`sx9�geq����
��!	�a������I5�?�0z�UQ>c�_��4|^2�N�Vd������.�)�'�I�9���|b�T{̍s�K���i�^��w�D�|�Z1�	���n���
1Gy(*��U��2�vd]�VT�*�ge�xXJҙ'���4j����)*BD6���`z���.�ɜ\*{��f�©Qi��;��(�k~�9��x��6�׾���d�SD����������0�'�5��9u�vy�׈�-�ϳ�Z�-pnb�D�4N�S����!n׫6^x�vMg���~�P���68�j=�`�Ǫр, �O��r(xS��E��(zf�]J�کb4qN�j�6\�Q�+���0����y+���(.�s��sOլ.Z>p��{AV��{7��"?�Z-, �^1��a��1�.5b�*0��h�$�;�v�jQ��n��튝_���z ��1i��a�o���gD|f ;�\��(?���.�9a	_�F��t�����" �4)�X�
���S,�&ZE����a�F�q��K�u�D���;����T��fu*H2��]��t��_
a���YF3�.��\H(��zw��c� δ��l�fsXlxVHYEB     400     1901�L=��k��r������dl��dp�e?��z'F8��9�]���n��Z���T0�����R��zd��z�|R(W���k�UR����+�LS�n_���X �R�%���V��,3�09@-'���z#a�LM�9���a�_~��YjZ�vMa���75����ͪ�����`��!��J̮���\ڄ��n��N/�^N k
Q��}|K��'���7eEp�I-ǰ��M�g��g�[�ѝA��������>��ܣ�&�5����"��n�`��e/"�'�A�a���8`y��P�����D��KǿD�o#��\>AD;T�vNU��Lr
r�$������*�J��`���_ws���Q�&!�6��e3!�>
��6�����m������]1�
���φ�^XlxVHYEB     400     140w�c�W[�A\Ҥ�_tX1��,��D���^H���ɑ�V�g̷M��B��]�ݡ�A[�D�)�LU��NF��.�G��{ �
ᣓ� )0��!������f�)�l��D)�+}?�XU�C[��I/-��NR���=������>�۸��ă(�G@�k~��	�����VR:i���7��4��¡�K=��2�H��ޝ8�b`�G)���2s�R��'��絼/��[*������1|G�v�c��Y���s����񁼗�NLD7X��
Dvg�	^L0�h�}_�6��5ɿ6XlxVHYEB     400     130���24-�e��aݰl�c��ƞ����M֡{U������� W'�Y�*�t#;N-X�������k �CMe ,3k��<QN�?�UJN"��5�侈���e�����'���j$xB׶P���ߠw�Z"��[�r�Y�q@���c�D��v�yU��5s�s�Y*����?���;��zTo��� r��l�}�����K��B=wG=9F`��D[y_�8.� �/�>qz�KJ��%1�@Ʃ�ddy��ǐRM��,	0��Al_vde��Q	ן�5 o� ��l���Zã4j���K��XlxVHYEB     232     110�L���5��b^B�N�VJ�/c)�7�J���J�
,��;����R2�Cq�&��������Kd����#I��a���\N�-ie��3t�s�ʅ�D��﩯jF�g}�!�`�����2gWQC��H�[��3���MZ<�/�k/ٲ^C͙4b���'�U����P0�o'(��w��(�u�˲5�u��NQH��HG���ʔS\�H�Hn c�>b�[j켆�"��b��ѝ���|�q<�#���r��-E�:>��A 