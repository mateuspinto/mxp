`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
eSpHy53ihpilQyYPCM7HaDFB6b8ywe7zxHlCROo3007tPWQvvC7SIeoA2RztZJwOX3SRHWmzHi6o
Bg1YWjqkl2MvdhvC/mrbQB2J1HtByyHfjeQbtfsG700AgfnL/LhE557tori4/3Uk8hChY72UTdSd
6Xwo637RAZUvGyXt3uLSJJrlBLKVFpGmx7mz6Ox6MztO4wdTwhj4yfJ0S13RZmcgFff8in/yrazL
HtPv2qgjoIRefpBg2kIszAhJWniVwDSoe9PJAWczjOmt+QsBxRiz60vyyaEsiikHoI4FSvBQziiB
67x4bzRSId3v9x2z1wksqAGD0v1qycFENbRbgx8/OAJM6NZK6sw/ZHDbGXMb3lWnFKlleIocQxs9
WFVutElDNvcn558/ruaFx1GOLg2XC1dtedXhtCNFFaE0O1WT5WXz7yr4fqXAWG/52rD79ckagHqW
vqXsAicoCiCHRGg+w6vn+/CpAZKWFwYEuRbHduoghoe0FrjR0ZZzQHj7hSBQPaAVrtIfpwh8Oh7R
d+DBRyMk9b4lIzi6n6269Byl++bF0aqPIAjJ1Xz8/CUriw5+9vSij6tm0vqymH0ino4rdQzMuXj+
yFXnrFxSErZNsZwXCLaln2LPiow6jAzE2NMyDqQFisPRtVgJkSy7FTOhXfagJkSUPWy78u2ON4MC
026hIuRPgP1LRwlkBg/itJSJLxodLPFL0E4bQRP8FtZBGCXNWLb0AHdipyhrz6TEQAiwB1uVgQGQ
xy8VZBOabEjm+TT59BymhjyD3b2IcbSR8qtq5e/dw+jsbmM4d92KWH4zc8GXGBQF8xCyPb45ZOcU
FjXnQ6pQ3ex86CyOzRQ5X6I5BqUgwVHVYd0i3Lf01Mq51bREgOlR6Trn2lfSVE9GjV7q0MG7PeH3
1o/LTWYFO9RiLLBX+GSuxZrnkijeQjsTT/FDZGCXJu0WIozvoBZFZaxTou64Ks6yA3GoGCbOK1XU
aTEXHsJ8o+m2jYP2ip1qV8eMpOnGkAv90DbWBqBliUG4N1bjOFesqPFyY4RXdOPoC27gozORH7bz
/GipAeEhytZhrhnYFXg5bHbghSjIuCr5RtH78BnytJEidLAmhXjgdVTKpeZzAnp8HwNoit/pwuHO
FY6vDtiyW0ptkk9fVW2QdbGjL+VS/axz5p95o565jH8U8Mh7t+/a40kzBi+qvhAbsIWBZNEihKaH
zTJz6GHwvUH4iEwOhDRS3jGdZesWBpbb873OB+DYJdspQd4/1FU+NmsG1oDBUOwcPzrpWPo3jaoH
IB6/wYeudFnQBsLn7UDEsekf2F85JzN6HCnxYPVVzPTR0vYfdnv2oSY4+5Kz8r184UnJLla82uPL
mHUN0QQ3pAXQh1tYbGtPnBp+NHw/1H1PrSpj7Ff0fv017OMrOXDY/5wMjYruuYcdqet5B+WAd1FG
Udjjzkd/9kzFjgs3ddxZaVIdJcH3IUSybnLvDF2N4L77XECEkfewFz9zAZarYdsrgZ+MTYHZEPEI
8yk/J2nChmi7bu+afiw6sz27nyQKbrsilwZzjawyEfqpYHV+4t4tKcEfQD4E4ZJ1CMvuA14fvwKr
QaaM8VLNRTc/O2BdC/lO+ttoMQS+7BQ2aBthdxVIne6YpgqjHb4dRpeso1OANPJtJWTFnjXgwmry
HOnRjAtudh8ZBLxvkbaij1TbRik/a/2TwSpFAWU3YyxYz0Qe67VHyYQKGCqahQX3eCEaUnmZcmYU
LAvW6LmxrVUlzpGY3VroYRLz3wjwZ7C5sDKNaF1uv7hYFoj9chfwWcM/IJg7YJdZ3rSsQBt5SP34
FjMVz4qh7pjfsyI016lDjBUmBW1PGBCFmNG56lgUDEJwFBmLTNRMapVmB035Uk7npzWe/NTbOnM0
wzmcfFCxd2e01Ttf3Yv/q4o6/lZg7HlUwNZCP5z3ItzIKtJqHNVofTwH4vyRhJyLlnrLKtt3/21W
bx4M0G+CbQvmfe3uLTiHZ9sCzIYg3oYLqLlc8Isy/ynwfWBxmjwS3WdpSKCmr6A5yg/8Hg3J+BRh
CbX6tv579peWhkb/vErOmN6DGTRCc3m4rFbFieen/a2HKyVF1uIq4AdSpSF55FZQj5LEKH7OB9jU
La9//As4YuzXNJSXOnPtaOy30rOsjdvihyA2In7Bf5iSZykjCF7YFHeeeATD/2wwYAVct6dIFIN0
p5kl1cafNq3hi8AyHa2WKGWr+kkxhpYqKX/yVEsNfmYBTXkSJ2DMfHZM2ttJmmgbm01L9NqohAEX
2slgxGHoPnyCCBj4wYk5Cf6PJkur3JsUdkKy+4Q5tqtUP2MoskTO+sij6M6kzcIcgVrbAX6kOefg
F0FoPJiFlglLoIqZufTi7UxVBWTWn7kss4/2Ug58TKdIsqzXHF64xZ/AbOlCJiFZDnHj+e023jFO
j+c7UThKc6QVUjW6OBfOht8rDOrJoLJVlfJxMHj2VQyCkve18yclvNbQI2PpiVMV8PjrFVWwZ0cC
0iwlSbVczy0i8mTu+zFRXbRpre2Ao9V2n6sQI2rphEJlpJeLVlHu8z8LZ/Hj3d52A8Ptc6efG2ZB
I5f/UZ0YoJ5klC7LWFxn9hmUCyEmdaBmiEeb1tX/KQVxz4YEkyv8p67jxPG1Cw7qQ7mDKPmmgHdX
gVgp7XquNNvJeevtQdObUehXrEuIQRJW0YrWa6HO9ugQI3dzk+grE8j6aa8W4gYjhwG6A2/EOF9H
t46MlVCvVOLucB4F2bD+ZFtFFz3SEdqP27MfjgJ5sxQPf8A58r6LT6EQ6cX3kK/AqWcnEd6/QUSa
ZXaNf5sClnH1czQbVi2ueTMexDbvxMs7YDsjYly2HdAQBECCQ5rkb/vlmGSnme1n4ys38w/1kwtu
BZc2tBWOKqgFW3obpYDg0su+3Rc+znFrXxk8lxRLvWTnSuOE0Wh/7OYpoSqJKK3dDypB9aL96Wsg
sS8BlDqZKPzTXMXr7vI48EzvKRzPgcVlUZyoZKOMuybL2Ge7LPrBitzjm+Nc+YRorrHOICWiggsA
kzNX96nT5v9KhDxa6G4kewqLAezem6LJcFHkWk4JhaFNhtjgQu2cAf0AhDbUo0y2vqvbCEcZTwN0
pLgOi/SC8LHF4tfugDdaSz7j217SS8041683DrzEaoFMnlsgFSPuSfWraS8ONr+iZtcMIEMofmMQ
1M5jNSMQtvizXxyuNHLhJCMRN2pyP8zEtrqLcxPow5P+RDmwgeL7nysUikIC+DTny+1b9sdLlyJY
xwzgEzySDm+I7IANJmw+lzB9NcACkB6FyswKckSJZEAY+U9h0tJfSr/udOmSbLOh7Ct7nHEf+MkC
1xKmOelX3rFB01a9DQQwiWpFenRoxkixaxQC0QCQdFfdVBYaFZCdnY4+JFzFgx4ZQL1e/g4sCrqI
4gqMnoCaAoYnurQAl5nXkcxKPc8p61OxSMo2H7aGWVwfwY9CPKzl2ChPFjiQSUo4L+KIATbmrqNv
0sxdZWt9VO41OH+TwIgLw1KwuDunjQYgTfQShSZkfguVguhSidKDznh9WHAYx0MsiJP28Hi5pI8/
7fpjMDQlZVT9ZmF6sSZi5jN4a0+IhR6QDGxgzeuC3fuB0tvhmtWm0tXUPxZSZk5KZw5rsT/N8uO8
dJ6vG2ug1EP68ayiDLyksOwcEyrTEZXtYbfnPzJ0i0294rcJ802FV6rUSpD5kh8oRI6178PK9Ke7
qZQb83Iy8F7QsfFV554/Yp/SYg1OzvuUoNv4g7kdLudm+l3N+OJFhJt7RzvvNnnbGCjPLsCzNSx0
+Co5JeczQhrgnYOQLneGI1VMwDFS7HS6b67MqD0qrrbNozzPeJ5XAKJQ6GFZm9xJHh2kPIM30cdr
HAKdPxovIp/D4hiZqCnzWPaJxH/7N8msFHYhIpk2c8SXQOQ275u+LIpv40Yq5NaDgTVc0XYCWGxB
d1rCmWjJV1OfZJpRkFKI2R0iDMh0VTGPOPhOt99tGIe5NVKPbdoK970QkXW02DrVz0+Tu9q7jS5a
B/vzFNpORw53tpEda3pfDqEKBV+YuBchraGrnIjWgKChAnwBOJNudpBJWHJrWOGJ2RAgiIOBc5qJ
MIz03gq+jxv9KlVDrczoJnqelOz91P0ff3+BFg541S5QZdfPHy53GsWLUHeYeQDxJBFuPfdLM/jy
7MSxogr1x5zcQx0n+Ho7xl2hXi69BP2WlBqBvBe2inR3wH07z2651nguZ7gm0d4CzKt1WxzN4yB5
nsCvcTNHKlbxzXJcTGU9u/8QTGnyIG3Mb3xT8bs0K1uJgdCgnWRjaHtgkV8TYiXP5nL2UvLZjeTc
iq3RCtyt3Ws5U95gt/7z2iwiMw7Aidjve/21bKyw1nEBNH97vbo/ClWpg8x/BZecFEYxL5UZnMXl
hDqtMUcqehk7ZohtB/KFCbEE6u9hHPoJ1w093lJv5b++V7m90cDfI8JMBjlqvTfgfzh5y2KFyzus
o1/tHgKunVZaacSiPJC4FpOIHIH0H58S8hKdUtBmHCftpFH1MM0miYpTUfHamncI5iXGA4ODFwEi
tJPvwChld6bXy/Tg00OaoJ3amSIqr1RoCo/sHhcxlZjosLys54MJjQ2QBk3KEqhMCen/hfickDby
+T3GagqqJfcbs1MC3L5KTA/f1p85L/bsdp5Ck8DNfTubCo9gco1/OlO7OhV4GCPpzP37/uivxvJW
1Q31ehPM+SOvGt1MYDGJNsUpJL5II3Ik/ZML2J3sAiVRJePT1ikPHJHEcJ6x2LVs/aUdbxyNPPXf
EJReOklz5EB8EWhTmS6HlDPJg1jGIB/db3bMkiUH9eRTQDAKVnHvPCky+sZ6T2JRDbjSOZgEYPoa
7ZBzfzZZE9OVb82nEgZzRJU6oTSC1tPaKNv1sxShWggR5U+19lF4JIhPWltSq/AXpkw/eKcpym3J
gfEsycEVpTVCs9wAn9Gl7pZ2PFCQJj/L4IUJjKp8zlWERGcPCN9hLVgy/5qmNh47Ab+7PpBmvQ2D
LH7Nrh7qQwvm9/XvCLxRKJ04Rk2/3AfPkPLGr2mtTRku3SK6WbEYvKGBjfG07XrOO+FTSxeZu6Gb
zEqrHVG6yzZdi1Id61Yrrb1H2hjzqXtbZBciTaf8RKTY/RPCFZ3moTDzB8+JJK9DDl65GWFylNjw
ZD5AGhnyKEpcXQDJAy65od3wkmZjvba4gVNe2llmn6zVrSlH4IOwKisE6GZKXcqYSUSpxJAb9RxD
5nWJMstJTkj0EhyQxBRtXgwDHGS5Mfv3xSoDItgytbmzMCNI5JFD1N7mSYXKqVJhvYLj6ZAzlC5n
6TJVxHYtfpUI2ptc6P/Keb2YU4CWjgoj15/JltxNezEIkFvB+r64YTV7znKeJuFtQVZL960GV4Cl
HRWQ/cU7DvyYzeO+4ay5FPPmB0d/8nmcJ1dvD7XuA+Es6BekID6G7BYJlQuqsoRM64Ibpz2H/jW4
TBLUETPsi8IpnQ3y1MoKNNTelNRKOHP2RrCoMOuDYXKzSZyO03BWBRjpDsAa9LjlGTDSXK9T+U9X
cDnRs6AyfV+XPc0RlmRZRc1vRpJo0on6ynplbxs09iNDUyb6fRyhsK4XREsYyFtf74T3SIhEoKgY
+BewoYDD/rYCU9JPG9k05bauitcSa7uClaGc+bk9/xUH7HWHgfn/d5muuLduLwdHae4NpMoil82N
yZG2Wup4kg3pLRaWUSPsJ2B/uk7s/h//b1XiqqMVc4odTpImGpHqDibNU4RimGpdyvRPIihfVZ1S
nj60dUZ4jpCDivcVmCOpXMnllbNztq3I1OBJvuWAfBDM/Wu9KalqQpAgIUt4UcIRz//6vjY9oWW0
BkM210B4LM9kiGHV/RGa54AScSIHBo9QlGk9kJEDDnqBlFLyD7HDe+jP5dQ6RqEHUkUe1mXdQ5T2
PAuIuo+8A25+UJ2O9rTdIqSQtMuuSxEdI8Yw2wCdmSHsPgRSr4a7uOzEOhHvvNE8/AQpfWP/0O4z
RGkt82+Sfwv5WbnDHutljwf+exUDadJbTVD+BMB2JXR4EEuSeZ1O6JIPg2ToaHfiEKAZ7/XfPuuV
1sZ1Zgh2xw7dPaJTG+MrEnNYruOSnPX5mkhJ4aCRbKIabgT7WtRnjCBDbqh3v0ID+UspnQQK52Zy
d0ym978m06fF9Rdc0o+HZZWt7A3DwTdrhFAM3puYrKejMS4CPfqf+8tCN/6vrSsm4U/wIK4eR0ET
IkOIBS/nU0NNNwSZOQjqpfavF/tEOUpQLJAXaIR1sOZ6K9GIf59CDOLP5vzI5B5L8yec3DTKN3Q8
g+PIEevp/U8/6OONw8nvHX3ceDDFX+HIsYHBayhRbHoFgaJwWUbmRVCxQy/T3Z2ARHECXGRotmM4
WYA2jniDlyIYU9sNDO18/IIbsBXJbTTjmANqmooR4LItJPERPBJXy9uCTJ6Jp0IA80YP6F1930/V
5BrqpAwqBxDm3LCnt4RHEdN5sFDVVqIk03Nz+bY9EhhzMhO9f203/MkoefP5/Iw5+ks9Rt24FVId
M8/qtFDpZrf2Flk2PBPtl+5RnnLf/7/7j5oRG5URsAITHDwL8JKJWaXDfTbvKNsYkkKblJZBMq5u
C8EuatflcqWFC2r1HT93Jy5G5zqO0N1QNSBXcAsNJfMltI1Pw7btfbiYQj02iTCmHeykehGs7j3z
+y/IaVOyChBz9zYEYB5z331qY7d8u97dyCURGsv/TeKuqx7svIeyVrhN4oNxn3JYYO3NpR2wwoUG
nhSa6hJLCwt347e8QXXIF7SsvC/eL2KKWTL44FAbtOagNkBW+9i5AC0QCl1mjV4+8xJ2RH+sl07A
U+tHm6rlKL18Y+50mRFiIiqg5EHv+7VoO8sdknoqtNNb+MC2XgTI/mZbDICooV+8zLgofZzINff3
nPG9qi5qzbQHjcF7o0P46rk8so5Z3g5xqTFNX8yQhVG/XdLGXGr961sI4lZwFg/OI6kXRn11UZli
3MURChoDmOtETcEwqQwYmW9KNABY9QfgyscVPhk+iC7vBxjURsT3K3xjbltTdBEPdSnHEy9/9Mtq
tLAiFYVxgxM7pnEHBFiMYKgmdBl8WUqYpepRLjrcJsurz+a+/PGdc1FdU14bfXQ8YTGhotVugeAV
2Kdfx3dQZpNCPxHlHu3T+qeJQbRZGPT4btP2eIBVpPNgjjvHVNmyqazi9kcedMvMUGqdPC5xEtmo
UJNq284+w+GVZHBZ1v2NTj2yWfJoXeanRDdZDRwexoZDbpPunNxjNS1UtSh3jczCr2kBiSa/5o4l
1FRipN7diyjE2g3HRIGUCiylMCApsGxGr4WHPqFNk0y+9oyx+DMFc5o/0iiDnV1dL5KppnzaoIC2
kW9j1fJxQPcBzWiPW7CifqG06RgVs+SzGrsDxQlYKgFahUmL5RYREq0XHM4Z6xShve6A1iKauYY3
/zMUkZANcm8oXzUTxFwy74LId2Hy5yRAHTuI64+bm7qr+artUD9Zb8OlA5znGdFfaQBP+lHqwfGU
9mo7R7qb0RA1kTDEmVKBPNC/STkSID5HUjkn9a80E0HIsLsn1HPl9BQYg1+6ulws1b5daJV1TLBa
EpoR0Dxi3HAAWOWhuWgVVooNTNYt1IhPJgGbYi+vLEVJcrQI8k3H9CbagZs7IO3El5+Xk8YMB+90
zzam2UhESK1frNydnfIArIFk3syb4V5Ku4P2cK7DkZtw0WVqjgEV167i6Q2VA5CPCt/XJ2yBNEjK
kYJM7GHQ6ymfTI4qs9coVmPJtd3PXtH6OnSPrTzaAJtxnFS5bEOIBEmIGAIGqQHqcq3Luz8m6DlF
88Sm4pqgCoYkggdxHKWIRCWzSERDSiVbDAbn/plITsyNaD90Ej/++v7jb/x8PBJ6TMC4GflrCse+
WivXuKZtWhW4gpoHruXq8ThufPkJbqCDVVmNI6eGNBFj2eyALs8cy7a9MPurnSScBv/p8JpkPQqP
1N+hdv2NmRi2IibzLdd8FI5HAVoITopCTyRjiN/X+tg0K5ZYiNbD4jZq2CSEjl6BFm78RoKT5owU
hl8VuV5iKr1SxDRlLNFMxhgy/oG29FMEXNW5GbpuhaNMrhI7dZvBSwpFGFAHXEiQnTJT3sDj7VK7
u2Q8qt6Ug7sxeHc2RkDK+yZrUA5/iJf7qcoO6xvYN9RrHsAZ3+HVLMB97r9rGnppeYmTZoOje2nd
OCF7pRRt5SSPeptjJiaSMNbK/yXZUSZT8I1VqWJ7coizYtKFGCA4t+GRx2hr00OCOhy3cJkI8VO4
DgJP/fgD0JZHrOIQA4uGQUEO20hx6A15oQT1Zw5TAAACp//3+9p5jSHeSWEv6YHawKSk699ZxCQL
hlyrxB3k2aACp/kn3ZTA7ORKIf//n9O2sP3PHobCWOZxI2XwwXAYD5X8Zp2vlT0N67ooiDQd1lg4
Ce1eMk/NcOtIUan2qfT8J4nKidIdoNScXNG4wIqqAYZgA6N0722IfMammswhKujO6xEd5HLErkUC
oyn8hsQx8yDqn/9wbqZSXBW6RbZ+woDE96UHLPrQCJXaZZPqhx2zhhGxWtyTVRudlLgZJwq/ORt7
4WoJUBqQegohrD7sBcnSzLqKqzEtyaeiuGz/MiWp23t+8Cc6KNz9+7sxjZnNzw6MqEdzOu9Te4Eh
RLW7T6oochBI9ofj1ceHSZ9IpOJQC8tSYgg34ijT7NXsrigqmMpV2zNx9vcuhvJC2g5iqwCKll/D
o6AMrk7i3bJOVhXjT03K9+z2U89Pr5v2r7XFpSkSPTML2ZK1NFq1w1MvNO/jYeo9f3LUaQfwLuYy
cNWCjF4zoHbvxyuINE1j5ESSn5VX3oZ3ywzic+2lvH5RJTasPINSFFVp7rsZj/Pj0w909sJXl8nn
Z6EXbp70ILcX4zoVRXw8bzHu1cubVyd+LKiP2Iluzfemt0NisVXRVwqczpteVE7PbWdtDCAa9wd1
aptsL1hXaK4o3tPQgGfV7CgupLVUHn1EcCE8Hfj5+SsDiGvZvPywWKNk/pR4BCyYLbS5R5/BPNeq
vlhDpWWmct93jXrkHMQRLv4edunU5X06N821heDkRDycqZU3BAa67Z99vyQP/2SxrBMkrHJTV4kh
G37PaDCR0CgEEMsshHOkcns2hdn/0htoKGIinEcAC7aesYmSWMdHKkNWYA/pYgQQhmWr+Rb3kMTj
U/hIH5nO7Wjwkc0mSX5aR16Bz1Okr9NYUb655CfLXIE5ugw/BaQu7mQGlCh6HrXmf8UZLO/9ad6c
HMbSpagFa/RpJkfQUooGei6mlIBC2eTfZZqWdoc0bn/V0ujTyCS2v8uHVkpk1IyDqWLsqd9s4bAq
n8xWYXPRXHnwcBDPAm+5Tpu38kQ0AtpcRATGJLB4pQV2fYQYZm+Ori2gGC13/jNdt/Bhby5skO0E
7NoD6XP1J9VdP1rPGJyj5pNHgJsVEW6mYqV7yV3n1fSDKf2+JmvYYy55T+VWUeZVAtlw0aZk9LAE
hubDZANhRVnrHj99Q122nhnDRf2IdaZMnK4r0KYuJCMZrpAManyVhaUjqt28KK9eu/0kJUFfECds
og+QLq/MEJm22zXnmoat5h5agcOEw2KJpvG5OUY4xoWpj63iwfs5GLpp/DIecQYiWDyc+RK/RcYf
W3rqK/sfb2EI9jVAcgmt+m/NEIyNfPxfvgWCNkZfMZQdWFFtBBauVKtL4eOSTU6cMH9RUSXnzoDD
Ajglpn1Zo3zJiJMIdMyRAhPWecV8LIZPB5FWCgoppkxpvjptr5sf8wCMiCv9D3u2AGa/e6ntxTb6
H4OiasnQAzL5ldbZkxEBRmXHTaQRvKRIMNHXt5loaIEmvxI+wwSxY6DjC5KQLfPSW+Hf7AJq1kUZ
YL5t/DpnF5VEQ5DNoEr/5U+C7CkT9y8a88n4FGXEpcdjupBghGBBzRdDl0BSgIBGK8yur3SEJ+IC
/9tCxVB/OGb4lbEb4i6l6jQC01z79HfJSIUGTD4Ca14JceV/B4P55HJdBqUJ14JqVrbmUX7fviBy
Rekgouuu06IrFVn/XITGMJ1FUTMPwDEZxHQrhOPjeEZ2HnC48oP6e1CXiPJ3z5e71/eUowQpplzs
lElXfhOJKzsBenD+u6Yz0gSjtMaMW73mqwVeCrC64SzWhoo0rmPJt2O9LRGlvC2lp3yt+umZV3gr
H7T0YNBO+lC6IEX2+bEfUUa3wxi60ZGbNo8FeOM09lxrSEhF0s1QgsH73641D3GJbhflijMtDm9e
+OyLOuMg0OaCEQXOCNZbQ55c9bZ2ZzknKQI9aEgzx8mUXIOoie4OASuSe/HSgR0jbDioeS3Ql+ta
X3zwRLPI/TyY5vIxhHYXcy6kZv1K0SALcslqYd22YP999S4F96E9iVZoSpgB3zN87iek5t2S14wY
icyC64AfBdlR3XPc8Igxsng9+/5YwwkLdl6SDEjjIBxFmu+ffZaOIfn0zHKehH5z/m1Z33zimruk
3agQVMmuotRyYvODAVmAs9vCgMs83p5rtoqXXueMcgSQ/y76gRYzkG6dwamcstWS6wHSGETTGYvJ
XYwytrsA9aLxYcP8fd0pIp0j9X1eN8juZsD/2nULlPDy8QlWKqjbpUtfxe49HsjanTwmup5+DXIj
T11fIrkpyIMwoJPG3yJulmJQq/AZ9xa6Ao6aqij8263tWrkmreSpzun20lTw/mPQo6pw8jwsVEHC
rdnmW5OMiaQjuuzy9/Q7wkNmf+8ID3E2BmpeywaXvyKfyFyHkl3X/Y6nOAbCQrsM++GwEA16+2KI
5Cc5X4vBf5uXaoDzH2hzk0qrPerDM6xhf+sWi4M+MOMB3ndan0/0tVAAmNTOixvcpHK9X0UPPNs9
G1pYCe5u7uQtp9qwm4NbB2AZed7DtfY/CKH0XuhNOqtdG/GfZ8qUxjuNVQdvJZwWIZ16TNzkRJjn
3tGeVsk4iPlauhbq9eAmLHMYLBzc8EfTg5RRL3ZELb5bDoZTvt7zLcDr726/Jox71Z6x6gF5fMf+
D44eNI5qabxv8ZMs5J+HqicL5bNNzTDL2HxoApbQQeQb8nbJ7NOXeuWNhmW+wrqBH+j20U/3rfq+
D8IWK7kbuRttE4wgw/UafkfyH/eTAO3Dio3X7aeJPXez5SjQotKr2JY9a1HUTf0UXG25rU28NsM/
N7cVGrqfNomvKOB5rlaDc3usZohwRkPjWKqTE/s929Pi/mgbwvWCTKRGjJtEHRJKcyx7CuJf4YJ6
zJjUFYg9xBF1CKKf/d3v0Oq/brrRpy9AuK1EHfnpuUSsJruphwBbal1M7puXXuu2ioTYOUgHI1zT
+5D9AS9yNnXKtWdHzAo1qzpELtPRCbsJvtu5DSW2BWjpruJiSu+LikLt/zxaTfk82+z/NDBr8x7a
O6QBoe1/65tE25DpNsA+s8poFhadKs33EooLdTk6Yp9XMRV5DIrvcVmBg+zZ9Vm3xqD70N+A4mp2
dq7uEV41xltE2rfHvMMtD72egbCJwfhHAHwwQlYfOOP+rBiRq9bYoy+a2344hoNMl+NHlYWdQFYy
bD4riy7SYjFSB+JwtCEIML3l5nSwnflL90FLibQun1T2+LOk7dnEDmXr1W8dpuwVy4QUVF9aqSk8
tQilIimASWBGk3vhfOfGOWFqdtCzpTKGBlCO3/DGaMXnz4CFJeMa+U77g5xsOsfyiOmEecMVuoIL
9dipaRr4ucuQ/orSBB2deQ2Hl26E1NDu7Es0PmzkEfeLyUHq55CEInGkMl8azAd9lpdioHBWTcr+
kYOxKRYYDxILdKl0nEfsoOypfmZjdpA2NTPvDyJqKjK/1YnemGCdJp1cLwByZ7p1fhgoj8U4g9bX
5ABkJiBARWZqmNKl65+fa3DiZqhHapOZh6BDjXHErNa642Aujg7jxd3bel2UBUBgomlx+/Ea4ac8
kkH+fBP5XcTSJH0/CFGq2ie4YaKButaP+1UXRzLOdf9KTMPJ5nftYRpQ48YbXYMujkkefaN9hyfS
yBv/q+tbOJI4+TqHowQQd4NvBg6TeqV8GYz1Tkhz2sd5ZYJq09zBB09f3guF0AXiAsnfpvabyQYb
THcFnLz7NMz3MIYEyf6BElLL0kPw6VBFaYhcowcQR3pW032ZXbz92xk4C8YaSid5fphVLx2Fdoqu
U91s2n9m5Wg2RUqCrY3Yr5NJf/X7DVXJu5r21JTm96P7oyUOPga5VmUIAabxYzSiXLcTVQVVzlfi
rkBBrutKXk424RJIvVJzv8Wh0A4qU4HSi3i+WOimDixKL79hIIrt8rWSypJwgmECe3b9Laqva4j4
H7DAKpgcHGtFHxTBG86gerRJn47f7jJm5J7AzdhN+DX0Hnf90YBBRUGmfY5jERcD+kv88guhPwuh
PMJrvYsBNi+Ul5bqRGGU2qTXFbrxPtBMq7TTa+1XbfMNpFV2BEHloSE9ys1I+/SMGXDPu7i21sFp
plnIv78fTObQbCFVjXgTqrGH/+ewoyyincQnuhStMqMuORRaZSUu/F7zwy98SiGXp46cQr+CCkk2
7x3l87PakS3en0BCxAQWgWMZUVnSyILbDBkFWsxMHDxbou7TzpeJoqjm49FD1SEb6p35mNt2UOAk
L2OhM2XwmzjNKdxy4yczzi69v9ftP3cjSFoXtfS4F9X+a50Gb4EueBoETW6uI7SzmyWywcXSId+g
fgRbMuvuMj6g0zuXUM6Jl6+a6hORE7OvIZELZ6GrJzmUm7Cf82UC31sKU6fTnF8fDjSpuMJIp25v
SckXnj63YsP9HHLND46OZSGJEtpPf4uqwiLGwVsNeIKqNDVETj3zO2y1pLFWd3VsWa+7MitbLtUi
uKL6qG7LGbCVJz3DMn2u7n0JcjeQRg6Qdb69tSiOaf4tK/RtuiLkAt/uhbXbriLgKWE8qDm8LIfq
F+vE+cgPFjDCygci0Jr2pFRYylrZ3AYhH3QLwmkiSK64dGJLGdgYB1sG7RtcrsPxtUG1kVh5j50p
LhwyxiLo4z2yl2EGngtqpA0D8Dm68usnT/cjYWjQysK7Nn+aFgqPoylOk/GFTP/CuaW8ZmbO46Lf
0RWbvP1h8g3z6zaVkMA6pbckVn4Et7mnUzjfXXJiMa2xyZ1AaVKe8gC580BHEPVa6gIWxV1gFrvw
+PeDU1g++Zy/TswCluPp8YNK0qLE+G5rApwpuwWJkWf/amyomS6eQmJfDcxX4J0qjJRqofN70glT
ST6vXQLAUhpRr5ApAaq9bohb0kYdod7u6BN9iud2lR+aPgxKVM1yA2b7jX7PNy+qwnwz8faGlR+N
3LjWg2TsLzEZVoZqKSvxpxU0Y8KJd2jOnzY9WJeBbTJHsYM0hcJGF2LWF6tvoXzpsNPE2kKjPWBE
qcTpi50IizJTOtD9Jhthd4hu1qk/fv5rbEvcE+bqftvFe3G1Kdgh2wNue86vC382P6UtvbQ8Q8Qh
/kspsfaCHH7/y0/9YAvVm5KN3xReGwu+HJBJijJrpLAgHZG5km8Mhj5tTj7uCDvqDn7sgpEyGMqU
lMl8+EWdVJWzEXjArnycGPhqkBOSvgkn2VcI+AXTeznxR14tKRG8D5eLz4JfLM7jSIDS0GMG/zhb
pMs1hHuj06QICnK9mQ9uY7g6ENVQ6Cy/hOEhlDJhP4cv5z8p6BAylNQZrk8OEIfM/Ap1QvqRQv3M
S842Hhvqsks6pP7a/+A3BRs+PyzEfRJC5j06dcwAX2OylkRO2LwBaLHZWOOQUwLPfZmyNAAixncB
dDDTLwwTazdGPH1ZTnx+HAt5XAqzeo19lPRXJEoRkJAs5KlXo6h08HJQtqKR3A78ZNh1klYImEC0
3876htRXYbT9uqfiVZklSWV++DwfrPgHNVWtJWp9/vzyEco7AK5C3VMIdIIVR41e4wIN7YUWeNk2
z+hHzwXSWKfR12tQKAd+B+uyln1GsJV1zgQe9nQFt7G+uFfvwxsdu60KjELSPWjD1r2Hn8+RFvP8
v/1c9C6WGzo4+d0F8bQtqpC70GBnZbRHpQ+nGQUycWODzcqswAQx3Z3u4L/IX4oCbDtTelFV3E27
IppWT6XxnwS1/1SjJ6ISzD7LUGUElZmmFMbHMQcxdqem8pAKPfmUPuiub7fDSRA4J/6S1ndpyYGI
Mp3A8phSgOPo++xBuFSiwZa0LoB7prt0hrQjwFF0U9bmxT3YRHpfbdAoUvEpwBYinKKZtP/UgmrA
993caa497MlcSJ2MdyHlWwoN3W3Vvni2Ghe5CfiApaXV1Y8Gqml4leOrqYFDlQzav4C4PEsTcAhi
+0vjWmKB2a/6rjv60+kC/IZhwXnGjvOxecEZn8y6SdTta5A0Q63eLQA+v9u2SQMYDnY1bXcHsi7w
HwvE67l7W+clyIVn6fLUarg9ZofbUlCcJZKOidL9IIq6v4bCWXwbssR0Td6RnalF+5iEmn5YxuF4
8SNaaJ6LNGWGbxrVsiryrpAVOsNFo107nvRn/9K/111qVKhq+CDhfq+cri1QwhVKh3+gZOiNopEO
IZTdNgS9qZHx7vH4AIKo4hVs1BRIbOLGtX5y/VKZdFqFiYO8MH9015kdMS3qzR31226o9jaLqSI9
JSL8Md3qtbKPCeNJZxxqeZYgTlI7c/w9UDJa5lLLzdeoQbOjca9zPB+9iGoyHhvxaI8ssFwApd7L
ehaWfw6MJawjww/gx1btd+A5kfiE/m02swr9f6NTwE8sz4toFnvz8wOffSiSB6HH/Os/55Nn9N0y
9/ZU+oVjTZ5x7d5I/uXIk6/vPnm6QIlm6sco1UdvuVqdUr/UZqv9/cXzCMRv/jaWUzPIbST6I2pY
XRFJd7MKgKvFZvFU3ME1cu98T/mPRYV3o3N069ls6aCqx1+5ttH+8dRIUl7u9+XfzlphmHLNrazV
cBAVIrWhhr99NvsW333RHBGUujES9wul6ODWYrY4XNlzPqZOH93M0Y7/yXYjGkWR0q0yJn0M/A7B
6cp8usrcAoAyeFqmkhqNBWRCeDlbQcDJ/yKHkFiC8wxa4qnv1UI8J+YVUMEt0cSVmLRdcIxjFzn2
8c3gFMUdpAc7yEj7a+1fFPvXDe3uOZYMxQMcqJzc0tzySA8gc9MZN4H9wf0q2l9gBZjcdThgj+ux
bWZJNHPoaqbVyeKePQePTKtYDXQrQIOmd++Y8wdMXAxisJ4jnXl3Sq0fPaqChcXYxTbWwtk+Y1y4
K0e1zTQ/k/ZPsgX2gwjV96itfoeJY50ezqJw1WvJ37IluLuwdnBrB35f44NZlGX3CouVkPl4WCmB
0PioQyxofZlHnPwvOSe4nQNh2CbbBXpEj+jx80emOjixKHX2q8tnjboIDbwQboDxlsS0n3oeoBQR
wZPWD9MhKhGcme2fhvDvv0Sda26a1Gb5MwiwSQyjnRP1zO35apHTfJ8BaK5hpRJwTaRMYu4EdVcv
TXWvtGe9ZiVvnDO3ZHVeq/h2c81ul8SjyfrMkD/qKpyxlSd6J7R++7bi98O1QWQ4Yc9fwwkBjs2+
l7LVLKWd3UeiHwWf6hXk5Zccxo9T/svExCY8+gZNFd9P+V5PQR4sNE6AZD02iJKPKOjdJPPD/2f5
ntzpbKig3Rv1b8ovUYDPjIeX8CUtW+Df97hXDCzGy1e9yPGe68QHw2hIUhd35E2MLbMhB/8mMKKs
XLM8nekURQxmH98BeXbUxKgUHs7R2G38eV5xbWnmi4TDiQLksVJLTaWT4CQ1/4qm2QPz5WRCqtHl
bqbNrbEofTK0iPGveWYedHcZ48FG+kE5lZ6AD+Jh0GJNhAJ+tWoR1VVcS7WnhQKv9TR6Bc0zkjqj
fXxXfwawt4L/JJJuDZPqRIM3WP7+JpE1cMoDHnog7c6oYLSsP9Hqf9oF7NR8WKm+j/xRbCH8BMee
kIppkHD7dv9aTZmniiO1QvG3mHpWDbf0WuzLgNPhufeWAZFX6Zke0MhjFRCIcVqS6G4X/Dwu1v3d
/f6p0s3KOTnDIPlCk8Tlf2EYdPnNJPypQ8HRQ/1zn7mkvIWjHuJ+EZH8xr07cEg8YljI7y9oWEH/
8NPkgv+MLFbXOr8lslAMFtJvfw89fzZObUeQsCTIGhXHTMv22m1bwyF19yUD24Vz0EfnrpkaFslO
RspPIyZJEEFAO5tMdtt1mshvbBlruM2sGi7j4bl0mKMwT0DlM+MO+v3vj9ODwh5eHBuTA373ADmt
XDZ7zQDj8LYnHftroF4kB1Ie8v9lwWtXeEtbv0HPg1swxFC0FMybGsPbiwFGAeKwE1pCqSxU+UQF
kF8chsXgSDw4/p7kxOwZ7X7Ft4Iu3hA2zr7DM3NPTUTjZHZE0E6ksX8rgy+MFrJRNn7AX1/9l31p
RmPzoD5URakYFfWn2sraJOVgjij0GMbGiCpQvhUpvOPPAN7pIgj+5m5adDjPDTazf4zHK47eanO/
ABpr5ggI6lin38p0TBBGE4+U7SyeIcHnvWO2/gb2jnfqDo5+NxKNu/2xMnnQGRBlKGehWwsmkl/r
bBjVK7ckFCld5sqOJv8Jy7jwviaflXsSfO4H+MAp64RHQWgXlQ/FSiWEm3HNdnOre8ou+9gjwhyC
roT12tSvlhOR40MNZ1yaNgRWZXqb4aTJ61hfG7b7ONYN1z6KdXv26+jR2rgf1N5KkIfRXVwz+W+k
HeeH1vakcZEJiobaU2rUmA+zZoVbsk8ZUZgXNcbCsDzb3ZEIgb7/8xFqUh4HNEyk25tE3F/EyOja
m3QA9LKHYDZ41yoybry6pXsXdyNH/NUQPGz1k6qVf7QHKSX505yrMt4b2PGBDPB+tgW6GVBk/E+4
WqnjiAWoVXe2cUc5M6WK7tuFr5KWlataJOYhfSH8Kds/6RyJEJ4LJEuyj/3aLxM62+YMROEzEh2G
ElhehYKAvsTSYpcNKGGOzfih9UrRK5kJB4FoCMDjtvAih2erPCq1G4X87RLSGepFE9KqTbEw6orI
PArMYpsmsQj5g/9OFy+vcrTMA8O0iOQtnhd4pCs9Umw1/edh8cbZhXV8AAPFgY5ItCoNHALyLCbT
4QYtQTXZlVO3RXOO4FrWt3q8v4jvkQJj38G8d+fc6ZF4l/ChK0mUkpdHn8THe7GtbEi8mnwDEBB6
UakQpW1hjUmGfUuJh9DjFMLgz7nW1nYIBrQkGULirqAvkQ0164+F5qJzrYQNuy8PsTyUL40baTHC
exlWw7Iqndk4ksYkRFD5ZamA/WJEJkGkqkIuoCtsD6uG+Nf8ad0T0CvuJyY75qNpK1pvEzsHOzPI
8/oEoMlrBC8pJDpJABDOvs421n6gHkAjL2g6qwQJSzothF06F+m6Rd9nvhJHvJ0pTi8GAnn/cLvt
L0I5NJGiC+zBOlpnYebZQNcgoiSCHdx9dzt8OXKbpaI8SOcPsZYVC1VAlrb18MhfSOwPDdG4b6z6
wyo6cZsuiyE5SzsLaHqRtvXuI8uErikK5h/o61GN/pWCFMfHsKWYRTw9z1IE2Re4/RZzLzG0NEgU
mtH/GEdnk/m98HW7CS2PZWN206hYLGuWnIlqbtV4Ob8U8wmns6LpN5JwRcGkS5tzxejjFmKH04q8
ZGiCkQyq9c4rofNvRzIgx8M3JnuxUnevfT3+GuczGpOGHxz/gICg120tn2B24qiyVoBkIsXueXVh
oH2Z69gcLQ9qmbReyb7V8uV/Xo7Ro/Z+/SgSI+SqYXc7b34R3g7R6TCm2qbnVpKDPDn8FkgbH3oW
lCBDrB2xPIXHGpXAX1tUxdKvLRhSazulDbZZo5aHUC88LH4UHeSphm+MPWuLHPEk7DoezXjjou55
dZ8p6mPAZG+0/Hu9kr6GCnVtaEzBhoo3O6UrMVQgejxIlpGwijJrhhsl24vndZz8KgpjWxB5pwn0
XoGxw4tvyGxunnG/H82Ir8hf0/FplB4V9zHKrVRTeRtvONN/9lk9hbeEbd/tt4W+MsQy/sEny4P5
I3E2uuOS8baE/nkWckQDGAQVpZGBfgqpyGzbTW3dEV+JOx2jsEYJtSUU40p7SEOlAzOTA4AlLYRK
VPa8ZXAO0mbnGcn7wZcot+oCV0MV8/7x8oqsTz3eE9jzw+5dEeaPWLOtd3YQYqLXfUoMw+xKqs6L
u8c7PkSxamue0LHDQSRNcnbxi0BL/oA7no+DkMeQKepxm/goX88irp49QBjRLB3PUED6hZq682PW
Y15/Q0w7qwiXb7k2GxBdhSCABezI96sdpiK3u/wFi4xQo4OBGw4APawjr04G+DJmyu1Adj1RPTZ5
gV0k9g9fdBaxJR8roRfsSda8Dthmu2C9uGHjJJkllCriJoExUULfqEXuVJMoFdxIj3iDSPmsF8bt
AcZf3U8hzDoZ2Qt9solBOyvDv8a15+6+Lup4qacLlJWYQkaKv05EP8OodI7/7slAkkaH2SPai2fD
wldgHVzZn6CykSGVblXNWThinMtWS/942cGOLC1vCsKIVpYenlJt9rLXpoq2GBbMB31pc6j993QF
lxsM0hK+Kwd6ewZgtyXPSs+GnpcaNQFZ1wwC6/XPPlbtw/l1CfEuw3A0HA9/t5UZPhttz4VWNNQN
Z89SXjDYAsGIxMQeB/A4EZGGwHshwZS1VVjvdB7anHm3Oltmz1DWfaSyS7dxYQAVEZowHeqJIXBV
XS2/HppAu6KyU016edYxzY+T2XMarN0Njuri5kHh4ukqHbbrQ5Hq89LSd9ZthIEypc3qCn0+Nl6N
Q4BbKjPjSF1GrQTuS6QsIcScgn3h6k1v5EdLC378Pn3VtXjOHxP7LHsxEVaCNMqSrYp7BejkQ8Ys
KRaXf/SE7eyfbjVADu+dMeQvMVsuX5RxqVBX01rumELesvQlPL0BG4SMYrsdraGc9Udy7Rr9ZD3V
6HOIz16zUOwI1SI0uBGyUNup5kkPTXmIaVZ4PPNrM2LxWGmrVTnw/S4sQzS07w4vwNUYQB+QeV5Q
LK/l/QCzqSyQceI7vAm36SXi3opNGJA5Phq4syofPObRdyvWRPOeWTf9uWi867FBik+OWw+dXGYz
Ujn2aJJ5S5T5VCgBeFN+2k1Uo4EPqOQoTZXGDT27YkXZb176/SM+3jRPcNN1Ou/3Qx9lqnOePWzh
jTT3PvSb5Wl7SoiE1NmlS8rRTqPt1dJaX9f437VJUSHpciv1dJ/RFu6nZUWirRPuhb3JLgQVtoe2
Md/1ZFoHVApG283S286cPe9SEJXUzge8trp1XVZ4wobhnn1SNNsw/72rVPwL6OJ8Itu2P0V7Y5zj
pE7z36qPrvQZxAERjtqNVDddiaIBruktH3k8Xleainu3ZWiMHvpPdnxRcHiuldsOMvGUM93GPmTk
lGyHRlgxxPIZNXmwqoxQFgeFhVe6KmzWC2DsD3eW0TcHExdaeyTpi4qZj4CqQ+6pkMhs2OLgUjtw
xcn4WXXYBfj/CgK+uzyTORyfXxCsRDhjF6eZxmb3uJlB7la+eatfVgM+pVOk7WTBgK15lIDRkFcq
ygPBxLoi6zzoAeFJ8gpA16QC0Pv9tibB7s47lgQPg546jNk0TVSMmpwIfZMT1kPZWd/8/Dq5NX1H
yyHlpoCWGpckZK4zqPbrwsm1EigHU3vLeCuH0PwJO9ZS4/vlFdFK5f2Tsx28+YyYZfYsYU28EybH
uqMKYf5KFYtJPURwet8cnu2i9cGVA51fomTaayYS+8t19K9Lpf4qmUl5h2FsKNwkFmHIAvz58khW
tatrdIGhaSeY4GWmxaMRBX7MYzTJcie+2rwyEH95QJnqovr2ddxZGkChdfGMlJYupsqBMMZyxxfq
6buYT0f6jGmkmE4vfofA189XKgroU6MMrutjyjZFEmTa2K3UYIuwoDNV8r42u4f34NOD6A/juvsi
2ls9epQH4C8XIvEwSZKXDnqAfoPxb7AfGEgyCUdUBshw/KpWG6dHaSA6bE8zIMqmtC8Ff6jPfIry
Uh/33zacIWW2cZRIJk2MNxg25Qbz/pt13YeMAVZUy4ny8rLz7FZ8fyUkWmDdV8bwGNOKwix1iMV7
lNON+F4Gav0DppeEYIaS/6wQAEyUr0L8jKOEgG5Fj83GW2QVHxbjylKRND6F9nEN/Ixxa1+14Uqg
+ByU2t6hPUMOq6x+ScVBUMkpxt/IP3BzmDq1Q1aWPUlZGYgNXxQyhRYECZ15YhFPquOJXBmDkFKC
t55rvy6pbxNUCgnCnHqMEmjF+5IO/W7wGdXqYjEYDEEnKlA4Csud40tKMJDg4VWdlO1ApYu7amAW
+F7PSOjV++5rpLYFj1F8+L855eIMFlLVNkv7BbuT+wUJNcvscUw6TMdqG5G1yfymU4DhtBzBHNsB
AsmmnP59IvAd37TiIxIUYA7mbssrRfMYlwHdLV4Uex2KRIVu978Ryd4VAOdPVgoSn4ZBYLZsba7y
wyzeHVnf+Ip8ib1AEnW1FYZYH4Zrkv1o0848xt/iqgG8XmJs81liUzzu9OBYsQdl0FPXLjG/ToVB
ht7qWDxk+omoNBrmgrc/8iIgU9icbfTK1kUz7WOAuYxLV9e8CqsKGNLKfALg+M6GHJ3RrMmYPjLz
fxHB5Zu4O9JEOxnXfEyCHEtqHQVv66Lqx8S+PT7MM5S9uTLeZ7L8fZ8BK2H9z49D4gy5CIWea5jg
zKCDMBqvVZHIoKBMbRuDxeD8yLRgHx23tabOV68UbD9OIMVU7jwXRmBxbXigEwshH+rHjEzMbHDd
GtR8HSKUnXnZtLa01spnYasT6QKBeBZP/TqYosIBwRLkqfLqlbu/IJ0jsDYpSg6PgHmNKh5rgrUk
DVo4VduCVZkKREHERl+4rn883/I/nsEXLztj14JChVHfM+mMNEblzkZuEu+JkBv67O0NhhuiPKxD
yyWnlPtNkxVwxTTWCLj5NXL/ma90P71OLPU6bewzI+/mhelvcGdCTjTHxQvX+wZEtQi6oWPsNt5i
9aGyLLSM1ZKGpA2M77294cT69puAlH+XSIqnFleHzhrphJKSZk5GXPS4mxQ9lVJl7jW0fnZDEu+m
cyR0b522E3PIZeEK5z2G6ZZldURHaKvOquqtRv2pbcCo29o4a72jzFvTBmrQmesq5doNuN5/NNUC
dfqrwqWYeXHlyvqpxFguxO5uEzqaClQfoXdFrsqYN+BHVA5hOBNEbAfe2r0B8cqDeOc9het5fXN7
aLZMqzR7doxdpn2D1OsKMH83j85GERGUUUE3YImzvvdat19B5x01HEgw+RJVgod2WMWE8y6l+NEH
/gFasdW5lNmh11K9O0EiRmBvckRdym8OW/LUDlcptNOrzaXkmEpWj3ErYBmlCGgB3CK81gWV5yhR
g0n8ohfu/MkHYghJQGzqU736nLq/QbW5g2NRBGIgZ9sUcn9vKzXc6Gf8USNBj6wMq8X3ohtATflF
VxfZW4ZKBn91BF/7NWJfRYBOa3Am9n9HB56jWnonIEl59bTgbdBp1PzcmG81w36T0u6F1BocSRk3
2FDpleuKlcfMFNXx9ruFiF+V1dIqkTNuwvgi1SOVOELXJk+jM1d3S2cjuBTpT98ZL1fGQiZxv9IN
5rdlzEVlf7xEMHgFzQqW0UmUaLhNYcAA9h13nLabh6gwmwqpoUTV98JxmfwG0PZjRm4hVIHc42Cp
Ggb1Lg1rsKTc/qDF1hKx8jjXiSV3tJUNE1rNyci/3mQi0GTBQJTVvjgmzd1/9GlYhkxA1UnYOt4z
USF3QFtoY9WCvoVe/r0obPeHXWhdPAcM+yTWKdF1CUftaioM9v5UzWgPobcHhUEllqQnuO+9LhHQ
y2hQc2G3BfOhaJL4k142fa7RJ7RuDn+1BOiXfHxS8ZV02GXiwgvcCZ6K3Iy7K6SYHS7GEFOua0wW
BkkmMbCbvETbFDtGMM245qmsCf+JYQzW+S6quJi3EO8mMtfc2YntY+jShZfCr1zEk0dXHlo3yiG8
GNEkL3m0vnpI3+L3nGOIYWzqPGCbTffcdXtRJcuzcJvTQ0o1cOWTHnX8tS3cou1ioF5EQyCyrGeW
yJLfRr/FGSE0RzlLmfeQjsrY974XbWImRxyskMy2g/y74h/nyt7izNJ9/WZZZ654pQkzyAPUu36s
hdZ4ZFEq0gLaboGLU804Y2qSleP4LYq5KMhqLaquTYMWQiLp4ajkBKXFt+o5ut0zuuZAGiX1bXJ7
jFEthmKtVGF/3/Jpnp9TMw2SWVZd5M7Us3GUSEaeIMauZp2vi5XDW3j/Xsbq8UI9Ut0/2c5sVgpB
Lh7b/UXpotZRKN6CLGp+eoLLxFMXYbjDn9ihLQJA/ehz/f8bRtYQnZwde6uxE8ygY1TOHsAtjLOA
n2tUKy3ze3UFtVkScddDK/qCpD9AkwjYiXGm0m8AE9ayBdGLs1snkTDJBewiYbU3/oHXJ78TkU8w
CYt7+2WRuGpCQOjjW5s6Tto7BoRi7hryOQzJCaAAhevlUyOSK+a8SO+0vp4L4VJhK2wicXlBZXf0
Lj+DJwNE9Nbs7Ud18CbKUxkvEoIA+PPxrwJHOTobdZ+ys3zTa752Q2RIapQvNgp6Mf6lVIa5vrn6
2YRwKKj2up1JTe7nlkSpMP6J7ApLhoMrUBdMmT95y1ip+W87ahgbNY9lTv2IZ7QGMguFESJV1mcV
f8VzOOawXGHlu1OY4SShoY//zoVZaf48otWrFROnd254PTxDyyXOl7wvY6Xa0cEUf5kspJeoCrY+
kpcHSi8hTW2QSQYXIBszMkODIkgkzbzvCmZwU4vdVvdzgnaGKNSX61yUtx0VHiMh+UDo+IIzJFaG
WLRu0NomMumArU8F4J2BBQgjOo5tKzlDdqxllGY/f83PGozvJYOgZhaURT2xV5ZpYHSsnv0bRCby
/JWF5F2IA3yffbYNEXxuJwBo4zcinQxOYawzqh83YGlTeSobNKsDsY8aTBmP5HDUMIvsxzfcqUJ6
mxkl4L6osHOzHMOcbBD7MTEefktSCuCQGu3W7JXVyv4fVeD7gbx8JIRQJIGjIdgbinRrcHq2V7hs
0KuMe3JwMRSHzqEgDXZgHKjQoywmCWdpLeR3dpiuzOB0bR2izwtuAYBVGxjHmd5+4V14A18TYe7X
L9s4BcHc/T51GJiRFPnJ+51J15k7x130xb3QHNddRs+l5QBD+GX5oWlAGNfvdfBcTWBhQe+LcMHf
B1u0SjyHvcjY4FOcv1IuEZuFJZXFNWUtFBM8KXcio/n9c17rHg7v3G3r7bceFHpLIeW1Oq0FZM9H
eQUMrQb/7vDgcN4p+tGZUG9HsDJmfLsteyYEJomjnvVe/YcgTDx5FTpmmPWKoW0ClzaYk607PQHO
Fyu9kDdw4C2q5smn8rHRv9xJFuxsNWzAhvFuYm1Pdj3MSuYZaRX3pyqLSnPEDVEKcw0Z2O42/Lw6
TO2EUsjF0dFssAzUOTfc4AxeGnvJLhHnvizB/52SZGLfa2/g0GInZWzryuMrC2xE2eZ4KJjOD4Cr
xIauTe2lSvvJB84JNUNQyEt8Ddb/tnocHX5KhfvjIs0QTlThMupH3UDakOg8e12PodVNdwXyJbOW
6ERGTiraweRDD1a+XX3KLVSnqoL6OhVLHGWbo1sZqyr02CBI2LukoHjfxQ9IKbSGn3sh/M9uNzgq
Zha6ejpqjI+Eke0cBiahq5o5SX01TfA38exFHjysmGZ9Jug8UJmbsE82A6XGpS+hdaEao42vEgSe
6OOTmQshdEUTK1L9cejF1tTQ5pr0EPF79Dqt8s1irfUBRf62+/zFS+EKvRmZFXVG5+pdxr+54VCl
pGkURGUYabH2KaY6HoaWOYG+4rQZ9kufxNLkAt/zABbthpdzw0RbiVS7PRhoCwRWYJ15fFI5ANMS
uR/e4zb1/UjUjjV7h24Ui5Td9JDg4Z5pUNCGprRIqixC103x3ShRCC4fqGyp492VsUSod7XpEOLc
pqXuyvtQhsE3JBj2buXIc5UFCVKs1i+4uk7fRpyD14HRieeLtmuSZNYgE8sqKY5QvlMWupR+9eKf
MEnks/0DdWrTbVRwgvay1cdlh1bJnrizEnnsOr2+XJVQpV1KGWZeVvA4tQ1wL/9jvJuI+DEOPhk+
kfbDGItr8G8J598JMkiwZLCDIUwUBYkBi3DWiYmjH9govxGXqQu+3TsyvArMqEE6vYx7RnmItnVE
cdswDmh3J3ETItw4EyY/Aatld6DQdvLHgoXh1lPlvjWYzOCNRdp8qQO/12qvxNMsVZVKQeBtXo2d
/XSGioohaD9NivG3v8BAFnw4G/GckkGIh+bJbagxqckjte58wW61ELxe0KvQvCKe5yxpKDbpPF7t
ggof4KEhDjsjms8k6CyePQYT32OHAPTOfYEnF0jU3CaAV6oC+y2xKcCwMNXI4ouageTFjErO6K6Q
Yd3dioz2chJzTA2rXbJYXgztbhC0p5iZkxNV7UDdgdI7V4iTRdWvxykubRdaPXr4FS68CoZp8LNB
+2blk2oranmNAeExasYl60Q1QNe20zrd47dHSUV8Ukw6CyaHiODFoFKXyO8NiRU5XmNlkBQIuBQs
ifNCqrgGgUmUzGy4AuYJO/qIh+P2CZfef0IQD6sycVyy/xFraoqg/XDG/3XXbYsQQ+KdMrCqTg0V
lWZsOuMiclFko9ovT8IhrUTKt8kf3aA+dmurbgvHTmFXJsD8q+pYe0a63NXnbpsMyJoN0l5hojmk
SzbqzZiXxFcWprJI0d4xVeNGlToRPfpMrZP3aEqqhLM5vQLqY6IJoaTube6vga8s6dtpniAuRMGJ
H6EnEhJU8FaHt8Lb4L7p8sLOoTauDlf80bcZ9sqHJrSCERC3f75cB7YMNiI6ZKCPIPIf3S3zMeJK
aUGj6B8l3k8Q6aL66oMk5F2XKnfzUUSNaH0SfVcnXBFuLHr6obrGfOWXf5XofyoSGlVNPCDjMaJ/
TUwxHfA8to3uz7Qu4ufi/zA9+0rfg11HFP4j9JMoaiOgqRSfeDeQQPPxggLonXaX/JGBKoCuLzlS
1uVC1g9/ZZZPuJQfWUguQmNPJMwUzgJt07ViSm7keBN24FXjyS8CwCwNsgEqo+xc8Kj7oLtUFAAU
xDnQ6uPBMyOBYR04lr+d50XTQnRmJL+jX+3LafWMtmJr53CPzD4MABNxUKx1tBCwJzjp4K3Bz7Hi
Fa5a9EKcHAcoWfT/Ah56UD5ygVaJ0CAeKxB+FoI4JdN/pzRdgIyn/FqTtZvdJp/SzsFSr7pMQZRn
VtSE/c83IHRYq6K7VRTGpLDFWFz+T5ysSlUa9jnsReFZ0EPSTNZ1TFEubXSmiZGv/HAbeR2Be/A0
3mV0XjPH5okf/8O7FEj9DsKpYkR3FhEYhWdMkcSdV+v97CDDNgvIIeocn1FrSoV0GngzFMtx5hPn
2D+egTHRGNg5ZO/ldQlj4BBk9dWn5UDkUGsDvQdonySsFPrtrYX6FVxKGiglMJ1dc1hPWa0QbCeQ
Jv179l5Hc+3Ya2jQl4SnWy6i/XLVv47SXHC6WCcUzGv4RP4/6IDVM9GoMi1R9QuySxhNljclO3Hz
pGxEqWr/Cd65vUu5DSWV/j6fHvdqg83xpOjJheuNgBX3Yrx38tCTgvVRrDBkQeylcoe3b4UQ1+Fn
LlIREkNFideQ5m5yIigbR/hvfVDuHSFuU+91fWY1mWmm+9DX6v80Wor5tGMZcJCIhH51Pe3GeP0Z
okjzbkhKWiCXb0bjZHD+HL1Eo2l61T5+G+VQqN8swCKNEnl6GAzeYiZQ3hi/FSF2QsnRDLyA7zVK
J3XarxE6ej2esLASD6N/P3xHmIYlL0/jibiQ/8+lPesr3Z+O///wT42sZznwjNPcjygX7KEK/hGk
A77TWDP2nSeVnrRDQB/194yn4lTTXBRtJ13Gc3CXFOdW57MHlwzuWy6SJcpbPS0VwqqjaC/Y+MEX
UtpPKPhRpYNjW9B4TELXQesTENygNG2PPOQepp2X4s+Z3hqwIf/Pv9t3YlWfQtMognKZrXrqQib5
amfbpgdrKBBJtCHgLNgVZQLjac+HorUxYk+9LCDLVxfY5TfdLjxMtNkkq9S9JXhydvXVYHKG0JrY
0oS7JVSdjQYHckXiBuklwO1PFqRihNdBHji0HUoOdpADpvshK6DktsQY2XAvOX+bVxkdYTCptUgw
JkxHNM2ZUpYjL18/WC+zbsaaLdLqtoHg8FDGXOv6jOF6K1EWwvdQxqW00RR7lQpyagqXuSRPG2av
VE69BvsA7VrQhFyQvguulrMK10NLrrr/r+Jin5UFzitPCQcvDVnggFp4zXhTQKaHGyhukiK1vly8
+ZO/w3jQYcU6Q8marA9b/AP+IuZBg+7GyUU5LDCuIBPGsGwDnM8RTeL+BsNxqj2yhy9HgOrtKtS7
dYS98iQJmHGap637n3GbkvylPEY6K/NYT6UvUneI3Y73WPxKM0kvXu1jO1NCd6np6UpxYVy6FBGz
NNLt9CBioAhh5xWPzvJ1Is7pu3hTLAFIIyMLkfmnSKelLechz0YCkfbx3W/jl8R97fEzbwrpsJPo
f1g4iHbiv78Cb8tQYsJN13bAGesMqinQ0NstgJw+dq+ESz5Pl8+IHW3DIluEnoSiP0aiWxxi87zE
O0WLfnJi4SVtlMz1xRlvTg2kPWGq4n9JtiXr8V2DVo0oNY/tbIhuQWlj4xHjdpr9Rc4f/Au3YEkJ
tR0amnESYCNoy4XVJouP6FgJf/IqxMkesEcUUjxnslH7DsuOmSAx/Iu5zw9aI1JwGgm97DETK3EF
LmGzYuCyWNg20Fqj3Qf2dIev4XxJsBQrdpNCVYZq3r4A0GRQBxkw2pnEFCfKhXLlQT+8cHWxtSdo
uKVeWeRVoxI29o/2lifHnaI5cFT3a+8M3Fh2z1gTwjjma2jccPhIeTVo7GYCP0Nxlu3Tyqy5Lr/O
GElSx5tN39yhSBWHwpFrJqYxYQaIQF/ZOyAdAcLREQuDQV4wiyblZ9wOeqHSICL3l9fuuEITa2N3
vrZhjcusaMZDjQ9MRtaUxmPPEDLtrsbNJSV9J9nMUQOMVfKjEIZabWUHAPIIp9h42oDPHGMQ7zg8
bazGtEFFqsdObBl6KcE/8pujiBclTk1PstFY7l22O1fXey0qrzg7gdsl6PD5kBg0rbRHqssSnobI
Q7BqM+vkOkAoiDkC8O4HpgCLnw9Ki9aiSF+nJXvP2nYuOMedcm7VFN9nMYQXLtWCHCSiG5eTtBJI
S1CxQm1doI/Vk/59EBo9v3pJQVnLnx5/YrJRTTnPd+HTOXII3AY0NjjDK199xQrnvL1j2fWvMpJy
M/XHRnl2fhG23eDNMvhSNigbRl9iJhpiOyiWybDo5H0Nh8TIqB0pRbjeRcGvmNsDPrjPc1aRk9hI
pfv99+MwR6QJtA5ALMt+5vEfHCNHMda2LCR8MzZ0fmP3ebbcXnATv0kkjRZEXfyMgYK/ODQ915da
J2NzKh2DPuAJjiPAqGdcbkruz3oWjj6pXI1PA5xZVFYHxk+RJT0dT0nnzMqkMzA+vmJBssAkiwOe
EKbMCD814QBbIkBBamcm69U7WilVoOBe9kG5/6lhQi0QswW/6ra2/Db79vkWOmM+gl7ssXipQWlR
U3iZ0gDDqK7xHLPGfUhuCVGSmt8jYM/mnzyHAJt7kTds9n9NZvaz4v211ydW8bftAcfuNq7Bbm3z
5+JaeFQH1vGS8PLHdMw0VndNefSEgL09ug0NyhBm0Qrh6e3DawY92FRW8o1dfUxFnu19UecCuEHv
Pd5+FsB5LnFNbMymlUtabHFjzHPwXUqBDgy3EenMwzKOR9NNWsy/u4y8FAxUxzibE8YhT91ktDpE
PP+ldKfDQqMDZTlnm//Uq0EM06kzjwsYPs8L99JRiURe0B44RkC4TS/ym7LJky6+BqV5wIK8EOyd
NsgoQOh6ul3oUOvJonCP8LH6NUDqnzTx0UICh0Vf92G/4GaNL2TnaSe+5Fksg8fkIOSbwlBt8JQ5
b9fBpfT4Ev3IeN59aBSMEk9mjYNUEpfAWB4IbAJ+5CR7rQmsjvwtvZbrR2+gQcy+Pb2+0nYAR628
Lgm/XRuE55LlcibmuO6RSUId7Kc9an2/Q6GtIDtyf9SEUddaXYnOf/ReofydW3NyGKQMQ13p+gyr
2okfuLpbQGyJdxt2EdRpY7bOcqBtMHwtIXXv5kPuoccFz6QYh252bwW3kleZmhJCXbxWbrPO4oPY
QaPKUF9hyUpw+2K7kLSGDKscQzhF+3Xa3zLOxwIINcRnQiViYg9kieBKNxq0UjdH18/DIlGIaTSy
HNV/MF51lkkEcAppQDBTGg5azKuXKnelkVkEHWKXRf1niJ34AUt3DpAu52LA0FVl4zrQhl1jIiTi
rf6XfeZhLh7CKa0hqBf420s1VOhmfeQjTrZrvdppNbJkKHjulEyBlxFq49ms2l+zLpG9AID3/EkA
4HjGLWxBE3dalQMfSWmOI5tVQtjSerbynb9QgFw5//ekxkZg8Zn50K6hnJ4XBCXHYxd05EeOIgzz
cT/f4PyfrY9WlpZ+9VqcWC4odSAGWVXRd/xHiVttdZVTMM0sUi2JS1QkXxrKcrNb5Izfob/IOA9w
jta++/pa+RRBzfOLril02M5y/+lBEYTzt/p8VCVrVwqtQQ+cWj0n79PLQfP1xabVKpt5HBE7hvXH
4d8fKrH9J17AnpatWeGNPm8EfArU7NDLDBtorGjdpQRhbEO+o05WUZDPGnIwCfq4ae1294C96xnd
xvMvJFMuURf67AilTDI4SPS7tI3ZspmbjP95nO7xkORP2gDtngaRT4gs9vPI0ScKzZoP11GOrtmy
+byrpMQ82SFkKcW9ksgGrluFdJPQEOCC+jBwVVsFe6SgX/ba3wbQ3QFej1SYgLYth6i1R+7FmxqR
AZGL05mdl7h5RRH4c0e0XrKiMdP8mu/j59noXxLAnl32BZWcOuhKE8K/TzHgPtNCxZPMov9OXvhM
QdV+j+JLmHzGe0UAPYpHJIqgjJOodZBx81POe1Wdzs8BrZr3KSJH27vUu3gb0VafMrirJSJO5rJx
KYj+gOO9k3DKSz4Mm/tihsboByBHajOutjxyfBGscrF4Lw7bH0Yc6Mdq92xXElIaFgePGGtE0/gV
XqIzOqe7MosRabvujAyxbzq5vbjEWHQBaC4UQkJz3mhBSn6eoiS4gmdznaMXN9edGjjLfqAusHAk
kBcj8/jNM1vSVq9jJu44Jy4fkLKig3lu1grpTt8/JHn37JkI+uv6aLX4KCzm89DFGUn9J+VL6bT3
P8Ukdoj06e/zc8t0/7EXLJ8V7mhU73swWtB4FCAekYHh071ZrbSYNq3jknyWEEZ2VLwrsuTIvbUG
yzF731YDzZk7XtwIkcC+eBA10xtfdzj/aT6QcQ4+Cy0mWEhlR8BHfEeE0mPry1Xtn7JP3oBzWNVb
rY/VSxbcd1iDEEadrgld8A6VYXWH2+5HnDdWiMfO02jrFd9DLL22cvaB4S9UCdu+0c9TfLQGJ3jj
eHOgkutvjxewauHt1Q8x/8s+MkpW7iSa+ujFtQbnTIOQxyvrXfK6D8k9GYqtwgwcgGIGwR9UVG2s
PeoI6nvdoxgTh4L6NW6Mq/NRAKQcIL5ITkGkjpmylYqdZ/vRvGINdn4paI+Os2oXDP5zbT2NyFhn
b07AE1cOnvP52/XGr8a+gg4boThu6XMk0XK5HK2F0H0h4hGzrRlpTuTmZ1GYbFGAMLRgQDGCkqEr
NJKQzVV+UNY1PDFsCPGCm0AvRqtwElB6+KWCF18lPVc18d979x4ZswghV9dSp3wgKwDM+KUhzO+u
KcQM0yYIM8hWvZdeX6rgt9MBlxTKEwQBCdPv3w9PTY4Jt+83hlQJK3hyrBYcm3IFjZLQhAlSHcSl
DfBWczn1Tm3eGhC4a/+sobze6ry3U8zAb687N+Tj5qoinHfI3N9nzHmygsRBpCklP9nANpkaHl+X
EwKat+Ux9TCKFYeCJGI/uNTB7zEiyTuB+nlErOFydAXc9HhnkzlTG1BUvM+LPCkfZQDulHGXVV4O
MuWTkf7KplpcuyooVYys6aXq57g0EZdq86KPwGSMJ6Xrnm9aIwCTuHLWupSj/gxLMnJ3CrAGnaLJ
/eZlUjeot4DH0HQyBCcHztS/lHD6uV3y8w6lNXK5uAvUPBVxKQcBqJTNiguwjcMEvGMCCIeJIHb4
fhncoSVfmRhqyeplQQ64Lsh03tRudUaV46Mbhv1VxhDtduAqXuHhRes6FPBMyC0p7L5bG29Dqgaf
J9LrNfCrK8+/aPpid7rWz8G6rI1vY4g1F4TKPPaGbKtI4nNwh9q/BVmGJiJKnvzarpy2LrHFgzOH
21Z1bKPoKTDGE135zcKVbh66wL0rMRJv1+YnfmB9VWSO2uhM+pNOrj5n5AboWi7+CktUfBRShPtN
yfjaCJjbVcDAY+DOFbn4U+RfhSFwRZTAJ8wf/DrG+lSEgf2RQ/Ew8d8enbzI3iGfdP74FUvVRojg
ftpnvu5DOh2lyYUpLBAKb6z1bhMFkqGfAPgh0RRw+fchX3nb9NMA//rK/3I1pmFO9+To4kgLgn5B
LX2rxcWdypRex6pHHmpRPEFksonbnyRe64mCuY7UIDeBh4FkLDrN5/1GoegdnwTfnjDVHebkscc0
Kk8gyHCM7DVtE0oE/Ro/tSM6bgiU/smxfmKR09RgSaYEpo+zb7zD3ecKDV3DLWfjLHrNJw/P0E4K
dxXm8aQWWA3w2vc/yeJ2CZ2VghtcsbMtwIMuUyW1l7AmvyRltTU1Mt93Te/fasrOOhuWoErt9ADY
QqrP23SFt6OFVv6TKbz+FnHl7l2WFMISpT428xgKVSBAKn2V0KoPdQuVCqDk0BP/zxjloiHcYWxh
0u+/Jdq3wqf6rEbwCiksCjJ+1AJuahLw9lR2PnsEPjRYkZdx8tycHvUyWR0l9DAwX7pBOTFr7Y2X
/MdL//YZJpR/IJORAtOY/7+CFg5mWd7Pk5oAIWRZvrOPmwTHhjivLnTveHLX8k21mv0DQSPSDoX1
h6ENyyEWXOE25XTQ0HxvRdTBTlSwHdiHAhqucYm+Gv0e0W/+Dhe7P4oQWlFGh3t3Q7saDyM10wC7
kyipEz2ZcKp1HdrSk79QVYpgeKd+FFuP98Kin9oyDZ3UB209lz/dh5/cXfhjIeCcfqnHsNlqZ3JB
i9pAj79tJVvNF7y00LSWIEmt45FETavVte0zEkCUZnqtf4ZNMhZhqrbMJGcR7u/c/gQGFDEKDn2e
cJBjbFPaSRgFAsidedknAN1u/YnPZK6WKf2+IZ4uN4NAfc285T7IyqS1vYDT6sPaGm4wn9v/xguQ
Tz9uOD94CDora8NiRsjBoZob8mFc4wrH2FKv4wwqOykSzub/65e3bLyVHF0nMHtmojcndzwHxtpG
9jtg4x7AF0gkDkDnn5y7FFWLFICu5VggaVLmDYYo13m8JbgWtvLYyyE+Z4GA5xI2qrwj4gGdCZ6z
cSzjJMZErH313RrK36Of8muKrN72YwR9QFWQ6e/tD4JNM0rOZ5qQZuW26A31Cqsl9H/FZMTboIId
JmsqnNwRf38a3Ssxd9xPchkuEggHXQ2266nYlUwzqmRLbXjhf0hHtqoAOAKmiXe8vP4xY5odAP0v
FnkHYNYvtC3BV66vqos9naKY6ggfnqrqJm4qmNTPBhpaT8gQ68ruNu3otfOWKeCUozl01qS6FJSE
z3LCCm/d1Bf6ujp4HsVeO+qVQiokSJzR65O4/DFav7zmNl5c0ry2qD/UlJ68gif+ScgDG54vPz5k
7r+nvUJTzqydUPc3TiN8A1Lat0mX72GkWDwqINTD5Rww3OkZVqCb218iWgzUM6MRX4OHsNJvLtr7
tuOuMEBeWf6Zee5hSN1+x/64efXbbpguWwqzwNmH2CSuTmWGtouTakdAUj/+M1BWSs73S6PeJMnq
KxXtbOT3nzxp6m77nQyAsO2A275BLZS/xh4XHIryAgz0le61PzClY7l7crbDU0VEeSxicIHT6Mgi
v3XkIj8cwDyPVyAIVukyXOJTvQe2gobx+rJJ/4SNHpkPyfgCU0dj9ZZiSDAZbBQO5igoLSLW3aAP
Uf5Sj7nTzgD6hyHYW6TFn7FbN1d0Lpfagj7oyp0d6sYbynpfbVcYMCU3j1Ht/UQIs7CT82G7HA0K
8+yg4cC4RhD9AK55Y2g43pz4Tjhvnf/tT34YXwHXxdbJx2A+dP11PbelgSrM59eaOXYxnPWELYmj
m4WQQWJ9L+1QofYc5WU2VnrksFsKawme/ilutGBySy/cVA6C/EsOoc3pztkL+G+lMhPDOUjgKgHl
+ig2WdsdSISPkI3qRgmzK2S61zBYSgtWf2Rt4hO2UL5Yb2j72y1rzZmqvPbQlrgGfWmDKCisk9cU
nx07E6fKAcPnozuAos9jYBvdhdCNRhJXE9aBu7ogPhFgctReIfe82q6INFhbcyui2JPbLlR+Piu3
DHwNMP6q5LjbXEqY7WaQFZuEe9sjkQsUzjhH1WrevCEo+y9vr86S5SQwB7K9sEmdEQJktm/lDQk1
yOdL8USRG1896qmGlu1S6ZNlm4WBrOzcpURJOdRvC+qVaZ+8FdHs3JI+LG5OODROr2+NOpNiwmQq
TEeL8JpNYUESRULKXao3biGg2+KgX/3pkhsFcm31CFcbSbGy/Gd56duNHFOpe+cvg0Z1MLZLrJte
4nQq3whpXZoT9MtRWYDcIibyTxxHPPlB4Yw662UDdLmlgRi3JyeTqCGrwTYZHj38KDpXIYLP/784
XVYjy4pG+nSe0sVPV1EGZ3ZUVzIA4fq+lrR/y4I8GKuDGpv3EtZ9iSo2ZkbaW59OB1f1dXEJ8JX8
wrjdhG1Cc84VMBt2Ircq4G14HgPB42Tzo0ydm/jtxEtISDVlGGXCUPNWb/Qux3W5zaqCFfLsZT1k
nNLT/k/iWAkDvEn7kYM4nHOUP5e0SX4vjiBGkZNDapIPXIe4sx1bwglBYUmpr/LNTyR6Um5vnC1B
5ge33eddmB0QuU5i3MZgQnZ/fnB4BBv5TNQJo5qajWIaK3Zu5R+PoGGpyl3rTP7G/5g3z64MV8SK
zHFkjw7PuxyeNn/YeL0brupMdqtibEzv15P0zrTZbK6WckZvflxHzbODEoIXHTogw63aFQeG2MA+
+YsGKAHxASzOrEqZLEVC6HOADQnKqHm91jjq1SvSm1AddKg8PO2w58KpdX2EqsZfbynK9yaLy4Lo
Ep7X4lnKnGcx7EkRKHL3PlBWqQIkoufQcE3dvegzJZ8LAKXz3BkhnKPHRV2Qq9xc7UeQaVSSNv6u
uj3dRKMD1nAP+TVhMW/OR290eJueNE+CeUyQV5aW7CPXPSrHvrA/4KHP4kxmQ2CYI9EKIUfIZzM4
9ysTpFXU4Jc7wdUZUQ3Va8SQKTplRbnl8X+mr1NPqH6d8+E3K4S/XqSw8EyvM+DquAAMS6CzRdCj
+ToOwKXQN+pKiEboiBCIwZWyPUs/AFePTP1B6NzZ3sB83DJVXeAa4zbDmpAQlWP1W9MxhIN+WLPx
domLirhax34SDuIH80yTunnRfMINhsDhpGsozW2iflRA99nDCzXmc+n8DCKgrDdnfbz5DNd9Q/DC
+O6p6XcWi+TJ3s9aqYuPwU8ihVCknvdstkr2bdYId4T2SmXpPMaGqpQMy6iX8yLDhbVaVjF1Bolh
7sXLoEOP+hzaKbIWoP7C9lB5NyfZMfr2m7o3HYwXLZZSCRgmf6VG1pKIgwff+ElU6llBsxIpxrHp
KosTiVXTq/unzkPnZ2P1tDK3Y2xzYT1LDoYjSMPqFlYhkw9nHFbtEGZx93hc+5ISzlm4SKcfJ85O
l1kFyO/8Eku21vj3mRWOC7tXLYpfhCdkmjEvvH4jFlhpjG4F4JfR+AiNGVLBFVBK5/LTqZ2Ega98
wSZAO3ogqaoSyy5jzGKkxGlhA7uWybsnHQ1vn6DnGg1iKvpkew80r7O5ovOSGPGxxAqU59XK6CZt
o+yEO0qHCFcOypkiO51Q02sJM0ae8jyLKlgmpS03aEAMSckszcDcPjukTnp9aenkQwmnC9lEoSjH
nxsRe7BoIZhU9kQu971XCoObJc9WyS/K3buH1wudj08Barp6biP9a3BDZzwoB8bunDXG6N5qlped
IGngsQb6mQbWbPtHywUedmgwXdz91p0W4gJWjXVAf8x5/muZExRR8bk+afk8PHtRa5fbzBqysT1L
PFqRjNQfci99ycrl4wDEHY23aZLi5cqJ3jias44oaaWT2QgRGLTqP/FA5JQ21p+nZ2J58ajyMLlG
WP/ofWc2Zl7kwTq7LTfpcpZDPLJu0MCXrtJIMmcxo7MCoKX8ReOoccdtaph9LcMkDehxacW3RETO
GiUvwXqkojcK76MsTh5UwxnOkihKFaLYgkRkg3tbD9p/ra31O5PCVCtffvXc0Bmwnf6SovkX/fSH
okPXLxgecRrnarEIpOlX2ao5qKLM6Zjgbq/3n0kE9NTTNOFr0MgHVL7NejMCEG7AFoMeP9vabqDR
qLP3SWd5pU3nfaKMaKuqDJd7WNBIIa/oRC1vkkeQyVIoYZjHmdxrwdjj6OdhkwqxOlNUzfIKPKuG
innJENiFL0YxVzBsWZpRTAx+RPjlOWMKpExGar6rDsE31E391/9D9VPjTvs9H5mb6k0m/YZCfO0z
NTi0aSDeVab65qv7KfyUQtwExoiEp/8NE7sAOmXLZ2PVIi9uEzROOHrn4mJvX5uPDzTS07XreK3x
3IvPx7Nt0Jog57tolngS7GaoRoAOyk0ZAFgxviB5JDX/AFEIGle/WQQnO9AL5ur9F94ZU1H9/2Lb
7N7rmufDpE7TdAWsfwEtKVs7yYLvhcjR9zAl2emlqf92hPRCGPZyznLtfoWTClhz4wmYadDDdfUH
tyuSY8DE6P9dl43WDzbp8MbNT5pYgfF22yXN3hGMAszWS27WFkkPDcldCzlw/r4eRjzV09x3XXZV
7WIL1QZodRLa77kf+5DlOBblJtg+fqUHcvmC5waiZ97QTiwCi/eeWU5WJTxmLMqduKby44TbBzgr
Gxev3PD+d2iHbSKjp4+s8IEuNZ1zDPYDAy3AYDO8jDDIlkJtm0D7U4l59u4Rj6ns778UIhoN/TeX
p59OX4AZulbRwuDwNqX1iuEKIPnvZtYXdKWIpVWFtAODKmE47yr2/JT1h69q0X905VSIQPRMmYmT
SSmXjsg9z6DRuo+lIou2hDavXYL1Uc4ewGcrMtKbOVthVheFA7R55XudW1C6tjwjE6m4H2PmmyeH
v/y5WBKl7fsYz+CMZiGdsD1G8wsT0E9qeztEWqq3FMvwLe/qOP96OGc+1FCWm+nqXItKn/T5WgfA
pGUK3I6dOrRHCADaRzslmF1F3SOU+pHjPM9LA9Wk2G6ce+cd++/EVFbVPkg1PMuvmBeUbqFEHoLB
MvZJJu5a6ZTU+t0ps23wY/K0XMJBeAYY7Uhmcjl7o0sl/H4L/ujv0BimUtC8jJJeCgz62IXEmRWC
wY+xAW8aBd9K3/KvcLmBrB/srnTg2dhQOAg0YyY1HgHrjF9tcHDVIcSBID/mWs7Y86slInzP+kE2
mxEizUZYZUy0jNWnn87FPKL5n/UFEpWEuktKBP4CEFtTgv9vW2l21WFwh4AZD5Lvx4UaxjUVFtPx
3PbafCR+ZqfGQeHn4f4CAmXBSxayWE2sxOpIu/7VdkOkAlpq81nn5+AJ5EpNrQjc+CpHWReupkqf
EumzYjtacuZ8m+bPinMtWxffSbPeBXiDEhNpe+Rj2xmeByE/u1/q4B/9qQi/w/lJ3G57mlmCNppK
gdq4VdvKcy0xwuUamprXBo0xl1rUEw8MaN/eV6MbZsbs4z6EGJxixRlAk4xRGG10jCHWV5+gOyx4
8RX3FqKGVEfJR5XR+96eMuhD1gf8BhyCNjv9Btr/+B5oGvrqKntJbfanavBiWxrLdSJAyC+RU9hm
B7vILQ+Zlt/hR2wGU0FkeoqINeTXetqy5Ve4eqCpnHzq0/zuT6bMPuL/4qet6CCl/iYmk4q7S7X/
cGRTaTg8YQgRtKaxCPj17AKQNWKaPZnJdR/5PHWqKTjMItYmlZT+ZrHKfirMd/NAegOI2VsS2ZTx
RdNtjX+V1aiQOr4fBTkwMDnJzTcUX7SfQiz6mr0WIDPQiLmXBeFg2eSYDUle8gRv9hUm5K/QfOsR
O+Vb4no0CsNV7MouId+v2SnS0bWOPProS1zzw9X8H8qmCYWU9ZvKBuphBJ1hHNLumT/IC2zSAyGV
8ypPfU1Hwr/dt74+Hmrp3Xe1lldifqCQsHSmjDHOlAM/KyTVygHM1Mxufh/Q3UxS+CAc0LGvi1ux
vkQuBP2OmhKRwzVZEns9c8l/02I2aYy6ye1puCr7XMJJg9sdb5PY9vlw79KAs9DkglxzmSkSPw/6
8dZDoAfOPa3araNZeyZsQPHFiS5M7D1p5I/3X4mKi/FnTH7LL/Hf7HzO80ODA2a2kpHDfuIT9htO
JhVD/9VvZRjtTJ4gK1Q0+/8mu4GOpwr4imw4dx38Wtpgj318pHGYTLtcN99ormsRs8VdWwbhcYYI
KbNDvCiZr0GiygFScSoXkAK9CPi/Cvp8S8/bicvUEtrl9sVyxO911vhuBw5x3hW441RM6SGM0mcI
sSP7AM0fzTlFtvwBoEm3MJ5cn3KPcI+LrlHxbt1kHSfPXfOuoN1iEHw4xKIHLVBtUPyy6Ml0VCj4
dafeO5Lw53XinYF8RUJeJKjHKhyaMiSoTa8MQ+eo4rCsZMIm7zhPPYsbPMxtIwIv8IdBIvQDwDkf
nFlsI3OqYrxf+BjPbEliv7qwysmL29uKzJ/61uNWyUx5LTH9cHuouVxary8+ZKdV+8QfiFjKwEwD
Caf3ivKB9LvfFXfYLwiefjb53JC7k8hVJqDcxELRHKMB+sso0T/qjo0YYkV/HUya8b3l306vL0/R
4+fl0ScivNEDUC8n/K1SmZ/QkgMbxXAOmN/vrth7a29gayHAwSYI12quGpbn1JM732knIFRHjFwI
mQtUKki54YZRnaf2UP6F+n7snfBF572LL83Gb/DBl4eUuciMzll3yIBBq9GUfxipBqZD5V/ZvFYe
tSAjP02w2+UL68vlr1V5HQAOcf5f9xD4HAAyPpHEJuK7jS5GcSSd+y5BN02TazJuGyAuQf9MhoTd
IXVwGrYjqY0Nxqcb1w425OT/wf1FP4rGNGnPi5grOAyQinNwu+dr4qPZIUudq8Ek/z3LOnkJZ3AR
47xhq1qxKPh27RkbiWFPPUf0quXD5gpkQP71sex0M+DoBspN+cCIlMDjOM2MfQeX8UL6a34xhllw
mc6sUTegCdpSTtNWExGH8/T5ftSfiFNund+EY65lwcPlJ8qGqJ3HbV67iUGlb//J/hs77ONX2HK2
KqKvfn1s4eaHv+8b7hdc22yCI09bcurBsWLeZy0Xsa5itU0o1kFEyYD0pPLirgHqyCM1HCFhxy5w
5gfE/V0Lo3tCuMVY0jiXEzZXCO2eQMBLWuLXr/F/2nstpHtuepze7wwNs5qsA5RJrQsdd8tquBFv
U5mszGAQCJtupizy0WZ1OMJg7CQLnkyA/mP9GcybM1QqC5EWgc9bbOgHnAqVtSsbNyILgS32uuxK
IzKZ2TFRqIF7eeEqn75NA7LZHLkjkQ4Wl6kH8KNRpF8Zyr806HQWJc9xkfb1fKbVm0xEuv+4YyUB
VF4fbjfIYC/OScL0tgyOMXy66MBEsXtFYkp0lWWMy0x5SOJDBHfu+E5LOPW1lUhiOLrhq435DJ0H
4SbmCxW490yELo4FIiaLsjbrQhsf/zMBuB0q8BnvQptIn4+obaeyqNa8qMi4mdXYxo1lcwopYBvD
srTop/+sI9AqlrIRdMqmRRx6X3cpvea5rmE2DRWza+RioIjZuvhwn4450zqGZEGnbtDw7Zjr6H/l
Js1qGXzeo1Bkt8VkSa1fzy+aXMyjXqkLKA75RCXrYMG4KiTNv9PB91CruKz88I1R2vqzt/inucGp
aVizcdNKT7vfsOfYwuLGVeIO/wVSNTL6p5dKAmQh8ENTcXdtnScmLuU5UF1bk6vjkPbEZZp0e+DE
RPgfTbzkIcLpzhQQDR2w+RjfkNb1/5en71O72hhZ4+7FHF2ng3rz3zp5EWRGAosH0M+NtqmU6tqy
5QaOWFDgaZE7Ig/MB1pQ9kIyewiRrImxEpp9w64dGPFB34ipi+LcZB54nP5n1dqmHgUJNF1TySqN
Px1XMuJne0gCCU2WWjMfJGBrhPMt3VpXqUHrsfqcR3Uhg7AZcgqXPuB2bwWVwrNaNgY8p462V+gQ
dkdPaAKCKGUtOihvAwZtfmOQSvYQD8dW34u2zk0RGqU0JYcU3thHx6UEdCa6mN2kQQi+g/7czaid
NBrL6/FdXyWh0nxWFzizgrfxXGvdp0gAmv4Wm/e2MusXRc9FAiixjfIKHJAFIGDRPqXZMdZNG2oe
bNeURY93340rKcajVBdq3gEFiNgYzECmTrmrRXOQcTED00vMre8wpw6W8FZ0eHL95erfsfzasGbe
PjogWKvEjX4ix3UK0XIIH6v01rgnXlVvVK0SnNWTnRDQIeBcUqoi6cicigyDQEE6+MCKFh9/VF+C
+4XewqmP7eosqCdcQpiv7XVv/gVyB72tOh97zPJT1ymzppRc09Ap3D0vDHD+SoFuWMfNpjlkZtta
wtSk6m9bqdA5pwzD8MMDp8dcROeY+XZie1naLNHiqbM5FGILfKe+2Cw0g8R1g0EQ3VzCpFvYecVo
1AbIQ8jX3sDeh0vBUhaLtF5azPM2DuxQiRjjb8Qv7oEJoZ6cYYxKwPlFaqZl+GBF9902cxgZDP4P
smi1MLTJP5qWWe1790gxYx72y/YanSLG51JKMQJsCtf3f9JxR7TJVg8vJ8Y6+lI7t7BR9KzF5GPp
74q9G5yOx3NROOexC4m91DoF4WiHzqpHt3wU7dMe+Xsz1nygQq78MW7KX8Qdt1TQDfI5JqJDUIfJ
Nm5Ta+xhZ5wQsZ2eCTY0EonBV36cDiFcK7xnw0E8kWzw7xFBjTOFxkH6yu0G0G8cKaxEzfroPeVO
0HlDMYCizPLinnz6K4zteIYoCxV9Zee1T9LA8jRuCE5QrpZfALoU0p1WIhTU4RT+F1z0RdBZQ+Y4
w8TKJdn6EiEu+3ewBoQCzHkiNrgtd9hkEuXfmZt62utLcbaj0bvQgRzkTENcc3ItXpZURiqf3ctJ
jzNruHl6L9LkFuNaMSEbHE4yz7hBsqexaAHohlVxLpLDfPyMCHRViBVcnw3ZBVTuuXo9tgxy+3Mx
c1S/f7+Iw+axx0fHe82HL3/OHIofdhklmHqO729W/jZgh9ImrpTXT34PvemnsDc7Ef9F9Vrx8Nbl
3rWopTbn432u5xVhGgnFLUr0z9Cb16dcJVaWwVtq0yMtNo80VkSP/qo2CrPc86fz930Zd9c62Ia/
xNLgk5QyILm/kLI3xqyHlp6RzvJ+8pCTEaDUelq7AnMGl57uUxbrjoi2n2orTGVQhC3FYB1LDsUD
8XZmz86xZVuDI94iLb7XbJk+U+jM6NiFsGWUv9+mdtALewYx3aPAptMZ0u0l5922Pqd0M1u/x8Oh
FzdMoiPQDN8BrFLgw/PEsu7MOlriUaEVfpQTHkh+ASlMmb0+69xUD9x/VON5rlroSJvPRQZfAXom
S6aeOYgyiXIQhe1vWJOpT2sgZm+Tt0LD1RC5GnDniXyDcyvfHvUaJizxW29cnS1+FZfwZshSbSMx
5b7YbHIVC77dhWBCGXksS8Iq9SHSSeYyFGBWjL/FxI6QyBuWAE14o/B9DFMCRkcd3Rq3TvQr4ojk
S4dbeN6M4KjWwwy1CFtM7FDjXOqSO1ObP8kOz2Aul5CJynJWGwVYNoPn2+Ae6GE5d6WWfFjwQDkn
JVbDyVrt65EZPZDkc3u3KOtngGzxwsQ4u/VOWmbGzkpZliySKTdN4OEg6EYRyG4WSPo7tcL3u8TL
XIbmGAxYlJ94mK4axSLPew/TpB4X6wuq18gFBfRzw4SQfVZ+gunDQq023LJM+1Dyl9N1Y0RPKltr
5kqrFhLG7ICaWAxDLoZT5yN1aE3m7T/fi84RaQPa0dAgBXyQlWE6tmD08bh5UU4IktQaDHu7la4I
ZP/69vKMMvtLubb2qaKzO2TND2zYgXxcteIlpN+4Bf8ZBWO4UVNbL5YlkXD/KTEulVdyGPCFANoq
Kmt7TKLa6Z81bCShoqRXSG5w26rB7IOYaRtaRtyXk6+pa3PhkVF+t96O/L2qqVkNQpz9NKzfq8AQ
VXvSD9Cgf84JCZ5KtFxf3KhA3IpPSCc4134XYCX1BV6x+vVtOzrU8JAgQJQC35Mq/SCK+K92GuDy
i/KOxoS7eEn/LGRbj5qo+AIdERWEygXVeTPNDXK03ho6GSnhTv9TY6lvU8peN4yEZcrozHEQJ3+X
z/rKWEQXsALT/n4WJ2bnO+yzg/9UMguTUH6LGha+IB6W2/haqZuZ78Yd1kkmTJY5j18xqF5tzM4F
tyfyF8KAQuheuFHGod7Y7V/h6FOvZewqnhwYiA7HYP6Pyr9MGb647lBkKz5F4fVYAlA5QEUh+JTH
eUvv8Hpcsm9zUZWgy2MYoaJmaSisq4znPAoq25VL1pfBiMT82kRTSP80WuOQxBX0PdBdsuz1V1hL
B857OPWhSpwyzxNso+FseuMdN093uCZUi/Cjdpn9nW7Bsogwa131Ac87iJjGyN2gBKYa4HAfSRoX
PsD6scUBqe0lKT03qpYSD2Hpr4YoSyVJMt+RT66U378hDBBN/BgQMrDnD4ZU4GDcP+jK1Vpd8nHN
UToPdrDTz6L8Y6fnuwxhPkXByA05jCGnPyU54vduzkrl0jIErltgxysHMBYb3szbBROg+iiUF0nz
twNtP0rPFqAwpysG5usdcTSqyHDP3CW7XLLT5W8dgghLO78sd2/lKs3tdqZo9qFt/ihNzcgrGpIB
uBOUmzaJ3BA2uHrxBOgM9/6r0eiGATyjb436wABR3VaXcVQElIHQOq8WUt1W94bzKz2v5A7JEoSj
73kJD6JSNs73FDk6uzg6KsBHnvvWW8UH064SVv+nI1OYpVJTY5rBOUUmx24uiUgEtNy45vSoEXm9
B8DwwB/zZcBhi67hd0JxTYwK9PU6xT/lZFTY13Si8NObqJ+2kwmM3dxVUwohpOSSvPvZ2Ywv7ptc
tMCrdop/FQj77dbq4b+CEfEFpgZ4JgSLZlOwrRd5Mz1jMgqb4mkISUeL+tQEeGGh12MlOLUGcpYa
9u4no11NHiYBrYZnJk8rHK18wQ57ZLDnfWT6P/Kfn9qxpVsm3I/NQHxVgLUCr97Q5WB3DOsQByx9
qusYkt/og4Uyn2KevJnhKVjCLc/3+FF3uXcBPXHkWhbc2XsuUDJ2U64uaxmGpZW/KRRVylbIEK+S
spGXiXXcy0I74hex735AFJzBrnlDukSLHikgTPJjhAXmvyeYz5dFRvd2TBG2a8PTTEC4AJA1bQdn
FFNuQTnv9nzm53JIrr0te93yHL+ePeDT4VMpRNFknpYTb3iMqG4vkqjqP+HjievUtGUlI+TvGNFl
rSITjdzpHPsYul1zzi5EEgP90cGc+hFNNpne3v/dEPybAt5wwH49auwpRroIi+WyVOgybUPCasjw
JMHYU+TtXW63iqCV05d7BvhotFKoUA1RlKVA+YS3qb6Co8sK8Pwiz1vBUIj8/FJQZTAQASAFJSXn
LY8TuDSLdqeN/Ae+KNVPdQICVJ15ia5RdKGEOfmUBeTicnrSNsp8NDNzS+BSoJnLP3fXNqvB3YVV
yAH0GbTiRkgC81DFN0Fu4d9hp0/ii2eMmAed0MtMOuGebrB3y/tml+icbqqPnnX6oKqnzT3K0KOx
bmn0A3Y/ha13eoviQ6niDUVWUedx2s8K4+qKNGTI3OYfldlmfz5esIuROih1zWLCcj30gaLMKVi4
3N1Vphd6mNZ+UtpCP5oYqD9JlGxEVTsKEs/ruzzRKj1k+IT3u55NHkqrd0Sp9vJGY5QhFR2ElhNv
RVyOW8xhmnBqME8bqmwfHkjnEcBqLHPYP2gQyUnWD9KmdgyiwPlIT4Pez3PVJn0yFJ3QAwe1XnOu
kM7azUDGZGsvx5tJYf+Eo87KKeZ3XjM4sQVCZBMAZIEspxPmCKxNdcVGC4Ltx3i1z12v6iamrpYY
4TkIzMCql0obcI6qQLzMN0T9LQ+XSkNe5qOFbUjLj+K3Sh5Ah3pY8k5sB5DpbDdTQ2qJyAO7Hz4V
JRMPOPqCT9KO1ICCyjADkfc+UQNLucF//AE73vqTc9GezuUR/zzg6SArL2KTmry8KKs901Vp6NO6
70/3omA0krzs5kSiAXUFL/GRVYx+Gxyp2mAfzTfJP6O1I5p9sWgQac9poVljRdE5RU6LSvXcws4y
yEu0vmx9oWe3fcVCT8QRM+OpVnVZXMxnePuHbxPbNELJKn2jT42NXgGwhaRC+9GeZubUVlirJk9m
1Mi8EonLp/o2DXrAsTCkZHWhqakbdeKQd5049QPWT2htOQveXKZg8s7A/Yb9acBHqJm8GL55LbBt
wsqjkPmtiVHnxQ1h6hXM8P7PzASt9t74nzbaIc4RVymS9bIwYLoegYyqAWt1nwRpZcLc8TXB1mxJ
64uoH/WpBA0UzrMRbuJAcx1kZM5SJuEXipHvWDTXkInnMpaAdMOsp5kVh7iGF4fTnJwzOjOR669f
kb135ym1tYOyGP/34XrVtnej3MYY/waDlLgJc6GHDHxkV10VQhLM24v9pJeLX13EViUpcaFpJt7o
5BENGDCgWv7wj7I5fOE1o7UO+rxLfX+u5iibx9cIemskUpEmsFq2aptKscJE6p33OzoqSiMv+Qe9
icQYSxlaQKyKup/bNJUi/xrTeHY//JYP9mjpELOqy7ShixA3uvP2JLnzPUjJeMEPlDgX7A4PcPb9
e+PuPyKxUIzZpfOY+KQpjQFFuboViSaa3Uzkzg78yIbSBdD1aQ76OY3+7xuEhnzrU2Yr9PBzwIAM
VibTNGQaGg/6P8SILqgCGpBusr5gIEp6aW5FH8e9LT8z6ZJL0Al7IHQJ73CkAjvdNc6o7G9Lw1gy
fksaFnJKXmwJQRtIPBSCVmFcybHQnt0RYip3gH2owfemaNMuPQyOGDTa51Vk6xL3fz/U54PXAWh9
PDhmiiVlCvG8aYuYtp9q+UYH21YN0I4mlqMo4XtLA3wzaNCUD25Dtv8VG8jgtIEBqBCin26CoqjH
tFQ2lDUOm6cJD9CE7P2AYrJDGiTkWw7PAV8vUcoBhzwdX/1O5SqvLokEf1Wr5010s6qsQDxaQ9n+
fEtQLlFfn0EBAU8953AogNy58hwmUv4Ro8yVdAytFOsN4D3DxLJCuGSq27vqZ1XJV79Zw9l9a1jw
q2FyM8L+u0Zykm+nYpMdy0Y70SFaQm88sIQLihaCRdwenJros44jrgLZkPUKRmEJUHtapDeIEWTG
PwrKkXJ9TjmZNms2drYu+6LbnhgE6YsHhcofGUa0Hn7n9Ahg3DV6L2tfFzoBX2F0s+vHvPSYwqOX
lgLN9nzdLD46/6NtLYyOaj0YtmsMlurFZsf8o+/3qcAhqVY8+1wHPjsNyarDAIUMAszHmB/gFIej
lNNTS/3Us2zYK9mKD74OrvqgYpqIDQBBKIH3VKCDP8SXsgspFaZMtcHwaCoA1S+SCZxyZJIm+tm1
CV4TzOzBfJjJBnVcljcczmDtTfi4Q3s7mLwmvCdGj2srZC86AvY8tJKN+Ic5e+/VfmhWDVltsFj7
/4jwNdxCFT/rRWM+SWT2UPzQjxZ926PsQg4avTgHcrVpz+GCXBNdj2pcJidsh1tHgBIjNKQdeioW
g74QH7wKj52ISJ9XugSCyYuuZ03J+CjuijXDGzzdV1cwIUDtzgyYnddIt03UkRMXvwrkz2XEKBFI
eoIILu4wBtd0r4zMOxkcs1B34RCLCunO+DvCvSyqAioD7nFZDb4ZitWUAsdjKhSVcZKgs5j+6DLk
ZHnoVPt1z8il0s4V3Bc4YcrTYXyroim0qaUcjldSGUdMkVmcDV26QxQb9N4OSyluT1tUV/asdC17
OPRc/ZKhD8nsA+IiVqN+I0qE4fk04p8DnvcgM9t2vCMbgGktkW4pJiezObH5S1p6Y2QnGQKaOPZo
9x1QXLMIKV7tUkwOeLs1KSq26iOGeU9wbgO4usxdtczOLCtZObA/Y8bNWxrKW2eD83saO0Q96xHC
wmcxCNM8K9cOY5JhsK569S4Rb8kcHoqp2E9MWJykwjBHsrwkl7CUhzYb8WMHBtTcMub4K5aYAgWG
7kmI8vmutbDEN745DdUrDSqFcwQCDzTXdDk5A80o2SYrVi+jGxe3CWO/748cWuFPE15SWpd/BST5
W0xGFlnyMR1X4fQgFHWf4qGWoW7FdTer3qASnikv9f0t1jptxcN0XItkIE2p/g17eCSTvI0NTjFM
r4kkk9uedxYahVmTWOtbjnGnBWquNw5Yrjg1fhAYa9SqEpefq7BN1lYejQ+/tpzpwYYVT+F/TvHP
hs48Jl/HcyWqbu/OzTmZVi+dXNllgHZl2zlyERGHlNk0R/VxllKAOEc1RXWvH3ZCVD7wE6TZnf6G
Rk9jMVOc7Slh+YAteNp5Be/rbgBK3/fEV7cVctV9hOC6zHNeUz66Fk/fPmx46q3csbLGAJ7ojuL6
tTiAToE9Z8m12B0BKrXCMePBxFmenK3igqS/MOrWYsJRL7YmVrnVTsQQ5305xlOi3SrLze/nIj+C
vABX3qOZSlfPa6oW8LDUnWIbkC3BKJslDCh3bm6Kv5CsBOUGWV+LkOsp2FnhIBEkcBU9TaxvqYLt
AR4+4PW19KzlYm+FQ3xwSQqTiwMY+ySWsJ8O37G1cTxELa7d4hbZ+acjYmsyfzyMpM867dTBtLbw
CY5W2iCkiX82ndl54F9C7ru7fKz7b17zWWRIt/fvenp0R3X4WKEdM0ILnO2EtRJAfzan2Jm3fmju
Y82ghtEXKjfBGC7zNJyzgFfK2uonaptH4QVceE5PCfiqjPoUjZxX82EbNS3lN39jiMf2PYt/gH8A
18+EHkFJPQpr1oxInwdbsprGND+lIXANtR74gOmBHhp3Mo4ekxCX/hrwZTxXY6Cw8XSRqwVP+Znl
nECSr39ZWSmBuzLaQkQjwLS71QTmctyvY4mR9GMvaOGnAIToYiy+yKkB2ChNey7DIDM/MY8DI8BX
/eUQI67KZD46vpi66RFAnuB7b+A0W6b5UWEdCmoZC6zP1pg9Weh1nzNp6zR8kiUJ56xPNcKy1nwq
zxzz7ucMDrwdwxlbZ4ovNOziJf/xloA4zwjo6Vo/gVrU0HA06hmpXW2MyafBRy3SHxT1Cz9qVOE2
17b0BCeJE1yqysiKiPYPr4G8jL8CZMiamyRE8hZGnag5e8qDmsLLvg5KqYyBhWLyO931dupuhdTR
T6htRAjljmq3/Hlx0TDO4p/cxPfZh1ajGc48s0yJW6h4BZhJ/gstfipKIUheEbH84cfFqmG6uUQR
2i7+WTuJKfFQqHDUWn9BpsD10Yp1Ex0yVqTAoZqziKAofCsoKdmWkLo0iwH+95LHS9fDvd3mTcFy
4v/pZIYgi4QEmwlaVntIPJLl3zDzYUFL5qxF90IrCp/zhx2/7iwNMS/v9mqO5u2a8SEpe4f+goKc
M3n62Vq7UClW0xXlj+BT3T4vN9CIvFFUey//UYYrFbpGYau7zhEPQsHCOmHwDkirx5dxsD1b0e+x
8gLwT1vFluUZq/YG6kydZTpRrhduc9A35KJlmCLazGyDMOh4hyo/8ckfkuFk6/lnESo0CnNkn0M5
PfImqA5fhK8e6GwUv0rESKsCDyuKdcXfnpdT3/SYhnlkfeaN8kSJIetYhks6YM/g8KhJvOuIF+PY
YOyZYDuAEqFWh9ct5ngRAmwDwPQ93oaey/qS9SeE29v8KUypG3hN9jMK4/vYavhCv51hEtI7NFOO
vTxb0YEasEg77slLu4LEfI5oHfVEJTczCQF8yRMEv0V6NXOlnwEcMIlh8+f797RnUWzZo3RmqSQN
twXE93ZEeCT4EdSZi10bU0r3SjllMI51ZHOtdp24IbCOR0Ms2m4r7uPvhYrOKvOaPOV9OVZZT+ux
K8+TYsGbmrFYZpx1DXehMbf7w9k/q8ZNoOsdfUzFtA/gZGEwL0SiT/ruQdawOjSRH5CLKiebHFhH
DiEbSBbt9CHIIg4FHU5r1rvu+6Szq29kWDVPmfZj+S6nuBsNDGTW1X1XrZLO01trYe9EPaj5FXKW
j3nIbGfM/364d42LgsIl4b2yawpZ9f3QQ34lsrI52hFWdgD+cv7sNk9TQ+M78BJVZp8kIPEkfxEH
tpeZCim4/sji0+0tg8i5Jd/uruoHVir1p+sZZJERv+dqlMc5ILdiNRJA0+gG5oRt/UxFJHrz86Q2
MKMhVvhIXfVzROMJ5TxmBihtELWUM6vkkg1lwyHNzzyxpd1W1yd6K6dGex2yoJtd8oR8FhwI68Cs
Z3ecO55RnsBmpLuf/xeHoo7N3hzfBcb8wcIsAp2Lcg8VEbsfYlzdWwhVyfJfZ8Z8ZjcyTXllADWu
h/XZjq4pKCJYjX0qnj0r6uxyiKdFBnOpYcKT1s/tvqdeno1ZzwBHWUqRdFvff8pXFPV2oYV6hj0g
Fa2qyEcU44pssTM/sG8S//zAhaS+J6nSXabDszvFEzJSdwlpiaC7FBKdxZ0zlJxyhYsvZBxVIx3s
yPLyNIDNo3uWPNCJcbEgvUv52QwoMPasxUE5vEssBLFXrRxNlO145k6lu+Sy94icu/M88FPlfVVS
tuS821KNUZU+Ks6ysIAZuYHF00LochIPbzUoEd2vrunmSMFhUP5g/P1n7kggCxULKI6v6jAMH9T9
l1PEt0W+p8Qm3wC+jnUUfV7kbVUOfM/KH5LZVcqSzq5rEiIAuEeod3/MKEQCR8o9L2rp8jEnbBxw
OzM4/aE+m2/mprPdDHSpYMA/1NvcEDwLRq6uAaqck5aTB4OBNMNUkXdpkD80GyEcPmoJdmjNxuoJ
VOn/Pqr3w6gN+ufqszTkNVEiqX1DZOmxARaFAnBzL1uRt6xlkfEfqyGodaXUE2sbbFZmC9pDFroU
e5qeK4dc0OamOtNNf90GZ7D1l7tVmVAoxhN41WZisatRsVgwALBVQR/DxlyWgrl5Q2qdJh48OYjr
/nxyxECdD6Myf6KZxVPhYdssMMBzJ7WYeXllCQns1IpV0tJJ+y0PNG6Gk56SJlwpsvDRS6WRmcIB
SyOemkW4SepHf+qFbxrSL7TfizhA5RfIQa/sJhWuoUwFZYGTNl7kvX+peuF4t46g2NayQbFRiiUF
9ynlp7TFXKak+8+S5tHnA3RFspCi7GiQOPWijTjAUrcCHLadQZEESpZI9IJUfJvt3FgohtRQLat6
9kKwPQaZgmAGVBVjXppAMqkQFW9lLr0Lsg0nX5vwA49wzJSzLaa+1kGGLVonayFO6bm0bBKSJnrE
TV4i0FNy3i9tb6k/1vN+Un3gnVD11mDvnt8fsekGUQaa9VXpLJBSV9afswq6et4XHN+Fs1TreepM
x/hgkm1VuAmuNlbvF5Xm+Grv3eFCH64zvsVyHhWNUi49/hFT962cYeuVH/0S3CZm+NHT4dQxop17
WmT/EGdAY4taMsLUVx3braoAQJyQ4VTLIL7rnON0fQF98GuPoiMpE3YwsfzFYxJPPQ9PakYZhqCM
WUEd+8Gg5zCcA3yP/nhZZyCIIdIaAow220peh4wAvpVwzT9N4IeMKruT4HkfJzuz5RIQA1ki4Zkm
QzEfsAWfVMfuuQo+ioxgrY18ZM7ymgHY1/c7Kx/mMhGAdZlqaTeFAYInwvP9mjgm1Qn3OOeoFO7Z
8R1CfLHoUAGarjI91OIDs6/6weewQKwnGMeJnY9J/hWXbCOHFFV+6d/8PDKnelw6GXCPH9mk3w3x
6qlvPRndYGhJ2DBirl0+iQh015xJ6/1JlyZUqkk6ZiYQ4Oz60L93Fok1y68q3ME0FuBxq11hOBNX
zKTpVYIEzjewCmMDsLzE8lhKWBggVdKaYFtHqlQaSaT4Auv+z1+cR2K1PY3uLxi9dq51IZruvj1D
mFXYrcJIQxQJfs03R1hD5o1UEQUwjUJj299xb10tJrjHGW2ax+fv09YbmHEJ4JOG+PU8xP0ry1IM
GYJGdP5MM/i4s1XpCO+x79pkkWT2dpay3mOxvF7FDoGmS/rvijF7X66fpzgph5hzl6OfYhEES4K+
UuTvBYUeez6R1N4Gzcufkcpr6kg/PDnv8mgAWm1iRSviBSRNpyhmNApSF9u4gNbZbQmWa7vSyany
LFCPP5qrUL9amg6UxFviqBKvq/PATjsCcM/Ocr8mmfS6MVQ2tEejveJ/lxr1T5hCHkjt8HSjYYnE
kgKJeeII6dLwmTjyDsJDelI3GhZRlVHISDH62LOD60ZShsEl2pWTRCZVaskiybuxgxDT3S2t20bs
UMFtSyUWBn+cMNRO4sm8HJgZugGb/P1IFzxQxluH967yy24ns4K0QfFqSm6bwvFq8rzZ2U5wDf6x
7Zzq4ssTjwmHAR6CYJOj+btpUErMiQ8Han1zcX0nQagKU1SYvvcggakNrSBPSACyOSdy+rQCaPGh
IdtacKslhFndkwrDbRQPiJuBBpMp5p6oznAeEgB9yoKVtleHLSluw5Si1RA4h8DRiamDQvi3lPw+
MFi9Fur31yey9oy+4f4rnjj8p8HSEJVvkYgSb5czsmR4n/NZDKG1m/nV3KLmvtKRCYuaU9gaqadW
kAcM0Hv/PAqRsA/v2XGknmD7Gw8iqQyVpejYCAGyKC7K7hzXTio5wMAy0NQ/0pIbbBVKLdq8iESI
vNTSA+21pBZlTQEcdDC6ysiqoWyXLib0LohnqxVrxBM4BH8TYNPPM6/LmL3hZNxU/EPNijFZWTV7
KsEeI4DESF7ztqLPm8n3F0ixQCegrKwMy1gBLfRHPtZNff8C8mNRbd24WyojrhmvhZ3U/bY2HK4B
GyQkuBa2LnJNqKq5CWd8JAA9aZfMdnqEswh6SL8DGeDn/gQ7UnvlhpiTBUwSruvHwTn4s6Sev7/i
KoRL1pEnRstXg5dx+UDIzc0HwMFG1CbLNkV//rsw0H4pktbgRNmkgIMDt6sdOnogKlqd3xu0XmYl
KgauqxiPTpZVeljdOpA2dxquLfCymBKRQPCMNGupvVKrSPeV6UEIl4oXp5BBnEEj6+1lowz9cM1H
mklAsqBK8Vm/k+iRPr/ifOtzSnCJZ13AT1burult5JYtRF2oKLAOAGOTtf+UfNwU7viYwTYaD191
ls6/ZBj7WiMJH+ojSXs00FhKPzIqp41kV5wl6T15w9ddpk849IQLcBzIphV9DJSZmSnk/B/dTBwc
tMf7l1yvRU5IDPGEr5IJ3/ZgDpdJs5RT7PXymhWX4nH2i3AtOMOX/HFcH7oIh3Y+YV7PrrfMtBUH
1av2DeKMIKUS0FhDPSEoAU39lybsp7Ziaum2Gc78G295EB1vuLwwzbUwDd6nc9JG1291rYGe+Mxv
GKKvivui29Qze8+9f4yN4Pj1FJLsId/c8ZMXOUysQPTcnW6R9ktXe1QqufOBREnjaXWgbG8Lx1kF
wa11Sl5KBeF0KSmOGrrGg/rrIilP01MNMLS5wt6nROnbe9JX6e4+jsUGJ1mx4mgB2/qw9+P6z7ZC
UJGD1fQqZ8q2HwEGowfU9gJJcz2nkbAsG3iusiNZMCG8VCqX2IhUx0YMZpnAj+CxBrtzKApKqvMB
M2mVSRj1gTMww02VsmjJXbgvSXPMzg83iR/EflcTvjggRTLHWhDix987aTNtec+yiOVtMdGGlGPP
BZGZYfGfp9MAOA3jjv31DPBTNv+9KUf4V+WoTeJhSEAAHa6eqCe/8z/GYgdexhfNtCG45yCq5ryu
rtkRUEADY+s1woG0G+b2e63LUBta+P6TubiGpgEpq7pREZy2Orah1KiNfiKjRZOE5DE/p3M85gui
aKmRABQLITLc3gupoB9YDUC9LzugIS92TVHtoyBfTLLqUeOiDYvg6NHf+jW5xWzE1ylKP0YflRAO
CYVL7Pr3Zk+yttQBuk1USLunTvGSRvZ1huWo1o41nmLX9Vq9A5nrAIwLFOtc6QNoG1wEMvZJLtiu
Q9ovtr3E0yBld50tDf+oNtgx1TdLSbSN2AbPvRgDWZ34XsNzVeNCof3y8n9bhuvxG28GT3aXSjo5
z7hOIe8FV4A/2vDzUCYwEOxzHw8du7wAjqQpOOyxFwYKeFlxy0kNtFYDXL7fnEGu/+cxWAW39lsd
jvIsYP9NiUIfiNyWt9ke9avlalGIZDxZNi0QQ8Jrq0lgKVnC5tcCudtYPTgoxmmZkOjHEVgkyRHR
yNz5Up6dQaXfkcB4tBUxBEEB1GUwpL8jyp7SuxdpTbtFfo3fapHEl8HlchAnGEnojLtQ8yUYbiTk
G5nqOSOq3BK/ibX2cc9IY2YT3SnIrqFDBPZttk0jKCXDlPs36Z5MrKfSux/9za7UVQUn4PeLFqqN
qFKy6v0bnjHTI+NrCLfTbFnsDqz8DeBCHmvRd5AYpAePlgGzmidT7V159zS+2T1D1IEjmD6GicVo
/9km/GBRFgSqfFpxi4n4Mh7b2P+z+RyN7HkYyadP53eGoTHrSspJWbENY/eQ6fDrfUdAQV16JdP4
OwAtvmsFa4Dn69d05kBT5pGgyzrdUFnk3Y7qVwLJ4nNlqA59UO/mYL0b6G/GWylJVvnH+98Gb1JO
8I77rc1nUR+f7mVptzMbVKDY2W6mISl8jziGLfXmlsR6/AzmlOIRfOOyyUbDO/ulhE7RmsYVg2wF
rlcF0qtdeub4eQjr1OSoBm34w+Cn5GwXG0VqVAkNku1Jl9eeyaWJSuHXY0evBk6Re8lNuIGRKgH9
L8Qi9Z4RB1q8kUBBzOKXme4LQ36V84zy4zIMy3pVeBSfIhKWugSK1Pzly5DL2wJyWtoahpfKYIUs
+wZK9jtQvAKviYWVY29Ro565TrD/nbRazo9VkMiT4xX0DVmXMUoNYfltoc2yFLsZJ1iVijELRkW8
KHHW2NWXuX+m0kwb6NwZpwcllB7vqlVp1Lge271RLU6wsHxbbPlXbC7hWeMJ56peG3jfAORZDgeq
AER8sfdfADDNm4+LTQsqM1ZE/bkdM3HyM2VrnCokZZdVSLPIpCHEFdFQJqltxqYeGBxQ2hJzHxFG
cdlMlbHL4c3SYnNPySNchQZJniu/+JH8eyBrHE7ibJLM+gpZoJRxUJiyH2JF0VVVojqml1HuYDWs
MkSPTS0LqwN2TiG4mdDrJFAx9SXMFsGi6WJ6RCbcf3AjAphOkdOvEKxJY2q3Eo2BtxN41Q3v0QQQ
s1b6r1TN4HcsveKYAvBogjjQkzpCM7ugJp+gRKdhSO6cRE+EOvpAuYwz/c30T0/nISoviIisWzPo
CeJtcsjxkPpV0CITEtJ9b1baWL9t1cNnBdRxAS3Qkd1J7h6uMgUYfm54NWu/kh1FTJ+OvSXDu6Ou
7hp9Rhr7ypdlYYpcA3SFkMI/+1TDS4dZfDzDMkY5QZNgzAfpTbxSWPCNntmC4WTjEtXJqGx7EzeP
ianf/Fz6C9TG9D2QFdXvZjfkFqUC3BM6ImY23IO68srA89avSGLpEO4JBbPyVdO4ohRdYfhPbTXW
rxkFYBsLR6Y1dJtaAzF9axFOyFObANowOex6rd+/qa0R3UUCWCvhLV1MhjCsRG4s8Q4i5Hmp9Wle
FIVxRnU6rlWtZBk2wKrJWEEfl3TUEUwCA0L1bQSuNxbu6pttoY12RrG72DxOoUUN3moo3znYklUC
ZWd39o3hSCL7M9gdt/B/iraoX4eWwKY9Ovp7kvCULcvz8WZhVpAMJvXl39hAtB+xYVckBeoXVRfy
F3p4XQ4BsuR9Fvnmjur0tmbBaiZQrxfzzQ9IognXye3EURrAexTyiRBNwPmLfyWcQsAJuMduZ9tH
tOPGoMWbxu4M18in2W2cpcCQRZ8lkVbi7qN12IWOjd+nqsLzRJBco96YoEQzNSuf8Hv7kWVKQQpA
Z2Rd6H+/3TarG3KdODIgPFUCzb8tSpqekROak8hSkDoBQBd3jAnUtxx4zUcU9r1IGkymTtxb7ghl
+EJX2egJYAhosHgG/MPa0hyWmmXGj8NE1d4n33FXQ9rxsIFnYWCPP7NX6BJuXmrkZoKfU3hyvRp+
FDsUAE1yLdsQbVT6gJuInaDy8tdmMTIQws9Y0BbjB9XvHuMGsIAAtykVnZqOax1pcNfaf9GNebOp
JXfwlj4TcJV3tUdaUzC/LItbPz4NjfCGzXH9BYyCee2k4U1GrtYD/oN4SBOYR2kK57Kwh6/ZAuUV
NQ6DfyWIRYEAGAo0rxp+jRhffsgS3JAV9S0QWaApFJvwrCgxe9CGKN/u7F8aE9VmyHWIpmWLD+pe
vM0MgIjvLHuz3vy2r9yNwL2E3N/sbhaFlrKVLDGihMSJGGKnizQzC07shPBCfb1HkZHnHnDQtgA7
EYk+i7d1KeBAJv/JhIGZwTSSL2X10CEq1Wa3k2/UR6CQFge8ZboN/iiZH070/+WK+o46NwrItBNX
pkGbjcjoBs34ChA+ySdJcYahOvumbrp+kQEW8tdRJWz+NVlEXcq+2D9CHxT5FUSawiTDhFfdCmah
cOkMLuj96+paGaGM+VMb/5I0DjbeLgFyiNzPTx86tnSDT/9t8hZ52+r0pTlxw26X8+IVlCIe5JwY
PKFSJp2Z9sMQ694xvbC20JlYn88HyqvFliR4jCUiU1jWHrs2pnPXAvgdc5x/I8EFX5MhtnUpWP1X
prOn/84gm0RKKuQJwIdY04bCmkPmDXGSZR3VkSYCBXVVUGlWtCvchQuZJw3zIrSkdEaPmOSnU0jA
4Vf2WcPu/EaHJ3gWIXo0vsc72et8VUiHBk7QeP4CMqrSDuIs5KVySPjx7WmJAnWx4lx/HJ/SUxU9
wibAfG/6ycPYAvJ/ZOQ6fE3f2RlfUprikihVKsKT1hDfVYx3hv+Olt29lCj9yNqCrpLmOtLYhF1Q
vObrMcqRB+Y8iC/pn8cHSBQpcEvJfvq1acIZqQZ+ulK3Ne2iH6hpRDtslKW8zQLE2LwbjWzJrsR7
0AwnvbCFwcWFjdpIDVH1SK/Xg222D4bkG3eDrw2Nvopb6O7IJ49zuKFeqTfW7hGqjBrjQW4WOotC
sr1rpmSyT08lD3aCI3MOPAB1tpzdUOf9MLFR25HEqwWhllxvqASCkSEvgQ7+H4JoJXPiREkrev74
MT2DSaRbUehhl96yHV7Zem2IXI4WjqIHhESXut9A8hwTrJhtwwmcMj6I1RImksGcP090rWE6kLMS
e7HC0mEz3xjgYSSYizQ7iuNFA7tTXrpPYE/eW032Fopo1LtdsWrXGYDT2wo1tARKLStSqYQHbHWD
ZTfLyVzQqrbKKZYUx/NtLtjrua+1bsVNOE9FGqUizoUtwJUnchQ+dJdwoJhKFv6bX/IZ30DhrT+s
0muU9EG3A3LYlCv5eHwBv5CRyTIYHbLgOGpa3fmpJDux1NYu5pLee3SZ7nCVRebRLbHCBomuMJbw
s4TsYrVrP/UmvU1kc1OAi9r7uKMhuMl1umAN5KetPnKIJILb54DHs/aL2VtcAmnkVUhk2hYG1R0C
2M6DTqo0tBwKqloLd8OUuHt3JjgC2zjgXXI2XfYu9gyOhevYcuScRTr2aA0ubSNaGZTd57U3jilv
c3iGGG4LvYhhXSJbctjnCaY8gEOEWfwZM5KUHbj7ET2bJcmZdO57OTfXv18R/lFSp9JSOr9d92hi
lbpnALKQ3x3r7NQQAKWNHy/MsANs/Q+uKLDcxGoV3UipeYKmfAeNHj0WikQTki22I0u60vWI3M8q
F8nl6/RB5hmTb/JigG1wFh+Wry1pN3Ot9TKEVGba9MT5DjhDXdxUnIDGTTuWgmabUjH72lZ3tjcU
REqnWxZ6rROZDDI0pbi/nQk/J88HWwL0luSckR9poAfuxfMxRsiZoNi4nFF6T9irAJ3YFyWUxiI9
EMV3WampIzSwL5XFv6ZTn0L25bj8i11kobEX2BzBChxWuKu1olFEnBsCC+r+BVTQ6+E3i+W0yxyX
Fo/Evn/tZhFtZyqoF709bQdvg8CLfJI3rEVL+WQQU+BEriTB6wpl+pU2MTHMxUYPxz8WuxOgeAK/
+eLIIq7Tmszte9ipcs5Ea7Uluu7TuwyLk8YSkYtCjXlBHCwx+u+dNZMb4dDaebslOEZpQPUmf+w8
dkdsOcyhgkGjCKTofsmdZuE68IaDEdjaGRb1oN9bR+mDcvpQnyakUM4UjKgO8tHFGwYGfPELwegK
u+iDLOc8R3bWppJsZ/vkzz5a0/in48CuQWe0d4FpuGHhDnJJfd3z1Z/e0hoW+2ZTAsL9BSSC2bLJ
XaXKo2+DdN79wGjLIEje5OqIQpM0fIGWg9ms2qLb0v7Y0YsiwL6SxzHNfs0OrbhB1LEiSMbEtzCL
TwbTTBe1sj01xqVJygPudd6M+tOgpqcmW40E5KLL4AF7TzmcWU2uPcTchfg1cX0bYDWdz3CeneLZ
6KV9PCCwOaY8MTMlcS2DazygtaWSwBxGrKxnQu/dVa0FOM98jVP47ThayYKFh4M92ZlZGw1qeZgA
uyIg4K5C+LtS3GE5ZCukuHRWsDvIP2EJW/X9wBwaS4r8ENknL4g/x1xoZnoUfIw7a8BWnhNthy5M
zk25VfJMRtZJt+o1Uqz2HQeZ2RRHpdq8aiPIUrtojotoisvepGE+ZjRaBnm9NJEXnhUI5N/ToAV/
XUXcpK9rNS0HSmsN2ps+CEZPxqTYJan8JLW4LerdDnqVCulqUHRkM7Zg9snBOjCIIo5l4rfJenBh
/dCuERy8BHaC0kYZCxEJCCSE0DPaC76KysYzrg3mTLZ2/p69Yr9uleqwptpSZM/+jeih4p7Ydtvo
fhWt9DBNKdcJ5gZs+wXhetrFw7Dr4EQBEwAtHmyAKuuzoWaoxZmSE0EgqoPQWVl0MP+y3LrdrzYG
cdOZPnDFdGZ2ChOmFEqEnUi+F3Niukn3mvo4sjd/ptu5VjtmVTOhnaRt0L/zHpvkUw4MqBmc7sSu
NJL3GZUcyzkNuilPCFnS0GkOkIFrZBaubkReINJnn4DX070UvJBZDYb/r093S9E/9+dHdgwqLwcN
WmkR7cvHXzjER8H5vZw/Yk7npr9PEd05+gTyFYE2/kP8j0/8N4t8Bst/zOrYetS/3OHLNHSTknY6
x8TXl6I5yS66J3g/9YYhENvPtw7hHScsn43GVIR19nahv/bKEP9ioWRZ+fdAZNHu/zrMHZ7kjQ9U
2Zr5Q2rBdxHL9wBYowFnbzUFLgreOqIogBMRGC6sKxuMDlv6H5H+2V58l5Ld5pc9KKDbAR+mW4ep
o97ONIx+iyGxY12tx+P1kHZ6a6I9D+y0Pk5kUYi7LVIqp6/R6B5ttuO+6hZqhHckrn/SMx1juDWp
pMorBCDwMQJQwsWZkEOkD9Y17s9ZQC9NWLvHWt0Nuxu2XmEnTXDCXg+QJ8rY5GDpZinHWYiGDC8O
aNKiGj+iQSk5ivRwMBX7pxMrmgw98iaDxvcvq4z07gNTBbXfO4UszIx72KDI0vW4r4Mc23TqAw+2
7ymUVSPR6wtCwZzwON8iJ5wCsuOxDof+N9KWLk2GP0gpkPFb0GMIV4axBzGRBBSKeh4prkxY871W
6Q7kWzRWBqhPMrJrDTiQ6kMa10IbAoMzeIGA9uQeumDhm2Ga3JyALBxn6F8jyGUsPUP75s8Oj/Uf
aDCe/HMZ9MlGIAxlh+eLnbvyaTPUlYbGBQscNpzx2PQ312HbJLpZjyr+ZA8IoPNEFQIZgHGjQWls
kq6ZGle/93ayLcJ1GCrqfK9Xw+dy3ir6PFHxROMgdw5CHRNN99h4GlasZQA1XWZ7BC0RjxMOViM7
D2qZ4UyDg94EtVyxJ86TJ/jdvtDeSk56Tqep7Sc0JdAMqtpzCK8KRpTxG1DIStCHWjPaAkSe8DkJ
slrFM2Pmx++4Pyp4hSRAajvATJhwCKn2PJXlkxNUlu/m2XGQcLfr+vfJf6IeW0T5ZY0SANrriZSp
4UKDeWni/j4qOaPIYgIJqJYEQL/n3h79rF4pqLl4ToY5B1cHnm4e23LBOzczrytYRky3bLEj/Mel
50w1DUa6O725On/TwEnpFGdSk8FRjDvmARRvLTUUfAfkvYRAxEn8Ru7DiUaRTIhVrggoKCA7b6X5
bbFdqvmhaVfj9dfx1GaWxdUVBH7E5kD1QZzaMeDnmIWA+eiw3axx6M9w1L5Q8AIWloiJ21VbvrAi
D00p75Kql0aEQINtdtrE1MzPtrjUiMqOEA0H5RsRrYocp+aQPJMKflSr4AFe9ws9T1mniuzhjc0n
eyyYgG9CIe1l7W/f/Ax605A3ugry7wPMlIQiq93eVEseLpYaC4nztCzPIAZLLvwonVHOBZw2wtxn
neymLor6uqrTK+FwOy1BExVsAZBYEDHHJesTeXIsqePbPdt6NkDzvH2E9H2nm7BdGtSEVm12CVlW
zvBR4mriGfqi2QAcE5/cZv+WsScutcJSBK+EVUNRgYUcKIHR81VaBv8vNaapY+mJDUFirodmNG/7
YP7MPfPRCEZf8kh9jxAMQnwngwlKoo/dpn65E2uxgnQ3NWR7w+UZsFn2RdpI/rIOyjdLUitFKs27
HqsJHSRq/FcuOvrCkpWBu8TERI0O/sPLuLok+hd9mRWQ1/WTmd/PewP4S+Cx6th7UX5CJa5BXef1
xBnl2cucV8mmTBfyk2fH8z1R2BgpBDsL1fR186M/l6COcalmUx7uiQFeR7cP5Ta3hdOQfPsB8l7a
GtjkOxlvXOnc4AGOHhREzXdGry1Z2gdA4t3a2wxuozYSgMgK/m3Uz9aI9qf/EgxJ52QfJWOKM99f
mcO7zzP6T4pI9djYPW3ioGRfwZ9p8GSViky3Ib5XoJBAUxoqZKf9hD1yf0dACX1tY26C8ykhnycQ
CVOk5ENb7PCLBJBh76baX1S4etmZ8BRnOCZWlHgt74BVV2rljBidh02euWy5DC5RYoBLPSb0amRD
EB+vbrUQ81vczP0BGoc+Ht6jG2pNsaAomqe+o2Z9zzz+HJCwYWXUD+Cf4oCFCZQgkqXEYwSP3VuR
7OKpswmETUaWNvfjqSXNHBSA9fyYvhdqqXg7uxaT5ws+ztil64RuQ3WWxCXQwTiMdknpnhtRtry7
KGvPoudA7QIB1FbKoCSlP9HTYK5vwCdHw0trA9zMXDK7szK9Eeut5PwdTTLQYrt9LcCjLc38zU8s
H//ctzGYhA1qYlCyKshMaTfsju9Z66ofbnOSE1uEKnMGUhP6EOvvct+Kwh124IEWBZqziGxlywTR
/uUZ7dZxI61pej94F6ENeL5gNKKJjKLjbk1SzFdBD8kNp1TwcUB5/ESIOwwCJa9zXf7gPRqEXagW
YjaIN2Ck7gz/sMPBABiMvuCKkZnw2bagjeWhAOoljnzpcb4NYGHbbRaIdW55bL/i0TdOqM12Schu
aAuRJIm9cHr2nuSl5y1+Y9VbYF5C1eOLgvwvqwJcKu5Vp6MQGHlx1ulY5T0IQps4xwQra17Z+fjk
21Iwhsfq2jBWm2quB+u9cyklLO+zvo9ZAmQqDJaUamyLMIncsqYEswBxRFtlCWyeuZq6zIqAdTf2
BkvgmKK9YRZZLsHOyfrNlPqF2DhTdbNkNtJL8035SG8m+WohZt6RN35LJg7Jy8t+kWh6a1eT8KmR
vdBIWSfTVLqFQPO4u3Xoox1yiwXpQ21WwBYcgZ5Z48zXdWG2uquZEImfe3hrLfi6Qn6UzJxK9BmG
qd9K90OEchZvQw3qvjgkbmWMsINp8Sjdf57J0gSEcuLUmfOQk4ci5di9jyVifbkC2RHjL9Xrqd8h
TKJa4JqcQMWeWoMHVgrb9EpTjoDzU7kLcDyGaG8QZB287ksZEy4Iqn9cT7AnxGX2ieuAjvdTuEoj
xZvSfsNOEtuoHhNWDzLtX/XEjfjw8QPVoPYAoK4oEs5ZNBu29XPoJ6Ke8y/k9rI4D3D1td21MVFD
vCp7HcKbwffvJT8iRhIBA6BY4dNOBRvaZ8fjoM3LFYRgWS9L1JimaVOGa+yKl/5kODRG4ZNdpyWK
JExAR1n5sG16Ku7o23ecEMLQLhbB2Z0Pn/HU5uUq/hMglQpcyJgV4/kWoAHvhgf9wJbpoGmX5wDQ
AnOK/dEsUbSNXU8TJebsHFKxd8D5IZJE40z9CQApv+8fuLWWRr/NUh9qvnbGIyqIp0H32O4WBHLF
mhDqYjEaj3TmkOTE1AfUVvOoAM1nVAwUqpyoHz2xtlmxk7hvnMVm/sDt3Zw7g2bFusZN2aaxB/az
fW2k6hQhxdqCGb1aWIEaZuEzN8hEHPgAOHbePz2c4AobfLwOHvk68SSJLLJJuukF/S/w5mg5aOA0
aYlylGcDD9f+IrY1o1F1Z0DXRah4SbXl02tgMaxF2n5mePWvTWLCrwAQfw6PRIA8zYDYnKfr/Pfj
tyMjSpYsv7tKjwIHkHyvSe2ZZELi8kJn6sLLUeTHEZGXqiR5Lk3kCvIj2+vAVvD/K7tAiEvDk9LJ
NnmUxMRW7JGPeifWSnhGiAXB4+0rsBdKFsZC5FiWgYiYatFG7APSZ3MJGczsie0ooMfdD4ogimQv
o8/+EmH1n9eTf+OEsphYr67Q3fHN0wUrYVSqQzdPRsl3Hbnk94BcBekTdaSyaOAZ2sSRK7CoC84l
oE8HB1htCsul9j+kfG/ycIokVYkW3ZxZ34Z5z3SJ030QDmyM0eixObxiLAsT5SBpJoIW+AV1llii
K3SvF9sQv2pC8ehQcx4QJuZJN9vsbDZJXfTCEiQPq/O1/CAGZU623E7AHvkeg4fORN8l42OmgT2o
xlLe3nYtrSWCeCaBY6Fhz2rxlYyNkjtbzMrEjFtFDT1uUN4JPW6SY/YjhhFJZWrZetRokMzz4oI3
nEqGMmQCji6H4AwtQZr7bCuRavm+Gf7v/SDmn8d9SvvpkrYH6SeLuq+smjYcohdMZ/EgBkL5pG7x
yR5BVj5PD9ctQCLgcfx34B+dIoHTpM8O42UN6VUQ5wsU8WwApDvOc29YnY2VOYbU9whoijuhsgUs
dgF/a/zqcnJTNYmSdKrBMobqGKF4tTEZda6wSOV1dnyu/+G3nmKrZlfaoo5F9SzCRjWS7uRXNnLO
5LNKXewOdBh3deQFxcNt3uwZUo/c0NnhnAu9ddth00CCpFSjp99VvlITLBW++CLRLrSxiZkbfEJP
euq28amXuXA5omNm+81zydh/zkEnt1F7DNyFg7V7kRZdET56dYmku1q+zmxKknk7f/bdOJ86zSnU
WeMWNnGuXik+SEx6NAUnUz/0bqvjHAR3aSTtVvVZ857b53LQfLzNyiuUUZPvAvko+vBpdFNmS76z
CWEtbTRoNnSkKNmOP+ejAXNigFnI16k+zDQh0wIjr4VUPnsDo+lUX4CWwh4oy/2ebl+1qOPXzp1h
Qn+GzcsA3ljq1pAYnHuVtl2PmpK+b5GhmVFVFI/x4SSVvQxCnw8i1C4K8+0ETXqbSCx78igMesB1
T06S1u8Fe05aiYyLzEJEY7Gr5Rc6h0RsTHeDRtIhfu8hCR2dPrSRggFGBpjadf+GID3f3GHA3j8T
hRaCglUSY7SZDNhTkn7VR6iwYmg12z5Ebk7efkxeW/WdpW2WB+d4InbRzf0LAcG5sbXyj07rJ2GU
e8nnpkydo0iREYEc21+5fsjw2bgSxMW7KyNnw7j7I32DmYqoev3rZ8vgYnKliCTUdN+IFX83Nt59
UUCJ9WJyQwi7L+/Jsm8G7gmL/e5hM09y2WADAKXxbo/C/OF26Kv2VymcNkxjue82LO2xtZir4kYh
IkNP0M+9vWaY3+oGcz91V922340oEUkB8SyxjMNrmpGXeyXEgU0RarVqZ26PuhvGGLenIxDD3A/4
vMQdWmUMCpXqbLPwepFZ2lZme6HNl/GZMYZgRaBlJCMpru9+07EX0mT9qZLAM31VT7KPpyU+JkOQ
iN0wWArwmgQ6CusWE3QQezcekE4gvyIdgS7Ruz2Rsbv4h/88TROi1v9H4Rq/ZLyrz5QGqpIZEJHY
w7YAaKG8yASlIGj9gcX04VivWBrZ8x+ml0acwzfvE2iH2tBPexRY2hVNA1MVejD3NQ0Y1mjsdyVC
tqLi8bFb3CDmLpu4GqEa9wmYMOWvVrmZwyUDtMKFVIOTsDpMujEytD3AgvM0IHPJglRShsnXUN6U
Y5K19WDbv87Q1d3fvSpVSXNaUuY+BsusxIjB/IpfRsA7pyTqeYCOABvwN7ZXWbHzQqLitgAhga1F
QK+GJolDKDrabecuHLmL1uFirbfxLDOzQ1nRUuWJQj5cFLfany1bzuceQ3c11GSjnUqQZ6/CYIjL
QbUeFudPR1MhcnsmXUjCdCySgh28A6gdZhj51coF0rydgPUo431zhxKms3ops7Fd5aKJRV+4W089
Hbd9LxnSdG7B2jDL0yGraica+tPZwAkhMkzecg5XvhMqq2OpuTB41wK8EX2aIXX+gxWzPKh7/R1O
PJreuYDyCaavVE9UIXVbDcr8LP010ib5W0ObP5Hme7WKwenuQdww4EfmEgeF+Bppil3TN/jjfdtr
+nuaDSMhYdk130RUJGnk2zuaW5jvnZL9uuBmCvhgPJAR5IgXJCRUkyA00JpVr21xjeYkl3Itn93R
+yRoGhymZxhsXcxMkoVK/OyEe1PKMI67BLDgI5LCftGOkMXhlNuKGBhnRPXbxZdKrb04VpNZxxtE
hZ91jmTNBr7s71MP/MqipYDPm71X88MCZpQl6wWX2sirbyofPiQ9cgITAJqzCKtf4CnvmOygBtNz
Q0ed6cd8gv9HEMXik62X0GqmY+ZCsFs++mnaDrtnf9fO1BnbiHktRgCMsdjoK4xYCz/CIilCotaJ
8wyrSc23ZLdpDACa3OUqT0RdXK0afplqqbsrx7mG1q9E5Ubk0PYgInqL0+D3qTZ22wKSBUOxOzhX
uDziGpcEjtgRCT0K40QJUb+ojJtjYjYy3HJqqLgj8/frOGFauzMXW6/Yf5smys2nmPgDrYNXaC4L
fpYynLLn+LsXBHPn5UP6u+Jdh+TPdd29keISulMbxzYadLAhLaGQQ7oIPQ4W+psxq0ETeXyzszjw
xHKbQU53cm2Z/SJaDj2u7bZm+GyqScWYto9MOpfkvdxRrJjyKw8ff3G35NFeuEOGWYtbInUGyGqY
wAig8zHBC1DeIOsG+AwBOU8DqviV8RYUeHPgELZWiy7Vb3QkgtEERfeP7tVXTVIOo/V6rpV6sVLm
CyMPw7ZkqJd5cSaxN2fITevNFjXkksThCvDTUZyepJODiUfy67vwJteLq4nATJ3sdgORqyM0xWXf
Le3ku0R0nE3+2ckoKr2yFXPmGOCW1K7/H5tDiFwh3FUmlxkXDt2AAQ4sHYjdS/PBw1HV5eO55OuH
Z2yN7Dv25qL+QezykkY5UzGOQk9w/YDNGtEn97y6ZqvN/vJkUxMhKE9ul48xTU60W+Tc0WQAbrID
Pg1br4FJyM0uyy7slPQap5tj82R7aRX4a1XxSnIK8muaIq+9lbiqkxtC7j+PrsW1U3wTLr0eaMdp
/qfu/kXLtUM20DjwkJp5U3U5md/yKe4FaMEB3ipnZlq4nlmNSFb3WAlMKly2vSJjHLr0D3+hWvs8
+g9ZrrOyXiRcuGrmU9vzatm8V28cUIKetcKnCeP2fNMPWFymAx646/CzY/mbU9N7HeI8V8L0GF5W
YZRjPqafn7uCKiu70t9YGgDnnvL1xBNKGUIUDF8qrbAfsBCCVy4rQhOTE+RcsxhriQwLvGAf3Eze
C45c7c3WguZWwok20Haa5zUdCk1b6LPNDH7hY1fICH4+364jv+GT7ySsbY1YSCz4fTBiwR+1CnYY
Hhfc2YqSdiDbj/jlbbLr2PrGmuPrjQDiZdBghSDn3MJFAhPsXHEnkUbP7gGN5b0Gaa+vkcZ2ZB1W
sADx40njs7y9CJBNrPKiBKNLcvd3pE5+xlqwAdcdEKmW/v+7djaWeCyMspQeY68JrXo/ua4fxMie
lLsghonMiy248YbH9iM+s138LE6zmd6TjPbI0cC3inDUSkWy2/8rRKsHJO6/tBQkASHsqzSKTMk5
LBBg0+idzQYKqR5LjJ3qzasZ7GIojjCiC9ipe+R9QTK7EOJjJ7UICx1ru2/GX0Kzhy4lTyFDvRu0
wi/0amWyXEldiDjExAwmF8+5xPcmLW9ThyO4zQQxVSeqlTfOg2xkwzFzBIjvIfn7Mtiu+fUBOjyB
wffM7zT+yDSfzR0AIDgaDT0aTsRtQOkmD2DVUypRhm5/qd9qgjxu6FTbCytSWpt6Y6pX6WUQw5l1
PSATZe+nYz5a6yB3ESxQMSemKt4/GAchPx4ERM4sqA1HD6SX5DISTSC0ny56ILgRBPwifrMMgPeW
UGWAqjv/AoVCs7WJ6p94smtUROLxxAuI6RCnQNth7cuft1mKY7Aonl72x7X7UdWfrNzPA8p7II31
KdKKufknhFFxlkGof+/isN3YTaLX7x4ex/iMFkqI/kW4nUJlCylBWLOroOadUi062rOXz/oR1Eta
+PhRrPLKKxcL2vuR9tV0605cIrK/L37OVCn27i6AVcD8FoRpsoMM/LfLHcHIJgNTOrJYEtZcPPm2
jOLMGA3M3a90hpRmq6b3mnb2a1yQKrFi7jf9MUCqov0xyLfk6i3OSCshTXi2+ay42hCXAc9mu72p
ekTi4JSkvuncNW7kIRDPn1OkYth1qw4yzF5Y5EvjU0MlUzU07f5XC8uc5FmAHaNHwORcMDp1TQci
+43gO2KbpoBzL1VD4cDNEOm6HDRUfguQr17qdsMNQROVQ4Vy2EBAw6tegCp6CEce57F+FTy3Fc4E
3nlLriaqil9URFZM9kuPONFXyrludK4ltWuFe7R3xhvsbBYTCRzTMXUU3fSLMo1WCOpfUesSDqJd
Xf9fMS+zc04cicnCqTI1JmZ9ZBE5ahjeOMWOHiVMWgY3f135N0Z8tZspvErnu+g1t5hLaEqUHRzx
NeiHsynpu8WqR8xR6M0LA0xDVTYXiFIDjWlgjx0ljZ3WTCBgNPcUlvaWiLWmRquQg90lUL0C2bzI
CnWL/ZR2U3R2UJQy0BDL+eGGE3b+M3k0dwfVNAH0kWFWmJMj3KwKIF2qUj6+O6a5yMeXsV3ShbEl
8BgaiPSznIXKprEwT+KI1j9KxZFgeWX497tlc1uqOARc1DOrOUKvz1tRWOy0DV9C2l9on444e2Ev
IDR9QIpqxW5f2GGbfJtQsbZUuS24nUxl8uzlLjM2u5RFwm9ol9SzpxpB/9Ieluql5iQkgoTKHWvy
TMPoO/XKrN7cT0gNZJeqaB1UdeOohEu+8JS3BqQiq34+DQLN4mgitIfNIk12lrissjySfs6rq2uv
jsY8eJSiYFzzmc51kfzbUQqbO0xDjrdywCVH6vzLmdP8PWrNNPZkujS5drU7k2LHbY5srZKwFGhj
cAZaiLz/7dK3g5sfdszU30tOrP2kHHZzhYlsPD82zvcxYixUVVQW0OeA9Mv5nyRguMuRWCTZC8C4
B9MUO6Imho21Heww5xNGLXHhWoEciTWZ23YqWmUhGr5y5vzI8MQ7mTV3otYUAu/6+pcsjbqNhQI3
AfjWrW5aKUSnlB1PwdTeb9DHzNYJhfFireCqM8c6xJ+zoZGkH5NVZjO7xkCGOMJxetHtkGMRwIHJ
PTdv6DBb4Z3V53maTDPa1tx99OAvVKZM38qi7kHZP80GqLVXvuXmEoqln8NwTC47KWmgee32FfX8
SCo4+5Hp/YCIyK65Ww6SmmceMuxPC3rRihbNZ9W2PvzQTE9ldjYZ5A1BKCop7GRj2NIINMzK7Lvi
kx6/duBHzrgbKgGFpThlxsI30C6AGQCidDXw8PW1y7/+w7/SMznyx65sIwgBFD4Fg15W3OcJg009
RHgWs7AHwqAeoOgXx3AFEBc8CZTDg/+MhorCuFrdLnTjQG1uiu2gdNMTdpwibzJGlJYQ7SH3eQ7K
vbty8ntkgttRhJkCQULWwsXWIjWaKsJ2fOUQoRtIBDF4xNL28oQuRDLrCdxUdlB/c29IsUPO89N9
Gvlh96WzLzgGEFI7gnKjYJ0lb4ZBFbNig8miqwakhanBBOzAueMaJVxmqy/oe2N5dQ68zSCEoUq2
Fzb/rnoxGuP1MeJ2jkt1wOrkf0NQc+PZgGxCN2fIt87OOmQ83HFr3Z+Zcn8X4zvTIjsdSGujSLI2
ALFcpvP5m5ADPIdtGD/XDQ2wpPsBLEDA5lr7Iww4xflm8Siz0rEO9t5/wPy0FBBujEINGDWtvg7h
zcBh/xQZWuQOkmVEvevcpusYP8W3/XMkbOO4+8twPVlJOOvY43LNprOpEeLVDN2RUO/NYbP74L0r
iBCYOuEk3BLpVqVot5YzQnLBY245ZproDMuIJ+/I/XuCACkAhOVaju4ANERrwsK/4LggIwwbx/ME
bY7N5R7BkTNfkAfoVsQMmI7rljJozC6NCWrVz016aGq4SVthmj2YlY3ysT464bIXBKlSKTuxBPP+
wUcOdDywIOFfLHj1SoZD/Olvup0ayXjzoMzwZ3H1HxZxbRckVF4W3OLoIjR4c/ktOm314TILuxyY
cMETadxVluCoAeKrX14YnUi1C8jYbYh/q3GePPbFJTYEgTUORmlNnkoJX3Ie3XLX8Cwb7SxvJYjv
9OwnWIsiNC48HrkLTHJpBXCb9qkpOKdfcEhCXzv9AQ/HkUHrUbE942VczsB/7iKAOYZ5UwG8Ggx2
jE/Mb7iTzhSoocfAeW/R1BaLYNbxQ92zZcm/Ztcn6bqPWeFCgGVC7emWucm+2htzwnRcWNSm4+Sy
hnLsA9PyN38rysV0VBgSYcz3Ua7x4xfX78xXFy98rt2vcQXt5Aww/j2XEK9inTK7S1C/LlPW9con
4K2sbk+0pYhWIXBHIscqh5xtVd0dbnM9XP1RPtADmeCmX93YcxIWcpgEYLjcbmYRY1SWBkZjCfMa
w+HCs7E/wm609LQKqzuH2s5PMIz4v/DT5o7nabUhus4aeyj1DsYIVZZOS3SzY9Km7Fdv2CXklLHB
CiwABI+dSg+N2JeSj+Bz+x/4jmRY8KGWsZdPHvWK4jlp64WxEvAIA/dofjnDzfWChar3OSZSBglI
GGkXvAhv8IFHkOJuYkOVQTMRWBM9hXbAQjCtmlVYYIuxsGJ617/x40a+12voeiQP2rLhsXoeRJMI
HKEJCU8ejqnggGgz5ZXz2eCaX4ZmoCwMUGdoOdl2k/LKQZGX1IaGa2FvRpegOOyOZ/dxOy73c0SG
dxOS67GqePiKjesOCUA1nTOPZayFhMFf0r6cCj7uDPo50IJu+xwBIDKQckd3rpXe4/CgCsNORe/f
nH7w+rpAuK3iUPFo9PabXaeB2gV9ESz9mhianKeIaolfNGlAW8wwI7NFY00OX231IDCgZ+v1L1fv
mq6WWZ21ylk5O63eBAVjvikRQSlclzGGm6MMiFOaxNPkmC3UNFxfvFYO+KT/Ja6klfuyYp7RrYlY
5b8E/4Eknbog1g5rs7SUuNugHGRXyTu/PU/m4KN9x8LICtITQV0tXf+D+IrI+fsobOjh4mjssG4/
J2hCxAFJyHs4JrtOj7RscP3fE6c7bPCXgZ+eIRhTv0rRKbGe/vyJ9HGgi/HoWtkO3JLKYtRXkxFU
3OVYkRyEGM3sBqUudhb0k+GB1CB/ETk4b4CzxxVfonZ0GHh7Yn5yshsrwkpEnXu8eOT9T1q/a6TC
sIFgRNPSJgdBnqe3cC3RlM7jKpNLNEgHZt6vFyLJt/cnp0vc2DqJr8LIoTC8RvSLHqVp1T7DO2ZV
6VaQ2uE1mwu/mySgorJhX7QMd+M2C2tjmtwQ/jFLdCeqWTuefPOckPQnE4a3JMqTtc+2pgryb2NF
pqZv6WcysGk1pA0Dbtuo53gNHg7wtu/Cn8KzMCJ6ATNKVj2hr10Vko3ij9uZJ+rLyH0G4MSgEjUe
kAhCcGDUomLAupRc1fLW6lrO8+ARKtKtARSquKwmUjojSn7Fw5V4iHF7C3tqjiAh40EwMjvzFFFx
dtCYscY73b5nbXd2fy0MBC753krW6ZiRX/balG+aTAVUPPLjCenPF0zzJork772UhCqIJXG2eO8H
9D7j1XgzpNr0BtBCaA5OCGLLf+qQDmp8Sa/6h0Vy7+NnY3nY/frioo66yCDBUEe6R8J+O/2JB0pr
TkxLSxs4Bidt8IzerqY8iopCI0cl6e5rA3cEUOuX7/n3ezkI16dJw+VZ8nPKjtUxt3O1BOYtC6d9
NFUjpyFBFrPKgm4YzthV/xqZafBsxFEpSZ4fHHCe6b7PL4Nnj6I765NHNGh0uo8t5YzAgehIZX1H
KRwd0n3tdmYiGZHRXtGHWkY/a7Pq7c9BeyqrHjKLTkHb+Dms+IcADt6Ath4YdGa3v5x8oZgmnV0Q
U3bjmu0xVr/ktYU+W9JRu/Dfplav8Hyg4hacPoBA+tUKGt1nxK7DKZSyOgNrhUKOJH29kwVhYuMo
iCqwIRxbVt3/+JzHZ1AII1Td0ObUqPEAZ1EenYhFWWOjf2BgstRJR08sIh2Lgap8VFM7SNrrOJxI
ds+8EEobbuMqtEbWgDYXxAOOpgNVhdA5A3tI7DKjeV0rhah5J822WOsD267yaVlOmsUCWC5x/dVZ
JqxG5x9DlWeuF9h99PyFDiA7qKwBlqgjxnMsMYhsr+ivMEeWydz6CPz7PVcnlsbOgXG3HMe5Tj+Q
Dz2qeu/XMjdnzmZNgd39Vnic7anKZ5yCsyVsKkBpeVkdChn+OyZf2vptDmv9iPDvaEeeL3+KF5AU
2le2VAU9+5/sV2pW/ZmPkhJwuGRZJ28GS+oNSNhMcR0uy0XcKkBQkR2wjayMIeiIj3UQDXto02jk
62dRx6MgXUJLZtdxZmqNoPgc0ELUxDpfkhyp4D12FXkiL9HHkn5h33Yb08O8q6hqHLmQ3fpvqMU6
UHkvlhG2s9V3WHuBCLjVHqymnjwrkkvgdMmc19yrpSOYOzjJqFgD8YRpWov9eSHoG1lZgjr2Mvo5
epy9M6nYsnOeSDQJxJuoiMpLw22OI8/jeY0xZQ3pTNp3tBgKrj+PGqssmRSPGgpgg8Id453u7DJp
cPjLpvaLKHvaO1RrUnc2pMgyExPplUcBdaXVAxXfimz8x4I5Fdb6mCrbmipbLNX9nb6YojMPeJ0m
pgsq+4CZEo99wAwUJT+4pDaMDot3mqkocFLK1sQk+Do8YhdRsEWlhJSliCtKzH4ydf8OphTFYZ2v
ZmaD2y1Yr7/z8FhAxVBxZre7r16OEBg7bmRWGStpsGQZtF3SSdG5h0qCXgJQMA4bSpkyQ9qqQ7MF
9SIicvd0aX1tYrOXLey4qWRX1zYHikLFwvYEk/UgwuDK/ITX/YFXuVSbLReBMWrzHsTEnx+JHHBF
EuFFolh0euviah6nFLxobsY9lylEPYrzxWzpT66NgK2eQEe6W46LKtR9lMBHfzHmuDE6/9/98DLx
j3NglnmT6Rm2edI63Ge8bMUrZObSqiM5LbjaVXE9TVuxsd0kudNwy13f4jF+ZdwmAzShoTtLMsis
FgPPKShH3vX17iVEmVOpZknzgNUT8Yth8hVS2OUSwHRB2nvwFOVo0uwe4gb4SuKLfs/yxyJNfR1L
EbD7hQTJCQHE74GOFITDmMTuGU8WExpbaK6iBLLuHARe0cStQ523qtDIdQEHdtnILX57i5OYHBZx
hD+17cJTmDZjD0zaoX2cUHjEQtfSSIAAMk8y1vXBvJzLcSUUxRbyMPbfKFESt1yAIrXfWW4L65h5
5hPgaADQNgiJirXxQOYBmd0BjVC4irlktsUciIK3zDybPAGeJQMwHHSqnU06/kvBVXhYlCkNLQJL
aYa0+WyfzYQ8UJH1rvz6kYh483HW2NIT12LmSLhtJ24MdHB7tqKBiLlm1J4Hsi718698KUDF4ZeY
71Ypq+uuZDSVkz6O20noO2tMZ1dSFNkR+PO9KqMFt0wrNDHNOLamEJX0YglmRESbGlVLr/VRtQMc
lSBPqI2DKc6o2k9m4f1zu/ZokRYFsXoNi0qTNPvAeZL/mnhhm7iZ/nGwgTZ19pT7ukt9Q31o96yz
nv873k9N8rW792ukM26DL07xC5g2hYfahDHRJjeE+1pYUqYdna+O2UTapVtPP1bitddLkFap1ddE
9BdnCPvhld9+tGpYTWeEJeEnKszPmcGMa4/HR7/GsZXVEwiVwjj6JVQAEsm1MIbJC/RS0kxQAELj
l+NAFCOe+wse/MeZVNDpb02yCNdmIcxmiW4JuXv2ymn5Eokqe5iSKlM+nCC5Qt3ISO+I+fk/yXtH
WUWprLZDD1HdW+PPJtgnd4CV3GssT2v9OebRxW0uw51ntpZFAYIKruitBI2iqlBHJPznEjM8GMoN
UAvsIr6ZNmStjQeTXFaElpgiD8h93kHwT8FC7Mwit9PgSDsT2mqGgTLof1HVb3jsTxwkSJy5oTZH
VBEzPRxvHT2jdw64W08trlkavSR4jGqq2+z5xGmfjjosBiZ+e2vP9ZN3g/IQwEwS8ewyDySCRtkH
CXZ6LhQBQWxpdqSfcvit7ThAsa8YKhL1FzSavZsDDuecWBO3oT2evxCh3njp13eC/K9Z1SsAZJc3
DZL4bUfTf2n+GtAghFXUEtT59SPbCMkL0NIAX517OwNCpLQ08PFWsN5B2EnnHqZBnFb0uEUJ2moq
sDkCr/UY80E+SscNKWIP2CVCO6ZZutOliGNhOQDpJu8ttubN0c0fOkw6MVECCc0H0Ws0GTRTZKt1
+zIkJwAhaFpEFsHSvl409E6NLNSdBjiQYBbuuTA7a1rV24F/b1peOg2pPqnvSz7A6b0czO7XdfX+
8984hFjj7i1HOaw+P4DMh2kkxFh9hRqrF+rJ1oRflgepqg5w+U5l9XwnaFs1ieK6cCJ4jp8VS0IB
9m2Qp/0IVTzZeN3qXEn+FfhqMuJxC5g3CUbdrEfnwQuiXogGEhdwUtfE41IotBabdejb13VAz1co
TX7AlDS92rzaeGsfX62SM5S93grPSzsUj+qpBZaY1xbII4+uBrWuVJfv6ARuYmh21lu3jba/5/HY
qYwP8w175epOEBGwDz7kjh3Ql2A/PoR7mkNMfqV8ahCP6ZbNusUkY7Ly39oPDrbeXkBmXoURWVV1
gCP9k1RtWAjRilrL7YflE+rNjtY9dIV2QfxtwrzCvj0Feq0FIZ3/5I1da5G/l+Es1OuT//2uu47B
2QB2z2lqrtSyFqWXg6AgXTVH5qPq8T0gdsAQIvMau7tJ/nKFaPCs+LH0/xiskDXQxb5iMEK9p6WH
FR28Eh/8ptZT3YdzUFG6KbCFLLn6QnTD2fPnQxL1KMsgkJ8VmS2uB207q4345/CjNq2Semaw0AlT
BoZMj2qUILLOlcxE5O4OcMN8CvHNjuVhg1ZaHYLiGEyKq2xgXMrly+RbznWx86d/5bLLxCRgUE8N
agm9gXGmH5WiEFibMD5cDHwqbKiYG3nzgrrBUwXHsoHqIjWrtSrhKUQiwsg4sNXSkfLkaknsixc5
8GLcL9PTn6C11Ru/0y1+oGDThznfpKuZJ6cUdWFROZpfK72+AgFeD156exDeXUQW40cTJ8yKl+T7
K/Kn9sl/IUMk1e6kD9lrB2eX25qJU6UghsypIgFjkOieSDkZNk50xuYOBYpvT52LB5ZGdIj0lyTt
QCQ3hoPQAxWVyTv/ARMpv30OsHnsersZbg3SQcKu0WBRL28x4dQS/WKl8Q2myhzri9ZIdtNomdOZ
ELM6l95BCaVsc2zc1bf120NcCZyfLo1R62mg5I+69rVzogFlMrD8Kg0KD0QDrP8atP830d3Z6uB3
BQ2psvGgpM253TirxbMmWD88YpmX14uyYnv+hn/iZp0tF/Aqi0+4JvrMuiKCMek0r3DhDlUo7+7Q
vaJ1/6N5sQmXNS9ccQQIZ175Fzm5mIFaobd5VpMm4Zf3vXURsOrO63ltjtnP/vpR+IUqEXXDFyX2
y9SI1Idze5iS7lhJVOMasSSV5gKpeIDPueKYsfPpypCOMiZ5xYk4y3TemLHe6ORjmdvuiZ9kmEv+
V2kk5aFT2ZjcaqdCD2xTokQ4rMumxH0lk+hEwo/Xe1DThKOvGxoV0xJ/06NHzPaOrpfFsX/Yn3sx
/J6QI5snvo137DBQSJ/mmuN7twmLm+F7mRBluUCEYxx1BJFpfcdaojyGtmVqEuXOv1dFAZDxKfYS
BxqngLO28iUi7yjLne/HF2qZECgTk7PVTONNmTb3vJimjpOayuaTR7iTIsctYPOdSADjUUfBx4dv
fjdMXLutHPN0oUT0xJUJ2ppFptU7TReoXEgMJjOHjTSIJwNRtb28cOVoqR/ovix2XyAAwSdEjZ0b
uQ93khUfhfOuNgK6/b8pv8Y36Hk/C70deLJd9LOmlPGJMUZtHzRntjnNjC7eyemItwOaBm17AEN3
gJIc1RC2yp9Kt1TYjtg0dn2z26385dQ6apoxLYKaI2KXhK7oVmg0aJZH+G+SjwhWKTq5eBSRXPb7
imb/ZjpAEsY+TeuqkyXy5aVFiu42LOTsms21cmwnnwWEHHlUFCSUpon9JhVKnNk8muB+l7A3XWKC
7dXDXDDwtJfcJYTJPSGWpHIm7qKRFzkUTSvobtsEHgkgMM5sUqB4ACOjIvdHUKVqG5ckLZDBmIQp
lzUfZDzG2jBxZl99n1OL14k0ihAtTDbSYcbhOfY1KT0khdSAdYok7O6aG2c94F8bCf4ldobo6T7j
/UnZcFjLLIqq4+zQ0xDfH1TbZjVlaO/unx9ViHdymNakuJ3qK/nRjOOhOJoez0WVimk0XzYiaxn0
Y4om+yZY3nOdCm9i0eMAijN0Ihvv9fAcPHoHbiQA4JD082Itsm8nImqmOlZkkHIIQ71fazEcs2vf
pxvDjGgQHe605IMXr6QwsguCjwnW91YbrjIgzeMIJ0C4uiqzL3TLcheU7jtZIlUWlL5AT9UMTJOu
GqLgDfAAPvUXUMKKtpRmCoxu4oZlL9BTCnIZmRGh2njXrE/oTH9g2vLZgZDL3iPAnT5roynht9x0
C2JtwngWpZAIj6AXFdzKRouYSqBhgVpvxYxAzHYJApcIxlHKkwY7rtF9P8YhEXiAGyobgIbkek52
NKKoss+RAbkd6KkHvr3Y3Lbv4/Zc94cIpM9253DE874mBzSiUxQ38F/sKLRj+WVBYK4qgemstE7R
OHIcRuvDUnkZTM5PIRuIfvklZmOGtcxbBV3g4zPJxYENHk4j0S2+8I6YKo/pzE896WL0bvW5yqCv
RxKpfnERdXM2fclPzYnvY/Lfu1WY15OAv+owDQIu9q/V622jqDZ92wD1yHeKNd2ylKtKVjo1qjrY
2YsONOvDHEAMPvzStdye3U7u34HMunJrcfTTg5yW4IyBdeefY98lN0BEx2dMWTpiyGfH7RnkZVVS
fOvIVVJVbkBg1TpktResIhdnis+mWwcg5xR+d+atxM94HBZ+DhMUh9xNd7AOXyc0LZbDBX3L//PE
f3dIngLj0V9eVTuVuZLePdcdwUSTygjYjwoGROdOhrSQ9srgQCax2x6aa09raUcb5bMgTp2WQX07
46wYqwqhwUG++w6MFzrqL6SW6aO/BAWQMsYyngLNAcBHqv2h+681Qbkv6Or/WWn7YFQCqoUNB5Fr
X1dVxfySr8/HVt36wSd/8TRG3RpfwSAT35YjxNc5JWAiNiJSB3CpjTjsUBNOeZbNtdj3cmzYnqE3
f7J9SPd5JGebw5GJWkyDgCV+tWsk+l3u1ZsG5PLy+Pv34d0vypvLPKjaP16pXyBq68qdgqQD2VkD
VgMjcP+00bcQEpJ7A6KhQoeNvtIRfFajKjh3FtAIQxfvWWGzdE6iF47cHFdVZXLkZLmSpODgRXyj
wTzVPCkjOIG7iZ3y9mQv0PtXnnu9bcMchNM0n3V4x4XpKKV1ZuPU85oBl3RDijYZR6xN5PU0kP4P
lQd037d7iuQsoee9Ef0iWMp3yWobVULa/6Tlu7uz/NHo5Y6/9ItmZ0jzXUn1lzz8wr0IezlCqs0S
1GVUojDBgnU86iR3WUeCGbZJ+PL0QfpELZLcUUiIQsc6c+9XimHOeTqn1I5RcLu12ZaTFTLAfaMy
7PB4/oY037iz6pBeN11MxQr+nk35njS0BEOQKL3xDsAsSeYcwpOExt4L9iSPyHWuJo406QMH9FjW
Q9ZdiI6CmwqQqdjBg5kqegG90NNRey+Vj/kJ9UJbi078iLy5NQU7wr3VSY1c61RhWUXaYY8CobQ1
5EzpFO/090EPJMHUZuwfXYB1lAcze7r1yGINmXjst7V8o3WgEgXr8hHCtoAWjad/5gftQv/Vuj3W
hc+ZFhf4iMVE2IMnZAZB14BTvX5JcPiDl5W8CPqY1Ifg0DIds1LuD04DBL18nCzRF1rnepTb8ojo
bmVH3rXh5sHzpy47/+Nwa/M4gx/j62IP7LtW/46NOAON6MB/Jhifg6dNIzuIRQZm9N2yApv4lRm7
8m08O1iJ/BcVxL69QA1V8jcWK+/KJLSf5I6fQvnIBF+LTVu5H5qGtOsTL7HPrMA6v3PzrQ9fjdg+
vX/XDcjd7nsrsxgWIE6qTo+3tPyX2wGZl9DDW+PToNZ2hth3YMzaLoPs3b23qPt/sru3X8hVZ6Om
OEogCZYU5vVrkkPIk54iGqNfDKUEe/mfrpJFBsReDt8f9mGXV+KoLBgA1InL34i6wMqkI6OYK095
uPaBPHADX5S+zJMN//dNS5SvJj/YQEtdA/JkzMj9LVPlnkYr4j1SanynCPW06hDIacrOBTVyXJtA
bsoHQqvxPAp2Tv3CRG94cWMl4ave8nPORlXn3WltRqADWy5ZC/avRewl1zzMx795jewM/2ZKmGLI
GIAUD6RXUEYAMFl/A2PL5gmwZEjtZqpYREjzBUmLC1c5d9WZ24XFK3hBMWLPG0xy0A67Mx6DAOLw
gcchk4CAVfGISY4JA0nlvC1j+d61zvbuhGXltw/OYZFJq7+tSncoUHrZyO0Z6wQ+dYSeDKkpP1QJ
3Ilx8L2WS2cMdLd76F9Yqq2NU0Ey1KtV+AQpinlTFXCAcbS47swKtOtQqsCOeGR/lUJKvMRyUXD7
8YgITrAGRF2lZf8sKwwtPEWlIKuzZFmxNE3iFqnkXOipq+JjIHpQ2aa811Da/p5PMZtA9IJUZqi6
UAuaDijv8DZF5sYazhoLuXeoGu5pavVF7V7YPicvcBczarSrHbz23zda7WjOqhZn3/y1icyqzOlf
r34ix5gzZ0cAdPf5cTLpZZKkmWaOI8BY8rynnwSLYHZTxeTcs6xQxEybbHrj5mAHuWFf06erKyWd
oBuu/SJn5AMj/wrBJ4A5EcnkEyb5udB8c122D1zGzLtDZHQpFJY2ygTGKgYsuFu7HU4CozT3K6wx
VO0ZIeqwog1e5CWp4Cln/PIoofiAoavzW+iCIGN1vxalBKP6QWDTFxNxo4pHjdhuwXlMPutt/oz3
U/3RtGV2tpNwWVCfkpO9FGSqb1i2TYXdiuGj2h3XCz2mFN13jkrnn1rarxek87HzTXYzjDhI9CQA
zNwbnBUQacVJqsAwAZGtYr3PzQmNDLipfD76SAoDH4wdcKRW9TsO05+xSpvUXdeiJk9UFX1yA/UG
DykxmOqfLTpjwCT1xdIkG4w/g+2a9otlwHAQctZu91ysvz1V5ofe9XF3qKjZWWy39ldfu3WFY8RB
ONY4Ri0TsjjFCJkfOuXyo8xVk+6ErVNpSUEzJ8cj6F4HkE+W2GLHOzftTqRN6tFFNRVVJWOU7SD3
kUuDbWwpbeWh8K9vhGZ+X4XVJNjqjS1vAFLab1r8/T3u1HE0rZmYK0Mmy/FWCFHXaB8hee4kRyXt
8P2/OdnkavULJaLwMDn37hhDOcXg2kpQwSIwM1D4v4ZucVXcU2HoV799SzmhUtz13FW6tUBkffvV
oFf1ay20Vr5letVjWZr+82TnwI/o4B3+TDThy6EnxN8LaLkYHRawQV0kPT4d+qHl91Q/oBi5F+t/
h9nr//UiqQ1JqRegfGlWddeuX/0Zp6xEIA/crKbni/xy1Sdm9cQhA4xSldhwF1QG8EYLTY7rT22Q
hmgiPg2mSrfPUgcdpR7E/slfAT3m1RTnQIRZIUrtfDDG2VixDggu+DJy4mtCMOLRWH448Xi/jFek
WP7liUFUxFMkWT9HffuIxVXiRj03bnqr4c8reS/f9UuRJyXBMUutWh4hcG77GkT/6Lm+XZQ0K/fs
RcmpFfYAQRBnWomX9CdXHh/SB725ak/hhQM/LClGF4TfMF6ST7R/118dFHGd2GN14KYDDKtOAYPr
WVcKY/dLpTfUsAld7XEq0f2X6o42KvfvRQId2rSsT6EBa6h0HL44oBRnsKHrEm0im/OLtvtungSU
jFsacY07AUzt556lVsJR5KYf7x3kP/F8BO3YWfEgVMJf/28e7Ev9J4KoMk5Ly/e2WZh2ryGmG3zj
gRk8LTNvW9MRJ0CHtK2ynPV8lHRituCHT5HRUnROaTcypPQvjko/8ayA1LnyoP7I/OGcLRqPNnxv
PLcZ/hxDWwxGrzRfErnnEF3c+THNGAUfNLNbsQXNvV08WIeIVm3nVDrLbD3QC9cAtiRrje/EAooU
qAfI3Wet9XVLaLyAEnSai6fitZtHzAnN7pkltC9KRmoUWlzQ3xIuNdgGRnnmSPmMB9SV5A/x9tml
g0i5sWIMsOSaCzIhTR3VFZAzEhSfat+vgXM1Q8Iz0e0kkUlgyhCYWGeGMA9H0IWVCFap02wWQmKB
RxY0V5lPfwa6Qwuhg2r/+7i78jm8dz+UlhL/mdgXDDlyHcvGYvmcHrRxmra2mH2LfnOoh4aNziZ1
XJQiOZ0sRzEbatGJiO/FShzp2Y8JODN22BEvwaPnF1B1CmYAfXfbzMIrwp6N8eHgNGlMWtRlbXFg
MlI8ykh44IGYN3JikMS3E+X3250gjS9841CK/vmkWoZvCJtyzM0Kr0ghneJGu6NPl51bobm4ZhVB
w4Cb/hLjnf27eOVvuonowKh8q1wRCNVfll/MaXyeNBFVgYDUYnmo3BkCJvFARSQTcnrbowZLL3JP
9TYAeL9sXbHUr0HMg3dWmC4oydjhmjDQ+KeNcIeHvd5AQs23jWEBhTEX0DIZiodqsGlMB2RcGyfi
USv45KQofq/78nLtr0rwWiHesAknXPf2iu5KlxIju5h82iF2IvNG/GIZ30yPIOcRnx3sw+//gUiD
Sfou/kMG2pBL3ERpOvRxmfIiTohkGpUnaobLswXKwBBoRy9/l10S46Oy+Gl6h+zkqoJoEWiEBdj7
HKk8JJQ0Xzc9lV84ah+Y+lHmyC/iO3M76IjR2NLSSIjEYSiUXVocZEKLxTC+8vFSebm8kVTsHscL
Aa+MifLgVFlkxWPMM6ZLXd+umR7WKz0oazn+u0OO7+/Gcw+dDQ+Ho5CAlFhSS9x5IfFxx16pwnfn
wxoZorCN4wo3cTo11xmhFXzfBQibx2ZwtcQBlfZcmg3kEUz3fOfw4A5xD/yAlZ0yMjiyTjv68Cjv
d8h63tHR5YfMiIxnqfQFBajL7PLiL+FvyrPknkCcgTtZNH7i6rf+KmO8fLBCtswrTYW/b2hTCcUx
Fm19acmbgCdUu9nff5B99gBUdjbEt3uN6utjnVILn9P5cea5QinbTgR8Y0nm/TvpGyV65YQGUjuV
b6u1atluiORyJInzAFkkCs5SX/z2hdpADsLz86+JfeY604BIb+hfGRxWM0nkjyt0kMGv6MeARCkw
JokPRju7O487tqejBY8NcjdT2fiIlQ4zIQ61SJpvDo6nO5gmmyFArlQ9iC5bnICkCNsvnjWmeG5d
Mu35DMqF+uzgEFal9uWt6X3nu01IXwVMZSUpwFXcqV401D5KEx4FtVDKx3CcnV3WS+E7ZbFoXYtH
ylNX6ybIQTnWM39g7o1lRERSDbCcyrz525wAG6QyozT9kOsg032SYIhBk7jAKoMfDA9ygr3V8OZL
SB5XXpZ4ataU7ajVUIy/ebLvnFkdfoHpi9P+BVzJieMHGBEPFyoYxu6izkL0fXtXKOu3Oi5EWQko
jiFJr9a2WpwRP5Cl31pAqMN1TSXk7eogIoZMaz/Bf4o6TzxZ63ZEfg/H39MsxQuNqEXkojzaFUpM
OvWKcS+4JIEg6U10HWEAIvkdRG4QSPHR7xeHSpnyrzX9yoQ5QPx7hj/1NPjtP9L9sH4tl4oeDUPA
F8pcm+6kHjMLEu5Io867XIDxo0GZSsbC8uLh9n6Gu/u9gbj7hUQOswGksEDUw9boFTeMHQ1YawzS
pjIBjmGIq0ca0h3MtCDinM/4hiQIplcQL1JIOdiPtfe6TJIGHyP1Ma3Jgsu+I7pq4DFfTt/QnAJX
DDLGaKV7Asqm2KYqiosefdK2HvNfzXjVs0X/+Vsi/gtM4ILhv+9SqrPrKqJ9nw8kSp2V0ezqN/hg
fuAPFZAmxIbTGM7+wrWSf8sx1wt8XqMo/w+i3ut6sTakPwFgxPVfZIgg+wv25JwI3TLNlvfU4Vtb
EjtYH/BqCl0jsLoO+Tw1doLMy9v+Bv6XsrQmAyMXT1wmkUPSdNLS1p24+DpdAVDwZpIcuqomF9ja
GUJ7DGnNYbIkj5kooo6kQ2mjBRysrtvf4mloxJJKiR0XwslcW5/BMyCbkqXYeUk/NVOUgMcjQXY0
MD9XPSMnnZEd/mI/fJEgyAP1Tyc76Qn8n32sWW2DqddzvK8F2nsyzHtTnNLjyeD4MRgfRXL/IteQ
mhTBN2aD8Xtylt/OCvryG/BXoExu+ORoYH1uxOWaRRM+Ruiy437P737Bn9HiaDGNZI7P0SaRN0gR
sNXNXy3VteavyTMTu+Nd+JXu+ye769zafbPZMr0gVJWNjChKdXCpcK1L29Jn9njEybZ+jDLXqpew
2IKBtDB9EofDXNR/ahHX4b+JMIZvICEzR/ir/+B6zxYB5kGxztonO8fuNfOOsKNtLOA9pPcV/f3i
6TSs96ZpiacIuPyHQ+9EzF4O5MQHmUbakzcQ7ovWGusc5NeMOhrIj1TyVPX0zRCruMSOSJvzR/xu
ekxgEkzmOWzM2wFCg4Xhz0fHtFndZauCCKmMyNMBkBcY3hWsp+Q8EadfAHOOXFg3m14fVIqOSWzX
KEMoL2z1DWRtd6eOoW9o40DqaoK5bwo0jw6ZA4NJScNmgdi8Ajeil2DXshNgG96j5+RE8lCx3bXf
Ae510/6BkgIC3TBqBRGwPGv/pW66bVUIn/Be+gFb/xmM8c2LwugRb68wtqGPNi/tEZgczlGwR5QA
J6iHRwMgDgJUugozfHEaBQBwzlFJYY57sct+u6pGL2PLa9SaTiMhPvQk2kY9ZRqaJF3bqKi7tAh2
qZlmZkP90E3SJDe6AHz2hRqJbUkT/XgmBenpBY9Fagn6asFmE42UiR4NEfMeHAGHtAG01p5M2Mcd
thW4//grUxdPXS9E9QuUBoXXWrK1+rAQfn1vUGdqhyYG+FGtF/bZV1ItohCr2mRR/BCCO3ZpKC/u
sLzz3eNiUkBw1oakO+hHJrvwBWVI0YcjRGge+5LhLrRf6K51UIDI4F7vOXQxozxiGo4H7MXmDf3l
+KIfu0zQSjLos5um+pklNo65E5Qm9NBWwD76HL+jIJTBbZMQtJZrSC3cuCbFBrwlDEK0NQ7wCEzH
FVcp3EVNtcjRlL9fIbZZovkTkFAZum7PEAJYDNc3B3WLoK5fvs0ayzujfJ7AHvde5BlKLsILqsAI
c12TvBboN3rPtz8NfQ/4h+Xe3VldJPLme5jT1fMnMxiuzQoOeuzxlv3tHYaYOd2QKD1nI33G+oAU
RdEac+dUvbRCrqtSyZGqmyd0hr7rqN1c0pjEZLPRCfJqYWD9zvtCUQgtJvz9UpuO3W7DfiQhDnEm
Dit5TFlm+r0yo58DpJIz9aHWcJfcQqroIpH8K5Oap02i80VlsKGa3cxSahXxcyvLY2ipVhCuVHNv
I6F3+7lpxJAXncGyRAFonv6vo4kj3SzurgNKSYc5f4J0xBKgg11IOEqkINZnjSs7mx6KGa5R3jZg
NPEQwZfYy4kFHZKlshz607qKadV089LfKMmfo4AKycqfyHp5BrJGs7eDDC9jKEqD7a09P+0iiBVL
mWwxw+U8raCc+JGEKTQsRmNVQE10xJLFMnywlvpLCvaq9nbeNTUZYvTgoq0noc9NSv4fQ46HTCf0
tWHifsBRtodgOzSslgX4fix62QYo26us+tE38eUwuArIQ6xn+cn4Nig/3SfYpSYHm06sGoUoG4Jz
NdDtaqHlHZuhG/G1mBJYLQS3/LVBVVWcx0/KajUCIWpRmsMTqBbnry5WDtEnLagFX+q86UvOtnOU
Hcek+yeaH7pDiiv+b1+XCwOc+J/KsWDN//jLEu0kTSgEcrJrIDmkMiPWv58Y4g4du6Sfk3/pNmAD
++06SRXP6N3Su80FlR1iJ7F0QkI2Tc2rPxPv9efdswwb1xvYOkMZPN1tF6kSWRE2J8K69HANEwWy
gwFBAuDo1Yw/fwQEaqjQ8UuDh1As7txf84zQifNCcfkHyvf6H0NZYSZcQxrQ2A3kLoJ50CqtaQ+F
ZVgNDdzrwjHp4+ZmFRJsLaoTxueYKHrkOObHZY3zGxYJa3VmusOAGhAkBeieSJ12sdIhxiCaD2ZN
F+g3SksAzPNc2jFa2FigUeehLxygu2rSpL/8tP5DkF9VQo8dDwzX7sfqYYykPdwhb7AqhtdakceU
I0ZGnrvbmekKxxroIDXVinLvq7I9WSNJI+BEyv1ffYMclqVUBlQypo/Sfiw7ZKTSMrDFKawFvm/n
RBIapobgks5lqw/dsd4e0qvnjval2tOSdpT20YM8X4B/2wSYxh7B1J4C/dKwMxVUkzpwowL2ZZKa
KyfA4G6dpgy/4NJ6mX2P2Zl3jrVKHBZC+oVuLQcVPihu2+t5uEk+SWN6EefbdXKNSWUT//O+Brm2
OpEMA4VNZt7JjJjvn8ZIUZw/gvVTLwEz2eGAg8lzOxSGwOO5QZuklWIQ3Q1A9NhueMwMHLAIHQUQ
gYOElShV+vo/Hh5e6QqB+dCqfMsXQt6jtU/YHkMIgdwUX0F40uXkGtZ4A7JGfsAQqtQAWEjWnqqc
IB0DxiqWvd4sR6rzk4/Y7kgeXTP258F6IsZnFHL4aCvA+X8l7e1me0hxkWjnHuWLUeIGX+yuAv7i
6OtHqjJmNT8b1/p+ihr6roOH+BECi0tfc7tLYvzmICMqLQWEsGNNh7HRNQUjUkJMDeph46fv6wqH
gWNqrXWEohuZN3XoMe2FZW7M1+METcmepEUu7NUNbaeFST3cHXX/e/mcAv6Ej06ANeOrLUwLTUxQ
oe3fbuRKNHLJTBZFzE/fufn3vnZ6awrYbil7ODNWmqx79LavLq6cn+cJE5QlGgr8Uf3Gsilgs8lQ
GGZX3l60AX9PgoPHOTZb1r4CYkiFErBb0fhxO8adFMqxoq8GZYb8FfE4VuiMQ0+FJ4VxQl+pSreZ
0hYHyoq7AafMtiRBCAYUdIPN9CxTf3oomFSepQdz0/Ys3qfuQjLkUMI2lYQiMfREgF154Ek2amhQ
RbWvaqHoUw2vr4Fm9mO58xzErHnsL/4kk2QCIa8rHttCmvVv3Df1Vh+J8KvUj0QfA2oVqp3uTXWJ
pQ0iHzZcCIrc0dlYTWPgkNBu4k7cx7FTr7Y0rIo922fUKRHhMQbwkIK0KGKPPFEV9IRZ2H2tIQIm
bZD7YHpcaVB5VWtY0AKaRTMwkWZle0J/2hBM7mYZ93PYJvYC1fdnW4vPoADqyToiYeRXUANHTvl8
FcmE3WifZ8ZhEFbOQVF706efg1RAdFaanaP7/5jwAjsd4JT40M1bzly6dBHHGF/o7LXJ/F6BfDGL
x/i96Eby9iGvh4CHaBVYA+ntAlN6d9kb4LblNNd1gFKgpWLs/SmL8hHwezlIsDLC9CtOPwq+B1hd
zNG8lc74EWbKLpS2HtEpj7SmawstGZYDCy7NX0Joyf91p6D2EeTacPOXN7+TVhoCCnwl1Z11S/rA
1ZsisdWclY0VteF/OtUIziasxe+5JDzCaIC75r7wjDht8PuEBy5sFnAktmyrwT8XU/OtqHIoFxUA
8bVF41A+dBh9XZfA+onZcZLydc/12f8ohx2cJaWPDt3MAWNnc8NP0IZ3pjmlHx8NHdrJQPx6yY6q
c4QXgJHnz/6fwogfnaZoV7PsFxQjnoIL8B7LdWeym348bC9ogkQCg87/lOngCz5pJPNEl+nnYtn4
Jo9XqjBq9sM45oo2KmjVrK6ZWewtY2rAVRQSS6N48r91fFE/QmYrbBbCtGW/U/8VmQJYTMz8hix5
yrPZXbl93lG/2jkrmhCcvdviDSy++uYzFimoqFgZvI1evSOpqvQc88FQM7cz+kNvv55ThAD5IV6u
Xlccjco2F9FQsmmzPDeYV8RP51WTDPRWA5tH4qF4rtvFRCv44vLDcYVCgu2Eh5JSa4Lqehi34s7M
K83xDBVCYl8PUgCPyyhvVN2ofClWuup78CT8R74gsHWpUqb7WUgqM99utiT4CWldSG6he8GvE2KI
yWFWpqeC1F+9UnAVX433nz2TTzbDzlrqIc0R5ertZh2dmGRHbQ2GtYOd6Cj0CDQO3/negcF4acYm
8Yf8zEHheEqoUlmdnKvl8YnkfAQuIPqLfHvw8v/AMkQ7rq+GxHQZBz+8//VmPBo4GhiMnReqQelt
uy/2ZfJ11xQiFLGrbEe2cy09+XsnfHAC/YgopzddpZnHdv2SWW1C0WB9cU9NsjyaxdMmUBJjrlxM
AOu66Nz1mAdTFq2oq7wseoQS6+oURnna6QzT6PJ8wnn0S/98VOTCeHgyC7DlwIg2jzXPorzdpKAr
6voXthMReR9orxDx9HCKnq02YnRRuo8mdikkJCIakO7BACZjMRRKmvMi2dD2KhKSrJZc1GriDfQG
L74pJTFgBcs5+eVXkTwJi7dTsRjw3RETv7Uat1CYvtGLZJ04d4jGrf/8FqsSU3pL0TOXt9pmlpAT
qxjdsrXoYSEQCr7V2MGEnTcHyqYLd60auQ837vx+X1/9wMAFx1Rib3jiGcqRxd0GZZasGM+/7eaq
oAGZevpYoLDGIXMnY7K75DRcBt3/NJVijXu5uU22koQ8htrYdhwj2ElBESWaV2qPLo4c2ptmFn2d
aikl/183FAy+gMfPZdo6/jNZkCNa0F1wqK9eX/ayEnAnl8z4AKlTQG/U8fV3GrZaGNm5SW5HItUF
7DuGP9kOofiKW3yCxlULFIab4yzuBoIIfxgLKmTte2Vr4/ms0tTsahKAFySpjw0NJFLpiOCNSnIl
XQGqiGzlI5di9qVZvwLcGXH/Fn1PC1wfmmH/IazL+qyZLWH2Zz5qdAuwqn/fhdTCi5TK9hY8uJpc
LwtGxgJwA8qBkFwYAyXox3zxQIXX2zVaL75dkKHLC58MtgZAZSSVoXEQA2wx0acuIn6Bheg1qFUy
sH4fceZAGrO9zT8WIqOB8iB3lT0Flzb0FitSZrK5lMuEYkPnZI8lIRXdykNCnoEjd+i7Ie5Vyna8
s9VmfBd5xqdX6IcJ+B0oRw338egBaDoBYdoIx7aDH/X4+AhZwEWsr0vKngJKrhqje54mukxzgrFR
DLiSPkDGI2qko2KJ326rNAH6ZhmIRxq+INmzvRDtDxG+QuWDQyZYFHgbMtGK8LIw5UVTkQ5ZITzG
WpaRoY1w3w5rD+Ne8kOUFhoGZmyf4GX1xUAviyivk5ma6bUfSRKAVegjRUX5ADmpaX3+z364BbMg
IPvWrScH7fFzvzwUwBwC8FSpMzyzKcHjYrOrjvy2PdJoNDUpSpetBMGvjtTnX4yC3H+Vi20cJtol
Y2Oq7zg6fpw6J7JzHV6OakqtePxF6xFrDWlPojygJv10zXMDQjLeU9X/UGYQhbF13ocJlKLM7YcO
fBXnQoaZT/vy3Ndw1wUGlIRz7NNt0Kqonaj/d5R49RxEVzHdFwO4HZM1FvzSsQKTkLOEpfgCBl8C
VmpncenxZQrgGTvCWnFTqoAPYHe1V1owAYAh0X+vfUmzvwVBBLZrJmcm7g1pGuOIC9UrFVaWzGf3
yvcnc7bp/mzi06nz0EEp7datJcJqp/wp6pWcw8RW17OWk7qT/oEPvSb6w+Dv24EHR28395UH5Bmw
IDugJlDeit/rcxJdp+PRadwu4wsh9HG2LueXmfuCq/gh5xoaS36VxEc/1PAA8SbkZzqH5WSDTSsR
zVKRwQcmBQYYTxizOztC48P6/f3TFkgleZxd/0Ir+pajEgcY11XHcdHFxLrjvQBAv336QoEZiB8S
sUyS+WXNoXaJ/72IC+0dRV8bWZgri31SPnA+hIT4m3xf/Q1/ZPUrHsu4UjeiySU1Gh5XcA+3lHNK
HTb4ZhY++xszEB+qYaJDHfgEsMmKbJ1+p4fb5wZNQNrE90bDASSCnTvPAdMJoCsTKdybhGyQ34DT
TZiOeEB1VNQPlVS8lCAAoOMU+5gJbKifj3xuWD2NlTf5cS0COHZBLYRmZSCK0pAyCTQFzw4Gmz6A
zHVCkmVWfW4dP1mzROLwA4XWCHsAJobYXpSRVo1hL/o/0ZhVjrpZ6P8YvUE85iBxSi/hjweDzoSN
FKAQD8W1FoDmUMve95tLvVK9dMKVjCsNKVy0l4fdn9ABO1JYTEpBr9hLMywXooDVIQBCsqOKUalR
qzahFLpgeyi2vnPwtKwndAAFDqYcdJljuBHZG+8y85uPP4WgA5jQo2F1lzC0p7qyPTekj0IODALO
JdfxqcM0A76YK6RiZCFShUN4425/yIO2h2N5w3qm1TY1GYzLgdrqbIOnE7qLImByJe+Ooc/i1/qr
q3/Ft3EuXoktdqCbTy/IJ33cxyXocy2h8WNLvBcV6acnDIJ68PfMMMMuvWzSn/jnL6rQzWPVqM0p
oeCaP5m83ODBRkusjJQGlObInuV6Ge1urBTEEp9jk4kpoJev4H9NmT9y3NZbAjah3rb8u+W/IKBt
Vm30syXxDyW2kvrDJ+zw/2l1dYPY032XdgPsaRngVojptCqwWu41o8jd/4NxJVL1lgiKXQ0XhVVy
EJYIJovgu7lSm7sMJXRjepVhZ35hQavBEGIw9VsY58BMGrpEgWOzcl1MBg5t9f2gD6Lq4UxaDWtG
W6eH7C7zNhr3hfGtA95/DmJoMcnNFEKEzVjNj/ZzLSZNRaqswmIv/lGDZnfZS57P2FUtPQWvBfjs
2+25ffVSLriiaW8t0+O3YvHhyZDmth6/Bqzaw2f+Z46rU3LEMxMi9Jf8F/P7V7vzEAhsgCt/KjO7
Gwjrm0MSZYDGax5f2w2aN1JJFF/WoxbgtKyBelcioH911FnisXt9wSHvuHAzdtVQUIgzCGGyjskb
EkCZPaEcs36C4wF/FcNiLOn/CajsbbH0QvENWAHcHIjkAE6mP9BQm2f7p9SRpFSB1lJP/vrZBzp8
VTj1QfMdoOB+Qb3jl0UPVLE2rRI/Qg+NJA1ilFRwoTU1BdgxMRvqV0/HQRLlWslkvl7n/KhLuF4K
OGK0xV3/FbvTlahHGTqRpoNAj4h9Z4RD97dt2XglyAU34uAkvDI4oDy6moLTYyAclBxK/PPaI0rw
/yIOnX8FU+Ai0EsFcKp2g+SQfAF90f7CNrQJbfSAtln7omZ5b79AGsxBYQuGPssASl5VZvkhrHzc
yAxwAQE+y6XtbyhsKa++4bRBcFWPffi7ELamKXRPxGMeqMCz6g/FhSXuD+x4YeidgfFtXoDPm/fY
ok21yZlUDJVsq367nsKjjurjmdk2VBDUBBkr9ral1FKVaVca5dG5Ayy1JHaWKk4UUqo/SJBTiDZf
dR1Aroe+DQ5BfHSyIoUByHklrEUDFrQX2PxYofgZ7E3VmT1MY5GhBAEq+JPDvG3Lym/QTmlEtF6X
rl2RlzYkiNE1PieEA5HZCgjInezi8+MV2I6JOe45xEJjiUvNyMSitAS4P2je6MIdxGp/mfJveCJf
moF4wjpzlR9UmjvxrTBSX3HFOHhkVi5hxxesHZhxU9H5eM2kYh1mra+EiqckayRaWFD+BUi3QmwL
QRRP37vSjipbXB8658B/b/MDsaeV+bF9eJVdzgN+yzWrIDVHcHBwwA1zQWpc6LQoCJuTb+1MyqWT
5n2rsB3qT6Okx2W4YmSeD0HjLrb5XUQaMWiausWVNc1UaqJjflnt3+UntLmyWXvsk/DRnyJhc5Mb
DzMOHrIRlnumVs/pz4XKXiaYmnMg6RahXps/yeVRtDgHNXxfkww8Ya3GHp7ea/pWGRW+vYKsHLcY
L0NqxadbsnkFYSr3hXEpXFJlxDAnP4nnKTn6sW8qSHPuSXvXnVI4cpsEs75ugMtaTyDMkJZECBSW
CVyvusNMBaf8xMqkCjpaWyL/eFi78+vynmOgwd/VUtugx5OtBPBTkxlTzlBOpahV8vG6BniU7jII
sBIVu3to+4IHIlLiRd7BBYcTqTTIQ5auIaZzuTd4JxoYosjppKIYXSRaxrmbv6j86eK9aqKebE7n
KhF2/GKZ6OjYz9VaN/D22MLfgc2ZTtkwenDU8NYPNqPJF/o0FcE2ub/ZTCFonxu85qVQqnwf1QnJ
a/Jq19jB/f85kJTsRneO8nqBYU1cJQyvTztC6rcnL3RwQXYrkPySg4IYsitglCDk2FPNG9f0byqw
nohF4YnYJIZiBwIRjjASnsN0XwELzWYCyDQtlGk5HBLJp3lmZoembibqwhsHVRXqBnp8a8JlUVyI
jVeKA7CDbABxlQ/9KUORgb//logPjCBfE9RLV3btzHspkqeNmOj5OqdwaVOi8XluWnDnc3m2Ba8d
V0tG059nP3ueNcvbmblrTvCspDUhtMlVpmC59/iOBx+QhHF/gIz/V9rLvygCyc/ciFXIKOx3Jyig
sF+4G9lQOF72bJo+ahiIW8VcAKYb7g+D7sNeXLKvQpWFPs7VJeLaem9+E92W+YZmURHg5VGwx/ot
P87M9ZHCh15f0CsibALLQwBio/fm60RgjeAPQ+jIiCocIE+pJp1bFSqiZlzw/FzlntoCtq9Loz6a
9ua5flRTAAAsIdDS69pBCB07fDS55G7izfjSP8XQlJY/Z5WpE+CZXCgZEjZDMP9NRoCUzd5VRDOc
09y3Z59VZsuuM2RH/lB5NQTgO9o5PIoF3Y4NbzdG7GRU2YDKi9YCUpP6v2wMAfp52XcvSj0I+YKW
HaGGhrdxI/2ZvwE4TBDxOGl+0INpi7egsW4k6AYMZUVLVIUzjSGFSdVJ+5CnZABx6U3913YsXD+h
vm0C/wAdOyHsPwtKHJ/hvFjOjxSkXKohrsyGIzIU8p1EarK2fj/NvMkLzL+bnZI6eegPyh/H21Tj
skXfnQcGDjE5ri8ipNQjA56QZiLgOq3E5vQMW84b8ANGEubmWUM2/odVe1/X+XKkCZjLYZePti/j
wECrGLEIb2rJiRRug1kfwkgbiFmNxag1rrY7xAGX/AmWXcrUB1dWZQMEt02ojKr7INDgQJeo3fbY
nR0lG+2+qFHD/hFykUUXB9yTI2XOO6n0T4Jy+IAS/v1jUsv/ougx4WIUyrXYwROfRtKtzXTBPPp7
UOzSde8v5fWUw02ffDxCelKeayomUqfONz7HEtcU8Q7Geu1hUOR8UfEmePKpwfqdZEuC8QT9txwg
Zu6PWW7gq9S2YcukEd26k/d/MtXGZMcT5hqcElQqEBkghTL2XsU57lcwFiOhaaGCtODC4tidoDm9
viphspG3vP610dyjyQryh9cXpJwk9QYqYD3Wzj5bYRotznJlDxVW/szKAI4mr4fK8G1BSzk5i7zP
x8+k2ZgqZ3s99/OZABNR/LMN9laFXeLbVSP3rjyX7QfzfIOfRH0dNRIs0Yfqud1d/gP3YL0w2P2l
IJDpzoY8tI/LFJ/hok9KjHWGem8BqFNCYQAQEB0WXk6RIiyqGRf65gVqA8F/G6dwVDCTAunPlZ1E
CNSnRePlsIR8wnXm3teTtix4iet171mCYYx2hL3absrL+DtqmqthKC/snwtPYZ/Rl580/2zgkvqX
f5/9xtLsLI4T8IFCRX7wyK08HBYwcoZkpk8WQmDeRQ86tVTuTWh+bo7/l5/Xb/FLQgyUhOBZkwcV
k+Wr/nnaPJMogyJcetgv6Nbti9bQvAUWi981lU7Laz92j+aDJ9xGX5h97XFByFfmhmFlAMN7x+kX
54WsRbvrmoBJij0o+l5e6qi9KV+9hkVJkn0zHZM9PUuZONwNumLatGU0ep2Z4tcbI15Qa8rheV/6
CzSZMT064yX3ZIB4TPL+/qtoElPN9qM+RJUIajnNA9rNlI2YdtkaAo57xMN44nC5TRnW1Qh5yrN0
sU38s/DPhX1jUCL3WDjBg/WSqU+4YrUNifKpLErrtF5jUfMKqJDDumsctc+FbhPzifP2UusN0eDL
3T7IzG5zZR/XiHxIoI1+e6eGXwwDZV18B7269Xt8EmTAHrQ3GA0yxXcMSN413Tr6ZBTxdV2BCdUO
W8TWwOk3FhYp8pEXSHxaCCmnAVd6dcFtEkVUW+5+tbCOYEF/d32JYK348y2CNUfmmCBpRXHYyw+K
G+SpqSDXGX+5AJ1ypp1Nykt3nS7t0/kW7XiDBmCKuBNuf+YEP1vPRcURuZj7XWO4SGi6hNBAzp1r
SpylLS46MSLbzznBneQesADleMGmSxGwDKqiA/4KotniMNH4j7mRrueETcUZh5jF3l21fIz71odP
MTMCQI0Fz5qu3JU2O9cNIwJAoR8vVAR5s3xc+QilIkQdUATZZm9oJcyCSC9DteFiZ11H5XX3kK0W
PvUW5BC9teGzytfUJM4okEOdCbSEJAkh9kL3b+K8/csRwWEwxaztZZ70jogE2OuikLJrD1Wr1eEn
F6l+wIlRcAoOFEUJFXK95JZVIw8tmYsmTh244F6XlNG2osuEFuSYrYqbrkTMFoa8qQVB+yjzUpUC
lDEUOUZ9p20LSsF5Hmsr4kaMmxUPhRIKmI1FfT83JbUY+lgAlAsnqR3pCnD80vsGn+JmFimyad3y
VIYyncxbGOKtEj5ybzvCfyq+mJ1iP9tDfxObW0Ef55dAHt8zInFI7MO+HUE2FNr055s9P7lYTRrF
0BI7G11ldgdBFP8KnUXkXOcHwlanl+I98MOQ9zHiPb/cCnOoBIXuiP9EceIGwZRaCrBo46pJfgqT
wg3z/T+Plq3dW2UNZnYEX97WW93vGwA06/Ca3A6r70qqi8AJCBALZ+M8BJc4fZr4s0g5/w9R5cPx
LLl+lOTR/lr8ddzgUd5kphw6Bxs18tEEq8Fu9PCiW8u6qoAz13wPaP7u9WxA9M/ZGSxZyHXa241g
uWm3vLPVNslm+N2pNZn6/3drigcEfSTnCmVax9HoRh3djeyH4jV0xVXKrSEtA7znoSPvrB7DVAdK
ClOonGlRwOUiLOzDeTiluBElze5KD//ULeeDRqWnd2ELLzPh5kmbkZhG9j/WGD65JjGZW1pN8jBe
AogrAIx8kKEbk+dqI7k6cbisNNtdI0uK5OSSPGYt3oTuFAu7XuGhBUOND74qCVLYAyf8jvCNS0C+
9jJNwVcH+8Cjr9RvGPxBI70TYacSVj2r/9pwOdk5GQH6pJw2Ja7UlgeK2/gJ82SQ1wyOQE0bmhOV
8sJ8zL4BqBs32qZqvd5y+1PLB971Pe34UmV9tmLeRvtaQb+/icZRboISkXFrod4QCsMxjphFOhmY
Nyc4fueRYZ+uhZlZmeA2jRi+HQHOSCbY9/YsMUO3r7ylVp9W++M+6tcFfNL32i+f+rEky+8sGnaa
0bsCfXxfWRl/JN1DUH3XuyIAFeXNM+yaAW+oAYeM7fGMqnyKKFCfxmOqKscHKthf9zReA9UTUiQI
S3C2hrOcWJnc0WMogHqWXi5qzPggPrVqIAVoSKdO/dTDm3lhHxDte2SU/6ORo9VrEBAETIot5WJY
QV35avAe/cp9YiLbh+9qcj5Yy9YWKNCBIZtJNy4YXfKBaGXAxaMZtZQQTYLcFBdC0+fa31DaXEGN
YJAW3S7FJLduLGvm2/F0RhZbGgsHk//WBR5ZIZeLZVsc7iogGffa0n8z19wfdUTtccC++YJQMlIQ
UKqd4KelTMupdMtAn7laXatBxyT1IL6Ysupr4w/4VI0cDEuUOPIy4sxlblrfhd2nmp1H0Q/rPzOg
6XeMQcyZGigFnsDljcT5hYfIZqDpNdx8tm1OGf7uHKF+NtmHRFN2uqX9No9ex79yEKFx3fATOwH+
Qel8IxGWE4dgxIKhtOK/j6GwzgPrA88ul+tkJZnx5nKTZjS4uRXH9p9ZqSiDIRh5POY1rYGNhdRX
sMQE+Oh49MktItMhn6kzjzVQ/n8wS4g8IOjYFv5cKWvLp2zLrKxBGLSYMupBMiujGoXkCw6guALj
yYwg3MJQ+gYglFx5L+DvEaYuUIS3uAVkuTC/04egUEgC0sswQvdAMt6HmLrOaQDB8ADOdpCz6S0M
wmgoglO/jdk/vTy6iEm3TEaoNPC0GcckZP5oRxpW9NtanYbUALrvNnEkMoG6Kc10mq7u7izXYEgY
bBVb3GQii0bc4m2A8aoSQ3tXDienYVEXVXvtiv1gcQ1n6u2lRfCxVn9SrZ/qscxzEW1bBxHvPz/6
sVaXl5bIxShtZtuTXCP1iKg9QoTBlVH6HD7kA/6PG3h8QxFgdR3zeQl3WAV7e28rDwKwkMQ/ANkD
vCMEs6QHboDGJnQbjK5TRmKET7/CmHeztMknbZGcBQCnoOCyU7y6XYrIb1OBl83FpjsA10M/ttCm
N/NBgQ5nb3DWrGTls9izRtNHzrbcSKAXymYH8lfLi2iKTWl9Cr+fuNIXgYyWvBbSuSzHUmDSm+Kc
lhikq3fz63vF0c3HTTJRvQ8EC2BqOHkw/Ce4nYiM3wDOKJ3F8InvZQwb+BSbiLpWhyHaQ10mFSBY
agPYrOn9qFSmDv7aWEKHdHNK4N2mmjcdunPppRuR6HhdaU7WEPobsqGvHtvN0xoaDLtGnGmmxL8i
n+gRtbBQwG3C1dRd4N4GINVfueBZzMm463m42eHT69/aRWd1kIj7s8rWXuXaxWlV4IDCDl98ckWx
N9OsWy+2iUvGVxDkWaWurv7kRN73ETlKZ7tsjCo1naoSQmxjfPSJBe59BjNT0/FF/QyhJ+9ELFM+
nvZ83cmhN9OqcGSPWznZh0+RErFl43kTQ9cK58LlZRmhMJGD9eGdYPfZBYYEEcLMXmJHoOIfsgj9
E8+mD8gGF/6X3O1h5hjgvE7cLDeYRdtNBTDU1jVgmE0RGkeWqzNtxZhbTAszmabvQoIIjZK/D1Ca
khF3CdoDMTEOWgA40shfBlHBsX6xzZHheMNHQ42tB1SLWYMBET2HfqrVgdNN2waKH3yCNqjg9aX5
OlwPRM2pw7ScYWC6kegYfkqEm9KgxDbB8KZlw+rSlpLK9a1aEEWvKxL3Y5FN0oaW0Zir168uuBaT
jNFsDjQPYshTBy8KltSEGqKTgvf/X/zmMC0dmXwTaY7TiDylJDRnASTR1eNSLFoukpf/j8HASByi
h+UZ4/r5cpkDOf4sKOlStJHWoKaNa6ehO0ns6TSjQFS2o+VDZL0gqxBwUdiA/XtRHatVUcKK+yQY
8mjx/uDVM329tdZwprdPyrNEn0VLgO8rdTxpu9dGBcDfXC8mZrfD8CpNLR955uuXAlru3Iluoy/m
yCC7vmJZYUni0Gqx9awR8gn+pB6+UwmdnAcZP638Qrs2c+NovSrH2EzAt3ZG6v1WnnJNJ2LRkwgx
Yb1aY9b+gGOKEsDObaJiC0N9+94o/aMCmudMEucSfLMu3E3+alL1NnP4WfidbOvZK9HDhmmj5Fcc
feDhUWF8v0UlF/tFNvlbYFYcql+zegYw+lVVNR5P58Vil/Bph1KFbXsX8RKQUhLtBl3SWUHcnpeL
CTwezvkdY+zo0KKtYMT1118tC2vlvVe5s71b6zkJeHUfiOjWIBtzbI9t7MFKGH23ZaOgxWZDP46O
cLiCSEk/nqa0F+SOH8nZUM05M2vUpRCDvlkAYEZvdmJ2Ybj/nfDZiShzXMcNIRjns9Od58RoA4Zr
p0NW8MWBJYfS+dGGM3hExjLp3ZpE8emFdhauzFg2mg8lEdDS5jnNT2EiqC7r9GnDz0KM2ukuSC5N
oDP5d2oStGYLniRVOK30cTllUJsre1WiQLJ4Cz5+BgSM5xLTz58N+l+1mTn2zfi0IJXc6xX1PAuJ
625A5/iPZ3PGCQkbZFKYEM+6y9MeLl0t+aNPirQ9r1iLx1f+nSEEC1GBD+9EnWuLt+R1To/KXy/u
hu/M+2OHskcNXXLALJPgClG7KQkap+jtMYHTZt31u4CyC0qSwG2OKKUNGFvwj+/IRLgFqJpf+o0V
rXP1098upZF6LkrbeRkyvaJlVJIBhZMsokfY65QltsRgVuSh2fBtABwK+b1kTytuwQ8iIZSW6tpo
L6rBobN0XPeXbkUnzp0r/IBf9FfJ2DeYucDlAUROscXi3GFOvw04ADAeLCa17thOBaNANr3uJcdh
NSV/QFBPjyLOFzLpbrONQ0Wgw0ezLgbtPFwZ81WhU14hO3nBJ8/C7/+6dED5XHl7h8nzwAlkAy6i
B9WIYVQ0OznChthxKUCfnZrus7xj2vRPW8eqQSLe+2a5Rg6qSRDgEUiafceZCuYbxWJZyKUIhWXI
tAhlDAqmbY8VdWDCjnXUJ4WydRlqeuRXYKd1b0B31gnEER60yfERIw3NJFxcRBHQLGd2YQmN3BmG
YrMgr25Qk5wnKgj4iFNKUI1R3qMrD7BB7HH4WZ59k/aEk+IR6wHrVaIrhqSVtEAr+o/IoGs04uHx
yRYJpQlEP2ehON/cDv8MtumWt+hW5gac0gC8hIItJZeuaJQtmTWghhuFlEKVHwP7qtyQy2Ck735/
VHuwiTetX1zmZs7HAn71MjRorKT4ZDWpnU+8UCrUlgg68x1SblqoXBuQO3mx9U0EJ4h1ncryPJPE
UWPy30bhRjHC1DbqWwyspa2SAMHTq3YmrUXhUZu5tr9rDy1iXN4Baw/rphuzJMvtHZj4G5EMVDPG
9IIBVhEGnDN7A7YRQ7uHHpAl91RUByWOpg72mJ1SV+RFmjQKKBt93J8ecfRpRW8cNvkOJdaB0k/7
BSi5ggfUOAy4Bo9P3u+WUcy1qUO7g3CN+ZKEzCHNY7+Gd9UZurnYWHkd8XfgPctFWSsO+1xqWkhh
Q55Qtc2UCjN2M1lBmSGxLkMgMr2+wQ+NwUIZUQSqX9vZbjydzBw9/644j423abBb8sDxUUDR4IMk
w9iCiTr1K6V2tOHJFYFsCK2NSr6JlkwKok/8TDjaOSARfEgkW82D8RKpaJWVmRFSWvn1zbrQg6w7
n94C4Lu5kuHbqKaANJMi705j4IOGsdWRMK9x+jvskPcCj8aacGctaxGOhoHEJwbU4MyxRgbVp6M5
XE54bm2Ls9MdAHL8cS91YYe19kSXzdB0egJraq/N5I7fZ0NIYTmuHJFSoZ+ADMHw1lOzgPKVQgzz
fbQ5wWYCnlLzjEbp8sFTWN82TpvltUl5V4TmJ53XBfEXWOQ87u/FyTZW4ieAPVLa18Gkq7gN8lZl
tJOJqVohkk7MaWD7EEXp62e1BAOpDtq80vXRNqm30xsYAfJzBhYlZBtHLYZBETP12NE5nA5yw3br
eDa+8Zo1xbXgjNNJdlg/6e2OJxf1DL3OHwGjOHrYZ6kVmKg42RCjdolgbcqaUErcgWEQBLjw2zHZ
tBKoayJxF/5htW09681AyKrkEHkqFJYwmnYMmSKa+qCD+Dgxy76nFveE+jf0oq6tCsM+urS6IldQ
77EMFYpprD9kur84SV+D8ZtguZE8q+DRjntxOGM1+Dzp4wt5iM9FFViJIVY2CKlwYBYpfd4CGWdg
jw8bmTia1m+7mOp1QrbpScZUywZaH5zCtmkAfZXaBoKkxL7FT+DRjQnrqVgBH2DHvSZTLnXC2/NQ
0DEL/6+6CmPDg/Pnik5w+HDuGtWC4aB2cRM+jCSfvX3djL/OfPdCB7ozbZE2CX39EENcTVH1GugT
rCd04NbJafS/ClLBdYj10zirfqZRqDJ+oRU2bwRRid7XIK5hivSlbfwpuOpE
`protect end_protected
