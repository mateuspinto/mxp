`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
7VKK2iBqskVwndpDY4Osb1btON9rQxED88LCXLQRPMepgalUiFWiKL4PQFYqYDEoEMiaagKApKE9
T8JwiPsXOCCSbVL1SFowDmhrAvkkO7Ypw6FPo982FrkhUXkaZrtS7A8B0iEu3K51yFmutcAAtC8x
4OK731BcjOQ1lVHM4M7y2DlIwXiEJ5UA6F5eTxXC8d2biRcF8+h1dpYUtanEOvflGbwze2bOdafF
v88uTwf1U6JBBH2bCmiXmt00l3ZQFcxjboGrHC6tsrCAkMdeDRJf9uX66Uvf3j1MLoiD4W30Y2yE
WI/qZkoQMzcfCi1o2xjbUGj2QTOJRbbElWe+W0886y3hXTabo975crggAjFGijvOS7XFU13f8E5g
iKg1puyHVgMoAD+dDxd1PVtCGtswp5XhJxUD7+kZRBN2i+00mSdm72wGJoMO6rEAy64byquY0WMo
uXXKrscTzhIEOqwGoQKUBP3eQGtZqCiIWThe4ZVK1wy+Vw6mUDYlQjygoI3jIEwq4V46XwkMisje
wUzw9gq6uxf8NL1T+kb5zD9erxx0MBnp7UPIs4pApU0dCaCc2d94tuBVD3qjxfMClq2+T3f/sE+x
RGKRYdQ68DvQyoY4pzTSaRStp8bgZxm4DqU4z4wg4M7JEb/Gnf866wBAVZMYPUgWS6AvSymicCgq
1ylZ5Bgfhm5A/xuO8wa+yp115fiX+skgXJrdp1fA2gFYGRMVkTrT6xJs6Dz+ZylSMaAi5Qhi4eoc
TwHHKzfs47/hIzOSdLfFJ8ZyDppqnFGOL9061llZXgsXdgtlDZPNrnA6oHmGOE3MVxXQpdx39Ppb
0dcJgyXpQmKPwYzSYzLP7dnopJE4NGGnAKWiLeD8AkfJ/iiU57YFrdRo5S+3y5eaW7De0jeWpYtX
1PFcoqSJQYPLdJwRoRYkDL80nR/dnxPw0gNCkwXHVAP/Cnh0wZB9S5am19TpGLaJfjYoUf9GYIU0
pCVG/XL+lqU0kT5kNt9KexF68wwqOlCLPXcgM+SLdGa+Z9lYIL0lz7cfi56jZCcbObIl0r7qMyyC
1crUKCjLHXWKnCKFNp6OaZPi6aOjY94hFqwA6LCHB53J2LN+IU2q4GFqiQ2ZNa04xhybMXN7XlUQ
smBTETxPEYQrs10N+ZlYRksx9Vpgk4UF7iWjNaVSn9uv/Cj1Et3wujIHzsEJ8KJEOARsFo6Kx1GD
8AE0EoN7XTcGX4O3Q4d38hY7x8TX61pjbRPtwAW8b+4QkMEna3AoYK7+slmWblQxUvfWJoz6p8Xs
tdl0mK5emafCvlps2CduSRHBQWgs005n6la6bP721KXPGPn3R7YJ8toG+iTYNYQm/O88arPTuFMv
oSwYsuU3E9KMbj0+Oj48AM4zdlvQpv4rwSGlSwMDcStmB1XoJZEYhTNv5NAyIr02Dbor6pi3FOiH
NVS0btu80c9NM2a3TMmQEFwTUKgl49Mbq8+d0eMaG5alHBIoFSImpj3tW0RGm5IjBjOFDOYnLpf+
ptkDwtePO1Kd42yY3qTE1ICuvM77Yz7Xwp9pOc0egAC5Uum+Rbxl1blIyzG9X5Fl8Ct3HBGqsYmB
Ogq4s48QAvucI4XA0NIL8+MClevQ1C0fnkWeTCEggbDsdtkg2gtaTLAGnwmVAYGpER6qZD+qE77f
W1pu9XZ4V9l48BHFdRmrXsho5K1AF0/aEGTOl+5tAcfLCrjS+RmQOAO8p2DuZ2atnzhNAg2MYRZE
eZldwr0E024iFQ4A8SIHSKlmzPBfvk3vy0Q0aNOlr+0n9fjS6rdHnl+V2qlRVUEXcT8hCpaO8fCq
pLQV8iK+O18ibfn/PApQgJAfi43zDEWCy+xfZ71SZxnGMlVmyPlyp2UUT69CChGTRgVyiJeCYNw1
ULUhjqytU3Gyzl1ENlp7BB8l49VZclUZ1C/7q1pRNZRYF0QZbg4aaI5TmtpuU8q2iIau7R9K0FIL
PYTuAU1si7L1gXXriJ3DDnuSmuAKFNDK7+5NJwv5WEjxjkpnrpjcFJwKBFxj7Ru+EJJrcH2tgO/b
LjZN+FuqXe+i4yAcVP9Hbi7ezWk181SpJTXcWNSixBFi3MVFA2cIPBRAvkX8jFyNe5KO/Ddn3lh3
crSIffxBg1zt2joDlhfHMYCzxXqhA/ZWFtwBvJhLoF+qNrYBhgsr/NR4zt3bA45FWS7JYh7Ljnsa
g6XT2/HopUlGa0DVUlxUV3UtroxNkh3P5LUOyIjUcASSywomrkCyQOcHKJbm2iJltf4fOGeoq0yx
YF2apyYnvl8WLLj9JeswOjXth15PjcUXvELyzGKIpF/xQogpTtvZjEoEyieA1EAml7pkzDeV6QzG
N33/I+cacBgIDazLaj9jd72Gb6b6+vo+jQXYHWzDV3C9nmUO9hdT+XTDy1la0/lvBY/WgRyByVox
U4Ms737838C6TVO5UWaRtD9ExTW4b+E7kSXjP35+CVoNfrJ6/8nngQ217bFqBBw1HGZ8oqx0Qemy
dxGHZMwD/2YbnlYV77eKqWWPH/c02cWcJLLDK0yghyWEnRxkeKv2z1/o7M4lhjDPHVOcun5o3Tl9
i24v6SrB8LF04pYrxxUofuzV+78aqwrLD0oNzHmX42rbV6/ilw+NNx9XBndRQVwCQr+lIq6YWPIL
9F+arD+RRWdW3v2mZZCKcM+SIhm4XUxP2B0O0JETQgTX5O/bA2Nn2pMjMwoW8MpwJsRCEN1WHw1k
FvPDgD0ZiC6MufvYk0CSEop6L1jvj5FLROWw6qoUf+lVNoOYlWG6lbBPKOxczvOKmXnODy4wtmx2
zaYYoo4Avs2boUVWb+MOtpWLY4+nyHvcurxH4am8vqjSttyRIhkkmQ3OR3qcTSmUCVcxOErgtgxA
9wshwFet2LRiubnN4ncdAyMcON6RSAZN7MUI0Gt5BSGVgzJTAp/PfBPLWuQOt3EpJdddpVKw2C6W
gdTrNxaNhts+hHXXV5nsVaLAeqY80ZjATbDXItOmMqJwkKaifpiQ71+ZcJ0p+G5uh9pV4e8VHf7U
SMafQUCCc0YbSH3t/PWpQQ+1SR3PzUdxaUUasbeZt9Xap7mXYJOhEy11y/+w4xBcc3QsFYN/HUm7
NQ8umZ9g6jfaYgCs03gf9iqYPAiebyTWnwH77tHopM4eV9Xp5rmhBYNJ3CSoM1fgttXy+lEdswFn
gDDN3ZHTeqGorzKA0AlfFWU6y1fgowsMllNgZReNHU08xERjLVWuYvfn15//v2TRJAT/z8vpWg7K
U6R79DPxD+f7xzbwx8BemGY/z8DaZfOEkLuiMgaP6DV2VvB+0bl7GCI6qSMey9vPSTNJ2jdtZAiv
pKJ6sCO21WV36djwUHyfpTffNcVmZiT0K2My/fxvMCZby2riG+WxppZn2KCC5K7NWvU7aoFbK2q3
jLCyIP5iPzr7zjkQju4FKzWgaF14eeLAmh02jSlAn5bvzw56nAwXpFsMPyPJMmTsqNDJC5mBm1IC
YYyH7AJ7FTXo3kUcD1wzvhBegjkJv7QhUoVuG3DgutLDdgSF2gBmjCg5j/b12O/HRPHXhoefD5UN
Oe1Ls8QVYefXgY6JVmBe2ma7AKuetVYW5r17RMmrxeUxER8CXXVYHdoF1DvcG7tqLGDeQebxW120
4Pv7z/plV253JnZ+ofE8CORn6TiPSe7+kpzaXbOyEDSJdSN7HHGXnCn+0NyeYVl4+ZLDitdHWHlN
l22EXFT9f4Fh2ndpc7fU9Wlknxk7HbsiPkDY+UcV8ivJ2mBJ3fjnQnugaqoFrE4RZYCYk3UHyhsk
0RP5M657w3ZUkvwmlsAzYX+L4b0skzeS+TYDGviZS3DpoERI9ILMxs3Yhf0XyiCtU0DRSYWrYXPe
+tTyzGndgf0EkrGmE6AKTnn6RV6IeRxmkPVNUxsHwqBElIOhgBoZ3CXWTjgGC/YYsQt4i8oe8l3j
DGaGQbIbzw/r70lmUfD9/W1hmIuIar0hS9KPhV9s5sX9+yZA6UQFDJ/DZ5v38xdMzSgOsXlpY9Gb
YYctxJbYCt4gu/41B7j1P2025CZ3f+ErCD6F/ELYB/S364k1UjjI+KNgLrif45p/Joj3c1ORTt3c
qaLvs/jVJpP8DPakQOO5OK2JnhEVZqZlg8CR4hBM65o2xdHD7697qf89WzjOCTum7N0SWGLk+LkY
qdSaeQrVCOG+f5bgNG/UlbuL7GRsZncItU8IBbev9RpYU5CJsPoTyqMm3y0Z1VrsWKp0PpYFgi5V
4M4KYNaMATGLzmvnssELeHrOdxo9qTeHqlTY9ONBadSlkRID8REp1tYqT0AmZkWK9//S1wOoo95W
LBpil0g3Edqv2OZd8Xa5LVQMRdfZsEFWi8+YFaRW03QvNv/Xg+QR70cqp6Zh0J4jidt0hU7ptWzG
Cks0sOmtO5TZ7UdsiPEYCMajWKPLeDDIYo0tZyCBdHhN2zgYSGTVrnXlWxQTHW5FS50kpo8eUIot
3vKEUsV22B0yLtfZ8sXmd0CqXnWo3fk/XSb+Mw+ZbvNACGI15sL0ZBpZnspaP3KVkQPFUZaMA8Zr
iWSaOMq+gCQIf9KhvusdEcqAt6mM4i63OmfP7ZnKZZEQazbUuBp1cAlObcW+/4WyXwW2MLBUaJPT
uBrTc4XK8CjiEAZ3fzElEI27ZVDQoW/Llel6
`protect end_protected
