��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����Z@w?�=;���:D�~B�~[��X&hd!������D�Ɋ���Uj;7oP*��Q��#� @^S�ى\V&�J��0=O;�����6��U�AZ�� CěT���ܶ���AX4�����d�����
�邆]N�!005/''Ӓ�ޕ�J�=-˻+��%-������p�t�]x�M��s�'��-�֌�H��\�ѷ��	U��;v�Z�Fd��je�O���/L�~�A�1KG1��a�)��W��y��p���3ݰe1)"G��� �n��!��4D��E����3ȗ���v�%�� �<rv:�uA%��ڕ^=����4��0�=��.��P�	��阫h�Mi�y��?���ܿ!Y����OkT`"X_U3�6�N"�I�����`n��z�i�YD��[f�S�zc�1���=U�J^5��Ё��"*�訁b��:��^(bybOO%�h�w�`7X��F/�k�B�k:w��kO�sb�׸�c�a�K�5���)��4�f��#�H�ly��\U�0uv�v։���L�-�6?Z�s���E'Y���x�����i�>�p��k�] KӰ7�N�7����3��ܓtN�x���,Fb��s���M�x(:7�=�̍�}/��[�,G{q�T77����wi�Z/v��c��MG<�:1d��*n�"'ݚ$Jf����/���'��d����#�hgO/�=XzQ��|8N(A��x�/)g�)�K�S�l��햻�[�u�Fm�)�.4(r�����K�%)2�NU��T�?x^ݻ���j�GD8���:?�&�<L?�[������~W�MZ��J�L|b!���P�m�Rn�ȯs���}풓5���0ee����V%�����$mi&N&�o����r��@� T�(��1��'��1�)�=����ƃ`,�~�|�Y��i_���iЌ9��� 5uS�c1���1�޶� o�w�4��ҕf�2�H1�fIB1F��	�3y+3;��l1����>Z�v�4����a'�w����Æ鸡+�o���]5�o�w���{� �Bc�"'q�MՖ~/qz�vc.v��J���>O��c��������M����m�
o�Tn����;3..�0��2*��K%%k�B��w����V��Ea�D�ә�}�~��0�!_�t+PR����o���� [ 3cj� �fǧX�����'q�.0�&Pre� �1b�J��
+��o�9L ��Xc��w1[4����'*ތ�l�!z�.NΠ~f�г��vBP^l7�|J��
r�D���@�P⡘�Q6ז�W^P�hD� �q�~�_�G���)��EO,v�E�sG�7��������C�Sa��S�ޖpy-�� �:�U��Ez���$0妫g��x���ov6T�9�+�k�:W�:|66elxc�잰�U�3�sk�xʣ��C)��-��?WKn�b��(h�k�R��������ᆻ����p� ;��B?�o����2��o#7qpjO��-��BY�?���z�*�����"ڝvMn��O�M-���W��!i5�*�%�G����L�-��7m��Q�{�ĪF��F^w�)yX�Xʕ�/�K�Z]�qZ����@�l��BQl�����k�K9a�}��t��w�LM0�Zq,o���v�p3�6)���������ޫ7F�LW��~	.���]G@o��2���f��%o�N��m�E���<.�Пi�t#Z���ź`_��/E�v�6���D���H�Ycn;��Ե<pڢ��)c57��{��YH�����6�`����:���ϖ��.TGa��{ִ���j�xd�UI�y���3y�(��G�N��|Ikdh'�swd<j�2W�mб������4���	�@,���Tf��6�֑��@��A�*π�Zx!yv;�*�LR�m�
L�;|���.��]��3D DR����>$�}�{("dkf��QO�"l� �'9_��,�V�y
.C�`���r�nc�w����H����dGp��u���%�Y�V*�@B�����.�\:���Ҹ�/�=v'�x����OQ{|11��^�!��
��K��_&�eL���ONX)Xf�93M|�Qʗ���>aB�UҵQ�%>4�.L��3M��*�v_Tǋ�������2����B ����mD�EN�����o�O�M�G�A�6hWP3>r1R�LܓxE8���ԫl[
)o�w�=P�u�I��oQ�Alo1Tv�y������#��V��b=��l�*.d}�&Px'���������q!V�P)+�%>������%Q��?�|	]�n{ƺ�mG�n���l)m8� .5��|*;w�D�4H����h�9%#��l�!l����r��ՠq���[cKr����q�U���'P����9E��N�,clW:�Sdt9����2��w�h�~kEG����֨5߯��JġK�E���&ǢM,%Z���������c�AТ��`����|�)eV�=Pd2t��*�fT�>���B�X���hG����EԔZ\�}C:fP=@
y[��u�Z���[��e�UFXI�c�TZ�j�
��V��8���Ӡ�����NW��-�d-
:W��֭|����]�}|����w�L�㉹'?!?VI��}Z�lJw��FIT�+-�
�z�����s'\�tshr)���24�:��D扷ftc 5�p�QT-��F���5��:5�YP׬�B����<�}-]�>g��To�/�΅wXM>_������{\c��X�$�_�݉Z�H��enK+Y�G�nX9�T26
�1&|�x�Q��/BMv��4�L^{�q�3��������ܪo+w�C�yC־t���ѵٚ��*3d��q��78����՗k�n�g��l�
�5�ZëDg�l��y�tLx�F�`M�B�Q$�"����~ޜBYA��>����6���"�֒t���to�[¸��
d�u"�<�k-
�╺���z��l�R�F����#B#�Ϙ��XYV�~RHa�r"������|�$��Y��u��|���C,-�6�:ۚ�������-,�h�����z�,���&�l���^�e�>�s/�GP5<� �Ej~;tk	�u!���zp\�$�n���"Gs��l��\���T��{�S��$ػ��3�Bź�K��}T<NlSJk��l�1֙Z���'�n���<��羙w����+2�����g�P��8v=�����X���I��o�@�h�
��]�Ȼu!�.?�C�Pe�;=�H��!��'�`�`G�<��-)c ���ӭ��X	E�b����Ǯ6����Ѳ�n���;�#g	�,e-�T��x�Q�|_j�=4�J1��0��=�f��K���Sz@�0c��9�;��9�?�R�o}5T~�\-k�e�W�/C�6JwP�D����!�1������Hq�e4]��V��;� Ώ��*~&1�#%��t�Z����0�K�1�N/�l�R���Q�|=8��pj����[C�!�������ǯ�r@��=�胲V(���	����Ou﫾��xl������$F��H�A�.�B{axs`m��s��d[�"@�a9����P��!��A�,=0�fOǭ4!��_�/b|�.�A��ӞY�ж�G��l���vz�~�ʤ_�5,B*+�Kz�@��c��n�pۃV����_��$�_��?R�\�g`�;�z�l7��4���x�Z���C�^]˓=��2�.�JL�bla#�^�	�&R[
ЉpV}o"�ޣ�8��T�T;{�L� ���Iȡ�����K�h�=�EO'�C�no,�,	�e>�j�"tc�{C����^.2Ӟ���j��B	�u��d�(�M,��A���l��^ 3�ٓ� '<�b`���pS��
;�n{��)|-c�rʠ���n�����%��a(���|γe��p%^w�������u{X_�!�bi�}+���=���7kL�+�2�#"�	�����~�>�A�ͶW�z��0:�o&Qj���I�[�����1<N�>*<��q�y���巫���Z/��E�V� ��P�N6#NG�Q���>�~�p��əɚjޤ��ݡx��r�M	��f�[`�iY�Ui����R��te�L�j�z�#6���]CgƏ޸
�d
u��N�*�nOhM�!]�s����X���A֙θ�|�0݌���z��������Ʒ�#
{s�6Z�mxZ�%[=gטZ��G��u�;��U�f�Ze5Z�	SR|[Tˮ�������V��!���,�!�  �::l�p������U��UYY��:��a����7w���R]�}	��M��^�+�z����z�yoT�"�S:�K�	z`,Hd�	qs�t@q�q\�RZ�?����1l�!T�d�=�mUpf�|�aZ��ޗ�(_�<�7t�a������Zb/��8�垖K�i��"Z�P�
3�S���G�3i"o�$�6�h�U���������J|d�u��0ȋ3��H�X=S"��lr�U?KE��V:4�ٚj�@�b�}���g�!sT�'�q�ՈZ���a�M-�|?��[�my���@��VS��A�v��q_���ժE�r��e$��L��D��h��^P�a�)S�.��M�.ƙ��m��Ũ-���LsD�aL�Ko�`�79"�����7�Λ�:�(��%�����B���Y���i�A�i���%�<���M�f��C�o�54�윝�y+6�蛔�^pw�z�C�q���7��!Q�O?6�5��?�}#�М�|�h�A��h�e�(����vI�h�#��Ll�x3^�?�L�	[����
�ha�X�6@��p~����|�c��S/�!*�z�*`��L�΍�I��BC���f;v7�kƣb�F�up�{�gؐ�Cs*A�pU��f��y�ġ\�����D[��AL��ʅ)K������}�`3�&d�9�9������I�"��-W�6��+�;{��C�!M�~xO��b�"'s��aQ01��X��6
�ŲMUD̱�U����8{����in;�����~�^/����j^B�]#��%0��i�,"�B�����\TgivSY��n8K��HIn���g����Pg�v���k~��ٯ�ݼ�8d(܋���=?&O�M'�]���V���@I�.wDj�J	�T�.�۱�xA6�Y�:#o�ob/A����>z�G)����U�쭖�=	����+�l��E�[��C��>���/�3D"���i׷�)st� (�����|�'��2���+��CY*1{�O������0Hz�oC~^|+��gzt(�}�q0PvU�*�^�	п�eκsB]܀��:J�`J�����x���� �t>ď�4��9�y.뜷-����DI�Wȴ۞���V
�"�5b��]pz�J"p�L?�*qH��R�-?�Y�>hk��m�۳Q3 9c�%��ndq�B]������05�xv�� Rw��L��c��:�G"ߩ�~8qy(4yZ�C��B�o�\���271j_�%�:�=��(so^�3�H��į"��@h���\n$��6�L	�:lI�g4େ'��8Vb.��b����w��.�=tfY���u�~��Q�ȥ�kLІu?���ey)3};�k��?�a7�O&܃��(-��Js�M��m�[�߮��6È�n6�(���H_�D��B4���B)�1����q$D?:PvQw�J�RQѹX+��A�id�?�ނ�GLxxU+�8���
�x+�O��O�u<�7��4��YMZv[�p��AM��g�e5@A4���\��>�"���w\�&d���m�#
�8�����X�1[�-!-�]ڨxw71���g�!�i��%�:�
y�A��+B�3�Q���e�W:�����j�I���+ݮ.;ťy����$V9дP��5s�@��6^��������P���},�Z]�|��I9��:��0�66�2(����Ѳ�Ռ���A)��p���
ln�՘,��
 ��	��Àj#����:d����U�(9)�Fw�������� D�?�����{y"����������k۽y��������lk6E����GS*F��i�c�B�7��Z�+���`�M�,��3� ?C�&���C �6�䆄�ߍ�ΰ�1X9_,O���!$�Aˍ�.Qkp��%
�i���l@AkWDi�jh��L��VM8p��݂O��-'���5-
���A�-���n��|�1�^o�نo'��c���h�1�	���f�y/B)Xe��d��4K����\`�c�R�[��k�c���(�-�y����Q��yD���rqU�WIJ�v?�9Dː��l���c��	�����~��3۽I5�ӤK/BH�u��Q�X_�	���uޣF�WD�l�	�)��&Ʉ\�i�[v�M)�9{2(���	?$����1�W�%va�nAû�kr�ϛ!��v������u�0�] z����Jꬔ9+K�
�1��2�Z]?��g���+�/@�����L��& >|{�����q�H�ކ�.��� �)�����W��|��i��M��׏��y�`J�r�)bA�ǜx�oQRpH��&9kH�ϻ���K17�ʞ2L8�=�=�@#��&��2��%t��?7b/��=e��=����n��xa��$
Bm蠔���x{�|���ԍ��Bdi��}ư���b�Q?w�#Ir��ryXp��\]���<������B��f=FY����6�����kYxF$��f�YB�O1���*�9'������Y|��c	�qaH��@>�9Tr��H��׽��{X��W���[K�쒙�Y�Ԫ�h2H<X�"�T�˛�R`�g�����ԴK�=��	X���!�$M������:H�FӏB:ྦ�:�V�N��m���M�����S��{�u����v�X�7 գ^&pNBy|��Ex�d��	;wYI��ݨ��ۀ��2�ț�Á�ì)�YtW��}�y"�[Za�{�ٍ�^�)c_Μ8��� �`�{u�K+�jޭ ����=��_/��O��4"t��������j��+ʑ<�!nNN�@� ��T%j������J��$�H�쀙�ա��4����@u�c3�bk9�:���y8#�x����.�`W������g4T2�m�Kt�͡�/U_Q{�ճ�����"��|.�4>R,������X��4�3A�a�.���T�u�it�v��|�@��<���N��ԋ��|��X�vZ�M>]y