��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ь��-p�l9qe�p}����y��L�Xݳ�,du~{�/�mt't��UUe
�"WJ�>��.���as��^�o�r�?�>��{�z0�2|K:������@�����q�����ev���@�e����p��d	���v#�~'w)�U[��P7��nF0eҘ8�^���S��z�m���x�/�����tn�Ud��n���jv��Xv:L�҂�p6��iQE�Y�� ܢ-X�����G�^z��Y��|����]�b��E��/���Bc��@�0�Id�@dQ]� �HA����VT�)Y�.�U���H��6�<�j(������6�Fn��,h�jj���hc����t�VK��iH�}f�ݤ^K>D�ia]?�1D� �0����X;a�&{N͉�	��~�M�א��lęB\�a��`w��uf� Hc�xv�p�y�<�~��p�	��3���k"�0q�UF���:�S^��ǦD`�s(���3��=��8���sd9��#���g�3��j�i�N�r (e�ɸoȁehy`\d������p@y������f��/�X\��b�R��7�5���7���{*Ȯ�U� �Z��c�"A.�"�OA���Ǚ���K^����1G���k�k�����J�Q�`��oaC�֠0�����cg����v|Xv]1E�������"�wr�9D�[�w02�!L�#RV����M�%���ߎ@�z���O|�D1�H(��J'G���BL^�|����^7�׹-�խ#�F�'���L��z^��<�=�o�5���W)� �� =���5+]Y}�[sR@S}�>`Z+L¿����V��v	��
�K��\Q ��������n���ì��ؙ�C�7���\����cbh�	ZӴ�+ �����I$�bL>���������NK	��5�0X�(�� �2+!�������4��(c���0�|�������[6U�5L ��&�<7�y�� Q~�a���C����!�-��	vNŭ �ƚŐ�G~�v�|` ���N�x����"�d���o�$q�?��	?����B�mFI�5��R &���8%|�������ۃ^N�j�r{�^Һo��5��=?������t��挏SRO%�H�AK���ͿC2�<����$�51��`��g�  ��7�=4��!�Ln�%�fP�E @�{�F�� ��$Aփ�i�gά6[�8�q�&��~�?����2�@�b�_��?�!�EZ2���g\טӨK��u��0�o��ͪnM���5��{Xb6h�ы�{��M!�(@��C�o+�3�Ƚ7[�e�L��=J*����F�0��}�
p�i$����`9z�-5�Z�
��gA`�7��ض:s+������)��P �2����)?�4A�|/M;k��7�ۮ'��k�%s�3���;k�T;���V�B��[�nǑ�X|!��F����|� .��l�(�#�y,��Y)s]g�%�a瓇e(��v>O�b"�N���Gp +�v$Ç��nN�������z��\���_^G�=��ay�Y'��1}q�;_;��2��j�>�\!G�ϛ4�T�k^�qt!����ze�?�Ƀ^�Od�%C�ꇀll��5�Y�w�K��x̩,���A�oFN5��j���d�֟L�|Q� ܮb�w���}�r�Bb����:CL�7I�f��R�,�� ��;2��\���k��+"'���z
�m�����~mQ����࿌.�o.j��?�}DѨ4���H'���&(I�'��Ps�R]�:�m�X���TTF`����p�)^U9�"6��lƍ����z�CL�ӿ�ʍ>V�R/P��%�`��s��d7�v];�m��'�4]d�}�U�ӽp�2}$Q�4`(*���]D�0|��~�GLB�s�@�^��m'�]�,�#-�h%y?�/U6㤙�y��f`6Mp�ٙ�s��A4�I��׬�Ex�,v߻�WY���Ы��٬�EvRr|ܱ}�
�m�03E����x�ș�N+����GX:|�d�'��T��)m0����+���'9y�J�ٟfzݑ��g�Ї����:&���|����'����k���FH�|���!�%��SH҂y9R2�|�\'�+���t�m�mRqӔ�D����4Dy���P{d�0	z߇�&⁸@t{ 1�m�AN'���1�ł��	������'�!��&A�W�lWCʈ���@s�}q�{�����s�#����[����k���^��x��[+vjR��!����D�y[��<�z�z�͓
Z̙@zB��y:ܣ<�q朢�l۰Py�Z\k��f*k8µ<.�ʌg��/��~zw���Q��"ڝ�v�'cn���C��sT���/t����r�脭2H�mmn��`��oa���*C��t443� �m��_�����"޾o�����i�aD{��V�9������j��N"�0@E ���Q3���֤9����`t_�s��.�7懽�PW�f�9����>���ד'�nY&�.Z��2������Y^������D�!CC��L�(��vֽS"�Ih0�%��ƾ��{?��Ř�?/���6��~,�Ճa�3�-�b5Js �B� ��z���*�A�`i�0�q�ݱ�Z4�۝�|'°���A3eq�Hg�E� '(*����Y�:��g���O'�u7~#:�h-�£���ՏE*�
E}ٺŶR͉L�t�T�
:S�v��SB]�J��!����Qj�Y��:�ϥ��r�YR�u�1�x�|gT�B/C�f/_�S{��y*�O*l\�wB���f�I���ݔB��dk~¬p��9oo�'c�_���7DԳ�KӼ��y˟���f�'�lE'4c� ����}z��ѵ<������a�l.pwnWOZ����y(�������I�w�tY�TLk�?�\�Ϥ*�����'�{`�!䚌4!��"!�4u9���6w�0�ʲ*��@[D�R1\��u��LX�-�,�B����� Zn�� ��p�eޢ#�>-���\��T��10��b����0��~c����5O k3��/�3Cu�*�wI/���Z��k�\����?T�6�d�[.��H~v�6��Tk�.��4Dќ���:&K'v&>�FR4�<������z��X%��i&�J8\&y���9
����� k��2�Ӻ�~�Vr�5���kFj���Cڜ��4�g�#�+Q�����|���cO<�����H�k� $໷������^�Г�ޮ�0�"͢��/R�E�bځ�%�=�L��r���KRέ(Zh2ij&Q�^P�)��o�_77�Ac]�V�� ��pq��V<
��T�'K��d|�Do�9)���}l��p���V�3�TN݇��t�?��԰�.�bq����u#!�,���L��Ma��-V�j�����0a�oW6�L�T� ?�:�^=�b�pÒe:�3N�e!dokL���<�@��ě��(K��YO�JM��9-8'�I�үM�?�tkt�6��SoS��4#�J<����S�9������`�Bz��j����;��*��7O7;���Շu��A� �C�/Z��!�LP���En�J���o1��Xm�����Wo��I��7؍���
{�������x��n	ɪlu4�ҽF#a�s?
�#�����Ss���C_j[d�!q�g⅄�Z����|[wCp2̚����{jK���2;�%��蔞�����P��>|Kl�/i܎�])s�L�v>䖅��PZ��O0��z�,�P�gtO��IW�3aúq�{چ��!�$�=W_O2{9b$'�8�Fu��yCo]Dk���7�(in*V�V/��iDA~���= Sٙ`4NƔ�{:1��uT�f���"`e��|l�&��y[����PeG�F�p����4��TȦ��~7"�9RS�DJg���o�7�,Ңϼ�������rl<52'VX �����$�qm�%W�	.,�ϱ�%�1�8��D��:x�`�����%+�@w6�с�&Vj��r���uR�Iw����-z#4x��#�Ѷ-8=Gm�m2��*v7�Wt���zz͢���ɠ��Vi�Z���KW/ œII�g�����J]�fgNB�����宇��"�R�h�x��)�O�	B���/�>�Q��q�(��ҡc9//��b��>�U5�>�q���G��B������(��8�N��Ѓ1�9�M�����}���/�h�	Z���h&9Tl�7�8R8##�_������m�>4@ח�I*�T����&m��V�#�oJ~����󱹢	BE�Oy�Y���w�L���-�+��0yAB�Y2>�X��08�g�A� �w�e]�V����	��4��%1������"�tH�q�u�N�䯳"ZA䇬|�<�(h�s�eR�ۿ��]%r&�wP��q`��}�!�'�{6*e&qۇ���"L)*D�(М��/���Xzj(��af�bY^���������~\�)��MA�5I} F}�e�Zǂ�|���%K�ԟ� p���������`dy����UV�G��-�NS�:�T�CU��.k�nS˨�g�>�����p���c��I/��46c{��B�A���}��=P���!��Iv���HL��Z1�O��^���B�Ai�'֫�T�f�� s�C��$$J�D��|�Q	���Lk@trח/�{�@|T��5d�Œ��-w���̥����G�Hx6����p.�&4�v�_���'��)�'M�)No�P��k!�[�b���*ȼ� ��*P3��i9��Y�*OOu�t�U��n��P��|�/���@0$o����E����,;y|}=�S>C�uh��pЭ��m��}њ���J~�B�;��:*x��ΰ>@�R��
<�)^
/�8[���q.�L�wL�����q��izs զ3>>�o���?Z��U�;�j��8P���~�!{ɣ$}U����/��C�>����[ �g-�k̕����y�v�����B�/;���=j�|���;���M�B��mqfOOB�p�ץ��	40_���~;�=y��">��dBF9^J��:�I�WT����v�}����8W�����k�`���Y���LJu	���H�R�\*$��M�slil�zi��jo(�G.1��L���Q��r��}�^*M��"'�������=Ǻ	�h]B
��Ӱ��i��]�`/��}�i��7"&�HS�uK���-���b�;F���Ua z�;� ��"�"�*n8\7	��F����R�(ve`�S�l���ڏz5��#+�����l�E���1�7.�/|�3�d�f7X�:+=?-kr��0��v�4�-�9���|1�޲z���8��,�cm�jL���~4)��]u�rnK��y�+�X�I<��Z4�gQ s����ڻ�� 4��������/���z��$�[����������E�||O�)5�=z�F�|

w'�X���L���Oq?�8�b[g����wB�m�_�cZ�$�{a���٦U�2`ɘFCS�&�6ɦ�$��]����so�����
���5^:$���x Ǉ9�tF�Zb�����+>(
�0b���zW���YW(�,d��,�3ɜ
�2�5rІAؘ���-�W�_O�bWcll�=�A�3
?oW��3̿3B�ƻ[&��%����� +�3���Wz�h'T�����g��Y3k?H�f����^�z*��Ha��Ⱆ���#��2� ���&zr�]�Y��|{(	�S��%����+mp��YL���:��[8/���<v��v_�3��Y���u�ޘ.�in��� �0�*^Ka�qBV�S����d���v&Uj�����֛CLh��2D������*q#�V��4�79}�T0F��Br^���xp�sv�����\�ù�U0/�r⊱�#�t�t�~���Ia�-�߉ε=��p�dq��$*��Dn���ϒ�#��4�o��}���[�S��jT��֮`NT�J����6M8r0T/�gɷ���j+�����̉"V��Gc�.�â|����WY�U��6|F��I��5w��8"��b�R��V��I�	�	)�yg�DQ�^U��S��ю՗vH%�3��Ŧ���լ�T]�r�q\��5=n(`���8�3ď���Z]L'��=��N+,�؟5`N�&�u�6��9�k<������8����*�B#RA�p;(�vK��g�ࠛ�X��+���9�Z����H�Z(Vr��T��	�7F9)rZ���Wÿ�q�1�G1M^�'A�uSdA��4�Oq�F�#�w��~3H���\��	s}����X0z2�X;�h@n�Sd���o�t�n1��Z��;�����9WGɥ���ޙ�f��d�x���� ������:��D��z�4��=o^��+��f�;�݂a�	�n�k8⌻-�5�	kqaBxy�"�$9� ��r��u?A�D��eE��m$X}��xsӋ_L]U����Ou�d���^����4'�E������r�Q*;�	�Z���;�{�9n�
lKS6�T��{t�_�p����Q�*����e�V�N����=��V�n#�%��DQ��� ���O�5�(��%����AJJ�h���z�Z�i��?5��۶+�?˚��� ��U�R���t�x
���s����5F�-��=H6��Z�Pm�����Ԟa����FԸ�4V���b���C76Y�qf�g����*���0ވ�܁����Q��!&�A����.�q�}�L�,84{�.Lp�X_�P�+�8�������a�%73�Y|���ug6�\e�/ �>��n36q�{�@F����؊]M �p�+*����2 Q(e0�+�,���
'����7��B^S����Ln?�Ȑ!i5��Óv�W�> ��p��փ��?d���֙Hd�3a�i����`��$2e�[ew~9�K��}�L�#��ǁ�#����5m&�X�W�b�n�w��,�ޛ�ꜹ��	�>���#�c�_�}}K��f��q��T��y�y+?�R�Y^�9#���w�ef���O����'o
�z{�N�~���R�d@H.�Vdz�������ȥϧ�}��Ύ���W���݄��M�����[Rҗs�}d�:�z�����NRz�g��zu��)�U��P��k/����==�S0����H~��j�6u�+�k�5���[m�*�/K���E�A9�ta����-%��r��R����O�D����һ����RA���B��N�zF1�O�Vh
`�0;>���� ��{��(�PZOl+ BP%Ǔ�c�jd� >|����X����3���P ̂�����C��uZ;@5 �T��+6^7��.�� s��8.�g�A���还����(�2�Ń)�k�S7��+I{�~�n?7��[:�
��jɗP�2�a����3E\��<@�9:�ߒ�^s�k��vW�j���Y�wb+J��e����۲��G�l=��Юa��"Y��ER��a�TY_��o���Gv�|��2�)�t�&͢R�IP��k{;J�����[��%����2N���k(��������'B��D:%�^�r>j�j����˱�d�;�5���?���1K���Px$	?��,�0����#���`��t���Q��z8���MqP|'�Ǵ �n#i�$��QR�va��(��^\k�1wD���e��;��:( H���$8vh��v��g�U��W�My(�^:��a*J�i]}+ƽ8Pv$%@a]o,J�v�p7�=]�)��.Cs�4m>���H�#���S���v��7Ԉ��������JXr�A��)�m#���g6C��<M�]��3q�a4޿;��-�_�!*�Up:e3;춳�
��w]�z�[����+���ù�pİ���l�~a�1��_Gbg]ߎG6�znF=\wr�jZJ*��"8�ޛ�[U�Hb���9^�l����o���~"3�̚)��ƣ�nj�r(yܻ��_�.�����]�Z���A�.��,��j�(��o�ve�_\V��M��溘�J�]�FA���kDw�0Br�rE.>YX�e�&�!����D���� ��+}��.�2)�E���:I�2�~'H^�;��W`����%(jezcb�el܊����^>d�.�J�6�OJ�Ն���$��RJE����B5��r���F���*���hEҼP��D*$�4X���]ּU��N A×��؈�Uޝ�PյsKVN�i!�j�D_�h@�0f[�g�s
v:h�Ћ�]:��0�;B��C����$}�υ{��#6�4e�25��A�+Y%	��#.w��2ƿ��ee��D:��7�VI�
�o�u�?R�~4W~(�2jB/�bK��{�ȅ}�ڷ���YqYmbd�M��o}�5jLh�*��%1�c���F��tA^n��g�{���g/k5�#��vB&v��@_�����%�5��A5�g�F��%�}
�Z� ~j�ݠUo��,/����.3�<�jƛt�p�3�1
M�_I��_q��?��M����8'�S%�G�/�~�}X{yZ?4� �"�#h�ja�X�M?G�@bY��uz��)�wAf��Md���T:���S��T˵���8ߐ��rl���5��T�b3�ڻ�*�nu[�!hM�f��0Q)ΖMa˷������+���Ɍ��-�KF��:��ax�g��5�Vq\�,��_��#(w��|�Lf��WO>'Q| S���SY"��Gˁ˷`ךG��3݆�T}��)��*\킁~�+
�T�a
�����HQ���7�@��Ժ{��O(�7�d}�g���n���8�|ʲfږ��<uY��e�d[945ĵO��TT��ȝ�U���doV"׆��:(����Csi�./!<۷0*�E\O��oTZ�O��	'D�BB�G��aT�%Ç���"�� ��`)y�����O)���%�%[0����q'/�[ŁD�@�����4��P���	-O�翞V긠�f}e�W[_9�W���Y��3}r-j'j��<i@У�d�rI�T�S���B~��_ϐYt��~6c���|*�x�S�5z�7���ܕ#���}�Kva����<j�4�J��;�2�]����_n8WpNB�>M��m��.YV�tZ�����w%�M�X��e��3#���ȉa`z����^d����+_W���bO1 ��Z�
�J��P/U��ʦ쑞��j�d=���cß �0�z}�+�\�=,�`p�w���>���+`=���W�9��E��x
��!Y�Q{�k9�B��6��o׻�Z����BhnCI�+W6p�>}q�Y����� �X��Q���m�tr����C���-���enB��!5B(pU���
OvRm�>)$�̀�ŗ��=r�K68��-�^񷪀�t�̫�����ih���ӣ���u�g*��!�M�����A9��)�U����l�ZU�k�]�rm�7�c����y��6�SI�R0p�b�	t!�6��&���t�W�V�bi�y�]ڵ�Wצɯj�j�_��]/�{���&�퀞ˍ����7�#��΃�%#�_�ZRM���%�?It�r=4PS��y����`��[�A�g�ۻǦ��F	?�k�M��d<�r��ufS��0��Ve����ܩx�b�K1Ќ��!{I{83^(��g"E��{ЮT���Q8�NT'z���%BQ��K�����PY.���k�|\��V<�������z�@�����.=�c]��~"y�� �nm���i�7���;ǻd�������ݿ�L���5�X+�C��G��Ü� ��>Y.y��N�+M8������QzNؐ�@���hwCA<�	�]�}q��"[?R����^WY0�NA��U>��ܘ�s��@���q��&�_� ]Afb�se>�
��+����s�hs�ЏIP�$��;˵��Q�DLJ��g�}b��#џ/���!{�V�A���œ	��u3#���T̶wPǰ�hL�����:��G�#���ߧ8��3H(�@���jlV<����[
���+�	�F� �����b�8PH�c��-��8}��S��7ĕk�G�~���#��-av�㥐�_����r &3e5���C��C�k�'��7�:_�A;�χnӞY2!�B��٭
S���D,���Oj�ۚv��R;�5�E�o�z�7���ev�̊f����H!�$�X7ZN�S����9Ly����QK*-���FA����r%�/Z�u�,[����s0L�%��V}��r�s��c�Y�溵 ٩��f1R��:if���ſ8����k9�z�sam�G��zr�`%;Vz�U�T��ɢ�,zyl!�n)�A \���Cj6�BI�=��El�-a�� 
hF�v:i[�@�hZw�hC�/�����P~�)�]&��	@��ڢV�ө}{���C�*��C�{��Ć՛�U��~��l��zb�諂�7��&]1�)���p�'֢/������zBu�je2d+�7�*�u�c�E.ϖ�|{۱|Q��|��+dѶ��0?�:|+?L���ݛ��ִp	��}�˖�:XFr���e6:���i#klP�mA31Z���#�����),���75�z�{/!�!N������m�l��J�z�H��q<g��������S�W�;�����l.7�M|�*ϊ'.Q�P\�l���L�G%��SecB���/��ʃAQL����tMc�l�d��Sw�"�co^~����~ ^���E  �΢P�eTǦ�^ȓ�E�#x�|3��Ru
(�!��z�����
"��#s���<f5Ņ[���J������H�:�4���J5�}Q�"Xy]�x�_�:k���#�Y�?ǰ;������,p�V��n���伧�{��2�WOʵ��xNu�g�\� uk!�K�:�)n�-�0[u�`c�f�0ϛ��p��ݿƈ2Pp ����]�e����^��(��"t��E�� M�2l�����9�۸ׂW�Qz�ro0����*"���]�F�Q���nʹ�X>�(^���N�!���gn��3��/�c��n�	�y�h�a%B�
�r��Y��d{k�8D������7�_j���Oƺ�2�#Ih��K�:��J�ͼ�Dx�����.�b���n`�V��Ϲ�j�m���:5G��h��q�l1o���m�9�Z�ى+w�w��qţ�TZ}��C?��* tq)��S<��T1j�B��C.T�a�4�`�ʭ~�LU����S�T�v�;C���:�0C�eZ��d�J�9@�0�/V�	��a�(���S0�3��/N4������S&YG�C�yZ�e��(n(�Z��6iѼPc4���Tơ���G��� zj����R���ۿ�n�o�A��Z��Yp(�``�+���ܳ���Z���jH>LU!<���o�݈w��6�X��ǌ�,�o�m�]͂Y�����'
Klu?L���P,ϭb�� �:%9*�\�t��l����}��]D���}U�#ٟ��`�BP�&�Wi����밚$�M&��)��_��#3Z։��/��z��ئ�ۧ-��k-��V�΀����.6i�NR�*W�l隄���\HMȜ��ȗ�y
�_�+�;���i��A��i�Sf
�KT�Q�"V$w�ǭ�
����wv$���<�b� tM�6�2�y��av�rc#u�-���F߭�����{���vJ���N���;XR����ޘ���Y�v�PBc�ֳ�Z��'�>��m4��X��o"J�b7��N}6�6l��W�ە��iP*~���5���)���^�`nJ�><җ��x�P���W�.�6<��N��.H���.t��~̯�w��̄��ivG��餌�z�-6Nto�C�ݸ҆���J|4r���h��j��x秹=���U%��:�&�E0�%`�[7�ti���F�5���z|5 ǅ�C�x%��*��ꖉ�?H��]�fʢ^�S��������f�`�R�K��x>�M�F�zZ٥�uH���cW��J�M��u5Ǯ���c{��'J�<�@���S��y��N9:PQ�yT��=`��Ō���^S��s�����E)�QvI��F�+�U�ςX�G=�J0<RY���P��s�z�b,����{�{s�P׵ҟ|�;G�&�C��wdsW���ю�\�b�9a�2��Sʜ6��칷,DRx��atI��DG��9{�|tOD�������Z�G;֧ȿ������R��¡h'j,W�� 1�A"ث��S�\��S�_y0��J_I���Gk�4�R9?;yS�a��(EPv�1a�;�D����X$2;{�n}�b�������[|�ѝHќ�W�����^�m	���v��v��\���[I�Q������0�%l�~�r>�rK�Y@��w3)2�И�|_��#K�Ȯ8�g۱v|:��}���g "��ր/���ȩ����(2��5���+��%���.;��`�ޞ		�	s�z4S/��|d�?���5;	�G���v�-ڷ��]x�|��G�IRe�B(`�)\��o������V�k��@͈��E_�����L��G6�:A����UȌ�Gc����7u�)D���#�ח˙��?����J�u!: �
U!Qf�Z%���ϭQ�HWSM+�gWt^���yl{����'��l�Rގ)�F��1�@��x�)^p�W]0��\�4��@�F�_�j�ʡ��	&l�a���҉wa�bl�+�u�zx���mT�ﭦ�X-����w����Ń���1}i� L�Ц�ݲ�zJC�)�	�'�;F�$���ԃE%�ؠ*iT;k������|���H��:�3�����c�hr���`%���ˠz5_s5V܅�K(w�n���O�W�ń����
6��YR	���iZ<��ф�f���հcU�9����T�Ͷ$MX82�cn1��w��O�+���u��Ҥ*o&z��o�+�D�h�y��3%����֪�5Z�p
!���9�)N��XA��:V��5q�f{!@�x}��*i��>�Y��6r������A``�G׾f��`t����j)�Z@�@'�BL������no����C�ʺKk��h���`��/�Hm�pFKn���gB�t��jx.��;xi�]?s��H�m�h�����z�x��mɜȝ9��_�R�߾�����׫v��tS�,�,�lՁ��=��v�FS����p��l�����QdY�i�i"u�Ӹ3EeX>�ؿy�S��}\��}�:���Ȏ���E�م����ǚԊ���߆��j*�j�"2��.�ZTza i Ha�F���qeȚ0Z�����<Y� /��m����Z��U�H��(��4�	]�m�I�d+���^@	��nf���D��L����Q�4��C��k����7��v��wn�BC�s���8ƾ;ދ"X���&Ύ�L�1!��R�[pJ�����V9T�`-�ҟ喥▻������g��:`t��+��^�r�Cw&�	��<6���z�C�:��~�6գ6���-44:�3�N�4���PF�����#t�FA���
+?�S���V�!L�NJhM�k�B^?�y�w�=�T6�e�G���c"��y��������C<���j��X�?�?J}]�ZFI5�<-_z�`���������;P3��%�G�����.��*��RD��:`�:�a�1-���s�r��|�N������.>h�w��T��*�[�����:���JB�fq� E�O�#�Ht~��C먏K�A�V�:���;.���v�=l�[WG�`������Y�uL`S$3T�A�0�@`���V����0f��m���3�]���	�M�7�ОZ��RWsk
ϼ6'�л�r���pG�����r��}���J�&*���{�)���G#�֊ٲ�	_���V��ѫ�f�=��6�ϱQ�o����}=�<�*3�H�Z#0�P�/�6����o,��(�LO�$��7�C?+f��v{|���V�g���f��D�=6ǳ^U��뱼URXs�E�q�����}�#~I��������d ����9�������v��mA�TS:o��ܨ��YB
'���_�K���42�xz�8�ɱ�s�v.�G���q�F��S���-���Zb����m����g�K\D"�fa�jP"�yƚ�{ק8������bb1ʏ�׷)d�.XN�0�E��(Hx�M
�`�[4nX�+ �K�=��iY#�%�I*>��|̉�¢�U\�QUM�ͥ�**�I���&4�"�����#]�����Zq�"I���u���mU4�4l>��bv+Έ����oe�k�$��pu/mA�����Bǧ5�X����oU���~�]0�m�;�lCN�3+�M'!\B��c�$�\�_Z�F�E�-���?E�����\���P�_u�>n�#����ھ�De�f�1�b��qF�w*��:�")�h�k6��`��gF��dI�R٥��Y�`�N$��)EB������Y>G�r-048��N�o�F�&`5=�鵡������BG�_ �!���ƍal�tC͢�����2��)�כ͹W�g��L<��:��	a�Tj*\�f$Y����N{��7�閟���-���[�#֫`�6�|xA�F��k��s@KA���U� �L���mM�q�'-�/Fx��=[d
��� �}lA	����,����K�%�9;���1��gW�ˢ�M���ΐ(M����t7��w�M�C�q�K��s� ���a��RL.8�R޵�R�a�����q]O�f�Fȹ��$�<�ˮ��Lx@�,��A;��GN�G�?G.T=�����dR��|��`^֤�6�rR��d8�Qﵝ�1.�����0����Cqv�^D��_�q0��W_��51���36�]���¡��>�N�-��(��:���]		��!��ߜ]�o��!�N�}-���:5�(Ni9��+B���P�k�y4`r��f:<����
��Ga�eN�ah�v�YFv.���疓�Z'���s�hB�P�9!�R&j�'�	��k�1�c+�Oi��I�q��P{�]o	���H���'j��wܱ5s�*�`ʆ���롖
��%/���k��J�S:��N���$�R�kY�Ez��m�q8���0��@�A�04���D�̷.�7Q�9Z�i� �Lp���r�a:}L|��s"Ԉ��"H<]ak�a���Lψ��-Vf���Js�t�]��.�t_mJ�8�Um��},�$�Al��嚠�w"���.ٿ����4���h�[������Ja�X������Zt��K.4�'+*8�ھ���$��l��g��;%J*��"��S�n��U)���f�+>Ў�JKˆdy�N�	�xxI)C/A����Zܯ^lsG���~�=�א��K:���biW6�5��J���l���qK.Uk�P��c�d[3�(`���hl�:���M�s9�U�C��fJ�Ō��F	������OKQM}���NҖ��>��ywC���aI�&������r�r�����Y�� �B��w��s�G��g���	�V�)�ƴ�{���W=���v��b-��D��y�/�<˔��0
Z������_��̲�u�}��{�YD)Uӂb�+�ĝ��]�.�W�M���6�W�����/<�hر�Ľ��7]�^k{�D��ѭ�A���lGp55'JJ)��TZ�F"�$���W���#O)�LE0��I^�iP.�i:����Z�	ݲWע��vƣ�0�_�YI�� �-�UCFy��F{_��aD� �	�]� �=��,ϫ���lu�2?���Ȑ^����,��$��ʻDW�ɼ��R�ʗ@�s☟�'ӹ���E��ͺ���?�����Ѐ/L6.f�A�����@�%�o~;{;1v�)G��ZI����Լ���=8m6K�P�3���	G>�f�h�K��� #-"�دʜ����b�9�`��3vHP�ȍ%�?�߫Pa�hM����e3��}��Z�`#KC����Ոӫ���^�/���N~��"X�0:��Q�#���V?E��\�!0�����.	LdM���24" ^�D��D�}'Z,�L�f?��4��1�k��Z�4�r������pɤ���0���zRp����$��34+}�='#����*��? �=���`בm�m��:U����Ǻ	��4g�	����-��a�2lA�W���H��� �^
3V�)$����o�G��W��ԽP�5�{��4(S�TU�\F�.81����n�B����zz)&^0��:ADz�����*���Bf/���X����j��m��p}�B���JC�������.��Է'`�-�}h��Ν�䭰a�c셉�SP�em�{a��|�I&�¿߳pP������o�!��m�q�g��CXݩ�i';[�>�<�A�w�̂�gC��=��l���3��z:6#e�^��$�{4c�BK̮� ���;o޵��`t���W@j�����O�V[Ř�P��Wkv���S4�9:6�Q^��ׄ�1���4{��Q"�nQD�~��Q{�>}��_Թ�Ӱ���M�ne�KX��{ч%��F� [��@R�_�{m��0G�+s�zH9���;$ �<��Ň`CT3򣄲�QA�ɂ�3i�M��Mւ�Vϐ?D#�5SJ�p�O<�p;{�~C8�T��|�(Vf�vz�-;`.��܁^��1�B{���ԅ����Qȩ�%/8&`'�Ƕ�}G�#�{E��م\2�5�Q%6s�s�~O��S�=��D��1p�P�q�fAE\Z��	.����G0B��UW.�ޅ�n�<��w�i�__�<�7���.���g(��?0�X��r�}*r:�l���ZS�w������Y����%�Ft[V%JO��(� g)?���)��5���'���0��j!~rI�T�+ �]�t�g#2	[�Ty�P+NO��s��l)���$)aՖ`1G�����)�}�eՐ�J�AL�Ҫ3h%1���pf�y!G�jգ��<A�DE�'5BϦ����*@���3[j3F��3�=f���RW8-~��4sW�`���;�H.LMq�{6n��6N��詧v�����E��11C�*;�.cT�<�&u���E?�BE����0R��P��>[ǳƚp���}V����{+?W�!�h6n�mS�R�q�8��Ӄ�nY?5���(Wߪ"�|�?Ӷ�]_�B��O�jF�2�t2S��_�pH:z��D����.tL��l�g��o�j=L�!'�`�Ķ�Q����a�O�d��5ɞ�J⑎�U�3W�\���qa���.Qh��W2�I�i2�����hmT<�jt��p�SW��-m���9ς���_'�+O��E�����-��SџI�hB���Mnk�����mG�>�V<; ���_���Ȏ؆�-�/nw��4�޵�b-k�r�up�b[ȕ��O���U�t�k�n��(C;a��ג$UT�U������1.�ct�r_�K����
!��U�֐��
���#�)�CX/�<)��Њ�:��R��O!�IK�t�۰��y�SS��{�ك I�9�}�W�����d��DH������'��xG��m�����qX��rv�H����~ M��	���V���X�E5��3cЅ��q
Ƭ��L:V���O��I�����C�j�9c�����*Yż�I�<ϣ+4��#��x?�і�o�հ�ox�$����8�� @���
��{.7��x:�L9� �s�ԠF�]��½F'5�������]�����c�l��5˿�J2�r�1*�I��x$o1F�M��6)"��r��K��}��2 K;����xf��#j��H��`9��~' ,R�:�.�X݅���89�ʳ��?ؗ!L���:_b���ap�på�~��;�߮^��W'��ƹ����-O.�'J��bԓ$��h{��� \�������_^��$8枂:7��^"��Ax��8�8W������a�)����O����Mpمm�(�̜Yu��V�~?�e{{�ۭ�K�k$�wj���q��hq��92���#�3H����U�Z��!PhנлWv��}%����"2�"��B�b�wPp����z����j~����ҏD.=�l$��Ѽp�&�����.�G*��I�� �쒆��D +ya"*�k�����H}������+�HveQ���yyg�:�āo�tF��zJ����/���w9>���b8QKP����6mg�K�3��0�au�:��q��>��@5e�)�.wTZ T:`bRG]b��|�a�1[��A�x�c�'�������v{�y���㻗��Q�냒��'����,�-��8�*Sm���'՚�S`���OK<|�H�q���<�)Rq���؝r{�8_�כD�қ���(eB�A"������%l'�b��[x������3#(�m��1a؇�������"ue�_���I���X5eQ��XZ�$b?�� ���ɜ�5M���.M5�0;�5zOZ�'��ip���0��Y�h�����Ў_�}�aR<��j�mko�� � Z�0I2�-{��?��O�3G�8L0�d�eV��c2Hp�<c���x����}����y�g�9ߢ{Og�KE��{=�3)�2wTՆ��}
3�C ���?|9e\H�Rk��ꃾ����P	MC����v]�Bz��
i6
1SBÉ����*���5�� � pi2`wo�?��!��\��ֵ�>���mZ>,d K\����L�A3�R�Hz^!�M��+id3�]��3�v-{���;�J���w�b�|���|��*�5nb�>�rKڪ�U����p�XAcm����2j|�PZn��; <F#y����Pm��`�7��Y<uR�[�8�pk=�g��z%F��gCv�@1��Lw�Q�eۖn�z�	Կ�5IY���t_�D1��:�4��������kêUwvM�^��6L5���E&�i7d����m`\k�M�޸L(�n�򾇮f���Hx8��x8�Ma�	�K�I]����#[����e�}���
Ԕ^X�}�Sbm�ߑV��:��ؼ��a���0�ʣ�-��r_��fBDv!�C�~�T�1>y������ ��R�9����d,D�U�:��v�:lf5�y����ܓ��J�w2@^����m�S%�ĕ�����rK�N�09vtWW'�����;_TQ�I��u���]]����NΠ
~�_�XE��#�;����+"��X��{��w�B��H���t;>Xd��F?���tZ�����D�%����co �}_E�V���u�O*�L˝�Q�J��ߥGh6�V�F��=.�B�����XjN�����y~+�t������_�"�jixz��Pf�[����o�釽�v8R���Eu��bw��?rE�T �o�CHw�rK�gK��%#�2w�@ʒb��E/���g��bĉRy�ڄ� ��ҟ3�1��hR+NLd��L���\~��
P�/�	�#�����Sn��/ٻ���;OK���l�N{N����]�(���h�
~��Q���+���l��g�+^��<r~����P����[�e��t/ʘU9_�K��;�$�D�i#��Y0]����U��=�Ff4�0]�t'�g��JI��u��u^�0���#�1�̮��5|�S�PLy �P�@6˵װQ|x����f�"����#vT�UhHa=b7\n0A��F�y$o�%��B mɤ���#9ϻѾU���������>�eդ���+S��)z]-2EH�A�E##6^dˣs�j�t����@Y�lET_ܡ�td���f84���FF�d�?�K	�5�4Oe�ѷ8r��Lb����{�܂�%���U��4�ȝ���/xf����G����l.9%���~��"^���2�0�(�>4xι�_ڶeCT� ih,��ߍJP�N���r�HFofl!e���yc�+��w[��L���6�"-���q���E���N��k�"N�&��־Zd�YK����������W#㩲@kc�i�G�LX���h�o�w�$�eM�e�!R�9jϊ`��|׈���F�*�&9�>�� ��G�Q|�*?��=��	8�<�HDX�����b��ן�3��g�-/%�y���U�t8c���
E>�Bfl8Y�]`��!R��K��ﴝb)��x�D�Ef H�����
�M��ռ�
�E0�Ԯ�2y>�WK��y-�J�r��׻��r��O�1c �~sz���l�g��VGM$-QQ�\OD�8�  �����:U����'�/ιT1l�����)��8o|@.٩h���C�Dy�N� �6�OTO�}5�P�PR���Xwy�������99Ez��Ax"��BىI9Um��'5�!�����af(���D��{�*��2=�kr`�0E�Q)���E��z{3
��֤������n�Of�fMt��$��j�(�Z�����|`���Zʶ���Mqm)�$�Rg�(�;gk^Cb<c���smM�Q��S�̏��	�q��(�\��o�M�O0�Ț��jm�}���~�Q�����١L=];�Y��x'��/!o/[m����S����\�����m:�1�ؘ�U��P�U�b��Dp�h67�Xт�s��7�m5�의��Ģ��ƃ�,F��l�!knp��l���CM/�$l�&I��L�sPһ /��~����O�6�̾_�?"���BnD�hb�z�s�75y�b��]�����cT���Ek��~�m;����1C��XY��� mJ�N�
' ��+h"Ŭ���F�F�U�/���d[�ϒX�Y<��|�d��m=:8�l.��;w�c3Q*���_��1� �-6��D���ǁ[�~��#s�@)y�s�/�D��F�qr�537|�ȵ)>B�7Ou䬡���������mН�J�%�c�%^�M�#��ށi�?������)n6hi7���W]���##��$;C�L%i��b��m�Y�o��任��;<�@���#�O�L�z�\����zć�1�>���!蒂�+2���{��J��-;��}�~���DH��/N�g-�&%�4���U$^u|^g����Fz;�RP���"/�n�qp�ѡ�I��F��N����8���+T���}w�Ng�2"�� ��'�8R2�c�	~�&�F�HYd�[��P��beÕ�\ j�8O�M'䮥g��um�^Ϊ1a�:��	
���O��6�V~˄���F1��E�Q����H�b��,�N=|5���[¶C.���s�"����R�Д����!��/�mhb��a�=U «����E�E%@Z��<�Hrz����h_ڮ�'���d�$m���1�Qt+T��Usz����?OVΛu툕���Ꟶ�#LW�cI�+K0�c?�O�/�����
�a(������)�5-��T���
uk�փ>&-�1�
Xݯ4�z�6�mi�e������1�+�r��4 ���&�i�����ҌYkJ��il"e�R�x �o��O
F��%N�����l�9S�����ܪ������ɞ��$�`]���~Qb-��Z�v��Z��M��ieO���Q%�u�y�?��W �y����
� q
���CB�/�P��к'��UzDM׀��l}喂��x����<����:2���oT�\{�\��I��B�M�&=�W�,��4����@��y�����W*`�N��0�r�U�f��/��˸���w�=�3`���'������q[��\�Ȋ̪�x��,WIH��kn	��|�>$���6qu	��:m�P���->�`�E�hB:&!i@�k�A;M��s��wo��aC�� J���x�W���.�������GK��e1Ő��gWP����/���C���k`��ʐ�ۏ�)�ʩN���oM췒@��������Ã���ü�Y��m�2�/� h�j^۴��3܅_�7�\Lϫ�8R��w�\ӠT�Թ�p63ַ�r�����t��o�L���r�qH&�;[����h�J������4)�_�2�����+I$�Pe$�}��*1�k�<ʷ5j'�����/���a/i�rZ������ʦ�'������뮞��n$6��w� ��K��5�.lL�6pN|�@��Cp�N�R�Ҕr3�w36�yt�_@'I��Ԣ�^�w+	�&H�n#�:�ID���W-{���`��}1Y������=����N��6�?�Р���04��YUS��-zN;Aj��+���ͭ�p
B�%}����9�S���R�G���L��!���t��)�3IN,���8��Lj_�+�w͂H�5M�;�@��-<,�"�rٽ"w9C4�Ϧ�#�;D�̇���t�����pZP_�~L�#��;(-_b ��B:}�|��H���q�8�ʹ_,. �a�3@M��-}��k�6��Ȕʢ�,[���-h���9Dz�`�
����m�)�(s~�6�2Vo ����%�.uY��! ���d�5�C�<t>��$˧��g�el`���tD�fS�l{\���Wl~���?T{�;n�c7�Mwv�^�A�8�(���Z�~F3c��MHж�k��5傡�n�N�ӡ;{������|S���4F���b��+̗(�>
���%�L3���ڢ65M��F�d�t���rKl�4��L��w/��O�HH�	���ڏy_{P�MMFo���0]�_6���y��Ƃ�߸uߒ��#^���E�Z�=�k��$�5�`_A4e�2���/I��\	2(�GZr�KՇ��D@7�RKd�q��"�(���{:?%Q�_��G)���v�WO�b܂������TK/�(�k���2)Y��|$�?g /C�i� ��Ϸ�ߋ�(�a�{��2�;E7�U���<xQ��Տb�
0�;�G��J���n��C[�(�c5��Ƥf��[��` [�M�B����`A�ȼ߿�8��u*Ƀӗ �����3�Ж:!��Y�� �s�j�\-ۀ��m���;-��-��X��"n�����F�&F�6�׉6@g�L�n�Y�E��#�����WKEB�6�/w��ѝ�������E���� �� �1��&�b}��u:/"��k��2.���a���.
"+�?�^eƊ��W*�;e
y�^�>� qL /�*H�_Q����skP��᎘n���}7�q4C�;~�a�ceSK�Y4�s�S��a]��/��Z��^G"���p{��I������ϳ�o��I!5�&[IF]����z�%��Hi��tpx������p�G<n{��U��Ra
'�U�Q̃�Loɥ��9L�Zw�ٞ���c�x�nl�i�1["�S����~s�''#;^����L�����U{r�ݿ�i)1AN C�Q���P\�:��z�{E�y�K<�v�EGc$ST@�>�}=t��;��%u�48w�D�6?�l�;[���\o�������"Aw���r�]N��,ĢdW$h�U�g�$'P^��?���a��$�a�P�Ǵ����)�j�����B�J��Q\?W��#�I����@R~����8DD����oIИ�+�i5c� � '�]ɥ�V���Pu�(�?�!Ӝ8%��[�� �C�a�󬮒�{���nP��_���L�V�=�1��]a=ߨ���
�wx������m1/����}tTaث�Vl�� ��'�w�液?�5�"D|�K'���d�� ���@ bk�L"K4n<t
4-[�:���V-�BF��Ķ`#N����}�8�e��I��
'3Cƹ�lr�ʺ�s��u��Y%u�[�8,�(�����%�Dt�8l�I�p՚[�d@CDa/���vܽ�na$�O-���J�\ܫO�a��֌�]&�+�E;��A?�I჋
�k����Ǽpԑ{7ޥj:���oqj� J5K]�a�yj�n��X��,'��� ?ς�����]�hԽ�5��ԡ�,��bT�^<˚���t~΄�Y�N�%K�I�n�ᵆ4�����k,-I������ؗ�M|��[/|^N�3�����Z"���</(���Mz�fG^��=X�����DN��t�������e�	��Z5�Fpt=I9V�Ar=[���,A0��b�iP��D�.z�@���?��קD ���h��)��2}�/% {-�N�NS��Ѡ���ju5�m��~�W�[L���^H�/2�������	��S߶�w�\�#�G�`��[S�u��ǎe�	BNisf�)͕\��#�X �}2�RVle��N�T�H��"���Wʎ��g�a�y�Ƕ����&��e ��m�&��$�Lk:�<-�����"9�S�);�a>��D�`���4V-��kU��]֡E؈R����R��Y:���.yD����M�7Gؽ��r:b�%�*D�.�1���|��u|���M0�3S��Ӎ�^�q��[�͵�䣮BT=ȳq-�ZV��_�^w�Va<d�M����zNGTj�>���셜9��f��4�-ը 6-���[f�Ό��3<�Y*�o�}�˾��Ir��mԤ��D&.c�< -g�ն�!��S���֭��E#7�Ps��"�g����_��sT�e �W��O�Ӯ�+ n�z(A�}S��zj�Xb��J�7[F����NVE�;|r�b5����?�$�J�(M�cp�ഊnlM@�����G���(O5o?�\E�Ò�jP��zT��Դ9�w%a5�D9�$J��9�a��KCqa�iŦ�F���1��g��L�����<�4Q�],�N��r�=��:�W��S��v�lzt6�<��3���3�� �� X'����3[�ں��/h��_���/������UG���o�ү�ۆ��S[�V�H�u,�ʞr�Sʣ82�"Y�C3j�:+5�Aż�/�8�����{!\(�{.3f!YA�T�o������W�
ۆ��W��)P���XP�'<�U����ɗO�7i��*��7�4�$���!6P�[7b�;���d�E�"�t��蟱}y@rn6�s�q�Z�0���\\r�.�|*�Uf�X K�"�I�}�N+IYd�<}�P��A�a���_vi\�a�,�G�`L0���!�����U���wZ��2������>�W;Q{�5$U/�F����?�q�G�z��ĝV��g��L&��El�6��3�[�I�>�i��s���h�a�9���2�C��(��}e-ƺ�Ԟ�cc(�����MA`S���OӬ~V�_8fv�@��%���ŋ1F<MUh�Q"+ż���^�OR�˲ $<#�c~����{�#؎��bk��3�|�����zo�	GEqe��f胡V�\�o�c��o|t����n�7�����\+L�lrͤ��*�]�sM6|��X�����]'�Y�����12������q����D�l�x1�õ|�;/ ����vR��b�`��EI;I,U�+Ԓ���Ο'|��g�Dr
��*�7��ǵ�pM�x��*�!2MO��"n%�~��L}@�U�x=�|�yi���!�4��!�bYaO�X(���O�G�����䯍�d�EL>?E��]( �PS<�y��$6m� �lo�M({��v3