XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T��`L-��8�2�3H4>`6�3$W���vw�F4���E��Gu��~ݞ��_�IM��>����� �,��1���jgp5'�A�Z1C�'p��������M�������|�kH�-'Kn|C$���1r,�翕��=&���خr�h1�! 3Z�M�ݺiV�c�'}��AW=���4�ܥ�:%��4���(��`G��J>t=�	��/h��6*����C$�vz�"���<�}foWR� c���������nB���z8���_1�?���1�������)>i�Xk��� �Ѻ�'|����Ɠl�9~�E��Ud"�L	��wH{�N�u���1���\;�L �D}_���)�<u��^��X�Js���P�KN;�]	���G�Q���םd�dPs�����JB�]�j���
��j�k�(�L�!"�F��?�W���\O�(%�+kg���������,�.��2)��:�s=�\ީ�	���G��u(R.O໌����?q]�4�A�UwSd�HwVO[C��I���.���3��g��l�:��kx�w~k�������F�XrG-���4�	F�?�:&��o��
��u�\�N�vx�,߉�;����ke���82#꼽��@u}E���*� @��a$Ʈl!2�J� �?��|*tTu/�t�3�?��D$N;�q;Ӭ����Ԫ�ѐH`���]~��uJP[��8޷�;�<�rȗ)h.�a4 3��;��"�M��hj�cp�2F[��~�![a�XlxVHYEB     400     1d0򓏌)���e?�&<?���\������|�v�M��g��p{�.��������]������V(H� ga�E:�ˋ���e�u�v���63�{H��R�ߛ��]��F+� �� �G���^a�[�5��}VA==����b�膉�S���M��eL������ش��RT�J��`�>k�v�V#�0x�Lr�b�S�&>�e@���V��ߓ�-Ĉ��)*�EGZ�I]rd@�n@t1�$A�ʒB|�����d�s�>gD�����T&���Oə�ؑ�B���j�lnz��ӗ-(��騮��c)J�e���jDξ0{���$p������E��	����w��9�&7����hg�E��,�ֿ)�e�-�fE?1���Vl��a^�h��EN]��!��~�\EhH�7����Ezk7k�]+"���������t���j`XlxVHYEB     400     170]|��a�&�Do���?�jG�Ӕ��$��j��5��{�h'ް�56�qVۉ ǃ{-
��i�dhy!o�-�b�'��>f��!�p���d�@3i���BNܣ{T(s`��އ����o7fׇ�����na��<�Y�(P{ӥ��	e�P�j�C��)��_爈�,D-~ʗ;�+Xg["�ձ�������/���O��G'�_�1��ø�ћ��(��:Q����Z��1��w{�?'�����1y�=j�G"�4[��@�_�ژ�4la�l��XI����:{*I�S�q���Õ(��򚡎�HJ��� `�#��û?=��f����C�٢|� '{k�U�T-������XlxVHYEB     400     120�=A�6�u���Xp���G�X���m-��Wϖ �����w�F�J�ޏ���J��wϑ�M^��_֋E�\���������d*����n�8���r#��΅��3@&,�a^Ư�ͭ=�5M�e��ڑ'��,i./�^�A����t��Nm��;�;����yC��#�O�m����Hy�'����ŤJ��<S�i����ջ̉�w[sP���������?�@sv����e���>��f��O����h!��gk,+�1�R��q��LK��Gw��!�X[XlxVHYEB     400     170���-\>n���veXsd�U�qo��AD㞵{&��C��zD��)84b����[*����%��#j�qp�����{�{�`���A@����H%��q�H�cG��\(`��b�b�ΫM��$>�ǔ:Jw���ޠC�LSr6���a�ԁJ��W��?P��~�b���)��C&�T� ���.��qPKgQL._��$�Kq���y�F@���{�8���w��9ȑ�l�3�3��h�=O?3@�Gl���*������Jh4Տ��L1F�n)8�!��Q_՜l��RCYN@���C��&���h��?!�W���+Β�ܭ:��b�횥���-F]�́3����e�4u�'����)�V:W�5���XlxVHYEB     400     170��j��agƣd�u��{�ËM��{h
�<'J&��C�}c07� A���Z������%�LOTo:)��e�c�E<%`�֟�˾��۝��P����������̏��x/�;!y�)�o�ɫ�T)�Gj|b�c���s"h����$#<�'"��0��k��,�24������Y	y�3{
�Q�O`h�TnȰ��mC�U��d��i��-19jax�K�S|6�(E�*q�y�HNN���J}�F�B��@�:���С;~���lK�F�]�D�*�(��v���c��ۃFc�%�EU��WO_�����O��d�z�ũ,��ա��0m���}��*4'�R^�a`���¤�'`�Y�hY���XlxVHYEB     400     140a9��<�;�
E��2�i��\�r�dO��ݸ�<��$9�|T����'C"b�uE��T��Ǐ<vM��}�!7�(�x���ޡ�ͦKXŏ�	a��N��٫`=��.���c��Vߋ��ڦ˝���/�^`��D�@j����z�&eJP�e�����Q8��٩����@tE~��V��B9�!%v�U Pg0��]?�tp�u7g3��P�`M�e�~�/� =�����H8�@�1l$
p��S���E�w!�ݐсT��S����Y%�.���:Q'&�� >�}��{36n+���?�ɧ�m��-��h-XlxVHYEB     400     100�͗"l&xnqL~k^�?�,hq���d���v���JYzs�mp<P������3rἐ���2�׀9�L�|Ue�t��;��K5@e l���"����y4��J���~\)1X�����l�乾�A,pʹ;s��|o�E4n��ʳT㔙���S��u+��)U/440G�Z�6��ڷ�J�׉��++)��߇=k`���P�� ��\7�=�/?z�f����������^�>ض_�w. �L*���,�XlxVHYEB     400     170ּ�̢و�Nlld�ǯΧ:і?�M�<�a�⿌rh��!?�,Ǜ�+�Y)��4K$e��x���2pR_�6��!�d*��짷�&��d;�b����4������l�I��.���]v\Ci������mg��NC���
�oC��`F�A �p�of1�t�����;�X }�=x�/|c�wg 2e�l?�N��uF�k<���؋��R�t����+/g�wxU��>-'�t5Gu5C/�l.%dF���ɊT���-,d�P�j�%��m�1j�Ӻ+�w��I0�8Ǟ�tyN/�������W�e��p��h�U�Ԍ��&IEP�z���;?a4�t�d�6��s0�r�?�����z�]XlxVHYEB     400     1b0�8��[��^׍D���.�kg\�[8�;ς�;��W�sX���^֝��q0�ϋ�Q�ڑ�����<V���'������3c���́�&d��5��ż+�鲗e.���ͷm^�Z�9�Z�3�����T�s��>��j�*gF�|6J���m~�y�Ȏ�"氳J���;ڥ�V��n	���������z�~M��&[������k�T\�>��+	��Mh�wX$2��es��NOg��R�	T��s��=e)R''p�ܦbP�W�����2�R��+A��P��B��R6�
�:=��qufՑ,m��{S��m���ŹM3ԛ��i�~���2�e/<�@�i��n�/q�r�>p"9~�걛�!ĢR��{����hx�X������wꚑ4�j� 1��IhQ%|a}j��:ڎ��\��ݭ��ȸv<<o��XlxVHYEB     400     160�M�?�ǲ%��߀_�!^z�A��D��7Dһ{�Đc�]�E��Jh#�����੎��+LS��u��z2����ebU���]}$�TH(��?'�o�G��9��<�r�'E4���mAL�{�z\3'~R([�,��y��,�T(a��{�ѱT���aW�D�'ԟ74���:��4&�_�\��߭���ZX~���lS�������,;�s8���]����'�ҀV����.���w��ES�/^q���4�T8�����9'�PR{���B������}P%���B8�*�����@�Btqp��<F.���m�Y�Xc$�;l*��&�b(@��x�5w;S$����:�IA�XlxVHYEB     400     1d0id-�Q 6���18!ñ���k���>[�^'pgXW`��(M�H>��1��߫����ѵ�gI�7�F��%�J�����}�R�S/H��㈮"#�U�d{<$0��ks:�.����L��"t�E��H��<��D�Q-���e����������@!��
�Vx������o�o�O_�T^=�~�E�H���ɡr��K]��V�B1��ܟ�?^x��AbU��(f�h�-�B:��
�ڷ[
��$�qPP�N�3xhp�U� ^ԟC�k�lE�RT��AL\��WK�(._��e��)K�n{E����Yk2jfv����NQg��\Ǌо0����dӇ-ᑽ�f��V��_�g{�h.��� �|A��R�jܥ�Y�谼�t�e��2�x�Q)}�%�3U��fI�7��_d	��5�[����#^��ޜ�|@��8�G3���`��e�&��P!���^XlxVHYEB     400     170\k�k�-�e�sr�N}�4��U���qʧ7�K-v�_����h��{f>��iK���H�Y���eED��̩/	AWT;s��EyF�Uɷy5�v����dhj�#�eŝb}�a���zx�v�7s���d�-���ocÏ�Z.G�.��ܨ�eP��&����&2�U�p2v楌����������	��&�lk�ͼ�8����sI@yM4���7��M��*�������퓿^:.$�U�$=�'�M�Tp"lC���HV(�;u`����
�ŔQ�fS� �tH���9䃁�J����>��Sϸ �q�,�֟(�?���u���u(��$�	�I�]��YЁ�=G���XlxVHYEB     400     160l5q0��m!'2��u;����$��Ic�,H\�P3��+n(���]��������m?"����;�����b7rf�� ����n��"�Ok(k�'��⭿�f.�5��FBW�6hʊMKT�K���c �'���9���ae�á�!�v��k��lsR�S���!����<��[�����	�T��6�[�`��O�U"q�KR�t�°hƟ|�"�VMp��m7.(��5�/��}�)����H,��zb�%��72q,h�I�	m���0�Dy `c9{8L��q��܊���u��W��dW�6�����-��5�����_ȣ��s�b�v5������Ȱ�%B-���jRXlxVHYEB     400     180$�6��w`��Ϝ}�^�xU�mܕ�cIȵQY{p����SmjO�uC��u]���RsB��O��`OI�"c�.^�	Z�K̑��/`1�IN������?ɘvU=���l��W���v¢�0pί)b��3�g.��¦v��y7�r.��J#A"@���������;,?��5�9�Fe�ZXz�sW=���x�I�s/��+�8c���u���C�\��}�������8�if��k��;���t��E�9�r$\���L&�HP�:M:�#皭co����#��p�`�c� ���<SP�#W�`���	��֜ؔ�����L#xM%H�}�6w���V^�<8�_ 	f�ʰ��E��,`$e\�]�����s '�NP�(
u���XlxVHYEB     400     130��<j%n�G����1jQu8������� ��*8v�.�,���}�W�8�k���ʛѥ������n�;sI�^s��7�p;�-����쁞�������l���I��f�F�5��h�F�@s�,�æ��3?+�f�eQՍ[��4[�ұ|d�����A,^f�VB�� ���2�$BLK�*�+U/?/��ߒtPU�М���" �K9Ο��(_s��j�7�i����W�;&��'���$b�=m�$);����cUk9��nԞz�l*�:S�_�J{�����g��Q�ȼX���XlxVHYEB     400     160�:&��}�	���_�@ NFN,�0_J�Э�+WdG��*���öי�	2� ��v�
jf+�#�o8�����8\�{���U���kb���4'0F�,�J&��J�W�v�i������sL�lI/���5�m��l�x(���a�������/��ߍ�I�4�;��� ���?�<�+6�Y�f>]P�i����*Ꟛ
i�L]\�;ܥ�-�H��ߨ���=��gώ`�W*���۔�6@�I��!��\�@���}��7}�*ezﯿ󁣢�	d����h���Ch)ݖ��cN�j� ��ۂe��7��n���W'��i�kT�F'lwޝ�r�+�#E>�XlxVHYEB     287     130<����vi*�۪6s�2�pN��u�Q	���W��'YH߳��"�.��?C��A ��qc��|�C����������M�;�PMb��J�*�Rr���H �-��5��oBH���h��)B�Э�l�j{���5�)��(�.�u�#v�u��]��"­�9z�q��o���o�cm�*�k�1pH�h$������~bϾ0D���Qx�F@��{/Xk�F�V����$ ��������0�e�#�Q��Y2[GF�|��Lc�g"����,�m�Y�7;�\�`�����o#����