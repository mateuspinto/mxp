XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`-)�x�:$b|Q B�����K�t�vh�(����z�(5p8�		����)�N��C�+[�I�_2�d�@��wp�<0+{h7C�����q9.6��I�|�MB5��[�L\�a�o.*s��6 ��|��	86jj3)�ȆE�-��_�/�p���ߜ�7Jc�z�/�Fj�N'�!�Va+e�F�L;hQ�oN���B �t�����jj�B��/3KͿ�@��nv�.n��GG��}O�����o���#��=����A�U���8����>�S$���0��,㪇M#�cw�	J����^�bqM�wA���D^�F��[ǪG7�%J�S��X�A`�t�L,��VAfp+ǸΞK:y�1.�W��Icfؔ���6�KT�F���D��l]�O�u+f��z����jמ�S��jw��ϙ�,:�<����ލ�8�j����<V���[��%h�އ��;9a5`R� ��	��d^�p�N��q�i9f�l�+�?bT���`�o���2y�������#2����`�����s���R��c�w<�xpf=6fA��)����Eŵ�����l9��2��߸�Gq�㰭,���Y1� s��p�Q����� �w	X\�|��vhxf�P�����u��.C��°�HG�S��6<�"u�,!�y$��j&�(H͑�����(�V�U���#�!.�7ۋ��%&�fX>������~.'m��=���`��˟�b��%�:i@Ha��Y�1��J�vz�+���
��'-I9"�(sn0&�XlxVHYEB     400     1b0W>5���.K��b��e�k/Te�#�'3o�E�N�gg��1�:�p�sm'}�e1]��r/��X�^K�H����$#"�Ї)^с� ��}g���J�DB�@{��ᒬE�����n9��$�����Z����Q�w��"y�bs�Z���0�B{�R&ޛ��̈́p@t`ԏ��������a J�)$��׀=bF�iH��Gh�x!��ЙeC�1��o�����"0;+ܒ���=+*��+�S�}����C����J��9ɠkA�����w3�>����6[��:gv�?���vXaR%�䟊j�9vW�!"��
��<밓�{���*�� Ƭ��&�-���57�8�m��/���b��f;�[Ӆ���\�?�`ܣ1�����s�u(��ɭU�:^�C�<�m��T���=�,V�o9U˸XlxVHYEB     400     1b0��>��㰛͈+���8���'������d'��e����ٴ������6����4�fӔ�'	�8?K�ZnU0�#C��p���#|�uT���ۮ6����U���&'G"���a�c��足O� FU;5?l��9y����u�,��݅>��rw y�������/�U��FiДF�LQFgk0W0@�s���P)�]�����!r~Y���������T�L��/�_;��G����{���?7n��U��'&)ϙ(�&+4��"v&#e�~Ox�v,�����D��x&�X��=@W��(a�F�8��d��bj)�t�}�X�Y�Z޺ b�5�De���	�B�ȁ���sRB�M�-��i{gz
[��_b�\^�F�NAEJ���[�+��dtpd�
;�ϗ�:�6���Ҕ�XlxVHYEB     400     130��#�k��t��z������$�b���nޘ��w�O�U6�%�[W��������ؾ����|��O]|=Afu*%B9�t
q���7�W�$xm� �<�W��+���xX�A�>e�P��a޲�S$��YK���f���"�V���=����ҩ&���!)�POd�և<�]i�X�F��	6�e�9�r:a(gRw�l	�� ���ɋ?���>�Pc(4��|Y�J2�j\�p��ǂ����6v�(�ie{�u����r좯�I��r/��w�`Y��#R�dFo����ۉXlxVHYEB     400     190�e%%�Y�(cSD�}�N?�g�ʬ/��hB�d��R?��H�/���y�KԗX����g���f�I������+��{#�371e;�r6c�<e��1l���G�-�C�`D���q#��V�S1�����:�����4]k~�
[�{����f2)4�+�,0���v�@��	�R�>ô�W;H�~��EM���3��H���t���T��^�*�7U资*�3�1�:fPr[�f����M�m�Q���ҁ>�@f�A����H��@�s�"�l̹�ʤ�����ȵ����7>�����0���^��ƽ\��:�T�>/!��@@�F�J(Sn����;���힜� ���Qb�Ib��T7��S���d9r 2��C�^��h
�%֘��XlxVHYEB     400     160���bթ��r��]�3��ӄ�'A:5U����V^�w=�[����	�@7HvSV1}�ذ�'��~9M謎�0ve]�.>��u�C�>��]���恽p�w�TL|���`,�"CDĔ�^�iрSld���35c���N|nw1�4�ʘk�k`'z�rL{1	3��S��:�T� TDG�xff=5����d���9z��z��
<��$)m��˼A���t/'SP�����+R_D�Dʼ���}�q�/���u���5�}>���n7B��*�ǫ�
�H�)����	�;?/�ۃU#��!8F);��p�ۣx�u42��u�N��3�:tZ�넑�GO��#�@XlxVHYEB     400     1b0N	v�0W�s���)�j}LC<�F�<n-Q�ÂB�x�t2:�bfln�![~ Бds�h��O5�嘖�͚��Xѥ�:�ǳ���;���Wb2 _�������q��"����A�Q���#�q.�F���i<�� �`ʿ$����3�%���^����=A���͈X"� ����y@	lpFV�P��p8Y%�Jdf��Ԟ�.S����/�����Mr�[��֒?�F[i�Ԙ�.��\��F�VU$l�P�B �4kV��N�/���(N�q�3����M��o^����n�u@d� Nq_Myn����z�]�a�e�YM %Q&	��q�\&_�S1[��*�?�c��bn=���3���p���H^m+]�S��-�[L���qw>4��[��zu��*��'OsiN,8f�(��XlxVHYEB     400     160$!�X��7�����:جT�	�}�9�g���A�1�	�=�(;�N��^�p��,[;��f���lBYg������t�m��Li�mJd 	é��R�DAet+f��~kɢ+�LM;h �&{�a.��qm�6�)GU2�����*��[���y;�ŃJL�rE�H�lh�|���l�(����kpP���_ߏĭO$�'.����]Q3�@�YD�u�dT�O�u�h��J&�p�x�0�
�vD¼��T�Y�1D����O���Ft�G-tЧ�����>=���Bf^�z��{�)$�Rչ3[瑮S�
s/��ת��į|Z2�_���meu`��?�e6�XlxVHYEB     400     120�
 7�ޔ������ 0�@Z�������܌7w�'�i̅d�\���rM���yJw���ibZ��$z3,!���r���2}(��r�
�`%�d����W����,����x���9dw�k1�M�z���œ��Xm" >����5J@�Z�J��]L�F�+�f��ñ>�b����D
�MIn'�����.��&lb����qh�/�����ޡ!;�G�N9�g�R<æL_/=d�!�����Ǯ���.��d���PA��.7�"��)XlxVHYEB     400     190K"�"p��WRI��G�є�M>~I?�^;eي��J��:�k� ��u�C6��8�� /V�_���u3��O�B������1��G��(x��85��J<���YB�Ld�j::0�9+�s|,���^�I�h�%�M�+�j�=6����v���(�?�����M��X���WY�L)�7�݄�Hat�/N��i��o����yߗ��7�_���������
E��Z�Э��J@�F5X�*���:�4DL�CC��Gf���W"�)� Iե�G��8vy���۞��G��;��Ҩrɕ�kw�4��+�`�2�J!=6;i���T�SP�T�k��^�#c-��/��'h:���Ϙ���uz��	�Ò1܃�F�ʕ��W��<�XlxVHYEB     400     140[�Z�n"z���et��o�^N�8
���|�Q��1|���H��������������W�{{1�,Y�4�2^x�G�i��58i02B���3�/%1��
}d'�n^e;��ULw��4�����r1�NًF�/��9L���������F��z�F�v�Q����sI�c�}��Dp�	���7Ќ���(X��tM��i�U�41G2�����N�J��|CH��a�n�ٚ6s��������m��[=>��ڤ����Bħ�jY��4�t��#n�zu53]�#4��e"��Ju��%Di8�Gz8�Zs�ªBXlxVHYEB     400     160��=U:�J���B\�ґ	WR�;���7A����5�_�����@[>	;�]3�!y�4c��]
|��;Ke�iLfgg��r�d�����Kt�N���Ç(#���n�-�^���&���1�0��� � `���ݳ\g)���?[9R�p)N���������X)i������U��7�m��?X�Gqv�'MMh,� �n$��)��wǦ�rl^{!�g�g�e�uM�:��މ���c���v'l���ƅ��>dO����lʊ���]�+<b-<_]�K���q57� Ǹ�I qx��~��/jmH���QM@,WS��k�G/��ٽ����![s,�p�XlxVHYEB     21a     100�ny�e!���(Q`ǌ�{#�G(��$18�ΑnI��&8���~���,oC�2���A��7���'�pK7��I�ްF����/�5��|l}�]YaʉaJ:���۵ �4�u��>�d��n5$.?2*�;֭4ң��+���``��/�,���pX#ի6���Lj>Lb�>!k��x� ��U��c�i�Lj��0�߽ĸ�ZF�l({���>|����D��Ko5��q�Ud� ��:[E�w\Eb��7�}