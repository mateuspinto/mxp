��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� vU���O} *�(Ӛd�ڔ*?�x���*�m(�e�Xה*�Y��3�z��J���;��铥pV��8��,< �J簒.����ÌX{�����=(
�`t�W�BilmV�n���m�J����v���/�%]�I�Wf�e�	��)ZF����c	ؐR�)J#�e���z$Fɷ>䡺�Od��)��	cy�"^�b>�0c����z�l@�|�Gl�3��� =�HQ����+:2�}����@u�!��E����Ę�A`~�$빰��a
����P-��Oe�w3]�`T�B���v5�#��4"/|��cXiĿ��!�el�,��|=.��%
��6=���.�4`ҮѬ^B��gV}nd�+���e���MG��*�
y���3�ֻ�\��&:�����˫�1�E�q[��T��60q���^7����kwV8���q���H�9�T��w��d���vyt�R���1�;QULG�ZΜw����懵g3|�Q���@�_����%�v�
��;8�h��~��6�rCI�2-ӽ�˫�N�3�(����Yv�8gShc�؀Ư.?���	Lӣ��
�2��п�?��$��� ��5���[~8M�H���ެ��60=Gf�)��c�
I���}h�5S�D,�a�y��h?K�&;fXµj#Њ �y��t��6+EO����,���D��t�Y,Xg�ȁ"���`�|��+�u6�&.�;򭩲
44���%�c�����l�`��,&`�#=H��8f7��w�N(�N{z`�L�I�Ƚ><�<b[ke0\���cp�;�wt�GR}�����}��>%�w����Ҵ��f�mM���z�Z��v�X���8gW;:a�3�Σ-�ݮ��$�R�|ڎ5�=JX���>q0�'�!N/>a�т,ORnࣁ��,��$*�@a�2Tz���N�O��3qj�t6�j}PB�6cd�|[#�c��Xh>�c�޼����(#��2� �ӊhyc@����v|j��"�I޼�aP�I(��.a�m8jn�Z+�؀}r�/`�b6�i�l�Z���	d�]j�A�s�� �(7ı���~�0����C���q{[�=���HO�Y����a�I`Us�u.-͐U"f�P@����`�9U���Q,,|'"�?i}���HLT$�X�n�[u�U�BJ�>�P>�+>J������ԑ�N���?�2�����O���MT��]����uf��kQ�p��dY��Q�r��D�F���)G�W\DkG�G����vuB�U��OB=�ޙ���s��S�cu��Ҥ�\�Y���ء��:K�K?�������A�L<0]ыL[Z�\��/��l��I���v����0-*�4���� 3'Y-�,->�H�Ż}\}������E��BDR���{�#g��ڸ���+�4L<:�f�U�� ���9����VI	u�H��`��Fa�Ri�t�<%IAr������2��L��ގ)�}"O��ߋE���D�b/��{�߶l�:��(�m�������^�Xf���LAX���bC�T�K҈�!�gֲ%+%)�XV�s-�p9�hfGk(g��j��X�pd1�����:�������tʑ�)�d�a-db�	q��
�7��%�]�@hˍ3K��V�]̗<�l�Do�ǂ��Rn��Ϝn���*Es�_��_�	Z�	׷�
`���E��~�"��y�7���`C ��y|��J�'�.�T��tb�=�X�s���m�z��L���tY�Z׵@_��{�n�av��k�c��vе�yLx"�#�Z�ob�َ��6čP��u�ux�r���'b��c�YwL��8O�T���������ʕ(�M�R�l&��p-���.�|�E�Ͱ/�Klq��Qa��De�yA���PmE���u�7�q.��2�ݷ�T'C��<��� /��U�#|1����fí(m�At[�l�������/@MO��>wZ-�o9�F�rON�q�]B �d�AO$��G9޼�k<w��Y�+��j<�x��#NU�~��d���p�%5ʗ�3��u�n�=*��U)��I���7*k���G��9)�
���W�R�j���[��?χ��a��:�ʢ]�~���`�8N�L�����%�w�Z3E�F��Ix��Y`�l)�� �ND��d� 7(���s���4ЪGJ������ /�4 �ʾ������*�R>d���k�g݃�1���������M�Ռm��'�VL-���i��=	� p\EnX����C��Z*�;I�DI�^j:~�:M�Θt�zWcL4߽���>PM��rpf���rRQ�Z��\����n�Z׉,��({����0�&3�z����oF���Q�7���F��V�B2���[g�n���T1}v~8��KD�Y�-�zE*\�d����z|A��:ھ@yO��-	�<1*]o���Yߨ��l�-;k~�I5Ej���q�k��._�fCm�z�����P�
���e`�%��W��Cl�	��l���"Wx�����O�K$�B�$P�t_�!k���bB�o ӕ���x�R4G��_8~����\kx�a�(������7'5��R�b���I�!���t{��s�j��4��p��-?�2�?�-r���$Ҽ+Ĥ��9¬�s��/̢k���߼�tHW-<��u��`1of�k��Hm���<�$��.�!#��ӊ���Pi��׋�̃�][���0�װtY�"Nx��nW��a�P;+]ki���6�
�W�~ ��ɔ�Aj�Gy/_��/�]�s�qI����75��ZBcW[[�y����,�ZM��=N�.��4��/q�M�LD��VM���ҕ�b�h
�t��F���V3i&��$�o��~oEd���+L��쎓k=9(I��r"��d�����J�;�F��	��D�z��J��*"��2#L-o�NDX�efrX��6{b@[�}(��-���D�o|�����