`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
nVANgwUqfq72w+NRRS3XRetV3tAoXgn8BqgVCj4oByJNodeu88jXFDcCJTgc/gk8YgPqdOzw4MKk
AEsjvlgvrX5TaBZUQcklmRYtwbmYIgPR6DTecNeN9/1yvv7hFdkM9UkMdTN8CZrc4Oi8aJGc9xwN
T6EWrCKvD1siRhVHsNZEmGi2vZ4VT3n1AVpKDNomOkD6ulcF7Hh/69VQk9lTZQ0Ye7K3WGXusZvB
RdRmlsSKlU0WabAQr8t/KLn99OOOnKDp3hahAsVhgIIMlzw4NA7e7N+6fCamcdWVgvtUL4E9DvkV
75MIkhJcxgS6ouUeuxOVO5Y1v09lDFG8CkXZHA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="XdeGOyPRImzPxgqxoOO8rVLZwUCNmAjeBTrTo7FOftE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
nd5/TrGCIRrMkhVa3fGd+H0LgNES3Ru+3J1vTbqizVL4+FkYmkHwhgWUoMa3THSaxg7Zza37fOTz
fIfUkS9m6teyF5U2qTJTXxM1/KbRq2iBT9Vc6CutewpE7jqh16ZZWVcliTy3ZPw3/7/GFgrs7yCo
rUeJgIKWVMvlUzDakUpeFyEcMqy5FAVuMR4Xn9I4meBORJUT9bahLl9upaencKbAHR3inIsk+sWa
OPLsr5XSZLmvbp1hCfQ9qGfZb0BMymbY+q1akIGjJ3juSHbb7hWTfIPQUMswtMzv8B+IduSoaKte
wC+LMm6C89KPfxrNCkzy0BpyA5xMsPfAzb20CiyIERwva/mr94Sejx8BjLLD5e04sBq2s0RnBuah
JVDvsgJDI55DR0D0LEGZZsdjcwfmVN4vlMusXG9RK8krskrejwQ8JTbdeEm5RHDCDBNUJSrakMgm
VUo7QOYh4cWIMfZ7OTFq/KosZZNPDpp4/qZInHYq+A7bXN4VSiFFNkO+OpOYfTBT3zI9+KVzpJxV
aOdbbRyjfkPQ7FU3v8pxBX2PYZu5t40ucEbB5uot2t2AsPCy2uahfNC13GG1q/GA4qNKG3ztNtFU
b7v+N95W9YI+urQ4J2k9i0kLZSpV/pDZma8NcmPoZlwPkNL7uodoEVUQnS9qkwIOiFDFLf0NCdua
pf8WX1W4oqY95BXVoemRZAkz+nXbwxpJy/vlc08W9CAUNmoFf51szHtzC+aBWvMteC/T/Rf6sqDG
AiJQ0BujUKF+muJ9NYDI+hWcjDw3izTjIJslRwCNW/HZklWrUdEa9k53Kq4/E6sY5j2TJ9B5TRzN
2qFm9v7x0T/JxNP3csyQ6ec80iPWaB6HMCMSxVMaXRYyaRAgGlYPBjNnRafW9L/9GCzqs59sfNw9
SUO0U6ZZykxPQMC8x4kLzAVLIfcU6lfpbOVe5b0JGgXMxGYMTLNB59WtpWtK3tlFs1SxHen6Tz8i
pWR232BIDaiD9S/6T4utGoH+MzoJDyg+hMk6y9gFRkrjqRrNS6UFSf2AROxpbU5IXj43oVUKYb7p
bfYv5EGyRNfYU3Jo/vKXOOEH5fWzqf6SEKCX/S2k6dWygPm54PQXzM6qhbiS4ajCztlS6pwDq3Id
2nplHFdt7NdCyA7AbQ9MUjHiPWLqHEyvuBfkv82mPu8/MaWhqN41F4ogTCkbxi0/Ok9VYalSPwUQ
yQy3YHy79qj5AXldsAGxj97JeQg4XcbE/RjoZ7SGdqL/17plz7HTy8TUJVCOvuSseTyk9LErt2uq
V2JivrFJwKcPDgVLpDFXKZs28qcjeUn8yL5Xf4onCfTeuM0pBIwYNWLESyX7ZRPCcSWxOR8bElDr
/8S1/hg5xh5qgcXiwR9kFLxO32G+nF/d+xm2wEiP7NPN2z44Dps8v5Lesk+QrSrP5Ny5nHFhiFeK
zmA21pIXmCVmSC4quHWELY4hh82BGvhNYv3LLjJpI3/ZntGyO+zibNQknvFdIZqsBdYYl8trLVQW
5VKVNgufbAqkKB0svnZ08yFC5EfbvqvjuhomBpYEkhFxNVK8dWmz2LjJ0MPIncEc/ioJZg93AWar
BMM0XT2JyTq9o+akAdxGga17o6W+I+h5BwXOf6NktxtYobQt+uA3TV2vBIHID2+1CjC2c6x6ktPa
XNR0kqWy/qWZuBXMB3pCuia3rFazZzOnv5g5gf26Zj6Y4QTXElQ9iQSBNhJm0QxKjtBP8VEyLQcy
A2Nm0gPQn5RkjpiqS8CUSXmF3pdzfiBw31YADZQnO3hcAuWes2KJEjfr0fSkNb/KfugEhh3vtpbE
mczmoMDb94+zFWkRRKEIPoxP7jDuWWhch/cJPIc7XI3C4mVGvrQw7O59Odw8W3bZeezxSgZJNLs4
Qkn41FAroG7pb6izE+kd1QfAt8UeBtE5K6K8yMhgd8/ecNiwQzLwnidRETnJjrgZitSROSDf+Kz/
13KKvHXKBEhXJA27tJPHhaOD8cIwcTfcyyR57xWka1e4McjZh2u9IMwAJBc9QjN1wrXbwxAVMIHo
uZ/9EKKjAWUU8d0MjjDDg6MfSCNwuugtqg8UoEmBEt/12y6WuwjeqehlfuqbdTyEAoyc/TB2tpdu
Ha4gLADbRzwsnKaIl4K05T+NdSZuwlvR2OCD71JYaVSDEUpu5Kl5YgL/jag5Sk7ipvvQsR3kSlw/
wPBkDYMs6gN70ciAOpvT7+J2756UeEIxshYjcV04RjQdxPHwAF7AxPstBq1gMEN4mQ+I1aPOdZfa
buU55HUoeKnHU8wCxSuh2pFqNPMpmWY5h1HZ21f602NWJsBVRKCN1B/ymUUHNmcqiYVbvC36GKrx
GN19iR6xaS8JMZU30GRARtYPl4el/fHrR+H9VnovLPhUfIw8zLcAvxsUZ1IQfyDgOzTIkTHBaFVm
nVIrKKa6pFWyDB23ddb6Z0QqWkixXgekmzmTJlZxkIWF00zRoG0/dTqskpUbbRKFj7FRORT23qKe
AMrts5GqGyRUZhkeTWB0kYbvFmUIQhZD+25SzvCgaZ3+AYO5E07XoJ/75Cy3F5G291bsil0aKuvd
aADW/PhOP57JkP/5X93qYEID2p+puhneoYsemp3Y1s0zRCL8kfk50PdLmLwJcfNIRLQVi9ocvF4q
kidpygqp5QyY5f8rPc2KKtS4USn2a1SPZ5w7E7Ha6mQX8H0M+aCJIfV/lSPtIOghNJVXxJosSCk0
1ODSW2WoYU1R3dCJi2wKppCpW4P2UnzpVJ5hRoV32F9UfHhd9jKF81vgzhfUaLi6pRw2stUyMcPg
jjNA5zgHApZKmkONdNnr0TlBr9JVBNM+QEa2ajVTncV2Gr5aO8ihMZy4NVct3Hrs7GFPHUy6AOcm
RvwIQVr0hFvh7uMkig5FYgLP1RDYSVwrIWmeo2yuQmEAZVnxC86AwutcwYBNJC7oxCiKK68U1d1z
L8OCnlxI5PjyKdP9RtSCx7iThnbK7/1z+z6Za7gQqUssGWkZDhooN9GO8bfi6QYkyJvbgV4TjnTv
A+hs1xbGHXtdCwXqIhhSspmL02WmU/5rsT0GCJMdop5o/EeHR/SAJ0eFXMepxBqqD1GAWvzyk6vm
LEKHbqWBqxYn6G1djM9V0lXSSjd1hGaa39HnK5/cbIIpRsAthJzNM8Ih2kwff787JnHhZZYH+Ox7
Vie52XaxJ8y5viKSFiUGtTG0xCwNIjBcLfgABclne1op2fTZ31cw74XIfatLECJUYvtK+BTduddR
dY9L2dumhvFKHYbMU/PazjQQ4cf6G+V5AqufFYSe9aZf1UO04YLfGl+17s5mlb3d75LpkWZ6PS6d
QPrTdlQFQxPQi2Cok2VzrgdweoaEaDdLO5UoBXR589eOUWU+eeTlWoB97+I9OmQphIESzscYOAJH
3azJDk/P9ktQlLUTeha2OLgN4id9GC2kj2yaIvEXnTuT+eRUPlIVcO8keZnI6FYEMIMsXBUYlZYy
oQRA961oAOs89uybwnHunHChJQkSEWAQXGkAhywAwVuDefjLQRX2snomcRdPmXF3QisBQ1aPkcOw
ZtX/i71nbI4JQAhlhdKVSHaLVRAgLXpJXzFsgGfdZQsZk/9kNM7fGHJ+3SOfaGuaGJh1Q7k6OWg/
prLNJwydWvZlnIvaujqJMNXD1+ITC6KdZtU9UbQrj/eXXZp9pI2MgGMv8pIDj8N2RorLNRpXPcjj
c09Z81SLNiF7tgB73ooUzm0D0UCbFAvqYpc0Di25Epmm5eQ8DklIKFSToxvz8krbdWNPznHjJqTd
JOnElzU79qhiLaI3i+sIQMYpfdvqUzr06QhQ/HBAkDYs0Z0wQuTtIHWpMXbWKkMIDYEWM3k3Db3f
253p5lnFCaWENN0A2OtpzKzq88esVp4iAcCa/nw87hkJ4iqlVptlWGgEbBfwBtb85opam2/Y/i8k
ZnswhNz19UpUlJbKMX1LBxDBFDrZ81vzBvLCHW2WH5aZNiy469nylyHlTFjVwTq2Y1CxrUCyQm76
0AgqsGhpWY0XHniBkdkWYB81jfbDKTg/CowjHh+PdRbZ/0eIJb9LoGYU4FrzRddxKYljf2fO34lF
gWBcTGsw4og46i7BqqzCA/jhZCgACmRn1Y6S8PVYEHDyLcEWKCqief/Zv+2g1uAmmN2THE0eceNc
/3WDz5JeaK7W186H2A5peeZvCsLjAzadVRAnJb9hUb+iim91p1qfJULPsvmP52QOiG+FNQR044fu
xl2hZd5GE7fEJPV4mxJ382gOeWD1K2UsuzPRZeDIfQGf6zcKwxk7+uQT4ZjVQGxILyXnvF7SnQQN
YPEgH89nZozd0qTzqz7CeDyzs+3RRDTtJbTx1hRDYFp1akgp0Ov8Uyp4Jzpr1bl+JwASjWMEDkI1
vi0hto7UzYEREnMpfYalvnCOclDFdumwTmbkSfmZ/ZAZgxvlu6GJ5xobZhpERRRcUMlcX9F5x2YQ
jVe2SPHkPI7iDLPlH9VaVO7pHpaRaDhNPAdUe4J06oNeDC3SSIlHaAqCYO9EDP+n7xbxHkLabXcs
gkfCgy6AUjXQD+gvFF9MCvyc19oK11BAl7yq1ExQ3NBl4IgKGd1HgFg6gNKgLNxHLLHQqlPPFg9h
EM9GM3BIcBhVOzmNkvZCRWv4pU32hXL/13v0J+GX06CcQgGZaY2Uu1CHZzF5gSnJ/nSJIxsu8x7w
/N4TOhDgaGlwQvWQmZNVRWvppOM4SZiKhwGyjdL3IbmUJU6s+RN+zU4c0V+zhiADqoOB2pnsfB6H
PXFBv+tL780cGzjJJrgW8Jpg4i6WRhbhrGVBsQjo8dvoII+qT1EYqaHhLfe78/ZABdDxlajQYIqe
OnF/o0ueyTsFetmFBS21RWc1AU14e559BLT7bNfGuznV9hlT81yh4UcZ1qsVyhegIqUQLv+lJ81Z
vDmDnAIResnALgCOi2vI6lBwV9RqsausLHeLuj9XK/fKNf0PG6aDUWgliAxM4wtfN/8yLsbLCeUV
wspwFKsAHQ693KIAT+Rb74MMJvJ1yqM3jyKZQXd9N+Pm1GwTKGk7GObZKOHeuElGrEj0fRrJiB4i
4nKDYDmFFLdGP34BgaP27MulJ5HyfiVCOpcll35PSoDwA4zXIhP0m9TYNykHwadQ9c2Gg9e3GlGf
ROrjaY012g43yTw06rFNwaRyU8a3peP5C1uV4/BPQvqC7eB4DefmZ7rWi3CzGjxNgkRiPag2lqjd
/tkmTH1kEVBoK0B3Q/nmJx6YrM8iag012cUxLKuBfc302P46GVKF4VX+YfXTP4hiy1wgSXb+4tz/
4rBGLhiwsAYcQPBRRmSPdpeD868nv5gDTPsxs0XzH4m+fnr9YqTyWti33WcM7HrKaZrUgk3r0JeI
LSBhmH4hyxoxFF8Z+OfxEE2rO/RmXiMurdkHbVz/AaLo9RXqfkorRkY2xD0BPMbCOk8TsUBbdC0S
HP5Bnot3VnoGdNS4bbf1lCda8tp9ZSQuAWDnzSIZokByolLAVlf9xB2CC7/ukAGqiQghrlX9u50A
iO0yPc+OVDgXdhKkVI1eFDYm49DN7G+IPA3j8REeQBTZHI6MytZcpBu2REC9i8pBuqzTqmfbVBqp
2RsD+yLQneMVqOxjA4gyIwnUejhLgZKKxZ8tEzYrvMGehUd2oJSh1nz4YpIIegqsyeNVeLBMcyo6
o207culUOLabph42oPLsInoQTbcJMvzunRgoVsjUbeIdF1RCHcg5IEcNZQsssz1pR7cuUJgtcYcX
x8SQ76p9t9XO+3stWqc7BxNsyOmc7T5SOo3A58xZVtFiVmv8loafoK3jzFzjygrriFm2SDerQQBP
xe+XONC+QY/DMISX9nggFg0EaIPIU/iuPqHsomfw0bPoBzxF9rclIMbE8yOvXragUkHx4Zj5qnA3
Dd7sJGQ28+Z0srB4XmLeUVFe2iJptVSGXrw2lpw0GECzymLTwqpBvlWRdz76lK0wVh1OzzoeBVdT
XBJWFzuwozADcjn9hkFpJsaTEQF3jXPpmRZpXp/PamVt4OA8/3cepAFvjhZ06lCLu9Bhx6k44sro
jgtzMQExXRhI5JUpzIklELqICeLIS2lx9/3vSHYaY7Qn9ikEQJ51YTD8sU00+cznvQaIuiOhVAAu
QnCooln2MSaJNav7c9kKfN1RYrIapLRIIoy/XoY7cOw7PezLZVzamgNituvFH7duySlJUYKLfrdT
FUECS4kum5gVfM0HJ6PJxgkcvnmdAUGrTuLyA+NiRE0ssdCn9wW0KBsgEAblIXwdEcfMuem6mlqb
SLT6mdd25gcGSEK0JJ14hxVmxjyMnVrhRu+00WkRBG4sAc5ys1jL1LSZrjevMbnVhF1+8e6+5Z0b
TCP5CT4LsIvDcrLGGD3XO+dsSpFMH5bkC6eukECmgnfRY0/frE00TBXjn4A+mDUlsaFlzvKjXVUA
eSItoN7/v5/7Rmee5m+OsVNwrKcWTUg9t2HpK5Y6HV8Mb+598Fj5vjDLTPPczoLdV/oxlMq2DjH5
PP/PsPXMTzAHUfbE+poQcgK/h0+nu51WsrkudgqKgW8LW0vdR1PDlKhZELNBarD6KMP7I76r5NtK
e+L/ohKBw1rlF5U4nnfgh++eOvySt7T8fNjUI3FbtFBBPOF663flI6yUbRJ2cE9ngTfLbe4Hu+fr
uuihFkSdoxkg6aDnsKrzVj0BC1dqQ2g1IM1+79VQM3XXqYW7oPbWitYzl7HkENUkjShTGSrJjI5B
O/Ro/ilfzlVJZ7FvBXCYIzlkffmYhAbwcFcrRAKSjS37r7/o6JAwKn2Y/imt9pb/EjagnPknLhSF
2wnzsbdIDDjBMaLX0cumD4z9lcvBGGiXyxc5I9GTLo3MZAFLsmupkf0NKbxbLt3WVfO9uEdwC61p
ZM2+gqk/2F3k5zsUTRmVQ2CSZ1HAGMNkKuJiACGP2uPoTw0oNwXvoS5W73kgQqlI2kO3p2IATPjR
WYH5vlgUUjAGvj3xDZYZ8pw2mBuGSa011qgdvIV6qFEpAJvzj4kbWkzYI3Pn7f3Sf1QgWTuBYs77
LlvZeMGyGZg5FrkIYM9J1BU1Uy4KgFQn3KqXPVrdE3BxPm1A7rPVjFcg8AmdC84ELI/TLpTXJxox
bwyQTXTSNH3T4MbM/L20gURIaSl0EDD95RuxroU+b8eQkgpPphyIeZ0GTfhJttmwughM0rGfEEbb
BLRnkj4WvS/7AgbpdXQ4hhRUj9yLRp5Ltr9PF6lVBucQofLbQBiQzlOfAElsIkYIke1iy3XDbcLU
TGivSSbgx73V1ORoPeBMuPX14+3bA6wntsSGvjqYxNOEYHfsPM0m9TEeTbHFK09ULch9erb2Agzg
ICx7954Ui3KvzgKAunato5WTU2KPbXg/9fu1+OjTn28D3AChlSqEmS/ytRhVLMgiTQ1+ebvqpTYj
emUIGs9xMS+CvFXf6KYZ1IWShXgUnUC2hMPWp13JdBQ9uKVLcQVv6xZ/+9XWEtmb8YuOvZy5gJCP
Ttffzu3iu5XthYMUkCKKnIyGtG5codW9x+263d8LoIFGkdBOGTNI4LxXzHtnVqc+Egv1EuRB1tGX
PtI8jASMHGm41XtQ5nk2VqaxiYXtZ8xY+NBTIjdeqtMcHOGCt1SbtbPxKpQ96M7iIq0k180m9zcO
IQRtugBya5UWFkCMX4fZi4MvbrzWrnYf1R88komE7WOffsBt4iMAdRx3aoB0i1EZA2a9LM5Xt1oo
LHvvUnI4cS8GHRP75UnBzJiLFv4Nn4+Ov/AoAVBraVWcq2VH3yfFWU/IUKtIVfYAiFAGaj4Bq8FQ
13WI2oAUJc2erJSDJsSG3f8BH1CbDFktCY9h+NjR4NrGosovD9Y3pMv/xr7xr7HDeZXKHWj8g4Rx
JPvjijOGsyImoy2sD+Wsd3iBxl72z08iOB8NsN4v5dqNIMdaI5NcRzsgPTeVRGCIxubcxqv4rPAf
XswoWmdw4r7DATHYXAOxF1qvLb2dPBXwA7J1E3/+O0tMGf6kenWjI1mDnwx1guMKXDEFa6KJtSfn
uhpiU3KT4pmGlHdKUIJi2fF7Vgvq5WergZKhDtxE5GT9qNSMob3uQLfsiHIoHiz25x8Z09RsLYsX
jrW2A7xDLTbKkKVmeTFp9vsTGmZuXCW3ZWPSV3/T5oP/hALTOGy4/iUSUZzCwZkyJ6IvAHbg/UmO
nVS/QTMMNXl5eprLS/HMHYpd6lhcXOV2dNIAkGzOOOGKnIYUpUdEvB0DBxu6+GbBM7+jZJBxfEIz
9CT2bSt3UgB34qNAq2uZ6DebwiWfF0FgmwlELM0Vl/ymL7AvSwnSj9FYMt6AGxVBI43naA5VwMeL
OZZnRVrYoV17UZnVIabSXMVEwPixOCGv1GJvKuuRXi7Or1dsYUzV0BPdF5ccvPKyyhGtFWdepkKN
jlX9EMd5IFxIZKLu5AcLz/Twb7xVblbs0oots6P5CFgA2UDuDGr/sxTYiVRxpcDonDOekylUSG0L
KI1lW+4ToXXQbXTy0H+MEEW+LTwvw4iHxJx0hTvxsvm7E6nR8hEAfBWULOgVFDdJ10j4HMCFy8o6
9uYK5uC90CEaQx9a04wLZVJYyhO0zWXvVfSedSX974P0iH5SvF9VNl312zjRET0X+Y5xUn2NvXtV
gzzX3djveIluKJ46wqeb+V7JAwSgDxmKbN+s/5244Xxrd7fdW3vLgbj+ccqVxDQpl9dL/CXe/FQ3
UPQwL/AXt1i/hZbx/LPD8rXyFYJbIRdVA3WGLgFENjcaK9Ld7XMNjFUVTCCt45a8Jrl2RhwEiEoj
hNi6w5i9AXmHR5ad8oXmykBVj3ctl1Gxf9sOLBtx0g+GofOAYfeE96i02YOZuDnra9/gbLaOYjN/
+tEEBqZCUoNHmJF2mxq+QmLasY/VBbihx/rqELMfK6F2MG59aPL+g5Zpj+pKJ72+AsiCp9hJ41t9
V5fiuU6GVlJk8CXGvTyDWcW8d4Yzx/7yrmdYExQGlthw6CTx5XG7Fbw2Pe2OobVnjiNobPy9XvXr
O6WCuSmiPCRqrjem6Jouzim5QUa+p33WVA8LoX+4DkPz3qyVqhXjWYYwdmAgt0XYT8yCpBxA9XmP
03vIVj4mGH/7BFktsXQJepTBZzSIjZRm+CjtubDtxamDGAnS0xwdlzGyqTDgJc0tq3F3hrOFuxZj
8mR/LgmPcjpqeyJ4BP9pWKPKmOkUS8bHdYlH9r54iOHpaoRU3KKSx0n4i/IM2p4VWzwoSRDRaYHx
DYql+fY4/JJb6rL6uhTP8TaQgAv00XW7bJBs90vrFFVl9IKrC201g2PtEL/JXQ8ku/zJ3szVu0jn
9Jbg7YVC7ZufxtMVGFDxxCe3lWJAgjdHTU6fNyofUzCYuMTL4Y3e/3cEpnEemGzxkP2TEkjVwZaq
h7pvIEOiPu16Gqhyk2G4r4Ct8gOxXk4RKRewwPEQtwKW3Ep4VT2ekM8lOZ2UekGifcMviwDq5Ot5
10xMO+KeXjzILH78SPMWhnb0KGU8jkG1JNT0c60zrbghdKh6CdrJAkz4Fh2meqh3e8+KZIYiSJ34
rhk3TbN1oO31pNlfNaMM3lHj094QcSeexNuBcTvg7S8vOJvNQzj/x2uak9ohR7Nc6NV1nvfMtAVZ
alTgkJi7NYcw+3tvGpcPt98iINGpy9Jf5p9A5eYdi6cc3sB4SNbutKdTarIATgfRhdVOvZ09s6yV
Hpuscj6GsrodVathOQezPqv9OEYpFniO9nsk6ynXO7q0G0xN/dN31iQSgFllIAOLSZwF2hDI08/l
12RPn2hnPxShNaFLlh2TdbwncIjYx7beoK29UNUJaut7/ggWGfcmQqcSR+F0Dgcpfn9VPIv70WZN
V8N8tDgNvroouNTZS4gSjo1YaJNnTaHYLeXgxjhNDW+ge2ZHq56Ja1XUdcvxCPgy3hO0LZvuEtfF
xdXuYmRAIHYjHPpcIxmU+XQPwdBXeJlmyQGgnDG2K3ia/YFE3jWVTR0rUDo91dCw6yDo1sibSkpP
z+GKo0VqdPmQQ7KttmSYe/KGtyCGGsQ4i21/+7v5nQdtoLbpC+XKdB96p5xRA5D6uabaZszpSheH
Kh1EgLhVqiRH8sLd1zuipwWA/8DI//QtFGvF0r43hfooGXzy//6G67B/61dSDNVW7oUJHHDkKFMc
m2t8fHNq6SOc8nvK2+uH2DBK8Bi526RqLkNfCNwJXkJE/GWBZLAJmKyzaR432IfW7OpXMuhUt+m/
mI88Bth/qLJYM+biodP+8tVXT1s9cpS7zNIXAltGjW0HXNOO/KjOipmtTbuIf1PJj45eehXTFKYM
6Uc023YJJsE7rCtXOEIBmwyn2YLDpqv8RtdkJ7j4SgaUNPU+jYbQs+ulq3yoq+q+Hb2qX/Rb5tp+
DBJzlSw/ql/Jj6AvJBk4HR5G6/BkNLJ7CDPA3BtjcSXQ0kx6fV54LlawfuKQgyY9Rzu6TzrM2at1
ZNXFE/ZkqRkE4/EzxVI7wFntXWA1+sMzGse9zBCtbkLb9nG4Bu+nNh3v8mzpKivKDY5ZomJKK6UC
OfpgALs+4r+//JODyzarBD7B/tfphvZiJkRPt/eR1JinZ/64TBHTmJ5wBb83wSFdHngz0rHJj91D
4dll+2Q3TZQpuETfoG68HuyddGSs7o7wGaD+h2n3Di9epDY3vjfLuMvoVm+Wxay807Ml3cIdJX49
6LO4bmAW1mjvDLGXHdjh5LENLxBk7krLZKJ51BA9oRMzUYwX9ith+L4KyFiV6Fzt1M1z2PtMC/vA
oXQ9VSOecIi1KJ8ILYuqOCFiHCang72kJvjr0spIDaoYf/wEiyOIJi24YwflppuMSfzz82pbGa9U
FPXdVSYAF+1D58eAIY1L0LmINVRxRAR4IobnPo8DYqpLn9bOlFHJ3WSzELtpolZMXyCWeck3Xdw8
wsvOIjBg3CiAwHRbDL/lmPk8S8MbyuAyflAYk2IcYcq3T2BS3pU+B2DYA4an72hIv3FSZKA0YafM
lGT9G34ODDVL6iOkBAkK7Rok5Dm1OJ/oCI671/acp4KZt4r0+7F6db4arP6kgNsseTXj/tt2q7xs
FeiIGaHlVUnAnBR/BtdI4LIVedY6kPWa8pa4JpnfWUUO3sZQBy+3hji8K6y8PctscQi066HNUQDK
kyeldFC968wvsxsfOKRNVZPy/4VThZxfHlmyQoG66aIL2WFY2wiAjn8UG8kLZBZkmRGCCJDslhTR
AseCtL2IauFgE9QrqlHVYBnylF2EPynCmDf9oYDig86GP0yy4Lwf3Yc9rAYCZMYR4DWYZFThBpaC
/L4+qDthvKH+I89mf1PzO5AwjtyQU/XZnxeaB0hictvw0K5vL9RBH35UBpnPH/a4dtxYXBeLt38N
IjRAe4rjw1LxxnnONAyxOOS+X3QmEIMFUuAZooFHH1E8bAJtT1CFDqXKPjlvG1IXSKhg7QUtkjmz
p/x6eL41jehcHYlYydSKpRh5LW8+MkierDgLjmadVKU1HERzaJVAY7oEv1jUbroMilS02G1Wa4/5
vuOYCFOxoWnfIeu+nB7PTjN7EoVtlaNYN4c+5mOaSAmig7GICUbuxEiHaGKNbfr83ajVPUvjVy0c
3Z4sP06MHLaA6FUtu+Q93cguACd0VAba8EVJc+MWp2IUmtjbdKzJG/t0QvCCXu869fdybqV7u7SX
e7fd3cby/0BCoVRZBmYhWEGUePLn0kiy9HpcQcLCwApYt9trKI96K0aLWyOZrvtNVAAJmX7FBGj4
6Ir3WnAS2K894+5b5iSrCAgq6R9RRZq8sHtcEHP0CoB0vMv22O2kJZStIGUe3fPltxAYAz52iPb4
ZOTvRcwhQY9zhEozSxhbwGf0r3RVR3hL5Q+A7fOcsy4EzWlOmz+OdrzdWdNQlb4Qtcq/4zC9/rBq
Fb8YsCjBt1JkVKV16xvnnuabTgOO0v472CROQ6ib6xopH+1uqn1LoHy4hd8eXlgCucJVYunR6Hbb
MDhd/S8A8vypT+q9MD+NHr1Gv81iOqjHBzG8TdzvoCL35pkfkWU90hHyar7PZ6JV21kch3/5kFFf
BY2ErkEwooh4oIBAi66+7hRwn0PmEVEdystleXBDKeqpuVE2AlxXoNZ3QqXcYUjM9AIdzxIHKCfo
qBU/G6N6XVoLoyFflM9SSOFIFKxPz9O0Dx+nvEW8HCJftkSTrY3Don6fx41YxrM5vfBDli/jHkHY
SjJRG2XjV86eKcmduQVkgRZ3E8+zIDl0s97Iuxh1Ma8Gv4nfmgU5haCqPQSQLyv/NH/QbbHP2iXq
+hTrQXoxoCCKF/6gfd5F/s7Q8zSQIdc9bDoAAjJAm63oJ7IABPSQO5Oy/yj47Q5H/ApP4SgbkqrC
XWuY079LT2Cbf+LLCDWGfG+Q5juRNm4wyg262SjSlOW53Gi9RcgW4CJYVFOpm8nUNodJmbRkuEeC
QKUcSxMrLuwzJ9aQuNKzQY9Xux2C3fwxKmpaOR8xJfvxQ1Tk4ico+IItZM293XBnYDBYm2hK93wE
eqD6VDejwAmffaivocr08Tr1HKCIfAYlPKeJR2fGkSilxUDBwzKbw2whk8vgWfXRdqI94RIBH2px
gDSKKCq8gTE0LiYRoRaKXpYqM9sMZm5W4bZhTlstV5bfh2QrSOe3jHFxcjJukX0quoQB0+nu2mDW
K3s0OTAwH185J5cv0MEpfqokLUwIGH3/wOsZXSR8iAptqu/5L075T6gHs7h0Qtv5pa+Yf33A4Zoe
x2G8iuvgvetci39iWbKyux0IwvayrHOBE5ZCyofYcBdmOdsTKOrAejj7RtfiaJiKi0btLmOc5GQS
Bme/FY99vLOOuexvVFogQ0EYRTl38QsbS07KwG6WEcuC8Dc7zsHe2+A/BNaK8RyE2zhHgUxdLAlN
osF6vNUlsmOqxUz6Jf5QdFjz8SeV4gmwH0DikplUO2p79fyTh6J0JVQ8gab659TJnP5PHjkgMFPD
pN5vI/L+wztdERpQIBvTlyJH6BVwiocdY+L5nXDeTVUCH/zUVvYuzn9U3JzXBjYUmcvfGWPlD0an
nZhbNBhnVfv7H/XsXnZxsT00Epbme+vNR6+6C/0bM3jBXtrzu45JrdKWwKwec0v4VFxc92KY3uRR
9sGdR1ByvVMvYZHpxCku1RxMOe0u1Am2Ke8rxSsLpW2Dp5PEn/HDcYfblu2PBTNYz9fW5rHgfCxo
NOt06e6PGompJ5nELgXgP8KBo9x+IvDiNwKYncfwect17PEyxkU+t6hHenRbNbo9mjebzsK/MvV3
VKR9/gGK4KmdlbzSGBSe+FmDwcN8cJyWhv7KYLrCvWJqsFXWg6E32z9qGYc37bStqMRvwinILn/7
iwZ45uv3iEwFZr9kH5sNiTFsS3fsdkDY091sHE+nUckAmKd3YZ+i3wX2B/tCVfTDesDT0c0t166t
1iYqm8ysuHDAOd7ciYcEcDWp7nRX5bebvRn/LQHA9oWUBresg8duypYsIurtHxhuN77zb2s1aDZj
r+2AeZ5yoEoP/UN924jkc7m9FZ3XwCj+LwMWp1EA3bh++7Lxjbhc6BQmrX23fg2DymCPbDE/XENq
9fucBpfUtrngAAnOsPkPLxrZXSDPKBssLkuj2bY1o5sucUjskJdGl5Lz7ztrdtq3xgNHQ1IEXhpp
MKT++rA4nYW7SBbslg/XPDV483IuYWlwHRfd73GO/uO8JyC5GzwwbAH0cUI+wCawMoi3bp3ry4kg
yq0n+nGwQ9fejwotm5cFngO6b2RNj74dF44zMhEJsIY4FWNCzvnhoqsFULbTwtoqEyI/RaYQViE8
STBr5eZ2/W2AKjq/+CgZMqeedB9dHBPaNygHFO/Fqb5wJJQ2egXuR7A18FGVG72QQFsKyXl3eSNC
lRX89sMhJ5SYXqRWDLtINdyk25GrHyO+FT0Nfh+dvR0ZjmiGZEaPr7VOopNvzuOfFhxAezcnP6WE
LeqfcatbknmiXLHAyavcwUh/20Tg7Us/voNWVNALMf8iEjmmHErHUtkQrWD8gJip+DIGjcN/hMYS
9zlRxdCjTh/D+moeq2vMC9xVdbgdFEepNCQ0730EdEAp7TrMfZXHjcDRhwE994Owf6mnuGHvFkZh
PMxtPjEJe5xP1oym1gfv04m31XyrGwuPHN/DcP5d9VEzxHM0nwmchEt0DTeIlSjH2Q99Jzdwo4mH
lFPLMfMmpAxt0+0+sJ+o9X7WbNjHJ4Tgw8cfyZp84Slf369XRUBDDlueqUfszbIiO9CUkapu+bVK
0rNk7E4VAfe+m62ye5ZXSyXiTDm0acDpTh7/kHgFSJCA4R5fbpNLT6ajgzfP9IV7wDiwpBDNn0hO
v77m9IcnuqtAWKWoTYqlhk0X6StgyAzCJmfUrwW5RISaVDPNQwMEv655C3vTdzaJUsJjzEld0ijI
Y+CsgigDC8fRgQHcF03cNuYG9NQu2I9VvkHDZRga3+EvgagH5wo55udpW+k0zm5nPzRCebWMPbg8
wxx2Cm32VNO82ecxZ+94RMhhn7cL4/IzFxozBdo177WtMr6gIXtl0Ec6t5JqY4sS23Q8i0u05cw7
XVOJy2p3xapYXDGRfDk8hOCYepGtKmKsGRDeEXCQeWRRhG9e52DQFGE2mwrnsA68AZ6luFv+VmgC
HXKe7FKgLyOshbm/Jvt+BRexT216Xkxv+kNTWy2DjrG5MO7n+43HYoDpsVSKZBkwR+GZGZqEnutP
zcBnLJvTFcMXoAlZMj1kaSK6cS2jySglzPTgUIfBUWo78Jwa9P61X7PZGivuhNp1CISfSbjqDMLq
uw3HgTwQMuY1DOKV4oy6wPfXYB6NCUSs19X35Iu6ROnNJ6/fLyl0G28VkGoROdZMreb9b5GCi2Px
nyeK+J7EXfSZ4okMHIHZvl8J4jepRN57IwJmRjr+0MJzqHtdiVMJZ6VoDYVgLoSU5LTDnwKg1ybQ
yNjAOEZzHOYTFIi+KPKINu5e/b3WNsh7AgbAIDaKdVwtiqeOlYOjryTw10EqjJHf3RJOyZr2GnB9
fO56c1L/J8WkzY0Nqh+hCY4e56TQfC/1grJ5NeiwU4RVpIAXcKribUJvSxDAn5/5TvJc384Zkt02
Hnp6Nc/oM1GJd+lUNxP+zbqH7KzfW/JXwMo9JLhilTEHDn52xbuWvgs3cgoZqXAJtLy/+8gIoKC+
VchmpEbTiMA6t5SdM2lwJljldHMjSRJbRkMtAdPQdbU2ovsx/mKSlEQoBDSk1Dy00qitDBns6wYE
O4mFxKUunPEibV7eYk0r4O4wCAOy65BITwf2CTblfnDrckySNSXYbcL2vbcAYglIC4Yl+rudy19G
mnXFOhTL9IBOc/6Kz8sSNhM9MRWYZz9cFfqyl4ykCfRqfkzVNuX61qKjKwuvOX/7axW4jUphkLWD
ioo8476WLFEbng+1hGMUWJ/SLYt54xWaObZRBnYMyg2EOHYHRpteW07D6k37Ap1sofxK2KiNJtbG
2CgxxiNuFvLgYoeeZgzJdvyUi/A42jAHDylHTp4MNnc7cdyHS0+zywZIIqMrOmwty+tNUacX33cy
JcqKEEDUIJA5Zm1fsuaz6E0Cc6Rw0wSZh//D7qtcsXBO5K5ulBaEYpgSPTJrxkD8pnTSbjQtup6t
UCfIkeeCg8cey3kdC7I/oIXE3Irnqeowud8qAMduRsyNtmT/xUGtauI+2ZJFjvCX8i+Aluoo2uBk
GFMBJ1uFiv2CKPNPRhYB5J4YHTzV5LLT54nphXBrVWenvmTQ/SgYq3gtI+ccCeu7APN0SdztY+Z+
fxHD2uQetFFMRPp1Dg7/WtNclktt+3sNAIuXeaqgTFaPcV/+eDCD2rhuB6F2dj0inNWROn8OzJhd
3f9IaLfrQ7iqqLIO7KRv1kofJ5/nDFJflU8MLLDTKD6UJN4WmP9PHrXlyq4pkgLz5HOqwrp88jfw
Zx7l8zPdWAdNMzzRrXFpq8ZExd91Vg+Lypww4rmcg5O+aok8x7YuZ0vFONs2rN5kF8m6x8cAuISN
WiddelnbuXwOzkr0i1R98Z3fdwaNvJd+RnL2fG89F9tfumG41BofXpp2b+bmdftyNssBCRnIaKa3
kvQLjw3hOWNEUjYc7lj3pKuHqoS+ADoVMzbUIrs8h5lUAI2RvMWNKRGE95rWg07Ivctr2St+Mapl
iJ6k6SbY7BGf6zff5N9chSoRBUTkIh16nRJCcew7TTBhJNMUKP4VEtgs9MjE6ldSQb0IyE4UsgI1
dU+ML69m2+giQs6+nVPWXL9Exu+B3RTOENSgHK/YzioalbqzaUP7yKD5gucP9J1CqxaksmKff4nq
gcws+zEkWozVw3jx5IvubBtnNh/0sqEkGI2dcBf4J/UQluSe5PHb3dhgCnLrG5SCOMD3rK2tps7G
x/gWk4bK3eMsWgiH45JTCsJlFkKtkOXmO8YdQJ5VYbnZXtXb3e7HBYuSMzcUD3FUd1BHLbmYYH9H
TWye0+L8vfnbs4HChD4Qa/xXC5fyzEL5hfVIOGwzzFgQYpQByv1cm4Mz21DVyF438c0Yk+4EZzTX
mMG9AFeVz28L2zz6JvhJpVNnDzZsMX8JJY0xmIImwFQBdBidGCUs35lsJdFmqmgMDh7/F7RtT4bx
mwYIV82fRIJT6Z3bA4+bO8k6ITMXfTabCgswwpyRTD8pH5aoEtL3m/RcrcuTLI/iCN0iWaLCsECo
cV5kAUMSWZ89aA8Nw/h6+Ay54LFRHLjLwT3EtvULYOzfA4yzclxJdm5dUI0HnYKmBJt/zrV2CLV8
Kgqku8hOGZ+THPfFa077ubQeEkF/Ukg9IPZyK0uPCpWi+D51a2K/AiKBlWPL96b/8+qBzuT4p34I
Gx7nguBw8OCVNLqdyf8ZBU6t5ABFzhHYA31pRpEC1PAqN6Chz9DJhdpVd/8qrUUa72oruneoG6mJ
sdHdqBg0hWeWmASKBpVoHx/auTiimqfBDwHJfr96KK/bXUiSjXLaNNF10o471hBz/3op95o4JTgi
X5fSHXmZThngKFKJAWpP6jF9rWIRi4UUUFhIu06Ph6zLg2X2cdcYW/bPzIuK7BHIw2K+fFtE0UNi
0B6FJZN31Lxbx4/laKTeC8VS4y+/MFWgJVZKIIko8cYKrrWSOCdnXHZlq6A7ju8MKhNbiu7S/UUg
fDikc8KEWHyjXIdMwRyYsG1XR74v9JvZjOucvp1mGOumMZnHfibsNoyJeIkKvLCjeTBq70Av8HnR
aLhfDs4us7FJoP4dbPNAIoaDHD24195dLRxPPK2+GnsQr1bQcx9RG4UNVGC+Xlr5+x49eei30K24
yPWNHsvbq6uWbKCLAsAsFFuzxXlk2m6QvyxVrO3VDjEBIVblGM06YCTPmwZEzQg0n/3JxdK22Qdh
7MgmIF0QR/IjzQXsKszmCt/55TGRTFo2rUFuaR4usI2M+IJUmzhKpZeRa/60Q6KDSWF51aTnRVWm
jfft3ZVWmQi/E9U86Oqrc64F3HCMj+5/RgmP3HEcafq1pugu9L0We1nOhFg2KpUNmsYKIaKKMIo9
OIMQnJAFp/mnI8l3idQX1IWV4fVe5lDxetOKJFtt6ztPkwfcwpG4NeXP+6dHkP1WqWx8bmd9r+ST
bKp2MHPD63OocbhQUuc4/fOlewMfH1yKDKPP67Cpi4jtNqH3Y9wJ2qWc4/YTEavGRQ7sU8Wutvcl
BGBQIlRA4A72drdmzTCWnoidN7O3kvGkI/GNOU+UdRKyWpXhaio13mqcc2QHddEWyhfc1duF1CA8
QaEwIeq2ssgKCLLQYlIykBpgGp95MW8KAe9DWPO2bj9Fj+Q+ObdVKCDhy+dWoBZCre/8wDwYeVhM
l5tXwzmtKO6GRLTu3W31btJCTHz/afYtoeQw0Qykeqc0zvO8TYV+wqfPQiTKcr0VU53FEWFHT6XH
n5DQPVOQylFpTYP3y7RNkhVo4RBRSG3p08bHSpJjin1M8WkpUfRnpexHf1fIDqBhQe8OFfHH3PCP
WmA6HZmidGLfDpSiNmKthJyTo2MAFhbBq1IWTaacFbfZw9eC6WijziPRjqDyGDuXm7YcqmaJCdyt
tIAhmImWlysGaV6+AQHKUBFRMv6AaOleWHOmEMT1qoIa1bDWImjEA0R9DLYMvyYoHuNjHexb2CF6
qi1KjnSKYORw+vNvC5+CIuhoAC1P+gLEdTBBA6gbvDTo6qODGqyTLC9fofdVmkm2QhzOhHrPs0xg
XHcadyu5eoBbYJtyw+i3ZRlSmo8Grie2galADxIE1WcYL/j50f8D2QzgnEojFfN10YW2kUGLgSBb
LBmfq5uHI6wJt1Nwi0Lx2BSF5yZ9GTfAaffVIP1LrqPxLGlZdlfdtsVYz08tIvjMDS4m/wMlP6UZ
m5he+IZxrBw44n4fmORx1PvP385JVWFaI/kYvsGqWkQhEHWQo6ag1lt9z6Zd7A5ldeYqHPXn3tll
Sm2WUp3q+A1fXvUAfejRIseWx3A3deaw6tPK33rR3K+cEgAuLXiYwQ0go5lK/ewJ20nTrtNZ4XK5
gvrRp5ouuCX+HJBmHst3La/RrH7AHWyLGQYZMnisi28iL2O9ikXW2Ju2XPCB9dtkv0538Sqz9N4s
o64uOEakjnXUMW2NZi4D5o8Ro6kYS6Fo5BDizCQW+UehIfueYuVP87tfaDnyZvnwSMw8oGBf2Nri
OzI53ilgfdRkmYowAVb3Xro/hzoI5fr21NMjr8+T39rkypejBmK1E7aPGrhsh+MigIhbc450gf2P
vdN69v25iwcVWaUqnTjwkziWzW+KMLKQV/OCl+8DL/eqoCfc6QVVD3xDMUHTvVWoOqvsrktkc7Ts
BSqc4SvIxAcmHJukJqzRMvJhEE47E+tDAELbMEC28L49cvTWanUEI/B7hMAsWO4P0qNQPIg4pT9J
7o4TMwnqpV4zGqWKk+WhTSezIzW79eUW6BsJ/WiEaeKBq/7K3D06pdoRklp6jSSHYDTKCr7mtnTm
dR/stX2I76ibTqvvlsDPNnzlb2790MQyMCdv2qIVBk0wHJYEcy1XfKsrJL0uuKIRYEp8v/+bGkj9
LGiBUzkcu7sKA+r+5UCLDWUKOEmzvWaMa6D8sJ4UxinJ5COZwsDYuDt1pPJ9fSzARi8+yYkgRFOv
Y2AerzEgvCGbKH3eU5Ftic1D8PpxT23xQ2daYZ50QrfbcHb2ZfvLJodoj5MLLu7/6gl0UmSKB8Y2
yJA7siPUKOPB0NU5Khv+uTSwQpgVoJGYHIzGlxXNa/QaQaA2/jB1PFrEVMxXaAWF3UxzH6MtAoLC
s2qFJ8GCtDujlPW6vlOXjaNug2/tgkHIY3nJ4aYwp7cLHXn62kd67TswlwkCSPl5atwaKus/ShR4
y/tR5wfpid1LmjhsJ9KFCJCyCSi/PqKdJJzPb/8peZRkLi44T6AzPzG+eVgL09ODXPBJh9Y4Yekh
yOR8MrfYfu3j8YXalVegB7nLEn5oUg/MUSW6Sx2nKW+CJsWxYucaA7WF8oIxXQVeJB/vPAj6Qimq
08jvPcAMN1GtqO9fjwgHPBiUUeLmIX36hAE4t+V1+7JrxuUQs88ta7D+V3Bh4TP8Wcgqargb3/7Q
XBrWKDYzdXAvRBgyZkTyNX2IMCM++rV8E9MSkJ8RqXD5xy32AdNV8rA208xR1iEtNRbdIZAWL8Cq
lNoKgOo2NyaK0A+96VJ0TxULWJ8WNyKtlmDllXVFAr9NNaoxcC1XUUeAlguzuGvZEdu8jF4aZ5QW
VHg2GWtV94+ErsjzqqG0nR9vf7Gua3X10r1P1TXGotDd9NQKqdi7pDpfhHHiDaTC94/j/WmX+3eX
nTRr+abELpROpw5E2oi13571LNWrVqvl9MZ8OUcroeP/sWvcLqXVtEJW8P2sJltMr72oaSaJjgxd
oJdCErlL6GfoiBnbdAQMRUYZnQiAgbBQl2oEJcarIyjFG8p2pVJ1rGYGO49SLR7pQ2eZQy2zAH7P
UnJBeLmq/xuwofGMu5o96tB1KWKSCaMUJJ5AnC0GUblkzqwjBwVB+NqQly9qi39dXWMHLEPPi6Dp
B41k50tWwYsmDPbH8yP1oZSSGUx4C09KVwAxT1L0kddcdJOSqywGy6jbrSJyI5VoDpcTYelaBJKz
NIJIb67NC/WgcXnrfi6foOEpTGM9ohoZhh1arpWo29pEknP4Da5Ye+F08nQSizrBORXbzLkhiNsN
PFZEeYIaZ7HTCMqWfxI+cGw3OGHGSBynaWaqEBnbVxMwyFi6fAvdEvB524lm8jt0Be4Csw723o4B
pHQcz2S2SXTvjTd3MbZDL91vUSLWiRmk7b7ztQk12ad7HxN2XAxhtXHkbPZH3uu4E8DIUhscjD7h
zEvw1aBHsrMEd1hrbbXx+gaRFrPkNWFYbozIJrAUO8dqxzhKJEqw/Pwii1OFzGejcPBttfnESj7h
9tTXUrjsaDaYS4rRKOFnSb9PONUPYvhNofz0n+QuME5KSgL2KJiHqKAesss3HbnOLIZifG9aVjiX
Wm0AAx0IczI2oL58nwoM1BGN5oVjZY8ZS4sFPlrsR1YoPkZ3NQsQqBwH0GuhxflIvtsmVn5GBUC/
6UP8cMy+OqAiLSGp0DXzHYRy7DhQ7U4yOyVeTn2qSiGy21J13wYGJ3Aur32s7larQ31eOolvaTz3
7xhY9pN31m1hhDr5ZoZQua5j+5gT65ToJG07W/Rt7zEuHRSZKwQEsRL1ZK0G5RgJkfUPXLIPPbWq
Ne5C/RStMYej+xT/5F2KLDa4e1knhTGEDws+x7TrXfJpGEzyGG8PtYQPIYVbCawzz7e1Gc4nBfKf
lVZ/3qqpRHN4DIADafjYLLJXD5ooy7b1zuRZn2zz5r1sMDOGO/k//t6vO4J2BfYOMiwX/Imy6diy
R//1EaZVYN+zi2zLLgi3LLV52ztLVWFtvk554V9mcYx2v0IZwt/O/1DZECtlCEVVspEOqZ14MqVS
XeP2N+31ecPqk4ZYKNg8WFhlfmoVvzxPu6L8MAiLLEy5ugdoIuk61Ak1nIeKVM4YnWrzR1G2ksav
+XQk/nzX3HoFUO0JgwDyV7Kh/P0/ZWVnqlHhf+oc36fhYteSyThcN89XBwF1DBdRuFr7+bqrzt6I
Nf8NDvGCZhq61McEQSU4UI1+OEB/ZJ9kIweYEf/Wf5sROxpwo9AUN9GBSXybgCmbGdDZZhtnlrTJ
9XxQ/KzZFeS2Hte5RCbTsfGMGJbRzh3J4zK4LClqIzUUKp1YPArO3oE/t3Bq15CL7rCEnQlLgf4D
e28xuzxL+7CxZwjXmCXJf4HRogcM9j8hS/IRDcuVTwubRYpfnNFMDybX4Cdu1rkICXq8SfaKvkkp
NrTgP9vVYFxdlIah4NyqOk+as76bEaRH6FEjnQPxGm9JQGXNuuUHVh0Jfi38xJz2CXe8QSK3+pby
bkcOJ5iebVZVSTRhlM7JGwDa7lkY5ll6tph844sNyaScx93bpZL78/JYHEVPw4IXmLva09iQZ5o+
Gnlin+a1cG+JKDOEakAYoaNpcYOem8yCwz7ACJbsLcDkfaB6GuHZEFRN8vpFg3qxQKicyzEVfeiA
AG+ay6iGnnTC8kSjAWHZ2iyKyFZRc8l1jOD8K3d/xF2Yj+5VMBf1amxh/DCbjseoN1uALT5Tgdr1
BJeXy8+rWh9IqGaQX+BAZlqaFvHfLcWRova4SEVPbex+aLSRBWrYUN58jHp/T0q+qrHo222SYy1v
Tso/Dm+wUUUFuW5WX6QMQyjO6OF/7ok5M2/j1qiTbZhunA6KUi0MbYIjkCiwOXMDztu3rQY+vZn9
FaSwxHUYA0eEzmdEcGC/d9apUyWupOtJiZzvwMiaflivURA7nnGRd+m1hljD+hqM/fCyg5a4JNiK
9Op8r+YHaqRscfxkSknT0zJttxEPeEq9EXo8xZANUgxRnOtx0t2ZR1rY8Vrjz3Rt7P6sDLGhqsGP
pSAkRu80R0XHVmJfEoMj4n5tvs3wxch266k4B6O1DmMVHpKgzt+pvbsr1doikiiJHv0qJMLKG7MQ
WqpVglK6H6VunF53tPUAU8Yp4nLqdBXthQpKR8QB8HspXRNwrvemAj8WDSMTPy8JhR0QCubG6gqH
qwO48e2yg5Bmp2ysxVE1wA0sNmct/yNRrL73I646ox3PllBqHKxvMrvpg9ksNEK0jZ6ORRoHtcMT
5I3L2I7+JiJV0psHvqy8szMQHG57WWAV2hk3mWP6BbXiQpheBg2+w4hLlKhds3LfTFSXaWgUY3jS
c74AzPKk0FJTaNduhgYRLo7yNV4zC+7ekV4Fi77ieNTk1JvsqvwCgRo/f84pAqN58n9y68o/QOlu
ZHlJEy38EUF3XDOBZaftS+CkTrIOJVyQE6rlz83mUm4qeBilHFz+znfvv0OoqlZsWiwtLdmlOviP
dx0VAwn9BMPHvKUQ8Wm2L8PtJHBg0x27C8xfsiR+d34cM6o+Fbk4fPiXuetGUXRuBkZZ7nThosVS
AAEl7oOFBSw4uCazGUOTsmSOLXcmKSEhoU1W8M1h/TSLEsUFJd6QvgwbG97y0hVDAQQx3+Yp46Ff
SeSa92FAIRDB920tgz0SlaxW6gUoqrSjfqqHX/sC65hnuD6yrWdrU0761xNZd64wtmFjFWhHHIh3
fz+J3lQtEAZN9+V04tyrhy3C94ZcJXA/WGUMxNCuXdi+F/bL8dekUOvELixtoZPbBhZG6Ox0RUed
u3dBrkzIQ6ShkGPy3KyxSBN66L3e9rj4Z1mAF3uEqyAiL7FTB1ITAgUAxux9HsLGtD0utEOBbpeK
UaXymVDQ+8M4SogEvzCOITXu03NuUSWjfqeEMK/Vnms5ztcrXTjCkMlsgDmxvmZl7Q8YFy2+GqCl
5yQpsN1qY7sjqNKFdANxBCjMUghH2po2zhfUt53a3XFx4r4OhPAJbgjxeUnFknLrz5MFnQO4a7W0
7mj854M/jgGGQqyJHvC3iHtpZNSmPt9H5MD0bZWCNmaAzh3qEBD28PA8h3yy26n4UDpKeYBPYNw6
3WxrmMl6STcFeYNlmRyGzUYRna7UKmV+auZhEXLbDeffF8mkT8qcTO+coa5JFe3qbAQ0sKYTp/A5
+PrX5kapY/CC4fr9RBQSHH1KOZ7Vrr6QWVubmEsYeJJAJ6a3t56Fbmc9f1trTlJ/8mVLwphjATaQ
bRLuWMPa9pPUoljvaHsdVXMMmK2trtx53MIDAjLmsTmq4BVT0oWBk2Pm2JuIegC6tVL+ySyUvuTL
2z27SrWPjfNBoPNuldzxfl9sTaKfVdT36MdKadDAvKVG92wLAOo9dqeA9qGPpGBTzAAh13tPFNfR
GVAk51hSpdGywKXAk9Kjudm5o0t/dIf1DJj1Z0casiRsE64c+MzFgMwOmjbX8ba+vN/jSdJJABOn
9xjmEcMgxDWInUDasP2fUzrzMb7CAc7PU96r9H24AOHzXEksYpQmNUS0u32ReEDcrFigTHEuDx02
kZftZ+BJLI1H6KoxUjxryszite0jFY2WhCOJDRIZcVZheoFkQjalgsVgfUUdxOGzpPTmj8L5IqyC
Pn19jzZX7E+9u49Nge6kUUUkLgb2ZOvykeKMp14O+eT/pIvxeLKhUjc598Lu6DM0USlB+jdnZiXZ
k+V1HHNgYi9CHs5rc1aoFq8K0PeDT7Q8ydbguZhySrAveYIhpC5qCCFkyXWSyPVaVDicWcSqZbG+
TCmduWY/M2NTcwRKN7hw2nTAtYgxY6NyqlhlEHB4vqfhAMitKjdhV1TqmDENhsHpoUmwE89EwZhL
a0Lcexsu68owcPW7KlYc/LpSgyrdD+9jaXAW/k3E67E3zaDfBX+Ae/20VFLVQxV7uy5Sa01XR+WG
Gjrd5e+bIa5el36qdXq2ROrpqpdKbQ1lec4DMq/eGOJtnHOU5/kTy7drFf5H6FbHxwDayOwD6yGp
jU1AtwvolAdHPGx9VXlu5Xln8qbDtYCxmLOufH4P1AW7eZp3bO0x13sxxelf3gqXOwT3MD84aGjb
5STdF3DyJBytlLqRPmj5Qq8V4YW8vps87nVC+tW4r9CuKNTO7Inu/xMpfNQObwwRzesLKmPipy6E
TM8YEXkWjzd8d0fQnjpJjmP5Ori1CA3Jn/YyZTtR3U1mSp3eKP/iy+dPc9G2IHtGFUThunC5dgA7
Tk8YRulMQfa5jx++uqkXPyHaq1WKCriwtqtfAtf5Z/MKGGJhp0uYNI3PnAabWvHNjSIzHl7876nQ
0BvlzU1NyeMjvyAlnMHu18v7U6Skg01yTbJQTrOpj3UULsIB0oAaNIVsJDYQ/UNR5gwfiwNiWBIT
Gdp24b9/v9pQ+Ap5cy6viRLMW1TZOpYHMh0JUni/hAvZYFXCMhEEVXIlS9jKhi52GklCMDzcwoI4
mXtiyvfgp2q56MYjhgFRvQHoCoIep7Jlx568aYGQ468Nf1TjAA9Y1HEW/OlA9EAv1S1O1I0eneO2
prWCIbBuf68KVDoicykueuppxyesdre0fHA1XNiRgX46t3/Yhbv5Mzw3JuqpQnMIfdU5MiS0NOG4
Q12hMg7so+PJRFglwOZCFdsUi6aG7gk1nc8zPuSxY1G9XmfRsP86tmNDVbmMhNpyNCFaJtxp84pk
c/9rUpOyv3l4h8uIt5mAiR1gCrXhk5t3sfN4JrVMR8L29bYhWrYeGvAzitiQjlolefN5PaysHCiM
f9y5JdcdpksYar778U8p4shQdzFQCGZUfF/VCMn/1PNqjHf4KnYHZBklY4UGPqLnyfEHy4V3dLTY
CgMxTwyPgy7nAhswFc8wKbofNMzI57bPJD3Yc/rNEcux1PhDsHL0H0clxH0Cm9VwwpgTd7lsnRVV
YA1cOQxk81936waBFKCKyM0KyJxipIr9NpLm6LtS1kEiRdhNQxQ9z2o6S9ZtKPr1J4bIijvE0oMJ
I8C1YTuU54lmCZaI7HfDexpFbG03p5Uq7HLUlEvh2+hSTdYoViF/q02TsTiA9hWJpmVEn+sXhmYB
y071cTlKpHWKzk08czR+kXUIDR8HFeh/vq2pqcM7YHV/IYO1vIYxoXNgWL74yFqGabeaZrGVQ9cs
c1Nvd5e6bKtBece/15B5V1f5rs1uF8KefxX6Oz+3n2KG0NdRLqLA5BYvQWMbnT19KqAHYNeuED2u
N2KVoTaFFJDrOYGMtI7IKEnJI1dWNhTKyNVkooQ7ShYqSQ2H0BTvEW3rIKEUIk0mhbskdFbSbjUg
pl2/PVmaqiZ3B3o5WgWesQk2AfhJKrF0hIpCTv6hSGb+1ga0tSEFYydGDOVgIvNGuWSc9/WI4TnY
5zX/aMr+NmMcHSROEA4yCvCY16ahC7O11TVALdCJSxy+TE88+Ps8NUJ7tI4/jp/ENsNx+iVzELul
WRS5IV5LNLK+ATO/T3IHS0v4sLCYMBqi0wLY/RK1Bz3y4Ni6ZzPPiZUZHBiGU/UZVP1LK/qm6LQb
iuxV8v+Jnd85thWdA7mJDi6TsEbV9kadyEHbO4rNMUcsYY9uoRWDoMxyRq19eaZW288lr8IqgB3h
hv8ZX8KAh/IYXnoT0J1YRLnbYl5MIdfWmg+IszQo6cDP5YjQ8WHg/iG5cTwVyCnRlCKXQO4wqylF
halQrBFb6Lzo7au7fj7gYryZDfKbJur6uX5N6Iksbq5alY7aW2VxPYYglXS3GfNRRhve0cvLhIxa
ZHUpZhAkhMd8kjoLwtdcjzKdqhc7cIvfmVgoik+vVsPp2UvWpNjA4Tau2bqfnBI+qPlOpPWCvaLY
sc7Ka6zLlpI1xNyB4q79lpGbfIWBxvX7JsP0fvonh1tlOoZSPd7Uvyqz5UqKjMLXCBpJwz9fWPZA
wfqo7aBfl0LzM+FOmpP49ZHUnyo680iCTyqHjbLIaqi7aSV1M5RJQPE9fbsOS64GamA9BrzpLGKw
RJrhsHtRku7+DbRyZ5MqbUHcU9ibrwnWLaKEBpZ2YXV1S7IXvqeYTDZvoKwiBmqVehukugc34YOO
eJ9c2kjX2OV3nn38x0sNz29ZKUI3a97Qj7sWvsLRUqY1zzF11VBmGJwgPYaVrQkcz4wQBZnZs3D5
M/CgmzvmpbjJctrMJ+97ClRmdfItBOf4mYJkxQ4QjcX9tbrQAg7/82BjC9JbtpzEQRa/rC9ko+sn
RAj4eDQr6nPbxAxirl9BE4iOXtSHV6I0cw3krLia34UPZTzhcccy7r++Ih0PZ7gl+kOBEHV7t8H0
sB/D639iOXjK6pRM+QBKVj4lH0u2lsX2SImpPM6cJRr0Qk+Kfi69r2jftj3avq9+8zeIKJ4Fzf6K
MgtsQxFfqRD1gD3uB0feGAzFlhNovVZzyNYjGkG50bSkPY1xpjHe8tK1eu82Ydq14uJh8BSJ6ubA
s+dVnhfcQGlk6ruepg/+qkh97wmyvW+7mf+LENOR8m0SdW9ETvfi/8t0MwEri1zMRZltEGIXPE62
Ps6BSyiUmT00GVVwxMoeaESvYlZ1eyr2ntXm6HN4xE3xGGulWwvzspe3J+qE3nLELjtvGrjMeoSU
6AMBl2B3PuxZKNyOC9Ap31M/U2//wCW2INmWH9ixs3QBwXLhDIH40ERVujYUkxQ6CZP1F2Peanot
bKMr46s1+8u069t5AyGCYu9NVdKu+wuXx8AbuVkECFcmj7rhx4l2VAscpNy7GnYOBxqifmOgxUqY
Hbb6t1jfXcE+Gz2qjZoRxaqg5H3VxdGSMILlgoGhhtlIU8HdwfBLEyvFgiUo7E6CNFVABn1ycRJN
IUpw7w1K/5Xctt9YnF8zHHIOv14kSQMXjar9OYEOcy8lt1CLHzWFFzWunLPYkzyuALctOPDfC1St
L+zDq/nbeg==
`protect end_protected
