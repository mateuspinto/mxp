`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
vCxLNxq1W5X5ZFBrh8HCJ7lfNcjM9rIYMEgIrQ/2RAkmxe934uiVQgbqJ89I1jB24ucgy9O9z7rC
8i1u+qiJnrSGeDlJZYH03GBBfPd2wk31S46V6PUtmeaPjiYo6I2RWss2C9SI9xuUGGPrtwhZHe5L
n218Yu1FL03JvI46J9ap1aBNMBtyYs5uedRj1vDG+32p9pzptSgrs32/6T5KJU83itTx61ts5ovi
0DhRRSx1zgk272bQO2zFQ04QNi8JWIfkwf4eP7+TBgHyJbUiIOmPiflseLwF7sMicpMbecP5LhK3
+px3+DWHfZqjTkgZrISmbI6oGo0nBncnKDX3whoN0xIZrjOqiPINV1EnFmXGv66meavSimCmD0NC
VrO4TvRjDGCPxgGNfu3s0VO0PWyeJ3GIKQTK2GF9A1v3vdTs/yvBo7/YLLUZv0Ljbg6sjkcTuqaF
vGW6Q7VaJLTaGgqlXwpW50tK6NNXy/Lf8G1GO7TsItI9bmtxq4Ukx1ImMRT4wqMdrLOVGuwsyyvY
+b+KmxsW2WgFwrnyPadTKEyZyv9EA76+MUyLmiBC1KNGJc+o+0kQW85ankn+0DX4Ps7ukZWo948t
XN3A3BLpfiHIYl9q3JHD1AWdp6lAsVCKjwpldnp4LoqRziFukdAp4sg5XjwRUfr8uodCXlC0gVdQ
rkvzgAEQR1EAeSFL7xPZ+iLCKXev32+Twrd53EFRHWEMGuynBf4iFCt3P05HqHVq2uW/q+FlIwwH
ZbytyW5UqPkzVSEuVgQHecxEfSWAumRTwEtPfIsVlCe++JuElg5UWJBQAfEHtes6PDdUlrWFtzeA
+ReYv2U7FjelkRhkwYPGDtSmcf95s0rqwGbkq5Njh5xrOYKbkSf3laU4PTFk0G95+8AmnZa2zlFQ
T3Rs8GijIFLqOpnUjIUquPWwZyyQ9/x7Kg+yut98eNbwUYMd5kC0UW3s/gz+8WejIQgYzgD90pyq
UovaeeRojDQlPfm6n47mLW9sqE0SZsmfKpIEQAPTY/rb46jvmXRD7eitJ3vkEvg8dqYmgfcZkDKP
wl7P2rqxx9tZQ2cjj7pOH3DEFFoJ37mnfe2P2nT+Ff5xckgJ7Q0MbTuyYiBn+hRBoOLCD1FODpOd
gpYgCwblqSQdD5lnTrzsb6tdEid75DzdaChJCnOc+6mqaRU4QpGokDeBZJeyV1Cb7escU91EDOI1
W8KMu7R7w+TlU5wq5xjlbB3lbvajT2+zK2p31z0zsEplO3cqpOxjuB+xpfkTeAcWtx3aWjGqnKv8
r1UKZPvh8Hs8MpWIYfPdHqohjlE/WSLOSfKz+Q+GyjHWVubE5uAhut3FrvX9Rg+09DW2BpEwBnX0
htKVIarLshT1h6BJ/w+3MCLuB9Ojw/R8loQHT5pZFSvpDrGzyiPPQZf1YHo2xVm19NZkPCwLNG4H
6iaDud++UVUqUqbAwGkJ02eVWd54OMiKCv0C1TuixL+D9r4cqg8HDu1rjlwYnmjV8JghRPYKILC6
H6dn0Ms7cnS0pop4QR79IS08XsATZGEnNevv84Dm9EeR5W9twGuIDnGDZmVVlDeDzfDtmJuGxFoi
6XIhowcUn+kfebLApu+t+/+H9R8gdWTopnnUTncuXdKBrnN3ALN+iDf2RF6sOC3IycnenB3KXP1g
P5Jmv9OjUVVPTUjKefEe+HXAd4ING1pR8NmffjPzruyo6MMRowtyKayHP4y8R97ba0juwb5ek6B9
o5Cco9X4cSJ6FauLDcHO7yYQZRKrV3k5Y0oj2bq+xizG3qZ9vhm0fH5ApD4dJ7pNpXiVkNyyYef4
O1WyECrprqUa2f5VWHnrbMLFs47afo7NwEObmgZcq3DcDoYAUoLea4YpOXOCcLRcLK9N5LsQd7VY
U7LdGyNr5T02v9lA/PQqC/BS+vw7U4E5O5lrhhgIjjVT2Y7WqQabNaT1vMxi1qrF7kQLfbfPAuhE
ypx+NKMbS88iVMXx3mjpcpcdk1ASYFUkFB3nRSB7P8K8nfBzOFso02VH+A8BeD0dbcQJ58A+u9rY
9z9Pz9RgHlF/WNk6moV8rvhdKz6eXnROm8L0eBW2+HrXlfYZlgwR7PLr6HT+v3S32yeqo4jv8eOU
FKJfU8rmz5XDqHoOnZBxYMY5/jPoxG7SsUdVP90rFrqnqBP7d3x4SKQJKM9QNxcheBCrUCj7CACN
5atZC+XpgOFcr/Nz8ym5qEWGzvYqUzTchbtn6yRcI9Lvx/kwS1c6Vqcmf+UEYVfjTo5bnOvy5E3H
oj5hNFKwGibNm5fPYVRf8xDpkRwnKJP+2vm/i8jBPuU8mlXPNaKXbY29mDt7dIH7txgt1Y8fo8NH
R0S9LLgezHeG0g10VNiW3OxhfKCU6TIYwueooRyikn61TmYOILHV/kYzeCoHfGdbVawBkUQRlTbi
u4nE3mrIu+Ejai0Lzo8r1GhLFPT1mtyZSOKd8iq2HinAz0IoNXC3TWXpTGKdby52ZhqkIg5hkTG/
RVNLYGYKLkuT5SGBGUKh/QOJXRD35Ak84yMAAtlHrlxhvd9wZfS0RUYq/WZL+MasLpaEvZSY3teJ
1OyXMogs5BqOFXkhPVEIVF1Fc6ztxB3BO1/jqXK4bUD8kCi7p2t6WprRHTetURjQEdufsgw4dXp3
Di4eOrtKn6+GQttDcRltGM8hIT4sGH0nCR0waND5w8bUaUf9VfYswxZMkR9RK5YNus+IFF2zA5db
Aie6CyfXxUY44mte3piDoSBKQIYIzeZRDJJSMIezOwo4UPsR8sbie1BzY0ejIZYkB3nqZngvfxfw
6WhuBine37hhdHPkGOH3S46Kh1BcYppv2sO4i8jTnGOHw7dfW7UmqdBQZpFEOfiHcNhsnEynGiDR
5Y60HIyKMaPiQd3NmfHPBoVyPhbThYR6ZVqHRzkPI+Bubrg6HX1d7GxgJO3miD5+rk4PL/r1WwMX
OubyVgy0YqwppxkCqxXxetTaezLvIjIE/vjzsiFDZa6yfDdrPyM8qYHLs1akAhi9vtLu45GYIIqi
R3aR+oidmwzMNFP8DeOwzmRKQZikCb6E9LV6AfPyQs6tY83Ld8LsIt+HkPF4k2EPUAlX7OLi+J7x
TYvMXWl/XK2s/1iEBVL9QNbxOn5PY/LzwOHJJ6navA==
`protect end_protected
