XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l���Ͽ��F���7����,��m��i�gM��T��ۂ��<_�B
(�iOK��˕�N�;i��r*]]W�17E��!<Jc��%.��ڰ?���T����`��t��ↁִ��c�]��]Z�#W{�L���Yj���?� _�j�$9:�5(��-�Q@fp�'~W������:��_�S�C$��Y-����GaT4ƞ�l��E;��Nu�1�M���-)�2�h��3�v���.%���"�]����y;�%����})RL��Z�eԭ<Y��[4��^fōP��s��t�[.�l�=���� �饩9�U"��(�nC���	�D��6��̗;��E�њ
�C@e��-.����/��� BC��sZ5�W�����"3n�$���J�W��:R2�
g���s!�7�v�����8h.#Q�nJ����.p��t:�70Q�ڃ����O�}��r�9~ѩ�em\���c��  (%�zn��C� _��\d�H���	�t�@�ג<��a���7���]6�#R^i�=�'�����?���eT�����k����!�oYd�>�ܣ�s�f�no���4���7K"��:� ;���HL$����l�s�=���'˺ZK���^�*hdIX?�ag��wP�'DUjLr�k%5h%�W�A9�����uFe���I�l�x{O��e�p+�-Wy�|���ؽ�������h�'_��BQE9���_�dQ��1�(&�����.��L��HS�XlxVHYEB     400     220���<���US��Yz��'��Zg�sԔ�J�[�L�z��-$)�G������2���4���z�c}s��IwF*Z��Z�]�+��R�0JM�<v��.NΗ&c�+�'�#�@fo`�π���܈d#��C=�p��<����oq�]�*dЬ�1�qr���|E��c%��R մ��WW�¬j�FA����_��a�.�A�1�
Yi�ih!h���!��/�UƏ��+�H#��f�xG}����I 8��b���Y�sꫥ�t�Xf�Sh#�(���Zpk1���B:��X�� ��V�1�i�SND��G��%`�0�� ���M}���]�Y������+-poCUэsMs���l��G�G�u�x)�tC0����S�.����m��Z� k�g�\�ƚ���k�A8�+fD�c=��h�w7�-P,x<���=��Xlk4pFe�?���#Ŕ-=�,n T��P��p���s5��u�iw�=Oz�˖+��M����H��d�VE|������J�+�#k�LgU�e�5b��w�XlxVHYEB     400     220`���T��+4("��rR�I��W/����g�^Dႝ�;%��g�b.��M5�O���
�Bn��p� ?0���P:;F܊��x���F����4��=`p#4���<�@�0��J��Ǟ�^���ҙ�~�����*l��@�&�K����baa����$�?�=�7�� �ӟkz㵄z
��^K:f
�U�x������d��7�ɑG���p�*���,6G���˰=�^�{�wAx+#�j�!�w�5F��4��SY���[ �ێ�C'�+�[�l�sx9�J��V|������U��`}��Σ���B �B�V5\����^2Z���讜��m:�T���c��O���7>��~v��@�-�0���,���70G^G�T1I� [G��(ꋋo?TI�w�~�.��Gs�}��~��aӄ��Ի[r�{�0fM��pj�V��gX�
���X����5��OHd��{�fXp�h��I�;��1K��}�+�H7�B��%w�7'���N�(�mk����N�i��U|2�h������I���׍f!>�.XlxVHYEB     400     1a0�������������Q�|�hWi��/�>�v�l*'!�-n���3M�%�u\���2�.B�ih#��g5b�3i'���X�ӴE�Q;�gT�#<�B�NfbH�dq_�ef� �5��~�T�G� r�v:o�cI�yxnH��}M�꧕2u�E��:�+�J��ذ.��{�0���z�-,ޣ��F;2����ޢ�E@!��IM�@����.[2�8�^���!�"���7���2]T�WU����p-(�F�ȏd�Ԡ;B�p#��P�}�gX�
�4�j�s5sC�K��7����9�Ơ!᯳�.�W�ԍU�����*�g����蚲a���G�Op��V���0���ʨ��8N�Z\�^4��O7��.�"Ǥ���䵧.x,��s={n{@Ŗ=�_aj��.�r����.XlxVHYEB     400     130�~�NT�A�|�5�t��W`�E{:9�=�1h�j_�0����D�a��s�@fWX�R�pR2���%1~V�����a�$vdd��_��38Iu[Ksو�(hudcX�a����-�93�Oyb�r�dԖ|"�~+��Hrث���x�zBX�{P@�6Qw���8�OX�B3�'���n�ʕ��~p~�fG4
0����K�d���� gl�Ω�#ض���E�a�bG@�+�����3	�2vͺ_�_vNʰ���ZJ�;��ʽ�Z��^

|����5�]6I	'8��-�jڻAM���XlxVHYEB     400     140���:Xx��N$%��Ύ���e��V�	(ê�x���*��Z��dqy$~�?j�t.�"n.v���x-+�����e2Um�1$˅�>��N�[/1�6�u�X��<��k�86�a)�9f�l�s:�$mY���>�5����̢�\���e/ťh����?;����/ƺ���N�c����}��wr�	�9�\�&Oe�]PX"�"���фp`����r��#V�%Ɵ�<rT-'.aJR�:P��Mע�xp�sf��OR�?7C�\^�J	
x�������Xj����:��v,8�\ナ���W6�6�I[����XlxVHYEB     400     1c0-5$��)D�`�gȔ}��b��{� �/K1'6�?��0m�T��E�T�<~+O�X�.�^e�>?Ķʦ���Y���(�TakDbc�`���c�?��^�I����l�S]��������fW����z��6c�OX� o5���G� �|�҅`�nyx�9�4\-8 o���Q�H���@_������Dx:$#:�s^!+�!$/r���@�����X{���ȃ��+\C��=�3;.�oMNU�5�jV���\MuJW�����%~��Q����}#ni�j5w��Λ��1@�B��s]�~"8-ː�jG���)*ݢ�(Zi�]�{�����cET��Lő�~��ۓ�1���Wf�
�^u'*�4c�x(���a���ɀt����O�,Г�hؠ�<�q�/М�Zv*���ರ�s��vPP��d(10W�엹�=�H�����M3&�G��{_jXlxVHYEB     400     200��b䄵�M��nZH��K��\!G�*�8��P��j�,̎�iK�Q��_�G�o��7��%h��ئ�ق<�X+�x�7O8�ocn%+~�u��s\��MH�ִ�J���(�wU�|n��}1�i��LL��C �
����V=�{����!�f[�O#��d����GfNW��ǟ
W�6�_`b!���a�\"	����Y�h#�`�����bQ8������3Ha�����g�p͒��݂�"䬸)[��J�A��g���S6' ܩmⳇ�2����@��W������֤0�3<�r��\�M6"�Ʈr־J4 #O�b&ڿ���L��!-ג�?�A�C
��W!/o���7#{|>��Q���(��X>[��?NI6�3���M7��"��ҳD&o��2{g�	��[����`Ǿ~roc��7}��.B�߈�-���/�Q��,i���5V�<x�?i��=w�]��G��-��/��2�pTaD�XlxVHYEB     400     1f0<q�H�����et~�f@}�j���;�(�|z��֒�o9����iuBd�q���2���!Ȝ�k���<r6hJ.�H�e<s���u���x���p|-�rA�!jE
���N�����]dݤ�U	�	��ۢI>�]�E���ih&ا�������ٛ���e�� 7ل��S��Km\��bܦ@ƃ��"�0 �Ȏ>��U���R�
��M^K���T�׏^��s
�M:��06���y!��	�>X������q�ߠ�O�XH�����d�h���nV?�M��}x1&�k��Gx�C�)t��U�jx7��me_�xFf��Dâ�����n�fj��!"?���ۂ3y�Aj�
�<W�ub���զ��9 ��#p���.6�f��l	Xx3�t�$��wW��o�%)
��BSfo�>[s��56V���Hj��܍����KX-�j��T�2�.�K��m���-���t_���!�r|&%��YQ�������XlxVHYEB     400     1e0�����ߴ�yȊz2��z6�T�@/���S�:7�;�Ӧ�-.q�-;T�gd_-d>r=�J=y�}R��τj���=��rwd� 
Ş�Y�I���[,X�Q>�����[b ��_��&���p:�9���Y�Z� �-���'�n{%'�XFҙ;~���G���/�������bC�Y��Tt���,,������,���4��/P=ô�����V3�����S��@{�d�gs�u���<�܇�1��5�8��P�,4��.�U� )���Bpx�Q}8��ilg���v����b�>�)Twf4�	v���N�g�U�5U�`�No@gdu^�.d��tV���r]�Z8�<�џR;���|��ߠS��~���>��1���]������8¥�bL�} _�����:{t]pz�\߁C�[Ϥ����s4�w�;��42����A�SO�K�Y�g��	��������XlxVHYEB     400     1c0_�U�K�~��3���q���2� A#\'s�D�k���,�y�����|�!��v:�;]k��e�^]B�6�(�l�bu��m(�1pE�Ϥ'��b'k�� Ŀ�.����(�&���L�˄S�4%3�.��qNo�J�ܱ���Ӟ�xe��+��8�R@��=tS̫}�����oR�PKXL�
#�H���.|9��˓�s@��Ǩe�P��Û��XW���/�;�؏+B�Z@(��]����4zR\-&f�߰��"�߫i��
<��%���/vh��� �>��ˋG������m-��QK&n��G��:^��³롘�6��)A�����=$8tEu��1���[�x�k��u0uuh�IJ��C�B��W�X���BڔY��89�MZD��֦��O,wc��x��f����HTy�>ѵEh	D�oT�~`�Eߟ�XlxVHYEB     400     130������c����@2���a��nW}HP��
~���CL�I\�a��܂5=��iJ�ww
�x��j�c^V�&e���J���M��Rg��8����ߎk���\�а�.�p�� .q'��p���L�A�-��;��P[t)@��UĊ��]���R��)�:�kM�\��Fw	r�]�,��~�T�		"�66��]�9S����׾��sĄN0<�zI�p-kN&�q^=<���w�9�ʒ$!xt������Q� �"�Z�g+��g�Ä0x����)U�'3�*�8�rg���U�5�8��XlxVHYEB     400     170��ĚOnn'��٬-D&j���1E�����i��r���u�=�T��.w`��_��Q����꾷Ǚ8�h:|.m$!�~�q<��L�bo5L眱.N�6�E]�8�RT�R1{+{cK�Oq0&��U��e;
��|cX{�BCo�@��˦��Qg]��N辎�:�|�3J#T;��a�������+�i�������#�GNZ�Q��⒝���7?�i&D���0u��^:���U���y6���	��.C5�,��a��Tb
{F`����E=��>y" �ПR
� c]�V!���<Q#h0����-J�h��vm�O<�%�}�Iu��c^S&<rѸ������s K`O|m�p#'N�XlxVHYEB     400     110�
�3�_{��^��v�5s�_�M�:�N���
�\���`��"�}��;\�_�:�.�H2��H��K�Z�#��	���pPW(��B�_S�� ���q9��A�}Z�4��mQ�ϥeձ��%5�LŢUf�V��e�m*�j��BZs�-��GfHC��m�BN� |�yV�:�R@&qî�)m�ع��V��Z�y��h�n�r���?�KC��o����D�x���(�w6)��̋�d�&��K�^�l��2$�Ilw����;��ތF�S��^XlxVHYEB     400     140]#���ģ�p����3X°�r��p��sa��� ��f.��j¨��E�M��4[	�?3�唹�N�y��*��ЈZ���K�-�V��7ա�j���h6m؍_���MY�y��)7<t�j����˷���2I����'q�X��R�a!�2h!��=r�l�������]O�E��J�R��-C���V��cRU�P8��4"�e�b��W|�C�!\�ix���w,&�����{�a:Y�X���V�b�6���҃Ym��n+jhU%�J�!R6�>��!���;o��g������0����_��R8�LԢV*XlxVHYEB     400     130��N)�WC��k/�]�l7^�tMƨÇ��4KO��E=�&����a�ȲJr-�WՀdW�~�m2��||ט��h�髧z_�r_����6�49A���P[��s㪘?'�~^���g�^�W�R�% }DL�8��ag��
��\7A��y�z���6�z���Bh��m�ᩯQX�~�ґL����,&�(�M
��������J�Lh)���q�\G�ph1=ؕ�;�?ń�����Z7�����]+���b~��o�?��p�Ol�FDh0�66+�JK�r����<R3Y�XlxVHYEB     400     1309�˸>V�����[�����t�LdKg�^�DJh�ƙWl5�n��J2o_Uw~>�=V���<ǠZ�ў��� ;Zr����D ?���-����w�jZ4(/qG-腄�\a\���"��W_��Gy�%6�3����@�Q<��U����ܫN��4-Po��z��sʈ�"0�F
��:tKɆ�6}�n 4]��c�"�Of�r��"�]�CMX�x������, C��$+���щK��P@��?d��a�w'{~�Β�6<�&d"?$�<#�ͬ�Nџ��4�_l�x�8u�/&XlxVHYEB     400     150�rO�[6��#�lMsJ��ߗ;"�Q�'�ܞ������ьŧ3��o����g���Y:�k��ǎ^����D`+�X�����;p�#9k��4�+�]��0T�}��Nk"�о�����>����k�P�G�q`���r�b���P[�v�Ρ������Všk��f�&�E���1�,�������aG���#~+��|�WP��@���-�ߋ�5���*�v%�K���zεh��&-�ȥڥ��|�-}�0R���β�cg~��r�����Y��r$=�݂�f�������+� ZA��9�ā���2�u3�H��M�o�k��QF�L^���XlxVHYEB     400     180َu�ic=���3�b0�%^j� =���O��K�0/\��p���b��GXU���T_PO� D�́�t՝��ӈ�Z�
4N+aˀ�=>�v�!���ׅ��Ry�V�~w���I��`|����	�>l�RӬ�������g����Im�Ahc��'��R|�sI�l9_E&Pi?��|��yCg��ы["qh�5��B�<�L�-�b�f�_Z���%L�?NC�a	��6;�̓���Y�uN` �~�,P��F��i�!Q�o*��TAC!Z.@ղX������+
 fS���'S��s�]߽ˆ��;�?ˈǼ �L�&`�YȽr5�4�Fӓ�Cz�����<!���=���h˾q�S�R%�I2o� ��;KU��mXQXlxVHYEB     400     1d0o��b�wJQԔʽ�r'@	AüR����^ݧ����`0P��ϟo�S>-�GǄx�eb��xe���0����9L���b���qm�F
����7�[Mqr{��_s�J������Q�Ż'r*,[۾��	���C�`��A͸�"�{`�^��`��]g� ?��"Re>]��R=r��g"tu�)yy��%�oB�m��*��k` s��Yί4�m�i۱�����oi{����l��l��@L6���լ9��8�ˤ�B�e�:����}Os���J��1KZ�d�����ᢓX���?��Y4����Y�����7�����J���Ϡ����x�j�'�t�J�#��iZ*
�`0�'����$�Lk�Ǉ@G��	C����_�BM��[9d�RL_K$�5�ž�Y��jAM	^xe���ϐJ0���R8.�Z�L��uiܺ�sXH�tM,��4�>YI�;XlxVHYEB     400     180nCK.5�ׯ-����U�!��� <H>���؆U�u���m�U��K���[�GM���q��<9�%��`X��G��YG<��u�hyS�F��'��_�yD��o >�m4�!e��J��pAi���4|�����F=]^?�+��T�r�o"��w��eI�J�mM��r��ҽKocQlD.Eє#L���{>�ǖ�g�*�`&�����fF}��@Zy��a�Atא�x����$�<�n�O_�����L����kE�ǒ��7ˢ�����m\�txO�?\!V�0��8(���C�.B}D���罳 ��Mh��J��Q��1�>���,p���:�{�z�{;F2�x��8o�5�R�fO̹��a��W���.�C/�XlxVHYEB     400     150�[U����$���6�M9\���=ޘ�0.y1��N��kF2[��D��	}�F7}���Jǯ�is�=S�&W�- ��`���9�������A��e��8�+X E1<���F�2P��cA�1����*Q,��q���M����|�Hj�l�q�93Qi6�ZA�5�\�Ω6c�YG���$��U��ppL�$$�H�cFt�]�k��_�T�sECji;�>�qj#ޟ��N�+���n*(���ꘆU���f���SO-��t���Q���M7��
���
��)9s�M1��%��?X?nc�D̓�5%}S?l��(����<#^<���XlxVHYEB     400     1f0\�Ҩ�J{���<_�=�Ԭ�->�z`�/R5�%�f��.�kn�5���PQJë�=�WM.��O���z
����f}�����
$
��ظ��C~y=�OϗH�y1�2����G?�KlX�'�vg�����wGU�4�^��o�]�qm�g�ӈm��фӈ��tn�ތ�^�эHOv8#l�G�#;i� "���������@�ګw�<k��A�M�������ir\Se ��M_�̹�j��ϯ�|V��U�ϏI��]4Hσ���ӰМ��	���d�*��ЁE��h��+�l�P#�4UnM>R�<�]Udj�t���� vY�@u*"Rh�������V�o;I��>�����FHE~��5H�L��e ΃B������-K}�W�h�>�ҡU'��A;�|�-��9��\��1sG�bz+��&qܳ�P%E�]HOaww�EK?XZC�i����[�o�N���6�2]`���XlxVHYEB     400     190����|�J8�Iֿ��������8��s���������gN�B�7	����q�Vn���
((��Ɨ}���]�ED�S�����"�tS��ԃ��:FmӔK�6�>z �wp��-JݝKWl���F�����qI��@Z���-�_i����2�D�1���B-V�c]Z��y���+�s��yo	8N0����	e�?=���Lī�c|8��͈4=������Q��KgMg�f�ώxC��2b]�ӢJ�;����w�6-���0�xɲ��߳Qi-S��]�W�1���R����C2��w6�,#��R��D�"���{��y;,t�Ǳ�T���u.����]�h��{')�����f��TNs��c��~^]$c<�#�S7��y�6�XlxVHYEB     400     170�&�p��M}4%��3����� �'�CT��Q}G\�"���%瓢���Ob�#E�W+ypY̛��;�$D��5�|��`��u�mX+�����R�Am8s��r��+�Kpv�:�^
mF5���q��X$�X��z��;�T1[��������k��e�w�������W���e���@E�����[ 8>N5���4S�uq���%jbs�g�=�VrFݸ+f��n�����!�|��KUԘ����s�Qʻf�O�����PQ5X�<��:���<�����x (���ע��E���X�iun�S����S������+PbG4�~Mq6{)r���j�_>?5ٍ9:�a�,dCg��XlxVHYEB     400     170�B���Z��c&�m�g|ŀ�ۼ���TO.=_d4�����X;#h=&����~/=Ţ����2ooV�s!��/��6C%	��1Ճ�����H�"-[LBy�8�x�t�����>`����櫭u����e����^�_���r�|��~UQ�K�x���՜��R���K���H!s��ٿ~�O.��.�g*h.���E�I)��dt�Z����_[�b�+7rܜRT�����V p��
FW��Y�&v���ax)v��#V^��&�3�����#�Z�©��+JKa_���:̙��R������9VM8o��`�B�CL]��T[E!5l��~�m%��qV��� ��I�]4%wRXlxVHYEB     400     110C�<��e�3%����·�x�+UE��j���؟��
Z�$uR���<y��p��h/Ǫ2�t
�'@�fq�G�����O����E��T+N�~Ԕ4�|���H����܋��ΦS�s�4�\eD|`�v�!T�e�"AAݗ�䮲���=��y9��%w#�4�kKQN%�|�̮�$5[�	\��)M�m-�j�TO��G�m�ŧM�u&`��07�SL?N�j�����)x�]��A�"�����d����"M���|��XlxVHYEB     400     120	ۂ#s:۔
o�Y(��{��vC�xb���K߅��]��R������*��ov%N���o˹��W�G��x��zF0>k�p�&�������&�&���Mkѡ�A%䳉���t&��&�c�� ֲ�۳c@^il�e�J�wf2��g:��<KD���"�O��&�a9���[WP2���� "L'������mb�V}7R�b�{?�yN����=�������Z5�q��r<�9�h��a����6��z��4KF� �lG8�p���w���z��N��66<�#�%�XlxVHYEB     400      d0ӳ)���a�L̖�i]��oP���4I���$�7qm�I8Q�.�V���r3�z'�՛�L8����|��Sg"��=�y�,�/��r��
k3
Tŉ6�r"J��^��~w�h�j�����]�0e���=�k�;��M>�U0L�8ƙ�7#_(�����;6te��:�%>��� ���j wuQ-�i�9D��c$�%i�����aW�5�&��TXlxVHYEB     400     140��!g�"X���1q�y�|�"$�dK��,]̣�~�(p7~�mU�7�"�&\��bg��=�}���jk�al,uXȌ�[ˎ���#FS6�B�L[��E+ت��,���Ho�����D}�*�]�Fzp��lk�E�����1K�y�<������k}�*aͤJ�Y�ѣ����f| ?�O�ʩ�hk�ӭ<C�9t%���Fe��J>%��@�f&��0�U�i���WE�^9L�-X/I®+q��X*��&c�N�%\�O��y���q'�Pp*o�����#��l���)�Y|y�����#�h 
��XlxVHYEB     400     140�#����g`z�k}��Sĸ�/�G2����
o3w즁A�;�ZW�ɒ|���:�+�X4[�+�3�ܔ���cjŜ)@��@L�^OV�<���usZ���8xAi����5'�� �����A�����6(�A|9�ֻ!���zb�
�u҆�A��C,��j?Q���Γ=�S�@�'�����v�d�W|�g�s >��Sz&p;?��5�z�њJ��ug�� $��ȷ���|(;2�hc
�,�-����#\��� s=r� �Z���Md��'!�:4<�t�j9d�_�$��4'ͣ$�Lwp�f.�<��XlxVHYEB     400     120���N�"qnt�^�׸K���S!��G�M~3;tOV�It�s� ����;�n��|����R��?��]U��^���y�-^��WU1`i�6,@�Ua�:
�
����&���{�T�e�aB�Ӷ>�&�UVkH��"PI&�ݱ#�����TU[�33|��	b+��w���?�@�/��3���j"R�Z� )@V�OÁ�4�s�j�	i�.ԗ������M�	d�[z敎�x&�C��*_��������P~������¦� ��d��of
[��;ji=/���XlxVHYEB     400     1a0��ifhv`�yLEv��x�1)��X��.�m`���=4,�B]����� H��m��E0G"����6�.K��� K��/;��?u|ƒ�xn����9��ջ�z����'����Vq��Q'��(��^>P~�	[u"![���6��ޙ'��b"��l	�_�9����oa"C+���B%'�h৲���ٝ���څp�OA~��f�� �Q�z���� E�����Qx����B����ہQ��; �i g1���2|���\�e��K���gD=����>�o�g��5�e��"�F��	�ȹgn�{�<z�"[�g��$���5�³��BN~@l��n-\.*��y�c�˺���l�m��t�Il���ζ�ưL�����A�N+?0/�b��t�XlxVHYEB     400     120RR���� ���Qڇ@�؂����Y�f"�ޯ;�y�� ���������Ŕڲ6j��)xn­Y���ԎשRu�p�Ə�F��@h��
��'�kE�4,$��ܷ2����r(���evq"?�D��l�.$G<v��H�p�C3Q4�.����X��¨1�`�4Rj�Tf�y���/��mz���)����+pfӧ��ƆW�U�{���m�ת��g\Y�U��B-!\�������/��4�Ώ����	g��hƙ�cݍ�<x�Wvɛ29�SXlxVHYEB     400     180�ҹ&�i���m1�����a�����^��A��̄B�4��b�@����\� �)Yt}�bO^AV?��&�mt\m�4�M����f)NK��j�G(P�96|�ȣ��(]�"�H���ܺIb(�����?Lyip!?`�4�Mm��%����8"��|��"5EL��y@�%�j�ԚNv#5,�zY�wڬM����D$4��ڨA�;���eMH����Z�,`?�4�+qJ�A)A 	�tj�~G�Z���>�����4{뒀��#C��^�
W�*5���jc�����[���q:�1���R?/��(��o߷ο��ֳ7��RY|�~�C6ꦟ�a{Y# o$�I2g�$�m�;�>��ؖ�ϟ�4M�&XX���f�XlxVHYEB     400     170�n?NNl�O�N�J�+}�f[d��̷��MX���<�z���q5b��0�	�R���π㸢�L�!�}�O�;�`gh�1a��k�0� \�v�n:�����ژ�������_M���*�-d�ږ.�I�`!���7����f͉��T�m����k�9������<3t�+SE�#E	�9�����3T��Q\�� ���2w��X��#�'º'�[+���x?2E��p1C�Yg��k|���X�ȳ�C1��Sx�7�#r�q�?��UDTZ��.�^ObN&�n[�����4!�;2�l|M2�kyw���*"�O/�l9	L� ���.~	&z/�wJ: ��W��hU�8�����|XlxVHYEB     400     1c0)�I�rE��|�,r�R��s�.b|I_��*˝,�dGl 5[��!U��R�Өa���ul��*�NF:v�*���Q&w��b�s�+WטH��p���p�vH����[X�X���:�2g@�����l�>ż�]�O׾�%]?����F�'_���w��иOfY]J�Ō�ݫt!�g��!�W�k����g�bi0�յeqk��*7�o:	������^.��k�~���b=W�d�$�l���8D���3) t��'{��k�BX���>1n9l̙�m	ݱ,�ȚP	$P�zfB�4�� �C��1H�b�tE�"���߫��*�R���,T��;{����[��OJ�Eg��pM�(P�&,�F<TbOkX�Z�Fe���D�F�Q�F���M�
t�>Ŧ��Ov���
^���Se�7�1�L��uf&O���(��[��LXlxVHYEB     400     1108��e~N:��e&~���n��#��D�}��g*Y�p�3�y�,���V�E��\P�0��G�����B]3��:G����v��L���&����`r'јJ�̛0�f��Lg�ˣh:���98Y�M$��-�%L�9\TĬh%6Yq�OEEP��|�(�6�n��������p
ǹ�K������x��ѣ�|�5��s ��!�tuѲX�P˭��sx�.�����9Ξh��g��}ί*��B47~M���; `XlxVHYEB     400     170w��N�p++hA�)H���~r`�$��b�<�8��)bzL]Ì�����Cω ���/�	���!y�����N?��}����_Bs/����e-���\3N���0g��
��L��7�M�{k�������#?�� ѷ���2Z��z�%:N�!�l�s��d�-v�����8�a�����g����
�
%�/������p�|S=@��jk��j��R�U\>�^�C|���������+���@������o��s���3oog����Q�yR�G��ED��~�
>���x���S ���2gź̤�x�Qlw�0r�lfw�G��XӚ�][)�C�.V> ��^uo��0��քXlxVHYEB     400     170��,�"bS�6WE�3؅��Ni<��=�?����;�2�W"�o�E<��QH�A�k�pF[=n�S��Eh�K�6�S�_LjM��ނb�>a2h��>3F�氮����:[nsq1��5/dx���Sez�����r!�g���6Ⱦ-�n���x/��]���`!`���5M�l�����}1zo�l���(��dU=%�J��ߠTg���ד��[�9F��(������Ɠ�����\_}=�෰�i3���?\��D�?��v��@Z���7y EΙ f���Xy� �@<���+��9t�S<�:�^�r~�av����19�-�c�s������$�𞍞0��30O��u�����*��P���}�XlxVHYEB     400     190�P��~�d�������ю[�P��ɲTt>S�"
Cp.�B���wm�|Vͪ�mP��. ^M*E�_��L�̵��Lk��8,��4��Be���y^�=�iK�g�An^w:l�Չ���w��?����clb�})�`��������)D�n`��?�jl7���|�۱"�P��\;�c�;c�F�����������Ţ�xx�ۚ�q<��>�ZZtY4��ѿLB�$d�ZL�6���{�,��mN��O��^�����&��-�'�?�T=V��,�Q������k��������cz�~|�Q���_��㎔�k�
�H���v�=� �G�M���"���C��"tC���w���u"
�y�Ҽ/��;W�V�enW�0�fD�XlxVHYEB     400     1b0�� �d����y���~�cG��������g���s��P�5�w0�S�:�'���xͼ���
JJ�E�*OuqZW����q)NZ�s��o�l�73n��z{M�r.P�7W�Gz^���l; `�~�t���0�W.6�S��'m2�@G��\���6�KUg}��3�~�=�l`�(�1 ���"�$��M��:Vh,�DVy����s�.2��&��~U�jΏ]g^�ikL���XH�����XӁ@YWI1�
R�c��|�"Nu){�wYvb��=Y����lzn���P��ڽ?���n�;�_=#s�{��OJ��XD5����h��:k"���T5�{����3�3N<g�9��1��,�vۗd��*�/�����n���Ƥƀ?�
M\mA�	�5})7�x��+�xq\,]�XaXlxVHYEB     400     1b0{�#�igh�� �N���'8�:.cy��uXګz��8抎Uhj�מt��8���H�2k�D�q����^��^�����ܶ��v��.��zy�7W���%QO��C�Y'����_��X%�~��ך�~ ����p�u����j���E�� �������Q���(��e���xIQ�tU|A��v����������u�\��G�B�O;�[���\8���Cooq�5�Nr\��	�׺	���p��8��a�0X���[�F������N���|_&	=�A�l��f�8�d��~a��}��.�ӺJ,lⓉE��/�I��<->/��2�D�7���蔤��c�L.�k�ufn�¯ U�si�9'��W�@?^��IJ��;�X��0��;�bY]Ӏ�}zĘ�Ĳ?�'��ýl���H�ې�Z�fC�XlxVHYEB     400     1c0��.Ƅ��_�����@[p�Soԏ�@����|r��~-[�G��D~q)��@�!j��%.Pn�O\����\]$ևp�;�Ж��������[�d���l~*�.�Wv�(sS�rK$���n��. nc!TC�!�A 7u��D�G�r$�^X��ģt�F��=JY�B%�3�-%�P���vs�õ��݄~��6CM����y�a�9O30�	}��[���=y���ZĬ����A���g�����A0�0�K�=�c%�˜� j�9���I�E�����0��O��G4K%Uf]��MF���bǀR�˂�AB+(t(�X|y���K�E?L�'v��
�w��>_��O+���%�����b������ޔ��*a�|�� ^)�C�?C=��I̉`���st��x��q9;��ϝ�H�#������g�ަ��EXlxVHYEB     400     140��f��nwDͨw\%ZU��IdN:̣=;
�WL�2"���-KRDs�֪�4{���Cv�E/.�f����ȑ��1K!��#Uv#��#���+��5BE�Q������u���w�K
�uNu�g +�����L�>��,U����|WJCGXb.�F0��p��>�ITm� �֌��`4�T��R[���i^oE� �{��T�+�R���<��|�5�(��ee�ll��<�&��C9�w�0�!p�klm�X�/U,�e�W|�՟^�~����^���׽)���=A��R[Eqy��_���)e��, �K�XlxVHYEB     400     190s9��R�×�1�7)b�u!Od�"����96���M��2*&.��H���g��k(I��Q&���D[P�_,F�L1}�']�R�2�(��H���� ���*k%��ϓS����N+H���e8��ō� ��/�$��f"!�	kAM���qi�i�$�9� Q 7FO8���jj�-�Z�K5��4��D@V��V§��s�u ��Q�8)�q_(X�UN�#�c��ɠ> �8S�~Q�k.t� �)��������`�[�uT.�Ϫ�z������ޝ�;�8��0�e��x��?��h�U�jQ0
�~J��m2!�l&�;����x�W�J�or�9߰�\��X:"�D�+T��^��q�D�VFyc]T�Ķ�oa�hcJ+��.źo�(�FXlxVHYEB     400     130�Ǆ۫*fRn\9����A�����c�뿟a�:Fr#=�\Y�\��zg����J};��q.K!d�	o���.���PErz�)~ ��(��"x��B����	vj���(���G���v37�Z^��$u"lq�L��\}���.=n�/����k��-������c�&��m�r�d҄���_!��tT�� 1#�\b�%�6�?-.�I�}�7k^/��t{���i�ߒ�-r�A+!�:�3#mM'cd���u2��80�c�t�t�'�l5�� t��T�>���thN��XlxVHYEB     400     150w�"�M$�tOe�Ɖ0�>G��}<���r��b��?吲ѩ��ڻ�I�=�a�tռ^�.���x�b���w�j0��q8�G��0��"����e��b=����0�7�+p���R#��^�{����A��QE��F�H����/B����Q��&vz
I���TY, s�����F���ˁJ�m	М*�"����/��H�%ah��� o���[����"!�4��ݏ�[���K�|)-��/���eU�CD&�V{���~⛖sl�n��bz�k׈pǞ��x�;��	����o]�F��UE%����]1�H����4n�kƂ�y�9kњc�Y�XlxVHYEB     400     190�0d�y��^)�ֱ�n���
��#>�
�1dtZݯ�"��g��ɸ~�[;�w7b�['���g�0��r���%5V�!q�Z��H�-��d�W�=kb��۾b�ǽ0�����Y�=.�mD���|R��Qh
M%�Iժݙ?��&0�`��;ψhޅ B�>��d��+QX�C*��ͣŝo�#@H�7�;�X���J��oԨ�;3��]����497�%�%R�q�}|y����LCf"�0?xTI�e��G��%���M�$�B�9�R��K�Pw�.�?�����R�1)�wX0)}\�>eLO	�I}ϧ ,;�e^}�?�ѿ�Ki��~`zI���g��cϥ#�5�Ɇ$�Z8<r�tϡ���d�Y�,y|<9}J�J%OI�y�!�XlxVHYEB     400     1303#m��˪�^���0�z�����W��\J�s�㚾�fE.�����3�Z��ã�И1baM���d�d.&g�����3�e�C�?īί���(��T&��	D��խ����N.����օ�O��/��}BG��y�0)8u�3�9c�"?,,B��g ��0|���/S1+�MI��qEE���L�=	��p�@n,����J�y.l�Bd�%�����!���{tp鍓X�9�a�6�5��ʷe�cFH��CN�ȫ��Y�L`/?�LB���$����#7�?�c�)�����#kXlxVHYEB     400     150�|�q��m4-B\ë��x/���Λ��� I=*�p&�zbw��0���ե�<5���=��,�v��gqi�r�/�'�(RyF52��a�U�a���E�@�j�>m�*%n>*�]��V>4k'<6��<��F�;��>WB�����m&}I?���\i΃C���_3�Q�|a���2R#�����c�ك7�ymw��=G~:�]�L��O�i��Tt1�˖5 '�2|A�Jt�)��]��)�^�z�*����K	��^��/����s�r��k�zt�:�暖0LU($��*|;&��|�ovC��Ę`�
~9��I� `��ƃ|v�p$��}�I2XlxVHYEB     400     1b0�b\\���?�i��A�jJo���y�,(���O�o��~$`]3���gYEhˌ��к�"�	�^�C�kJ�d�����tQVz@0U��Ƀ �)*��n��tЯAR]D0{�1w�l��=�e��6�Śr�O�ܴR���)d D,��-�"��R 9a�T5�r�O�~�,��o�Zu�g�v�17�z�>W�y
�JԀgj��a�@( ;��*}�M��"M�Q�����Ō�'z�X��0�~(Mq��1��N��?uXm%ߧ����ҭ�hR�p��X�0h�6������[�ԋhe݁q�ǃo��}ǉ������Hͦ��h؄qA3��ݐF��p�9+ߛ��RغTx)0w�������G�!��׽�.���5)��c[��>��ש�֡^�Av�OX�1��0�(Z��e.$D ���՝&XlxVHYEB     400     1b05r�.��hE:��t�"媅n�EJ����R�����'Gƶ���~#�];,����
�NUA7�̉��l���"|�4y�ިAԳf�?�7Z���H���9��PN[��L�#"��ܞ��w������Xn��Bo�x��3���e]&秏�$T�	�0O�l2Q��
���F�R< ���71�;0A΃�٭��~��-�M���Β����E?�&�Í�@�,Q_7�Um�+B P��-O�u�6��r?���'oc��^��K�L-�������,v�r��+�TBӑ��5��]Y�GNl�+AD{��|�q����8U���`a{<~;J���O��=f]4
�r������A@��a��Â��N��Wː<�*f�ѵ��i���ⷍ����^+>���0�(�$��6uTOg����OCoXlxVHYEB     400     170����96X�.�`,K��k�!�1ِPfy̽sb����xa��@�%p��Gn~~Cg�o}~�J�\���?�~P4U`��o�����R}h�qކσ�
\}
:�2�088�[^�<Dk�9+%� 
lЏ�g�0J`Ņ���F�;�[c�ޞk�-��/�)mg�<����K;����L��mI�䧶2�� 9wDZׇ����*�k㲔��m�*԰�uG��հ�9~��s����\	����?S\��#t?fvu���Oa�1T�[�V�mxCA7{LT��ƒ�>\�x ������1�LdP��%�8���z��x��3�40�L�ɶN�KE���K��ϳ�=%`�`i.g��w��p��:XlxVHYEB     400     1f0Ɇ)������U�p'<�b�P�y��(K�p�۩� 򗠨5��|��`��S7U�lj�|�~��fK��R��E�P*!lܳ��.��![}K$�
��ҝZ!jzОO��n �'V�\����z�FH�Ţ����!3c�ĉߨ2�"�Xˉ�6��
�>�I���ȗI�1 �LRA�3�����	���P|g��C��\�>�Fa�5'�g"��Ҝ�aBp9!�t�7�(Y9������`��&�a�bx�2��Vw����+�,t��7Π�uT��k �7D���(����D	zA��D@s}`'�h.�e]<���W���Z�uZ����xv���S;�g�a��$PvO�n	""�n��:�"ը�_JŊs��eϣ�%dl�1����C�n�"�a�a�^��M �<���I9����N��Aێ]���K������<5+e���	��-8���U2���i�B.fk���!��w��4f��K�XlxVHYEB     400     130P=�4&,8qֽH:J�1�Na��
^�}��+�*�]���#C��]���"<��������'y� S�N5�q�B������G]������7�j�ռ_�n!Y<���ݍ�;��:|�<�g(,��s���{�����k�k�}�����*JuR��l`�g�����CZ���f,E@
�%so�F!���$S������4�u��OƟX�������������ʠ�Snp՜	8�I2�q���잰p�̵#���} 6���c��L'ʑ������_��W]Gš���6��j-�aaXlxVHYEB     400     190bQkM���Ӷ�L��0e"</_�Q�B�ҋDy�l�8�I����A�~7l)e"Wg�R���\�,.XC�"���$�_8�`�~0^��Ţ�pq��:mj�;�NM�1͐yGq�	�e�؜�=Ǯx-OZA.�&�0����P�:�%	�+Y 8�s�Ɣ d��q�)���_�mT(å"67xn���D`|��c�#.����#Dv�fC�=Fx�خ�k�˰A A���n�ܴ^�^���<G=u��^1s	��^҅�+��n�' ��y�ڊ��&%�}'�a~��q�Ѫ�&�'TM�%�D	ɽV cC�����6��,V	X����p����w�7|�ŋ�R;9T�V��
��Æ�j u�TB�@/N���]�_�Nz+o@��>*��b�XlxVHYEB     400     190fƳtࡃQ\��j(Z�"l7>ۦl֤=���I֔��=P�=���#Z�.�\ń,Y��oFFv�	�Ɂ�}0Ho��,�P��ܸ0�̮9'�K'�P���L���	g:)DޢL�Qߞ߀����{����&f�J<����I�?�Dy��E��եu�����{��^���[c
�md�9��4��?t�9J���㪜8I�G�"��"��iXȵ�}�Jp,�b}ƴ��B�����#��}(gB���E3ڻ��Նm\k�N�z��vU�dtk�"������6���
�aˋ���L=��(��A��"�"h�h�EZAf�bq[e�C�},���>��h��ve&~��}�"�w7"Թ�@���ć�5�k�˱��/XlxVHYEB     400     120��X��:��R�o��b�� ��\V)4$0���L�]�I�0�ڈ9\��H+\Q���@Lǵ��i �X?^pN��oBE�e��fKZ,1���R�����h����j^Cf�,���S�X-7d���4��v2K�Y�ʛ~�#>.���5�w�w1B%X%��M�;P� ,���'՚���H$ה.P��!�Y5���gu8��(�NZ�G<o��0��/~�J"��8�HhT2h�.p��v>�aWY�`j"
W��q*��������GS�iD�7�w~�����XlxVHYEB     400     1709�M7��F���"F��̪Uk"����O�'�{
��h�͟ϰX��d�;{��/�>ꄀ�/�L{��=�'�nq�_��i�.�X�(�lw����W���_卭��FLI��PpJH��	��r^@h��ţ`�Q(^<c���4����,����FI-��.�+��S�I�\�:Ԅ�:��+sGL���6Q='8/����u�a���U���{3�9oc;��%h�����fam��]�E�+�WR��ѥ�k�b�ra�g
;�,�%�A ���<Ž��c�ӂ�����a1#�ͺ��aO�ʦ�ߚ�I�n���4�h� RI��)�uĨ?��MHt�v��f���Os��.$،���;�XlxVHYEB     400     170������Xt�n\e�{iX���0u��[��E��������CB�>��G֩�g��]z��$���|�:�֗�%��� IZ.����ucB�/u 2�_�j�e`0�[�D1����;��?��%0�[�2�	�n��b��֜�T�D�q�ܼ=�(�tp�M����5�Wk�����OLA�vA�ɮI���ʮ����X>���0 ~ҜhoQ2u7��%i[�TŽ�������c�΢�����1[!I�a�dQ.�|�yL5��"\83/t�� �(�W$�C����}�=�M�u�[�d
b��8�B.�X1X�b�F#�%�±PU���+YI� W���g:?� ��	����}C�%\@;XlxVHYEB     400     180j~_�	��V�6��lǚx�pٳNB�@�3 ��m��uA�{���Т]��tz�;C�Lo�QB�����9`צX\+�r/@Y��r؛*��uT�_�.;�7�0zt�7���ı�a�$KI�%Q���u3�6��V]d̏���u��.!���: 2%��ڑJ.ȑ#�A����BO�d��T6�c)^���@����J��h��pKC� ��{�\���
�{���B��d{���+oԭҳ�
���2-2#pMz"\�%oW���D��m�x2�0�X����sH����f�e�����Iܺ��Cx�w<���n��004���t� �0��2�0u�I��ݤ�n/ct^ʦs�/�
��4��_nUC�T%�mXlxVHYEB     400     100�1�E�Х	P�2�p-���mx��p���j1C�+�sU��h�(]̐{��~{�q�%�#L��q1ꝝz������D�� �.��D�r����u�����Q��a�'�<�3f�A�0�O2]��FڪF}G�P��8J���̷���[*l���0XW��@-�1G? j9�stQ���]b��Ъf����@}C3��~­{ �����x��b�cM(�PYcK�oc��rB��t`���Pm]3W�H��9RXlxVHYEB     400     150�l6L�3�4vJ�m����EX���X+]'	�y���M� C��ʰ�8����8�r>�)�:!��Jh�����L�\������87v�՟�咁i��ermU;,{[Y7�H�l��jO��u6��7 ci��f�����&�����'gsD O/Q����&���"�ӳ,�	�u0}�Eʕr?� _�����UjA��Я��e�t��S[^r��hO���)>�����i#:����e��d}%�:�0eE*u���#A�@���Gf�� ���/�9$d����=ϷЁ~�q�K����3!�8�P���'A ��B��XlxVHYEB     400     150�kZ+��+�>�rm|��L�ި7=�Vɒ[;LjBk����a��w|����fd�A��D����hA�vl	�;�d�Z��UQ�c6�ǥ��6�J�m=N��]������aFV��}R׏$I�o~u����9��ZF�K��k�XWao+��&хG� ��Qi3K�j��̽��v��n���/E�˽CX*<����A���/04�@:��_��1�䟇n*�1��c	>z@Rlھ�?��r��b��r8�]���B�j�!����ڥ�v��m}���D����h�w��o}"��U�jfF(��t�iNk^�Ϩ���8g�c��;UI۫+�R7�XlxVHYEB     400     150�ȈYS�!�t6y�*Pv�O/̈Y�g�8r�ϙk!�C�QeF�?�ǹ��2���A��WҞA�*�J�����uc�Ѳ] ���
��n<�YfY��g"c	D$��М�(�݅5�p֦� ��X�_ `�5aH�QϲGbR�@� r���q���[�,/J��jg�5`��� �e)c|�:�v׷M�ˑ�ٵ�N%m̿���1���t�j�}�h�ׁD/�GH'����-A(�c���y֮��+$��4ڤ���!j�	�ז�QY��&�Sp��j:��q{0q�=����3�@{����]j�F.Ҟ%��B��Hg4�|����Ȋ!���XlxVHYEB     400     180!f�d^�Oˤ���a]i) /Xm�
.tt蜟hYv{H�nc��=��k́����o�ߋ}A�!o��[� ��mz_����Cv��&O�?��a�W/b�pƨ��Rk�^�m`c��5$KQ�hV���:����pB�.I�����P�6��~�[		�$W����y����i3��w�i�(�OW	�S7ʔ��J�$�r����>�hr��RiDa4�20eG��gq��D[{HC���e���aG��7�1��s����]�Y����"���t�S:���{�9M�v�@A���l�A�-˂�N��t�_�?H':�>~?��A��(q{.�q��5oO�J��S���.�3R�
l�U��iuka�x$yE�5|q5XL�0�1XlxVHYEB     400     160�Z�o�EƐnY�	�����XsjPj���Ji�`�;$���[s����Q@W�$���L��"��S�ׄ�0A���:q5 �!�`0��#��B�hg�
�=Ls����4l����x�o�Ǿ��w%:BC�̏y�����)�z��_P�Y!?��Kr; ��8��7q�V�N@:�^t�)�4,��4߆��`�q��$[����\���趯���G��pݖ,d׹�QS��!���J�#���E��SMv�%��0���;�;fc���7�ٟ�z漬o��iF�k�c�/�>�lk�V���4�,g=0sKR�����}IQ0��t%(��5�
u�`�	[�y*v��3DyImXlxVHYEB     400     1a0v��C?L�/���}����rb�/�ꆂȠ�ޅe �@���Z�֠^���Y�E�r6`_�od��0�d�?�p3�O�Oh���-ӽ
</(�Ȇͧl���bt'Ё�M.�!�D��"��<�A
�a���1�]�>�Ca�.6tAq��[��g�۽���3��_�q�]�D�$3XԵ�x�8�T͂�>�G@\�`I-\x4 �
���`�E�2�M�ƃ�#�;����2�aO8;�.�Zi:e%0�Z �F�ϝ�l��f�r�hL31@8�Th���� j�S�G]� 	�歜�w�"-����sX��zUߑܲ�>��1~ <�(Cauɶ�SW��[�A��%j� ����9���_�Ɗ0s�&e~.��t����T��>�5|��m%�"%9��Ν�뽖,���O�,�6k�R�]XlxVHYEB     400     1f0
��ցt���޶��}��ЗʹS��ʥT�Ǻ,kKu����`��Z�[��<��~�=�Md-�V��k8�N��t}Gǔ��.U�������9��_�t�Y@��<A�:�����5�&O�{�!�E����l�=F�@Ίmݒp�!�Eq}�<��& t^����֓�U��՚���KC`��^,ʐ$_vƔ1X���8X�٤����o�h�s:��L���
#�3�l_t����nx�f�^�$�D��`az�Y�l\���q�?,�`,|0~���rZ���S�3��]5�n�u�u)+>�Q_G]�5y��<�x֝Z�`f)E5e�I�8ђP0t/��'ۦ&*���%�����glO6��X=x�ekjih��h�U� sS�E���#�����v.3��?y��/Yjnk\�X�|��^�?�
�f���ǎkY�	GN�v�&��9�Y!F[��C�	�����rʇpE7���>��%m�/�yV�p��u4;:�XlxVHYEB     400     140\6�p�V�H�B��L��q����#~J_��nT���|��td�s�b#�m�5 gP�V�%�Q����d�?�P��zo�R*^/ʰ ���i������'C��&�:N�l��u���,�}��d�O���ʤ�������8������~02���Χ��ﾀ�!RЩ��ޙ3&H�IR@0��R޸h'�_�� ,��K�w܈��)�	��l��b�@s����[�hD�n�b�9��"bi|c���7؎�8��C\��E��J{�A	�G����� Y�� �{�o�����G���8e2��*�b��� ��7�[�XlxVHYEB     400     140q,�Q1`nj�l�S�f� ��$��E���T�~����ބ�r��j,��s���۞�Tu}���E��4��l�k1=��؆@ċ��/�+d�nM��'Ra���e NW.�"�t������D�]��ͭ�i�=o�	C���XE�_��pO3�8����pѓ�w�KT[kv�����k�༌��e��ř��r3H�����;'���sOI���QR��mѶ.vDE����>�xk��p�/����6]�����#$* �
�vF�yŒ[u�ÿa���o��F�G�Ot`�J�|� z�Q6�,�>��XlxVHYEB     400     1e0U���Ç@�J�4�� �H�>��z�-��U��kj���R'��J[ӱ���W�736��x�$��E��B	IO�y�T(*n${�fh�mwT����o�_B!1����y�Q��,G�a����>N..�����t��Ī&h��R`�,�D�*3�J��������;���;bFQ4Ѐ���̛.(�jS=��?֗�u'	qB�ᄈh�լٸ.���L:}�,}�̟7�$����ޤ�I	N������ ��̭��=E�w�<�]%��nk�������@���YK"�;�>�_��D�A$ͭ���lsC7�5r��{��D������a�����)o<�� c��R?�-��D�����"��s��?�)QC��9��;
n�i��;b5�!���6nK��D���#~Q�,T��^�+ݱNكjo�̈	a������p&���k)3c��B/<<�uXlxVHYEB      90      90���nvt�Zx�������(�`(�}Z�q�=��_�/X�p�O�g����F����a&�f�����=H���o��I�QBAY�Ʃ�h��
�2-�ë���� ��h��`ğ�Ɨ�� 5���m"��$�Y�mm�ŏ����-