`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
uMjuzPY0HZ3vC95H+Aygq1nKuewQsbhDm64xqgO2KaLV3cuZ6wr+m+o5cRVTvhECDhKZjMN973hN
d3Dns+Y5x2TJMdWC3cumGUYznefZHsEANr0LI4IB03HGzsshx5sCLBtBmON4INbRRkqxxI7WAIn3
o8IhHGYXLNU9q0RolgnJaCu1FSnFdbIj03yLIUX2n52PGMPeuF18rTldHnHLh4xywxe+IVSdQj/2
6U8IyDou+B6hgqUSiFJbMaTDAHYpZVEo+IBDmdMvu8QUeK1gNo13+Vx0cgh4DrLVWCbM5KbjNA9I
Mo25dlmcYV7Gt3jIL2TQKF684gbG+4Na2L246g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="MbujOblCV1m8V0YmoBz5gNhfr6uIPHjsJcypgdgV5kc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25808)
`protect data_block
sMZMEEGf7j8vXEx+oabZ7/pZhKCnxrudn8O1ZZd3QGk4VCBMXPUcBOsJXMupLrjv6fUpDxkdxzih
4d8mDLJCNCBF7KBDud+sSiskpDUzn1o2asEfUy5K9Pyzz+eFeO7PbT+5FtyPehEl4lHh1N3tInVc
W6IBC6xJqZcKqfCJn8MyCfD+shac0w6zbRiEdV05mJVmnOb1ttO7eHDW2ZtUy0+XI7w12ogIVJwx
sLM+9K0Dg8xhVWfRDlbN+x8DnrJJSY23srxfROF8bvj4lsgDq0JRHLPpBYLBm5tY45vzFaDgcPSu
VXxkFvE4MbIxra60pWVtlkObkIZwpGTaxUiebKDRvJVgn+TP0AxURGH6end6yTM/1cgQAPfyTrIM
234VX+dJe48j3On4BDvWxqGcenilb+RhVL+0jwZBv5jWe7psSKNPk0S2R+V8kBzp6/+qFE/ZQwyq
q8qExQjRiejv1fpZKpMvw8PIjaaXT08WqTljqjMD0colGbRRZ8eUxRpfhsi1Zi7Oq7QSotSxHESb
1w5tB2ZG6IZ55Q55fO5A2FlUih8z5q/guGBAQeBkM/d+9kpK5oYVCNulrlnO63XeaFn43wx1qvdP
UDDAF8RSaXGo/eGOds7FUsAJ5Lkfpl9KSQiggXt3u9950MRxJ/9mNVpE5VDGcUE4Ju4451ssYGp7
RzJe9JFzXMFl9Fh9m46Mm3Lc7M3LtJ9tQIhSl8HrDgbUuKLyrEhXNVEsl5+1bs2ZsI40IKmQkSdr
jbxLErmeciUtAM/7aLYGcRr3HGpaxfp9kvxll/Alx0n02WmmEVaroaq39wRIOyDIVpPk97x0Rnwi
Mr/dCt7XCIKVlFZ7nFME2m0072LpmSTwesIUVngkTTCmXVP3F1CkT8dnDKlyYRKVWRYDC5aJzZwg
MTar/sHI5pTZbKly9l5RAzZZASN9n/d0BXde5Jj1Q5VzWRLrcFvcdACBIp89VGXNSgoM1swwd9Yu
lvC1iMq+aWDzvB/Fjr9HujNivuoxUDYH4ccqgxn6DhBAVXSFBwqVoVY7zmoobPDbtf+zFw3gCt8J
gOb+OY2cHsyATL/SJLbH5eP7jR1TyIIiS73ysRdRmct4jzhD/CxqwjXeDNdO4sH9aq9ofoOec3Ei
ne9B1QCbOzDkf1pi+T7bmBeK0Bf8TsnBePGkfx+gFcsT3FiLQo5nLilCAKJGxbKcJkv0RNQE8tRE
JJnC/ootsPSrkSthuMCQ5OVGOhZ6n/PwiS/28CNVb5eKb0t6TLfRfsLmI1JJ6BeVAompGSzBQ02I
qs+xeUuApacgRvqiqGKFSZ6BgFhxruVd1NZ9YjF2jIwGMgmRisXrRfkspl3a4enLVxzt7Q9frWkT
LjUZ/QCDh6oUfN+ysYOwkkk0mOxTb7d4xZ/AxBtpz81iYtHmyUaC7gAONM2ZRFGDLBkdJ9ZEB421
IWrNrOHH8v1VdjL3SSQJw+1RZqRMgW4RAeHyn5ugtVxr0fGjSY2J4UiWCz796LUi0ei6Z7j1LTl2
Z+LCCPk0SEsKnIpjWVH6jDqL44DVZ5J+ASK8b79AMpl22jQBkJwSMsGuIG0sksNNcYt+VSCbDIIq
utWBKj+lCs+tythtWhU+8M2JjQAQBrV7ppCr1tRPgnndmUdvHzqUsNtk0hxemppA54LD5dB/+0nu
gWeKFnra0ThbTXWQ7fOPzOQpfLyKzbDiyXp75g6n2/oasC9RM15cD9p0cMlsQ0fNCwaYWIiaT3FV
2gIh1FoD+e6ClIt3hTTryz2VPObnQtkWlwShaiPMQnt2NTNfwfhgSBmsK9ZAGfYfoPvk+QrCHjSX
zX0UXcRRDfYkIX55ClTHc0hG+K/mT3rcwmsHqONkjcHpQi4ujqKv9MsZUrazP/k32Mcry/Rgo1tz
0GITQyjG5lQXufXHbgVTk2wWICxv6qe6PDj4yglViTY1QoCLOOxXbwY33pGYR1LRQZglHZeiCKnQ
IBupY5NdaRqcE8sROz3BDzGzBtPvuoPcy6wnwop47LvvvhMV7rFbS2JoFeRcY6Rjj0sniWHus0Rb
pqACNWzUcYI5j9ACQ01WGHQK9syD8cZQqd/gI6GJG7Nm8EFCL5ZFL26AxLXogUWRXEZLczOxe4PU
BwBKFUDVMb82quNfAkhXdnV0fjGJe+Q8Yi1GpoM0Ew9mruH3nOveCjO3FCsBsFP4vAd+WvHiiJiz
NZj6yHCJyYEPVToywHOekrfcfEkJO6JmrzY1Xx4w7QVC7eKgLfc76dxB4QJjZqG0RFJglkczwaOm
VZHRtMHCsYAaXbElcXwZSEFQHv3uRnEBfZQbrY+sTxf1hMMMWtU9ix49A4Dixda3QzzBmgwiFU4o
Th9pwKleWbdJMBAmZ9Q0ahjS2+E1PGf34PUsPxRD+VPVMtV5Y4qv/xeEMrCHxBR4Zh/FCU+Vf8KG
toTIgtIG/99NFOxR/LA6cujTiLz46/wz4H6fGQQA5nlTc63Ss1OrDJK8U6VDgQYUUUCLP6MRT8Jb
ASJwoMD8VwPyo07LUT+6NjKfWptChj3XIPiF66HMpk6u8W87Pz5QunJto8Asr4SNkuGgCahjW0Hk
BPrlXGraAX+Azj6rUa33tyHpyeI16J2uCrCXacAlHAkHUjR980EUnxCxj7yGSHxz/62eqshZI6Hw
VYEsjrpgfRH+30F9cFdopTnHDInXy/prDFMSMgfrgrdSGgvRBy40VKoWoMA94h/drVh2FtA7lMOW
gSVPcbf9EAyFkb4DgaOLQKzcI3Ny9ZikP8P9LZgyv4Woy0RWcD4kobl6DxSrGiN849Uo1910qxNc
EALIXvNCqDcg2qnj9Po2wO9yT/a46mAjjmITzbxTCodiLmJ0XizHfr1kHJrqkQxFXPU8eV0gB42y
2/Sx8Y8qFgabPRbJ3vT64hz11zfmHX96yYRi0jMK7Osqbx8PUO9EzPETXlXFcmaDg4VDIrJb+zPJ
dqRw8c86rAGHdKCqOYhy9KULGHkdJyYEg4xjp+ze5nx4n5PnSg/JuHGkJhKXHFsKijULS+2eg3No
t77uHprDH2r5XjFOU0YisrjYXOs/aLz4WcowD9WucJ8/cbeilg61rDC6eNItMdKT/v0VaRhy0i2B
P5MY1Dc1hlAILZbDuUsv6I9wibGEt3eVnPnoNM4bOX1dLP1ch8wPvMi62QT5JSjJhu7ocRVTexqw
vLoOVFutFeDQXcQF3346cB1i3W9jU+HGMu7oUzg9k6/JFxNxM12eOjGtvuJCD/WX39AsKr4mYfK9
okDh+CpWklgZvGZMVeU4YeT/GwH1/mVhy23LbXy5/p+HIuQge03DxB7ahI99JbB6WXUFRavPFeYL
ISXi85R+h+LOSNDP97rO84GRCZfc9YHpjNUOhrU4R/cpTTJ9gimMiOuW1IsrbF0fPDH3FRVAy0Q2
0wcCd/6BDaVxHgwzPge80s9hUYJjewAnhHikgGKcs7GbOZnoZqHShUQWdW1UpWqhZgJXg6KKZkNn
LtmeTpY8jtJFzxdvPm010xKbWujwWrbTOgStjqU0Oi998MPsyPT14m4hx8UXyKrG7yqsBEx/H1HR
GcUjo4WCvTrw2VjwDPyud+lANgVTdtTpQ0U+ap2iO5oxAklutCnNbNrkck7bitMz52UJ3R4xsFbw
Xv4PohM06+jA3ILnYCdhCujh+fBU0lmsz03eNsPLa+7uQ4f3v2m+8mpDNa0NfiyIP6dNaB/QINfp
R4wifaFhey9JqotmfpannDpwcW4g7v4/38K6CAHFqgrjF/zVHX09W6ahb9EUQPyLXDx7VoX9Hr0J
2Ezx8PmeIHnq4VgFnzWaXEeg1mCssb90sI5hLHYWXjqBSDzdEPvoi9Vlq/g0tDDAVNbfOv2eAgY2
cHVnX4SECa/PYfCVajXbdYAa/YAZIGp4aVdoEO/sfQPx1zVJMPq5dEg4RZDDTJxuJ/5VSYAnGvv/
pExUt70+l2c9zSDB83Q6AWu7ZZl0KqGYHJH2CTDmQuEQsr9Q9E6Rdc8Xnj2dv0Ew5qQjPzr6leJD
Fh1dKHanTCM1JGWvvD1ZFwDmchUkY8dixNyV4XO8fo3XN5Lsox6GZLbFxw3EeNbqvk7g6beMsg2H
nyw3Kfv/2a6q5QoWDpI2b9KjtSY+elruDaoCwQy8k52vgv+m/9Ce0tt2FPUGqHUswynR2FqN/GSi
QW7dwxZf3rtX9jk3ZKZG0/VeBktkFpZHluZvC/hoh3UOB6i50zfAwH8+D6sFyfrWTlxw1qZab/s5
n1DFMEjznKhAZm8tnuDWOlYkiQ4UTDXxMa3BsEXzvGspne4RdnDqkU1msXIchYCmphc20FYjM5zs
2i1wd1avAHKu97Fjb2fS+VvjIoAS59jNmy9kqSjoqzyVDGYH2NsLBz9b+eEMLPP0keNTdqRpsWDH
S/c4OxBD7EF0WNZT6x1uLaYwVNKSI04MGY1XaxXWawUQy0LeKVafBCvuAeH6OWxE0+R/gVC20/PG
GnAgjcLfKohBOCh1vtFyZScehqYsxnZcqDaiZnGgbx9wzGJogPqD/0jZMe4/WmABd7VfVSW4ti+G
8jzdvziKklDvj6JNIxLheVjy++whAHNkRPAiPB8bJc4/82rE9sJqKAbht7FksADVS3opiwWWT4Ho
tWOifn0T2HLg7PPvyCg4E5SYKspaipEDS/MZVwGfoXI4zCEo9CE60eXQAq9LwwMs4dOYDNSYBcik
YHG47En6bpIjMqXpWoVzAXHzB+HDmjoI2mHIp68Dzk0rv5sxaCM5ll3RmBK5sbmWjq51iWs5EY4X
F43nZJQeM9TEfjVsqfEHeJ6ht4wltcxbNflhqUsTu5txGQtecFPXhXa53jBePW71blEqiFdyf3fc
GSUCDkrinv+fGomP7uVexarnNwyXQPZPsJKVUSGRxuw2+qguA/frM5F1xgXL+SX98bJh3r6vBh0J
8bev7V5nHuEplrXA0igwUQwCti8ot3zx7Tt4msjrcnifiNoDKMZgq2sCsjuQ78rejN21Aj9yeK4H
aDWRe9YDJqHmWMqCN88Q/g6e0lFSxY2Fn/YkBkIEe1FdpUmntujaNEgbTFAEl9uuthddFMC3kXWc
WnHFoMkmQRCBeCvhWT8sFJzjozQ4vt1ONuv0+pe+GZA0UV8L7knwGlWZZbejWwXPUWCd5EHrCpvs
32mi01chWSD5giTw8kYLwoR569gLKqfT/l/8cTfuR8IB5gW0j08SBIgxDyu0GqrT0/AUhoQGKfZx
PK3yB/5tDY0s228w5d3MPP1m233cCefABdGOZW2mDiNNn2ChxenBNsr+nyz3BvLknVFPvuuaf+qt
YSKV/qXOoIjZNR+PzbH/Mhl3cFLRAzc0I9yZOi2EwUe590Hk9UXsFi5VKXOSfOPw0mijvCW6fQZW
0ANPy3UhBOeb9Jd3l1O2szCJENE1sESH04GEbweJrzOqZxSND7KHdaCke8b3p34nFxyImrqNNYnC
Zp881r5MInfQ2MTdYMhIJIIrRqQxmQTWltl/RkUZJ7/BLbxa0VU1u8Ii0IP3+P0DJ0oB9i8BK4eP
EqjnoGlYNuX/9fF2nPrZG/ZphDFAeNhCYQGChY05/tPIuz6SyEEyUP8+XTcAKJhIHRvUJrdxi+mF
cTiIcj9n72wiRXgcYdd1SRGb0eFFlcrjbusZcB2/aiwm8VAKToRHrQSJeLZf77ApcV0qu8u4WL4f
ejxlWvs/r39C2g9KBOli/v1qNsfvjfnCY+322IzPRUdCJQKoTmAmCUNguHh6Fx+6kYICdf219fx/
lL9PhrCfsXEcA285Y3eMRmzaqEoa+80we6yxAzISD8fWhE+BZz55FuJnl0flw2TZ8u9rY6kWaSjd
kyEckIoD8kFMD4iwKc5Mhfn46M3VxX4FE3Tnqe9Qe8kH4u7mZD89C9EpGuYg81vnU7O53bGr0qKe
mCKgjyV17NpjS8+j3zJUtEqm9AomsJuP7aW0EgopXPKqajVzRK699yr7X5OqOh+APQLNp6YcDeuq
uuWLdkxC5HfglGuKV1NLghT/TJ/mpUHROUn+aiD1CZ0ZXZVR0LCIz/mzzhDFh8g8m2fzpqUcaB22
IN15TwClZDOt7P2br1DecSd488fxglA0e94ScDICXQkVqzYpvwKqB2bRc9ocCvEZoNa/p1D+Bd1A
E4WxvUYVIft9afCxG6NhTsRyHmRwf6JLfXYAVrBqsH71tAYQYuJGcIqFwbQPtZjKsFN7e60pDzgj
Kah8AL2pqnt7NdTB9lNBGU7eWslWsO9gSFRk9P+rU3aq0scDW6E2rA+DRgVxQYP5TXgpoEnC+i/l
uOFXbKgAWbWHSnQMGMBGBGUcmB5AsgnLH5VB2EGoTArF6r/1wptmrezHnfsfhiZDy1XJTDDFSake
ekgBTGTMMicLWawZJpgFmZoEBQ2NUvXRMsgrs5SqCUMAhtxsQAXBYuuQvG6+u/r2wuHYt6Z9cV37
37qfVRrC/bhQptJlfUkM76VROnWRWptEENPga6D+eFK7D2rpTAA+pBHkdIVGD+SEK8AI1BMiAOyr
2QY70D2hshp57u1uKhYoe+1I9TDmGG6WIAAiwlRqt8rNjcUSVOxzBqKM0B8xcsKW4Ar3V+Vx+c07
BUTty1GRFmR6UZb96oEOujtbVa6LcSDjlFRRBqqyBJo75BjjHLwQKPElYNpztaM/I9dNKgCsTBZ0
54SIv3yEZTaS95UA9GR8hEUozkoWfmTQ/LCh3b0ds+LhNEZAmaqAzR0vTZ5wmGl50A3qckAGZ6g2
Br/yFwck2j3//TXcAhxtcl9JvF01ry0yYRtxvlWkKNR+ycJfpeaZ3L8RT/59HUXkZmgzTsfWv8z3
tpXD0qUH89Xde26UHQ3whM/NFslVYYFyQCSoLkQNAru6L0iMxXDOwD0qgbOv/4qn4S3fjzbKac0P
pplAqC+eGLFpU3SNfsGGubZs04EW4LSdS0Gq87/OBdu+xx8V+S1LLQyWB5NAPGVB5DNew4JWGFIB
li0jKSfQDHA7EOhYnU4NepCGMAu2pYu//wTlKujR400LK5DAwMJxoPXNa/0LfJAMEYTnmAzJeqCP
xxyYJmYwTdiM8d6qVfmrbiDKqueKTnqjZevZF3gqBzBBYpSR2tKcBZ45HgU8OPKPcafvzo0j1aV4
RLTKfVUL2no8NYTBvxPch1aVg/p2qFXa2RP874UXATZi4HxcsLxuXKn8L+hKsqmeKKdxi8K4ccpl
eZO16UlvK9CfNb7o2epcrcIeEx52g7Po4FpFVyfurqCrmg2qX7tbtmL2FbutoZIl2qK9E2U0YuMn
uwq4asEp0kXhUbAF/y7VlcnU7rBQvVxMaIZU1frZwGrwTE93viIuf0sGx9Xozh2SCcnwcRylxc07
vUnouhFXzr/s2hBU1fr5f3RI6l5eHewSTo/hCqQighJYOnIzCDTglgj/9+Y3ofHuI6ZV7R4xGWLQ
YnnaDO5MwZreQBhRNcsmxZszpu+nzPNaYjLSFhlaydKn1EsqVF5TsCL7ZWW23zJCBuhVV0iX15bk
ldDsKtllExzGCupZLPcR+7kenN8JZiYz7F2GjxD4MKun+TXuzqvnSBqtt0eWJsoDpGNtjMjE0BqS
Jq2Gs8JVSeg55UnTjtwCCTmoxw0sU0KyIlivpCClsUxtZRRiukb8iyuQNRWVIW+6XBmyXFTozBjd
SLum3ayNPisS+bCgEIAxWr3bwJD9nRtJW8d8uNCDLdo6s3YcPmdXZV28b0AFFNIjyZuWcfGxSk83
j5PKZqkszoEVsPl/bTlUuDdZPwxQxLpAePK1VicZ8AOowWYZBZYGK8D+syg2m6UnP6wFD+8NLH5z
wQ9z3Wa4YCuAZlePn7oEbOElEN30IEqz5kRYbbsQv3KD9pMYLf1uBNBkBStucPYgl1fSq6A7oiDy
uz3QenPPXdMQ/fWorvme4e0GkhITpFyu5Twx+maRoC+K+py7z1RNfAswNZx7ui9Og6iQhjktbHrC
vLd0d7TGc8BJqGdrOgVhhGQxcmyLDFo3uW+V46tbAXDDWppR2RcVpPeTmJMdU4dnw2jyn9FHpbnT
FjDn093ZS9Fc7iFW3LEN7JzyuAc/h6tRbUi1pOoR38M1gApKINldlnOzN0Io4UqCZ2+u05CY7eEJ
2NLDSvZ5A6R4HNr6YBl/3Z1W6ymoDyIBFG//6hM/525s+SEXOLoxMEmj1eE01kd8V8OT8EPSXi+P
1o90wbD2PFzTPBFHU6QrnEmHYpAMj/FNdnQXjkkOT4JNCOwZmu5+an9pNvd27klGgwCUUDUyip1K
NRIqlgyNZuCyu/WfOHjh3JFOwKHdvIcXRz4VwyfYDiv5yH7wcdCZTMPNrZXIlTO7XDccegaV4+j4
LAMYHwZJ1rlTwHbjfGslTM7mA8+biGNK637txObWrKA088IywTIyTnHoIJaPG6vKLpHnsnjM9JTj
LWds7KiHUWx34qXMIsXov0V2pE45BQsCExuEErxOkzVsjtv6jNTitXnPVUNqDsEzYvG/p6+OXXxl
d1kSGJBAp2PjtWImknixpR2UPVpV3PiMVNuOAMuR6PYHSPLskmDnFXgxDAkIrvhRH5glBASht+TD
qJMfO+6WdZNKUPpe8Wi55Zp1zJe6e7TH4W913hC2VoVz8Dqbnv8G4Nwgui4LXyRnm2TyP98TA3uu
iKhRUVzR5w7B8hIJrfg+dRSMTL8n8dCM71iZU9iEOIUyyi6bgoQJDOv2N8RilpoeI+59J0X32XvH
56m8H3lcYtaWN2oIqB+38zw4T3/Yr2huQn2HCd5GCpiLJSP8jtBvvYpK/VSBkfMXHaF6bhuopseq
0cuGeTw2A3y9qeqcx5b4e+ea3ZhuTv4AO0/FifpjHDPKvScz0g2FNeBeiHObo/XZ7Yw8X3byqvk1
hbWi+HrGgqQyHHxv0GFQGkQd/QVwR/eNNiazuYlVXiBM/Z+wEvjofEwoLljBhhJjq+X2NiXfvHe2
ZAyPf88DteWS9y0WP9C/FPpLjpSsdOiJSzdHYgOYPkTbGH5i+PLWMrbNAPSOMrI5esCzMW1JXviG
t9y3toIhWYa8avV+ybKK4OBtZzPmwRXWItdkMUFPFLwahdoVr7MXs5FQsbEbRvG1JcUPKxzCv6Zc
0TlAgoZF4RQKCm0ZDmOhVWwTGYEVFbxUz+y5nIe7azCv8nKLEsgK5NoMftPeNqBnVFQzcpcXbltS
y338l63kDhLZG+HaHEke+f3KHM75iUuCr7JyHDnMxAHp/qyS7bPc4CSpV+RGnnb2P3ymK9fkFaKH
Bjpqgde/Ru+ejMrntCj2VC89A9OTEkogQnE6X33nDAmwlw+eoq22j7395Oma3L3ttuOHFGMeIIQK
CUOP42YPLcR12FJoYHn0X3+aHE4O/1lpeW5gYiU2dxJFBpBPBUjIPP0f5H2YL1voY4MOgPf8V8rC
Y+jf7bvHrhe+dBCfnFLIrfQsmYIZkXwSime2AXtm19aw7yyjnQNqDkCeK3SpE+nYeZP7tcqkN+oe
pL+UVdOXszyUTBrd+XFoBTEZOXORWu/XWziMsk+oX0oZB+rSVlKwySgg6tsBz5u+gZD/MLL/UQai
4vyG65/WU8k7N3DL97CHo5VQrSBT8SGcGtrLDiYRa14MW4XGkiXFMgnIOHJlPlaYv7a09cdVNoEc
XwSkQ4uBOCF82hU5PCkuSWPNzZmi5fjlGtvYmmB3EeSyRUfexCGReoDeFo0CcufioWjvp9Z4U/Qk
aqEVFAfsTLhRLQvem/2o7v+MpOXyiKPeJFY/4VQl9NrrY3ZjsATBqb7Y8PuekD3mOEy3vhduWvTa
2NZcioK9vbUU6dqiadNEdze+CWz/uUZX20m2fvjhh+jiMXv/wU7CQiJ48FbqH/MJRTaXFVk1Y9Tg
RNH23BvtjUAhNayLVzvDA8/AQIUXwwlrQrFWPN7JGo/rFBUZzzXrEHfvMamWuTd+tkirUfPDP7Pb
Xkm4ehu1bcHteu1kQDtNfMiANdFrQtxFlpH2MH9PyhjAtmqP1PDSHMMLX3nzEsDQswNLMWCFc6lP
o1djSuWwroL0IitCzDgWczL+u12eJVZWFBStMLfRQMxAEd8zWjpIWSY1oW1825RnnWOhJINIAa7T
ZfdDarXakMr1rpQYjJjPdQ2N2aQzfH/AXIZAhggWlGqWTSpyEswlPCl9sSNFkFsrpB3UjziwlZFF
mVVQ89byw3DCF3JPUNmHr2gXHNnmLMOim2gkxMpgZhcSN431O+i9/NagfVpMV9belh7yhsxwNDjP
HXKwf6Ud9GyqX6gFQzSRyQ5yhJD0YucYhOd5Om0PlwZdsSHSiclb0wxvKKodYECoiD+85r3D+HN8
5GfydK8ZUJJ2AqKe8g3va/DM9Xni7X3nJdVuV5RCW6SttZ0O2rswYfFjq9f1AA+CZ6hLTedEBZgX
UufBGe2C/RhBAQe7WZqGUbTdZDhqV7wi41PELlyoTSt6IrFCht6QGzLuRncvnJJNCxf8fN/19FAI
5nmNhfi5V3KztL8NOvM8L/ENws7KoEDkVOUemXXUx4K24YlkfHtAQrJYpJ9k9JTvmuiWvxdOffqM
fqNXtGYHzNucw/G7w553MF05oGhKknaaa+o+RBdEgIXmQ2geMkspiqWyBfDDQv21vkOnTQZTVM9a
VcuoRqDys9CLPkX0F2eQwlTzIqXas+/dud6LiaCnUewxgU80/hBWHAU1tR5gyp8GXqw0Me3YU82I
30O60Xl1YdYXr+yQO2olEQrIgB4YX6Ygb9KVv6hj0oSYUBbV1ezzATbW6jh189RjSNnwB8I+pvz9
ymEDEhFKP6BduUTmIsRj7HR0NXdKJUpnpfHGcqZnDJqIlwOi+mfhuESYG/YFXN8ENrPhfj8IyW7b
ojERJaTtIRs2bNsKeaVoU4gdsQsXwfynEyWonAcJ1D5K/2hnWfi2mCmupmbqM2PpayAIrNnYM6PQ
NajplY3+D/YlqoFC7hXxnQu/S5bzJxzwIB+EbgpnovRPrdJD4JmM1aXXBzoYzzhhpQGEkqekxdWY
2UMnUEoDt5pe+RSEGyE7XVKRLmWxvtHhUjJZ2QqwytYjaYvstzXymxJeBD5oj7R5LFR+FcSkKcDM
t8wht6m/FerQ8cuBPJlGGK/icbKREOw3UZd5IkbUE8uVEuCR20nupATTEnUwZlK2X87MzHwTaoo7
4K1WrvkskL6XqB/HFRyaY4uKm0vjB1zfBEJ1tfVDsK2vPkz9uaIHFxvyM48QxLBnbBthS4iv2pc7
ih3Tp5qbtpfJLZJgsaIvVY53oGtZGyMrB+WCLdZNGh5+pCYgYsFUwiDxooWNG5nMWbL6KTfI1s8o
4XWdD1rzsBv0QS23lrZ9MfqLqVO+9fPLbl8RN0duwvdAQYOXIUypSdRpu8FHhdUtNPP9mhQWaIh8
Qa7PB2ygmHdIEIsW2B6SLXJ8Bt7w+Haa2CUPFYOetmwt90tbFASaGxlqLo6GeIbbF5smrBAC32M8
moM1ogylbQnWCTfajKrkc+i6sL/spI5oAJdFsFpcxAhwB9amioOS5xs5QQyFTrP94tSbCslk0D7V
QwDc1getOLpOTKv/XRmyn6tSBolPzO8qBS7AcAMKMdCch1SVmPHOTyTNbeCZ/sgm9DI4WKRg/yJk
NEF/AVvFZ3yybwn1x9mpU0Pf1YMPSqmrE9J4kX9UDqWCmwpNL1EYp/ATy8wKy1ndA54n+hO+7Pnu
Yb3wT3TNat368uOK0oDSWVoYr1Y1FW100GzXyK5nr2wD50eYad8ovyn8X7CjOUIHn0F6fSfHuAvG
izpSG+yL4c6KSc7RxHmTqXnMGcjfS9B7YwA2DmfOaDQ5+QA6+B7Rn1WfZT+SU/fk0XtFUbqkh+Uk
SDxgeDImgfzuc0bvR3j2dzj4T+b+tdWYfEGPuinXvOu5CfQnP4vRNCAPyJCIClfxnZCbOD+5/pI/
qSmlIc3B8VjHRsXnCyHIcYguTMP16EDqL4s1vaNXkxLrnRX+P1g7Jelzd5SIPOp1on/UiwIu7X+o
TRePpCIVoEPVU2C4Vc5JChGiafKFcEJaKYJ3Babevrue0v0nDGpRr6qwUXBoNH+23c5vMKllLZzh
MTqHPxw7Bp3env878DFa3U3FakdnCJR7NoN5dNjfcjHn5VU31gRNl90xBVVJfo8mPg4W7siPXXPI
rqoA40uc4XtAQSKaoczXLP0Ui0YN/S8hUfZyRQY5ioyMJTvp26oufQqmPO2Ss6r1J/mFNIrDb57w
3/CEM2ZZWQdkuhqihYAhcem62TwFKbv12Xzgk+Rwr1Jk7sIGDSS/wiB/AY+VBoYr3XZVl6zbYMzo
YSuv2LnpnOTLUKHNuc6BH5953l+qfQatt0kNyLuxD7kBv68/wkppXdhweUYeqcsA6t9Fe3EBKZd3
gWA2YgPfBj03tfFwM4jMptwoZWK+ul9we6U3LfcypMtIFvYVDAshSn5dTQseeJjqRMZxF5dB3B3P
GaTi8b1niWSF1JHexv2NXSpY+yOmj4/PPuxxmOxlPOQfTGlQ21hYrRVrXRiRoFIAitOIw/q1Lc/H
lO4holmbffzPTtaDB+6C/335uT0uxZo+C1MlTkCdfHumVhGfkdt0PBu9/71eQ99Tgdh95QFjOSgR
MNDjD5H6d566Ohf+YO3HkwgnF6co4/i7lxT22abyPd94c/U00y1+4m2GRIWVCal6ZdJ7L3sE6TfF
uXPllLANVmA1pioVuWyLWkbazVojmTCXKH9CH4UjwDKJ9wlKvGRNOC350K6lOVHe1kh3E62jI5vA
xchiLqNMtwAnkMQeJxdyFirNCxcUY8fb7ptQKlMOM6gmaH1qyPdH2OLunyySR/fcEG40DfOjYRp7
+sPUANOenvHX2utoIyjfsJ5Ey5tjVhZx2b+eQuwL85vaJK49AfotXerTd0PV8q4hvb+N8TFkgu04
MrScxgCnIG4W6pfwXukr/k30QmOTA5CMy7dFljqFKOCFzYmJf2/ZOWnpsweNAIcD30uQ6Sf+17rr
2mTBzb8vrbrWxrhWaHBhACDclAje+66+KuFnH0UkgjZnA2YDRHMgrhKThEXiP6/ej4AVt6fCKyGF
+znPS7z2ubgFIxet0QWAnUT4UAwHX3fyTugSHRmNSZ4QxUXPjh0SiQs8env9RyDBncaWcHxVLqLY
ssaiCxYYmMQcAqdfBUUmQP6GHNWcrFASe6QfQbfy8VW03RLZ3j1sd8d4R8faHEsoIIDrAmrJMut4
4kBufFqHJ0U4nv1TCoLcQpW/f6Ul1f32RBP2QLiru1zeUvjPwQLMTsEZUpKJ1O7rEu/Xduw8Oou5
DfHTgzSYHdO23iiCIEzonz6N/fp4wwJ4NVa+Mr2A4rdG0f7SJcwWqxyvAMvEIgNImZk4llAMtHe6
x5Dr3f/mnEZAxRAxRy5VMoUE0svKRyCjU7YeWPdvmC/NnnZlx88JRRaI7waocNrB8hRItawLxB86
EFcR/EAFXeh8GLlbOqC9QPHr4ahxwkqXUwHplZsKhZwAadzOZMA7pgZ3dA4CnwT7os+R60drbafh
jymSCNd+XoVDStY+G6kE9MJCwfaQekYPuzkuFzkmdavb091o2QSAVKkPtg7qhIArdB2flUa8BsPY
g9z8QtA5hBzJdt1BPAINz5Ppw/ciQLBYscTpGkGp051TahXC5Nf4j9FaAzQQjYj6yG1sL8G8hHy0
kgQm6YKN7Q5CyTwUUgA/gp+PBrKXIaH5uuBEYX2DTwSrbwPkPpfKY7fwrSI6vm0gkI3PTsB0tODo
i9SUVfXNfBXy/lQFufgY1LpbItZrbck+I1sujSZKBiSy9o2u4Mn16PNz8YuvtupERe48EzieKItc
tMaCAZW6DXmPa4Wml2md3eR7LU9a+vFIsUXjNQvxxb3HYxXyC1YMbABbMUaAUHpjwyldLUVq8Y9d
UAXVE+ANjKmArp+MXUSzLOTb10LcnxVt2oxS4DwXYNKF0javorO9yrNmklEae5l0jm5eJ727XYm+
ckBQrd9c+oX3op2qSbKngB/lG+O17ICiOkyb3X0cqek/3V4s6iN9tBjCzBmxluH0YQ+8sGNjf+0u
bFCDF5f4eVx/6ChhJSJGm89hb2EG+hDVUf92S9kZhm0ffC8EAs9ujC05ppwUnr+CUK3ykhZUMIMU
gihW78cJyQY3KbuPtQZWv7NRXpA0tNVp/iz+NhsXTJmaQThHOYof18EToWncsCcYGKjJ8m2Dp0zY
eBJVFekbuKMuj7epRI8K6DgI2/LFiZRkq8wmm9Ugk9dVrKcwj2STbbmLDk79sA0o7BAmi88Tx1VT
nf2GP/DGTk1SAkwSjngvSKquqRaOlRnuUZHCl0BtUADc59c0rTPrkiJGWBmBJCaK3U0ypRI5tyUe
Ks6LLT5fRYNvokD5di/CwnZxVC5AcK3dse+E9R8ZC5OZrEvj5PvSoe8KDK4NBbXVPxKi/3lsKnDB
47FeasuEzFsiqjxNUS/XL82PT0cPEUwH9z6rjoQ2WTC5vxerGPL1f9J5ta4RX8xwnAiCG84QPAAr
lbce/yvhdmFFGDnS2neglQ5euU5s1a86wbADcvXYFQJIji+VZynyvn9uUoH8SGd0tGR6HpoypCzo
wWcn5RYb2PaCp7rbYCTACIiLZnOCZxRZ5TfOYr3ch4h2n41ayOe7CLKK3z7H5eCZ4oE6jIgvcoa5
32A6ZsGcO5CSLGHH2OLx/e3P0t07EbRyz1v5PsgYuLsSHWY/Ruy6DnzKPHG5lEjheyn3mganKNZh
RBi1Hvhs9mw26RPthdP1Mr2ZqL5tJAXO3w0TfOXzhkVEIS4Z+8eP5g+fJsCOiJ2zHwIbUJIjePrN
X1kHUqmS6iTznFUUlWeBA93ytcbV4ADJsTeFs+z2xug+3Ax39uheN8Wj3n/H3x8UZ7xzu5ulXRrk
3tcpciMM6iaSLS6tkFWAim5rMFSowH/L5p4YmM5K5fXe+wDlKlcSqEhwA/XDuhDSv55BUjmTnn94
Yz2hoG6oEQ12SDpXuaPCJHnLkDPEE7R2NZ6k1I9Zl3oezMjhBFsUBJ7ORZO24fizLRgPnG+c4Ixk
WwqOIzd2rWCCHzBCCPVnmckp5Thz+JBrO3eYus+X5bF6B58Qcy6PBILlTDD4aLPVLW6Yhet9JJqw
oxpkt+GgkSmyyYrFIfWhQpQF6JYPPNzyu15KhH9G0m+UMUf6012UonAJmcc4JD82ajmVUqxiOgtu
z0JoFtfOxywmBsUgN5KJwHWDxAawhnqnWOzN2j8fiqQDXH7k7IZXnHGGwH167ITBQwMpHjBbIQMO
mmDYMQahhuobT+5nFqdPbp0k5y8t9JoGxgjSU7zc296PIZofdCckI7Nyou3al1gQZ94yHW13xQNV
YNgZ5u8iUw0xuj2FLRrCxS5r6/L8uXJJLdnYb+UbHtQvKUjVejOqK3P4SxRLzL7YL1ITXKTxcfw8
6+8+PZlsyNYSPWf8edtIxImd8/9RUHuoI9UKwkXODdf2P25+S4UfLTAFsxHvNyUANzBHzHZjlC/m
RRfu9jBdBBaYeXK6cPgtwO5ltfJ1A62/r091YhtuY4/rhJMYbVsZS6YrdQyUzUp9b6m7EDjLSoRP
cEmgZDro4MuGQq79Kh2mV5x0AJPUaV0FysRZA2n9poF0U75I4GhFfyemTsyE9ItlRrSzxlrJMecF
lA86jporbX1WI+6c0bjLhf3FcgmQh6yz0HSgovV0ExmDpYr5qgwP1+4QuBuv9n88FLWQbvtmh8J5
PAORV+neFaF299NrbYlekpOjEnWn+rZt0jIaav4cNHuaRK2B+anNzMd6IFVWocQYmfJJIhWJNsYN
NvvM3d4/NbkGXFPrP4NEVy3X/HsSHQ9ytewGJD4pp07INTaPTc/MnDmk/Q3N8FzXfxJMoUvddTOv
KY1vDk/lG6EFFytGowEYcsdfZixpFCG6tCD9xUMZ45irM4v+0hYLQhDixiIOVn5MMO+5DrgTdcci
w+KOsUrzy5c/jmZwRANfZPcLjLTLn1PyWoFQDVeljUWm0Mp4s/QdgQeH1Xzk7JUmrxOlsqA6GjZT
s6eSkgLVg1cFGFe/QD6/fVUEiV2mIJqIuXG0ZlYGiYlEE3xSchA1Za17IT+2ogS8eh6gE8br1J4p
bDtqVrpDvg2DunGMm8KoIYDcgkdorx/LIEp4HOjS6XyN9HdBTi3XExYA4/PFTEIu7DHorPcFeUch
ghSKQpKvrqeYvvJLZphk9v6nkM++A2tsRZNajxJZB/YgsBC6Kr4BPgso4DH7VOqL1aIEC3g7TNSm
/FGOeS93hFSfpsMv+qpjIH95OcfiSZ9Hob0z6yiStU/deDbeg/MjxCK6qCy8FA3rabLJWSglUDSf
rotQLOiHSxm9N/upF/BEEJCOdD7Dgy9PUbz+CyYILw3b5eNUXltQ/TEP5hnqtZSi7kbRmzuHFORJ
6RFYB6PNFHHefibKiCvtVMwUP5neTv9eQDxidOfRA1kn0368hD2glPMISXevxJjPzi1fWlcc44cI
9FFWQQN3CuGc7TwSXWwEwxaOqex5Q1O9Mt5U/11Qv2CoAasI2oiasjQA+AvkbuGFipghI+nzlc6n
nYxA5m6Jnn9YUSU2Z9BAZgDrBuKlTyuz8hYri/BoL+85wpS6mwGB+VXS0nb/ffViFGrKsedhGUyZ
BdWTwTE8OauwZ+Qv6BOsek/iUU6x4hxtjCD7q3ghwNOUjKzCRtcSiia2j6nusHfRms/Pwr0I9GcB
v0os1Lzcej8mmjcXkX/Cl/mDjBWlbDREwzx8OXICmseLWTWeBHZkCB6u4yDOszsKx7PvZ/WyWJCu
71vjDlUPRtB7rm9QJBI1+yU+JfPnjqlbhzNYn+vLqG2+cT7ot1zH1IdpP4eFgTpy+vgfhvpe9qbj
fm2t7A3HlKx6J82JpzmMsDnFS/QL6awWN5XrVFmYBNxL6DhoCkwD2yJhMv5tTQchNhfTZgbi8FDL
+OljMs0q2S/oAVZafK2cp3yp4TdH8WnyhimK9mEHRt67Pcw6O/GhQ6h33U8vOTR7BSlXAdNuD+3L
s5NH/XWRIQA7YtdTADpK5hWoCS6RKrObyBl4u/D/KcIrfyt8WdEvWSSr9FLIIt3vqebdEj4YwDjp
dgMK/1aAYkrubDImM6NoP77pRS5KQNXocqZKXD5k8xLzFXV8+dbcsEMRO7AOC1qzrU543DIiSVi6
PFpq2kPvfwJIrNYHO/rdCaP5XwGaaxZ9OxzBsH5hEjWSccwIynXXUjCMaCKrUNZCqM+l2l83407O
efrmxXQ/anAYzH8ywpl7hs1NsCw43kt/yR+609JqSTquxNuT83oih4ddCAl2FqLSkKPI3nP97HvH
KzmJl2GTA9IVuriZsRm6qufBXw3xeP++Zj+egzeA5Z6BhmEOGZAIXSn1f7Dvwip720BBS6h05+by
03ZvEjiUSxpS3qYjO8yXv9PPRZPY5NLEa9x8K1bQ6t2ZhLloeCAgDZJjG/kg5viyLS3NcmqkMTAu
j3Vo13WH1KbhQcudc+WLePXoeH7kGaDA7k0ZvSwKvA3lyKCu6OXpWNTAb53hG/aGdBGaxVRbrXQo
oRt7t8ARPBNjH2OHKlA56wuSI8S6cigQg2NDZToNkFNryaU97PwVYo2i9TYz7kQl1ltxPKLll/fU
dPo49oe7zlqV8ieJLwr+QFjwjkDSJA/xyC0DRMtXkCrDdWQjuQE0Uf+gmHocMfLK1gAmy1ahof9y
iBW8LMWq+AwgRa6lP4BL+ekB4WrvYtzBXHFaZO5FdSUr4hGKxxIpfsT8hC6xCMy8lq++su370chb
2416/0xba0IGRfRCZnpmaUojyACM4juNXTOUwK5oOOS4RDlJw0TSJ6+i4aNtnp1+euYYzwx5WY2Y
+murqUO7YqBY8W9Bnd91JwsyI6hk/hXO1wbJUbOuXuOj1XVnpf+Q0hBgUEqbUE47rH/Gh/YcI3sB
GkC6SKOcM6ebHzYpanqDc4576G6XzS+mrhdR13Sjj+dztd49rLJ0WbXhITxz+Sc+M5nfV8dPcYba
W9P8pyXztQZ00iA5cHb5WG+fd93inwK55KeFWX85TfzyOS5HlTzDX3vhYlsAb32VUprCw18vPQqL
0duN+pcbzcHne249wZE/GxXEf5g4NFeoALRRC3D8Ygp6RshT/qadoXe6xJA6HDSoxYGAgxqYFsUF
0BCXG2cYUO0AhuelR7DWCH30CGe7UzurhPj/PnGteKb5pkTny/7a27MMGsCWzJXAuBhuOmQb2SKU
i5YGrgEL/XWhJbJA2Wt3j1kXsPezZx+zMqJ3/weQHZX0FrP6nzbYU+a9ECwtCY39/MrOW0s65Dmr
SSUo1rvh7L+8g943EWxXASkyZW19KtfTH1osxQ/WN0KNgBsuF6E0qeReqHEzUYmbL6n/rnDmgaVK
CQmlGOgCxzasMbe7dlKeglH8QHr3hFK0lcg3e4MWf7I4PVpMthEEHs/GUYZuLz9xeUDw2Z9a+Pzt
dfTpYnzG2H9lz/0tlZgqgJ/uMqRHDYXdXLs2AUOqZTI1JvNLYgql5pL0Xu9tyExmFMz0Z1K/YjRm
zeetuEqZ9M42zX1OysBZXgoKrCz0tzfi/87FX0xOwvJn1/bQyq9qp4wvriN28jwsfNjs7o0E3LN/
z+ETyrQ2TmfwQvsZmNHJh9ssTfm7JBMttRHdZQs0u+IFOBB6dpIY6QRsmJ6rtitkJ8Xeg0Udl28w
OtTwwjwtOoR8GUym1DgC/uZRMCLQoH4NaivrKgXqr1Qy7h9IIUzvle4DEb8g2YrvejSkEZZDIq0U
DLD1NdLxMQ/JkrPif/VcKo9aR3meSAHu7fYz/lywPipxC1TSpiirh3Z0bKMSYksz873EVPqUd48A
nk+BmaoK+DtTfGMxDX2tyqjwQLhwLPPJEmLwNR5YIjRIF3C31B61npFM5VlMqQHb8OwuZoidOBPg
Dvl6vBmbdhDZzJKYfWH0Ml4ZeZReITVxv1gdf95s+YYtHXVrvGklVcC6YlqGd5ktTxagK9dH4pry
V3zmUtVIKgvqMAXvhd6ydLcGsEXOfaInAcxb/xiOfMgjclEXqcSi5TLYYZlEkIp/bonoDR5awZy5
7ANZLfTw44pvayh9HKiIWF32mfGlsaxKAHOmaUSdVK56yOCO9aEFkBtVvbP+GkORGKKZlEWeP3Oo
pD0AvKq/Q0WIgbe6vonbUBcWZep7ocuDxwieecEKOckA3Q8BBAnlCI9cAkT76pgu7U70XXGz8fLw
b7vk+kCAL18qIn7k7AyEC76kJUS1+b7IkKvaNynw1uhv4wxzRZkJrbUy2TODt1Vs41ILElh9M+TG
IhepS04Tbp8bywK2+81CpqfPVE4Asnd9LsIZm6CqY6DgOoEhq27NK/5Ly6234WoSyUoNNp2lS+N5
F03cU/nxFa2Bh5dGiwmY6Ne50i3Em5TaLLulOsSaeZ3CJV6gx21hOmilX4R61x1/WKhY4RoWiymt
Ve7dr3qCF1sIgD/Flw6qqCOKvWqCG2gqHUo7jxPv86D6u4CE5BtO3v852hMvBBWnD1sbxQYEMt6H
bAGyuTlfpaetAQOUvBa6H0FMf8BwUkzDmnQu2ivTwLmi09snJyBGUaWLnJZqWGpgaq/1ZRL3cehK
Bhapf1OloSUComxWrenRx6MLjicmjx5rdNiVY9ng2iQR1DhpdzPN+8P/UWMHirpHDIjJXcP44pE4
M8tOFBGfiLIGBNIewOIWtHZSn49S5FEu0yTB7YT5RirUnahqwTvfMf61V0YZHQzhp7ODdO69PE91
yM3Lq8LksxY96Fe2aqhXxRhDDit+XVqRgD0uvMBjvFCiQs1btRvX6SMnAvGgMwaiI77YCWmF5kbp
KyzkZA1n/cmc0rbvQggBVmutsoE5Bc9UPuG4yKfGh1q4iAmCUOMbdzjIpgSpxkw8KZ3CSrWCU0FU
xQj/6JDMpMXxhbAkw2TD+mUdnWdgQklVD74e4koTsae62prhd9av2vIbba6WLXjgxmBRwFsMc6t2
Za6qXzt3nxLAHlj84gXK134ogIFyLZ0r1oOtCeqcgTf5FnE3PpfOGOc+tJzaEHS0+J4xTNhvpQJl
zMEmVeOLN1IAYMTF0E5IIRpp5xFLbMbBr4Zd/rrp5zvJrJIJyqMCoAJHiiQEFr+xUtWH37ih3198
kDVU7LtOfdc2zKUNIbZ4Ibgm5xGjVYbNm7k2wy+SfNE4HnjysycSLVjTkpHiQM6zQ+83QA5FSMAZ
cvZYr/k7t8gd0aaIaqvWwpRWglOAxu6Qkn48oARmzq1/RHuLdIf7wm+/uyOvmrF2PeJKqpzW9IAm
gzwhypmQp6ptkdYRIB3MBKrlYe62ksXkXpuq5Df2iPupcICCI1Y3rNZly5NJ3NZwOM1/ZKMln6ZV
ymYbL2wUhVyZ0WuaDt2vU0+F7ckOKDTj5kvP/RKWn9AEIePr4XMRyniRJj7osXNtyfroZ/26NnQv
nmXEIs58lnCiGsRZ1Oeuo905WJSpD9DXZTWYMkxpoXzsSaJUduHFKA1ohXbQ7o179TVO/SCgwrqP
g5nTn35q8CXhU+PxG+KO1t4hUgNJEe5/ghV02ivN28ObhEIH2iuQMRcWUicW9zACihL6QLZW5eks
d3qZbnjPO/Ix0NweEa/njD2szIsVJiGQKetYIPBF9lJEWENu6qhKvXbzL73snfJSI+09WtKK4bqg
4hstrrSrtvXhFA5+tKGY36EYCWYtnxT3FkwWy8v5snsQRwZ9D4dBiqxnd/MjhZCK/KEibHPBhFXP
c44e3KEEwYrXpfzRZPjW523TFIUjmOojwXUzBF/g/6pjKURcGKZhU8jcDQzGAnzvsyC0hZvRqLaO
xV4+BaNq79U8A1NxZttEk01jmPs9MtTLhsIqxj5GO6y0i1nEIOubU2qToeGs9sEmZy6PJMdtxXWl
NZxdBU153S1RRDLmhPgn0HySaiaAoRK4QGP0xKRBNrKnZ9WmrrcE+3oTAvZOEmNjrZseOh/f2xT2
0hGbr3ER8RNtENDIEpEsuHyh+sewB4psZsod8cL3Jj5Ia+rYbpuuzwtXIm6e0EnQBi2b+Q6wDJv+
sUW/5ylrt4WOrETj9ORPpAW40/puvxP4DOE65hgyM0GgSRfhgEtuvfvbx9oAB7EJzCPT9BQ10XKi
GTjJged48VE3pMtBXsPka79pzVNqBr0YjnyzpacEQAUmPbQGTtE3/RtwKW3eqF5Xq3hj9IEoxI4I
hgZAML79GFoAcxa1bUCqoMPeskf2Ie1j1We21Rp3qOBPIMG93c3YjvshoBdhblAJd+2oCq7uilA7
qrZLaN2YvK+9tbtazetm5UsqPVcpZ26GKklMyqi7ynTZHAxMOf3RzcQku6OEl8Q6TLBttoXiqg/h
1COsS8Tz3LDkrStbtJMj7PqOaDNOCzXI6RzjGp2610Mk155dkIZZK9djiT5PfA0VT+8FOY6Kx797
0218pnIVSboubUtQ35eRO3+uqn0GYlb1qZ/bp5NbBHFC5UPOMae3AJhmHBHcQuDs38A4HHom28HZ
YS15HZolLDgyjlF4Lxt4JhB9WWCJwEKpZF/D9yKQ042gzqe7vo3+uFqz6mRDfqDprocnFjeZrHp7
J7yJiQCCSuIIR5yqxuZDzdE3Q97ykYAtoeVsNMwPE6tuf9cktnhwnbO32lpY0W89aWLb2hMGJcPm
tE3Xj+0Sms4KvvaqxULMqvC3PzhS7mY7+mh+9rx7xHSb00ltijymy4yXuPz779MuTKNAb5lsRP9o
fHMa9iBxMHqnnH5Bb9RmTGIW0mAgauxmebMNQpcQGRh4T3ApBWAdabz8Qm1vh9sj0NkrLNOaWeZ9
RGc9n9NumSgUQna+XWxc6iFRkXPfjt3Y2njc8d0/bd1xNsE4LNJK32tHHS3P9STXUqQAfLvbAU6Z
U031GB5aePfA5JpEq1SQXztSt0+RLM32Hi2MKg9WUDM2ujRcn4fPOne3EvQc2dXiySx56Gkre7L5
68Sj/z7K8InTkPQyDbKb9MBpDSMngDkTB4IbU91hvhXFhXKreOrkWemZZG42jlccVBASzoeINPFq
BkbCMJ71ve1NlbiOO+LFSCs4nyQJrHFPm0RxCo/Z/9CDfGpc88G43kW2pH07U1anxWl+r0a3MYhM
2pDCGVxZ9+TF/ri6+V75ZvHa7y8pbPcRYTZGFzDr4MUoJnG+xAkEtgBWgZqsHIIk1Wy3n1KBm1m1
npm8XItFopUCTaJbVg/9OzOjdqZTqZvpSf/WGmfVVEWTc6np6sd06cdI0YPQkK64pOMFFs1bQOoZ
SM0dU73PfbJDApeRbx1zoBmKlu1VHEazfLgj5Cz8g5BTB7bOx5iJw1Dt8e6Ym1+uKf+zXJnfHT7i
svmJ4Xw3gUiqrcpOL+tjFxiTq2N2v0+F91odktjYvw/q2JTumZzzYBZkrRBD2LepaKutNzF9EXVi
w2Ot9qCyHDc5YEx7sYM+sB3yOih0oOnyYWwTQTQFGwD8fX2Zutle9KXriztWQwdjdsvPdWPPe+/b
TYA3I2McHPJ8Cd5liHC5oKteBbTyXf4ceyexb1o3tOmZo0QAG3oiruyngHfCsSj+Nwl1/dKZrgUh
vcVcq071DsazsbAP5VKW6ddH5+qla/y9yCA28etwqGIpsz6mz4DwMc8PvbVrdPH5QuvU6t3SWyGX
AxuoOA3wjdlJHI1wzg61Ngqhx0/mxE17ZJAX4dsGq3rQ77Jqy9wWd6npGR0i6ygkIC6+g9qF3AIp
jMQXBfNE2BMwdU//dDJr4C009u520hntwsQ/MOhddJ5rvGiYPXIGK5rx8rmnTX+7d1u9zrB3u+gy
TrhdEiEaEK1BTLKNzql5TTKRi+fxXBTX8lMJTBB43dYvA+XycBem1c3Nl1h3JYS7ZFMwf1vA4Zt3
dGrQuFOZl+1JRarcLXOzt3SHdUglaMW0fmkQaRpNZYyiqubwOH8G3CyrJOM/JOiW0pfnjdkHSY7s
eyqgtZfVe6IZWYN//rwjY+ym7H4l3hDEumm69VxSAsz16iGnbYK0NyrJ+uu/Hh63gFminCKkJHUQ
+N541eZ3y0jybwgfXF2Ag71iGJz+BqAyJ+XdXHX+sOd4skhosWpF0KQUgcOh3HmPJnwGJ1GE0roz
ZdSsJMOclLii/DxMt91azFWOHIF5wA1S70n6Jl/VgeaJVH07MZCSqKd58PH8ZjDQNYjJz7yxz25B
JTr21Bgq19p2B0IM5FFhpRRJAlCzII7dECR4rSyXTF+TfsVArY9f/8sOq4o99a7uMgHUonM6yPS/
DmptKfemSbyrLoFFeGCSmH+7wiLN7JhtvLaVezKH7877UHF6boTOKs6rgWtooZQGjy7PmlygQbII
5h0B9MAJou7XrasELNo7Pfjb7hzy5eXeqD+LPRMxU31DhwZvRLVc+NsoLjt+VUegc1m76gMrUGUp
UsfPkQCg1exifUurbRDlg5R0/q4VHNA65+AkHx/sE3tCBKFKb2xZKIXUUI3P7QzrlKEZ+6fOYl6I
i0vpOzlOu7ZpXmHEYsWmzaf7n78piSeJCgCDxAqyqB6dnWEBDIcDbPXkSzVngXaZiqVwCwPolufD
cXjkMq2jpReJmzxwgtfQTDQOJ4MwICp5o4Wcbc4sLEv6Nh3uXdL48bb2LKZj/JYx7F6kYiCcTNEY
dc6CS3kafGpsLd4pchb3lzOLyN9NBqqAdVnHmNZp1ChDPUmBg0WZTPdzy13E5rWJE/h66EdJ+Kcy
g7lIJHzzzFHJ3aAs4H87AO+ksxtXzuPOza/rPz8ZMzA8yIPvacwVR536Jhz0aY8qnnym1pg+SHl4
EmHicBIuU61Hx7CD7tij/FN6yEThS7jPgmCmY1nbraUPtVQCv8CkRiv2p32ZoflOfsiPchYToVm5
RTRugJ7UPOECQRMDsmyAzR0xl+k3uQ++gxo8m2vMz8ZOGo+W9tBXnysn7ob+2zvxj2HToXDOmd2B
XUxaXEovABuYm2YqVZkgWPX68CBjK6yCj69txB4twhkCS9aqvgUBbof4vMOW4mb2/dhOcz2qo4pm
qrK+RFbG7dEv1/Lqo8zh2Pvd4WNJMgCgZvzcosX1U29C9Zwg88GR2abh96LAO8r+4BzAh0HlzGGH
hEfgVJRjW0ZNuLjM6SpBPV4uk1mJvXC1u4SnKVZDX0VKInsq8J3WCwYWlKszTr7F9wUdS4+QQzck
WPYicYWMBGk4aWn328CIaxjDyj/uC8mtxHk3ehE7r+UJHDEh/cNwS6vIx26CWaM3f+uENgH16M2A
dtWTPQY8Tfosp9/TfQRIv4ATAisQpHu4kEcs8r+tGZz0FzgWAUQY1cyOSfmTDloTuvupp51Gj0Fv
5BE99TrWKxMN5TcJW25zq3Y3he8kd9mz5x1fNDPN5a9Yd9/07pkXzRHp/+hAZfOrk2zdQJtAfmSv
HU2pO+SwtTDypBvG1IeXvMZ/y6nw32IuvrBWP3lWTp3iS0c73K5tUpccLScDhHIeMCgyUHqVpTKG
2biLrFr6dBdpb8i1POSR3Bdkhs/kPDZ0j61ciJMylK3y40W2jBPF2du8/UcaGVA41QQL5gUru5BV
9zRbk1zWOREeUgADDG0qGGcxU03hUvApJsm8HZyXs5KX9YWfLA71vkp5uOgvvshSEk64tNzuQOv+
0PvwXAbKvo33bTPXcw7UV0p9xOVlrieuiuZlz8Kp8LWsHMs8XIe4d58oyA6DxZOtSFEU28M7tvDD
Y9M4dGS/mjy/ZVsPaBe4HtznFen7aiIewI92bBIZfzrULg6UKoUlkBeMx4E6TtEjvhMLtULO6AoL
ZowgeDOhMWMScU+cDJbmj+mgjY+z7o5ug/CqgzmGdWmGhtZvH0VwOca8dkqljB/0n3ua4dQGv32k
DPpxaO6YVbBJ1iOxarCCOMeL39vIBRiUJi4gEvnZBJU/ctCEeCKgNSwOT8uFAuycR9YJTPcJ0LJ4
tp79Q5QnKjUzIYw+SPb3sWUDgh2RJPoKGWzPXm8wkKTQF2BcJRGu1zSdVJNhJdhWDT0spB0iMV7j
bQved5NipasZWZPqE7rS5BqlapHLbcbl+aM8FnxRiqYxXXxJAKUrmpaGBjMXn1s+kyG9RDaOh53b
wW3GhxSV9Ptr+8hiPj0EDqwZW0E5cCjvM/5H3m5mAV9/hVNolZHdrq3GI5L1eK0+U+oGsUwq/HtW
nycm1GM3hPu4Cx7uJluIfDgID7Y+HWSufQQb6ZHisuY2F17dVRp+U5ofwQn2igG39LlHjuOo5fRx
atpzlMI0xYbsmukoYKL+lwuivIXzXh+irEPgMYUExq1ecuzsGBCXPK5kKaVdi2+DTkWK676xXGrD
ELm8sFzMYuYnrRhvBMES3qaqntfTPusfTSsag6l7sBjuHaMabAzyry5Ho5/RQ/UEtxV8U1ZFglEF
RSwcsx1dulwWlCIWyF8EGd7B4bt+hqeiCtMr8ENuTHZtE5bZI3HXtdxwmsM5JXRx6aPzpRsEpAG/
OcmpBH7OGS3M0go4MWAlQIHl/HQrinTSuqBj8n5iralr+bRpQb8a2bFu5i7ocWv53CBJ31+Zq1dg
yPNjTnG4HKEwoyfqT4mQZAeFS34zp5F+nQINfIVcoLbDItAv+8c3UXFqI1d9nfUzxy3X8jlMkUsD
/c+qMCs7HpeBY69lCs0s8pOAsRw0xqOnYGOVSiuOLhIojWDYLsE2t+OltfJrgGGwn2uuEmghFA0S
dcEBG4D/JNG84I452TIbNsYAnWKModlBeHCvMjuF8Ty4F/4Mq+q5zzjukjILVwun+1OCIH/hVB69
muG+7Rz25/BnY6JgznMvnxZVFWn2pX4UKCNtYJG2M6vM5Q/e+UwwDHPmngsp2zDzqHIZf1BvR2El
GjVEOadPBwGiNQTMDAwVriBSMqRUFm4zPYBhZItST3TwWvs6xPRBDOxW/nB+jPN3iRYjuIi2mqgy
LRXFVD1P46LdJZUuMcuiut0mol8oc02bj/dT+8q0ryTVGYsAjGBXydc7Gk2zNFcJn6UzkFpsQVNv
bfUBr6xLqF3UtngaaDMqNulhvSr0IbZiLiG1S0saxl+ZK3CRAZwxAUbAIH0g7pD+wLnSiMiE/lFH
hck9nF9pSvx+xKFeZSvDhm2XnXiZRuEwkZ1ntZ2lFvzaJtCxJ1vGOBwHaW82jbR/6n/sZb5DGV5h
7wOvOaslqv/lkbBjLtDSvHwucfP667liYzDaLc2/rRKepAzzwIsUVgWsgAKL9viNj2aWbE09GuAR
9xMEhPk5ABn/noQ/QQRpolsbhqVVCwW7Wk55qxPRqN6yCvL/xHYgovj2tNAQpKHAf/6zLh+vqTor
BmrZ5BDJpc7Rx8JkygvSLifhIWnBSxC1DkYmHDOhzf5fmX160zubLlSxmaD3LeFfSC2Vrx+ZeOZf
1KGyvuX/pWdOl7hz/EfvLAVvDWSmyvbI5lF55EdbHWkFpb+jh2qorQsfabB7LIoXATLxx1A9SywT
A1e2CHZCySAfGjDWawotK4M9fRPVOGkgE+HrHHN4AGNlzZnvRoyP06rqqnXxVtOS35MCAmyfzEJO
iQzo2UKqw/TPWtny+DiXM/932LvMrcry34x7ZNsKbZytDToQjJx+bjw+WW4OS1HevNS3/2zlvNb4
xwQR6V/EZRNTeXqy6V8327uLziVixd/yF7O7daghDVXeEBHkGccNDCW4HVsfdglCH04fJDgWuHfx
373B5FyS30+WUmtsaV0XB2y/yr+kkzQ6sR6XNKP88ZPk6XOBrPcnFso/xWD0vN8j/yZAsXu4cjlL
WphF2+tx941r8J5FNlqmwEl9XM9nMGB+mYnZFyNIa1LRAsWu91pXLCdlNa/8xMm4iVMTbvl+a4Ho
bRPkKbyIuy8IVSCxqGrv8ycIu5tW0ALtXE1+atv+WPEM5befwZbC2VOzTBxZajxXj2vBY829vEA7
RZRo2xht7x52QZ6NSqcZ9rzOfTli8XAQgUv6XKqdagOajVoioUe6VgCyzq7MSKer7J7+dVuFYGE2
WKzDFQvirRuYIFSCOanlHt8+gUaGPooHx6c8vi7vcDUZwPLfM3pli6PAt2SMnNvi/lrW5aJdCCuQ
rhT67dNdfw72aY+0NXPmXPRoPpHvC8etJH5rSOgqUvrAWgMHS0slR4/5d9bpKdRIX0FaX//6OdTT
mLy4H/1UaroJd05DcZa526O9/1fIn4GcQb2BXGTkVZKrfu6BZTeXsiSlzMwqRPMrZagKzR1lPEfo
31Sj5Aa1mbuqeux4IEgC3blC6KBkyaBWsKC3/AuWDTkppSWX7rtm801QuHsE3pJvGChJl5j47enk
juLDYxur4hh1GTAKe4rwLq9qaTQy5bOCbHvRa4J1/jiSjnEdYxjJIpm4EkDkfKb+HFM6Jmqfzfci
wL3qwTMHd72l6AgxvcI4/voguUf6B1hEKDqbzoDf29qrsLn9+hLrCteJ3R2mY9vdqrM2+Q0NShtT
kPuVdvlSbzBU1Sir0ryQBq1uFKRoiOBP2b5alPFntq17s9QZEhhStAHCv15c0LJlIszgk5OTZB8S
7cqjhHR9UPaIqg8dZey96wAJM8YG/IQnZHdvR0YTtoAwxYgK+euxd+0TfSba1m+W1f1v/xo9RmN0
hufy1nriAgLrVeu3sxvYXhDsM0EW3t1FuPtxtk24MQGQLGj8e05qS6FmC3CKodFH8gOLeB1PdkKx
/0Cm9WKchrKb2CZa0lFUVurl+GmCZzMY9QuvsVXjcmxzCNtLoWBAr+ZyYqshD3j+SYV8U97F8OXA
miMnoTaMoiylzGd6AKxlZGzAylGfNZlnwT3DVnnEKBUXmQLN2qtLgRPHAGqmoMS/HgYiX5AuyS1H
5QNWsmt3A7lyp3Qxv7ccX7f9Mwib0O06ZJARXv2PQQe9dCzqHnY4iEOCnjL9jNnSHC8q/nBpSC7t
0rnBEFAEJt6dRz9O1ND+R1ePcQqzx3Qee0TtEo3zb9lOgix8BLKgYNi4oqIoGTPWiy6jLwQ3EFGk
KaX3FkY4ir2X9uN1/cHGpF2qnn8cDxPl0hwE7Uo2yRcBHdGaov8xb8kRpSChDsDOb0d8w9J3y9Ai
qxQAqIonT6rnGKRnj2xeTKvnSOstMGAWUGKoFfr3Vm23x90DbNLX4ITa0SsfzEbi8MxPnKiUe2y1
RR++jkIfyVwhBwBusF0A5eOcXjXiLL0NVNen+zqAf/et/AJtrKZ/P0o2OaZVi68lRAGo6qa0Bbjh
Z5oIpM3bTogg7EO55M7OD1vfDtcj3RxvXaDrKna3Q1uQTtP0B7IJDjV9IbVcRuAUZU4NG3/qFZNn
OQ9wb+noXl2PHzSBEXdec0Z71yrx/Xll3kNGRz/Z0HxkVisV0b+haZf34vl3z6JX8BYputqGoP5P
2yxhLXBAasqIlmB+u3Bfg7O3dus45mf85g3PduA/MtspjVY1qglHTSnnuMEsJQb7K6qsLRl+ILN/
9F1dYu+UWv6diuS8PVsMgc1rm2uR9ObbhwxAyfg82nSVKpxUh5bgWqCPN6yv5inUkDgEEuw00Bj2
asRaIuRf4YiC2aK420JS6twn3f5v7qYK+c0GMbDNednjR4qA7zFsfoENu4f9UDd2/GoxiTovcCsQ
Ssm95QoEdXwoMXfnZtmCylMM0by0md53HAwjKHxLC64haaDIWHTJKhPNk4vJMnypawHS+OvmxoEF
ZPdMNs0sG5GdKm5tzclgOuGzuk8o8q48cgt3tUmUxfq0erZ3Nj5iV9I4j7j1m5Tdgw+amYIcrHg5
lrYnUCpfQd532QnD5YuN9w2ZqGCewxZCOU9oR/l0/f1KTSA5roDSKkKQkXbTJBuYpDE5SyXB005g
vH9CYPeKblmVWAJpmI1kGGDObgPYeAu4p61ZK/0z9ppth5U/tmIXAtIZnAenk4yVNXnUocduIeqb
IgzqKliRCujRaDuDRmaiQZEDibjaLFqMNDfuBcTnfNrYvUws8dxyta7w22UbXMVd23RkEHZ7o1kH
L9gHfbKrT22SsCoGH8n6wGzM7Y0kc72feW7cowwxx6t1TbjLIIEBq0sXhxHnheF14lOiXllBWQ66
0oQnQzdCR3XpqNm15FHFDvxhGLk6x3GJXyKHJAFveSsFzRDU44KlUiXWdRuXtQTGkfBMuFzEyT8U
yFu/d9b8iPR8yYzXXlunMCqA/MxiNuCA3ISinj47GuZyaGkJfBL9/82apdKsWLOew6rHLLYag9Ze
CeAf0HGdge3YP5uV0zL8n0KtS8GIJ1LmLWU5nXW6KpD/B9u8hNITi1qrC3Eh8oTLfSD3D7gxk0pb
LrtjYqnPhLevdu4ee261lVjlbGCqgQXr/9sR16/EdG/RTzshd4te3Msps2n73q19CwC5fHnvsAR7
5cdyNTLuLES6g1rXsMHYY10HYbHup73CZSpcse9w7E+WqgR7T42VoNvIt0N4VxriV93dpwC+cxS/
LHUGzuWcK5RtAnGWBqckG/uuKqaOt5Ww6/ZYoZXG9dHFz4yEOnUZe6KpoLndWohaR5XHxrbjhfs6
T5O2VRSI6jbwpj/zj9WYw2mOSecpYepEVbKnsLNhmfs/TibHyjxZNscniPhGNSF2K9tI5s/1s9aH
/z0+bQGZ4AY8yE4m6x5Sp2TQTFiRGZWk+L5GI6I6HMqyXN40akpDDjbp3f1Xt4BIGeh3e7TtCM5s
qTBWp49qmBpjKKMWCNn7uQbioNbW7A1rLw+PuZp9MCK901MhgZC4G4+QSslth7zM73WT1ulmbFM+
WUeDkh6wVRPMzb/Ditgj15YDFysEVnCE8xIwDjh7h7aZAdnpBz/3a+gE3Az8p7Va1KpG35BEdvYH
U3UAz6hx1Zu5LDY8rLl1qsGJjpMgBK6PCsydcxFMw+13MqF1k/Zo9wThpSKlnXImYxI79wG6EZCK
O849UIwu/pL559wecmW0vQ8ZIbGRFslHFtk7wuDISeI8pind05LgRlDutdgLbjRiMFtt+rj2Cf1U
rlV597SBlLB0LHfzoBjolwfSIMO39L0zeNP1d2N+HeZhkIic1UBQOAkdLbXUDH74JO3xTBmeJkEH
eGy9GwxgTnYZlpdFAJDE4Kva4z/13rib0cR+yot1L8oMhCC5x4mX8DLFL/ZH3NQb/03edUrb41bA
e80s3xWW2/1X7HurI0ROa1BO8E76XiuJhalFVsXUJZfD7dIPh9Kw9BdORaUL14/dWly4yctdLGoE
QEszc8uAdB4AHeT1aExv2RZHYpWy23r7BBJ5I3GTrYDyH3JgRaDTJ6U7siP+gRgqhV9wrCT/uW3H
DUlfHdVAwEI8xVE5hq7KmRLUPPeG0jr1EmEr+p0PNqJcmWHv4KwSs4k+6yny1kvZ0tN/XyaL94Yw
M/ygbhX7T2hCHOybVVm1zmj2O5wqoXN5pe2v/iZtY0qi3XeUtgrCuScjSD1VArChw3let82Og4Io
eMhtYGAZ3XEEdZMEN/71XreaYjJJItHQVrcp0HqFHh3iNQf0vf1xk1R9rrDsvrDsjNUZLS6C4376
cyu2UyMdLxH6MKAVn/Thv0sL0zDGGmxVcxjda0ynfFAbrtFLsH0Xvk70/xkHnh/N9qEyp08LofYp
XHzZXtLJvHC/lhC/IIg4/nER29+9UeMQnRFoVat0rQYGIekMH+jWJdc0neLGsfv39FjMymBvM9cU
8d6l3JapF1YMH9k3vL3Oyq1+R1Bxwzk724kFIoWu1Py1Vo9/66iU7IeGZlwKBE8DJqwevmazjvtG
UU1s6XFo/mPAUFUO8o87jOnjkjAYywaoI5pjFSm3G3PhvR+2p78+moH29jfCDioloWw9c4Iy1M6T
l61mNjsWUr34W8k5ADx/13amm4fDNXN5qXrCmO9wZa41Ur7E3YNGXwt3Dx4mlGaFfVp1hpjwRnYz
H8DIFtobsSr1AexxpDBuPPRRuhItrtS6tCEeNFlIgrrBpNmCz1ycA3W0iDEVge1TNmTVWWkV/Lg9
vh5dLtQAxGctyLLBHsWPaTxxEFoN2955Few3pSL08/s4zGe4FKvAh/zLLOSmMiySTyVFqvzCG0uG
Ob3sLbmbxuq9zrCy9qxlP0wwWvW5wZA+EMG8U0BBTtKUDKMzdJ1PAUcO9xjAkf8LoCkqD3sax/Pb
ewFcH71olnNgaqgfDQ3FT9rd2JtIDex7D4igS5JqtMmfXo6gVuWonpG1aY2HIZGl5jbQOmGhqxlL
mhlvbaLl0g6JZaQuzwNUp5Gbd7FUFiVXjAhql/LKop3ZHNfvlqZoYfuH6ZoJxGDJmCAJzg+p+jQg
+aoLFjaaWZIAIgpwFtwhLJoDTsFvwYasGgUBeBiCsgX34zooGoXsBFcG2z+6wPXIkPOhPEKQre/F
tVhIuuwOYbW1PSH5Oug52xnlY5tfl9vBNCr39pK/t6UuIBhfOHyZmModdreKksCRl+odIilO2uDX
fGvpGM1DpIdCWYwczVpK65Hqyp7sJeLYawMLKSsjOulaisyrJ+ztN+Qo2RuG4RI0c2T2R3AnXvok
xbyIbueNRSPO7akeBNozR7F8AHlgwJkmhA5AR5MVysOQNpTlaowTBrtxIFR5C02Au55NI5ZgiyFh
s3lHWwemNA6/tFT+26+Ej72qy+Mu4eTUXYjQKsK67L30AaBXZ/Z5fMnRlQpDIBin7BYlAji8f7L6
QVghD0PM4o+jgGtOkPQzgsXvS1rVWTxjzLdOtt790+E3XBv58sB7pPdIG47pVrEbPT/4fPVwrAGe
QJ77y8mBEuYm72f7lj7UZEY44N4Pw7nQCrTrZZob3Kkm/f0ur7JN+eL2seZj58XokMKQ6wBqDdvg
H6aMPH4An266UKJeY1IpBCtpwTx0QG4ZmFBu5ZPhmfOIF4OQO5Vn9AW8ocfgx0Jot538L7fBaniG
t5Ur2zzFmni0aoxINMyysvTcQ/Y3/2CQeOo91tbrHJR6HjdX9kboYLZcoS8lwHvXPF4wN/SaWdZ9
KMpbkqjrJytnYi+20uzq9B4YNoHyxoI7OkyDUIQ8oQ6fzQD+/m0gAyspOXgwf27X7bG6vnOkXobV
y8Obg3Irh0vKbKdZ0HtAr21+drVLCStx39nNv2qQrKORHhiXOhSR2sFI3F5QrSFkDF4M31IuROGg
5uxnq1ooy0hU/7apVcMn/ebdwrzWVO5sX/+ZEMWtAnFvYhm1f2m9yVp7CKjyZCmUtl2eHgm4Dh4H
mCIFrD7JSq+aCl0ofPR/Zba4nHmLqPn3t78rMqcmaN3xagpa73J65rHH0a+rvThXAFotxWqGIm3t
ERaxJ21Tyc8uUfaKdtJBHPYYXgcyG6YQKEXUp4BoOMZ6tgz4aziEhfZPbQpJ499NG1yAtWbD87Wq
/M3hrDIpabdPL/Zi9B5aLrJtWpujt8xnitWXkp6m++bGL6BUte6PFlSkfpVIdfItJt4Yfhz5e8Ts
wXjX/4FP3Re4Nq1nQ1oImJJfgC+XIQl1v4n9Sb5pw0RpKgMeVxYQu6ti5C9v7w1ReDaC+E3tZh50
2E0DxXKT78LGRa3FSSllQFxxh4nK3T4uQKw3gCYHTlQe+AJp8ttjo7p/o+CvGJoOdOpXhafNsSeV
78pNn4tVdxZX3s+7oxM6HWtr7oFFB+S9sfIuHNmYcF7H2NB8u9su9fv3t5ZEJQz+eGmr2PBblR0T
FN7BpvdZpBZe1l9eHDNfdiANE4w7igVQhKnLNPdW+b/By4AntLZ4uUXXJIDbwK3k1PZbcX9e+RIp
H8ClF2DB7WS8WyMSACkWQxYEw5A/pGyjy7ITPYBI/qt9BwZBGbxLlDUZTuv6Edlwf1Y7LScR4WjL
DI4Wf44xhV9OS217ZqmcLHuw8MhHxEH1qaKB/jCN01S8Y/xcCjQ3ZcExeAn8LSlxs7mQiTJhH/IT
V0Z+4UIi7OpE2Xp9LTjOeDzhecSHmDZMyYRjIWX1pofEWdAjlJKpKVOREDkNbapQp+jjeueJT/Hk
YHr5jB/UxTqG16hbdJ9Jncl8sJ5J01wE1ffttz9ja2gP1hwGfxYv8GcQQ0bLUrFHWUhw3vgRJ6sH
IVYOSkx0MQ2QZY7TD/Kji1VFwisB3/Gwi4Nk2UdDhVT9uyau6QXSLiZRmB1W3LAg56zXvc9o47iH
No7znmTw2yPdoBOJuHuavh34wHCLKIU8KaXiBhMY+TImJx2KD50BWjKNwk4C6xA0DMC3Jq65boVw
bMGNngIVohnyo83nkZNAFbK4uI7tbTT2FJ8+144LOq1bf4SX2MfTLzxjYuhqwbLMXvxEki0HOUbu
6p7TTtJdSn8vjx93MWoA3TTtWcgSXrov0rbmAxJzWcpoihWmIEygq2I78U4CavJPuWXzIHHxa3+Z
X3T0t4me0lotOBEgynqkkzRXeswikelEHxn/YmfrbATwJh6W0k/8NhYAIdsBTkW4oE/8zeDmu4Mk
ueoM3Tgq23gCQU7e0ix2Gm8GQXzxl6thaQq7U1wQ30AVArhCRt5kWHTfvVIp1+cA0uFwMqmQvJSz
GcTaiIWWhQxr7ueXb8I97DeEb0j9j4oUro/B9oQYMMmTpQ9NVmkHTssZMO1LQjrNwHP52zDTz0hq
lRLGlOBb1SixqCLEFS9PBz4NjFaxOX/MBZbx9/tEe/Wq5uTuOsIk0elv/VcwT1VBf5gFUjCaFGTB
+nTnxJvduDbPUzsvt9xyspnqlku1Q2uRVoiRiKFqZlqhBGDy2AkoLWNzHLOzXovrmJgJNi1jMfQf
NcSaHrIi6Q/a+7SOpAhkar3O62QsOweuO+Hnb7k1PXHNHCEjYQb1WS5aUdAzBzHEmNsZt7/KYXhC
NygcBeUhBlnlWhXvVKTKYux0xkezIjWQwFRajUhQ+JL1sbxq1TXYNKT8vYJc7bFelx6rfKy1WnGX
1vtLFlYO9OeLAKeifRQNhxs0wIrqfnzxBsld0Xhw0PCGFjGlZ/Q0vJ1EJSf13pS8VfS5y8993/g+
IH+4gBs3+2X0iy4WR0CBFPddLMpOCgCsItJxZu37KnMatef0C9iki7F1AcSEGoiUqbavSR1Xx+/X
Pps2W36M9H8U62GHoW/akYqN6psKVMJKhsM/KXXXcM3fP77M1+svvVKeRS/qcDLnD50cVMoJ+AN5
nTDnBUIIrbr4Y89JdRtYMF9sUm+IebfMewnJTR436UXR9Guc3qRfHCyvpSlQ0Cu3T9MQZFtfKl4u
EWGTNfBzg3SCQTHWfRY5wnl6Cz11al/B698GmjPhu1+3WP9iwp5ivfxcCsUOfzhJQ/Ue1v9/6FFg
HJOohzoPrOExAaly79R2yORvqwGcxBT9AZOBRsEn7cKPgG5xaS1nZ3lFKf70oRwesYR8n0882pd3
WsTdvxHw9gk7UvWkRgkWoPd5dRET4J8IhSlsnlF7uXoRnNMpXZF1Q9dGjo2IFC+DUqscq5bx50Jq
t5i++qJRl0SQ9+iqHojpJwxEsIwbY0yKO5pKSfI2uGzFqBCwPlyF8SWMxq0=
`protect end_protected
