`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
eEjJxT2qKte3LFVnxmMKd8xUUNVqct2KJM7rS9FOKt6ZTHUKUMbSAYFSPfsvamvaEh7gwS8fbfQj
a7MYJ8No7yGPlLA5he/lU5+bpo5e9EzRBwgVpywfVzrFgJpjFhmm1RJSr+AMDz/+OCSF0LL7yWTF
r9ElKOYsCuihJ/beMzvQLIEIKsE/1xatF9pypAQFzj8ILe+7E5FjmwobqDix7u8hQhMQ2CHcyMrP
U4Z2s8wNTR1eRWcUuYdA+wgwnEWVdT+DutoUYRgTJDTB17bbIHL0T/HnoVohLHlyTGDE2GUJNloO
d+lXvpkeA7Frl0OUae8CHzz75+rZGDvHQfIM4Zv8axQOp90vsjwfi3ZVLyIv00tU1M3UhKlCtRdx
lfoNIgn4iCQxDGneNwsuDzqDK/VE5jNd4u0ngb05ktLdhdqHg/XXweg4pjwCNq4UjA9ZoL7/cnmG
+jC51Od3UDnVo2HX3SNMdWCxiUH9jDLh2EjiHevznSnD23d84SjQMTku7I+UzLFXbJCyuEsvdTOm
o270k2lY3sT8Kt+CHb7LpYjxSRPeq0nJL92CYUl/6n1sI0VKcJXmBznpKvV+crGZcmdxw7sTsnFR
o8ZAVYvpfON92jo6ajepNG9IlIsopHeMRHh9f6z3xJID8XavjAHeS/NWCCPfkfPnqLBRoEQ1Yo9V
R9fzmgaEjnPqwjrt2wUhzYm1bYYoHi684l/4PDAasmmLqNo9pJz0ikQkCdPtouR1jIlXfYvtfv+B
19HfuM0uj6QglS82Uh9CjQNBgYaOVj7+XTG+A8GswC+UeDO9XhjKnRv5df0QkoVe8fwC+W201udf
XMPzQfYaLB0Isg8Ecy1dE7sz2xblHEeT3tpxcO0Xd16bN99BCCEBIoDHn0t2TeJaGR6xezC7sFB6
38OgU5KNuXMiwF+AzlF72G2m8+62UB27hBUiMo133TaG5KkH3uHBhYPO6W/PO/SAoWkCZ1Euq9PD
GMo9usEew5dK3wUwn1nMBTGjH2XY2sFfU4KtNmDVOnuDhggylnVFwSV+FrHM9Z/FinhxwtVMDiEm
AkabCBVWU7O7r6sLB7UEgP3H7OxFJ/uyrLF97GVk3Go7zSigukgt0NulbkB/KlYFCrhJHoKJW9cM
/55MHsM593lpLxDnTdstdcY2ITrCSVJVD37kRmPCX8jtOK0odL614Y1DJM4PBqPqxK+UE/eY5Yy/
mzeW+2lbPiGgvvZ2LZ1hoarTCqFga+lHfx5iboahRRZrsgm3WcB7l9eFrcfugo6AJATdAa2nrUOr
Izpau3CyUeaS5J0yMhYJqi43f669U7YPDhkoFKnVEnM3n7lqlXufi0XvGBLeWrePPa7z9Z8U/Oj3
1h24bhk6Ne9riAkYj2cG68t/MjRZbq1Br8sw9fAZKkOFVINuIsh1rLNgU36H4FsVHcVBTlya3lVX
Jptjybo/eduO3TfUN8Jxy/8xoiijkMqQDv3lHwRVCZKuCf8+0SzOqQpRZNuYJVGQHmnq735FwKrV
SGbzjqcghnRtmQDT5xI9zL7QtMQ6twUkIFCk3ZLHwNjoJ34HtJymxyMx0LEBoVeL26h0V6V5F+6w
XoipMb5nSlQppyG9kKXiK9UF6AZwVsTlu99nuiM6UCGRJ42hyRDTz+r0fxHRhwAZ0fSucpV9nCjA
caIgfdisFfbWFf+BagChfD4ASL3iBiokdoAg2VVaHdoE0F3+izBizZo9oP77FBe3qaEyH+9M0IQ9
9zr2rN9NddjzYMS/a1/W6zABy7eJNSIzgryu8fIewxQijMiLYoh6BzyRTBA8NAzLuP8PEImjNk2g
GvdY6ZW1mFepUOnpWRjHIOELmLI39La4toa2Y5SDoaAB808NUFdGQ92wtc+KVZcVa3FjGqDfmdFv
BDaLxH2BAnGccAJEWFjZtd+jIUZ6kepRqI3d5vqnqhtCD3fCsCptjva41FwLWpdCzvrLp5NLHvwZ
4UCp2Tu0E0JQF/cwyDREMm+cJE0HVntYyglqVw3fRkhKrckXi3bpFgNGML9yF/rzugN+lFDWLIiD
sQZWjwedZE7kISDMwNHp89g0bd6i/4FIHt+FaSanYB0Zgfj/pt7WvWhcMoLtUaQXM4hU3VwEKj0X
KoNRA35gewbHyXNzTHdZltcpIZ8bsWq3RzfKJWJOAy9UNrJjHB4JsvB2A2orAwZ5KAx1Y8rFJ9jB
h+anIeUUaQIgQ6FSFz0hLGQggWpe5RPq3yWzSaysN9EF8mhiwywLtMe9NfEwGjPVQyFvwOFgZFUb
Iio29KTmk7b+XbMsOeShcYAVZyMLAhLIaKLhopiJV0Br7I96zF7iugRxvtB7eCzb4t1WdsVSWp6o
nMv0lx/QTWEzevxR2ylA69A/MJfTAlbnpDN+FRYpgpt+5xtDgV7RJGPVzn5Oe3nTsj5vwL65x5fF
rpg0OBQhK1YLzQP2YrD/poWe4Pp7dEptIkDrAalQtoqxsiXmyjMzlo15Fqs7ixxUJHTvGZSxTbPE
HfT+1GGqNSIEtzCkOLZPICxRGLKWAdD0mjWO4udsqYlhL78+QzpZcvvpyxcvRCzJXRMvfTuriSBH
Z36HcoFekT8BOvHY4eavgs9qzxcfYHss5Ki9fSVUKGJIkQiGfqf9wMrk+nHggasrg3x1v29o9scC
gBx2zM8Yw9rVnYJA7Wp1R0k/e2+AQ/ZOFdmzesDdXr0Iupwi407+yzlbxQRosxeiloCe7Si9pxDk
yYaPJm41Hv4SyfkxVl+2fJPS0754F/13cIX28xtPMtHFvQ6ncuwktnOzTF5s37D2miUDIPPLinsb
fZjdJcBJ2KXu1Xmlwm2VpCnwRZQUtp78arqW+x76TJmHcpoX1/86Nl8BA7mGhLvtaZoyfs8SbGt3
hnBCTS1UyVyN7zDVQWfYr9Ie5Ht/W8+awSmDyUnL6OEmtu9QBQJvI6zOyk9zfFMjsmKp9FvClFnV
/1QURQrLoYWPiRfTVASFwDNqR2tsuQZJyrrCBm51VglE9pdCDNS9tlG2Ac711vkBhSu3nYBgdh2G
k19+HW+epLvFYfCz/EDQn5lnaUnztendIJWQ0VaWLDE948DfX8qjsyJ2M+eA+PA6CDr3Em5XMfr1
YrTBf0jc+0FTtlJjIEb07a1cTFsXvABb2OJUknxpjoujVwfVsBcJLW/7rt64pbslEAc03hw7XhZC
ZbXYFgW4415C5mWWv4RZ63Gtjdmp08eHBbXzMbam8Zd7kChQsK9B+2JQshltuxxlyK9CGS2Z4bFJ
CpePkKcB8ux4Lye3+XrkNCo6F2IrSxLo1HRML2OFodq3DBLEsqIwf+sKEWqRdV2sSxzmxKv0TFZS
jtgl+kGjLZ6j0mbcCjYCMLKQrh1GQF1Wqofolz4XvDjmpgogp1fCTtzuGmnKMPzmywGFoi1ynvuY
UQhWbI6Qa8/Ea7r5E1JxG9Ef7gjoF7Ys24p4sBx4J1QRRsu405m5+BfnvYne6+UEDBWxcIoZkQVJ
Ux26jug3F3PGDBdRM/h7fylxuwV7LwO3BqfuIuvn5fSsR0uRGiv1hObScbqW7F5ZA/LSOY6D8+wj
DmwKgnACNv7d5tABlt/rDT/CUE8RHCpSzOC2BmXcxqXK6a0PxlbUxxmPEzBQMOqHIqqs0RSiepeg
YTg495XieWq7Wi1Toir80L+V6j8HEmEvYvcYFOEiGoj8+K7Y7SJCHO6fEZDexzNeNwDsKMtszIRG
G1INBciNYWUl0/dZZQSVbPUIs3ee/X/Ji5AgITjnwJpg6MleDVcxvZJierdYLtqG5aV8r4p8cTY8
9PhojYkfRIP4vd7IVvYn6wQDrhXzckhzofPtf9gCQF4NOyU9NTQ1bsC+gY1BHx5YKCBI2WKc21XT
HS4cqlSCjvBwt1M9lWG+Xjm4nub40jp13LboiY0/T1CLM8Q1Cpb9jKQ4Yqy8epES5lJvvyxewMx+
g5Ql1Ojw24HXcNqQ0w57xg3L49swEaPbWep98icT8QPLuP7D172AiFsWRbFQje0mmkEmyRujIRvE
o6hZqoObRdJxW4oMVrIXCMQD60pySUCSl4rJZlpTG6RmvU/sOFyCxN+541xyMF8P+q7G65CSn0h5
ViXCYfqOixGZdJ2no5KSn0QPXSuLHBIpRa7BeT8brr5mME7iidUnXvW71MBirlZDCwZu2bIgXNvP
bOQgVIrInJMBRObvOhA0pl+Z19aHYQG48M0l6rs5GRoo2+wA1s64omXj7FBJ1QElz2WO7j8tOfK3
g+UhbCOMg6zeGR3cW+Z0z60LCxD0Nrft0vbtj5Ev7BmBYJ9WlQDmoj7WzOYCjN0rGQTrDlV7IsGj
Q4ev4QslVKNs4BtmUSEZ/UWznOWRfDhhD9cadenYDJTXwGSsfo9VY/k9osZ78GwHQYLoQImn1qpc
fLrlzXBAKnGcxMAFNJvnUC+gQ44P7ymNVa8y5LPqzRc7kTI19YZdnl4fFej/zV0KuF6k/LQom9Zf
CowCFeN+T+u8BhclfyM4pJ0FilbCbswCuUhQQA9C9Nr7FyhsAy3hJg+OOdtyWzd3UUhrONrXZmSC
Zeba/GygW0G8GncMHNUoi3Uhgz33AJutGg98m4Gxzz/qVQhWu6FMiJmYaN4n+YwxsFKDykVwhC6t
w3Z0mY0SS0M46L3ZzoeIauk/yg+TA2PCTgADOrYGc2F5XcZ74+WDmlLDsGPKjiuQNPAxbTbsJXsf
XpPbe+ItERGC/0kQR9WoQ/IjCoMygcJs0ZBpEXHvFAzw07aW2Vuw+kwGbBSR6XIDOZyGQzCdYwA8
jF2i5UyjsmKgH6yB+IbGfQlNi/C98GmBRNkQUBBeTkJQZjqggdiG5wrKxHCCuTO393TccySLV/Kn
W6JyEGYbhOhLsobt+uLz+UFJc6gwbpVVpg5aIVbWaicGO//a/MlcvaUCE2erK+p9Z69Y4m3jvKpQ
f89dJOHikYxgc7Dr1Va4pftFsAXx8UU4sIusSmRn80G2bFCOkrsHzJHR2cpP8he8ieTLUOwVAnpo
Xo8FiN3kbb7vcaIPbmONx+FDik1mcXzPYRAWdUQ7HMOY1EPu1bdNe1MtVA0k5I0xE+4QWsGAR0Rz
da2MFuA3xcpT4Kq2pA2g6/KMFeiVwNSUug8UGpyB5r06HaCMPblWkfhNmpKV1V3e216WI4W1VyQU
KlCKpngeSPYG/l3iTvCjn9yeX3lTuj0CcPmMK2NuvoGR2W0wk+H1/r+Drl0AKz81vNyoMNVlXBsP
bGMRFGmsk6a7bVurACXgouPNeR48V1cqfAOlD9TFJX6QeIBXuSvph4r0ocJzv+IoW7qpQ3VwdWlh
px8Hywpeh7fBr9eBjTbrtUxc4PCZR3lnrIi6A2DeEQyJ9IS3XjvJs2MeawyYiKBXWlVAqKVeWAEu
uP/deHlLeIk9VmLM741AqUOqWB+/h4iTeCg4GdcMHlS2qFRAAKsvx7zflJg8pXAwZTZNKIzTDg/v
f7TnS/DKhgfJ8aHL8J4qBbf+qdO5o0ePwQJyeBu8CECayoBHT2NGwaybXuKccr9d9nyi3qbu/TqP
PQjGhZG0z4m5Fxnql+h//n0GZgkiyBXLeX92teUclRDCrvChVhry0KSKetzFGQQokZy2CwLCV/m4
ZOwyJRYrxviiopgLQg2l6h6SZHTL4JYDbuOtZE+K/gWNUn6EKbACo2QzcXAS3CY/baP5UIagaacv
Nxysh+tMzkg0ZPmQVJ2cAbCIwwsJ7Dl1/2b33v5pm+HpmvFSZW/HpzpBZrFt2szo8AbCMw/dPMW4
XLFiC6MUyqf2YA+tGYEh3KpF/FJBGbQ1GCAns9A2VUmEeE7OysjdVpxJq7rHp8FT7BoMCgNw+neF
c4V+uzg+qOzxhQqPUngm8yIZOUwA6XctAjEcd/85/D8Ou7Oj5GIe1NPpZXGv3FUo5cxa8MDSI70C
asuPqdSj2AXOrCIGP+cp2i6Hn41eviMAlfteyfqATVQWdRhK7VRhraBhfqOvIaEhToC793fmJNqj
aJYEAE9kdoKk9G+Dey/eV22U/slnd02gC8WtVzGf8kp3LmoRUv3CSaufJLqOstOd33uCVZPLOZCF
/Ip6IgMRaIRGpWnwn0mGB3WsGniSAjAbR4xBhLnlig5voDOvVN0lY9ifm7e/NUtsJFcheJQhxE1p
Pd6Ai4fBgy1rztKbTrheHhJs/fbn7xvM9rcsBRmN6mXvgH++bsxvzA1CBAhsawk6eCHY4uxiHn4t
U0DO9Ow4uO2owF7YLmNXzDPbGFbRysthOqBa+CyD4QwG07IPBFe8nOT8DJ1W+djV8hmrpxUfwyvs
XzjMbhxYyOnyjw3pQ0G2ciukh1FW9iA89iVDGOiB2ESDKdnp1bNp8xA7Did+9nQSiGFxRc9I/3wy
vRT9RO4PQr+WQmDh3/pWn44W7m3Pch1bKb4xGv8gbRGI7hEFKq4kNil3P03BF9o2HzEjD7Wfr/PI
n5eJ95hncx1dPODiKok6OBswa4Q7XbLpiYHhHWtkzCRrr7xAlFlRrM7rSgFfbuJzGRV/Ldmte3L+
Q+/cqfxpLCcOXYqsoe3WlxX5ROxpJIpDKtrsczEunODDtNq+XdEHT5Q/evNk8Gwe1oQMibX9j/Uu
YMVbLnOErxkY7dWupemhlwWTKcr1wD95TQUL7MF9xLt90LhAzsM+ulBMKGvkEiS44FZutednyxJP
8Z89NbBG2E7e+CY6nU6RfC2QCCe8DaNE5E/iTUC3mHG3xla+0etg0DCqiBKm/nArsNQ+gl7IQPF6
jHbXcJ0HIAE9brzUbMy3Efmc/gUCPlZF5Z55NJVdE07iQ4/gmcJYeTcZ6mrhDINVos+qZ8Rx9yCw
yLHZymG599yhiZZ0FLwGb0MFEajinm5HHjDuKDhbRcb5lCX18///N2fCWXsAQe0Bs/gCnOjlfMsd
YAFKciT6d9ZmX1blsTaxoimKxeZs0X+dwKfUJwmwdkYB8DCPM+SFt7MsLyZb3Pl7/l10oQ3mIW/Y
TkoOygaU5FX+SKWRtngwNr+rme8DPCh4/wi05Lu8iZqTphRYHxZwiNJ6zKVnHHPcsNkhNUBleL0L
OfKbc48JBJwGcFP+QXjwVKOCxRC5xv0uMHiU2L8qbbNrq5sNL7hAFMoH/Z+EtZD3zoDa3dgyTCJd
YbHrYD+BZgMmZGpqEDN/Yn7gyVNgkiCPrglevWaTGPAQ+BKK7sGz1b1zxRfgQ8Zdbsj3ufKb7B6Z
XmY2JGvNUgCkPDjHwOGDcljALfWUmA6NpOQHgqvei5PKcAb3tb/gf8/NVNhAwRKfN7UjXWtZIrgh
5gGw6hyp7ayBokJUgZFQTp4bqDm9+Ynx/4ceMwezkD3RzivrSvHUzrH0zTS5qDFphN5Kq5EFt/eU
kcofRSwrtHyNeHOew/mXvfLZ4te8R9MqePGEgaYlE5I1SlgYSTfKb2q2piuyQmB0OPdCfZwK8FkL
nJ5lnvoZmqtb02paurGqVAAbQxybivxsSqg/G8Lgu8Q1Ll8aiD5NtC5pPg6zAJc6Mro5wu4FQB/1
srb8gYg8jLFYkO1kRMXOPhoLAsHgBDnvUjHJxgs7kNRjIeVhLEyptEC/9DfzMJecaSQC9IOOfCLr
umvVSVphY8siChfIygR1vZ2Fu70OoKYfH41nweGmOVaoCIkVTl5+MVRuy2DtFKvGbj7IIbIpQg4V
3lcotco9KI7CE4yBWYQlNfmSe8IvxYiqhnENeXdHPEdl4i1frPUwiYYdGdIEH6YnI52R9mx8Ng+Z
vn1dfRtjjF84//cTgaJOgv1E7sbYc9wCJOjB0AvKh0bulSRoo5SokEyXDVz53MTcOlyhC/A1mY7R
1/wMxqxCPdF9E6nzbnzUIr2SJaqkjfdX6k7PgtKIo5yzd3OarEPJ5YjQfLaUkA3rNfNUFEr+0O9C
9iYaBDR4NLQxR5OVxl7amO43c+NggUI5fb2FpBD4LCIZM6XPStrPUWRCIBwDkJIg3pXpsLWVaz/N
ufVXA391Hc8i6LGNjyhqjBu1zb3AFHIVsd91VCBIRk1GrJmHTiBpcZ8pF1hpcl2heNwV8hr0fxEZ
aXV5Tf1c4x8DxST+ZXnL9taWykM3uU+7jGIgtPJ+FkA0sACDogGRa1N54ULXl0qtyIF8GwIXOsTQ
Df/y90mpdK/NM0wN7mPM/2950K8AzF78eTi8yaomWNhl125D2BT/0142KBI06tPACfvAUGZNUL0L
NXVM6kd4FT07ceULSB3/NhfpDRJNW2wgKfRc731PfIm2z46xK1Hm+u06Iza3AjJN37PCB0z/SqN/
Iil4zRZ/e1E0sF+Sf5MV14T8+LdcuHN/M6L0YTAo/D86Vdaj5rm/Hry6SByXHMW1gH45Bt/hPCie
KOxr1xg6Sy/xAd+Fw0j1pDU1wySuDj2Zxjib47BezfH27WYWd1S0I8Xb7g+Dbf5PQedCMk6REQv+
nl/H4VgOxr0/u77D1MVGOmrxluUysbPGbMAsVj27RSO/npd2kF7we2O3eRBN5CF3vHHOTrf7dfNS
HyjRJVFzQXmkqZ3cxk/QwhYTNOe0afIcEGP+HNX0+TnlwG/iiEP1S7wUHf4jK2oLpRc6Vqd50B8G
SgjVGRL3a8gHtpUP3w3kU1hf8fsPv9yy5ugDqTRXGlAE9mjAOwqJONpQXlbvWJp8QA3ytMUNeimm
Lc28MNZy45DxiNQwR4qefMKFwGxESJY48YB2NIoMIrc97oYbxUFppT5VjCf+fwYf5z5WSxkgm/KQ
Dc89uCv+S0Aufj4T4ylgbl2HOUAr9zYsek1zMOt2eO+FWuochN/PnNu7Vqzvwd6xVNGjzDCU6yWA
i0ssUQn0Tcie7BLCMWXCGFdJdmVa9QgjfraxWJyXxWT3D8Mj6I+zHTfBz505Ka8hzCz1rx769xB9
l4vox6r2+Bh0S+rmSn6fc1PJ+cIlyqllptyVrtwCDCI7+qZ86UR+LmRaGQfovRDGG1TYMrl+1+0H
iqEi43Eiq8OjwwxUU/zXzowx8Ykb124WksWfYSJFeV+GMXywc8IBfV+WsFEPgk5qN4yKPJQHGesd
AgrPdM6OO9qTnWlBdpSLQEU98gJpaEfNQWBTT/Unz6j/vmKS/eMGZheUzprM8MuAlInPJzqObwxS
viJ5D7pC8rXhGyiu/1N2wGEzTCdDM7kjlBOlF3kS9MEtEXDqnL2iUTFfnopkXnSMgJSRpZPziIBc
nSX9ix5nisEuk6xZo9r3ueHPZC36EGmQ+97BfN4sTvWOdWZEsn2nCHPzFXXRxJ2npyA0BybtMgzJ
gt+ofYwe8lLQZIbyVvtfEXne42nRCXWmWgDt3LhpwjKc1oI/ni4rbq6fZmwPyn1jZ/mzdIXwR3Ud
f3JRT9L0FmY8KQeY7TD7WjUgNQuO9OyaZMq9xqsaj8gkFbxs0Db02ucSUfd4EhY6LUoMOLIeXVRW
u8MmKSLu1SXWs8UhNSJ//VSQd/BW6QR+HLCltEoBsfWy+tIHLhV2P6J9eJjzKsEOV+/5jcjrAKzz
ecHl0x7H7uB3jbCASlDamNM/NWUqlpTeryC3XDPzsh8COCfqwJ3WdOUftbk8Ou0Ro6jZ7GlY4m+B
TJ3fCU8Zj+mzPKBrehR5fLK7Q2RGHWewY5/+81xFJr45aZEKbjOJz30DPysjYXB3gVaJjNIB9C1U
AnDLew1ZhOGlfaTr3QJN6scDLbcf7ZDySm+pfvgkC+HTxfvQtHehG5sDNatGuEHRXV3huE50b83I
qzCGOZamry6eOU61snPFCyA697/W264qTuQWfZlSEf+CuQA8Z6WmVeToQTjwpzopELxK4FQAWtzN
Gn77plaDu4ZRdwPXO0GPR4aGrykQCx5qs6xhOTA30idCfKKpNN9YKAjOnd6VKlZUf1uqEKDaqu/y
mDPtkDr80AB4X/f+MUPecxkfoDAb+7YOlJ7iESOTCiuzvw/MmrcUXCkf/ebLAzt630ZmSfB0cGqL
iMtnkqbgn9Vj9o8jMOkTw2oAH3wUhBSMXhquk1g8HNHN34tvliyVEhe+yogYGhEuntRclOF0DMhr
PPH+xQJsRmJTS8UAS3X6Z3A8oQqblfTQwzhC/JBFk68DZmGvpr0gYCiaZNt2fheMZmAHGK4swLZk
PL9mgTvNh1iGddNJkFs7Y1ZrO/fx4sAJaWBDB24Dy5GCeo2gkAJ0wwGJ6omvqePbNZH4GwP3K4yf
ns9++8XaQfw88zZDp/q76vj2HRQOgLd8VnNiZ+26zEVEFWi8Ik9I/hmsJY0HvyctV2qATVn+0k6O
mY2C6+RRKKfCyNep7rtOuzPh28rsg6EkfiHIfuLnw3CPEDUxFS10aIIF3Me+JjD2Losh5oOEjfO6
U07Oq2ZerwCG1r6h2fAyHgUZ0IOaIk0uw0hV6iAdEBgwhhRM02Okl7pFFtGSLxxooLGlzKf0O20J
VC4tzYujIoRsILOnFkLjBkooDoOEaaZLGU2VLJ3FaH82C2cenbeTjV/qYNfa+5xnVW97fOLKGvIt
vLQZE0h1ir+9cb/1DaBOpZcqLt3KAuCKxcjGaHalKMRSLnJlvgY0WbngeG9p/FhdrqcYZpXZAIwj
mTSlAkLvh1PXbgmeVj+UchCCaZ90O/vvR6IhpbbkIbBoSrbz0rhRxAZq+vnWnP0dXesu6UUqWKnd
uxbOeDZ8AJA9cGd6ghlKvouYPSzUjNrXzhhtc6m+MmqhIy0if9URHd1hROM2A1GhJg4dfmpCMfrt
86E/tDMQU++7lA7+oycJiLH1cyIBIMMAOMRXlVO7Zy3dzErQseKunyPrgUK62c1+zKr1/527Ak5L
3rn45YwIokrMMVIgoNN4NXkxxh8Egm56VpofailZEhibAanDKBHMAGQI6dp19kxpKN9UKyaviSqU
jIzQcXQpNRq3pyWgKbsP63nt6kiLwmbUxXEpTYRJstMEpXVQVwGYwD/e8trKLpxSg+1UZNpdJIVU
RM9UcZDaV+/A0q3qZThYhQapqC5+JJsUuHNdbcjoL9+ROR0h3k5DAcPG2z4+Bvekqreqlydx7vv7
98/jVvdSZAhM9/SwXYzh02JQrd0ejNMLlxGyqIJB/lrtSfaopTWGYVTPcDtnR/tyCDGizx7fu7xj
SASPKsfyQCoxgIIizdd4smhoPh4dW9Lg/9sCkpB5C/BDwAlz3vOZoga836PFkwQaGg3LUkZAByDU
9scJJ9LQLfVj47jFgKgkfqi+9rHw6voqnvNSKfU1IKudMzY3xyHTiEzMai1y32DfrGupmCFzjqVz
3co60eCrk8LCt4NZHiiws3cvgy4VqMSFJCongugonyZuEpx2TdRdleykFcveThdRfHE7CLTTD2wR
n63HfQ1eRV+2PH+88j1ldd+dyQYkROHTRsKuoO1QV6iM8piSzxZFo/P2tQjS9c5W9fT5JlPMOvk/
vkwhVRu6Di3BUtkyMGw2oOq0fViwuTxoMSy6MJdKCo6HOk9hqERDkWpRC03tV0Y3GtlGoYT2Miy2
p9DyJxf9ZboWO+rqO/6Nk0k60r1bfe7FTGauIiL/cy5YNX68u238LSgC0JxaWhNd/FhNivtSO/+6
1jrdz9AF7ACgATGYObWipX/U48udpPxIuodl7loGJMBKdNGApt28odEjP+/Wd9ZuNRJPy5GSPz+Z
/JD/lH4cM8zNjePxibMjomTsHt4QEnOv6NpXDYsuQXtYXEWtyyTdzIBPIXtM9wP+3RV3HwuAGfre
BZuA4BL+iP0ZbqFanO0XcKD3wIJr59grDMmghkcP7b//6cm3PL7NFeajHUXIL129d/WIp20yqVj5
aifXXxIz9yQqeS+Lg7/3E6fzD+sy0BBQcmncnkjKsCzlgNN0ljqClNgsHncjAvoqPuJAB+1KlQvS
Ns0X1C+UNN5Ul+rl/qFc42f50H7pqtkeogq0UcqOQBXE3uDDFUCQfpiiUq5u21HfiRNhsswr6qEO
D0ydhfSNWgmbqrrveowivLukITi8VLdl7R6cEcA1/I+5A6Js2dfmW++b/Qd78JM1uWO+nPBw778Q
NPjwIZjEhOaVWbxCWq5fBeEtf3XizsoWjJGncyDdqRnwo1/un3Z/wA6UXsDZnCDIAY0TDoTzgrtN
I0UmysLWSYND2J8aZOZ5nAgHGgNuOgkxNt9W/feWsqZc5OHdqoGK5ag/6lGb6h7gybz2MWZylIJ+
ZYXAAXfH8Jwkwwx+OjivGIzk76RA6neo88W66+PkRnnayleR7Tt5YKg3wT/XiAoNfmEpDGIWHJkb
gs60GGpMg5+1vYpo4SRdCUrX4As7F3BYT0XbVvm1Yd/Dxpng6j/OQE3NMrO/YcdniYhhFuqqwdL/
Mu0ed4LOFU/VtC1Fc4VJxA+t5/qqAY+RxxQ5SAxeKQHBknBwir5MoBz/aW8V+GnYriEyBA2O4UCl
Rt956cvGLUF+JjRU4i9CtdROg3dNp88oEyqJMdYEire38n2xZ+tWEAUnGR+bV4HxJs4dZwcDDqoj
HDaIrpx82sJpYeyCaHxmmLLrq2Lo9E9UHTqDshc1/2Q+YzF9nWsuYScCdAR8Ri8qbV8e9U8DB8id
+rMIh7dd4H/ZW4+CjSwXHqht49Ni6VC+ESP0H1MREwpuOT2godJ8f4P5bgk6paQhiqhqORsTPRCg
KTahtaX8Vauv9nLykFjX+C6de6TE62haKOCOJhaer7eLr9vLlXyAoRi8VmWTmKNkZkj1XmoELytS
4+/oXXsT800xRWvx5whYW4YNFNFRDnzvUtkBZZ/dlK1b1471u9prSCycxCdRdVLv02CWyYe0DRZU
ElkfC6KA24ztMh5BtRAFSIzZCtRgP2C5zlIZP9r0QFzp/bwbzbL/X8GYqw8nSnsRpErVoUvsOG8P
+P9dHuXnvMn7ItwGgfaOfHv6kiFnK08FncDWU2TVhqe/ysPV7NfMtjIQosaTvNIZ3Nx/Qw6uxnfc
BXI6bBWRrW805XWbAI0qcOatl/TvaMeFfJpW0cZTr4afHtGyngYD37CwQ0udfuub5xgcs1iHCc8N
twtEvY+5B80u5FYGkQkDHYMV65lp+Y+foTRU8YikKWfSq1WqSSiEd8OU/Px5UoxEEqXGVAtl0Zk4
64LcEBYEKY6J7ZLpkLP+dCxBxpKtM+wpPV2AbFDJeUuvEOhYQhb/ym5CvuAQ+xkoVq3yaHIT2CUI
mxH9NxMlhad0SgnVCvn17S2teTzjIykpMIDffL3WMstA6cD2jn/RPal3M9AttMwmE6drJ7CZJ5cz
gnGs3xUPDSLSFAovZeQeLaWqgrLd2p9gkONdyuyF/8/3AA7QPePMhdHA0Z9jg+R/Ji/Eig/ybVpA
bs5jqJN/HI5PYnbcRtGXxLq+/Qt4abFcriR3iXGa8YOye6mxJSsLYMNFeierDfYXXn/H1DIPsFtW
mqHFtPD90vAQyI1hjFKsqCz09d7A0fZNa1wOkgdB0ssls7jTtxEdetrlFm4ktduCo5fEnu0fIx7r
8LvpuDyF+5T1mhKK/l6nMzN6akWw2XUxGQzO26h2e68tlPZb/Hwg56tJQPAf/rxzgX3jEDex0S8D
QbxzlFGKJK7Iu1EZ7x7shDMTOM9rUz3iVM/NtOPDqIddi4WuMHMdEYhOeT36C4hPbHRFca1koguX
KaYxP9EI0MNMdYIcVAGZaz3VaN4Wf5MBWIvqOu/pFbZHnt3KTRlwDECc0u7Q8z9zyvUD3nOJh024
aH8sRsCnt53nXhYcxN0mkOc6564CLc6QeyhVI5f9qIV2dRpCtMjkDTLUp/X8qhseP17SnkjqTipj
GHTbgUJ0QNuFuheTaSYpGQAoBms+zVgtUo5+Xd1nQclrv28kB9FjEAvw4Kxbfu5Hrzrz1c3d1gZz
TueE1iHvqkTXIZ5FZ3Phq1h8j1dSNsiNLTix3bobXkeNR20gq8OFcfnrH5yYz8vlDDeTV0iKBhsg
eZp1vEo3JJbGxfJ2hIOghHz+7LAYQYUdZoGUlZ/P0f0jQPkjVB79/2+A8gTHLGk2kC0t0w9hSpCe
66fczu5MESLvZ/km6ADkhBLN8pK/hgz6pX1nZPEClJJsu2Fqb0q9TQoI3dwbYfJuCF0tDiWLnmf7
Ank4TrL9vl8Dyog5ap5QBRaDKpMWaP/PW8O2tDWpADVNCx86yo7f5qkAvuKsjd5EfWUXRsfQ8sOK
BskpKyAHVvVfadR3rFiR8rV0ImExNVPMyUo8RwMElakKl+L4j0RpBOEBJ+BHKCsJXCSY6jgdVBfR
jbLEbN0jQZhSnhQE3enk5PYDzkN3/5DLiFoxIWTzaMwOPVMxdlI2UfTaQ4s60ib/RCyt0Lu2ZtlD
7I2nDUBRnf39ga8eVtpis5XqmqqEQ4sRBsk863Qgodm2gCMXe4zGzH2FlFvW/jxjf3ZbYIr+N9JK
Y12l7f+M33haCX0eF0LZRPsbp8sWhZyM13p1gNZ3HL+5CIp/mB/EQeXqzlEJP0Egt88wVqnJjspC
6xdraaLsS6IubCwlmbcC55xNtS4F8G5yEfLPjHsuM0Wd2cHVxmHb2TJ2zkR1BLJp+W/TsH4ylELH
k1RO8JNGOQlGcdnUblPWmiJbX/TROn9LkxIQlNXX10FngCY2UUM2YviXoWb17nuwbOM6Q2+/Y93I
6Fo7lRVo311hW8Tns2DV1cjKtsz/uV5SK/uUtjkvklKiPmqHfPRulEZY2dtKFFTk1ALQe9L+SGoo
NUGLnLhSXNQX3EV8vl0LomCnyYgK1uSvr93uvg/UCtxYtxSXUe+GL7qdbJSBbgGyRLaPRyKjBMdk
CZ35QONBrcqvF4T7Ntc8Q6O5MXiBKXvq7o289DzLvzhQ9Mrtq+OdxcJSRf6GTn9XCNzHKJngcJqR
Y4qf+NtBJ0Bc+WUV0GGDgrKPICZJUXkkcdAj5W5BWV8q89qtNyNoq27PtKzSNXQrH7vWdsycgUSQ
KoBX3V63uh7FK+3YaWpyMOA5DyQ1i0GwocGk7GYIBtNbPaF6gQXxaX1OhMYcIzLIyUpFzuNm75Su
N7QLIWWjlN6edRVq/EUP08BNRr4s/CPRnTBXElR2SsBZXctBQLZF+GK4V+D5GJQd97Y/nNvPzR1B
l0q/vEAZagPF3eMeJKA0QzSuom3h32k0hfG2RoPf9ZwCg3FCUpQwkRv0W68/8RC2e2ntSKI6aDWw
C5ysM+Gz48fkFuiF8f3zxfM6tgBQDkoEdchpv+LckIOJcys0J5rC3IzQWuGdaBQtrIL40jaqrB1z
Qv563hBscrkI+rqM7MrTrdMAip+6/9uE5/twpoiyyLXiRoYTP4E6yKJNTHAQRjN0P/DAsORMbXrm
erm99LXIZ0lpDuesmXCNXpCrnNg87QNGOPVWjzPTeCcy+2JIX6gz646C6s1u5bNB4y1lc8zjc0wH
cMjop86UlUQJki9bevaFr+OYrM/kAph4WiWrbNcIkN4qOV1Hb1CM1s9YYh+3e2tjMABvWTVHUyMw
cttIYttPY/brHPPQHUrwk8hi5zoF4CXgkWk6b8N7+IPCIzAUeKIOLI+Qut1nPqMCuRooniEScIC6
7AKHi+C7dApjNPm+lXoTufXxj9tAYBySdZk2cMMFbzjdMvd57anF5LlPdFOIvynAkIFXBlnp5hGY
3IcPtolYL0QxpjYf6sp8AWkx7wdfp876pSFysh8/wG/k7FrfOF200u5TznahKcWGFtQXVFYSBCzY
tdtDqM6Yvjh0UPeJUYBo73OqfjbOm9DddUnVDgWM89GMjxyXtI6XzZLotjWzlnaiE4duP4IGGZr/
PkW6KlqIZjlgCQyfZzlYFZc6SHCtjzYKBDDyE/bnY6DbjKA5wcoSDSVenfajh/EkGg7XzeGZSfdg
U4Ly78PeKD5CYiW1e1kgTp/ook4CHAkoLu6ghDuQUern0hubN5ibnIyVr8JiBnYl7F7ydMTvzf8I
dRGXdiqHkHvMqQVwJKFqvpXyQs7sIR1CgutgqfdJm8T3Od6pdRJLDV+dqnW9tjD/euVlnaBHLGQ+
wf4eyJpE6q5mmrbVaR/xZavATvk3Bq++WQUuQ9nsYFyzaHNngljB42I1h1GMuWoDfAq4bI1WOgmd
X3+gS5SLw/lueXrIXi2yDoEjqBGl2AA57QiRV+EPNqLkknzlnktMXZ6cdsM6vgoqi4VgfswMkbgc
D/vVll5uP1IOX/J9ogiYH4w+b+pEjDWEX+hio7fCsnGyPEjAjbicjGznWlSmduTXHivZs6hWWUSo
QSpc5kGkUl/F09U4YaM/HuGCs1AllwfPBI+nnEh+89YNcmhDnEuUj87hyutwy0oXDru76WfX+2z/
rN0860op8/JyMFo8fW74olHAXF7I3vccyiQb3LdJZW5XAmp9aPjpVX7wfMG2fozoo+vwohiWpZEe
gz4pISZ5hG+eVsxxKk1sl21lOIwRKA2bQJ0yrBrkWZjewIyRuMAVYLhIzRIhJDGVjATXPaXz7RSt
QmHJT13+t6ZPSD5Dj3SZN7A1NoZ1ONohw3KyEyHuTyqOjKBEQWZqeH+S06IYJfFsWJopvl8djJga
j1oKJI7o99yEvUz86+34lulHr7wtPxAdVjGlPnJo1rNDcNzOk4VmlT6qj54JKNAdQCTg6vxtG3cZ
f/O/2rGBJjapkEODbfwf5QWgyBBCym8zAAChPA3ds3PVKtn2EZrxtwFVX5d/KwZ+hf3/DnYxzC/j
Q3tIXTuitDABboh2B/meaXUgvYly1zlC0IQzEflhfvyXNNo91qO5o1IrXtTADfzklJI3+o5E/Lvl
uw6y3gem/M+yy+kaweqeQcOv/uYgrId54hi/ggFvMcz63gLZvrIXTzJxu0Qqk8qpxYk5yzdfDQeo
EtQcjU6tyoxDVHyiSWE74988q7W6fDidW7F9yKG/sBCUCyqQHNM0FP0PtNIcO9Jt5P5fRAssJSNX
JWbvrkPFzshMzymHFDCrnYExVEQVwBdaQy9KKmMSdHRH6K7okUmtsxyttSmTfsyWeBrGpRa7jJ+D
xlVwv6hLgVLnoZF30/VwA6vorc5UplyHxh6bhYYOfEXNv/JrgOacJ2vmVb7Z6mQDblhhyk6V+WJF
Y/ZqQuStOfX4BDEpBur6vilWMcRztLFXXr8vvSEWlEVbyQWdhSz11UieFlh4RoW+aT5VbCSg1Y0R
EQPQsb79uSpwJ6UABWEBgrkGFnXX5QoHFarOAp0SIoVQJnuCAfnpRitgWeYcHfEvCF2YGeq1Mb2X
0qnyyZGUo1I58KgTLIAPTqpNdGiRpvnADvphn9lMvglw50+FhlmXflYFexm+JMcwlZOq6Y2QpRXg
2sId8JfmauXznU0l5KNq4HNVIBmzsKPw0Ww0oE1Gb4vdpk8NVmZ4qDUFXAm42cblaardwL0iklK5
VL2v1JHohkfQADOvQnM627ALY/XaG64uaSZ/Z7gllN/GTx2e1s47lXCTHrrUAD5/sJCJvNLsauqn
jBMXgGxJpWAsHzL14pth1vQ0DtkwMgmHlFm1XOl2zb5NFpmQilQmyXJOdqDNncdhSxIhwfDF89H4
MrK1PIPXfckjHOz5p61Ru32KblWaGfxc/FFeQmyXQszLMlkjbS+12l8wms4Z7AD3xA4ln4Rfvhe3
WReavYZsSAaNejd2FMTydE/x/Ev0ehL5YDUNlM6UxnOwqvmzLowqf30L01QyrLuwy2BTl8YqhHAt
6vr/bXP0Kii3Qx/cxuzFjYY2MbjQi30DlQJJhI3yVQwxVr8rtlZydSsQCa0N12Dd4GqxZJ0Jmuo8
t+1ODAnmKlH1YOGHgoxhdH1D1ttBWmP3BL+BYXCTEa1x20cZ+AcaByQYyr2L0VMzcgSv5FYwbHGQ
LClf7nK9/G2lQtAJN7UYOYxlOlvHlRwiVCiqWPVh8k/grfk9ELVr0/YnvrI2mbPD1bqdENzIuxtP
Q42vCcJXlmXUKG1qjokcJ6faH5hdflsldWfjpZs4t8qDbM6ULKzgq+X2PetNEcx3Zq4IXBrQq3lh
xNURS7WGxx/LFns6N5z6CLl9dRDyFpdfqJPYa5O6YcnLqHhUNnVApQBESy3VF0m6OT7ktYI/zJOo
6OrPyq5mdRUseC3NupQ2RGylbn5TOWQkx/9fle0Yd9oITY4MoRZVCGiMJJCAyOjc7d8BuDypImXr
3B+OfAo3xQvZFkuy3pS38My839ADwXVW+MDob3redeJQ/3vn4rdpyXaZndD66d3VMZ5yDZRLi8ws
XRZ0OvKji5tQGAi+boqK4fRnM/kx2xKWNYM6LDyKrw+dic80zqSFJ7xuyNw9F+BGzDYdeKycFLu7
04cSOA9dW7IeKNGyPYQJ55ktYzjisK76YdR3YA5o4g6rHqJJZFWCzRkjs8nvVad+BnRCBITHwosp
O0TyGIHPjRl7hXSqVC//yLhFHNnYBCuzmxE8pNWPKH2hL1gEq3c7DmqPFze2B8hv4qpqZxjSv7rJ
Avuq3/XcLiV7g7LMM56Hi7M18SvjyiPT9VUS+yxavSQCdXtrQcA0Sp8H92ovSNkFZVBV+GX4cvoG
7KYNv3uvcqfWCxP1JaVZw6W3ujqBsyilPn52zdL+OvLeQQ2siPNHaBubUO1OVxAE/KGpWoBocQG6
cx70qpS/wVV5A6/O
`protect end_protected
