`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Zx4YoEI91Rsc732oUi+/7sLzZeT7E+ZnTmkBNE6wo9/46f3/i15d6xUcRzCLCfN2PHS9J4hIBeKQ
14adx4ypJlNllz+H8AOhfQkNsOQPxqNcOBlGZHGhXfY33fl4GWM1MqAmYpHG1AxhQq7/5taDPtNx
JGM7/Vya0F6NWhLemayhGN63mVe2qYGKPXM9oWnfXK9v84R1UwqDASLVrTS66nhaPfcyR61+zYPj
rGL/nPhfnkusJUxci43YKkmGkR/dv9HksuYO7A2AI4d0HQFIqOHM6r0NzX9vERgWSYtcARbGY2CW
yVyBR/uXrWQdjKd+9LVPYrRWPmDCqVlPugwHeg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="V9pVIaJGWvK+m5ZPFuaBaDh4nCBVQVotH7IxGve/01A="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2960)
`protect data_block
u8Zv4tGxkY7dib6hh7AAeQza5Eu+4wahm+NYXwUzhrm9rUZIbnaUO64Iv6UHmUpG6O/i19scPznR
H9jN3gzj6JT5loeD3hbAvX58yjwsBpCJQevlKzsgYNu38BswzUCWjdFWpD8S/JArQtyqzsrFnZEE
pOTQgdDzLQBlUHRr3QFTzBHsmCP/Lciutud9sMswHeKCD4QmiPBCgY5OH9Jcn9ZfpOJrDS8JyRPx
A8wgv9PY2En87fmhd1RwLaCW7xfNLlj1eSwv9D3rro65HAR02PwMxz4Rf0FePzuz1FCV4R2tb2zm
uec61bvj/MCinUnB9T65leT/4OmSPQ9d4LtPRbo/ziOMOYdhR8QlC5G2x2h/5qkaw4QHTyHnYN2E
BjlKwgq9FpeiHvG9gx4udFbeTEm+w4qJJW7EOrs37TEdIQa+BCH7RLBvHYNxpGECmn4gVHzL5LWW
MORtg0u1rmAoIw34e69eJDV/NWrmRbjk86QdJQJe+TXZyUFbmQtmq3xrXNDtfX1ck5u2r0A5Lpay
rkVJW+NkWyJuSGO73lerkVx/z28Kz9A0lmC08psDeED5FA3eDalDAHwwzp9Rw54RYs+mphJP94Ix
ftzJ8YBh8/yoiDUDKbTo5RXRbFagWdsz5OWCJLeevQLLeQ/Hj8M0A6rY/Tbd6AD9n5z1/zZ6Ymlw
l0oL4R8KrqfFv91lGLDunL4a3XGva+se5DxWh6AfkgXFwXpsCjZqxUHI1vc5F3EEY/QWQKkutT06
3GrYWKnDrUK1F31EKWzo27cImKnfSAvwyAs0q8OL5GQ3NZMxUGh+hWRDSHD2OFkaAejuGIhdFgsH
sqOegZGQoNcggKmT1utb+cvsU/cGGInovq3IBlPnpUNLsrWv0GMtpn1o9EWwHE10pVtAlXCjPM1A
8SokorJ1CUgl/jLPKcs5B7snt9fFBMINVHzNWBLBrzrnIioS8HTE4UE8sgyArL6qzpgdVV2apa4t
2hUQB5rFnhVBKLSCEeEcC9wD5Vck3VQaq4jH+NI6mrZBsahMpWX9RtrL6IE/8Rz+VoMcF8vZhux/
PiKX2H5xspGhEQAF4zyPChLUFje06iRC1gecLC1cIVXcuKZmr5r8e6/oM19LwjDoOmTgUeSFlcgZ
dfEQjmZdXr1Al+7T3V/ON9aMW3kV/MapI72SjdFcGdVJ1Vbg3flxejVilZX1E5ZYl97wPFm/rwT7
zvcMyykeWtSnQGsmOc9da4DpTosM54Qe7jM8BD+U4rUnzgCRWUG4OEu9zUvMG+2utLMs3cpKiHVL
GmjMQH3Eic8nOLmto1svYGuRbgBhCHT+lHCE5+c0Rf5di3dVsuZATZZ2wpClZElFmICiScMmfUW1
EC+NzZ+Ort94ncXlaDu4WqYr6A3C9uuoj5AkhYmHYqJTWAuI+Vh2JmqDkv0tW3VAc2ZosNQU44Mj
ozzHKLzLnOwL5WRw+cVwRSO3bjo8SrXSDNF2vduND774bPaaAn3gLXJCbEUDWPp+f5jbsivdJaYR
mEvwZxAAzlFIaECyMdRA2X0LPtDCP25CrltUW4dcK5iR+c1/aCCUGDzQwj4AUPHxIX96ZI4/1Mww
Jsxmm8OGy34rltNHt9gB39hCb9HMXA+baAAe0rNK8HksQdJ7kaxedeHmTUlkEWj4mnDQPL69DrX4
o5NqZW7dBFXs6c3cAF2W+AcvTzy9cR1+0mW/48ozKGrYlsHwNXIY1lFUB6iklYpCegAlkEZ8FTLX
Y0VFJLkaL8SVcSrokpA+R2QBIvnW1opxi74AU6SzYPQQ9Qd+BqB9tDdXZ7ZNljR3/hGhRNN1GdwX
ZUxcF2cakdUHW5prdN5YuvpyU7VtH6CH36pnxxez3/2pklTAMTcwG5Aku3Fgw2fHIKbk6wXEqk/X
L3rZ4OLHFR8EEjDYYLp2D01YKuSwZaCQ2kqdY5lskYX1kD9RoY1DZPLW/78BqwV4M3z2NVNcluga
El63JvlSq6oZ+0Qq2rY8esOINGYAumsavyNaE8OKAhzekO3MRO6d+/ksTkNBr8qCb243jYAKuvQV
UusB3PTpAvAbj9Wx73wZAk6Z28VSmW1Qo9JBwdJ/73XT9SIh5p4YpoAWnQypCjwXDvoN9UNRZTZ0
aC/PS1vAvyOaZzJjO2xuzL8E5RyvSLbcEigGRasKo50C7PGFSoisei5ULYJf4+bi8w2hS0eGb+XZ
VBio0LpQrG/sF//ZeyQLBKpV9GuYTF7dYYKv4oOQIhLtrKyJFHnDrUa4R7YqTXoIpHL9up9kPnrL
b6ygcCudGXI2zuviCScoywNceKIRove0YLprJ01XXagC9hDOoo55waMtcP4PqL2yPnU7B6ZSW3XW
gUehm2Ww8zCC5e9o5v/zTvxqcNWn9eGuNpWdT0ZEUjLV9kcA6o+z/2tigrmonM0bVDAcUqPLEf3L
mjic1t0k9T4sAQTILji5XKMhmLcweZhcrYNrBkNuMVNlxV4bphYYENuVI8yToeyPyE5IJ71xFSRa
jhvhxDX5DMKYtDqsWSucM47nXhMBCuQ9JZyxzaANtoPofOhR49Jr3LCIhK4NGZhnd7ttG6xtsw2W
4NGEQHLHTt9w0NZ0IA9r81HbnNN8GNsuuy5s3/txKA+/R0O570lPwuIsF6z4awJKzCdtS0m6i5iS
X0PeDssXEX4jZ14zMAclnUqY7rKLeUi2JT1xEc6e4AQIbjBIFA4RYkI3YsiU7w1IRLW8fhDBV/v/
yeM2v4RCJtm13QRH8LwBaPmI25VX4Gf3Tod4TwDUFoOrBFbLrFmIYG1JUhJPnlzc49L2CR+1D2K6
9F/6ya7J1OwszexKm+NjF+/lgdmkOL/fWKQ16yx7rYkw/tLbN0rh+qL19tzeQfjPMPL+8RxonG6c
Bb5z7m7WCCbMloPV+6QtYcfr7jl4mbGT0g3xbjC2gAfTVuG3840mdlI1hI+dyZGBfVJ+GFNXEeRE
BUx64BSDv5WMQGiBzqc0AzmdetuDUj799r0YQdufIrQMC8xBML1BAnvfHIS8uQYc9FwMwEVTXoJr
/jUeluieqZhNQiGPN3I429G/SfkuksUwhcuKLihbk3xoK7uxvBobPoOBQqBO6La6LlJYmkUuH3u8
1eOfFT5RvVRN0CAaiRRDwGdwbNA2k5I7/zvlZK2j4NthI1N67qdsnAHMIjWNr1M7jXgCdwutulE/
fXDd20TpZeIJ9chSiocCSqRus982zh+zh/al3DIPdXitqzLzcnMFfuwRl1tXma7L+4Snt2/8ClFn
OC2BW2UnVMrugSuc+C2KtBT2gpt70p7Xgq1HLQZsnClpl/4hJTyMhDNTxjgt0UAvMvZAGmuwtHcj
Pewn0/0tlMKMrZv5tC5bF0T249cG8I4wE0gGoou4aIeLHb8wuJUpBU4d/pddsTsBl2yu7yLVL56e
7zXRAdKxtQAaFswEpuy//eJTfmiy5a7Q+dCIPj0Qb25TIUM+Ixp6v/NIusg8e6pNAMbJHctp1PNK
4CzgQCdgKwM2Lv1HgZ80CeFppfo16v7jzJfPuun4CQuVmQRYslnz4NASKH5+IQdtDnc5d4SFvZY3
kACm0sA0coFVncKQsBofO5txT6rDj+yN+xmw95Pif2OFnwpTjfm61B5ammPe0z0xwZem7Zqb6S10
nfRJ4fdsQHYsqI5LChBkBL15Vp5tJEMTbe2U0Sd8Ou1iRQZZWhKo1l0a4sfRehDZEgZaoHg1j9vL
DFFaEsvKslyJMVl5YxDk+K9uZsC9X7v5b3XvC5YE+S7+G8+w6C93GOnD6sGD1ArQyrBAtiPo9QQ7
Y2+BSwZwbQsIfGfH+OjV6NnNivL9P2lrQOGCXvudUDtBOT6mYZZ90ZjDbFgtaFIByqXWykZaErCU
kBmMKzLR2/sMD/c9TRAvuafkT90or5tG1IodxS0kqN29Ac529BWH2zRxlZff1CLvfT1eHZI=
`protect end_protected
