`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Dc3GAZr3HtYvcB13eC+r/3Ka/E0FcFB6AhGurVwCS9lEmiFUrokVGYg1j086lMIEsj3Ij6z4HgBa
NLZ6aBBL8sNzTAaGqmHte3xRP938PlMwmhaDKu8/4mmJn9LW8FfbVAiUb+Nd0vTKkfxLvRJzq4aW
1Raj2/u6ptZCvILCxaiQcMkDX9cMxGsSDjHF3mXrRHQDo0OO8Zcl2fYFoWtG0OD2MarSnbXda/ia
4K0btq0GltOPyWOmup7tiKm8TL8Hj9pqf+j0z0J00mv8EWlwLR1mDdY1nNNbz9yRjgTnT3w975UP
SVGw1Y1zXnXTdClOA51rYxLqr4jujJmOahOjpw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="S+oGzY3evpv1eW17usMc5vqhk/Xv7dRaSuLZKRRl28w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
5RPHUqTVnAJIYahZHzzWWmh5rmBL31guI2KoyZqUBat/tGrqFdnsIc+6boJZO8xzoeBoqPaiw/YR
RUASz5C7NOdns3NeNcT5zEb6ydnNFiyS7bQ8b5KQ+fGcQq/qvxCorXYvfuRnh8eVELk40bKK5iOP
o//CeRc0dpx9dsyikLNDRmobv45TNi8YiOQ8WZdzaNhow3QiPtZUPmCWXq6+ME9j+NN4SJgjorVa
Q56myoXoG/7MPZOHhEeZRrq6DFbQjW4+M0UhVEFtsjAgtiRsSZUDlhmOzxDazOVcl9RmorehOJao
h999qLrtXVLOoh/6YiWQ0nRAIdwSI71FjTtmyKtENe8S5qn3h2Jea7BYZ/Pzwzb3Piab4jxqaTD8
MP7jr+cY/UTsA2LooMQmDPPEXcIyAryD9cWC7MV4RKuFLd9Ej1JJagIWQVMbWO+Swt5bw6IF/1qB
G4fzo/hEbbAIppS6sg3wqcLYZNj8DVJFuko5HydYuMFXaKUWsIR6sWDHSdLFjxDLdST5Oo99TYSG
AXD5uN4VYYg7FlXOeKyMNJYe31EZx+nZJ9uUhhJ2yrub6YhDmhRwDFdUoVfmgLtNFoppQjVItbM3
QbvWC2vyVGdIDzdoY1ROEpJG5yyEP8F2GsXtD9dlCZKnRzEVMZHQNjZ++2eckngUtBrsDMguGczW
rw277kd8fvQEaUTBSInt2OIsHFM0f1HKMHw19KiE8JuBaBYujB/3w2vvE+uhNO8FBNI9Z7tkYQfv
Nhl5tAPFWEBM/XNlfXjDH6mh7FknG8Pe3vN4YAV/ktl9w6korsXAxRwMiVURNy4EDr6YI6TvtgJF
/R7IczFEgaHdnABd5ExCIdMZsiFBF5UIW40vCU16CAYbe1nmprxY6U/fE0HKOTX4eGXvAaqZJmsQ
gO+BfmZuNc5LQz5CJw/6q1C658j4WrSXQ+2prGHk0Xb3b+OJk29vo24aQzkMeRSCCqqzF5Xhkj/v
2JgG/XHTZesuEe1K6wTSWw7VgOVyZ1l3H3Cu1UrKLRX7RIWh6VSernOFW2ORd+VEfdBGT8UpPdTr
gKxaxujToZUq7aBWkNwDfLXMTkw7fE1ZG8JJszOTnASN6JQ52X+1fLg6drgoIv/bD/M9+0/qEQ+r
nzMtaqnezEusllYrp2zH9nnxBsHnqTulv6kDoo8ja9xoh8j35DmvOUKNumQO3X5jeQ3tzhKSggP9
xESKhVmW/HlxHz1GJwOG2WbnGubmHoF+Oo+GWuG4UKO5uylvjB5jpArbVVc5duR2ItnVqfBA6lxQ
udZSrQJn76e2yeo6A01wocuqhFJNa51RG5J7SE8qmsMOeOaLB6+eoCE8NlTiYoqy739DMufh9cwd
2khgK+KgA0R1252h7ZZQ2UfIErqd2kcs6Fm3FKpTmlOmbwrxQ/sironU+YSUqe7W0snQYvGKJcg/
zc6jDUeOA7Clei09c4doi5oo7IddMRH0TUHzRdD+3BIYo4LVYKf+L3o1qFrwBAs+CG8AI9PxrD3l
6CrJGeX8dkfXSZAAonZp1NL5UkWLq0qiuMJVFZiRTJIjTamznDlIg0wDMxWYt93K1Ckzmt9epaXc
XCG971WsCVB1vkmdhkHqq7BPDtfK8dWSI50wO7vOEl6wuT8Eii1JMPCjcJ0NgocFPq6OzxyZDfl/
IFNXjOm25uUMSTd6xBjgE6ESlc0jVbRyFliCVw9IWZpK57SVfwupHDD1hDg5l95YkxPpxvJbGV3a
6TxdqBLgWSG8o169JjdE+WjR0wMn7JgTKGSMifklX+Mix8YbzchzHFNol1KVu17XVHflJosPsX/K
GNGOMzyYeS4yLx2gpi0LL+gh22KtkHnRbkZTQk35vW0/705Gvzozq4HwzF/yg60MZd+v8tHxuHyL
Gd2znB955t6+qgrffJW3nZ+0meDy5ZkWHGCvzAufrPYVSAwwe4FnXbmZBPIjRNY2oeAEmtgO9C0+
TOISpsA4JYcvML9Zq9KusaPusfg+8e81Hh9Ovc/GUulfZK4F+FhDgz+DeJJIftKWtvHbSMIlYJ/z
SEU0CLBMTR3muqGiG1PjpJNxfJCdLMtYeN28P4R+ODeaMPxWWUUFEeSDRBzxY+LRzZOXbhlt4lh9
fXnwxgygrclvuEHExGo8hOogl395mEx58n5Z3738Fr1hDftENnPtJPmrAwgA+8CbLpBPa3v9VZIy
1BZbuJ7r943lFhYBiNVy4LrA/3sE6KLfosUWCse50EtiRf0blJOpEQMu4nlj1CiO7TLzhl9h1pgb
hGW3pOmT/VWJ/fnnIAPMSmM+wORBoM8d4ZwX1HceAYL51HzB0Cgb/buZR5YBioky3m5rk7SuGyiQ
FrAvAwX1/VKGz+wC1eslahlnv6De2cDNSiBWBnX+S0FXtdwH+Y0+yVcIMIaimNHveBXeMyCJyclQ
eRPOS4wIbrHcLJ3AyvWGDsyJYfOp9y0bGES/Zq28yUH/7DojzCi4P7tiT9M0n4E0X9SEZ3kEnmAO
kJReRsfwny4MyCobrlzIwklqPDyASe/Upd8J/n/n8P9W45TmEbYN418UI8OOk8ZsmkW2J1C+4d3L
UDsZDXm7LSU4/UqQcRqSdXFDPxZAc3ALmSBP28BRzwjhviKwstHKAVmo4Kadt6eIAa3d1uTC4zqH
mxdMpjkWeEQkrrb8O9zbN5/wzmkO98scR6olw7gTwQNJi0sY1VxZU7PBHKzdPNfgyRrgBnCUoyiz
aPGWnaXqdhDmZQ3lWDWAqjYMu4WNsaRtZEy87yQSvG4fRm6OE7KUP4JnaFlieEx9EGwm3NA2gVdc
ail6ACzgMTmfymOT+qxk3exm2FhV5r6wIU/g5oG6XvG7BtToigNVggByh/v1K0DclMacuKG7u0Kt
VFKEAaeE3UeY1JkGLdR7ECz5BKSg06Kk7KEXsf5QLbm4QyEu+K0JhtROdNar7qMOpb4iIQMAtRbC
OhPRTjnYhG3ktZXGhuRWIhFyrgTv5l+UnS0gOY/k74zsoCAKe3bPSztltmco2n01fe5v2YA6jZGN
QDpz/RRtupI1mel9rrQdy7VODCHNEvAQonLSvKuauSIQtCWkR8fxbS5hQ77zzd7J0cLJbc2FL16s
9kdWceWzp7iJxbXpy5UYYzqU4XyooD399JoK7fmF97ub4p8G7aOYjgNbLe/nGt2nf2leBoFyWHMq
tWks2vc1cmu2rmK+0txicmDEOcD6RhxNq7tNfZ2PcfK1wyw2cMPkScOKG5zo30wg3N7njuTkzcjr
AhwfE9KyLJuensU0gZV5GWr55eSdTcn9ajFV5jHj9rC7YPyJgLtUAOpYGNtbfdjKURAq0VDIvCL0
JExE5e8N8Tmsz7rRJTEi5KEJCvMiaJP001jU02/4YbIa9qDkhVEQka5V25/pJm86ZmSplDGuvoAX
Gx6HQLZOD5U9h89EtPoTmhVsQyVp06McboLFgRL7FMQZx3G9olXA4iegx85QJmEtzd1uS0xXA8vx
4alXn5pC/YP6l4i8U122WsfmiRfXP9+dWMjpx/PptdXJuwDi2ileeo0tMWioIucF6s78gH2uAeMR
DUZ9i8CRdzeDWjLOliSTXi4dBefLkkIZyqg3aYli0jNi8wsyxlJCKB34dXH9virxrcEXBxl4xMBu
RPB/43liGjKL5g+MsEKsSSRoBnVT77PUF2K7cjzyKLc1zxCeY/kXcW5XEqAcT3/w1mcssSLwSKCq
PRJhGzQ2YgJuhPa3h0KjdiO6xRUCbF6sJ7G5o3Z9O1PmJWZMvyfuT3rOIaybWtkc+fgoD4BRTHWl
A391/0KJQLcAJn/REIc1Gmnnwyy0CtnrFdzgo6nb0LV9Ol3pwihFJ9ehjwSw1J7aZpQRNVhGO34h
0NEk/JN8kAVGZFRFTcCGVNcLbfe9EtMQxP2wckFmBg1RFn1ZYxoXXJtXtOfTu1/RAGCQZbNzkeTt
m6DQ9aNIZzRmOwuo+H1t0iWBTZKQ0LLV9ySfbd0SNYvB2HarF/dKwECF/SpGaDkuVjCA/0mAk3YX
irU7HAvm6mVvCUor4tDd0Bk0CjXtA3PsgkoSOr9M81OPtpgBEkUnXWsEDAUZ6wGjtOArwMNBbI/7
oy/3WOiEwFGwkgrbTi2irP0849B2ndEMsEdJOAt4b4R4ehnoNZHxIp0/8FMk0fAGlaY1rXH7gOSN
iEPs0kCNeZGqt9qL3wJWpp5roMPh7zupugeAcS/SF0YThQDasJivASHCjuHYLNnZAuJJSDwTa81T
tx9AWVi57glqdBurJ3ChgRNbBsnE+J54xKCFFnbT+/HIwWN4FSiY8MENo7XHdMTFhUdTyu0GGAtw
wCKcQVyJpMFQEtBZ/6aSyzc9+C68OlgAH+NKYbV5yTf4yowL0X9101eTZex6S1RdGbNIxiQrJHb4
D2a5ZpbEPWbRVBZXWC+csMBozB/MOiaslVO/MyKZzTQ+B9bXdBU26sqJTY6n2EcR2jP0xzwi5An0
/WaEAzjG+vGeRpBJwN9eWsk0O77gc4/+CL0vm8xat4ssy/YotuRnS2Q0V/EedeObZcKU1er/Sf0I
DCtM8dcYndi7BcUxaEzFOjA6/mLiwL2tC3j+9kV2AoM1rWo9Y4YliKVyktL2ZbPafkhr6J39neZc
pB2kSUQ+YWF0TYK3FbiGDZ2T0oavYcS38JEI/3d2qXEFjfA21ICsv4MrcnE4g4/bkFPKfRKFV1qT
LxGVAfuxH9MBu2VVlP1Gih3vTj83BiXnQNSkyHqtQGRCriDBxEqpEcupk1PkqmBuKmX6fxU87Zv8
ulj0DgC+CXSSwOAO4cTkFjNFicv/kGDMqe3r0B7V70Ada9pXDbIrOp8Fs1cyZNGkcDU17U3s3KOn
Xw0OD1pFWWNQZoshIC408dR+WmIe6zGKHlbX+s63aedzaFUEXX2ieciclCIj474Mq0L29liLoOjS
bajG2DRavzsUiGQ2CE4uXJ0T5MFBwsQgvFvepmmPxHfJ4JVxgYMoeMQIO4M7OmHzxHB4MB3uZwnI
l8M/sm7WvRHeVzn5bWA0fgcg4duyIop8hN+oantXinUyQfzVS7q0Mv/ztQQXe6qTXi5RLbmG9beR
qE6jmBWFU6EneKmxvg/2fZGhHvML2ZGHOCx0ewIIC59AbCzaPnta/jlY42E22+MsFAs1Z7xarDWh
/8VRM9CqyRBf8gaozzwS+aMKwYjCiMtvRAxL7ixRmLLTrnsszUHCGHn6u6Wdo45Ry0Y4sVYYuH32
ZzlONWM7BybtTaBHHDQ3vJbuRTdMRoPkmWWSMlaAYsOiPQxzdcsn2l7M8p26scZBsd4RgBdkJKzC
XqMGhmdNt4sEsNfybkSHsUl+XKdTWcCQx7GdqbUklbXNhW6/cHa3DNVJuIQL8ig07BsYKjWdYZ8f
g2W8miu/0n2wa2QfeFnIiD9kx8B03ndrT4l6XaBTZ/GEsceARSW+fnv5sHWEP1QloBFnA4xbuYD+
13o6zPsjIWHxN4BC+zwK0iYxrUb2FUTkV47HWNn8y7aeyng28YF5W4aDHOHkgm4ygZZAaNryEWD0
von1fJ2taO/OXA4laGA7fhWdglRAkK7aszKO61JDCsqWG+m8wUTx8FBKZdUY3GKrZqEMKjgM7O8Y
F65snC1qanOAlnkfBpvMN7QdwLCWDEvz9iC2nIEGB46iTFTVcYJNrc8/lSxJrLhkQ+0fY9rUExqc
pWuvbHYEEgLhEYQuUQUQXEnqMzcb9wexe28E7AfjxmXkc8LbSWkUvye/32vxpbeiDx6FVM0UjPi1
3ZgCTPceT7E54M3TFfP8Kbp7uBL0bFG1bLB54fwMk54YvkSYwlE6ef4O/MpMlxsHjubtvKnwRtTW
/ld6q1xYrbBeN3G312vkEN/fpyKM5/0BprOndGoTV7pR+7oCJXhYOvcJ2zHBSs9XfQamHawvE+6a
ZasxazIDLez6uqkXEDRq/5pv99nP9UFY8EiFIvn0NsEBLLfN2hOHmpeGwcjdQ/wqXV/++AsejUj7
jN0sLNRwwXibvXiNljHhXcxk1TVs3s3x9y16bx2Gdp+kA7lHlvPFdZI+FTc+EKOSMrAY5X1dFH75
UyzpAENmUUd/Zih01uv1nLvZ2IPHNUyC7e/XeuArRwIT9PDqN6TYTR+AcKtCoVHEQQz0QNFHTsWN
Fa47V96iENl2vKvyLY07tMMZ6Dq62v1OOThR68Nr2gVX7Byti+r0qbY7gaWZcuklYN01E51UezpF
Z8xA7XXFaphWckBY1ECp6A+8Y1UeeuOydc052JEoRBcGew7u6RiPIBiyYy1wCH6mTTMHdPF8ZQ6m
BIUlzR1zPC53lR9xZvQjLEZiyOcWCm/H+WvBsGVUWYbBMuNvbs3e8xvwWeDdlppZSVe6mPdhxbRQ
p5clFkxdEGbNJPrxE8qdf42p7HSF/csbSrrnQ55MEiSkl+uPXum2FCRjrI8zRCFNEW8xBln2s8L4
RP+X0BJ8ANtkpjt0F/Hd+4DKNPVgAgreFP34VX0emK6qYBYHc5rHsUpzmWmldt75DZiXjZl83PKw
4KYZlEDC+oq672yGKXl+0h8pbfRYvhsTjkG9mTiUKQezv6FyGKJ2MwKHdU/Cg1CM1t0xPhcklCLc
XpAXkJgZpyjmpefh6OH8J3BBUhVwUhIRf5DJIFKTgPvKhipymTMkawNlqR+qrltJfz1y3Rvz11TH
y+0xVH41tl4sE5Nkm7SXJQA7NLd6rklufkD3Yrx0eAuScbZfZX+VHt/70tP0LteUWSI8ci5UnUo8
3iKENDrLgAoNPisfSxRypuxYq1GHkuYyAzOpdu1KCdRMAalzaHj45r7Z6t3ljwG3P4i18v/o1BGR
2GXXiYN1538kcPxJJRNf0sm0G4whqNNo56+VxQ94Sf2NrnsN52EuoT/sYzKSF0pdh+n+CzFfS2Sy
fmFLQ/cNFboiKd5c0pCRZ6yM0Rn5YbFybICwIa3zl2El4wqO9WQSe0MkgQndZWC1ia46pQZ1tE0m
BChyp+Etq9ZsZMiKhbrqrmtqiFTx2ljgGzm2gli9HDMGLnrQxT4pUK59PY9cRJ+IhLLuQwUSO/7G
MvRxZ+DrMglYLO7TxJR8AjaYTEUDBAPYuYmLbLzCrhVDb/zbijTSoJbI2QFCJV8+PGX0VhtYSii8
yUytKapVe1MYzDAacBX2aFXM8WWyTrKYHD1sKBa1l4xFOab2FJmftKzpERxE9pcqRGu8WUXKjrHx
m+dc8Z9gmQgzXx8OiM0FOj4hnMnSQgurZInmBCUv98TJeOvzeih/5hrir8jmnwGCqGQz3TTmmI9O
SYWR6EoRANzQRwBB7DUaMn1B2UtvEMx2T/iD95v5KdJptoWy/iB5TutKl7itxnWFTcInVVH6pmx3
Bx5S3JqZlv2wfKNiugF4+kfrveexFtfBRN7qpYpVGxXmECVxTm/pIaTuOlpDmpk+fOK7H0GTiXm6
XcAmiQo9Lb2wbx3SrD0f0XFkeOrCs/6DH35Ip7X6VYBBSgl6LmQuaSCoube3K/E6Wur1ZMfMTobX
rQuyJYPw9D/kjqNo75lCAtqTn6Ue1WSVbW8h4arguqdnEZmgrQNzr2RgGVQxSIySy5t+VfOloadM
8B82xkp/DSCZ115nO3z+QeBZQ84NuHoDTF4y5Izw08ackSur6Wu4DHJ8pHQTUd0FU4/TLXl1QTyh
2Ahx9TWTpR0Pc+J/sX2trIYt3wBpMXTK8eDGJBuMtSefhzr/BDG0M/8mmKKNRR8aa9GRvED9mwdQ
kgx70cXU6Wg+KEuhjrnkRjJsqjGiEVLl9iMCMilaci4QYXBjdDj01o9IrZgbGE+lzM01KtAYgoCs
5z2Y0bXOOI+WTxeQuPWaLByTFbY0oMTiN8ls7JI0fGPBMcIfH1pt4JS72sG7pHHaT5eGKBDE8OKO
3S69yXv+5OwF5LcLTqoaB2k2402mFJf5+TQeV87cUUCigsr90vsaiKFpjFoRw6gtHQNn11gPkuSB
wXila0yEHkKw3en0QGT7ABKuk0XuleOWgfqGtLOzFXPlLFxo/+KAa0lw2btIqYDzfA9jgeNSgOz1
tbyQ8wq29oTqwfAgvXZwpv968Vz0NALhHU1lLg9xFDxH8A+HLb0bl+dwTKHFJnd/az7zj9lBWugh
gyiGuJ5oVHYNKKY13yVCgtXQqC6nOX5R2nJrjCBjtY6IlWPjCZBYGIa6rlCobxeuTydQI8iel/Yo
eETQfUUXd/CTDpt5frx5WPSizZlaI3YPSBIXhmNamiurUR09N97wkTPx7QgWo0shMzzy2qDbuB8p
3MRBctd6Em7spf3ZuNdor9XSwLwcckZy6OviB+FtA3fi5za0KepwNIrvXHMvr9CxhtJLyvNQbQ86
pUs6qpkLutVrxpmtmFqeaROaB3gIlHSu1JSokF0qUtdhD5RZb2VaWywjtNkq0xa4P9ubKET11N0D
Ouu8xZgrxf3O6LE/J3D7WnRhwPX4gVuFIhKWEM3yGyqYYq3/+FEhkWfuVuhntNM7atZFk/IBu2ms
mV1KR4mUL6dgXOZj0j0jQXzAZj+FRbA9yJLjvYnmLboWiNuAaP/KPDWGjFftXub/8IMvTuOWZke0
yaLFdCmJhVgGat76Dlcj7fXY1qvWhkMf25xFbI2SVQOyYOYy/g9N9JpxCV6yloa5NlftpdwUoE2C
x17obwMtTaF0T+0z2tAwudutPsjQ4/VCQkqUYu1+w8+3XHULZTtbIboif7MRt3CaXUo72JjSMR/z
fBTIDFyeNHD9N3m1oXjBHOMbvBm365f4D184OMgVRDvc4tWKJAmD2zAyiIkFx+D3CTbUtPfbYfwW
lO9JobQhKwY+FQQnIfpIsAgc/aUsIx8YMxKN8Z9rz3DxKiCWbEixyUXNYBX7OOzWxJcVSaAJyvW5
UIlSqwNO2aSmcn6bOeQx8XVao2Hy25uMxP5QZsg6vG2c0/61c5ngdFQf/zJUV+AhDjZ+dLFJ8Cwy
tOxTfpZXlRCgvw9L6HybZLQl/tXH4t0CKjd2He0R3SYoZAS5voVGkZQOgZhIcN/IGC+vWZlF0l/7
Ek9kcd6tSGZufT89IslQ37sZloZVeOePyC7S6jXboztWr+DjjQ70ToKi7oEP4EVBd8l9xgoZFdEn
yY4BtjLOpzvLhfLRoqRUGi7RqAT2o64SOoC1Y0FSPRpVvnC4sg9LJyA7wrs84BvLwXQQwJkuGho8
jQfXcJFKH1lu37Ilj89FDo7EMQGd8xh/Ykc2gyIZsJfTQ5C7hV5zIx6pTftV27GveQe1cm9mrss1
+B3m5WUkZQ+WkY6gPQTThrqeU2XkDiFhYHmD9DDbx3YM3h3SNQcHuDgwhzya2XcTs28Gh4p6qZUM
85jZ8ccdjwltsq1LNnLxq293QueUnEkQURUTQT2I7owr/WmqrJ1Ut9sVFgSJnTm6iLuWJKZhJZjH
30ukpkDW7Hb9E9l5awsbgAap4GzcFl4xjajtYQjKcGK17rA2Zzpg9/W4+xOo2ftgMi3KMhtpxpYh
fmcKC0eWThIuK7B7qrLgOhqaX8fNj70M+csDB9am9AFHqvI55rqg0hkspb7bzdSfLRfJpdYWfrrF
t/z0UN4LjtGVDyhuo5ldIJ+2exZc5sKWHTWmHh62QPLG+4einQyZ3Ne2IPMk3JXZPv6rY3ijOESS
vvttFxuQwy+jjZtHFapBR+Gfk0VdFiqWkQFJ01HkcEtGMEt8McMeqDVbdkMHuIE2brsqcuERrBFz
UKN8hfblRoijsmMdozaIs1/OdpxPc1W/i0vlaFm4BD+XOUXERiVwOiuPOc34i+UueP1wdTr+A1wS
fq6Wt9RqQ3IPfj5M1repB0xOP5/C3G7DVOJn4hEOFEselmt5PXizy91AUOW8ch/4I58oK6lZPKBu
QQkTmZP/Hjgl7dOujxGTjnVXIJpa42hJtzo3Mn0Lv7RDBvuEDJQwRoCb+OIbtPcVpfXWREx/TNd2
OKbSNgM=
`protect end_protected
