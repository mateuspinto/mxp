`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
yzfwMXsDQzFHTguEFApOvi0AQO7DKHjALoSx+bfMa5AFk1x6F7V3LJP7vH1WRpcn6NCQoMybI9MH
OshlXJbdBg4A0knp1uSnAnX2bUVLbsPZHqUciFpaNVbSJVoE5l8RtaeY1bY7ik2dLxlxbnjrA4oK
UoSZp0nu4MdZ8GTaMnlUSmgHj1j3MO6kqy8L5tnNv0Izvb5ilcEMTk1GYr/ivgAos0EzKi8rxJub
BUdPJQi8mSzGr0o4VVOLnc1CnMpGH0tfzw7MO90rM1LK7fK0ckWtB/u9Ptl9sNFavJVuC3vz7nNk
Qlk1STvqcPOPktXkD0HelVhfNu/KwTqLclTyJH9RLMzFQMDD9mrKLxjFTNXrn5osJ0EkNOtvdtGE
ifhDPIflzoxmx+Th7bWP7O25D2jLx1iwjeYfOaEzO4AD188ZkV7kjgR28+tlx3DVH7Df1ECT7+mC
27Eq2MiyZQ8KQzdiDWcYTMDQFKByhU/QTrxSiSRgniAO5KIkgHwHl82ThKF6lm4yLeJNpt5jAMmr
/pNPyOUl1jyUhahd5pibxFzyxLYo9AgcQSpix0hW51eeJxB62vQE0fgGJC8JZ6uwCviDW2/rNFoQ
1NwfhVO+deKxTOwrIF/Wiebm5hksWQ8m9upCBIypFbU5OuQCqaenpV9bMICTujPc0OEUSFQo7JFQ
xsvNsZTso0xkTTnS3DfADMARVcgmHKWzrol8nBIED8yB9m4QZMkU0+M/QHsfU4waHzQSZxDyKUyh
4Ey1v/P/EIiMzVPWlXEaEh+zNH5OVBZXUlFOUVkc4qSkMUXTKJUspDnTIIyCGH08voKEJngZAj88
UGS+qJnH6C3bo392TXLXuLDx7HU8++cw6foA6+3Ev70KeUBtUHCHrymwOLODe8s8K1yJmUI6I1QC
ToLs6D6mo4HX4TQo8p6YBHA6eyvXwV9FBiSDb/xypajNIBSFaTvkrRhhjROpDA4i0y47jq6fMUH1
b7SC5EHz3zEvFSicNLLnZfQYrSOP+hyhw2tclvefnLS1G78RuUsdsxEurLfwtLRlcOVhpNTmOH8a
0EeDjC29LFvjxHGBCkhp/1blJVXhvNF/NiU4cHFXO6z1lkWSy8o2ASeB6Y/kK7gHWGrow+nlg5mg
grMglnpfi1M/+y1lPNpSuzFcOPSvHT0KqVHUGRT27edA7uBae4dKxRIK+w0C6UOD7y+lb8f9vlsD
wqo8CK04oevm+gxt60SyawPKHM7iFBcKiLTzGCXJItcXxAmtl1agF5Y6T+x7TIThdaZkV/tn6Cdn
gPf4dGN7vxPz4ZZdJb6J6ELQnfpAt76Lkks09gYqhtpAv3UgRpueVadF2rV4yV2eQqYOT/n0594E
EBYX2FqCPKrBiI+41tMEz1zg8slPPsQ6FYzCVYTcSFVmHq5hLLoVK//73MOR67rGYEbAvzivR/58
JRIXISjzkR/IEBMr3V1JZEd1ZH4mBRSf0uFVa4U+6ppisBwuHw==
`protect end_protected
