��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���`G}Ftv�V\˧�\�4x��F�g?�y�sr�D�M��g�oJ�|,���a��p��Kp� ��/o�}�`f�=V�6R�Q�6�ߋc���>r>��E�EqSJo���{	k�����?��i�����w�A8ɋ�.U_�a�mq$Ba��F�B(��`�>7&{�D���Q�l�|��\���#
�/�Ix�A]�x�5�ؓ).�+���"H{N�z%Ԯ;X$f��7�z�~��õ/0��M�@;���>�;�Z;�<��#lb��r��>\m��J�d���"�ߺ:���{jh	A�8��5�f�\?c�im�*����\�~D#�Z����&g�W�E�����[���O®mp�t1
y~�3u-{Kǲ�)�����B�0>�rE��"'^̀+���8�)�K��z�Rs���C9RE:�-q+�߶�������Ե���g�4/ ��w��xKf�����#0�5w�o��1xa��O��.U�u27ڦ��*-T�K�_��q��`�����X����)6��֣�ԤɚgLyI]��
D�r�ze�SP
�:2��3(3U��G-�_���,��G�n?:f�#S�����2 ���݁��$�(�j��^-KY8��9��0��VY�,�^G�i�
�} *>Z�T5��GS,����O[���N�Rϙ�\��K�+O�2��Ydn�H���n|��2��& ��m��s�(]Md��)Ķ��h��.'�W�"N�mP��,��R��*���N��L���c.'�q���ЃC㨯D��թ���}�zGѨ:�oU-�+�Ԕ4C�K����p��V�|>����^
�=���?ۧ�|����C  WSD䄭T�>k�_�S��\��3�*�{.��Uz0�:(a��}�~j��v�H��og��r�)up�N~�(:��6������F�O�<s��ux�r��	_��F��f�R���O���j'F k���}J/C�竁z�y�Ch&�=�3� ���. �a/����7~��ŀMw�(+��K�
���p�j�	�" ӥ/�ܿEx�\7�@vD��:���C�V\����x1<�<����@���=\G�y��o#�G��	q*nEW��cʵ��-Z��	�'��bf������4�&x_Vh����E�-�֠�����c��־3�!���K��9�B����'l�=�� ґ�q��al�O�G]e2tO*��l0ӳ:�њ����2ڴ��vW@��Ʉ��� �!�d��h������Ճ�V�&$S��p2iD�X.��V����몟;&�j N}f��{h�����[�vT-�N�	�Z_9����V4�L��[VoqZ�d��� ֆ7�m*���R�2j�\[�E�"�!���K�՚8ۓo�5�Ĝ�F�ߧ�/s7.��F_mԶ]���s����!q�ۇ`Z�3�4[��y���BQ�X�ܞX�O[�U�R���5�G�~�`/�Ʈj�2�O�&�Ose�aZ��W�`�ǎ����z�������y��It�vx�s���1�4'�&��ƪ@~qe��'�p���n�^'P0�+� 4W'�y�?^�Ć��$��]�w�HZ�TY� Kn;:)*`��ե���S���.	޷Pr_T�W�3éy�ֽ�^�lvRN';b6a��@��Vu�n�x�{��T������E�7 �quu�+��xs���g~���&�h��|SR�n�u/������2�m�/Z�-��ZJ~�'����4��4����)�/X�\>6yx��
����o.���wr�s���U�e폳p��Z�TJH��K��4���0H�:,Šb�$�X _8��/�i^��)�׬/��A[V����5fYJ�i�_�çD�)6�i�Rv�V���{Y�]AUq�d�,��X�>�9]����(�ƥ������E�k4��*@)
�"�r/���/t�~��1�}��gLj5vyn���iDq>y/s����?Ǒ4���+��{^�c��G"�B�JM�{�'=z!��0�oJ}*������nڴd��IƦ�0�H�!��t2�Y���v(P��C����C�MJ�o��^A�M��GѼn=]�c��m�<T���N�E@ӟgM"��ԓX���j:�c��^]�9/���s����u�2��ؚ�lJ�c;���%@ȋO-�Y��덒|�_^�<�#�n/gβ9E�91�"���O=J���6u�tg�j�]�����t�!eG3�rzȳ�3�a"���BmM���]�xR�'/������8!P��V�<��)�]�7(��J�~�v�{��?3K��=do@�)��$��ܑ��ʘS�`-��<ã���[N:g�2��6����C=�I���Bl)�tI*��G�e&�Qs��N�����8w��=���!fa0����T*\����q%��2tc�=D�	=�!��F�� �*�h���K���۾�&��=���t�=Y�l �mt=��HCw��6�vb�Vw�#|��g��q<V�`�Y	�� �င�m�2��c��I.�^:Ǉ����=�	�E|dM�9O(��$��7jLR��$�ה�WeΎ���~���D ྙo���֨|g�Q>c���1��a@���pwk�+����<�����F���Ϣ;�%�TAc��}�m���|%e��N�c+�r���8��v�xh�1�(��C�ܠ�9@X�wSc2��J��6�/�`�8����̴2�ŲY(������ծ��V��\L��� �Q���tl%:��@��]I���@߫�˧�]��glR0�V>MWXg���84@����J���4��h_N--Ec����V�?@TD��������$�\ө����с4T*��1�0/���Y��wO7_�h�����S��ZT#V���7�
}1�W$P���}B���<0pc��~��	\R�/:���-Y.�b	�#푧�Ru2K;��
:�N}=	�x��́��M�Ҹ/��ۊ���;xn�,�������T��$�U�@!���f�#����c�T�o��[Dj���c���ⴵ��R]fU9&L���"-���Ӡ/<��s��.͏�)	�a�S��D�.'G��n��k`aM���z��ξ�U��LڌD�}�k�!s��.ɧARe�-���TZ?��D�>�atC�������;�b��z׌�ޞ%�1���}��rJi-*�Ïc�ǣ��hV/=i���e��nj[n���\��XU��ʄџG�6o�6�?~�n�Q������!K�`���d�e��L�=�F� `�{f-����gՕ�7��P�i]�r+�ln{.��}��?^��E�L�����T2\	�٘�ܾ�T_%����xՋ�k�4:] c� ȫ��[n=�t���G:h��a�y��SA�����,oHr�E�L���N�R߯{CCZGrW�]���7Ҿ�U�ŊC�dZ[���H�/0���OjHk�1�;L�m��t���Y	��)'0�b�悳A�[l �m� ̹�jXW���,H���[������#���|pa���TlHKc���@�3�d���7��'N@N��?m�!��α�ȗ��p�!e߫��G�\g���L��9��Q��N
Q��D ,�{Wc��t��RS��.�C�0��KȽ�7�7�M�ѷQe��<�IZt��L-wbr��U� v�Uׯ^�k�D�]7��a�����>�Q)>uN7J]�4��=ˏ�|!�m#W&��h�V�D�Y�H��=1�X�p����|��x߁�K}]�cU�@^<^5#Fx
C�SE�NjR�4�!�-�D:S�c�o!�v#4���̅����8UUw�#��#�p�$���K��ZN(K4q?�.휪�{9����ĺo���O��ۢ��{�k��gԉ�/�Z'6��;��C!��#Oo9�#ꊓsJ�d�c��G��V�������J�}̹�*������r�.�g��2��
-ʾ��!�����lĔ��%f'/E�����V�۸�ۡ��_Q�"N��3�����<?%���sƞx-|�XM�vW<j�y�H�*�_��V���2�J_�L����<��uG��J���&��,:�
HpUPc�5%��0Zc�u\�w����O���r�g���5F���*垍�Z�������yS6[$�o��O!�Mq�O�W��)8�j��hnc�\<��_�YЃ�6%�r��8�N���HZ9�	V4���-�b
/9�89���$�.�����3��#�L�-��c����I��"����K�e��M�>i�7S�\�3���)/�f�9|̘B��!�,�?߅\�G���rꜻ!�������K_	�=c��7��9Z}�1sw(�q@2�A{Uo�c=1����O�&?�����Ի�B�����F�d.���x-�6:�� 6��O�q���g�+uF
n'����)#5������k���Z�]�,4����p���@���å3%5�����ï8?ݎd��s�Ej��N��NK��4�j�檓�s�;�NJQ�1�r���L��?�Z�c1�@�Ih7�U�Y��^����\?�֢I��� y,�E�sB�* ��]{6w�]��~��X��!.�*���Y/���ǭ��S�թi^U����D��DC��ac�2��qgn�B�=ߖ��g-�P�\i�4R6�v�9?1`%8��.|1�$&�.r�uΟ���n'� ~b��Z^f��lxa���1Iy�?�	k@:��e�S,���e>g61Miں����O?�_���,��8B�Pv��u�@f!�(�@L-�0��0O�4��t+�8�e�n3ٹ����D����c��ꉯ2��c��H�����o���.��K�����#F=s�N3�KX>�����g	����ce�ΝmU���ТrlM[�f�#�~��H��c��#�f�����g�SN'�O|bd�4�A����i0��5&�he�����փ��BC�x��\���kFJ2~&���EՉ���Oaht�����1$ҿ53��`8�0dq�5k� +#��ܠKiC�H`��G�b��G3����1��w$�t�tPHd�䄣H�z����u�]\x��F����R@���T|��9VA�O�M�ёŠ�رV�eI�;�����x���4fqn��>�T_�zO��_YǷ|�X+Ҏ�	_���&�+��DÐ0��C2����B2��RD0xp�����B��	�<	�q@|L_�r%xf������wl�$;���~��h�$�!69��Ԣ�5\��.T'�Y���a������F\��JX������+뇰����YFa�Q�����y���y�-�j���#K7�v4�^�����u $�>��
��oR;s�����P�j�L���Q�Vj� w¯��x˹y���H�6�N��'!dy���������6���T�&kn`ڂ!^�J]��Bwt�hec��N  O�@�AL<��<���ݭ��Z�i�)o�3�tw�]=�v�$�4���D����A�f�E�j��Zv�r
���	2�������/��)VM>7�rN�`�����a�Z̸�<�Ky���ah\�+s��Y?"��)8E,�("�j%&֚]=qT���M\��nm;��p���k,夰v�VI��,�6Ġ�L����q"כY�l"�a����ܽP2�F5�����3��]��Md�/֢HеX=��7S��cR�u���ջ�׾�b�)l�L �\tC�f���ΐ���wͣ��|�bh�^�`;�ʄlF��!mě��lXN��^AS�ɺ��ǫh�%�?�,$�����V����p�T��ޔ�>N��9:�"�� E�T�5����T�E>�&{��PW�DAd���D(������ܪ:�H]�̉��0�ܩ��@@�����N�y��%�F����������\�_�s>-lJ�F�����k�m��dP:�o�͒8$C'3����Qm�%ҏ�$���>ud�f����94��)i�S�9��БmX^�+Z���M�������Qdm�򟪑m{�x�����L)�?4���)	��ߠ�g��&Fj�Zs����᪕w�,Md�eEd b\é8�f��o���=�S����dj]�Y}A��c������)���a��Ns j=I7; ��K1CL�=�%�nC�wO���З��E�������^O�r��f��^&~hf�L�!�.�k���RP �X<믱#��t���m�!,E[�{�Kۺ���7�B�SA>��0l��(d��%"u�?�p�Ue~�+~S{�l	����������ӂ��i��b��,�O�º��^��P.�2�]�
�F[nr�?�e�Hl�j�MC[��.�YV�ً�I#ʒ���`s��
G��H*}OXH}5�{�%�>]$j1��F"0
 �i\�Ŋ����3Ì�ɪ�!F0�W�-_��e#l{CS�`���v_��{;�fT��AQF-�����4�,�	e�`���Ŀ���tpz$�{H'Y�ܸ{#� �����V:��]��Lo�#`�RۏZ������ޮ�b�
6F8����F��pL&��0﫜��ڍ��<(��f��M\�:���vY%�2��a����FW�-�Հ�t�',��F¾Y��[Qs~U�?�g���������~�*_������qxL��ڰ[2��MӽW�y��>�5q��Je19|M�K�N{J�y�W��VGy3�M�[+�r�bj>�?xF�嚧�yF���8�v�5�~31i�/̔J�.q�m-T�+D�3Wu>�`2����J^��dv��k��I�D����Z�=m�3� ��f0�ն��c^�ѕܒ�	���;���3�8���b��<%��'b���N������_W�4��\�N'�����ĞJ��nC���ހ:@ON�� �_�k�Ι��M#��u%P0[��e��a��ȼ� |��eI�Vݢ�ݓAQ�~�ݓ$�_�q�G�\v�Z�"�����(a��*1�xwi��Mm
���F��5B�E+����x�I��&�Z��l(��O���4˰�[�1?o��+kk)50�k��W�?\"O:�E)���=�GE�́mpa%�͏�MT@���m� <,^��FsI�.�lND�ޔ�/�L�^�1�{�C����|����D�c76�{Q�]ǽ��BO�M���/��Dq�D�ӹ=o�p�뀱:��&���R̰����'l
�_t-Z��A��N1�*x�R��yP��<+�Z"V���塊���Ş�k�[f��gO�m�����#���B�0 �����{'$L�/u�ZI��I+_Ǌ1��I?�֋���v�r�L{Z���G��@wX����&�����3ᗷŠ�m.��a���S��Oq?A8Q\	 �|1!0��3:�%��ag����ʒ�Wi������5�QM�=�U��z��}i�:�����Ɂ<���p4Ѣ�[�Z�i�Y�y&����9�"'?$~:�gl6j��<;����P��7��[� ����RV#���dc�������=����!Gu4�� ?���קD�³���ѫ�pϳ0ʸ��Gdu_��(���bxW`��\G33��|�0
G��s���&��s�?�>�1�g��eRgy��I{F�r�\f�.���Ȟ̱��&F����1.h��RĪ�� G��5��uԳ�)��U�DB4�1��aD%�����n/�0`��7�Ƭ)�Ճf5J@@S?F1����:�%�N�@���D�7"�-�*��^g���]}� {��Fp@|[���<v�+���m1X�+�mq�V��C}2]�|�d����:�Ut�"��"c��H�^�ò� l`sX��X<T��>��8��E�"�0��tW;�(��\�-�9A�U�9�D�����k�c��'�)�����[_���+u�UXg@U4�I����"��1���Y=�i����Zӧ�� ���Y�0-K� �D!���OY%^�x�MV�.�K�Q��ڬm I9����;y���{ǰb�A����B�Icb�*�t��1�\�0��Sm߻*�ӑ�'u��I��5��,�Օ��[�U�#=ވ}�ϵ�wb\v�V�R�T�Q�=��2[0��:�}_����}}�zIW���v��.�=vjjv4=�(����|�}V����Op�5Ysj��3#���G�r.L��r}DO�\<-�ͮ�� ��:	ɭ�����\m ��6/���O�lᔱ-`�+�~�HV�j�E,��fd�O񈋪��G�+�0�6t�ApŦ>��y�;�45��s����;�:�_G$��91�s�T`[),C������<�&��@�W`S�6�L��1 2�����>�,9�Z��f��>l��20�� (�{ge|�J)R�F}��Y���m��<p��G��=�����N[ֵ��YRfƼ&��`ᵙL�T�Xͳ:��]���ciY�a�����y�B
�H!J�x�D8_���HF޾|��<�-���B?�2 SV����)|(����ÜDc��+4���\��&yJ�l�|Q����_C��'��=�_K��ώ�418a��vI�*�u�H�Ӭ����\�f\�\ZH��8�&��]%bO��aI��<C^�,��ٍq�G����z���������{^?��)jp�eUg~('�l�,+�UI'
��@�{�e�i.�� �	�W����v���M4�Y�E�`���P�4E�� $��x�"[�B�g�7&j瓻A�˓����I_��aԁ�7ɷ���<Lv�5�-��_��
k���RT�}��{'�o�fj�kꉫ��>���hߧ�� ޞ�Hb+o�Ylk�<�+	(��P�1��А#��ȃ��"��_z�X���o*C�98��Zz����_N�l�/����Ǥ]���'�GEF��V��$���6H���.(��%e4c�-N̷�q��1�T�ҜR���~�\�e}�$��[H�6e�j�P�
Q��፼���'�Ө��g^��à��,��$Y0˲�9��QeC�H-��ݭ�}�u�n��Eg)�_W�����MA]d'R�c9m�Ad���ˁ��=�\���Q���Ck�<m�UJU$w|*���^&q�+Kkk�h�Eci�/