`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
GYvATpvL4lWNSRdCp1nHgAzwBp3dEEuxfowsM60KpAOKkVeHEcIHcAptqemDhp4WDP5QR5Iv/8aD
m7J4wa6D+WxIxv4YUmYfuxeHUoS8Rc97NRCo4Grwum6qz9MdOY3MZZYtimDiOFObsinANRKGcyrI
Q1x2IoPCc0Rsks27yI4ISyl3jUBOaydEZ97pM1DEJoK5OOuJAcVYM87i9ipfsYfGPfDNSUwqLyUB
FU4DpPWPpvdl/QaPNbTcdGtA6MLiu4Y5DRBb07rRep6/nzQ8T7T/3V8SpSyb8yzinPdn72qevVaZ
WNNTyPBQCae8m4fkZ8mnLAIQGhftKMBXifR4CQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="3554XKrqbIAEhwz0g4Hax1iUpMQ7XJ97BLSqF9wMJ7Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3600)
`protect data_block
kVYy9JmaBy+EZr/uf73ChBQxgXpiLtqNgKJUlGz4Gtx/ceuMopBmyC0As0ctRDT7neHk1xrdAN9b
eqCZxi6FBJxcaiTvzDpL/gWFWcLGyoFUYvNQsAdeZLMrcXAjpjHyq/Kg7WmcvVbJN9eYmrEdBXjO
WK0AP9MYDrrjCDqrakvif3A3/yomn1YcI0ziVrLvAaHcH7YeWp7IjmaWRtTK9uc10rNhwgz2DfIV
dXsplQ5ewYNC8p4Lv50qnxsbHU6ItKrk9RoONX5VrkN3qaRT3qSs2Oqom8+Akgq1ncLm5rKCs0X4
CLJkpYqHjdsoJZTezlUny7hazwL65NOamI8lQ+twJo8yl8sEe1u7p6TnqkNE6m1nO3pDMdF7kEMQ
ijPpTQoWvZHvbfD8G1WFAxXEL0au/sRGBq0GuflV4tgF8HJFHW5O5l05kImUA9DaslE0rij7rukK
nTfYHQiMcdezRIfC+KgTwaiDTJiphJ/jOc1u7eCuRruN+OTP4CMBzfAQMP+QdwWbOo7GF5jGJJCd
GYRYj8Cm+q5dHPkbc15iyJM/w4GDRdLY/ADaPUrTdQY+qljWiMdrlpL+bGnekEFnH+Gwg3LWxx/7
Ll23hcjbfxKoVr4+iP8c7z3lo5Rzl8vzfWFW+wIHq/OZovvWjNCrPpBxwYb9he89H/zzQNj1E/5y
4ojLXK+gTDPEZnaFJI7soPuhaVYPvs0m22MRGwWb3qaBeU/ToFgaj3p833Y1Swk7DuTHWaYjffxe
4kMzvatEFH2x+LUeW8uHpgxDEADiMz7d1Zr7Pn71rLNRAZCUWTe30WkoRQYzYZnSdrVQhzgOnLZQ
14ApUIXKPCb5PM1rJWj4RcOsPCSbqUW5Db0wjZAhFbkh3ohOGkyYwrtaxBkVtljDp9FEamT5MJey
JDlRa17ichPsOhLOIdqbbc8dbP6DpDSwQ1fjKrz/qbz20Fi1IpbuJGO4NfRTYHDh+pu4VuNkYL/A
XxxDUfHxT+bj7fCeSZ4DTt7+WBiXAuRVEUnxESkFg6vcugcs34JJiavxyXlzyTWusf6ZWYtngVC0
kOlt2F/vCm0crkFAmyBfMOTeuqOlXecCvXgf9RHyqtn3viHgX0eWGE95JxZnlMggOpYB8WvmUc+A
0u12KkFxAFO/WbZ+td1I1DD7CE9IpygENvc5DgzKLj6lhza12ctQ6nY2EWsqdsaB1D+6lM2WXqiH
PccPwSQtjs1YpHFxgKedv6Wp0+sOrBXIYgKEHIL1gDBtnF64lJsrwlDpdqHyj6fl4GxzPzN72r5l
u4H2i9Jz9+H7os13kPLHk0B1TNuLN8QQo3Dc2LhPvwoTDDkTwHgldLRMn7bDIcIwwjWzL3SPYbTr
adlQcyjlP72OWvsinBmQgPOhp2e0C4+a8dcZW79GcUS9vstUxvpCeChPOb2WwcQ2mEAwsA9bPhjt
9xkLaloZXpS+KzVbmreLgLeKvtx5r9H4HPNu/KNnI46h2LFTf/Ve7a1QuFARoQrfflLb7RKHRfnx
5Rvoy0jCw1DFlo95g3NOGKn1vQzSRCb7CEDJz2adKfjrYodWFz5TTYSlRCP+LlVOx1StoiWDP2Ht
v7GgKdJyeXZxllmnXSqByfFWyArTRvbE+Z45XI6tdvvDSXIY8JwsmVTruHV7KWYjvqdv6WdNdk22
BaYD1SPcjUHEirEx2DZe2dhOMSJ3tsszAYKdvkn/h94MerK9GXv1Zo6Pr/CXjgDCsO4UaQPtR3a6
0LrpLL0vcA8neuhlHegi4FyEfOrxjVOFonMlE1RN1Vo/crwMgb54xotzggcPXnQuAucq5IPciuCl
/ZgIGjhCcb4ZcKWEmGn0PUeXRp60i6XbwNFTFKeqkiM4h3F3tdSueboJ6WCBK7tWZlM6/4hIDrmY
xAZ1jUJbYKwVq/Qr5PQpmFwBzc6U+4/cA6Tbyq9asTkCznhYJhLkn5pJK5xMvUbExOCLzypobVgt
rGpvwQwth2TUSSUP1xjruxZVXVFWcb+EpPnxC7ypwNPvJH657MF9OCO6XwM0F1Xo1DN3LSgSLYQX
ccNOlicGzMobjbpus8/XiBbxyQUvrq0QOJZd4C+K1OZoyn0uX8z3qz45OKfzesDuAISVjXKRf13d
W3IPVouNvOxh8Vm/GKFcUaZ4jzXwk3U4pT798vMib10mijHNB4SL3DPBCIVpoj1O/WHV6cDZfV0Q
Jaxn+Frhk0pdWI1P18Ga9ZrgEH8zEJJJ1TTCo7/viD7BckVjOah9F/7Wy2n/Vvi+MQzBCg1UHoKe
ewRbqUs8BDABJhGBy+OyHN/m2RmqmMAjBXdcAYh8l/AMPvNQMTw6m9LUdCW6Hy94BHfmbvIyMCGj
j9sdh4/ZuuCY5lU7yw4YK9I9LNF0hTP5qUlaxpUFfFk6qx3VSFzDwT5rT2LkwUvq7tTvbKoC6sfm
X3UoPopv0nwnTj3BW0nf5D7lIrIzmiRUpvmedKStbQ3ZLgFJHkdYuoQbwdKljsjkSYIoghDPindX
V2w4RDhAj5n6ZULWlAvqt9X3YdnO/osrGVwaTnYvoxvTiZVS5wycru1809mOjRzfo6o+CCjoZOld
AOuLQHDOw7OvUF3j8+/8TJ9tBhSYeTJd326cu1/Or8WBuhF4jWTk6Yw35oghUh5GBt5xZ/Btmd+s
gPnx0U+d0nrTcx1NDrNjX4ODU87IR7NUfmASZucEWRUpvgAJo6MvcXePqv4KFb/BeVnoje0X0X0g
Kr6AvfbyB7P4Qau2JMnaYC2q9qLANjUdmqe5Z37wohbpQ6Tgc3efo84h7YS5Yd3BKVanM0uwf8IX
/Cllfgx6rHVxknMIlIaSXQNIDrDIF+0VcvZ2FH0Xvb2ujadGl9NY4QtmQtN9QVHQ2oQOJ8TOQADh
xf5/lyUDhqJzQn36zcM5+9hdSgIBYL/+bPL80FtBjFMouKzCEHz1K0jrqOo8G3e05RK/XvSBiMj3
UkzQYsO0z5CxOFGw+XX/OJyyHGCXDZitTcLfCsJUn3ki2qrzLUMzbeiquC8CEuxJcKPiAC453iDR
cAxD9FYINpsavro+Qa6m1Alm5gzt8YVZ2oudqi7va2AJQp/Kw6Hs/eY8P6HfF3pkDO/rOKFCDgNO
sXZEYCc/AfrxNvVJd6OmAifFenxEyihYPK45CDmrxeiWdKpMZyTDGrjrFipwOPzH+9tShrAShm5I
4phaAVXPck+xaCX+qhQGI/WomVQJ5Yz/EFkO7yVfQOMwwy7gubLB6x7KDrHFU2LWhqvcyATgS1rI
zsX5yEUIcOmyU3llio3XqO0qvkbocmZZDjNNPUI6wtWoHQ8Hto807qT+e4E7MYySJW61jD25tf1L
salzizDd32j3bckU9l3O2tmZkk/Lxe+5x8Uy5J4OEm9SV8ENMYPqaiLC8cNEctxg8Bi/CUD7fO6i
FTpBuhZHliGlnLvo8ParB4LwW25kxnW1mUUOr5BePitNByCk1qvMjmNmON0cbuIEoAYFJFse7WzW
lSUD7wJ8pwmL6A05hAuB8N+6YWek1wOQe2MpavWN8n9iPJVA6twLfIKUZVkwEM0FxHON6/ShlNos
mdNWj6t8uuMVeszXy8E5FbsqaD7FQiEVD7P3XaTNWHi16G3fd0DkD3Yj4ATAESxG3Qtu1XYWzjah
wNvWqSW9ZxxSWlseW/v17pfcSbCDebgZuHest+zstA7nLTfiUR/GUS8Gqqr6iPnmVkaOMveh9qeH
3JQvlbd5MIPkfOmh/X1e6tF3Mdnk+ce9/hJ1+CQ1zggmreCpWQnz8SVrHeRtKy0KNniusefAyvz6
vr7xu9mwYSNs8WUrJgzj1nWtcDFs+xtu440zrGWZkfCNAnSzZ7rVyau1QxxiZgbLQhTzxvn5nSST
ATcCNV4z8gnuC6YMxJVz8a5Z1ddN6dIQbJJo2i/rP62jPUb8U7i3gA9vv19bp+m6R00ThKazG8B3
wv8x7AUOp8kVMpwW01BGQgqP5IPcx0CvkmwC61u5PZykA8bwhFELJfuX9WG5FvRFV4gdUnKFc0Oi
PwEwt2sI07mSWaGKjZz4rCXDgapAfLs537EVcHLfdyeSsVfwBVxPr5Dmuuaac1qJqHn3/Jwh+Maf
3uOCF86uoy2IRecN0ILBM7mr9nWTViApfo+u13pdplibtMlSut7J4Mk0mGb/OGJiSNksBSNzNGcJ
2qGHyXEKUy6gE2piyfL/vKZqh8OO0WWToRP0bFuUJo4kz63z2giinUUiEKVx6CHYWThzTh3eJLId
oS8DjT6A+LhQwvohhCEAk0tXgKuPyuu5sSFUU62BTtimdNCcC3Eza3l9fZwQH4uIHNufjFxbQMpb
OGxt9RqlytNOXOY9Jq8IhomS3GaS0B/0pg4ivNabcZZ3gwacO/EAP1pp+FIY3m9MPtFnoGD5mKuX
tuUkicQ8L62f11hNFmJvbV2p6o25Hg18PvZKQm2OWG90V024bSMGU5nsTIxhxb/GE01OslRIIrSa
ZFzXV5YbQvGaGQiCXJMY04cScfgMrhjd2aHRfC3ZTqBYDiaEFsGQC8JLxdE6SpEwUKbZcrYQ5KZ+
HZ9JKB+PowpbXYQd83jMDFS3tEU6EmJMgxRohhUnmeKgKgcaE0/evIsDosd0Q6HcUrV7iOptnNp9
45GgfmMnn1QhH6RmIUMt5ZFc1GIip3W/+AcVuN3aPly0slSIwc9C2nvQQsBdx5zKX1Yhxc3AjJTQ
+jMUuYCRLsmXz72Fv4HxR39A/BWcTY4D+CkuybkdVdVHOJiUdlq//99XFs3dmzKEc8o+VE8zQJ9F
CZQyUb0xkPI9
`protect end_protected
