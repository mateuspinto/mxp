`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
i9DuxHcNDnb681kuQ8051JXZhvDgEk+Dfs7eyvHg49eZGSZNEotagt6hzke7n9SRgliln/A0Xm4N
riM2w62f8g4jA7v0tx2YtiPMSs57rIQUhsU7aqP1BApQexFqttA3ZHoj6CXLtGtZLFbxYCerbQGS
R73IsGv01b8iDmqYotCJ9kWS+c5Zq0J/3UFfYT5Lvrvd+ZdzlpQQ3NkHwfLFvrZuS5iAz+R9dVfe
JufM3wQrZbB0dwuseca251rMTM0Td5zKvmkTHWBy04b4b1232iC6g5kPqrjZy49900xeGSYF9UHy
j9Y5woiOAMCO8nS/rzWcM84VLDfaE99VvFRkooO4L4VCitpEIX4KeGf4XlAG80Q8KbMYbgZ+xCgn
W46wSTmqAUJtrASE26SbzD4dnqiDxlhxQTmaibT9kdpBU0eoILXEwQKvUXqrHCHEwbO4kvpWTws6
q3HIOcpXI0St/dNS6LeEm4+FY3PVRgJPdIzqB5B/2wyPd7WtMXOkrWLn581IBIwlPmphTg2+g+PM
D/LdjxS0fl2zELFD48wJtfpec7NT3heBWLicJ5uvuyF3CUo1Xqbkl4seoimpSJHiDhimznf2OwPW
KmWt07icx3Zc1sZ/9frt71No9u2n6dNjLtvaIO70NGkGEzIvRfhv+qLCdkr7jWTytiB/m5gzF5YI
viYwKXObzxs+offzy435fTw+jaTsFm7Bs1obqd05ONnAKBVGKJCo3vDW26WDcnfpzqN4wvRNY2XO
xWuJ2l7v6lE6/Uzlxy1b2CPi8pGzLwvPlzy4F4Cnk4+Al38vxM47e0V42de+RQ7kCOQxP7Wq+WWj
4DS/XWIzPdWCFxHxyLtvr1ir6DqVu+F6VEQ45VE+SUXPZrQoSWeI3dvxwUpiCiZl3ml0qK49j/UN
u0cG7DsolAW8/oO6Gyi6D4+qY2ENlZTKP7kIqn904iNpOgyLwdsnDkCQWh1IirN0ZlBptyO60l/1
uI5EDykMBNYulYlVHZFBjZauV+aoO41PIpcVeaM/edyp2C+nHAljWw7z3Z8wpLq0QxQBLkf3/T0o
eEPXplgwTMslIFMoCeqbJ8S+6ut+7jpozCgaUKPx9/qeRnSAkF4dpIS/t+ZV0DHxVU3BlVNB5GvV
Y+G2OifHVHNjcy370TK8TqtNXqU0kRmUqTuwGA/UyDMvw7ismrQYqqzHLLQEPeCmtNgqOAs4AQ0t
Tl7FFju5ECJondPNRjpbUaF3E52KasHhFpFpajOGP2ezCL20qanfKJaOnjDBGAm8/qDxWELeccuR
W0SHmMqlXAg+/M6oEEAi1kz0LbtUoE54YiccFCET7yEnUpYyjv8MJx3ZT11aujZ6ENlU1zJIOllr
bHjZQNU8rxpdAvzJBhjUGo1iCttpgUE9mpHHxMe4y6cBNuBDpB87NmuiHqqcyFP89f44HMpzVpXv
+Ibmo6UnHsmfbKhKRLaduRCwJZapKGWLFaYTrUg6WAwyn+D7WDB0auVUXL0Yv8S2z4tRFNkffyGA
87boGOHUN8mWVmkwLcAficmt4ieSf0EHw6wWcGR0DJXk7oCRkbu0O7QMfMXhU4CngMi1eR4Zs+2z
UQuc0idD+Hmt14WO/K6kAEKEjdVHMYJeA/yeahRJN5AUfzf9dyhUEIa2dldwMjG8hEp3sSoqCqHo
IW6qERZRG8tALTJ9kz1lCtbdlJ4txVck25rqjbY1BHXuiaqsw20oAT/SNYypV3kOKt/eI54FE7E8
TksaeX81+veYJv33BB7Nr34Nky96e11Q60F+d1T8u2A9bymjgi21JIAtFVBHsc6rVgkqj7HZ4/8i
yDLDt4LsHmRSC1rfl23b+HXLXM2sUSVAKML3ZrjZzzdcaPBCrC5Vvpl7keqNz9T0D5jRtThEL606
i6XwDmPhza7Lpm9PqdLle6qUueG054yGGThBlzMi02MQRBhe2zHq7OazG08bvbztSBcc/RtKTeeJ
NzalACCQ0lG6+scMy3/+3TCuP4SFrDD/+fiOvX15cwZWKnsBDB6amKs/kN1k0e69NdjJ5SH7K8vs
HKDfTELb892FmN7xTn4oIcOcMAR8BtSXU8EdJR2JCRNry15WCzIqhbLhV+e9WGoUmtm2mFmQeaNP
+0/Pau+7aub4KfrbMNl0sHIt+GNBtIj+rwT/B0ZVwAdKMo/LaU/9aW7p+GuV8JbwTfJmUD5y3Vi1
PfHOChMSHrstUXWs957QIlZ++0Lf8Bxonynyq/HX/1r1Z55A8FQPTjv/G3ofDniIDXohMjX2yxmp
iW2EDsFupqqxyfaZ/VXsF+moacNrfii8QX09G1x5J3UmtYHilRGEP6VGsMQXISYLEqhv8fzRGuBf
psLX9NoihG4GQ1Q1ihNjX/uE9zcXJFxxrNN8GKVrpxNfhvQPxI/5CtPrk8ZaliMBwNYLGXbG6/rq
y4Z4FvgNY+aN1IKNLHNFDNnS16L5fxPtXeTLBOA+utRBoZFixSllyleNdy21XQxv5xSWe96XjYJj
rkgBYvhsZnj7KrISQs7N1oNcU80J3Nm6ICDtnF4bGE1VqWK5gP0ObNwVyTIoqPimIhiMyUQL9CfJ
rYz6ncGH9mDwFSt8hFk7KbMfW3Dmd2Gsp+E4q5RRu7OVpoG3wJE82zFKB56pHBiYesCC26CvDc3h
ZWAE4Yor2a7351cnjUepilFMtkpHZRHgQFcyc/rhalfsKGIq3EX3Qz5wbbS3WjHKyFghQwC3FErF
V7NkP42EzNMK0hDEWRORyr8i3IHv5qR0DdVZB2MzreUhPkTK7bJus5GbbzL4ahiOT/i0H4U0oxK3
TjDQd84ZC2cAkVSk8oEMPnEAWj+aw5Z4MuE6FvE+3iZ5Lk6uIjaUl87rjhxrZb42CIj5A8KpcybJ
9r1UMoeaGcBdReuHK9ZUigy2GP4K/tx3gwF49EY2N5ByIi03hkfp5EluCuiEi5QHO3+DVOioqnu6
G2CVIAKGTy31NQrAKklCL4GLDaXbpvTVm4ug2a18q7aUp2xzotMbC5ATyyM9vZq9rw91bLmlTQ+C
+OZi+KWN/QSbvXul82sbrpa7OvkJui1Smb6oUM1O5Kdw+OU7+UXXLKVhjpUnFoJOB66znsjrSEli
a66v560diQQAZPd8WWaFKDAkhtI4WT9gpOjydCNzuL24qgEVPJd7CE+2bIHfm1RytWZbwi51vfUK
l71hKYB51QfgRE1GDXJuz6MUi49Op9PQsskNo65jBJciSEUBvxp+yBDvngud48mnFSI+D3YIuENc
Ch/hN3mTPmZHE5TF17/y0GCURQJ/eRPfhiEZ560nlxYlN55WwTCcW9gNZqGJDHNEr740NF6nOrl8
od1hZE83bcGtyylEAzlYusBwV9c15yB9qHaB3x3mJxuKg9jwnF5nvXE62CXbzH7oCM+7PPXQVVHR
wNcjEQAg3s2fPb2f1lT0FAVM9N1lxjE/evAzWahVEmgxn1YNzZsscMGd41YFASUQB2Y1EW8/vwGq
lks28o3txWEP6gkB6cAkWIPuuQacm9T3bA+maNbYbTwfnj6aUu8QvkM3oFJBPcwRpAGs+dJDHNi/
g8OSVn7a5wbGG2mhb0Yq9JOc05IP+Uk1wxhc1WxErJs6NZ1KHrXpN1g7JvUCXjS0ZKzAhbRgzBDA
eqGeGdMmtoLL46hbMktKtWwKkc3jcEoSOD0asNrfWN4BtjQ2GT7R8osdRn6VRZ47NpidZbOfdJFp
37UWYqN7pnLqEPvYHJgkwjX80paNHLicp9uzskZYzFZckv9mmDYwsROa/P4FObZsQc4RFplhbEXi
2r8ONFpOylP5fqT6fH3L3QxWSixZhJng3qZ49mhnIuHlXPuceEaLueThMsAqvYNbUXj5/WJI95+p
SwGrVR0/lRUZVn+2IUFhZ+utS/YbjF7BEhidOHi1r2wLsiM+DzrZrm9oMy6+wZrCB5CG0P8o0LN3
PryhUmF782BWoypqUUq6qs9hf4Nt4IvdO9e5jpnRztrKEOTTdyM6mb768lB9v2PuMQRbvMePYi6k
C9O1ibF/WCiRngh/tSlzY5K9PPMWEOyYO1yPaCPxDUREFoZVMV6y9lwk0HU5dNcO3oasah5dUJLf
M9tHPmVJFZQiFRf8OP9n8Su+mv6RNqjLBzcKy95uQ7n1g+scvFQqp11CoBVHgo1ACzoz1JObePkY
H7wSMZr3/e6fwxfduU8M0Zorddu2OnKVnnqhI7TYake5pKamE/rODCuGtRmu/9cmlaHEJpx8MjN/
DgfJRlrbZiUYbsFiRtvGf92juGqgNmiw9iN/NXD2Yi6KOa9t1oaSizRaz2S4/K6Xdza2mPNtUJL6
VMqaSxa0DL25Lj868GKWx0oeBliuS5veMXCYhjhIDZJlhVYBN3C2BJbl00ScT/VXHv+FFfeikPFj
v9jrjSnzlIG/QnTJdGPRgMcSRM3ovMuQwn6AWgywqJwoxt25GqpPS6ok0J7ZISELVAh/eic51zCm
m7sW99Cqlo62ck1PbCmmULcrCa1Katc6MM0GLKG6bMBb5IJPhKwrBEx2w3d5k2njsdNY0bYMj5Ei
IopRUxDW0rkHphoPRVkBzbrq0uKK3ePej7HFVnYQRwPs/Lnym1lmCFK4aKzucAHtJsU9vhjmISRe
vI4roG3HWdpfPm0G6qEmZVJPEcF8EjbvowdkiDs6lHqTGSyoZrwTX35TQpoGuyOlrrsFK34GAZhX
nxehQyYwJnZrlV/yF8p3mQ2SK5TzYCrG16rg5wVjM1PiLcHtHaMphTxEGUxEGqb1N1OAnTaRoMz4
A+AZ4pDEynpx/DFmhFPVx1xyIJSosSlEKHLX3U7FhY4LAtLceBTqhOyn8bBNGiA0Ha0ZZ5Tkq/Db
6qZvbd+NO3Dyt6iqqGsvCUvmQEfpHeH7fIWZiuV5sLQOVjlXukyv60QQ8n6qya4QSL2HM/837GbV
0dLO2wzGQfsgZfLCdqRcnrPZoYoGezW42d/PO1EkVnRWdB1i3xVfTXkkFfoMx+cv6uzC5TJnyiP7
CQEJLaU+j9q25en8KPK3D3flPgWSJg4MPTpTsusvRWR39YQwBoV3DmmeogOEBCzfpL2kWbQJKsCH
S6d8iv/VQ4ThuEN0T7dc0yHRx+puSitYVPfFSkWT0FXFKvJGiUfN323ml66dxuoh8tIhNrVdIPFI
xwyWTzafJ9RitG4xIndVZdGL6BPpUOKIaWgREVap0DVLjpTqYH+WdT1l6iP9Bwpy0KxHmhO3K3wv
g/+Bty4xcUvF4+hJrHnNZa8hEO+Or3mO1h8P1mkTLrWL2wm7xhRQmzwG1k7nEb2WiXBPVdPzeyiA
7WMQrIn970jr0HHebbYu+OtVazL+eOiZC4MKw44fPBWrQcn+zx7EV7aCwKcbTaqEUuMba1thEAoF
0nJjHgB5RLdlkV0BW88Uu398oQjNFU27F2HLRrkrqIIoGDGnqLIS9lhdMJx1XgyX3zKYuf4MaFih
18AnEWSQnNsa+F2O20jL17Umv3nwy+E260eR37GhsCd05ijIZBA2TpVVfQchEaaGpJUTXcamnPrl
eFKRKvM16RCsQZFuAEeUFLR0qo0Vw44Ay1HjgAHdzT/9WdU7oryz0wtMOQ15hM8P4SManzCRLb9E
3jrk6pT8zYlFIhLE3bkfS9fyEfRPmI2FVfBI+16Xp06+3oSgDtxXVTDr/uX+oCtHjf20ncvRVtpc
ZxHsnXShSHyvPSL8gUmh5oX5Dq1xZaJtSZ4EVG16TAqtP10UaCpbdteViiyawfsyeTrRQo7BUD+y
ydB7tqLa2NBHNmjwji18uCGyicz3rwi3/pqZzIgA/tD354voUcLicR0qI3nTD9YPVACI5ZFD0Rb9
8jfl8Vv1KwbnGo+zzhHDVyNzXaozui+0dNY0/tTuSzLhBunYs3FOyfyiU0T0azblOobWzyc3Yp9R
d/N/hlzrCJChb72T1ExwABvSv/t2mz0rfBDuQPK3F+in3xf9BSxRlklKSotojMRdfkPx9TL5yz+t
eMs9m8WyHZ1cM0uBeXucBV1RM6mbHmyAD0Vvq2WeqtM9nWpRjBlC2Qj0a2GNHgTpDsqh1VgF77U0
k7HhUI6BOwyVU0aIZxGfxUwxuFi95SX81Mopd21rviaAETwrpZWPekN9owkVGKLSFNxhDZfj7ses
nivw+fxvYnHO6ze/3VGbNrsQFL6VEhXcXbrBcShJOKQ3IMoUti6HLoyIp9l3JfDySxIwiEd4sWSg
5PdMvyxjvF/WDZnEEYeiRZbjWIq3oTSnew+LcUsnSsLXidga5OUidwNV8dT3msLNwaU4lFAZUDZP
9rPE7h5jNDO/qc9dVk51q8yek00d9VnOH4ySXZH+BS1FSq3Yw4f1huBbiVt4HlMApGtq9S8zYDm7
iTwjt9GQFieiCK7+fkyML1xP8nKnEblNYmSUIeLhLdFsC2/hOUsyDH/x7m3g8m2RypC6o03hpm81
br6434eNBWy9FCoQ7FI5g9OnjG7Hq/ETLz7Utk/wDpLfVYfxKV/BotKbA3wtmXssercBSAmN+zTB
qeQ7NSGuz1HSu0kkL7LKTR0VC3PeIIsttUiBxfY6CBCqEotSLVrFhb0GlMbFR4S4DqGF6OmuNJSX
B0qrCuFf8rYxLoylaZ4YQEDcdEktEoALiWc53ZnzbWc66VHjY2G5F4EWs5PegBqXcmXB2CvdsUJD
0ZyArgb1ZqBbZkIs2Dv15xmNjkPnRqOgwo8WOwUB+iKJTIlkNySWrRqilbaI1UiHMZWJ+45L0GWi
KIh2FhL7yn/onqAU23Whes8rDwkXehWc8VQeeWW2luEZg34HilLe3jt8ZjhOo2V/7M+QVFlpwEV9
sd+u67cQfkl/0U/TW0qBZSad24yHDCdrLs5oYMekArt6Sm1BPAVrdkJi/qKsrTELSLDb1XbvWr7l
atutAdDE78rnU7WZRmHPPo6jAqaik/yqswfVZAondaZLMyzY31l+TMIhh8aoi1PdwqGAQj5BBm+H
67fSBXGPbfWNp+wN626o2MpWKSzOsmucWDELN4wIub9VD5B6REmlArueETSQl+KfNBxJgfCQxT6i
4hB7w9mL+mKW9B6dAGPM4Uzh9vFAEjMJZZ0VWBQGo2EA6+NHaxRxWp53dFhywe1GosSEWYzePvns
z1fuClycHVpBq3CsYEM/iWwpZjUaRDuyS3IilHH/tNG26loKdRkDjrZkV4zr6uM5P43aWX2ZascJ
pCOIP3iYQDMn2moe3E9ucSj05S/UnwsQWgpZIIB51ogd9hwv7koubxU09fvYRtQu+Otj+w2eV/OH
/iw4l+gICUcE6TAribQASJG62qg1Yi1tpARRFPp9ckLKVwL25iKh5dG4456FobwFRT8wdjrRIBPi
klz7O6/0h+9s2be+L+tla4ttEalotSkAAdF885dLmOe45Abi/BQkWmFNluZ+XptOGtAnb+L40GIz
DoXaVSJSlmgRMmUINsCFqkx382J2kDBYDJGu5JWkZxf9bxY8ARLppu7kvA4LiH/9i8gS+xQep4uI
jiJwmJdImDXRX7AHtvssNb+4MSPCXc00zG3omo2DDnIKl4MqwgMBHhfMBa8tmeQd9P6MTHVDN3cC
B+MT5O10IDscnq2Gmdlc6wwiUNqaD/w48Ii4XUlrCiQW/8La7IqzfFVFCAOSI6LVXkoadUUAHYQT
y/7CGKsWR+sLx2PpE25pvTr+nqWe6NqqCoIFX5foeEO7vKkU8OmjWQWf4B1doLG00EVopSoQoJI/
vGuB/Y4kx2ofa29RHvOFsiWiViZlPZHjTzzWgVInroqAaRzYEcL7GfhFUiripzwq85x0IXeoDTAd
LzgI4hCXpnVSh3hibReSIeqhxUmqN3HtecgNh9EYd1bo0PNIyqPC2G8p3toySwIXSnJALRmc4fe6
ql9q8Vs1zBntf0A7XP6Jw0S3LlB6thoIx9sWF/g/Kqgk9lTLRcURHfS73M64rmp2h3LbXmKznpKi
O17P1h1O5d6vK96f2nc0jvbIKKbMEchSTDoAXD3mONUqF6Y14z08q26IBs/JOv+AfJGGZYcl1Ej1
4nuujDA9ahMN5gmLFBGY08X1gnE/47UxIYRY5xyKeG8ZkqKs1zW4+oqVTrMQ1Wwu2lv+05T5pxBd
BKvTwcjjz5Y0q331fS+t0KRpuiC2ESrHtjhkRcenrPMZX3Pt/1LLc//S8votlqvn3J9bz9iaFVON
gPZ3eeKnNOlDDLiRcGKTbe87F4ldTGFUBBoAfyWd2tPGhVBRmT5D9Mpra5mJSVU3fh8UF8EsIddk
nj8raYY8BE9InEhzXqxwvioUk8NASFqMisguF1MO2l9JZqiOdNZVY/4UsR66hkwuyc3zIKZsT+RE
9IY264xrcY+vVjgRjvdOW4q/OqSCEsRfjvxMTmEpUdI34at5myhUZ6X27TQD7/qeQf5OQKnKARSc
IplITLM+8bbSAtnpcVYgc/T1qadyh0YL6o9oVRwGJe81F6GjhPHe2YBeqprJBeJerXtMu2WmN11N
o+OskEYVrHMNxGlnhVn0DZjKODCPkL1xuVx9nYWlLhAX293171shvY8rkZ7ckqL/4i7HaBCrEQyW
usD/eKSOHFFBEsb7jQ6n0Fod/CnK2ReUNdWLe2cCa8ChatuFxoIg2YXIOUu3eErIscaUtcz8aFrJ
l8srnTqFWjklMNTm/UP+sq9XXaLyFBvll7Bzvw4dmtUxuaa0UyZt66OXt3MgtfMLnWH7e/9oVAyB
bjlU78fVknBrmyn5ZHzLj2mjMPtdMTo6X0HVznvQcbMvFkbWvPZlpIXM8gQDiCuUp1TrqBrN7ous
eHUxIb4WGlU6CjkvZeYWd8pvJCHh8cMOHOYTfs9Yxh5t1bBbaSieY22FrZnrLcrc1G2yTCfNDFIs
yvzUV1upBDzX26lykWf5uALZJ+9A8iWt5OCGieuTCNS1bgwX2k/4YcqxNj4uc/+fmkvOM/v1q+sh
8/WzjcdhkY3t9BWLj5gbtBp1mFjRdtc+IuKVo+aACelCX/T1dKJR4kZapuizNHNMbNIiS36Qw8NL
M/TdIMWHvy7znkcxYlJNmT9Tj4Yfu+UEExxg5pSOc1zeh4HqHtuVZy7vEYS8PyyHeDHgFh0VloBG
gkXhFoSxUp/YBSVwCXFDzWx7Pj0vVsftgUVKS8xX8ZNW3+0IA/sbS0eBZXH9OPPuvkH4G4H+NHqM
bKFsxlcDKNgk3OvKVbq/kUmx08Gb6hfZNys8rkW06Crsqy0/wIezOyBbinny0uCw5gy/8psELsRa
n+aRgDsIkcEdgo09+44J9DCqtzHOK4Q95aIHcjFpCzWcvRgj7vlafWaksQHy++0kLP5sFYX1TgfS
mRyGDIUOpIcL3tyuEuq3Cbtf8hVE4AZXF4rri1RXDec3+UzCYyjnGZnU91V3Z/H30wsUTbZm/tvs
9hYuJf8dkwyVGlvaVC50jsy3nTdxDHw3/OrWjWwmTUK6IY1v0w0Z0XgtwZzojBzQ4UTekqJxgfOK
jgstsAUalPUq7JTBp+sUSIDYRYwNPuUztWKAZvLnX8EenCu8lZpVuKubVcAFfBEhxkG3AmQBHF89
SdxT5B9p4CLRBzXMwsfgsJfDYsfA/oS2Juc2fBQtPy24DLcJoH31hwjj+9v7KQZScxe41eI/iLtJ
WMQ83YwX0kRlLEExKtm3+1Xgqx0PChtuzDVPPMPPqyNP4X+ZGVBrDI+GeCnZXzDXRGyQrsTFS6yT
cKTsPz+feL6EkHjMd7f+hb4Jd8fCyHQkThJQzs4QE1VHUTnkJtXCeh2HBi/2s/i48RxIIs+uf17Z
bmewcEr1qoETTdbzAhlTENQHFHcKWlMcmN6kxMeIGOFxGHxyn99ZotJPKePtQOgwVdZ9aYy41bNy
qZgXLTtR8WVhW8hrDDcWCPIpdmgkklyaNEJ4nr+ybr9vqixR1G/S74EvLzfLhUP4BkibN6zaP28e
cDoLnUo+NVxZmx3jsBQjsgLRq4IIEuGK2Giil3Vgz37/1WpnKpak+elU7AdTXureZO1Ahl04v2Zs
SmvrRoLML+dJldGoj+3XGuamg0HO7PRWIBL3Ph09ykpaft3UIwQKG5dD3kljyljlk3nT7KfowqsM
cgJ2OGaClp4ZpG0ItF7i1cnO/LybUxfATSqEGYSPzjbVGoV7WN6EIZeg/OUILWGwNpySKTQuQt4u
fPv2oVq//dWVOwlnaSJ/VuHOeOCFBQChVu1b60+JIDmezRVrF4WPfBfVejUL97kKcsCDHXYoFku0
c9GKkC99OISD3OS2bDiMBkEVssWYz5SCkCgCtl2x9YjxOQI+mQs66cESnzB8p7uGbJQOS6kK03J/
320anmNNQgRJ9IGN6vIH5kovWZUjFPpkyqF/RHjp2HAspdNP5jd2YnOLNEbKLHfaeIW1ZLccn6lR
0/xfCYd7wJUIyqMxjcEGy+U7qb74Aovz2ONY9B71UbLcfaqWtim+4j+KCIKphXjQq1b6Lla7IkNE
zuABf/tp56jzwGrtpZaz0I1KWzGg3NR4afE9Nykr+dqGP1b3b2SzERn7E9OZRzAhSjOooyHBDGIX
bLZFJg05hHwqHxEIIjyv1XxTF7RWLpi0aWwyB02Hq5bZQe5y0mYPILDZwzupUnaEQtJfoxyaNNuU
6jU0ATZuP15wYAUgic2TjDdTlK3EibSURR5nVuMAfsaoRMJLsYN85hALAorSGeS7hE1zugOFm6Nl
Pre2gUwH4NK+NM8oifHClK0EqaefUuKR539o0TkHtImRGORvAH+2GJM77wQty+bg6JVvXK3ZIdl1
DiTIo7bzdTM2Et9eqbBNBEvkE+j+hO5mSMUEYibucpYo9/bByxcfZnmkG+3/q052W5GP587ff5x2
ONMy8igbIIFaBDwiMVvLElZnptN1viepqeCp9AaWH7wENbGgR1G/POhrWos6uJlaNN5THqaRARFQ
7gKZb8puJgJ4Z4F1LFibfx0EKbze3u2ZDWkxPRs09c07boZBcCwd+zY6UDktwanwtdhwbONZroSO
H9h6qnuEfZVwKH04aXj/cWXreWafnvyMFe5NLKFkJhzfzG/FA76UXPNooYpBQ3//dQWKJxFfY0OG
deQBxnZw/ZmgQpMov6vvidiJq1AyaupFnox7EqGQsebByM4rMmhgqoQqZ3KaszrsJUUwIq+vECNk
gmY9Xeecu5eQoOhR5huxt5lvrUYmy3TQWyg5lUhwD/s5J9K77l12bpItga3g5WQ8zD9cEbMz3Sh5
Ic14KQEpfuI6N1Q6bbrvn9lNSuAXbldyw6ymhryNlwBVm7st170O6GImwNbmmgGewfUrLc1EVgcE
FqX26cX2auGDhgtytItEaK9e+DjM/Af0xDdOtJJHITTgzLXGL7+4apC/rvqcdYwvxeK7lDBtznkx
rno09QB+UktL1zUsGJV+DMrhliM9n+UnYBRgDuQTurmLJi9dfrcsdsR3Nimu2szL5KksVpzDxgy+
KcJ2lVEfxZN2wdhEijUynBkzV6jKa4xFTvq1HGBO7hi+Cz1Q2Jou3P/OMMrErqleru/Rqk5JJMWe
zied4xWW+cnmMf++XM2NqhKNOUyZaZ6toknCOvtFnbnRwgpHuC5+x6zD4OSv1fJlZFTk69BFzCKl
zJwSGk8q/c27pXmE9vX4ragKA5qhzDK0sIWqMvgXyq/adV6Ba9egku4SyxvP9Hx7VMCKaBaPbKNB
v7b4Kjcg4pB+I8Ad38i/3TT5yC7L4MopAKUwhg0QpwpXCrIhCZ6DLkxrGvYCZQk1SbUdemrk+W1L
kLiRFd6I1HBRRn6RT23MsrPIMAJIuvMeI4ez1VVIWxqZTdWHh/ftqxBbsFY5dldiI2nDJZ+mv6E1
62cWVQu5QhJADKu1ZwoH6NA8xMVuFtpnfqYMpgH0J0XbAn3JvFkdPtC4xep+0PYd7TzpblLlfYXN
AdXpuc9AaNFGaGHwvcRsUF71YAT3KyuTiVvFD9SEAysXf5e0nb48FT9CrPdfPnypWtvxBhelTzf1
vUEIUybK/5pxdQ+WIVpaLk/igAFyu6Nb5kFyAWHS3LbubJ17ww/YmghyBllBdnKO8BY4c4IU6INt
kkdSDIMhucFjueZkzQzsx6PAbV267kFooS+xXo8ylpFRxx7Y0yCtZp6J1biRr7+BCIETcs4gYbMp
b26s4+PLRzL80srEBu/CE+MnI7rJ5WExYgGAIb9evZMPpPSzdTxwPSWouqS7iGgRuuwin/bK9DYD
6tIweYwZZ4OK330fg1aMoYKfnLDblEnffwqvr3JYRkuiGZHvOmJ+EXwTHyS4RrWGnBlTDDyK1/9R
XnYIj7jjp0jqDM9iWxn6zAwqnVq2w1TMgPSPfvxODLpE+91g0NMZ5dlh38b/vGWBo3tDMxIx+lRM
9eTdOBONIknt9aEeeLrt3VX8UABe4BwXE/AWj1FXUhGFVLZ7GH3lhDn0R6nMB+YSO/y3HdplPchG
ytO9mGvr9EEVRQnnj629jLm5yuv3tWtIGB7M+h4oPgJBefPVQvMwoqnw+WklnVhCz13JcahFB9l3
fHQcC40epHgLHoBs+FuKBYRIf4WO6+56QubF5ZE6iPaOwJ1Yojiiiz38f7Eyw7azXKmmKkMXe5Dx
MvUxhxHuYkGvl64ePWwyQRfScB9Iz7K9/tLEYZ2Ifsl5y4z21CZn7Z++wT1kGjW/Oe2Iqz39jpNu
T21s85ebkRAbr894WrhBvZnu4U8k1ku9Jr5G2MWLqTNNyxo27x+2PhgTfDZPc9thkpFQ1EeaGqXA
klw6HV3F4orTlX5L/J2XrGosuE81P3150JlZjGu/XTjBvdj/4Vj8QZKVvX5Uq+AgIVIn6/8R4Yji
CVSGzZWylZoXZmMULDEZsUwPAyAIQ3Q/6oN5l51oS88LkAQsPJq5NYm8Cv7Wsy4gtFYlqqJeT3Cm
fc/C1S7ON66xnaDJ5sLlTgDKZlr7tm3ok83he1AqSZODos4Sf4Oy4dlEWCsM/mHUtUnzEPzej8WE
QFHKdVPQQ0FdACoAxWLPMCYOR332McH8OcYqLDStnhzmoox40wW+7pkQ+NNfnK3aAtgKKZY5v/oA
CYJnoyrJlQEaCHCePud30nL9DpGgkoc7ArnaQJVxx5JtQqdiU/P2T86bQyfFZa5Jk6warJ8vyD2d
FtxbyTyZXErVT4+crkmCuMmGk4MB4ZxcYSPF2aADQlCrpFvqrYHQD8Mf4AhDFWh1jkaBDM4Snxwk
s6fPLLeELe2sKzKE/dGxHfaJAq9e4QYi7MrTkVICspXY2cOn/OkFHHoG1A+ieJgJQ3hG3oumkoiZ
iJlBui8l1FBO5NcEMjf5K6IaWqHxBAc5Pubbd8mbS2GrBeiSF2Dy/5bOaWl8G9NQ7+exX/PHdUJk
9gXl3Zs0sLdtXeKTiFuwJNEnxWxeaj4gfOTENMvFixQ46ejjpFYnW1zEnGmabXmkK8j3cFwoA23Y
O+7FdSKUnKA83L4MfMXuJzXF1TC1QhouvGjoiy6jX8O/B73F5vuUbKuMLQCpAUAYAV4WtzzpDzEY
v5QsgCIUqNekLV95Ir+u+7KMFEsRvGTpT/aeHSb/ZzO/DnoSjrsd/bWGahrUoGlwdByY8l5C9Rf4
5YHTmLjpaMDkUe8O/Cv5oTdJKO/aKKTfCVDGB7WxbEHKR0NpVi3kLWfWtQN6MR1u8cna/GsSl/P1
02h+dtkC2hhK85Ngu1r0WzYixFEhLZeqRL/XRbfbIW4G43dPRTVjs9Ja/C4krD0izgY1SnIkEwUV
1Rh6EqcmglwoVFJflBpMo/HtDR8qRpkWOMsjwPXGHK/Em5pT5n0Vj5wY+juETsXND8EQsb2tloLD
s9tod3MsVgn6oHizaDcL9Lat5yMKx8KxUq4nnlIsN0qOOhLUPmKyJ9TnKkUxYJ5GjSy0Ty0mPXQz
oIn/iUIrIgxfQOca70XpZyquAWcTS0YmDCbxAIeWkdYLQfeSddMHCetr2JNXN9cBprHLkZ87WwSX
p4lP/9PbVTPzjr9GFyZCfiKO2uwBkesdb+0y9g9yfW7xa/dU5pSXh6sHkKYGbkH7QKGS1w0DvWd8
Zp+QmuVlWtco7QjvtiJdm8hs8zOJA0VZNvhxHzSQf8xOsoOKEMnmSn/ojKDZtEOEB8tqgyJuOVDQ
U5vrXLn7TkMyaid5m59XSRIKgC7mg0NomQiHLo8ZrUy7zhibU93syGK9nzC9iYCZA7onyOVOqkDm
CjdJlTyCc8p51JkBNG7yVzNFj0HToif/jjO9XFlKbDIWlt4sCeNst4hd/7COgp0AJ+xeToVr2UjM
DG1rihV0AS9Px0Rk6+nSimqa2n/aKj7Vgf1pY6N32kj05j67eTbnuVCJE/Uyq5XQ9r70w3e2EYoH
begPU5EVk7EarhTNoU6uXR+V/xdwF7zc1W09QJSngBth6e52Y8rXlHYVO8iXFyGjb23Ml7loLqTZ
J4bHxk5hY0Shh9/4ZA+sst5+insrJN78qFEgJCsF8SM33u9PdQa4bbAKRmGB27tPkW9wM3Env9v3
gQzzVDGHH1eb4+uvyxiMBg9jUErzpLN0pqAB05WHIcl5lIoqikeBdXqISEvgfijTxakb7WUmWuEX
5oI/owplogdIu+rBPd70KpXArvUxXT2g1n1fDW4NNwNxGKYPZaHccTqO/swG+rw58CDjYQDWHot1
OpavHJDaGUfkoSBDi3NTR3WRFLMF296ixu7rDs3sayk2ivVF59iWFnGYkEUKarQBQlY0O9VlLHkZ
ZECXO6Qo+nvOpjE4JOYbLHiurBS3nX5CEE1XtIxHV1E6yKC0rNJO8LjlNmYDvjfBNlfSyprqFrDN
UJn3YfwR6h+capKeIvFPbrcY9LKKOTIL3q5c87USTqNqBc1MSWCRjZqefDdMrc5bDgq93whr9ON0
Vo3RmrIWgDyn0xw2ltkhv79xUV1KlOwqVKXYDmQzgB75TONuV41RxzcPKOFMyaI//JuF0XMTt414
XLKDgPPiTo4iCQQt1EITdV8q5AkZHIFdsVjbvTcb3PPozte8hV6gcZuulo461TE7HL79VThuBexb
xycLu/2skufZAtKi0MAnRAn3e+JQ7XejZoS1rY1umf1ldOHjayyg/GM3hTeDMIpWXMHcW0dhMAZB
3QtRqQwiREGq5OjrF0rL3pM6Dy6LKod6Oy9+gFmKdZ8csbRNDI8sSEZ4r1JU0M+lsVFG5Y6+4/tC
6oQWB8ArU1Xue3ZhQWvRDfyGvHRRFRp3ShCqVzxzeqcLwhXqyyr1HtYX1M9OAjqRHJQIcLltmOh0
fB5MR1hVHfWs6CQgtloa+CPbZ4yu0TYwT+FzBl+waw9cSv1w4sj8wpiB4vgcyhmb1dSqW3v+BtNw
YnloRhmPK3FjqcL0gl44hmep4YFuHpRhqgMhuuQvyB3rcjvO/GM+tnoP9FMIKS4AYcrGuvIjN3bX
F3r+j+B83FCKrJDUlHUHNrEAAd6m0WnMo9rlRxKPKPI2qSKOEOiKjYN3L839DEupfxN/vcxGE2kX
FsU2zgx3pJQDJ/r6f54djV7vxztZiRjMbX9xDH6ofiOxWI3UDRvRPeXBRGOD/3YddL0Tw8JyrvRt
ynjqHvE6y24+F/ZPyr6dWdqMn3gqmQq8jHyUPuQTOOlX6xaElJqzZAG0uAc721d/g3FucHYl6BZ9
X7SeVrsMA05d7zkKttaHANYy9xd+ajPEkbPfIgtpG+zobQkGswmzFh0tG0Grpk+X3ntVXqUlCnOL
o2JrOdws8y/uba6ebzEsDHmfkgB6D2mK+PWAjEk4r3lpqpxFvVhVNvkeMrsnBkgMJ5sfer/jO/bx
BqVZSEPvogunfNQuXc6HP436xUziHF8kefb7HGHAR2Xgidv4QD/hCoMPjLHoB1NEWWwE9ioV/Y5Z
zP+FAH0iwcgueAePzH9eEwlg2Lf8/sq+uBIivAAkYZaiY3lPj4nHMBsN7hJcferlFrBoaiyjyIhL
RPIJFmD6rBR5V1mOnKDHISazPg/0lBVUILRO+DqZ/IXxHgmcG4S3SDf5oFZDBIXPgVTEilzT0q8A
sjaaBV1mbfKQQlRpC98PxL5VB1EOMnpTnceKHJGhbobOHalPUOObyhmBaIIfAvC7Zy7P+hLaAtDU
l50WfNgG+QKkEVShYUySFtK5PSiDHjSEqvkyrz33sg9MIKMyco+vKu7AiTonC+xsqChO/6/x1kc4
MsI+cwsxb+OAwEeBRJkCkXubmfOhJaKIqdMOs6mBKW4zMw7T5Uh1W3W2g10RjGAJbIYYmUAlEkQ+
6StuSLjlGtlSRWhB0oIsuyQPMdFJxd83jL+eoXH0FaNI9Co+C7pVu6Kzf8sVZqkE9RYsCRjFzwA8
qvHm2WzRjUPLl97WDQc8VFaWt2J4Ee7FI/7g5WvNOMOHIMzy0ygdzKe5vtosnAyXLST9A8DUnVfX
rzZaDAukJmAIazW6x7dV8F6QISVUc0a6bgceAXJZN8ufGSYt9ZRbzzMg+mxjZ8YIrAfxnwQZThDq
UUQ2ZH4+Wdwdm4IluNp16VjUurFTIIyevh/oBx1zUt4JD5glnRU1OGkg+Wt64DMDzkbh+877vwe4
z6fn/v2K0HKB5/SYfsN85Nkxf34LOOvd3EVwOUxtz/wU/fho/4CNPM99MOEMH3Qqgx96OOBElye7
35qHH2k92YBLA4KitzrNMYvglQcp9p7wCd+ydm1cx0Nk1LUSSIABhThOYVl2QivABWohGKQu2D7P
dSdcLYtoGvgmI//vGTHjgRo8rcduBp7xr0mQYtblt1zWh+iigRCRJCGqj/9gF2dKSOeJHLIfTQjK
qFtp0F3ZGItnSNrKzoMSwsqdOwwcZp/KN+8+D7ZQCeHxib4hztLM9DPikDkeBxqFs/+31JctE5P4
NFn14k84MxVuGMdGOq4RTwZd/+D3lCt+rewLAxknl2PiJTRNAu9x+vzUpP6r8wshM+xEDvsKGGoc
CohI/XxdOadP1Uc0FUXqW/lU5cr1rvzikTErjz7MxGaLY6hzqTFxf2VhXzvfkgOBznvVLnKgbO/H
HJlrKgtDR6FSQgKi0qXJsogdhRH0fIVXT5sYUnhAAM5cZjTfpoV9JWX3j7xGRHvv4GwNtSW1lUjD
p0UDS1LzEQkPmOfGy30rQtt2AS3k4OACuQGcdWWpNWCa4Yv+8n9IqdK9QY/yw0F/q0ruN/0FtdUE
0IcxBsEZ2yTMK7bZQXFMsWnWHy9l5TX6evOwSmVSVRf1NELU0xzsFPaHKNLyU1d+isEljRjlmglN
N3z3zMVZMoO4q6WfRiQpNZfsrBAkhYI40XLhD6LyXmVGLCrsWj1n5rS88ie1rhwwhPnBN30sZTLu
z1khBUBpli3Myify4TXV8PaUisWvjqN3tHyr5J0KL4ifrgNtLQZCNEcCp7t22diu5wY9qzBjdXxc
82GCiI9WaOxIXtNC4QAPfqRWim3zPHLb8EIpA+LkNHqKaK2W7YMZkvIpWb2OlPfyy3GG8FMmuF0J
J/yKo0e8Wn7vGwGVYWamvE33zZatPP3Cwi8T+/+jKoS7y9t2i/8or6rNaxrmZOP/lFVHU6xekyqD
FQNk4YdMLBxpyP2YtPcFcYh7NRBO4GgBFjJe1lWLfAUmkvpV/OPVh4Rq6i7mjP09v9MPhqRgGVBc
HVnNVOjGB1SVgrNm7kxrZ/hh6+QFCDWFLRP/Hv+ESvnS5SpHqacpBX6mgyXl5dMaFzuUpBDY/B0N
ZS76/PKFoMf5v4oganbjyuuZmj/BCVpbTVi+fOfFIbG+917Mt8fi0WyRUzIHmA0PxHSkR2VMaOXE
lgh3BJvd1CMKk2KpP8IgocSP3B6a9FW5VQkLSzjbAu6Xbz5x+ub81V3NRq87tKMe7ZfVOdapxen+
l1aeR0wCSscAtAnJPL3IE44dw2wsOPVIpQ8j8ydOA4lBmMaIGK2Vy0FxiPQWtevMPsMuA+Wf0qaX
pBmDtyyqG60VsA3FN8iMaca05T2jMZkZO8UNeSaLbjt+G2HlS/+UWTYFDTBTujdl6fS3ovoWDIN7
Yqt1dkz1t7iNqbpTWeqxoh5K9JhZZrYTVyAAdZ9XzWwPd6PnRO0EjbiwGDmwf7xRA0gJdqFDjYdE
qg7mD7cFWc8bqVl88u4N/b4iAn5ZMzCPq/ZcOgCO5ojdszDhSEiwEl4kIdJoPf1VPMlGwLu4Fr77
IRjhb+PWrjmwJc5at0uLvzXoDrwWGOnghIBSaE8sZ33dHao+aBoKsT3sqBujZuy/9lYAmqpY0c+z
hR2MvOc5MZNQNfMwn7ERcSBaILScZiCsxHJNvxOh2omgD+9QWu9MgYA302zqPvIJM4ejf1hYtdvW
jXNv4zeobS9jPCeDEQ5vOy1A6GadphG6SpEOjBLsJonTnAly40pePN0kK9fVgLUGCzTPZ+FvafI1
rniWmrSOjB4MtUlTyuhK64nQ/b6iPY6EIkDifQDpEjWmnXfWczJDTE6oz6nSuld6om//bXbLoTTT
3snLMFHSrEhJFzXUXVQzMeY6CnuW3HOPzCBo8wcI/5aQoc1RQGsmyAXDrO9pqbOf7/uSSv5diQYT
2NFm0HZHWjQNRo9WXCLH6iiDCii3QHPh9035O+qu7LPMyKRE9gvLXXOob+o2wJzwaJ0UHiWxgMWu
muDyU3sfzcXirYY7ZlJ2+A4af3XvFlxtcKKwhpYo4Z/VbgfFxMP2Z7tg/QAPYFUb8U9jPE3Cbqvg
9J5hrgsWtOw/5IuE9L/wV8XZMDYRYPJT7BPxyhoYeJRqWRtRaI4dCVP6CXX/1vMn3tKEKrBOoZEF
WPkNSDiaZXdTRWTLZIeJ6EwMUVzCNmy1G8YsQENUCYMahtVIRvtAfjLUh0OnlBG9CheDznhfRjrh
hZ+scKlKPz1D8FzoRte52cSa3Fqk+KlAqX5lzzEpZv1xeOvvuDlGC+Hw1sejg3m/3FbLN+dp9OTr
vrYLSLEd+TiZe7rH+CVvqHJBapTpSIWMMNHz1R0juxLJBBHEs2RW9sTEtTQAyzRvyrZ1mnliOuwN
mJsgEpgLGdFddbyrR88/qfK/lJcbHJYJ49FNfWO4TBiXvJ8OM7Qxs6xZk7j8Z2WI2wpagFst5sBg
ng8upbLa8kHh2+yUn1K4224qxq583/gpM0n9zZq/uGVyzAci/hu9wrCA0PQu0v3YLDOVTrBOSb/q
QwQN4osQBGAv5T6YL57E+M2BaAGxEQRXNeq3RFKMzBqg+njeYB09d9dGovvYWoz8fPjjiYzIjQmW
2AfIzaC5RQBAqPAdg/l4AES7ssgPhCzYBV8TMGBJXfA31JalwYawEZ0/5avjSRcohDFy7pRcxoRX
c7xSKQ8hArlnUSt72C6+LXjHNPr0NqJlMa8F73Q5bnZ5FYpxkRF9pi8t0Kx4LmBu/FuJIgcgofB6
K4hsLojeO5AZd1GMMwnk9UhoYhhdN53VpE4ZW6agRc5ejqhgs3NJzKAIzbMRCEpUaw8huefxCvmh
4ft0C4OGHqQrray8NbVaZsv8PG0T5XfdNMfaYdSpjvgtjs85suraLdIOP6eVAnjLGNaI4MiSVJaS
V4x/sC3wyAA2K9dab8ZhLbZEJkjwNgKM3zU19C/gA7vLDCimalYNcdbNn0hyVDCbbZtQ0Nv1X8Df
I+gpTJtDcLqPtMekaMMXhxN9nIVct9k2fQv1KtAu82KDQdespqerss+DmVJ/wAkCqHrGoWp+kNdH
kyrFTZoRQL2Owuxsji5M/tdUBOqFTIZcmdNzLMV2YU/J+Fq4n2HCd7y3zXJuTFGb3jLS/PN2lIjz
FAlHdyrmuDYdFjZpfMlpEaGdXu18+3zJjlE4MU5BNr9MbT8IoyUOOW3kn/bbrIgwSsUH6To7BaOZ
ixJhpTBoVG9+2rLJdoqsKLXmOqJ6CD1x9YuzyWd7M8lBcSLycjxpsVfSZOIh8rDiBHF89tWW5zBh
OTnYSoPZ5WeoFA1joujlghcA1jsCZhMRiSC6C59I1lurzR7iiubh2D7DzMU1rR+7rXTMWSm9caN8
GGbKj5fuzogsyHDTsNVS9FLKkdz9GoL0lq+S11WIWAe1aWWAW1subGcWF5D2BoNrhcQplEdg5Ie3
m2lvlDG88kuzxFv+KY7vCh690r4nkGciHri1KnHUAj5xnFZgKSCipOgDg5H9T4rbLq6OCzYmbj2s
kXIk4NKP293k+MomOLYSn+esIuFlWh5VCk7x3AWRsKXsfUXsjZVh6fOAttZx95aLCB5SdxKJvj7w
FpKIf2GAzOHwS4FafOfDMdPco6bnnVrAubSl+cSCwhyBCh0eJavTCzS1JaUlZTqaz9/j6ENlo5pI
xChIWBHlv9we3D516FSmW+Mb++GqqSvzKCkH/Cfi2Q1K3f16jgy8lWVQUK6IWO4Rv/2+sRryC+YO
0IGUia0u87Kyfdk83ghYI5zSFbK8zN7prpOV4sAH7RMrL0kq9KtE9a0xHBoDN2yXlE0E+UMivOXx
JpSj2alAvtQ2fhBZWf8Ikflw1ti+CQEwdV+OaRIr4Y+qMd5AOwZZztbH20Hex5wc+Xxlk86+U3gG
Zla24FqjPSgEU12vkOtTbWYIKezIJF1crz5e2/IBNI+4OHB168ju/hNKrvOM+zwVwkbcQ6Yk5By3
c7zBu6kQx0y7VhYr8nBPDumzJtCdFWm3VrC6+jMtnW6WUtFRTMTBDxovBdx/9bL3RdBSfb4jRDn2
YgILSgIzVA/ZVDOQqfpUL5CzafmnpHBY72hpye9pzSAR1vwBxwMWf1TKI8oY31wXqa0mCIRk8OI/
r2CCK08Vt+gWZ1bTrzLBTZtpxd0yopie3Kzl0GWLE/9qd/3wdIfKlXC6GE7dv6rlw0KbyJT3gQQZ
8+uhbwUIBZybhQRl6kTtjHuxqcb0jFbSPbcw2KlT3bjbYFv6/x4g76pDamaI0HfTPp30+JAFXc7f
rJMBcRX9uZD9r9bJCrwCRndpAMQlbFbcHO/zX8xYk4s6yLRLR/svxzj2tGVSBmNXI35TFN1YRgxb
a+NI3Z3CcveAfKqRH482+QqhtKh25OijUpA44eMd/S/6Zrp3Q4l2M/fNq7iv7RPOJ2GOAsRvLHew
PpayDTOVWj+lxxqwrORelkIjRl+brX8Kqyb+JXcCsLtqJHgxwFplMiRptPucqL1nzulMTvPtlX+f
MCRsasYKLkpOuRb1WZvUixRcB9fjfiAWroJRiIchcRbaH/THHh9PzbVyQcc5hNyVTFq/OIktt0pH
PjBuBFUVB/hOj8yaDfMi0/YbHPGYNEgkDXQZSSi717r/wzLo+mCLl4PriMlSqXv3BWSs3Rmxxpvb
Fbw0blkqsXMtRF6HhOO7ai9qb12Iu1BsruhpqWH7C2PLE78V48qwIn/VCZaiRi8ZJJKZPEIf4EYA
ZzIpcCeBFgq1HwJR9qHsDbD1zcb7lew+jpzBgDJHeuPk5LmG4fUIqYNSbNy4IB1emcJwQp9Z1w+K
ONdj9GJBFex8mHueZEd2Cx+6OnUmlXAhHc1onjG8UJPu50DapnueTcMSjZbBG2si656HtQMvE3A9
CrsZsjdzD1XZZYBcj5dqAIGBOAgIhSAapy4Zv5xZvTLRDJB1rIo5a6xGy7MVpqmIj1FvPnjE4SoI
DSTlOo9FoQRYMcpBV+jDpd0A0sS2T7Dbsm8uqM7uELt9PYBkuuK/76f9iqqseovdr+5HBLvu3ING
GyWvdYZSd+82qP6kEh+15hKUoetsnAhGyWxcWXZfX6K9gJHlaQO96NrzBTmCm669daUzZ8lM7/dr
kQe7OftRqfM5XYT2a9YlpSLQUyqH24fZFiitv0HWtGOHXV1ntQ/qgc34Ypb4Y/hSuzUCpyHNxspe
rBAELss9+RtAdEFGScJzxIgsUZ2qP5FgGL8fcmtyrE8l1eAxWBf6hLkr3W//QbelOGHb7biCG8hW
OX1B0/p19IyJZk5JHmURnB4P9ERZHTdipqP1CFaKBmOyEdhPWmgm77Q7B5VwnJmj0HQSRiAjZ25r
ywnVztPH4JvXlCKngUDq0/mhk7zID+q5MHWRNS01NbagtRxPxw/ASl/IxkVM6VU44YDRw0wlf0+v
ccgXi+BIDGovR0QSiSWFSWrU8i3OJnbNQpNc8W4yqI0Q/rXCOxn9mF/lK/+iqUZhLcjzwZPzKT5I
LmbNc/UCiwQiILq5eWeapdH3f2JKrvi9/6gfmInUlIOn53KaVy0Ip1iiqvOmGgpGA9KBx/FmkCnU
L1jI4f9dbvRxCXJ6qrmmV3o0iKGRJ8WZsc6MqvcmYD/78Je8zYLIsV4IRN/lHMy+W5p65KBE0QHf
oDx66UWnfjAiDYWOSf4drfOPBanNzV3tTZ9d0icQJwFbqr/Qe2k5Sistn3vRCLllMj68bv+Y1TuL
eBT9bomznnuhn2PlvNSgzQ7VWfRBedH6iRlaKZNr76NANEcb/v7vCVvuVm5hQmZjxLL5/+FlUjTQ
Gmywd4MnI97jXW2LyrtPDQ0Q/CkV5/OqgAQqtqtr1tcXwGMBQd5pAFFpnMuJbXXyaPIDorO643uK
3cZLhtew+5rKtIDLCBBWI+n7Ivqm/w3dx9ux39AOwxX3LewfZk5y4zbd8LxxTd2dpfBf1QaUNweF
6fJ8mEy2Bq7FY7ESYTXQ4o9hgQ0h4Po8w8aUGWdaCdgHj2EKl5SrfBtQ48efLi2V1ZxrW80tt16J
8ZkY8Xd1fv6h4fntjyjuXT1ivg6Reks7x8+TL6X1Ioawf+RSkO7JpjLy83xkJ+ciqrk9tHVyOG7c
sfxHqkf8jdehwH8s2SPXH7kq+qC818fgHYHQ0uryr9VyhG9SrCkQCuzmxZ9PeXsaHV995sy9kB69
tFYoS6a1WMOL807VG6oy8k0v+YxoEowb+gnF/Ao9rAZK0saZHV+psAsxHosqVwkGZINUzTiY3zDX
3kTaNMcPDbNQu7SO3C+/eBa3tMIng3gTFLM96/+JHT5fnnV+iY7e9vUAbFAL/To1C66ich+P2yB2
Pp85jYAuD+wVvpoEaJJAtzDUxNQlcsVDhKfaWE5ggrseEZ31bFL7ne/5rL7EmzHAqUpuFD3I8Sbp
q1/FPrGTLsoblG+dMugoeYc2ySmEqGq1PSD9iLxgbM48fPdyPxd+TJtA7x2MRGvCMrQ2XN+l6qE9
jwxajMrd79jzy7bAUxuZVGMANRMuNCSB8IOt1Tu2lrevNUb01/u9ms+7EGbkPXoAINx2Zw1WQURs
ZgGs6czPgcjCYircrBuWa2m7fE4fq1WnvNb/KHANluvx+wpYQpWGIGoMkdD2xwBTljU2H+WTDQoK
bmtBbjzHxzosGVr83mD4SnJd5SPCpwdCMgFEq66PAvYL9lXUqv/N/E0QEipVXkhm8Obn8UTwKT+L
0AoxcHJyDFcnlYy5vMcNEg2GNNJkSr4ZN9ZmczXIcvZjwzaWIfmdw50uQ5rOSOthG9U8b0uNxetq
hhWMIHi+qzq3P+aF/bYM6vlc/HpY6RZFW05mrop76IEyiA9D8q3cb3CtWf37RcXQPY5CQ01NvWyg
smac6lBXuWECaF7iDzcU0geXWgLuGpSjMU5HY/0kZtCWL0lhdyQLRBDUc7aUDt5AuidDUhSN2tny
MeYSn5BYEujZc7oQKe0KqejGKMyzgfZF8tPLur25BySD8L2QxMmb+2sfaibVvQZjdAvqiaDgh8fp
mNc9p+Sa39eKEht4ky+Om8RmNTXZcPqNVYcs20sL3enSJFLb9tEndk9jMaWlSbCFxIgRZQ09Gr3D
bE7e1q3C258dzZUs59qb65qGKdkgx3YfG/g8M3p6RASDxxPr0osXwJMv8w8H7GLiwhCvh6WSdrmT
Lm4l/C3ttyL926/527NGNVl6TrMGrOX3B1SKp7bcDFC74uOd4wD2STvGjyfmAwaPipFYYG1o9AaI
MO3keYHfn/i4HRjluwSHKMe+SV7NsD8YrKQSwvw7AtjmB2cVNE9mWMkNm1s0iXKVsWwiawsY6GJV
zFdNIpRxkIk5NjehfHiAd3o2DP9h2t6KYcHl3BM=
`protect end_protected
