`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
G25ZkPi+gvmyhQyFUThGoxXQqRHB4tV+E6/CIXeRmhhD3cLpmC/BLtsDJ194GPbF7Kl51EttNsOe
mM3V1fToO9Z9ZGPvFsnHfddDSb+0RNxGkC6UhQo4YPxU5vu/qHFsEsCAOyj30sSaXqAV8S/ZIpNw
3lQxfG4xIz1KD+TAOJijUr/aYEl/4+VgHGRCWWuARioyR96gczbnWmvN3TMrF8ehwcMASJ5d0bcE
E/ikNnoxA2BpElEJNLEjs71PD+QjrS1EeTsnA1HWWhsY84U3Y5X3zWsPS8zzv9GvjAEm4T8VU0qO
CE89X2itSoboSnoCKO+Z5pPu29u7shDNakZrcHbpeInlrH+YFzx5jm0hqmsq50FJ1rIPujNKkn9u
ZcbrpNl3K6lFckxJ5KQrlQKC13KECErIr+B52GWkf4lFBrDZLQHYg9AEuhq2eDYSmswSsogBwAo1
KrF52HzLDqL+H+tSQGnQfhV5xGEZDUU0lpmfMzSQpDHtjI4e7+uuTgjL/kALQiYCaJhoAScurWWW
g0Wkk5XmiId2Wd0rGPUmF1k/a01nf+QKA2GMLXJ+6Gh8dVMpcUL3hrPP0+CB1ve9l7mXbpnT3NYA
l9L7EETewpsRQP5G6WvUv7/V6/rScKymV/lLUCH/ZYCoYwZblbZYS/o2Bavma8TNpovVLkwJF/hI
VowRig5JjTtGj/FrrFAyNc3i6+MTSoK8jDNToxOFYUOBFqgAOQtlohk237FuOvd2GMF9ekEXrm+v
4nRdW3Ii6+o4YK0AdVaKMkmuMWG3uTWqmgpJfxRye6QodLAFOJGtsnkUBn0Z/98S5XF+ewErpprj
SJh2k2H7JI+zghxV2evV1oYVaKreT2jRQNiomhv/fvF48Ukdwl3eFhnfiEBZC3DqG64CJ1Y+isSh
phbYUgqPC9LQMjdeqxhockMRDdAn3lOxIfNRwHSN3e1HmDw/ZyIo7Uz+Bj4CU8MukDiO4Jz+x7qy
NZMdSHn+8PLJXwMjquplvuaSmYHLSwKE2b4bRMwnu48OK2LjzZ+FqJiEyzZTVMTHPwwUWjqYxRws
rF1stsdT9vhSZf7ZMAikaR0h+f/JDHkTck12r1Zx1c9oPUfxUhMg28nbCBpCjf3dMZuh19RDGagq
E8WGV0OTpObRudqj2q/9c3K0S0y/dBYTW56Gf+aMQDb1XuW1vnIaxWrkbEklZd/T81ibNUUX7td3
EJsLIl0cusvXDSAYjjN/xhdWt//1h1XD7Jpq7dQmKf8pn1VY+BQKUPuaFjWIY4lQQG85JFZFw6TP
37osYjszhXomPd6GGu2H3DvDbWZi6Vw7v99zlbRkA18Ut7gg6H0pOCjTHbygB9lZ6NK4GymBOXOL
FPh0lq75DuVOptl1E0wo9hawbuHSnXUyywljpjCx6QGbCXV3RvClGkrKWwDmrOuvUjYKRBio9NGy
dDTR3Fk7HDoBHfwK/y6Oo0mG8dzd6vNkv1UizoxXggSs+CA8+kj5KnnneSC8uN4tLrM53AXV1tFk
rRvGogeb0jF0lIkolq6htdkrH2qV9wbVlZdejI/FSts/3t1i0TxlHFoog1ztbQkHwNGnrApfVhCF
zAf07dYamCTbo1aWS1a+tgJdDEIo8yB6KBO7CPQ4cUMyF8hcpViGU6Y3RZ8mDEy7+hXNatVxb3nX
uTGxbhbxhlgRpffiWzRtedTXmcGhX0CwuU9TgFlhfkvKGWRNNPREk8L8Dfx2WFeZlBXcTq8eXdoS
t/KHKyNqsKIt1kCQjG+0zTfczxcpvElpM2ZF0jlbQDK6kzt0geACD9ruaWMjnnkJ9n2VnxR6awZe
ZkZFlpKwB91dnxGNars5xHQEP1+4W1RWgBhQmupYRHy0CSkVvN32ITx5rAOvtx7CizczqDyZJh6s
VYEmhf/CSjKMaff5s0knwNmXrdnpYNJkikyVY5cs1Z/erLPu+lj8uOTgQxEVFVb2b+N6C1Zb3Mqo
u6TLa7tDTe8WIGUSJkrSU26lB84BcnQhLorPgKGDqTCCy56eCusHsUtsi3Oiu7xFmmh1CLmkeF/Z
26Za+Cuedd55OL8CHrHyd4DRjScg+Pp068Cueyppc1zRjXL9/SDc6OkESv7+b19qZN5GQcKfV1SO
gd+PgsihpEKHNBzO09B6zHd2raRdZyZJk8k+UelQeh6uVwXo2QF4XV/H8s9G9I6qpWrgURlGKP4S
uIxd5qCzUE24TGeoWAkLElvoD5UBMK//YIUS4QbkJHAVtrXTVac/UEMJJ6UiDZlv/HAO3AunLgLP
fvsqFpCvN8nZM5YFcm28WD/9aHh91ytfcTQ87QABmmnL5ov5PthrW8Cv7e+Eow/qAGS795KBOtvA
o3EYwSQiLab7nNthIUDahKpJxF5EgdRSufFGRNuCtNI301bNIp0bF2KSeNAyqSx+if9hr1/gXnRb
LvuN5XlrjFbgHl5wP5zdAWOU+NJ5vcOBIXpIrU2bNHPnmcojVIHGUUwHg9/LUE+Skf+2NNG4Cbtv
B2uRtjfSzpM2nZSuOtnge6xIPLdqAQCjhA0x45o7q1qdoth8V/nFJsDC4LfSrX/b+1fyzMyDfIRG
oRzQ2j/o7/Nl/S/jnPVx5KJLP+07HQQp/Zr/WoiU0Nh6LQg9X4ojoA9O/H0lyssw64H+2qh9btVb
NMctqoPjL3UNsKYUNRSbwmGofTJUz7pXnPTInyFa+X+nP/P3A/sOMU4oe4KChlC4nE9MVSmp2cmM
8hkHXtnEmsBEmxkwqMG6SejPs1YGxE9bBOWGlnSIVksAkQfz66s3ttJSu5f5+yFAoYpCzbCncaGX
UcZVBZMhnbZc2Nnk4xehWWNI6M8ZRQeZzQor4z9YabtVSZ5WhF/8VjTjjyObV7t6Gq3Cm/ctrD5D
nh6FBZFEHRKyk2+SV6zlOfXx8Vld3X0C3YIn8zXIKRzAKCEX4rPRkRGrAhZ7+b9AasWhc0M+MGU6
I9aRq+Nwg8NqWf38rouwa6CQ2Z0QLArSFHEFAx9e9W6Wg9XFdyZ4xrrDgdU5ghVNFDG5pVbrXW0X
sjfpZ8XFH1PAlhmGa2QKtk1aF912EIhs/G0gXc4ZJHbsG3dZJFFFu2au4oW2gwNB+wP5QeFH1u4a
D3Pyj82+QF7g2L3FVyHJXn8yeinV9Upp1OCHle6RAz/AUaHeULrd2+VZPrlgxwEiiRRbPxlHtDUA
gfGl37QN70kzBsSozuLsEi1QoK9L9YQxHXBXilUHFUxst0EL5sIITXR2Cz2t/MWRDv1gmWTVKGHN
foOYC3lD39Dq/zbaNw1CaGAhObMEypD1lezao09TVYcxv9V7023842q6dijYKbN28Mp4TkB39cmA
4hFQW0bj1YA525ffQpPyfXWs8BS7ME4rGalEbtU3iN6LIgbWWLAq8MbNTkh8NCM9ztu7gFuCGBHv
EMUFxficEPMUucBHWBA7773BVW313oMHWAUTjxmkok1zOXCA+NlBjxTMMSTOtoukJXS0FTBavIkf
KpNP2LV8LN16gb2emxzKprBfdM/5CniTbHHFN1YI3O3xJNaiZc/PIauozZQoV9xU7I3h3bBMCrju
bgXZTIxZEQBk5ysDv4/lIlY11DlY9ysNFl7ox+ioka7zn9pwA7xf4ZN9R6hpjv32JYpW+rJOqV0G
i70+WZncO+fGnP0Axj1WHpZAaI3nIvyUv0FoueGMcDYk8xU6ULhs8/bFh+bDpIN10TAeDkN26TNl
YnL6Wr00BxKQq062mrLT+DnOm9ZdjJg+0MhkWkSVs6GjiSzeaH3722MXyRuC1wQzjw0mEwIAW6q5
jmEzBy048tt7ebp7I0s67XxBnKR/vIrfE9iuwnqBeLzUIV+s/ugXjhHar0t6r/m2JXcYPXxLLJhI
P80OcKCmO/yvIJJciE8rlwWILaYa8gK79Kh3df+f41fgKi6aU3je7tk9ANb7fQwnZgC4auBresN1
l8RJPhk9wFZG8FgZJ5JeS+5ICc7dUysLwMA2TdF/RHLAQeFLrmxH/8dNdMLOt9nnnN7zel7MKx3x
9ZGJ7w4/K8b1E/u735X3VM4IrLMOFTfgYuukIsantNWbxY/w6yiw8GoZubLAGzzk99z63BBtnBAt
XxIqD0IcfvjcmOaUofqDr4OOqB6XnMl9M7yoWqt71c+r0RuTwNlfynJ82WkHh35wO9ns3s4WS4Y6
snedGptPWlk4sjtanfe5fv+id/ItK/ekIbpwuT5ck8GkEDfIJhXKNHgPbpKLT7DgVSYAXjlvl1b3
7Uulp/KSS1cPsZUZU1jw1C4BW46H8e5aFkVodzLNfw0OUv4h1mEj1IqFZBm/HWPx2K2Xvk2Tijte
SWhqluqxsbq+oECsWX0zLlFHTbdNdxaZIDYMVJcvW15ENYPGHpfkJnPYaKlcaIXomVCU7d+Z5G41
3c3v9do6CYda1/9pA5rEzY/Qww15AHo9PaR1+1YOs0RAnh1MMcCVWI6iVq0PujNcqR7JIAOSyyOV
SNmN+huIbGotWkfK4T3HRbS/p2NsHWCD8QLz6SHWahydeO1/EQW0sg6YmC5NMYQL3IJMfF3WoGQQ
DEWQB6PGccFJoG7ZwKJAwqxvwYGB2j0Zy37Tilg9A+2oTkIte/xmxYwlomPtK7xER+EeA0WoBgyU
rFrku/W7m8Dw0PqWGRAbCVUAQmWFR7dwOC+SLVgX9jJQMYzR4NNHerI0Zz0drQyXMMPNtqAddnAp
+EM+PQqCqELvoxMb0RwqApoNAOg1hAVNG/TWZXyOX40LynINnwfl4mqcGOL3WVm8BdiKab736l1v
ru44oCbR9tKDB5Lp7hW5wnGdmIMqGcSpdpAh2H1a59CNMErxW9LiDN0NZVxTi9s7EuFOwhlLo49h
yndWnVQsblO394BmF69qxWFn516Niw7CPgYws0MYTctByVAGflq/7CGbkEKYVhAdoNx382Q+vJVW
XhciXfACGxM2gVA0iz2iUSZRIPrfSyd6xa8KzPjsiGjBO2bjmL+uMKQ2mr6wzBR0nbPSLHO2ngvu
XWcDCU/m88QRNp9iAKKTZyYncbvG5UQZdDoyoxia1uFvA2mTKOzgQY10EXytvqT7xN0Pp8FyeHnY
uN28HFh6MxHr4Cw19VXl1GKXkRxWZDpS2GKMs/506d6wAFqIkJhlTHr6zxDkYLgpxAOc08k9ckGo
+HuWpUtQm+O5ZBBy1QUk4c9ScQZO7CDSWLpF9pJCMRl+hRhNpOaQFbbafCg9Ncb1/O5N0SJUQ0q9
gGj1RKCaUJ/IH+Jp1Almb0wrmQedulfI2XjqiS2IPxWmekbtXh3GTFrXyvYCjN6VedOeBS293ehy
04TTtUoBveZlWcVBJDsqPmJBpwHaYS5+Feqf6eIqOXDqJryq7lPnlfoyYgTEP/03c814W6fyyCT3
e0qfH0RTEetVUGaJSwVxQSbVTY5CEJ/l9umFY8Maa/TxtZgdxnVlLij/u74xx41Yr4hcJOp83J2c
trlBw5CgLevLql/JC/BNKhs/RwJMX0rHY28DA6uL7u/pRZ4lIiVhO27GTwvPKIekylPrWHeDTN5N
nTnaghJmx74LyoxiZbDFCQThu85//66vctD5TCLlf7Bx3aLx1I58wUSltwSYOuC4u6q348Y9c1nD
wU0a9lhxf6/XIMMPvzvjxj1WnoxZ7lcOrJKc07fQqjE8J9V5bH9xhRxmVw9pjm22L5525KD+/b68
V7oY5vlCC8wkfceboYR9LGaFtfznHtmsiTGSwKOu4/nqbrkGfSsJpefKoBb7YT3Mrp/KZMXQaJ4f
pmKOEtQl/STvx0NBOV3rDw/iJpsbDfzz8RJqY72kIsaNhVynQH79pS7bzqqzF7pZZy9/BzvCoUzo
77y2Sf/fAkuhWQa8ROowI+wTe3wVCinD/U0S1L7xJVkErrmZhpS6ugvsJwQi/RYuEl/HtfzfhWtr
M2XUfy5ULViaq0YkLVkVVfKJi+So8QIv32oJElPSftxV/Vhcj1k8G+uk2K72yKLzBc8SFppGVVBv
braaqNWHivt4pxYTs3ZY+7GA4fONltZCDa1sh+NLl8Jh5I3MWxLVaDSQ5aD1rubwVAuMtkZ1HpEf
WYAJukWnjwNraO6hVQ7caqJGgIZTKw+w2Jqjjud5zMDOhNjAviRqrFO3Hb0/goNggfiSNeJE6PuV
NoZDCFzorubZFrKNRo/Ddhhdi4aMDNN6mndLIJksltEud07bAe6PW7B53pIuqZx+caI6pxUqcyCv
Tr8Nm42j+Hzqba/OLRVJHmUixBqsDYieAlm1koTbseOSYr8Fgk6jrJSB7t4gMeEmwWjMYRc+rK+i
m9+AXe8SHN9mnUMcDMPmkjKQitwvSksHTCHg6hBSBPluKFUsUoNaN9eKqsaHMvqoHsTF9gO2tLfN
pYL4ik9j5PmMt2v70iSabxdgSf2lhaeY7FSuE+Yv2XxA9sY3xq8TV3Ubo00sXPS9R8b38V9S5ZxR
aXABr9soaOO+uTpUQIedK/ZTOJy7akS+MUNxJHxvb11X6ELJnIL0e8wFpaYlyp6F32tm7Fv2aZ0X
vUwCpWqtuZvBMOscJ1JWJGDpRp5n2vOlhvnOzHsvIJHu9uY3l3bl53GpLs/nj01/5fmEihdOnQep
moYEtvunmo45rBxFVjRe8hFTSoFfHXKXTn08yQaL9IdH1W5y9lTuJ2Uzh8Vqef/NZiUzI+3JTTpH
OPgew1bsiokG9vI6vc9Y3Hsy7KWKMgHkfbuBE8ssp8WH5RNLuNmOiZ9RpGba4ebu5V1kWvAVsAtc
JrBQy1nZa1pj72hbQqOmeJo4M1xT8/o6Xjbr1VJanr9pQnD3wfMc4z8abqOsuQrpdR7efoZ86mYc
JuhnqRp7YPuzQ6FOPnUpNFvZU0WdKjM5eBXu0xGPPoarMFi2Gtg6cORgdJXWQwGfFY4SyP86ASDh
JCcp8bOoGSpt4duZ0S/PXA/P5TOLq9b6Kk21F5lPn8yZ8H63rgMatHR8lEmFfPDbMM4yvuDSSIU4
59ubU6gtYEzFVNVWsTx+RjtOs1hgOKtvqgy+TXI/drfXw9zWUUczFvzz5rs2S3G4qzLTseM06vSp
1gqU84r4ck2FZaEBa+4vQpu0Oq2D9KWKA9gia2LNihsm/gEpJpv6Rq3p+9oLZNQQI0hQPETtaU6E
tqOzYpjJwZlrFJ+WZRKNpluIYostVDXwbISrJ6ZE2E7fuFk2/rc1pntiZK7/zg6l4Swg8Rz0V3oX
svYQygo8plNrhSVb+oshVW67HHd60InuL0DL/VGDw8j89DrozKrt+qxkCfTnTGWr8Nfb2WDWpqXa
Ohas0YoH3XFr4sUz+MNdszhHaKAkvB8Eq03i/z1s5y/vhIqXSw/6m/4AqqdVtD9+yB50x09P9rLh
JWV5QIkdZlEr3KIob4MO6h8hWdeqxaUX7n9N54cX+MdZr97DK7jAjYkdGU6MhBUj9z0RMwOIPmF4
0ornM2m6venVqOS736aFrNZ/N0E7IhDVtZgzXEWTJJe+ODRM4z2TjudBjAyri1jsoeJBbNVK1uL1
iWalXZOGjjH92coBWHuiqIIJk8bPWIG0RE7Wn38kDvZKjq0+Qpw1qN1clBMyMtmRx425Nsi+HizP
lNo1PFLOAyuUjOkz355mNNm6JuRSHv+aXZ4u551AHYeun8bkXADLtXIXHRFy9n0fWO6sUIAS+aBV
bwWU86nlBqLafpGZVOO1awdP8We3D65yKwE2nY5WHHgu4+Jt7+Pe/M538ag4PS3XA38h41RAoXrQ
WQRaWVVp+Ny1vQPIONuZpQRlZ8ACrSjMArt3L0Mgpg33+9uBg5vY4pbBc0VRZyXm472llDSMhT6d
uFTHguqhi2iGfDIZeqfiISxgc32E8OlsLeEVjCUR8bu+FQl5/9VfBynO1/Ll26xvIeEfX5sfK9c7
KZ3t9ieRZONZXABmZFKPWSo8SQpWJZBpldI/GyNlSFO9ZjjCp23TIiJAL/+2Y4c/ouHkdRCYxg/+
YZlIoiTb4CvpYV7TyK8cAyH+YMBhBvujZLT0W5EaxyU8Eg81olA6suNxHq53VmUc+8aCblf8GwTo
j67m5cPiK7OyXxjiX2pY7SmV2EpkXZumbOjjKTsEpIVBe34Gep6LiwEpq297TJXeJTdZwxzEAVlz
h/6C6/f25vwbKgb12lXN1cUGDUoBsnzmm8j4UDQdTTT2QtZXEZ2Xo/koF+eOBZPKM6SWX9Oh6uCw
vBr6wZGcrXniOhE+eYESIJTEhuBUjUk152LUs0OSSZ0A/TyzAzNwgcnLkTo4fqWflPJLGRvaaLLy
JX2cOUQWC9aMixSPVEhfuhZFJxU4QPNQmxon5N+w/HbG1hDYujqUOZi3LNrQabfPzupby5ptVjC+
MWjKvANFYJ6QiBq2VUCpV88Tfprvv8+Rz04CCGIIoNHuLQr15CzDgHLl++nK+NqdXct0O7a6lW1Z
G/JHH2/wLJpfoI5CqwWWWnBO9KATIaNlhfWKC8wXku3IQN5rtP3eiFga2feQ5+wilpUGEnpfSS4X
gpOCXf9yRRlzAkM6UnoSfwM5cW5hKnZYQQxt4u9HhXojuABwTQrLgPx8/xVUp3e+h3I8rdvctMo8
9T1mxGOEeoQTr7ubGQWPmDONco/EhXUgnYY1Te/+rSy67FqdWLJ1YGyIsVXuh6EYMhhvnWszYyZF
FvMpYmUs09CTxEtOtFXhLRVATEK1F3ZIHIoaffG6pG+4Zp6A+Q+cjVCc/R8F/uSeeu2avNI9CcUN
ZAD5v7iksC/JHxOlt+4qkppJJPNSPyhIMlLrcq6flHqlOkyW9M00wAbd699XeUqB+ie2bALBB5IJ
u5oCkjfsx6KccTVaHa4ZEPqrfaBHMj50cF1Ysi1SWUGZ+kCaBJ84VxwyaJPSSgVbkgdT1SjbZI7M
sMOWch94Xsa0FoyLvXabqJgRtBGl0k2Jh7I+7zHM/GrzAsEs6V5LaLi4/6lDA01nGXw1AkumwzPh
mJMirTteBYWdDqnbY2L/k4+V19gipgJApsXU618zCNoGMHAYWr/XiOS+fFeX1kjg8ea+Ou7MoYxi
cv9SMNxWGGHyRE6iTGakOH3Sjph2dB3buFlEOfvns/Ds0XjCw1/FZee4dHsRcWrSHln9R49C2IFo
gwavdZ5J2A7C0wVNZORLzOyYhhSxuImPoUL0gUxppvOidg/OkBEUzgDvNbv0SpFhF4ENo+PNIIbI
90Qto2c9jGl/sWWCuq8EAAXXX4jXasnMgGXPUX21bbRZIsgGYkb3G3qyhXddGlKkjJ4oSA1nUfUC
3ijA+ot/Q+04KttfV86C2RWN+OSspxrxFJfgUJYNQjoT1sv61FlHlMJYaHFH5SECcNOWA+DEc1sb
tb7/qBxPyxSvurGNUpf2WOex/F2F8LJnyPfV3FyUEzgpBey+5WuD9zgXlHzcelDfr3vfe/fZSkpp
0MpXWFdUM4fo2SxYDWjumlagQjiQabscTBeU++mzj3XGlwqhOUx+fiol0HvU4uYAQr6wctDy865M
cl9OK2s5oRn/dp1y/U67u6e3ja47YgnpMwlqMWvBx1yRhzHIr51aOf03yM7XDcLm15ZtqC5H0Cf/
RfUwwAnbiSj7zYJmzAwikzsat8whTvlABy4itl5d4hKnUOt5GL7Paz2HZoTN6znYhrcWfWtmZEwr
ioNMMFLeTHxeYEg+3Sk581uPtVYcqTzp5tDWYlasAhIJ1iicWJLbA+1r24enOVvuo2xCZIUDvjIg
rSCLgYWJVYmtnxF3m1KAIkIMrdrgnDJet2Q9478sslvjIb2y6Uw9hx8957F0+T9fVZxnF8NaHUqT
JvRbUteWzS+PROswRDiMCcMvTy/oqqSdyTM6yPGB+6iV6iLnqw10nfx0Q1Dz0w5yrQt9oPm2rpfU
4rAn5/Wn/RIB3jsS1CV5etiLp10+RdjPOxpXhEoFKxBOVselR8XrgyjWlgqnM0OQOChoABt5bPCa
JyX+JA9J1ov0mrS1Dc+EhyW17WZfS7+nMMVrapITIZcx0du/Qvfhdn8pFEvNW/H+4YugA38a+58e
M4Xol5Bt8jxwKlzqUbun8/KPsR6upjeOs6oaXZOgzvA/cE9eVM0h50h1Sw+kjMW04ykKUJAS4JXd
gJ4oBG0iZm+4M5T+/MzKAS1pt+o8GAtfrXwGA7eWXlfyuaNToh1LaqyhktmefN7HuQcGwTnF+WjV
kQ6BO9tncsejCMrM8R+7+y0phnNWIJn6Kjl+ecgCeyfYJGrkQMog2YQdV/MDvSqmPzOyx3s/R1WD
AjAdqYfeO3g4ZSdikXqk18nwnT79G2TS96eRWYx9wPu7731q3MHXkqQnMv1M9ng0Q+N/aUUm64iA
XMpwn2F8WTU7k1+Esci+yjJ+5pc8WariBpiAn8gY5KyEKKkMYSAGFTxdf9pScmXJeKMoB9WavL8/
hgimSu7RNMRf18iZmW2xU7OeDYPJcSbhOJr4D8Zw/0ZSPqLk364LTE+yZ0OVIhPBj9pvgzaI7M6e
weMuB4Q0x02F/+2TV+VK+ZFU5QWM+xU7oNobWv73LaJFPSzq39K0AWwTvTZnFlzeO1wt/+vEsyjn
OSZHBXig5ZXezxvzHht2CSFCREv5xY4wZRf40iIutN7plyVszADX1fkNirit/XcmfYW/uAtAZKLc
M9+7hwiVbaQr9gBw9UVSRfWm848Pkk6onNByGCwsFHtrNOH4B5j2k0MvvDduzXtN2qaG+/CTrbgk
/lvk354vFTHiS/0fo3YBnJOA0JiaSGe8hNDDFknFM8Fl1sAoWBR8QkL4Dvi/KrNPVIu/R6GF9yUm
L/x9dlKBbG3xZHm/n5TR0B4TI0GtvsF7Y30DbfQ61B1pTJAacJo8edqsIBpIiIWdD72Y6p3rL9+b
6QRu4/9JAG3mjVHjDkL7unpzmnN9J4zc2CsjYR8ZU2LTxrfT/MyUwUj/1pr06ZFrqldwvk0Gho1I
5D9dWPXAhUPuFj0vjhdGkFLiPYIjzr+Nkx2SH8pPIwCzoPJRfs+yGWbmvEDGbM4IfdVYvcg5Snwl
uHJUHj2bvyD6oien0VJi9iANj0xTaOV77DTqP1hjhvffSJ7Al8hEPAJI3aviR1Sx57yUOM4145nU
meoAV3lzc0c5rtgAc/QRjtN1dA6SoNYx9ll0WoI6BltdYs2JWyGuasX1CX5cqnZnrnXdvF4jalil
50d93is0d1G3EgYBrMaS2EX4eobwPMxJ5q0pMgI8maFEBIT/VRJskB+SaBbfbOB/kZEGStG4mXoV
REKRJR1Sw8LyYLPaqN3p4ddP05/9VuMsRz13bFsR0mSZ6MCZhKHbtdEwGCTOSqcANhrzN3CM7omD
Tlchv6q6uLrEi787+zKjMYjtfEUyO1HJVAD1Gy+IUWB1oC3arv5yJMk076vMkR7GW0CEjZUFByHX
Fk2OXKqHAXnjsuaOesjta4ZUKsNxSXnpA5KCp12/GHlO2XaK1TawnN1LDWVN8PU0SGgsVR0F77Jk
uDxDhMIJOtDpBzwnDM29QmdxFLe45tZcuVe5+GtRoUdlmI/nfgC+g+1U71RGjNTc3CLqyFLVuUiT
0v8+X0Gbo9p1r7Qy1LLG3ku56SNTSZ4k1HnRYt1FN6cbvvz2X6DyF19Jxojgu2Qms4XfKQxJIl+F
xxpEQwRl6eUHYOcDuOIwaY3G7XyvI6t1yBEP9EsSj25X7Yi5OChb03emzn5C12nU3k/nYpluhes+
V/vM2d9ePO9rc6rnACWHDdiIhh07FPySs1KIueDY6llsw3B6RTGzzd+jCXVNvI5RUqnxjNySoe8Z
HNz2Ukcw3X1A9dV5RgCpFymhQuWkteq1v/g2G9EAGlkdbaxb6olEvj5QNzkduN0Zw1rPoQWSXQ+x
0W6z40oDQ+dmDhbEIRHREkRbAkpsW445IbUdZkCaFoSpNR672Rm8I3J5ncCyLEhrPKrsbTuw4VyL
MYrXWUs83w3PPaWC70k7uFyiQpAl1csJwWCA9NIT51RcUFWlvC2aFeQ+PlXgefja75C2moKo+jYX
pkf2y5XNhXGxIKs3v6ZZxVUfcksk6wWKs9vcES75zoiZ/gDjs8EG7pq/u7GQ+awSe8Fb0s5UxVQ/
YgH7KdnxGaUnRJPd4X5gArN4x6Y8TquZEJg/ICn1knVob0lftUZBzklu0X3MEMvgJBxJcfWG40Fz
T88WITowDfYH/YnA13M/coqRSZ4APFTj3rU9/Cwl+e+ucrdr8706i4IOR/OUcgNW9NHd/tz8Uhu8
ItMGCBPlYG4ED6OE6CgubhgB9Abc9csaGQmD2fPs1Il7lAf5Dd9t7UWz8qIh5xPE/qHEB1sPF1ie
wFYHIzo9TGXLLuRjyKR21NfF0O4MtAPtuvWCqsHW9ZWPC38PSbXpCrn3RfnunsPmacceD2/+YvZ9
2MNDSSLdR25bz9QI4FT9SQbhqnlhGsDTXORpha50Ix+R0oDAOSl5xGV5tKfYJuQbyu+khylMJnDM
v6VEWFAzPqVt+ApjFZYOtG/LdsjHYWAvOzWTzk2V4Xsmu+c6n2GtlhO9zrVVLDODiNZ/JDnEansv
d/rijuqPobRsLdc1O22InT6esMAiA9dJBC0+N8qw8MpKLDbcxAbZueM8cCTVPY3rpV9sT13gpKnd
7gWCDxSCCoTJVNVB3Yw8h/Ec8UHI1zurr0pMKpUTudLdNZSe71/npudhtHp2olBWvt4WpI3pyfdf
dK3YzCDk834Df0lxrdJo+pCY3uA4x8u09S4AZy68SDyPqrFxBoeOILYPrU9YNmW+0/Kto23RWjvk
xCb6izmCQzF7IwECzaS3eL1yc3od0v37jjzHP2kejjsvhDxQfYFyuDqnP5KfA66RwzsEiaDpgtYj
Tlrfxik6PrCQMCzz9yVFQ/E/QXsrIn9a0T/D7VgmCUYJMZaWlW+Tq+gUupBxwGJCj1QORY+r8A9K
krVYhJsqA4A0NvJxs5vTf2TQ+M4BGDyUqDbyw9nQ9GYCnSKdBApqWpbnxMyqXk7HmAFPgXt2/3kk
psaAuX3WHC9hl9RUMSY/pS266/0OVaRKFplWgDYRKEUSDrzl6wVPUwaLl6dAo2w6Xci8+lZ4v04r
V2ld6P8OVQdn5FsDC58rTmIWQRe0fJgcQ5m0v3mzlhHFcCXbEWHJxuAC5jw7jgPie/ud5r0CIPCv
tWXvvS2c/E3xqpPJmK36qE/tL/Ps2ux4mkwpZPTS9pFAl1B09qdvLJd4wUJQrAxdw6CvAF0MRGtL
TTsA5cDGDTXHjlDk7LyAAeRSgTjbi5o3FQftIt1t4EIy89ccidmBbywCY7uPnqrhbNtU3bElX5LO
5CrMUNcnwUAQ+VOGHqwmxioycgRIINkUd1m+rTHr2e+gwmqKPSLsy0DKCKsA+uKZ1CUl+aJh3Epd
4CVXKUKicxbwPEViIU7+vbaakdjhBgdCapteGZjB/4qEwCBidUF/5iOQtodd45NI4bZB7AWM/waw
1crqjEO7iZ/8nIyU+mEGxNq/SWylMkoBQ6RVINLVIpwHrPXgC+Q7ufmKOPHq9XVPxR/LJJ+SCvjA
HGJs0KM7DDMO4+hlR6g40xVoCz+lt/R/lDoFNEHCB5CW1eZG/E9PP9TwEsgzyTHmEUh3ixpmG0i5
7/0rk98Ysbz3mvKROc0vF2v1StU51GxiUIMGLZY+Iiin1mIUZZDBnCZl96vTkDcSbBiz0aOKf2or
qiF7511lLJM7xx0JjsE55Ommi59t/8i1OEc/ry71uVZSYvZcSoduow7+YNsWb276lP9jG/lSz2xo
1zl0KzXImRoSCrXQ9uKse3fK5Hfde5gKcM2tTQipJdSdD5fiuIyO/vn+VXPK/1C0rh5kCbZM0gRB
UOggXykVz+XD+K2NXVhRjtnWNTkw8AEDfZNZlQg22edTJbcZXnNDTqUnAqeQBP+tQOP3ERI7A4Hh
4jyt85wDHe1qWxqBgOsnpYsrqKDGINNoyV2U5mKqKNB0kb3RdycVHiE6NtM0oxLOjWkGXqVlFSvE
6dR05/v6rEdfaAwrTPPEIiYuaRZGiPx387+IWvid5BTfjVMgu96TyEUzv2q1Q4y0PtlAn0H1dK7c
RdpzVqIXzFEAdM3qOwIvGJgdgyoZpiYlh29x5XNKt+VbZFE0jeCX8gai2l1CNrxw4oZQjvMD2cKF
0UHffY8Keh9lC0epsZaaHOAqiTGdBbAeD+8fbt+Ne58xFjx22uA19ZfvSidUdU51K80YbiOKZrds
fUTMlmvb32wmjsfmjH9F81XHH0lZErG22UZwDzOXY5/EccuXNmF6w7QXvmCvbVPA/au1EMqmhchL
DXUiMtsUIz04psF+mALy485ZC0UcdfM/kzXavEebBcqfXsOadHeRATa/M5rW/Q8X81N0d3drKiVh
2BkxzS76ja5z7uTatmoa7cqaoV5cJYYrCnLB60rIVLe5rE+DFBIG5hQCIzZ3d5xt6aL1NX19KCsM
eDUmxgr5aopK4slQuSMpgdkFPo1+b9mXnfEYrLRV2T/BUyVjURUnDrhIZVa/8Q7Ecnd8gKTU9/Sk
Tv2BrAJG4BpmgysKq0E/Xx0OZF/9ZHuiIx0sTiJpX7rLSIkJN7M+3MWOq/gED2qFWfbzMPuN5gbc
JJNzkgB11f3TqQn6AlxosQc+QCv4of1nFR5Tg1EGObaxifhz/2w2lNotIWAfjmw02StW4MNAs4+a
MLRI00hXhO+s1LgrB0RKZzQb9nEi9cLFkfnHkAWfqX8x+desSI8ZSJhzEay6nwSLdrAnygOEwStx
1a8yQy2CIV0ijKJq8lOKBI5fNlG7WG/7V9PZvtx3MyMcMhTySJ8ipGWEJKLdc/xHV/krY+RDDx4N
Y5XxQcn/FsBaZYmHh0mLozQGGWhzQsgP6IET7vaBujafM1wSApe2F4PyzmosmOXtryTQxwp2jiJi
0i/QjOEdZ8vjMrjmKzWQGPmNuWykCVfvK1Vpbq10TIKqBWd2zt0pdTEIUZhBiF3V/Kkq8YG00b1E
53erSQFeuVWr+jt8bdfA9BizmngwUXGS8e8aj2B9A43BO+2ePEKGKQyTYegI+mUiORu0H+jVC6PD
rksvvTS+guj309d5gowA2PLAHtknWd2VdYpr61p4I+Vh6aGiN9H/5WnnWtX5X3lfYgaRyjQyBcJP
IqhqpSs5ii2GhB38hzm9cCCNvkTLGZeTzJKIYI/qDO0s3XXCzeEW1UYBOhhhFiF0XIz32NUTU3G+
qcsxwd+9NmpCoKSD5qx83NOEd9Wmo/6PTDrhlF9Z9C1E60Sl+R5xGJqnpWnP195Yy4OiDBhOchUg
Vg7FXyNv3sExZBdAp/8hZflFzftuJRMcfnP+UwsYXmNoq8jnJ/TBqE7lVDnoVCk+wuLy/7cUYjbR
J+MomWhjRzi3GtiSLn9oMfWgAYaxcEiqUKViu25l5YKjVosIS1MTSeRDf2u2P7JaeZb7eqU1zmRZ
Wcv1b/oMK7QUisWChV9i1UpUlPcYnk4CdCWRgJ1N+r8MgVy637sVla9HTpt96uGjjFL41E3HW0+H
KxEWYogjIDYFfLhoXmbHsDn8ra8ZWxc5ZW0EETKZ0bJne6qZCHJORZGqFp0DljTnzDSI8yxoiDln
zSEB5frLlrkbFQ4rQSysPbGp8hZFsKh34lVsT/i8bjIoGVsiPkoPrsPXHcrs2Jhkj/Vhioz6uVgr
niq4Qg8qx/wQ4nnJb45xyMvVm21wWnwV+p3tL95J4s29Qbuz2o35iGGU/i4graiMKWyyJ74vSJGJ
5CvRjGWMtGsavUWQi/iL+zvStTxTXa4SMGugoTq7ZE4FUy4jFU6aBy0YoCEqm5W7oyJMnwiaaBLy
+/ZgFcJOn7Q6mlKf9vTJP882PdZFdisVshXpZK49ktPgI5UBP78137KIQs9ifQmiOJc1Hjr087KR
YSbsG8G2OToj5xOtkke2sWRYn/Fm/IY/2tT7IGJgzie1eeVi073G5wCTnphuQS//xB7LTXudkBZZ
zKabeE2tOSMxmnHNUQISID3RsztptkLWp7y5YL6+NsZK35/lkMyHOuMel+X0gZCXfi54I/M8KO69
1izsU87OadpFZjREJtudw3soBisH7any6vWoy31z4a/yDOWB61KjGXzNbvzHYB4T5h5E48Q3Y/aW
FqypK4UMifQhzCLxBnUex9P/TVe2FpBIsb1NR8XLLORfzrdDKvbvfjZzpUJX9oRk0fuqPkLg3dHP
/elZLB7y5VoQn/VRbcyfI/vOYIXZWl7M1Sp0eWI7em+SWc1093XX/XKC4Mrc//cb1Xpi7ZDSvgwX
Jzmw38chPjF0vLBmq4bJfGniZMMP0XepwkccafegIoOXe9QS0re6o17KpH4NXo/DgwMk0zkh62an
BPLW7uYn+OomVXmQqPwPjdjFMZ3e/tY1eEQamWbcbJ8P7YwRzjkMxAOzTyIoJqPFQ10paucbrvKY
/gEQ5OxjY8yKlexSio0mkJ5qcZYSRTH3Adnrea5fSZ661HTi7I2bYdNnLWk8uACyp3UKXCgq1Bjw
nmL0uwmuLSUWELjoEGOH3R1zlqsTMsBBC6uDGvjuKABiIks/n5OinbRdeV+yXWoOcgE+bZYfQldO
Vfo0S5ssDml5F/ae6NCbDj7hmCCHMGehDUXcE//XGneEtFUzDKc4PNHoDLmexoiCH0HW/7LOVNLY
KUgqdBD3mA/iPPBKQDg6c//OwRZf4Q1Med6c56s+W8AmWtyncNLCIWXEEGvH+6n8P2+pAYQvWUQG
i20cVgC7nZT8hwE4mTc+QpF0uOc6cPegsJvjWVIYiYZkJdu21m4Iq/+Tj4ms/JcNSvrDz7/nuD1A
78Jx4sR3dZEj2WtMuQrN4LqqAOadQ0UJii58zqDZ0eMOuN4tiACjrgVU6buF6xeVEovAzAAjhtm5
yw7xWzcfN7Y4cYCeE0KjXKGcvSIzz5u3GPD9CueThD6DVUfU9KAlg7p1cHXsVwqfs3vG6VsDw2Kd
bvgj791qj3kxx0wA0JgYD8wiZvI3RteYxQHl1MtlNgEctB72nT4asvngX4bEoopyK5fcQBpi5dB9
mRskJBNu3dxMK7b76Bm8e2HCyxxsiw5LXzO+TW4wYQehQtIQoM/ekjNi5UvtLR3GRFy/CR9Q+L3a
MQ8sA4Y+O0jWfYLsUBT6VEiyJQYgxPFHnp9ZcSCclfOOwHHCvyuBkpXTlm2N2y/pdUh7xM97ItbY
cHP5G7l4ACXU750Oh/BSHtrxgidEHIVnha/+urjGgtG+AtNWFYAJypzorinvl4OkYu8SZ8rhooCS
ZMSs6aNFsgkoq1qewSUrsoT9YVmw9hjmh/mQcUHzHY1mUt+yUlBcNjtCZJtIL/V3Gc+zdyJwS53N
LwemSf9CGA0ftcYds0Lo/hPsZR4GvjH2F6R1/MVB6HncJTVQ6UOn0/QsrX2IRTSmmZsAeCQGhI/X
0HijWvyEr1z2xqR6yY6Htzr2QHoXycvTOICBexO4oCsRtiEnYEdMfwPQTXmRI6qolAWn/LgYdwY+
ZNfOYKJK3WPmWRTHsq63n+8BUuBKTMnJEhPZCMmfHXNBOgG0FzXl7/0I1sOgmfuysGiupj7pEKsT
QyhUv+x2JHN3X/L1P8bI8FaowHPNk+CvC+YMts75FRO+LFdVEs5Xvu+a3J0SbsJ9HQ2jwmUZVsNT
abBKuEOuvUHtkCeWvscUDwLKAJFrlfgn1e/VQ2Ne3wSEsxT8rTnl3oeOHl4gL09++C4Nfc/NESCv
Y0/TDAyd5EkJUnStgU3rhURothlagKMVRhSSj2ztyiNsOM8TFLh7fIFtWyN+6CMfq8W+pa8PPn5E
80JAL7HBJinlINnZVFWml3KAiqMNmfcaRQFcORKRrIKd3rWw5X5Uf7gdOiSgAemrU3fQ+cNQQW0q
XoRpBlJNr5RNnZGaGCI6o4UirBPweSknU7g4T5G+T16cBTsxaFrt9P6hWMeFSB/ijOY49c1KXr22
mP3h4xslOuiaOaco4a6JafkUxmHj7PsjjyzfsZdzdtEca3QGW/BL1n8FvAROVMfuyAHe3z6wnqx4
069uBMFoD2VvIGzLdnfv839mMjCL1auh+9ZsLCQuD8am2uFNx+AKLVKEY3DuAjAfSBwNLj5wp/qU
R1YXhj0IUI02N1g+cgQTGPl+7qYrxO9rO85tCNabp7kVqeQtdYhPae8KwEenCx2a8Th3kt1NjF4P
LZUvEHGFuhiLtWPSCUIM2ikjo3fjnF4afxuvlHN43cYFB8ta5UW9RKT0eAla5rc/X09Z7H++0oHv
boVK8TJCYNYixBO8kGYgL9oohnvmkpALtna70MZ064OfPBlVY5rmn/vJkZ6lshaEdJJWok8QOmHT
808IoHK/OpFbzFO5cZmZIbXsXUIdEhcMLYAvQ/ItatRFrqQs5aM/jRgON0hlyD2oLQC6U3XjHEyi
wdqdkcHdzfYQlOtMRlezO5ElVqrN0quSkj9oklNugsEEmtW4pfEdMwy/duBYTxdj1cX273l7lMPL
EOmirfcHbSO0ur8p0URTalz8IUlsAc3Zd2YePHoccM2tNRBy1eEhVz08k5hDJgx+FY+k8vAn5m0H
LzU2e16EkT7T/PEgsvsdEz6mYfBtiAIqO7eH3kuIzYhKYPmyHGXmgag4QJ+drpfsqeUkigDY3Dd/
mB1QY7mnClV3eepaIr+jpCGthB8fSCXExiVmqRCuxVJQZm+8qZ+8httqgJSIGkm03UBXxZcUJaC5
Cl8P0ScKmGCgiZVKTr2ssGTv1crJ+vjun2dbSnUdxNg9FyB2UmjkRV0NRX72MbafWJvT9eMCCjPg
3u/ASnIvtLHF9UHC83UJkeXuL1wNzYr37YFSZRBiLmP3Ze0Bs3b4TpJjXfpuyI3ayzHsQKeCMclE
F70JbZnGOlHD7BntZCcJHEDm9qNJT3ZEFKWelvqnUTfpOmqHuYhFmgWnGZdahC7I4fJCX7S7U0eM
FL0e34SIoJHjIIMw7hDI/V0ZjHhfwxqjuxXtkJQyDf3pvKINu9+U8gI894dcZrhu2DzeaukpCrvL
7u2Z9ykDQ4qwC/xJRZd8ZlADxU8p/VxCfO5Iknqk4d6mEXUEDjRyi/P2p8eOYR++pSfs6O3x9/VT
cceWVMeEGDzO/D1AtOtwulULPwAWntqmvHm2NWHBpbP1zP7tQkcdR+ve6bqK2ijVvPgkAEyQUljb
xFQkFSuyPrgHC2vHnErT3rXz/gm0UXkcBje7IzUg/SpvIxLEL6mG7zQppdqVA4++2+XgQ7wol9Va
9wZ5HKau1DrOezZXi1sPgsGElWB7IO4KNtWVroPRGgjb08r0ATX0pgTnR9dYZHnTHlfTnYOFBDLg
zMtIsMgg3OiaNtZepIhOJtxMfHxFjfQy2Mf34iLsjEpvs6HoZFMZy0n4aciV9gwRFjh+cYNCCw+/
HKkA83l5QQ4QulHYllJSyQvWtYjakbz/fZZgpsCcJGA0EK0Z+ebdd0uqW7KSEQZA8YxrsXMVHfdh
tcYNkuBHX5439SFJHGReh4Gcipki2GHs4+wc07n1hZhKpMOXEZ6wV7AswBKNstOX9ZyZLlhv6Cvj
62quRTu2m+8uS8dXJo0Z78UsyLZDF+KRPYYtueHhJSlCFR/pZGPBVDlCfIegas4R74vSi1DGKpv5
FjcxIvr/Ke8YL4VELsCdcMrp+7JDPVz5qqQf2Rxk8PkV+C847cspZUBbQWzEa+OTKzX/eDd9kA8T
RA/upJgKx05gSBqmfSVFBBwdW+ThCMBXVCDYxnTJPxmMcsbU8Ehhb3RsyryG9776FsCieq6awtN4
p395AFVQT+PtUvVXr8C7YV9iyijipNGHTDSIB5BwrGdvpNGJEN0RTdonpX7SooEQcQTsAYquha0C
wbB7XZ3pcyU1KpKgCVpDM10SlW1K65G30YpFTTYDQ6PJ8xlNWBh1dijnGd8DNmpcX8TAN1f/StgM
LT3/Tlo21p4+pdVF7NhJLedJT19McElAqhOOuNZDIW3hM/wuoF1CpJtWFsoScWW1w4FJUvZAUsul
ZOPkEvzoTzgfEXkU3QXhNfntf/qoxMf0qyhzMA/FucZh4x/UlQC23F08ICLSsB3oKSKZJet2u1A6
PfybS4C8CePt/xYx/u/7TypKo0PwGbVULNCbF4U+XGSeKK+TX3QFAokpV+9CDSMhcFtY6guhaPFd
UsCPpguL/iopa9XVlRV+g5ksocezAq9VNl5qGdHSjdUxtQF2Q1wOJ2czE9EXmn5PH2dP3O+YnDN6
XU+J0SLa181Xlp8ygihFrftnn+zPuGq13Sl8mc5fncW69BbAvcPJc7Qycr43rs4XRxGvZxL8IOmQ
sbcZunBT7ynIicVAqmrF5G5ZCXaSQsnKXISAEKhQ4NndVm157ZNd7duBBIcwqau+MX9huQ2x+2kc
YDNX2nrCrDP2YpllZwoimI/9odUBeaoOgtbhQvPKuZgwhD1GXdD+/0VrJMbUdXHzT3cXvFn+7WoY
pO0Ia5I0+SAPatej7CVc1mElP0d9iXtulkEo/qtw5lwpSIM+VhbgEiNxgojdmsCvlT0541spByvx
8PQlX3kJMOOdfv4r41uYFkTWuicxxHD5RIUB0VpqgdsCwX6VFmHalPq14eDVMVsxL5fs1tX/bZ/y
wpDreoFEF8kXbiQHbAUnAe3/dBBHVLOB1IR9SJ9++becu9Ia+q8HGeNxQ8kIH6A2Yp0ADIBpkGJk
7X5B6XDsx+zih1lmh79rj8FKVn2m0t621L8pZyElf7lkr0xD21ibMFsj1Pyi2s8wbuOGSNV2Vxly
Lj6huoqVNQW053GXZTuVAA9x86cg9uCEg2CtrRVLBJzGMG+aLZKx3UxsGHwNmqFPQhEy40ot/28k
AWtqPDr4U1mdsMQp4v8DN5edtHckg+i70AhTNXuHHEGYuT7oP4WbYTIsn5nSPITQkzgmp3CcM6mp
+9kb/t6DNKBRnTJcseeXcRgzZvrTS84iG9Cb+uW+5OR1D/wT88YUOrNDm2lNoiorbMnkpQT9cR1T
/+/tAGQFgjCDzmhDiab2aQFolWf69HhAqqU+qfRaVrTdOCtmN5CgxSEfIU+kYLkPZFQZU9ZEG3lx
pIINxITo9AVequYxVEe2w73vHLHj4TL1Ij93TsHwgxu+mU4c86oRixqySrWPMArNNX75Q5SKnECA
87NT9kwkwGkepP7QxQQZw2ogOQuBb6xf2TXlQotpn3P3OVL2a2xahD4SVXiBni/bvKuaQdFL9u/J
3wRVuInIAJw4EgkrBUWjfH/TRNN7ONQXRDCEWn4gfx5/s25k7QskPJ3o5JuSdorWaPgiX2nhw3av
NwPthMdAHLQ/Pz0D66F7nOL3cI1C77scutWsfhejLZXS0gchyJGO6qCKx//hQaib0wQ21Gfm3bf6
556e6mA/xKoqOr4Mh3wjRjH+4J82O71IUHp4YSl1+iz52q4DOTZBpuYI0N8CdfxLwxK1lStE8df0
BzFmY99kEuGyVqul1lwt8iBng6Ldjbq7L9CECxi2u1XIPXoomVF+j02G+4PpH/H81r83LXcEDRE7
QBHDIPzd7rS6tKdSc4rcFr6Z9cGtlOfYo3SzqbFAGJt0DlwZMAXnq+hAemooqeUO2r1EH313Bqwc
Qma8BkCQlA1nwdiXF4Yx3oPB3AJ4gDUoY8ZYC6ezWisNB7u3+Xa69368n6Va2ddoQQsZzc8cQQmD
PhLUErQdY4lzmumrBlSif4a2akIS75jUYusCC6/s5znwJqP2CsPKKKfr+1zhZTVGo7EL+tB/L+jB
Po9GBEGzyeCOI8bIh2FhbpfAzuKLI2nnc3pRyK9DrJ1V3vaLrNXlYEzBshZ/ZdEA/bfVUdWXVRfQ
4YMPS7HMXrx1vCAP3JK5KbT7MVj/pLiFD8TMqiXt8fzPD/n2Ghy/CCjYRAsNwAdSWSqsOXD6xjhx
1JeIZTqmfeGJ4Nt/PM62W2uFAat0s0ds2usw0LKonwKNv3KU5KbT2nNGR+qd6uS6rxkSb3JP1wBh
umcOapzV/4p3KdTzZQA+eCu4gNQkrRre7yHx6DlcCO/f11Qh4urvwHP/cehUIx7ygh4hL8LuXZMh
5spYWT19f9M6LJ48vdGaRpwNpyVgCB3u5GJFXC1Uf4HCFvwxwXYdtLp1aej7RqLTSlZI2EDYM7mv
11xwPDQ0I3xBj2LrhD6RfMOnNc9q1mvdBFwJqX+ZZo6kAi3d9/XqhHg/jcYUntqWSu5OyQbKgVNt
cQi92Ta990pkU1OY6PwMcQfX/8tKk0TSFp2+wD3lPH6C0kCJT23QEJYEZZo6h99aurVLsOqLSwM2
ni7CbbZDyAfh21UR+qGf2LFY8CSqLEr0oIrpKZrxOQOOWjv+Ca84Ou7gzf7vzCmXVWO9GTZB1icn
3GF+htchIi87XFoa8BzbBg/NoVBLRFQFD9GiBPcb6s5GQkGAwazNFT8c0Hrx/bhr607o0z07fpDQ
wE8azVCHApCsAsGDLsHgv6uSHikhFCvvzmsg729JLevmDcfRJPeCbo9NWYKwUZPobtL83q2EWoPs
q2E7Jaahli4fB/yR6JboaER5A1g9OMcypZ9wHu/kpQspFQFH0gIv07vUcUms/0qheNigGbIezarW
DTS2ROa66yMYtEWVlJkyrm+RTTTAX0Iy/L8g/UVFumISVp8V5xiLDBJqTIp3FTFR+HvsRGjS/LrY
iA0Rd1/OUUFQdvanVZq1ydHJ6q/CRm4MX5K5TQyNh4eKrHF3ggSzjJRx3Al9m8Oy9L79Ts5KgpJJ
fBBh/epGvCKSq0zCDA==
`protect end_protected
