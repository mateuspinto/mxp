`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AmsOsK/A0LEpz1jHjWkrE4bqibWxKzdrtuIXd+t1s68ZmTtwrsMAbdLSqgAZZXmepvanFYBF5ssq
qTtpQvfUWOsA13USSKZjCQVUZaY4SutPtozI+ywnVxikjXeKk6Mx2TNUICV+ur3kLQwVuHgVEZGS
nbkXj7ZEO3dAN/MhK8uKhGZAZLm/5opJxDZHQFSP4ZdpR2o3GrwbQQpDLFgys3/Sb/3H+NpBhOMB
TTL2/RvQeZ7YXoCIOY+zyMpMiMhU2pppGd3EqYs7FRmSRYSKHLddTQHNtczZkcqWiQnrYxzCu90c
kzNA1NbN3jxOqgnxbnzUUpACgem1i57Wg4dg7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="HCSZYL1mau9bEMcQiISxMP72Whw2agbwcsDD9re/qY0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68736)
`protect data_block
JjL8/4h0odlz2fwPh914Eewk/P1lKJOQh+iGm5Dtt98rFlKR8RPl4MGVPc2cKPZ0sn8vEUnBlw8/
xZ84cQzcNB2dcWm9AgMYUM1bCvCxdJNdUmrVAeGOHpkJthMVj7D7j7x63mxsSFL0J8Cl+D6lVsvI
ADdBAEsxPfMtNYM6vNsHPdydV+i13JrtuXHTUQndjvFgpm/C7/AXC4KrmOayGUxkxiq54Kv3+Pha
DtsHtXnJFY4A3YaunNmxqUptAke/Iruk32DTOsJBWm+0tIJIsOmzEG0xY81+egKrmsMQwDjEEjjS
0sygXSSs1J01CVWxcQF7l4rKt/I5bIpf2AwkmukqpFh/PFk4UGJkWIkyDJ52szmSRF2qJACykr0x
QWFIZPSGmA0CM2nmwoJKa+1a0rcSJYsuaHKu2DGM0yKSBnKEmNhxiRgJJXfmwX3sQ1NwsI3O1yBp
GuciDhrL3bEKxSGOxc9z0XFSyIq9oBBKoPV0858/U6YpuPfSbWqr6pGY5cLfDERoFrpnlqubUd7V
pU3F+brG+spsu4KaZraj0eDWW9aknQPcehoNPKa8qoX7n9ux/OzXoNke+CIiC9a+R3FKElmT8FYn
pWPTCM+aGzgb5t/ldb7ULj92QO2owUGQXOvQj/iYR66Yj1Z28FcxjXfm0gDScr1p0Vlfa8sMicQk
cHMpnJ5x8rSP2cgUQlV46X6vh+DunOXVsg9lk6MLFgkVSXDWhO1LulYrMpQ/ZAK/L/iFFx8lZDGz
qLP+NGm7cE+Ynt8AapyY12WriEiidt/oT/Q5/Emy0jQok32kn3itx1PUKcIminrucRlncU2J4cu2
L8mpN8IlWuMu3j2aGUlJegJAZ92BijTlS1h8wDgB13am6DCkhGv8um4eAU2rX8W2LFi103oZupHa
36tAc+eHDAA3hObSDFcx/GZ6R/OZmDEsyHoruqbklOsCpFf1WqEo3/ri65Kt/WqTeJjY/T87geDH
kM49tPmm7ClMuzJmYdeWrrtaHzSCrQRJggHowFg8nJ+z/UmlovaY/qRrb/ygHbmoQjHDB6QpN3gv
G0mOpF5rpjx9ROLtNp/zIxS9Jjc2/yCWbzrWBJYpgl9pYFwSnvIlHLFeiNsda8+ektIIrq31rTP1
UaL1Zc9fMNHWnuk+lyeWyUgn7hvJrGmqC9c9l/IPp/BmVafKTy3QeEfCpnTL8LhZpGxGmJfBxFhu
jdmxTPxSnMOvSmzkSvPBtKbTzPiPHb6cXPh8Tr4Wz40HfPAySeU+Rn2Ql1yLFeRSw/vzJGmnvh5Y
ul5cPZx8xtTkmlcboeeWgvR8AsE622EPmddTCP6Ti9a5uRxqT1QKQEOXsv/XEp9jnxMSbqB+G+06
3Opkxe2GSUWA9rnDBRk79rS63XMo6js85ErEX1E/n7Nsi4E1sHicirhzbW//quHUt90ANFj40Xoo
CjrszrPd9ukTNRAJ2+utOXeAq0+w/elLPEz8QjU8EBU46hAZDkrwNNTk64itTmKOzuuWsWXKAc8e
R6ZAEkHVOX1kxyfqATic1ZSik5VOtjlPGjsT3NQ51ndBGlufNXsuhw6t5VmKBf7JNCggE7pbmCfk
ey1t/oEqYmHfjftUGH/5FXupLEMqfVZZBs2/9Cc1ZxLF0oYbTI4MAVL09NaAc6O0vvigYNw1NkO2
U2F3x5PzAVzQPvNYOD1olpE9BvOJfHuYbuPZyWbKEgfIJMV8zGBLl+0r4A3P8MK1uSRKgKQWTyLV
Kobhdaivh+6RRh/Oj8KwEAk3wP37bXrN3lx7j1+YCg0NyEYYtsjNRVpKbacsZOsUCzMVYd6DSBJ6
8NTYwEaz0LSvuzMbwlwr1FTSaCo+zVRdsMfgxdGvzjfd8eJjc+nRxEbdp35cys8/2kpfG2XRvXSX
VZXAltksJRHpBHk+jePQ2TsKPqzURJiLkcw4WRBOeLUB2vq6//neZKG9uXyE4A6iiZpsCyHLFyjV
iAlxZnChiVWAJ1YfXdaWTc6F7e7PhEX3GCzP/RVIbJv2iAB7SI1rS65YPrXyg/hIkYQa8taGcRoX
PLhM9Yc2GMMzFEumx9oO0Fy8qFCqXIdLwHQzxNUvM6GXz/pu/8Luktk/z83cHHsJuJx2BuBA0T3s
1ZViGGg+num3YOachOGAGwmPPWSV5f6zTm1np5q31T3nspoXQ/E7QWfmn9WCxpv1J1wxQGckAHB8
uqVJ4e58HE/GGNaqLsNqiSHva2KCey9Ba8WW+ISbjIrnuA++CaGM/c/Ouv/CKqis8/ZEY73LmRkb
ihZRPJbtUPz+MAgYUI3L6A3ysm/UDMyTRfZzhoferV7SLWyFLVHybm8/HlJ0nxG2L6c4p6OAqlWE
GW0DoFnPLZstLhLUzNGdqiVTchRQnbx4tG9+wDVbIsCaOxg+mIFT/N8eMlGCJ1PP2H2RRcrEpTPm
cf3gm/YNUfuAfNG+wtLk+oNHQgRNbkCLRTYd3nQ3A991lyw3UyiCm8AB8xpT2tKUrSwD0/syYI2O
j2X885iM4pYrQpgx+pA7x/D3I1CgxLr4FH69FFVVWmiJfGOfj6GuF/8/634DdENxx0lMr74HNw/z
G92g9zzpx8zzcwcMYwQmegJ3sh4otmh2US3iP89a6U+5HFgAwJF7xJBbkY+bj59XGqdOHESZxDZ9
C0QdUtPRVhhJxSOTYKI4c8k/61z7U0pmLnk9foBPwCIGU20O8BRCDKVMNQ197za6ITfDR9TqmhEf
0h4tUShFnYGByCygsCIoh3hSrIhjLOTVTmo59vaXA5qsCYubyGWeAVROEscqBxdECLE2ZAn73rbv
xbghC7RJ4ZQSIu2tssCE7sdRcL7MEgl6OkVCf3tfBctMrsbgxnWtuDoCNyXbxa2TnWjg4Oay1MQJ
EpclaqLqxj5aZamMPEqxvXF62nd4B6dNCFQjBD9mUi5ctju98Ecbiw2GEx1z5irRJf1XnmJiCLyS
hnvWz7OAawyyJxbdzcc7aw9yxq/BkPTtOLMGpaEGbeC9EPIqPRD+n65P1xl10OAjVk4JqZ6vkDPD
l29r0yPa5Qlu22SYFScHhEklkSt81ENdlDhsrlgGOi8mS7Q7hbV5n7/hqEbPecV5WTQ712gm3hDN
QQmaIJbkdzM6JxLt9pU4smgMCK4LhN93tAMFwsu2gDBaKif9sDXgY+rRe7G9BkPS8ujMUrnJBSn0
q+M4Uvwp4U74fokNac0lOIoFBQEx+ZI3uTjlYKLIGsD3yiUfdvaEb7CuQLcD+RPpOhBPKdOPzPsn
uHTki/dhHiRB7DrVtYwifblAN/V+DCu+09jHnZ+nILpmrqNXBTV5+mwxAP4C1FJA49rbiPQw7pH0
d9gIDWCG3M4x2tp8rVblSUu8xG+ezcvOaPmh70lp3YRL46SjMUQoFGCiZFilqD4ndjtyjfYpo0hk
dW4T1uOHtxtcnKsU3+j110c2RwrcydyfNsvGoml4pUk8wjWQC42Sf6aNZE1t1x9o8gy/epIu63gT
ayrFfVuS4qLTZau5QjHU3jpDdoWAVLmH4GPkfZRq6QAELYaJCf9xkCdkJqiDqNexmM++nDD7P9hh
AseNvAazH2NjJsivChp3UKZbrtsLTU5atWgRB5pf3nAkfvnh+uB9o7bJLOejYcDhGDoe/nMDQSGL
bBVN9kApFisxiYg/bN3jI18s4S3ipPgTZzCbbaHJfZXtL2M+g6WW1FYZUeVOzpctvfvrRUaEnzFJ
irnPtc4d9KT9PelsMkz3WPa91EWyTEMq2e8+uaWavRNtSLIva2ayUlyllBHD0ZA2lsm09ofvOc7H
KxbE1Ju2Zjunsomwh8g6Iz8hRSKBdJxqgIWozrhlQDp7tssY/pcvwY1fZN+r1emuh1bG8leCp3Jv
S6rGgQEwtqrJONUCPpWW/76CyVanXy2WFu4UJFNBVHtZ12K7B08Jj/4u4jMPD8OqzFKp8qQ2ga88
OhD/oWSgKuY17448wzpR0kjeFgRTtcW20LaLNDAGxXtK22hyuuftYiwUFOoSCp5fmRXLQo79eYVI
bNoFhcfZmKWEMrmdUKfLJo1coA/1YVth8eEaxr68DBmUcxZ4WEaO7FZs1LZ7orBs9nvjeCdqNrCY
inrlYDJjpL+66XR5RkmL/NqSr6dMmC7sXKKEwsHhxgKQ4ISfg/IK5SXddmBLt/n3rLU29uH2uj4b
ZXV3euAc5U1kzrmBfS59sAA3fxA9s8jB35ummk+Y8aY1iQ0d7N2OYAFcPFcyTvSXF6NL1Dj7zkZo
z4w49n/r/gb0gSMq5Y0Zr1Ucw97+XgJnfn16LJSz8SShJCsECtrFwOEdqYn1Aak6NO4ZkxMxOCom
PiDZGgzTcSelsDs8Q2CekDxv8nA5yZqtiaOXilCvkHnUVbs8NRCcziLenPq2MeV1ZagmCBw651CE
dpEjBVZUFVb/C/35fBCPn5GQm8S8H+CpGMioySjPUe2O2jbqCEQYZwqRwJMpTfQuXSO+HsNZwTw4
T0a6z+rlgRZinUK4A60dSFnfCPLhvt/htVsmEtMCIxsOwLaOJmo14p0C6nPPL+ZfLNYAT6adfIgK
YguA14wqraveOBisTOftjmBZmzkjaPS3ESZJqroeWNUVh5RlHCS1tLlxpVUME6CbYZrTDEWjXPVW
J+80krcdKkIZFW8Pa/8RxRtL32t2JkrXnUycrtWtjtyVQgmiXdJ+BVlKRhAvaTFxwUF2op57VR8B
IhemeJRorG3lgfc1m09vGjEAPKSmLHlmFMso0fVpSrACkdXH1bBbjbUxQ+b60Rn4CcLp91TEYPhB
nDWNKLD8JeRdmSUs4oJz5RUMDkr/CZHmjIEOZ/U2ro0fvHIMCsqtWz8iJ7QikBzNN7tu22McRRtI
ETJVrK3h3aaNjU9I/TD5wxhMkiu+pZyAMNZTvJ+Rk9joxnjSiLmkLQMocaDBW9lSg8aUMNbHgVCE
5pPFVi5GBnrm9Ctg6JohwP5qYIdt/RJ7YHdfb5GuUwZB0gzLxZ+S0zyk58yI+hi21ikGPoNWpXAR
VhuLlu8XtZ/s4QWCkuMCf9ozmei4m3TI+BQ/fTzL+GnQur4ldnnLctY6ZLodK1fdp2wrU+oeIErU
FZIMK1k2YQ5Hs2EsI67lnISRkfSuknlw2pWrxDlLClFOZNTlg44Rynpnll6njI46rGkzenG9Hl28
X3DAHHGbGb6FQKcsPl7xqN8qquZbP4uNtw+xCMUD615XMuG1XeTw7PsD6qCRO0eFBcC/k9FcI3U3
eOydvpB6FHU+OUOShoUXGCoIV/HrXkzTglpiceQVW824tenRvviAOJcxz49iASn1Z0rsizPFNmoF
rpAQDwYMBPsBHp/Fd35hgSbG97sfapWeC9M8JxEpOJJRojqDITBJTYn2lc1VcWkkKq3TLwHqwN6l
UOLZ1I9ynJPG4/boj1uqFbGssetU9WfahaQRSFJXtYq1WNnqaYpFrYfAUkPSpEQug4RIPqNnct59
w6xfDjTXUOYe396xY/FK9QmFbBDgiiTe3NSfMcAr4O3rxRVFfNCLIlGrdDRQCejv/UgcvrMD4dxv
YRffBJlKp36oZ8W50EylNbTq8akSHqSGPgs5b11JM90dMlAJrHMK/XWYsRQFKdxFJm9gGqoSFeW/
56Lno3kseD/mzKPCU916vXGDw0pPQvuWVeV5faEe8ygcVl+EI27I6Fo7Fn1LmnFFRwMMw3l/XID6
ed6wRn+uc7ZUY87FWkTKPUNIkd0vNErXPocxU6he3+sqMpOqIbsoYZTixwXU88DUj7V5erHp5V58
mmldtUdfQIx285oYJnq9+4oivUiImW5A3jK3f7REsYiGXF+zFXyUe/tZz3zfqF29GOv6KW6fiiRn
ejvLROkIuwjQ7FwMvGvNitSODKb+QSvW9m0CFSeaIrAxeKHBKGlfJr3eYgI/iiZ5SCgUq0stLdIm
4IfWBwoiAqwakM9VSRoGolX38qvfd5RyspouuKLgdAIh16UEwb1nufFyBslhbEM+zGS9hob2B30c
MLEArGEoxPmI5ygPup21Exf2bLvjR4ZOr361IDmHcfXTzIBgLNTASLKqoTZvSPjHpQ8xFiSCGIeV
OLrPFXf7h0CuDW8VUcV0zcNhmS1Ra8WypZDJvEBG1Q79vD1BCkRa7/bkRRQMel2gxnEgIP3mkHhn
8raToqkvQMeXUA5Mv+hZwK93bviEpAvjr76ViS8ewb4aLl0ufD/JDkMjQbCPOhGesIHq847Jlg0J
V+98V2j+OxIay1k8uglzYmEknxnmIW/hDFVFD5bixE3krSXkDS93tlbs879Hh+Pcf4XtIM5rkrQg
eGIECOuuD0ryZlHVF7BC1tlv30NJ/AVksdllLCGb4PF4qPh1g4ZDL9sGYpJO3dxUvIL02YUgLFVr
B+8hmk//f4JeT2vpDeCrCWkwj/IXE9BtWkKDTuTe+f3d655Tc+K4obJZn/PjpIeUB2gc8xdnfAJ1
BIYDH8A4Qttfut6NRvi4R2rS69RttBqcFzHFAI+JG3jtuO8gOrqDmvwssm1C78CDptxtHc6XE5jv
OmEFuqfSU2RvRRv+xTGR/fN2kH1tVhXo3I7JQGXEbkukrvf7xd7g6vliGv74sc+53jxQfiZUH3LJ
nJT3G9xru7ckM20raUvF7AzISluqk9c8ixuKbsVBOcNujeZzJNptSolz+jaOfKr3QjjrKU0/Wd/5
pcOreI+kPCB8R8X33HjdIWD0XAay8RDnhNNof+bEazjxcbknYvh8/qBJkVCoPdhhnmuP8/0J115g
Z2Pz8bOvTdI99IkSRn9EY+W+e+stHv2PTzmjBdTep1+fT9WJISITSjaidJPFG1h6ycH4+yN5NDNZ
Bo4BCi9OkybnjoqeCXSQ6+aHTh7J0q1c9RonIxkN3xUPcS5zbvzSzcUAGyaDm8MS2LlcsbXQ4vRQ
CuIrO4jrMv/zqUyBz/CR0VZKtUOjOIlmFfqCGg9x7J0d/VQsbDFzqCrbCa/qxWe/NDwBPslhWUfA
sZ5l0tpLGGLSGS+8dI954/kOdPSmsJ8gtjvscolSZsP/gbDp+EJAIBDAPhLdChInWsmlBvxcw5cj
/zP96aTQdny8p8caI36zVrVBcSXA7eD0rRL7tfpG5XXP+QfZhZzqjhq+CBLvXgIoguMAMGxoa1q/
/zaUeTkSqoC+m+oexh3/4e62RYKibsdBLzOsS7adaRysF6YoiIEg8f9f5vAiE2d7++jWrdYtR+MA
3VnP0KFDOAqjxWxiupVzljkoy6VbzooW/R4TLrJwZnDFkC++oVZNTAEZAEpg+GSRCZH4wptdCzGS
/Z0fJGVTSQVuIP4n+mlNjMj+XA5W0EleurD3f1LxEcMiAbG5F/tT0kBROdbn7BcAOygv2VHOoQc5
/5zD416+imoYvmif8vRccyYOA+L96p9wwaUT98RGuNXPKCF5F/JEDG6WIZTy9HagAbeYHWvp2LDy
/345icIta8to8zb6M/9OVbJzQR9q2FE6/LntG+a4lZBI0C8lK9Rlp+ZOvu3bNCER2/qC0J0KnEOZ
rn9ew8xPHcWDTEH2LSx+y+QUqDimpE0Z67r9ezxJniPWDEb48xdG8Q8fL2wWdN7m5Qk8zoJhmnsu
N1oJSspDBWMIYdz0CTo9RpofdLtC8maTRC95zjcRGcglr3zcFXaklStibHTscN7os0w3/6sQMYy8
qtXM98cRo9IJisi6h5MoPnPRre56EvLaAl2CzE4ohmj+KqiJn2vVi0ouIqH2nlThdSOm4AseVnoL
suYHzoniB5ZNIQ5M06U1FLiy7N5IMTsvX6gtgZCJM3IqxtStuG5YmBpCXTqol6MW3zeoOTfXpary
KGoDY/0LUyKp6rJa3F2QKVQMT/vcrtzY6FBo2de3OTao1Zn7xw8BRhVAXmURwIXXJi5WBhNmmS5j
pleY6ncPbQ8j3lEmMDe9QVC5qQpZCfnt8GhewTmsSBbizbBy+5C8YSXkaIGLU91EB2F5i0ETehdb
PrrESQY3gbIZbgR+yrLKgRP8qmRiz3o1xaDo+CaDEsQ8IvufjvVbjc0vIPRv6ZXsnVBdyKnQSzF2
Xwk1JPSrP71NsYkgKbicKT4GtBJDfflgYgN5d0JN55sSWPCtb95WxsePJ/vKdfJyw6JDG82KIWNd
B4JELtevXhY/aslISW7Xv7l3mIenhEMSBVA3W8HXcU6b1F21tL8z2vo/asYD3YrzyJFuEws6QUYY
YxVLZG/p/M79QNevad9TDBBhFzqrjup06UdQ/BH2bpWg1JejWuTrrY4YUDuAMXRkR/7wrXY91FIH
8L7woJIrtJNIQ7qhpPuhAAgJW01+aGyG62ot0+AkPniRp+UILrxUN0Js1Jqs3XVTedg4GLQm3uPe
cyqbzcoFHTYkL3FLqvCRwNVetp4i4skYCYj7cPD9H+T7IkBGHZSO5eaPcxurtnZ7aylq9Au9qmax
Jpaccg/iMh8vCFGVPjC7oF+NlEMbaabnXxHr10H1Rgt/HOLTxuMVbA793Va8ewpwMlXp4PnaWQO5
ZI4UEiIFRcA0Vm6fq6ljMm6zF8P+SjzpDmiVLo2gln49rEjSqIXrR3nkLJP11oqU0GLrPoYHokeZ
jxGVClkm8dB5zJNJ76BoksjRgmk5R/YaLcFKSXabWsjYS/4NYiU0E0Z0ZG/MHVRw8ZrbYf7tFitW
t7NwECAXlaNhRP7ZzDiBXmycS4OsDs/uLz1D8Bgi1ac+LE/upHQlPlzeXokY6pdnTsuJz04pQfgs
Ifn90B21I7uozoXBFdDbgPzJdkYbOIbsokBgf3TJWt2u288uTDPMR8CR/OXwB05qsr9fAUFe4/vT
Fq+nNiKLyyYSa4G0FE2QHqFtDAkkQMcP2c2GA5nrPOiwF2V+JUUM7e1TtKn/vbJSEmnED8s/V7Vu
OZ+Ac7BGMAkR/nLMQrVoLcwv+fwN0LBTX3WA0qczoxBgwsvNKfh0qDQ5juxBCNDgEH9rBxenF/h4
HR98uy/ZpWCdfl4DNNLmD9/mq4Um0KqTPfieDg/sfsLIwdQ9kPgsOHra4l+iEkY8QlHNxQYRZ64T
YKijixyy3+o/rHGwtzidoNNtZApNGtkZjd5kKBkLdgBtlIBS4DWzg/Td/OFavxc/yOTQFMZi7SN3
YIAYB7K+wXWlIan32UN3KDrIBScBhUsGIcpmfQQl5htbqS6J9dGriuPAj32vUTiM25V7FVxFm+Xo
Cjj0soEy7uHwGWuVPxPhc7HUfVve4JuAIdthGo9z2QPiUfTsSvk7EaRmfCDWIkJ/oQw4vJ1+YCjp
V4gkMV+AtDRCJ/XZH/BgexuEBuLjFC9hbIEE2yeOQTBgLlk0o1OeH6o1/4u65OAr5q5wvCSxfOX8
HPEtJ2Z8i6rwbr+54rmXAfO75IgyuPHBsG257qoG3VkA969wS+jwBGBvxmCWpnUYiSABCzN7VZvd
hcT7J/4FT6K+GdQbaJ0h/oBBghI2rPJhDt62rlhsK1PpWjtHHyCtiZ9EdGcpL+mVo9oXf8fgrbcZ
tHaVIEQKfRNoino6+enGBwOBTdA0E7p+ftinUPUGRQwymW7100es++PFXQZeg+OoD3O5DAow4Gxv
NzwIjgoFzpxImvuXFZx3G0Itkcu4gY/0yp8eqAChOgosAdlnFji9Vr1+1kpyKZZI3C1dxO2h+d72
ZHZQiLDgzTqsWupmaCz7eNDudyQZvgSXsI9pxbb+x2iKqKDE2JWmunsHVsk8P3tPrTcXO1uoTQRw
odosFKeNdH5L0EcjgP2azyzEyZI4mY+BGAjkH4W7+WQZ8q3LYiKReikowRPyuQ/ER4ro3SjfCbBI
5xQfPHhJ0Ud0aVPL6Yt8v2YUrK39nr5cntg1wdb5zzYI/iqnEd6fAdDpC/sFY0YspF9GpJlpNR6S
FFuS11bFdUOn6YbuNLXo2eRR7NWfawa0sSI3GaQYUdBwxa2Duuy8PhKy3chUIsgRhQM6wKG8VDSn
zdFcOLN0pjMLucG92NKRvwaZV80kf89DkyQriFopowbYiucyATPwx2fXy6jCOF7MtX699zuAaRX/
NzL38BJJ0a/llWjAakgmVb0l/SOAMQSy/aayRLZUhuFENpWpqmg6sQbBBpI7E22nBhZ4EWqdNpWn
b8Q6h7TaOyGNkOO3NDcOQ9WtC0R6rnTn4YTACVXwGhn2COs6fa1khIuALWuOtj1e8Nq3WtuJ77kb
2fuulHQToSHUyRsxUw78bl2/41adXBoxfvqdMUacOBtmKFoIvZ/aqWbB6rOJkyyIIkgQw/q35nbR
JDqS8nDezoOmOOkfGnfQYuS5eOp3LD5u6M9SVOJeU2EyRxTgRkj/i6tQEzN1o7uWoAFZoZrRq5sA
zZiDuBUwMUyvmnXWX7FLV9qB586csP0eWw33PeylaI9bJiMeeWndQqechxKaq2m1WPGFT/yC936z
ZJD9hjETuVU21IyOYXhs5sBGidZ9JMoyHHN8fkJNnQ4aQG8h/4l4TPBIFHza744NYzyuJfKLCWD1
px92vV6d5jfrwv83t+0RyHyF7byhiWjgaHld+XsJkKY/3ODjkLFukXi49s9yeKJTVa+q7zOw2cPJ
oCItGE22TSOS5HSc3SmJxI9hZ2ynVcr1+FOK/3ft3dOqLrWHxA+wZrHpJETaFKirls3opDsC8MNJ
ibvFjlFpI5snIK0jTrjGfC/P2AnLDq0K+bvOaKlVRbc0X66YLHTRgKxOsLS1howm1epzg4OtZZZM
2QNGg6EsbgylTroyKc/nwSLZZBXXiMfFAIJFriMFoUZfH8i+UXbPBukSY9mvk6sUvaOSK4M6gprX
aHrC5N+poHBSG3IcqjY9Hv/78yB2cLwPGVGmrBgtPNQmPLq9vOWwUk2lGkcIOzFsmCSySn9A8aDk
ZvLKLYSy+781b7lYhu5AG7tj1HpRe2c7ieKh3333ti3zxHiSjb4YPaVy3JJgHDxKIh2gVzhrdUWx
lzP3TOxW/xm1PyJ0ej3T+gJgQKzJKNNA/IyrD2fKUE1+Cdw3LZL38QQpfVM+/iskqpvQV/vQRhOf
sggm8RW+kIufOkqI05cN39ounqvsyWsrTWTcPfimvLT4J60Qw3YUdDwiAmGEBta6L9z1TO5fstI6
xvwI25eMY3cHZTIrd0gdeWETVtaqGPxGMlOVyMbvjd/kykrCAUsHLgzpgxCZ3OIzLdz3ThKyGjoI
feKWJ9+zJJCyS1MlbL48GmYxQGP0/8n0qBQpsifUUwB15Rff3FqxjhRM8p6rpXAjXSinIDxLj7Oe
xMnSyOagwloLnaE/s6WEqTgnq8xJaRyG/lCpOXUBXne7jD18jXWnZ5v0i9We1yaDbXvS3NlKM3W/
N6gWOBvv6S2pyZaLR+ltvUokmrl5aK9yRohNhPNsXFEwfggnRsFa1/KsfApMKPResnm82HzC0GNS
TnlK9xt9XwaN7BhpM9lZXnVmgUgKMcj4PWZhUjevvEAw0Lq5v6YwaksPx4n/P/q1yRxwoumQBsgg
sYFE6dCJ21WT7eCb2U7ZeN+FQegMLp+PKWG5lQtRTNHcc7TyfHKg0kWzHGdW4j+V15n8fGUf9GNF
OqPbDF4FFNZtm5FhBnYi3ePu8q2ioFZRfyKwNadKFhZtHdUlJG6fJavAZ89H6y2eCvS7Epb49G7S
EurB5whyFopLCYfzI+Ljt8bOk5DhjqoRdVSzP9bg807JL+xIhVnZPtg0oLlSOHkxFqFIHndYhcEs
ibXgHzhKkghWBzaaEntFqF18HaPsVI7YC5k6iWmTSxE+2IEJYV76QkqXRA1EFtXQ2b1KniS0d9BH
SSQz7k2E3O2XMjxX0DIr8dgG1Td7sXoLuqOwHqmf6ltI2ovAC0jF396PiJdkQMijWIO1BPvZXhlB
3j7JzU1ooSL4iYt2SvHtZgLZU7qXaJBQaxSgjWzLuax5rLoOMkXwtJ/6QDGiLCsIDg1J0zNW0ia5
7ubZi8jvoBburQluFryHWrrQVNL/rFonhhO9X2GRnis71ixYOROJc1sIRDHDKYN0xZijnkZMHvO8
xJshoREYccCf4FRyFfw1eJ7xp7NO5FIwu4RmbRvKOPoMkCD7YaK+8Vmw6rJ6P3hNWM+oWKIZ6QTZ
0bm9AkCZOS/5Ec3r21IA2LaAWKnl1mGntHtfc5CMR86OYbpnMi6wL9GmYRdfFLJbDhTICo0Hgcd0
reen978ZANK2sCVpEOPLkJPRPhcKQSS/6vZVOyQAl++PX9nrBVLS+yR68gA/X6AlugqB2FmXa+tK
/v/sFNWZpUUR5xIlMQ2uugScm+JbU3rUm43/20CqjPQgiXzLsR3ksio5GsadtBfrYyip9X0xdqlG
TtyaNAbdMPmrwm3GmEqHHvfa//8AErY6TV7ZRipfnbZHTXH4/pypgbNwvodBrVpwkriap0jFd1I8
P4atnZndeU07pHoVx2yGPtf61wYOWdn2sllgw5p0eD7Zl6v0iRuqF/Tiz4xJUFwJDbgzye8l5j1K
KeV90ncSpbNbSQXaadDZFQzt+ZcLRwcVoOguYg/Q7yir5uizmJwgYLlrmSNnBe7cBZvYIYQ2dcfF
ZRx9gbw7RCD9/4p0w/cGkk7kvYiLC07Evy+PLFU7TywE4l5pTvJnJHelxRwYEGcVW963rIW93/5I
+fKqS7rHfjswzAD+FsALjF1knh4/z4eVOfjurn4hga3eWn/eV8SPuoCMVQKueMCJK1J5OD7NU96U
C0CQ0eYPHvV8irj+uee3DlfLCWHwgRtDCrPacYOmqDn918gLKhWaAquJ2r9utfWszmBjC/mEUfK3
QiYvLVBl6YIWtwjYeSxlZi9LzOXnTXYgDUreM+H8bdB+WxKv/AMF9Vp/ma7R8SNCJjs7gyP3kVP+
kdrSj4wL0bYK666YRiXJkBlkODM3Mp0v8kNAC9uF4p6/lShimyvzH7N47s3j7QbLQS3VdWIeHnMG
h5bg74I6CHmSNQqDRaquqeKrCvVXBpM2eLR8okzLzgERoidLkMdHTvDCZgpus/wFhxyxaEB+Ev9A
gM6ucxVwr32SewViWsbYjTPb0D3oBH+w5ABnvxblPECCW/V7a6ZUfQMKsIc58o7rDuIYzf9jBpuv
tCe+eBgWnTTNawdCMtBMHD5zT96WvAzvt7LAXaV0RNKsGyOO1AwHQh/kFtgAM9QexKvIRS+nde1S
PzMbVJVOjvKMAGEPBcszqsVjljU+UVbkC5YhVyps8Nqi5nAzQx75OGKcfUFwyVeE76DuLI9M/+VO
EH9J80uxwOG8CwQ/GBccxaWKrObyUdTQCd2SE2HTMs310bqCXfDPKqo/Wcs0yBLRc/aKggL1pSZo
AgpyBCTCSyISs+Q4j0iSKxAx5E904GqCkGl25elmO3OqcNJXCmjcUZ42/5ANjDPf7HhPWpH96BLg
LpKT8fGjnXWlhVYVY/7tiUML5LGRGg7LlCJ8fwdyBrP+LAt0BPhBEzzSOsZpVEJZhAVVCeJkUUyD
JEEpT4uXJyn7S52D5z8hdpno+TOz8uUDurf0oD4MYDdnzKd0Ffpfu7KE02s4UVagxG8Z6KzyFFAH
RdQlsSJRPQvzUF/VtQjqVTue5rHAIkdSDU3GSZzeeiCsoo8RuDtVfetbRYqua87vG5Ew7P9qbsxK
/GqbmYeY0+BgYiVKXNeLKdwUwzbQBTCDV4R5YHI3FCvVF4m7TK54wbCCevphXcFA9QKhFod1MboO
W+Zfr58b/DhrGYFFybddqJSi+kNdysz/t1z5r//IC/AoZnSCcuS5TTXGcI/VxtO8jHK6IANWmWkr
dc3W3qppeFPdN0C0gZIkU7jXmW9gtuk8JbHABj+xrVbncvC84cae2ILikTG9QQf34TcrmTccrTAS
FYPXepHo4v9uSDfpIw8xLIG2Q57+5DJ5oY5HL9+94lwkACa+oPmoVVPvxfSbaQu6v8Y/Zhgvgjn8
6QO0zS6OFFJsz12R/cTcP2rF+wFTiTZrfSq45srK4EzgnWegG1Z6YAFLDEp+maBX+vdXC7WUCpyt
LH3+9pc+tyo8N1opJCNLdCpuc+s8boZx6/9QzlQr4UgHtZFjiK2+njiWbgCTK5pmUthruoFnO80G
rt2mD10jw6h3GVabhS0P4Xbxax9VD4kL0Wwa0IRhntxjMq8DOCNyqneH3ESbEcgJ0yQewyuugnSB
Zifl+TUyL0uYKGRFhe0VR496UCbqm+j5h2QAgb8BiKVoCQ+uO6KSzswdSvOhAv4TTjjXRTCQvMDC
9Cw2HAX5ClMbAUDCU6g37+oTm5+/vN6pfQndPcC03SxTx0ii8DyKHKO/per1pXgQ3crDVQc9KbWe
Art3ksI7UX9OcZD/7e6GPUbl8osZ4XaFFUuDgKvqOc4lNd6JqOmFWBR6Z9Bllyin45YkYuXaLV70
P2VoipXhKfoC2OYvulffDyibTfsfX6k/8Rl+RZiAqge1cCSsEKRCuAio8MfDuTXCyG7BlTkPhHXX
dcYYap2cwqN6pVFlxLp0cEfFIG6I/lhdOd/I2wapISQmDIYGMRjEd0wU26zuk6jiXydrdQUSCZS/
ycwOhDe/KFnczYnS7PDHlrL1aFkThNM4atbJultjhJiY2XtX1EE2c3Mn69aPLflkh+Q0GT12PYfY
LJRyx8aB+cIQhZSVHju9wTtASeI0z1bKVV1D6YtSnO/VD7yBRtIjRC03TLcD+EtQSGCjFpwd9roR
mGzEcDOxPOqf0lq10JeDyjyMa92RLeyTBzGGss3c73giZWTPL3U8Z9bjwf7QlZBfpIlDYw+DedCn
/TT0S99yoAJG4+VF9Y0gOi7EZ4i+tMlMwCcNR8xDX0CbxgAa1tnawmINxHZbWDjxXyPiJtxaTn8I
EhyhcDFPpPU/cim0OyoYUxwPbARcS2W7S/qYXYYJ+wbjIiwGm/6cZvILwOVFIZnLJ91TDtwdus4R
wKt1kmcPrYEo1w9SnFkZoDIMTT96TFGvogDDaeyHmdfgcr1Fmv7Za0dvp/1TDyqWH2HPhbZX3pFe
OFghnf77qVl8KwuPhF2Uji8xL4itaq4BeutP/+xfDvfQ06mB1BY7nUGCU9ER3oxzf8QL0P3dXCcd
aRkbw2W6nCGwiGfwvi65uykHytNWTaXAvSnsFvsanTRcGtBKgPdkq3xw/3+tNNyK3ls86T7X2dEq
X2ga6rkIPbQ/4U30vAKukxpL1+xYp4S25pCjEbq/MX3xHsMhi6iZINjarE6qDui/16A20Q0z/yG1
ks+8qImsaXU2Ln37sM05Rr3peoqoX/ZGawA7HNW13Xtc6tFlOjKWurEkzGzNchiVKGuKcQfSHz1m
964weZMPgEs/qntPhtAkbSVANCdPXEH8al9gFBz7BWwrPM7ocvOoYp6YptulOVPnCvNRpYbKjou1
9Sh68c1RQRmkIFdwigFVVJ9Zsw+VIfrzih/yb6X6h5pKFTTPqBmWDGmPGkcwsJbs/TFM+k754zKR
LvQNMJVyG7PyMEVirxfQQOtJObp24Voz2M6utLIUoznitR0bMrawSpyvyFNJVFdRkT1Wc9Dtu/tp
gvCjBT4q91VenzhmFaPH+sb+CgUZY1hWEnhbXfdIFu44+EP0cSL93tdisAYW4ElIUg2H5+a0PoIT
gqx3xMS7Ku0FectCI+UNU1+l0zVUD5UUvMjMBS1sfKsAy+aufJWlgp50S70VmdgUR8B/Nl3E/+vH
SAkWzUCFWGRScfKJI1phw05mDGk/9u6O4znk2Zl678cn74RXCk+AD/Cr1w3TKZADCMLgnY8uOURK
89JRYldQ8nObj+m2vrs4Qu+IQ5HuZHr1rJPtellNehj+plgwObjsA+0pNIWAzUOvCz/6DgA8fYyL
cHHgTSbDg1UZWQpqt9e+//t8U9efXvLkSwpxvqokFjHbFA/Bz5iUbee5eUy7Izn93UjKZciI5ZZ6
UBCBVQdAgvKbDOjHVpRiT+BUrlZxy3m5W+YiQ1qWxR5qEexomP57CnjCCz9mqTqAFpDcQEhI1YSv
shlbRnUFzh4WFdQ8ZiXB8QweROicfcyxoWlaV+OtXN4eVaSXhsbQudIBcAnRQ/Mkhq+61wnWzS5J
09wDSsBSOMjGYTMwuR9JUxhiuB7g3PoM7KLAHzTiiSd44IwzL3htKeaovbHDK9k+u+OwUyA3o/du
JcCQAmiltUg3IDcShs4w7ACDcDRu120TtPgEpHdg9/IaLqjP6cyYFVp2aSGS0mXjfOusbHfMKW00
R8L/1zGM6ULwUpr3pSHHxH8a3T+AzwMdz8XJaI6hgTsI36tsvpr4DkjdaWRJFHM/gs6rGandpd/9
T75nQAwqOB1iqvB754u/jqbrB3pP4QeB/6nRtcJ5E2lJfdxtEcocr7a0PW+UCD1btmUU33orl9dL
Iinssbqa6absKgo6EoXrC9qMmxa7zkhFrwmLVYvERcKjoNc8R8RYTGwZICAIsBgHT46RHS+8ojvx
FRZIgMc7ItMhMD3SGQGMes8blujzwJGzsfDUyHs34EiMkUXLBdfHj2k/Dkv9EqoBma2ZJsaJi31Z
ss/MMyUVQX5Og4ADNCOi7Ua+p0zeoqJbfCCyZpU0ig3qdpgBaRZYOVWEZK8YlWJYo6wU7p9haf5w
Kqy/lUBjzezsgH322ub23P647aUqPDhjkK9TgFT3pgPICNOrYKFmpdmEwkO8KJLkU8OFzkg42fVv
XoYdMsUWgzVDhrasVbLnkoQsA5VAbSZbi+llq8rJ0AeoYFR9em1QZXRpNVWHnC+LJ2lCsfySbvFm
PVq8pugV/hH37ISM4ZXiLXmhdILfYUPF6R8pCFjC3TFkBS8QOgwDSHjNFLDyULniMiBAi/4XTXMI
sjOmbMFP6CxYqs+ozZpVAumh1GSA2cKoL+4sZtQOPAOiwqvPZGsYnOA7yRR3ZkH1AyB4s0GG0nTb
WjZIzefWhPiGIFs9TKjjulblv6gBkAOHyPpVFD+wPy7RQiQBM923v54lXsTKUBBQ5KRluKJOZp8w
+58+U2dX9tYskiiMk07TsVLDn5Zur7wFx+SLJQWrmUoAIv0Qazcfp2hfCaXxnlISiSypNsg3Io27
4KfDWD+IDbwYcEOfD9gk5K8g4g/crQYAvDD4g/uzOFBKeS9L4uNlMHxAn2HWRZ+npfMlRadpfyzy
EYiNIkQhNcsCTg6dKbQO4ZjYTiqCi89+Mb5m7ocr3ArNotec2iOGOVu7squOeI/l6H37Xy0qgkHp
najMHLBk1ksTB+6X45I8tJXvHuIo5es2PkSTLjZ53Ojn2nyE8ZXRIPYzg/D3mbF5xgGZQ3ihUpcY
ZZ5Sqqj/qJweH521xCeaKyhv+EWQCGYpirpuPQdnuHRGlIf0yfW1F6yAoV4grRB+EwT7bHBPQCdD
r1n0InJWFTBwBox84F0hgSDhP5FtHLih4WLkoxbG5U+XJQYxBlG5qICAQMP0VfVsUenNzs1ICAJD
vbRGurJIXadna6ESHQEUt9Lcuezt0MZ874GC8wXI/zKv1qNh/n+qggTylRtCBt4c2EZX00/FsKqA
dlNx58YmV7ikzg+MrGbc4DDwO7U4iGFwRPQH1UQt5hnbM+oc1vc3atlqJTNEdmfWrMR5OeLItKdo
2J/ufxtMMr9nmOyw4GujARc+JYVjza0QsIeyuz+0JHRkldz7smWtLa4VCoL1xH+p0ajiwLOqNHee
MRowSg1txcmwhfx3517Lvlm9NIn4bfKug5n1iyK7CneNwspvA8zTOLZsU6cIGAm0oDUTY1kNhqqA
cn6MJ45SGrRiEc/IIKeeBwOpzArU1TVq+ele+Gqk5rKGUGSP3ycUMn4E15zD4mTTGviySTj9eoQe
/VgfzrsPto1Y4qpP1Yrhqpbi9JCE4l5oNpFLx3NUfOsd3bJC7R6SLVRpfUKbP+zVitvzwi0sO1XO
GZ6noYAPkOL9Ax7/4WVDckSxoyU3QfM6uyZAtrfQpWtS78Fq254X6nWKN00Yvzn8XTDJhY3Pg4a5
aCZOHa4x+Yz0nm0Ey5pi34xDOxykfUdrtctXDHXVQftMQauglwcJbaZzpm33c1aBAKdHREmW8FQN
CaK2pq69R/HSMzdcD6HHC02IFL5OXjDFa8lLYKRWlMjxiwIAm58I9IeitCte6oXR6HrSC95eG06Q
PbRG5wFjrtgRt/idTkTHaDyNjdEGXBvG2t8/PBH0e7lVgSQR1z4p2MwZMk/xVdXNDhBo6Rsiwzcr
EF8Z3014muBzUL/Ow2ToPQVdxLl0UKMK69/6hJio3f6mkzLQiKgpkJURn7L+u1AqSK4BIWpuWTak
fzzFpfxprfG4OqprOP45rHkhbk60b8UMh7hYvaLC3dYLorPkmgjMEYbcMSyc5R45ybOl6jFqxmfl
Igkz54u19fTIGwJDA3l4s+r+5VTYHpBbYHnvPA3QotrVaQyOJYu5rBsKtJ0yW2mvBAxtgFI5EwXg
MX1xGk/PO0MVae0CMYEJ/eiQP4YLGIJa5zYf2iezt4WnVSzYeKqxOiHU3Wa/nCjxb52Ka0c5EPMy
6VBn+pySVmnvHlMov7RA8/UdxVA7BvthYH133MBCaHYT62UiD9tt3Q2nD1p9M5rrk2Pt3kD6+M+V
C1575BwbuEqQqSEIrRHJqePMxOKSN7n8uv4H7g38CLcO5FTBP6PizFRUE+yxA4KdUbgoc4320PLP
J8y2t92ndqOJJs+ZMLfi8Cse7muhZ3kUoQn09kkwhq+iYBAcJi70C9UiME7g+QMCKXWKkC8diuKe
XSGoYq9erbQSlxfRwt8AKbb2iAq/JvQRAwBF05jAwsIHorYazGvdi8jOfAmJ0ezeVENv4XNBYAvq
LHOYQI2a/q7TUCBe50uQG3FHOgDt3buKk8OQC88b/YQT5y6pQ3dGOGVbvKr7Y0WCpwmJn9PMaTqJ
7R9X7QfKcjO4ARC8ZUeMKAhF+lDyAsRNjP3qL8dWPW19pK78/iUrWxQ1FV4UaeQaPcHKxBkVznry
MFRTv0CxuZB5kajNJLmKUdHk7q55szKR60R4sAYuAU4OhZKYvGX4F16rqmJGbSP5ZYOxIbWpqSNJ
bZTL/b/gBWCILZ9VD6NClwd9uyIfnxDHmYBBb7Qib87AYU+GrgTiwi3xeE94o4D1VS8+AMZ6Sxzf
tgrBv4+S32TY98KeEgGJRcyjyzgoAh7DIB3xvuUewL94mG97KYxeuida5DXMQkym2XB0HLvwNHEk
FfFijXvge1OpEhRpVp0IifplLUKxquTJOby77Z8OsJGWhFFzMqCpb5i8HlOJYWKSCwtPEgwU1OUF
kJm7S416faMYEt1D6dOY48HnrZ6V1R/lSUm6eS8W+H7dfzXqqkrFbtjZbf4fQyjDOpxz5iJo4vVg
7/1P31iy+zYHiUpKk+1J0tc9PTCA5SFVihEkaPt1LR1JjRksn79RauK5vC2iLRleiCdoQBjPU1xM
Np6Njmf0Ky1BCYdh6ZXbHU0wneT2qJM/wg4Jwi+MbmNKipEGfEgt5qLrT3d1I0v3NWcgvZ/9YWGC
rItgIhMY1X2aOIoy6331JrZlnIkUwjRgTPYBvnSb2cJT8sHSnvbsHTb6nc2ojg0d+hf4fSuxhCjP
w3BwEYhMTTA5jtMDjoJ8zGr6vSr7yYGpBKj7flHf7Jadh9G9DpE69I8/5KA2XhravjEuchM5V95x
Bmw7VqeSvP9c8Ijf6hxXok+YRQEhLNQdGuw8DCmcflG4P9wxnYdUg94HOcrh+3jNmemz1W6sdPXi
kVwsyMFUk+3NinZC2ELYa7lfsOwO2lSykrpDwhpZ02XVSuASssAZWBsd0ANKNVBG2tE7d65TIfDp
T63wGJ1vHxl5HbRIIWvVQg5G6pS28v5djGN9RWQYYqDiwv9KKCGR9uWDk+2A+zrtAmLMCZQGRqmW
A36tGXa+JMv6B20ki1b9rncW/ZIW+Bh4MgVJrBXWRjdt4NbryJsxe+XhwnCTHgVQsjjyRDyN14bn
PNcJI6GjyTmaJzK4kdPXcYRA+wCf0MMiO22Zb7lMzF7xh3smdlXCv5n6xM2oxxSOLsjwNb3zbWea
52RCGoPTDUtF6ngy7AGSB00gWy6Q72jbwlZqmyWA4nnfQruRdJmdyAxIsSS1o1B2BwHIACDfAKkr
bn4O3tvnqlnZZ2Xur7/TL2C8Jou2grlrExBZN55HtJkc4wCMAPxJi0W3vhlcWS9G817DSo6YkgMR
eLu0+uppm296n0nO0Uvu5wOBSqdXxaeAArkERxw3C6j+5BiDbMg2G20RLRHa4/7qzp2O4WQjlLP3
T6EjBZFpSN26MEga8/2T1OAWssQKJiWNjG3cwzN8ytsedYy6E7larHzTLON9F9PPIolMWtccxw6d
YDB7PvmWjfe7S9lcTlYvNj8NLNDgqgeYg53ua7Tt54n1k7nzF6IAMGllXol45zwGnxJ2qqINVo1E
mH4jhsLwNwEwoI5EPG4+b9LtUESS4Lo5N3RhqQxi+tejQel4OHL1qTJqPNqJrNE9S0L/8CfE8Z8P
WP9tc6k9ys/z+3x06HaI0ZZ6wRZ3nbWLeqKllsJ4rQT2of7vaFrWS0Vb6Zpz8GxiFXs1JKFq+iaY
X/jAD7Oc9Bh+uhrGDrEPyvS+NVVnbsy+e532Gl2dNl7AUQ32Zy+ENVPUNjnicWZJ3aZ/ODVnbkFh
8ELudmvR30Ih8t9Mx8vL6xsqQosIPAOYYUeA+6H6n1V198yI6Y3y82qk68hqQRdNcCEQKuDAPuhy
RR1FlYWkKmCwLew5DjN0AWczWJTmsfVVkXi7T425JeSNEbSO4zYOi0oGnQ/f4xE4f5NPq5wvvBdA
VggUSifAoqq7yaRpctWxPoBEBIhNebV4KStYazQTF8Rf/htkuVgQ1eq+gIrP2pprFfFvnjYbJH/1
XPM2lAE9tNQhGibcblYgxwt2Bj5/r7bfO2J9sSuoXFPBl4T2MqfaQ3J6YWLuL1B6hLYRB9UXdjsQ
hurf/Dmo7OqDJAG2ggU8LKy9PcPvrYJZvc2ziWy/USco0Gp9Zq9SWsYV7dSUeq8L15psADU8oqu6
ZrkXeMx1JOXVu+m6+8FMdWXoV9Cin302N5pmeo7ljXYN5zNBrSLq2wWlMfW+4YIp9qoy4BO1/6pd
AOmhZAlxg8vQvM6BBOP0vVuJ2kdYxs4hLEkz851VDxwNGFwRXySAi0fBGvrFGn9TTKBLgGSTSqUI
B2lbg8Oasbcqd2nSvD0X0BG2uJzTcT7MqC5kMrJ8melq7Js9PRa+OGNi+wpBAtACc6bMVpeGt+9A
wkLit+wGZsahFbc3609rq701THsEekKd/roe82ZTQ0rBtod+iSRgADx6cb7ScvEJKQBwv6XIajji
8fa4DifKVC57YVedaGIhSxb0LQNSWeaUBDvIhuEb2ccHNLEdl5nlCFG8gzuWEu33+BOAqd4LuLwC
kbcdnyKhSuMilXXPrTOlV7TW5mpqiZlYTTgkOOWjeQKqfwrRJh02xVIHN3nDTi8GfCIMTj2mp8Jr
WUp6ZGTk12HA4aXdKqz/A9n0AZwws59PH93w/1ZTjQZOzkRtHbaQy1YfIMh/W7uaZfwQQA8Y/NSP
doImaWwm1q55Zv9PDVbDZxCD94nLDNlOH/Xa/HF7TvDs4ABqlZ2K/+FIf3o9AB2P7XxbA2kJCGa4
MPlXXFG9kzRu1FJp7tIdu1sYFMpqQGijUCXFGkKuLCAjvkMsrRN4xGlr9Ni5mb4j2fcE1lPGdc+/
wgkgsTW+rRM8MonzI0nLrxD27o0Q4Gwty86/5bSLrnLccWg50u7jU3kdLj+/sRAImM8t05zm0U+N
KhHuruX8SbcvggPypQu6aJcdBOrFSC+bM+WHUdnJtSjh2PrkWneqyOmXTM3OHoXRqfFrRBd/PLzH
fHZ6ycEl8y6s+yiCII5iXIIOrq24RbWA20morshQ8iWTdrO0I6E6aEHr/WcA1uW8Ql6XZUDe6lSR
eW3WoIBtNWMhLgDDrAh5of9VoM3u0rOPRmMQp9G9ovA+8PEkpWv6MQRV9gNRL4cJCvOwpUTj1+9J
gMoHDwjHt797TYtqXsGJxFLEHmDnS4yWPphxA5pPHXEjjzpkktZ5+WJ9H+4lQOM6ZWeZ0qh0Ut41
+JiKtxPJs6Ru+i6D3PbxSndWCahZPoElP2CXHBDdQYBw37gLB67Adw1qgVCNjT+7pUAs141bUN/D
i2x17/TANQzgfvqpQZ/TXSJUViKx+gRO7qvgs4m/nJ1bA4MlP+f3LN8EfjQUkdhxLib2KQ2CJ0Xj
bdwDL5AVRHJBkPY91A4OI0FUld7JMmtbgMs3D0lA09kls31alGj+urZ0dDgTsTc1AlgsjBUPkRVw
w5j+3d/GhXFZPgR82iLHRuKdhlyG4t58bKBzMo4fAnv5YIZ7lAoymsb/tN04Ogai7qsbOL8Os46P
14SF+SgrcgQhZVydeTj9C08gqP1CxonH5xwTjX5JHmy2zrC1bRycWGLAJYHlHYv44VXZEcG5VLai
8fI52acb4KylR8pv09DvdZI0MQk3RGlSmffsgmk9rEDySjoPOt0eqIXIt3SkRg9tm3O+HXe+c9Rz
4s0vo0N/SS7Sb6Oum+1vLUA0Nzmnxy3WeKdvk8XB9taq2usdBL+naiSsC+6MHCPNMD+6kg/ZG64U
qaEc6kFgTIk9KDpcDzHk9cwO/ydx+qlHtcXXdsfkxv8Er67B4V+58BSBZWAsINYRkdYWLdQ28Omt
oGvQi7II3ODEJJPMhMLsikxNDM8vtVIcg2wEj6ZjuaVuDBua01h2NiFBLuM8j3UHojRND6Okic3j
9HoqzZtrakG5uuuQ2NTAOBJje8nrgSqiVtt1v6A1+m1Qd5N8gt2IN6WUyIyWm8CqlS16y3d28sPP
xnF9EUxycBmn7VkK76rBdS01wlu1LQkhfN5nIxLH+8tu6ckWW5C+S+vZZjEaSY8FYsacJ+i/K3ZN
YRB40tmi8CamnbFR3EK5yUmgeMjpL9yOhDrhMyEUJOiZ3MbgodHfdBvj3Iw7DhpLkLQlzFjQ75oh
uP/uGIxd+6c3bP3lEajcV4obzKPRmiVvLlOLuphPQnXUahujRc6vsFMd8A0mSXrLk1Kmn8rlyIIN
wPMlqMtU7ltH8yOXm60RsXh+mAPFrSC7BZ/osFBIn/+WuuMsubg1rjBemLpxmz5wkUxPPt+lQM2F
qDMRwsR2wQHws46JZ0ePwH25Pqkk6gD2Rnal5ZXt7lJGv/4qTp+FBGRblnJALsj0LOSW4R136R36
KfGu0oRaOGyDbWC3SkprLqlye1wPCvF9oB5d4DmUTh84sO8csOW8hA/KTrZjs3e5yWzv3OLFMG21
VutY9o/Uh9Q3mYUlmvYTg/PL07DH85Fr1tY8XfGQ2bkBj1Y4RnC7/hil66EWZ1OoOSmJFkDpO+HS
HRNDyd30FOzsjQte7bfMkVanG9eupTLoNs0Pd69kFDz3Ht0YNw6msC1gkIt3IVyZNWEZg34aZ8+b
bvaAgco5fJGTskUrjgHt3Vu18HTnkn/NVOabupULLkizG/gviMS4RfZNEguyb8KFQ8xZHF7Wuz09
u61IyeQx8EXekbx3ZoJ6WAnQJEfUuJ2PtePyjJ0Bvd7lcZLVkzWuzGC3GJNRuFI9viCzM7vjB9Cb
xsCeH6/fsdUmJfEstsY2gu1oBuJsYf/8VkAbgP1hpJoVip54qD630KMDCcK7DIvl5NmJ0vsB1BZ3
6vqRLpVd1LMS7mFCadGvIuvEE3uekDmLcs+ggi/QwzbvOawol8Bz3oW7x/pk2H+VwQb+O7pL6HGU
31UhrzUM+5ALng+m9VmTy0CjOuaCaQZYOeGAY3i9bpZ2E0OHDW0ntQsDVWzvNRvhYexrtAF5/on7
d3OObaNG0hiTyjdoPgw20aSfDf3zWgdEnCrxK2x7Qs3fj08msIf19O5e5nuR6pi1+O3XeR2lAUJY
O703mWQthJfGOFhEr4p76CD+nxkisCwncEFXOO0ZtlmLslj7hSLNh4dRX/4lrjMh02wQlVzZlKuS
PIvG7H4IBUM5eF9HW+lednmznax5/DcmnTeRDBryhgloViv317a4eMI+EoS11aM2gyBRMrBibnLw
TOc/tdYtVT8S7MPWO80nCdrS77/dwVBEBmGEQryrnFbOlrVIcq4cqR/WOC5CMhjEOf5D871R5q6Y
hWNZQC9ju/Go0Q+UJMWkERNkoSWCxXR+UlksCo5FnCmZccsJaApXi8OatzLpIwp2+jR8KgLOYZwQ
giLlPF/qXMXthZOz3O3L5kjiXs5OGBvMxfL8MXqwdI35cWtpfPpibfYf1KQFzKUyddKNmI5jRSP0
Aev0/r2xV4IpDGPISl/s7i5HeBYJ1ZqWvybmUUikFkdhu1ZN9szJIdbRE63BbUWhI6TntbdIJRG5
vQxgL2rx2mRs+n1Xnb12g1Rm9cIfBg3clQPxcTZx/o9Vgyfken6Dk3B5jyj9QG6LHXW1eMIvxcmK
GFPX/xhsbO6KAJig8otY8CpL9zCUrgtbc+xyxQplcPl0egRYXHo4eltmbuTqCtlQPR6hgXNglBKo
c9heARhOwA2M1MKYRP49my2QTedF+WSaRgFtG9zDYX0KbyObUJauGccuZy/3CRhTH5svxZpRZNxe
q0salN4L49Qu88P+z9d0lb5UZ7pvsH974u7F7Bngy0JkeW/PcstWlW1cYdtNcKZ9POxVf0qiMOMw
3XABoxU4z0YMGogcfp1BW/zvqyHoCaH6YhcgG1gI08/UiJ/08cPGGsf40ACrZgzGWaC7d9bc4+b9
2OjsHVS/LVGgkrrRJo2YJBXMduo8loF36l7JWK1G/m/BVk+Du3MtF0aSF4Oe5M7qsHi2rD9yUR7r
2KUPaQjaimbsBxxqHLdSWYC0/R0/NUCCkignd3aX21Nh1Ye3IzwDi0TZSvTRg64xmUqs7cnHBiMD
KVrTvTmmJHlJAX02mB4RH+xKNK0ZASMSIzKaS3dbJe7vsUhrcSOSheyhJD/iKoAw3lC80LGBtzbH
rifmD6+OiZEJz4n2gOIuZnhjJy7+nF0Jp/bTVjXCqm65Lr1e1/MWH/Rwrl97lr+Flh6J8Uifju3+
iuwYJ4T6ftcQ4olMbL89T6Zolafnk936tB3dbInYJP9Cakju1X1IuE4kYZ70zpm5ZbFFrx/JQp8C
fF31oeAnE5pIh3QDoQNCmIGMvujXy9y96GUPbvrmT2GgATfoI5kkOs3ihx7Gpt5csl9CRPT1GLzb
aoCO2Cax/bMAjULGUU7oaU+KZ0YW2z+pxWm4p21k5SGF9cLXEI2Lf1xfpFtNj8zbf/mGQ+BXHwr6
8eTCjcHWLx6gUqnx16zbxYUxVmx8335Z4thdiFJkGH6pgNJj1PlKonpTMDPNAPJp86VEYht60O9T
x4ED5/+OaEbyxZ+6HzQO8uzazln9H/+argbkvzmjydOA9KjcujNUrkniAEiHcRG07nYIbEIk0kyS
CYi26dDVFtEbUhjmv+RbudPjGlGDR46ycOEv3PzzBw/jfKoXtvH2TKaRVgbvroiq/AVetGCBJ4XU
MQ02SldyHnzaooSV/7QejiRdomltQh8VF4pwuLeCrJUVW27rWkPe0Avuv1GCi7zqG35Ol0rx40Qw
D7MmAi6WIIGsaaqOTj/d2PP+NjxUEE6W7yi15zuaNI31pK+2EvT9InNv2l4UtX598KYPUAoD3ZBJ
+m4b7Rk2dzWo2TQv0BwQbTtQZXZnT7xYBMTrsHmzZmYKzmVWTWApHCAIvFCtTuS0BJLnLbjXj7RN
rc0Ypk3l5bMePPi8dPE9oejjbPTKdLTuJ0R65Y/WTSStXQmrRKoeQR56TDblnFqX4ncdE+lUwppx
zkcl0934Ro/Fi+15KvpYEoFV9A3fXXP70op/uM87yZCwEpwoqQZ4HwvvC/oczyjI4EoHUWEGHPLF
+1fnCHgko/Up53UwpW6mclEyL+CBxbYFOdrG7rI8ZZLWsIgEBSeRp0bIojsFZ+Fql/tnx1oZUprz
K+Y2HYeEU2B7JtTQa9NAeWC3TofXitZv8QqNu81mg0MeETJjgmqjzbR7Srafmif9mvRWaX91+Crc
8RXd/CGAngXKrmbJ/GEch5fO0FMT+F2hwl6QV/OV9sXiEfxdZe5c3Ff9xXlhtxxnANUXKhs6mWtI
VyYr8rrJeKylz70mMjexJxvn1EYn/SFQ3RgC7z5BUw7n7equ/dhJEd+n6HZbTVL5IYmx2g5iInRM
fpdKnOQFsaKeaSK75xyaQpt0gRf/OZ5oQNT/ccWEeO98qoe1MiPHxgrrrGlnNOq43LzI0VCkZlSN
uDSEQS4l0To0t7OsKffPz+/rmMPJ/QPx1VxZGrJhlW4xlTueGujcyp61IF7n+IaLMpyvkdg0Bkn7
MypU1UNktnxd6e9CBb0IcVCkoLD46ewY8+KLfRjaWN50DVYeND6KvqNF0dzVctKKQLB+0SDgzHQn
LUFJwMbAKEBYkNDlg2786801nYaJeJD8NrghpEwKmbgQRqqqsnO1SQEXRc8YLSvfMyTcxUBnGIhF
tCDCSiAX1YZZK0mFEFplIc/Fyh0R1z+k6yVkanOUEF7uQqgsDnCagEFDtTzG/ieDLHgoaokISNYA
4Qb8UUWnG1gI0ksSVQE4xPaea1mRm+OYRmmBei7jC4oxbzX0ZgsKzv1JEgbWZ8a0cf67+xJUmRZN
UpMt/BxSfQ61/gvvil98iSnFrA8osAExCjbQClbFYpAJiEHSnKpZ/oTDVm3zFwlXrZbtkuGhF/fV
YXt1fousrQq5u3l2rcpOvSzISv0qIpAAGo13kvbco9+0308auwZ/lq+fvl4YN2LOhxnq+bdyC45e
5XGOB5VcogEUpP/Buarocn7UDa3mEVZqxrXb5Qr5UyQnKVcz0Lz08wyarSaEun1SIipkw7DC55MB
ASU3Yd6p+suHpn1xieFTSB5QBw+fgPd+LDMV8CczBFCgAn77iXsfeIhd3YgnRbD/6LeUQIOwWRhz
mz3qes5bSH14/dCmSdcqCcNcmec5qTn1KvGo0uqjWO7nnbMJAo4ZRLGmmCJx9rCJ2OXz1fTiUrUU
k16GjM5fqJClrMrdQAhDPobj5KKPsGJcv/95ySm5Xog9SR4I0tsoZRvQqLr1nFki2O9ve3vv1dcY
5qs9ihtbMiXrOWqKsGzSF5u6/n5PriceD41Iu3zS8t2Y1UdhNSFj5vcVWiDcX/pFoHM+gFEj9Rsf
8KRFW2wciX4ORcKLhXqMi3KPVDmvn9r/fbTtgT2fYSbGDV9o4+gh4ZUeY3VCAYzpUn2M8ijwfUoK
tfP4ZeuBZMDIfK25QeFKed7kR7bT3ODPUR7zN3vhHGnMHOPlcgXLg+ECXqG8CbDKFLKRt1MvD1JF
UhE2TbSpJBcrbyE6NVEU2CJdVpyhLPcXJQqQBg+3tUIqq1uo9A0vcaddi8nX6F8ytcUShJGQ3tRo
4+gt5X+fraSBk49/ydugvDKFAk+IDiv+cOVZIkF7ot6IYBxf719w33Knli8kXdXLMB2Pba7CkDpE
8zSa0yvBWHYXV106dmhjribU7whfMBV8ic8zZnP74b7LmcIqPmhAr3CSXXSXTyj9CusW2dAFGeee
eKrp7cXwwFKgNVbVOuIm3QB0VkwqmlRUW3jCU4Fy5KB8D7C5EcZWZGML0zG9VN9FNyNJaciGjnaR
qhbiwUG3PRi9TN9Kv0k8w78Zwl+1cMT0bxhq+GeuGjVdb0MS45BtzIB1VfXHMmhp8STNAQTfzuFh
PePq/AyTbP9ldZ4qZ1EkZyzGWraD0U+NV04sf0531ZOgskUfInDPiDiaF3N7nscf4EyH69zClchQ
6UE4LLMRWci+lE8cQI0t0dt71JGcL0yaSS7oO1TVaA4I4fnPXXACo8My25UKrtqmIEbvIf/3ikaX
71mXGRSeCTtaLgLrLlUjinuNXJsbVT6B/QDFwjiE6ZxdtMBNqy4qG/Unol3xncj2iAFi9vbuhK4n
qf1zet6fznJCno6zZ5632+js9jANKwhPSTCOKmsweeZKthiVhFqkmqadMy+a6PJBzqE6OOYaukE8
6qF/VxUXdg4JyPqWH4XVoDq61aEHCbwZgh7/xSMRyV0lFCAnbjKeMMBQTdTKtQiWfDUwZZ1GSGZE
BB3xPiW4aBtPbWcfYO+IlEwDGKsyz+YY2xFoblTzeryKVZoxIcjcEokDxkesDWBrP94rvCuoPMV9
s1o36+rM3qM4gY4A+HhDRQEnwQ63uhBmwcHjpYFqCzGS5+oEXC4G6IDEqFqKKSHGJEF9IhYkUK1G
P40xYobRiwSC/jrkW7um+KU/64StFpgHZzobOPcgToCHJSFewj0HDy07ZPflTVNm5pg7sr79d7Vb
J/IQ1qtU0nOi5A0j4fnnqFpn9UnPhwcqridsitjCM62K8Av3apAE4PT8+3Hqm/PXk1g7iKYgojHl
J65JXvlZ+54JlX5FhvJvSdziDtPQf8kutFpS5xWOdVBjYhQq4uyGATzFYsR/6cBntrv9fzq+AfaT
Ers3w+vatcQMl4LojcS0bUi+mBzNw0bblXu0Tle50r6HinDetRsXqvg5l+M8GlhIqLpVAC5TWnzB
akZQO/D9dbv/shJdTkLPl6QL38xHfM1/9YsdMZ5P3Gy7Fka6SDSDwlOSa2znkdPBNl7fbDzYBgJC
DKUZn81Gx/xAjh6tHfJ3gWsxxctd7/N3ZktxuqdVL/RME5s2vhkZdvyVXeFQwL0UTnCRZDvdsKIi
yCfj6Si80MkYV9RQ1KCouOy86HyVnlz32pUc8ZmmaIp5+1lX1wcD71DEWRAYXTHCzNU01pPuK+xt
TOGBQBt+tTt6XIQVbKFisHWLOmyyxY/ajHiaH1sCeVbBYH7S8NqveXY0p44AGVR1+XVEiZltiznN
mGOka75/I7nGQfx4WDvlcjROZbiHD/wCaRlJLzdyZvcGPXkeG9CXnASQgeRWErsM3BfmnWa+ZXxu
9e/QCppAl2OJHrvMDVL13NSTA3gQN1MgtTun97t0KQ+hFqo4oNly4OoPpB/ec8exr8uqRhwOLuWU
vvwYA0ihdT92W6cKj6P2FnRg4nNq8aXeDm+L0bI/7siKuB3d87aFvBDubLVPQf/BfbZUjxZwBD4M
oW86bV7I/+5ZWyi6pE8rNiabfnHRzpeDOC3XwZVIbtNZdH81lkTQoNz5MOurXVLHMuHuHSZZmVjP
yHz//HrWCqSdDRvhl6NxQxBCuBV72YgTiTUzMwSadG2E0ejWQAi8tcsAymTP6WI3KlSZgZEkcPxQ
G4OziIG6Pz7Xd5mO4OY7AdhUKU5CsmC+U6sz5fsx/nUdo3jcWjQJodGY2U4TgJWsfqaxazM0a0ed
KkEAXg+/Y4nMCXUgfHEo+Zcy8M5UD/eaCW+Vk82OIU5E6NGpVvFBBeuCUR9oWcnH6u/bNIYwQkD4
s3qBxxPd2SEvnEBXGUlfBKMwMpZOv4n6nyoJDE5bJNzBydrVBOLDvkhxv16UpmNq7COX68JlACQr
FX3DnVogCw6StsWDaF0DW+XXoDXXpmN3kQ4/5fJ01mJzjdD656K5yWMuPKOxYeJBg6hDsIMxtyMl
Kri9jNmTsZwMe0ALP60A6ldIk1E160RYVrd3Kp+ItcDDlESBioRZ55Qfg5LDYDKo+lSfY7v7jgau
IcxI74qgtSsX0oftfaB3Z4mpu+5czZRvVywsuRam83Hurdz+3SCfvLkWp01hoEmtA8YKy3X+WN0g
MlH3xllcIEhI9I+Je8aMSu1oXMSlHlmMLGO2YL/OEjQcMjbHVyeLy84WDCUezSGteKpQSjHSnVwu
EAipK8e3SxEc1rwrJn8+Ky0FXzQyiGboCmV+3RLzcIV9txKLrKAGK5GY9EnN7scksTJVx1cXDqk7
YJZ8r9DvW4WFOeqxeVuCnwZ8mnVPrdfSdpURjqWf76N/H4l76YNqOBTaAf6mnTbdu6+4kOTzrEEo
0v8CSGlD2JZPfvwoqQJhbFebQdMgAmUhSnw5nUw8r0pa7UVSJeQchw0zAfYtu/WlBdOnjZhdLIau
bkl+jesa0zA+9RKVWzk/l/3I4pfDqonJkGiPTq88Q0ZEoVDj5bgfCeE3NZo/TJanHCXiwaDJd2EH
hDCDSGUwem0uJgNCOfHDby/0uwZ3IL/2/V9ga5nwFNTFDAk1IOi1fTBmSwbq+6CDhqI/5CKsVd+K
IFZwkatTuSjlS4jqWjscCVS9pHb86NoMWM/cav8OzJ+3oNdP6QUigqqLfi7kZFDNnRaA94lrdYVh
w0BYdXi0Hab3JL2lJRqdLoryXnpBXVPGtMJCqKaLIsC+wKiRfLYTWCxZuhIgNGqhLE+ZuuzPvnw4
5cSueFELGzr+KrgVDpQW9SWTBd6wGAZ3+Tu8tl94CGEbCetppw2ZZhZYVarO7ap8zGbinbeO2nxj
xWLulYsTmCVqF45TV1HCkFc3praKU5inH9jbS3CYnfHpE4s/2ool4Li7u/Y2Rjv48neknHfauzA6
gh/T/DVGRwOymiGqbxqHtshaeL2VInETH9UTBCoVyR4aj4vnur9nOCeUG6Vt5xLyJvavU/Nb7xb/
Mt5hA6f3pStOUkwZfsIIsOzSHXnlVSIxm1HqkrKyMBYVYzkVfC8/oJHkP/ueabwNiV7nLhw/0Is4
H/yuZBJlgAAW68taFUj9/p0/G/pV+9R1D94zMjHDqJx0uYwLRcXXO40ZENGuaH6cM5pwi6Z30iyf
hdKl6Pi5kKi2Yd1N/6i3Gq2SR+ZKdBbZKips3uYeMz8uw/gpL2ewJDFlyIAn4Ok9kLGaYq5VGHI8
3STPTxzBCsAHkozeUubmmFucGHgSRxUZI/AJu29UCCftMVrRLlewsSOit3ypWWhn0nr09tinH41j
RoeKBe6LHCx0U/8K96eaY54rTAx/UdMmCAXk0DjSwrZfjA+1Tez1vpnhjv5dbrlqKYut+S/eqoG2
yHxxL5E9PXxsLngrzkop4JpRXDj9FDsGnaOow0ahuKprE2u1qYGhKHz2XfWhIv3qZHo4hfO+iPof
/6gXkxworShL/DeXvTePZ7+YtYZRi4y28IEzNtFu/MGmVRIjYW69DefeHvMMVC7A0lmFERUVKxv9
Z1SIyT+qZfNi5cKo1xkFGhGt3APcRJyPWHhIHqwiWzyaeS2iFjgWCGZqTyP0Vlxc/eqeatidIbuJ
gktm5k1EP/iDJnIBWccLo5Kze76KUcvJ8qU1Qb2nnoS/jelY99sTfyRqoQ8cGRGSr8U0vR1Ajvlu
nd8a39WvCxjQKwJtvToaDHPChxSwfcveivgfsTWJAenqNP1cNtZimAts/hVNe5kf4xB7wC8LyJ5t
eJB2VyiuAghSjmKXHeKYwy8NmF0ZE1+dfFaJG+ED3F3mgkP9/PFethAZHih1UKsKo5OEHA0wS3qh
wMuZbiwmjv5DlmZa6bKBZamLOgG1lJpjHDXlCrATm570j+lnUHknJC0pfx+BeKl4+0wiv5/qu9HN
dCbO+Qf4krqe7rnV4GLnAmbAdmy3dK6gi3J+3yHIoS8cdcwhSBGtDYNlrK+JE0RmOG1IDg7lx2rr
YlauzSCs/zO8MkNQooQIjxmlqQkW5OsvFI153qQ4j7ixpi9Q7sUOuDK6FigYyGJX0j3uWqnycnFP
BXZ2F4Qgk1Ssqnf/A+wlCfKPtssmKBRro2XH27sCoFKmB0KHpniXQhC89bIS3CEVhPyY1OcWFOHp
W5KSNkVwvAzJluiAbo2AHAi6REpBx67x0diqBp6C3nVHTWEB2RGBn8fV4nWCx0AdKTnSOU9CoCwZ
DEgVZbeLNPpQ5OFgh1b64FOgIIw5XwBbwJbqLKypOf35QeStSzZBSjbMTeRpejvAAkeBdibpqCGx
bOvgAwdhYfIj27l79e5RXWar5xPo4dbiJWKt3GGfqn7GLRU6skffV+fvUkm1HutxQpGwJiIJU2Lq
Xud9f6tJ6SqHnFhNC2raK2DsJlv+vHR0aKwDOHn/BcNoth6tNwfvjl0GdYCYZAnK+YGOjFhWC8Mv
WRa7O3b5zSRLk1bAWY78iVvbYRvA1+aAoG6EODfJvtoIFu2vSUg4KmFj+674r2N2PgrZvPvhPFzp
u7zM3PcRMUhBZLufiFIHUKOqn73C5RxMQ0x10OxH5YP1AsDYQ9EaP4F9TPPSCLWYbOyYLLlUWBYu
bEG8jgICVYCwUOhXoMx2J6sylI/Sm4z/g/+jA3HxDJnnOS2dNQESSAZNH4ddgs7kK+UM0VWD0awB
LpH5pkgP2pjMJfykQhJKYUekcC19lDccnlyS18YOuNScAzWRII2Hg7X/MYLYOeLMnO1+SAC2JvlL
6t2qOnP7oXAaANPNqCCRJm6IhLfbKLTmSJ2/VqiccVKwVZLyxw6MPF1qyCZscAqezRiXw6L/QsPB
Rot42fk4Z1rEX9rT7KeJjl001yOaqhylQBsLd2NJgkFN5DMPlCR99z/D1oReaitwfwVODc1vJjlK
tVKKFrR+Uv0S26BxpUSFotMBylMfp2Ye1n1EJr+gxrl2kwbylqkHR9A05vziagkB5C5wMDPd2tS+
WQsLki0+KPBqqXgp9KpWyv8rELe2boBD0LOQj8dIMYMkX0oKotcOrfq7KUP1dpcMZuxt3SU5dUSl
GwB4AxrG2V1c+OvnHr+9vNA0kFpw11TG/mgkWZ71mhiY72j0unSFz2qCkgjdKp6N4urNvutMX7Yv
gxPEvE+2YGd7/GkwbjqCeHT4FxJVHG+1soQUp+9FcewUAu8dW3VU/WuzNTfSAHTbDBHlTRxzk3lc
iAg/Cs5l2mYBZVHfTxODos2tihaHaR/C7JNGSIVU+MpzYtbyfJUz0Ot9jnCDQaZSkygL68eK5eJG
0goqZLZrrfMLquETAyNRW+cee7cnsRADIcgfHtHKcAoOErjEP1g3j1V7/9kfFReeIeRy5CrnUM9P
hQOkRSs4iWa0G3vzaC/+Mq1P72AfY94dNrctplQvBD6zIWFwzt6YnDblJXIa37TKRk7II8w9ajvA
VdyRlB+fPjcWNukgkyqsKZ+ivyNfkcpksHr6QYiYNpt9zv36Auo74ChINOnM/Ui3CApaWKNIcWQf
ZgUiKAfPXfzJ8xfh9E3yBNcaYL7gByBfIRc2qf14LpQIqhklSI6LZxAhObi9oWXC5PYflAxu4T9h
BOuN5dqf01INO2C+ovqYgrpP8+NmH7OJ1gBIdc4bs/FbJxTYWee2mWpYbRScqiL00X2EJejCY0QZ
zwbiRvUnxRW3DXpA+Wf/hb9c2ZE2/4mB3pn/jFSWaEsqZc+/gmB8uFDWUMQxYid9B4S/ZcYasLan
AQVXeXZsKVTI5tjFedyq0RRAhpBW9hsouegSJm/nGpmf8hNA4hGwJPumXGEsgwmKJbQaqT0UiLzS
XivfWhQfu15TR4yLNMdI84uemgww64GkQ8rhLTcQbpyhk5qHx8er/NOjDd0VYylxftPL/y27aSLF
MEoemGH+jvvWSgr8UTD+qEEZbpIapldXf9KuOxYMqluNj3RJdXfY1+FSd78gkeytPPfmTfxiCoIh
uADRBmi+Y7E2ckAtZzYxLxTZkXFUy3PLPinLzsE/hg3UxLduUUgwFTDdfmuw8ae8Ggfl4cUASPgB
VILif6Os/b13hd6Tbv8FX/dAZVAKh1wtp1r5kYZRgiOtzXUZXLWy8qmQuJaGoWXr6SrGbw274Wk4
IoTPJP8fC8TzIMryBd5rOj1o9pQ/5Liw6aKCtq36uAjy3VetqzroYc1p7QCFbbaU2X0bz2mdJ+eb
r7nZ6rI7PjGvDQaEpnV1ntoKN/dYql7vDjRJufW7ahMH5Gbtmay3QahIbzvnlbqb2ui6JlCs53zw
1H1NC51OXHR1c0ebKP2M785jAnaWP1eoGEAp45End4ru2asblRmDLh3t+3Z2HREGZ4DH7wXfpX5l
fP/VkHwET+kuSnEmRX57oZ8wpXJYqgMljw/NetCFme9q8lw9fnMU9vHr995OpDIxdXfR1pdKMygf
CqCjF42V1vGwroVODQnkIuNk8w/lizBjlZq5z+YVJbpXPEBxba6UhrXvYUNAaol5d7lAQhH8H+SV
JXpW+zwHyz6cDjww6EnG9UIakbymU1lwjbZ7bFiFPvkfcQbFOeQBARgg6lvbr8fHQM78CHDJnQoT
ybTbTYY9Wqen9594HzFKr6f2rX1qKJz55n0JjwcyiX3qGHmiD9sUje474gfqjTd2cFvBHPASfej7
hHo6ATk0D9wmCP4s4d25zMjwb7oOxhHl7kQn2csG0GPUTehpSQhJIFfXpO47vq+azA2kv2j18ZKd
hyDhPJftDyYpL+XfLBUcZI/U/8uABYGa/zyPkEZwIFTT9n4qHb8jfM+2N9CrbfhAentrNRTosFIo
SLf2MVDbwECp2ef8mBT5XnFNvRRWXaR/XERXmHhvUExZV6YytfShtqTfKoUprC0xCmqAI5DSshqR
zQtKEC51dwCrpwWo/BWaHwndYyn5aD0wA9GHJSzVVOp/NS7K++KnMaGkNZGYwjo4eosDCjSSsnVg
6mfTmyxl94bEDByWBaztThaTEC+A26za00SyTsPaaLJJUucY/5jsYOrnrajpB2BhTg8c3x9LS7ch
ZjLJiB5JEkENM4nR2Kty0PlzdfGhjqtbcuVWdykFBRaJhlHXyIrhLqzORLQVny2HyV/aTWGVWQ10
QR1zXwwrckKlCfEVQRc2LuwXRA91TmXcfifl8Sae0c0UoNfEgxUFSiYaYyUONcuEWgnvBzaSKg9M
t9f3F91QtG+EneukWYj7humGzem6ZIpgCtkcBTLYtsjLKexS+G/rauQoXSef2/VMM+STxRnA7RVh
qd8+H4LFmWHyWNhfC4VesbQW2cpMAL4uK0poIlkGT+mt3KGBfMcBBV3gba0s6jzV9xTV+VDt8pQn
y87l8ekrFTKK8KAtyuF5D2EnnwLH/fDL+Nrm1KLEg7OWuXPvvWN4Bm/IMZizj7e3amtkvoVaNNQa
3/4Co1PCAc3TwWHVRzFJ7Ata0IV/GQKJyXCJWKQNgcCunIaBUbf2eMtovnWrY6NpjKnxxtu2lGp8
2N4OrmUpzV7SeE8snjpZuGnBxY+/dMArJttjvC5uwmidO3R3bUHdPLh8cJlVF3sBfzx8VJewAoK0
+WOzImUXPgAfccBJ46kbxI0uSvLq46/pGqzyTiYQWRSLLd3NptHGG1CtZTgSXuZspHlddXseQGRe
0+JE11aJBp2hCSHs50ArwcoqmeA9lSTd6YkiTKRd0apleczMgvLGRvreN/eZnpV2Ug2R10YHc4FS
97mnJzPuKnLFIEsYyFK2bcnA4Q2xxGKQzPvHHv+jYclpPmkiWl1Eu3svoad/jukK6/NhgGdh/rH1
AXr+3ECVGOS3PQpkAG+pgXUB0g/P0YwdgZ+xUC7GFkX57t4rj+71eXzSMNDxltw8k9DQtC/E/3L6
Erk1OsKWsL48ZGkmXL2xhp0tT7UDi2M9OMBAhd/g/ehF5BG6LAYTxTA6a0EDCGUK45aiYSffYt9P
2dQl4P379rzhol52xY4r1OqyxtG/Tm7GhlUB1YX5gyRz/vCQMN8GUrWf49niDOnfp4Yd54HAc0RL
6JkQUHH5A4iz4RNTcsdd0bCvlE8O7hAppW5I5Ui5I+GZZjWba/+W5zbK3Y0bk7XVf2sKHzhsL6Sj
9xfP6p5JurfUotLVSatOrqq9UOrTXBmcGvAMugijEa83sXJvqZCSeoA+s6iOr0tQQ+EfhevxhAG1
zo78W02tNBSs+GGkGKy2F64a7jZRUwTf4FlzztzpQ+ZUg6FRfikRyg6WYjC7aLvQcdGlZTsbjus+
/aLDWqQhM6t+iG5MX9K09EB39jnE2Dr3PQYR19Js+xYtIrulmjK8/OhlBP9xjyAiCDceNxbJDizx
14j0+FUmQnsqhZxDUj9VpbZ6VGmRzmSfoxfJsE2EuvV2M/4yj2o4escwdPZY116YV3Gykrwp0lN9
8HCsVZC5Cfx1ShT8YImR7YxMI/EW0H+Z6aecauYEj55BzzJSoflXjCK/2GdUEsZDHkMyARikJlIl
MwT2n47dYPoFNZef5TW+pSv2TW1qHHJvH1mxNahkDk8HQRNAb1pNZI/ywYvhpt7LXWN005/n8xeR
Lea1buTb/8vxGsKGw7Nfz3C2fT8efsOV7p3PTLBCevpW0hCjO38Iv/YaovuNeWOgF1Wu4adDA3QE
s3eOgRFkm28qEfLoOFiNLGHMCEQbnRStz3voHM3txHAfErNDwjfKtfro7PrIy5K6G9ZrSaoa9G4F
4Wm89dV16rtrGoa3KDBUsKI9gaqN3jhfnrzdKUHTVfT3C384LKLL6vs9zdHJU93bJ3A69KkIeXI5
RuysQdJUzJnig3c1zP38NGcTKrfSuPcsYDelpJKZiZ84lxTbBxCJgyUkkIA+bT5ghEZ3zyXipGqz
8SXv4b4Hv38IEifO9o95Ozts/TvKfqrrBpj0uO8U7LkjKQ6C8R01VTBxWT2eXHZ5XQeXZ1fgyB1a
w3HOWxETjwzEyIwKG8RG3h54DGkCR69eycdavh3WV8RNgf8pzZ4Tgjbq+PfjMkn+Y4z22A9PTopm
oyeQqf6tuDK6587gcbxlic3LqxB9jckDTfYcdnB1i+98Hx2eI0bs1+WVFkN8IK6QN7SAdEU6hcDM
sKlGkF5N4Janz1bl6h6Vfpc7zSUNN+6exYXRml3b3tn8JAXnKTg82Zkeqs/w3yWTDje1Jfhl1oPE
zyhY1DUwlfLFdH91js8UEh8nLmaUPY490C2dkMBqjxay5bYFX/4MkO4+Oo0l8QMmt3Ej9Qa7/S7t
iromVi2ZOY4K5xeCI6AG4mrutg1j37QPnqiPFCE+A+hAeAbuzUXV/hHZ5YqhL2awaVv9ZKKVFyND
KZFT3nJmTrRtTUbAL5G0u/P4tzycl7iug4p3unHHdWIKkGNEncjVA6D4yQToNL+jHdYobhdCNdRu
kA7qEskCfEvivV9QIzM8ztFniGvkRRf8LZzt9wXR2h27NgD7J4U5NoroW+UXaprO/yQhHeDSSuWG
ayNoek+S/iSKgqcRHe0Gq7fVY7pR9GL9/lP8M3OGaVjuhWXLfKHIgcxo/knckYkC44iMyH8xnxz9
MZ/qhQf5cYM1qfyydnCbyk/+x2+iNGDhWTzAcefwJuXaBV1lfFGGzQpPXEBXyJwlK/7ir9b0VzKh
pYB8guNVv2JVaY+BGNO9cvTUuAbMuuVQJu6NpHiV81LOS7Z6pAP9FczDC3EcyVvJFqlvso8zDYf9
2bMKw/mWqrpzcYBA1TjSqbKdue0Oe08hhDz1de0S+LcSIby0ILFA5LwtpWy2jAAU4y5LXhhWatWR
ytpBqAWD6XrLkDKqpDz7N6AoR58Bo2rSL6UT0Ran3gBWQ7BxOhAcUJj/45lDd/HVMMG/JjmozAQk
uaDukVjE0jqy/XeawELrnvyhMYX7Z/oZZMwSd1PPav6hXy6BiR+av1GFyGW8xp1QYo6SgTCqhEYM
sUlTxJLleqytIPKwKnJEjlGjTP1g1ckdJhk4fEgOcsiQe1uKFBMOgqzJMN21VeUhYmzYRitT16GF
UjOMyh4KfIGLMZveSfU3dppmaIGnLSFRG2El/lLU+bvVzr4WZKD3RCqIoHrC3rfWYwVqhYwO6FOx
gO7TwlnLgvXCo+yCnbIZG2/agThluse2haNJnJ0bmezWnmslZx5DS7ENZdUEDBsmgf3TlQeFbYkG
6BP69B21GSwLJ3gQGvRpKfEuUKtxCJBcCzgg4ktoYV10x7H754RiSJiN0/4kIy8S4V57SemN8GzX
mwJ+fGqePAmVRloa4Ij2q+kei3VN8HoSQdYDaVC6iIKaYiOtsIOl/c31p5oOT3xbztigAsfgFdYk
7FYvtq/8+GbI9K64RSlt2JT8kqAQA4C+k1Pr6hPLMdDyDsljOmI5ApizUxp0CXcxTjtmK+5a0CY3
h8/JJfN/IcU/FCUtIXKpPqjb/ctZAYwQzAmpUkGUMWjWdzXG2NRVXDZpCeX4ibHavrvTJQAVltt1
Ml34Auj23ZDLZQ7m4KkshSGPTOagE+Oe5XTtKag6BzgzF++iO3cpvbU41EJPZg7hOZzNrivBLHMt
mfj00zzDOeeTiaTMN2BnYlYnbMBhos12ZW7FCBkuLjgteretAGoYoPMWdGJls1iM3g5R7RfqS/zw
HpTijbFIf6QnuttlLHFC/RwnMQnZrX9ZoCZAlM9huhEYLhJQ5p8erNWRRMk3vfXxapiUB2cVRtRq
zinMGLfVCmPlQU07CkGN6BoEpO7mj4gnV8Lx10gJYasYO2BY2ORbbKXGKHPSkZBbitpP5XMw1l7b
LCA2JDEtIx57qV7U7vxb4Mn5Ozldsigpbcs6xh2QKYI7/EiQ+dFEtFpF19qrcpwYL/4EWOy+T5Sr
T1vH4hsAlUNv8APPWnbtl9LHXeLZ1sPOW08MOcyHCbacwWsxNEB+axFIkXVuOHPYhgdNYcSqlSbZ
43zummG9/hF5eLTBIM+O4UMvBESlU4acPhGYGu6ge2L+OoF4yq66BICU4dyqvdjifkxXufcn94wb
92Thvs5rTmyvmyQnh98ZHCm2fqwgrz9E5ArY2MS78KMlBREsVbOdVPF8WQTmcX7W/hSTRs5oN6JU
nKbhdK6epPdUe7vNx4lQihaikI4y06l81wgTbZklBHucTtsMY54FZuR/cReabxVCkvZ6s3A8189g
TJlxMFWY5iAWpHofZAttt6CS9ICdWj6/9v8GvtALPGuaAZFpOWANB103h++PBtkMrtg6JLt+VU9g
QczCWkgqPH2+9K+bn9cUdnupNskENDRtQhA3+tPBZvWxOOX6LT/W1k905XtQkMv9YqzbIgCAgOAo
0VDg24BIOIdVXt6ISzcoIEAoBcJXuyQhIgtennANnFot9Zkq6QERZ4e/RkoSN/dYzyKxqLgMwA+U
csJZkjRjkv1UJ1snOck6w80zxRk+9hU9muIRQCKmXgj4n0HUPImpVLdJc9kTKf4Nd7z0E+fUW0od
TsXdzjssunwt8u8sbYq10ciJmJgz2lVbm2ZDtlDQgFaM05vR9TQYzhd3Byu/Qx+9gNkKQKmPAINe
BsxtS7nBBC7vHY7ghy6QIzQ+5CU5CqhR2UNVPbKuxh5uwNsJSwkfUZCEFNke1r7KjioLuea8WXgJ
9lQRqeWizEoaJd+dbDjVOJEaOwRkgq6OFsTkfd2ODZkL6SttAbzQALxKY3cBIXai9xnbN1JVvNKd
YOdr7HBS8DszTTNio+pJBcCmQquKVQEqBxg81RvnXJVmjEHHo2y0H2orqDVoUYWZ5cD46Xk62GzD
DVLpOwa1mt0mBoUYIF0lYzDom7N7Irg+BvAXH30eApzJxfudb7yXFLgrm8ttieZ74CdcxZDF2JPG
VKQoTQm0dEFmqXCrclgt7M4DDayq60zgcnj9kJMigp9Egi0R7Q1qgAjiCzUUjN28FEW2bwrXlJSa
DSdlriOkhI5N12nlAKfbWDhepw8/sW0PqEhqNpKtNNa+EIz/aVyWk/cOauVQ9J5fKndebsP8q5T6
7qFOWvLW88742WBjDFbdZ81JehVautYNj9F9wUzsI6LH86k59VuQxXMcbmIHj1jO8UQJR6K6c7gk
gG9QfwkE3QcYRri5GfVPFL7S2fHigE6P8Z8H9tV0PX3jMi5J4mWNYcRvqZwKJX3RDBDMHMVpAWNo
8QT2NkalOdE/By1Hm8yJv8DDhVbgsXy8OYYm9kZO+au5heUn6Mu5ncsD4vdRquCDkL3L9UgVnWo9
RD+0CbRSeTJkGTSQTO4nV6JeaJGezXVRByIuBzTLMTYsRs/Kn0/AMQNHZrI6x0jRnrQnpd22uj+T
OLXqp3NSkOBkOQnMFKedJ/75hrMnlSgcAOsy2QQJW7gsYyh8Ttkw9TW6SRqplqFR5zjVr28CNphZ
X5dhVAU3lvsfUWBaU4WqTkuTzm0v0NvPOiVJl6vW4L+tWXNerx4/lqHMQ/eesucmdsZLLQoUJZcM
xP4GtMGpiU1Xu/MT9EzMP6pKSjCL/bcVeSL4CvAz97qBGvm4BMuOwJJpd07houXIfY89++b/Hug3
NeB+J6MQof6hG/V7aJ7lpAM09CXf6gIUbzz4LNh1BDdNXooA4YFa6ZejMZAEGmsoUkn/yUzv4h+F
sUjvfOaxYBKSCH/PqYUXXsfOSyjBj3leqizflWWR2e/pjyEXJ/2RNUY9s/6ed/OfOtkU92Ja/2uN
twniHlJu6RTD5PZKBTWEYuio36KeVTRcRkGxjkfipAdjFeGFE3ZW4fFGzSD1ptsP8SoNJtrqR5+a
fcIyFejC7RkWVMHNHFJleaVPFsvhplocoKHa5TZygOImNnbYou/DiSST2soLJuv5qYV3JtucwGUG
Bu7O8noKZffWT7kRzT9gCBeKrvKKm220Ta91dq8cksyockN8/H/vojITg7o7vJqAEePinBaEhecw
LHFNp78m91qLxGiQY4pkkC+ghtCWWa6qp5M86FiVSwI2mCn5R2wDKEywynOrjQ5tRB6t0bMJLcZR
tEttqcHgxvN1YAx6+FhTcaYe9oxvoLfUxOvkMAi74hkr28nrUdcz17Ll2BttaJX3p53WKtZJPm9g
TO9yemGjW5SHHlrT5qIOd+MIaAmvJ4L2/hJeudTe+FZ8qighjM/fHF53B2mvXXIzRBFh/tUCHOVJ
YD2bi8EqGZscHe4gTluosvOoKH01G/HXABXMRCsr/TNdJahoTBhkUkujOavVxac3mY+pSuFzGpCM
gTCyfZLc7UtbO83kIdRhEAyKoR2YjqVMUpND3vE/6De1rOpwEccbQ6ZL0eUeB6o00c8S4f8pHG1S
t6ubY4vGFp5YFtHFT6J8x/vp9XTRxUox6uHkmHWSQXxCkhNaQ8YMGLzsQLlyldOljJsE4C/UYA04
TxJCWXDs0FT6miC9SVQBXPI6zDUE2FJiZDMC1WC2rhxfkRrMc2/SN+AA+acaTMITadvBDfvU8FIC
0F9C4RoMGezRmJ1KgeazoS34OSeu7mTqkEryJeteAQ+kk6WsGRsYq2czHudNOaeSuAXiCvdsJuCh
6wKuwzzUMUy+lwAv2ei3PNZdK3peYm3k7U0+NDAdyKCmm1KPUYA47oc0UlPGakuInT0xg5Pk0trm
/3kHa5+/NWzwEnwt9jjgZD6Rzdoa/jSt87n+I2tIPSUXckfbJz/njuyQzw0meMNoeNTOXaU7YM2R
TwoFFGsS2PUetcvAGYmNAGEIICw1whbBbkK/wpHRpyntvUgT76ZTWOj58yNXRmoazUiSxnzwUdPJ
lPe3ByHoTGIp7hdi1Dk6P9nVg0aC69UDD/JxC7BBdBCpKH6DEmqpix36b8JcpesiFuvIOVRtlx92
t42+OQIp9AqfUge8D7weIfus85fdyiKlSuEbk7QWue78+n+KGdS7jatQq8N3OA1XcamjEjJ2PW58
dXScMP139g/7YpgWI59ljMrIIuV0G+c9jqs66wcGW++P2tJRZ9/oD6vsf+ZALwS66yaC1MOSPh6Y
cQl7AtnEjqz5HLOqY2kQxTrtA0O1fMmETtQeLpWMc44BoKEe1KExhQhcJQgwzVVge7vUakWEhZ0S
Rg2tCT3JmUg+etU8SBLB98VWwl5eLfODOUTEsotlFz14UXuOeOdGVMWACqrDjKH8sQWDI65v0V7V
Q77rE8LKNmDKCM/FePDk1JUOIbbHcLdXVFmEd1e7cITnmdh7DMrsQZXNRB+UtF4ZGJrlmwKT0+7d
12IBP347vIo3gh+QQJaz5EJZrw8XtuNv8yyrv2trgFoXKklTSPPymgEYbphXfiwiLBbKy6HRMgzB
3gGBHWLCz4CV9KlkDKQK1lqrmIaAW2PFnDqVbzcW0AbGuL8PWMERSkaYfMnQf//htybf61eyfeJs
ssCH1qc6YQjWaEPFROPRBnAfMrJb13R5O3mZdkhQWj0uqQo30tWhIr6ycoMtToVdsgHtK4j/fiMC
yU9S26i4hMYbeX+64v2WsP4rECqXN6IBYB/mJNUf4mIhwLNcu1L1JwUvlq+WbBfVyBXX204pUSEA
SAUW8lxcHHuugHkry9Mj5v+qDeT6L2tZ2IeksXZuAB0jeDyFpv+hsgiQAelSzJxXesZ2u/jxXD1k
Sk6WGwi6+29BzbILBau/JCVlYy3vtcqpVu13+GvLyzs5zw5mw3qceI8fuVfi4tnxbq6n+5m9dyu4
PXDNmzXTqYMYnRTX71nkqETwJAyVU5wdWv+IYn+DNG6CiDnKXlSfH7ccqGi6wAnk2L+4SzRBFhJL
aEiJV9fY7ASip4nl1PA/v+np48T4UQFGLatcUC2Kzxukvr27sP2RSmn6GrcFTKS9OhEN3y7nK6fN
MOs1vhOyoKyM1J8pw5Cn/44FkDx0WwIp4mlpNCTpIc7/i5dn21kCTxG4G679hnrwh593iqmlSL8O
CcjxZCqRsEQEhZXX8YLyUKv4jMaw6jJqnPWKiuGHiy4jfSWgvjF9t2VZGXAYiFtxZPD572KkdcfO
BZdOdJVzW7SZeK2oMPHFCRhHtVnlC+LHWj7X7Hm+vX6toREp7TVm0GgFwH6NKCZ3BhB8uDHCaeKQ
yl1c9DISB+rUohXd+yY/kZkZXB1SeXtGd1/H7ZzKBqvOXoWd2JkhtrLKWVRvXoQX1zkmScKIC3de
N+SUQcuhMs1r9/Q8eaRh2YBO07x7EaNpjbIyy2uZC8YFU99jDyXY+3hz7TmqPL010q3NfBNEMOgN
heWwN/FJRA0TQbtciEUf8Z2MKce6I1iWuPknJbpcDOHkuNa2WHzo9ttGJ6fV0baZUrjH99e10Pe2
n8QcbWb5FB+OB8xHEYUPAya/UgBMOo1u8HKWvwI84ZNnXp6c2YgGNyjK3W46AZiKrtAhzFpj0maH
TzO/QC1ak0AqX1eiRyi8eYPDJ8G2rJTvSQwPGA2MBFpp4xd9mfcaC8URJVu0gpoH6GMgwj3IuNOk
gy8E3ysA5SrD6KPi82RATpPUqsEkEPAZ016CYRmVzTHf/I8/xJrmRvtaDx5vJhTf+TWsCXXHav6l
6E5nWIHFUIeMxmWBmN3uHcWgSyu1BtZjnz6XheNdEIOk8Oo90G7Yd8XlP/BFpK5o4xR6iCkdbHzF
8Y8QNB4iIvRYLDhQFa6SAI+8fwKU5ZAfAGG7IeHCMBpSsMTHwy247X4YNT9xXi5aSy0inFXdu2NZ
bHndbzXzpW2X5Qmrz/tO1cEoUUtcfr8+oRMW4MHwC/52pz8ZKtzxyifgsAPI2qveAAixeI/H+TqS
qJDakgES5dvwnPzC5i++gICcr2wbD5mghBoq9taYeB3H0DKVBQxMrFtc+GhVs5jNaEaEnaBUIn5o
gWZ5L1szOG1GiBIjhPtTiMMcjAn7F8YJCbsZHoLalFCp5rNBwc92W+YO/bPovD+DuIjDRkHg4SDV
/cVS2j2i44XTcZ8msMSY5AZIYZ2Qt2niw8VuvWdqwDCDpSMu2vpdjz7jATC0UehypnieRJVas81F
KswSMalkqChGbhx3ZRsrMMsJahrYE/WPsz92P6K1KqYAoMsy6fXcjkn/voFLJKaJWTFs2QYJLI/I
L/3/0UN5VP0DgRYfTxxQjh+jfryJTvayg0CdA0a8EjmDWREvVI6j3HFt5T+ohXUVrf/lTFXfBsfv
eII2sVWhGHRVVBFPdwKqPSPDQutXDvWGR45l0qjij/lGFNPT4ERgJLMxNoVo+xaaiVZvGqMrp8mD
SNob3GKXqW28jqTzIUIlQUdV8t29EvjCpYfnYXJ2jpQhLFS7y//SdJI2xTOoB/TF0zyLpbK00fDj
bE5pEQbUdLs4wb7iWmSj4tY1F3wRXqBw7FDK86bb/q7h+VTrv96pS/DwFn/xp+QbIvCYftP8LHsD
g4hxI9n/H7/zja7KVu8f0RpkuuiBzbXyufMdlB6/UywjeqEKJE4D8IBbFW5VxBupB4i/Sp2cS53O
n+3lMnDc6xGonnURjUQQfIPu+8hxP/eCHifx7sPyexIuwsy1avw17zgj6EZpcrohwNR3pO+DVQUc
c2oDuWTNdc6sGxLKBIROXo0DanHkoAQHbD3cA9wY8bd17cKK78EfsEamGYJ0wZIHWAMZsjUZMJkr
9PghraHMEjX3yxU9BewBGOjlIklINRUdySk1q4yOL1aTchUEJTtT/CK4K391VV00KRPg4qVIkXZI
ctuKfeL7JLgX75Nl2RXzK6hLWgeoafj0oD0PB6RTwr4cgnRhT8GYdIuj7iBbY+Af2mgE7GsGGiC+
z+4FvKYTNtifmHIAi2H6HC2HolMwSVlDNykjlRxcNDgbJmi8LPZnoeHE9/0BBjcD+2804UKLM4jv
khyyXo91vm9xNHiLfiy8Da6DmHCrl/b62L1LU5UBnPWR2Go9RZ+1fLFjC7ZZ1YDSwmi6ZojNfaQY
Vyr6D4HiQF7cmcaJ3Q67H7zW0hIE4fYsRFKhVoL8xrUHOBvHWyc27lNeyMJD7RBFj57URhbLBHpO
ZgQ5ICe2rIeBxlClyxTaMfMpDlWtc3uW5j9LHHCHLIEWOGbt3rR5NiDdEBPr6Y0R66WEetgKVqwT
kIgFFMtfFEcl+rF6gQZ4HFp+ie1a6Bl2isOdI0C0OFWpz6BRnBPNOf7bOSU2Q2ERj1lR2f2GPN/Y
4Sho6PM6suT6DzwN6UVxeaOBZXvhloUShqxeoTpRNBijzrabsT6PclLF1D+egW2M7V2OgLMHmZ2v
XRDA6TjQPmDWr8dKo6QuhrmwhMKgUMFD4KSTQe0AbjyLc2FtfuJZDRIaRNKmdjp8dOAB9HYlRkoZ
hEKljRNShiInyUuA+FT2E2nJ5Wun62PDy5gJxzuoGoSKnWuonjtR8JzPI1hVMMgTHDDNlzWP07nV
37r8A7wTD9G6Pay3ltHxCy49sJWgbMLK1ths6aZ87G+s2A5F5jl9RpCVBm40O4MAtuHLJP3lWdhK
QODnddNazsdyQFcEC5UlkEA/cW8jkPQJjqkptL8X8ii48HoApNF6CvIpJ7zYbcOrBm73Av2sQva2
xPvf8Gwacy0vM+HWTTHvtfvaBAuestH6hK/pafzf3dbDAsluGFbAZM56kRfg11pxwkw2fzNDrJTV
aWV70T38S5VZvSNFt0P9ZJA1BbxlW3oR6kD5q+g1RXdrCzat0+GMeK9/+RRxjbNx6u4ev4XXX48v
/d18MuvbJDrQA/wYI89mRrZNYmDjgvHRjUuAXru74wb+Iu5QRScKgp9Y6aPrFYHHvHlsr3Hnz3Ax
jJ8vws1lrMHkoBkZHhN/sRcUbg00tqiiX/M49D3p0SKbRk3HP4zNU4pY5CXh5kHigb9RM+4trA+g
h/US8cCiFqrP2QMFMzWC9p9zgmVS098TWQg+7s7vJessReRuFb/iV3hrxxyFoCbuVnoayAR3jaIH
n56hGbGWIigjpmnidHc153oD22Ery0AfTVOJl4z6jlRAtVg3rkHzmEuyLodOlMUynKIuKJvoxNgB
HD5mA2xwyFgHmU2880gs6eV2qtZhZdpy9+86horW7sKhup150vbyklqOJQSY0rgSgOJFNc7kSfm8
1Z08Duy9rTxpymyhdIaqe9LyTM8kNEHgpnTlTy+QM5nWYuUOowmcoUOtYu89V0HtPj8B2KgHkaXb
5vtnvSLOipIRcWwQogfxLdmBOVqNtg8yEElouTGkKBEsItcUpuPrEYwghz1gMW+z+PEoP5lN/163
fMUoYAsWW6Hgt+RTnJONZv4Pz97x3YmrQ13wvD4swMYBlEGOEOfCAXQM3irG30XHrgW6H2VKIwat
IpLJlxpC+UZ0ty4DQwAF7CHpMRGfEOxJerO+6Era0nAIPg63ItMxuzF4NhrKVnM50DJZF0Z68Zx9
mFPD+xk0bmoAz3cXeHIlsx/8qZZq1uejqu4vK+O56hmzkWfzJPB62+HwHnf9yJRRIPphNsNWMZK7
U9mIlTC5bhTfgdPaBIbWrzpa01lcyqvixuinueVRB+LDTzp9Yh1ihOmk1TxAb5rzJk/7wiw6Vs2e
S0AtAnbXWdQMl2BZebMoNRC9m1+G5D+b+ITLKX6QpdVXhkUMYTh4ue0NlqV7C00XggnCS30c4VZ/
0TMt24IO6b7dnpDbRgFq3KtRrVcYNusqzifpLzgge0laQd1LbFEKjLFCET2Blv8av/IcCbVSHNwT
k8iKRD7156MHxWDxb7DIbXwAMLOdY0outJoPxFS65oKJSaLQ5PNxGfzrpnvthHs1jiA901YecjzW
vteYLQ8FaN6hB2TIpMlf70g9Zp4FLwH4/4Ic227ptlNxON7jUTTlXyqR8TxoBTGOzA8n7hqcZro3
4FRqYuFg44ZlMqS76DgX5x1A19r6FGQp71lrsFcJ+j6+MRfTN50ZBdnHFx1S4CuQNo8Z2+iEkRUT
3vK2LttiaZbjLYLNvXizfAd/3ufm6yGB96L3VYItBH+fXQGumbVlFkgVj6nFTPedf/pVb1zdYsUR
j2pBRN7GrFdruTVnM6AFTt062Q0IVK4diQ8KSmmHhIPcX8987sEADMc6uBhY4j773dlTRGjXV8Gm
Yf7bB/Oo6fD0ltk3c9xP4fvyrphGnGKeJKnIFEfeJNE+upg7nuds3bQGBO9PP+muAtezqXkzE4UF
ESjRT0GJx8kjiGeGFcrYQXnZU8SF/IkzEbnHu9eWCFSd0wD8b/usZ43FxR2oRezXD4TZnq3YRd6u
sfe2MU8kZBbRcde1Kmi0HT00y0S2uvLsT3Isdkq18qakFgKelsvh0kP1PXGuf/kYwBb15LODksZf
Ak4OYtJZaLNi0MzNe8r2dLVOxnJqlyng6S6L+UvwrqkD+j7YeaTBzgyLKdvKqlg9wvVyxjga+53i
kbbWrfxRZM4lcP4FVWmnkGtkV3alFGv3zpTDbJm0wY8SGp48DRKaHev48J9VSzp8PX5GjQTy4beC
NQNTNTczQII3PGCNHgWwyNv9oywACVcQ+6EV+jBziytzAgQR0WgwIkgoUAjIVvDHuWNMuDmLtGfz
p7o16pgSfmucCHODrqak8Q7KeA6G5DGufwt54VegpSdzSKnzOwKDJ5H3crbSfnUE9TevSUEJbtvR
xFHcJPntSwflGOLiueZTRpTGsU27GuvvE3Jw/smxOJnTSSJnI6EVhEWY8um9ayxAurYLg8iEk/fk
jaYl27X3tp+3NQgddUHqOlA/eP2B8LPSFmT2szYV4CTOoCJ5tDpuWiSbYFCiaMAG3SJtYOgPJBGr
QDsKOb49md89kGYFf4jK9Wt+nok9O+G4iOdhkVfAkNdPKLM3QlmV+dyzIm9Nf81l2tlnQppAecVy
h6E2l1lQRYoh4NqE/OtdqBCI4NNLstUhMald0t9h30qpqioqcKz5TvVA6JISW6a0lr6Oi2N/WADY
1j0K+XXqCAg1lqGU0fQY0gHh2R0OKkrqFCi5vdVq5wt/ytSOEy0VicOTmPH7Mv/2tS3VyOyfKK1/
oc5uTQXexRmkKdObmj5Bb86rhw2/2YA5HclRJAOSxPcpDcSFRsRu+v2WKz9MxUpYv7E1iy3Byl+4
b22W0k/znIECTCj7uoAl4e8BesLc2RBFMnYddSR23/KBr0Y9LKNUCMnlvzxo+km7D+hMa1BHHY6I
0PYpTtIpPhamVZzPFLm27aWBy89tm+19LFg7sQHKyjUQY16lokdOC0RlEhXsQJtBB8QuA7/+Ih8a
ND6rSBgxFCEcv1B95AG4eyXHnFaX0qfe3VMSqy0e40bWyiNnJ3J+dge/Lv5Z4Pi34OCCfxkdcWlb
oYGTY/kKyJ+9jNU7q8OY3gSDCU+/0BbDrJx7xEZWtJ821H16lw5gYv3kEca6b8E1ht1Ihec6N7np
JOklZEvbNgGxDtjpm/HExf35Ybj82FFACSJ/u+52i4T0TKr5bwWlwZ0GhXubxJKHPbQA8boIww9P
p4PYt+QVndg8hUvevXuuPMwqzLwRXt1BvrWh4XloJGT88httyJZsip9Kp3051nxAE+rkqgjCCjxO
8gIlgGbrjyijPFtkpIDhlxI57umEdmPqa9LvU1t5MA9ua3LqgiRn3hkSOWWQZPsXKbdPm3wtCkkF
TwEzBkQM2e9pnEOf02Y4eD3aGMfH/RAj80w5ctWfsfBBhru/abiukMzQiEFv2JpFPXprVFWMqQvY
H6UcLOeSwnvJkg9v8G4Y01XSxxppkLpaQNVBHxntD0RtdR33+nSughGg//8bmJRg+/KdyAySEQoe
/vJMCFAWvmmXHImt+zP9NRVg3Et5nCtLNyZ7S6v4fXMWndyH5Qdc9+H6kyqs2fuTks5q5hvWEmMJ
SeqmO1X6nUkpO4hlbNrQnBHgLBscH1YGdgT1EO7tp0qNg9/fqvSrN6OjlgZwDdb23C2hmLb7dKQ+
RNIc7NFfBVRacX/6NhHxB919jQGDhYhEdLXp5Mnc/Q8XGZYjyyTQR1FwKTmY3hJHOY8gv8G9RXk5
/P6Y1Jeyo6JKTxyIGZn9N7DoN0oVrmSVKOvJNJF0gw309C6KoQf7n/95GVRYYdmEeiFNAIp4XGFY
qpfQQuUV6s0gdUduc6lT0VPdbPFELLRnUX0yV4JBKe/239FG1vJf0fYma/pulocRJd/jQe5ta8AG
RPsaPQINiR6gatjsiE7wUUEX7SFPUu7PEa+kOD7vL6WXy+pE4bO8Iqzm+e6ps4bRHtqNR6O7C/bi
D44fdGNHfhSqJFkQGZsZNShB6E6Nju4GkI6logrEsEozSzu8URh5NkincYmF9pbcdA4g8TmN7YYD
MVBSs349N6rPjrhVXAB1qUan1mf9h/xLiKbQCEOP9t81XwSwGG/RTganEl6kO7iJGUoA5UY9fFfv
7kbfTtiitn2J5lTVnQs//VLCz6Yx/YwKVJLbNBlW2VmdXLEOODsTxy2d4F9RX5dlBTVdHctJ20tY
7eza0XN7vnVnRUhc56h/LfLO9FiU/2jH97cCkbp1jkPNW8FD5otWuIOAENjVYNbT6skATTrW7pCR
k++rRU5K9Jro8yLqC8cy5BqE7SHBMydmLiUDoPKAaEbT1t/ztJGvscDvsCVgYHwPQY1aQKhc8PPc
FwowiGU15Ug+Smw6kpxjf3sA1x2kJPEf9T9ZY8/5xJT8qjmrgg2jw96hZdd8iP/b6OGvXlRO3KHC
EBcLy0D9Y27Ym6JKh0fru4uaLDPAinFS/OqHf3USv873kKQCyKLZOcEobPAl2y1KeqxAjpRm8gUa
1ZXbiEcqbFpWdLVy4QWCRYWhcw/GoETT48jmvT1ytUIGv2dHFv66EHwVfuE6B1JYuhCQyP8Gl8cN
I6kslJV8yxOTI0kFIFmkfRZ2A1gqVuLxvbAwZg1S1LUnv9+4OuBZKyh3L3qyXUMa5i7N0zLoJ/H6
QH6qXh5hkOdbxHn1Ym6WFv9dzNBlyK2mH7M0SIdqSoUGD9yLMI/0TKzOoDePf3XxTIrFl06kNthS
GRcDDDffJqxHZsCFHA1r03I/XVAZ9/rn22ykkBwDdjcFACFBWWiX+HDXbFhoRhBOu+2+yWVW3/rn
z7fYTyPkXwwndUVD65D2i70SgqwHNV2/27Ja9njAx4CER0IwenBnhVb4XWM1RGxc7UMCwSn0GXgh
j98px8pNXDeW9VsAEHky24Yp53zuXi8244FdFnc28tmLWqrx7W/hcxay0CPne4Qh7JXOaUA5GAr9
cEyoCEW6AtNsvwRtB94ZSgVpvBFtGYVBtxhGtUz2Ion2Du+ltVfbbLVXKUopXiULNXKPHCqFngkc
8HBBOO6Zn0Y+dWBvHIT5A9cp77BYC16d1UNMc5Hs9G/yXthQdd+L+0ME06DVb9IpARUFlz1qtYDP
lBP33psL8r4ohs5IEMG8dw7xuZTz+Gt2FlgKETgi0z/ACzeIxaFglXYKAlZrwkEzmsgRbEeIwJA6
hk6hkCbqg1mmGKZNB8Se8ESJaWgvgzD85iF0MjrGTgTy7jbPVFqKcG8bxXHyRL8a/DsOwh5Y82tY
ijTTwKlrCejQKcjewu4BRU1CISXR5Q6VaeX3kKHHk7q+NoRKcV/rPjGlzRgpoEt+1uNQB0gBxuXk
Q3Y26LMe9Nk3aAfRYLhwr6LXTSgpUsuX5Gork7U+/VEKIphnidPXb/4u8ogXxR3waOLB8L7E4AZ6
7a5s3Py/jz8ZU+ScOpLOpuW4N41FZOwIkpb81oqE8WPrrvFNlA09uuF0cHpQ8H96bghvDU35kJ6w
QI4K5FjCANNysytFfi4giWJ1PE0Ql8vBwU6blx56yUYQp90xRQH1+swDgwmhIXXxZEaRJ22Un/9t
5HDKHK/jhXAVv21PpmzR9K7x0P1r01tcUyAmnxgvj701KMilN6ck16F4wUO1za9su9F2n9zW8CC7
kkUe00RNSa1Il11mEzkH/S7vhyhRHyhwocPqgFG+oa6wkMvRmYKXH7TcV4nGxP+r3IXp+BQEmXz5
mmEq3tmtIuWLqLfY97STVW0E3RsmoyZAhSOjc55WTVz6IKYyQCMVcpp65YsqxseatpJv6CrHEKOY
IboTIjD1mdr2K8EMz0D7KVnWNw7Tuz1VWk72Su5Bct/5ZEkJ8lflQSAOG4FJ8mgJFMcPKXdb2TdL
Rgrg5gNvxUW2judFW8sXAoP37HyW7fg9J+JgLRycyz1FPzTtx80ML+dFcsX4Bie+1h+Je/ZUnFNA
oFnCGZNWhr7hMfXPBvUnENdZkx489oHs356K+P0BjfB7+Pz1u3tw3kX2KkwGyo4sxGrkcE0G3QQ5
0s3aeh+/N4baHjuUoE8mtDTZ41lhnwKalh7YZMrNbEi03umSd5FrdI5nuzonlKVg+B/UhG/Xp9Uz
oNZLSu8vVZFe6z2Yvz7ADo7nbAim6jBG3hENRRRCE/e6NYxVwb6zZm6Z3R/XKrljnDlyjpjzyTVz
VuMd1ISW6aISahRvew2ciWOcdN58s9QwWoF+smXPjzkhAmqLYAp/o3mL/zGso+ZNdY/RT2rEJa9J
8Ac9J4kXda2bvPtLFxXuslk3oUs2bJHqq110Agsf7he/uwQAtaINFuyFHnxYg9qObmtecAUGFb0S
0nG83Jn/uPmsDQTPYrf2vC0jz/NFZxm2myMryPo84IMZ2ZvvJl2/PB34X8QIgW8PwMcE/3LkT62S
o0bIyaXt4oXXKI+LZ/sEkuzlmfubOislvYIrJ0KPhNMyNgzJ9G10OPwT+FUrEQ3S/PpCjdMUHHdl
2lD/bv7SfIroEnOerAWXHBU5C//+Ma5/l78iVoZiPP3ENLIs2xCwicFjkVynF7xGJEq7BL3V8/Cv
/Lzij/DHEI4J98VJGDOYRx9fAMjKwxeDqN1bwSmbmuRSNckYEws0rIvnkZH+Uy9rhjqgrEFjh3st
qYstpgCIKRLYC0dcZ9aejgucknXVhsoxEmoriEVhAeg2Mv5l20GQitHSmiluRhOQPnWrsH4nGD6Y
0vjv4Porw40j7rbu1Q4lHOuE0bLzuYNnyXWaufCmYZ1mSnMsh8vYifMH1CjB5ee0Ksp+X/Fbb109
iM1nT51FVWFgnKn1I60PW/LTqfxO3J8O831SBjoLX0nmITFsXf2a4jgA4EjqCqR+673TYepUm5pC
uxsz2nRsx7Pb64PVVq3Sbhz3Pp9riWaqkec83zLg3zJG/11MuYlXSnQgfeFdAHgK1OPfJW3cArYo
OWbbSRWIwF2LkYZbSiu1Me0YJGaDITNgkxV3Wc6HX4eqBn4v1jdhPujMvaw6wI0kAgdiGXEgpu8z
5wqL3SGDk3qLHgHr/lueR2xd5CnzuIkec6I91MH/wMxWYtGNKxu1U9uYYLktPpmdgZ4YoJLBZY+c
33P3EtsEpLWtFO/2co3lCGc0qD1dQ9bkVPsGBt7prnmDcRCxWnwO9eRlvH4vjgdN3pYJKfwItIiQ
NnvT4DUHHs1s9lMYFyRRzV1RhFgJWZgROg91HWfpnXRl406aSqDuDyq5vsz+3lNSVbVuKaqxQGMO
F4bP4NbJKAQ5wpWGSb81qn6SaqbVLb7Hp0f8SHT3iEm1m/B0UrDYnN0zc+EWUVMz5UTrkP9tQ8Ub
+FJDbmhcgfJZenY/+Vjj08RigQ+d3Pmmmt80H6joQCrd1rqmgBYgCExScIbmkeDi4pCPKWdb9Mtr
WnaBBDSZBL488DEsGz3WjcCwZ08uIxT59Y5pRnVEyiyRkSSHjpN2c92KZ7JJUQnko8ihOyCww5tc
t7BY5pRTIfrx//7cDHhIWo/kKeROpzXec5LnO4IChEnWiB2qUL99H1eYOJXLtq2GdhUrMSMn8dt2
bqbZ691kYu59o/c2LW2oGpo1uAB9MB9c3orwtdPYoHhIakFYnIV+AoFG4yuQf5KfHH5ATYb3EsQO
kzwmzR1TjaZ0fSrsOpWiMGkQUS7aI1dzVUezN3js+XxHF3Lm20me90RHSB5FibKRKi+/M5rrzRdK
1CUdl1ga9s3ZeKQJhvsuMe5yBBMdoINQ9DbJdFl5ekgqp4ySB+6987krO+4acFtBgx9u7RymbZ5v
aqZPMEabceazpdJ31ETEVoIpfh6pvNAjojgVmaZJ02+3iR9plbrJgb5eDY7thFJzmW+krVUhFPyv
355FDEGtKlgWZlv7qHoXcQivwD6Bum61ih4UnwuL0GD/aE/uFc9m/MVmLojrV6yu89ilZYaTu7MO
O+8/Avs4/Tl26jY4nh1c9QH6blTqSakcCph8gZXVhM9Y+WZKhSKyCvKs80pTD40PAO6mROH5JcAY
GIpIZk4AikHHWWneU9IpOouEPcZVDXHUyHM2heZQCcAW8uLjoPx+sLWz3aUtIVIx4f7WFqFWQ/mk
vcR2URD+iCIi8MYjRpqwhaHDkXMVXLutdu7HynYSeCRWaMs9oWBLDf5c4GI3hIB+mEGJ7CQCl2mg
xfxtVCGkPS/5VhRuf2Rk57UUkFPx6vagdgevqxLOaPJlJ/Qrkx8juwaYPlcNXq+wENf2WweREtLV
whvesZA2zYItjEYqOSsL3AG9/n05HLUQDcWu+JN42WwapQ+gwS0nyK4Pe4druaRFCwVeErngVSPu
cbbh+ycczBpscZUTvw52JsgSHnokbnilyjboJkaD7DOF8FgyG1ppc9brsvRc2qZreHOFTbkHt5dV
167kXl3zq26SzTB0I96JOCtSuopVvmcQ2jZpwOTWMb9IBuN4x7bH52rqmJ/aP27rGxR1JWh0z9bP
fnQbTFHQxsCLxTUtMLjmtTAokWVrSxuRHWenQPRHd4chMkEN3PPbCt8R43f/miVt6HhFxLmFtoD/
mKBjgp03uz8KqTd/8lgz0RtRGg+8UMrfKCaNXBkwc6Azjatjf2Z/Y3ip2KuG1XJK+tnWKpJbIFpR
DRzqlzVYl1DUGz03R8dZ5gUkvG4/P9L5T4H5GWnH4CY3LYYJPLJhzXf7VFaNlyAFyNUZU8Z5+Z+h
uVKspDk6tqiSKA5n25xZzWLBNucuztQKVGbuoLf/gOrJX9B9FOOY8fGSq4ELOe5PVxGsyvP15y/Y
jbcWuaOoW7Wx4XajJkz3MlJZf61ntnFBCT39L9m9ig4+jMttgQudUl4NG6aEGzxXDk6P8HLvTQ7R
Pit2W/p0nww8fCFUUfLDPQmP8iKKUO/NwL7z+QUCRKfOYhbqBEbd5zdRf9mIF+PvImAq8z9uudkq
C0+Zs4pJ0qeB82QBqYGENfBqY6e4f1iha958BDTzUnTDtwk6brVgeKIJg/nyHpz8V5Rw59pO6vtC
c84RZX+EXzEqSGewt8c6XykSip+C0imvtnXjHHcEPtQfR7RJ9sf11pIZAl1ZThLr+NFJ6q5ilUtZ
BF7BSBSZAEjbdVR4W5Uj2p4CjDzDVZ6Q91/lLLmhDR6d14hRfiowXNVum0QDLomOEE+m6VNmpbMo
VnqzY/fMd5Hun70BuI11l6uqlUxnT1UdlnVz2LMuFz8tC5Zs6I98GzEdfZDH0xhXzIkc3pwhE2F1
wINk4pyhVvrD+ixImEWt5VfLN5v+/5z3oEelRQG3ZhxREm8ShpNou/6TEuwyZyTjVY1F3VKM2240
49vocb9S4m0zkBudBcYdRtjwRyvuagO+MiEsN/UoVN7UBr6QVxuAUb7OT1H9ySiZ0B1tg0epH1zO
IPP2q+6gUQgzmsJaaIuQ2hzYgQ95pRh7ueHYi4TYXnrCmcO/tgCHQ2Mk5KcJf8SYLf1tscZ83ZWG
gmB96t7TtxGwI2+M/94W/WrdRDH38Ao1B4Btny4CmzvCvEFVli3RXo6LIylcj1tPJUnN82fLoBVB
moc6gdjZaOcVvXZke1H0P5Nk6fb7Prwss+F5lVf+Yr4al56Mq3CiGThkJXFxIDstM29X7mlMEGgF
YE+HNvnB2LY02ee0uD74WEjR3lqAu7qtJPxfoBLordZQIqUy6Fn8PRW8+6sLxq12nuoTCLw3l6UB
V1JiqR0WObTaIZvia54eI1gjbPG97PsirIJY6Ib7Xx+ZvYEqa4IuFrc5IGpcyllAd0Kzp7KQmCYu
AdbCQ563w11L9l3DszkIvvTga4wP4yBp0udqX20XbBqACW4Zk9rvwEYj/6bdnGVEb897KUcMks4U
4VTxtod2SNTxVOSsPusI1SAOCVSqLLPWLmmTY2i0WC7392gyORTDIkO/9/K0eRkDNjBlGFxLoy0u
AFG4o3n5kGPNTIb9tjugY/46DFL0bz/t4YL0ICVonrKlizw16uNa/8bCt4k6GqtlfCUxeQwDc3gv
cTIsq5h+uxYbpsTwYWbbeBTqn8A9xFvLZEKP3/l5xfazZcY1WAn1GFABl/sfZJRDFJBkJPS1JCHs
5ty3yX7nGw99xbI4XXvuv1MQfoOJLgyxJgEQvIE/y74ifoWWVzWy0eCrJPN1jimPoEJc01AMMimy
9u7H8Ruh1eQstB3IRzApPrLPxagaQn9wY5VlOWrZnh16ygVoEypO8fuGuJuOy2a3Z7EAcVWm/IkN
VDo8lL5hS4w+EHQTc0KTtKUGML+N9u7qyaOYiZjgdGsOcNT5nFGtOUtBBNeQM/kEcg/aeYnbss35
/lGo7Ebc7+d025C+Zn7vPf3fEuu2pSwb1BAoAg0jBc8ILPPhsr++kmwI2VXpwS8ZJWOpDdGEkxmW
0eBxGaPObk5pr2h7t8uvaq+FDvo5nkeGf1l3uA/+eYXChalKU8IZ20NM5b4rMJmH4rRpVFAf62Zm
sLrfyNewPUB07TFHo3F/GmbAAaTaBtEAALznhSARF6xO4lWJ63BXANO8xeR9fXfMlo5g9JXLkNVs
dRMbnuOsVIGan/OS4eXDXFbx9NMWsv4D4TSYYJnY9Z+6s6VB/yCjbVozPFGw1WDsYfHtXKAlvocN
JvnJNv5648QQktaDFzVWswmiFcAIdaOem5eUVqQNWQLeKra8aCLQYJjvQvLDExHkCerlQ40jSsDp
oRjZg1C/tifyZBxovzdk0RCusH/LY0lm4Mw1YJB3Cvq9Jlp1Jopywk5dDmEYNDRFEc5tj9E+XKWB
c6Kb3qe7Y/nTfltVWJHFzfytUGIGFfN2fKLaRuesi/i4ZJgkE4oq4hvMcXaj1Br110rsvzNzEytB
tFiuCxLjtrMZnA8bQCQtGTQEzqOF/rsPnGpVHLDhT9dQrosM6wKe1+RGA8PHhnCB3WsX3uExx+/i
cF6MNH1H90nLurrjw/awB6zZss7iUC2APOAqerNmcdWfghkf7gCEDDDUsK7sBPBtaJwE+6133YMH
zEj/CMiC0SoRO84Ud9Zx9fgfPrRck4TZxQJWdISLiA6I7MFwQAdM7z9hx5VlZpNOD4cO+N+ZjesH
1reEBqvxDeBpjd74p791Q9qRr4C5DNnESAz11wVR+klSHA+2/WrMyKPfvASLgY4K9WaaOQmrsxIO
7EXjpGqQNtR3WkEvkQQ/GgxMeTU4m0nP+zbviAaOCPVVKEk9z2w2sXmtfzmD4EnZIrgRRk6fDhuP
IU0632fLXO5CfjI8+gvxjcDtE9oJYHb5UiTwOZW9kIIGU1zq6majI6zDCGzKHZTHIUDpJyhpqSPp
cYVGd0nDnBokmuWfnwly3LEpAjUH2GZPScMZqDToz0gR38LGsZS3Ke2854Peuaw1v2CsUGjtSNEe
3PCiHaN8B6BunrAv9o/ywOr18d8/DZnbhKNzgeXcSCXQUFedoJ0m2lJg7LY11MhuEtaWqX+uR3ja
nN71JNR0s0Vm4ekadUCl1PxglTZAVvErK+yq9JtrndNbCwcJEmZiC/iQmbUp4etbB65+Td0x6kFN
d4LXiyWs5alDuGHCfG6HpTSYx9Xi/WHPSWkaNlipzbXXaZJXAk4VTyz5VXNgDzaRpL9TYr3jtSLV
i/xiXA6d3W38PkMBZKYjtLYw1ifnGEA0AkDQAVJzat0hpwhf/1BeIHxlwSHAupSTrUxJTjfgmemI
lAvNaWvdhB7GISImKVueqpXNB2Rsx/cf2cEKO5jKS/rXrdFQoTGnLhj+tKEiWw6XZUzvvX4B1JIt
JWrRdMbxPhWyxsp664y805APsnoPvQoNtUqDn6hwBf6hJjx0fAkMuFkhNgkgPGkBM+IZgoqAKfdb
RCa46sU3owozXbkmdlcx8ZlVYqfh+rFSbRHbsR3cRm8enqCkrGwitVri8vZRFt7nBH6FCGOzF/dZ
yVH4vqDAjxRloPFO/zZT3KAniFfzXSpSPp+F/vX3/RjetMG74WGDY8144AF0DoDEyJiScckoaCKS
ka8/Ckd7Y/7LyWUaaYBqt4H7tp0HjcPso0pfYHkg+tr0Dk5ua2ftQFwOV3I8fRsY6XCKmSiUqCVA
IJWbVn/c/fNGffrIiBuHyaUIHMbU8RB6gUXAgPaTBFu6TXw2+FWhEyqREGuGUqxLgtXWXQi5MwUs
IwjlyT3pynEL8OazFTQSyfWBn5Gw7Wil25WEbsAY5O+PKlP9aquckwevaCaGfzwe3G9gf+Aozrd3
NiqcZm08vBckP9Z+WphQ1i27ZnlvPXCRF3DszG0MVathfzo7h70GPhUUeeB5dZD3o9KstIW/OSzO
KlGkeiuyXL/84kyLDGzAkCbplvf7NCHufOMEek9py1OHyGjNnJD6viS4NjgrxBQtLdD6Wj39PUcL
2SAVTnnKj1AuVD7TQAy2UtkEzvgT3MdZcwN1+pBk2mK6xnTunZmH/Yg35W0QiMmBkA60wxVI+0+r
agEmfxxLBfs7MVV/zBJcYSlh1/cDatdjeKjRjvH/71UL5fK1l6rgZ6woKojtwaWL4gF2g+wQo5nm
MtcZcMjMVgGLwW1/YQ5xh92qqqvnyHOkVPb79kT0CU0BFonQFMbk3paZU6SBanGJwY7QD4elxGa0
ZqN9DC27X4X5djnEGiYmlv6rOowyvPw9po6ZyHMo1iuercwo6ZpuPi5t3qiI5NYToBVzXlVi3mvp
PC56KQEom3ZBRZbkk2g+GuT+CeK65MccrQM1xWJuTQH4LlVDguWfpGY/k938iIuWEb0mcdpe594N
S0Lwu+K42NaJYzjbJywMTg1624rbzf6+ISeiHnYulLaDPG3NPgD+7eZUbPqemykQMUbUQ5MuLK9p
ayY76FEmB7Y9IzUFYYKwel41J0hBFe6pZPZYcdPKroCY6g3DZx3mPBMUGojXZqmIMq1+YYfEn/P8
8EOyelm+qxHc8K7WdlPV/zDInowDffRRsWRNuRUCmTBVXxVq5B1ll0bY4delXQUyjHAfE5H2yZX4
6sI91DMsFAl3wAPdLeF8c2nJMuOBU5CNoM7QdnmwfkLFnB7CKqNurNJG4PMt0JjG3y2Z4WFOap7g
TxkA0vQf5rO3U1keJ6otziAEqk+de0t7CC0oIhrzu38H4XV1bjqDzQrrTHJNF4EZhhZwws42sFBv
wXDvtydhe6oDhRSLR8W3W8RVoy34iQpMpv004DAE6DSI3hAx60Mr6EQ4Ur4RcndG9qGOATU30ayw
4hATgaVmPFyn57gijWkVdPcExu9j8fVk+QbNv2cnCp+FcWeksVwCAyhUPtrGWJwi2uCfwjP2Egll
QtbNVODJqClRUE8OjVgPHT08ZqfryTAQsRe99RxnIg2zLzvplMkll2NEipM/kaFrCwjd+TlOw5ok
OeZ/8jLAdw7tgZCAzxUL9ueFS4Mycb7LdT96o2m2ena4MTk2z4tPBWaiBHEUTwSDWFQPkwNjRhRP
6aIFZlIP+wIMLqomWPfECB9nFLkUyQAqTjODL1Bx2uCe4mDayjI0KgiS/e4VamdLZWRbjjIcyLYg
oxGDRJMi+StcIqdQHeyUTJnWMXokEd1T77MDufjexrwPvK3X1QNbCG5Zpic/bgk7ysEv5OMmSeU+
i5VoTiK54pqCbF+DTSlYyXVT0tMmx4D0Z2ttgVMoPtsw+2RODgzB9lTUd8XfPRnant2pNEai4WeP
AsbPJXE4+E2xG/FZg5yeFK/viG21kCzNbWixf7W6JZDOB0cIEQMNCpjXCZxY014EOsZ/69x0GJ+h
ql1ZY+2m3tzfFHurilW6TXf7hLIeu2gxfqElgsTFKYtf71yOM8qu/TnVMP9seOGCABgEImHi6EZC
nJGfHDcPdqVOjNXYJM5TU8xGn73dHlRLqR52a4LoFJnpBZ4BVXUpf8C3zZSVeqMY+VAXkl7PjTXH
427o52Y1Ik4N3XMr1sRv7fJYWurRGtnzX76Nbk0NoWnNalVuK1eIw2yqTUcTTQ2wX8DTr/ARDGam
FcrPdGBQ6OxovacmON7F/Js0qtJfzoBhb/YPsyyMUH6hE0kmTo2N9TKGR/sm/xXx8o1vDGo1m/gL
wv7fow2renv5aoJjeBXhrlXjJqK++E2OxnTCeYHBqR941V4pDZK7Xm/ZX+Ec0FSQXzJ9EBN5iBJH
xnYaX6eHEaZM562jB1iFMG5w6ZXga46OlsUmlCD6gORtnzlhKo/G8M7JNx08SqKY/GHaRQTw0c/K
VZ1mF2Zt6lZIIpHTi3/YTzUN09rb0EsCDCjpMA7N/ynMdjoH9MBkk7OTqHVDVStfMRNJoyTjOpSB
3B0jYP9pOqIi7SgiFrJtZg9EIVB2BC10J7BkS50Br70aH9RLVbFDkz1HjMSeP32HN+bqQPB1I9Dy
SARgPxvmhL3RD33S7R+vRgsJBrIdtWLU/iRPoCGFlqMO0agt9TLDmled5p9WUoY6KDd5eCNpvNu5
MZkuMpWhnYlNDP/w27NWX9DuuyUBcM8dumkBJhGhEhZ38ARJPzxvtZQU6LalrtOy94imaqUTSz5K
K9AcSebKtet/3QK4O9LATQiOr1ZW5JjZNNdSE5BPMz84PLsBTZbZNo4KOWsyGWnRJmykqlHQJ9Fm
irE0/RTEo28dhm9JD5i91bS2jY2NhUERo8vr15B6k4e1BbwG+KOH1ydBNjwh5nkD+A++SYSH0iWy
7526k0ScrvjVdO2nx5I20YZw5IBq2BD3fX0OsxPMgG74b3UYg5gzmg75cK96JcWVXenfy4QaTHXD
zv9RvsHvD96nusPwkPpEJ/gIRl8ehYn7Schdxku8peGaRdn0l72Q34x30mvyzhxMSwfaKCt5uKFU
+vkrahpVpkSv7fEe9m8e4VTS0kVaF6NDCL/wQqt/LXl68MGf+xrFWfkpzl0xEMCsV5FXxw/YwK2/
jb0aHt31Xa+2vfL53H5dPGWsGWolhBaZ+OsYc/3AW6DCdzk1tsl/8ijOfwe2qDxirOuIwLMwyX1r
5zKbVV+t8uFVE0QUjtFk6xBE//yq4CJvHLh/SlBdL+2VcCCTz/QrFrC1KZspAO2qvlAs5/JHxCuw
wP05RPR7/2yXNMEI4KzHjQzT2tFuFSYz3Nx+libWT/GI1zgzKu+BdrqjOMWdbWGlNaf9xHp+11yz
u8LAw3tJ9/w6YC4IbeU67OpwXoKs37v5V9N+NlIPreVnSkcZ+dZnXiTehvrP0cY2ieC8lwC/Y8QF
G5zlcCRWqnYOL1G+5LNBUsME5A7fn+1Te6jGNl3dbPGpYzG+Vtxkl+YXCeD4lLTvrV0EGmOlX2tX
kSGUUTLzIYchy24B/ELXlFdPn13YVl2POwF2W3dLX3r5ZIOZQZVjT/rumFqmwpVe2aqR7EzcLcDQ
Kpp8QjDMR2Z0vFrAA3Wa0bdWPnwfcg4WmhjS0PPkwUkeBZ462/jni3JGUaOs9sM+acrVPX1N7Ctu
RSlQB3mphPArT9VvfbrOYafPNQeW6UdQBukzo6shCI+mnoSOBn68+JuJEn8nEIh2PDiwEdjN8D+U
PiabOsc0NlCye4G3m3MR9KXHBKU/xZ9bFFlHWkUcxAUK6Bw+yf/WtG2kZuLC7ISE7x4sDsR0NBKe
Bz4EvBqEYkVaQ72VeEQLT1VUDzw54cIWdMoABDBozbqVtjLgZJnNk+JHyx4PR2w9+8sQ+YWTVys0
ZpnEXIJedwdo1yNcJpSJ6IQENUTMGyXfMEBOG24CSqRdwjamKsZTilGGdf7UwA8eDKqhVwh4B+th
Pmf6kc+RwZcUFZDKyqUWBq41mgDtKK5ThBtV+wgYdXNr+uKhXLvGrRXo6EEnGI3oQx6ndXkd+fFw
txuoWZ2naRCm8RzFr5Uf4mxDh6x7P6YMLNAp51lzG7xp5esZ40ToUJ+ulCPDX4B5x0QEaPDaXdvN
WqEyzH3LciYlSUbvA+VdJIpjjsIadgP6MkSwv/PpTNqMP5yoYcolB2Z4r/HBFiityKD9ziT44ziF
a30Zh8YhOE4d+HjI9FiAanjyhI126odeb8Fc6ZCd4QEu5F+yaOdIQOUZcuR2oqjH75g5n+GF00Vd
iDDNr7SkJhpzibffwYxrXmkbXudwyyQtUI5iylsDFj1s+FbsM5Orb7T8EOLF93mc8QpIdmyXDfuQ
MoAJ/OTOh/1jDAaTyTOSutKvL+/6Uy1DKdMfGuiPnZwPxVjyTkM/HREnmXIc5kVZLJYlQM65BhA1
iVwjnx1xYXWMgHXpuB99HJf2jiz/VxkS9aI6goquyg0FmaElugdnS0ORi28hrixf9s13r2w7iWvx
p1uKxkLXF6LXWs1HCDijM4J2duUc6ds1Hj0uIyUEzhZ1+MR9j0nemt2kjF60+YG2m6NIBt3YfyTa
KQ24qSOUHAozqi1kU6xh+7d4+RAbxiiqAKKZHFnrtmrXa7+/LRCcSq3z0D6hVI9Eqgt/zjxGIs9J
YIKzeQv6ob8vQyt0E2HbFAqxFgXfb1G1BFHTVgO9OBKvXMR5y/4jKiK4e9NVBC9hecBqRNi0+jr3
FYydCuhBi/TT1bjMtiSY2Tw9wqNiw9keclaYm+je89A+hFN3YqwbgTc7NAWUaquFaxH/ovOJb7X+
oH84NPsLHt6DFAJobUlJbYbtg9iOm1SMoPQalthvjBY0By19ALpGCchlgNEsVAV1pmZnlWc0+Z5F
gqV9jqAE9H4jLM2IiZb5vTMn92QKOOZXRd50PkVlnhXK3eNWl3bqfvfWtJOPT4EuArduSjetmFzH
Jx1nMdc5Q6HvDXT0rFXtnTs16qfnKqb9/i7vMVy1QtayWDeLR/rvmC5sDqhR1WOmqQwlkV1Gyr8V
hebtPUikhoZDLOnMnfDkv3VpEsByaQMKAr+TDigZYxKXRWS/CgddPTsK9SdXLUqKa+MfCBCpa5sb
dKrO1vFlO6Sdtl+XrXTNQiB7wYTCU51hdilVLquVQGW/4Tt2OTyDNVQIj+Jgc59eKPMlEJq2bDS+
T/iSLAPPeZK8yC4r4zfvXtEb6dH0FFaVOQml5lohUh5R9PJBnvZi+A+9AxPWzIxSke0CNBpjxWPd
Heo6HRbuUBq1PO2m5MjxBsY+KDwlGPIf1qcZ5LS7vQhdPJMegD7u5h8zrM5MY42lUCcmmQ0Bj/BE
jMuaI6+nBhEzAHF4Jsy6i8EBa93G50wNd0IFVfQK30UsMVOEEo+31vBCKKHuAMdVRalDivKngPjx
2IFA8HfSHngJ28b9+xCt8/BWxbMulyYZV/bOHHAUBFHyNxvYF1ctAjRDfu6C+GRc+nl7+kgf6Vt+
iZxwft1OUd1o61SFSuM0zcCbgFqmCDufuQDxT+R7TDVZE+EheHkH6QOPssQH5lxOSBvZVNTPM7wn
zMMS1bCyCayfVa6G52kfQtsEonKY3edyCdNKXAsK28zpFPCkC5WpncUM2S/ta91x/b3xzvm3evkx
a7Y/XKOeAdT9U9I4UMP4MkKTTJWpAEbv4C8P6aua1At0zRt7bRi/vbvOz83kAfrkPILvZ5Tyabcg
WT/lRU/gdExicv8Y4FCDQUX60alfgOHaT9S6NXSjNCTJ2IxIpkISTJCXLHZgZt+6QaIOKiIPu5wQ
uUJT4pRAvYMQtU1YpNvMPlEhmJAxWepZUldwmhVzb0TbAtUTYHJfJ4FkSNTbFF34bNrXpgMJavGi
POooF5+DuOwx6lUw1wZlT2uxvruwp7Q5J/Nv/YOdB4qyFTkp5RlwHj4dgXmjAdv/L77GxyCWJTCh
g4op3jocoXgTAFNbmlOTgKFsHc+lDidXimTOD1djjWGQkRXOiBUu7gekEhouuCYAjsnnQZWBJRSy
CMv7EnM/faXsPqGSY5A4sz8qPUrm+f7RVI7cuzsdvAX0P2EYTp4az9wupUM+ZGapeRcEhmGFjR8J
iIl9hqFUXcUS17iOyNwOd+sFAZVr1UrrkqFxjgjIrCrVzfXgIebSuJ8Gm+6nB5vvmSBU7llfhT5V
J6bbSmoViMvTOTj+hMjn1v8Tjc/pEKF6zTxKMdOE7xDwh0cADc2q6JINcxs40AuOcIpyjeZlwKEv
OYfvCVXdm3DFsqHfJA75WjsARjtJFgYBcQVNwaGj1zF9fxGCh0Q5NGepaeC7O4dgf1Ah8onBRHgD
ELRwWf1PsGgsEdIv2l+rsNU9qK4YBiy9iGhK8TkLqFfYb7l+PXeAeWZSToWvxouJqDhkgdHLly2m
kBBP0ZCgY9FxHtqi3ktrhQgrsVFZzhqjRxyDdUHk1G1pRZNzgCVNw0ke4MWXjS4+FMfAaMgQeM2z
C8vW+jC/mZ+sR9ZFbLGqd7e6s6NryiFbcI6jmLQdVcUxyngPrvtfeoWb4jwCs2/zlYmb2ogSYpBK
9i/0SSD/irCDU6vORiWCVPbhgA3g67V2yLDT5BAPmIvHprH8NaOWvJdEgpZw54x9ULB3M9qMnabe
9UxngCF2biahpDaeYrDKs8zK//XCxkJH0KLINc7yROWoQRNvi3Ys8jANgQsX958jkNjqO1gpJTSz
i3wbpUphClWFb1ohi8y/eahstyPUQQBkjeHZFU+TB3jGeesSLFUfp7BFN9O/Q/0mXVF1dd+bzGm1
r4k5aQQi1dk49SZmnHBo+TcQH8XVMsA2r66zS35XWOKxnkK3xh8NVc7e9GsnTQ7iFEJ9qmviEDPn
+5mZGZcC7eV2/y8gfKeiKMXR8CzOHa3OqVB3fa1zD6lqPoaNI4sGtekEiDyxAZakXZb9G6HNvnhJ
kwosPWoHKiK7pE7QZNuLrBVHYSIuJPsIuSfFaja9tfAmJSbQ7TVb5Qw2DWbpICvYf9pktUgsvoZx
FjcxFpOz0pZqDbgV7mXcb/SjUl+c3nHZnqTHEod85YpuJAIcaexGIdFBd/A7BTQnNmC9gaT393KV
/ofnJIc2DSfTxjbzTzByuT3uId7Z4p9EO430N3Y0xy7o8Y3ogMEjk5R83NLfaKT3RJOU/pi+4TP2
1PR849UbAgUTG5IGjTFsVj4HEOBjBJsM8qS1OJCovUg2qFcA1ohbRWa721lu7tRVgY9hTBMHQLxY
BmnT/HwXXqVMa8rUGsTNXFPpYbarA8GQyuuQCUcsbMCH37OnzXehKCvUQxCufjnCNPVK7V4bTeKs
Jj2T9uRkIKasZvJVk6lUf/YZgdoM7VZ0gGVh+O9/vx+mXZtSlQFfvsA1ZzXOKkLOMjtwLkSPkQwE
IckVD3+zSiIyme5HmQMiY6qRUxjE+FL4MI3iPiYGbtRrgq+pymrCALbOKeySGtrTUAIke0yw/rto
lIZWLD4+7U3U+a0OyUsur3T5QygbyjwXsGWCswl8eW/weXlSjhXyhj3FMa+b2K2V9g66bX++mejU
oil6GDYKMBLitzTJr5l13EBmYaA6UDDnWEqC2lhouZSFlgoOVKCCDoYyrRvesGSQAT3bYSDyzM1I
anUspoWjz0Kqad85GLOLiDM25vLHcrX+1veGZlJiTsx8+ia6hA6rE5Lx/7A4sMoA7AWBS05o9UHq
M6rxE+vbvq9YxcaCbaZcMT7NL7pXM1EJujQhqZQCyAa5zpe8MeoPfvts4JPl1qybbAiMq79EmuHy
MWI1CzKOZTFqOy2kya870myNgd1vWlGXgBBB3Oc12s/FKwLDNIsRTpP8Y8+lVh2nAPB0H6SSC4uF
Us2C9oQtr1ZqRnpwMq2L8UET1ylHujfffm4gJZYq+abNm6aCV5j0fiN/NAYtyJT1d+b3n2U6qeiR
WZjni0Uyvb/KB/dg+3sR1qD+K7JhgEPNcnk1+TlbkfPDJobU/AzehIhlLnvW7zeCwme8j6CkzXv8
Jc8a/k3Yg2956Olgi/mGQ8bg24WTG7f4gIrGFR+Scn4foOTKjge0NuX1BEJVWeWuN3H73k1VblsV
Enaw4MuQ4sejsx2K+mvXu4dpVGFnysm3if9hvgvXKwsPLx75JGGDreCsV6XFP7EoTa1BZSNCgRi6
/RZOfwNd7U8L3gWTuWQHkYhLcP1pXkZvDBzN5MevQOQxiviDwp1ckVlZPHQfSmQgBiwvoyDm+kTA
serRH8S7m7rJO3Uva48+as5Bokd4KN+I5crKcmcGZr/eEgZUJGBlUdZ3QWXE0AcAbQbi0y20NWmy
X60OPUofnSZieWu3CrEtx3ouadmEda+Dm2KZWYf3qUw95MirmW7fvYApFlS/12Z1VtnpSxHHL0cv
hAUATXvPneIFUoPiEcWb1ZhehDH//R6P/YGpWl2VrBhh4xjjuHj12rGOXv/DFkRpGuicLFmofBmq
Yi/rCXx7rCK32zv1FJ/FEUA7/6C8L5ZZNiurxZtxiqre9N4GIvXesVuMEszOvh/hXT+OAaJsGKzD
R/q8SOX1ErV+A47WyGM4vbmj58YV6WGjTN/IsQ9LjQh4FD6i/s4aaGYpIBcW5ewgQ9XFmlLBQ6xP
EKgcudObwrawDYSPyGnd/kXDMGvIZPCK2nLditq3InULYwkOkdW3gx/L2pgkXhSVFTcvi/Okdp7y
svZW9ce/x602LtClkrWIlg/YcYVmK8rhDcyy1tEfjKWgW0UO7K/BP05vQzorzZ4YBED/1kZXj6/q
C7ilO/oL/JJ2RWdqb6YaRa8D+bwy3U04tAxiYCbNuNWrTUm453ZMbociubN/VTSj8z60o2h3cKeO
qwzM6TRqdjNGQjB7T3u+x8aSJizXav6ZcaSALi1KVx6Cf7KnbUAF29PDCeKcKR0CZl6tywALakta
NCK5Pul+oVN324cOQlDs983zBjYeJWmkZKNBcy5Uq6CEqLeevWTPRbxjjbZgM8mW4UOpYn42Vmp2
fmZSG7sLsQTYh7g8wogxpzLmD6gc67Jgk1CC5vZ9ckpuKaJygS7Fp9K81Z8CsqqhKF3wI6fxSaN5
cLowD1+ClIAFsMLoG0mjfWe1wSDAVe/nBuG2OEobIZt8Z+MftJhGHBuj5OHakK7NSSsogBQn5WBf
Ua8Kl8WnQ/0euq/DGX31piy3fO67d7kQcgwrWaUhpVyh2ipi5OSouwdX3Jy46BW30LYVzGzXl2Rp
n3Yk5iWyIQxtFf/6tycbjwgUUEwHlSP9UVODc0RhW3vI+kPr5MwvPTOypYQ3gIsG/zTDHl7DGSEj
4Lzzp8G7VYJv0ZvdYsBL/cuiGk9+zgyF9wi7RfY9iKaEdvA/qMg9ikqtJRYgisXBxUQGr6OC6frO
xfW9o1XvcBKJ6XcpcoogHU75ZOrSwlrFIwebbJyKLQbc2VXNHQoJlpVEClgfkbPtr133G4QX5XeY
91pK7UH1LS2P4qzIcicIH+wa8PaRDTQexLR50SOecMAIgPnq+YImI8/+ma1doMhtDI9PG3Bre6/l
JHOWnja1QuUHs86wwMdoqIvZyaaupFNh645X8E3/oeAg9V6ZXK/OlrFYlezhpECWApYugeLdjUsN
M837k05KJHmjyeTgG9IwIq6CyvyM7THPL/KFIVmXXUPm2vdXIoLkmSGbB/SOZKZ9uK4k1PNlnR5P
5Q6Z+6amfBEZ+L4Adbuw6XrIUkQpQ5Z8RzLKRW+w21DTOHvt9s67mEdG8DAZilbdsc221moKkIcq
B6YJmmTd++iUHITOFeIQE4wTwoukpVC8h3TMGOR+iZk7nt/Z1zzUEj16ikfQbryAlXmaXOlAVMNb
GrrsIdhinjIKIzSPqQ+tsBipO/xmgOd+z/t+dhEXXtWSH99pErJ2C1Uwe3ODaT5DyME0PYIsJRON
zope81vz9Sk48wWtUMeCfvQkpvXMMRaOyXtLuSP29FhHca2wWupJFsiu+fbUkrRW1Zi/B22NkqiW
53igb4a7UTkXJ53niquLDW5iEa/+jIZPuG0gmeRC6f6BBn0jSpcA5lpIzcjlq9llCyYrKKoz9gqg
TcUNdIO+TLjB2Y6UQ6Gn+KrXlSBW868vmKW7a0G57lGedVJMiDgKb+aIp0HvMpg/lOSoj3ougs61
k06zTAFrn85bwnneqCqwe6BYIkW2DU7m1QpQcIqnMJEfnwFt95oRSdhCBbr1Ihck6ktAEAM9481K
TPqSDkKbbBmTmqrzzlMIHTTgtxuR/cmoxcKkAvIgy/qpey+2NsJLhwQRvmQtmgBypG0H2ZvLXVA3
0w9u00HHqiax6sUfknAie1GB3HnM13jwv8LSYyIC/a3e/h6WEWreql1DMCE0Z0GsE0b3Qkw6R9fi
hZDVXFsvF/5N2Mhkyjxh7rJ4Wv3R4gNZwM1Bi/9a6cGYPhgY/0Ge4o9mas/cS7MZZn7Iimbw5iBC
C0XMeiHD/oFpaZriVv+ZeX+F7QKHB17Wc92vDlxaagSwye8wg+RDNMs0XM/RmJl8iU8lfykzym/9
eMCvgXklUiVqFzWfZVykmORd/+1gfiM/82FdVmfpxqYDh5JFv92zvv/c3VtYnVu2A46jyPAt5W6S
PnBg5BbQABJ59y1CeBUfzFzPTViJH2nkfSd3XaQxiOc5kVQJARiUDwd9QDmLet5BP3mmhD5u3B3a
BdghoOpOtEx5pax5By4rc5EN/3c6AeDIU7unTVzTNyijN9nPb9niwy7xw6W45gmO+eb/xqUa9kbB
VnHXlDp9enHjkO8sevxQH4g8y50CXT4oqz6urHwmFKs13dt/Y6P6d13G5nyIrfHfr+FlzMwWfp5n
For2kK6kRk/6O/JP1ufWtsHO1b/xh3i0MgAD4MSo06fW/88Xtx2TMZjf6kHxChP+ak9+SO883A8Y
4slErtD4L9UYs3KlU5WfkK8HpLQaq9oc49AtU0llsUWreHyxSY9SnaJ5VS4ILc7hF8rsVs9ch4Qd
q8chX3tnXgPJ8W+fhAEFwToX+wBkJHbEDQtm/LYEbUl6AfLe1kMc/O7emsbCtFVJC2L+9sHFL2SA
JgIISIkdyVFj1kiUed5VQ9t0I285MHyoSwcXskx3yhR7G4tOurd95hvLpnpjugCd0e54xUuv2D7i
sY8/foRz+qARYkZGzuD72k8XVEDsDelBXHQ/WpENsmRtu21J+/L25zH0Kr6P7PyhvFtT59jbOGWK
JowMy/MVBD1sXxPhAtqjRCpzHTfd1SIol76Gt8ptEUNzu5KDb04ZOzgPcQu/sPSBb/CF3XR4AYe6
JtZU9Bm9YpuVNCJftBnF8L3DKiQazcpMqEiMDUuZFSNwBKDzMcqb7u4SL1dLa8LIIOl5imYbSwPa
ygt2vxpGbUE+ZXrJ2U5DyTEGJHaUkoQPbdWDAf3+J2CUZUxaEAhzN5nuV5lVS5bO7ok5TQimcyw5
e0peShynwLapYqz3X7UrHutqvKI526Tw8RDOf2vp99ECc1bQXFMMKg/HpVldkV/fjvag8q1OyEqy
VWeKZdxOqXJrDJW7s8jGQhM2NA+thAxReG9iFZv2NiGmRpSB06JvKWvsok8ukYAlESVwrxoY8mNr
hSFgqvzm3e/Isl8OOoRthmSGUfbBRc3aIFF+PU/NvHauMSjTBGPZHnDRR+W0CyhoOD6k5gztazJ1
mvrJP2+nE8HrGFEc4Pl0PH6tC/T8L5AsmKUwypHNhUtkoO0VbU7BfJvpzI1JKmOGJyJ+4Og2kYnL
YWbT89C35NUditmcuvktmpB6UiMHjMEA4UO2p36BPYBSaakLse4EpBBsv8nM5+Mc72sBQ2RFT8ew
gnE+UkW/ap5pEaFHhmNN6T/ApDBYXlKL6mTV1IsVc2iN/nB2EqtLjUUhBCrdSHGzOu+UtIQoNcSY
5Eso0xxUDuAauAxgvJCeqr5CHFEMEKxRKSKTVYbOo25Z95XJ9xNS5gAZ7KEgHxuPNJyYLE0ksAcw
EknfyBE6yJIIbMaCCCtOEBvWkuu7Sgyk3OlHZ4b6VfwWcD6CGzqP6ksAMf0XlmW45c5kHGXQKZv9
knyyzZ9TZbBVLWRKNptc0feyBosw25suwm7fOV6cPxrjXV86tSGp+Y9jrz7t7eyWlKNRpafnS6hs
po9zxH7CTmMTR25I+jU8j1H/Eiir2XLHcw17pGEsXvlqz3FTKEM7sGrD9HYm8QytDqzjjVs2lXIK
+RBVVJ5E5+qoSk62Dwvrd++d35YmspOJahOiIuza/Q2JsVCNost7iGPa3Wzb2e2jbQXclakYVMoX
9hR8vd1B002mNZBGlBr/i9myI6Mn1svoyfxYusn2Ob0SBWZB498X7JXcySU9EQ2/0gNCsgpGIfzR
6sZQChyuDP6rc1ngHL8FF5JvLu/gv2LDSkh1tClutx44G585y9+qMeTX/y33sNmsg1ktghk95LZP
TM0GbjLJyshBScSeeZ0ybU2xjalVhaPXbQ1NcLK5l1K3xozaMHSBHJjM/P/exmlveNG/cN5wQYa4
ljZodsd8fZ07DbYCc2tXFq3I8oyRtirNhS80K2OnqGRoDp6kQ8X42V9+v2U5FZeA7BOwdY1Vi7ZJ
W2R5kYyYVQ1GYyJImhtSIL4kTNsY0HJMPFBjTl97mzOClFiJeSV5+JWjZU8HR1sHxEcp2JHtpRJM
fnJS4uFuXucUbIjDm2Ikd1QdzY7fEEHE7+lIU04VKVJIk3oGtdNvslb8rAgk4FFtJL6/uIscBU3K
brv6l2tQgK70/h0qVgQla/IkbXgjJXQ5I7TQTzCwXXkxoGubyG/zohDpHAehcqgz9MCvDqp4kA73
WfI5AXEaR3sQ0+1A4VaAcyEA6LIUxfgp7kDxmiyhSKnYzuFbfxAtYBWyDs36gztpMzXS3Yb1ymP6
koUyjimJmJkVkFXZ/MCm1jTtm4nNvZ/TqlZpKpwAXDbNrAw+kGhVt2Ep8HIbbZOnWpFwYw5IY/nf
vgD6zbbzEcjVuZjT3DBjN6Ke/Lrte6xZyupUt39z5gp1Zwqic0ga9HpzJSuxyKuQkdrmmokaZPd2
w5MT9XRZ2SwKhtsDIv8gwltO5j4/3PpYFIVmu12+wMPMJOFw30WKoTJBMMaq8Sl+kVehBsDnzCaJ
uolhYsSiVgnJ2Hoaxm7DNe+DoMbMXBItQVGULcFEeLOGwhyh7cMBSvjyIu6Gd3oQ+n+oQ2C1MynG
q60wTwFXw3lSRN+5uNHtp6y4QdGNq9ilcAiGglpbOa+SQgmAQsAyNF9ifHRTa6OwXHZ+88BLnv6K
0JiABWV2OWK2zyGCcDcmNGC+IzHopNw/PIeDlKsOyetGHSPR3a1MhJ8NERRgjr200726i7VwVhdI
OobIuh3eNgVpv3IPtbNAluZatfsyYllnfT954eiqSkzFCw93ypxCWKByvZeF0tRuRTvIE7oN4sTQ
mtj1kMq3BmloDDm5KWL0lHaU/LUnuQ8sNl8I7lZ9ktFQCsRGRUGoXgY5c7zWZyKXq+qlXe9bkJXH
yQjC1vKWLbF7nwSJLq9sURTQjlWAXNQPjhgMMdnS/+6UDJG7jVeEZlEJcn5hAoPHtKKOVBKl19eI
Kzjc742jDFxkFxRRqKydDy/J2j6ZvU7029g/ettbJb6NZQs5pE1IWbdw96AynPb1V7O64vXkZ+mH
R0i0fJ7X24hDwIgJAfZMpIgrffZaPt4SACdYRJYTVNrf6rp3eoOE3anv5R2m8RI9cHCEuBe6XQjp
VSHY2DQawuVEL7phFZL2M4Rptjr1qCxo+3FeXNVtF5tge3x0x0o9lQ3WMxKvwZbNnKBhwzDP9jbS
5D8aKNDu3MTDGx/26kyt8bA7qu7FtBT+abkXhVGMxBCloCGNC9tJH+HsXO2gQD9hvc0LZDuZKsCc
CLXLBuRtC2YcyqO6sZUp89DJz4P+ayLCvTXFC/6wzYkMJb4IeKV5pwFC5Hc8swSUQGqUJeHaMdAl
7v0rz+AKz2J2Ydloun18TsBVe100W94c4TecG+XnvYzBt3/TxjI2Mg3bH+fNI9D3DYi3niL6jEZe
nSL3dQ1v7AoOIkXixr8D3Iu9yXPyUw6HdSW7WhHd2eb51bou4CJ24i0mHdXFrvvOVIqYOKlkrm9e
+XO/L9wfBqA/fHrKPFSWQ8nJtdg/ayyPwFyE7qsj0H+8tP2BiRAo3ifKiSBYVRxmTzWybzKaL88j
7kmwzTAvyCQ6YDRBosCOIyb+QvpI+V9vqEiLuxcXMTHBJ8oPPBxSWcgSBfmkhV43M7vvyOyfGztg
a336NJaKoSgg7tUH9864e2todYdRkiacM5xYRRE8YKrcoqp1FMySHGTVf6nwxQpFnYnmLdqWuR4o
B/jqMy+58+fywiE0Ix7ws1jWwAJ3nVTeoR+F28ztOQY1whSCR/G+4rhv79SdEEFsNmorGkkfyH4I
wZLVgbF6+ugQ33KlvXngUGcSk3kBAaWOjTwUCD3xHx8qI7EkjM+Pgvfn6o9inRmvqD1xnFU3vL0n
+qhQB+ORLbHSGjVsK8noKPF3yz6p7tanae/EqGKjgo9n4pzPTt8evBr2sRFTnS828UlrGPxmr/pF
tyjqU6LxsSShmFRI2SNfqV45VD5m8nSlsTyKIC7GS3V+3RSS5k8a/FjoxdIdGX6XXh29yYbDO9/2
CKiN0q5HDphw1Xnzdb5yMr0qtb9CcB9Hu76j4ivJfVnKiD0cETWMHFhUGzQDJ9YwVNE6ozIX5Oyf
gsO4dH/DTaHVTlqB+chkLH1boRQcXKI4P4/uMdQo8WqW1ZSfON/NvNH+d51m/t4/ih70MIKwd/VW
d5HChuyEjWrfnsBlSx1Z4TglOxPxMhfDCxnfr3Qz5z6s8W1jURuU3aVTZ2cqgHFtWY8n2QPPS+SO
wMGhGq5IAWMlU7W9Jc6SbuaSsC6BkqKqqemgkyw7RKiwGIs13Du/XJyt1wCvqqFLeIsNYq7Mmrnx
ituKRuWISiWPcR7qi+DJZZojp44FT3h9nroZXv+K7wRdW71djzh0yW/zDB1uP0gNpx0FYfpEqqq2
t/gDXIJEdp5jyoWbAl85+S/XQ3EcEFpVrA+cKEGqaFujfTZlsGGfE1zsC7Uj+RP4m5i4Xqh1fj6H
ey2R5BWEuRDYK4qeBiJTCtqyCLmv993JO2AuEvDeMLlmtS9xW9rWOSUx4AeRlfzSAGfvOidtdOC+
BWZQmJxPKR7lqL67BO2itZe+KKnnxWCsYe4iomf7oFURyumkc2J/YNxmDJDBlZ5DV1jG8f5KLhtI
3tUD9iaYHs7gp4c/K2Gnh5GOYOjiUB7N43mMVzWgcuJkB9NiPoVFU38XYXqXoQlXNJN5CEvkxpZg
aorokdJ2U5OASr5NepEdfg+PG+8DgHpMOogMT15FnoZ5bq+hGis1jNhZxi1BYq4lTI1movmHJJ6S
GRGzXcNOVtBRl/+7xQThWGM7YUpNH1SrZS+CrU18TnR94cBNZjcUOst+zd7o5RF81AxurgmgyR3a
Ip5wUxLCLSp/FQHZqRmQS49HtrCZ4L9pKGCUcB8mwho7G8fG4umaxDI4CQovvDkWlakpk9R2f/VE
wW2Rfx677U2FTGNUbk7zR+iUjLor9fYq4fH/zkLTf45x20cvJCEyrOFWPzCsferEXjt6YAo9p7QU
Mkrz6VXXd9jXeal72/CevIYbTc+fXFoeYRhwat65SI3vNeY4LQz0xs842lQxwBKKVl1ykvOImouS
gOa+MPzAukDx84MFVL+sesgpNBV+sMfnBa9GePxk1qCCxQGeaxkIbdP2i6Jjg9etvSRyj9H08r1N
sW9TyvXNPAdaKZQ3DlqIWtM3Ht7WHGH2b2C0sb/A3uXfJeCBJ7vUwOqcl2kGdNer2GfDfTaRX94F
EHpL7v08MOTl+GTg4VT95Ycd64e1/1Rp00dufKROFVYBCnCRz/9p/YYCOFXCw7+iRRmhePRz5nfo
ilKACyUw02HaSbTH6FyZEnWy89vlNi/NU8s7ZV9aUQCmCySp6VXerUf7QWhOoXCL/fZL8cWReIbn
hIzGhG/2aTYOn14s+ulw7SFV4VV5z+YsFT5/V7Y5rwRlqfxmu0qmAUi7aXBQSMOveD/inF3b1ftJ
D7BBHPMMCCnq5Mh/12/kJZuBQbhspU91xHzbVC4HyUpSx0srrjfKu/tHE/sCUNurP2rYFyCIdbGK
sJWQ29bSos1uiQ3gFrbko3N9Hh/jOCSSzC1iMyN+xw0mj6JUNagVJP+Sjjrhg5k8pCOVeSD4c0yN
qcFQsEbg+/27PlyloM8b/0iJLvfNO2kJCm4y5fj+pes1LbGm316XPcitGR+C7h51ULeuKPLyJwaB
LHc03cAEx/h4eugsznosNVpSZ1m+qyEgR+DI7hzRHKcvK8F7+wGPBR3eme7n8McwcFS909CtuIzw
wMnllm8Yo9iL9c7DxrI/vDd7B+3a5RTyPX8EcNmrnz40mXHyE4GX8BqrNCG02ePKkiUbQCj0drN2
jBVjtlLQp4ufWC4musQuZ7BpbbOZtnPI5yneD/6wBwHoYdjXKlLjZenF+SnKHPal7LyFHE0/8UCf
crpaFN1CeAnxL/KdtUSbmj72kcH684n9KqSiGQtYIhZ0k99ydGaZ0bcWsX9BjHFXDYkUjklJBoge
sP+ILxBqTycXAgsktiFkYjTn6e2qSzu4kqA2d+5wpaOAe6tm9fCG2j9RPhkx8/YtF4lzIjLE9Dzi
siIHdC+EdsfRj3TkIpmm2MGXLGMI61dtbfFYxcZG9nStdvxoXjpSbTMm3aA94waC9YjOOmU4COF/
Oi/O1OQZW59rHNFWBFiBSpHhNJpu8M1ujIO5bAkBVcqkQP/W8khfbvZLIudq+Ov8uLh3BUvm5hq+
FEfExDmOQ3QBnLMy75cnfhqiAxi+bbyFau+pNNI4/43riZFjsqo9N95yEF6xLVLj83/jAluWFqQJ
zfXmhGpLrMvkMvMPX4UAMyvTaiFzfgOSjjtLEmkPsvfRHabwacS+kt4Fv2k1D1mbJwiksTL3Q4QQ
EJaocz6hZbo6p4feTRE0GcWSPfGUkTKN++7auUEu+D9x4qHTWohD6Vllpvtze7fGGv2kZ5BPMp5t
U8bGI036bZWS37V4kTGIain5rdUNCuCxPLT9xQE91AaLTVBvwa4fUjw4mRlNH9A86/E6LbW4iCyd
8efrAtTfy0lgMZXNP1iHfMGURN9yIdVQvbdCHk05WXgcIV+hZlBxWIa93N5CNA2dLmzmtybWPo4y
4slnyBKsQUrtHBX/iWAyI1gUhopWYQZtBFHMGwa+kzqfcfVQOD6DYLjMOWlNHgfaX8ixH5CI/v6P
RlOs0emiXzS9HScYIWecSzqfF8qQ6SMPscZOpQ4qF2bNwAB9lSigBp1cMUdUWyllfy9dybIh8dew
mVJzBio21EoUlbhHdIhqRwg1wItj0QAWiSPlDDKtp4XiY4Y8EJg77gJFXCEecMHPX7x5vRH56prs
sYvqMGgbQfSfJ5NQ5XBYTjVGaAQn+GwKySJDsMMOTRBpeEjkjZcDZ2iG+VHb+mTgfyyc6x2sY23d
u0Tq/oI9fWqkv/EWS05juKqOdW3uJPTdcDKW32FXvZxSOC2+zyVoa7I7kuFAasQkzEEmh6XJdaqd
5ys0SGlZNlKKm4oA4dWFNa9afhVQudn7qHHhFDDCeab4O8cufiE7zFEMiyJ9tvI6INxk+AqLM6hY
q1+gyKVYsgwveyK+0iGwrfI8I1s4KmBs8JlOyPwlSNevuVx77ZIgStHaJKaah45l73C/WZOqloaD
EAga/sJW8QUThisamAXQRp51Cf7NkB/AJDtPs8VVJqCndcflfXphMyfz691h/+S+DFP/FhtS1/rW
q5Q0CwF4Bc9l+DD+ZO48OAt3idaze0Ac7s0vzx/m9qxdegCkNIOAqhrQtgLGZyd8B6C6DVemoWi6
m53MmS7Z3HAaLp/Bzra4iVyxMDVfWY6RzPd2Fj02YaMlJpuk/euJ9woIfBbYebOSR6SK+qRWSPs7
BmoV5we+0aU8ijOcSUEXikdptzjwDWVZRIixSosPhaPF4vIHHgFb5GcTZ3kk3+/F0phHG5J1LVq9
MzRV9JgH3DzJzbfd8RfR32NS+a8cpW06d673eWa4BizpFKzS5l9aDokCdt/LvuBlj+JccWdJox25
Ng1UUO304mtJnmS708gAPRTk5QNhQQ6rciLsReRraISIErB2+QUb9etsqdo6P4SLEbt8UihwYuII
68F+Ow8CeOI8utJAM629SOpIdDhaVJxaUZSUsv9GsaQfuoAjcm7A7NHrQUD19n/yW33/5VFOOyJr
rXLk6jtBp2Ebk4xYhrnGD40M3Qg7GfGdGwrLutI8/Jmgh1cb0faTTX0/EldbTqsaxYFprvIQJElg
3ne1VJP4zSCn7azlb/R/60B6GurZbF0IOmYn6lhxzRmiJ89mkTo+/ZA+G/4p1n+IirysON9HjtIU
mSvrvf8w3roBQGH2BLtOBVsWGceKTHy8fthge0FJcv3NUzBSWX60Jhz9iAGq4qReDYFcewOwOsT4
WksXzQlm0kkrh/Jt1XS4wLC5Uq5w4pXn0EH6WRd71967aRv3GfSb6uo5vIA3B4ljYNyfuk89gi45
o0iunnPhS5WBK+n74kHFVdYMp/mj5dekwyPOPazVPxntAZAaqfD3nAYG3yzbDPh4MZK5IHeQV+8m
fG7292fkd5LwXi8B/RY6znQMU6JNQqFZk3km6ubiEQ/Bs6AOdrFQ3PBoWzNgWgxrQyIGhoH/RNaX
EkWYpLmQUkYkmXntQVjCLq0BNLpRPW7oIKom7MyHTwODkmJJEG8Wg9ZnTwqNvepPCKKxNjbqgB7u
RtqODXzmwIovF+HzzN+hETBWp2xKEC8VPlztfBnBxC62QPe0+B+zzoSm0HoF5l39MpxqOuz5ikhB
h+ccOK+OEluPDAWGtAj1lkLNl9RGiFfX8Fs694w44+6TeB/U+T8myMI0i63ttJmZc93wTmEBDigO
CUxXzEaXrQPobuQ3neUGX0HRL6lUDyyR2AYIJ62mzmq3Fh20yNif5AWdeB33YKv21nkgpL2gMMCu
SxpKUccYmER8FeGjHktI8QTM0wIW9Z//BxVUras/1/sKfwtnUJNXuA43xIlkb2RnqlrU2rHImjPb
d4iDJvDxfUskxe6xhbccAOgobip589amj0r32Oe+MjlGnNCdrHWgLGgTP6ZflVBQa10sXQosbUtu
Ub9yOl5sacFVqJoM5LGCCC0jNZbfvmEqggEiHFIS+UB5kemXZPOQ5I/iXdl0+Oddj0eIN1881wom
ssIPF3aOwMa/qxRRyG1Qc7/QbTPmVO6GZSxCIkpi/p9Y4dQ6tVThn6u7RRZyqb/xtE3qhj5gGna7
RiFpKWommVAw8cDET55i0V9MR0o7er2p7FQ6y0ejaHkPq3FuvjCNtqjUIbnHPHnd1mH4NNjDkxpo
2oTTeIxKHr7Y7UxWNo9imfrmluFU62ikbA7JdUcZ+Jvf0fkGbNvhsrDHP0NJlZLH0Ieqm6wnDO32
xY4bjyWDCDErH+k7GfAZQVZLcofQiiSNTWiTtjReuQA7i1KkoKW2nwpnvIDPEVJ/oR/8l3wmbqLt
VvV4XZRYCoQ9Xa8yFtOAE68fGBbMhmw/1wSXchSNYl4J4ICKISW8qwkboOQn0f7qDCHVk1u+rqKs
8DXNMF1igcM4/v60ZEbeqLS+E2TjRZa2f+eLzznApPPD6c0ji5LS82YctQ9FqS7ofMvfexxVw2xl
8YYFGG+VxKPU7KEpjYH05cYqs5UmKTgE66LsGKw3d9n7Q1drZjOVR6X/KBQ+9qPmIYudGakE1VTG
yxQ0pfbPr5599TGbO7/AQb1RymFPX/JeclboeN0D50hCtcTAyN0o59mY7QKfRu7Sw9LNCXjxx4Hl
aXF5t6//VfwZYFIzq/EJ0jPOpJlx5PqwnHkvyVhPHZSkciaot4t9CSNPkEEey4JWOnD2mT5pLfb8
gQlTkhZLOlyN1JCfzhD9GwQ3fbt/RCLtNU5EuJNseRTnOXUTAWRfA9APClwJBeF0pOaUkYUMe8aP
TYuotL2Xfj7Y3wHvjTUnxIOMlxuE5uRtyHn454iw/ALHmjuDnXfxqtTwOD5Tkzfcv7adUri8BkF+
uAACgVygQns6yYADz5w28ZQCBLaYh9QdPr40uWAcbc4kGLayQQqcW1SFWjpv+msaahlMATdrOrA9
yJalOI8ZBCub4jY3PN5PBpiQaTF6BL1ZSEnZR+lxByQmHfv+5alqYEchcQT9C9jkTemnvhNf9Lpf
ZyPzBp2tohLSbHIWn03oYGomHUCteYPvMDthiLgQOiY/C3274qQKvHO2k6/gy19gqFrYp6yzZaFN
WuAqqsdf/G4UqxWc6mmP3Hi62Ju29nbEY9UycGjTxU96UzmGanjkLBQmyFZhlx0pXzWNJkr5Sq1Q
UhhlnbFyTc0xTkLuWc5SA6Xj6hdcf/SBSwFpPk2H+WKPc3y4j9OdgvfK/1Ktug78a/qMBdpGQo96
G77re2KBbO20tA5k/qZPbbpRftFYgbCHmVKEZKmdTlOuKkSJlviEwhYwqEDCYHiDau1xh8UbAVRb
I2mBgAsPf+08v/DaT1mSFGDO7eIgRgRCUKe5PT3ssQ4Rzvy1onoC9jGi6Buer0FvCGR5dBGE++A/
+di0HmghQ4QryZoP6VZxb4SS+7WllgCjqvyVwrPgU8U0KsZZ8A0LTetvKYQZ4AeXmqT/Gy9alnBK
wnKqhsjc1xeWZoRpde6mx9pfbXICy/Q7OBF+YTsl0L3+KvKHnt74PWdurlnrDISda2wXT3EVhdAr
39+nAm0YFF/ANsq/R3MmNguvREAzKx9uzap9OMW33/M+yVLtA/k4uor3ctAd34hKIPjQa6SA2PzM
cxW6EOsfTRKafjyKTiEwJmI3py32jqIyhNfGoEciM4tf7bIeEHb9etxn0It9Oz84nMkfFJP3e5tJ
FSGokuIeimx0zFSmx7J/Mv4KzHHZMyr6y07gPrLMVuU3NY6aNll6p41+WsZGWxBlMYjwpVl1dFOQ
aeBtTXq3/+6/XxuZ6kH2lS4Tcdybbq+i8DFZmamHZXuvoHSLaKks8f16j6J2o+60RZKntxO8JC/2
rMUMEL6NjHhJYATHm19hi9z5izC95Yt8t2L797wFt1Klfd5l0QtWPoFBEC1UeW9Ra29rPFIQtXcW
alEDeu5H5ZIFWrODTyt8wil1Mps9d1fCvSkJ+6n+4Nqye0jCGbqnEYgd9MwjHjgUevOm/GM6Mmi2
qamKHEgGEgjPE+/X5sSdm646RnY0eNBthXBvckQathUFwlSkDn9xD0g/7aHpOfv2SvgqSdg2TJ5z
anzWyILkgF0WjdfpJ3yiYCLYaFiuf6kSQTPnnJBigH3NzpL+lzv++Cz9EO7VnCOamAJiADBUZIP3
Nwl24RHX96WYSP6cc7C1amv5+ehwQ1guhIb4nSXmIid1IVrVTWo0CjDnu3rr5AIviuDDqv8qL7Fp
qxsSkec2V4pFEjg4CWsi7/SIy+MFISZ46fB08XeZN/zzgfHD/eM8Acpv4hbwwQKebc5ZpberIwa/
g1iV0cXCM9bjB5dhTtNixE3feTjw3pQjfx/rumHZC8zki9R5tN4u4V6vTIHq/kvNQB8zjcPZh+80
OTqjc/AmezEb8jGYjzwr5yHUaLwCW/NG3c+8WnfyB028dY1UFQjFtM5Dzd+BmDTHI7yxjP6xSZfY
Ct++IHzs2YntfWGsXgsf44KuznwzF6MKR1wyumYyN0AcsTEN3pkUB1uuV1KgyiEIoBY4EbyBiqnv
3QtZ17Xb7LwOTY2VeCJoQ6C089g8Hr12dLYIaNL3euW3wSRtLQGN92eVs8LirO04UzIBDDKhZ2WS
5bklJOI95D+I6zyPvWg64/lYrgF06O8TfOUIBljeoO2w704h8RAdoomUESYNkb5PDKrv+Op+ueq1
xaW4KBoySIsyf94K4mRqYJUn0c2dUVC+Yxe5qv8w3BykhUHT2nD7YFLbBfvK1Q4Xgsi+vpdqTdfK
JPAV//ArY1jkBoQE3MUWKD2LYPZwpIEvwcA7j8FNuoKu653f8QoAO/vuNwHZkPQdGbuqtUmlYSNC
PVAYdQeuy+RIAhkoJkupyN1n1t1oYMmcGAqCvY2MuYKSQcF1P8jCeiJLrO1N/lQPD/aM9u6oXHI1
B/EOOBpX9OBY7uqnc3n5RBQy/ts9FkjrX9rpJbs6rQJXi3yYKbj1i8sSYPmG2zTa/06bkMrk8wRJ
uxJ1AlaYKoXJBt32swIjaa/Cjaih3SKrC5WlrWcj7nwFJQSKdFTn12bLUbtnK8ASWI8p2HbpwEVc
63AKfkfkwAAN/9KsiZn0b5FOsaNk1OS+Q4baeM2sqs4UjTD80Bc41h/BJJwKsXnPqiUwLuOFRGLj
9BINz7uIP8KxB30dgwAUWQAFyIKGgxL1qzoR9l2YbOV/CMkCi52GYMjR/C7UJ6hKfOdc0QFuWZQp
bkLlrkTEInbGXnjLoZGcs11rJp6rT6myajOGodCGOZcECJTaEMP7a3cPLZ223CiUM2odfvsSVi51
NPgsuKOEU3DJ5L2sJDGezpOZ3t0r/mPMqzONk0FpNGqBom4RYXZk83IJy2myf0vS1OzuIkZDNor9
bPJLmET3rCq1TMg+xw8JoogPsffx3ngGsZsufy7WsnBuogfdZgRSqWhY40gKJerhXGhtTf6+RR5m
r2q1YHOPlWBZ2mxSQAF9FKcFOMDpHn5BMgc4IGIpJRx/gswr7+fR0NXdZy2O0nM7EdASSTAk7ncA
ekQ144nPQA+fTEQRWnWR+WAXkfsOfnAU+QalpL9UzL7mwz+ubcy0U0VReoodWBKd4+uVKhLjaHPk
zR1JQ9uj3FhrrDejiH14yFeLdVnnfrKwG6NJ4fOZc1el4zsIVElb65a2KcBr7Xz5Na29m3reW1gL
yMvbhejkHf8/Xv4I3kQvfkCPhNA1unK7ZHfixmrz4HYUsHe/sUPIxy5AcRt1LadpsR3UMYc5v5eo
c3H9A8F/eCtATg2c9+klRbijtW0wmGfu+u2tJwby13tMQlgp1gBlo+hYs2VHltGvoonRKAi7I0Nb
4DzThYIuXuA9WkzwNA5ZnOaq6m/zZRX85DYBjbfcya96VRoWHWeKsGT2O75hyatgTc2Hs65o69Vp
YOA7qOKA8zHGR2qIsDrmKX5klx8Pw2RZUnqfnSBP/bpfBXOJtx9doLu7mP6GqB6J/W+8Tw4KWbHA
PSkxMyDBGpK9tL6omVV2IoGca/EB1sTzZqPKwZfxZoCb6JZj9cR1MR5fLyEPYRYdLl8Q4uVJreRp
AKKczis5WjgghtzUwc1Syv6ea6IoalLSLXmWsFS0KM5ISY1UrzRRlTGq+xFm6+mtGKPJtBr3ta/+
M6RAB9q7gETWQdIOA/hAbu3b2IJQTJmynTZXEYk4y2gjuS47BNbfnQ02qzJ3CYOZV5ce4U3ii3VD
WC0JmDI8mklMcZc0xct6mjVQeEGWFr6lHBaqiEFHSPmaB6MCbwn3gjFt1o6azf+J8UKkiya6Fu05
DSfLv/9gqlJ/dQAPzAPEN5hQT/WR/uiNG9kCHN9jYoQGmHPt+fXxsQQasdzezbbJ1/Ozk+Gt+IFE
XHxAM1wfPnz2InkOLNo4dp/txV7q6GoDcTlA8o1JmTi9vYyv9Arm9mhkgB/BbDdVnYfdCVREA8jq
IymTZW33uKkZpIPiv6eRir1qU5W/q5AldMwvx1LZNNfHR770D0yP2J6H6aiwXSQ2VHrm22YqFPat
3wB9cMtI+XovW1p+eJoPnjvNFtb54j3hSQ2n+sbG37nGAp7r1eeKIBtYO37ld2AtoA5NjuwGRZlY
SbotnR5CSv7FlnqyHJnuoMstzNY2vOBV4lWKupNeu2oJuM1uj9WheuTWpcrI8T0r8x3L0C/V5Otx
jQ1Tc/A1AJsSwWGsgL67OMBHzOGsdyYw7FjCU+VzRAwcXt20YDg+TSu4VS3P7/A/NkE3Qhqcc8Ur
HQGZ43v8RYV3d7tSxZDdsu/26Ud/QeeGlJOQ+l/XVNEKkn93Wz8tDOyFNEUbdlwcURkCtUOTQJb0
KyIPd6iDP+InbPxJzOjJbYBdCfMgOL7PXAQrK7zO51YzYu4JW5Is0lzc7W/8+ala3IX3Me054VML
T0a8NPSKaIwdGzZqZuO4zu1Oo52PZiyVCpgWOsHYrvueAIgfF46pnhL7UDl5swnMEpBSy6xk4Pbw
ZH4oahaLdvuwZk7MvfSuxfvH5ETlSnfpRssYjix4ApKt11R8ZDraT3Q8VnrwM7NIrIzy/requo0M
jIby/MKx5NqkeI9M+OO5dcxcU1mAJ4RZnnyRfjbpFG1PdMFhzJdSureFxCzImZJzKOk5gcr7a+aT
eiuw4/G0P+p1Gijv+PSrzkrWb3iautXil/tWigvhosdJAMq5GJN6Qjj6sCBOmRk3MJcsvO3lyDhd
wwfbcDiGYo+k7rTjw+S+t5h1SjL53V6iODtvWwbVWWdxMDMoOev1NLf3FIUqvwdiqt3WkjWewjW0
B6DDkUxplR09cTe2ycL/lyAQdqPCSt8au6n7uOJfDTMuQ0fy/3RBECISWxXljL7ym5KHJOKowlVg
qQ7FkM52E8WNGj2/XtK9A5CgBm89cKX9RXNyiyVXGJIWo0KJVFWevODAXru97ZluaMg968fkNuhu
alSCxZQKcYIaAVlJgrogbWjjIajZcj0EYLbWo6j1EqVRM9AVPbtfMRYOu49VgoogpHRUfrFhfqSM
wrjUnNPMa94yUDm3pIZpUznyJuOrv070VrCaL3hy5OqUB35+8uzTJbQkVNphMdAMvzL/8d+J8Uc3
resgfQXIkEZOUY02EENblbgccrTaXcHboiLBpF9xyF59Nk4Kv+cIbOmSOJlRNrMTQkZHU9eyYbkW
+AM/uiLru7DZars7pz4zIZ0yJROLWcSKPVwXAffj4mzFUeZ0xkHZDPUmFCH0xIJdGVV7VsN6BHJ+
ICuphe+G3DNXAIDUgTD2AXELsnhJ3Sz4CjeENvDsxBt9wI5YzZTqRoJU9zR+c1KQcVH+ZIdWq4+Q
V5sXp1Qx8Sn+dQP/ILkRa3adBf+qq1gr85mXln9Etl90Sl16gcbVFlxqgc8b+meLbHfiLd2JTlGg
GTVciyZGoum1nMqTlcEXpmsWtNjQXMx5qYf367vQHhII0j2FSIw5l4KKwGZt9JkBnq7hf5VP6XWj
pftWDspGoG3NuSICaNlaR7E3AfjYEj1q3L8/6wyZZH7nMDKNbpGrsCDrJZE1HqHcWRNYsehpIWut
k8peVYqWlZyebfo44EdB09eY/O1Rj5ifnLXjJpL0XIKvEQ8awJBmX+07PXgz04j674I+HcAyMqKd
J1uPp13dXHPmOHD2PveWFQJ30nl2bNdT+QAkn/xXHVSbvqDXXiZkcVUM5cMU1BFQ3W/Lr8uxc9vs
5yTtIzAKqUGWSJXy4FQgR7lEqK3qjt3ZfFLDX+rE809/T6R4nWGxsWWjdooyLHAM8u5ZQd/u7Tcy
Tcu8UnpmncXn0k4k6Q3KF/wyxexv62jxuS7FAilVNsq8myWlO1xqqHnpwvHbGcmGRHVjpOuoeYqp
OdOCbjIr6P0EwEfgWhXPc5v6UpmYF74tDbnRooJO6TsUUrTawCeJ/d+FmuXs1+HHN+y77J0GqtOc
d39rkvyvGn4/hpdRDVUTfTDa2htwHIrwWWqnxkYE7lq6MZMUbrjm1UpH9NCKf9VFzZIg1OENY7aR
lg6Dp3RXw45OmAtQH35Tv/6kYuHNMN0cgbyAFkk7lY0R3mI1yDwq3Zq/NRqRFe4dvF6i8jRhxXKC
Z7o4rfAvba5+fHshpbQsJi9kHzGcTQlncV9B+epgtsJDUckAPl62NBQVzBNMvLM6ez7A2vIl6Ca1
UndiAXoAbGYBBQbAj6J++AilGuTZ0muEsXUTC0lrbsV4MJYkpA3DAUcPJuL9L3k6wiRUblMuWytv
pAI2Ymh9FTepAyOnDZ9JHqpvCiHxdHXDauXE0Ci0MItRexd6u77dXjTAneverrtXJYmeYH3q38uw
GATHcaFD2agFGOVAH5K7bzADtQZECd0QjjwmY+F4dLFLLS++pZmCcZHAXU93CBXgm0zH47AUek41
g/vKhVtALzqkhdSYrTcLzWmWjV70rX555K9fJuwvcrb40S8b2wA8qcMldWR5MKo/gGgz5DrCkmXx
bpQ3UQjreTJ9pq/0/kg1iaal+mC2T9WBc4lvXzUeXIIWneITiS/C5CXeLISziHQr4nJfyQckVFFq
FNl0QCc3NGebHwp9IPc/4T0VFBuycgssYM6idANMPosoTzr7LmAcMwex74bOx8/cLV9T87gM2/+c
e7gh1a6han2QDGCjZs1Pb2aSm30WzfQt9ZBNy2K/y6ltQsyqD5M8gc6WrDoSn8lUkYq/qzmiT0m4
B7MQDnmnEyUh7/3RcXVsKqpWuFNqTsu2ANVkl6wWsIOph9gWuQUOl66dsWbfoUtWjVSYxQL1CuIl
M670ZJmQ/Iq5BQMSaynnKjidexR4KqvW3+Z9AONpKUCXVTm5qNb5dS07fcexMob1Vz1GDNl7JWfN
qN2p0njpeMla978sjJURqJnWahH/y7/dPN9cJUcUHiRkjEdEuv+07HC2Tlfy18Za+VDwzKSzACoc
eHJcskQCOwpS5H3z0CCjku+k7ev0Wri1pwEG4JGwTL1162O2hONMsJi+HvkAnd+H23jL+ZvhSKEI
29p/sp7D0UiESOmO/k3YWnhqGtrhGZEvXYnx1s2C+COWwtTCGrGhwqMwxhqesUyGED2+ZHnkzWVJ
tN+bBcNEf9n7m3LDxC4rJkDuiV93lyinZhD7/aFHbMMIMMwyzO5YgEdl4FCU4VWzrakuuw9h0w33
5GphHqOBP498dDltYUwEa7zKewEz1zEVZx+ur+lOc5CBdO4TreNQUmpAbXD/les20jGJzkavJeFK
WHVrP9Lc9dneGiOBie/m9W5HN8d+4vV/cajAXYdSV9n2jhjhiDd4NHg54fonasdSdPbcxMj4OUSR
Im3TCQwB102fCoF3rFNuHxCqhQf+6n1Nh47g16GoERsY/RiCloWYrpa1W6e+pYSUYDGmiSNnz7KD
LjE6XuaVL2bHdJq0znztRogHbO/mCiqaPiXZnjn6KoyFoEtBYDrDsXURfhxQsxW0jHiWhrUCwMPn
JkeQOprFbubkjqsFoU2DL5J6wl9TqOShoC4xhkQL6HdvwE/3icE/g2cVJxvIrrZvUQf5Sma/F39e
nN4C1OOr4cR5Af/XNnhixV2b30CIrSF/+02SsIL/mC7IHPU+Ro+m2GzVRvzCwZ1E2uYAJdmAlS1D
hlCRBEA1L6YufYMKj6321CyhpRARsEOafCwODuaLV3V6TZrH5OGlOTuJRYum0ZhuzmDeZXo5mFtj
swjWUCAlq+4+t6M265JJqQn57aCibV6n6g7F6J8HUIvem1xViN4HRU6akB9ymq4MWAI7cfgXDLde
rZ83o/PUFhEg/MhcJXFlwhBdMg/jjnAlxgqE/6/FlfXhr1lESPqdZkq1QGSMvn+PuGtpd1N2arxl
47oqktzOB0Oj7MFRM+GMCS+uhOQRPOOYJsGUnN7dJ22TxvYJwUIezg4YCaUIzzNc6vUQwtxZ4TLN
g8TkosocvuKd74s1n5hRjACVPp45FDrNFNME8pkAkFwBqjJyb7RTLmhu7XpElsDtgJ5n75Z8cqPy
UIDz37+ACzeNdTXAFVUXOkP2ejdjAywsPTeO73kisaXPdoZvNaxI78YI6J1glG55W/a8wH+BxMWO
Xt8bcwUZAO2rtnirgAA0jdh7/QH67gAPVr4U2m5arVzBuHEkDtpaSMO0MG8KwNMySGG8P8xtxUcj
FJQOP6f0/oaCJ4l0ck6DAzkiR40v7ACmHJs75g4cj9+32E2l5r511Q+qk1zr7TCJrv4AqfASpFjV
DdUdaLaGW02bACJjZJTaDyauC7C13gUUYt1CcRerwpZ+K8JOj627KtHdHb0ICEkexvO6Q7LA1J5F
RlMVK3yxj7/5+s+nPcTp7v1q7Ih6L308pHy/BXA5Jgl8XfsaNzFEC30ekwBmD88d+INZS/Bg4BX7
m0rmp0leRHa1dLzkj9ceCwt6bGC238/HQlfqKGRlkevqaZ3tKclQXeTmFKeZo6itfH5iYoJcSoz9
XoeyXNo+0FPKTKr/S+mAUoTshdYtkYCWqPlV+MA18u/3MW0JB2oJ+sGqx899emkubb6YmLPOPSSE
s8QbAUgDkjb8LgojDjeQwmyTfAMZ1SP+UiT5spRimr9Ql3Mbkx5X2ErXJHN8vfZ2ey46bgNm1bi2
G25Gt8oXEQMyJn9/mzVzRzoMm3cUqm/PHRIE2AXznZQ43iFH8CCzWLjEqSllXNQWDhzB93+ZBh37
WueBhRW3pV5DipA4bubiQJN2iEoRngfn8FFz19Q1vDcVTZCx0myY0WdpRHhZWPwyBZVmR7KnK9we
Vr/B6NplpeYTDUz2lnFAHkQbpEW9uTczJSeW8+7DYgCEcibolw/jrp+zBsHjLmBk3ruqTkZn4S8C
Qqd4smLp6mXWcxZiSCeWbPccr5Rki9HDAkwRYdcW93f3p0TfLJw7qJl3UeCqx5uJAAF1NdG3fA3t
FbBr0KM8jmP+NOlBTpSkp9oYaMZxZMXyTAYnCWCw6g1zuBPwvUBy7AroeP3QUr2SCIIlsF7A30Ca
7bh7Z3/uK8g0O8I2rlF2yQrgfjw41WtQvh/j8DvmnlT+f7RUIVo7yd0OtP0k91C3YoqPM8hXxprL
oT20YJO/e0Tw5ywYIa6B7na35Zieaj7aC2RdY3RAl1Fji+UWFeHmZ/ig5DgDDbN5nFEv4ywqxfkV
kMSkGxeieh6+EtZRKuYC/Q07RQJTd/aLyHxg04kpk9Ni2Q5tKpOUlCcbsWzrXFyI/y48WZwW46PT
cbBlwfWSF9PsEnm8zqzLKzw3ChM+mPKPCMnigacrkjysM7R4DSDEtGll4d6HijNQhxzlNPgPfcny
wtZSffJhwK6rCoNzfQFIBc8aqdqX3rTuN5o8dH+sfXotnQYHXtxEUaVZEpXe7Qu07/JxFhAjZbZQ
aoURiZTYq0wqjZ3B5HNWhRzDzBIsT3e04y5V9sh+boFqB9nSs+JXrPEPces1N5pOWQI3AhvB1s2E
qz8zbpZeSUvmBeMpiZhHuCGFTZFHZ2AVwQuoG9QwGjcBSds42XcyRkr5OAav0sWZdMV6tZ9R+CPF
y8+iOA1+vMzB+2VIpK2eNy3poJ9fj/O/kG9qE7EMnG712t5TBWaUk9kEI7Oqc7KlltegsJIcYFRK
9qEgipAuXxHlOAwax217Hw+GQaXobPa4S3B5Zjf1FTKKWD7O/tUqKWNavrMJkrDyXAnnksfwpz4H
kWWFr1rDfmWGpgVUfxt0DyXsgraRbWTWxYKn3bIkBSVS2sG6Ml07Vlc73DeLcFY+7AsE6gVgc7rd
TIa6bXzwExVOxKCAJatfRta2eiGYIQlqlTztG/FLGf2i8ScOpwKlsmXSOT8cs/rvQKBFw5UfgB7u
RCNqBul9h5hW9ZpHbAFhkBjYy7O6pOeuiu2tymvp6dA8vZEuGTGmuT48ktDXpOyoBCmQxeaoWgJA
PNTLUTy1RMSx6LrirOYCIGv9ar5pBbOtbjt63jBb27vS0GYo3y4REvnbU7xt3weL7kg23OP6OrD6
15ECLq79sFTdmHADTnhrICecImndYf1iv6WvG5p1SkJsht1Fp+bQGBY9bKHobFNc4bxY7+t8kM92
YhrqiVq2PtmFL7fBm/V1I+5GIoYLGwR3SxmeNgJDiF2exOmbJysQtumjXZ+dQYw+lBk2VYkZiSNv
ijg9ZjF4VjGscPblpYKqATeiNbP6Y6n0f62t9nna8q+L13vp0qMvMt4QgHE+xeV68/z3PI1ZTpHW
c+aSDPO3A2EVDLrURGMUCrJAn8jZvjMJLWLOOD3NJ9eOMkUdER/UFvwORc9BU9TeQcZEdJIfNccy
dx4HhfntfnUHcVQheb5ThbgkJtkatJZFe0wssFIJ25/LLfHont6z09UXd9FpWELas7Ac/T5cslJI
EBcE228EKxiWXf7xMvA5XY61XPB+AGKx8QOiqNrhaOpmnMLS8lHu7HRapsYOTwda6jC4Zc/EhBfb
6roy2UPRU8B9StnaXpF8BHrRV5dGYzcAwECaODzdKSuwspnmfmudVQWkGn1C8/8tdnIZn1EgP09z
QddlMnYxekAxlcoilKBw6CEl0Kxj7qfdSJ+mX1od7W7wDm5nAxbWBUlurt8kmHLMrvT6KPvvp+qf
V2bV0ctewGpcwh7NFhW0RrSZQcnbNWnhQz2SrdbeHK3IIFgHtGj7KKluUFpdXuNxxYNe0BCnSnAt
lxQnK17QhI1eT8xoXnoAvI+l8GTbc4nLs/y6HnoWFRK04KeT16YiONQu5sZB8KbHJ4BeZUsUT/Fa
3tWfF4SojMmxSZWsTUeeGI20yMQldliMngUg8qUd4lLiy8I8QOkf14mecy645aFlKWr/wORNIZi4
NyVLMwSk/gMbkhed8cgMqfLUANEKXaYAi20mUWSgAbVz6u38E5CQ8jx/NZrntvFzKITnfhuicoGM
/Z79ushKv6fA067J2hgyzdeZ0NYyfsmPpfmg+dXE/EeuR4UUTsmkjSAGJ/OueDr90TXifmd1bi0S
CBbAZ0Zsw6SeYFnv50Mx3THVE8ZZEhjqeOQ3TZBNHATYCi1VaSmnrK7QZyHFSTkyIhPr/1vvsu5O
dUBi+JWzWghgCaEtquxgM7qz0aEV5kffxRWk9wYiVPz875DhxgSz/AkZIpXfrZdzmEjUffLaJtfI
rNJzgB52Z9sH1v78F2JQ2UY9bUU+vB+Ig5Mxbsv0gw3+S3DTy9wvu/J49WAvTfCqzYgFSqEsg4yD
qTqDr9V9WdOi4Esra8ibVa7WoayhzNb5hd8kX+0iQ0o6IUPD1hVhCUMToU1CJ1N7g5fxC+FuW/JL
wrWSlK1CbW9caPNOYDKSpuYxe5x0/yEZ0k5cwm94fE+p5Sh47vOGxVsVv3/AM5ahjAoRXN7dKQ2i
9S3JN2FRJUTZv4S+6V+vc+cD7xtMN1Ae5gjiRrFmAsA0WwXBLaTMkyTLHgHPGx7AGkSRsALDWL3r
2Oe4Kvqwl2wYgxmvPylRP71WwTx/4V7v6+qB0AlE5SnooxKV1Qy4yRWgYswafVVBxAm1UrdX1hN3
3I7OLzDGPRHRKyxCTJKTtuULGDWnH6KZ+Mir05E6mC6iSLae/Hfu/AdxhkPvXC8w+nYyRYDcJ8zf
BuH1BjYEGu4c+G3WSBAzOcy+gIBl8hIWXg4x+9nWTXGgOHxwD8LiWxuKhlpDSe8+Zbz6blJXBP0p
eRPnlKrZaCqVA9yrOjKdKmceXM/VDoeagO/6ICSdjyZCwhro3fV7yz9j1zCa47+7gnl002i0nE5j
f9eQ0JrOrqzf+Ik3uaP0WmDg62A7xv116b4C7lKaYC397bcjgfey4W9YmnJwskfzh3iGKTJ18GDg
C+sUqzYUtMag9kkqr0hV7ccegEdVoOUIp071aRNIw4yWVXzPYZa2VgtYVXDs5khavvP8+CCs9U7I
I+XJjz4uZNDCaXpOP0Q4v/aCf4jfmNRDgKLD9PEMxWrz8Z7Kqr7Xf8H9E1h2tT0W61rsyyUN4GL+
lNcBqXK1jMmtQ9T1WyFPu3V6Wl2oQn7aiTyiCxF6xSPFkJCVuPCil5EanFviJV4DiNx8J8qlyxC0
L4o6eBPwlgfpduQWJnc360IHVP9saRV6dPFTf1XAHFAhVwZXoyJHhFi1F5Q5PUpiZliSiOztZdo0
ICZ6wftwQqXiNuL7SLbju+RbKUQFS3H/+kN6wXgP3NzdzEFPRu1Y79EBviQNC1Qh8pfvBzCJBr6L
D72Zhc2l55c5s4JuVfgFvI7M/WvxxdbOF2fDiKHylZK2aEwYDivk+wwnwr7+6KI5OgIwUzdlCqvQ
sdoxX1YHy1L3atckEwNPcXAdAUS+s0pBGFJO+h1dgRwxbvjM1IywP1A+JMbokeEDO7/H/r1bE4bG
v24xhjlfllhD6aoiDcqbinjiCd3SVbtHGYBO7EHoCY1FV04vdh1rA4/B5XjY8YLEoEPltV+kJFeB
iOx7DjPqXHrCgPV2UFzsRR8CYYaiLYJnkcMD6qlym1m0nLD9x65VW/b4XzjmjUaZjvHhjr6VI/58
o6H0k7R7J1t/dZmWkzDW5te4A+CYi+kCHf9xIpG8GwugvQuvQON8nCzZZUYWavZVKX0ZJLFxtYY/
j8qH3rmPm8TN54OXAgIFLGHT8a0wies6UyQ+PsOPK6PKPXVN9Qhgsip6JXYJ2rIMXsIm+OTnY82Z
jjPzfDDnWHBjh1un83u5ENSsUdsGlzYpnBwdJyUSGj8/5k28goJJRttFFAlB7jkKKxhtpkRY/bAt
zE9l1H5LQJqT6f8IBAcs4ONmEsNH/bJwo/aACkm3zmWfaKOTDU//u/BHZsQn3i6QBIG3QnCge/Qx
Wcv5EM0SvUK+LQOYk3lBMK9cIwxNavoHeHy3O8WS08JStg29epGCf1E2M56Lgm0CA8oyq3kp6D3Q
O9cMEpy8uSR5mFZLQWQ6LRtqkdsgBwUFzBVYnlpqGeeZleCbpWfHky1/4K6Pz77PhNbPAJ/eR2cf
rSdT2AoXfG+oKSBH3ENhzXkRpBKjA0TxDxjOL71gvpo40YsuroOsYyywZp9sg3H7Re0IfNK4gn8u
bDf+DfDNE4vtXcWXN6tYAaZlLJ+lkWCRboHsJYxBNYMYLSmAOh5PfOZ84Waosv1NENRZTlckZqPN
sUsV/qn/zkO7ZS3AVDNqbS/brdEjG14IOljv9NVgywHDWYmDSwW3+XQh/3OrqwqgIBL1bxAbXZ9Q
/i5EbYhkvjNfx1tyki/dCM5UVl6iWgPkC7Ht0OCF5Hj7YIT/1zmuWZjjT7JzXsqsZSZleTZkzvI0
xdHhoBlEwyh8vyCyxOKR+wkfBzCc3NO+a55i2ZyMjmPWbzwJiBQoT5O9sBSGQKHKhU2J3xoYnHoT
OxZvBJnNytsj4cxGz6kiq5Jguulh1dpzIjUaQeHJCuTcxyD8oncSmJ1HUySU0FGJDadK31HByHea
k1Tk4tJHjPLRzVJKxnUGfMezqkzg6d5bfTIvvUq6WkZ1p4QK2pwqLcK+R4pnsBjygzhVxUYsO4jV
l00n0bMpmr0YQSzeKMSiiKyyiknIp3MpyKJ4mp2dVCU5+Gofp5hpFKj0Bp9NVA2Oa2QnNaXSFD9y
jE65DyfOie/VlRVViqzNB+05P8AlqI2ikbLGikbjHrweE0WRTeF97BV9bO5BNn9R0G30Rfx56sub
sGt9wX+7L9jg870cniLvWVVL6CXmPbilJNZGm/vZH4AR6nICx2bQw8iJvPGDKVGT7W9sGOANj9zi
YcdQQZB0WYIB5MByGpMg//mOL7F/SIHz+x5k5JfBuaoTCWseDe4iT+tGDLN3IIseE56aTj2sF/Nr
AkrOwVKQHcyvR9vkgxVA4Kww8tOOoA1QPA1ttkp0lKJQRff1nIDFxvXHDPEzHPHQn+yfSoGOC2Wk
Srmw0rWYqsGKzRWR9AEUVTX5CAYYkcHU7NuuzSJQ0OKkZQhP5kGyrNZ2aVc1nIPmNBJisT9F5J3I
F18W/+2fmiigvRZiU9py5idY2hYAs21XP/RnhkljrzXvAvIYpCOxRC8Hb44k623B8hTp6JL/hENR
zRR/3aIIywTH8FDBV0yrW/R8P2j8tY7knhkBLo2otZnt1yQuyNauQq3z9zkC/jkidpkGERAzAdq7
H6fDcTLrMlnIzAL5V1WGkRRHwERmbZyzh2T6YCQVjQlU9csgXJoOpb3dzn4mJ8TgD82Hfh2aJiVl
5NWIGTPwkLmxqqjkAs+t47bFRoX7+3ZycYtj5MPQBrKP8FJiLnNjmkTT2Rk5zbpNgzaje3xkySHX
lePuIdwnArwGylv6OerhF4JfXBUhVwlFndyyPVWcGN0eQCzQwu6E1J87acf9FRVmpO/LHts1sKqy
ma/X5alCd0gEHjAy+pdWYGXDiUanKWUiooGWyLw3KtfhhnTc9yZ1RYJiHAg6OujO0Tmp8nr2g9lk
4dWW/URTN/OoHpSipJ38GVL8TSlDS183iLgk+/NAWwjZ7R/0L55+HUIYe68wa4EOMO2zqIRVHcVP
R3jZXY3f2tsm8m3bPl9mhaoh6Dbx8hZ9by0v9PuMB+a+8Vc0MoMb3157apdWs8WFLnYkKeIaGs/O
v63gilBhQrv+xqVwaaD8/zQvycTcICkwykrrdmzMGVqpTy/oygDTZLB/UJjE8lfJcrb1mGEyHdc4
Y/nz6lTWui9oMp6xBjKAFwI1110Fz00NFr0lF3ep8HWedN74l7lZ6BIP6nUKzcQw+1tehwwWMXy/
d3RLw70SPziAN286NnwZmyYG9NbIpxovgfuQd7WnjB8C3oNnZGxRo/NpQoXi+ERa2YKJ+GQ5P6wF
DeHb/HdWRLpFNwUfSQLf0FgYCP1Ltw4xQNg+VArRAxbLfmHMPhG5oSsj6jrAGjPPBaSNzvqPS6a3
HgArT7Alwo5vciC8oMni8eOW31W4ayzJhGcrwpq+xETX+vXu41AOfr+CD/CntnTMNJwwsU2kuwPx
DpDUlxvq+5RTQws77l8PhWABeIx6Qv+ICezk3K0PvUNBZ3xzMKFx0nfDGYgoXB/Myg3RCmkXuylN
PY2jTpV4nUJ5nOs12sOkCJqZQtO1mVjusNZiS2JSsSHRA3IwR78dt2S3giIMqWWDMHoEFKN26nyJ
gbwIhH6asdHIxEKt0tjfBSE+8RcCyUtje7TbidBv6xu3yrye3e8HQD5KU1Ior1bFBLIabL/+ilkd
jkL4/2eMApaCHbvvhcxtQdk2WvngaUYSEHSv/DLBREY1km/W6BKhLsDL19uIq1hvjY7uUmKSeg5V
7GS/2uk09xSzpTjTHy0wLHhbPl6cOfXWETSXpacwtogJ38zM3vTwHDG5crzoDkj0Ae7W2Hu6vSlS
x31X8VmhRLUp3rWVt/QE8zkp1w9gRpT3utDbeX1WrUWu/iHhT5DULxi7VQrhVpw4ODLXDBCLUi32
4BUAyHMigoUVXrz/9YDCN1AFF5M7z/Nen6CtZnxKpSFEww/bAMJcRX5dKml+9vaVKrCX5kgzHHqZ
uB7lQRpDn5+u0LmgcgkXsJjADYfQwwYyroV5lUedH+mPhoid8RJPr+0nwv/O+QZejfzi2OjL744u
m2BXpzbe8x92IfrKR1/y3a+dJAXLk1/bM9LKqCJclqN2kxx3y1wFmsUnRObVhXzF7WIHN3sJXt1S
VxkOa1K6tQMw1l1v2V9Lpy1yxZX5vvQK+JZSxKWZQlvJ7zRFU4f82032s6CFZe3e2IO5
`protect end_protected
