`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
uoemCA5K63ZDVpLu/lfQcCkRpl375712M24F6/VrodVt88sdBWPPHWuwcMdRLi0LMTY28X2/+1bI
hQS4THO6pJt6GsyAzFP3HMnSoS1cylrQ/I4AFdd3E6dwLyJQsxzoCe2Gajo17m11mwbK4hd9gG6q
219UziTitilWR6oqubR/JBJxRBhtBDczb44yxFeMI2FcdH4Q06xGjAa2Ody+wW99EZ4NUTsVIwRp
HLt71w/Q6FJq8FcgK66+p5u62VhZHgq5m++6vaibMGiZplBPPRDpp7sQiX0J4J3fyLBr+v8aspF2
f/4ksc7C6L/kVT4kQsPAhrvUL0AQZ5AhhwwZ8lq5Iyg5VDqRO8PN5zQ/pbZ2c7h0p2+/pKMFNSRu
az7GLtBU3yG8granvoI+hAqrCtuxsRADtH4rzetgIgR5FivqiGbzTIWwjZZHnW/EzdOpuPWBk0MC
WpVwBAPCRj5kYHdOrdIvJNOO/2BoeWwU7Bb+1B4Mhnua2hXAlw5jkO+ehM0z7lUkKQYTH5CQwZiv
LdmfXNaLxCvYv02dnPYsDRRl72EgQt2cUUDHSeqvR0AKF58I+XVyty3QdRgeiHsc+xrcDX+U85q/
37x4HxKvqE3s8m+8Of/UiUOuqNPllp0gA6mSj+D/fVeMacViJuPkh12b53LuEOOiXFI4WAU9DCBD
gGoXqKZOHM0TGMQDS9It6+Xut4f+peyNV12XGXOf/8nsujqWYANRzDDB9iEGH2PYuYxMwm1k2GiQ
l5Yce2gqTVvfKQG2k0EtZeHgP+lpv7nx+U6HYiIdzTsQ7nO31FSDeeB5AzIsfGUOpednfgBHm1Qm
iEJ9fCDHrhXXZzWX7iXrE0PLktNpidHzq8fztulD+I7fehJ986Fxp9+kOpSf3Fqz1O7I6r9yb5UH
xPORuvMs5KOYhS13WIhCoEyonfO9KkVn10HhgBvpUQwirGgnr2OzwThXxs/4LWzJD+il47WV94hV
S4k6JsRRhSZSCP804ROVd1H6JfYNVgwgyyABVeqUzwj1Aabr8i4VK3Bhp4/pciPgWR1VpXJNJIiL
ZFYionOYF/iHsXjXZtci7ZpXZM1LOLltKgOBCQ1Mw6R58BJqB55MowB0ii3rr8iT84l9CvAsV3S5
HLtSbN7EGGCnCpUav3uRJxUD1S0QmM8kKh8F8uggrdbVPTQXdOrLdrdI9mCHlXGRTBu/f0G/HzMq
66Q1cBqvyKj6zXl2wC0Rofu4mLvjIg+Mkv4sb12JPGU9W4IInJ0OaaXT2xX0hdhKOE976ckaptEs
1UQcgmpNuot2moz85g0YGWZRDQ+2ruKVtAtU5y2gz1Qr6e+c3MYf5bLEbmqE6CLqggfunEXkpqHv
ET1wAI6h5YEfOhSTU8XDddR7Y32duoFHpPXr+iZFyxGqLWTckKQTdPeNVZy82B/3wFroUrAxneVw
vKGm/PDYDK5XI6JmsSuV2xQJeBv7k9/IdWJrPJeGueV2AiImPbXBO6cNIR/64DPSRHeNgivm334R
f7Z2pvhOa5R1HEHrWGFLFI2tIivJMnXymjjSlRTW8qKN2+o7yUOmkreKLiDkp4sCXTSwJcEkwyyE
lEUW3cz0KL4YcInTuhf7LFthvfjdnCW7oEA5MmNhNL1Ch+QYo4GDqXDzg2z3WVEMADSnxuHBXT3r
zPChhxtFWfhou4a3PvLPKlKRxZ/cqnqyhqBHvS+3wK4HkhpJC5uw+CRDy3ldo905ecEZXLmrQpHE
0GhxZwjk+ONAKhW0B1SpzAJvb38X/YBx3uXc8yr/JxI0OyvZooGcZrfeblRDhFlWv/L+W6Y3HGph
Q/vwYYRVkEBjEi6YrbkH96WreeCRMp7J6TYUEyM6Kpaw4L5609iV5mEHjElZjYPQJlh2xvIKy5Vc
A9P8nPDfKkzieN8ze3NRoDQhaxpby8EZNh5KRitKgZgx0xVQj0y9I0xVrVLkmsWZ0fi+OMKmSZPb
VLAAuE9VWw2XkTrhNU6AHFsN1hkxNLGiD8AvukudWsBmSXm0JZMaTAjiaDw6hT0SS2i/p5zYSG/8
rMhq4bO2NJYwARdIorJFAdQv+kkQOqyHfvZbggdzelCSX7S915TTHy+2QL2fV8QT33269mUlM/Em
c0yGmcc+CaqfImTjWsXpOE5Zt9VDwiGNKuoHdOeIBUnV1l4WCamMDSkjw4LqVZkJLcqgW4ovXmfP
5kOjVMmy8KdgUhjSCXLO4OtHlzEC6yz6tkBwvOfoNd3SThRYbyY3KxEMHoHjVVMRJS0yLwVP08Nh
eXRu3dZr2du4CGZg52whHMVwHAAM5rIpkuZHcGauG41u+kixR4tG0VRCifwMpqwkgzj+vQDPePYI
EbWZPwZca3uWuKnTNt76KqGVDCC9n9oBvqHmAJZ53dLq5nYyHt9K8ZoHT4/Ep1lG87Ic+XAPHwcn
1AeOOWm3JL+z2kHYCsJmqtC78SCH2dpabuRtGI4FyaGzSZaNoH0g7x5v8K6uUnLdXTRkpkyjYF/u
4N1drYe6XiKdBTwMZu01B5PP90CXSohow7SGFrbODtuQxcLTD+KdjbWWfNIUzpvfZvVg1I/KvcCJ
AWy+Gp6jmfiLNPFPpQkfEWW8djtJno6k45OGmKR0ihYGg/3ytoqUnYH3Zhv3zS716R55JDvVYE+A
sOUSIta/DSSeltUTOUp02cuKfTdI9rGRoARvm1CH1gjDmsww5AQCRA6u9wANVYVkJAfXj7oe6HpT
tcwWoYsDYTvz07oq6mhhoXjJwmFRYWdYMFRK3DHc08TglzgRbhJL9vOIsxFgXg3tpX120FkqFlTI
bvVfQKC5SAZOyhX6BASxdIjHrd79PfCwZFjag9bK3SJVGzxRKDrFl1p2YY4n6NZ2fVf3qbgP+WYa
eYHmprBb1YhWILW0Othc8iPpW4Vw2ULqey04VBAsfM9bLi+x1QoYHl5FkwxW59cv4qQzJtQjE6Gf
MnBhhWxz18tVet1N5LdQcwjT8zJ1OKzpx4TxgEk4DTFvo7NSPjG5J7cQ72VQQcXNZpCgDxwIu+hT
dPniW+ruciWXqbX+pYyLHjvu4edWYQBquezqsuQNcMEO5No0sGc0M1mB8/VzkO2duwi1i6hJkFQL
AEKJz84B1kQihmJfd6ejtjo1hO6KEtktUa3nYofpeHn6X2kF3kAc5S4YfblHo/gyvufhbxmDZpp/
fAqgcSY9KnqCWUjDi9PtsssipC78xPAJ7oqkJiqTc2R1lyC6605neVom1ZEcMsIhdUVccwpW9ghf
lANMg3jFBz/hBBFlhSl8VBuzDqLcnein5GdSCP3hRoStu5IevmRSGA1z4+gUtBcsmQfxL/uN6g6w
G8vGuDNF2ZJYnHJQRv/O6S8nyae6GtBEvekwBqfgnZ5skmJTqcFtE7HSx5gS4HecO9zoDQqz2b93
DHTePca4d1lrRURJkkIp/hz+q3pgUO2gc3HVBc+m2HZce/g9zhScVuOTt/shX9tr7876yXk4T6CP
PvstiSCZvts0LY9tvBxJgSy1Qj78ybDV3w/NLIjpuOK9OYiT6Ev0xwm78rVWQpjr74nfUw7ckazm
81C/LSJCLfCshpo0J0dw9Gl79VfRbfmCGF4oDdA4wbthpa3ywthguFDYaGLibHrLWo9XFaNc+tzP
hxp9+5k43zZrfBQqLWsOKiQtNRMLH1cwa+4zTlsFikM6pLvgNMREaX8t4BFg6239KP8TDJIXaXRy
p7hyEFlgAPwQMK3FjMgM3tM4/6J9hueGMxLBNHL9fc7JPIagkqEy+ousAT7MRg0g3GB73dzF4Fz9
eYuH7bV98jlEW07hyHuYPCvH+1CA2w2wLY/DVa7GMGoPEv4VtpiySl149onkCPJ4gYkrxCKCOLSh
VkvVwN1hWSXVo/hShH3HLh2OhbyUp75WAaqSW384I34w9CDJlD7SzdxzBZEXelM2jikcWiDeFqRR
Mt+FUlOQk/QFHVUzsE8P8sLrSfOHb+XTPQ2aBoOFG0Nd1Pd90nCx6OP2FnO8Qn4BoLzIyccdOUEd
DfFUJXlGP6dCrgPivTbVac2Wca5m9ZwjlkaIzen2kZCbBrYdjlsFg0Knzt/vLb0NrJpAP4VK0Y1C
bCjzJLh4te/CNEaitGZcqXp9hqgqIoFfT1bXqy8FiHmnH4Vlj1TedunOz7AxMXUP74vz+MX06W7i
6Gb0JRGqNqBbLSqc4YkBBo/AGfhWWuOSkcPVLJFw4MOOiX+YeMyS9ocbIC9CX2WkdqKqY48LOe9G
n73FpwcD6P2SIkXXgMjVZjAo51YNiqHz6e/BBnfX0j3TVFxyS0VOI4+XWyE0e51KBQ1DurpJ9oTQ
4z2Qgp+htbYWpHoxblIClnNA/SQE6UJeFieMj6DT4ux84S41fMHfdJPU/+9qK13YLaWpMXlOgyIW
Mu6gjs224bKRIUb8g/HQbF1qQRcJrtTzyVnVoypLCFoamb4oYZWHFDisA4+Bjmr4+s0R4U1C5Lj+
zYTbcIT//7B5KJVyHlaId9liFxqn2CK9g05B0Dv3kU94aal+kY+fhaxJ/SHE966XwbWkFFvVKd5c
t0+aoZkMksINs4HnckYiJZHbGicIympixHbqh30IT3REY8vlvqnwMhZGrjzrE5wWcVSnilwQKDzD
pqnB28z8LLwj4mTRjTZEWh1RjAqiungbxve8kk/B/KowIt3homEjbjBmOtrvK0ArJ09yCIiNQ1z1
jnHjdHwOAEfcotXGrR+HHwhLlQ2t/Q9cH9BoewxGuWSys6fFy2SiUZtuSvib8tAKrbBCqLhmEqgZ
Z2X/i0UUA86NxLEk7Jquk10w94jIF13+GyekNNObxItz1mC+Iq4cRJsaGtQ0Dn2wfZUCbq/9DdrA
Ak72gV90e28k0B9F0JwniS6sm2Gto7SWV4d0cQ4CeffAJGWqJLk8AM1o6Jkxl7eYIpc49V1daqIw
8JykQjUS58lxJlnBwQUvr5JhIpkxVU3Evu6//M2LOzwrAN3eK29kUqVM97beFcjVtNY4OteEszsw
9pkXse6nC/TiiPl53Aliw+p1sgwAFQy0hJCeLRazSLmbmzYi1IvkInd13SCLdzbP23pw43Qk5Czf
MBhM0NCwHFelpOU9o5/nmRwgn4avCGG1hoBNHcVTK7K4h985lxGvkvjAIdPjq4xjFCECh692mRdV
lVjLoCbgYY8pv/LFt3TZM9jRRF/uTTTQKQ7lFYD1TkO597je2DY67sRAR8mnWC1kk4B3ZyDmnAeW
8vhxPs6JnUG2zy/yzrVR4Ty7Qc/G1CJxJPqlZ4nxWc7Tj6w0j1WprqZIZSh2l95AnENGf0s8sj6D
gv+VL/VCC80pSil4eJXGOXDFsNSawMpMzE83ShoG4WVx1tfJcLsBgAV/cOS3fY9ytrBdlNODD/cq
gY35HFeqHNUactCrJ8z6DzfiO0PT0tkXcbPqvs0CR06uyQQqqv1OU5w8s8b5D+7Nbvnb8ShyBPVg
XSfSfS7YScfA2AHepWC4ihcK+sTGQBoVO6UzCU/pcvUdGeVcaFWRuOChbGrLtPQjMXDQ2ehqX/Pi
5Pk0Fje1FuPiuFeURcxkRhSyV/D3+sf0LCAa87Sn+RDBBD+Ij1c1RM/9aS8WsEM5Ec3n3no3IS0f
bInANH4yUFv2dm5CZLlvlc/gqcYk/Avy/dRAeyOuGDD2vbt5e/gUrmxevn6iKuUFsAQpOVPnRKBB
uES58vccA39Crf+o2oxBwLm/LcQ3ZckEMxgxlxRgO0IghkYpAVAqtsGTGTjBmUU25zhb9/CSu8OC
Yi8QvbMO54tYp4aXhcG9eEsMwo2J9+pi+GlACAl2bCpw0/kwTT9M+pJ7iIqSnkTwEj1lGr0JjhMq
/OLINNdkFH7v+YElGPHrieTmOKCEzkEaTkPTb9piswJjSZI3UclPI7zswSeOUMEw/dwr2XBHR6JG
RVo+ZHTTqDzswTp931mld9zJAzsB0aOxVv7YUFESFFdVpYe/recMalknZ78jpHq7CgZHzpkcgQpE
lA/i4crrx+ti297ZxtsV9b3scRdNCSgif7cz+OtOsjUXffl9TkLQEUG7UPhI2oasutWOGWyHxf/s
GEzVQhFvSACzqDnZmbn28fDnkEL6qTcXzgANViiSw10DV9FuvbyBSzhjYp0fSFVJ5MTopOzAkrX+
6baOUCOFwVtxItNZNhZCYamirbN4lybCatFt0WnDNejpYM2ivPgxP5kKuJahtLk3qUDSMxt7taHt
EQX5jJwrZjZtbI7VuSUz4teLaeYmSOFbC0X3B3t3Egdd8PHYVB7rloEsVCxiRnm4+Rv5rC9UkR0W
16RaLbAutWSpTl/D4v22+Nhrdy4LgTjt2sDzH8kdOvgUk4C54AGA/9oG86Vd1ur9Uih3r7S+NLmQ
SWqm3It2nsd+oJma3w9uIaT5qIol3n+v3nSKDHtm04gaUdsngFEYlzIoP3EIhgf9fOjOrXOy+XPe
VwmdUYmouAfmpdgEs6B7SnBtD0DMSvs3ZXdmgdzKxDYiVkjSE+ZXnhBLPMoLGHeKo3n3Nrh+ck9G
LStTJsUVFuNt2XM1LN0AP+cjUdzHp5Wl66WM8ZxBmNCsOcpZOv/l/JhKsauoYhWOqEikY7Ijsovy
l/hpD4hhA6gzLCsVGGUqX4YvqBEkGZ3BrbeM243dT7B1TxN1cYaraBmajBKfkN63lb/jeQhC2TB4
S0wsHqelQduDGIiub90uzS+iAR34nCRuxLjGsZgpUq2a5QV5H5RsotGskkuqbCPCOOyN7ynaO0HA
Z/EoijejCwWBZ+NU6cE8QMo4bFDlH03c+stmREzVg5fqv/NvS4TaLlyJV6xT50HfUfYsPnTTbc83
J+Ka6y3/AbUFzu20+Aqg2CJv2ZDeVs3QlMVIKSm/M60jvFiAqXGdn+yB22cVhQfdHgiaZQkzN5FZ
jfeBgLjMgrHbMsehj1S1/OJCuEdD7XEkSYQ1s/oZdxFd9VyEXkckR+tHrG4Jpl00HSzfNfKDQczX
nc/oOgDhpyRTHom1lxhTwq7ibFqhDyvAPhrnRsFmBQwEc64ZlNf2KB9bRlkUENgrpIJ8QZQwX81j
LMOYtkNoyX72/YAAMNfHZFNrQxiSYWeZI74Zn8X90uxAQ72kHCxWVZM9IHfXJ9SbYrAtu7yECoGo
lm0mw294bLh5IEsAVCjxfU5CRhfFh0Xx151OmiIbNXexlAbuZXeAwUFsjnD9Jwqey/PY37yVxMbe
L1DFRzPNTmDz43zv2ciG5ebASyHlka0GL5g3+t7mTxbHfeVTPsCoWzJyn1dLXlW9poGAeB8QugqJ
A/GIMWyji9yFVwcuL92+Hyw/mNAPvBtuy32z9aSLG5RlCQNzB2tG+7UVapgML7+PKPED3plPVxqh
gX3ZVJ9epETuxUsg9REjJGe8/gGdwhdFLmzXkLjGbwEqScRx//iipyroyv4xWN0UMEugfnmSGrz3
QGDj/JVIdncNqolfkcip05Nq7VqsbxfkAKvQuNjll7NJZk3OsxZtg4ktv+jtNFwiCxwVm1c9BWez
ly25Q4pLn+3XHNoCUzxZnN/U+5JtCI7XgzF4sLsAcTbwfJ2zYElet5XaOdo6W8PHiFa89aeVrnZE
Mlvk1ALix2NaVYCoshxB3CvZnoNPzniuQUlUA1vH//x5ywx5GvP9n1aX1gBnaYhin5h6Iactb8qF
pn+vd8bGn404tEJz3ZxxsTXvGEQRg8/fwLZtNUbT938td351jtfWBwq6qOOpN3QiTsO2mbvO9QUh
IwXaZaVD4XsnYJPxMN+3kOLf/7oZjQoKzhhEFX4smSUZlQfDCDRkNdZaBIonuuf6Bh5tpL50dB3/
hRumoeTDU50rbbI1eXJGyv/6couViRv0pkBwLts/u1AYOlaVOahVaqsObFU+txk/zUjPZLCoWYOx
i++vTA/+s/S6oPaTCHhrLndHbMhEyPQg60yX/JsVHjVbry7cRSph28zm5wEQHrk4g7/V9SkoqpDw
DwMWbppuP4ZvnWXhSl2rIgGcdT3Yjw+A06rYAEva5MlwURbVonvWUW6qH7zCB3a7NOp2vCDpN1TN
xXdWhOYUT5P+KF3Cs0eshcIyifKONbic5FmL1PIApaEe7JYFRlCdW87chR3ku+vlfJGYUsFeRlvw
+uVCT3mO/npyv9iuZv5gnAcaS01WvOO/bl7CzhceXi3J1NaQUNQKxjEUhTlrY7fIVrlPFyH1czJd
w3Q6TbRXxHpizWW0o0YhZ0NIGwlo1pvFEy/ESsv9iq9vdzSaUjgW9p1vKT3Z9V12xHEI191eigLc
b3GdwjUT3NaPmABPr0c6GiGSiUbe1hFl1134TStRROofDm8FMRgyxevNjvvPWNtDrGpCnpGIgVnN
2OXXkHOay+zZa5PBn4Sk1xvPO/syx+XRQ6+v40BWnRZCLMvfznvbvyS3viCADWcIJjSQTn0RZUhO
95y+TiR6GGcPf66Xcti4ASLxVPqz/ouOdzuKS8UFWwIwoD4Lz1IoRpeZUu4/R2U+FAzcsguH+o3H
DI1C0myFHkSWVW+dQU0ouZTs0ju1CdpytUCoRBHK2sr6XiGEnyrwfD1dhQK/XpnqrLErf5TRRDVr
ovqxMnPAd4cWcQZUoeAb7NWmpDXkmOTTHYMgjQvE/CWf4ZySzQwTLNtnj2ukG+bjJ48uQpmcVTdP
gsJPCILFGOgIooceQcb8Erx+wh7wuDQNOrxh4yKipxLw+0zp+HIHjtGnl2yeK0ChvdJgCHpSaDzu
vkLyagEngq3rmlZ8ESqFMY0534qQlGq0frSOmK8WjB0a73+qjah/FhiW008gqxXlTaQUOx+JbC60
3S126Ys36zdso/qrShSXPEj+LSEA2UfMHXSR+NVl2UTZzYDuV7DB5AiqiB4rXfLUk38p4nw3LMX/
VK0ava2ja1fUXeFWW7Vx3vNx+Cxj889hoe71Td1rxLkGH5k1wPjU6RhmwUB9ABuNnM8bok+x5Y+W
3IzdLE4Wk7zLeLFjKGqvbcXzmlXCnRgdJM7PFmT2No8HUQ/DRPeHlUEQBIjW065ryMppieZ5Ttpf
xe2mXToWawNfUJ4aL/l9B1yKU0i6VHNROCLwUyUQWH+yVJyxDHYOXGJXHOxUlPih0HU7Nlhn35pb
o7NM6NQlvzVI9sXHfGTH05MUm9ratFld3VqAqwrMPZNooxS3icW/9q0epZwqrJ56yuDdpraTB+Zc
DsVNR2TAqYmpoeMGOIvqTOI0/IHymgFEbU2qYaDNZwrJsJCpBMYY4XyLJQ+aGs70oYzraYuFbpEQ
frn0FKYlK242Hzwe/LTyl8wkjwpKAJcxzU9gMP72TkEBX0w9auFw4eUkDrc2gYoUIwe8U/MLkv9c
5wdJPlAnEm1RsBhhI/NFr9G8PssDXov7QSjG5+74TN8TWpYYlesWVLYOQPKA9AuYwL9l5ivUW5j/
AafFGpCygRAZqMAaNj0s+zfDjUyAsP7wgjzOi9DMaFn4Y3MU+qMuurjJQEUJced7C3lb3iifzOzv
NLmSvTB2UExwss6qz2nNkLXPVlSmmkIdntlGKe35u+naOW4h87gtmWL8thpcOAMPvaw5/3kA8Kyd
6I7+j4BtRrUPQetofmUla6/l61RwmLO9DoAZjO6J6Txl1+ZJx7H2ZXt4w9LZ89Tt6NO8RIPGXPGs
kHyeT51cXtljobikzDcxCJ8nMp3IlhGUoQqLLw8jdSIiVjAHBKiSXzNABjpLsGK2H52IDpksniMB
dEx7Hvgj2LNlP+k9hmPOW7UJICj5aX5086BmG2o+EzLtHY64joIt+dvIPAd1cwH/L25+iZ4yeL6h
HUHuUbb5icE7wqstZffsRc1VEHEpsfwmLS9u7c78OVYpY7LBEa4+cRespeeKgyXNDfXHvoSPugeZ
+hc83lp8jVNa/rozdgAToA4kj3fjHj/jU4j0fQz0aKhQfbEOymCqE2DdC0z5+QYaBapz1vsdpcVM
Q8ePvzwI/KuDg17uh4iQ9f2J+T6xJhsvhMaOWKGB3u4/HJEaRgluo8lkCO6YlxkbBWQxiass+WZy
bJCpHiUNwCAFeTOZTbDAKmGh7CKUccQOGbfmQNNX+6HXxXQEw2/LCNjs3Ucpu1ZUkIBzFnLBn1fg
DjFezuGnlpxMj3pBG3zas4Vzw7nADht7I0rHMJEysF0bFkHcBuW6dGacdKgTwtLIFn/9J4KQ93Vn
aF5LYbsOCfJzHQkjDBm6hZmm5QLqpnq1ZYmgG1oNtlWMl2urSaokr1PdEANgLX3IKIFzbxtxGuWc
ojoUwFGEC0HtyDuzqT1oX0Y8JvYQWAU5zz3/3KOLjEipMigl0oBFYkJuAhN/CfnALz0qTxOStu4b
1X9hCsZly4Sdinpbz/mxQOwAMQ/w3jj1YwB9lD/21CwC7IUqGdmZSO/IJ44yQkO3axvu5BylefT7
xVmuNKYXBpXzghpRvy7jaed8f4vv7yKGoiy12Y5dSzeXuYmo/NHIZbaSpbFMKCT+1KmfHWKF24Az
6paRC7RcUIe5sTFqC7RvOLsuaoOzUy3PmjlneYAm+t5Fj1Fqd7vhORY/Mh+ZHlVqK5fhQQVx3Mo/
jdKtn13WIrMJA7BeEa6hWCdHHVebutU8k8zEhmQlwcN31K3eqxJzyy+ZD4gPT4ub9GuHjZVK5X/2
4kcVDlTRU1Bc2b1qT0XRfz5FNvIlJEOqoJJa+elwNFIr1HaZ/BePtk2fNcdmNbQ5IVJh5ttbpfez
i0rs6Cp2wimNiuA/kE7FYy6AxBeeQrM+GARPBbjnrP7ce9zwWAU+DfQSi9NQ4O538UmVzRP3EKCJ
WSIrQ/Gtdpe+mWYtD0jylRhz9w0HbGek2OoQckuVNbu+N0xNZR/0rWvGgLifW5Pg5dK81w/wCX+j
6QgP5DxL+0kwjDFOzTtmND8EZ6TPxM924X8eBuy4CA/wdzsFlNTMd+xPYKqoMt7YaZRAmpCfeV/I
QgSD5lwMOckwJU5qay5m7MAvDVreYUiRSIn0GY72msJqlXTBX6KGgHUmUMW1GiQ3hr568QWPJVxh
RW6i394Gb98lK2uSuPu0Pnv+U1BXGMgfSyhtMjmLM8NLFQgvbHvT7L+J/UmhLrBX0pzNXahKnWFo
NyZcFOVyk5tZiMAyu5r5VSFZK2FsR+p/IxsSv+oNDTXtgvgnTQlJYk2KYTbGdu9ohNxq7kSvNt7a
rOGGaiX2I2zvY69nBgl0/GaE5fNWrL1uw27HZbD9a7ngkHTKX8Ke+4gWU02RjVlm9W5sbcm4QY5T
ixtS6zBDgMshaRiD4ATcY9s39RRmWl8bs7zWUlMSOiGNL5e4VRDjAAdmpM58UMld6XxPltMCxjd7
WkCDLeO9DQX06rS7NKXxmAnGHKH2DMikifK4eesUJs3ofjuBfu63qSJ5Jl2z05C07mD/Qe8ci+xL
RH6aOlrxUqLZ+fYuzFGJb1Gj+bceKDVhS9Vcr3XkWbRdEaTq6PrmHgQmX9dSzvgQU98fNiOBb7DP
LE3+LouqtQ1ONcgGwWwEqCszACq6OUbflpcSnXjgeDQhyKZsVrbbV26VUJOlsoD3Tm4CFSHFZAul
qPczOcJnxu6ROViDbAddzh8mp34JTBE1NhjylSHV1QJy40pKl2WOiNYRjgSU42hG0oia1CclwSsL
ZursITLgsuGiVURzZJF7/blUF7D4dDITrMxiuT+PZi3/hhGz7mZM2Xi0RFyijNEGlSjZ76XBq5uO
Pzi1hONinDN/FIisuOYUXtiFUZZ/HQXZXLeTS7Glkq5UpNSEyv+4TJZGXkxHY2gA0yXCRGIHP1lL
4R0x+kD0JZbC9xpFVX+lvRZ8JzIJpazbLKtcbEv2wHeAD/Zuvakrmx/vBy+BUv+aX4yMSYELIasD
vPnUwgebZhT5Kdsx9pp01X2DfszvLiwuU8b/4imQezBWLWN8fcBMAEPuaHVEtzDy7G/Al5EvwSd4
MMUvQdJY51027uzFf91Rpug2ejNQuyR6SzV4VUWoHI2U53eV1k4LsgYIAx8Xq2RPZUQeajY3cI8v
kBYbtX0LFPXC9iZqsYhin09VY/iMwGgJWZfyzx3ZqJ+g/mduWat0x6sTZg6rGBUvP+8ZB4pymSGs
6OaioEzBLUvbWsQc/Y+uoOS4ImXLXOsjpxk95fRDvpGqHLEzRJZAvfh6sRH3nBJtcpJpO7N3U2Jd
BdUXQy3FjEe/0Ue03YWjGnvgdj9TzuFO2MP3sdjSQcWxd9fTFkO9I/FbiT9e101WtPmQrIa5qDy9
nGonkPhd6kG0imVfsToANLMC90GbqpDOCph6KCc2iSPINVz7xEhoD+W/191Xab5bZCZVsok1PIM6
2inxQKjHq8b1MZzgIbLpQ275nspF74z3JIuewocbbGkQ9Xm25+gLDckJoBcZ/k/WHlI0g1NxX1hk
I44VgeONX8LjP5/p3R0nyLcYahFSIJSEdGUL/7FYmkIQhUlEzY/I9MZNWMH9MGoLNzDmvgNydtYT
0xgwUpMU5ncQYihUVia/FcbbVaJAzrg0cADahISHi3U//H6diuztRsy9cCs24D7q36G+tq2ge/jB
X45rw1odoLyAc/GzreWMGDZKVWetqmspStYzyOG15LinEL+sV5XyA7natYwQQ8zMF8oRca6TSlDN
NGSZJ0qa6CXY+Y7NPDxPMT21KVfkwDbY/do/dIkGiaGarl2Gj7jNJM2g1ic2UGqItVrD5EIsFxVZ
NJ91+LOCoapyTV+O59mBT61yzaocRWuUkl5q0Ci6mxvg+MxTXqRsFZJm+RXCZUmo2TbtcgDPz+9y
9mFqkOlTG9+O1k6lkD6qxYYEIMlxfPA2sQXIo4lWhHUqqWPZuV+B9UIp951VgQTrpX2snPfQdWZx
xa6Ku4WMbiZqWmgUapssroBoWaXzf4BaqNqosRQUoBDZqOhjGA6cWbb7tG3WnJbYfIYeJGYvsHkX
PHfFv9UDh5dzqjuiEbeySAlLq4C57bCxSiN3k+F2mxcKHw63X/YBinUzwlwvIKCohm+PKPQfJKhL
3WYYUVubMwlrZQZD/pA/1oYTfBOGM5sRph6IXArwvotcGx7nAy5VIoWmJ/iBBcEwdSO/hUSL+5O6
Et/y8R9IoPLTXl+Snp6NElRRwyJhYHyaLZwU+emuXeOQV0vmgYzjqgKrfUNQ+jbIRFcKMhiGPiGw
m2I3pVODRnECj4KTALCYWRFPmgh47tECk0d7JtvGK1t7Bv7MuBSEOHVcjdgF/JhrwtP8xwMqDVCi
dh632gSrTtMgwOxmnhba3x7dBPnU0u5ihiaDFyI8Q5w7QjyRsTYKjzW6l0HnyFKrDR47t3Nsj+t3
R6HbMCztA8gHkRw77c3Ugp2mNuU+aQqPjmy1A7fjPPK/JDFDZw791j+T0kQorJtEDd+ohn5z5FJx
fRJhp6qBqZc3aS4fMgSKlMKeBw46X3fsxguMl0dP7/vpFpZTAfleFwwUqzUmuQ/c21E66+bDOK3e
TyXs4Db7sgit8KclMvuWBG1b3po91HNJ8dT11uSuIlIFl0O5itS0fwIGRg7MZAmMZbdKdsMGZ+r9
Ig399FcVocQKaQQqB3OzkvE+NfzX7SPPvLHw28p37hhlEkZLP/FB2aTfStJE+GrKC7aIAk8DAcQR
zWOkYIXygsbVhgODFlxWR/h7NDu+c0h/j1YQKCAG1lcqIlMGniyZuljdn4iv61Ht8/phEjajXfT6
FYZQpWWxiNeNMmgAH9xyaqdkHXOyLLSIRM7tdBw7TNh4E0WbH9j2v0ru5bbnVdgZdmunTb8oVLJc
abC1ag1kH4PxLYLP8g5GASQyXCQ+wUvrT8rLdSstRf6P7+eY456ixgofgexk5tOkbzkZRz0hVUku
y+tpFOIxplP256JzWlj4NkYy+a5Y51DEy43w+vfaiABdsvwJ3Q0aXh4c3T82bn74In7Li1ssB+2V
IQKoFEbST38cVzwAnOFelvN28EFeb3jK/jpCvu650AfLD3Yv7B13fsDyxEY/i9hh7jdArAaHqH8v
aiDJIY17wWxgvnOmW4S/gCtuFqf0znLAZ7qlCHaIddtDr9hWG/3X8ucMFazbewG0E/DiKbztsEER
23rZ1j7D0RQbGm9VTCx37xJ0CgyAIa407/LvdPfJi/aKK3j6oPrMTdKAaSgHVbxWgF1QvnRhYX5v
EaFiYBwSoROyujVs+HwXsVCh4bwl8r1ZnvINbyPFpL/YsVbSbM+x5sR8kZscIv5KcojOqx5JamH/
MfVLexaPDem8eslXzdXxZDv3qQFc+TfZPvNz5cklvkCUQILtubPSNInq7cU2YOmBQQ017WHEnHuc
keJnDz22DpTBPhNnx5Iy5rS/m6nmCJkXTNygvfHpr61Umf3NkCLEFQddBB9kNGq85wV4sd602OcW
0XnrQ3McAmWviVpw0hpAVht8Of6mILVezFrIUdnRxoMCqMj8VNSHpwTzZsBHGfEUkdFJJ5lOiekV
ERb46+JcL9W4LBqbxavOJbJky2/BlbaPQatDXdSpBjQBShhMLW5H4mlj9yyRbxCVGVl1IJ3waIti
JnB3/MN/UjtY6Znw/umD2US86Lr7darDqKAcdmdhMhSDA5FhOiTk4UXYRDK+BUv7FUYZYfjJyCUL
aBKNO1gUY4nzuvq8FLg5sJGvAbNXqh2v8ySEMCv+tyHVw9umdysO6cZYsL3Rjcy3e606kUA8wyKh
p/JMRvXgrBTi8eqGCsKi8EJ3jqZOMXXqojAiEicg0Ow33i+X+cUoz9b3Uu+OsfQIo8jm1DcRD1W1
tn+UAhC3ydfq1cw3UFfS6UOGhlpQmmywf7vZHthTkElZ9d5416mkgkcbjR5Oa/ufXICTTfpD0jjw
MdEIG58uOskL0pGsFB6xbpgv9cD5PJJedaPAxgkvuYjolSYbkKXTfOYjTcMCLC//63qp7hiUCX7u
ByJSiKvjAj8w/+SiqMwLHLXzLk/GCCX5dr5nVgjmxP7qUtL2plDYJOHDPSGhHGal5O+gjs4ccXbf
h8IRMl5WYKximM03H8Hr2klptgETLg+t73dU76xb1G2i6pyuGL0eVayuUnz6+y5NcwoZkAOr3e78
/Oe5H6OfeSmUgp5t1bKCv0VxjYtdyKs4K5j7h2Uc9X+4+Lqunxw5YLRygpnC4GrmKfMuf04knwYX
Rkd3mL2rHY9LjHJPVe9+Maa27sCgbYzZLPCuI4e74bhPJ0yh6uT40V/59jGKlRW5PR2Co3+Gs031
JSaeHWnl+efXixVOkniK+zT5wA4vGV/SbGTwkkaAZJ+NhxyJPda/cdwpYcxR4I50+NL3MHpK9J1u
hpXO0l/1C1RzStN6o5ScrfaBI1iD2k3aM2QHIV9CvYFxPo8t26hxT49eXQajcq9b9Z38Afu9SgOR
uYQJd+FYaPgBjvsU2cNgQ0wB5x9QuKSypcEA8pJEEqFmVOhYTxK4fs9R035kP9pmXHoMOMP81vn5
iKBgRDeYoI4ppNTQ1D0QAqymNxu4krkKRJlzx7qMBAgHJOr14v0x9cAQQoIbtRYUui43DTwZ+ckY
vow6HRaljw6yLZZ4MRsaasnkeD+Yr6pOaxwyN0uio/s810n9Z6SWkQEssxk+UZyzqsQDyX7/CBec
e2bfMRwIxnb2qhwY298BrTYcVWy+9UhiAcX3GYT827YvVqYtjPi3Qjwg8tm2FAvnYeK2MS9aU7gu
tA5Ciu8Wi7PWS2D7QEITnU/tEUQwpfveLK//E3zgOTtWwEDqA7nex0RoA7i1Xh/nFO5CYbK8fIt3
/3U92K12egw9qeJK+iObkQii63zLihbme3O3sE6hD7aNU6KeghWNnGi29HJvyuehbudrhFqORt0G
FA1k3Rw6pjzWAmWqPv7K6Sp0AsnJiTMZUlTYbLl0T0I0+Yhk215YJx956gm6Wcp7mYqB5vGXgvMD
zdp2C6cPAQQSkUnMrV/Eg0tcgp3x+UnFt2mHyFKtjdo4Sq/xxilnO4wrpPSV+wZlUqa2p7qyaM/I
/GhJbli9vI8w8OGh1ytjMLYLEIhT12//apRNvNQR05AzW4GOEBZH0sYEcEWaPpxa570rrwnHAJrU
zNvCDOGF9Ow25RlMcA+8CBKAawy5Ad3UUDyg0YgdV25QINe38zZF0AL3fwLwD3nVj+0LARvkt+zX
fjw8NqKP3lR3XRjMLFulAsXdCnG5h3Pu2Pwk97aXFaxyxK0dR7pwP5Wx8cgxgNdCaO6O7PXcSml/
zHi5Ulaw1UnbZ35TAicwafUhPz0UqIZNx0rGYvinB7/hx2eOSGRsnPJeVz6r4Ug/FTs1UGpv43Pm
HqhyaFG9i6NjjPq3fouWbsR2+ipitOtziowGF8Hk20CCta5V78Gvzr2u1Iy7K42SlmzOC5QO06uK
YQX5RR8MfsQdKiXZX27csH2iA4AnizOFTWTt+UNbiF2OrprzEEA1gdFkXBEE+JAqgaC01VGClwAL
FctRxyehXk2eZYCjFGSMnMB7rc/hJXzIzbgTh68vCec8BDqflqXt+624qNZdYBG4CgTmkpL2oS6M
VwVNzhZHee/iPP+TggWxYnZJh3U9vSGKJLVOEtU7B2fNRKi9GIdR15apVSZtuFYDORdo5IQ+c5yY
FXVyDt8bz5Ycs/tleN5sjkhCRj/l0Aj5cG76ZzL5NuuZr2J6kSzbfiAGciQ0+CCIqFlkpG5QcNqz
AtTBhcS0Mk7aV225/P+zlIt2ERX1SpU3ow7ybZaIrLPQ9OQzp29y441hwP4BcEr/UKJVNsQBChfK
qskPgt8yep2DwVhLecC0T5JT5Ujy6MZPy6qI5iJlM3r8vUeB0kTFeKbIZN/dL3atmCY3d6ZS/+/K
G1Yrp9MLlWTkYWRX/EvLiI545A9K+rdovsYc/bGQc/kmcr8NqoPJ4aQx2biTH9Sdege7sej5QPpj
RNqzKZ8bm8VXVRH8LWLyCQKVx+hJm938P8K8jaOApj506JondnPElB/FYsQ0R6Rk0udvc5em3ESx
YhuqPFtYhKGVWWFuWl92teFOkTqCBwNAHEsiRDx9uVyGnmLwDCp1UHvo7SXd0EKVAFxtYte+r0qH
eYpYzNYYvhgLe6wRj16TSS7bsZKI5T3OS6jY+sZAL275w75VEsANX2UltJASsybf9kzGRY6V+Pwp
jzQ0yokBtUZCL2eYJI+EEN7dwi3KRYEUBUyn7FMw6bccesPLLR0bgagSvvfSYzbj9rP8Frjy2xDy
2mFjqpRw4ww7zHbe/AINaSLC5UqrwSP7zcRqM4p1TdzQMOhP/7KZv/P9d1YmFNanpcXA2cr4dkSh
uponF5/5w5LuuL+NwSlgkymXRmXm923D1/FhfA7ieoPz8yp5+eeVnXEH6oAiUR0kBGG3dQEJRJHp
7Y+FcT7hRqgQAL2gm6nJD8O3ycLFHvtI7q8n7nbQrn8kjhvjCc67LWxahRg0klBC/W+0RteYDt6J
ij40dfVbQvY00IIqMY8+fhxdir15g1Xk9jHbuk/VvYiPxyc1GmcoZ1ULNQTjPaRbrsuSzSvLQA9y
Qz21OB8IPvijQXk4SuqoYoZLmXrOEcnYyUwMnArhQpiCjVcJVF8s9iYNjvqmFdMvBtK+l+ahbVLS
Tiypwf0QoEW03vdIwnO9IndHQKzM/Dg6s3Frl00TzdjMjM5fBVAB1kP00qPHSalMYip8djVsvuFP
knlzkXxhbFicsqkKfLTU/GJs6HpgegVG0LT+5pi9Yx0TXuNccrMRVUYs/6fFo/CyM9gGuJJDWXOd
eXZedRuffgRmQ9mvzUAEQFdnbJnvqCrr1oUSYCS0xsur+fiaOIEX1RI7pJcOAWLg2ImNWDODamFR
HC1PtzCe1rF5B1noVK335gTh9AEF9G8M53xDHfml1Qr/NuCFOHbjYOyGvX8FfSnkpkUbKkmwjZEf
XNENyAO2BoMlukjFYQMefPoPcoIL5iwmsGy79JkzaBRVO4iPA9hAGDGCMkkC8drHIjeJj11f/u76
g0JLHCKasZFP6/jXNqa/ksiAn9++Rr0er8s013hthzmzzu8C/4GRgZ0eOjUX5n9pc4z9u5sHpLsF
hqe4DHlf5BfjqeOy/9kWU0z51EMvuoL+YoY9teq1zhm4fBbOUO6PBTGof2eP/ttGTkc7XMnyKaJG
NCuQCNHe1fxtRaabr+xG1tXRkmuLMTwn9UeP2v6eXCYVFetKOrG+olWXBnod+XgBn8K8hh7CU4fF
pteMcvUpA+vUsJ01bbhPG8kl7gjFQHTiqxMy+JpCtaiuVpyHf1aM6ULXKj0Zgxv7W1atIz11eW6O
r/hpJL8DVY4UAdhVqiC9YMjcdqVcb86ji8Txdjdp7xUMCon/S4csO2oMftjTSZr7Nm9yRn68zrHH
GlSKkmKYOXy7gqHru9BbTL3o+Q7ysV3hCVHZffEXJkqZcBeMhbUHy3fLPtS7PHWSXCELqVmDP2qE
y7gkB0NV011D9b48TPKBVHc3uEA8m/smii7gA9ruBkmweXleEXjMyGXSOwYL5FzPALRLqd8ttiAY
SXAvent+uh6SfxGRExraskbClyGR6P4YdYsRnSPrqlOwWgokiyPPOMlOReyjLw36Dgcjrw+KVFew
E3esplxdpuMjYimTbLAFXJxjk7VXLRsoZwTf8ynEnaIxouSXkilPOzs6BZ53LxM+3iSwf8MFeKMt
PCec2AwhMZFwNVBppl1iF4fov1igwCTKx1dqSKoMPg8GdVFSu812HNo+N4rfpMArhp/2bPbrwoCx
S4kolC9psW71wSR8Yyt27QgvHstNHo655mYYDf9TgKoXpV3VDmsCBzOEfqV6z9Qt2OhB+Bhc1RR5
kHP5UhRcPBWWYDjculHmUZ+bcaf+S51JnvG/GztXQ3vkUchEPcYpnsdqKPa4QNFK2WyBzfvDt/O2
WdLIjagYAJJeSj46+40wq8bT9qSPZOdmUmPyEuK+JvNasUKCUE9rRSrDZEpro3PTHqE+r7VmixEE
75WKrS08kQLmyE9Ic3HnmxSIZ7txEB0rLhaeabrvgd7ROtgC3rarGI0Q9syBqCptQcUKPnh41uUY
Ac2IlVWDmX8Tz9OFl9tpXQTaeQxLYlHC1kCg2Yn33MtiJfnwCLZpQNgm6C3pL65bK5kNGxNfenvw
MXxW1bMY3W0tgpf7Mu2oviYtJ6gIU4uutkfSDUf4iGnHSceCtuKr8qBDlhKlEdrhXs92PuOZEhCn
NvE+ok7XB1PKxLUqAWONu1Y27y8fwxnDSw0IkzA24PuRGt9Cdzhbn9nPwfiORks6/PNHjLzfwx6r
xrD6du63io8TMBhbgsTbR0YR67+GFvwxnv7ozmQIbH1iFmj1d+T25C+2XKi3W+QNbVxQtK1bUyav
dX79sirFwdk+6NKOL0RhwEhKMcgbl/CSDzzoF+AOJsEly4eptHCLLxiU3b1jxmqpw6/NvLtmZ+0b
lGweFhDkm8G3NUq+XbTVdUevRWRayxWufzQdtzQ081hTMO+EPfdiYvRsBMtfKyWetvEq3Yb7pQrK
ux63/gyxJI06pm/QW+wRMNox0Fa28kr6zYorre26aOutHTXvUP2Y+OBHvS9mUZynCpGXvCb0Q3kn
pMj61Kj/JHuMlEuUmhs7cvSoj2j0xpDqMheNGipeOH7mzx3pSMbXcBEq4lQlV8XlxeBZuGfcF85j
FveOCBir12iLvUVh1vIVfUpkuxHdXsmeImLe3NL8ywiSi6TtQMfk2sW3u21dQaPyW2CPRMmXyKto
9sOwe/vV1HRLMAfsvLfS1yBuiJM6W5TpQTkJxHaj/qrpbj6VY25fMpa9zyYjxGlVE3Dn72bfXxPY
W5+daocf0u1UfEalIDdbkN9GoAOMjIs6mMYGfkgpOK9Ni9NLWhkjBOIIz3wWcQr2OK9c4EvAX9kv
9sdv5xN6ywbnlq3uhByDSZgMKQH1BUevJidQBGxFXUFHVL6jTi2q9glKZNyeqa6BouWni2Mu85nB
BWKCmE6BwgLlN29u3ICTG/Z8CjIqK3UA8gUTW1yfycJ6CoRHV4mPP/dF5MUeoAT2CH/lcB9GuooV
CyuxygRIq2CbGFMH+GM5IZ2pA4j54AnQrtz0roCtYbbiJ72t/35RlycNV+U3QD2qUmGpzJooDGm7
P7G4zmPQ36a6AauGGc6GI3oXXvLTv7KH+8bfXXOmxvUvmFDWRs6am8n2OIdTPCcZrZ+EkeeSCJ0M
2EIPLOH26ihDbegYl9JlCxJN6zZxSTZgfcqs82yRzK7MDXpIFEmVXpSrpoTawpA5T7TT9ih7Se+1
ATPC6+MVuLbOvG77Gm+OC4n53+J3MEfLq3UtdRJeQhmpu8duzIqSOrT8v+tlrnsPn6Lwa93/YONw
S8g0nOXeeguK/uhYgOGaC2dksmJ33X8JwJeBfwlllYBrozBUyYIXDC5CnGsdxjrBlqHabFiBp5Db
5NphfONp8NNji/6jCRBHW1hqQ33U5WCriimTMRg30cW1YfyAtZkhJTNoYDI+C8LzKEZEpO83K5GG
TLuH+ybEwywb3Y+pcH4MZH5likQ1E193nuQ/wenNL94UGO9VboY6YeRMtXByiis5TeMOJa9Yo++B
d9W61NTBbKm4OujiqQnPx09jLn/PnEZqkpKdmv/JPyLAYPHwHkzw/9mHXeMGKrnRkWgbTa2Sx919
P77UPeV2WHQggdwWZD/1O7hFcG+ZQw6aK2NWXs+UJtH1emtrh9IZHU0Yj97CjdrmbUWkX0YPWfWA
wtF4x/hCmOzQaDwwit2auPSuUePalSVIQ91kWloCh7bnC2SlFqPIU6Vnqil9qRgI7Di2KTRXMEDQ
UoJThp8QOl7bKFJeviSXhx5cmrzHbHZ+MTck7S8+1EhTsg5T9WFGqi3haJ4r20cDVy2SvLXaKMMy
uQetWIizu3x8Xabj+8rNgrjnWfW0vr/0WaOyiQSiO0O0rEj8olU0dr9PW32Zsio5Fw8agGcdlZej
R0TAE7WervPlZPJzpWX4CJEJDzwED1uf4FduENr6Xn0nbLtZ2hOxnYWieRdzxRRcr6dnH3536F3b
dEvfilyypx+2Hk4n/qrAbKtWLLzYHk7kYK4VaDo47QINumWqfbDZxUVPigFjBkU2MYnDv5DnRRb0
6iRi5tsWZEbqfunZ2JKXReg6F9Ko7gYjLdUpCYUaS0jI0eA+Qr/EtXisIkiLIbORgGIoQz1mso6X
Bk3/g9q8dmbBFwGtxJHRj2FIXJcKVQ0ThHp0bs6xvaQvMllA4JLR2Rq17lkPA3RpzPw2U9Iih7zD
TwVCukRF7sgnEuFjL+w+6AxTFpDLIqKa6r+LQ/PvPjQWQ6az3HtIoIu4E1/W/qCV5VZr7MvKMzoc
bdiuPoFSH30XfkBc0YX1JXw/NmUMOpBgsjYPL8Zr48B6Q2kZkW7pQIiLsAQZ5Eq9NeWUit63rjg7
bd3Sw5T3XJpdtjhiBoopVxvML4RrkREFg87go/hn+nW+Vlwy+AJneX/PMwZrZlGzAR/qruKgfgY7
HwOuukQI8j8xd3y6zXuff2atue4sWWhmTD632VdtbADScVKU/0KrioO7cc5MK3R5QO1sBmhkMeJl
L0OlNYapNi+O92NVEYOCyOgT/JzcKvPN/k3AJYQj5SRiEJPKRWcyfDBBz869K/eYlB+dKnB7wY4o
UbMrZzZ1WFfGg665MIBn7nW/9pXaifg8CBZSg9zdv8R3Ss54J5wRsqHZz0hLYbLa+r/5MiVnCc17
QgkKwPpIDpF5swNJyCXIBlE564Hr3b5a/M483t2AaLAmlG0HQkmDn+ODfPEwis81Uocl46ir40RJ
x24R1Em9R6+Kb/V8F75b/AGKxRiR18+86Lb5J/DQim41/FzLcHezI+Oq4RTyozDxzQXn2LnUb6q/
jX63fnbxF4my76bJD1bEZBIISXtcf4ecLvV/g7PXogfM/SpQ7NuYjNfNDnJnvUOTm4CVBVvCahV3
yQ4sZltf0mBvYwB8ZCCGiNK5CZ69FnTLbOguvPQAxVJA8Ah7qVLKW7Zw2T923AOxaF8YWVmE6l8Z
b70vlIG1gparsyWstDu0Kr6mXiitw7hH8vOmE4YkmOWlXvN0UgLcnv7m1XzCx294y3XexpeH3C4j
sK77ugThKLerLvpyucex2XCnr+WgO9VJkmJJ1xSTJfGS3E1Jt98edtiJQduU+J1lyUr8EhNwpYOx
8aBVbXRtsg8AoHww5DzfzeO+SeHcYQ16HEjBCsE9Mq5cAjA+u527yYpS1o8fmH5YDHR3C1R+LEZU
zEiuxgMwO9k+JumNyOWsLbTqBnTuFFiK/ACRLz1H1cyc9OMSQuUHAYlqubyVQelZFwnqqsZ8M9/k
kYqD+uUt/qMOHfKPFoDraoWK7xECANxYbRs6OkASYSAZo4brxKzSv+i4y7k2f5DpnhldJ3WzAtwe
gNFEbvd6ywpukfuL/N0ybNaDRVrR1bcXXJeqCUyNDPVC2Nx//JIjsyShoc0xikdqG0zmhybxHUU1
Uts2hAo99zhTyS8xC2pDBw5znd6pTwKCbvp1jJlbao0WXXHfpJ/7DjL7SBOxi5nHoy2ZE08crmKy
gsohUhO9byhGaSOhQDAdhoaOvLX47IVWjFD/7JtS0xIfzJJcwhDynYYxNQMoJrUsGa+p+ZtKwiGG
QWRZf3MQd/06KoeLpIIWfKp1lw/mbpgLm5jxMIOMlh+1+rNOF7oKqK2All7hVNXF/40zNGpPzgB5
48ocQhpfRGmxw5gK3Ccm62zCUFXCx9nju4H6jVuq0aUmb8tsJW0ehqkqJ68XTmGoXJCXCtheBmHM
ntrAbkqvQUp2a3Lb0A==
`protect end_protected
