��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����ǎf�@�}͚�|ET��xW�(����2u�y_�5�ɘʪܼ*�\w��c3&�c�zP���^��G!N7�1p�H��AK����s@To}��]�#U��Σ�$�w�*��F�c�Wf��/�5��Ca��b1��[��b����Ad�|R#�O9B��̓�5�+l�f��b�to��q��x�V$8�����={�P���ڷ&�i�K?pI���w&_��TL����;�O�w�pQ��.� �Z��� V��jK��9��N綷+��[a�C��S�2�?�܋�0�=���΁v�S��+���mz�/A"�v ��-K#P8�}O�]	�H�f	�?ʞP���up|����?��ıN*N��/s��$��w�"NY�N)�.�W?uJ)���Οyշ���%� �	�����ZK�
q�y�dC���=���8��>k���g�
�*|���!}��T�%��Dx���P9:�]#�j�	�9/�ǝƼ#¨���}��Z&0����ۤ]orG2%�"�R+��qU�q�(���/�7a,���i�2����+H	�4ɹ.�E<�ɉ��m��P.�`����z�b�L �O�"}u6�^xe�S!����.
#�jkXՀbYC����$�eH���jz%va|������k����S�聇�tNĵ������؋�A�v@��@��1^"�}�xf
	��3`1B�]����"]��&�����ki����ΤuvU��`>�C�KO�$�� �ӂ>��
�nG�E0�.�t�؜K�h,�	?B�Ix���ƴ�7i�M�Qe�Ekˠ� ��c���f��{�#����'�š��v�4��R-�1%zA��l�	?��RU���3��5�|]�6 ��T��\$P>��)7��Ly�m����m��U�ѩ~��m��8� �k;��9��7�C-XL��8��3*�דL�eP����Xx���0>��>W>h{9��wM�'��_w50E��\�Z���c/��T�,�G�Ɓ��I@Q\hYP�56K2r�Z	�%m�E'���Q8����>g�-��b����E���c�Q��
^��<������Xi�{�I_�.nT�R��PtE�܁�5'HD��83lq�|T	\�4�Mb�~��`\>b��H�c� 0JX�ċ����H0
Ԃ 蒫Q��T���,LS�jS1�ec�Y�r4 �}�顬}���C���CW�Qs􁃘�A�w�V^�~�.<�J�����_��M[n�q8�L�sp��|�yXq��4�kf���xӿM�;�T�/�̑��:���˅��8IGdr}��#��p6 ϓ��mX���g�"�N�>ė8���e:v�7Ű�]����s�F�f���LH ��he<�_�S�4h^�"��C���!�-*��k�h�r9*
��O=���CF/�>B߻)�.m���p��L?|�v���"Vr�#�L����wvLJ:2
�L�=�v����ktN��'�ҟ����o���6��5�p �����:<R8�5�������4h����[ ����L\�fՏ�~�c ��ɑȽ>���Yr��a�&�V�	w���-<��R;y���Փ]4��sZ���|g��ԗ#��ju9���-^��J�4(P�4ʎ��V�#���C�W/%i���b�kR��U�;[sUL�+/�a9��;fQh`z�8:�.��;���z;Q�>�
r��+-f?CW*]N��u퐹ڝ*4�����;y���K|�<8�'hYǀ�d��xp��d#�ې�����dC���W̥��d�f�$o�@zy�,l{wN�P_U�]PT�og��d��+E�c&;#~��Ā��>|3;!5J)&W�oϏ�JИ0�{�	rkRN�e����G�;�K6�&&����1U$���B\Cz�<+㶸�Izй�I�T��`�j��D��� 2b6�����'µ�wC+c,����x�P��2ӆY�j�:�< �1��S��B�*�U��aGw1��ֹ����@ͺ��Ğ]�\�j�_�_&�oE���tg��a����[���|��Sz��y8�q¡ع1���1~ja/�A�<&�.�Q���N!�Wj>Y���t�J�X�t���ĊtϒI��0��/F�cy��%��F�����մ��h�?F�b��_�MA�4��"����5�q����W~>E7�>&��,I]_�}�%����q�[VQ�D������{A�ɫ"�3�u��|SY����Y��^���'sΊ+�V���6=qT��XW�.6r"F�˅3���b8͈]��뛃�ic�߱\�:���=���+��e���k�����c��g�]�~]إ�Ht��J��Wc#��?�{�}Æ/_�3\O�/�%���˄/$��y�����R��ƬG<ٓ�Yp�Z�#tf�J.�6�).,͍6A�\F}"Y���k���\�J��H?�����~�032���&�)�*�N�#9�Bn �	�̓��BU�tߦz�!�9R�e��Դ@�^��o&Q6�`�q22�]Ǻ�q���T�k����h1X�|��5w��8�BR�T�3��|��h� �/QZ����th�@F��^\�<7���y6'ƹ"X�X�{vj�'U���:��0g^�7..3���� �I �Bv���U@����uW>�=�p�*�c-}��H��A>�$�~�W�{����������)�hlZ�ҝŸVW�(�6�Kb0�h<F�\��-v��@��B�>a��M��S�`���jG�_�'%���d��8�<�:�Q@
��E���a�ʒ�O컻Bz]�|}�]"��\�yIs�U1%0��Ю�k~���Z��K�эny΢׃sE�ܦ��ܳ��}��u@v��LU����1C��ju�=�@N��'޸��Rՙ �+Mh��cF35���ԇ��,J^�;�A�[��UZ�?n�P5o�\��(*v���9��)GZ�����z��76�����F�,P�NOvּ��+f�}0#51"�&
-�xV 5Iq�w#N���2�@�R�ً,%p.)����u�c��P��r��FT	���/�$+��z��r�nV��[p`M)�)+n����|��TU�aqt�~�}�ihx�TqrC�8���C���ueW	bh̨���em���;_l�z��x�ȅ�� `S�����6�MF�ǌi���w�W�)�R@N�5�(��[�ɰ�V�VEI��~�Hf�fܧ�Pd�&+I��Q�|W �X�^�>�,DC�&�9d��-y�-G�����Ϋv�?D�Bt�Z�����=���O)�+N��[���¿�F"�!NtO;�w������?�e�O=t��U�k�UQ{8^t�`�<j�/��jm�'�W�ZM[J�b���/�Xr�$#ֱ�7�9��o�}�.>!4�Y?���(�� �(0)�z0s�F, _Rd����p��5�|�?1x+28Yv�n��2�$�ֽ���N����O��I^)%|�<}p�8E�ڞ�uxaf9���W�w1�\�J���i�AO)"f�14\�m�,�м1�2:��3J�X�3����I��*��~*oPbz�d�xU|�����	̙�3MCk2�eH�+��ڛܮ�f6�==�����(�n�u#�������]j��gm�&Qj�YY�<���7'ޥf/�NmH}�r�$n4�ZS*� 	Ը׸�h�4��RY.��U2������A��q�����������a��=�3��s�Sv��He���Iٰ�p ���%�ӷ�@�)$Ġ`f���"sL��:�
p�SBߊ�m��:)ϔ�j��լt`��2��n�{�"7D�{�#_��R�*�����$!��釒�W7�H���i��pU�� �^!��\��o�rv�^l�V��,z����p��Z���F�G%޷���)�g�o�
��g�	G����sw��te�em�d���e�{�=����UI�A8�j�Y̥�� 4i�F��G��'%��R~k�N�wv� ='1�';��FXp�g������𖾯L*��o'�9D�4�����#�/R!E`�=+jib��t�.$w|e�3FqQ�-��e���k5�����#�25�Ï�D;�I�
�v�cD�V�@�q�gHw����/Zy�t?W�`5�yF���7�~ �܏l����r��g˪W��%aӒ�YF5yf嘱n B�>*~-J�.�[���_�g~}�p�#?����]z�~�)��TƐ� �ڛ�W�Y�E�*TRe�gI�O5\��1��oُ�&E��ga���,�d���D1f'��~�>�k�3��B�{(V�St�!���"~~F暄�9O�u]x�A�~`�p}�����0�3&�z;Q�O=ձb��_��X���`D���"�a�����~0k�Ij ,*��#�4�-r!'&���\#1
�[�|�S�sB�c��N'��ϳW�g45���V^Q�O�ǃ�k�Q�M5��;��b\���6Q(\(I2�B�a;R�Y�X�W<0���Y��y��ǿ:r&�t[5��/q�8��.��\(36Πf������eʬ[�cta��;�ä���3|.�3a*�%�S��(���R1V�������g�:�v������\�w�Z$1d��q+�[B�V,G#�bh���A���]آ�A��+ͧ_?�l9r�j��x�;&�����{�y�Y�a-�]��VKn�B��f
	�r垜ΐŶ��
��jtT#Vj��,aYXc/&p�9�V���;ʗ�#\v��oA�M��0�쏢���8�� $L�)��"AMU��T[,&g�o�E$�7�������� }y��{��F�e�⬍$��{���¹=U�
��I<�%M)it�V�El����%��o�XAQ@`�~�-��X_f�
�`�-�5�n4&������][x9���뺊B�,/�B��k;R��jt�r�||��9�
���u�A�4nx6�D�� A~vo�c��"k��������	�!C�ڻn�8Ojrk&gԏ��9�>�H�84&*rA?0ĩ��^�|��)Ƹ��WwC블��-i�}�j-�s�:���6�-N{E�IW`���Т�\):�7�ۗa��Dp�Q#�v��֒Φ�q�Y7�`�j�Ev{��P>��:\��?�����1h,ɥ\��Uu�ܘ��I^�r���)��x}*�<HS-d-���E������Z�¢�v��2)��.����l�k�JZ�o��	�xMao��ԀHnL�,ƒ�c��-���_��S �3`3q.u~:��p��g�C�ti
�!��{��;TYR�ἓG��*#�4<�úZ�.��{)��4����7)��9K�O!��G���f�:g�YP�y>t^U��I&)eR1P�'Ʀ��
��B��-ht�_8��6q�P`�`gȑ��7�i�RmZh�c�	�Q��g-������db1A�s����B�q>�gh�*�U|�����i&
�!��h��a��zK�XM];G���5=f�K�t;�,!���,o��w��͜��	��3[�� ,9�De���L,V�;;��󪢵�k3����G��e��"�R��j��7�&wE�	�&x���[���PZ�q_$�%�M��o;�z�R�k!/q	�g�w�#�o䴵��i�3!.o!,�U��u�j���m�
��^	>�>V�6ER�.P�طM�̔��N�?�!�2�0!=���C�s�g ��	%�kG�X��8_���]6å��Sٟ�&"��`��R!�7�9�WI~&��l�����"HEn��8�����]%X��
��K��
9�Z�=8t3s��1G�71*Y������z�%�p>�4>�My��V#*k������?{Vբ����D�K��9 ��"������O7R4��x����81�D��>��Xؼk%���1�C���,e�����>��զ���$&�W���9]F����͍-�'����;33�p��Yp��:�%�%�&���AV���:���U�:D4��^*��
ݻMn�߯�.��$ˀj�M�zAp��.�9�&�A@��H.i��Ⱦ��<}O�c}�Ԧ����X,��hXf��������}"n�|b�*"�>W��:פ?`eG�L�)���[岃�� ��<� ���R�3٪�
<`5(c;�li>&����� HQq'�߳�)>��R�'
�G�f�7��8���tä�ȧ�@8����c�`�l%]���Ϛ�H��;�*������k�!Ȥ�ܒG��s�i[�|
S�D�`����=��t����hW�����(��5a�H�\eP�c6_��.��f2�{J�jp�v��D���n��p��݃E���nT��������8��Hv�c�?�W �4&����d�
-8Ǟ�$k�%7Un&m1�@%�dJX�J�*�p4N[��s*���'���@��Z{�,���������y��L��	��hr=؀���>V��Q���55�� p�L�4���z����Ǽ���"w;�?��s;��4�Sa��7��A�М��\+uW�\�J�8�Ĺc����{����$&8D��Qꆩ����AY��GW-��zG�~���<i��s�z:Ք��)�)��ǭ��F
�'a��kq���e�*��uʼ���`�jB����oMς��
lhD�ё��(�\yf���2?+j���;Q,�6^��Y#�q� �YL�&u���~��7/��%l�GJ���}�%�Ey��c8ǫb�(�dk�@6UP���FYw��c�׆�-��Z�����j��w	)���� ���4ǆ�d��by����t9�6��c>j'$�Ŷ�.GZ_xM�C�a5��3�8�v:����<���	�VM��n]I|����Ԇ�a��@@4��6��v�BP�\�I�+ҩ��VU�,G�i�Je�'��\<�Ocظ�V��d�r�T!o��c�>�X�R����,0Y�^sD/�T�I�fniRߦ��[J� Y��� f�*���L��Nr��Ψy9:��8O���>��שf�'8��&cuy�ieN�o�.�x�Eh����W�I���o�Õ�en��${�	�43k�=N*I����9��k �c�<�m1��*|&X�7����PLW����ۂ8�mŃ~^�:�d�4���_�H��9�R� ~����"��xl8c��䔯Y�	~	�a� �uũ�Zb��6��%�yL:��;���L��U��J��4�T#V65�*��nG���C�SЯ�!��P��X7r�d��m榫1�6�RdM�dcc�X��K�
dd��y^���،#�wP�J�n�̹K�G��L��A�6�^�	���@�8
��v�ŷ�����9o���o�:�!:��R�����Yr2`2˫���h9��C�9�����,���l?�E��͑�pKw�|)�f�.���ʫ��\�v��t��t�
�������x��4}����lnr�f0�O�9�Ǹ�>�HxS��Qi��c7^��$&���=j0�S��}�$�s����l�Xn��(��f+>]���+r"ܦ)R�w�PnHW��J�=�Ew�C�$��e�&	@��nVM�0˫��q�p�+�
�ʈb�HN ���Г��S�.�&���V�g&l�����Q�<�y^\��~�[�_;��|]Y���Bh@�>@����pW#���Q�B�(�����L�7�C����s��3]�q/�K��B`��+�5�Ŕ7rR�SJ������.?&"bu��#�A��
H��ވ�^_Ĵ+���Q����}��κI�4�Z^_���vVreP�P���lBZ�nt�*�c��n���t�_��{���A�:�pI��`m��祿��R`/�K/V�i\`���1�V	�߭�qa_2�r��>�Ϛe���>�;�tO ����0��3A5$�^�кuG݈
 �-�&Jȼ������!�ҫ��v�{��v)��EQן�<�#�-(Y���Ma��0��9 xb��V��\̵�������7%p8��Å7�����y{�H"�U)�B�`����U@(qd>k�r=����Κ�7+?�h���sR�[����2|"M����6x�ގ�A&�h�P8=�O��4h|��M2�r�k/�f�$�n�G��\��6+����) �����A.cB�GO��r[W�D k�xe=D���f̻�{�-Kz�0���B�8��-�Gwf���iL ݳ[͸��f�w%��t�Ec�,G��|�H���/^Xe����i@�%H|mx;�A�D]�#�WS-҈�K���Cv�7�@,"�H�|�;�Yy�M{� q��ݩ�N���F�33ޮô��99� >cOY=�����!E:�{[P�}�e·�=����:C.�zw��Mc o���]m!b�9�6��;������l_���U4�����TU��GT��l�y��r��-K3���vX�>��t���[W֪���f]�|E�oJ�����ҰC�ظ1Pٛ~T�-��9&T��xv�}&YW�K��ӯKT�o	c5��UqT���>�z� W�?��[�I*0�>2�4öy��Z���2��<����+Pu@<]u�y��ʦ�B�m���uS:g�t`��+��؞�]�?��I!o2Z]��pƫ���(����hez�jk=�e������F�z|���f��hbI*rӉ1�����)����C͹�!����}Tp��%��dB�<�����G��6���C�v�:��Cb��0�QQ��H���0rW5g:%jR:�5o����i���qx�7v��-���&�|��H\ᑮg[�Os�$�R��O�Vy�H�SC�`�gG/���4
�e%����^:�����$pf͑��c�r�	����V4%6���'�y�ґ6KAp���	2ͣ�q��gv,"ŉ�����oJ�fX�@⓬�"95Bl���!�c����H����5���lOnL�����K)�9��92}Y 2,�i{vs�Ժf*�1n~�;�E��������uPg�ƒ��a��-����:�H���1�H|i�Ͼ�3��{���o����#���a�6�3��mG�T��6�r\�*�A����>xZ�oԐ]B8�Z ��Ry��(T @��Jx�.�Zm��%˧�tR/�, Y��pd-A��
V�Y�V��9-�+Х�zz
7���
P��Ő�t'vlb���B���M|��������v��� ����r;���F�ь?����9.
�3y��ЭͻI1��!���x���^je�����P5<�n(�|0!� k��|��'�kڕ����T���}xY���u3��g���H�bW��zf��Na�|�e,��
�"��m��;�W4�]��aT]������d��VG����q����b��U֣TK� ]��Y9��⥵ab(ΫF�9��$X����5.`�u�6�����[�B��{ �/�bp>�v���3-��W������&�v՘N���\��s�;7���#ޝ��YU�|�0sK�����y �%0(�I�s@괐���Ԯ��jI�स�eG�g�0-��x�S{����l��ɐs�N�[��qC�Jf5�R�1T�XI�1�i4�{�h��D��QH�6lO�=�F�a�L=)��	��̕�+�]ֵ�^�	�����In�^�zet�·�t<�
;�]B�u[�Y�Q�l��Ɂ��65{�C���'S��O�Zr9Qα�5,�i���[��9��e)m�$��~kxm����Ѣ=���>���{�6ٙ�}�������?p��� &��=��=�X.�aTMH��T���c�� ������M%�&7ۘw�H,���S���ki�zSMma�*xݼD_�߶At_�Q�K�,[�K�z�?G��S6��=�((H�8��������'+�����2�A�7�7<�&<��H���ʭ�!�}�i:�R1<��77��1�~w�;j�Z�,��?J��B4`ny*q��8lL�n���}͋^c"M'7(a_t�)(���	v�0��q�0��W�nq^��>�_e��Tm�hi��r1��E������E%��H�e�\����{���/�R��a��x �<��p) =R��FR��t>�~|��nn��̓LL��j��9���A��&�'}�t��-h4�e��c��<2]��h	�˔^�5�a��k���Z� ����v�Ԁ�3�q�B8B�mBj��Q(��Iα�n��a�i�Z���� �&GW]�����;�lLYn"ױ��ޱ��D�˙���4E~�ǻp~s��b��8 kˌ'����+%���6��/ַ��f�˨Nc��9�Jӳ,V��y��ެ�D����f`��IIsm�4�\#$̣i�"C���<�e�o+��z��,
2�v�L���l!3�%`
I.u�͟[ް�o��p�+���A�����s�b��������\���F,�9���r���o�T����ϟ��7���5ޭV>��u���?=[��������g��f2�.�V��j֣��H�S���y珕|�&^$�J_�3�ƻ7$�fp�v��g�E��>��dY�%�ld`����g��6m�h�o�$�^'�����)������/���cW�Ϸ��ո��FQ����O0��xBc@iˮb����1L0��y��l1�#�j$��X���
c+u������7X�I�t�A���Lԅ������kq��}߳��(E��T��	YXx$Ew�R�R+�7µ��#��VĠM�|*��$��E��M
���s��'�D[�	x�hi���V=���Z�X�F	ݐծ��Gرs_MW�%���{�\%"�c����������7�-�Ȓ�{kE�iw�H���R��B!��<|���-a�'~�ˋ�:'���.8��	����� <[e� ���C� �0��+(�j_�a��/�����\>J�[T�}9H+{�����}!�NȒ�P�γ2�/M�����R��4�Q�%@�I����?D�v@^S��M�?����	O(����A$%�L�H	���$�ͪ��|��C�;8Xil����k���S�B"�O�6U��*c ���W(��� ��m�u+F�<ZKU�s1��ʼ�)�f�+gHӄ�a�3��ˣD	��^�e�?��:Ѻѱ��}�F�%)�Ũc�@$Q.��M�[]R�PN�-��e	#�G�j;,.<����o�S ����r��F�x��4�"���}�㭍�4l7�����,�X7�h�"�g�I���F�.o!#��%;���{��7���K�dCy�����q=@>����#�#HbГ����Lأ��jVM�7F�? a�lx�1��3�jx*v4�96P���s&%�}���/���1�_�h�5@Tm>I��c�,�Zx�� ǐ�[��o�Bo$@q��M�a�ftam��&��7B����C7E?k���R�}P}��|���dFm��S���u��o{r��