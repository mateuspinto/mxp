XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����������Kdz��X׷]EVQ�ܗ$�h����W�ܻߛ�ޢ�B���zD'!ȋ��Ѕ 3|a����J~�>�m������M�A��ht)�4+���w�/(��l��9�2��z.K�'M���oTb�e�<(�1��2��Ҝx�K��u �y�"��c!XIT`�����Mv����o�/��K�UW�"g
woTp�f� ���5��|�7:���}k-�5=,�.��W�xv@�;�����O�w+�<:��:�H�b��U�޻��%�v���tl.rK<�����J����eoC!w}ڻ` � ���K��:�(wYڟJq�F@�[���zY8T��,z��Ӣ\
_a�SMZ@t��n����܏X�a}\��Ԁ�	�akΡٖ�$>�:�I�E����+�zq�l�{?}�j6��Õ�_���o1��	��ڼ�H�c2F���	�����s���C�[~�H������؀KAȰ��բۖ�u���犚 ���s�1r�Y ���Vn�)iS̵�͇uу3G�#<I�f�Kn&,9������嚥d���*��
e����%A�����fa��V��"˕�ׂ��	�j��f��6n��>�~D3#�hԘ S�Mo\�ji'T�,޸�d5��hjW/g�Ao�D�<��4����E�(� >������+J��C�T�g�י�������ΟV���B�~�� ���}HkW�	���c\�a$pE��u0TOE_P_s��� ��H�XlxVHYEB     400     180hӈ��AI)�!ɢm�����5m��a~�S��H�5H���X�*R�ȸ��+�u�K��e`��K�
u��PuO�Y��#�ʚ�7K�e��&��6���)�w���q�DC�Exh5=P�,��N<D]�!��)�D.]=�/�U3^u@��	������æ췳;���:������u���iD���忐�0�	Ȓ�qP��s�ʳ�r.���� JKh����_]y7���f�g�4��w�YC]f6�ǡ`�j�n'���r��ۄw6�v�b��2�x(V�����ED�{)d��6�##���6��kb�o.��1�KZA�Qx��ɏ����rJ�q�y�"d��iz�>�ȔS�+�qx�\3�Y���6�����XlxVHYEB     400     180nc���-E��AňH�����N����!��Be�	��s ��v$��������)C=�{�/a0��GkDO�_ܰh�E��3�WR\���������z ഛ�l�o
pPenlNK��FYIN�x��(��]�T^"3��F�쇼�v� �|hEے4�z��� �N�Z0��g���z7K�Ԕ� �@f湄L�����_�����"ZYP�w
��v�(��$�
�T5o�r�"�6p�޷p��an�����m�q�q�?����X�<Mc5�43��
篗SV�f,��W1I^�B�����3�C7���ϋq� ��t$��L��]vF!���p����l���@z �P�]��\���S��v��XlxVHYEB     400     170>�EB��G_��	*�!8���'B�|[Ƚ��;KlAWa���+��v��.6p�F���������΢%A��l.s����s(�ŝyn�m(���2��V1�K�]�Hv���&p���y�?�H�e$�K�@�+*�y�'1�� �'Sz������k�S�]�Vz�������/���.��!K�_U�$�2D�F&��;a�_Ch��F'�.ޑ�`}~��x���ǅv��H��J��̅5?`r��q�����F�K�0�{�5�j��Ƨ�8�Id|����PT3��	%� ��h4����fkس_$4�/-��b{�V%H�X�g/��_��k�ݞW��	`(�5�m����/S�iZ|]�1�g!��\P�TXlxVHYEB     2e8     120��u���/YLg�� >�;Mq'h2�����A��zTu�x��B� ��/
|�9���(;\���
��b���z�Y�BQ&Z�,��򬢒���Z�����KIF/���G~�[m��'��DrxN�w�YWꝦ��|��)S��EG#�dk��#ɻ���� �*eYۙf@b��) ��x�=���Z���)�<�a.��6�|�*a��eA���|#r��M�ڽ�A�kUz���֗? z��=�B��1�Ͷ�s�v�1�#@��!݋���Wc�)�@�4mݏM�