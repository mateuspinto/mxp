`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
hWPMsSHVlQQxQpy4MI7ZcVZeDQSSAgJJKcsuy0CjQ8E9KNCEkGpYf3UTJbuje8hkq6HkRWmX1aBD
sh8Xgd7Xffu1dRSIPRd9Z45HAgEM5LocBCjJr4mqBOWHL/7atTy4u/sWI0+YH4EfuLMTS3dsyWYk
chC9YWkg5e3t/rci7rFKr6zkRGX7QGDE1rZKg9c8AjvkV3z+qeyKN3uJ3STWSyNhz1L1PDjg43Oe
s4cKs+r9ZRg9LykrfAzWqczLghVgPIBEY0+4BhnML9NY6rKntenH4Mpn1IgHwPwrKCZSswzCs4Fv
oSp1jIo9LJxQHKpZLSqiNffcphG+r4qUvw/Mv+RJJso6Gh44QoTdjdsc1N6rVXArD5zspFiHJkfc
yurte1z8HgIkhNBVuUt4AA1b4ZGX+7ReNEsKewKHCQHkXJEAQSEOIsbOu72aHhGlNtHnSrqcIQMz
qKLfzsJLbhgnS3gevpty8kkGJfqaDtAgR25bZ6y8dnE1l7OLI2Q0HdvwBXdDWOL2JBV57LOeOzpI
fGEL8FOhMfD8957Xffs1B9jmDi/EMhuTTOHRQUeJT4MSwmNPf904WsysFttnQpY1HxX9RN3pcjIg
6wxWCyUWH4+Rd1AqpI9PopbJLxnexOFmKCA+WxB3qqAHm7UjTHmXhpiLKIsO7Ks7pPvFAf4N1ZsK
1Wb/Rnf8b/x5IZDnoS81XIw0Qkda/O8o8UPYBhajT1cIhEi/zWWo627ktkzzpyS86svdtM5l4clg
1RDG66oTY5+O5BIaUneNnojqDP67sqcloNWMkxlKammW9I7Mu98tnyhta/t2hGXWjwzRW/+X3ZxG
yo0qJLcEy3cd39LU42xQ6BTzAVqp4FUW17nLAOpIwITKZDkLY0mUGqUlE9lUmgJdCnK9e8v5kW9I
EEnuHqe5mZcANr87ZiefYMWV27LafhVDb+WN3Mx1GpK+z97kIv+NontbG/E92Ns0v8c0nYsbhfa1
+Wz/D61Hs7a5vp6sSkV8j4iYj6DgnZc35cqy4eiDxieXA0l1d9C1zQYXJ97w3w9rbZdTEl1Hy3LR
sUlu6N2ZOCKwZq07Qnk8+KC6mJEBZIVOfQgGN/59rWKnn8lOgYutF4yWgzpFwFUmg5ET3o8HiHsj
0Vv638LL8fUOy6ebIuf89argp2miEwLM8iLPKjg/QY/HqQTLZu7lvLiMIbeeP5bq6QUU512pfx2Y
x4x2+F+eSABsctFlEcDoO1coo2QMfbkjoalgkKtNl6GTaIPPGsSvD3YYX+U4pw1MAwnsMgytnJQ9
ZsXAM12NSwbbgAu+mKOt5B9b2vLIbtrjT7oO8GLMAtYDQP270IR4gvvLlqwpQZuO1rxF2krcmSHn
9ylyJxf0Uu9aJB/FF46MxrjW3noaT9Ua06qMRK3ssS/2r2cYHOULfsI/mS/0XBDGl1DcwEakcWas
HHvZb6A8WbO4Uh3GWftTEkhBZyizXbG5WHaw8hsux5KqkLNOmk78xcoS6Z1lO4DcrxshQoCy7rC5
z1+2TynbPxcyOIxQLL8KppV40tLHPRwGnPsgkBFysRovnn5jZ6wPhe5b9+IhhQFUUte3Mvyia6pS
vfyV3p3D2bSPAo+zV+LN8FucKbd39A08kl6BUF/pzAYyeGTKMNfCpZeZYf/+4AZCdFEstAnqTQ5E
M/OBPFMFWRQdDuovHWcpfAWU3Sn+aX0yBNs45YSjPc6tmb10vlww7LitDTthFYF3pV1FRlavIdmT
MXNMrWBXhreuzJR5YL2q6noU4NOmUW1yA4TFUHzXefVlLwUDrWdaTEP4RpJu47PhE95N/vQBnYYo
6c5wrXr33szWi4rp43UID2OIHDPfSEf3H6+bKqNi8DR7/HfLcv/IG7I6iTVJavhCZLXUPKGvP8wH
qICNZuIS9SizCyiD28FsGGenDP1AfjDuae00cNomWzOH2T2xEly4sXRq/e6vX/76PyaEoS+hlJta
NaNSsjSxrZgVZ2ngbLm7+JFlNVv5naHC70FGADQg4QT72rWskppRngfKEHR44vR71jzdXSaRusU3
1AmR2ZRDTvzT+aj4pg24t+0ZaiRNSE6CCK933GFTXAjB8SyPe4vI5S7DH3Oe/++v4ylqkFUnYG1J
JfsnfSrp3J2jrhRBMc41rGrrsb3WvPyNhImuKpRMf5meRyeRdFY6gD3Q9F3vJx1vEgbx4GWccC75
jkb3d+OkD94OzMjcLtwVy+MVoO3tIv3WNxm9oH9cAIXTok3K5vnUQgA7X2xRX0HFMJHF3po+SGKE
2YnB6bVZE8W48WXQHac9t63X9rm1GvgyEbwjnA6fAMXbZh2GBCWz2/Lw71ekm66SsT7ckqrTx9zC
/FR5rS1FgWhCwJ+VX49Ox/Ao9v8vhzdnJ0nOdHUdJZ4YXr2M34Zs+ZzB/Th+guM/Gw7E8ptdqknu
to/nxz6D19pG1svIwB841iD8Te3KwogBGDydHm1KBoigKdLGkuJvMLpxnW+oOyiviwJNfD1RCWdA
Yt3mMAlXab3ONDblPOX9ZCFrMj4jks3DdhRPMRO/SF8w7nGjdkVuCmzvFgz8u+LQWu/kxcdwGBUA
jsIbo7ZiW4KCtuqNBrnHjbqNq1NT3Yz/7l4DOhe/f1fwNrfLNcMAMFxIy4i+cKYXwjHR/XqlQTCW
YufnZ/E7/ZAOWptRhYd5WLw/FO5AHNqaIsWyVPZuUyl7oDWerv50YZlsyVBdtwVC969qRuOMgnyi
hCG52t1RSx2xH8+CkZ1RqqXg8PxTSSq7KULm+il7iEdRu77zG2yIlWLOAKmPYiOC49yfW+ra8Ui1
0Hk1HEGKyzdkRfEBziJKBhowO/FIL+HYvzMHMoPF/8vy1pRoI1kcf7AyDmbQ3Poqvl5S93M1orqS
MDl2j4qE9UyIGhccUMTaN7GuI3hurUBNRvJYZ3dfnyJuxfhYPDMFWILMVkm5Z/ooESrEVn9/0CEY
bfcTja/2Wfqf/GSmHV6K7iM8D4SWuJDiZ7aatuynLjwsyytrTZuamx0m3UhFoUjYpTzRS2D2VC/F
z/uqEVNww44/FDjygqmxKBe5gj9Lnh5ddRmAB7z/lTffoKqqERLTOrwHHZ+y3cbbgcJCOmuT1myP
2iUX+wIWpDc8u5wAJJO1nRFlIC7vArSBm9Y6feTvgB5V3x0jH77y3TSBPnjyVRHG6Naz/S6qa+mQ
2unJntevmoQxr0aXCH8dmI1KJdKbG3OaZsvYAB1SOK3zaKzYEyA3FM7ePiEY7gCtDxuoG1OmwROd
KDATq/MiRdO86i900bWCPAfru7PHgSOt5+3WRaNI7sYU/AzSC6/azIa5PGAl06NRyQIwDZ6lgbx3
VrJnmCmDmgTvcju6LRRydd7umqJ1wRGlRCtli9bqu5GvW5Esfj901+8kGo/eQrplJGBX39ie0k1+
lKBSd7Ac4cI5NbUl7XD8BAZqODfjdivN0TXzmviVo0yMwWBbN4gZmkh763/x5nGC+XsVdCRYu7hZ
wpFf7Sgd//g2ep9YCE7II5N2rJlY/MCV7r3Yx71E0JwJ+h/5KUGHxDTDhetVhJT16/wBY7R6bAZ5
XwNAFLsziP1D6/GMMMiBZxeAYPZXiRZTQ4We4ZKYJR07waSKP60Wy4PKOnyhUXyWv0g+RJUgon2g
jnrSsSkCoZvp9OxnAkWwhSYLzGsulAakqcvycdliUlZUjBS1sklAteEsnBHxJhx9EBMnjd6MFL7q
UcspAyjXrikT8IqplqaPz6xFq4YAdXcgUi//UgclZjr/aRHVVCQNbgl2vCy+ERuj6z2GNXvcBqMc
hDcUb7lxRA2X4Q0ZMYZwS6qPlEBGr6fgIaJJ4nhhILdV0894R8R5I9klnB9HvMJQKGS783NaTV9H
vMEYs4ACk9Qe8KsLBirbcoFbh9lNXuJpKVy9wznunI5eBC+IT2eiyjXAvSU21L+jn7HsfU3s3QaB
XbzQf0RixH68HC8lt20wPH7IwdoOpN4CmBBc9HKZ1Us+Z1jcC6rrUjJndDa7NPp4bFfnOU6DMn/1
+ft63CzmIfS0wcBiRKdhb1C7s7uvSUXj7bC92kt6LfrMYk/BTP+0uhv2DgZBYXN6S5tEgXYKpbJd
mb5jYZZj9R/fuPQbZdMeG8wHqFoWtilbxnAqS9gLCjYg/d37gMJwK0I+ch70aqvyYSF5tHmp3TCc
Za17a78U0X0VSG0Vl/a/Hhu28mKkNZN/zS2FbFL6UeYrfoRiyq+GYnauueSQ+NOH7loEBNN7Vv5j
DrYmgeP4k0homP0rfIpWmjU+1VW3e3pBVA2DyxEfxQ4+Kh4ERoZqDGofGiMsx7p5cXKkZfZC4B3A
19+UTjKs/fYAdLaG9Klg+iuwCe0OKYbw+roSqgrOJXP8N1rHKudEDjWgTskNlUZhMJ5yJvPHFMJL
ybeEwA/I4nBapVQc/WygBBFU+d/XdKaPejPx1re+YhNheFraooHe43aebBuvTPMKadJ616O3o6aA
dn/a7cCTFVL9L6JwEizFM/+K1mOPK6x7vFUCsAjil8Q3pASmY+IUQdV+1/1LJex62exMsaUbT3G6
jowU7ADD35a9zE7I6tqtD90URQe+UWJIhnSOk2PtmTxao49I+nYOxa1s1Obxh5mK80Id9bN6O7ks
1jpGb7jcYnri8k+0bNENmwfxOwrMGDIDACRWLY6XN6XpHQ8/5S9pxOYuFE/YHFGyKWatPshHRuxG
9N+wpOu9U0pHeiTCxQSzaXo6trzqbIKUkCzvZByGuapy6tDZIWVObofkgeJmpIQY0+/SaNPRzA70
uce7cryzfN3NI69aqpuJHX8QMhCPxkfUgKZJwEnDmQnX65lQ+OgQS0ip7/fJaZAh8E3ui6m5dpNR
ILFq6RRm61T7PSqoe/hN7yXWN56VPx9xGHBoUVEaConDzt0HU4jkyUC/vEjnpMsmKbBTseJd8ail
LyK4EGO2kfkV+hTPoRIG+bkf5CS048fxN8mi6Wgw6xejd2mJ0YuYINyNgUBG1n7YzmRbg7CxVZZ2
nS2PgGsyFIipmUl1hROnqru043b+8b6l/Udvvovdn9EZ9GKppkx86Y/3V6LyOL0Xsq8F70UFxeXx
T4Ph70mhQpqU+oaMu+9rO7VwGXtM4DItJjpYBN02Q3yf8nfLLuCiEO57mKuuvBNXIl94fryxRpYS
hEmSB9X585BzmgOAkSwcScsMwW6E0cunKKxm+XnnqRk+PUjp32vSJc4nR1MeCsvmdkBPyrr0BivK
vlGmvaozyioAEUcGaFh2C0mMQmW1JwDQQARAedHPGA6VKfQARsxiMCXztMw0JnplxiCTe2ZTXPDQ
hf7tKOj/wdIw5QNNxlVw//MvXKTR9kqMA/RL3xENXg0QHhGY5tiMwJLyNgHI1JZTbna/FM4B7H7V
CbOnfUxMJSP1flW6UIVjEZRrp51tuG8TrF0qzY/YHuij++13dGJ841SKl4WNaOvfyK2/LIZyZaUz
b2FB1+LP4u08jWVdhnUbV//kKH/PwbPE+/U3S1Bc/5oyb2PyK1NqNW7IH9gmrPdtZ3D//Jzxjh4c
PXvN4oYMAyVrCXNJYoBnNGk3lxO9w7f0SQtSzNt/J5W6coxVsr8Yu05HNCcxF4nwTkWcCMvobq2b
b7oZpqSn9NpAn0L2E3yrHDWra/FHUJ4/DsM8iWU4CQCG4j6QCRdbmbWEui9BsGwv1ga834CHtRTE
cT3Nrpu1Z7sP/yTAhDf9h3KmPAvUkYvYyxnEy9kAiaQ9b7JOhU4mIBMgg7ZXpGP+ZZYwOBmoAY40
gfRxf5B+ALD1kL6H/mdi3SN8bK9Fj5uGspygmeAIApojovlb9AFBAWxkIJ+F2ojys5kUl/22Vphd
KeEfeqIIU0ay9SX0n7xKs/8bqgvhIpZOGjS0Mt0EU+EGZGZgMV3auoj90Da52lnY2Dcuh75gbpMX
qyPc5I+zAvRJT7uhz0ka0XZNw16bk/wxDzLThtOJttPXwRSYIa0bTOa3AC22Z33GYcsAVM4FYsTt
ETvcHFtFQ8BdIBCXG30g1yZPefaqP8kYTz6RRIQ701ArryY6RELdTk8qBymSGhXU74x6t+psohCG
t4/U6nkcyVMWrrCT+17j4V6xMdHUcYqg73NO9Cj20YcfMecfB9QiR5N3IYh1rzgjNqBjrX8f9PQr
5IESWmAHzqdVY7qz/HtiBwO42SYRSnXhY0Z8bskGXfdi1I+UxMGeMKEQm1Dqb3b/lYBVrXTfWhcB
ucyPC530xbnvPrwagmPJ5uNrvRIVLbW3LBAvDDLNIV44b7nSnmZtLXUx7eHheOYuw1SESwfpY+pg
Saarna727GWWe13uTDDccUEScd7pVKRZ3HEpg6Gm754mQ31pNj+x7EBL9wAHtAR2r7/ku/D0nQmO
aZ/iOYKHmdcoOqJedMC6GVwmLfYoXJIdAe07ENqeC0bdSY6T1GgBxQVtT9RI++KKxIhnFLXwoPw9
MLwLZf2KYdHpLWoxuCMVKGCAEVqbVBugY5zYDImP6Cp31mbv/MtEFLylTJ8TC5+zCxHXPKRhgwfP
UXG4Glp8V1YFesNLMXxW1D1NCCOhGudOxCqeL2P0IPfDvoeIUQccUxiLdIWateDCRTcfHkE55NFt
WzVizjKq0H+J8GtdH2rPZpZqck1A3xuQ1LufP1vORPp7Q76dCTuqWsw13Ll6dm7lDdlzoYql/UK4
iY5/9dg1GkKMzMAZ0IBCTM1gluccgDQJLY1KWSbf5m+OWKn1zIfkcEF1JE+YhjP5N+nYOhAouZq1
yE7uf3lB5Di+29VLmDInzqc2GJwHHtA2pwrvU2O2WhXhrzzS/D8PeBemrHhzMQ41eDira+FToAtm
jv8idQc+p6GSrDegE2jvDdfpSjnplzLfUfLzI1T4ifIwlJSbJLktprFMf8+gJ/NiSsWNSbVH1KnS
G9Qg189WtxymLb5P31faekokdg/Tsz8Hs8zX33ufAJ2dK+fZEtrlFyZLT4ZXRH6uDI8XP+ACXlt9
EhT8utNoWlbe/a47f/22xSkmyLewm019taQZx/T7aNdtTct6M4RsJWs8bKwMSxYyBS/foz2Ahlj4
Rw5NTw6mrLwvPxCYK5D+aEq4xc7s4vI9IOS5cXleQIBadiyb6DIyDcu6/eHvjNDSFxS+HHdu9B5I
0djyFNIyiDT3ykdQe/BFM+rujHOjEUXpRdrzooIM7VNhSl69PLwVhS0M9CEE5OIxUql+jjn2KndZ
UiwSqdsgqL4BSNR3dX77fZ03hI+bbvtkOqicjypsDZP4Z8gX0myR4UVW+NK/d2ZfEBoygujNfh0o
RTRUsU4MtsyTI/nb4dDa1n9ZBjTe1w4+2Daxyt/fy7FVLrsnC00Jf8AQ+pukoXstUfLJ54JBTTVN
1zoWGs32pq+J0jVmfvcA/AFSRw0N/dDZK27AutvMMJiNB4BWyXxFaIDtuzQzz8yIT+SjZi5waQ5r
/Jqdi5XCRUXV6lJ4kKR4KIirGp1D4BEw9Lb1bns9ORrtyUrf/4/AEAH2E8GseMQT+qGnSRTy4C99
6P3Sh5Nyl52feqeG0zjq4K/OKhMH0rBB2DZ28yXkSztjh3Q4r/stM5E3/hmvVCdMEYH/ofEQ/zNC
Z3sT4XZExZVI39+eOJ2UfsEQQLYy6TrRGQdLiPc7WqMXo0gZ+lyL3fw6fX+FcN7Q6hL+yGLBRKm/
TPO/WwHrXc03ISLf2UHugWEgJ51Xbu8yVbKAIwWBMzwyeaJrstS30yQbOR50yVkfl2zp2p6VL4b+
tK0+0T+nL4uYH+aEgsr5x85WWL3fT+pQYxSJLs0/HFPBnhhgI5uyMSouejEEq5ezztcqdGNnu/e8
ky1yWVavDyacVaDXiwvmDGckRVP7kvFidwgtHxAxUDgW8EB8dJDjb11/Ofz+sYiU7C0nM/qJQPp7
aIOtzad9SlWsKdWSI5N8CenPdLTENRXXBCHnVYppYYDQve+PxX2Q7RqfhSQOAB5jkA30PhH6NchV
gd5v28PN0pW+V3eTkirNBeljBgIsxvPz8OvX+nqDMCzN+guJcKngeKzrzy04USCUe1YIacxwVr5l
CAPGu/LDjd7SKpm2/LFwg9rfU926WJgmbR+WJfSh2V+P/sCH++lDy/kqx6HuUXXf+IihULeXBKCz
CQwq2FKF9GYgKovIqsPB8eclQIrBRSWL/gokVC7QqGFOX79yHba3s9Y61zzFofIlC53yNcaNnbTM
YOerPqvg6Zf01JXiaY1VrqbdiRFUrdXR1fnYCQpzRG3YHaE31AHX8WYUgzIC8/H0/9o0jUzBLhXz
e3oucA0z0O4i4L0RcnztBGdUlvhhcmSi+kDgNjSjWEYoOrY2PdYHVuSxwI3mJ34adJqVQOLRbIJO
JBh8yvRC/fKgvZ4Y7OZAU4ogtiYOd5X4z5cOmTg5diPNFwAHxf5oXRjATA4PXdJh5cJRA4VAt+Cr
xYCiy4gBxKua7cX4huhWmGrNaINN8DWonmn2BJMgUvIvg5BSAtb8DROThCPiKCweDVWuQLOq4hSi
W9+EpIUndbDY+sCdPPINlx5ZjYQBHkyVibybP+QqMrZB8ptawoqbq7vKobyCD5x9hwdOwomfmLLf
RCmQB7kZNHRd2CE8aXMjBiSru+Ch3vwFwJEQyZdWrFDF2TuAFYr0tmuOzVAFUj5VolP7mDXJTkQb
f2DyoCIcR2ISQzDUaeh3LiTFbcoXhg0Pz02jBKflJXuURCfMX+7B3baiVwsdbWT04AybSnZKI2FO
nqpzUmhU8eAnFoRLcMRClqRY5f1mZ1oUbkWsouReO9iYztQROYChs68MsVzHvOQPlPV9+LnQNZ+H
VSb2MC+jwCfQHvuvwsrtpUUI39XpUd+/Ewi+hUnVxHHT8taDy3XXEOgNJTK4LN3FqqNrZkLBjIjF
elAoYXefWFDL4yT4D6SY1Kn7FAalhoZSHb0cPp0vjSzXnh8PYm2gHhB/KJDg6FQDb/HV5YN/93en
TIUS0LPGewDNwO10rbN7sp+r9FpvlP7mWbRIBrRCWD68Z9s3Gs/YbzUfOYTSCAmRNB5ME8E+PnqR
hZVUhTi7JyQ/7k7DgzfiDRC1wVMcoLvDANruvFhPLR4Rft1rei3+JAfx0xmju21yGZWGhp+X8TNY
2VDLmcUhHejkMcPWPwosEr8DX4McWhGxC1qfZPpe2JJ0+Q+5KbqWj+BvbJnojqIFkhw/s84s4ARE
xiHVPN5Kv/Jg9veZ8l5TeOtqBiCOmdzwQ4SuSWllnPQpp/Pb2S1Gfyss3njZHbgAONVO0Pgng4m6
b2ns20xr56JEN0Mvig7KoSFZT2yAHrd5uLVmZooy1CsZp9cuWe2XBK6M073fQcmjiJfaJbBP+1UQ
pmgKRbhQNk1kPEXTzqk3NwGJwFV0xfDeJnP/Wgfeqoc/a9Ur5H/DI+ee/hNQlxuriVr4t7rqfm2B
L+yKpjEwXbjDf66qa92KuNxJoOmAlA5zaKwW8P01D0kBhhGz+oL8KF/mtwDLu3qgUduQ467ePoAB
fTIGvgA2z8pzECyBqqKkfH/a2W/8rWjLpG+/jYvrX41DDpqjOjBBlJ0gBzvh6tUXBDgGoM2tT2ak
BMTtXYGQoi89RYB09iow4g+it317sMByI2IpDTCV/eFrfNCMrK4jfneukDzRTZ9qyJVwtZfAXPT+
n23TVHIMVJWKuS3OXRSLQeZCcUac2e+6KWz8dPSKFbw1qv4L0PmSircjwa/tELNpZYtTnr3G8tKL
1vRefKDpr9pbuxgWFXb6D3dRZAf85vrdK+5JrHVmX3zwjwQ3j8YyuWsYIdwXhKd/cJNVx9KRWKv/
o+DYrwQZF5w7XIULUzhlXRmf1hPSyp0Dj8zIjxsYLvh8HhX1ZHANZO1KAYOf3cjZEU77iRsWV3oE
9jjW6nRA5pBoZ0go9eRktkrFlJ9G3nmu5R+A3b9oTUcbjfKxGY2R5XYJKnAWA3ODo6fOE9PoBMfQ
e1oSN7ec243k+WZdcjsstoaL/nsbrcm3l/IWFmw1dnlkK+kEQwRRGn0WNxPaogIhaLnr7EQfyYlP
XetutqiZgnA2/EpC3zHklHjLjauSlAH8Ot7U2LYlt8YyCwPyw0pQNf54zLg7UK4BJVHAbpwApH79
VTHIz7+7XupxLxSPk5/81bFcza46pNg9ftnw3ENg8MfHH8WfTM0sA8d5vDMGWhC11MevAuPbY8ps
z86eO1P91L6Pw3AltpAU4m+ZPh9zhyZelmVbN5KmomJ+otbVqzVarjZ3Ht1DUGt6r8Jho3/w8vAH
wyjkiahjvVba8oxVUuVEN5wbvnn57nBIdkX0aAh4treV6pLTr39G5YwxE5vrluJAwTC28bVGKOrp
dul0xjyqOLChCSbl8D+ewDLHQFxEV03nPDehlEz2DmSGFzTX6kGtoM6wg/DH5SZf1rnzEqpnt/fJ
97gb3X5fpXTpfKK+LsUtzHCCgKgkCJO4QZnqfzeil6fJQ51En8EMwWc/qNtDSOo6JjzAq/XVfPFl
25KcZ0btC7fKJV34YK70Fl5hg8JIIrwpRPpad9do8pZJoE8S7irNgyplYtt9iHH3/yyG3AvhYXXT
gd9+ha4Ge/wOYuXbOv8dhKkeh9i0I2c8IsqXl18g31g1tkynFSX7/2zY+fyB2x0wzRvi9mH6iel7
zN9Li/n2Y4LKf1CHrnHFlLlATYw5Z4jaf29q/MRv5n/JaGaEbOZUNbFu3bkcBiRvaYi02vszdgl+
jpRKj5LYbc01GfZuBCu8xWdYHRQmBc/Px6Pc9LbkrUw5zMa3WenModBwrqn5DX+1mwottp13ht9k
ENt0X3XbZWckISaUVpn3RqWZsZA9RhtmytZcDc0wCnr5n0bMJx05oOO3bsX2B6q+2vmG1gxiTluF
i8VcyJV1aV2kDrR0iLhxPASPNucz4u8xDeAQCo/U9GbE2vLn3m+v/Y45DHTWH7+5QIdCEJtzlLZ4
sgfrJN7mDKvj0WQpFkra9KRducUwCEeOpraMQuvDz59gJ+euMibViBR4CGl01v4ZiIoawGSxM628
E64nwDwc/SdrF360ntMltzv2UtyYXnaUbWAYPxEfb252yczwoCAsNWBiOWM0hiW5uLgBXQETGIBe
B3hOzsOYxSD6BRawsA87C9i2L7PEglUstGcv99rchCo/1QH0OB+7qWF2pAH9vE3M45ntdnnOE8PS
APlUOGeVjBz/BvNcLx+WHw+lyjlM0Y0Qbz4imnxZ565rQ5tEYV7Vn8cAqSWbGdcDvoKgEwOdxeuh
KUu6RWYmDu4hVBP2vAMoK9507myaUpN0nWHh5UqT1a8xeSJrKHqvu9UacrMm8utsOr1GrFMA/z9g
ZOBkqufjHfQ7/Jg5qAr4oD2Vj7LY8c1wVn0bGDgF6xEPLe7bUIKLeaRiN2BG69jcOKawM7ji98rk
PItK9eZEWEZ0z7CN0mKIjgh+dE0w4dLds66zXCg53Jj/agz8x9I2UZUOuKTX2EKhqgDND9X00V+A
/I82mJAaf6cDDb8qLYHIVr0D5SptWyv7GT57EZSqNn6brZklPblvf6Sc5cX1AWMFreASz8Y6ahyi
PmCV0hQyXdbyU3jZeG8lgYbmigJz8V0rBkxDhYH1kDc5zBqn4aJ3PTAH1GWq3xkNET9W4w4qOSU7
Sc/l+6QBEVpHEm4MKEL/gbkx0Xefh18yGjwB4xQD/Gev/ay4vx2aCworSAo6Tmotbwsiz2ceTMvm
B0UVMtzIPYJlJHY7fl0sJXovuIGSDHdECPg+eG53xM/fNDtfa+dn5zEssemLxmQBFPposIcZtJck
0eirUPs9aAkSYp7VOvmQ+ilK+adVwIb8OQmo8IMotF8a3yJNDHBkw2MNwkWptBpPG/mYnq8U+59t
1mgZSDAYJHYNal6Brs3zBCJFpnakrLuZZ+8jCOlWoEDY38AHrcRcvCY6l11vVL+X3Dc7yXF/Vnzu
aq843UyNE7NCQTlp+UJooZiGbgj4fQ3oTWvG2Ab9YGv0nPiAydmWzTCqtsptt5BfycahvjziK1Yg
V/vS4qtpWXTP5w+lmY2Q8IRRk3aEst22w/6UsX0m+kR001MzQ9llaktgWcjb2rUqS+XjD+VwjPy1
+xxZ94U51m4zdMT9v152d2wXhJCdNzntROcHLuQ2KO+CArcpZkpaWiaQtyIGpFNr6PxRJNgZXMqH
H2oXLE1yfEUbDU32a6UibugVkjJ4Vmdoqxtns30N0s4fwxb0IdHC9OyLXuEuCKXztnRRPZd0sA7A
sZPmeQ5suyJEXo4yYqGLhhugsLV8F4AS2Pta1H9HBxboW6OEsRsujs8yAJCX3M7O7lvgFIosZdsj
yhIzx/TjuLhrhWIdw1oG9HG5wqJ8OG3VSFN7U9mletdtxLItZllh1o6Gt9MzRaYGZl/rh1+Qp9mL
94sSTaOXeSQAmpJZ2CWjbxvfDoIAQmAYcUSqafHBqu0EmGZEUz/Vye3sQ9jCBprcOXxofSrc4c0x
rMGsEP0mrB8bLz99lzrRUm0OP/EvCeueQHPVY4VFu3GkPyqjk8tHta4dpHJ37SGvCp9Wdj0ovUc/
l8RrZeKGRj1FNp6ZdCx0E/jbDumw+Wg260ubaF8mvdmRwTR57mHnew9kRJNSss42KGtgsyrylWUE
cu16sEul3GA8JBAD39fkEqXP5E7u1S/CIAwpvMMJ+Fbg7vd8YkjnJI93AxvQV4HSiMTH4NlM6uM5
IbCSypRyCwk4XvkJTnx2HJZ595Lnc0qGbUQSoSMd2UVlVDA7L5qDGvDPcfYALZflgPflZSjB8wNN
Gm6cRQZ8ocL3LYFzM7ZryVq2M9/0xxxOwcGso82m2ROePg6FBPHfrEkLY5DEWWNXQScez79404FJ
ilqfnWMONJQBI4e/SD008iJIAmN++S//9Tz+/qRxLvyo8+x8SzlDjRu0aML1o0WfyIKWOwTcb+NA
c2rqj33QIvDdYLiO2irygwNK2tA4sMSOI9HlRt/3MmloGDh21VIl/qGWaUydLmypr4/P+V+OC/Q+
YPael2pIyjGAFTxb1HR4QW0zvLZHinZfe31Abc4WQw89HD5goM+di8lGWFE4fSqQFGLtGMkP2oOT
tYmmGojiGqahhFkKAqkYB8xuNURH1ubkpr47YixhukXf1+qRSza23TfYAyjCqHQNcuGiCtPXAZCa
jqGY6QfXsUm+XJeSwrALBz4ui/DAU/sc3MVB3CfoHo590kQEgLBilHJa1GS38ssgKxs7OhlCLuES
QF5/3FSfWm4t7bWKYHj6QACpGGYUby1InPBbU1pIREM1yNJdryJGBcUk8a+Gm5BrG+vazQZNcI9D
rC96IGGop73c1U4B+l/W8qYQsB/RnraMaQYzIPPNYCEaWCA5BIpgm+1FxJrMRuKsm1YafVgAHhUy
6Wmp+Bm4OrcvdHW4maLdwmqTo5Ix2UVruEnzB/XxikElyHAcyv8jHz4910UHfLZiGt1tsIPszon5
U7fiSNhrU0/Sj3us7xmcjr707kNpZpq4IWNvqXcQhJmRysrBtG2GK+nYEgNeeXDOs+y3O467jLeS
DUeAJVEfrJGb3bcGEkjPQHVVvN0Cae3V+5fJyltmOcCvC4X6ItkZg+1GBVBpSjejkXNhDz7mzRV7
w2B4/8pl2CysarpDnVpUWVnxcus0RHjm2pngm2+XGAp/qe3PjF202Nbx9cU1c5hdcaxqtucQvpXJ
aILLLk2Ve0mI2vAz72njWQOo0axMVEtTFO3TgDJAaNwdr9yYTC9Y3+47cOMYMmO/3H/Fpe68E0ax
Z36HxxRfqEb7XADtXAKHmdeiEguKmHbCa+XzHcPO918DlLjznAuFQqIa5MuCjBNH00FpRoAZA6g1
Cp/k8pwSMqBAGdmJKwMGsDM1uzEfXtyCVF6TLTFzu1UKkHbHBNPmkjmvjdUQAWs1jDfDvbBU2QQD
Fq6QkdGpW04a+T67ehWzRGBFr1kcJOxFicE7nqD3Snx3MN/aqKHva7Y2KOh618U2Q7b5QjIEGFuW
KKOcSsiQDqpZHd+s+OzxK1rTeC9DjlJMZDC8PYX0kJQL4YZvmY8blHC/qmjnOmOtyPWe6yUiXJrl
PLsq8DvnL1n1gq8EIIJcHS91lQV67BfhnMl6fNsxPSW19l0ueqqRDJwE+7fvwivgqO2gQ7x3Shur
mWKMJDHbLXCUKh/ldH2Jcezp21nGXnz8oZZbVAC6wLAw0pnIAxkN7bKzn0ZirEkyXPKa+khuwo2I
cL6OePOMDJ9PM2+VHHUU0viPU/ChKNj1J4i9sDLG6sw3YfNYjrWWk5u+Sa8O8Jh0znHygNXTbae8
KIfZ0lNnhiCYIJ3iTWW2zs7j5rNGbSWknXaPB5X7j4fBcguT/+FvKEqYgdjNtQz3+0fO7Bcfcm7b
Xa3OiJU3IrOw1WM+R19wcfp941Lurywin4a7T+wcVWCfmMgcN2SeRsn5klKR3fEvUzgxBdN7Pybo
8NspxL+E2D7m56DeNtOGm36QP/Onf6szAHxwOrEGPQWTX32mZxknx1V3b7KfjRaPrSBHp1FkVhF9
dHghzAqMI1EVk8Q9EWGo3eB/f1jMdvQ2PS1TLxjZLoipHjtJI/laItXxCRUmIQCuRAoH1oDjpeM/
jzApwyvg3DIeTVnCW0y4rwypqShQsIP4vxV3bco3CRWrkNBX0IPAAWo4uLWxobr2q67h0/7xE6jl
RaLDyadJ3edJuuAzmnL8r2IPYBNSF3I/6auM1PdcddARt8G1gf1u9s0fKdIrBIHFZfvvfPcbSap3
LMSGzUnTlb6yc5BWRV+Cv7x+F4qNUeaQ7mgB4Whwh3qqNHUEuKKOsNQwS1YXcmMBSc4OaV2uEjbV
9u1GpkpqiE+zamHrcT4rkZUTc02Eumxb9y9JgqibYOCS4hy7Tp6X0FJarZbdzNeV2w949ydDoY8T
6GuaYfNMCOneoRw30BXRKd6zaXW4C5WGaxCqrGyIjjpa4E2AGknbiil8vK15vkQCk4ciP9yxECgx
sqoezN123o7M/TqV8mWWwMjw/rtXm29f26JhubNceqolrT3c/OLdDmCpo5M66RZ4p5vC9/uKdoYk
z2Fk/uBqPWJbeTcj1Jdezi5PPVGLYYmYcrUqD3YjOG8NYOuP7rq09pcGDD3eTCqMFkeEagu8TJje
AXLpIqxiPU2UlPm/CeVmtMXY/nvkQP5jphBZgyFakM6QQADZw9pFT8VJMeWOnEA5AaVsmd7l7F07
sbKKwS301cckPF0qFz7lvZFOhnFz+oEBcM0iWk/Ypej0BijpE0hjpHoLIldHvklmh3DcqfChFE3Y
x522imwV/DSg6wBpfUBbQ7MiSwMaduw106/9a+paMgrKStRe/Q6A0pse3klwiUjLXsf8yWdhn14T
H5MjePfSD3HH7GYUqFGkLvwpWV31CAyMgO0w801aLbrVIcaJJeoXWITMvE4X+AvdgbvQOuSgw6H7
pokPZpqtCFWhoPBH8BFryokLgyQGg9bhAy0dsz7mEVTMeXOBd0korg3KTOresjB+Dw2C5NDL3F7F
OsjmFDrdWUC/1GqdJ37kyI9RO5CR3WJKByVIphTFTDvpJ212+OjDtAb6INcwSOy+WULKLJmxpo3P
Tx07S68UsdwrI+EvloPPkqvW2FaG35vbdRvf687OCfksZRR+8OFqaNUuVcWiwdCzD6z79bEYsMQ0
ZhIoXMX1ihKMLat3q3/c5Qd/w1BHCGBKz1pARIMFJhvcses3wO+jj6VFfs1cKH2FmAxjNt49kWSI
7tEzIuJubS6ijjNzIwmB2JXNPZlWgZacFrebJG19tKDeEq8CMiHOXy53Cf+OjdEsqAG8ljW/ulzB
CldiXkkLaq1tnmyrUMZ7dKyXLsBMVlevtQXVl1yYK+cU8TR51HU/6urd1ExHrk44ALaWs0pVtNX7
S1sGb1mZjdHl340Df2ACVgYEPU5wNC53Z/L86lneZ17n4ddQ42UZguB3hDL/BAwVBSJWWszFMRC+
0WKHgvLBB9hcrNXMxdmd+9xvKb0PpgCItdFDpM0ry1IgkLI6KbgYrcICDn6J6ucCSqMIaRlIhiFU
Wm4GNm4caI6Mn8EMVuHyPfc6WgYsGNl3IeeDUlrMd3n8fBN2ZLfsmeEqCkd2YRb7HXELS3Urs0a6
fexsQDpkfrZm3IEXj5TIlDgPscN0jG04HHKTEhAX/tZW9vFJFzyMswRdM7hRbHFQ1IiTRtC0hx+W
QbvJPpc+RxTh8qo0G2ui7Sh3jU7h4BVo0ioW7LOiUtIvR1X6M1GTwtfAHL5PpgCK28aDDqh5a4ON
kqCtbp7Yh/RUAVaU0AjOX1WIi1MV82/QIWirJ8rQcGBEqVIxb8BkKpUKicK8hNVKVffedYJQaAkw
23WcYWIpFYZapdol6rllLbAG13nWaTL8QYDj+M94Z5Dl38SQsc2vyay+WK+kH+VsnHzd9NxALcG6
DbSEyGcPxNdoeDW0NDasZZqhhLz0C6MFwb4bUVkX3FZIfYxcLx6AjVlcTs4tYaA7QLRhsttr1qLO
1S06aj20N+PMbRH1Rgt9okDyEe8JLQDEnve1pvXAYBDKA+l4hlu/6bSJr5OO3mewK11fn2yd3Azg
oTbsOE7PPXR1rOHv/7Q0h+yNS2Mm0KLTbs/Xm84F3TmW2TNwiu/pQ5Jn/LUKeVoQozsOKCF6vU1J
xd1pqM+GSttobDckZUCviKWcv1R2k4nrmYwQqtI1g9JdgorL7TZrAJuBtFYd8JHtIeIO6UgePPzH
NYU0zw316UatPxvr2mn8tLbNuWFQ9n6dT+1ByE5tPm/EUA9vTEIZ4qAhv1N2PDHgjhvSli1X7iu3
0nA2Xlc81NJLy/UE7zn0vX0gSIIJpjknjVHwHxWbMj3iE/biizG+vs+FZ4TRhRg1lHPBzZ9p7Rgy
DpWEt8hSAN4SKyLxkcVEIz0OHn4fDpvEs07uxgF4FDA7wWcLUAp16GOepb0kjNfEAg66G54UkNIU
hgYkTKf4qtBB/3X1bVQehu+vOw6Ww1GbxPq1V7KvEkrZwyq1ofe/8Ak5XDQ69q6MJrPg6Jtpn6oT
ZIhF+4dsXOuwuGG8nqKa32M/XjcdyS3JspIup3OuuBmKhhN4pV2Pav7X6ibvfWa3jZXPQVGO+79o
3ztv5g67OGucjLCPZGh5bIxFWZIlGq4ZWmHSwqBx4gUuUqg6p365WjPRM6p/+4sFmDKWSd1nXcfW
NYD5DHwBVALAojqBBcqc8exxDaipGNInt3CK2uL+kAZ1jop1kw0RzZ2snDFzxG5Y3Ts+d7UXrXKw
rE1rI2sGz2tvZBhk3RwDMrirgLElQgvPRaq0D9hhyNhyFtPPDgyClSMamGFWk/G+CYIwJdVSbHac
SQ7xGbKIWoWx0twP1Ou+0Q8fRSdrCUvq+HtI0plj1JsDwtAd293w8kZJ9BCr9Dl6cu7RKkDmLgS4
sbWQY9VNCmqM3wm/GV38UGzpWXUNfFsIA2ScHqswkJL0RXNpGUOQM7eslth7cNq/CKfr99r9mvLc
ErmR+PwPcM6ZCGHche8hHUBZoX5Nt/xNx6tOEbObdX95R1Iw/mMDcd3TiH3o+DoeTCMsIQJRp9te
c5vblw+7AGh6zlh4lZRIaTu1JVtYhHkmXsH5S9/13IT83Kq5eGrMypOPxnEGC+AVwBIRDYyvXLo/
Sn4WavZeNHvgRo9E+wapUXjGiezbSmi5yH9MaWwToibxeRVtD9Ji6ODY2DhoziGwUfCMDNh4bThF
u5fwODu1eX5E9Cqa6zZUkIaaa4G4FumxYw9SBQpTIU2DPmRL+I4dZPivAkRYBXKyhP4y4lRkslwu
6L3Km9ZmUPmx2i5lNYcAhPmvsARpmVsAtxXy2Ru7EBC+6kLaLoXOl3WgztN8fTYH4tA0j1AJsxGJ
KbxL95Jnca0XoERDXc9adKeMLTGH/P30Zvu6Bi3WLq8eKGupg0ma2rEn3INfDBWfUJHIP9GnpKKW
pFzLKtQRcIvLAAnSViPraTlqXGuzCcLoPfeKJugepIadsRVWU5pdiAZqlxqGq0Y/VXYstBa66AQ5
jisuFORG2gm0vnpJaCKJQkFga0m02bdxgLFSKuXrFuehoIXGJuxRNvqNYUcys0gjKLCVnGCHpktI
ooMDfMHeHlhrk/e4HjbUVWJde0DjsVNbnrOakoT6K1fPtlLavNFKclSeKPA/z1XcVyetb9P/I8O1
u1fYtjoDV0shoFhpNOcEaW9TZnTQAiJQ+Iq24GmwAhk30E8yg0F+CUr4HoQWFB06Y7J95Id6SuF9
nhmU4ABbo35JfZF/mTRCFR7Ui05f3jplpLV4+4wBkN/baZlA4JAu+9GLfQJLVBNzbZq7cDjQuCT3
uXkvn6k+u+H+mrZw3n7sOvjqv67TznKbjrJWwBduFS9rhRLr2eP0cVjxhB/7hQmj5/7JtiOByBT6
+znTFL1pb1r+xbXnAbFunp9Fk3alAnrtEEzaBmrwcejXiulPbLm814qs52S4e27ZhnysxkgqLgDm
h2WhOF9di6ZPrTa0rYAIbkpVsbmrc7bYxZJFnqif+o2Vi+yYlBuB+AO6ghJGJ0fMB5xV0AUL7Dwt
Bdk6J6KVf9jearXENU2aNHEEwNW0MB2+FVtJkAdD/M8l4m4slZGeF341+dKq3NIhSPUqbw3b/ZSo
CP3vRM0M2ObaaELm13qfKuJxqr6RBfAhXmxAAGXa3px8KP5rmmPJ7RsGXmqYmMisafXZeH1nMkVB
tkp2HzhwodAdkPMKSa0bP/WPFUncbOthXOW4lusLLIlziuPRQAsq/UiayEQCX2HYfA0VeYOXjhWC
JAhzmsz0w9wAcmzVHzgX5vLPKwaZVUyWryqY7MP07ONLLhKQT0uOGTDzYsLvlG1zmq0TuS48qqhf
hP3Ck+yvynfX799aOpD+0kPh0eAPBQZRT1PdDzRLquy3dYR57gnTLi8BLTd0CwU00/i42V7389Qq
RlK8oRNIvBDICBqfhr6bjsLWUjXZ1gZCIu5Hejjo6/7DKJlVstSFLlCpb3UExt6UHxFTH8B8TwZO
zQ/Gqu21TBuhFBzSpmcAmRs93eXOxY1gJ9rkE5b/HMj0xxd0xy+vgJUGtq4yMC/Zbf1ePzSSo9KS
rtz1Wrgdg+q/7JCKwMIh9Gj7yRtvApqU1V4rkdlcaUykooKeXLjzPjpTIVXHQnb2AEcljj35oo7G
TrKmbHxK+DKqDH53xkXVdZboWu+QvgPXXQrOVK5JSDb5nOytbzAzTrdFWv+tjuTsfY50Sn6abvn0
pBq43kyMnQy/f2TlDvjGo2Se/e4G8W4KKJmKdW50W7redlMkmrrq9SRdHVxs3fPubWCwABUkn87Q
CpSXjGXbe153PV8PMxyINEAyssO4+ynZ/UFS2F21l3IAiEZk9s579mJYGJKG31msMudIo2ljd9Ru
wPDWWlLC+HnqLd0BQlC6HHivfuQ29RJw0BtY/RwO3CE0cuL00BAnI7z6lzl2Afzb/lVH6EP55VYL
tesSu4RpYMJdw+jCP1XHK+FQZylGLUrUMiwWCZmPuxVRdMHlAVv1DOW0H6XUNpFfNuTTWf7SC40b
SEvxLeAdskPFzd+Yd15FlmPo8OJ2lE+8w8tdVl+SHTkG5xooeYKoDjcMnfQyL+HjHbqafsazmCMX
JnrhfFI56E0Gvi2wiAcb1Op5K0pL4DgHGdsO9JCwP8QhNqWR4rY2V0Z0J5IxYT935+nah5n2bYq5
3gOUvLxUyBkJD9RVraw1OXqh/me8lqzb1GFcNK8XP+x4ScQAJxjEVHYvaip955YiqJLNwk2wnryq
s1rqPUYqxMLzD6GaarDM8gQ3wn/KIg1hlkBBhw2oauctO8J0TX0xFRrUPgT3W2qjU+f8dyH9vjgj
KoXxDizU78eY7ttg+OsC0V0Sd+nOzSgj0RPTgvkFfG3GXr1hUWapQaeHIMXBAUKSEmqlB3TugssL
eVljMLBzhcRIuiZxNExOI/TKABTCc/UZvPf4k/umaj7D0bwJ55wMaomuh1SctT/2/2sC6JSMklr+
/DNu1U/XWdrGCU8SDIrylQDM9Ie4Us13MO106FEFCJLc5eAkX3QkwGYIb0b4Gc4GfCTL6uYZaWF3
ekcpoWGj6+UsQu6mcC0uhUgrwgfzQzVpSvn+rqq/xb1B9ZxIqm9W0l0Akczf62mq4wX58P9cUH6l
eqONiRuDgit46RjNO9dkZnGmW4vr1tzfeIIyR/JK75aKRFViXlwi1gs2Hss5mnavpW/IBrbwxSVt
rY3zIR/5lytNlzxOtXY5uEMwrrbEoavTpHGpbjT3baCWrnjVbVoQfK9PS/EiBmiofTYLe3GwuN85
wVKkMoMo07dnPGIm1VVHR/3EMWt2RCDMwWFJVIZigJDOB02g92AcrkT8KTV9IdFup94dGj9Yd8YP
xIuM08fT+JEstfOjmKty8LrJBO+g1/67t5RRP5CEnAGaCy7QaeS5hz49Cfm4/8M9Mp6K6p4k0f0t
iuaILSK3TM1ilaKOK1lKuLz3hZJzTrmTmcgZG1gNR96OYkszm+z/2M8XEvY/Snf46d3hkWGyqtyF
ulwfDXqFvJjqu8lvGQjOE37E5onxxnVHRYKgHqFtcek7Vka1cMeCABqkFk85N5rcTmjoWxwSBSGJ
4oR4kW1rdAwcIcmW8vmCnxUtsa8Gj85m9zvAjiyhZpsnf0pFN3pIRplQX85tfVBJqr6QnoPyAmDK
moEEH3zD8KHkmYdMcX+08iAhAtjGXVCAAYLSB9zj2o7xxc711CCd2+55tYg3/ZxSgl2RzfZLol46
A9W/fP6VzQ2r2hCAdpL9J0sFSroUpKoldjwa/UqHnQmqAXXjo3xr89fNIW4gwGp7G9As9kipj0e2
oEiRljcjaVeyvdaL16akHzTfcav37N03Ahr42wH0mQ+m9PkZjLRri9fgvrVnPR+qPE+UcvK7QCAP
EeH7DhigMnsth6fELSWHMaLPLqZIY79krNbxqnDvNj9VXxEXw5FBR0Qz1UbL5lKY7eQgWHu/BWyr
jGQcGFcnW2S3k1iKTWU1siMT77VIvFB1IPzd84/CD36ii1Xk7ANSv9KN7mxh9v/TcHNcCsnmiKZ4
Zxi0l4yBPzKc+ZQ7T6ZIhsGgrYswAqYvTGyFNnfxnDI4R6DwvYddbbmMfNlQK2oYjlpxX3se4ZiU
O924mtGPgSzKqtXdorIOLAJHPibpZwRc1z7WXvbJfYlRuTTi0u7sW+OQ6OwVk+J8bPwZkIffFs7g
JXBMJcomoYDEaFIagcIKGUc4yKFOgXM2sWfdBUnZMVPDFErpgJB6LjttTt7Uu+iADOJoZVYWCR+H
unBsJRokcwpE5mz8K9exYTVW2+2Zd+eMuSQUBuKASgjVdhjDXs367Xk+VAYPxmfmsCJZkzh6JLOj
pAXX0jS0pDrueGYNw/yPw5qtODCC6ZUqiTQ7H4yJrZRwcf3enKJovTvYdnkAivcApGm5BARb1B0s
BHKoyuLVDEGFMfKS8u+L0kEx3gUAM1Evma+norF+9bRUzAcgVvLBryuZ/I6TMNh1QsKAsApHsnjh
B2VepCcHe0JNdndZWwj3U5PuovoZaCr4s3DmLHtGLzO5P6rojRhgjF8Phiaw+30VUw479U4vAOgn
79B6I7ubX653rUTK3gA8gxMyWQ6E+oYSRcMsy9QEliVS6XZCImb2MfGlX5qmQDHPNbcxWFRsxBc+
LB7aS5slIlATHS5c0+iMNBuWXQGNvZziM3DJR+PKTfLEc3Q9TUw84OHTRrdijbJfayQoqb2paQzZ
brQpywE2ESAj/oGjQRIb3d9yntcOw9o6IYrUMYKltjSI0tCzsD4hqz+ZxU7QrXdz5jD2d86a7oeP
SyjjOdemaMqXQv2naHJHHmcdErdxBoBrr2LXJft+CPk4BJSia5RZePxoyRcs6WRmJ37S92OoFK8E
2qr/eyuhcPeN250yn0uIxlsqMZl6KGGR5C4N8rjF/8P3wpiSwL71QpyR2Btpz9iSO9vhmk4OLUfV
oiaFRDS1Y+2fpXOzRU0CroeYA3HNlu53fp5QEdeKg/J3fDy7QuFpSvOMsTOg2oVeGFqfFmv5Bv7h
tnaIwijYc5UF0+LBQYZEjj4Nlbvawn+gSDvOzw3YadsiVuyTX3TlH8UuOM+ddVYZjEFgPbc4bD9O
OuKAYn2K9bNnoEzIKTFHcq1EYO551ACiv167fW71z8Bpry/5+YhCCFD1rsdhQpq7L28jcw4G/Pfn
XXyBcvPF+2ek/QV6waTrRUM8rvxs1Sx+EipD8xBYYR1kVM+qCjxYeL+f4A0fysMzGBk9+IiSYes8
QFA5GPhVTtcduUez45AGXtH19zPxNiAGBrtfdrXBoZxO1Cza30Wa7lWcdS9g/wgdZ9Ehn81yxN47
g5pGcT3A1N/zq81kLl84p32A6DQ8Lls48zLaU4ZjjC41mOhhJnHMC+qbECDaopl2DXUiSNlBmlQE
bCQ+ES1jrd+2SSmgLm7/+nckGXk64n11HmJ9wTADGSzcITW0rdwq9clYRvDUZmS+WQchn8+h2cei
G7QzfQZxx+2GwwHwhBnY2BJh2wsMEh2afBdzUStrOOacWyYBcyIfzm5CUsY2eQEEKrN0AH3hUPnI
Y56Ku0+E/4X0CK2gbT/+IbICG6yWOPzAsrw32vGlWnUVUmSTVma/tZs8v5MTMbS5Zf28nEijDaWw
50B+DKE77G5SbN/00hSLeDHiGFG0RA2Pr4sYtL3+UBX2uGQ7fclsUQS6M1IWyWol49yLe6CpgihN
l1oTYc5tL7s/e2CFH5OrD94xVn5rI2SJUcT37bA1Mw6cKPzbKAAmdpgOrr5a33hwhlBQW2zzyMPS
yo+dA2vquchosk4Ra35fVQ0yM5uXSoJukd13Ci53q58QgfCQ9GT6auCZaBn9JMgBuobsAJKnqCfl
aF/Oy7bgjZCpDVtrxcEdsgCPzDu2JJF2l3UcqR1wtvnjGrHLE6D6aVa3cn4QsKf7vFDuyrvbvrTi
RwfHGJsmdKMnW3Zod8CexIfqK+rQPgWZNKkDZev+Qd0ANdbZFm1b3wVI6uLE18HQ8eOCX3ZAv26I
BCUX6EXZ8tkfHx5r7+aBV+kFdVH/f3/Ns8Jf+8tdzduZQfpWY9wXH/Rd0jgpCf2fenheUY+PDEDf
IG1U/CqDSwBi1htACk+nRsRRgSRj4AsSPrhCCelIKNEj5z96LgJlx07RUL/KBWLJOOQXIfUiC83G
Iqwky69bItNMV1mAOSqX1g9P9KoJN0Vzofn6NR3v3KTToa8SDw1u03sJ7bTG8Qq31szpEa/lwl6v
5idb4tEALonzJCISGZjGhXX7l3d38zeD0uHYIrj3dfUtTUH1IaByDku68z0iVFnynRP75UontfH9
aP+pnzMaZJBRG/+TvvrxR2gz3WMeBQxlKZkY7LRgfEyPuo8Ufr/rmLewJb1xqsUSV36E+ZcSlE+F
ZbcTK1eHiKXvuGIvHWcUAkUOs5rLRtoLfRJ/yNQf8DZW4bnqQ7n+C4HgiEJ30AXX1F3vPc69F4rE
K5ZmY6g/sPcUJZbgPxCYMN9KS0U9NkP0JDqbRVOXTPcmvZefgQQqooJLbfrAUQvaEomoWCw6qpVk
2boK1dqIzLr8uRFblN3jzmYeZnzYfLuuYAhwkGKUhdWtVFfAR63UjymgjaHbA06aBqVVpPqrlUon
5weGZ5Ss9Cy0072BfDgU8j/oQePAc68qYN6lCai3fYKH+Xqgo1vQVa6nMjOkhp3j6Ryc+6B7z83H
TZ24/0RjepbRDOlsYHroenzUdg5sebdZRkQrS8KH+xXJKmqJmCjb5JT3cMkfOInTLO3186QnVZ0p
IT8YLR+zDEVFGgc0TFzVvVHoPNi0gMQLrvbVIlqQe+wds11UogktyOKY7oBi+VC6EzRCz2u3h2R5
3GUg05vrTykiL7eKPZVanuSzMDVnCs3M/Z1Ti+Yj5IHESvyRyiqvSwZT+skLdr93ayIh4GknvaPp
lkNGKJqz69YNQ6lom+3HW+DBFA3GBtow1Z6N5hDICnAg1f3cyR6k2ecSYiNzBtOlmMk6jn3oOoxe
rFB3zw5bDorwLLgWPWmBv1TzatxTrOYjIhzcg4dkLn4X8RlhXswERVEEcadpsoJ1CX8nrWraUVR5
F0i7x4M2FtwCzyBnjaq75HfiJBvsBAsnKZ/v5q58GBMqT/TqW+Nczr55zsZDQb47BM1PhTOJWX3W
ofng6bVx3o0oRON3kKPaxYS/HhULFNlQt8n5mCAF8VhzwYtcl/wTs/kIdk+1qoMPGN0oo0grj4aa
NZTz2rY0Jm/JLSxNSuTNiLfpHdb0lIcqDEmIpBwy2ZVg153L5Qjr3u8CDut/PuhnXqtc9Yk8YKIo
ngh0ksIUhYdYgKHyoZMPRCps39E5pFXIHsHvHBpEilLTlNxXfESuHhj19shJn10kFGbnvEordqtA
6/hpT7OFdEn8bw/d5L1gn2jcLwwEuozr7HuOf7M49yFnGcdLSc7wGEZ3KXmgBWtj8dHZGzWtJw5/
vt0EH08rMX67vhapv9J/RO2/vbs1vKS9a5azGowyoG0soDufjdArMLfl9G0pUm+h8cMiImXRZbE0
8dpWzfmf3qIXJz9Mkl59otq5x9Jb1xS2jA5FSODJbpM30RE5svT54I0DXieuWAA3e8mEke+9J4rX
lQ0/KK8DDQZq+QtVoAmdrMrGObYHNP04fcWrzZHrXau8H5uDWwieKcfdmuUWuIrDDVKG9SM414Qs
71eOFoi3lRCQPXiqGFq2Y1JbhWnGtatgMZmJfuBVUXnC0qqNtd5SHFJH7q4yhVH1UIv1WHNQwPi1
3eIJ658I/MqAzEswDuw/psMlsv6+Qa5lXL8PO5m7+sEO8mn/SipMehYqCX9Ub2xJhHyVMxhgHjQP
/bxpt0Pr06BM6GCZIJ9XvqWEtNMGOJ2nAYz5holKFUEX76TmD4/xDF9rNw82OcgoyQvTZIwCUycY
K/pTDTMCU1ZHKWGPv00YgcGpm5OjDdd9hhF0r+t0E0ob+USJApBO67NtzHkMHO3pWNpvQlfV9oM5
H37PqX0GzLdNP6nqJGeMpX5n8HYj/x5oBl3qI1jFdapGY9o8Diq9wdIOcMed12mkalo1TYkzFxm5
r/myQyNtFxV9zrmmD869ZABROTN4JpwUpwReb/GN64AZk0/HMzNreOcFRqCUvjTqXN/I2AC9UR/V
juThdheO13ICceM3V++ADE7+laXOxP5oIpkZGEHmmyUpkTZNvAD5jsy3lc2dni6aF0RS45SS1uZ8
vdj7d/pDO2tW2Ry6SW9SvSBLLE18BPM2WBi2e/nrw6R+GlocET/GgnNeuFigtpDAL4fQ2Sbvd6ux
Iv/32x5aVQ2HmPza4RS+8TRoDBdBJcb1rtZpO1uzCvkDgsKqw1+IulVdnqcLGoJ7TdGS/8JYXsRU
pwRghDFqbQBxGKdlLse54boDyWmvsV2DGig9SKsjgPEpIIN+r8xyqyzpsVIRadjR2wRlESd95F23
9o94fRTVm+MZw8pKwMLUibAynemdO4qY1TkeQouYdsVvCkvWgWRUes3pVFmtKyh94dnpekmw++ki
m8R+yhZxIjnzqpxn9+P0MPwzM+pUXWIbopXjDjeoIS2H9m00A4sCfeleXHBxmcUZMKEKXEs7W/RP
++VQXwKbjzXYJqXLcit0JZf7uJKsptBKsiM1k+sJOfpR+ShJrprPx3dmc/QFzuhfCOXeHDpSoGWs
ardKXNYfJmUOtRatA4tU5ofaHzXVj3nTE1iowApUsGpuqz2Y7ZwjCqV+47Qps/Z+JzvS9ADK9/WZ
fsHzz6CjYTGZ4i+QM058CUQl/fn1zwYVj/yIqUCt5h3+aOFNTFrq06IgCXQ9jQRQRg00/eRGp6qd
g7OBl1v3o0IMb8AYtQg5HYPmKAtRxg7cNnqITq+vcdtOkkQO8Kc1+4EMb/5EXHYGSSnKWDB6xeWn
oqSxorWb28n+TMowMoPK4t8BF5d8EOjDmkp5PPyGyArtA6V2JnrqvUvxdgVBQRPfNkn98fkQlOD3
3DVeNebfIFXTTwOs2AqF3rDNYWQhP3Gq5yAPoxju1LT7naBOBSxbWvmq7pXoPAKlNjsu0dz2qkN0
64piJD9rDNvfohZt7y3GszJqdwN1kkKmBCbp95/KOQHg24bMDseI2ERlvA+KZdtVTb5f9o3Et8oa
ObwqDcmd7b0Y//V9TP2HXVdDI4k87HYC7IzTbF0rBrkd0irou9mc+O8AAcdVMURHlm7n69/ZBUOe
09gQIr1jvAckAQGiDPCAjT/Q2bU0lGIMLuzmP/vLjcNLT8ncdJYCiKHgW5TauHOic0x7a5HCTGV8
XW48FUjCVbsWI3fjV0AgE+T7zTEivHG9yLMiFO9RyT0IDQr5A1a+bufhMM68gURVXa1kHMzUJaKm
QvHAdohvmzqv2basS2exEKJsUbrouY7C7ftlSimBpf0t6b4FCt3FT5ZKnJkX++2cvk3KJIjL3y5T
gRtlRt2x3qqlpjPmLureJ0dowurEqttwDE6C8c6TESNk5joIFjqZvDN0CDyTqzfX318hsPeH+OUU
eHwUCxq+RWY3Ju7D6WxhRqadWjDCOjW/6TmNPd8LXfH5PQ24re3W9Fi6ha5e8dxy98ZXUGioVBYq
nQIEM410DYdy2mMjX+6FkCiXL+FbHMZjQpxupQthqjUKaNLy/HLQ0Itw3+uhpFEOjqp5vJDhXK0B
qs0vZ2Lmku2SECKfWEbNVDDHBRQCQliNspHBMZwEVJtFgcQ+vcB031+CNc1kKgaJ/xYVxw+u2tju
US+WQnOSsppr6QRr4pVVITpiIEKMfsU4G9zmeXyxzKHkO0QXOj84NPqulpzdpUukP0YfHur0Ibxq
SKhU3LWsGSqlBrxcZxIDplhCL2MHZp0+CYVDpfABjvJdWbXFTWk6/IaT5Eq5hn0gp1xqcL+CZkdI
fJPKuKs9cTXPqQvxAfL2OsRoH3olB+PgGTWZuFgk28wX42PodZKvlIUGA8WgVs87U53FS5dG4py2
ExJn4HijS4/TgoJ+SiiCv943PT6erBD/fC+hD6l1qd0ssB49gm/zIcAk78/giJPKQ4e8tIO8UfnH
LAXzdv83zD7RgOaKYRPdrZ9cIiwzyKDv7N2COvo4JzRIcJ2SuC62y+o4bNhHv4t0B5FloABvYXI9
uGe0gKr/1sXhX5ua2NGlWl77R1Tr1kPlnpLtRywOL9W8IFpIBPNAzpQU4Ohkw5VJuhE8TC/QjvPy
RbnkMGTRDrGiLlhsWQtsi1Z6Ua/hg+mjh/VxwKvXPxotr9M7VWm/l7tVUSRUMx21wf2SLPy7xLkr
S8VBY0rP3l/ZxF/YR87XAdhXZT26zz51CWZiziDNgJATqBJLXeDOjjaxsA0H+KeblpVjMJEicU6S
JLCnvvpxYicgmPbiS3Pvr1Z5qQevFducIoF5H8dL626HZlsiHqFZjryYH6pwLdoIGu2K3hFWHIfP
JqlbQant7Aq1Z/kBZr6vObM25cpxALsCXO/56prUuVWcK42bj4XJdGwFsOYkhiDZsqPO7ferUr1F
dMqgo3BjfmcsSAZlEaspN2LNlvBMEg+GPZwqnZWal7pcnyWNtWHZMXOu3hEvqWjOJ2p/qXFw+2dO
RAwwXTQvT9MQw7rRtwpKQKehH04S9Tsql4H385Gc7JBaniH0BbUQ9MYTRdCUWpjUuMggr2qh+X6M
vNH/2L33GDie85fXR0fPuboAfdWOIqsTo9a0mluMg4EYoJVT9+yOtfnJAP2wPNtnbo3uiYY2HzE8
6Jq7wd9s+OVchv2PqqbNfEyChYj0iMCawOGchdeDTT2z8TnWtCowdze6CvRR7Ex+UHY7MAQRRJTJ
1rLZ3XjfPDPgEUsKyI8htLJX71E9haC0refl0NwQ1hReLb6Bt/0trsZ3JZi22kdivvmcCoPSZrgV
xhu37XD/kMitMPrF/qs9f/G8o2p0/1rC2jzShIHsGe6XGuECv4u5Vr9KaINUd5XDLVGmTOamrMYz
LN3XNieKzLpaRHkSjVnLIHt2tW7oWzYk/+JCIHNLHyxVhFTa6oLtExPwANhWtCMkzXUAKc6KfQXf
siWxU9nlcvYvAFrzUeiyPCtaUilkBErMcknb9cPbU1MMqheJWFns32QxTIhGOfQQp3l9yJiwpeyZ
emZ0ePefT8TYj6frV1N7THeoiM4FX/jA/sFL2O6lVAbLVat6+1LgqqaG5E4iYKGfRILafSx4Gf2V
0YuNOQrP4DdL2ERxjY/nzLd7n/Q2S7CwEdVk5pEMvRbOTLsB1xIbc/iVpdnUDqjgWrcaa61F1RXI
ReedZ1G2EirHGtDFlrW8NtM1OJRml/RZGGVOwE0x3GDiFKsHM59XQ/VmObmIoPPH7/7QmfiboVbh
XQLWJnX92qJaNu5fIGdnUXqsFzucaxw/rQ6bhgezMKEkNw5RJuHBzARHUWTGOAEE2Pa89o5dnMh9
AD470yshWmawVshJjrlzNVAXCMSTuyt6ZyqN8EWcIkzCoBSTmyJw6RrZ4l5rmE8Ve33xKOLCgBut
eMPuxpe5RuA3mAW1Zc6q+gJEN9RczTe6g6w8Oqe9SpyX2LVKio4f+2dEmWb4Dk6qYwfguyO6ws/6
4KT0TIQ3zmOCd26+1MUk/ZBpmvzaHP3Q9ch6k5fiCFx6HzAArtwTwFH8lE+4drdiQU7lEUb5x9yt
9717fVFCRD0guSGuKiLKjl+ZkZTwl8N33FXsp1Lg/ZMgu2nnnEzzjzLV3tAXvzopEiyKJ+fiJq4H
TvDcq2l16We5k1Z35b3XK77WxvyoKI59pAMp8cMvtjpdyIy+WUnDEeUw6mcrxVw2vyDxJQhh59OD
8EEzmYDzBa287mjwJTy7ino8prItFn3Lm1rJHaTT4RUBoUAfx4TkEnHpjnqSroA3qFmoP4915Rdf
b+NFxexoysNWs/gDpC/F9SKapYGMSCHSiMQPwtQK6vFuMLs2BZ9BjagL1JwxO1YKnnbNaCTrBwRX
9FKSFcdI3cjMF1J57kG0XD8n95VYxdRUigOaxBcNF0/qnC8+qjKwS0MNgMwmZsIiVYDwjhC3QtBf
Q4+VduVEIxlQs7A97cAv1pT683NkMsKRisMVqTy3QjpEO52L8gD2dMg9qC5Tylx9/8SV9sQfB57Q
XBMZiyPAskFF66P3IysPqnwSjB1IgyK1logJnXHU0T4bPKYaDYsbOQddpoSIEgbxGx2fD90qMNJR
YJFgIknUYTjS3k1SBgaebdbkWVtLF4EAEWXXRB9dGBBPaig0jK8NZ8fWDmLcp3k4OdSj7joHr+zA
mKMt11gRbbCvEifDC0KzmNWvU/D0ZH9OGJyF7/HSFT3lFoueC7Dj6MKPMJQS17MR4bfRxHWPDO8y
gxRdIBtjvcqlOJGtUdxSNmQ1QWE8KRMnns0E2d2vQoH884FfWJy77NORQfcDewWkSVtE2orVcf1b
zgBBFNuQcDgHdGrE/ABT5mbgGxnTcPoj4xNGiN+bddV7FqQ/sPzHohHMN5JHtgzbTNBdSplECekd
RDhptWtgKvbZJ8oqUwtU7ddkU6WvOeSSvZga4yOX8lsQ7wA0W1NBDcM7qC/hirQId2hBVIGQFdk+
Rf+Y9ITp35nDKkEkhEM1+trAJdX57e72nw5/qH/8NZXPHnBC7vvpFmJo3Tk0eJDkTRhunAcdLFF7
ffKgk4Wng/Ek9x35XSLtktoW3rsqg2m9uf6jzc8bQtoudLyqWQiM9O6z9jLxacsegDKLti6JIdT8
q3+kuKGv7zTOvlzvwfHo9iM64fzpqvj181rkSbnGzOBDEJCfHkAIfpGWeHgMviia4t8vRqeoPGyQ
0PxFcDt3AMpr2G5GVF6hEFJ+ZiZ8IpWDt5UZRTuzjPmrjBOEux1mdfpUTUP4BtK8aqB/PSnW+LYm
ik+/5iAlJWVcaN4CAhFsYR5PENLOLQoC1C/Y5p1v3Ap3cft3wHbLdv+36aIwLNxoQ9lhCStLC1yB
cw4vuxhAHhDvMTVZG0+XF3dC1vesJivgbLj1GcQvbI6sitcqI0IIO6OTOHFpUQajGBUhyYfd0v9t
R/g+PV5jkp47S4pD7sTgq+E5MR0WTzqN7Vws2ahGIQ2rcX7SzBzR5K7BRVkv1vZXvqpd18onqOul
E+lGHM8KdrFgC6y6R98Vi4OAx6qbJuYcXx2Hrgqi+YFHysxl9WSt06y6ZqFrAdrBDwzvLreMvu+a
JZqqF1jEH33ZIbtgFd0f2rKxpMmNiyuaAIFDDO50IH8XiN6FaCvZZgXkEeg1Q8wFpyPEUzHES3C1
SWDS2np8T5EUeNjsT/iYjAtS4UXYgsG+I07XH27Zc687dG+N5/1QDzCzChiW1Nd1mEW/GVAVYyAP
w2GvvSkzAe+sIengDvaG7YJca5UZMDtOrxDQ0KjB0wfzA890l+cfL0HhbJukuSDN/gpIkdGJSTFl
W6F+WPMCRbfArmgoNuPC5AyrsCPAJrlI+YujIH/qg/WFEP2GurzCJ17EbbPNTnWZ/2hNdV7d8jBo
Lg34X1PYy8obFHPN2UfkE8Lzq1tEwa8k6qt8gvNWVPdPCwmdCoonvU5FBnQOo/ryyCocnUQ059yk
zdBF2n1x3jR+cCDyEUAuWk9XbhhMYUzCvsq9/0nfSu1mLPLJ1vQZexbVaxJo4V6zj3yEOKMs7OuX
/hToRP+/UtNWDnHnC0ykvC32HQ2f1cOngokKoqbMTUp6+fDFR0H2lwDfK2ivifGz27DTuA7r+O0u
zCUxxFdXM722Xkfza0gBrNRGHnZTGVutAF8pKgnP7G83cR/7/VGWEOFts2CBqKXmd7J/RiFtVDuW
jhsYoMikksnI3/+lEGNQtfNlMYELjOdczLs30mRIk8/b7oSk69sSkTjaTbEkK3cw1ikcXWHMdJHj
rX2blAtizqG+Wg4pcjxwR913L7etvL9ijwAQax/Jk8P/ehOXHThLfWDGIfF2loN5eAAejc2mVnXx
BbCV/4VyYn7cU0tEu4GkiA5SiyFj87RVcMRMGkc7nKXuzZ05/zCd+E91u69FfBnqgCL0fhQiBf7P
g4SWzO3rOXMg9meBN4SZLaEJzPQWsQQTL2r/N9a4i9sYNNcVaT/jkXAsJTvf9NLrS2nRp4h/T94C
FLcF1+q/L+/KiHtc+IFUu41vkS40SZT58F1S+tz3RFJKXmIRtXzm0MioR6eOd5cqVthK2EXO/mY9
z/jeFQz1INx3Q25MiVJ9W2UsTIDaVFxd2wegOOrHE8egr1Iia5lZ8zrHRBjFr3cYM7P4aEX9xNrO
taO6CsvLVRZbR29hJMu2xU20Id1YQKVHk3pRsCoFqqRdqKhT7dHihutrUY/nIjIPn5DooCLLjFMm
4D3gUYlt2EKMZIsYTs/xh73zHLvtmJmKZ4zM+wedwpuRLxAgytUtDkKeUWHzovYE++QURxeXYHH8
EJD5NZvbQw6QcqM+XqAuxw2tGEaQePxEZ0MK3TdIQhsowGfzFPANKFEhettZYfkaSBofQhQhrfmz
1XwP3Wuw5u8Yn1v3LNpzNKTV6NVfto5VazlNj7oW2vKpHx/c5NWZLF2VfPK0wt4eUbVnW8y9Agzx
7JgjhDomBvsmSbfp6r0lZ8/GiWdhjoSIwfexHYmfqBC0w82UL5pRr63JwqHFmMBzlpKz1rXNhoOt
foThp+NqJsn12kZuvc7+1KwHmVjQWVazbp7/A/LAcOcTfixZAFe2tRqjQS7o1cENGmkUX481zfOt
lo5DGKpYl0gVIRlxRvqqrNjtmPY25nTfS9GqVsT5HVUpagz1YGgAvS/uhyx2Jd0e5k8rGPSiDvYn
jU8dGrS4bsL6eHYBEly1KGX9X2F9hCgUsp8HIrvlmtp5IBan+VV9W0KQ59WAa51IxeKrppGeXn6Y
ci4BxkxC5UoJpEocRlIBt7TMBEUVGlpMQc3vXeK4kqo9dXToSHCFZmXSk72FIvNR8VpU+z+pZvRn
K+rzgyf+ZrwqG/nhw4WXcH+CJQ9s1I1L5324Yk1N9LF06BZW5XPrRv3hhOYcTbxh05x2z9fVssYK
v8oLAe355TLqwbHJ0+pHdzuoFxsgof+gv9gnxG/qW2NYwHfxcc/LT+VnN8SZ8GZghRfoRCo9sNiM
pJOhQCioCCumTSvjjIq/F3gOAfagtvuOw1U9ieBRXpYMinB44z8mOC20CcrnsYVnQ1EWfbqVDGHC
XWCS1MNWEvqWytJM6n1SAf85KqAriZwG3ROE1PQvbggar6xOZpA1GzZTQY/B7A/3HEiaUVbkR9ME
XpIXSGiAmBjspwi0S/wf05BFgrtJHv2b9NWaU9bLaln84VSTLjGKEnqItX9CYlH1T6CpEQYthwgs
xUgefvC35VyDbKHazBcNYBiwqxdgpSY2EMkaV3cHGG0hxQ8C6UGsKtVw1bKnbGvDbZEiziEGyRyq
hU6CsjBXv0EhBX16DsDhbvI1gHqxu5fls8mjSnTELvLHOQl57RlY5mFe2U1rX1cYMbJtb+hTB2LT
crPn60zFCDdZ2GvqmYsG+KoTyHizPPALqV+xW7TNMCkOKf1rfptHODfkmSaYA36asYT6fqfdRCKm
GpBGk3RRe+bpfF6qa/ff7G3g/X35AmzynQUSva0hrO5OTqp1MXdyIGBMsXBge/lEmluqCc3mDYeY
xDZVlDm/QoaSG8pt7u1xiM34maC8XMc3JnBwM0q3Q6DSno1wethV5iAlt+7aAjfNkImy6rVKlFU8
ZxQoUMC/9sdHIaiRBlmu6a1wR7EptGuqfQzOZtd7n2ZTdBF4wbquvl3vHPfuwlSC1tX72doo6j5z
6gdsUxiM4gjig7irNinSc1WauweroyOTqOtrH42xPFRsICFbfEX8DWYM/nrG+TKxvSyAwb7EdKYJ
xk/JVQSzMWQSbAji6rZho+cYekAvx5jlWBE/Go5OxyNAZ6A0PARlT8nsvdYwdnYlgxSxL2niumQG
WOuzbnNZ/xUakx724k+479gCNFVIRR5qG0SOn60OvMukbvMsdVoVDZFTteBlP2I1VBdlvRWTEYme
HkWjxgqGe1WWCCXBGrShZgAL9vnxBc9h8p1KN71quT+ZDtOEWxMnOuNeuD8ivtZpLlUuHpbXFCaS
RTpr5uJ8+1hNOO/O44vToYn77uW155wRWDP/1Eahy8ctYVGk8SBWNhS8bFv7qm2yC8SLyzo2nnre
QMelhc+DTDyVtHuFpwlbuh5bBm0H7gaLrplzWkcyJgHTEUt7u4Cjl5DoHLnAUBzm+/h535CSW/1D
WTZK0jRUrb3WfKkhD+WAnL7/iBNaWbEOL3Hljr64R4WRhKLPKsRPx3NLJY34lQzFzUK1tlFhaAZD
YG8edBzkChMQ4HUkBGSGjcUayeQuD9GAZMZPVOVIBJlVsTEoj8O7ZOxokiQvU5oTdwv0/yn4kZaU
WUWzK0TZxnDLJra7GugzpQI+whsRgG/wpKGRlq+IuohrZShfH/KJ1MuA8DCgHL4VdFJMBBxx1XKh
ZVxv4qSyxB7bKUFm8GUsdErz2CWyJsLx0/+fcGBh96nSBOH9vRKf9boweDXCXe9V03m9BM1TTIrt
Om6I2akUt0p4XAZ8HlOoEjkSjNVVwaqnInHJ4lg1YI6DBzJKMAiwybXG7/upqpgfMRE70MVT9zbt
NpOBlFqBqgokmhf9eDacsL5HAlliDcT9B/0PvNgC5OCH3Hysb/iWN/+HKmxGP0bRhD2ewzjmb4Td
3aGQc/5IJdA6GuAGtxrT+O/ESCQBB8B+RfsBWhxuC9/nSmOeu4lOhkQy09xFwGgzax6TBpD2MT23
o5zYa73VnbwDgjkjCzYab7q7/x3zFyKx0NKStpuRpM7Yx5fMnIWwHScABKmy4FYqseQP5XzeFGkZ
yB+SlkeW4nlZg8NVg8lhTxONEHbZSDW7RKWRMZuHl9UhnDMcUBB4NM3FCYNI2v23ZBMEy9eleLwt
XZTOboCmmp0EvBzmV7JmKMqu6v6+WAe0DBKObGjClMXAkaV7H3HTe+C2FQ89q7dE/9CJ2wzfHn/D
tbc/5wL9bupSyd7Z2oRGvuSKdajie/nyPWoO9vsElZ94pWd2xXChQwnnH96NE4E1WLlCmvSQmDmh
0Lj0Z5ne6aoHtuRYDeRdIiR/0ZgmD4BFizmwV3fW55ZkF/LQAvX7/+QoLK8I7DodZPe9aQKaYjnj
t74vJxlwUXhSFZe/+3REpyF1YuV56OQH95JqYpQGzHhrRT2LwgSx1NY5IX35XZoeMpMAu/yeSV+X
sS8aTlpd9DEqhovFdOeEJ1FNq1+SCAykNhHz0yXGUxJ2UaEEa0kKq+96RyC6nA==
`protect end_protected
