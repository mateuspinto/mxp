XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���HD��P���bg+��+6,���~'z���ł�RPNlS!��4�j���Q�8����u5�]A�ʽ#9RQ
g�@�
�A�׬~�i��$TM@��!?�1R�	�����O�^�d�F��	�������ҋ�*�0_fc�����44��
m�b��Z�̜x��@e��ǜ��>��gGN(�Cw�>6����K;�A����C�� ���1�ON�i�j�/��}� �Q9������V�f9c�Dp/���r�G9�+�L�~KR��������`R�+Y�b{W�틿%�!�T��ys�(>�N��˶X�]�z7;	�^\!%j�{�^�6O1���(̽��ގ�H�wu���6�۔���v ��J^:��ؾ�V���!���W�hBF�i�D��@$I5v���!��0mI�;���8K�r��/�e�ЀI���C�(W�/�S�����b�0v���A�	���ʈ�-&P��~wA}6hl�qD�N�6'�?���Ov��$lD�R��bER��~���>��v���8dV'�o�~Ã��(��\d�}�n�����r��l6cw�'H�r���O3�B;x�ę[���2+�5���$��Y���8��R���O��QyP�M]��x)��4���L�� ����p���ղhŕ���d����r�z'��8�}�w�%~��3����ۮf�lz.S;���e�p<x16/Lc������)-��%M.���"N	�� ��Y��;$/��gV8XlxVHYEB     400     240]������y�o��	���៹/�MS#ۗ-	#v�m�G׷�fjmoQ�Y0�8U��\�
��*�Aɾ���{�� (k�ŉT�W�+'\w��.~#X뷛��R:�'�*�ia����U(nW�"�QcԿWy����o#o?�2!�5��vd�|J�|��H��u �2+j3|�%�t��/�������Z���u��3~�+<�frĔlN	� 2��[�?%q���%�DqBɛ$�{`�Q<:���߶ZC�,����*�ų�T倪SL}����N�O��] ��/Ֆ����j.��1�e���޺����D���+|)'��}X��]K���b��L7H��_�H�ϋ�7� R���������CyM�e����g$�ak$Zu��b%Vl�E̽|$��Q�X��/5�鮍���zQ���#��H��c ����Z���T+����fQ=����W�����nA�G8G��4.r�����mK�5͌�?�8r�3��M��t���F��\�7�=�)Jܛ��v���&h���.�G:�i��N��Z:XlxVHYEB     400     210���W˯����E�w��J�*'�c��׸�����@�~�q4�ĝc��@��41�Xk�-_�'���nHƙ39�=0�ɕ�t�HQ2Yx,M�B���P>K�k�)�ϸ�NQN�&�����m�$���s�3h��t���U��+Q�\��-p6b����}/J����$�;\�sfrd
g���j(�aL�^��dRͻ���¦|��Q��q�˟�o�M��Ԛj����D�/첩��hGF��j#��Hs٩ ;�L��ʑQ���]o�M�.H��;����N��a8��)^��3�?h��#O=&�]�����|sf	��U���`Q������g��nu�?ˈ;�7mз���ȯ��#�ab��[����˼e���'�Ҫ�xHTcU�&�'Xyd����srz��n� ��V�[ ����X9�8:aZ�nY��LbT��� v�k�a[F���He��(�3��m5F_�����*8�r�����V*�W�n��H��DQR�vI�p��lo�꤯� ����}e���'��XlxVHYEB     400     1f0�d�Km�����Q\V妠�ܖ5tz+����۴��i0��� ��3��D*��i�������F��naU��K?i������SX�0$K�Ud�@�{�âO�E&��-�`��k(�(���p�
�o�Ǟ�ן��|=����
k̟�r[D�F��/�]� g�\��Ʃt�4�k[�Mf��8y(��r3�m|p>6h#�� ��7�o�`b�h,=�L�}�*� �Z"�TdV�.t����J�5��O*U�J7�l=������-��ɓ1���:p�����_�&��`n���k e���G8�l�i��@�dG��wN`�hӉ�v3�r�K��f����ˋ	)2��� q��r���)��\�^0x�O���� �Cg�
�	�M�f�j�p-��WBmE�s�(��r�@��_��	a~�VC$��YOp�١`���hv��3%B�V^oo�/���7z���5���(�H���2;���iO8��*XlxVHYEB     400     1c0W�����F��������B�kj�Vx,����[i?" ^�i����[m��=�<*�sΛ����)j�o��	"�Y|�O�&ÀM�n�S�*DI�0ǣ���h�s��:qW���u�
��偷 ��Xݶ�U �����+��΅�x5q��̳;�9���e,��+b&.dӦ3���Ľ�><��W�����`�0��1:�Fĺ�@!�HQ{�>.���}J`��U�2�u�Um�WLjO��H6�>���!�<�J-�c+	\[D�ۍ��a�\?���+�O�Y	3!v+w�����Ǯ��b6וE[��fp|��S���ϝ�w煢yZb���om��e��k��,A���_���y��*��/��hgY:s�S��!x�X�O��P5���;`��ɥj�^zW��6ة�2��H��c5[���<�觗m�z�DaXlxVHYEB     400     200p4�%���l��F5ڕ����յpB��x���.�H��/����Z�Z�k��*�!��o �÷OX�ש�"�wt�����7��lJ�m}�ݙh��6�_r]�d��	��!Qa�k��Qս��b�#���R�-���+/��oGt����8k�42�����3��3��	��kE������f�Ī�_zd!f}���TL�E�́5�R�L���v���&��[.�ܻǫ�Jw=?^����ą/���#�����@X+Ň*C��bw�A���[fW�4����SpI0ą ��{��f�{�H�<8yTՄ0��	6�����wЇ����3��ɧ�y�� 5��2�4&�����A�'�n@O2=��г3�^_�A�7�l�j�e��ÿs�؇\�#g�Z�K^���o��q���S0V�l�P�-����1�+eÒ���6���5G�L����n�=�X���u@��9��k-��1ҚfĆ�L1�&g,s.��U�CjN����́�^HYBֺw�$_v*XlxVHYEB     400     120�ʙ���%�0�B`�" �F�ep*��kD�.��m�\�h�֌g�2]��f����G��g�$��W�cC`��B>S��=2���������*6�ċW�
�
�^��(�^���9}�#�j�iu:�݆ˇ��	�l&nX�/�B@��RNm��"�a�'�g���.�%����7�n�mڛc>A�q����[ ,����uh��6�T����f~,v��H8�R~��C��9���,�*R�5�b��g�ø�FLɎ,|T���F{��L�س�/.L�/�&%�^Xt+�#XlxVHYEB     400     1a0Lx)��8Kz:t�~ƶ9�x�8ڜ�lhVy�N�X7�M6�@l���|%�c6���G͙3{�rȣ�$�����	���ő���d�?�v�=h��А�N"Nwh*�����Vv��J뎭IO�OV�@�X=�^�m�E�C��1)\�BqUj�^���$`����6n����G'���偮Q7��#��8��pY�;rs�3���-�)���o�x�t~�_��S#88�ȋ&�w(����úb�9��sYn��@`��o}}�_�j���R��Uū�(�Z�*�I̫�_�ܰ����o��le� ��[�7`��m
#� �$��D�t�h�*�v��zg&���cx�2���?x��y1ǹ}qf���ݻu���������㐮��'�ǽ����-��qhg�b����J���XlxVHYEB     400     110:�`[32B� `<�o�Ey�1x�2o)ڙfU��f�����'�0����W�Ղ�[8��k������Ԁ��=���4��=�o��|�n�k���|�+���ĝ7��Y��,u�T��1Ն$gK�mf�d���1Q�#�õ�2e�,-*1R9-1�28���<��Hz�/[�5a�Br�vLC�w!��a��l���4��4&[X�����ɍh�U���5.��L9C����\|�s�'����A��{�>��@�A�C���@�XlxVHYEB     400      f0e�.��O�q��	��A�I΂J��ă��ju�8ѓ�����c,��ӡ�f���͌��V��W�Xn~��L���
U�������'4��8�߫>e;X��8�\�M�,5�̡Z���9�����_~F��N`(Z�pp�݆D-���DRR����K؉��������C'�̀෎﯃�d�[c�l�v�-��,ņ��'�ŖH�2 �o_�{����sZ�ɩ �h���H�ce0�6	��XlxVHYEB     400     130��1�uG³l�Lo�,@"���DWk�7��������z�^uZ,H��y{����!�B����MY�7!��ʺc
�"�n1p����q��5%򡋨J��-Ŭ�Z�=ѫ*Z�	�rW��!�C�'gb��^��|q� Q�c��� R�W�j�`���.쟴x x�Rz���\�ۼ�2���7jKI�l4M��r*�A{φMQ[�v�鏠����	?�,_[|��Z�Ƣi�&�7��'F7�F]��%��AW�C^��Z=u_f	5}@�V!�ԏ�����ʷJ:Q�3�ru��'�
�K9^B�	Q��݌�XlxVHYEB     400     130�,��=�&���*���ct����,abt�~�~t�Ġ�ݒ|D��I�	����%�i
L�d�D�A��}f�!�sAz�:Q�TnK�փ�!LDy�FDU䁞Ii_�S�ĜH?�hL�������m�߶x�j���:áq���$Ȱ�l6n���_�z�ǀx����d*$�����3���؁w�;`,���|°܌L������G{~,�}�|�ow�<EN�!!Avv��h
�dBG.U��6�#�ٝ�u; �
1�%���-�R�4�����H�T�ӊ�>�uqq����p�%�XlxVHYEB     400     1303lz��)�,*�2H�4xU���`��4`��[�
�4-w�W�d���K���'�!���#��eI��h7�K�J��,12&up��1ǯӭ���P)R��v���.��0���Z��T���=���y��o�\3Cͪx�\*%�fZ~H�:L�d1��ډ��0�3g�(6:<���*��l����H|$������	[C6��B#4�^��xS�TX��	\��>��&jF��]�v�\�6�έujd�o������eMr�[���	Ұ�eV�rC�3��K��dz�)A۴ve����V�;�u�*R<XlxVHYEB     400     190g>�7B;� **��Z!>A"]�Z�����uQ���0��L���܆�H���[B�)��H�S��jXP�.�H���l����]̟C%���څ%H�̺�>�+�*K�D7I�DmS�B�aM���6�f,}�YxMi�I���ȑ��G��'1-ƫ�d��@wݨCG�Xq[�j :=�%�5���\����0��ǧਧ�z��1���%(��N�[jZ�i~��Ĭwe��ٶ��f|�.\�{�=�n	@�S����?~�_�)�N�H��t���,`(&�pޔ����lc��;������.�u��y	U
M~H>�u��a�_�&)d8]+���B(9dn�&����?;����=}2�3����Z4���+��ǡ��	���wQZ�gg���� Q��J���G�XlxVHYEB     400     110/D��Ήr�&�0��]���D+|���T%�h#�����O�?�B���c� ���_aBp�q��\�XL�U-���ч 5�r��.��@�P�L��8�B�L�`��6e ���>����0ݫa�,�gBFZWjO�D	'y��"B}*����J��Ԍl���d������MfKK}�c!�#@H�L}�a���`g+q�-I
�ڕ��8���@�e/��%�	[pr�W�v����	u�;1��-�~�1�M��. ������H d�L�=XlxVHYEB     400     1b0�7��Jn�yR��s5��f�{c=��7���F�?�Hӂ<N�f��XrV�J��"�P,���P�R�ooL����ZGN���\xP_�[Ᏽ�f���W��5�E���_벏|�w�e<Q��G���WG�2�~o�����w�m�1M�A�a�D�(�5�����q���/(	{��`����y;:���,�Pt�0�\b�Q'�I>ɬ|��á�Fw���e�W��Y��~b��Ԕk�5qd���d���m�,x���*Α\�d�_c�5G�"�&�X�>�Ѷ�>���d���OF+�����0�<#�"��1�!����;�Ն��i!�ܣ e�w�[�6S���6!�� ��Jf:��k=w1��y�^����O��$�}�����AP�q�?ZV�X�Z��2�\Y'_�:5�1�R�r��k��@���XlxVHYEB     400     190:l�D�!�))��i�i�!_o�O���5&����9H ���#)'�XGs�5�z�b1���b�	�T� ��1�j7mg��t���_`�A��4q�US���Vi������*L�.�J��7WQ�Zk�*7nA4�#|��$�i���4��*� �n'����2��ڻ��|��>N���=$�����G�>�b��}l�rP%䚣-� �z鬆�I���6����K����i8�#H/h��v�>�3RAe�)=�����T�,��#�)�O+/�Ah�q������	Ά&����C-A.lAX��ѐrA��5��:�ȥO���-z3�l=�"@�oBOu6Y�޳j�'���!���۹�=�v����њ�+�;�����;�S�s�� ����;؃�AXlxVHYEB     400     120r��5�-�a�Q�o3ܵ�jF�s�3;����~�������Oj��|9�(�Æ�
��q����n�yE;&$��Fԙ� ?�]~���0r��Q��]�9���F�g/��ZF9̮gs����̳x$�|�U,�Σ��~ɰ��%-�����!�	�7;^1�����f�@o A��[�m�y��8��B�����L+G�A��o����P�?��}b�˄�ÙBj����4.��A�a���Z�x#��{�}Yʛ�*�-���6Zo$[41p�z�����c����+w눍XlxVHYEB     400     120��?��D퇪�C}�Q
�-H���*�8�	0�u-�j1&�p�4�$>���~r�F"mn��)�h��:+��Ixt=/Z�ޑ�/�l�Wa�h�_���LZ]xxqsky��C[Z�&�p+E઎����'t6�s�b�T���?Vk~*�Il��I/ ���rP����xKގ"D>	��5|=g�H�6���Ƈ5��#H)��-u�]�����@�y���^�W��![���֪5�8�BPXRVXU���t�@K)��i�]a�qD�c�^݀���D�;���xXlxVHYEB     400     160�u>��4�ȁ��>�ƍ�!bd���^W���1ؖ�y��+x9�p���&j�K�.6N�PDNT5Z����'ǃ�B��|�t����vL�����ݪ\�˃���|6@M�5�CoX�In�s�,;�%j�co��\�w�������*9�����=�܌7�E����=�����*+�&E���dNI
:6�՚>w��'&�O� ��/�_9��y���F��o{'��幪�@��g��=f}�\�(>�"���[�b=�cϴ�+"�"[�8�[4��_�&�#��f)�����+Q��q��s
�������dI0����0�e��%��Y�n��.�b%�q��g�XlxVHYEB     400     150�T%��4���O��K)�-+S�i#U�Q� q��1C<����Q*!��g�4q�C��ފ�6H/���^��x��|�.`�z�S�6���\a\���������!����f�Z�]>�(߲�Ǎ0�ۊ|r�)(*Ѹ,�{���$�F���R�V�=�zr�Z������i{]6:�6�>�z椇�m����ui�(����uF
q��.�����ّ���Xo:w5�y��*���綳�N�G?�4�����s.��Dz�[9֌�G�G�ê�����K�=^n\W� �����k����0o6�0¨���4��ٮ��j	Ҫ/�{�(��2)@ ���/U�sXlxVHYEB     400      e0�x�2��[9�	��`92ߡ:�c�t(�<Fq�_\65<��	�w����B,�M}�"��S�,��e��{*�q�2�ۄ�TԿm�����Nϲ�o*#V�{�I��8�ւ�e�/�����B��] �M-���͵����--~k���h�c!����N�4ʲ�X������b�Z�f�y��Ʀ��C����%�ⳣ��eJ�x +�dDӎלXlxVHYEB     400     130-T�|8Ђ�Qq�+�O�I�����j#�>�<I�G���qq�Ᶎ���Is��ݡ��yq�h��B�)%��wh�0�T��CA+|�ˎ&1��!<{Ї)v�lW�=��G��qb��&~W ɣ�2�cc�����'}��[ɫ.�vu4^ٍ�HuX�wr6'�^���\���F4�!PR���\���hϧ�b}��W�._��w��z]6�0zD���"�D�+\A�dU"����xԢL�U�jh�l�n�L�H�]f��,�K0ĥز�����l_򺈛޵v\2��-�bbʑ<Oa"�=�XlxVHYEB     400     140@V��!w�!LJȚHJQ|jw�������~������_�* )�-�X�K�� K�]�L�Еp~h���c�fH���6H%���<{D��I?��~�֪MihS��k@~�cЬk}��p)���~���_��mcYv���LBp��c�ShI��
w���Tj�o�9�N�0wQ���n`�[P��Qp&chUҫ��q�K$g��#Q(������I�g_h\�c֎,L}���tQ��⹅iGN.�LH[~$��-�$$`c���u�dF����ؼP���#�k���E1]��[�ҜE��x�:�܈㏔[3XlxVHYEB     400     1508�M�n�0˼/YO�#Qa��{Yif(����_l�b<�I�Z�M�9T����ꉧ��f�QW��FL�=Vl�h�����cixV���;�D�rl�쐾�K�׾�t�.��>ޛt��7~����z����?%��2n��Л��&2r/�z�vA�L�K�VS��g���%�'��"�$6i*E/�A�C�̌;�-��h��8w��]��m�$�D�s��d���.�7]F���a�I���(U���j�p�*�2"<�� ��G^ΗY{(ou��L�Z�Q�#Td�֠�`�i;X�!"m�XC�`���Tuh.~_`Q%#S���O��?Y٠XlxVHYEB     400     150׿�[	,v��`�Գ,ݳ0����S?8��- O�~I��,N�$��m��������/�g�q�H?��O� �1�?',����>	m]���#튞"��ޜ�?�Y�]���Fģl`U��6� uq�<����1��nO���Y�O��-��j����**�F�hB�XN���#�U׬���K����"7�f&� ?b����|�#�1�be/n!�Ȫ��})f�g�ӻش�����H�*:���ҷkPE��}@O�0G�!��d��6��I��٫���( ϙ8��]{�$�$\w��$�i�%���{��i�+�X'�
 c�gXlxVHYEB     400     120ͧ߾ aV�%���K,��#�&�"�?��Tھ�������cQ&��)gJ�19P�`�4�sP{$&Bc�n��,�����!Q��em���oZ0i��b���{�b�1�e����11��X�7��E��)$iX��9���M�5���O�DϥZE�=M�:x��f�A�-beljw��F-�����?\����`��D&=���������y�?��@��y!�wJ-�C��M��_͚eÅ��X�x׷��cf�"^�b���	Y���w>jmC���s�[sJ�(T�XlxVHYEB     400     130'�*0"��}܇�s�{�˞t��^/�1V�G ��y%��H��9M�%4��C���p�m���^��ﴘ��/�s��'V�w�-���
�}4���$=υ� 8]��%�mL1�k���o�T߹dmzPK곋�&�np��(��4����ʂ�Wb�M\[
�A5�Z��^_걅�@q��y5@�շ�Cz��:����Y���ߣ_N�Ǳ"�v0�k�(?���M���Y'�³�K�`��+��ݤ9x �|��v����,���`��@��|�g+�U&S��T�B��pIDċ!�XlxVHYEB     400     140�Z.��'���*:�`��@)桃�	mL�e����x�y,R6����%4Wd,�Z[iK4���I���=d�^��8uD��}��q��z�084�]o9n�s",h�)��*v-vZT��Fgј�kE~pO�#~�Nc�G�jG8��������.a��H0X���x��\���V�v�˒�#�%��ɻ�8��.�h3�KQ�֫9aX��%���S?+d��#�gzC������
�VR�kC�� 7OT��t�������dۼ#'c1��oJ uE��v\���!X2Jh����A�&��\O�7��
�pf3��E/��fS$\XlxVHYEB     400     120�Z)�!w�xm��+V�2�@�@�i<#�c���;���ݸ3�*��'�����z[$���u{_O�cY0�"Y��;�Q�`R��"�\�4�'_��q���3Q�Ͻ�9�D�X����Q��74 Q� o�� '��ޜ��Il,6d [pڟ�ld�3��
cx���ϰ�l�����L��1�˲m�/A����Bbi�Vr�1��)y���ϫ�hV�{�m�,�>�����[<�*��b+�ɯg���. >� ��kQL9X���WuE�dIIM4�Ac��=�XlxVHYEB     400     150�ʋy���6�n�ྣ�za ��ٹ������WY�����(�E|��/k�Di�HNO���Ȁڌ����a�Z�7-��<�] �̐�aD�`�3����[���z�A��S)F�n���I���� "�����t���m��Ȍ����mS�t�@��d�̍gY�u��z�����2`4�����R�e���A�7Ygb)c����Բ�,4��'�?칕&�!�V��^ϋJ�q ��jR~)^h-�775�������ER
±���J+0ݧ��@dʚ�O"tï����;���K��8 ��	N�R?S�e����4)Pj��sз�XlxVHYEB     400     1501\e-�2���H2Q2F2�M]ڋ����81��z�Z-��X� _�vX8���xVW_,Gc������#'�:D)�����1ٖ�@�B2���N=�E�@��ހ�.�&^Nx�[��4n�g ��}���Է���BED,�]����:"pʼk:�g�.�n�?>6�^��-���7�o����~�����F����^����d?���y�A�T���b6DqCU�� �>SX�6�4�b^��A��	�;�س=�ȗ�e���Uzv_��e�0��MJ�> ��J��ۦ�b�e�ˮ>"�8M��
Kq)<8�����%��:��<���XlxVHYEB     400      c0�e*��o?��,�^m�-�_R���i��X:��.�T"a�Ō�5�H �r�<����jv�0CTm�k�c��6���IB��z�|��aV�͵No6��bk��j�޷���Lz���]����|�����K��La��W@��,���٪u�jI��ъWݏ���%�V`Êlk���/
�IX�0��dK�XlxVHYEB     400      c0Gs�Tv��TN�ú���R�Ң�/F����8}#�i?D�CI�+�h���I��k����x!��*\K�1��F�c�Cx���%&�����[_��-�(7t�KWw'<�M�h墉�e�՝����J�����7m��X�:�9,&��`ʕܵ��9����p�:&������r�`�z��5Ö'砟�XlxVHYEB     400     130��BC����U �D7��+���ŦC[�C��h�y��n��;_�����#��"@���߲�e���e��Wy�~!S���D�b]��䤡r,uCD��lHùڶw<���0�����H�L�c�Z��G���2Fo[�о�7e�������Wnr������*N~��p���	��KnP�NQ��!ۋ0P\����6���}u@��"]ݴ4ҖDG���Y�.�Q�2��we���p���d�f��BК\���z1MN� R؝z;�聴-�Y�p��;8�Å�T��m��rX*��uXlxVHYEB     400     120	Tn4'��c:�$���OB����,������(A\r�?R�-�eI�V2�5*�]��zC�B]��Z .Բ�]V�ϭFt��\v�u^H�)���ـ�~���z���vG��#ƕ"f��:Ļ�6�n�+�e)PJ�Ŧ�O;�9)PN���EK�x磝Bݞ}�{�=�)ƒ<��F�ؿ����)Ȋ���s��E�/���KC�Dm��.�đa�����r�ML,ۍ�|a���>0��T�\~C��ی�L@�S�l$7���:Ԡ����:��ƀ� ���	XlxVHYEB     400     100�/ɾ�����1?:������Z2��Y��w��g�tς_s��M���('c^��;�y(H���!�9=�7��֯�£��ٟ�����-�c�����P&��x;�ڧ�R&��2��O��E<��n���s_�x3�sQ�3����K�q����F�re��� ^>0j�V�hY��A̠�[rQ�>[G��\
l��klM�6�~��:��1����z��U�bf��X[�aMʅz�x^�#�F��qqx�[}��s�{XlxVHYEB     400     160����<��aN�6-m$��!_(@]+������О:L_�}�b���=d�Xu�5}� �3"𻿫g²8�����"j=��`$��>&L�V�(M$�k$͑�{3�Y�����W�mf5ʱ���pq$�Կ��V?p�+���4����_i{	!�rτ{%�!ܝ,VV��,)
&H,�)�\�ә�_��	"g��qo�9k��I���$RޮoI�ݮv
-�xv���%��GS3�&܌8(y��s���er̜E��/�Gߞ)�G��ϟ�!�	�H3��A�"%�&��%<��o�m'�����F�劻b���g��Jn9uƏ5x2�.J�0P[��Z��tߟ{3�	%�q�XlxVHYEB     400     1c0���3�Z�o�A
��A��?�?=>�H��^O�agI\9��Ba�[&OOH��������y~��b~��`ڣ�Aμ �R��2�@��r�H-dɑNS!��B�}V(T��㲃o;^j0�@MsbLOyŸT�+u��#���O� �ݸ������Dh�~yʾ�>�|�$>��|�4�~�k&$�� �.� �1Z�x�t�|}�A*��V'�!���p�yK�H5
0���I9-wT@9�ݙ�?��^�P��;J��	4(�3p+ Z��}��.*�r�[M�<�K���]�0�����nk�� ��>l�}%���(�An�U<���D����_���NҖ��I����P7�8B�٘�Q���ÿ}�����E-Yr��ٔ��#�����k% ��nO��هI��<`પ蔅�4�Sil��U�zS�+KG4R�k�GXlxVHYEB     400     1d0ɼeTX��P�g!2�����4R�z�,z:|RC��3m�:��3}}���T����"[�fp_��\�M>�u����`���&�)ܢ��8G~��x�t�\�9�w����SjKCcp#z�Bxr���f��P�J�؅[i$t���&���X��hf�p9[0�H&��Υ�X��!	���E�c�1�x��cX���sn�Ѷ{�"gU_�a���,��f��L[��n�z�����O�iq���FZ���jl�9�{^�'s���
D�~%ŗN�����a<�
 [>�Ia�.%iF�o*�Qe֜�	��.��1�7����i#�����\q�������U3�#/p�툽)��yqdl��ɍ�o��� �"���rk���*��*5��ٱ���p,=­���r��A&*6��)�O���h���Zɨ��Cl�B��:+�JT8D��3$Z^/��� �XlxVHYEB     400     1b01
Ѐ�Z�f��S�G�Tj��e�헩0j��za� ����V󕓝>: T&�7��d=^�W����ҭFiH�#F�Ľ�]Y#6��t&[٫;%��=���X���T���ay�ߧ�JE��<��L�'���b��`� -�'��d)�S)�]�_)�5�m��AՎ���#�ח<�:��
_VL�"��hN�anj�ws�@�Հ���l�������!2��%{�=�"_�����j4��̴a��k�m�db��X�ٲhcB#�:��⏧\���_GNU%�k�jPppC�ӶNm?�ȓ�\e�my��蚗Cݎ��-�#;����6JI��.2݉���;���
�)=���,�dB,�-��aD�^n�K��_���lD�������
93(�����ya`��n<���+����L��],$G�P�PXlxVHYEB     400     1a0e�1�H�.�iV c	>l	�6s{k`��E_<����{A9�,gt��X~D�#?��S���	8oJ���}3nʽ3�آh��J�yU�s����#���)D$:Q�F�� 
~_�#�6N���$�F��]��-^Hr}2�32�z�w����c�	�έ.-�C��'� :n�￶'d���6'��_����W�2���AwEf{}��Pų{�G���rɧ*�gF�s�c _Ƞ|��������~p^�={
�Tv����7��`r��+��M�`�|�\����"��WA���$r�랴�����	��N�6�d�b�(���g�A�T�C8cr��	�`�Jʟf������=e��"��"9҉Љu��Q��혍W�b�Y��r
\�i�Z /��8��I� �@N�%�g�@�=�<XlxVHYEB     400     160b�<L�عL%�e_2�"��ӿ�,�gb*g)�Xr��b:�m��z���
H*��{�j>��Q�Z���������f��9«.EA�'8^�7�w��%|���$O[�_�d�'O��;g!:����mP�~��gEo���G�R��8�a�m%��ԓ���힬��g���b��� D�6P"D�7��|6����'��B	��c�T���^��E!5�ߵ}3a���_p���"�h1��V��
�����at7�
��ڊA��H>���>Ńﹴ~^�Fˡ����0�Е��Of�"k<%ʈ�XM=O}�_�(���O�c��A\T	7���i狟�������*bqp�iXlxVHYEB     400     160��>����_+q@��� �0��7��=��<&+���]������w����i�I<�<�O�1�>�8�1�DHt�Y�{b=�Z
"
x�;M�Ԯ�	.B�y-U��Ț��^�ZO�q���*m��.�,��%��Np�i�X!��Z@���c�����^d�U���]s~;�vC�����Ϯx�D{]d��R��c�;]��?����@�-M�ڼ^sA�Yh���
�]�e��l��c9:	��Ҭѕ��Q0�����Eb$l��@ FmR��O.7���N�O0��3�Yʙ�a���SU2�ۺ� j>cK�~u��L񥁄'̣"���{���lh�*�ɹ�XlxVHYEB     400     180�W�i�O�ךбZ�z��X�`��Jt�ا"Wkߏ��ՑV��ʂ�2�E�n6z�'E�߳�81\�1AG�RW[h�`|��LG M6V�2�M}QŃ��\�oȎVu�?O��(� ��[���ʳ����Hb�L��=ۅ/H��}zJ����#��V\��)�}����IL��r\��F�d��y�܈�4���SoJ`��F��y��^��W�����R�D�v�q%ԭT��m���\�h��͌#��<Zq#H;D:FئH�V��n'�Z/���fx�nay�bA���Hm���y��_#]�s�y�mN@�b��[�_��[G�?X���R�\c��~$�i���_�����t��+.�}��M�P�#��>xXlxVHYEB     2ed     1308�`D�B��+���e!�W�]��'0Ǆ�P�N#+ɟ�|�5�;�(�)����n�*�)�e��ÿ7$D�Թ�NʷORt\����B4.����g� �}�m������Sr���{a"�B�o�iA�:x�u֟�W$��vS�+��������/:ߴr������k��H�n�g$��~�+Tb�3؋2��C�?u��|xojp	ĭ�`�#��N�zA]����&���]q|m7�Xf���,XoBJ�S�V��%�3��-F5�*��#�_�(���\v͞&8��aKU