`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
vqMcB1ulrI9hmRj4qw4zYNRY1d/0/onPcR3ZSfGs21X+bpUkBKqqQyVCHJFH4mgveM6agw58kTiA
XvCwxUt/iJAD/X1U1tTE4h9Uj4e08aEVjJcl23yPxpAiXBnxy0u8JLrjgdrLce4W3DBrQlDEpQ8C
cEoOt/DpxEVd1OWXE6qNvX5loUxQNnOHKnUYFoylnEulGLMEl6Toe0G3nqC9TOtpoACsVNa532x5
MZ/Dfh5OjM0GkUBsMzCDN8OfzKiNwJoJajDR8IVPOSVSWbSW0qqxsWEPJE+QfjzAYanm88NMA6X3
kKf3mkyO9c7ZyCcen3Wep2H7bbhgF7+e+EF5Kg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="SnFGl3BG5dYVzLvdE/TocU2KR/+EqXWmslM3xtmX22s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26208)
`protect data_block
ONN1AvX8a/mgjBOgwnyTBSplFmfruHPCoJ3qiKQB8cmozTUYpeRNvdjR7IyiTEmF1tpUsV8rWjQq
37ckTIlUkh5+GAXzmTyIqnWNDtZND2cen/37ExX7wpSPO538P+LDTPEYv3uJhXH2+xgmOgvhgT2M
XeKwnOHw6AlpJHhnJsDO0LYkOxfjFBD3y007n8p/i1LZtGP3pHBvv+IyX/WjHUcEh8nRZq7s48Sk
04Tahromh/ml9YGhCpXnwxSRLODL1Gt+BrAspXei2JLgO1fRyb4OtxPH+iIexi6cIx42b4b31/0P
+vPcWGcD1ECoGdEri5bMw2IOnBFdH7WpD08gbJ+VvTXF1vOxlYfwJ0F+5W3FFZCbtZZmsAhFi0j+
JH9r+/zKJLiuiXu8Zh7w0ipF/j0g677tFyOQqlu+y9RqRlXkzBvgbxEgQVjbhOgmCdSdnaQEbuGw
aEOjHfUMyCZM9MONMqSwjPRqHkFI92VJhUkKq7qlcAaw2Ul81LWSuB+Bu+U2Lnq9muDS6yQEEzTm
1dVNMp/VBh6iW8ysZutSVXWTSD43ExmgB2pXxx+ReEVAP8u6UJB0r6+5zz5nYMJRSOZSFnl1XZ4X
UM/iNLHoYpR5FpITW6w4K9PFgDPMSKjAeq4LALple6dfKNI27SiEfxklh8ZohGX0lXMtHiI/JY2K
THopZqp2W1SwNNq2s+4wtPBMOxQYk85JZvwc8oYB0UWmt2GLbequ5J6ZX79gx8XPIW7w+Thv+ydc
E/LFxjQ/HxS3BqZM4MuMX7iJWRwL2F6ydm52KFc8ijrnJay+q6dnLXKmkK1g7cRP6s4+bEGns8ZN
yj9CE97PzZZcYLni+05gOX9M+P6Awk8C0TM+Haq/3vFBj4pO6SMYRRImeCyP6+ZOKZ9LqQoWMCiW
fKFVtTljsBLso6C9JjqQ8GFPHcL+TIgRdqUx0u+JfTWCOkj6qNTodSxbMhbTVlBz4fuyktmMD9wD
x1JGQ6ZAiE/zGBBQdqOOO70HG2/rnPVGsMWmxsYsYA1vvwTldMjPOvuXBRpZIYgoNlgpEJeKxWFn
+zEvmaxlq674EHkZC87/cR2x431lxIrQo+W0WfGbXEKsObf10n4ajP4YQ4qi2GctghWyIVnlicsi
Anx28g7bX4IgxPwwkxyCCGKxQtBVbCOe8WzQGqNg6eaWpAteQhdY5GEAzaa8pCzxu/aDJl1cETZT
AzfzQKndKPtMNL6xwx97n0RFL22mZuJ9Ay3OxSgX5MDInlT2meUdNA7s0GzAdZd988XTByFEAmYS
YM5/PSsrgLOw/OO1mqwVO03PEfaDxhUv4JlUun81iYbKi5dVH4DTnAs7dQgT3LxEq82FTWr+Q4Ym
RIER1anloBkyC7kWnnliZDhPZiXsR18hm5XDpfigVEFsGgEMzyy+yA2pMxOxxwtWmpHYajOxT6Ax
BbrbEpJBwXMh7Qhfzy3sgWpmHC7XnGZF7IUBRHLhnrDoX1V7TtmJEigdXUoCG9tvPSSm7W7vRqiO
exWFCouEhC450R+CTfT1IMLgeDk3GK7z+Qa9Nq2uEPaf3WBPfI3GyyvR5PsAg3fxcqupS4axCi8T
ghZ1yjHN+AQBAItnjga8XoVmWWK+HG708uB50MshTO3mFdzLs/0WWurAOKfUWgqzrcR3H+ZGT1/x
oPUNK7E+6A77wFh6NWNgN+ga8ANusIP/cnz9JixNmCIuTBjJRqOkhx2O3DTHPdpK3XvTGjwfuYA/
moSiRQIAkHCgGoFO4nnLa0XxQcF3zaXfCVWubXXWj4FLN6Jaj/Fze55ZE/4CMXhk1sbVZhF9P0Fz
YpOey7qC1swqcgaQMq7DaicyvIH+5EucrgsqKEwPTXmuVwhPzT/D1D/zpw6H2/Ts9HKDt3l+9BMU
Gh4906zR4kfwvpB0vmimPRKpAsz0Fa0Lcz7x1zFGcMyss26Fbgm1W0aVaPy67HCEf/EyYBbSXeeM
dGWlq2vLgQ1I4E3/Biuy/u0xuBbdo+Tsdy6AiTmqPgj+u9mQFH+5hjeipGxIAPo1BdyFdiMTvC+N
Dw6W/Pg9QCPXGpO9qvh3wtKnYurq66/5MuNiIYVc51UsmCbtI9NDZdfsQ9yLBHDrAw5cwKpetJSx
p8mCkpV0ir2WJY6X1+kTXMjON9UdTj3mCnMa2ALjZQepFk1tQfPg2XJGGi6IIGqOZMwnHDZD/oWH
6dvkwNLeXJPy7Hi5l7fyNUaPTKX7/fs7RLXJ0Q9r7uMoR+WMxXR4a1TBVFU++Bu/yX8yFnP03V+c
oAKSH/8xysrXjBaLzvqWSvSdn6E2dwy1EbVg7KJ1GKWmpvs3eRtZsxUwxD+tETiycAya2XH6jC1n
eIIPfsZv0gKy0IzV/JzrCSBz3Jzi1A7588ulKcifWB+jpJtzQHUOKmPkPo0Uk2GtGob2wYyjp4AP
PD7ZJ/u8MrCnyzvMvITTIE4CQYoduEWzH8h/YnYLdzi8sHYQEZRi5JRQI6GTPBTsix9dVwDIAzJY
3fwE3GeX0tF9QqOrhbQFRYeaTEnxDyFxxBeojHafo85dEfiifDrdRmHtnNk1gyy5yLrFJ0XbGnqD
scF6iyLeJTYc5/mwytxI1S8ikVzwdNpUAJywFbBOh3B5CTV5D63YeI3TXlImT2RamIr5/zkZrCnO
dC5/awfFnGL9l6aLhdYXTPDWoTLop45rnHPXGPIOiwX19yk0vB+Srn96z8c4OebelbCoQIHqUG6e
1Ykx7A5C7jn91GOnKtWfgkpSbslDqwkR+eBsb8qi5jyZiZfW8SdCB2CZ1gJokxn4Y3wRVFuBIyzp
pibflOrcGIiXTikYxzYgcHvjiZixSjgHmC1DT6rM0jG6s0CbCaI6JjJTVy1PDhJe0eDTdNhoVzY6
CF94ts5Hty7N0dvQK0CmM3YoYm60ysAwnKNx768p8gvyY2d+vSL9TBG/tl5PioHhRC3QsNTEhqDi
16KZ52vKogaickurBMG5H1K+D9VcZ4S80V2XHHMcu+UwI2PMIQ6arvPvCUTCjcY6+PtDejVeMr59
rhvIPXZJFGlEemzRXZd1DMwitIgdmerHZoBANnXtwoPEdEQrq/CMfGWwjE/CSokrl5+thk79+wLb
GZJNjNXp1wOTd5FB7jvB4PYekhk4k7ZiZWzGX330TghDO8ROWDkgiLjIMgEUzmBjxmKM+WORNdPP
SJKVezXB4U7Dgz5iOHNlHfcTsOE5K8fIVIyZEU+67m5sVTMwiq7krGN0FNA9yutIaOajfdwPDhOe
ExCiKNF8oGhxfSMSFGB1DjdsCfJx7RYnFZRx3Ks6sJ0BQ1sD1oj2TwUs2qrI0t1cvzDllt9gfbR7
IStNcVM0Giu7uLRds6cs6H+VwgDaR89OnBbF9u2Ruw6tG3ZwBDncTnL3juIBia82OrXPOEhHBJq2
SQwETm+uD7lvIm2qv0vKRpexowsahlEflTv+k/YF/brMKry2FSxhLTXvghxX6na8GQtLAIPefF8p
GYpUzndToo8LYHLdMvVU3kRIDPfyrqMoBnLCMYwmARu+UW5LBX38/g+xhgtLt7I/sO6rqPohqgkM
lV7Z8xB/1bdEBVG10rNQqw/O5JwVeoI1Cz4U0aU5P0vs/psOvtviz7B7Xo6Q4xbPy7qniTl0FCqn
rdjRfeNsTOaIDK8USsrSRIrlieZPjxouT63sOsLlFSbRYoJXQM47VDTqrX8RZdDU5+XldIBUBIU8
lnFc2vrpNArB+fxCauYuEN6y9VUzwo8HmSfH24fd3xVT9cDzgKzrWq0pkCDTuzPD8BXRfHjSCNPC
TNfJZ5zh3/a9/seotqu2kK8uk8C75diCp5LF+GOuDraGGJmdw2fYR/F9n2sqEh3FafI3YUMJNUpY
iWFm/FvH7gaIvAnkqJwFNHSyNcJ+oy3RfZYDlcBqs0XAFXW/aoGM/UzQk2gDZhYpyQMD+hOgYTvK
ksjpnw3YYetb86RlBeCluaQPmfWsbSwJhBKJ5l6Z0iCkf8eZmn22xNwdKytkWnutHJvxibTT9b7m
h9iUnYYMhg8PmXKzVrl0s5bPXCWUWQcbAlV2oCLMhrDGrMdn5CXc5XeAwjGRK3806kCXwR1bQM1y
kl96OpNNY4qoF22opHlOpHFswGTlGc+K45lVzk+PPi2nd/Ji46sz4a2A2Kj1ANdZ68TY94Zaj/yt
KBbz8fKyGLQCDXRQtRAto1pepPF32HGKEDRYOl2JI5ke6DOro+UIvkC3C1i6ghiI8upWUwjyd873
wwzmMijA6Z3+noBIEu3EauqtkPvwACenaqIo0houyMgNCIFXRadeCWyHUO5ocq3HUehL673BE7en
HWQ05c3p4srd0T7iaLLbXADTdFHhiQGWMsfxpCJ9SS91nnfGs8zM4cC3iMd73cFM+XyL/HhrBbJX
CrE+gBCyxZ3BVEU6GoI0ZjxyMvZugyNiSDpWBaK51Je9KiH/yqkL9l9265FYuBjWnnpmIXB7KRTg
1ZISu7NtN+6wlviw/QSPdVFG2UxzU8cnhB10CbDClOQxCDmFM7r8kFVne+5hfHmWy4J6lBzeRaNn
tT5cBtrRzsr28hGo5Y7XkNTm0TVqe62dUIiyXr35/GPfWBr87EnOF8FjDwo//OiI2jE0/fuGvWad
HvQeglSpZqH+AlfB5S0BTkvsj/CITVY8UOPrlR7P3X7hlZ0mQb4LaqaWgvHPc3FH+sPOUpijgeTX
gqzdzerueaqps4t4Popx1bRlF7HUwK+pOsDNRhwgGV1SnWEVlI1QeP259Cm1A1W0xUiF8NYpBtc1
ydGB/K/ZWoYTplBAnt/rGQvB3PIPDohGA8Tc1yd6Kb2z6YFzS5ui2gXFt5dj6vg/ddbVA7wIKjzM
fFmh9Ry54P7MtAzSwwQvuIs+tmVqP6QO0B1EjYXJ9XO4SVRDxZbNit8p9w3kJokA90Wy0PLdz22L
d6gpX+ErPhUE5w1wgj4QUSLY8jXvFn7Xdz5suTociZPc0CHem+Y36+bqXlRlWoQFIxLrsYaLHf6W
Mz4LvhuP+RjlpEigAvttecphUPVPxjJCNCcXfPGUMDCHTv+XIzhiHvB4hwht4OabTXO/EazAylY0
bksRRm78MnSuuqdSZBmaw+NXeK+dNTGiUokGX2dsam6WtwaZWKNjLsG1BCMiE3VF5tIF4yTFyUWe
cIY/M1j/nQAPKhkejOgX/PDVbhCfjs2EssWpbKM/cxF1vIV7uQJ/7DVMQIhddHSrcneXXNJRZOH1
FTAOfH12UsPeBRgeYuP22vtuUSDov+Nxqctn+GsJTnuL6kGZVWDmpg2R1Ls7wUBal7wucpS9myXU
PHOnw2FPFl5yQfCQ/qXqbmMIZEs/LKvCjIvGuQ4CIP1mViH23gayAVWj2rDY0EwovAov1/g9F2Ji
T/DTXjBOvEILeu/b2fcdUGLf0XL92kaASmvyVqV9K0KTekCO6AYMwN0M1j3IyXy1vanhcb4CvJtw
jsZQ/WY9ONX9iNtNiq4eqS8aLJhtyWu9GL2sApZEVYqdF9I8qH6QxgHb52lik9sYHaaFQvwGYC2Z
j/GOUqR7CW9pvO2zZ61YRRW18Tvgt36A655tjxWgSz+f0YIGwuIF+ZS9t8LS/UFF0RzGb9n78cqF
avYVElH3HS/JDWCG3k34GM0DGxNwIn8hyMP7QQusjs7Z815c8yt6d2hT64G5vRIAfFsH+Jf6lk/L
YRdhPajN2XLJ255owDDZI0wnXi5tacBNnb2s2YOIi3xXrLwZU58SlNF2de7oRfG3w7R8m3d1be/6
RRzs6X404O/896JmiB6tvPthMmAz/o+mjhT2YSttiv32PSUfTd5YGnQF2Wxya/UDWemlDWHFuJCl
IwriAO4rgH0S/wN0S3pKHrcGpXDjVkkWhcw1RzzkFYTXvNm5qqci7H2dCfPXq7HlagQCOulDrk3g
vl+HQrPRVk+rf6aG3d17XCgA/bd9DYS9pXiFHYsw5/8l93/zQSEm66E6yAzRTB30Gtods+Fb/mN5
64F2zDmgbJQ53FVUS1ixr3QMrWROmX5AuHrjglcifgLx4L0b8MOg1zY2TeWjv8u2bdsBpePDal+/
0AwdgFSdlaqyvqxaShjcISzCpMC3cdF3IJB9mcryI9s698Gb0dKo4AuHYf7rdYAimq2pyxQQvKDt
fpf6I3+tLr8O+JiNDbdd8ON+1JSJfeSNQ6xUecS/3S7dAhyIjdq8Ybrr0Pjofy7LLToim5FDIDYv
7G/hNpcQbLcb30b8b1bQhOZ1kUfeOAE58LegvSZyV9fAz1Pk4+S8LeMRbjYmWjbjUXAt88qgfId8
rOlJrYPeHNgZQbbWCk1EchxQyuRHfjfVVA8AFIrk5LyMxM3EnE5g+Z2wduDj/RLEgb85822NaaXR
MHrbZtjBLxGq5fo3F2DdgN6n78FD2sKD4VZYf4PeSnDNsrtQkoBXkkFBtU8EpNaOZxcFPq7RhVX6
5dqMlCydLxwUy7eOgW5vbXtbM9dSnfMj/oTxSGgmfPWlzDmpXSgTJoOGq7IlekBt8SR0UVT87AJS
9UN1BbZw0lmcGyGckUD8mT4u8SxCb+BtXFjFMY7AzEnVhq5pPNPM749gVQmy9B3I1VxyghMk+BcJ
uALn9jPSSefwVFm6Yvl/kQxiIL0523MWFfpBQvAFDQAYo9yjsOhpTYq+Xbo+1g0UFqb6mDev1oGm
8iyMrKidUFsklRkKF5HSygK8JI6qKx0upNyJtlaF/CV2fdwk7uCcXBDDqni0IixRZTpsSyTfTxX/
Ww9Efysqp+XuJ7cHNd6HW98J2YDLMfeHo/aZo/C/QntYw4taN/1sy+jPVbwcODPnslgilr/JdLnP
I9Ehxv6iUrElFgseB24FAqdGsRBYXV6q7zXK1c4dTshpfwEmxL+XFr29ySxu33BuQoiM0faMBTea
TyG4+LTwl1cqr6C0a/pZaR8VherORUnwhysqVxEiV9Qnrbz8Ex4YBBal9vctXvAAmWDlZfiQreY7
QHHrGgNGm+YMnUEXnUpTyXPI4pIgjsgooDIwrGukob0uIqt8Eq3YjqS3fcE3/rX/rYZdbfRyJhi0
nT/d4RkkUqPQmZSf8mcyVAIsPxWtyuTw77qeack63qxIRGfWV91wiT9h4IrHr1yBS0wIfYQw8qy2
thIrXQJ8+C/N9NFcqUUp2ucHdLDIXN40FDHfr3s9BDD8cQPTbyoCmjd1+Pxg19Hl2UmMXIG2ETvV
LvhOJByY6rxsktAdaIYG3WzQa45iAI3rypxuE5WvgRQjfBc3OQme2UBe2DsTQv1qet13WmflwTps
o6vUI+WE1oiZBvbarbiCI3SHChcosM0zMzriEO/fTkZ6dpkDI2Xdt63ZgYDs6/r6GANFXo3AaYDD
EU8QjgSTYA3+1qanfbFDq4E5lADy1pT4RU4TU/d4vWNUm4/Gmyx+MgajrBo4yQ2an66eEMLyyN30
rsf/T1dPGdhyrj+6bsSRWiln09ufmcAHJrOPn1jbRyDxTCfiJxU4ub1iAGnWlafe+O8pMXptPYne
2S0vw4Sx4jsnjy4xph0viNQJJDyiBOaGOO0cdXfOqJ0aeIM+LQ2sxcokhZqPvVaBe1yN3j4ZVOhq
nXDtJ2vHPv/Sn21TircPAcbJ4hoPEN7rBSfRc1n15veYFNQRdr7VPnVNoqJzYYC6FVeOZ7H1Ih81
nqgjEyyyFiHHj5pp/3M5didnYt8yLH8go9RHIZNVWw+MGFhfh2YLTOxT/fyCIAuQpe9uZ0dLW/mG
gMIw5H+7BiNIsib9joCVFc4dOx2Wn5M6lfSly6h/nvWPFYDjzRRhyjDENu4ItthIqmWkjKvAsTk9
IvFOnKGSvKn+A6Dik+Ddm/PwC0NtQUTGCKcSbQQE1rWG5LFPqjtqyy/pwdgUuoEb6XOsoSsbtS21
shmjQBGaO+kDChBMBM6spUa/KpIMcq/DSwqM87HmMm+XYtZXnU63mIecZDxjO5zJrTQDNtAi4+G2
1M6zMAl6Y2GdefnRTRvnJI2/FVVegv+WqOSHRQmBdHkHxWuilS7HCcmbJLK5TA0izN6AlbqxcOCu
K22lw05ggYHXe4q2/iQePwePnRJaCJho9y7FiqnjO5hBmnJFZpSrfsDe+ruBmYxtUGp71YrYXBoh
DgbDb+LDJ9mho4j3VNuprQ1kULb3WWQSxl6Udv0Ua0QTSfFXAqVnjt2LBTx17TfU/2eBKfPjKzDE
0DoB/KOTVEp2QQuy1dcuW2ZphgEVRn30wC6/ClYiMvwiWKSUG0PLzhDMA6b58+8Q+kpajfO0UDrm
y1zfzlLkEw9mCbkCI5tj1rNscEPqDRw+VEVkqg7K9fOSvF7R5zprgiKiG5zWwgEFPd2jORUjI2JO
477h9B8vjD3Vbuts4Sr3idWi8I5g0rfiQkt4BaXIcruoxKql83PyBTHsgen+u08Upqfm/aI0PyGa
S7+NqTJxxe5Z+LgD4Lmfz7lk5N5wIxBAGzecuCTsVDOxNMCcaFWsoYlwMh2Y1pJdRH+/qnJGbEFC
QOlt2/SisM0PDXTZC7XYEcvFGj8jotQ+JfvJAGoiA8lUO1umQgHAaONhEFUmTOhsRIwA0GAHzuvi
U1dNicXjgFfxdXen3Pc3xEgC/QmR7G48G8wDZJ48I4EfVF3JDXZIx8dYtY4uVg1bZaosebCrGgLc
9O1nh185PM/4nR3r9GbazBPLCZM1efVYxv8uwSY52OZYuesIe1McT66kQxjZvpYMle/jes2v8U85
AnBKA1MEaKCChj7oTwNLxoHzv1kSldB0/bJ17J41ePiAt/q73UFFGH880g6IXDC/Q89cw60zXfSL
CSGlwZ05r+PA0x52BmhBhjEqKlIw0jbj8TIUrCj/y+nYLgIMvU2zAJE955Tc8Y+XLcDLKiqkx//S
SysgzKM9RTm53AZTXRoY3zI2RoZ/N68hdFf+XqqisuxkNa+3HreNeg9XQ7OS42Y+ioPX69U98hwo
MMtJgQHrmqmPu4OGmG/L2nlyznjG9KMcwoOM7XcddZ7eEqRKT9NsUb4xpmPRS4RGi2vWtzV/CHGm
7i9EQKXDdc4H6t99ZiJMlDaDbT5guVBI3BFL+xAkooe6odf8pT+XXWiAI9jzn5HhQVZvGIXleWPR
yKUrlnWdbOQhw26weRgQabnGCj19Jzb6gSHhea4Y9l/PMQjFWpkEaiNkCkc8YIiN5mkZbRdVdVRd
m6dOO9siLP71rGGJJHD3YPx1gw+hVsONwGbQPQX70xLGkrgfH6CoyckAwW0tGHX61JE4udEdl8Iz
Y6Gw6YgjLQDtb/wQ6AP96RJ49jY7vjpzDQoTuYKD8McsKN3vCXyoTBTsAqsLtHDBb9a2cnuJ607O
H1d7WVCDCjhjSSBoW7Z3uoV8BhiO0VjBp7Xn2Gsp16EBoVzheEecUdyfaPwcyKjnHGtxqkKN5vkM
dS1msz7be05EDCpZAOjZpZ8N97ulSFIw5Elm/3mF3mfESKSd+5wCfLls7zy+gABGzdzLXeJH0BSZ
BaAuruoMI2IWBDsj735kCUsZQZSJKWA3/Y8dwx1IvkUMfb7FVZxTj12wQk83RdZvOgkVpjYg0Z5R
GibzXd5H1SAnYYwsT1d5lw4zKIrnCmAu9Q36d3AfbaiCSZXnKL4l1Z/Ye70zpBcbGXYvhNpNvcvB
C/kYI4C8RzZys6Gj9UtdN8+xI2a9ohOL/X1U56lHHktr0RpIrh9V+nKvVdlWm0xOMGoxkiD+Sk15
AsJPMkccMBzpPI0hgkd8LbsKsdIPd9I8q0rKwSCuf/ZakGL2P3/1AEFMeCWrLNYTmcBomUFVeVTh
WZWB2pAFmhG/1VxXY/w3ad5C3mjZXz67ctl0GYd+co6rOcvlHvtRvWC9GZuuQXBmR7YOT1gUUqL9
QsufpglHj22Mk0doCKUse/V4NBxkkWWBeH4sC1cH+BH2Sl/2dmChOTjIFd752OTGkui6JXdzYKma
b2Ru0ZRYf+nCuKY58tkVSb0YuxLm/nE5HRiLR3U2KCBAOGzmT5AKcHdc6pvIUSmkx5owMV6AdzmM
QGwF4gJ650mZd+pczBIB0HHPyeVEFQCC4+0wnMjBWH8iEADY8uV8UUzWAxmJZfajr4nDW/LO/zJZ
4X+o3BkHDYIx5sx9oNmqtdRi1+ZCCRzZT3eX0Rv5eTaf0X03F24aK4eP9xy46WIstv2WdfbbCM3U
ICY7jcgDPoNEwPqBNdQdLDGkhyvkOGJShX1KiGqIbT9lwY32XnI/ljk28QUikTOwY4yy9jBwitgT
PHaPvVOd23ji2oNJCVkOFsWVArnIJUfseIhENGt7bD0OGpM/Q+uutdIhe+QnU7mC7yuoBzHgBUr7
N0YX62bx2f0mExkR5umKVaa+IhigCBYlbhzUC95jsXbeQfuNEyL/Mz3pQH5iQ6L5SwWkbQgDS74j
Nc51NoE5mpW2pPubmPA90kVCVew233RzUG/qaqERYgRHwwPQW7tyUZum8ugVZ2Jt8Ba/cC+E316H
OOBZjz44GKJoV2LBe/lzmUU7kTjB1LAbB6Mtq22QpQT5Hyb+8+6TVlciP8x60Amka4Irhj6MHAJa
6bzid+Y6dxw288Oq2LCy8DZIMxyD2dszxRzLjY08Tj6NXBGGDu57siLzpYFEabD2YwwJwASgc7Ur
1Wk01VeznQnAWKijxs/sRb6BAYU26ytkzIhAFAA1YDfVkcQiwoa322x4cqsI8q8rVThxmgOWUztS
Tm6yCPCW0cKYS1r/JhoAARF8tSG2GUXFcr/744cyxHve0FaTX3lni2aPjf46MhMXtnVNvGpKQSy1
HRbeweiq8BIiLDemIQEd3dWhs3BrBMUxAt77e8v6q8Nq25mdTTTTs+pqbT+FYbbYZqQN/NkyB1Hw
m1bklk/tSQIMIVyn6KomfCwsoUjAdXBQapo0nB0CDgCvY9uWjCOePuJJehyC72E7Yk0L6QJHN5bm
UTJTzAQ13eO6+14aP5sRipNFULJRtJ6SrCjiBzJBVU+SvlWWTtqfTN83V6lIrYOoh/NqXikfs4Yv
iuBmDP3yoWH/2iKdRhXlmwjCySyHKGiseMmWdqqVr3jCivynJEgymDSn5BKflKeqWdt6DVnf3wu4
tNpiOjBLMmFsyjtNhc0dyxLBwI38biw8pYCf3fZgR0hgpyANuhSTskpR3g1/1wQ8UsjGgvBCbyb5
C721DZJx9Nl15ppK0MX9DsVNWiDueVh757NzkQLUVrY56o8+lgaUxYDduy5WXbpfOKlnT6g3IjqR
lUBil5tFjfxAqFpRecyoS+ljVQ5l7rtEssHAJqbnlxxe5xdqnybjfxzWJQhIeb9P00bmj60dNST8
GUl8B+rdmX8AEixhH4FwkCyIxTlAbe/RaouvIUfzX9BcchyHaU/goLcN6RfDEJCoKHgT8PZdMnen
fS7rckFyCUqCI+GDURYW8QYbW6kNubxBawmg54/T7wzfyHmD3cCtvi6JxuSNFtYScRfh/lgFrWVv
xH9WsOekoBULWU6CiZRSrbKVapYLLc46kVuwqtwXvDF5e2x3yS9ssBO7TPdxQ1OrshrYbbP/6Czm
kZqSBu/vLgCy6iTh5wyOmjNUlMNoMP6jzU7hZ+8PL2iObrc5Q2nO3QlRnxcmsJP2C90Me0+y10T/
K74C/dPNXQrDuC6g5jHPTQSLrBEoejRiQEIrqmb+x1fNwiKoHJHdf2cqcBwzEQ2GFj+v2eLd8eMN
Opoe5omG+Uyii94vBzIHwqOl/p9MyZZZ7D45dTnnyyfse832RICLX4a9Up5ZIfxFVsi7g5bBccjv
ZA6op+DqntgTz0ikwGBqYm+PfAYMO9I31Z8oslDLad/qf1lZToy+YxBW4qxObVXUcV65lPwZqABk
WF/xnR/mNKGjBeTd45NZUY0Sg97oKGRtb0rHzBhME9SqTS6gt88gx/baAJRNNmOzeDPoIyB2GKmA
3wUgPSVnw1z0U+9Sgujcl3YEZA6hG91feM4njVzQ8nqB7UeB5aXaXIoobC4+HhSMD+zl5jepN48r
5d6ksjH0Z7K/IB7bDtafMZ5XZGtOOoxgDwp7N+UyV5bShjOsTdCroaF2ErrJlO5debx49aXyWeuF
fCQDofBuSrYj2QwqB5EZq/e3BVwD6xAoFtrwpHw7SbI8YgLlTZqC6fxpbavIMro9lK5Yn7vioFXq
NhjfQABxqY4gFmbnicBC56EOsZIpAESrio3Y45ZnXquGAuYqVhdKbPSZ5XNmDcvn0OS0gkgx2PQs
ACcFbU+p/KWXVhcyPROSJuZAeGChNDohFiKLtnQSLBv99/LwNxCmHilDklmvqXS73gV2s0Jim1t/
Txn5p75Hp1kR0QnYpvos3zf/zHmqxX89wpW6ZR2I0S6Nhmc/ZT2pj/6e1+OlHMRq0sAihnQIpv7c
+uYb6myWMyVYxGlZys5GZM7NP9Nyv9cCjXDhvnqZELSikC9viQicQYliHCshqmBbAG6nSYKAPgih
AX5ty90GbLzoP77nHk1gnVoXQKFWjovNiinFUkTO8X34ZG1plN7OhO190zCumbLkWBdQKRwnwiRJ
2ivywS3e3HfrB3W0RP4r7kyd4qaA/DTDkWVcyL82EXSnXkB45j8JicyHBVKXYcz1lLSB5xvX+yoP
hxqmKe1I+q666eZom9haKQX3ij5rrTSjUWPhJXMfqJ79seOM6uOhuAV8HI0+G1/3VahELIw3Skrs
F81RbADklhiUKGJdTRPTkhhBYiqi7+Sji5xbU8PQhkzNPywJbBDe0c9Ye2SalgZM5Xw9QRlyTXRH
SN1U53p/+v9jQpjivw8ifm1dfcr51mled1o5PHFSS9kFoEEDISObSKeeBIQJcIEjzP5ux/ti+xcM
3LY0IJwlGF/WhSWz9uqflzl06kvycYOQz6dnvBCOIDck0NMhLbPelKZb71MOlU5WDETWwL+9ecW1
zl3vpktlthSKZDEFvHoD634fMd3ph4DMdH9jF9gXflJyCs6R1L23F9ewIMCGsVLvLi84iQRwvJEK
RqRy3JDDzQjtqv70GjcD0G5Q6JpfQTTS2NPIDs8Icw/ldfDGXOR7j/rGJp1YwNyVfGKpJ7BPxt9s
i3uXOIEW6NWYbXKXg3LoPJa9yKGmPMT1FCqUM3Zaq1BhTzrjwf9PU6ORBzCs4WUbMiL/48HNNk94
CjZhnriNJ8SiwjuayfMRP3JX1b1DmdBnFqbxTaBGU+4TSm3bMMl1k68bu3mm4nGztfB/w+z6+mQB
p/sDvRG6YBA/H7vhks8YRLTl0gj3SjMP8wgcfyEolTIEW/jLT3t8reSURpqKr9wgUpLrA2s9qav8
Tvf3TzqOyuNWk09GV1iqRFRWb4bT3kU6Mu10zh2NMuDuej6iKUN7YwAafGaueI+hWOgdxDQM90F/
ugw97a1p29PIIU3s6awoCkpD142vjYvLfSjhPwrfW0CIUcNJKRjr46vGQHRbtQ8hHUY5OIwxL5/6
2HBP8ZAePSi/GscYx+kCEP2S1Og619uZ8bNuxMixdXZFVhuwMHaK6BF7n3QLcbdcZ0S6vhY0NCBt
vpzyDjpmq1P/bFXwX7hpAnx4a6hP1QLk8VWycoWuHxRJROE8Jok6auSo5d3bE7F2eP/tMD3xgsv8
6f9EJcbS0F2gOSf+R2t+os2LCujuPxUGhE58baprJwnB2nMYlnIg+yUuYh1+O7RDoj4q5MCI6IG6
IZj4csfaifphq3LeJBmya3AR4Hxuy9cqihIEsfDFtlm7TockedICATdJO6Y8/HIE4wSzbS6QejS5
kHMsKdEDjkPIQU1Yod43/4udr2vzHSYm+JcauMpEN655fajy7wTy3jvqPD4UUfbJaAeb6CRNNAfi
CvH+A0MeIYsV0UOM3y0Dvu4qVM/6P7iM9fmQMzyq+1ZbjEfWV/kbYV7tziRdTZbNKoD3pQX/5j61
URvcJos0klngjJMF8Bdib78n8YySwsjkf3t6yvdsdVB+xsoSXzTxhA6yJfglrFfYkPld3XUkLp5f
IrNTVMelrz9/B/U0+wRV1Ju80cNGib+3SSzfZP6T305C0fL5S4lUbW41ZoPe6XXbVgQqRwTI4C0k
bOy9KBC7mmzxDp0ZFickXnggPX7PqRTe24Fwcgsth1Tzvfj8Xde61xL96/vd+3MhVS3QG/Sgh9yg
e47iZ6Ue8yFxeQnINxuhMSI7Un0McA8NbIgv9LOM8CMXlg1cbJfavc91ZXRgELesOSqllAhHHUKJ
dbTdnvPZgFsfRCe+HB36tpSb+WSP27qZrQ7hGz8D7kwzXVzEv5T9d7nShaSsUroR4JY0G5qt5Zpf
d5e+H6w8Dd4XaN/E0pTNNOVpVrXot2IJ2JtxxcTbK9Xb5/5InLuLClBj4JCciRmZd+sFp8I/CSwn
/zYRDUfNO1CJORbZbeT9MmXO0wyEtO0l31fHrfwig8zH0ZO9grlIlrkKpx0f+Ir3yE4muViIKHm0
oOVaKun5Z8dzXvo9HEB5jfbUQbF29X96b6A1NImngVEupc3wokFokoOg6BZkA0adVr1uv74/v5Uz
XxghQ70PFPjCUsdvHrRjTnGLrJPqgOMVsept8gSs92pItnmmHQ4IukvOLf8/gK7Ct8xKLR6Ib2Yv
OyluPCcYX20Cee0xbgk6AMoZe2xNshJ3u8m8DG5ijpLtdXjLzrpJtcNvsaaeCYGeD4oZFB4pWNFg
+UJjGVZMsX8/gWgEsi7A4GI7hk0WpYtPyO9mgGWPjKONsDxVMX/WUwszQn7UKd4oyHnvwVSKv4p1
+XYvjUHj1FG1NbK8aJpHSMh8Ff5bUh5TGECYnOEDA4NOvRZbmMQH1S1UPmv0s2QwCSL/WraUIJFn
F+W9QkfoSWc566VZF2eGyKu6QoHaQ5009/OPs1RWjYJXapEzJYEakzmmcqyZJK3OcA+WXD04YAW9
NQiqjLm9Xt207sG2Qau5M0797pD/sfsLJX8ARITIMXgOzCGkxSg5ooU+JYihZXmAbsS0dskEatNR
8UzbeaO0tr4N/ou73CJIFxko+6M5IrevN9rmCnp/8i+5iNo7jelA7N/5Zme5dj1+T7osUQwsSmRZ
jXqhuqUnqpakhRFQn+m0RTKtCARlth/6bLdeN8o+gv7JENUxC2KJwIJMDt3wZYca1seMvuHFmVnn
6w0QgJW5NvQcKuko6NNHlqkb/R9v/zgrZPfTmojSNSkdz/0hzveiivpLTt1YFXAAwgDBEcA6MeB5
RUgbRM1vqcpogB/szUGA+XFgMNCjvbmAVa/CuWx+ePZgurQd/A3Z9nPKZLlFvPXkUEgpeYQWye0Q
Mo10dWPnZv7XauGZDceLaI/XZoU2Rf9QxtWQIw/a5OAFSUQue868zYDQBqWPJzMcyzGz0m2e1u5H
j51+1sRmdet7OMrO6uvWC6k5XK3BLQ3GPtgKYA1N2g7zgC6cJ4W+TsItwKcjJAFL+gITLPeULS3u
RJTHf1IiCVrNi04j6fpHhE7WkEdmMIyefpNikeE4ke0mjHTPwy59sA8Y4Uwg1joUs8w7mT7fgUk/
Hor25ekfEZ25PAkuqHZlenKx7e3g1m7E/7M946qcLZwlAviLOBuPtLO048sHyTcd4gnlp2ojDxgT
rzUAF12IvttMVqNOSnUCWaPoUcQXMM0C16Uwa6ft1uqQrHP8uZlPh9fFhT9aKZ2NogSs8QSgg9BP
eIyU8nK2LI8wr5bVX+FnlXh/4d5MNwcJP4j6bFN1nFgu/cO8dKVAuk2Wx7cWqpFhZBCOkJMz5p+3
yf1rcGqaHgh8cLEO1mU+re6w7jBwvtPRDG0nwILb6xv6zNeKdcwc9gVo0qfU66I43mspNEtvHohc
oSGYwCxYlKz8Mi2wt51GT388ZvybLm2agF/NJ7JF7/o2LSsuBMTeGZRLI5RAPZ0WZm2GuCcNZiuW
7ytFi1XLuHCqum4tFKcqTtcxGa+joAPzHP4wX4//Am1m9hY6/fgGe3JmebyqWtIsHeGXyngMtLvr
MViwb86qHnopJ/6dP8qryaBcd5DLvwoxYAqxgEt2ICQygEYKD4lcweY9eaksIDjAXspXHqcFeuuu
W2+JUXjFIaYGGAvp8Pk2TQP2It0kpAVDaHAsBQkLqCcAG4ZZJTfAKHkHyNfdNR69tVaSZxDlqdMi
wALmpa7o0UNbge0+8TfzcZHAYRkPVxLf5keG+CMV1CPdKZn9S57D3ShuySNM5OjlwQcqF2MCQBhP
lfUqHEDbOqy4H3zajnRYMUn/ftlT0K30IZvWPR1K5cy8mSUJc7Taj+WQ3RQUqPp+gC8UpY94x5mO
aErdpqUqgUBy4aBxzYeY9RbyUjUuVk5Z8RoHVHniugFryFYB4H0ErBhsg99WYfpqlu3xE/S5zIUa
+e9+iiF0nFlxAvm1npkomgFZJKK3Tq6buWo8nxKW25ecLubhxkOVw8vc7YRXJCJ9xt2R6fg1Ahrv
FfIuwrg3Q9la9Rvh/5Wp1H4w+/m+MGah1DuinT+5scCX0vyAjNKzf0yfmmybvK7/qg9UbEptAOH7
qZh7nd53MgIFJddeXhgJ79l65EPQANnNNYL/JdLWxTsopxq18cSzQE33GCR76bTd6UyCRD5tQEDY
Bu5qOFTMi+B94KiHqIgaWAqsfizZSxX8DbJzVpTZFX7Sc9lzvd7huY1SkynD7Ce+Qm4yitCoy/1k
CAV+Jmy1/ZaoIJtNe7h9pYl5UWDu+FgmfhWljCw57dTWWCceIm9xntjeWFWX7WPPEdrL4a/PFU41
B6xX5FVXxhQRMfwP+Z/4BeTzgrrVj5yTWXPGd9l23oeohCojluCPt+7rnmfCq0s3ZHEgIjWk9+bW
IGacJmt25AhfZg25ZCCTfMwrYS8EiE7d8wFkfQkkfQ7XvUgQEbTKEmA5ko3TQWYzdb4jjTh391u4
+c188zm9RP4j+zhdRGzw8FiqzLJaK6no5jBsbOZFp5jAyo6RLaW+f10izYHSMtDW/dR2g+jgwHqq
LcYc6x6ID1gQEXkyz9QIuvZemgifJP/dVl3c4hSb9HNIcryfBuou3fyKdeqC992t1BCnNdVsUZq5
p8CDddWa1sIJc45gnNZhNIK6jhAewnhbC6DrZWC8BnfFLZhpWR8P+JHbnFNcmx9EVyII0lCjHSIZ
wtpqJiW1msw73z7lJcfpTetmPi7nSsM+VrDPjNkxiUFPwOOoE3+XUU0fKTGq4uMg+r2luB9n4XyJ
o/Ucf/GRvL740HMfuuvow2+SWVaKIsBv5SI80/wbuXbaR/V3tRbXstTL/2bkrheQGKoffCch27mv
Kc13MJinHJbZuXiSMuPGJQd2hLqYz4wuM1bC16mmgZm7mRETzdVUgDfDNe+xdqklvyqbcEvwiEzW
oJFzDedKBQj+nmY/mhR6fVxrDfa0xGGFDAnX3+6MFO9J+ISJ2ikjjCpibdz5Gh0kM6MfcV9Y4PoX
2sRF40RzrQowyit7nXBDpFtieJXjL8Mw4/Yqflxbap+hrWCMZfwlkemntawE40yGAuye7UyDEnzk
dKoWx/pkBznoprttcv+k3kLKDNIeKfOyThjHUokz+JIGoFhwZt+b9fDn1VwOLzsFd0SuNb5UbipS
OI6+VIlfL+dDEtHNmyHUTf6MLfnXNOb/t/OQIoH2eKwhEEArjLUXHvA6dN9axcAXnKSSSUkC3alZ
wirKB9Y4pzttduqOHciMAKiDRVr3JP6+Kjb0oTFZ2RnfXWT1bFhiqpLc+Al7mP6rHuViF6SWnN4K
35N4cSQTzjrELvMuXBYdFugYNDhmj8v5YP51bTeK1PtOOHmb22ZuxR3jIw4J4C1fIJATdahnIZDI
Zn9AHeCFLW15YqDxojfLxYEjuT1CykHTV1xN3QlLpibO7wrq5fNd6Al4yPvSogXAAKviv9v8yJjp
Sn6zOMSfCCgSV8MY4J+/ibe19JqFmFrjcYqVu6qPl6qMoYgo32c/VQP8BWAqgC3vagRg+Vx6XxFT
SxOu+dxKt9RdZXPsJU5fJ5K4S4sUGxTeBTLQp4wKPipajp1gtmoPXjRWaUowHrZiAENNionAnuwU
uUps181mqRJ9PYm+JxOT2phWS2raiOSiuiXaKVVcZ30nwXU65NJ6oI+MW04EJeYqUl/8sOlqsTNH
oXGqcGW0l0SzUjxFgLxmt5vBbJosHELGV3A6oew8SC9Bbx4SItSD5wzro66MEVTiqWTpIu/YkAFt
6VrNLk4Cvzxr/ksI9CNlv2etQOZP4Ayc+MPXjzLn8doV8d/BR1xbt5L8YxC8EkMLHW7Td0edpYZu
KQD5RZeVD+g/Ao3Uo1E6OONKQ7LuD1oMUonKhP9+JFiaEDyg7tST3I3Rq83+mGzgUYpkKfc5bFBH
3IJdNTB1eT3QS6AcOdXVsZ7r4L0NUQDqlSkn9uxe4DDSPM8ZlL/4f3PDaZxMx6DFg9oZhE9jaUPq
jhmU8NJBI4S4m43wBRul4RkPyo5C48jD06em9S1KBKNtVQZYgS1toav8nHaF3ZecPmzsRutt8TUI
cesbXk9j2JD7Tp4XdT+6J284CWZ78Pfy2UD5RC81xcUrRNrPJonZMmfTYcTTFTtufkUfL5proqSf
0INyDFW8QAfPPmJq9FNLXhLcXb/543FpP/nPnBLHQKFX0A/rVfZng2e8f2ntdGrBf1/YYe3kvrqz
pd0lB34r0et814qDrFUxAmy4Y3tD4dCh1qcx7LzqQU5vLXUcd06LrWfzBB4c6Hbq4/m/u+QxIV51
JpmPavwJO7kux4oBPmwHORvvD5Ks1a8sDbQYId4UvhpoikcWrUBX/L4dD1am+f9VkuH321Q3xHcg
MokjfVklRG93VVFk3HrdMiJi0lO/A78MgoxiJ/e+rfAb+pwWD7shptMLFhcinSMFNAxSzTe/4LoH
gjdznSAXQnEAJJaHS3uwcvf2N+/CfRmxF9doRzmOanA0KHMObu/qBDWqaJf6hd47AOsP5dIJmDJi
iJUyvTO5ReLB42SVTtQaqeXn0aRN/zRGArPMpvLN2Zt9lAhWqtWe6LgKP9IbPWvN6ywYXCPqYLq7
tlzT2qv70G3Q7J1zsSy8jS9roFD14TaKK8IN0Pc15CrC5Hkb3WG3022+27WTWND/2zQCR0K9TGkJ
O2NWaRPfrHYWC43micIh98nhAcOEOj1635m0/KDAUsE/ycBB4xwuqIUsqzd69ZbJnB2V9ApzgdiF
n91o1TjssVBOMCd+NIxsVyPNico6T254f1uXB0tBUCZY6BE/f8GBI39FTSPjroQT5G4F0l9lWJCB
9zCCGv++fC+qBkh2BM5YAcoy7IaYXbaFrh1EPw2FCYOYv80CTAc8EPbx3RYVrUyVR9RXw81fk8+4
PcOAtxDe7yAgeQTMy4qqfvK6ic0L+sZxix0rfL2tdOAB2b4pJmFNkqkq4PWAGg6ge0WOSDXlh9/a
18qEK/K4UpZBgtaAAIzUl2wBezf6j3CuX5CC4+jzr6ahRG3Guud9P6HBW06tviGaAKT+jIhJE63G
DjF28yKI8jMY/nC0YZ+QNRy2ce9x9qKHM2zDwFyMSDtJwuxtCoJWhi2VVtQ3LDtxp00M6+tXA1e7
RaozZrlltYLjiYcKEP4zKiCtKy5xFVyTKB0g1rNZussYBuNsgD/3voC36iorIw4GJiNlKVjVqDAT
W/FR0DJd8BWW2GC1YnqS6gtKVtkqjW8QKVX3UObw8aIodOW/g3KToX1SKAvfzuEFF9wXdCf7QAdY
kxO/eqKv1s3uOrMykURnX40orgrdX48WFLcXkvWBPL49Pg8Q8O4zDabCYpSjDG4S7MyXztwKCtEH
l1KvpwGhZl2nd4s7IlAl2ujqefHfQFuTq3utPAWNJ3kMqCCjmC2f2N0suIRYh4BFjvYg8HDvd0vD
YsCMwOyMgTDLaMBANvTnbDH89OtqnUFOisYDa1fLrhWg4pKPi/e6LekaghuD1HwGqzBSkcH1AVqt
xQsJI2pBtlh/237+pStMqg7NkX5uiXmjHlJxZAxpgVYtQdQCe5nVBDepowe3mDu2TOPm++jYkFbx
OD2mbNl27FK1VxteCIDzLCoAHA0vU27y3FD/7SdZzxwWlKN+37MLpHaLiDfE/33nAI3080+1z0Wl
F32U7OZmkZBF9GG6YHJqJuCQd6oxdu66y6ZNdNWUhSXujGfORrfRDeW8giVOCJ8gJsT/erXm0YPP
lmz5FY6YFObhjNSrKVLP0V97Zdnk4XPpJU9POLK7Fy0tkU1pqpYlU8Wr0ePkp7lCDUIVQOOa32/W
xodfON8K7JQ+cOhb302vIB9eFmUVYu7rUof/gejqMaTBJ8t9PeSEHR4nfMoME4Vo35kBSmHxiDjE
8ODbot6MGT6zl8Xo6Hor+odeZMWQiPoDhI7JMaP5YU2U4cvBfFDVc4B3GlZi5eQ11HwI0cgOjQw2
NJf0q+eRbPysZbgirPqtGRJIPhLCl6I9xt5rv4W9r3Oemxh3t+pgo9URVbBZkqgew4kgbeNcRR58
zaggKTyU8o5E4RQPA5+sn5QNGgstDDOBinR3RuqbCvYOskaUAFVE7cF2KOlqJRKEhJzTz42XaovR
4Mkxqo/mwypAXYCAZdk62NEph7lvhRvwuxNAfGX0KCQfDyj+VgkMOxEJfVcE4Ob+ouRmhbVllHvM
HQ+Q6WxUr6DzWCEWHVqBLs9x4GPER8L9TUuhqkgQ3KYV5n9tHLNgXSYmgmpUFZZTM9HpfhJxCcoC
y1z0T1UGGZ/IRUokG2dQ943qW2MjCHbEfRc00XnRl48ShSwtTVokksWOZNb/T7ZmgmIWHxLX/KHn
+vXxvBXb8r3HfpU0qT25LXSoQPHrYJSBtHLPWS6fZvjro/E1V/wyedm1atZBX7KDoQjhqWosP/Vt
kSZ0BdnF7hFsaexObyB1n277Zn2Sqn62AO93gelvi1P9Ijgkz0ttvPWYdK0xatGG+zdd0RmfnW0B
SL8I1dPSCqnlUE5oSPmHvuxUsWdvzEAtbtapR7HBCuKQqiqaqmfu3kvTDgE1foXzCN//6cwozHGd
cTmIbZL3IPDmx79N80WKAHcTSdBKpkys/YNOjU6ovm177uy8yu4JoS57DE25rsf19yWrJv7jbrel
ln+BZ2LlTcxR3PwcPPp1/dQC89lH4pvo0qzxJyp0kl3fJyypCANjaW7YTQH2aU+Nx4pHtr5oeDBB
zjh64Uf7BlegjanOSqiqOtfYqOs8ug3s6a5k0kY8uY1WQXnNnLoCp8Hf4MzmXEWV+27HYoNRcG0a
i6rplHbSdk5Y7xHBaPzx5bLNo3I29TC+0ZHk7kqWXSACqy9p0FGqK4+WsL5Q+7UpBysD41T3NeOO
lzSn+gYI8JUNTEp2NftEVLQaEeaBfFGH5HAZfrs/lGA979VBSOvhcqCs8EkkY+dB2dZrzE3mX6rb
QtPQ053zDJddQFGT+LKZIfW0UEIn5CH3SgEPmWCBznGuFD1B7S7Ohib1bLNVxeXMaMfsZmq9I8/g
vRWWE9qRsYVvbj76v3PcoAtEkWQY5aNF7IiCJa1XeuW+07AZ2OA/07+uQkceZLP/6p5uCqYML9Nj
/KmNM8LVCzSo4q1LsMpaXXwhufPXUfzXXPdqo2b6ZS4XN/6NBxeC3np3/KGIUXnk78o2rkRKfb0t
1EJPwAIDfTU4qtXRdXEZYNBb5yQb4xHJnXqj0pSjC39vzcQySAfrAhpEPXsGg6nY/64BV8zM/zy1
ePtq+XiITDi+GJBrnKHdNugmEU0gVAmp0IbZ8PlorWdMqUjCgB8XdJckFOlNj9lmwfXLOQsJvpQb
7mPlSBha894iNfhnrPlmnOqnZJBBGzH8o+pkV2mwJxcLI72jwgSPb2h4hVvEWcVkaRYXvW1EMMyV
6wasEmmb9cJe5cnQTflqvVkInLmIqL90pFsMJ51F/0U4bi6GDnhpSy+Fij+kOVoccLQhWeqwYWYz
n5GhoNEhqiNyMhZmnCPy7MWV9VfX2PI1KaJqEOgfRz4IyZ2iW8O3fg7JxLSUCzQLh2a7eUKV7dUw
xbA4kcCul01j8gb80inS8q+BkC6QZ0xKMBb5gdTD7luNpNR7kwv09+p3igE8uu7/sBKaGKGu/cFN
ODRKG/rDB2yohvhUgKtTfubLWySlnkbT7sqL1cCLucZXnkU1X2PM0YIuH//MiozxGfC2ziDVtBZf
f0RAeMLkK+sAepIAIBWQ46DMnpPHWJLJKUA4GZC4CKPx/yttM9CxE5iLU44EPYdJcvqVZQz8hPRC
w93593bTwsXaaoX+aLSci4eAOtQTsh5TAI4hbpfQwSdHwCAO9E5R61u7Zoaz3N7U3WF3X1FWDIAz
RgA9WQh+Wqg6Nzt+u3ioubrf+Q6Pg4j9/Me1LHuzULrZI2N59ImkjXAMlLrET3PS3lyCRTvTnQ4y
wqbo+g7kFhdF0slQ0T4rYT1YDWi2auouTjKRHcKCyfwfLOPnGmKRFnHBk2p1sQHeksA9RydllhvU
sFEy9Bp13QXlQojYp3J8HpE/rtc7/+idYqWxE+PtK3NcBYcBqWwqLEM8vO6/rC4tE8/UHGO4C2AK
18dEHfxmRBA0nbPcuFv3wZr1Kj7ae4fRT1eBdo14sKwLWuoee6luA9HxSYkP/rF4rxcyilf24Dg2
6YBoHWZes4Ov2Izs/LHRO0Vx1RGz4gK+lmHRGwZr3bZ0pxvOxrAKrvcs2dSrSTZLRLrVAm4DOuiI
WM4PdKMCzmF4DptcsjnJhqgdsXVIZ+yB45qyOJrJYc5zQurkwg2b+oZgSQZ5EKiqKVCx9o/jFu5g
/VbDn8cRnKp6fltScpR7830qG4Nuf5+zJpmyp5hBMqyrmLHFlc5J1ySRezUh+NswoEp8hGOsxaBW
1ZlgdX+Ofhcy9vY/L6+5jMHYfa2asljv/E5iWi2uq3IqQypoCkjxW8YbafDa3VjWmC9FP1xn7fHf
7hEW4gTS2IFInGuxhhUnmyeb0nqRDQAiCSgfkajeN0J8gY0hlToDiz7ARPa3w8cRGO5xf9Y8uZ3A
K82wXHgHlNZa1wWtHL5wzQL6V8GevwBqeiUOiDH2BsMwLqiuM0GhPdImddbeydTwTXWEqHqldo8O
SC6TxkUl43LHbA14e/6lKk3QrF50CNKudTTqnl4O/Ll4j5bMIgszvb68hf0bq5NkTktHtdh3n07s
m7D8QsgyUeX2F8Ek9X4amO2gRF2AfhApvZ2bycCR7oXSiWOFH+E+KehdwSGCPp+NuEsS1vk71F0W
9i6u2ta4PxC4xjuGbiaxnVOk2Cw8C91dcRGlr2AOI+nddnn7zCmYmepJBfMLuAJhO2pSSjvOXoa8
XTp+iHbsdaiUr1Ett5AKCbQyo7OyEvWgfTVgVxlLiJD/Yp5ZOmmXF0kW4CzghKSYDxVdnGn2Yq7S
tl8vofozIzdtTVvXtwzhh0JmDDFvBzAVEFOTul86/pzWU27LcT4OSi+b/Rp2nmDXF+Jd+J+8o4w3
JKvBz8VZrLr3SO3LkvBiT/A16mbSo2+qbAXvEnVmxcRbIP0T/MXkQPvJrrEnSCf/BhqTICEtEsay
rCsQxbcxeq3Et+mlsXhkHLxPnJI7oJ077NrwaTIw5Xg+94UJQCQ4L31Rqv8zevtlQNE3cVVP6EQh
/7n1rkEHGb0+1k/Hn6ZcirY7wchFxgbcuq75kz2YDa2wJCBC+e2TA94En1nV4OGVr3UFlymkBLW4
PUnBFEoozpP+ZDVg70NmzdvU6EGn+XwtUWp03jvbz/eAjKXcnEz/lrPg+qR7VibSxr63WXO05bts
plmuSSVc4MRrHrxYugqpGt0omcuHXvPGtoMGCkmtCP/eRY+aD1Kz3HLh564eNHPvzT7pR/0wA+S3
jqPTRK2h3mWnt5QLz1td+0Ifwwd9wTAbfTlrFRbPVnghQX0jAL8K691f6bXs7a+mynjlovNUj9nY
4+UaINK1Fo9EvvYqQJqQHERmRtnIhFuc/AAk6RNJcwdbb3NdsjDAlGCSJ2mY/qSHSNdR+YhpX0f4
a1ZmTASdILSYkohxxXKKEpmPoaF2dOMPEvh7Rri19/RqkV1MwKio9NWGY9eC4W9caEkAsajrCt20
cS76H++VhPhNpd8aH9wgLUFBsCFVYpCCEs41/WKeoL/sI52/RXrrQu+yCcU3KYbbUC+YuHR8+eJP
NJ7rLKI7Yag6MsY0TZb2eK0gONLbaP2nui227aGdKyCBvnmcwFlqM8L/YDja2lxrSm6/OMcfY9ap
mevub574kD2KOJpLgpx/wurXOZpGiK1E4CRDeHPKGJmQPlpZSGcevPZ/hupt9BsUEzWFAagCu1uq
ikFnr3YX00qQuPyBSAIxh+jClFKpE+3qk0MFxzZWwKSPuKBcmx31D3Bg9JwvsYd7uEhwYLS4hHo3
QVmbzKDOY2QZC6gK8P83pAFkwm0m/QtmzYA8bJJesjOQXNqmpoTuuHzboyk0hNP3nKU+KkP3ZTfd
yA543/og3KWG7CmGZvtRNBvBoQDcVlLbpT2D9C0bnqB+xSHT31vrz3kuSh4KJ0wkx9R8lPxU1gtW
LY9tD1hvI1x5YSFsF44ndkH31UYVEFgnTfFf4hefpc9HCWSI6onnzUwZNrdqSR2LlvhSCyD+GXAD
/akiYwj7OU3LQyGLQJi68N7jWUfWyEu/xR/XNFSWpuWNLUb4eV/u4JQi/zh3AZUa+mb6iHDPnbXY
/kaAZw0YTat3iLknKKIc+RlK6DJ7n6O12i3lD12b99QNok2877Fl/YI9vijjQdcNeO4MZysAtvK6
TVqVff+nHBzsH7wAMMcgV5yokU/PIfIZNXlICCS5f8qwxs71iz0jXEwl20wgjucNh2vZMNw+8std
JxhHY6Evbe1bU2Cl/Cw+TOOkFb6G2LTBgCqUnKPcJFpC6Ux9k2c89aupxcOOoyWXpkZ6d5XXPiso
5TILdCsuW7LEsNxMVhSicNx5BJw6oN1zIQe8Gu1XUdgcCfiC/h/wcrcUK5BISFrgfAc7aK61VNYy
GcW3B0pS3982a6AVNSedarjC3Qdr1HdRJkQBAZcMKl/rm79zDNpPEmndFdlRSr/kLrK0iEYwPxZu
zZDg3HKigGpfYfDMwZGMsmAyeOZDnXiDmACc+/OCCC02NTacZwh8vA8/8+MZxkV+iR/UcgZ82lrm
bcVXNMyDDqUBvU12kwn7yI/GaeXZhB+CgIlxE5O1R/n2jDg/NHNrigeysUXwiphXnX5EJiksE9oh
BjQzQgmAIGgflOX5b52As7h2jPubH0mvQFkFfJnACG7FuCkvYLv6oBwICHI2vPFm/RR66xZ9trav
a02Ys3OU6m6xIDFQyX0hRiAXeO/YxCN/+NZlbFIGv6SzEv8ZQfrtUBiKdFiGCYHeDsBTujNyWcA+
8sYsRyyFcRmvbJJezMUachbR6e0s9P5bSYsO/RfIQP550wUU+z6khr2tRwwFij+nROH8h+uDnmO0
9W6egANrmXWxK+YRZVhloAsuxGrMXf6n5K/vWzY3pQWJKK3G3nAuLa0lKEvoagNfOXaErxPbHIru
+9ROWloxqxoahTCQj5OoDAB6FigV4UaY4zLLbE7M+LLIGuX9L2r3wnCirgTI1COjHatRRzlB/5o+
r3l5ilOan+FPGJuiEOb5GPmhcktqLJ1yhwL5aciCclWTwq44vrzfFTRxnrLewtGc94j3bCAXy05x
t45I0Kf3zEQn8EvXjWUR/bviWRtdFvqSf72I6uR0nsydN1x8PISN4o3CnMacIaouuJdkIS+Ndgpl
CU6eF7GJOzghzs9rddbbkH5wW8TZUplfpQX/aipX2x7lt8Vdxa1qdCw0ARi4/CefKJD/aNkyCkx3
mmeNKvfgO6BSNrZo2tlcrefOwbUih211JmlTbt0w33ULDLhYmuEIAHlaeKeFNTAhoz64e7a/spmw
ndTdkD+KZ20sHCubYk0Z/Q2V++fdHeF4CjlNeKhsA5noCpUVqHBqQJrNqRuQz3vzPHbLWdVwa1Dl
4cf1jK5wcu/HFEMyI53J4apB77PpsheYAD4zBnh0M/aXuI/AvJ6ekI8gRtfqh43D6FbLRDlnVmQz
Ju1uesH5smh59hzP+eX1TNXBeIon31gix/F22BXQUEUshFwgm9dQxkOg9dmf3VaQumqfz2Fcfowd
4Img+/rAH0ipshGNQJEdW+VCPs+uRBKW3vlkFeA5jheogzalsNFA9onQ6YnbnovQL/jO6A72QOcj
Ggxs0kSuWgklrlCWxnPWm6vnUuDFmr9/+Dcw3aQMzUG4fpxF/ZFYffOAaX/Jld3tNUUcIsKln4T6
kSYDjEEO5eY+bcyrtcFPCEd6GYTm8Du/EwYuWbkERvmMpu+h8BH9kN9GRZSrOUFzv4xB9nob1sG/
L+cmRREGSMlPHhYbD6tI4ECRDQBJjBSiN6e0rXweo5KlxNreaLlReCSl1iHp9KVJ1M5ODFiJGqhO
z0ABVkrHmtQr+T1Ef3P534webwt3On7xGTVZv27cs1Z8aREXjgqvHmH6g90Z0noRepyD/V5/WDsG
0s2itWbqZ6geACJOOwMxbZ0MvaCbZ+KyF1VYrH4RM6fo/pwsaGlIEWO5YPWc86mBV0rFfdu76MrB
TX0DXTHS0ZX28Xk8ORGMpiaP0WTFzj5geX5IfLZTh7XGIXXd5g3r9OES4LS+B7VDdMpwPhJKVjiH
/D46acZd9eJ0D4wMs3EXkDfrYxPbzHfZNe244nNdNpf6+OV6Q85cIqmYcXiaojbE+7Cl9HIClAV3
Ji9I8Z/Y92Lhh8SdYJ2g6PHYw9ylWPgK4ijF38By6RIEi3RstNOBDAKsRRKaSwWtZzfnhQXAhFz7
GUkGX3kI4o2NsW/OaY3rEPROrsulJgHxLF5QyExcqytpKMk/Z/kJsgg6eJnLsKOYlV6IRpxrhDkC
VkiY4dB5h5mBjON6w2dkAR++DtbVlfNHhzXNHrSvwMSwcGhbU18DgZstVHGrkunrQyjO7cDHkOo+
VitL7DNlw3YU70S1lF9esO2HjImbzBspQYL5qUVdLU8pKhsr/r7gWGwkBMitCb+Srhm7Jp4KqqUI
sgY0HxpOtyGWa0ee9l+340XmM+B9y+8QfqfpERwAQlu+0bDm+xPyJUf5F9WNVu6zyX7H9TkgpLqj
N1D5p4MhjxYIhtomyAXCT+iPfKqNWgHOP3DBSzxrhK/XJstlSGG6MfVOqFqr80iYB1UdXwBYk8Ix
v/PqNaxvpfpngCBks4umv2Fs3gCRv/2h7CGLF5oZhR4F4j/hx8zGMal2an5+rh6mGFxVNDkrxGeK
lm+bMYlshSqBRSBtaib+Ph/30Z5gEz/nAMKtkM4xB7oYhK4X3oDUB2Re6x20rq7LUfvKIXIEjqTx
CnOHbdiq86XgHAFOuV3td/c56vEXn9jSya0hJLYExDWP4Sy+qSjmdXs47yoZPkic00rDI+wOUHpH
bHiHDciWwT9zyEKCcIpud7Yx+54bLWuQ87zDr2g5G4C37+sXoHm8XuqeaB1D/3KsSL93M7/V5Rl4
A1EMSDzYn0WPtesHeeuKCnniWeKsugwDv1CoVo1zgo03d4dDo1CI9zFy0Eay3Br65ZBkTvzHhorN
AsgRgzJAz3qj08YX7cbAjsLaxH5rQaQMH2WBxQrLh5xb9EOfECuJMVUOeAjfFbHI6uSatwomAnds
B9nmXysVOjzj5HNZNp7MJDqbJU180E1tLMaYeFV5HHMEQ7JRc7lgnaRQzpxZYgHWeiVncFCg49K8
p9V3N9pGf3GHnVK2A8h0nWuZsH/O7zuS3cjuXZEemch9a2tR2udu20530vGegn2z26V4g47+/9qR
nIVL+o2vghrk7SFdUAgKichSVb1Vtt8bwxrtq1YbDZglVY6t44cNKdMazajXlbNjjIbdYysaGNgO
//oOyJAxi332ADg3WJCIW+Ps3otGsuNxjQ+LdefsFDLBPaqa7OfTCmByDEihmiXPBQk2Mpu+Q4lf
87aQIXtNf8u10lJ5EOEnCcQIZ/UiOaCDbiydJEM8foGSlPb4fUUL2vEbHZ1PVMwQ4o3yEn8Cltai
8jGx0L1yzFzuqyWvEGksluUruWU/Ea56MFeD9q0jKmorlF50asbeTvsAv77Y5EK1BBNNmN9R/d64
hLaj4jUZUk9hKziQE6+rUKn8/bCpRfaQxvQ9o2lj3ZZphAiyhiBm+NwdFhYg1EkUwy1c2mEBEct/
8zCy7vmUhKHJQK+3O5XXN2iIs9ZvXXmGioQXYqk/0fQfmv0pWBOxWXvnkC4rXnNEoBtGNOzdRxsw
5LswFKiUMgL6EYd52P3s+YDMVGClME4sv3ig35vDg2HtuIJnVbX2foqks88/A0RlNmbpG1cVnbkV
0kSbKeCYU5xNGo9YeCGtOsBRLJwoy4RHpYxWmMReO7tbDP6BzG8OB2SzU57GjIlhtJwp0P1IFjs3
ubz9Jg/5Jczgr15NTSO0tlni+4HcfNIl7SHNJb4lugEQqSNLb3QkWbY8khSxyjIXNydvj/XLk7DM
5gvBsPDkUnuuUVxf+2lwYQsizeHiFsAIMVcIO4EQgdG5r27317NtOex5DqFgh4N11opyHpFMDkjD
XYcLNjDRYijhMeGHNmL75AbL2oZFAvRxtdIsqk75CdVu3c7Vqi9avMN6k2wRgaSrly+x9GYlfsOX
piCGIEW4qS3q0SdsizBVcrD/OMfaCDjkQg7rZ80Ph5QI52SKzOBE/0W8oKKt3y1uiRppPTjkvgTM
M4aecF5P7X6P12+76nZBm74C+fo2L3UNaz/OFm3PfGYHTp2Kyq9RMaSSNH6QFs4jyO1RaTeCExPQ
eCD3VDZDgr4D0G2BYyPB7KxaxrrTBLzYJTu9Vsl556nR2nVMATRXzC23o0ykj4Xse2np+lw6SZzV
TnyxizRpdhpNauRkLtRj3EsXATm9ZJhM1MLx5s7XNUXoQ8eJJbAe0iWP8jTyYiCwvk2FvNvlqNWM
az3nTNr7+g4is2ssAeJXSRF26uw3r/OUC97YEMaHKKoB/9yMiyXyV6EjwbIZfb+lK3ehjV8QnwWi
tzDHHQgEmJqZi6hz75BBQuwO/zvQk14dzMtQNKo6uUEI+KhU0JVci4SDSk6AcPqm394ZTC/ITrDC
ch3e73MnF6WbWTiWVwKHVLPtL/BcTVSsyLIuXHgCt6XKLw1+hI2PlPclQH4Rstfwn/JxnEmMcJOF
lhNYcPMI7fUYZ7gYTe9SCIDW7e86GmxdluMBPh/kGnRw2fSRrBmxCX/aVssSZCvM5AquVVjwn3su
ohgizNVuYFXQ2QRnsTi7leCA2S6x9bWL6D6Ae7/LLpaevOxPftedEdCHloM7jjg7TRzqc9fVwN9z
eXUZCm4ScyzeT3H4sEiEeQnvDR3QPBhFlVVGP6t6I6Twoaf06zSljWz1d4LhMzNn1U4dx6pdD5V9
LHxbASxFVtTc00hn4epebx+8o4uHihXR8n5SrPNBrL+7cYaW7Ls4jPyf2N3AopHUWRf7Z5f+jNRD
VoznmhAABMt4OidjhUjELx4Ze10n+VdDPwTHZBDlj/eATRwSFxT/0MDIqABQX+BmpnAjC7vfDvAh
yLGazRE4og6+/1LnigdOD96C1Yl42vBIJrJzFTQR4UuiqCr5Ja+qzmQdv1XCyq88uBH1ADU6IUNr
xgcUf5o2/i3KA6ioyNUPR3GZcvBu6fHye7hub3NPyZdN1LfUZEXip6rcPUqt2CHqzuHds3Gxi3Uy
nxIsBsFjJs+D9IcGU1nGL4/V07SxknUk9gSHZx6uL4p4yoPGYqsnmRE5I1wc9qORbQRhZzKzN8WY
sWJQB6F+TU5h1V3/XJT2zJ0FT7j11OqqpmLLb+KA7aqwUsv29PoeikyYi3JSFVj5d+VvynMiJEsJ
M6MY4pOVhSM9Us/SQ7hhMEIMy2NR+FotBMyJgBACVn+73NFIVAsNO2HUWn2x03I6vGs9QixjmVJ0
tHu8a5J5aELMPASfiQxWeAnrbeQMxY1c0NFgp+k1fV527abpsK38SOoGAS/XN78yOijJACxx/vcb
fKoSL9/Wd1qktzh92dLCJY9uImxXJGFQ5ACIBBReuJuat29IB4NPA6RyhSOzgGbmpR1ya/pw1SjF
PQRauAlLRN9qXmg4tSuCIZGRocsceAd/cPLPfJSRskmGK2kr6az9TfXgjMXpkf29APx6Sxp89bfK
/nXnX/5ubCaRDt1ONDzD/3v3RNsi2GFG8ey0FH3/S3AJif2wBbqIZFJfZRiVrntUxepkM/pvi3we
aI3Vptt58M9dyGeAbFnZQF5BITnyjdQNn6DsVIwhL3FFflzrPq9GOB7/v2V1tg7PiD+B9gpBUuTW
fhXtnoUXNcAD+ADiDRRWwWreDHtd9iU325DXmgp/A3IdsP1okPdKiVL2PO8UrMulFG+GTVi2UWCa
gmC1FmtCVzPB8JwaBqo+wa6N8BrBkBfDRpukZC1UisJ3RgunBFMmfiOrFrsWOWqdIlEQFcCVfjfj
uwcZSP+CArn8xviaN2AnxX4hGLeaxK5ZqxV9my8Ry1teDs1YK6SI42+ZrwxmX9OxauPNI6bkakza
61mIeGCXiYx0te+ykWqdG7J6is8pgDXv3qdI55AdYMSHUGA0uO1ARt+TTKoF5ZxtxSYHLCBL5EFt
SMfTsbQY6ehLJ6y7xxRnDqmsCHhqNwBunWI+YFv7Fus303HlltTXvqwCYmg1lbaUd+aPprfsgPAA
kLJ5wve0Dh0IGzYU7zKI9OwLw/Zy6z6nAIyo0XrGh40U3YikU5Uok6vcOmWfmvXqa9a2c5oH8E/7
QBLUPI6EM+Fb42PkgRn2bu/wXCy5Zf9voCzuQP/cf5X/9rMlbZ5hkyFesOeJzQnpyZxj9Lboimhc
Gp768/o4X7r3uP9iC9yptP22puKg4QdEdt0bsTwfzk+pWHSdtoXFjdsXmnFSqzs+rLShIdOpmkEh
AFZ37nIv+3f8QePtnc4I8QbCx9O7AgO/34ZTz7YWSB+AfpYJkkGyCkxFptwoqom9G/Z8CXAMM+M9
UM8f10tzPi+AUY96NBfOm4PIYCYZnQksf7Vmuuz01VB704CieVknnIsn1h+JVOYWzx9y1pBs5RMa
6yd4nFx2awTMEdBTip6H0Sw+9Qa7chWz8pkEqPTi/1NsUfjsynYdMzjCCF3o4esOgCg0rYHm/p/8
Xmuf3Gd8EHdWqI4Qt8B9Fyq0E124SmpBCGuj2Pu6WPDAPldkCOCS88eG1KH18wYcbo+FCINytS7V
Lrmf50qh3TcALCXlFer4CGxpyMU6d/DtujEiJWBanXNBaQj7O3mFHQbwazwfMT60UD/QcHjM2z31
gG0LI7AaXOazbQjK/Xl0sKRwq4kAMnmJye5Gu3ap8MUDCiN7egCtJlvjMVrcAuxn4YGHuKz3DHNK
bXCaMEC7ZIKeNLREPMAlso8nafyAkD5ULHGrA8Np19FEa8CdfV+q67QqM0+SYUfpHOiJLW3nNdk1
HpB13t54ucnAf712X5o2J2gzvul6K0VxfxBKvXvbLCtEDtNH5Hfadcf1VysyghvcCOWVqltkGzBT
j32muMJcAKjNIt5LPyL+4crOje8by8idIRVeCOtl8DKerC1x/tgATeDbIE3plmX+m6fz47clN9vX
IwqI1Tsefq72U8XifY3HFgoT74Ul/L4nm9Uh6UTEetR8E4IXfOkd4bapHtHp7znaNcmB1tLfNRzF
eBth7R/e8oRiBeBSxxOPmCV1b6XbQfLSZrnRpDvPOrjWZaVtDDl/gDj1rCi7VxSCIMAcnp4xHSSG
BwZp2kXzHOsoSMgSAgSCuawk3U0jGPhP1Bp6HQuD8Yyt7UA4SPQqm/bnE7HnmB6L4jWWb4FH4kKl
ScQ/SLv088+0KGX63yqnldktNMPpMM5BQ1MVRJqq9oTOeTTpM+rQ2LVXFlD20ckGYzqINI26ABv9
StssEV2UWUK3hQnDs2kxjMuphBhhuqyGlMCgimeQ8SLyDdCpVNJpbQeXFbxjUhw4QTSS2nic1s8y
SzjZCXkBhCSRJ0+yp3ANJPEbDfpZlR7QF72fyH8X7ZlhadB/1UBFhi2xxmNgIhmaioCb69hfTCUO
ng1mRGHoGP3BRCb0ZEfMjZqfUsf09t0Viby1LBojlixGg4/ZoRiEiSnSb4olnC/gNeab27JEn9Ep
1N0LD7RuTdkgOGcFsDGb2EmH01UwbDn4Moxvao8r7prTQkERe8fxLDck92ta8bq9uNhS6BkMfUM5
frzkF9igX3yi1YNT+iWd9k9rPG1Lt84U7ljqaZJde/MMvpMmgPAFniZ6gmWjWu1kuOwsAsiwZAMB
CKHD8enpuYfs63KZPK5caIuW9ntXdJr0PmK2eM8OvrGAqSgZ+GuNDMEmX7sTKBIrriGbsZ9qd9cJ
D+ioRaIfSqJKjtirZS8QmtRQz3SqLfeeYcw86sE57IulNqPPvrlV7h4b8XvN5xmrPpuTXoZMUmB2
NVTBACVH5JMfWikCITlZv73tM4rf55tfTerZHTf0cInVPDd7YtI7VmMoF7pHVYQFHpq7cEGoU7rF
dgQAmtBYEVb5Lg1AN3R6a4l1IQ+VyAcXMLJmy9WIPZCpajM7UVoJ7Ph3TRWb5Jez2stB/Wm6Gqor
jmxd/jpTVkMaDeIz4QcSV2VyUNrxNPM5mX1G1GfMf1vh4si6I2HkLT5+ybMIRVdomlL+rSClCRp4
zHmPpf2coi+BxaDq7t5rD7ybevtXTuoHA1HW06XAdVk5wnbF0PsXW0Ma0wKBAHnISSYczkj3nR/y
YEo0SlQgDmCWsTnpXXQvkfcpG/1qBwLqNXeOrUBdgnr8wZVDz5SdxFDsX97vROyrZsshpjgiwxid
FJY8g0IO2h1vF8crYwPwRt4jaaegE9uObIy1OhBiDkttqTnNZgO09ANyhwWHq7med9DJPPBPN/Xt
dB6BCZnljJTqENVG30ncr6O6pEzKLM/APsaxI/po16I6tlkxggYu2+UTtS+xXkgYHy9Bz2zx0VnY
oIu1dMsYiq+YkY6HSgxgziJ5OdeBbX+jSTTExsTmwb6plVVvlgUff233pwkvsiz3XAjHbj5wGFYG
O9D9JUCy2vzaYkXCphn/A5hkjcIQPcC/GmNbTSIWlaLm32GYkzvqWfJ5Pe2K3nKUK8nU3QpuZcCI
1GFnjxJahFZFS8xQ0mQ7IAfGiHd3tQigcoFDkArrSxTi/S6z1IXJvm81msnrCafjLsAsBsEyLeHk
GP6jtOILlzoabFwWcufE8wuXmu0dPLDsZgX1fNpTOsXVehiOUeBY44dkwILIPcud1IRPgxVscb92
TK0OgEZNVhttc3EHPig0Rk7omur1hmmD+UQoPzs5lc5TdxNBd+BCEAM60rl511Sw4Gpe0UMKbGow
wM3TJ4HdbieRDWPUURyOa97soZXjB+l/J2wisKob9Mk+5uB8TEdbRp3rlkJnhY9fEZqKFvgAmiTt
fvZE3d0qBpr5qbiR6oQZgJVypWDlFZJQxoWcld1w7EBS1vbqTVgIA/Z8Jlxo+HwqUZHJeZfmuWuy
aAX38T4Im0SJxU1whN7O0kkLNqbEnRhToGGG82kYPZZwqbyqOHkIeiE9AmdPxXBGz0rCeuzKE9oB
Zx+3ulEbwWApmADk713OxXbfJpq81PrVPdgO/M4kfMmKOCu4dNyH4ykiJY5t0w4kEzYIgj4e43X2
X/AFTzb6QuKLVE7B0YsTwGa9HJE4cZAsSlI8yuBCR4AC861plaQizlMEDF7XAJS3zS1a5Dr5HfVQ
Mx6s+usbsU38eRp3zibn7xjCIQh0fy03/JrsYNGUShPngvkHJKFtwf/IoQZlX/KU6LGztuccCCAW
A8hnZeVai9C4vS/yXn8xW3q5K+gRYFrdQUagzFJisQ3DMbe4kGOb8fygzQeZThmVWwTuxwbtTRv3
TgF8Ba0hLonIwVmvgwuCjayryqgNaj023S43OypspHLdVVQXwOl/CMM7RJSBfLDrQxKzYkfkzPM6
QXnBWcBapF53eCdesXHOBH4SqzBBAGF/HVsOez0O7JLCWaMUP2Be6o2nPRwL6DE75TdhhF9/KHgE
wdTZ9ureB6v9OqGolFKHFguqpRiumYTgT6xJCzSIKfkbFtPnEyB42rm37JQ8wqOjZ20dIt6Nv1By
U+cNPiy/P0+kQXZeHR9J33GQZJWgre/sKCQ4oEicZd0nKBSi71ITkhnCheh519rvLVMlG3Lhjlwl
DBi76PSrF/s1N/Q9epny+JQhtnL8sxVJNbyNdS18X6YSexZ4CczV4DC65KWpSstRTvWf6j8rmqv9
3Y+I1FC6PEg8mI8nSuo4Ya/nWmZoHu5/IzJTgQVZYOwGVf+B3jEl2qTeW3D/iOsMmw/43lBRebWx
bT80N0y3YszJ5qFkmlnsqWkRVTR/tcKb2vDFz91A6H6sHRoMRBtA8cxXSn1GqzUXX4MgyO7+RQ5A
BqVrplrsUNoBAGioiRZ5q9uavDiArbA/dbZ3ik4EIi5FqU8fQNh5dFSMR/V95eu2kJmExtRsJp7G
Rjb6W7Xh8f+P8u7ztr4xt/adTUTUm9uEm0mx1n/l+vLMtHwRTkuzwiUM4tvXkEp79arcZsvDAsR5
LJXheQFN9LdyHvvV5lyIcr6aQLdUZjaIT86cl+EjPoTplJAZ59+24tY97cEw0QW7d1Hi87Qjok08
BpmbjLZgqnFj7oyU5GiGbaaJyvfVl4wk6bqkmoFuAWPy7u7EgReoMOGmspq59/fcZwiwGJPVwRuO
G4dmJNKjyl9RIQuvF3W0j9qhkPScArEnSC0Wa11E7rBNe9KpUCK9lCeKWf7/1vV/7+ttq8GPqcyi
DIoeEH9uoNaKiYxaJZF/0AcOiFG9zbKRIaTuWjHJfbbV/o12THHHi6hb0zqb/ew2J3tAx9suGl3W
w0FaMy+EvHW7l59mIWSRb6ZJlUTH/Cq31nsOUpudaDsSoet2oVNN/u7f4qqcN/2irVCHr24nlyL1
5zmNasgFMicSuHpHy4EHPsQ1b2Fg3NuQL5fPesRwtBLI0XN/2sDmobxzIQ47
`protect end_protected
