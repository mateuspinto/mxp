XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oGX�/��� ���?��Ăg!�1U�2��7�>R��^#��UUU�.Dȶ�qWi#�B�CZ��͢�~i/��׌k�O��=N�LtCW��Q�Ƨ��"��pkA���L~b�%�\-����Ch�|F0!T�2��+�Н��Fn�l��h��84��7�A��&��V��7� �n��d���o���	�E_��?���n��h�o<P3(6G�[^��~��Y���+�!t6�\�-����wӽL��B�������B~9��g�
�ӛJ���At�Ӧ(|�S#/O����s�Ut���V�@����/��GS���0�Y%5�&៧˹�/�>6GG�!��q����6�֝��7r��p^�7����akv�۷����RB�/���lbm]x��;�U���e��̌#���[�(���~����	�`s}���6���8Z[��?���j$'I�KO�p����6('|>�h6d�#���mH6�����%r���=�P��?we&�#6"���$.ܻ�w3��<`�XC:Rݖ�}u��z�y^�OA�(y����dYڝ��̾����f+L:s/�����>t|�\���ډp)���(�|��7�ӵq<��*�+S>�$plq=;�&�W�AN<.펲�m�ٚX �����Jp�������Q��@�A��-P/��%��Ir�=uS�E�?�H���t 1�嫉�l��^�'�e9��]���M
���AM��:�e�~�c�˙p3MxjH�ciֵS�Dj��MXlxVHYEB     400     1e0�t��s,J���9?m��m��鶴��F�=S��Zy���}@p�5�6kΐ"c�����`⤖�3������0�B^I��/sp��N�h0Ҹ�6��-ڔ��;0ΰ��
�Aa\:v�4� 0�w��Ď�BHկ��g��]rǸ���L��+��_�9�~�3��6w��0�P^�YrP���7��R��� ��LILKg�wJ+����cD�
�e������mb��S$�;��G�	S�;�H[�Z�h�G|ӕ�]7�����梪,B	����=�������(�Z�~�ˏ~�!&˗&�n~E����U�y�����fn	=���JF�΅�o�翤��>��v%}���PT�x��������o��V�����3�]�=�+?�
q����L��Q����+(<��o�7	��t,�y���8����bV %-n)0*���z` Nʱ�?I&u���H�d ]���nM�tXlxVHYEB     213      b0h����6B�����Ugˊ��e�퉛cч=�Y�~���l��fZ5��?�B ��ǚ�q+u�|��Q�L�8�;�E�P�1��%[�E�us�m��
�����S$M,�$����Z��&^SVS9!���!�r˯�0T&�v��?�6��	U�'����N݅MVa�~�