XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����QA�d#�V/�T����F�WK"��h���z./�N7*Ց*�ע�u,�v�{���4����K���5��ʈ#+�6��^��̦�_�X�06�g`��༇��8��ҥ��m�R����v�Rh��%&���"!�Z�D�7�p�5�����dt���,��wi�d� ���U��(�^{�����u��~�0���L�ܚ0��T^u�=���n�+�x�����<99�/ln �{����8����Q1���Y�K��.���'��*�d,Y�8��)�t%�'B����egl��f�FdU��&[I1wz�A�vh�����x���߈(P�y�4?��YlF�/Տ�pm	'+��(G*�T
�I
��� �=�'��y�b��}O������zS�+ޒf,2�d�Fkr+����|9'U�K��T�p�v"f�c���Gt� �ȴsJ����(����TӒ^�F2���9�8мg/��(eOګF�f�*����Ht��d/��i�dn�@����%3R�����2��l�bb;���+7L�H� ꭻȝ}�R�9�!?+�jn:���P� �tj�kĕa|��R�Tɖ�P�P�a���f~u�2oS�Dŷ�ߩ!Ŀ[&�� r굄٨5���O���0� qX�Y�j�|]\��j��|gs��9W�u��e��o�64��<֌�ͣ�"i�n7��H�|h��5��a$s;˅Joi��PR#���������٘����>
��Q<���XlxVHYEB     400     1a0�����Mܭ���A)J�Ǵ�`��Bc]��� 'H�H?�b$�4��،_�B���>�CL�ا&'�X=����SҚR}�	��	�X�n���+�x����b&fK� οq[�ۑ�ⷁ>�v������R�$\�]A�)&]%� ��ɦ=���gS�Ae��~��*����י<	���jFQ�Ŝ�W1j��w{Ɗ��#�o5�7;E�Թ�x���n+�T�<� � ;у�/���ƽ��7]���1��0��+��-�g�7e�n5n�4Cl\5��$O6s|�7)S�J?��C�=S�h1� �$����.do^'�,��ڹ�&"�O>�mv�w�$��
�0�ĝq�����3��x�5P�����q���CYq2Әc]�ίJk��-G�� e�_%484���ܓXlxVHYEB     400     150Ʀ�4�y畴�_1����J�Y�Oc�x@���Аnvt3��+P^���2����ah��[B<�c�P(�%�:�l����W��ӎ�{�vԸr��%Y�ɶ���B���HZkwMr��'2��ˏcI����U�)[wb诜) �	��A�Xe��2��e��D����s��=%��l��ᆚ�H�b���܃qq7�X��{�>t�a�'48YÑ��5r�����Q�-;|<�Nq�H��V>Fp��	���O&H��Ȕ�!w�/@8�4��E3����`IK�=�FCz$�׶}Zeĳo�^h���/b����₅&�>����B����^¥;XlxVHYEB     400     190d�3���g�?[Z���p�3c&����b��R�;��!ԋ�3/'iS�ǰ�V���h2�Y[i�?��?��i�֍��r.�4ϳ�ç_�Z��#m�	���d�I]�D��"�@�"R��_m�V��J+|�;� �_�V�b�|�A����W��U�2� ���k���.�+l�_7����Ӈ�?j����V<���O�˹x5f��� ~$-��?�<�WF�H�l8|�
��췚���z�ި��iةy�ݎn�<��Ɯ����M ޥ��)/���5:��
�rt�~�|_4|8�W�f��7@䰘P2��zd��Q8y�a-'C�3("ɧ���ݜ��bc��Eox���K��v�lWD-��qB�"!�����P��y�:�;�N�1�!��U�X�a{XlxVHYEB     400      f0U �����23��L�&���*C���_�M�}ih�]��Q%ả���������l-?x���κp���2*/ɲ�B��T��`c�j�d}m3\���]@��x�K Y=J^{����~�7��V�:�}U��(ʱ���r��=P�l�����7��݅)s�:��1�/�����~	�lE7��ʈ�6���,�?���~�v�������c?��҄֟r�E/c׈���km�������XlxVHYEB     400     120��&wj�=��QU�g��}�3� ���#�-�v�}ڠ��o�=:S*�4�4�灭ܤ��u��-��N^M�Q�ضL��+�跇��Z�Ť0����L�mo�B�_��z��z�"Z���E!���(۲ UA��c��m��q���	�Vy�%�B�.i
�|%�e�M���(yV]7	��������R�`O�f�P��x>w�駀�O�5?�T1h8�@��Us5����N�$Ve������j�|�T}=d��*�af���*�J�pFR<;1^{:���\#�E������&!�XlxVHYEB     400     150Ss��gK����&O�!���h	�H���&2�y�0�=:FBt&���NHnm� ��" ��Dƈ,ݭ��\/�A�O��`�h�`���m^4~��4�[�(T��4I���M��B�.QĠo��z�6O/�9�����vC%yA�^�����i����� ,f�2Dc���XR��I�>�|ĴxW.��}�����dJSvoU\u��n�����Ef%IG`+|䭼������hIv�?���I������b�~G���{F����aB1�A4�y^������"Z
t�����@�~�LH���:�Q�I�4>���d���z��+�"�3:�D ޥ��yXlxVHYEB      ee      70��d��@5�l[є��cc���F\SHfq����R̋���5��Y�uJrZH��o��[!�F�����I�R 9$�w���_�i��PC)'6tWÉ� ZU�~ա�=C/�i��,