`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
jQeYWZyaOi4Mh9L4J512KlIIF26piJtnroCqR4kb2H8PTcUtLIj4plkifjIHh7lLo30O+Vy+ydmC
XwWseC4mug+AYjxtV1+mzM6vjsQXPGQJOW67PTy6scgA0StLVCM1LCbKObf3fMmXmjcXKqNAZczO
mxkQJPthMj7b1stFwGNnW9TNBgXOxUl/HHcxvr+BlqO5sAbxqnZO8c7sgJqfE1cEjplrC5s+Lh4n
LECQw1ylk5wD0TkH/o9SlZshIqbJBEBQDlVUo9sFu44EfePSuEDTlNIn2cMx5n8VyDH982TYL00O
Ng2iRoSwxFrjE5Ev5nI1TR7lxrijV0VYGE+dgBIqaxG1ZiHoyPBsaHLj39Cr8fmO1oB56Nzc+enb
XgT8YwB8qXZN+I3n92PXKf1edPXYwMhf0QznmrmZwWcMagkykTQvRobYLvJ6Qv+LEJptHy1eullI
n92JgguTtnhDpUoP5UnCqsMd4MvboZaeFffkVzgtJMWPXqriJcu2uBAjpRJE5zLuXLCcZhj8umMV
w5fBZ3whWz3helQLa9DkKBIwIQYX+2wS3YCtdHercBNAH8iHgtuWW7Wum8+fhZgpqAvSYFIPWzze
BsTvX1aqnMPQx7KOzViuWZRZIGBk1K1KkQbXM8U6ysVmdad4vYon7fpruYvVX8qWj7PSdXAYUl2E
NgW3VT346CF2/JcD2tZ2zacMk6EjkppwZDnBOjBajG02scl3ZOhaKJlPRi4MCsxErzLV1Xn26f7m
wepX254ASUtw5PlA4J+Cs1UvbTLiayj7MWUh1SrakAkpI+jk/yvwy8Y4PJAgqpA6nPRU3GoywgQv
Ld5GTf+DkkBEZiSwQ9a+TxJjxRx9aHsHpns77dr39siuHsmzNjiRI+RRYVNWuTqzZHZZySR95r2z
M3vvonc4Cy9EpOmf65mrdukfM89i9eD+TcJMl/igH3AsarJFtcyZgEizxMxKoRuST6nDyweLL4Qk
0WLIVwywzYRGr4YrZ3aF1Gj7OTjp+hy4y04Otq12pMiUTqElaDfIHA1OeO9uyqIJcGPjjf6z0KmG
ISTdYOxddINKQGD0tMk2ybwEHrfzLeKQb38EakfJN3M0d71A1gCr6h9Sp5fApjThVdqNQGJ8itEe
EWUCs2kaRO5IFLXLewGeV5lwMpYSAeudxByQe28BO2XdjDQDsJevB86jeCSoJotBh5PE0NHc7qpJ
0oNd2ub66Z3MJBNH9qdt97A7RYWL384QVzKguc51OroY4+rTqco+i8UGfSYDl2QhBgym++v0CAet
x0dTeSrxriQiLUF1mlroN/i1a9Ci0bVS5srvPPqqcZBW+iY4JhTNbqtuGzcbfgp+rlkp9wiW5N7B
JhkyCtF08DnQnkWhaeFDBWQ3B7sxajI0VPBUxYr00lj+PCmbzmYyhWGGy8aR3DNC/oIgy6OjrLTY
5rm4w25/QUtQ414LxrUdMtBZEfybBfsGgXdEY3F8kR0tYxdvYSZE2GwgClO9wB3IipYd51/uOmQ8
yflAfahFHgdKmxJNq4wb2LGVt4b99UH9IdONinVl1OUUtmcDFIEM3LDPAX1ku0iGj5+esmSClMYN
XpIJ6Zse36Sa8Wp78Y1/kQWnQ+BY7vBQfl0bFDs8VUiC2eDX5mGp/njLcvhDFlN6GgvIcX7y7jCm
ZehDOvSRESsMK3FLlqxyeuwOPJ7coY7F5rr/INvuou+RyjOnCUVTe+dCuyzlU4WsoIW2898XAHG5
f7LKVgGvlL4OnMGyi8xbHRR2JNc7jUFr3q8qGPddL1O65Ra2OchhmOpc6P1ky8AD8F4VMscYZH4z
NYlj5CNAYfEUyAziPJpVq6peZa2DCJbOYth+UCRKArjFSKzKMuGgOj29SD9PZQYvJvU3xwOyUOJz
bvYbj06TGl5P6Ce0HrqdlvnK4yMhMy+A0+5CZtg65n+bkFs8UfiyeLMnj0/soukpn1p3YOnysUJk
swFJNAEP9UCrDkVcAAVcPDN2GVd79TB6G7paT5saJ9enLvlMzMWE2m42O6yCdXjehwI08tN1QHjX
6gAPo06YJQ1xXSD6kJaEJLnQrCKxPnAEKSc0eMOOtJ7wgYWniwQrioJsvI540anoyWjwVl5uMswj
dlVsPM/UAKoQMsxs3IgGQTvmt/iyTptigCLFcwmD3IXA43xj8E2dwpPBm2gDksbvzNLuoz/p1lCx
kXBxK5al+BjyzAlNznTeGww1GuDZwHohfDu/XLMkJ4eJ4fMoQvPM8DzVT/uD8HiQk8YwZL5nSyGC
vvBm96XRgiDhqM1CVFmBBqENzzhulCWTBfgPObjxtrawU3yR5BGjwYPTQQlcVrfZ+rVkceAooFzW
kz9aCdKyMdLbkCI15R/PuGp3xcROJhLX91OfYcPM8skjEDFCG8OaPWSiugu3Ve9bPKEH1uWX4soO
rynAnnGouTNg5vhUTkj6Mrhr59dXfk8Ovpmp/xDUo5M9eFUYRoQcJpLV+3L0tr2mNK9V9zNGDr+P
4oFq+0UvJo1LMI4KOpQYJS7+I1dKpUJ4mcS0F5nAwz/FLZdxoWA7gkz1WZ/2EtPjChQCxQQSJ3Ea
qwyk6GmYC0c09UX0+sR5nPDfKxKW+rGSt1d0V3BJbvuCzs8xsGvpG/0cPkTx1aM6gyhefqB3HFgr
YHxAevCcOWhgq3873AlaAyO0uB3UuChupzxY/whvAYgVUhJ+Imk2ULrwjp4/DD6EyN1RiagyyZ0x
YE1Xb4DhD0eFeu7yqz5zemBzbvz2HPLKOwT5b/XrtjUMrzsr/YUuIctezJk36+pnRywxs4Uuy0Mv
IK9qaJB2yc4zYyQrx3GFucL4L0H692hmO0rn7b+PUegZvzNFGNTtd03/8bYOmuI3xI4X8ouy5FVe
xoI0r5ZTRT2sZftqFhg8FYaJBb6dg5pSRhIbaGRrsoCvfA4qfTyV9SnWd94qkqEABA49q/aljtOA
qOx3BR57Id0xwUXVwcfUWMZ8lUZ9jQLS1zAutzUNKpfY94mnUj3AYuto+fRdAHUx6xUSySzcsxte
FlPlf73IXcJyfexpOw/dI60b+UzfcFQtlwVcyJ+IttjoTw/yWz0O4z6ZRimQolrM5tYa1EKWq3A1
AfCQyUecgxg2un75a4QWkJs/HScLKANJOr62O04GnUal1w3PVXYaU3V49U1L5bronLmP/PZG7El3
BZvutDiGFZnrXXPSuPwXg/Pl9qHoHs1orUlZGPsT2CKxbjV8V5PvKjASXxbH0EueK7jDyE9mohof
KMeKm5iUmSk12ZZSFel8/dC9PHl9cmxrFmhVIKA9w6VwWDk9yLsV3QNrSMh7hnq3OTqmTKYgidFl
iZtC/hP4tdcgPRjNxJaYZYBhcZ2Jz9FjXLTOVzXesyaU8CVmmUi8OjClzlr2GeFTlvGravGzVlvs
fmxMbDJsYLEnR3boK8aE7qwloUsPJolRP18ClUgiY7zAGrpi+bxxmYI9/bEe3/TB6ty2RMd7APo8
YuOIWIuVyrNxsmdKdzRzaRlDwbrHXJNPQo8+xuynuLKZe7an+eK7UKV2ScQq1C2djABBMB48U15H
ud6SPLwuuta82Fav/Ia8ecY6QrGwTGvlJ3VY3q0WbWjohOeMIGxkKuoxswwzskyD5pjYmc2zWa1T
s8R0UF4rHurqNRJwS1/N1vsu/qJYVKx/6W3kmpmNvWncRiU7eAOcFA8YCNpc2lCHYjE68lEhF7Vl
7aP2mqGI1r1vUkCkacT20y0cM5CRpzEqhfDF1NSqZ+YcDINc3AOvuy58Yj8PfvWiY8EyxVsSj0+F
WKAQycfWVUS8pnU6Y3XM84jg40REwGApKbILcx22891v2S9KjRkha5AruOAlCWhujz7Yfurq6Q/C
jrDdYBgqBobpRoKRkSGf8R+unng9WBshyRX3idCOez8Ippc/5MMU+nZckA3+7mtw1rLypIbP4GCu
Ndskj4ngRsh2QHgwKAlwS6Q7hIQMhDZZ/NAUHB8oF2SbHpGd1VzdKWbqL6RhfLv40F/UeVQThKFi
Deq8ObDFWhqGpy4d+difRCA+0I4ybkVUhUo7/gvXpY3ey/zrsrILW2qh3Dvx4cXwxYXv4hmKXLzn
Rtr1q6UsVD4admeykqgV3ZHAiSjBukubtlPfb2dzbXvoKeFYLnSouj0ZiZlZyEjKsrPZxHPj3cnc
qojGxvz6GsuJvXeeIW+9Dzvdnjuoq3NuPXPTRX4qKmUr7KhQKXhVPyi5DFscMJPSml3AV/bQstNN
eGFxklIku025NPRCE6lPoykk32rOXbQJwsX14GtpIqHxivLEgP6Ew2ce57kc07kQaegGD2APQJls
gPx77Rhe8Vd8sv8mnISLlOtsh45pBBSDHc68y4loxN56RTJvkLYdpqM1vX4lua75tTPujYLkHrBz
znHVwf3f9crRyMnn22RxQDzoNa5Vjq2buscbzibDO+AQkuwaBcEeall4G186huqEE4GX32t/KbDo
5pSKB6ao1KmSWt5p+tYmb+ZQBnCp9yTRfp3/liHz8A6UkAEtlOHnNrjQBvLG0/2THrA8Gomw3bmY
0SheFs7dr9k1Q+tyhc8QCa3i20oP2loYMwWirxB7yUPSh7Pr4kx/gpDDr2oXjzuvivKIZZP2kvdj
zAvwsRjCOLEmcabJisCG/ekwqz1IeuOHGQ4d3cG1SCBLEw0DndPc+xA8OLCfOmpVh6whnRikxCyW
gqDclhBpT9WtLYz8/4SmeCKIiEyaJDgypJ9ZbDoaSuJya3vf+OzxBxwCIewDiozWuVX+O/xb/VfQ
XAPMCqsQsBRjFa8nhaLqM7kjG/p99xwRGDqcRssj5su+pFupKlB8kAmj94BzhJ9oBdLv/Uyh/zUi
ok+JO0xs5h1/eAyFAvkvGEGdJaul6aU/7rJtLsgtQY22kVl70+7Ji2rtkzxkbI/h1ya5VoAA76Ba
z9p3tpI5bk4iBu2G4bVxx1DwJ7/CuQdKN/xn8EzHxOqzTnZvqpNo+KoY/Hgb55weqE9GckTPS84o
VUkLaJpSKvURxpRd8dh9jHWkq/SI5Ul5L7rKjLsftSpUvbz0SjqxtZOcOsY5ysf2dvwhDlIbDxC6
uIh3r4SBr0M33e0raLRxjrTX7WJb0xZ6PlKKRCHdxF5ReVyPNo8ubiiScyQFke9ERsPO4V159Ehl
/ErYYcrwDmE+l8FtxfaudyxMDUstUCbqX3rJZbTarbjvNfiw1jdKJoL0fMPb3mGdRPHxlWQvvooQ
3HcgVKIQnRB7/xHH+iWp2OO/WT0Hd0E2BuBJLOecIntrvjzo69WbBc3qwdB15uAdGgr+gQn+bRt4
Axi5AJWB4DfePgmLU9L7JfTIkICypl+cogjE3tuSQ19Jr/mOeb/Ri62zrB7DCacWafiaGq8CZmy/
Ax2h6MopzhbZLiMVaD7xYPxvq/YdR6h+ZYfzElA7GqUgz6KKpFdDZrda2uTFgItrTFMHGTZ7qBlJ
kOolbWSXIhnJ3vkUgu7R0RAcWNVnfYJKC+q5FoZBGGDwAHdNuLaX71b6Ht8Ik/3cNBQyyyFUBxhR
f15nIIkuFNkQYxS2FFWKpP+Na94ygogu6gPbKYHyYDt2WXzMcI8HH8jV3/9onAsLkkuTpRlGdpyA
6BgGuYDPcpdX/o51mqnjQUpleSB6oP1B/X1xMEhZZgsLFcMjgUTfVISK6hQcQHPo70Zdv6ohBRIP
aMu74/aXUrCRsaSrkSjTS+38AYrILhOPcqduUwDopoA2jZDJYGlPyNZBPETGUAVTiEOiECRToG96
+bXk93jMDen/6ZXfKh7TmcnAHE36/6B11N2xDhTE4hRpGcR6EqbLE/rNE7JpGgZg5k8lLTxi3563
1nzr15FuSvs+TuqrMjTVB0eXLIG7Xjja79veSrIcJXgbNoJxLlS1USVFDLrNmxCT5N/7plG3Nk7q
GASuJYHl2YGljHlfZMTOgw55q+BNO1Y6JLr6+LH5FtNabbjmBAAqpQ+yKu7svZxEz5lbrBqGJ0Dy
S+4Stx/iTWdlGdMPAOtc/XHPlfVrDr0dRpYsdfK7hjQVGTjB7EzYmPlUTY6jfbwg1kM+V1DwGz41
OqcBx/cmvcLOhDSsuXpFcwuSm67ZMoWPujqd0cKuQcjUuQujnxDrG+0Ofcr9JiEMKgWrCSvhTBhJ
Z8V5lLsk9wvpyPuriGMCteB5CzKrvs8UJSy/DueK8DJlFu4eTGcjaesDiUyK3x8wsMj0fG+TrtQQ
hNfZxsQztmecCjuKbhdxsJm0hZ8aHOhWxmLmzib75jaGOFywHzIiwrj/jvOY6LlSblDRedYtKcRn
yU46BJeYc2WdM47JQOv+av8/eyGzKSG1/ZzSw3GWCycHCcyZ9QkBDWpac8H+0EvCT+O9J0qend1N
iAsHyTD5e2WJF9TLDF45jXWFkf0XZwM/iR+Iqgck97iRBGq+VdxSWEIY4+ELMfpUCJ1+KIFGeOOy
yHdWmK9VGJD8uYphZHN3uLse5viNO5HNfdaVeN2Z+bwJJq7NGxNMDGKmJJcx867iPf6ZTx2HHWAO
tyNki2+U5eoqTVtnSXa6VQFW6SNZ+HUJQPONYxRm1gHnnCBrHKTbOJ6MZVIrWW1Tw+75RfZujKR4
Eo5vHOoUNBbbtLOt9KZEvvL0yCwdNktGs4k2RWRFU276vxWGAoWVMDNSvsLEMhUnjkmJUyU/DYCA
mpHXp6KcS1jOM5t/MxwzjDVf+t5lI9dOeaRPbTqacz8CuogvF1omaec34PoGWd41nXBAcFczWmMd
TAGwuRktz4jGl+npLoC7MksESUrSxemb3ElWYUJJlALJR9z4j+NGe1kIyqiJOm5R058/JimXrZ9K
Ja2tqlfQIPbcfv/Y9vmQ+hpPJXf2zj1QPcZz4JeaeACjtpIDzEWPTXkjFRJy2vGfs0YXnb3tn6/S
7cAnWAvEpO0upVwVt+eg+mp+1NnhlFBZGxAT5FR2V8/tl2aJT8+3N3ZGBij/vpSRAJjurKs8eYZ7
Z17skfZz3FB9+3MNYTJqofqzxCr2CswysWO8jsYPdMqkrcyB90DprRFJqcfzPcJ4lgO5rZpGeE6a
B/3e8z+IoZK5g2LD6WRhVdOBnFCrK3Q15D6tF7x9ov7v4tzpHidMCI5db83Yx3/ltLieQWDKiWOi
EM1W00+Gv5/YOFPlTb7wX/0RJDSmIxuc+5FLBk9YUUt6ptFvPw6NN7XBZPHFNAPPDLJ/X/awReXS
/EM8Grq5/xWbbjWuEYypRQoMNejWH6gg1xRuNzS5znTMPXs8TUIvYeZoecFydwU/lEo/C9Z+s0HK
FC9T9h21gcEeII3IFtJ3uB2tDhfc7eCtgrZDzrvIQvfaGXljm0wwcyaYmz+Sy0s0CSRHyDhbknD6
0yLTXoGq5yJuD9FmunuE4JyYOQ12snnqq+gBCXaVimLPeW5xvm00aNCtcj6XXT7Wks9TLbZWAOqG
Awsn6YB+YBEMeH8I8L67itHrBaz2r/e7TLLiKB9XaToD3V0Qha+USZWtHNZtz6bzAGmnG6cfFJwd
Ao6TMHRkpdzYdZo48ZFogZP9bzO8OjC/S2npB+e+B5z7g9ZA6coOyAi8CLgvYYDwIXZ3YRzFkZKW
A0DpLQE5n/fzNtRMGuqLZEIgMtOH9rjQjbLRk0ggaGqJg3mE3mj3MYQw9Yyo1c2j8qRSBnCtJIQ4
EUcWUBkS/6QgtpPRKOuy+80bWzxKqR1tdBdmejpFLljBIiMoo7lgdibn7Ta9h/RVFpDHAKQHx44M
vW6LT6hIsuBZ5IZwRX+VmM4UfxEdaaRCK75E+/UDo91ongjmQACwdn3+z0N6eiMw+1yD860NLWXp
I5oUxtoQLoKQyWjF0nHomJL8JPGorBOMinZDZ56KBcX4WoKZGlyL06RM7OKmxCEHgozVu4lV956j
vmU92nMKKoWH+RKzlBvafktTIrc6VFLpURzPrRSaw892fKtz1S3pk0n9TLYd2C1SpvipTyqUBxU6
27Limc8o0CPCl5wxIjVMpF3K2yXGfFP2YBRC76gkvK8gaSDR+7tI8ZtjyYr5QDK1592K5NSeQE/V
xOSEdYagkn0m7J5AQWOcIPDIaNt+YNzxQKMS3F3jVSsYCTatgYriYz2j4x+2gLndY9+KUbiJqECM
pwTjmUXsdIFQNElyxYO3V+4NLbGIF9sqwbvTbE8S1/kVW1VOOBXxswu2mBePmT7aWTgfMwYDqdy/
pNkpbvUCUmdQTDPSQn4sLTv4idOf8eg3PK63Rlrke95GV0rnlC754gGFXYhZoceP0uKkQXUwszSS
fcemPzLYf41sNepfTuS9nA3JTVtXId1GQBRv+v3WqH8NqtXL+lERWkNb05b4WFwEOMBHtiEKMbv3
ItTHaqvYC2AL9R02NJuYl7uE/hrBfUqnc3TsehVW5FLaNU2xD+B7XNSqx/bIc6bJkvrjLMxRM6ui
kNI1eepY/n6L/oeFhBU/CRJZ7fGyateinZIcLE9mt9/tsguaIMn8tcvqU19h+cItyl7YCfM6uGWm
J35oNFl9KEbXRy7GtnTxU1u3J9LJEG8bQwq3Z0UdqLd7t5tmxYgj7bbqXpzDAzq3pJlXIgJgWxHl
B2Da4nwjdXiuwFVqtQLx14g+OmlxnKg9tucaLitW6Zuw0K9RHGJwZXzkOYpSBD0NwsvGqnoN3baA
PihSWfEC1A0PaoLEeunsMgYf/ODvkjkqtTsd7ciO+1Ijm1xsFL2CgxB146hcwxsmjaG0cZ6ebuLx
+bgn1LGFazOZLgkljK2LfN4Uo0M2FLGLYvHlQeTBCwnm1UzCHu0ucaSngDNLGxYGWXMvB+P1OER8
dNqUb1Z3kHJ+YWsIIveiBhWEsCsxYk5cDwkEpXrGQXTDzoUS4BVuGL2T3WguHsGvdGWGR7mnkxNW
JWTQWE9lVv2K7NUz06VKMyK6Sj+jk5wHhF0DDfg/0HP6VBEydbFz3dQfWSOIU8mnPTtiWStGE/vd
8NFvPThcOUS3wfz9aH1fyDU+5TMk5zgzzelS+83VHb1CTyaJROrL/UvV20jXB+aBhU8jA8zYtjqA
4/hjIg1LISgMdQKrtO1nVAiksnfhLF8lwpAIl1y4p/b+Gj9JmocS/ZvcuKCSfGGMq0c0q5/LDwj0
Y1TaxAY2h4KYrcrE4Fydpfxcfj9JVL8lqMRdqnDMqmnhywSRcfuNKHIKWDKMq/pFf3JXhytmE9Oc
NFIgljZSvcNFI4LJa2nMrYZ0mR7FKqNGL3Aod1wXuGwPzQJ2hFarqV2ytQF58m2q5PwBWOYE8yIJ
q0++ccMs1KSnmkNtRG80pdpt8FSBBvN9CYvgvlFLLqmSIXX7oE8tskH5j4SAa7Td+vFrkym8SW2O
EZpBxYev1WjOS4gdsP0hm0amLdiwnhfq7jOvnOiF7vT86Ddn/2sqzm34diMGHO9kKzPDJbkTMico
/5T+mbYfmwpiM/dLgD8Sy+OtPFMsgGD6Wps2idvuxjbyGVL/zGUTwowv3fhZiYYr6em+WXrLPPYZ
GUW3Z3TalsGBVEEw7EH8csj9qRs3QqffhgAvjZ9l7Vv05vS73ttoWoo1eVg4inDIoN3J0Rb9F6Tu
lr+TeKQIxwj5WCV/LQKittwu+6xhszNbfMghZDDDsHRU70JgoB5BZQvEIB7Uh8Co88uad63mj7fZ
GTaOdGscorpxFPk0Uc8Kksj7H9l2nEIZQwZkFaZyax01YkGkLC6w6o9psCMFyRuf5eco0wgTSwwy
M3/ZWHpEFeg4reV1v41WLplSmJlyJni4YwCSsLbSj/lmqDTspePG9dp0q5nPhSoXY68Dj+NfEkJp
ctpePL5Tda0f4o9ILiuLYERrT5Q3hSq47sBa9Gd3cER4n5OQgl7BGn445o8tuq8b5s3j+61hRF+X
Q2bXpODKMBD5Lux9MverpQpwkQWGWFSDa/Nbbs8rwB2Ran+YIUYW76pdtatalqFzGEGr6qEiSql3
zlzPvkZpyspYIB2QCihGR0LQnec2NkEwL2BP1GwH6I1pJN6doranXuN/G/Eog74JJSfGvJTX/8R1
5AOc24FC/zYRaVKfiKYoPr+owMOMgtBKi9eCaubH+9JGT2pK9s7kX3Q2AeWFBNyUti0zRYrCSgFl
6iZeHiAtqf5fcu+XWUntk8Rc9fQQA71gpYAx94c2u1kKcCa6p2AzHrXjEakYbwIa82G3YkAyX2PW
darCpsmHHFRqWg1389VdatuO7SUy0R5HdssD0I8EqU7eRNcZUk3+Bs0IaIfPy+Xrm7ZqVx1CVloo
FErcD/kGe1OVuEQEfVmuk1GBbwZsy36oVxg2lItwmV8jpGXZ9X9TzUQm6PVDM9zt7JZ8IgEqd5Iu
t6IW3x2JjJIXEBc7fOCWJQgSVcmG1g541kiDqvSF91iYaYZWeINYCIYLB+1iIkU+acKDcg+cm/nR
P1jwTN5bk+44qqsCdLdRdWmOGJi5rhEjoXHuZ6pXAvO5CX6U69BdBUDmcwZiEegg91r87Tu5hBcb
tTNADdx4mArlPtRIe78dZGw9I+LEdnFJEhonSIzAkMmtvB9QM3FE/kzsLrbmVE2LcZfGAN6LDIdb
rij7UbYjK7ILGEsG7k9vKaQdVEvCC9jeqr9tK7ukrCBoTNky4UAaWqQ7757tvTaVhtxIQ3ZhqTn5
/qfvvCZCb2KwvcyIvv1RqKuQk9CPUuexSnVc0MlzelN+f5Br9EkrPtb5nPWy8odW/aCSjdb6GI4c
LliRmtc7BL3BAjWSVUy5GeErAH+hxrAWQQil1tevKQ1nTvgX8Q33x88ThEwqfm7guze96kN8WhBo
Wj6P0QFYTHmQYpKTKdIvaPAmk5p8bOJJMvrr2fekYmpGc8UYh1VJvT2k+cxyLmJLevQkFNx3tpy6
/nc91TQuYRzPB+77BtCdNBtHJjZ8nKQX4Kep+UF2HC7q+99CYIZmAQdFTTNp9siQJ9BwvaG55lRT
XiEKyr5fifodY5mogN4xEX0Z2P//4z0Vb2GfE9RtNRAyt3wz9sxYDIqII3erOsGJLMzTXZAsX+Dn
DYOy+NaXYnu1A7X2VFLRDqhModYDy8CEfvUKOCByHsPNqmPWjidRQkK2s6KldgFN4CJtVyEEXEZK
UnsjwfDc5xkLLaKXM2RpstXh5pGVEQ3wkSq01g1LKudNpX58wGRj80P2jiUsw8QAfgjP0ppNm5GO
m3emp4TpdOIUVTqjwbMfxkrIcP1WmYpJAMWw1M1OvBm/IYx3JKnkfV6S3eSaz1oNCjP44ws/WpcP
/fBNl8VPvO1wt8f//sR5BQNApLPauAhHrKbSBIE7icEWTTSmev4xyow3pN15+FZActGUu68HsK8/
9+9ZhzAwaCP5eu2sxX365GT7sc4KpnlRiYrE1yhYliDKxKnD5T2xgDTptlDG4HrrFH9yegFgmZOm
/9DT4amsAS7UQ9eod1OY+JiqzRkqZ7S3ZBo6jEgTp6YD057M0GRSddRn4pLgtWJ/q4wx9a78sMR/
jJadi+/46Yk16io6i6WkHrkZ+iU5cxcUsvlyhx+0d8VTXQhwVMLhnATIdix4X+SC480SmTxhKc3D
+Qz9B1M5j8adgy643hmbTEBfY4ODj16mDtz2EKpUhlAmfAqtd4p72BUjRaTUFFKNgMo2Ea3dBSlv
diIXOqP88Sw0qZLP2xAPTDh8vdYGkT2tYFQNvyuHwvYFLg1g1MmAK/OvcXnp7FEIo0ywU3r5MSMI
sAwQivZx3LYVn5GuKAMQQhvBZtfbh5OtaVQAOdT7gH5Bko/0fTJUS8hsdbu23w2UHbi1WM/RG11F
CJvWf1XO4lw95XC4rC15DYU+y95/0qOzhaZbgBeLuC8uzegwIfv6hDMWGazqimNfYCyxqD/kh1Vb
1qSimxuh1dR805LQdSpa/U8XV90LbY/J8a8V6Sr1wzHhHYjigxH0BlZ/qA2EOOuQiKkU1qaJT5nj
2p7BOFBquMk41TN8roHxAy5JVK6YTciw5WtKk8fRSb4JgW/0ciuPu1eTOQSHEDquByoUWiSP6RrV
+sVMOSTrsQm3uDF8QmsqLD92raWIHEQ16pV8UqMM1hmM145rW/VPEjzgWhqXH+6ABE/ivgSHVStA
c5Ma6QqxwUI7macTT2YZR1rDiDwexyL1MP6fCwE2UL2oclMHkHu/ovgFO+029MXLdKAlUQe91LV3
j7+wiQxChB1LNh8juvxl1QzuOGYId7f4jUp4tkGgDjA=
`protect end_protected
