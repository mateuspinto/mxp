`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
AjcYQ9+24vt2yhnEUYOvDQ8lut23niDY6sum167BBV/r5aBdUxsW8ba/Z274owq1lfK8TE2f/0X6
AUEuR6Hue1dEtnHLTXQS9UyKcFyrnBTDW9JkI/+pdMphCIew8oNY7+hJ61edgBwA8sZIM2mmFRgt
cTrSZSLbl2Ptu0UsnYd9fi58aFwCglBmt/n1QM1l/ZIzUBPGMLnZVePUpNJK/Vk+MzKVlm2Jvcb9
NNIhlY2brrs3Pf5RqS1YUi/EUcpNcwk26+cWDFFpC+VXAvY2ysht9hJYhySjOK0Yz7rPdVgCHb2e
ySfVcNa+LnbgJ/bR15i4Deco6OXhRFqEOfsT4WED4FMkPpn2gEG8/z4Rvcs4dRNVjras9kFQg9f3
CimhyJJq8jq9blpxIXSaAj3HjE/ZDWgIm3HaOjj/zl6tZmn0S4Ca1Yna0z0HRJG3+fTvFrWnfOJ8
+2wSST4lWlvxp1Kp51JXlz0SC0TGtQw/2aRafFhcvrj+Uua6BnIBBB25Oo9gSWRZT56ZKR8o5aV4
raMUK5GsjZGPhZl3xFDrD77lBd7otydUM5SPxb6bf+DmflWw7xTUmV1/50mi0YPhR+DmMZhtdltN
OC4qJTjS/TetlTI+u75XWGhhnoaa6MWk4lw4xf2NyDjaaBaKM7slYYJZDRYNmD5NLggnqR4oRhBN
MrQhm0DFsNopRzsjxiAM6oD59MbOeMqC0v3adZfHCg4n9Vo62rsNqZjIduQsrAMtPboiENKDyjsl
5e15acqfqeHx37TBAWWf3+81Am80J5fZnGS9bwb6rMHnhHaBY6UBYU1NVtIc+uULtCvW6BF5SStw
zysmWrE6Xe2wwa2Dl2LDsM7aXFLO3MVjU+OY6sO+x7xkKW3glC/G4eJ/9j0zWQX2pQlgBaL6TW9V
67/s/qCbSGrZML59yuRvq0Xrc0bbKFKDrAdsNEysaebSaDmFuQcErSKLRv57QDHKwtK5XZg603Xm
TyJ8g0EKYJpDfF5k34+yiPIhslpCmqcspvqD5qRJUvJtW3wSUsLN8wA9GQgDOmXY2+Dez1Nh/XEM
ozytxEMj6EglVLFcgl0lN3eYFCSvrdQ9440ckl7E0nf74ja/S5Xeu+6vL7HzOac75ISpW21DS9wG
ifTDeuHLyCXNT9dQSq9hnepC9zebE3/Y8VvklMF7Hpt9zSeU5QREEAKLQg6k0yeVt2RDTxkP+0E2
SBhZNJJySEY9HY/N5uqrq0TTLVgtlc4rRO7xmyrPCNLGo6mgIvtUEMuS6UfhINUddAVQyU+P2qXO
fNDJ3CSROY9ZbrL423yZQSTUxndWzxyw8pUoKXqo6WgQ/MKRdhFKRtwELpG5ZLZvVB5rN+lNqlJP
qCXmHbk9MTZRtAfp3CVG9/335bFq4Cn42QIknhuIVCMHb/d4/shWj0Gv0K1mpVlCY7cejcDIxV5g
+B2nglf03a6ZrXFRyLfacL2bluTtxCqRnbnKOJZF1JCOLRwLUqQu4covkqcpBf2HO094bzsZKNSh
kuFaErUbMYdtgdzVkvQSVY31KxA0BLC70AvHu3qbKRln1Rv8V6KEKqqp41q+Wrf4zqxsi5bX4XSg
503M/ayNA7RfdMmM7M2Tx6uXc3h2f+rsV+g2OaxWKUsF0IcjyxD32jKlwuEnTv7uMUp5tr0J7IId
FhyID4zAI8PXXQYBa4jSa2F09IjNgsC0VD5V5LuFvRGRYvPih//Hw+WNn1EohgAqd0NTQWDKZayg
DYusMfP+dwdisX0pbfojRmGV1vmc/qnHTCRsJ8DXobEJ+/qEZriUoqwYXlpQCuKo6tuuv54g+7/6
1C2CPvls1+aFxDQB5NG6ojzkmzdo7bKjsozhZDFioz0WqC8tnCDe4PT5644twsaEQQRjUGofx2j4
vCCFN1kdbMWX/k7UReXBWpTguzMF3kYx+97+OFFksyp2UDGjGD2GXTDe0i4EJErWdFlshRBKBTna
DDCAP6lytEqQs4XPAYpqKAuYIgqUf/XSJunISgV5uEXFSrnWtkmrUIElo5BzuxzMqqC0nH3oANvy
4WaKqCe4lyKEP9E4YxKprVILNHM0ckldgLd2sxIuhvKZKv4BgAnhagQ94cr9J8yRTANvhNwuKhyC
CH674T7pWRFH0vARkvuCytbTUG154s7SHQDaDXlA27Be4lp+VpnCiqCQZqppD1qjWm1cF2Kspygm
UmO3D+euixv2+RiDuWM/ViMIWtHj9SbgFk12n90TgMzRI2MavAVMo6OkgCWKGDMMs4xWxkDimq0V
xlhYlbek/Gl4nPUuFzoap0x6fyc0rOvT12qJiwzoT/8azh7jnFwWspevNSsQ2xE4IbGpeGzQR/t1
YdtDDLVYXWh/oXr2zd42QHy87q8I1SSI+XIWWDfy4KLvWTWYlxLuR8QDHVVg3pgE5ZJ+FSiYs2hC
QJgXlQ/DXxHGNak6tp4f3R7tz4+133WadkSDzo9tfjBejwvWaM/l8MrXscEm8glFQvVI7wl2DIso
lhK911P1C1QW80JUGKsuAgmxYMejXoqDt1xGCKN9uQUYilXiIXdarifvj8Iu6e2l3Ve/4aK9c7yd
U3SMNqW7zlvjqmichOnew3AtXvrScXGXRjszSnIX1Oc6BqklWp1rYhn1OcQHaj2smv0WL/gX5vZp
VINVfLVUXkytdVQ0EZhstMfiZ8pZ28A6En2rspWtSWDH0bNi3OH/a7v5mwVrVoqIN+RPxsIU99EC
ss7eFjYFStxshSHZ36sJdTAY+aTfC8mc7rdqGKIsEMaGLx1llarYqSfAVMCGxhcX/xjRd7EamYjX
w4/nIoorX8VLVeEtbc5yOHvAZcRaUqTpDxY4AwIXwmrOUP6H6H9YI+5tE3STslS7j57dbr7ztm5q
tnT8ApesWvkIkPkyvn+iDdaK6rBiiBap83jMF77Z2LgNSekTRqPlocyP7dvGWjjLbctLXssFYlIW
WMwihgzyDBVdW89YjJwgnaw6BPFqsWZDI5dgITmt0RwvRQWsEeRhf6zfMC/yi21SxzH04+iOOMXk
1aDA9jRGU5FHwUC5GaGFPczbcCGPRoiYjcfXTAioADis5OELt97mkVI5Y/48rRbOEAJTYTXbzN8l
eQBDqdXdIbKai7crc0dWc47hsLp97ZwGgtISdyAjrdG7IIslnjF/WFLkST5qL9WR6ukgZdq8CiVe
fK2Az5QXpKH7HnkJYM4sl/0lxkLmIyOkitYB3zl5apRsoPKbIcUuULW6D5h86+PlJ2eOmVwFUZuo
IbLfdeiIKu2uq6j5hweyQA9EEzS7D/aTPHZsby8GdK+riU+oVR10xTDk6jPd98cPZ1BRsJCvxdgd
ys5BA69qRh3mFsrGUrhvABgC26Ei5iIxd4J1F9KBeqsMidLmD8O2Rq+noAkIPmjn4arbXhqIzrkc
blZNfmwQPI2gNaFledvYvhHS1RLjH+JP47rPlQg90zPd7aWtaclB1BsSx/1dQ/x9iHVg9Cnwited
OHw3xc/wpQjOfH2b8mHnuPFHvWsbM6zi5O9/1WBM8CQJ6ylUdD/m+egUCs3svs0xK86zS5UcM8kU
D9CfKs4fA0E7W2N2R+y28gt5PHCENJ+BkevdbKbeUx4nxPx6M0LsLwxXPDCZozedgXrRE4UvzXCN
oUx74Ulat1eTEkQKWep6I7hXWYOfYb79gUDoTZt439MaW8abvwpJtoxMqatSEubavhMwiP4ajaGa
kovY9O16dDk7s23WPEIQGnWD4Z+jRotUlFY6He38xRgVeUs1Se3N/9Y1A+Zv+7MTSzs+HExYvrbr
ssIWnx23tGKzkfkDAdzNONSgF1XtHmm02cbZ9Y65A1utv40+rVlIe3meAGQYMsuOJnZQXImDuiEA
uw9hqF5/kcHDnVorJ4pxxAc8OBefj1Nda+kQq+B71hRv7FMUYptBVgWEwUQZyHXHNfouiQBygSy9
k6Txlr6goRCpkKzbdH46MhbtXxg45MF6tEsKXXohDKCoa9yknaz/Yn/Da1NSa9UsjfAsuCx3SmS+
jgscsNjr+m/NI+YzBjN3Hsnw0NWnGQ0rfUnE0n7NHGYBsE6g16ibLDZ1MiTf63N+5PAZnBGia+ud
jQj1/C6wJcV5S9TKVkv8QHzNgNOSdLY8uvy402/8/7dpBbzX2UfZiZBiDs5O2cYJbSAiIgrBf2s0
WhU1HuTKc3+1pFJhIqhLo42P0elTsVYWodJroQ+nMKwNWuLlXNqrW4pZquYbFHorcF70oWUKZymf
F3KKD5aEO9hCzITLrVPhaNZHg8SoWaKcsEaBNThJAXCk4sel8kGL2EAkyfe3JfJ+yaBhJiEnjGsk
SkgBmXBVacn2d+STvAHs0CE8nVW5h8EHNVIqKQycxosIS0u2wciyCS9bobXkSk5gfxkpxEvyZJiE
fndJMSsKTeTIqPvQJZQ1oHYfXdje53MSBTM7hR6ySPGkexbyl43hsynADisrIB2UqqNO5czyRnZW
IRvQBAFl0HlitoyJdDfVLyajYVIRijf4zIB2ltDH8XkVo2OsK3QF56b5cwOSNd3IDNdqm5jQE07Z
DKOaL9/NuEEGlr6bnIoAdnC0rnQ0W6jxOrZ7BVMJt+3Uh+U0GUSOoyrRIlzAAJSY3/LYtVBDsHRE
CxK9Amq4udYSL4kM6av1+PuRaLdPKZ23Tj441H+20IEX2Bwmz2LAEb23mz7alBP80wr8Y/E1idym
OgBMCMFC0jpuDDEPAk6Fj18+DxOfNRAiHdr2LYvA2Zjv3FG+pTmaGXO3reLR+IGfNKurGHdul7rm
wmuPFA3Z9bj/a632RjhMpZn4689ua72zPAVmFtMAdIHO44krmDNPMF+V3Em4ZPrrO7ChgJaDiiZv
sd0qYaa13tCjhlwrmvUmD8zwgSVV/wuOuO8v8Dy0BWvN4apwG+BhrOYhrcjT2t/JrKGhym1eBrEs
yACBbggICHm+cAMafiSMu9dEH+lATrPgPQhiP4FY6JDu6NN9pAV9w8md0jWnqoXOfJ5jT+iu5El3
wDR2NyjAYIzn5Hn0/erSc3/ns0OSXW5aIA7P905/QsjP9XHcd253Y15+poi/T903v0OMG270snvH
xMKQBkSG1Ftzr6i8m5YHfCN9UuU4lpC0e1dEzm4MXLfz97L9BVCmVqXUQXKAFUYdICR6U7/PJwFf
5JngbsYjztiIhB6v89mA/q27xEeGHZrZAjeqq23ELI/qOqr0xPedahC4/nsL2Ug8t9wqOOzjlVhB
GxMZYvk1/jFlFOfLYWha9Rq3UTNxLzPozCz273ZQ2Rbu76wf/+c2qT2cyVPTCKw0OWfUoWJC+N2Y
HCR90isGzCNfRzzDXFA8PhN6tPj5PmmzR6Fz4aasIGMLyABMwxTC3SI/IbFoeeO5vxm4t39rKBL8
0qye9EbzrDDu9JR8/53LttwxzztFE3lOfzAF5s49IBGYppBO3QW00IItFvLUnw3U4vu0/h/lcNGN
gqH+fRpgBG+tcEsAtrf2KkN1SveqJrKPslyrWqRQKvSAI2YEMz46vxzy3B1/i9qRWcrEYMHWdp0x
Lr1eHyqeuaK0GzGAnR953G/hVwe0XDviBDnNTnN/AsK56I6PSJCIk08qtq3tGq1rEP/XDo/9lCSk
yadfxJXQ/QO+44z0C1HVrj4FHgcfJPLFYLwWItDt8NRupibIr28ZzYZTI5J032kcgS1+kzaPIfd1
pCfqN46HdVmCmHDFMrfS5ixkYBsXpVdSuOW/Guqrdbqb+WRix82EAStWofg+FIwMnG/ZF6ytlZmg
OO9SeblErWxbirHXkQ2wCpCDT+wjnii9lQl8Fn7SGCyxfMrsguyPJ24nSZ0UqS9jkPyPeSxytmrm
1XcRy0+dN+/4QqNNk8BFAWj4xOQRdDg0f5jpU9y1ONZBJNI6OiRRjqFsYbnS1HTzedtkZugZMICc
mAym6jdPbrp6FuSCpDOER3tu1+7JmAdJmAiw00/O7Yr/F/gzjANumS/Ly3ZcbyxNTfDicIdCgaSq
M9HfQf/qni3/sPWANZQr5PEwk4jsxshxVA4i3VUvhOOo3e4PAUHzpzAPp55RApIGQD3g6WaQS8RA
ZNR39c+XnxxYvAbhSum5wwXMrcYW3Io2irLjVHOGvJb4JoWkey08596dGVkqPeL30RYzEjI2jzo+
7FfQrBhRR0muJ73yNkjn204au/rvA97CHn3SmGXrz+14gYAeWG/hagmpXR53ZxO3ZKsL3UrynuJQ
AsK3DnU0NnQX7/z7mH+lqdf5YOAaPsP4nF6+YIO/L66ebzzh84dgcgwv/XZ6pGXNaGJf06dMM89I
V5OlWhTHWV3MHS1fytRchboKUDUDC2mq7qaBXKoQjcAxx1ZH6+BSGRwmMF9tSVVSRKXbaGyIHFm8
PN926THzRHVqtCRtILfQ8PmxgrGXgSbQin40oxoOIlAG3VmXpnMpl/Il5GK8+QtyjtbVJ9VAiwLa
h1zuG6m0LKqavuCmS9LXGCx423a7ti72Eu3+SdFlki7skva7HZxUme6MIgZZVfgq5Bvk3PwirQJ+
GBj1FmlljAPhR/L0UFkEUGJHkEFijhK9Baij7WgYHDvqRNtcfL0qwkGG2OdnzBjiibQqPcVmJbUC
7lQ281iFjoEDyKYw3pdQ9osfIOMdbikoWFuM0u41iT1yasL8VhKFlVIQ4Q92SY4Nfm2YPlBBPy8e
9GiGPoh7FFGNxs1dzMPFJ6MkR8mIk7nqFw5JuJKRybKJUnDMOi0zzVW7FMOp7Le6V0BM9rLNBNDT
HOtlYDjQV4rf5M9Iga3ET7Jf3EiC0VltAzbYHZBdTkteLIzSrzs6CJehftojTb0OCcViqWGz9Wrf
9/WZ1Tm5nB8kPrJXtfWdjgHS/87rXtv6JDMqHkoGFbcvzQkx10dGYb2nMyHnSNA2UgLLK+4m6iuI
c7cLvewn7UAGHb7FxxHaqwfY0WOO3/nIOdKSPPYgm1qvb0g4tMnxsCjJc8kcib+3w8H6rH+bupYs
otXjBkJmGVgEzCv/8aMrrUz1R3LjhPMCqLMgSpC39n5H2v5YJgSTf/5nWpjbPKg6ClTjjil0x0e2
V1HJbP+FCkNDI9eVkJEY2Ex5aER4ls1F+U8Q/dJTqF1yiFTbIryO7tVRcMGFHqmRSgFdhqfBMpd5
uriNG29+e3OgYUKpftkJE4nVLn2nJ/lN29X/Ba2LgJkovSeXxSM4tNCk5bIL1U+BWtsCrBngL8QY
3ZFsglGONJaorgu2bU0RdhHg+Q3MP/oIHzMiM9Pz8VijS2FqgA0GfupzRrVqdQRNXw9Npuu4pSTh
eIg9LqRU3Ghvf7t0DFcvvhleUODTiGjrvQJVx8vOmYg54u07/eLdLClubjkUeEVP3VDJFp0KYXAE
bjrjjJ9GSAP8lCKoEph0aiScSIzdx13s2/NQM6f6cFSjbQXw2qgndDB4RMl75p+rJPgz6a+whEIk
T/1IjoTYAXml9JvBKedIFZoCJJ5e3tONUASYXYRJm3xajtSC4KrkUXZ67iKlEEid/08CCU2UWZEt
fMuNOzkTmzQ1poZCUW9OABCrOBLXPKSZvMHsThdGkTNIaXfqN2EoZaNLiHwTqabPIPElqW1m5krz
+nSiZizHGxsW5c01sI6v+Sft0M1OeWo2EwlmbIKqgxRA+3ecv9faATFBhi4lJX/HtP15ALr3KZo8
LFWLnM6sfGrKWrp/+hlw8np0/2Jt3HgMveeKj3IKgLK4B+x7V6HspshnAA3/kXqcyMjV8afqIqYL
xGd5iQokTGDkPVtUmKbN21jJUu+hAdvYz/FnlNpaMW/RH0/neKhfeWqLX6ndij+BEqHO1O+8d1ND
s6+gxAWdlZN8GtLcdQKb+R3QWZLjLSQ6Caoxesun+9KIRwDPDbDhZiEHFsLpTNP102g9PXeArq8q
7jjqFekUZfL96BMjtVEDJUppAyULm+pziP3iaQJzIOui1NNzyD+PoeRJlei1bi+pXq6PQ++t2Aro
3M9AysWJbrmTngwh+8Gsy6uYUqXg4+rHdEdoSlJvFIt2zydSrxQFIt358pokfbZ6tyJa5h/ubGft
CF9+sAoR+550QML8whuVIysgmeDHLMLTR+YzTm/HDMCXc9NhT9vcAsxth+MryLMkHWAX+8FpIZiT
8bvLza7M7y9KbQb5NTwcrE8bqka3gzRYnRKodfpQdT48Qe1wToflxeVJq6eD3a56c4AptDknZI76
HiM7Xg2MVCyGKW0efcWLllrNw1AUyQ1Leojejt99Y8n4zY6v6ktWVoFssAD9ZnSzz2rLhhqXG34B
qgGqX2YZo1CeMomhePWZIixzhHz7c8LDjI+fLW0mzEoXx6Mef7/JXvbZFwjXyDJY/7bIGHb+Syrv
l/3t0H8bv7geub6Y4NepJgHw5LpZb9FoxZzHMvJ/7FhVOpkqSECmLrEH+XSHgkY6YaPQidLUQSQ5
fKxnG/ASmq+3DsyfCi4uGUYBhVJX6tXDC0P4kkyqbDkbE+28lkEWSPPDAgWnDuuWT+pUpGN9eRS/
NnobRzZjHvKfHD+9FjV/+JDEet9bsmPpaeQZYR874RubAwaYdLa46NL68LAi+Q4sbX0ecKb14qTu
hwdaib42MxquZkwt5Mj1lTWrLlVgvwl8qFmobbFVhDSs4z3LGOhMJnWkzHJU7cNi93K7UulaM+Ya
f5Q+8RNvyvkqOfjqG1+wWNOjzMp+xZf2UItH9ecgzvMyS9dyZxxcbExOneEuNtMFtQHvRaMFFOnn
KC+B8slaPs7Pj/ontz64Ueo34EYsQ7NEhKKBVLifVL0rpXhbGQ3HBxZfhKfSP03n1I5wctXC5hPg
cQ4t1eENYgbmfwb3ZksQ64ea5Z1oG+4VXWsVY7r0s2s9cqjRhdh7qNUU2Tcqy87PDFJ0al000Xft
UhpySEPt9Xurk49Ve16gEIikZp1pMao0oQcobvR8lL1P6rxWHCejAuDTLs9TidtWL1krYLFHijM2
eETA14mF5Tu0E+rSnGlOrMjIXGwtYEICMasDlR8PkPTjZiH0NKWHqf+7By66QwyITbnRT4R7ZO5Z
Z+M7tAEbK5PtsYkzvaDBvEqueXduOr2Lfee3m9Wv+i08mE/6aaMpmPSdJlkBMp985oCaBnOl2kft
CwtJcth+ejoXwRMrguYCoD9opugktaUzndFGj3DVwhjV7MpuscSyoruumGuYzLSDneVTb1jC4z39
ZBVivW5Jyc1m1zSkVS/L+tb46TOEXkyn1aIRqaNq9+wuuUlt7nxclNAa7bP8GFdT+17Y/LBzqTgQ
xDvBjvxVJ1oWm2DvEf7/nFlTng7PZc0MiVoeOqzMIFX2s5HB9BqW5TAslmkHF3I3fMD94Dt0O+iN
yjKNGhqCTbiqX+zf/d5nStLbovenFw0vNOtwKSIeVIEeRRybcZA6S1xjw6GBm5Ucx+KyBsuTtQFD
T15dHybZO48WhwEbEb7jT20IY54zOLD2tciddCfDyDDV4DHyVMrh2qptg/+uaL5ohyhDx3v6m1sf
NXxQImO2C3Gva4I8ykTW43zQz5HliSHGkZwhcKA3CaMNrTvo0C8qZLVq+DpY49TTGxfo/YdDk9tj
vrQm0V0khJgT6Lj7ncGZaPsw/rHAk2uxJnZuHzi0WfFwIS3RKNbHgqdyjG+BXsQ3AT2Ol8sud/Du
5RRZJwH8Oayo1Qj8YQqv0LS0XWzw3cb835rxuiF9UfsDMFVN0QvODoqBw2G4rpoHxb1/lDehi3x4
7xz1n5q/91nlAg0GqHIaoCU2FeBVRIluIb01hZ1tAL67uk7ezYTidG7uNwafsFIGNjemVmOEJ5HJ
aQ6QDrmVwp3sXM0gBX0su8eF7C6WFIv/MpB2kmkVO88ELOXzEAqPN828tMtc9x4gW21Tjwn7r/k4
ZgH6R82AUEGieuNeBPjIGle09adF1E8frEhyTk+tOb8xbTdjbIKXCbNUDg598LaHFfyy5aZM9OtG
EmH2A1t647qPEAmdNxstQUFCnOQx34OHpKjos5BTHyP1Nr+wRPsapUaEXuW2MTLD1njy60cYyMdu
XDAm51AhgTMAGkRP2zh3hpGZjrh54bRA2dmQ0jG5pkbjax99W8PW3CDY3jCUdMN/cXTDH5wPEr66
4KZqOEfKUSQlhsscahpqv68HRoQx7fZ7qSmbIi67nvvG3TzgvlrNDQ2vmFmaZgQDQDxyETOrxpva
X8lU/bVluG1wAEXPr/fVBGp7GpOIdWsvlx62ZaYCRH/VhwTsOVT1JjT1J/VDiWPioAdjtY/8y0Fq
ijg4ESowDEydjZXxApf0ubAhpXgulg69jbLdkm5UMmACLR/bAxhmAYLHBMxZxZREWx1e9aPbKVTS
8nhTR0vll5wNkQEQ5uZxnaOcXhlnKSnbSYUumzLxBizwA6mSK7SIuMsZ81sqQ+bwmg8loXCgLD7F
vKv7qnFUw7iYx63sAINgB2VJzc361aoSl/DpBGsv1W54mzS8rLGf9E1rbHrQzoQ0tmV7iojIHfR4
7AJdtWneZybh1Y/qwUhkeuwicHGL77SWDBiEm3STtdQbiyC43Q8mhxqcNptymf8G9HU0587O40XK
CFpz8yMMx3lRad2yZ9QeUF5f0N1yaY4SgwnPEHgPYvxA5ZfIgrcMhlZnyv+lvRjK9tTsc5U/07E8
IR4JjVMxcPG4uOCj1MZTBnPa1q4Gnkm5TxAogUfeYrIuol7Ww+mZjsn9GCvDoTKS0WuBabk3crGY
IbA9jzVHirpVSqLZr2T2lGBB64Bmo3/xmrD0EvM+MM+y/O4oa2ddHSPgbjUSBYbUp7ysuqSS9VBa
is4YNLxa9gVd4E1qV+lh/QgJCSNT9TUQEHBpNmumjE3mhBRDyc0e6nmi7KLISHHn4XiqnlmwlEO7
EVUq4i3nG43WnbEIY2mnc8MrNMRHzngpYpU0gmDyFtscx9Ng9+8xr3L8zxFF0w2cW57/EKDa5wml
wSbac8KbMBfLHU8MgE7l0+3UlXYsWHTVc7QzDMExzrn9yH8+2NuoZ8YD/hkv6/ndaK5b7lwVolP3
61MTSFsgd9xW9pmL7BxSV49kUKCxi/W50FI2GCf45uhaUPANVfXz0jUdTKYfV+LA036LwudmNUY0
SushCzTa89Xbe4n1nRTX+YTcjpeeUr5S7ZYKBKPs0qSTG1OYnWx4oPR7LpJR6KUPr76cj7sv6Cfw
YCC/rZzxPk0Sr5Ijoe0DhWt43AXpX/kYHrIvGLytAVrwK42EbnN1ZYiHk7V/ltxy4D1RzwUUwvlG
JQn8wlBodKLXnd389nqErh/rH4D34Jqj03h5jolbJ3oIgLJ7C72wCIoMsQ8KhOLs2AGXYqtPkKAd
03dkDd1d21Lar2q374G6ofsvjOneWVzXOTafYvosaLwM4CEDk+Epg3ptF9ywI77sxIBwk5p4Xo1Q
aq1bGg3H2q77fCeqFHMIh+wM6r0jHiESQ12FigUVbs6Kd+TEg3ZDVXwquBngFgxcp0gkIdseoOdE
HSY2Qphg/g2/qnZTiUnToGfV+aShn3Zfwf0Oyykpge/h+gMlcfq7EQoGfUCXQO5RyYEmyqLSv9WS
bMA/JMZvfVbJsfX4vW5vJzm85xDp12LPLUuFEvg/QibLsNbRVcfPShQR3hkfmfx2rJ02HFGFsZzH
moDuZIEjik9kHnyS3d4iGPdJYM5hB1GL43RMNhzm7UqouiSpxXhrcvhpcvkfKg+Qw6XqaWHmW6QI
IaMApcZG4Yc6cHE9tsnhNO14lBpBQqW7A4By8aLHjHeQiaJWJ892EqSPIkWFWg5SEyFCJQx1YWJ7
ZNqL62lO5DEl6QBcId4h65dK42DccMdIiPyXgfiFu8iQEBp/TS55VN2rrp4Js2P/F7Vn0BYCjZ6y
sS1IMDf2tyHVYseqDZqpOTL45/G+Wdy7F6/aj/Lw8Q8Pvhn1it4EZim49xcZXqhNOYH2PL5D/HAD
xd7EkpVU8ulBQvM0QmpA2mRguC5hj6opSFzw+ND3unc1tR/hCXyyUFy1ANcsnPrsTFY0MLCmVEMP
yXD+K1wneShxOQdpHHbQwFoI4E1GLTtjHQylNX/Nf3c++m3gR5jyihR4TSiUP4ulMqSCBHe1O6gF
2Ph0gC1emCMG11MrzxK83/rGDBrhDmHxcr8Yb0adQjwyJad7tu+5MhnWANB+IO8Zp3tZOokH+ehV
Mx0BaMw9It5t6AEXVWMwUMouUrvTvgJDBzI9E+OGIUCTxdfIMxH5k38VVNCKtMRZtj8l5k7ZtbWB
c2/9a3By/EeCJQ7Wr4tI8uuNOwzNBcUm13aw9Xl86uAP/8Kc/T0KdcbXCYRldOFr0y3BuTi8Bdwm
j+rJ2eiSF/NYA+z8XhE63qQ2pdP3W7dsLKgpSrKmsg1d6tu9qT6zbIvrDtCjIDL4L2wCL+EkIv2M
zULqzgV1aBEHXzLsMiYAXSfq0eXZhtpaEVD86jF98LTTxR8AJD3+muO7+fGVmkZpYa3s245YFFUt
fawSWQqFfh8H6YfKwUZ8A9w/HvqU+9yxsYkUp1/Td1z9Zoywa3GoCDoqGxNl/01W2E4jNVdxuF4H
MhHJFBRNuHKuUNcwAwZ4KEbQPiN3WYJOy9xrvlXZYDZyggzE9dyDybAVhGblX1iVqrWrelveEYtK
m9pD2uhq7DmSXn9tUXAYtJPhMHf2W9Fv66Z4cSeTp+LWCEFA92nRlUz1P8TdcwcFZErYTf/16G4A
6iMOfQ8M9+qz/W5kETlzv/xVzuZFILjIJzXS4nhkC6A1vUq01ndHYphgdXCPfkZ3EFQ18JwP6rEE
dVKjCQK3uw9ZtAJ/4KOz3VOPvtU/bNRHfawEq8gMo7r2vhSpDRnXltxN5G7NIkRWCWUhLoDP3LXY
puXWRasPv9quDrrDeTQWQ7yaoG0LqR2keoZEnJwCzbBt2qHZZtUvjAL/BsS7ahAUEkqAm3YXwtez
Ls4aHs0SLKFCIrcCCQNLLIYLTLXt73tqlGV28BLssstT/xmgzqrOr3kn7h1nI73pJ5qj4lfT2Aum
zavzA68oajFnrCWday4UIV7dIFM6AZ1HuNB6Y/LNlSFz8N5G4HVcQy1O5D3sqtmmvME3Hhfb8B5V
CI/gjj3JsQaqSnJRkKBSX8kWv6MK3bHaEEBysJqZJe91pu8UDJMZQQdbXzXTjjextt3TpVDtQjTY
DQmKVKQz3xO5SZcNUGW9E7k5VEMfCzGYI6SwUHeQe4jqQdtHD28gf6uz/gv37ubkSovOLqciPGpp
MnIFNNriNSOfjjTm410AuU0uJKDRCN2OD6kx6Yj9y1CjjH8KzrBPpmhFP1RG9t7O+vk7QKsV/7MP
mDu1wt5jj+4HeQb9+UwY7Xln1cyT6IliYZGYo0hMS6SuQznwHPLB3J/xjcRGEzwrG+lCPguH7w1m
gvFqXT7IoqNFPoFOJZeSyGObJxSiAriq7NY/HLDzSSI4tne4qih2Ce4yG2G506wEsPs6GCaR0s/X
vaxVaxAKYKMbM/cMnjrFPND2X9THkQ+NVXdgBoImtK5rLTU1StLF2BqX5cayTGx16uo4ogN10HiJ
+EWT+1x1o4Ar9RnXCRmG0CP/4AVCTquAokWy+ndHDDn6nJD2qwe18VSuRFGQvfYDz4JcQTtEVdXQ
7JLeUw3r8WO8aJP8GmPd5c9sPDeFExs7H21vrN+HLJcilI8GeLKVw1VbysohLnVaWxYPTvgFfr2o
Ke7f2f+J/jjYBt1GGIKx26o7DYWmvLGWC3KZUkCpL8v2XGjSGeAidVGWXbEnch9TNt6Uzu9Fzb66
jKqaOirNKzavHRRGYml05w21HCEC3KLJL17KkpeKpFa0ppmdkXrKGX5+MVJJi/w1TyVj/xk/FaJ0
EYo4PZvEJlzZV3NJTnR3G1CcV8rE6TtvuvVhcJ5OAcP5d9u8wZmJbeSP8zDXn/mjtPMKSf/hgloK
IipyYNpCX4VdF4LoFugRwECG29t7/nCGVpTbsfDTdDDOqNQbBMQdikmEM2s2e0w4jwqOkbMzlNQ+
SDbt9GS0s/1IFGUKWj/mjaYj2RONSalCwE4x3HdGQVAGsd8MzSauDY5SczE3bLjycWTL/RGyla8B
HoyiBOnQTGH+uzmolqKszXCk19hBikNhz7TAhX1molHLMSVeCPeVYz4eGGsdLFcOfroGro0AC16t
cqslld5LVjfDiD3Nr1Vf4taEB0JZfeETcr+5/wjcYV1Nt+8iScYwEZV3RqaP5eeoLEa+vDLXUqwY
EWvKHeYk6W2jFPVjKaQzGX9Kz5s1wrx8ceLXFWKa/YEs1NsAIkWvn3sZAV8RxDStKFg9wRHk4lWC
CoSU+PYHMsLxvadgZixiZh8XkEUeAtyd+x4+Y+Nn27v9x7J8wXBY9hHNUyewtKxU09evwbToq5wZ
TYEQVKgK+MN42w82g4azIRYZx0Fcx47aTWRizIbumHTURKusJozw48l4C/WJR/oJzLaGnpURoA2A
weKEojx/UCZ22m862NWcccVqEnVNzf2YGP+MpDaAWaH2c35muAaL4ZWcu+sELtXV6/ShD7bSBxDG
SH9eTQcFJ5mqT2GNDKal8cFqp/oH53tDFbtxUahF4Bk3jkSnarKzzxSsWaARATaqOxVjm49/JC4q
0lZPEBpMagBVyvJLiKnpZqFzVYufPikJseX5KsZRIAa6D2+4LeK0D1fWzg8axBawT8fMghIFeTRv
HNYE1/vHoNUGgS7dMXRu9zJ6UNlPSvXeNDxmROYnrC+7sK4RVDwHpg78vyKHNkSVqcBpRwFJDh+y
ed5C4Gs4933vEMUpusqhJu2/X2gBcNCqBfoRbTYjKHUo+/zogpKBDurFgFGAVvEoWEJLg/z1WT5A
/eHWycPishwrTw5f+FGQh7Lp7B8ByBeBzV7UYAp0pnquZ1OxlrF/slTnIWG8w1LayDpiyhRflzTF
rNEBbYn2k37BswQG7TxnC5IfXws+5bs5+ZU/JZwM24IA67wnwUA3KTEQcZkYOvmP9cUMmWaeaSoh
mXlq+KjaldqEvmmmId0wTdqoSW8u5LF1ES0ewA6fNWztgk+KHZQ+rP5YUEonaUQFgzd81qj4GvKf
xCvgiwkQnvAYDTbX3NyUCgSkrUu7u54wLBQ8H3X4SPq40IC3ynNZykmJOLKZ/bRE2FFOYJ34XhnO
kkc1IQ5jdrfTUNbPmQph4gigCQbVaer+964//HDITawBVxp4lUPMr6xayu65KE/Rfs1cXas5E3M8
btveeJPFKp5YTUUc/H93zT59yjXmkvwA0uS3jYNSZI/8zyAjj7vzf3BDZoIp7QYWdnfsgVWrPCeC
i+i4t0noi7HwAKJkdzr3AhSW0IOWp+eLJ9yU1nxR2wQRCe46V6LSKxj5hCjU+s8HVNgwaCq9/s+C
xgpouYPaCzx20zj2XnEpXR9sh4ZViROcEiD7aaKFHtMya962zWjN65rAphBJT+C+PEM9vEEt8SGZ
M2CuhWCphUFFWA03EQQ73KxZWHz2p5bn3WUhPHIFJkqRl0+VsBerDfXicgntzw8boCHzPXqv+cTs
aSkQVpR17UP5pv96lhWrD4G6+WQuhuhX8WAgUTLoSzzvJ4IUWeVxohX0B3WFvxOFgavFAe+77HBQ
QQp7Og+2CDxFQfeyPYz/0Bj67P2NQ5sxd8aNLH3fRpn1oCbamV768ZWUng3W1cDTsKi+Jo02hA6N
shHIMz/NPcKZnaQM7RHtwPuEdfMd4kOAjT3tUxUlh5sRcKdLQUXD1YU5KX3DJjk+/oCvjVUCGm1k
nWfrX7u5cLJKreYHLTvccE0udcBwo/XH+T61lcsg1rxsJjniZCOGbCVEThMPvQaK+A7ZSB5pElb8
WCp4eRJV8tv49ZbVJd2RXRzuQP4ezW15j5bgD2JMcXUgy4WP+8svwLCp2NkkiaJvcX8jwjuueHcz
Ymd6Zmzz5R7HbU8WEbNceyF7Prozk7g8JbpSUNqDE4FDJakFgBr1vvD8XCCPaQxDPHHPjmpyjMmN
kakoX5Mpvv8GCweHzopqfMRymdOvmbEX4Gvxe5prFJfnoa54rpyMbjN5RqCk7Br5huUG/bnNPD9w
UW8LUp1G6woBFq2Ue8iBOVA1ZnGwuAiVgLA3kWyJMhaOkoKvngYGUdaS0yuF4kVtjooiJLmyeGNo
nQZFoUexG62XiJSfvzaSh3PxNUiE5YL8sXFshhA14x+GVqui+sOGdHFnbI2/MDuYhpT2UlVBIrRL
R4aiBmn56pmALQnPLrqaVzrZqI6HFFEsLIT5+cJr59ybBI+EQGf0JwI4KQ5c8n1A1nusUmcryFCf
IbQ3ZhZuD0mIJSONj0KyfTCkObsgNfuHxxyDPJtH4uAitZOxcKodiCnPPxivm0GIKUkLdnyIVavm
EF82azYLCoz0UyHYKKjAYHeL6KIBB0UpriF++tBi33MilQRF6sLpf1lwK+kSnYpEWS9rD1Mtd3Fg
RrmWZ7Im6SHZdIrbpv9aZ+Kf6yE4HZPFNfmXkPtWLUujFJSTDlTh6sdjoTxgW+uPz69eIgt8lx2F
8weQvwAD8ypSFdGhw82kxUMqAy8QUTnyNKG43HWNlnPnM+OLwDesfSht2fIteg0KWvuKKJMHVVHM
JoZWRaG3ylyrePFPiVNb2dWEmwfb12pCSNyhX0Vyz35luYMkjhYHTdfuJpfZP5hyh1zNdOQOCrxM
fFMglC6tLfuR4/XN6YGxojcC6cigC7vFRf7HzwYM5QNdd3RjHpJObp/s14ZRUumPxUDfAx+L7HWO
UYOv76hzCg2ekBxnwJEw7cSU+ItR4rwY31TyXGCpiMJrTjNeZ1kFTwYiLqh2C7+8/HzV9ohS9q6i
jsLJaT1NCnYkII9ftTg4DhsH/JgyALs9LpZ/yQEvIpMHuiWsq0ID6gPYlOnCowbiSmaUegB6o+Mt
ES7aDowmJGVW7XvAaDNV9G7MaDdpxJr9oRva3I/r3fTEuoFxYTLn+HpdknneL78+5c5cZZSSqrx9
26xFy6/jq+uHTL/PZcBtccWzHjd6wl5VjhFJDHfjMFdps7yh241lFNTuu7n3hTN1Ff1nWOU6Ye+D
4PggKHux3lkZd3wh0hj9YgzePT7eksqXfEuKiGNSduyTG0+/5KI43urOdkG53bcxEWGB3FQTgZZe
uLOSLq9kI1FVxPoBLnor4q+YT5fttVnXT/ApecqB91ETxGnCLjAEGJ3lf+DcQ/WTcnFBJ0NkjGIT
AKRH2JjAGWgmUBi8Mna/mNvYfD6h0i8Gy9K2EXI4Hqge04nGBy3AAmkVA2d18/C2pF7TYHfnuydl
IA+4k+8D//PFXgNyOZGdqvgGFrldwCpFpQD7iHbwUyarWeOqyb3iO2b/Fu0FJJ7+JTN2yjJrq368
hAHbrHrUcxY09WUAAQxbnGBYZkMVUd/SSgX4zhz1AUc93Lbm43hnHkpTPAPv7REi4WYtV9JD718L
kk/NGMhrEgsvvcipcIg3m+Obm9s5GHhY7uvK/2fp7Y2X2gtKnp1ymyypTpDDPVxQ2/GvQOVCwp9T
HRIgpC1M9jdZJI0oS/hazLeLPNgjhs3aqvH5eNjZ/dadF5xv0a7eNFIP3LgoRg/xgp/sAefYMzKP
johtNgBd8FWkNpNofQt7XI9yLK6irsoowageas5GHL8Kkb/9wkAygoCkyjX0MsDmi/AAe8uZ2ifP
ux9CPGmIQ5l8U/Mtou/a/peCff85zfMzhuCqAosBRbtTvXEwguNCgtZmOCFXnc3CVCSOjxSDXRbG
Ma/skU2TpMHfq6tTDuuLDenu4fhkoc+afDQRyH2rzQFOF4EPsiox5SeHtI7i+lO6Rfw057nPB10Z
9xAQhM2E8XVmu5FsbvN2WwSRCd0837/d+bjCNgzBfuPUM0qrjxnGA4+wsDCOymk7rAW2b5P9Ngaa
95isPyekTkE70THLKY8LTnVPlJ6XWBn/ULmn98CgT7KhzPbKjAI+8Wxha4ZaqGs+wkkuj4t0umHG
tfNySY/KtNEZn5y9LXbGlnhwZTiINx5fK7EWZSaIFUvdJF9cAweA2vbJ4HG8Me7qZsJ3mQTILJXP
q+zYMDzyVAhAvJrSDzKS0130Ld2YFLOoLfTRUCpf7YHqy1sGh1UBKL3hPsfFhi3R1duhmaIsYtG9
wQBZeolldSrCG5DA3RlLEjQzYRHeO39ExCMfp+OKbDW/bg+YmvUkVz0gQbb6Se4W00p2dkTcKo53
RTOLNgHbnNGN6AfQOkmLKgtcrkbqUjP6b707+PFETFj2EGaj9M0IijZl36F504ajXwopnioI6R73
zf2tEqR678V/FCvZ/2SHL48MdYvpIbtzziYJFjnxvemOBCCf0qiik4csrzp61KQ4h+M14YYG8xeW
vCe1rU/+YEYkg4r0HX0xWp0vc8h8c+OCDoeP5I/OzMOBbb/u9Z5aXgNSXingz6HWnAUbW48aPs+7
oXMOajrnV62kyYWfHrkOqMpB2LStFBWbWjYTdPoQVCr5dCUX4GB6HPutuKPUkd1iM74jWRbONp9z
OqPK/eu9jGNzOs76tuwcitlH1jtSxKSIHDCiONw1ZANOLtrNSfOnRg/VT5b9Z/eet2vQwk/cn7CB
qxhNSJg7b6frKAwCSOxIhgPQqEEBpXE6n/47Wrcm/HNV59SXSAg0EJmK5zhEU6o8ISClEpmoYLwJ
Phkk0dHpnN2ZSRXEwp0yGSpDGUYUbjVKY4ehYnzMs5yFHo8H/7I5hwTukGMaANUVIPjWFLxZ/mtz
vzAvnGOTGQemddxYrW8F58UBLaTFLvkSl2ZETTYb2yhZWF8VKLDyZLta5Ij2Q/M3FWFIYw+daD0c
tOfaugGopWDC5/WrLN2f4P++opCC0CGT4+KLVLk8pzikCbwpRzFs2mGIh30gnxmkJLK4gH3af6lk
7oi1znBnyFnU6QRpTdAG/5zv8NiO6H7eP9kQwJh6ZM5x9uhWNUWqKxfZwe+ByQmIymTGQZEHBF1l
Qn/OgWG5vc4TFnDEQRcHkJH9s/S+toc15W7Y2qOwOxQmEDXS44GZ/UbvchUxe4UxlAnRYm0v42y0
eq1vpvxHI6x7gNxeJtYWsFu7tmFgt9FqwU0JYVQiK3X7y0PgR2vCOumeyGCPGxtvTUzgPluWfcRq
iPmY9R9AByJZPRkwxgCT/XuI3W91I9PRUKR62Fhqu7cz4RpgsGotQ+1cJszHOfgmESFzJqd3cTVG
he56dBVnhlKVFhYA8PDS7/yP0f1yrZpsAxjqY2kLOwGESnQLCHy22cZcSinfBUKRE7jztIawE56P
G2Gk7wA7DDqR7fjfS+hyGwVFR+B/yYgi8IJ1x6nH36gZbqtxz3i7PcwbrjaYYKPPO94xWhYwWEw/
RK2LV506kXUqfDEShyN8LGUHDRM8jfnWocQ4VCdb0XbICQPAWNIggmhP0nkYFyitdL5V5n0948Fs
QeqqG2BrZfoa56NTYSFIw06nG8VWqJ1lAHKl8bH+6X1H8KExeb/9JKTeit5pPI5PyRyiu5wVduMg
Gu50vwMK+zGyzuaQuhnT/QrIgBVKBLhusVCYVOAKl0SmwqbCo8bXhwNJUSlmQp1E32etBGsewRBs
Agumo56i2645WD6noiHmtcvrtr+qZAsYWpX9jv2T9jiiFm1NPMJ2BClxawNW1uFCHb4iUDOn9JT5
plP9tMc2TgPP8R7IHlsfZH88VZYz99FpFrPNZROHw8Zac38V+OcEW+aeAdC5pu0pRzGkuc1Jk1dg
KAL47XmQ3qhI4V+1xrsUSAgISVvDnH+otBp+xZ86WblyGUN0dvqnE78hkCFpJKe8hxBNYl0YpsPK
GcRkPnlwzFQtyj1fV4w3fl/Uy3D10WFvwcmcJk6rHqD4DiI05o93UwBljJq0v9O1ZJC8pY2rcSmh
toQ0NvAPYBY2zGLSPBP1hCyYCHFTPHHyfcI11MgzkK3aSyPdNJI4AufCS1i/b75x4OWtAGLq35Xc
V62SNgt7b068c70VOdz+jcercMW866KEWzSpYdOqKCJz26dLDhcPh/RIJrLKL8NzdAGIzmowlj3W
RjUuEpSHcMA/+WcBLYJMUDwc/07LN0FFy2JWMmRL8PmCKrltx6sgQSlofSUc9Mlms0ZzOEB/zyRW
T5Kh7aeq8y7thTLhsb41Hm/5ZrbdGHAdILnowG1gFB210XqI8Jpdrz5kYsKjM46iUBZsB7XMcM89
Wj4P3mKG/cQy3og9uIxK1bUdIt9IokMMKdKzZ+qAcJssUPbAI8XEaqXCZ1Xy02dM3Gm9kNMZw8R+
m2veMHMUSwwGH9rdJ52uoCgp+LMNVdqe7CQrrPfTdtPsjXDCAD7ELQTRMvGk/d+kK37Ngw1ZwaLX
KbmqpUBXhbd4BdVT+nFHK5QMSuqkgMgj2BnqERtbVcKt+T2mBoOtPmTbgrAvTfZPi/zBgRlfjRO8
2FrI4lfgeEGspCCXbPa0NsTG0ro7pFFmV+m12uqwJTC+mN3TyE9AuUqBhrQv31QHm3Wv68zsDSW2
1Xq3vYIfryC7Q2R7L6mjd+8N5fGfCsXMeLYf+ktQxq49y4LlpFMH7KieTGq2o/XQ/kLqrsBqHQ+O
urKX84qXgseheYkbxxsm+8da+fvM+/qK42vAZJtQ3u6SA6ZEnO3ZLn7pjHdzMkvARUdERtS5EfDS
OPCNXHB99wuDei+rEHCktogO7VyDfqZoICMb5zubMhBApaNnlXPz3hZoeeDHi4AL8BgQHOXfOWay
73aAhpOQ1jOnuXUpvtw/po8r3eE1Pjlnz2qI6rXsju6EDCXWnvWr4PZL+LmaNlXva4CZUcBa0GK8
e2+UXN7dIbNHEeuKLWcEThUYluK3aEEOp22ZUlz/noOJpErOmTHA7pmLYDn2Q5G2stkQ94YpOn58
LscecYURW7epNmrqGoRThuwZt26WUmcoAAmE3LA+PGMH7Rc3PTx0UUP8CgAVMvmmALVRVEAkhvCI
RjcTZb7hthiTGo/ChVs7Qe26A4WsfuAhYNnmqIvNV9hyQJ2C4VJb8xjxjau/slMmTVGQJPS52OXd
y8Kdur87uGLaEte2AioJcmOnA46EyL5cQikUZaSODeEU9q9Fmc9GnGg+uPZ6D16gv6rrxrH1FdG7
PKsGKM4BHfZjrpL2pVezz/3HYw1lb/nshP2fNgc+MVOEQJboMMkE35GMD7CU+/TCgPuVkLOvq/35
qHw/gkDN8DlAHeu9OD88zfLooNKERIPNs8LITQWNXdCs1KLCKsCCHfYc+o2ApDEruGBHmqk6Nwu8
1bUQ+6dDwYrIt/4YcaRpPQNET8yiH3qVOxbR3s2uxe5uDuqNXIlSEKK+gbtvT6Ip/qpXasTZBbOt
bzt5TGkM4CvjQitOJRJ6205EX/v3UwYuTmaEF8uJS3WSBykikLNWwKnZJQk2HRrOcGklkpM6o25z
Bd/rrKqn3DWwlKDMRLwwUV1lFOl94uAFzoHWOdEptjOdAtQvx6xCABy8l8n+rDGvCVxJ3fXE2T0C
gVcZ771HmsqpyNWXX8zp1seS9Ki4ARCWCD+d8Pyw9pjo1g1ChGZrgL5WdeahL8MT9EiO3XlwqIkK
JBv9dW4hCi5jN+I5P1TzLvEyksjATZbsns0qE9UfgXEGCjUbqogHRwGogvvwqSe1ZDzXxKNzTE63
AyzbYPXyvqm/OR2GPzDD3fi9gdxLAm2LEnhc6kah3V9X+msH4euk9coy6BbrB0xz2DskxQ9BwEWO
fa3bTks2GRSmEPGEllk3YAqi5qOxLxLufveXzG/+X0qoIhsA+A1dJ3V2xfsTJ27yNBkl8lg+ENrk
8f7LDvUxEbJY5KrOZONvrj3L3rHbsR+hJQNaq1b0gOni9fuEsBfbjwv24xAf3huGS4kVDO6fw9N0
jWtVo6uYY7gAPljHUzrKuFOeHr6QaUZuDbqhVPEeeNoAZawQ2R+q7IDDfxTtkDcjBSagq5c4qNym
ve+EZGDyOhkI20GvxfPMwqXtQajccPlHxUjOLC5N1YITZTy4OdPCYyx+6aJYkjVsG+B01mOjcGSY
NBJpIAFuiQ2PKEST7+rHmGjgvh+od+1Al0csMtMKhn3VGpkzBtmSnHRzATeSmzE3JbIlRzazY6mG
fd06mdh8DTk2/lHVWRFJv3G89KmxJ6Yu/qtdO/vnP66RjzbjayDbSvs6/kRvfhPTdRTsRL5AFbqa
NR/i5fIEzvg3P09t8uuEP6bqwzUpKgvdswqZELeYsjosLMuOlFLOSU5zYPC8XVWeuu3GQY2Z6+xX
JmxkhWMBqH3WgUiQg+TNsGaLx+WSakxoujJAKYpdPAyMHgqZqTBNCM6jce9+sBsp6ntufhV5YKZe
70QAXUqcosMM1s823WHbtia6cdDYpGN930tiBKGcF3h2Nmj/1yPC/NIiXrfnfUVWnhl8jjiWOGIT
Fw7cY5RrCgXUuG6yeGVWsOjGRLlWq45oYptIInOteccIPj1rfA/icJIHjIintYJfXhK0MK9NZfsE
dvMlHxJyVzOW6bx3TF84+g4E9wey6V+Jh5eyulXidOoRnuu8eAGNHFk7ZKXmsyJs7whQwP7etK5y
WQNbNsG/Kcl5UL7jIzmLKleJifM6ebF/OozSIAAacfDyYjApXgj/bKtyBiJKFtYBF4WJV4d5TOXx
Lw4oX2ZvvsgE6Pws6XVe+WpM7Km4O/nFRcUdXMLXWxbfhiXadnCuEnFEHxgQ2THch4TuX34aY7hy
GPVNArfxnoF/i1t2eUbc8/5dWz+L+IPJCuqEdI2AdbC27n/K5wMSxX7NYAHVxqrUxUqxFKdvNS/V
Iq7sN/TRna9qzEyvf0J79MY892fIPXCTjnAbwgDolQLEPUdiiSdQOtlhx67fjPJx0eGoPb4lzehd
06YFUxuN2mG6x8QIrievA0kYezGZF2irctJBEoabJaX7sd8KIDIPqIs7+M1EmJCNGH56cU2DoOKc
ufM23KDJX1D7lZOu0qbQxCRdtZMIvrGEJnat/CVpBYnC3YgNc/wPx5ZMrHTKmPXt3wMsZjsx5umx
F/vRBQQv67WLnKTlnNErtR1JL1EjdBJEgK6Ifkx+OUgaDKAaEK075MbO8yBrH3nQrSZla/JloCdI
qU5CWiUuv43tBYiIfN4nvkrTPo1XXjMceVTzuHSkrIj3PU+3vQQ/VcnQatlo6LusG97Wb9Yl4RiB
11VxIU4/rbT/2fJ1iQlARNIrhsdZ0jZ6XfBlj21t1xp4YuS3yINf3HuKR/Ax11PLHa8Kfv5f52Ze
gVxnqyfBHSxXlri2bPmcorCAe+M5mAfCJ+puFySZbe+Pajlz6dFWmxTn1gw2o0cmS/lsljRSRW4C
167hvq4MgvQzuXL++pnZcJxv3ovRz7rwzdvJMcjF
`protect end_protected
