`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
nW53WFS9E30sz3Kp/SGdukU27NngHG6lXiJ+zyVMl6AdyTFPC8hy5gHaanJ5nDA8XjbmkK6kXix2
bOnzY1sbCtn5xq/e1Ds/RMm2WbYIZpLsLSDmxQ0KWdPnOvGI/i/KrvTBpbALPHc+qG+vZ0Mq7wlY
yC2XSE8UuWCetA3+ihA81Ak1X/AuLKPxbRi8i5O43marcktrI6XZVLx/Z4hUl43zAYUsqp+1ijV/
7JUBRgYyOZT+ip4N+OaIgxvbWenhKbrUYqgg8MR3PS8KgDgRUwHCnYH3Ld5xj6y7Et8dyldYMNQZ
3DuuPpY5jdSEXwQXhURqae9H03U0x/0hUuiQXlfFTTBeu8d1/HD7Cu11SuoUnNPTwct+CWS7wIlU
cmRGHaGTdtDfn6ZfP0vc2icmLQt1jck8G/iDhO2sm/Zv6AxhaPJn+OJyHzOhnQ4fTIctWCt1Lx0/
dJYCl5oCA5Nu3M5rBXUeQ0ZT99AmAZSnVQ1woGqqwEQ97iuYVsV19wqA7opvHG5Lf4T4lV5vFHV4
lkWH3EVNkYCnblB09iTuP+ILmlq4m3Ob68JJY39EgsD/lQ5Zdi7VUYSofDm8AMPmGzLj0BKXyG4H
zVo93XSEEZVqt1qS2aeXy2XX5vz/hachtOTQ+r4Qud5SmDSS5J2DusxKR/18zfQzRgI5Muu1pMkV
V48+3Wbc9uJ7yU0QuwRce6pPQiBG1SIWUqOU9vUs92TEutPcM2ZCq1uwrPOuH2saSbaJUsuxJ+6r
UatCNYyZI89wahrJi20wEy396dm41WxTxoSz0DWWFc+hRc4fimuX4ZIFMqryrpTVyesLn3iwdn+9
oo460hg61bIe5ecW0PTT1dPahbRtcg402eIflGoHsfWDk55DJIgVONk77CO14+gWcAutKl6yt7TS
2jPPrnFe5iULYo6eUxngO2ybh4xTEWRT3ltxrjuHyLa8SaM+Ib2b5Szq5Efmm6y/eKBaXzWgYQJQ
PIDupIf0jBNww7Gbw/bdo1yKJUn1C+woVs35Lnrd5svzgaYchnX86qF/d+xWwUAjIwVtFy53sqfX
ptp6DXTSXDbqn7agjME3LukP2Ik1QEcINVikjpOOBQF0lah8QxGBffIz63DXohHiGVSocU9dpYNy
v+T7giofZ31ZFPHug4QsNFcfnkRFxvHHpoqtFasNvwSHrgas2bMWgTn1u/bMxDzi/ntkUhtR2SSL
bC5ecAsT6OvT3FGmDAYjtocZWr8wRHvF8XifthuGN6KuzBV0k3PZf04atyYhzjAVQhWXy982pbPA
Rj4BixZZ3rOrmNtw3nedO1UKJfAoKOv9+Uw9ToiULdRR8VW91m8IzHPrX10O/ifoEpn2OyJyaQ7V
TufmKcq62J7l8oOEW4+/fRXlaehBWO2cJbAR7SYIJ2EXGM8+3BnKNHvFeIEUeT5kUGD2e1xsKIRj
5yOhmRMKL1VBftfiZ2kwt+a2LtQ9DoPyf0mFZlrLICL3+/hWkcBqeENE4960yiMrfObELmHDlM+O
d6Z1a4zzJIiL2zJ5Pa4l0CkUSOplX68V1dUDroLO8Jxv8O1lPiiU/oSGdY1P+5g0QglH68ZjHUL0
AfV8Y2bda9Ugbb7HE6lZ9ZFmTU6TmZwFJMBRccQlo9YeSE1rKu+mIbzt+r8JsOoahYzJXee72XzF
uDOoUxVhd8A+qdTqrOD6WnW3KMtpbqfhsKDYXcwMg8pIE6D1wJABv5KZXVODGT1UhJwkpc7VEZNp
LElF2MvWOaNqvnT+06N+sb5mOYC0tldX0cz8cNvWxdxw57mGk4l/juVs7fK6jQlCVKwyvmrdAF3J
tFZIGFBV7e1J+/1fA8YSb37jpV1eOGUbNqXIxgowST9a/8zTHv0DpZx7wbi0QA1pd33qQOPcAJUM
lgF1zxxQfvdFjgftiw9J3HK3LvWfIV3v5KRoIOhFwluwE2WGSJnk1N/8hTaZOtJJOFBYHx29Kmjz
vp8zNYTZ/I/C4hSnkjYXqJDCG3InMlGOHIRo2n+Bf9MTAm5ve3qF+3OQB9ajEpciyy1IXvij6cDh
Yw54Y1kq7buqCLehhY8noPAp1i3GexwC3uQPQGhWQ3+gC6y+ywgVR0bGLIG+DVaMemt805N7uh/4
iK+YpCglBxwQDo3+b+bkiq/DeqrNaz2VGtAkqnTa98PYvRPH3O4ePyIZbF36rOeLYUhormeUW+zJ
5U6/VWE/ndu5e9So+0nDdIHCQHJakmK1JrtigOMXbpfiAulvDxF8GIofDfLy4goHTNgfJec3ow3s
dZHNWZ1CNIEnQOmu17dxgF/cejrli0Ujf/X2Rm9qR6nQThYtHqDC5NRwyKu/my1RDIifamXsrDYy
OTGdtWq9zd+stJuldGiQCgL61wvowUkyJfIVxs7XGzscJUImoekwPQ6BwVsvB3m7gmc1KaYXQbI0
fZVVmKCMl+G9pv+M4UpVoSHHxRH1F4ZxZsrAgwtT0fIAOiQe69tBimOH1VzKLZ5R7ug9x4OdyaxU
znlKdWlSO0270oRfnuZfYFazOhnKSinTUDMhyDlebjUJivC2vqW1sM6h+vgxJPsxXd5sXYtWUK9M
1jqGAPgXlC7opkTgXpdUJVmRQX8zoYJYPMIdr0G9afdxlI4wIwxMYJxGWa1/wvFjgWaNLuS0H5Dm
EPWX1sOb/P3xYjMOVMDHn4bp/y705sM5dplcZ99hI1rxBBH7I2EcgHRvscgL23ppo+t8V8M/Rjfy
qbfA0rBUHM7fkhv9SYu1JlQ1CPARwFsQpJ5LTtUwuB0H9f+9An/jix0q3DwlGgzK+0pzdDVtRqIf
NVNJpN24eEAr1CKoggZx4zFST48BfhyfftUN7b5XYbiLaV80b5Dofo5TNvcBfdDZYfXUaMzU9oSS
8IUMLHDFSaAnHG7rQuWpQeT7e5qx4Df/aznXiYAO68EHd18g8ZRx3uLvon7G8kK020p0+o4F9wYz
ewwsM1qJy2IqdNalAJL4yWz4tg/Y1cLGBWOyDlvNZSC4Mmr1h9xnBubs4h/qyW1JYITD/Z4JS0+v
hlNHMPnv6SIRxonqhaGUMZn0Ywdwt37pGY/rJXVoEUbHLvp39HKNgq+Gkn+Bm5n+SfvNAfq2ToQz
Czpp6WG0dYgUs/GZr3nEP01kbno+3jgk7c6hr0a2wOHQ555iwYUUMQOQZBMDtOpKmLV+rkfcULgn
dEx7o4e+hWCaCLSY6WFiY29xKRhMhcS3kWj5qOO4spaoGINk6rT6MNqqdEfOyp4G38l7lJ4OYV1V
yAdCqqXGMN9Qnc5nRzmtknFj5S03+huHESqKIaLac3Dq7EX93DuQUmMqtT+ZvK4uzPD/5U83Y6W4
Vy1F1IASYkxeT+QR+dDK5+dg0SLhOCOD0VHD38c5l98LDzm+nnwvE6RmVcP98GyLWZ39Jl0RJAPy
+i/HMiKbGQwb690QtobFlXseZus8yGHcFRPMr6EJWppnl08BxaCwtPLEo9DwL/A7D/UZsX/wo35i
dsdDu3BQfL9K8FZtlEdHM3g/GCvnQOXaZSH3HKHYQgACbKmehUyF02M9eHfoq7EakSTRyaC5G/lf
91guvVRfTV4ERZKQxdS0SY30w117Kh0O/atIcRJpUn5J14wwTTEWSos0di8beA+fgPBAeNmtH/gL
HO9LGZSYMUSAPgL2f3t11tvyvU9ByxE661S9HZmlwDavm1vEsh7YzmU7O2AeaQcXdx9VqhGx0H07
UJcP7j9sS640r6jk/BK+xMI+XOWjvGEP/jL9/iZbfKYkxr/EhhYZaAr50ury21ZpOyW5ycdkVL5g
fd3/eGJbYq0t1eExgP/kP9Nup16E+IaWVj3zNhd8mTQb4FQl5sYZet0xHCVdLyWftAMmj/2zOSGR
s9C3725Tci9cijhqBSK9Mz6XafDNBmtKx6QwAuDiSipPjEojbenU8dMJKcPxrYJtmsYXRgWudsTx
e6s4aIwHU8/L/B1YyvNaizKVvFdh7RxT/LGKP9PQRHiuyRI1xJ9c8RDQ3mY+U7GYkDZgWvdjm4bM
UwGkiCZeSGiuzclU6Yy+psFFFOmoMJ6ayO7y549iyifmJyf+deDUWxPSZRAQ9CzSJN3aIHA9+BRm
k25YzMp6sBfAy6ZO5XgUBJT3b67yMhra47yBenyGpfDqWFnLqxel2KgEN5hVp7wd1fSxPe4UYqbi
wHxd4QZhhfZr7eccnoUQ4bobJIsh115m24+kqiIPyyYQ8xDwT/f9wDteFFKw6qIgTsfJ5efSrnD3
GltDz9Wkfrlx6BmWHyJONmEnkoZyYkoQuCiDipw6lZQa3Z2XCqMnOyC8jg4UU/C5RnFjcrGOuunu
NlwyXS0KW019LNHUJF7yOvKpU8deMNsrA2XBKS2TbBJ1trWM2IePFvrzMzumtYJnlb95ubmm3uN9
E29nVzdg31IJpu3lQ+uSyVBP/0tWgt36preBr4BCGp7bPhjJ3e++OBVFtRm9YZUKjkAHT34AI7om
R9jKu+pw/oVYd6U4H7Zut8moVkPerbCx1x/udBci/DaXnMXTVSV3SxRSx1+j5sF0w0WxLnRb7B/W
0VEWxQEQvIlFYR7mAfQP0dwxvyAZOB6Dy0duS+W0FgSp2MvVD1iIbFThSH8dln2PQ4NkJmnPTc04
CtfXgFKMTnvD9FccqVgf+AmN4nj00hLlT4jF5zs1CadJyY31j5BUSCuZZKtZ90Jug366ZZpSy+On
TCVDn1fIA7QcayqGpLegysdXk8HWz+quD4vbsk+ULMGuMkikPMg9Ih28ypmy1ACROzzWkWtSi+nn
SQmR3+GpLL3upsCZhxWukEdw8JW/Nnd6ZoB66TUYpuQ16fQ6rYFVaVmSUHo9PZrn/Hg54A3oScX8
FFLH699o5AZNvk+IzezAr8op+3HJXPaIhgyMO1dw7q5QZlmxJ8yHi2BOYCF9LBSlLQn8GTr230Sk
6mLYGgN9x/ti/oE79QQxKKukwhXwGHhFdWzYY/QCU17YlXQB799BknA+3fxcL7nW1DhCJ2hvQ/KK
EwuBXb/N3+gKpv2NBlYU7zGXafdKyYzBuhkxF0pK1FjNPv5l51Ll4wmbHVWRjxYFDwMGnu/BGJ1C
SagoBCG8gkdWnuZqtyuIJAORU47xhKrjSJh1Lk26BcUM3/gjNlKvmWUGavQi5SaBwmDzS0ipsZm0
fBPhf0CZPMc7BQiC3K1y/Lme+1ZZfOd+L4Q13b1bUmCFNiJyJYlB2KVBhJMg5eN/a7t9aRkfQNM8
EdsWkIR67nvqipqv4McfGqAir4DofyYd+j16RQy2BpgDHgVOYstjNe/orcff0LBb0RPa3xAjVqUY
H3QVu9gIbLdXo/2Wr2GDw2QO6ambvmoP0dkNwRchJmZJMjZgPXxEHD3PxK5amZn30YDpYHXyj8TF
sfV8swLnSHlxEvST0knIzcDUp9agDJwAO9e4TAmjGT0nTtmjasx0XNEcKt0Gt9s87SHeFfODW8OA
EW2eqNO1K8RGrz1qSKspQuI6ruIhZusVSFW+7V8Qs4/fQKjwuThbS/blRP+FOxRfw0RAn7NmYUM7
q1PGQkvjZVqPh6hGx86Zk+BHTKVP4zAYfqY/oo0M5DYkJTQNhc/iD6Y+7fhRFSmLGMJKf6+TgYZ1
eOG/iUE1AKmxzaOMhx3nXqBsdFxqxzgH87pO6nskRsMRIUEkwwJjy22r0oiD+fpk6NMhGiFiAr6s
TWQRLdb64B8WhQaPv0x7aUuw17rvqOiWWPqat5DNYkHQm2cOYbBZvN4ZtFsxf97PLYJp2hs7KIw3
GfN+/Njvi5nZ842NiNpWDo6/5Kf4h59hJInEJkyqLO/TdBCNZei0qCPm1iiMn0gMFRSdUOJZk6kj
+d2tG41cEprlZ8+yM+Wq6jNyUMzsYz5cHkbqjgtSgGlI7EZBU+GsOq6wce2ku2RmhEdxioFPH2bG
md2c+2PGyjwZ1I2t1rfBY8QDl7zCO5ed7GvZsllo1AJjnbYDYmKX29Jp4sXvw7WtGCUCCouY8Ljf
UHGwMnWMnRxXECZL6kJXQVtDQTizpOBONlpHz2rtPFdT+zblGb8dAEp8jA6Ivlqlsn4Lea6wh8Ui
6KqSprEapTk9Fk8UkJSacekCB7/qcgK+eK05rcwUNfd3LZvz6E3S+bF709OyLZO+YeXv2FotR18J
vK0Pysixlzlwi9i785DbKgRENBRlbER/LHlhxsHZAysBJhujBdjZVoY+3ZbtjjgQoTjNLOTrUXLZ
xN7nGswyLC3pHy21Rrr3pPBgFmJlg/hRjUXyqMsgsEKmlowqCbZomRYditWYrdZBxLOfF/3pTMHX
/OrzrCySIeqkYq96I/3s2vAAnq1P+okyZBEpBB8ypPek0s2mzAZGYQvFKAL+TWaGhAWsi/5z9o2i
/Vq/7iLHOc/rdXEC32SM/nIBMsz2wqLoClYpLXFsQaf8rVryQm8HR4ad6Sgg43KKYRk0c90ThWNn
hChvFRCz5nrMcWnkVVmVMbHnTZjz9n/2EcByP9ocAEiTBlkgXoSWVkldESRcuBQLIahgt5Ne4fFF
IaYNgF7D9z6OJvEa2m3Q3ZwFj1L9e+IH3qok1XoyySyI/Vok/dIcxLsWDY9MQgBJ9odGrG5zWKLt
bpGB31gajU4NikeSQJ3ZZAXMppzxVDiWhcLk8OYtePFsww2CZK+LAwtJ3vydiBZ724pkQq6Y/8SO
siPqsBobLvwl1yFf0I6GD40TbUYKvu12p5FBOTY+e2UqBt80tPD5R4kDL7aUvPCdauQ74DtY/TPy
+KZNSj4qtXchAlQM6bgPeiSzvW3EjIWkf66P6hlUds79coBsNNNkyA0Vy64GIL6e+44Qp2EnCpqi
GbRBPDAmRhBtL2RW99wB0IFt5VKEcvo03MOS+cjZ5STIvAxc0fdNXbw7Pz+4nidcwoS9Q66YOFAN
eVdlzI9TEJQjUPzHWVMSzjWmlen1K8W2u+Trkn1vv1sz2NkPlobTnV4sPmajfx0ifNNZTfdn0V97
M424uA8j5L7sonV8RSvkXwur8MLAxKAKH5NzQ0uaYyVIelc2R4RGTO3peThOCIsE/ZbfQ8sBI96A
/0QA+GMOl9rhrYm17cVEHqkgVp32oRwiFJ5kNnJU1/HxNpushcybIW7GhjOJyn/hlz+qIhzMYMe9
l+mbMrS62vmJnK9Re6L9zwSJX0U2eQv3HsDL17w80fX5YsqYRDsQ6ROQhsqrN647jpQkWBLjBhxp
BiVX8g7J3lHn6W6mmr8Yah4IX+EU+u7uVD2+XypTfr6kinWYqfXKm8lfwNaRU1RVW8Q3H4Us/aBh
rIkDf11E4I7tSI33ipKcig2zzSNMBQIYkP4azjF1wqDLBPKx9gsOLM1ZKT8daJUYFWjoWwgTTGO7
PWf0nRyJUr5xAD25HcQT+goK2l8Yv6PAO6P5GSHSDbcK80b2JyMjuygwoiVs6JRDDMb6wgvk2K1/
PB9q9PnEHzjhhtw/78UFPrCpowqr4N+e4tNBNb+Neu6b/oJSFhQqOaldY996R8T+3be5RWw9K9+F
r8spjdBk37GPdO0CoieG72kzQytcxbTghbPurNCiYjgoNtpMfF3bmzplpB//MKa0fkWEnTearnTC
9KR/6x7IO7o1p1h90D7mMhFv78mqNlSZya5idF7qGFqP+Bzbsf4vtLPLR38QHEWpq69hPao0ikxK
tlhatfQYV/SF0ijisPd0pQN/lG0SOPh8iJ/1mbVjKxnkEDA/YvXCyU1Ivxl1pkL37oUeb4Oszrek
1Su5616fTpW1FM+IVCTzSaDrFIaJlrKHoeukAAeFxswjspKLPpcOacK6LR+KChdpbLhhI+cqS4vZ
t/gg1Aedn4WdiGgHeiFsEGpIjMcNFPQkZRijudyTvKdXtqfqEYVil7lS/ilS3sIIK/HV09wi76uK
m3qLP9yjtWf7snKTt8JoBhsW+K8im88JiF0Pnw/Y+Bhd4HBrqpQ8xLa5kQ+2pm3vzWxqmtXUuAnT
EIVgWYEtnV+GfX49/nHMG6BGhzmE8K2WUlyXJTNGJ7WtJtoEeOxGRv2YgQD2echshlJAJDBlmTrB
HZEceMn2fOXHkWQd9M83v35i0eCHHzkY2NbMKUBGaQrpEx5X5lFhySexzsTbAxwFy0jBsIhUzERB
PUGX1E1B67KjS3+9x4C6Kwpe8mbDfrqySPkOzuDdGNsZ9bZEwDdGyT6a77oCpghIIRqhQRsXxSsY
6merjarc5A/T+6QjCiTIw+1RImy7jJOCRuc6FJpi4OYwq5WB5hKZ6jSulAEfGuGbdDv16GU8d72l
7zzbXBU3l9g2Bti+6KXsgiDO3xlHR+zM/2pCrGKBcfJSs5St0+5JL60ZWHJhfPcCfP3yCV9vj19z
tFqDO0NuHjqd7eMXZoQVPZrqR+G6XjVAaDm6xutc4Pjpczn06atf3lvNOaaG1dE0LnsYcXHzj5jV
CTM8LZbjmnbhWDBVeKDwlbPsnW88gu0C/MorV8rcxoSu+L1QJDh+4mZCpOyhqE/T4EHh+mKfDpkZ
52OzNrdwaqbiYUXbZc4A+Wlpu5NQDZQNhV4q2nZZvsLz4wImerntO+e3mnn2DoJRfjr3wjAh7T4H
AoMHDef6H5THqpPuKVsmw/k5rW9UtPEw3C1DBlSGXe35/phyTMBYgIZnanQPVYVXkI62T1grxJ8d
X+kd6AZmVv+Zgxhz8CHCIbDs05qmWcofq2TwtcxEIpow7ngfPrZmqwryNKx3VGMb3COuEX6pNgI3
LSlpLnC9lfCRK3KPTRc3tw2u28P4t8FAX0ARRpBZSB8HZcBByeCE3/09p6v/VgsL+6ZFSwB7NKpo
tfVnQlOY3TfWA8wW0TONFG4LE5H8fBeVbF60AHhF/rzm+PZn05cX2I+x7ecK+b5P5xb9FFa2d94P
lC98BKDqhmSfA9J6fH304+8eHh7AFq3snmdoQSbyHOwvbpqmVXD+ry079uRKCiVMzMTVxTayK9bW
4ZmoW0dBryM1mNQoE6jN343vdIxL+d9V3lV8s98jMaBtvffqFHqBAL8LS3lzt5wgK9r4Bkk3/nzl
WG+Ssc2aF7IcT9I7IRp3x+oExsMqoyPJgDZocGv7mBdK8XJSZ2S9S8yIJsRChrTfYdwznaa04kL7
5eH9qVUrNGdHvi9xDBw4TbfRSviDRKnK8EDgBxAHWtWaJ54Of7VunN1eNEcjLfAUUYPuibp+3Bte
4e0PpqRe/xcTdrlEUMHR4tciUMnowxMo8F7yB1MUajdFERoPNp2vq56u9GGrTFXi0ugJ0Mk7gBAK
TBY6f16vE81kPGG6H55Nyz11Qrog8/myKs2b1gCL83T6Vy00prqbWxTLIJDkQQozv9kMiGZ0EOSe
X1eN0UeWEtWRxLBystQLd2BG7+qC7RDW+STeQQZ97L/9UDOLzzEjk+WSD+NEKt4vePHhRd3OYEM3
5tSv49EsV1Iba6i4uOdCd3z6q+PYRo8eLm8jOnfFmGSap+d2g66hteESG/EXbs8kTN23z61yZPtm
5diuNZaA4zYZX5JvcSyKzX//h+oyRWMWLjV/R6QT/T82mL1XDtWcFo79c707BwDeU8ctsf5IQk33
KDhcGydME2VPzoMTqbvWcESFJP8UfBch8AFRQWQGr92zaHxktPGc7ZjC0Uarnz6Gbu7RNAixwwLt
wqNtdqFfNJFLVuhxEN0WyoBrgprdEgy8F/p54RxZtaGwQAL7aeuojO5WVhxb4aflUp/5QNReET7d
haIt+2vEJB71oKL5wvsx9se6tAHbyHEu/vqlu+FW+WRUJmeGmGF8JUNpHImupeT1LTkr9/Rtjz2p
+LUfOGayI1iCQDAtodAkuapwYjCMDF7VflvgC8AeBgRvBmKHsPDk70antv9NttN/fmgT72xzYVB6
UXk2SetfwXpoaJOFPmXSvILvtjKnVorA3VG60ZiPIdLVR2RZmTpaiJWmZg6PUt1s1RC265cVE3qF
/LxJDgFhVQv1VGw2o6tnQyECHl94Ri46ew9T8SB4tFZ8MzPE7YMH6vaOBOvB83Jq74mhi7X/3Zc3
j2vIJ8zUI7YpzWeKq/k268VUj7AYWWfHHFQiTcnw7jM6lHt6lJg8rrBzj+EcUn9X+mOdqN0od1js
PKwbRYBkQhZltJyUwL0MiY4iesQs54HEY+/ufsWzfrLq2q4Ia+0Dy9FKLb40kIKp4Dap05GyGSrr
aVXJvP8UwjBpNrctLTWkLQIgpsXknUjTEO/BTgcLjM4/A4ombn96b6h175oKlNQOvE8aQmACoCuj
HCwMLgp6orM23Uru7jhH07/DpPTJXH8oJldAfTDe7oNq5w8WVFl5tQ5yYlyJPRoWP9b70+nGMPoJ
i+H3SALAbAGd6yypnhTNJBtE0BBOwryGmBhqRKdXnrMPvt2xCmlsusy7HntJw/8isTGjSI5btwL9
qBP86K7IGdZlTqYw4rUO5lXIuGu6FpgWSJLA23YAiqLoWNM6sb4TUi5pcziggqk5PYOrOVj2D0A+
1hFucOSG4kuWUqv0rnLteRXGmcCTAiQ1yskYoXDWbzDn6CAl+nCkkDPF3GLo248tDeakCcQBVbqf
zOMaDt1Y9lMQNsz6jRdQ1yUU7SXBqzlhrP44yWUdRt3YwpHkkge3lHOETfKW89GiVW+qB8Zso8H/
FIsYFYkFHalspwYPfBeHbS7A9ZOr6c9tn9kIkWUEnbJxMPmDweDv+rWKJgUcTZOT349LFuE9G0L8
W3s4TQuwP6G7+j85jywiYrQmFw1XAYzLdsPeYfULbBIP29cBUHAU8YMujA7CsAaG1aszEYdcwUwr
ZtUGBIvQIi3Ms2m/jzRbtI56RXZtmlkWlZ+o5H2OSOIDnKZkUDZe1gbI5S3LDsWVl5TVNuZXLLY5
1KAdC5xwEeNjYlzESVgxtjIvZ02qSe5Pq7y9bjFimmnVOoOA6+G5FA0fP6OzotYMlEFutwhfw1oY
B3cPe42z8pyj5F0PsH/wlRX5M4xNJDv/jPoTnXyoNXcxeLP/8Gkg0CmCNqTGbkKBmNSq12guxfIm
sVtYgqTv9J/g812oZ+98d1Th2mNQWJV1GmkdilsT2HLHpzfXceR3UhG8+VewWsnCo3YcjCN7aB85
ipQayiIzlw+S1py/BKhyt2uNRXCpg94xYQz1mghZOSbe4sdbBOYrDxerUnNHpUURoSo8IDRkrHaq
gWgtFWmwogQRnprH1S5mcddOdR7eGTdJkQx9ima6XjOLEQNUT+VlewJub/CIVI9bevQPi+fiN1U1
nwzYqDhkmz13azfL4KEkB4Jo7DWp2wy4jjE+seAdgiS6GqcCIqy60Kv8DC2SCPtKgsv8rRHJfp6B
4pUzlNENVKnta410fKnehfO7hGiOmk4z6e6iwhsXJ0vQyU7DTVgWCof1uz/+/r0MnhSD7ZyIPcCo
3KRmAXhglr4tyPwwORdbyo5F7ipLt7sc3ZrmfrRRZZPKJIJphcndib6wzIFmGjWi3nZJ8ostMNPv
cnmZnA5iv4Kupyq/NqMXi1iyGYeoyab05XCuGgdr7qzzeGq8GKZheJUvZSUPB8RTk+Eg71pu2l33
89aG3aMbEU+lznRuD3/fFfjEDI477u4tsQ7yCRXqdb648Nw3ZtNgBrRRZK7KIaoTwswyW2ueg4/K
KSUULCpxPgnCVaq3mg8RNdUNEaoDGcAcSJJPhnM3HxrRQj4Up8sh58DsbEDZFAA9f9IBrZaBSho8
9HtK+h5qRiU22GKyJX36O6RfrOxITt9HLzdlzVfSbH16MhZlR0113ahqVFeLX6i5zaA05l6lJDOu
+SkvM/eQ1b5dutJDkpvzGHucBB/HX7f/hQDt+YkzRCW6umSUIZ3Uf4JSw9GnWDU2rMOjkeaS65I7
ijYks3xZqiyCzVbW+mZLwkoyztds7yqaXBAXkedRqQEQnmQ4Hj9GNrM1W+nR0/3OFpGgYY13kYQe
OW/qgaPrvm+r0ltUvHpuVUJE19v9OaZuUoTZekmvoGH131Rf07BznDvf592dtnPQJuOmtat/5l6C
85oWCmSPmxYOYl0KLEJ/kNdLbE1wGKtS5yJKUn83xoGtTRgvSMThuw4Y2CPfpN25y5HTw7qMvsJF
BY4IM7Rku6DYznvFF0P2GzwWMVUYxb4BAFPUyHl4dOvXczNQoPLRZLwo/axe0Q0gJxBHjAxCntJl
VX+5DqiNuJco2aKfUiBMMx48krrTFnIo72PENuGav0PqZs5RjdXYIoGfwQ5MgVnk2+K3yyIT2zBx
Mu50PyjB5vxQFpm812J4j8xr26MOEnv0LcytFEXo8Xz6xBy/n230lrIhgqm5WzvZiMtLiOMLQqcd
e7UsHSCBU5I4o/Fmdve+aL9riwn0pVmoZJhH0oddT/3+URNQi/uxDQ4UIFG+hvrtiJ4kw+lSNQ8M
Z5W8g4PeLeI320JJ+mTiecCVcUwhqL/B9srwNZRsiop0tECRcpZNDEh+hVM6QQdYWxWssEFdG4Mp
S0+tqW5Ykmwk8TX09roEfQpR83e2L2WDKZ0C0ObvRRvfE76EQMfjOg43QzcUP+akTrSh1Ltgfl14
EnbcKn3cVgGDhqZHgKvgrG+zMTnUU4WC5uioU29mYIBVCQoRyXh0j/4GLsooZsdUH5UmwDO3BZXR
/oy5kielr8sOtZvc7wLg+nh22XWgpESrsaHdD/21tT9T8/6qknwdojWuom53PxbgNfxAXld+poO3
uc1bUL2jG+Cr1YyaPCgig8NzsaB0ISP0wJy7snAOszbulOgeBwl9iz6njQCxhSVL4q71J4RzUz81
5gNh+nQ7jP5FTjjRwQ0kjVaCy8vreriGom5o3xD7mNgzPFsDYiwjjCvnlc/iACypIQJKkrzlUml7
gBtSUT2t6fBGKvtTdEZfLJMGnmLrLcp3Kg1e7YvB2WauIWtLjJvwvD32BJ4z1oEhk4cmOIJlmk21
A7U0uP9Aea8PtbwXO5GyJ4eKvl9dloLRvRAPEM0yCXdsG2h5YCXdhSMNaI74Kd7bTLpaBYW4WmuP
dl90hmGvXcW7D/i9rUiq42/13IRw9gGD2RI69khspVJdJ7Wfb6tEHfIVKF4PUN1SvPidOhG0fSuL
VQ8p9UQoroXEKWHHmu/S4eAMbPM3j2NLJrrEsIQpXUiglyJ3Mi/Gt7aYXQ0ASpfWgXktFtKfAEew
p8BvMY+SBPpyqxMQPwdbKtA0P5jsev7CoX8qPddfCop51HBpXfQ8jZv/0iUc946h5hogrL5/w/W+
a86dlzsSdXpOXBUa1t8+fKw7JOXTeJEAJtkmqIuApNpVD596iiiJ0g5lkmJ3soYq3e6dLxzYkySv
jy1HQxsW41l5/6B5nJobYXkGNds3EQllIO8Nat87Xm/bp4kXcqMHSXXSTMQ4jRWTsF9jdPS6klWT
qQkUXLfPFqAaZSkBrCYOLYN6Z1IFq/0ERB5dXfhbT9f0uit1SyzPyNhienrXo5wYHsG2R/MP4PxN
Xsv0Y7lqKnAPf8+kQIHdd6mcr4oTybYE+UUhYefv+CP0LQDw8oIk69sxwQ0VARTIpcxzPVwmzL7h
Bw7PWagFCMC6wLyJz6CB/NlSWD1VoVbfcZGsP7IMvjv2w3gV+aoxf0ERcF+ian39oPtzpXbG/DAK
VX4qkkXsa91x3Kk5lmeBpIsH45UaoeMMGAl3skASZCrT7KVWFv0B/hJvdMssCMHCNjAwegtFESkV
2i6Ocz9Yn7f2+ctT1V+SYFRpZ014df+ySLP005ShScZ4RzoTJyH/KeiiJTgS7VGweX4RhLHQCOKW
mkauACQWZsVqaVq/kNJHKdPVNJveQ2Lf8wGvqCqKJXcLxWJVORHM6yC8zjT8pRM2NtW9lES0vETr
YjuVmITa1VEVoMsTwMjOY70XPsvh3wdv7Nn+AnW00nsDD7FytnK07BHQ+bpY4fyDfiJr6toEu0l2
0upBhkBT6ThHUmPaCbSbtyYwHWOd3q+kwY0cEawopsXCETyMct/qIimI/10c/pZFUmJyYHZlLFm6
1kvSKaiQ5bSxXb98+Q3DzVXcDPPG1rK3eGILrscX7BnFmklgNffotstIVQzCvDawpNAt7SRMN4uI
C4jDfThUw1vQ3eB94aABbBvX/dOM8p6BrZn0fhfRQxz1lSc0E3/2EyrbKjLaLWHpGIGW7SpfE7dS
KDxXtz5kMvHssKlyt8PyNz810TPlNbeO2Vg2LTM0+o5YdZ/Rnr7aVxN5071Oq1cYzt98pht4EN0G
gVsT0eS83DdfN4SqiZPzpssB0vGDb+SqLYFXQbkbr0N2MO8Ponpsv4rYlQwdneNXvVuRtuax66Gv
6mFFtKyQEcrngvtx5SqwYd35XZXBRxBWBfNc4JC+VCY+e0ZYqoztijH9n+jYW+BTTHAl7AE+EERI
ljmoPOYFN4bWBmJ93ddGqkGVRTiSigmoDL0waApTCmRLscJsjGNc6Nc+bFipEcE9i1671hgtNA5p
nq3OOdZcLFJ+YXJzT5LjHPz1ADXSQqjZ9p/E7uBGxxZL4hB/yJ+EE0Foj3icWBlshs3FPtiDVv5a
tGx+x42baLHcMqpzopWL4UqzczIYKhkLXbUhGVAGbxHX4R6VmcMiK6oYQVXTSflveYmt1TbPcd+2
88CcTHsF/HVEgUMUITjHkfwwUVETPL9et8S1d8mgCe8ZivIp2j/9FbHN+qLFSsVb9Py+GqTIP3DD
TIziMHyVXV431EDMKJzXBnLy21BmQdUxMg870bH49hBkOZO8XGHTsq7X8/j4y8/TtUavReNXgvDv
gZvGIeM9ouY5A0StncCjsIIfyrFyp7WFEzHw1oaEOElfk4IjUePat1+XTRbrhfB0lOQrtoKJ0eBm
FAS7n+lj/8wY8HmYp5FSD515HoHx0g1Kn56PdO7Io3qLmaoks+IC8UUwf9zc6aNI77+NQacWNGaw
6k3uz7NfsfUqkXmP/JN7RIm8V6ddZGeE4yw2cLtJrdzhtiYopZzyj6uGCULzUFbOq+OMX/tvw31V
1hyvC6w4UMorjoihc+fJR0H12yWFDQ/0zHJqJzZHIujScdqardTJ3ISMGUhtV1ERqiiAnOzCVtl1
kgusQfOMga/v8d0IAk3V0UQZ3+TIgSOnRpmZN6k/i0rwDubK/maOsJm89/DCLZSiJhTYxjV+CTcm
0qvfMsk9KyJAE6nu0IbhP8oilqRuOzZSBE7UIZRQ1YzaMkBwNQefKsL+YpY7+tCfXNAxrroz2BKR
8SV+1Wgs9OMDpE+iZSDisktjcfdP3mOhglVUiW9/VG1RqwhvILizs8ZBDjGcZeTMRoBS4CHPhv1X
q1D4XKMzNgLVGqGhBwFb5OOel3hBOednT+mxEUmMUQFMV/inpPvvboj2009ztiLgn8A3DmJqI+Dk
5pi+l4iajgdgaECrVpB8vmh83YSjEsOQM37gbgEjoDopEbhX/AgFvIrVlXm9vj2ApS11HX6TYuki
DnivVrVM5bFqqAywClxoodxFWDtxLfMSyBsZTXW6O6TpBh9sn+2wPaxbgJnUBO+3eT7lCR+sPOor
dCAvcwhMdr+Heu5KJSpSFYF8eIWSQcYTmesfwxlyi6YSP9BLntfqd0bpOrWqRtofOObpRrrocs91
D6r3xDY44VecveiRjRfHTCVe4I/QYHk6b1xgsi3iF9Zd/43lSnz3KZ68j8ByI4wLPee25J6cuCI9
lEhNPJQAOlaabkVWahgogKjbeH/bVCjy0h1KVYuN5L1BzlILHJMsHjL7Q+O0bZng51umxgrQ5EtG
D8v96Qk8B+TXLupcnYGmqo7hJBkvBLdb4lE3GhqmiKWXNuwVbxllYfdZp8c4A7yu1eRuWMOVmnyC
WTRspbydv2W3Vkxj4bBkjdaDVzKOnBNVGI0PgszHscNJwGcPY6Wpdt5JthmVXSQBtpxqV2k8peSA
olAjEEADtG7RWJ7apTvQB/5OiT2lepBxPxwowGK2PYnO/bpKXIp3whNtJZygo7t50YAX3DGMR3mQ
Qgkq+0IZPq3g2OxzrqP9mal/jHnG2F98Uaw1R8pSPEpVMOXvzosWwPLe32o+dE55jO5YQFRrYanF
mTUIULTDOk2NtL8FhroeFGAOzquBEPDL03BiquYI0r+Jygp64N/mgSJFb5Lj5GbFp2FKX271Kuky
NsW6s8fJwdvs9gY9B1BZEPSxq9p6770xE9xs09U/aofN+vpG9ix2Wtxk7ybAu9P93NTzxR8XOt+s
pkhrsqPNuUfPGJx/Xh9lC9hTRZhxzI/yAqJQ0LSkdtFBOTPpiZYLCB3xk6OTyJD3k8YCkzifOTAO
0Rz15b3FaKV8qBP+jePUjCp9P+cfOzde//u40OHTk1Da1L9GpWHLqiOj1asqKKN3MVI5qWETaNci
TvxGP7/C+sbwq0sqy2yg/YiLIul7ILSj//V7QgMxZJ3cPezGObq4rAzMhlbAjU8AP3otePbPE5Fz
8oLp/461PqixifJIMlkKT8fVxbIVho/wwbUNRrzJPaN7qc91NghG19X5R7G5lStwbMa/7xhwkRXC
G3hf69AVT6AUS4X1p6Fmy4YM0y1pjEXsvicg187zmGQWC+F959oc7Jo9x2ECpo4u5uC8UJTPbNf2
E/2ptZGW4BpEge8glk4ryyUP9gqaRIYrl1XvQWVDBgcVYFP5YDeFy/oCy/qSEJZ69jAVl0JEWPg7
lqe4uy+aLasDENdLEfB2fQxlrR+ebfIBa0zFAYQpwTqr1iYeHmiuc8P/ksmKaGkOvI9fdifE6tqC
j3H/yZG7b1FTJbu7Kx9iag3SYLISbhXvPqf/vlaHIkRI368ObY64AREInUCFHXz0dbaMB+ooihdO
QJpgqFeKfKW4a0oVjTFa5a3iju28vEAs7HcIbLLjFxxYsvKRpgGEy9AEbtTOMBXi6UYuAjfqJhwv
tLJkBmlzy8h5cQ9FRPzdID34Frgwur8YfVSaaZNmrOGnx4FMg6oRBjUHUUa9xVdi4qktDeED8ojG
spGO0hdX/IWAjYDGHsnbGxuKYGEbXzzuhYc73yktgVPkI1O6gIsnLrpG+4tLDv0ARwHIjKVD0g/g
OhQ3QzJS3WKn3MkKs/guRjRT67O9T4uXYKcZAVIlFG++eR3QVMNTPDrB2U3ivhJrSI5OVKdxDTqw
INK7u+Eko7ItjKmGbRoFFx8pevbUt8j4La4neXzxp7IWG8Rkb10w+s+6UaqE3TzzmSO04M1m6Jpw
Ie/v+5rB+p7hkvgD8G/p7Hwm8aWMhFSx5opKPmJ6ED3Jnr7yrZuE20ZHCoayVJj9kerUu9npM8a3
2N9bH+vSwjN3KDM0cNFzeHHMp2RUDq2PN+NIEniaoT48qnyaIH+U7iH1tDnAdKUoBHydhOPVvn5V
6OlwPO5W9pIjezcIdEX45n/T3R8ZkUPjIOD43hwgSB/tkXrtip6AtMa2SjHFzLBgP/efH94o7Av2
HRHOvVB3Jez7TRVFfarIr8eGd1meWLUGQlxwB1E2t+J1Ha4xS/VGTR5kxJ1pKCg2wHq1yXdlGXgj
tyt69VTlHQdsKGzY9mOErJQqCLV8fLYNtWHVPvNiFsl9fDhCc5fBGr1VZn1f/29tjc5cUsp6zt/x
guH23KsD4hBBzgoCYLVifS4gHKuO+d7zSb77p8Z2EkemI75W00QtVLGMXydG9kSNREnlbsT2za4+
hPkyUHDHr4y+6vRiM/D+mPzGXr15YbNHfLMY8wRd1wL6qLEL5NhKds525gyyl/DVef5ZQc5/Zlcn
y1mTYbtQsPH3Ficx58Fj3BRqGwU++mMna6iAZOlxFMd0o/W3pDcGy3lzmDZyggZvl6pkQjmsLp9o
tqI80TFqbOGXsV4QGM01o58Ou5euATV3QzoZk4BpRSvN7QxkxtpRgOAb2ryAaXVNsxjPNriG5KL2
J0Ko4qnk1AJ/aURFE5Q6+vjr9RZlOKRpcHOq8qqwwrMPnGpGUwKZSHEdJysOXH6Q6Ynes9zU3OU4
sblH+6Tq8BPIAuILH4XRn29m4DXQuoMjdhsUiGq0lYZMzHkRTZ/Khp8o7WkSEb8B3oG4HPqRNmgE
QMy28MUjCGVUd7aubnY9OiVh7JIJIt4j14uNhz7eRxLrIcOXnCqmoZiJgy6GqjP/QLt511+1ozh+
u57FT/aIwhkMByvkhU4TKpNqhGkqxmYHR6ZSnvld8MWZS9fW4hcCqr0ICnr2EGCKR9ERX20unTwa
i6i+LicuL2Q2w4wdOlWIRxMlEwCpaxffaAfVXm6QMo/+8L+DjyMxCM+E5yx0zYswY/NbtPYIP2AK
/1/8P4KbPC6R9NrO/aBC3b3Pme32Dwi6f7BZCOY0wE0fuyHj/hqblUyjek+cBEV4fSn75edaAykI
hhBW8trEfRJV/kH7Df2yjCZ5xG+bDDpZNxN4ODSvdXGrTf+nPBjEFQihVV3b0CooGH+GihyNf3SI
w/E9nVQ9uV9d1my/83lv+6qk9VND+B9QhLRbjFrGyiF8ZeM8nLFdRpPKgHkNfZRIq7KU+hbrMPgl
XoHOwTZf7F/0b7ggNwu/Db1xBk7YzPwszW1ZymmjGm7uabLk4LKkQ2O9JmqiEnsx2Q2pKmD5aunr
ZHBOYMBP6BM3MENsSk2UlK1TzLY9K+uQtP7nu5dzdyfKplwACGzoXxyu7L9phkWNngduQ9D5LFEm
vKC203Hesfn6uqRkwgUEmYpQ9YD6XMBRaIpS2Wh/nsxA+djBMWhj6FJZdt+cVastV3ImX5ymaAsy
wcUfccXoOUpbz4KbQ96wJnxeXzk2B78sAST0Nljf+9i2kY3H+t+ewXG0B2fepNdCFunmcOn4sMf3
rUpDvjcx4v9FopTnyn9PsB7XNWR09GYNyF8XJbW6bETrAb+K/66eA8bLYMShWRg4TwbRd00/sS0+
sqmjIdXezDJzgCLxaaAhRKbw44M5hZ8OmCBXRcl3qNrpWsAZRMgaHrIJp0vWvI/2xoCNnKk3g7UF
EjD44cYLlaBZcjtd6SUbJ45bkJIk82eqiRrfwil0X5nBee3CN9KDb3ywkC+om1e/69MyiMRGO10Q
zrtWQFrdY6negvS0YNM7KcOLiSyTsSsBL/dyHmXQsed+b9Fd68WfXkC5jHyEprqMOIayw7SCwXHs
1ToXJPZGURHsSpJgfKPNPJRpQgvB1zBI3a0qb9Kfc0zcprXmIWL3Q/2hj/Vl0zk/faN3+AuN0e0U
8TOGoyaBvcabF1Ujkup9A61ZR+jgmmnDvhL0KC7EGuEet7JgKv6QCNwRZ64gMNKj+uEhFtq56kvP
DCVU9fmORwyVRfa5ivh3jhzfJLXYQZuUcrAgLYD6DdSdXg++cnu6HaygxWw+jDst1MMVLuBuck3T
uMnR6wF/yVsg0dqPrlomdAT2XfLJg8StlP1nKippv5abmswFsTZFGxlpEdXeN1AmDwpIMLqtz4aM
NKHa1XamSMR2cEJUak1j8hbFOh2bQBe1gxkD/tc18Q6dh0VORYazVowupq5WnXCaAHy3xdo/E3k1
yRrouo2OzbBMpB7eF4eBr+tGlpHmnc3NVY80mFhk//nyxhnDHD13WW7xVwJz3pApHsS7NQZ8fLAL
IIyHrXUXMCvHUNZDUAi0tssE7Fb5kxlDSJhf8vhoiHIrNHmCfIbrL6YYR4MTGTB+i42w/DjNECv/
NRLA6mDdKADxT3zagM6LSFVx02h6r4BLUQyhKuW7Y3T2n+x2kbU5q8r6Swj3whecB0jU/hDh5OkX
l08roDnM/iGd/pzoR4Yon60lhk+5I2H5YDrbJhd3YnJPPhRDnpfM51ApaTD3MN+9L45vTb39Cn4m
NUOZvsqcOjq/5RRctKxchq9q1uppHI9mtkNNMv9+FzFd1RRq+umyvk4wLjFzK5/YixlWuDPjMN+d
XIqZvLt353RrDbwjC7OJaUxNBTeGgLme1HSFInDwAQTH5Q/fNzIu0kn0INJYCA+3uPzZBEzBGurh
RECuZP1YR0SgUgqZ8/U2t2vAFDSCwPRM59qTOXZdAP9LJl2m4pRcesXSntdRsEXuU/xJeZ9yUOtk
v4avqwugSuUnG3W9XhdQna6F84dxW6S4delSqBsalND56EAPh0CrbX71XGdRs+Gj1e4oPnEFiuv1
jJX+RlNCcUyl6hZBZVHugCGOTKu6AJ/xMMpVJBaMzqnl6Y0yPPXYafljZJCROojOnhzl+W06I6Kg
gmwHaTR1zUb6umM+H3xpecHmSjSoTHI1D+lfIYwHT+fXlN0iM2Tx7hCpnkBl88RoY/Jr8WIyKqya
5NVN8TK9APgge5aZL/P7ZPHjzlTqSiSgourXF0gtjvi4It+6plPTdkB60n7kfuRSqyU3tIXVtuvH
kyUpBJ2LHKvTUBdlgukt705cNDdgcrUXbXy5plgkpM5hri83YhFRzTLGu1t119ezdmyc2tmddEPK
P/67oEZRmccQetlyf3BkmjXi+/ul9P6tneYTR2oJ+l7Qw7VfiGGAxL5O5VMfFiXNeyTIlOrYm5b7
WextJnzh5Ouud7wRwoZqhDRJ26zKR9pbheFkhepUsc7s8WMbqPRWRIJq6P2eqU5uCxmIKzwKGRUe
OsIIfunBXNlIwjHE/yI4GAUkScqiM/jQEvWJ4LEpQII4TXlTHPvsxsArik+WigCbOdw8QNYVKzBj
7kvcf/pYo5e1oBVi+x91l6mdrUZRzlodvRtVcBSounFcAd3UbCI1Es0iRdSK+m+1ZDrktMuIs7q0
kGfSnJvKWoE3xNLHQPuAOffsqByY7qHY6ox3HJjyt75pm7JAsOJeqPZy+KyNIDYV8q8DFgIcwRu7
syfOiKxs4jq7QB8JCUd6Spk2uHT4AmAk4ktXLK25hFs93Yaoh4C9oOj30/qQ9UayQsIV0O4OvjCl
9yyJRpJSUUzAY/LZCc5+npqwYbOL6FkBb5zUWxGWEkrFiV1GGHBcmASAPZ+aUEVq9+luk0NORjPS
9CpqV/guo5AObJpHKsjF99eV0UOcxI1BegFSaFR19Mcl7hO+yj6ilZ0j0ZFjDpLdY1IWZahaa9Xd
lfxKP6p5mTcL0WoUalHxS84FgZeiCLZSqSOX4IBzBaiFBwzcXHFqykWTIxJxIZAcwkqsIzM0CK1X
PI9iF6NkiSUoWbkYhMuyk0e1ZgY4NjuliztfvM+5Cd0WGlW/U6jXeRSoG6+N1shG9/sdxCQRJaB4
GsgxzVucSRrmIM1+4d3Q/WSbbwoGMpyn1+xO6pgJMuAnj+950LDZZ3ajwGJHEilwe4aIRjj+qoy+
egd63nqIHIlmaXjygzt7PzB5mnUALeeyRfe+1dy4JbbwxTCa2dw3PI7e6Z9DgTWoB5Fb4ePm5twD
FW0hAVqBDl4bUmVFgMdRgbdFxUjV8wOivJOu6CW9hnJpatLJq/EUPWVLpYxD2jclO1Muav4TbjDA
Ct1Pl/nlAiWTcjdbMPkTZ4jJNlJzVbrsib3VEXIDRUIRkOCiHilHZisdDfH4kuUuP4a3LCHw1t2j
LoPolD8BlLJb4d324Hz3E9FGA5wm+mOtzaZxiwcQCrcF6eJKh14NvtqgGxgaPeGZmek3O9p+Wpnv
7UVzuIazoZavW2cx79aSiOGmUBEigHaAlNYe0xRgRasQ+rd7WiIbvC8txt4UikI4StgwnLcC8e70
oRzXsZoLnFaw6omIW13ZmOY1CCWn79RmdosMNspuDWll1A9T0JggtcWYM9vF8CcSlsuSH+FHsyBb
J2P/G1HdhSAoqCZFgI10p5rRvC6hod9x5hGocQj8WQLxL64gGEFt2FrGyOOMuzELnS1UVCYE0swx
K7ot+lfPbVg5Ib6O6JKRbEMxAfLaD+YMY24Ua5UF+q4eYL9zyTUmxsJshvSDZiol0EuBb3Ls20zc
QJP/aS+6I02NZde4ynX9ZEIUHIRno98bM7ahWIy8saRp2AbiKTbWvkAAVLpe9DaQQHqgt2MR88Op
kPKjEXPpbt+I0CM3RPfvDVKDm08UN9Ir6AZFUUjUxcaz2k3luqNNzpmvCFkZK2y7+/aUWO11Kp7c
FA8vS0Jb/EYbmfvZjCHmfWxNieZVpIY58plv+D+cGYVtIQ3hdtl614LvWiqnUtshEdMLzYbMMtG7
xwzF1w7FIXOLwFjuj8lwUtgIrb0otmKyYUhyOsEvPjz8FiNM5+Wvs2Sa7n/uD6FoNg2G07tcXzVd
kme1tWxSZ+L8Dc69yTBTmtYgqe0CLkbCrcCgRMCtXva9xpsXltL+8VY5cUYhhjYYfYPE/SX9p4us
fSbC+aHbcJi9Rks3gq8zFGEs2Z+J/WMpnl7assP5yOAO5m4kIHmk+nm5KzDgr4NpxavT2xTMdmHD
G/OjBmOhWppI+rv6iOBa0IjhE+ehAos4gzvw06SNbs8mnpobBHR8GDdGJ6yIaZ8bNNZ/uVVOEgfQ
Oe09BwT5/EqJT4cSxKSIGo8q/AzUXDv2MjysjoC3YNhXVdTA7l2OqPMvgC43Nb96W5tm7g017MjT
8JbQTWRt3ndAQHileaq0R16a2qWrW0Ycq8vxq8eZ3erTnxoIr7qsWGBkqQvnp9Y/IL/gvEenfc03
NG1YHLJf4J2SgLxyMl9yPPJcyannCLADCX0gmwNlnGZ+1LpEF+it9XnLqLO1l7KgXBMf70iysLor
s8LNq7TO48ZQIEiBloRA3w1hJ5pPTykSwERN5GjWH5Y9kl8NVAPGdoJ3yrJbBoftAMk3eQz5q5wu
zim92hOZqY4uAuNMj8WbysnryGC+zrlY7HDK2Fj4k/6k0bno05v6Fa3tlCSalfgmXqrFsPBvMzxx
jUJwKriH4MEjupbhOv4YOR6hKJz8Ns3VGjdwdcfMNNApZ+2LkpuA+QpoUd46F5Jf4sUzk7PzJ+5+
7/Xs207sXMp0xywAI7FB+6k94cSU72iq6SLk6zj5mGNH7nXHafPOn/g6j6DckiHwYnvEykHdmXX8
dX+g19xWbe8kBHUTr5anppQ1IXG+xEUsENTm+hboixYU2w3VlnHynLZMYwQFY9qmU6FCcPDXsoWi
xgDYRiaMWlAgP5syNt/LSoFC07dKW2ESCFd+w/guyKP3uwcbR/gWttOn1jbg2fsAUbCHzJDrUfDf
ARg6lpAFtrJn/wLFn0PDryLvUAPSuys+IVqemOmMtyv286hamXbRMu/Px7MgtRWfI5jFOYpX3bXt
tmmZ9Ha54O+HUog2mHo61ukkerPXGcdAo1pH3ceDxP33gc/kvYVBKl6y9MlYh8w2WBfOpfS+Xy1C
XwZbUqhu+iLYodeWtpwr5QoPI/3b2JD/lHXWfdK/KkWo9R5R8nNkPI6+0GJ53kNI7Ps5RD759CHz
2rKAPtJIqgSIxMs42Ux28FB4NcgyZB6kBweKALNpZLT//fP8/OMXoPuDCWqIKPw6n0pjt8grXQO4
/4xNEXvaB1lQj0X3Z5jnb9YcCEmfx8Kh2SFXrNtYRm471aYkxkVXMhdORbIB41HVJx1G4v78OL7z
HGBca6FTTaapJa6V9Esg0GiBXfifTVYONz6ZTdCrfAhhGEBClI/GIBicJLkhC9tdXT0UhZjok8f1
PRzcPKb9AcbrjXxdSSv50Sujey8sC0UHsIi3UfaP/95OjexPxb+92U220SlUvkIXw//smNN5+MsU
Ynuh/NuT3moXBEtUYGzQBtq0Hl+xiRierMS4K+yzmLP9hjVqdBtNJmK/c2cf0B46eklr/g8ybfOP
xudlEyLpJxfcgkW0Ed7IDIEvD9SnQCmzxugznYDgRKE53ptYTVafoKYnBDIIQ5VLAuJGZaL6hra3
Tf80+kJ1vYOZqisL4UmZ4g8c/kWKiCbFxIAfu8mLhYFBd97xyGQ8WSrkR/b8F4szwJWH7ycN6mRY
93AWEIGbyiQ4f4ZJjZB6vJAcMxtbfjyNtZUYO5w4mSvYJnpI0t/FONwLuHuXVvvNmB+bJ71lTxE/
sXcQAgKjkbGppW1dvaoRH7uUjIopaODe2oLWWK+vk+W2Ppl4CWaMX5kRDKF1qCr05Xqo5sFgrqhG
B7kQlezf+veej2xjgClOgHccS6u4ZGJzhDY1qCQgxmwS6nk7zZwX8WHVu8oWfwKq+bTWZY7uWgzD
MUq/4ZC3Ttu3V5UsuCwj6ruILkvFNXE4dFFoFNI63imR05Lr07kOKW1DWJGECeGDmGFoIwrenPKC
GGri9sVuiR4IRYWf6l0SY1KTAcVQdWtIapHoPyk9v2Nm5k5JsqGd7k8q4TitVVL03SGsweawwquX
51w1uIyUB7BjIJYwGyXRAsaf7FQxv/gSmehnRwGHWk42CP3fwMk9mWfV+si7d9m4ZoRaVgV27YJB
Fmaf4ysVrHdFcVqS70hUiCm6qZYGNax1/t9Oz70TQQ1tOLX/S402cWUH9zoSkDX1l9r5U+pa+YGr
Ndqay8995QfACekUToLmpPzqxLx7cACfovPRkiEi8wyEREIFgFFAxpD/9bN5ukERfLjapXxl0r1q
eZXpqAK4vFQ/HDQFo7JAXZQBUZX68METDPzHOF/DEF79xRloCtvd8aj+ohRGzRKSt5ov2GkWijyn
qIKgaYuiqFNlx6rWcCo/n1fr9gSqJalYORPlr7Up4q9hNCXpD2losGeHnTBLcSdpgLxT0bUMcPf+
HH52r3O/QEHGXHvGyxppHuHlb2AHRO0RakyjaZtsGz8N0E+SDWdXHC21Zkx/aJZCKWtyb7XCw719
xlRrGEhVUVLyu1kPEplmP4Mz//wMHhS96ZgW6gciTCiWEA9eXl8zpSZddKn5b8+s1GmtiteCUENI
XH5zjPsx8KRqYo0GjcqRyJS8sG93tW/nVOXWyF/F5a7zWUYdEYNxIMRMXTu9R8sazgdjOa/ShA3B
tsWTviyU/oR9Zbo/mTVyOrG+VFK0iWYd26UB5SbfSgsZ0JFMChXrROEI8FkSnUwbWNW+xMaAdjRz
sHj3vA0Z0En5SmqeDkCLjUau9mONBkU96KpazRFiJMv556pvNoXtWcClDcNRhsl1Aa+n1KXEr+Eb
u1Ouu0w0SvaQjO+q10h3YD1+JPE4ePjUAnIIlZtc7Y0PCkEaHBGOTK76bETL8SXtyCo1Qq4loNhc
t+8F1FpzBW3ujBEurtqe4kgz9cec94JbXLR7ROTJqYzy85mfBhrkU4C1ZA5MX2GUyvHUbD7GxMuZ
AvU+QrEsCq7Fu0oABBnN/J3FQlCXl1fJG6OR92YOESs2FbvpPpJg+g5reqZDfJXyzgQx2S1hUR5R
U/p0SQubTSfsqW5+mK3GJLqLEk5zxywK4JMM6EeJxBcwyfC/Q8jMU3Lo5o7FZ0T/c52E1GKY8oDv
VoIdmh7nAbtMZFenmKt7es+ATRkmw7t9sIjNz6GgyzqSJ0fwckp+nlAFCzhgVhxb3C/gAngqIX6f
DEkjneVevT3z2uXbGRFDSCwmWtv24RgEFfmskEuNCvdHHB+f0AofPAtxT7YpUj/oA2vEkxjs6/e0
HTS9rCgiFN4/HYm7MNXL7SZF9P8xWFX/FCln4U2asaN0Fl4ALG/2KN+VvjoCTL9jRYDecL3VY6cG
7MprtmqFqqMY00qWmvXEV168CdaEtBgPZmGA3t02PeQaGoFxc752ynCEoXbbzt9MBBM2mc1EHusI
/7XW5f4ygCKUYi0BUOFyikVF6gNGP+sZF7g7Qrf81I2MFXSeRWpGlru8f/JLU+JSGLhDjM4o8ega
8y0VMio5F2LfXGObHoThr61pQY30U25zGHftigHWQ158qubV8/MrqluIEUqUscvTPR+EV+weYI/o
0g6GSLNxH4EjAL+wjgbgY3lFCd/gshUA2worDckoxx5VXMIYjVFQK8waFXCq6K74FpkQK+B/npRT
UMmClUSSZsi49F8q9UqNja3tO9gQ39fRtspAUbZ+Wn6aHxy3wXXI6k3vQiB4BfbHocCfeaYgAjxm
sTHrDqOQE3gx/PR7zCqvdw4IfZs1XCagjETPNrpQDTQ9GgXAXqCxIrPdiIS6jtHBKhmcYIHk0lEu
+4BVrtQ0/2fpuBQkXpASebkpoS/umsO5MbISwxjCJlH3DHJMz/bS0V0BtWFxG4ZlOnnRA/TqlDa9
rDU5hIgLf7HUWhWCI3bvD3zuSfrOQG9zebmz7nj+gUjMCUefJg36BazXlpoPgmqQIFOdwXnO3wxH
Avp2l16tm1Buv1T0mWiST6ojAyZa1cg3YABj8dcsndgmKBLcbXWn1YEioEe+Cx8Av9gYMqx3dWoG
DTS58aayTesnolslhqPkLP9N6KiVr/F95s3vcx9iQEgJyNOZEJ+oXdrKf7tTyeHJIZWC+x1FavXJ
OBxvt185rNsfiibuaBRqOXMofjX/XI/Sh5KNFJYkVmPCSwIFkjI22g8NziQT7Tvni4EzW291EJJQ
Vx3kev1eG8D3lYJa8AytaeNTkY+d6fPOQOmnceCREPFe1WLUEWsvKYQI80bEfg/nccoHBmzX67/H
hix7YFna+BtJ2CkvwrwHjFY6HyiC/6aWO6p5OYUHkpbOMtPWBWanbSIyXzTgIj8MTpW3aBNazHTX
4cotbp4qBvqk3roywmlIXX9tmCQXkBU9tRdtWCeen9b2u5XzcZgwUTKgxVDNM6WiMMP0qhb1M/Cn
igQkswPTrCmLFCd5kXfdiWlPByOVt8SgUzsA23K7WQLxXIlBIygqc0AZ5fxuaeEFCvtHR+qq9Bdb
U0A8FUPsqnJbmk08sy01li9WY66i1YLP/f0ckP8cv91xHbwtaGsVtUp/HKlQQUBjBeZizCthQR7W
dTHOsseZEck8Zw7ZywagQotm0YlWhsm4Sphz28ZIDFHJMuIHDJHp67SLvkGrjhBhbJkdNpmAWnFl
VEDV8oy3NIav9hxiq0T7RARaxh/bC4QiqiklD+WdfbFLKyN0r3Mci8b6C1Dvvet5PV/QUiZrsPhh
FmJfE/44cFgREQdhZQDrHA4WxbfOnh2nqtLcHI292YBJ87S0LCRhVYcYLgP8iBS8a3tP1ad4rVJ9
LoPoUYyKTWoD/kB++Y37R+FOFwMe/gxruRc+Xpc17gQZSIxDmF6OnllUJCDJzERzFiFjgRX0QHsT
oy88bpNEIGiFJZiLuihK8uF2cCri6YdcQr+L66QbWdSPTT4MVPrxX4utHd5LI8nD9XDtI1uLAE2L
k4XKpCw4xLtiMgoupzboJx8PmIxMXmgQHKwIdj7fzCBGNU6GS4C6z5X4gD6/sBK0xvX3emaHNFTN
DiKwbAH6ZSC/D55TD3e9KVVV4WuAjQtdRFJYcG3Dq1MC697QXZn4WJTHb+TiEUnBf0mCgNch/smU
+hGn66gFy6/siCWMvVTXa/y/9TVkSmBjfD/Ebuo6jPwQxf0pphZUvbYeU1eFwxyA77YdVEhaHf0x
WbYtg05lzvsaM9gR7x42kNRiJ2QenpJzsEB2nr4oCIL034vYA9RQ3+pJCWpvhx5nTvrGgTVohNBt
sAgFbPDJOqRDwc4Z+BVP95orOMVeZxJweIU5sx1zSYfLnd1+QN3KbzceGBn/Wfvp19Jpo9UaTIfz
JGb0OwZf8uswfOkhtlzq4W95bNIfdR9qBualzWv+AWXTZSEyp1tKlB5GeIl/VxvyRw+pgjfzK34B
VobHtx4BY6i30xCFlaCa72uuokvS4yTRySpfI9bGuita+QiHGgqpG24IOfYy3anZykP6Wau6faha
YLl3l//tj186oIInXQaTUG/2tzvWj2PW3PQuJFwbB4Gv4qfRXGZ1sU0ddaFlwd5Z81SG210K+ynn
zsEu1gWZV53r6rLKEV2tpCbkzo+eNKbZbyYQ3ih2xva4twJ/we1UzL0BGO2yTKbHvpPMYVKS87II
6vDeGfu/y2DOn3OyzjBpUPwDtnp3RBPSSUcZks+abO8R74L4+7U1dZsQgvsRjfOXbJ0xbKsgTDy0
cTsRZecoO55TQ2ivRNBzdSjMPeWTtOdB60BkIgS09WfYlE2EuEw1lW2PHdT4J2CYdre4TUvm/wfP
nXjOI3qEb75vNCNoE8TI/S/caJviqrlyreSxbMIac+veMR+CTdQrZPFi6tTtHkIyLM3o1BxAUzg1
yGrkzFdoyMSUtn0QeLi80PR/7zBP0bBLFD0ABmlKkyobUVur3aC71iLLnKkVb8mmwqQhxxzORrkE
EOfS278uoTcBC5ehJ3r6pq3sXiH/23jiq6GKXds5VWnoyGG7idtKrZ5mBCNsTkI5WR0NdbaPSGEI
/mN1s5moU2ijJ7znXVtTx7xxa9HQNCbsrT/YMqHkPUy1ZF/kl6l4bIk1NIKkg+1hOesbuXoE1w4e
8f8hytexPYljqY+psCA/nmdbqMfnA88dop3liX0cKzympGHMypF8V9tmzYDKzn3WkGJ6OUsV1V95
5rOTgZkxbWW8zoMfMPhokhZ9xej4uPJtZzBNUTVu2X9wh6tTxyXLYaeDCs9r4STssVrlN5MvV0Fn
9VJYjpzJuDXBBK0lbtLsSo8MHSbYnnJ8pHQRlJVdW8iz9zbC8L+DfzJzMBpXVNGznmYFiOtZfGkv
yJay51umTzwQT3fAIjLF21pNkNHkLweZknaNf0JrlWXlqiccgWOBAij8Sr/7dyDyYEQwZowTH2QQ
JfNNZFnhaJSdAq4AfIM45sXXhM3Qsjh/tzpY09YlegNEuOc3KHDPNHG0mCj7SWDeetGFmqIeJy6o
59On1LU93aooJOSSZRUEMGfu9n3LJ/nkP6e9hdfiWQapWusd3cCjSCiF4Bu7Bdi9wMg9tCTuhfXp
2N7n9/1mNez3lnCRceqk5AGOe5JmavkdXLX55E1XwXxS/4Ajs3HeEG9zi41cFIQgz9BVpkSmmam4
SuWK4mZMf0xCaDWFt9x1CyGuxJ8Pw7+mSRqcNbsRqdtJkDepp2t6HiOVfg0GB1OTLK3K5kSH7DJa
36NfzaJCWxUec5QOG8f/YDth3lVpR1ZH0+j7ifbFSu05xVO3YkzO3cgLPZIbWFSOhZi+V2U216Ak
nfZL6CbO57DvjTPV+U/qKhwYgb9b1repSeq+g8ygK5zFPtnD35XvUtEUGnqvd3ggFQDDJcfPyLjp
56bleH2mVeGQSgYBJx9WcTqsxwOZ5W82JuBBspf38fW0XiJExnE2arLYN9NKavsxLC5FFEIdpqRG
YMBPGD4/EL8MNnec8m82h+04QzffK9zz78oMKhGwbNlcCcaXAzvB3u9ozNYi5Y2MEcK1OnFUigdK
uCZ/StcDqQ37etNyGpuPD5+JXQpOpzcwZyyDvHz3qk5OBp8FnGGaJtapp6eOZMvNmD2iw+xKYxMW
/0uc5JdiYg2qZNJWpekCWbm9ya4jB6vTo8Lzyo1GcFv4rjoCjZfvLYFCUfsCyuFwKNr4Iu410gs4
1ZiGBG6MCZLeG40OzbUyp+cgpgvApnl7w5LMHivObhhXFfiyzPnNLIKUg9phCBbWOL/bw3NEicc/
cwIxF5Dt7JiyFyqcTZdDhuD3HVKdhPIaX4G8QJvEhrPv/FsJ2FCBpw9Sq+29Fj/9pC9xYaI6u7eT
S/RawK6xa5tokNC1I97dhUt5OHgBweh+lLXKfurqC9/gEAhT009DooMYTT9cxggXAdktzWqWyuk9
LRWwug7oNIltkst0VXZTclRZMG3oDHUPTKt3DdQrn9naryVLREMFGHxv9TPnRVzCJUr2DuZ8N8rv
58iNynepJy+BIfdUNBkYadvZetNoqLlBvBs18i1dlcbZFF1GLfLIBL1HEG+8QsV1rn777MOiRh35
7jYaGL+ZubaGiXanM5KfcxwSqiIJFjrm9k5VZu+bnfTAO1Fb0uPBBjutyvwJSTQNgaeQ2n3kCsA3
UzNEb3Uqpa+PwKfBk+ElzhPulp+23hJ6r1MO41KaqF7pDlbgxOLMQKM1vx56IRZm+3LW+m5CEQt5
j2HpetPmANsmP8mro5CvKzUJdhhai4aX+w3xkcwAcVx/vTIyIBJTPDdrkKdBW53NAbyt2MPHwbN7
gCLC5dCeE9dSLhaO+TkviYZF/D8XXyRUS2U859/nsCoOtoo73tTQyk3w9gpcFMPtQ9M9mPDBB185
HgVR5TugAAQRz/cLxJpjwSiAzTbQMcfIeMo9KtYUJkMWZmnm/UTMQO8BIOQeeGQiP8VxEL446F3n
xq3L7QqGXC9a1K14AjDF0xV2iL5eD5Bp4zh+YaS4kLG3b7vlf6HgvNiWS77pt7PX1ESWpttQwHZz
e40R8JcfvCwp1f1YPMyJQn7+BOL8r95LuG27VjWSHTo0fBVlW0xm3xOY3Yy9C4zuMVVr+ymzVMLG
o1guZU5Fs5zw8QRux6FZ2B2jJKqKKD+50YiM11RH7GaoJh6lHRqvS6Wtsd1GmRV9hvJf5Qz2jaPf
KzSyP58RLR6/7zVX1Vea/KhdEhfp2V3kbOmNkO7dUVrfgNh6KfOkvkC/+wHNSXvQmteXGaHZVUpK
83RQgg8u6eM2ECwXrdWilKmw+R9i/8kZEHcCHrGFC2YqemyCVVdTZUmiSKQb258ntgUUHTeXBkIj
ixlqRqN5iv6AM9+UFhamBLqzH2fwKy65+2ZmyGYdeLPp3lxLF5ntUwdZ8DpmYI/Y7M6IxRbKmZ/a
OTV/4qA8JWRr2zMOsswKzjPj+d82wEw4Dk8Fs8MpwtSvO+mzOi/Q2/OAY6nSRcZSfXdrhBPCch92
4gw6LwWhEF8m/EXjKyGAF5foCEg7mToe9pj5KkILdbINxfyuAuUeiHkYAMecRTrysoXO+EMt3PsN
xoNigugPXdWfO+oY+49ZzGJqVaHTGWqOiYa5FgdlcAcjlQLLt2Z4jDeR4eeI2kS7SboMvX5E1UDn
rdDlR7gyARzl5YfLuFb1jAZfe+Q3+dk0eJCE5yqodYC2vsw878r7BToznMVwsfc7ikgES0wOuMJl
FlcaD3vmV38FlqAE17qGMlwr0WreUFfOEeh1vWUDoz8Y0RhpX+E8p4jBRGu0yq5ymWnogDgLgBFn
vVHR0FoWfHc+ZgVrlXjuOVRDQyqo7XQ7nFULw7rhJephi0xeQhFm/Qu+zf6L4c19FGrGApt1dLNj
yJqXT4lwx98kdSH42y/ptubnyn0EmDZ1R6UtgocSK9SvlRfr2LOWJTDUTGZOdu6sd9Yq6OnvYkgu
/D33TVHDbQjDvoIBm+wIi2kv7fTfP4Cqkzg1NSfXgxoLFhHGvLO5rlNnonFQi9Ct/Qk1QwWNj4h+
akyuRJAF6BvmInQZYnYoC3nIq6fUNc4nRWqFpZ6YcWhGq9afa05TgSLTvuAjlJltR+nqeAIIYYso
ao7T7XUSyOMkHp0r5NT6d+W6QxC2W/t+zGEFjgko8cnfSG2xN3co2m+K1Qo3VVZ695kZxFShcEa1
DSAUpavClNzb3Pn1L6H1mdx7A9jo05i7T6Iqkd6CfOxFWzzfrF+TpA/sAK4FLmfyNgslrjl1Pe8k
6vqmTswP1UrPh2mgi+Cs2oTQ02HyM/pF2sikmI4iVCb0Y3G3vEr0X1DISzGpQkMGtqVbz8caNpoD
uUnCT9zjHuC8WuF0c9ruYE0zCwb2FwcuXsEK/JEX2se2O5fe/gjRL8db0TVbPfg34+aNGAQXCE1v
39odb/XGbkHwvDB+zp6RNAYUinkzZcdLlVsf6rafETrK3x1GYgoXjBX9jXqgEMcrXQi3ISviHpBu
3+axly71am/UXgf8UJh8Ilmek0EMQ8dLvCKUv0WL8MSV+VqPGOp6g2gJYm8N7qTVmYyltqEFiRP0
Ahme/jnMwzRlDMi+I+/O0qywanrSYIFdnxCyIZrd3KBi/KSw0sZ2kcgl+b7z112nsINHApN3fCBc
ix9NGrGdmnosUym8lNTCj1VTYqeAIE6DYN2Sq13HDPhTUl1ZBBMxiAuTW9Gdge/EklZjm946Ep8t
ANFEMmZl6wURF6/huuBgCl7j+ozu24crtw2tL+0/mG8QMkNWUW3aYT5QJ58RsH5SgwvYYaKvYEAm
TcLrIazCWIOOJqEIaQips83QYKNeQSZHKXIRsqOUvnoWgLkxQXzarTdPzCBbzM4oO++6glFizYOp
XYW7tiHCEJo8sTl61ohSEeOvTPtMgCjeHefH7u6OG/uHvHMS3NgvgzJdyztjk0ZR3izkDKol+niG
8TwEch1UYo1N4LifXjcNRDIgyW/HzKMxYhKcXwxPmvzpA2hS2rreiK27b3hPO/EF8FnZSeIBDGZc
dbPTP4Cc/9ErSjPjeIdV0FfR0w79k/oRh12W8Oz9zrwB6fioMjkv0X48LKimpgLR/Dy9HhBjZf3g
GjaNq24Zv0T+oHB3pJw6RGlM2XGQIYMwYvHH2uJ1ufCZixG2M71wNbxbl72l4aHc2vnGLcGL/QUc
aejiQMd2aFahjLEaaW+tbIo6ycJcsqtrfOwqeOzhIG+zG17YxBYkfSYWZ2K4AggpP79KvPOx1IPa
3XyznnmE/C9WERGp7fifhZjw/zIBOMUe7kXy8K0X6fXL3w34tLyUAyiuakgnwnz48eGrHwuTPZ5z
RoYWCqo+rEVenMnQUhlgqjNINiDuUmGQbrt41/5bSX9/e2xUqzxRScCL+yXY5FIMLkPXjp/UNhzi
UocrnismVNLwOWF0PW0vooWy3ibBWsyQN8gjzmIMlFDSO/WwRRLwW7iaE1DD2QUkBQ/5LAOsDS2g
DsYyHzc0NTPKESVKyqweNQ5ux2I6vXWGcebB03iEXVwEa1gvxqiQPPtq+auC4J11gvPOSX6zebXH
kXZDHKA/4oPWFY8v8xW67jGbx/XzUs0JQAmyBrQxjKLEfnOGmniQmxUmzmT1A3r9Exgr8bssQaGn
5WgxGNTG3bDhS0dvkYzzseR4TJwCnF7XkLmvwlWIw/HVLPmOzf7MobKZjuUHxu2WcvNpR0lJbJu0
eCSd8iyfY+C+UuFpJnqR5/XSq+jHTAAIkmkeIsYlUXXOenmnyg0A97dNQVy+8VL4pZrQrJE8faVE
tHGY/urlC/zPojEPCZ2WmY1BS3G1/8EDIOw3VWZboZx9XX3GnVNTZuH+RVp+ZeSTI6mSrxvDxibx
X39tkBC5onlLZ9oa5A+bqeHmp0owtkh1MHKEuCyacPyV7nktoKj1VANYlrh/cE5iQdY3F4Ei+AGP
KMcP8Et5l1soHdrmIzITEDPK+/gwzxgogHVVx1wAPWxKX5EaY9Z4Jd7DliM3VYAwfjqRKGfebIhI
HJWKGp+nU51B/5kbGJxtu2ejlAIG+IVaAI7Gh4InKPF/ZZ6wovBPenVQq7cBwlPZ/UeRH0HaDa+X
zsOLt14a5zcVTU+IdLzI8Te91rc7G6b5Hnu/pKiNIbWdUAZtg0iXDTs2UE8g3CwKFk3exyHtFVyo
nGIsBTvN+rucIwhdkxgQFjnh2u5evaMQiAkNBizU9P1+dFkF1ZBVq7xjiuZ7VDHWv05Pc9BHIgHM
DeKgMsyBShHh8q18mgfQTXMs+AJs52VBxB2HQcYZSU8bC9pU1/Gsd56mW1qLB06EvHxXJgbE+jkJ
aHv5IWETaO0IgR12M6GxwTYe+TluBv/eERgaiTiHNCLZGqtQg4AwaW0+kru0nrp5Q1fUIwiU1DkI
pRgC5ydkfnnhYySZoGO2bWeqwIsh8TWNnBjJAYPKgBupT4YQOU1kuEJyaJqTcNsUNg/i91jK4P4V
j32GiO+LeXt8zluMaVOnu0nIIUH7WlV17hoZvWQUVlgjmuyO0CQu38eJhkQatjYsjyi3aF8ccd9M
Q7XwtuTL4iHJoWZFovuygygVuuWVib3puJ1nFp0YgoAoOjtTCw+8QyxMNznK6NyNZVH0vlooTzSS
QfX+hGq97mrEIQEA6JBrRsNUgFnhfPGauzBBprTLyUNufMUuRbxBQfF9EK97zcrfUwc/Rop5F937
AZR5ueoKir6fGApdtYrtYqaFhWo24zwXNTMZ8njgrW+1d8yYLq0UBTTxh66BUjlTggC1PJH9XFka
JLIE3j9LbvHTez9dp6X+Kbv0mh/m5J+cD2G671IMcQBM4DYZffe0uOHnLFPi2YsLWiFaSCb3rcgO
NXLv+qrriJ9hA3xC8GUxw+8XL0Wo/oyhFwMylVTaVqHJd2ZTsA/tNn7eAU8gSV8iLhXHJ5886BYt
0/oDI82FXL9DlQFi8f913gl19yB2Mq7W8CQr3ZSikJC7eGT8j+zTOIKtMDCOOPt1Rso+ZoMOv3PY
ak3g4bkYqUfTu6siZ1yPuyU7G7E6mpeA/cKMJOPhM5HPuQ6OFAhelZG4bP5opSLpLvNdhiWTmlC8
adQ7N1QDlBqzTyy6Is11HYFqidIbdiHRJfC9ToHHyGIiAIeD8apiBGkuoVjZ+VZZJBKWckt3eYRl
/b0tskpEUJgwPecqaZC2YlFdEiSklbZTpVWzmNyQ7/jbpxcBzn4rMvZ0/LlJbWOH2nc4A8Da9t8J
R0v0eP4X6LtTKtsWHdd0h50hHnOkBsuNfKsHcwAccegv8UIyC2azkA45epn05fp6Xr+m4J6MtlvC
OENwzvjf8i9Y9OcbGJ8XRS6ej4NVyFIbD/TntELenyxuJYBBm9j9BqrJzjC2Qv+6S7IKzQ9XIjzp
xHAgBFOUC7ShJNddVgr273SUYtNUZTrxmycu3oiFVel0Oju9H+LhI01ZiHAtWYhxg5t01NCx2hIu
bh+RYzo0+OufrABXLBsH0cuGlVpSPmhyfmAmxtOvAfaxRZ5ovBAYLEHKDRCNTlW63luL+qc0ciaZ
iXKAaCTKqrjw6qAso1xhyIkOC6P6ZD8g9YgbWtLXw2KFqlnP6QVSz67SGC8r+BYEqIEWH2tECL1x
3wRFi4PMzJiSYirwY4J/ahSC0EABiqhywgRmW8OY6giUmS8GTBNGH4Cz5qMjoKjDnb5w71xHC+Kt
iuv+e5xmd3uKY9Z2z3tWovcQI2Jc8xjJuUUERA3qq4oGLXoif7nrfF1E0SWqGG5DjfWyzvKRKV4h
F+bjKJlKy5KoIVFoHTjtNdQd83ozzPZM+NvrTJqJpWEAzwiLsuhdGXL1sGi+aPoiuOnKpWXHGAjj
ZL22RAHUu5zf/oGV3xASl0hU5hCHjVfDjuHaUwS52zOTEdkT3diAOzcKQF/sMGWVDgwVOrlycImd
RH3jLtoo50wzewcDIwc6r+qbmGOw1Sc7Q/Xqnnp1etWt+WkeKfIRtMBXiEwihxEmT8fgCQvHbHPZ
82W+n75VIxm1YXm5O9+QWFZkYS8ZlF9CtXq6M8HTVvQtwZaxawn1eEY1C/WXHnKEK6oQiPK8k/oK
dRyLBRJlOMyXUsnksooVj1prNyrlClSmrNIU5bFaMwNP7V7gZQIvv4MCr0BV7KmFPb2MAb3PccZF
fh/tQlRxKcx+kY/mFo6X6sP8EKgK8HBzMyPef1cJpw0Hc/6QcPrcGy9V6fV5rQGYRhmTLFYhnzZn
qQJqkNuhRt1KlCL95/yIYpXBJIeN0TEr0AEHo37zoBREFL89MIBY8SUreO4zpOth65ZHGH4u30Vr
/qTDqhD8roV135m8SagrnPHmS1pYE/awy87J/LU2ogdxHAetEhBRRHkyKK25er1aPYfd4U0+hsVX
EMS4AnH6grNrI4vz9eeaDQLWin/fpFntwOl/pVUyNqVQX5GepYIQ3f18WJtgRKYKQTNORi9S9itr
p9GRFMzGvYI5mG1HEMM7LYv05OaCcC3g5MOPbzTb9XyYPHImMPLcvT9mbnhR6j3+3ljS43pYfsEV
5fZToxifIgf4uBgoGwOJbe3CqqbRSYK1fWHPTKZmQQvIzujoE+7HWvDWMNezZq8wu2slwLUXHfNU
fCreG/bcc4Hbd9hi6VeHJPkLCiz8btQJeFqR76xP2mSL8VQy8lblmFgc854lXwZUqOZXtIBvtBRE
bf1vqAo1OHZyxigNzzk8KyoSlM0ZMYiiRWK+Nv1kZcGSZVP7zkcMHYWh3dO9+BPznQ2RZZSnq+u3
0o7EjnIsRGnCtrMMC+Nk1SOHfA+PIuDcaOFMxQaW1ShqHFwYWIa0hbsAWCmC1XkwKD+TGbiKSGFg
wszyWuhceYtVWrwuCR/0mPEcK4VopmfLETLiq4JOWFdNyXdnFVlqMXI/0e1lpQxytgnT28xruyQe
v8CiB1o6bO2Iu628Cz/87mtLEgrQOmiIuhr4DarQbkfApcU7fK9hra+ikLQPYhFuiDpU5DoQLKqg
Je2863otBwsMDdH79GdiI5YnZgVAcSc/dRz913QoJVMODMrr/ECaT7M9zz8ISJ+coq4keGQCcDsa
EQoGuxoYiXiCLR0cuk4RdYZzbaw5g4nqP8ptC1jvFttG1ieoF7aCMKQkDlMYRM4EMSajrrwqBru+
6JEHAC5vPiESJsHP4l+7ZQYy2GAaBVyzPEdSJMJyu16anrwloldxMM/bRNvWfWEWtQLaK2uJV0Lx
UGW0vDZCT/+ntgR6nqM20c2M+qfKgAAVLNgidXIn19MFbjXD+6SbzeufPq6zNrV9OMHU0RfEnChD
rH3dOmeqiQ3kKAuvXpOAB/OnEMUCMI0ibn+BiXxJ6InFNaBH1UBNEOEhaxEEx7iI/y42Fu2oL3WR
hX1SRvkrFDYc7DjmEMOjtnCozNzaXAitFC7yj3dNJ04xDwQ1QXylPtgW/IO27XZZBEKNrXF4l07I
7Gwu6j5OZ9f1xcLk8tGaA/jKGYgUj6A/HYJhzMk1shhwyMIvlOHtvCwVzNxV1HkKp45Xh4Mij/F9
g0dOzc9XcTomUQhnUSfp55I9naIBHePYdOEGU19Z00kuOaKaLqnjbtz6t8Aw8HE4R6w910FqKHgJ
dutJVHYWUmd1CjBOVIJtOPgQ6hPXT7dN4OMPeogyUjGf7PsD5nVD8g94exGeJ2V+lhnx3mEZmN61
6lgp+HtMruAGIh5KBEa4M96jSehCiEUCVSyAxuSwNL1vQ1gkHbI9gsueJD+uiW2Luzv1lPHllY2O
P3weOQW3MmUIVJeAKj1LUzrA/PhiGrfDeWLCC0pTokgpDGEocide8MR+oSz03aAUQnYVBYrYR7oB
q2sk//6FnNIdkBUpHBuJ1x9cLBp8VxfSfZik/whc1dgHaIzCG7yXBwSVKWgltBVjjX/hpHjAup4i
+JISuEhYu/1UBbjZ7+w5Gga2Mzb7bXhyhvt3zvCtN00tweDhIQcr8YmeMg1Q6J0fAIqd/X/KeQb7
6fCoTaApS9MUwvy4QA1HoLrVCAIrg/gAJcBuawY9qD9LkBfM08ilCvRNxPxjO+I9cZlmhqMW9ebC
17wjBwbDFNR7mcrsduXOuFlCHJ5D3l7TNUW3YQx64Vcgc/BZB+WozQD4/KZwzULtikWv2GjjvI0E
nZG43PVK6VC07OulkvI8brxxfIjMQl92jgca1Ul+NioGcTiH0R0bmOkDnsdwOyMpy/I6K+ovevF0
B1emBJa7AjOMtUr3q4Sh8Olm3/Exw+9wan1WW/XTArSl4P2zLUkYzmi9SvEtjzVnBCt2QdMJXKuw
j2tbFKVW1MFXnTNJuIqA6/8lyyqaa2K/vH60zj3OF1rGZfzTmgcI3yfTsGCvg9xUWaVbGduGdJqo
/oYmwpaEbAw+EFC+TCgeHbqa1g2naDVHz0V39cYwCEazod7VIlX1BeeIXOHuXgxVOtWDYL0ZsKK1
UqBLk6CYe2SVA+dd9LNraN+XnY8/7TRm60Kst9tSnqEtKcseDyuHiGSDfMkKTvS0T0xn7e3hD7eg
Y0WEl0lumv7pBJsVkvcQAOR3Si/ZbVUo2qmgKUPYbQitB4zghFYupC92F7ihhdtJ1bs1/hVPnWk6
bRVsEFGWb7KxZoDNcj8H9HoylAG10lvMc32y1owBxigLkpXwNIjaJSOc/lv+K3hWsBBvdDEXoROF
NB0O1JNEVHph0+QkuBEWn7bW34x7WlYPk31loLdBFX+BbqkqwOM/DGxxOeOUUl9lHToi0ZFB8zyy
6vhyICpRnT+hjpNoGfeSkFWadgFLhACMw2tajkO3s7CcO/A84EeSh6KismBPnKQke2PwCtMeGEhb
6FysG6VxmzlSpBlFLBOlVy653jck0URtzEY4kqxcYd9dzugYsP4b7obziNMToRqKtmM/G69sy6Rl
YEYwbd4ab1FBZxzq1v8NePiiQyhWa1ayHLCg/Qhco5MDgQzPRvqVjXXteXLNnwbZXseb53mOeptL
KBk5Y8Uxi3aBJNGD0eghpyxDcAxWVibE5/zHGghA0xfIDqCVgnV0Glgzdks6VTNskE1l2p6/+OCX
he9M6sjOwzfriHlK51X+pO4wUxEw56UnF5yKvvTLYjFtaRuVvBXkPArLUkxm/t/Uq25F2auc2WEx
JmZXNSmvBIcRQ7CGytuzeAH75Dc8kMkkL/V4XLpR+toXHnVW+T1Inw0Vkv1wyhl7CitmvmPnIlaz
Nfkg5mkTIGUF6vOzP1AdaEivOnMslXkwHpqlkm3efEuE7ixPKTtwwnRmYoNZKc5SvCCgN+rzJEbI
hTnVppxGZCNYYD5x+wtSUvb3LAaVLBqR+l2/67zk8xR5N3cOBbkbzTxeIdn6ruT35C5Lm7Suv+63
euX+AEDfAMhALKk5zqLZ2UTFG1yngzgaVy82LJFGHdNcJnxODQOeKmbNnaYdDZdhrixYfhMK7zNu
6vRL6lp0A6H8NeuQVPUBQgZMzwdcxgCM5pgF778fqcCQ272xOlGMXZPpR3aaKIpLi28A0dHYbvrh
aKCbaujFkfl1KmL9kzXmYpU9DlcibwXwb+t1nUmT9xKovK34GB4tLobtpPYpbLo1V9eUhO8tTnSm
8Poyh+OLpIE7gmx2pqGQgqHqIYYc5fIUjbDSdF0ODic71o3NUkTk/jmEyZVoSMDq7x0C/wYUO9Ji
0+v6ZrDBZmMJCGZccuip4pPBzOdXKwiriBmkeTNkqUeNU7C+rzkE7YU3x/pcuvkLP0uN1022heqP
rGVWkUvXJcUsE/+nfp3s8AnQQekqEdxMbcrbPJ1jZBHZwMvDovJq9vXCBSBVgpetQtV55yWRiKaW
ORVNGP38ine5cERqzBKU0Y4Y7BnCdLzpeOeSI5nMBjnIMVQo5HxLE2C1K0/K0xXFsGVbu8tflC/h
q2dr5vwlbJvydwr0AeSLM5Oalwks9E6Q+dI2iKJGW6IQ8mrRBAcF+RXjd3MSNuqm9RMlaEFoAPOS
Y7E0cMhkhAFzTuwSgka4DxqkMygEGQxkH5zi/UU91JLv522MavTCM1/aWi3EQPjlB2ToslvziQO4
x/FdMbuc8/U3M/0Z81wa1yqyuFeBwV8W/AGJq/VDFuv9E3xVbHWc9dsWD9NLM6Po9VvQ//VLK5KG
TMvEjyJiLPNHLxiEuadQ1CZL5V+rFm8K0u3LSNt3WvxVejpdMxYygLRI3L0FaSwdRVO64nXkl/jR
h7amMX8d8fLtDZZ1ZTbvcR5P+qUD6AtWwrTbsDbXYoGT5hJUUyPCCYS0cnqjnOvwF2p/k8PtLB+S
MxwII6JU/k9x5mUwfq7xBRRFJv3Brq2x1qGQhgO/iMvxcaV8wQGmXzCZJqlhd6vD5FDUFfTEd4EY
JiCtFcNE6KEHIyWGm3NwrW6dfrXQWuEgx89NGKte+BBCkzKD2mYPaj3rvWFSE05nRzDdIJCJKmSr
tAsBhIMD9H0HAOemyosL3giQq1k3opSMqHeJnFI/+1fVZlJYur7oSjwJGKh71EjRSxY3EGsGbUQu
vNGatn++yPoactX10r+whA4ZXcK925d5mzaVEHgiJwgj7w9yWeMsV4xP9IpWMhVnMiA4XETLbnom
wvM/2j597Zz/0K4y4be82qZMFP3MEviYRifcgnjMC212oa+sAteXr9/Yx1ityyPZ3Ro8RXWg3H31
XXqQoyENumSSXYka5FCBaVFVFd88sJIa7NAJBCII2JMAzM+N4e5pc5HxpWczhoMTKg4EZioJ9xdq
xx6ze60tWl84O34pOiApklZmETommD8NkLNSkRDGovOcWL4AemNyTWc8nwuL8zvxs/aU/tnIyO/o
UcIVX2KBWfUuE6kkqhmBbkQuQUxAdc22A+F8ThDo0IT+phHW6RpppWJjkIeyH35Va3Isfej0KOgQ
dBp1rB7dJE4mzxp9kqk0sJ83qAtRBPSCPIBYIq9bwNpHqzNknXmNES10S7Q8Il/H9UnDnkgtxD48
apERM9zc1PSSfs8HU+vjojaAH/sWf+IY4tvh5rTR0LsIn7kDDebGD2Exkv8Ib8G//Do/m7ruZ0Gl
n7TyDNuGqUA5rXPJBti+cqsYeXli7ZbaADRcriNImvYt83ClYYTheFsmQ8EfEIhEEjE06LwneNcJ
KCTsaFRtEJACpFTbz+FtpESB8Ngb4g9thUeJ0h+ddaUUl4iwNLmNlw+kmvM1mSAlWhtKA/oh5h82
5m07LZa0NtRB8HurE9T3G4IGXxz7/eBQpMJU6UlWi4DGMFDiVmNG8uLIoNy/brH52qx0oX2fy0th
YTJq2K2cVoMbXPoeLhFK87X3d2Xks1VksS2pp0nE6XsIH0/si6VjpJdDVxDyhsvD2o0fXHBmhERW
y5zx8cCasN9xa2jWD46sBbUkI5ugJ2NPbytp0QCbKEjBCqLxKmKWKT7XCLDVQT/r+RhKxXLkqdtX
c79elwMxcN8RVUHw1LdwXFISPKYpTZyjbaFHCND+LmCqu+ncC+A69twTauDP0emHg3rcPS3WXOdY
PAnsfI9SDBGHyOJiGAagsGRdyJBrFtYOT+D9nFVd0Cx33vNYX41hJ87tgMcVxHhqwCyyc9xcvm2B
oaxhoBJPPJd9bOGNujQg9lgchLEasvRbT9+hi0+b4/10QcT74HzvNzWc9mI+GGD3GIVvS9H5Em/U
rvNdxWFptworlRr/Hqv8dCU0N0y2OchMyicYwRWu8jUxG22e7DDLPNCautlDZLHH92vO4Gg7fC7q
RZQJILt2a02ixq6tNbhaDm1DQxPury+/HoYgwir8sKMVbZ44GJ6Cy+5Iv73uT1LLrN2mrxsXHPsS
Lo0zBxa1DgP7a3UfI6txbFMvu7fMDk2XasfZiL9bmx88hTmLU+dpdOkQNEgvtwczyvW80WWCj34z
lQ5+Qap7Oo6T34geIWNlpAE3bpmv+RPogyQEXHIytheR4hj+Ovy/1UYre7tcni05OoOoiUjIMU+2
t3P0/BO0Ju2MkwdhdrsgOhQ+qTDoA1g1QdNa0jwyKgGYa+u36Q8993+P1DasB6Hz3G5iUwn4gpFj
bothf+cv+SO6ZuAHFJZ87kyhE77Rq0jqYBSZx6Wsaf6BTOrwT46aq8DfyiB7fE0PgKClJVF3rhuQ
srpmgzKQCdqyzhYSaDCDXxMzRyI8F/8nix8F6bFETLdqgXxVRtjfw8a9gtZGC0HSz8gZuwPZ9IKY
jTC9ZcBxv6qF8GziZI62ZoD8rOKnWSmzQj50L4Pfu2c9CpNh2/eL9cGaTekBnrEorFsIP/zT5t7p
Budr4tuEFWRWthPO07Ml6o2uxhIJcpq46MCqYBxMKkE8irbpzHGYK3a+fXTRKnzI56UETB3UCYmV
3pMeeOJALwq8eXvECV8fsH80EiZfHilqVgv9/WcDFgT6NgaS52iq4lAQANlKqioc8xlxBOJJs07P
mybZURUa3JZW1tscSL2b1IWlxM6dGw7UucmyW4lOhn4fIdQl3fVr6GOdW5j1FhBWBsXKseLposi/
IwFhyiNK3urjzQuNl+uOwSsCe6OU0ZphILtzpb5lEcrynB9/PQu32nyaPp8HeCdf6LmORDip0t0Y
IlF7yiPTe1HKLbyyIUQxDF2gC93q9ZB34jrvhIJPZVwMxoeUEyajVw7o+NT3kJg4mE1dm1oiURBe
gxJJS/TBPH9SZg+XQqHhBuRTtZhHqIw+b/6XnvlNOwyrYpqIjBBmUV2rb5+dNVxZ/kNFE8Py5u/O
SkkIkJ0OfbqvZeMVeYhU2nRd6rrv2UmP39WHTo6vgin+H7obD2+C4WTMG288XP3ffqeZ/r4+aa7s
6gsbd9JhcO//5SQ5jEAp50Apiwe0bdv4vy1JgCoD2an8LO6PjSNUaG3hvF9BV0WykIAFwcPFP84r
poj4qKsLHau7FGpaNlgq/rhNUwyHOuWKPwwVpz+Hj9sgqvNgWESMv+8w9JSrTY9fiGyp6W9fwTV4
QQoBPDqZVNzk+RdyNxR+KMhCD9JzDt4NpIoV1v6OQnrmc0H39nvXWEL5ZQi8mzK5uY1A2JE73rjx
1n72RTUjoF+pl6IEBes3+21lSnK/ongPAYzR07xxzzpoRsCHIGQ2PP+j6wfqpY/xqj83fFgKDbb0
2791srnQGAdiS5ettqFN2WZyfTpOEW68D2OxgWJ7pLedpgLJSSbVD27Htlyd/lBfClsSPIsFNpib
kxWvk+CB2qQRlCjTdUnhY6VWHYbdGW7lMBC02yMbAVAo3xOQaFljIw6QxHsTMCgrnQYtGkuQT7aB
A6xlq8N9nSKAD5YiXwcDtwlKTTmwa94uj8ETq0y1tGaQWRJCF3Hv+HwTfXw7sovSKKCxehIb4hvJ
RtgYahZb7XdF2psa4xWf9pE4FkXRYJdnMPd6isxeQtiBj/5XgaUxoWBxWdutjt422umkz4SKJIti
VTbYmDTfOt66F2B+nL0GhbGRskg3Yd6iOPEIPArHGU4NSVJ669yH3DjnIXd+I7ocRk3iKBL09AyU
SVYRmHY4tYPbFCotfcwKNNOVmcghqhzxon5Tts4xHZFGg/3ePyDZVpszSzgJg0fFvG3+8EyZFlQS
OOuWDOazZA4fSdK+Q0wPHMVSAxI4Rk8r78NaDuq+ysgmnW5FyU+QzRiiaGprNv/MS9LdEp9MsGBH
qM1GA4acI7Gg8aclIYLKkCcOdHmbQ5g7U0rQXgAdaR+4glmQb8MxbtAFSS7R/8IAMvNwurcrdw+U
zeqVbzYuGKUfaSGUr56rZ2UEKta+5qCBKOuo4AUm3QPKJMStmB39H+5axIifAoj9oAtL74on9ZOR
VV/IUn9jNCXo9lp70YLb3zhyi4jvz12MX4mVslHH18CmJDnxz57T1XWHuMIYtzDEnuD7SX4ZpK03
Mjjrhi+uITYQteqEALCb1OA9+Zmy2Bcp0nwjGvLalBcHDkwI588U8ifSTsv/YyHXBSJojXtKN42D
P/71IZChOMcKzqQoDbmWEcWy91kfWPhflw1bRWHIjn6TV5ZHFa4BhFfdqxW9VgVBHXs/asVwo/mK
Dq7+nryaq2AvB2wnGezzRARVmRxhpxcdgIKWnEpkHb9LwXzdGscQLVgDC+NvokYQIIr8VBl9I+e/
2Q+dYtGVPpoz5dh3TE0117GwBCcUp/z8kaZeujguqH1iZK/DPn56AFng3/0vjneLeAQf1w1fHBBQ
LGC7y9zoNTefoksaVhiUJI5SqsAAQxdGDkKZmzz4QPk4lbSzhQ5uGPLF9HdKVAAYBrkNREV4QbW2
/6cJaH1sKayRKkKu8SmLTOW733/8SdVlxiK+rfA/jIdyqOblujjP5M7Xvm4z5ONXeSimi5Tle0ls
P1H0EHP+axUuvdaIhYKi/bJaOC7JCdq7cZLW5uaqXjmuP3KznJ14db56B/LjSMtYxeB2lcVjdbY1
QL6vVl9ep+uWJDFk0dvXw0HmZsb9MLuvPFTJdKlqybPz9yp2ZhBr95d+Qxsq3S6zLqwr0ZSF/clY
bq5/XRmIRUOGi+7yXQW+TOTyeNi68KeS4H/iI/TubT4nGfix/jIfFUak4Fm6TtSXsXvKPrW2/2S7
eCH7fQ8Dwlc12HXUm+vZl7N0LKz6hbvGhnuyNhe1ED4e0QI6qatTdEJRReHmEBzTCjWKEqFPn+8h
dWZLwqjXwS3485w33C8CwJ9iT/BqwSqdxS2M1IQ6o9v5OQOnKmkb0l47ws0vhBepnqFv+aXbbL79
LjM7tBsBDeDCn4H9p/Pr/JGpQc2EndKT/+UCwFg52d1+N8FRsYGJooabDuC6JUd6skqlYef61SZP
xZIdrhXbHQojNxy1gtTngpr/034Gz/i2DLibOcngfUQkCd0UXgf2jadMo1PxB5sNrHnaD1akOmlQ
CnMnzo+u3qic7UihvvqPqr+mpwr60XrH/Cvidx7VQ7VzRP+mUgph0L9oeaYyVjGLI5ppFtiL/Uwy
OYdoy9FmbiyR189qzmQKbOubrNHK0YfuLFlQbSxPNAppISYlv7+CYmbIMbqxuldIhZf2vwwJcUHO
RgnEVHmBTDxG+fAkOPMTioX5ukN/Oc4DMgO0uTJEhbwt6BV4Oi74ZVVKRP0XI6Ycx6s1kfYsmVQR
sQ4uK3xNWler/ZQQ2PXSEoGBGAI5AEwfPCLnORpibVcvdeUO7c2+8VzqpkkxzvI2MCoY3cMIzolm
GnmT8QWGi84FEReRNGpyLcK3VCT2hvyG1KhA1g39ftww3/gJHlDKpRkcetqltFp3vFvmOKU8VdCC
jFKju4XvpcwgyCXkG8VStQFOR8OfkaQAmCze1QFrfWBMWzTz2q5Av/UQHQE0iIdIMHhV779E5a9r
xDx5vGpdBva9B0uGLoYGHyo7nSoNjRzvmmphw16qT/kPhL93MUN4PTMleDTjG6BpFpiS9mZ7jlM4
qAZO+L0BE5xOdc7CCCTXionKUNVFnGlUGuPfU8R8G9rtTwcMZbhKB8nKONVmzVb2ZPy/kus5HIvU
vkLQe6CS1UqeubAoLzIuydbx5h27yerbVEJXWflX9V0IyCI45jnDQK3D81QX0kHLQJ9bPRn0BOx4
x2mxdoHDo9w36GYvXu5ER4cDLrr8teVfJm8XRVKNcXvDLjfU5OyT0CJHVLXZl5MaREYssGcOhnzm
lNwcJ+2i0zkAhErVQUPvYo3KuZUR1lMAUPAg0lwzA+EgEvoDEmgkzcdpZvpTmDZeZtBGwxttvQcT
ZNYzcZYPGWWJbrSj/3hNofyvGyZSYo+WJfXp6dnC4KESI4VDF3y5jxQRlTOjRSuOoxZIJBu7YPPA
/71i+6hfbUQysUADD/javM6k30R4bLuiJDZWDu/el5FH1DDFix/J94RJW43IG15qjYz+E+AnVENM
09GGjJYrzFSpnbEFM4mTAib+hmdnqBWARNsm1qFWDjrOb7qFwm3Dke/YBDcl6zpD9hGuXy+MivDD
OgmNPqNFyKG9LZtZI0pNi8ArQjhF9it7ii7F5B4tKl8swotVB2moTqd4TYrDfQ7igO8cUrZerkGs
qkXl4ESJFP9XLS56G9FdM1QliDdomzPxQbfL9oTN+1w+Q4Vpp7yjvC5SqYdw9Au4/tRH94FT5b8T
CoGMg9lVzyGto93/f81ZVR+KNPOrNARDooOrrDQCURnKis8VGjxHWuZ9kWlWVyX4lulHfCxkHNth
0IDe49RPISqSXyLtEmDnbuBjHzYsBtiIuPC00xRLrPtT909XDUjsPC2HH92q6f9EOVPy6yjc/76j
Xgoh++L9A17BtUd1WP4CXkRc8pdLAt8ikZU7bmvaFbEvN6WnS9W/qdt0oZHXsZHdcjF2b16pGroo
zf214eneAxfcn0b73N98tteE7f93Hg/8BfdD4D9DNjhHRzAaWnsK94rYi+plNNFj0zzLO9USSg6i
J56ZZAnlob0zMAxj6OCxq2sdDUPGw90NYVJKz20KgvUHlsJ5IeFX/ySmL6o5GBFNkzyyqTO+X2VY
WCeAVuzryDfPXiMp/3ljBuQfe2zUvTFG5EBTd/Vpdr5D1XLGYtbwV4skvHeLoOFiwT4nYh/A1t76
IViEFAVm2RBaJ2OkzLLbbX9NuQLG9k84kH/ppmImmPCYCAu4OEutiszBmKHRotyfPVpCKUu2j8rJ
E1MVztM3HwL8IcgqyQAlnFu3E9oK3aQPWn3R9xxr++feVcjd9v6w1DqYj/fH8Z8O9nGJMvJo1yQY
6hIqaiVVoow6PQ9JvLUI5s3R/hB0dLhGs4zmgBc2w7HKcfsHzlyx+GtKYMdkiBZJrhMBpUiOONtV
8blOwtFhOVvKG3zuDPjyIeCcjDlJidmc6voDyjSuj425UINyI1Q8sVz6sj463wdcgxoDHVhepVFp
UulIz07FS9uS0vCPEHozhj5mALTFl6wZCClxIcrRnrrJLqJvRxp+7d2SlwXhWvKG7HVZpcn/KLj4
DmaZV5Zxqaiud7fW1B409QpEfeQCLsk4MWTiDUrfIREDLhZ4pDsysOtLsqJsVBYOgucWfD+el8GC
UNo5Qne9YrZNROZvRl6UzgTp0+Pn9x8Jo9hSQVB8EqM5l6dzAbbOfOjWfIg/pjpuhTEEg2PokNe6
Z561QbY0wVxKISr7pp/Xbf+rnpT9O/i3fN10jSn1VtMOkE8WRnHAlfbHkmDXxVNnQ47d3YqyhwkA
tpCJaMfN/ukWzfTQA0mwbeEZbSOUE51NsZyKAF2swCSzOwlbKpaU5UNwGXTz83O1BU/rPMsPytT5
n1FrGtpr8HuwPkFUCYJCCxebgMDxOVjR2PlG0bdfXSrMfvkB+SPghM/oiGU2vIV72uclM4pzIjcz
dTGUa4BbpNfuLzKaMbqaSI4aeWllTbkAhWzv7OklerNYJWx/lorVn3v3CGylgUIAz9dWmryV963+
iBXCPag90Kbf8RNVQ+zepro3uvP/IoRkJNWRiN90yYuwHT/xxpQsmboX1X78xPyoXm1Q2vKfpcc/
0K0N5Fmgo3eOO9k1SIj2sVV4RZK37JRQLDRdHKqbI6DKMiXx3m+u0t569GWmP0rZ1tQD6WtWbb72
6N/gYLp2+VNdAQeZzr7sou7hQPWk77/1IFz+P66EJz5dEozcuP73I2ni9ZagfEyTRDa4KFLUTAWI
yXRmDZ1GpxgO22TxXkGUXYHNrBQ9Ck0afYXgxk7AAvyGDs5+BDK5tDky/sO0nXPwcXjtKtZ3r57E
8e36EkR3zznhL0ZB3gs0OnytkIZb52tOQxFBRnx9NDLxUFjm2vBQg93mDyorrphhbbnfY72cxr5L
uBZse4Q7GfwQyiONGniXrvq3+dCLCB1TuZRTT0KU225f34RoAK8kWc4QSv7NZn+DEQH/UJqkAKPd
jW0F4MXib+M5iqRfKkpIoh6nlJTH5B3lWgcIq4Bq2wG+lwUBQ27YbyhTWL2hoBRmo3WeHARLIRma
CNy2TeSbhYn2fgpxF2JmlCCPflN+ufHFVPNP6y7X5kug2B6O10/Ecu/uTPS0qyCE21j2ZFgxywZy
pLxQI7WxCJML1guWita64nQZl82zNNk+z09yv2wb9hBlNhyYXv85JZ9cf15h+Jm02WhpwLJQLEnE
If3kzwxF3sntv6xEZK7LOoAJCfH7JlnbRKeBteYu2rNf7DqPSTZ/lcZy+BoP1VsR0R/ebut1hg+y
ptt6x9qLojo7ukWEkJV3AcjN3LAw3vIhcc8D+pd7sPX7lBDpZFWfjUld0njm0swCAkgG4/pLYZT3
XqhjOpT6+KiOvbH0kHMgaQAqnBBElFcV7ZnwHkFMULNtQRv7NIPBxOyRUDNxQE+OU01H+b0+KEpN
equua8gnJ9P6hNob57+i+fjkj6Jw0sgB+rpcUYgh6J9zoaEbkaFM/XPW4B2zOGzaVGi5bL7yq3o7
OI3PXak3RQ+mYyidREsAph5iVBfrqW2Hl+XtxmXEL/mjbpNDlgP0Wgoq70W+6m04EJvjBB3XQdU+
ssTVs3NX5GeIb6VX2w1BNCZcp7JJXUb6NKNTg7Q/EHzi5EQ+vGf+SNRrOIlUhsdSQ9oP0ug4SJPA
asNPMeLvSAiaEJBA5mWozxRgGNMjA4B+iYbkj/SKg+eoGKlxki3vO0+ckdn+r58Od/uh8oSsYWpe
vD7R1v9Oz9Nlv3jnOO7coGM6OO3iaTJmbDcalVjaZTupqSq016cFOiKIwRQyFyA+dknqAaFdKRnC
rE5UjPn/+iDATYD9VVbhOKjY0L/GVnImUIWPbZwFDh4jWPKe1Pvxqe8OIQ2WgzkzZhpXZ9V3tIKE
ZaVUYpA5jwmsE95/O79BR6e6e6fAyRvsN4qCPvQWQ4cArSuPKVjwtH28TthLhBlkrQzI7umrB7kS
az0hr8MEoeUR0I95vSFBQuxfYTBcZet3lQQxDcgiPJIK377WzCz7jUDA5FCofWojo0BVm2UGZpo0
fwUdut0Ifn+eGqXGOnEV/u+wx9fCg6O7JR/xtM+Jq2ceuGrcmeps90dfxsom0FVaNyLPJhhsZPH2
MiFnJ5rVYk1h7KlU2V+3h9keR6Yfu9NR8CyASf/DOdg8obRILkqyZFlw7x+bDClU3yu7tpxA25b/
NdnxmVDL+bmaM4Bumr7d+TZW/hVoLiwjM1K4s9xkJF8tUsBlGqgOOm6yN4AclAi9+bYAhlQD0TtE
mTN/gMilTt3bXWtWiTrgZmK6LeIocx/8CR+xqiUJQdV7KL3aPsDz0GYMlLD7ySPs7ypUxXQLvrFO
ffPKBbJ6iwmwwcAGvW4xnJ+zXronlYSIiJBBsEp3M3B/vmj+idMqPbI4hFwDrTAiMxj0GHN+qtcZ
ht2SRAjzJkeOUFP33pq3dnZvsapKwYZ/qQhyyTWIXEX1qM+ZU4TVCF6Q7VnxwHRsk2GtbMfYfEoD
cpII4bbqLWzyM0floyL0AB4yjGnvwpbumZ4l/pxStinH+tYWd0ibfjMQkxROBRZKRm6YlIRJGs6B
TxQYEvNrJjnp/sGgP3Za7dMH/TEEA97s4mhPt64DME0ikxHyX/PSfGAB5CoAbesLzFctMie62xgS
U9PHcq4Ite8G6tmB8LoU0OdlfFCuuIv1ZF6PlfX4tF0wOGR9ZhZiB3PoSAhcUBU86fOgKrtqCkGr
r19QCcvx8n42lh/yw2tGOlk55s8UjmgcNFrQaxgzYPqEKt5CS3x93haHSHPJDvKBpCBDT9jpVSPT
QnitqrHnTjQaLhbqQtkv/DQ5DxLN1oxfDlLr9QDop3119PXAW+VoklTmWsWkyGgatbVnONuQZK9t
eE0R2lXMqMAMV6pifpwpD9voiKFf+ZQ4S6m3zS2KpajxFnO6C94gGbFUCU41l5U87CfKXbjnzrIs
zPQVbXvfCLGowhdE9p+GcN9bslklheRP90C0/QQYei4jxZsZO7bfqgr/3XvRUroa4Rimu3bCiV7B
1CSVlQqj1gSJq4nteWHl5pw+qJDdhZ7V2Sa6hg3kuHnGD8jBkunSNyi7sFli7CprDhqepsc1qzLQ
WF33R8+J6QPY1gOPjMytB+85FRiasJQaIkuB37XngZ8RHKDLA4VRl3F64sH2+CB2yrbLl0lDq05m
P2ooZnbX/2RUu21tsqSxbiEUbexDBvPnGd2PI/IVDd6RvWPN/TCqDhZxi9rrREqKBmXXhQNUlB9m
PRKoms9JF9BENEFOAAGHn3TZ0PMWQ9yrFx45v5TCXiewYBrPErdhpfs/UnxpsBnBCGpu9XujkDdH
Bm3iWCe00HpHZkTLv3NquobTMrlC1SibnXIPFru7uJlNjWboMWjpmxLZx0oczS1Nrb4zWzEDB8N9
fghfDlgl4qDpIcluxbMm1my4ebwRcKyRj9mMhRjd7wXBOevOcYgiqBnmV33tV1n5eUwatXAuuYKO
YzSPj1IYSkyYq3ulaH1oXBJWKLhbq4GvA1xRJSi1+sXyim7FIn4VspEFT7IWmmLlS4wfrnOSBchq
JmXgaoUF1HOr5v12cWaQkKJYriNI58FRXsk4VQmzo0iu/cjLEfylq4Uxrznap5JASj/QZY5++piq
pY5QkDgBE4f4L00Z9/snUgoSw6QEZ+47fQA1cGOFyicGi/ueVPuD3dBnmcO3QWzZMPm4X5CMaeC6
ClX9YVQwKC7d5d8tPW0j5avWH5vY4/gV8KxdtALAmb5VGgHo1Ql3rDDVs5/f6sdcSTUxPfuZQdZT
8RHLkq/4RpT6SBhmwWDDVBKDhT6kVZYd0NRRIKMRsCGMGYHrMHkuBN7chPNV3OjuZwC71rH2n7Qy
REpmtC0DRrSXn1ybBNlnT4xd5gN2l3TBu/74MDyU4oFDs6wfW36IUbQqdhxHxMjRBV7K2BobKaT4
VLHdYZvibY+UqbVWHei/VUDv/2aFKIX9+N3zE0l3pogjFas4kFlC/EXIkZcw+lc3f6WBAu5xaOiS
BxF15uT8upM5kKocbePJVt5/+7+8aBXOPu0alAn76sD8xXE5yW8UIyI/p6jBDIxPB7p4oarPo7Ia
V2ZvXN6ofXCXLsy+V3re7r8PPmhZq82BebYKvYtFVUyIkZ7nD4WtBKWVQMvDmPVuDqgP8Hu1Y6lu
xp6oE3NXOa+Un/HejL4AQK5UcFNYy+SvvtE9yB2yBtzl5Y61QM6QwxbO6WNOaVUQiyFlibEwfRNN
euLNp1KSsP1KvWAVygCMalPXklPpkBi8PbbikAra8ZEJ3s91tDyQmwn6k+qyl+1ycYSzNVh5dSRw
owgHYgSQBsIS1O5VRPCgBg+7wlMgX2CreyFa7t/+S+FA26JbUuqgiA3Fse+5lTl7avCcJnrhWUvb
wjbKwyeDh1ex/6xu5Q+/kr0KWeB0LwJ5JDfOR2nE4zp/dXTAWC2tD3nNolOmhihNQXbQLs1VqJlg
vFMMMvvvSGk77MugjZxgAl7HMcRQ2ve2UVsqxewymobQJgYHswDW8n2AVpHlenobRT2/iQij6ai6
Iv0Up+sVwDxKNcdDaWyRXV+YYPHAKh5oyfg7R8jAbAD0r5NBV1+7YJo0HUfkj0hqJRnP48/zxA7T
tic3v35PwY/2xI8y+FIVDGuHx8lwcGo/FcoO4gkrpG0VHpVJy5sN5pOFe7x9kFyQhqlBsfR3p/Yn
QnNqBeu5hiHhKj+J20h2eVSwQJxQScS9EINSQMGnZszC1gfPyzv21k3PkPoomtUwTzCNL0EVIBH2
d8wiC+zDoUKWWbNjAoyCImgCi5G88jymDRPb3hu1XQbT/imy46KwogcrtUmamV2kgC+SwDqcmmUj
x3za5etv7GUUTc3odjAcDAipw6oBvBVkgldRBdyoepOJHG2OTxiSVgjUCWxC/Ow6jHnH7vZ3P0ix
/vYHSJJYS5ZFJnJcHtzFRspd9yH30GM/o5FSFQLMpDuoUc8mYJkEyzR3hwBrEtc6MVVF3N2AY9/S
yiQjRFKJ0/IlVcyWTb55SAeZnaY5KIhnm4QCYjGCM6HrOPNzD+0P6oznOHuyQ1T1bfAl0g6QrGQq
3dzsQ7okkjSgTe9DTZJT1jvvblpmyL7w7oF4HbCb+eaMTisbtJVVyPmrIDTGaUazX7nKF9UIcP3K
OGfrFOHPK0C1QNtyEO1uhQqfnqgIeJdFzNK+hzPkAR8chQEwlCg7eExFzUKv2GqGHduJNdQ73mN9
/yKRXCKf/p4FFHxJNY0W8Zh17fRRyXKnW3BHYV0c2wGEj6ySnIBqAcbnnldConEfokQsrPSN/+XW
ysJNgi3s42wLY06tgmhMy+lQlQRSj1zj0LeO4LnavWjrXm+9SJZKOnO3h5TgEbAzCYiP+Hdpr5tn
kPW5ZoL47XcZ3ZTI2F8/CoGIoE8PRey8JfsBKohKdDplf3U9eIBph4HPAZ+EVnpHjuIYmg/WrLxo
ZNLyau+Fx8KS9e0HYUUbiHWYFpM2Uag3RFzxvWhih9JIbeIBbbaxLTf7CdthsuPLNcqquR5y364u
cIR5d1KHPuaTueWhIva0KZZm9C1giMPTlCaZzIk92V4P2U0rNF/G8pHB8nm+ADsjO6zTnwzC5qEJ
1w0moQKtrgOapNMwAcNEJVCoVxeE9MGVF4zD2LtUGKT+g+XqEtGRzyiCgMa4AAa/Yyu2R+pXN0qR
c8BdJqJkmYg26661LP4NbpoMnUXPk8m2fPfFEcP6ntgYfiJhD3mcV8ohrAYNVBANiJmnbhrn2tIi
d5sUB6VQDGQzJQ01URFqg8QYaSXlI2tYyS6YILMVTSq1/ahud+N6hh5u082cleyQl6bAUK2KAcLZ
iTyvoFc6opMt0gsf9VZqvtfLu39ZspvAtPTdxJ7kKnqUTS0VHAdE8E7QI/c27RBacsKuBOiUv96B
y7dvCQP/PqwDD5LFRDCKS4Xd9+eU0jtPnPA/2evt1rmJP5ChOlIxKIcjYSy2LpuppLjWx++V3NZX
1D2dPIgMLfEoPtJVIw4FlCKfwZgtgKutS76PGcr9i7zTFYpfz4GYJae59/bFHQBWVvHK6wEJe9LM
Kq+/Pr0PMeym+7l/ZbqtUSIU+RAXsvKsY7upWdzz2rOXl7pHsjfOzYU+1Br5H2VeMEhCMnT9/BEg
ff9oPSfOzsmSw1YxTJghmwPbtzCP0NV3okKyuz+ru/7B3eJo0P8atsEKlYA+PhPnYmlughFsZAu7
fP1nZcpPEpdGnGSezZ567bEjdgTA2jRdQGkefEtdwieIKaGv4POAp26QrNFXKT13VeV6Qx+clEWK
k/V6hJF2ODj1jcBNPGvFc2tjXEn7HVLg60vURn2iKoPi77xbqssM/xsGRjR53NnUpO/G0dhnQmQ7
Sirr+gYqX3RtHX7llmvuzljS6KTZ4mQ2NskQzLcHvwevcGLdM3kw/tK7/1cIYlx7ZCw9sXsjRP6w
obNAxVUS/fD7X8KQJ15JRgtxn2Qx4n7yGRQGGa3VmbRcDGrpQSD/eaK/Bww50b2+DejMZ5cnXr/8
jZiXNYP09io+zHesxj0ubX+Zujw4Kj69wCxVtIsZzLXgDajSe1ld4fFCuQeah3YBJX7ZNJFh2/Xc
uXQElgFB1zVTV4kfl8t9K2f23+sLb5tOs05YkaYENzBTngO5K+LveqzaHrxl2OI9UJL0vdtIy7wW
bjVQosQAZ58330Fq5BXyd7LSXQ10wlwxU0HDDVhP/XW/TZahR7cicSrGvWgm3MdgKQN1o03q8UgS
LQNULGg8rit8aa+NpKBupZKzNrnMRL6/j3PdIT56vdW3FndETnJFT2slCQXcJaM4JRtV5t7KCqxl
XfXzwExWJyyqOiV514HR53ol2/p9P7/Nl88y3SOjV5Bczq8VLpTEYjYyu3wrMMkc1mIbed0VGw2Y
VOlc2/KVmj2hpupYdvmOT3P/9focfSjK7YnKJ1boJhsxjjj43uGtdxuaTA4CxPryhsO4GGHBNiVS
VYtluSBJzWMaINKynjcog1+Lq699YkEmLo7iBTCUCIEBEKuOsh7QaXETiRv5Vd7SbmHiL4ItcJXs
MX0DhoaQ3kObuagevloc6gw9slgYC6xl05QRnbkzxmoHsqy+WOL7Hl+BTC/i3tTKGP3xEWDJ7stw
ldmiEaR5Et5U28PYfGj/N6GKQ2LBUzem1TKvO+UMDB6PB+KEZtpEeFzrO+FKyrCPrnbptY0umh7Y
R68+wSunHi/tjG7fb10JjYW8e3TugJT8xCcV7iUa/oL5Hpx3NGCeqAyZUt75/WIM6fETXHOqrdrH
oTqh9uzdSYykQvOlYpUPd66l8GZhRBw6qtA55DWN2zS5RNl7vcMd6KJShUlF8D2F1NcPsKJON/f3
zxVJEMM9S5R8LSm6pp2HSJNYraVq99OksI4uwUGz29GLNG+LUe61/KPKpwDh8CkaBpyKX8nU4x4n
rr2rx1d4PLZ5DQiN3CzHsNpagSy9hfuk5O8oOCHkFyCGLMaJZxw8NGR/4wfU8Ag9ixvp8Ud8YW+8
9rZs3IHgdWEyIR+c7ZBSKtacPQB9SWP5YiJZvotfEOWizeMd8UBKKoGX1MyBjZ6ahmH2jgBxM/AF
aMbX0eFTDIwQveM9HMJaYJs/VOsubjS1eMhtW5ZBoZpfo3x4B3szdvtsN9LHdlkJkKkc/kvHzwk6
B4XcmXi1/Z/3Bd+/e1kWUcRPVupBVWH64m2mDFEd2VpIHz5wc5x9sWOg7D5/mFMdyqdWVF+SEt+w
GXq0na9MZ6mL5Z8rQCzeviPeQr8bjqJji8iuI5dVYGRnlN6MWDIXr8QWDB5CmZWz/Xrz+hw0f+/w
OIKtmgYEZLmXrYtIdIPRTGm6Qt4GQdnx5wEmLnpIEjAm9ywJ0mc6eb5wKbAZjWy6X7T3d6leC04Z
0hsa6h27FAm2lsoufjJlpfo9TXeWiQK3x6hGzLRRCwU7kWzy8kFBOVOXulYcvOuUCKAMFrLb7XkA
muAjpBBT2uG73HVi/nOZyXInKNa3vVbC5DWjjau2kX7ZiHt8frM7PdvzcVEmcosF+Io7awWdBLG5
Bn/FIXzIXsEDQa6nEl/0AmwuNLQTXR3SwXbwAF+JaMLHfBsTtUt6540H/5QR3oSHheAvi2YBVkI7
haC0+o8xwo45qFAodJJDllI+nth50zEcwXKLImVU4+Lco81lF+lSggQqC6QiFuJj3/LmGtdyxwEz
U5q3B6bnCptsNrdjZ/lWZ7bYpDacEy4dbnneqN6P/4u35W/277r1Cjgtl/W4zvnqjynL90sQN6Gj
D0UyRTWTc05SJ1W/QlVZLHFun/p7v/PJz76IhPZI14IMVoCHdoRaA02c/poGaUg9iqlU0xW8foFq
C7yQw6avv4lt/CQ0gjuK2buzKRMifaVIDKDYpMydTJthh57k5r+671HraDiI5QMmyTxTALM2Ar9D
vqh/4Hm/iIiGnDgQv1AGne5UKRadHS2+/7DsowvJCtT9jdjRKnA1aQBcTdqmGPOqmKkd7yh0iA7F
kJ1J7JINPF31T4kW+7akm8sZOjjwuP6I8s/74cqv677oed635Y7Z5xP02cF9uU0O21TLzGX9Laov
V9sZDWQfFL2otXEnksTAGtHdZTlubs34AdbaQjm8YIPHlAcpmasseccBiBXBrSU+DAYMpJB05aOM
p7+FxiOsLbHXCrLNbzLFepqgDbZCjuobHwidOiWUSx+LJSOzWV5liWiEKcvWpCLZ2nCI1AWKrGE5
wz+AFiU4g4f3l2Ga0pI2cewGQLavSKhnufseioyUi7yP9PA4pS6V1/Oj77EUhKZ7o16qTT9FjRRE
RbRFgd0BgIH0h1nYNeJbrZmS9XwIcCzCHNhmVrwQr5PdS2iTgr2yItA3s7eaO3pf7+lDTB3H1yC6
0+3/yy0aLcOP4Dg2arxsN3Yi24OYwVSd0R0xwwtJE8tqT74YCXNO0C9X+atCluk3FvCqVvgxQ23t
frYq68jc+DxQsjHDfxFbuIyr0xLhEd6+U32JeoJ6BfRRwmuniZysdYPHSwB2/jC4XK5zR82YBNZD
qkT7arLUYTUUkceDJ4wvrr/Kdx+Ykk2u/bdVb0Hkzwxd3RCpuzalx7ewJJD/m28o6s6IhtxLyxeq
Q6TXzzfmV+z6MWask8LLWSo5Yh7W1F3C9634XzRFWIk6lQe2N9nOhuCOdMmjU6SCzySYGvDNTQvf
4DttekXcwARG5LT8n6YCXfhu0RX49ueBX+KVGGa4uEfqRbwm7GWZPfXlolIFj8F/UWRyGLxD8Y/B
wlN7O21CD+Dwgx4bdx6oGNby2bbEJcdmrFdFdvqpYOgjwL+srepOrYizHwLuhbGJaQbTpDVRhJuS
Y7oqY3D1el9KPYQ8Qk5TLXL4fay8YdE5sK9xdxAQHUjjZ/nyvHjbHY2W8XGpGfToNa4iBpw8C04b
JmjhV6uG7C5xagFbMnHFSiCLmgraFomYckl+l7T1SEFXZeh5tbAeXX6csHiq1a/nviuVPcAG8S3T
6JjVwo/GUzkrX2kBYr+wV/iRD1PZydFhM/ZARDG0uwvly3O4WN3Gbb3izn1D8ZUZWELeSPwMuWwq
I+iTQ4vHX3PkTsNojPbLjdD9w5hzH7/PKA/77wPKjUUvTUsdiL2xpuQxVEAUgUBQCsCWHbU1blr5
CC1O6bBDCmYMpjoAi/bbiVKwZQbWeGnTMQ6VvLck8Ra2m/infX1r1js4tsqeGo7VfowGQjlTAXCR
+mObjk9inebOOeNWjQYh/ZELIASuP4FqCyWU3CPzXTE6ACd64YlDbzFpCYecWWlL9nl0z4A2Ws0F
jjdrLQ7lkW+1IWSSVMF/QQMC5VSWlW1sgaMWl/723s7w8X6OALfkH0yAAL7BBZDXNgVAT8JlO8/h
B3GyowOUv8kAe50qyf+p7JNp7LdXCM9HiCUx1u5YdKsbj5Hs79+7LuPKuDKrIM4qznj+e5lWz1ja
Bcg/XkapS4Y6Iv+whjs7VKY57h4Av7whAu7hixHZq3yFBW6hoXOWctHKCHCov+NEBBfk99UC0PDd
GRtGsVL710HlwRpT97uHWixEkV4DFnOlBa1G6lZHq8hNdmct9phD2WsWGVWpoZWkAnkZD2TLcuEi
3cGwcPXFHNY8CwgPF6GT301SuxTQQJQGOr1YwGffpNssOc+OA8BgPo6w55qThM0pQRKuTmPQJqDc
CPIpQwzkVShBFlyutqdIXa4A0jQxyVZnYdO4fm0I0T8lK8JLoYRqlr70gwk9ZOLNNvCNII3Fy1Se
mq5IpsAfCo6ta+3vlDgkmA1mMu9HcZbKdAlUg+ZfRZdhxeZatMkd09XJL3kn1rp65aPhHruNah8E
IjEyFZPAhoLpwnnhB5C6B2+4VLNpaSjBCufgM7SSx6pyZrnQxelS0FTEauWbg8+PmZu2pf7ReG2y
7yLBjCsJtV4kkhWzwlnbEtwUffg7ala2a3IJHIRdtvvRlxX22MkcIyL2WfF0+jnzf1wQz21VPAl1
3ruPEnQ3pQnfmnF88oi8MEYMLbzOw2hA80EZWd/xMo9Lp8xA3/wxR3YS2b+wVl72BW5xmSpCu3Av
2owPZ0dL6hm1vQ6rVyG0ICNSeEmA78E8AT8VdaRT5NpDcKd82OM9tUM400a8YBJkgzghEmzjCvnH
GoPeQrfngqZbxFpH4IeY7u+nMIz2IaMXzm3m6btUAADVVXb0Rvj7SgLJORIcn6qMLFBj63IvixQv
KA0OEYzW8F9sm401v2w+xxPX16gPrbwdlQO1wcdwvLpejXj4NgwcvTqxslFfU9dzL8ItVwk9wFvv
MgOcsTTnIMaU8KnIZIbGlmmj+/ONtagd8OIHFOa4iz9D8aPhj9K6HAu6GfLtNdxw2et7OMSYXoXq
AuNYlmFDBvC5wcXQqgHz9jwnWC8q9Q6ysfattbAp88ivb0+T0l6h6uVveUTh0H8R4muDjAOPrRe4
ZwZvNMzJ7Kjk1DGZKPhBePaBRM9hqo/qJStBmPvfw564gEcwQT9kaRffvinlFVccSRR4v8flNNME
AtkoEBBY8j+CPFkby1LagonKDs4Fy+3tnYNiaRHx8UIIaLsSePCOS86fgmhopdWu940Js7FFlpvz
sbQ4Hye5tqLbzWyc3bpyE/Heabiy3P6nN/gLc7lwsQHmXsWVPuvOwfqFzI3TQkFrIbW3zaUIda6a
CncBP8NAUrOlFjT+l0vtBvzMLMdmHO1GFeYKSA+73+7QJWMcslW/7GK+9rRqRkl33U4f+iKmLgwa
hmlGe6SWyr+hhrLfdRmRts6aenP4fQoVx03vleXNkOTWmnlzCBoLuOVxqI6+/sD9hA2/bidgSyj4
l77p9P5Sj0c30mHg8wZMWRZiwEkbLS1p1DBRSoidfaT4dEh7t0CRn8Sd7/DgwvYBa1ykfiiDAsFm
xrP84NbFMpyqbkbEiooO+9geFdDScZlehKM5S6rP2OoZYpou1D3Jzv26nu9uS2BtLdOQr4lDnJ3S
c/O1Lcr3pGukgH9jaK1wcNtXliUjIDWQaYVHJZ0Zquu3M1e0ooMdBBmFoXb2TywCAxxUjLJoS39R
OzIBjW9j/yPXSVUmbU7Dq5r6xc/A6nFDipJSnKYjpRr5PHJvLhh3UGOPHWoK4BjfPg+bP8K7l99S
Xj5GhPzsoekOTSl5dAlCiIWdz6CUBwFg++fP6QEyY61FAlwbTq5FNqpqL4QejCVG4q5PB6yuo8cb
p4EP8t67Ex1uhQ0OQgGIA1VBBfCYpuN5Uocqj6+2a+XvuyxbxVLMlC2GTd8zIc8HcDzwogZw7/21
KCjx4l08ppJ/Zs7XzOO2y7f8peAhjBIC/2wmxsLoBLCmsqx7Ce1ohFCdYXy7z59AJGP3atn4+mWQ
hQkUdXBKxjg94JYsh0jWEnNkhIPbQUY5DsAB1iNKHb23CoMgLj7dlkQHXGj/bxHtKdbIZYNFqCnp
SawzIYCHfMlwCYXHJ6UAq2eYqiPRtMLSr4Pps8OFRs9wieQmSuUuMBmyuGKzTbknpewPRiSGoffr
9yt7f9XKmZ2unGrzfsaDEtv1iOwcxhDQ5Eu1gGV6d39tS0Y0N67MRSoa1byFgEhYhw2qPO6j4XAI
9Z0MmlSY8mypjGB3p/yAuByzgDCB6LdxkzaDS9DAmue8+YHwmWcG13WijD0Sl+KPEqbJ/yY60ftM
kfN+wJuZkb24p2QjTho+EFFWbsaZUDoKJGWlT2pcGp9+OyPHGV0UrsG9QEtZ+dr5rECvRJDdFNEM
w/F7/5BkWaLKrFM1KQMyY97lSBsMzVmZUdS911Ga9FVYmWt7DcSjLq1ddaQjk2QvSGjQtFGjLhXY
4xiQcuI/F3Xi9gpv4jVoOrgj58z5hyG1P6/nXY3hb5pjWeTR9tklHMQAbrj0eYS5NXQIYSsVctpo
x5m+ppxDTC97bTLEKT3wSuGoHxZVyIG6U5onk81WqyX8z5y9iQAJFQPi7igRyDqhNdB+mVzR7/WI
/3rKFVaxSaLF9jkkgCBRK8ZWvAiSksKtC3lRsrHws/LNKcOfj/Z9JzFczVrz8CL9zfxp+VtwagfP
2SsuWu41PImXyxbo+uNtzU2XOYmi5bwUMS6CP/kcxirbwtnaaUiV35Rxj+Fu3Q7wYzeCbNYbDe+g
R1Mta0NV4o+Q/VF1zWde2fSMriTXm5n8MMwqHG2H4mLfV46tj1BRhaoiUBVAVLOB8YojRFn6hnGB
sWPUzFQyav9lx1m0jVNZFwkh9E01/SJefgrgW2TlNeMLo2FpxeYgFve9PqF6/prvEx8pYA495Spq
fWSL0u1hamb39pbJujkqNycebHA5AlpPPN43HSugiYMw1O8blShhRLs5+n421r1G5/VXpoNTZVLV
pBt1KinjsDHVhnk+AjbzJ/IfW747EMTifBKMWouOo4Nv4HHbtMgsQ5zzATTUaAI3aIvAKjHIe5SA
C9nkfbYk8ePdjgsoD0pM4Vgy4kooE+P5xltjmdgkRSREy9hNb6XPyXk1uIgtMYtc/yu7PZKofHY7
ua+BqdqLlUHg27by+bzbmEpONYDeiIB2vCuyB/nDAJ2AwJkddmVVrffsFOb0U1cVcOtrNbNjQ9Qk
jFV3fL1AgbcCRekzaMPWN0QaHuRfmv7pKJjYLZHD/w/XpzRA/06nXvA89P1yR56Zk/wph7stXTyd
TQ4SL1RDLkxECDUe0S9uHsDOm3+ap5aEhdcLsVLVBmzTTn6LHmSJFnA9yu0ffMwp8VjQGGXJaRJv
8Dc6zkKxaGElhYtwvOhW7pjHj9YWFUzAJPnLq2VTCkSe0ZFAEa/WIM3bwds/sQ72NjqpCAbDzgMY
6onts3dH7l3TbKkzljfvP4xET7KFbk8/765V5ot6zFnVbylLr6hpcp6bEP2WQQW3qhd1/eoaKR1O
WRk46sivgabl3GCOIAh+nVqGpIE7nGs/W02GW4EOkdzZU+LT9uMiBXaXdqderiNDuCLeu7a6MCja
shUejkNC3VT0fIybd7uK30n/2ys5TaXGhGCYJq8ghKy1/34o9fF7+U1h8UbipURJ1erdSTSdS68y
018qdqhb8eIH+N5mZ3YSqPCEnMG18OmmPDAUCoE2cUCpg9KajUPDL97YItpYOBm44HkxHJlzI4rE
IvOP1p9enRRT4fgjOQSa25xYCjcaRCibH9d+Zi3/ZT/jxV+xgiBIEk4Y7y38VjlbgJS0ZKOaP8sv
FLtGUuWpCPbTeTzPzQh1RAytc5ko/7Q5oI84QmFbzoGsgHQDCbu/L8UcAo7lSxnFXFn0icGfy181
CYa1Qql/rh3P2rkk304jylIgdRIYBEWcEgmtwNDBwNmuRsGWrTCbPXSllPSOlb+gBZPlGlRkMead
p72MvJqcnyAqxgityneo5unXAALbx60o6f13phP4enq8OMRnyb8KYhNvQwFFUFnktTDFgYzXDaWW
0Z2ye1EJNAl3orUrPuKnaeyNXs14pJqzKa44LiOK/f6NkOaBQ0JBnltwgf/cgw1bKo4BhBxsoppj
7l2WnfuIPWsVxs5wF6d3BOZfWH6UjeJlKEdAaz5ZPWeTR0D3Dn4TB6xJ5av+SF9aXFxL64+8I4/4
gDZcWR15W8cZ2XVd9Tit088ihhj8c8NrvRb4EHfDtPzEt41qMxbfoOINhdBBPZkJid3qpUl0eMJR
JyOWx6D6HMXX5WcqSbOJFZcrv89olJOZfXzqIqXeaGbBM6Di/cMN+8ooJ2s3OAke7qPjs/vSJtS4
F0sWU16zDx/UUZWjG0Da8AhoedcVVeYFP0khyMj9ztrIIUU44axtOo6peY0OD9xCpYiLqTUkrrmT
lP3mFkW8iezCsOAU5iOfYyACe/XRRFhfSxqJHo+KMhukCOdFZGuv+0jk8MdV/bvnGypMdwia1Gt2
nKoenAiNVrpDVI7ZK677upmrsW42F3h2rM8H+2UYCHM1HR9DyuRBYQOXEQMtkiBWIzYNPM+UZvVY
fh9l6UgcyBGAUfd2UllmisPECaMqsfIG3UGUeIG/MMgO///T1xxDijiwKvrfCRi+iv7ejda04aZv
8zoeZHWcU7bmWQtSPUSSNiPmfnMGU+YWtd0tUiYrFxch7woxwe6eQfKFNcmbKMS7mq5ENQoplrZp
hCrfQptnZhFHisJaJFh+5Bse8x6U0r9APi94YQUP1p187y/gez+Ts1aLB05L1PVU9c/yWQAoI60I
KOw0R0q0pdCQ27v/aGKTKt1LgFn1mQ50TnexUNox5iQh6vHV45r8s1mo6ga7H4g2ExbDq3Ld2d6s
im8RXTb2HCT/dbTXytwRIn42Ddc2G4vx9tv9HD3ExLG35iW3dgvh0YNB62mWc5LuA/kGbksX0wlp
0dJfDgdMQdrb+cqjP0ipkeJGMfmkNtO7t3bkzDVXLOn7QURXoIAJ+/2omMy0PLJu19uAZrH0Q7Jt
hEicvt2nlPm7eydcn8BauwTjXWghB/dvZdc3t2sfSFHpRzHTlnK5rrPCF7RV0FzfZRooFcFKP1Q7
uN8BEKap96u7FKY6BmzP1CWH6Yl6LEOAXBLDl/oLMZS5PV+SvSNhQ38MNsDgRHfAJ1uDMXrT7/5v
8Zu3pTEoD9MhhQWEHuL8mXqvmo9KFuK9eN3ogFhE2zy/eGuTLin01OowoktdkF2i1sIuTeqZbKJL
ZJIN6TEf6VrB3VftZDOIoF5X64gnHaFhASWmQuZy6rBu3nF4waUG6D9YuGy/kCNUr5jK7/sBRPd4
fUQM3oKfGRTDwv2YbttcsFjAm7uTGDUiuDUKGYBoEjVg1c+UfI5utqO1V0a9zM1JKujp+X4=
`protect end_protected
