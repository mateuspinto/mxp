`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
OX1Ci8w65hys1/l+WMj73kmlCpklxEnE9vvP1pL8TuGNP3orZBiFbSbo3CwEP9xtMCrgC67XnTx0
X/ev4MtJnTT9ejjre7KMlgoE4Uu9leJ5mGww4rkq1NbAvyttlnUadgYTYKperdO0KFfqCZERpnKf
ABH2UT5+xJeY52VcXuHE0/FXSpZmFZ7aURD3F4jMckmIqAkvdVdLeiYvgvRsytMHwFKEuTvo05Ib
Q19PpDuWMBSF0juXuAdVkaXvLfgZPqn76u67HDkrWT5u2hD68RlEfIRlwt32OBlofg6PFRnshj37
SoZ7NRnsjfuk1IvGMKd+9O0ke0usV1BykQe/KQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="+cNIegwFpigqdWbCXWENKIGYtB7iowLo/dxI10wqpao="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 93712)
`protect data_block
ip9gFl8L2k89HyMhOrMqsonibS+J1vIToPCQVOfPUGZEW4IlqsRjkN/NfIWyH2VjoMYS3PaJioID
8SIVHGJVM/dyVpB+nUQKS59B2f7jxWJkufxkucZvmlrMNsUQT9OxOMYr02vKBsCg+hQ4bVENjnr/
2IWUR6izfQo4g197+BBxBXFOVetfJHY/wlor07VoumsBf5RIrraEEYXjmKv7QSU0yzKOz4qy8/HD
bnQw4RhbXll/bL+RZHp3mUHv51kd52DfJtUTGC0p+UVg0l9GGtPeVw+lKtTSwKOQTeWB+REiTWKC
Yq72plqhKt55lAU9nqTs+Bb8GIbLbpi1v9yDMAzFeHX2B7q9rt/tJLTr9Vol4MdozkDj/nmCwVaE
blze0/9FsU2tTHm78q7iCWuEw99+gvCJ/prWGPsUiwcwmxPyatK/r70xTa34HBFv47UNs1WLEDE8
Z4tySlTrTWDOEd9uUi4pJNd9qupiZuZbGtpAwXKu3XLIdbdj8nZOoe2kstnh8oxqFTDgcjzyqMKd
zhkJ/WwMehZ8K7cIlvUvYY4r1mM6/BNjaga4YGz041q5AG1o3IP5J7IqJzOjz5PAKAX+SgA2Vk/p
hxyQrXUTBi4k7/YKgXX7tnY8izaxLPwdJ8Of7EC+RS9dfspAmzHznoAGMdkyaBRd2E6GDrU2NA86
hap1j41dRDu1171tieZFBk49rgIpf29B6N8YmesIbDrDbp9TEeZnSuRT18ExgOUQLZlfzRiaQIX3
u7JEQKU7j+eZBAtAAKSbcXRi7LERbr3rGCn4VFwK7HyX8jZeiq8F5NdnmD77KDJDlssrNoSi5fk2
AcIiECKSSpXEc6+bVoyON2IruR7erIC81n4aPsIg7/P2aZLshMoTQThoF/Ps552SKDKhDNeccsrj
5VXOqFo+IkVpKPBmmFJ6lep+iK0Z58XEVg3edH3ILqEabCBMdLSCYhb3hnf0Eg5V8TkmyhJlwXUa
goaxLDcKKoJQeikNF8lyvIws+78G38AYTLk1RPjq9XahtOODXHuJ/8671ESM78MoRjKVrbiHLMDG
ja5qHrwZz8SFyQMEyE9J4L4kouYuZGgssr7MJq5ydYiIBOAQafO4NV1phdI378Gh6XkrevH5V2W4
v6L3kvIjS66oWAUi5XhrdkaAJv9U/2BYw0ibk8xuk8Naa5q9l7mvQ2z9JA9lrYVS0f3FfDHnB9b3
+gGZhK7stxdhLehLGEj4sCybftEr2ZaSGjcRzTQ1c6khQ9Iq0dRIUQZgn8zzykkGKPv9+KY6YHPz
exus5LnIwT8r6OR1FdQCk8O4ieVzc2wp+8dGQ6Vgk3DA4T7O7cz70Xto/QT/eOsZNKl3TueVMmzk
pnCuLeeAL0hpUdYJcxl7UelqKg9DUCoJpohzyDsGafKl+RZpFDjNLz8ZvZ7WpqxBo2WGSFItgVTE
/XNOppTEqmFuWXrkqCZBlvkkVpDFjsHljqnmvt4STW7Ie0BqsIQfhirZO/VAQ+wZU781MyCoo0cr
qDSVtzBpCN+AarE422Lj9d5v6HLetKSZLc5o4bsuMTcRjGLF7+DJw3pSmMa0EgyTd73WUPzRmiUW
7I6bmyL98RStXF/abt0oU36l//8XRjHSLfGSi4S3U7C9/52Zp7JLPL51kafFhk9SUmEEX4pJTMrP
UR/pic1OOWT/8czARUEAKaSJxdQ4bQm3Rl6+QH66YWidFNeuA1xuPdcxeHDgdCE+xQXTnGPY8CQb
93bRb4KgSbrlzhFeuZEHwi2sQa3PV4O279A6MQNQrettPW1/7q2IEqILHC3JDZV1BxYH5uSXJF38
T9+urpTNBaujjNprEgjuOaIfVBKz73IdMAkdsdrYU0pOqVVTQm/zNwnp277vLFf2GPJxPC96j4CT
aOsbfjwZ5IBpPZYC2ScsmOKSDdKEAjjJxWPH5flihofl250jr9Gk6bDgeLWwRVrdZC++Q7Opt0IZ
bAcBVVFczIicQBYaDFI09Ar9YHuI1rxRr7RoODhqvsXmTkUvoxFemVJ9UW7oTLE0CpmjfZ19HfZt
fOwoRmc7Zjz5ZNuQz35UdsXU2gg8pip8f7TzIxI/8t8qiRGpIxzS0xOmQ32cjbQJnL3UYxIr2uZe
PVAi7KtEOccVKZpMP7ZFw7Sg/3AdzNU8myatX0gPyN5ZpIFAxVZfw3foGvohWf5pbI6suBJoBoDw
PvZQeiA3QslDf4I0FrHLRl/zKMzzktD0vQZmbMQTNOcckuXL/CarlWA068NXNS6wW4KNfaGBTFxc
esqdl03OER9R49A1szrxuETYmJy5upBtT9X+8ZIbdQuZdza8f5nDcDp+4L8oWOfLrWy1cbGDAgyG
WJO0pbf1edouMatrqMxIg7fg/1syJwBOqvlcOFqm+sDUFqRffvoUxEPbMQ5jQSAB2B7am6/FHqiD
rjj2bbJDODHQ5iCoaRJzxN+LLjAak1D/RlQ2G6BcRJnAR7kqW/ZvgYPCv5a6UL4GYMe9DePBgD6O
pit1IsKPN0kyjvBhPxjlyKI7oAwme6BQN2AS44KujkVcVsDJ7Y10bncezw3m2vq9LAypF/9ua0L5
2Nc6a+1cPQ1aLQYvvkKcpktf+y9GSAt3clQx9PS6SAWGkDfdWXwlHJa4MLCHlTZvOOlT0TO7ckGq
ozDZUCCkurPKfbm6qePjBO/I4I6812avH9hLYFKx30zsAP+Ff19H1IpTi371uasboBP+koheMRQe
ZOgZ8EfkiLpEVIRqQ9euVj8uuHI0TsI9jCIuWRfJG/agqW52B5Hh9xkMPo9mDWUX+c9+OrVIVIex
XAwOuNSh6JOpO71Q2tqw9mOxNLO42bwy433CJScncq7XBqKVPhpbPdVnmaF+MOVtE+hTSh2iyism
gXO7BHQy0LIeTyVxA+AskwqI4/TmX2gZWyCohUQ2RYHNbmg+iM7LsivZQJAjCGxbHzykt9lRcWJB
W3dCVoH3WQzhYXjdP1lP4uXeI4UYVPhtbrGzylBo2hEV1dGYEKDzspQsXB7Dg0PnI+/pTaCkrSmV
tLPI2B0IlQwvJWy2+Pgl7AVx9BY74HvYfgrhbUUO33As853raRVjVAQYym0oOOHVTjob+kKNi63o
IbwdDhYwekOlSYdZzVfnEHzwtTd4svu/YqGmZeq191qKNVLrcSI0Ag1t80S5OqcU7adItjZbfc72
knIkqHVU994fbQnQDmJnCD/ircP2FsUqJmqIe5X/wrcgU9GKMnDuEgsaOFUuvyqEqi7rChZ5frUh
PWoP7cDblaQ4r+x83YFdCMOIpwe8mfaulJLF8CNOcKP1NqYLtzc6Wo/4pi88trEuExGhh8b2ROWR
OtlMdGxGZ5XB4rUTU3h1uuas0C4GRUWrt23pEacaaB0s4OyQI+Xycd3hVppTlSvdU6rX7Gxr5Pmm
dvgHZLKhxIiDt7GW0M3jMCwufy1VPZILFHq55eYwnqCn3KKqeED0sssWABOoQag3NmGVrHsxLUO+
WZllb79oRwEdIN1Yr7dS0l8PyaDPcbFlloKKoXf4oAu7d5XFT1ld10LBuUsngW2iouQgFRGdjjR4
+RybAktire4Sy1mJ+Z4yb0Iarn+WJwJHGny8JEabph5oQiM8Eu4EHIG2dahwKqjB2NCFsigmw4pu
SMtmfMCRYbItIG0YvfKRDxFK1krkP+NWoklPE8Cf+OZzevIXl02SGHM3gHVD4UgoJE3pJlOGiVVC
AgVFFFR9Mhcnb2tvjMB/xBKmsBQtL5B5ucj69TmMwLcQsVpisIXeOy7EoN/KYrDOU3Gzw/yYgtP3
r3Hwc5YPsr/G9wvIVM7ng170KN6mHMX+mGRwMdi6ETkGA/lra/84elOa1mkZNLQ+zsVGkMB6PZjG
xaGToxDgLgt4b2R/CuaCGLp9L8OnoeiTATvbkg8GIGY/sH8Xy54PXnrKRt9ruoqFfe8j31kaBDoZ
LJMEW3g2F9idoy22L45xMCMui6+l/A8b1HBYN6r8wj3I+ThVwlehOXQS8uzk8rp5pV2O9hri6W28
C5yDFoVE+oNj1T2M+AbRG6yzyS5eceC5DWnqxE5JsnsgyZDpX8zYSUFtgcjJ4euQmvatwf0BCJpR
Xpb3z24feUdrUjqd73ov3wUuwLQ6WF38F9C5F8kn56/84qqRFufKCvNAGE8dn9nvuQLDLKZVUFnT
1PdLaKQU/flrWpkoaQWH5PFrfUQC4PksrxSUv/XrViEq1Nq9J7G5F6/Uyf/4pNJu5C+Zye6dTFe/
PBjWUJ0TM+TVZnSebxraLfAWFdtSWeFf+8ERneqOLtF9ahq7iNwTAKuznkS1mapNbeEYhYT9m3/T
YYgCCtpsFHTqfKVy5BOipTntSt4QlleJ+W3CmCl1CKPElgInhD5CwCdLIOm0AzKwl2zPLABc0SPl
tJeFN5lXd2PhX8M1cFEXCtMZB/6Uvuu6EWpiGxG8wKEuwjuEcuf7N3FWIdCdIetPg5s21tTl1Sn6
c/FAugj6JC0rN4/TK2VF4Xk4uenNWVJUaZphimUBhihaRDdgJBZTD26iee9ALM0aGWbMITBO1vsH
TXx0MLwu+W0mVYwNOtlTKHuVq9bl7w7wt1xnwnv4j07nisj4XLf/pVv7uM2rWlfJBhZ91tQkrj5Z
5mV02hbqxLOYGBTCvZEiYy2+myGOqvBfY/bFkShE3kmfHurp/6sb0TWNUBIykRF3Z6GKFy2BhWi8
wsEMZCv/cdZbb4zxeoQdjGzTFevKSchY+IMt39SrxNytv1trz3HBWzSR191PnzYvwYmLh4kx8HX3
X7T/KqIU2rLmp6ebWZrLfbLFwJRchQWzDMyxLTEBvkZgl689sl/MMPCGeiHl85Rfy9Kl+GKyKejA
qL3L7rYg4PXmh9qQ6meplYO5Mib1MFLkUM1VIPNQZWNcz8DYWjVNYUd54wKhe1cQmFR7qjkYNcb5
eeyTKfEWNWeqXTYT0cbuKvh3QepzcUIQptNYfXTTDRpTjE9ugq2Z+kA7HaBb08yVprX/Df56Vzhe
4wc6FRl7WZ2oUBc0MRQC5lAl1c9m7RPajEwrk6CSeXN0p4Z1xx7i+LbVOyE3g+VHCpGWZrf3VjDQ
DeDfeKYvNRpl2XoPDwjDP17TDyH1BOL0OG/CX1fLQO9Bou9fOoUwGj1f7Ls55gFmabVJAtZMcdpF
yItO9CoI00sReUTuntIW/bsSsEdurqLT+0xmbyX+uMCDeFu4nkUEzmd+669brWDa59Eu+YIm09rL
dtIg/bin95tJbp3FuBwsSPUw2R0zKxt3Dz7CHEfR3LfR2VYDH6OGeoBehaQJLBDwCOD8Asq0n1Ut
mx4BmHzpiw3oEDwGg47pmn2FJWiTiH6aMy1dLdG4NmcuaGC2Wa/Mtd3rsFEKtL3IoMNxTIeUGRUp
9pACWG2EFQKxFNLsgVrkbnQch/wf38ex0NLhVCpzr+fMWG7vHX1krzNUVsXzlIQU0RtxLDRjVc6U
7WMcEb/DDL9w6XQKdmrVQp4TqMFoyLIs2YurjRvIQVqx6zQbh+CQBl5vCCubkFDJB6o9FE0nYu4x
ZJKi6ey0HZMfk3R1Ntr9/BPFSLPMSDHRb7lo0LMWu47wOuqcPQbodcKo/MIoqv2QsFbNk9l4k6J/
bc+pDAM8XFViCFd75KkS41i5m8vbwfjgX7dQDIzrO8l6r1sgkjCSRxqU//NEdpZCeQHkXb5G5bhZ
RN4thJRiCPpLkvWdJ4S9Xdsykb3jz4sfKLV4xe4Alrpd/OHyC7iArpud3XltsRJUAvsur2bmOw1g
dF9qwFxY/sFlNuu0Yn+bW3sFx2pZXK11RCGGSyTfnuHiGn9gxYo1nFGzd0gJ2a4Um6Pmfx5Fek0O
TggFaFN3D8HTa3KtU/6YcE4LwXbils86mF6gxeUm0frvwTlann1kO2Rsj8ZMCce8awF+NGWYGew0
/9JSdtQJMLcJmp8nwob6OQOqVJfbNV3Yj9wH7VmFy90X2wxwDwy1dwQqZpcAwOWoQvk+wajbTNsj
CD+BW2upQ8K1NVwx/I79ZUVpinsQ2lLecpl186y/eZVRYV1qmS3vZgGdf2Pq02zilBz31pgndbX2
OqzmtcBWD7SQhK91Vg9YouI5X7Hd5w438v5ush6JDKxCthNc8UpMP11ojise0TwgvY3gfKCSnx+M
pgxWqu559WBbZpVR++mnwJmiGx8MxnXB8RRqsLA94Wda1ZzxQNx2eDw7PXXDN7P5U/c/YC7seJP8
GfWlrLisG0kwq9TAQwXYIGAgzWYhTWxs5z0UXX2kq+I2p83SR/SKVLVRFicqAZjpNy50dfGpNodk
z+aCnXjyYu+tW9GGFskHzgI5b1YBnEYKARZKyNUdj5TCSKg5YXqvDGtVQblbCwuMG25odDt0VYPW
XMrIJZI8XUuzK34xCpJ23o+kFAkXhqT+Ic0WbeaRXtMkSlCLR/2w9C9ni40i6PU8VA2GJ1e6/fVU
LZijpERqOG7V7WDYGrpai8SEvPKzXaAHg/qBYRaZpdr+SrpIceFWFN/ZPnJq5AkWyWBJTQDdwNxV
WX3Yix9Malud1uaIy3EsDbogFaaXv4lbTFvv+VqHx4CwJzKyR9kUvqa3XmiwqKT81MHe7fSWNIQJ
SiV/D/b43BuWqWYRZlFictf9UVKU94FLuS4T1AKE3uPbjuxraSDwEyYjQ13l9w8ZwHXRJd6yjgUd
3ccM64yU8NWQorlMDojNQEmqxvGnKttLvK/ipT7ecmwexYKe6/pv6/wRZAE9dyh7WPw0WaydG1cT
yR89zsBfmDtZku5xOhMvesK4C9ppcZGWfJfTjaNIuAQW8y0sdWQhlPmX3p1AvkSUMfPOtU6Yc9U0
gObzbauwzxV4KfKOX7VmcnGAJuQic4hrAo01so7OtRDVD6WMtVvQzPBswEXLRIt+hJW7tfmzfw84
0KHSxTOh4hW1OOTBbU1Wtaz2r+f3flOlit9x0tse92Z57RfDbL21YCBB+6dqwd1Z/4aV7AeUP5SW
hEbjEGvK4WvzC3L4tsvGEUf9thDfb1RVzx9Yg8bMBHgjPVNkDewIJG4RWy4ldok8RQ+i6VVQszmv
lsQFRETXeG33WByK13xsp7nh50Lbl14C+F7Xp6dP572a94WaOzWw8rcNyi5L9nCTSAhNqVLFEHKR
Hp3jr7NXVsZgN6xZao4J6+WyOVZYqOuTKPYl6+HOn8Nc016xLwkyRvENt6PPEdJi6y/b7YEIqEN/
mpVPn0JnRbgJwwpeUv+uGELgkCARmNlktCxzkXGvNEIJcPbxggFooil82/tV/C/DUuYLlk7+G5mv
IrbcP87Jar1cbTj4+sM+Ga6mtFT+LoPcyi+5OyF0f2R5yZwe8WdbF0luEHyt8lh+TTgb9kTAKgoj
QX5PNmgCICOuUc+DDNyPUVqSCUS/EZe6nIoCXlWNKXJiUy5HbzjDNemIoAbd9ITG3VTXZ46bG6ZQ
hvtVo5zSJLQTOtpqkDitrgKjzhg7RMdcm2bemCjeEldrgjvZJLdMviK+SWBZq5LI3FrzRUy/Zhab
aZHUF5NBc1MgPDzl7pzUvanVlkNjuxfZLGitQNIihrk/dWcTUkneMKhr1DbmnOC6e221otceZvge
XkZtd0AwyajirG/NAy/Yd7yUtLrXd/QFGAeU6lUeMN3Y0sAUWouYzu7pMCOQ2JsxQ6S/G9VzzroE
AqbkYcyaJwnb+Cg9NbYVP5dFCRHzdz1A/dUuf3mdnjanl7+LNT5EmysYK0IlHFjKA1uU70EPQa2H
PHsCoYoh4pocu30BQ6dJ6joAKTsA30Kd8qbh8g2v2qv3L0sN5GtwGdhjs8mR7+50aZ2fd5QYX8mk
gsF3HhY0nsRqSAfY1eLlF/yp7bAGeS79RA9zHivqnfGJrW/0nnNfsKzObvzC37ci2m1jnsfdBjD8
06ItKdh+ZxzWM3+siVRz3MtvWMEA0nkbg8UE9E+jJoK1P8IVdC23dvSM+9Ha3IddFfidxAroxi0M
u6FaWU7K6ITc3UPUuC9v9QwMC7G8hXcOZ6W3ZHvinN+Coqk5GYlC32tpD+HYWLAPhLhv4zX9c2BQ
OnXPfmRX1Ygr/+qBiUP/gTc9w0J1h8rJr+bGjkPhwCKgCw9KQn/Zu4zgD9yWAaOU4f66rbpzZjoM
KcixEt5nA3fRwCsNHuq0nThncb0bamLUCOAIdHoTzxZ+0uIGBeTYwum9cGJfDVKX7A7zWL6iG7wB
RRbcypctHkC0N5E1DhDVQVDr6ZGwdnRmlM5BtrDoWbUIfo6d14V17oupUswQWD4q90R3wnfMUMC9
hDgx5+gAi0C6EYU8rFZcoHEekEC2aK6JaLjWsbwFdE8BnjHGwAwkjb2zdXM2Xq5XObbIGnXwFByU
YXIJe6kV+gOcbDCLzY+/4vy/gPrawkXGhQTkoxE/VNfLr3RaU+tzl3J1Ql4Gv87oR0SklgvMhR+w
r+2oEfu/GKAV+3qWUIRlz5RrWsuv6+3wenBvRtrThl3XLSPCJy5m1SSCzRwn2tThdLwBFJ3518UX
chZGGvKI9edszta7DaJ10haObGgzM5W5Lewso5ot2pyGfBjkDma9+uVgNld/Jn5a/GTkl8gLt4n4
0wOfDxbOjw54/2SH9DH22oEF3W/kGMAQeUqOmzCUiLo8Il1qdpF6DcIlJuqqQLcsam+Tb59Im/kT
UQjixwXc4h3zPHOvYUjWViwk7ErocMxVR6y7WSaSocCbwq4T8oycvIL5wlbNtfvTeBcOEv4Q2cwN
krisrX4/LP5BRYZ2le4QghbbbsDRqFSI76P5wfo6m4mfN5+HGGosLfbofZEfMF3LSLY7upY90R33
mgb+8reVysCgVApvPp6CEckZrZzRYyT5HVoeM/m2IUoGrcXVTHpyeJkA6POQY4RPaC94lLeE0M6S
RzIFxNyf9Jf2lSxfeiJYJ68zK0QcGKaUyX/hONsWwReGXx/3iyN+sEeCG8n9a39EfVMMI64s5Xq0
iGKjKtmQMtp7FC6EYhP22leZ4ZuIOAJjX8GK/Sfrq9fEKL3M8M4kN+lXPlwoaEVQ6HWg1cRJUyBh
XlVpUzjiaxKSR21mYj6lAWXPhOQC2z26kM+OgagvzXBxf62hQUgjs066c4Tkjbpjgbg8DZCmFdXi
EhgMeViGdphX8if6aVGXyIWXQ3BdX5vtLe3g6B/CPJRVaSTjJoM+ZUjDOK8fz94QJWoN9ZgE2C1q
z9Nov0EpQIQAsnTbsEPtNmB8c9ZlTizDrONRIboHKf0hGP86X5Sm3xMWdwf+8UYafg0lPNTetnSR
jlrgPtjYRGF35jUAdxjp6JkYmcyTfexxv2zrdRP+4KZ2Fz7BjA/5EOB+bxjY2y3hSqQzfkNK8pw3
ameEHGszjvz2aVeJXWUa27AH5qwPDOK2sPXWCkpQYw02qJOArL2VOR9XJmGJCsXGGR4C9X3ueZsR
cN7F5/q4Q0jY6xWvq0YZ1v1ndyO3v78vnS5LIDcPX3uQyJtLf05dc5h1f7cQj7IBy+rbbqnG5sYa
5HiyB8H7KQkJUSvlKa9Q9Zsko/V2NTZVIn6qji0Gk3Y6fAgdxqyJ5TUD+36Y7ysI3bl3uRbFZOa/
bcEIneI5Qt33BJu/l6LW0l57sVbP6Uw9N/QjBrWvyh5MV77F2rqWFs1pj+BY/QUrO6DQUzTBQLT8
gbet2d9tL96af5Mdpbt3o4vqFTc0tatTT20gWjwGqjiD9wuI9WvL+rpX1WAdtc3q6lsT2+HrOR5e
DgknmCXh8hNAvJrRJGGi/vpX79msjmxQopiEomy6eEYL56Y2lWKQ+/x4Jp8mLt6ovD97hiTMP5GW
SM3z2TL2gQa2E/plQ5SRLGePYerYYaJzk6LXi7DMiydL5uaqoOZkVBQNrIFM1f1EWttBCkKqPbcX
ajTdrWNL2IXIsimoRBe5sztxbNPQ0RYX05LIsl/Sv4R0zvRfH2xqJ2CeNd8hjl3JlXABALBsLnpG
S80wrsRVnvf207S4CFVivW6G3qYovNhctgkFsdIITFvQsRqdCh9SCyzCeUtnj7Dwr/hwhKKK5fdv
nti4g99cOip1TkvDkr6N8gElErlEdgYUBPFU03MI8jzVsMcGMVQOGR2qdg4/xvKwHNWQfQEUFHCd
U86FBi2gUeOmxoLa/jnXUBYO/JjB28XpWSSk5EnjMsXC58rAjZqjhdExTMK+xyI1Ktp88RvB0r4m
iZTQgAOlwK/GJvBd2asI4q0T1Em7zRzR6czyBw+Xfsjd4nc343ylFvDYTOhf1kV7LHW8At7hNGrD
SdUIvrQfT1RMFVVr3HHeSVc6Ng9RSidfcVSv6tx2/q9usr3GEfAg3hnVZ/1InuaTRc1/yZyJHOWm
wV4eXgs0QsiyvEOxr0xKM/5OMfaZ9vIzfwL8/ttYQhNbdQi/T7eb8Ve+ZPUqhkqPSEXmwvasZsRY
nQ3rg6EDslporEO0VHNw4uCdDSWvdH4fxeMGUS2XRmxmhRm/2E/n6WV8B8OK1/zRQvlk/A5YuMDD
Gf89nl5NIvczmuU8pLUJiuT1mPlM836ij/l3e1qi28DDU311OueKS/7YVeax7TNfXJRLL9+HOD6H
vyedyT9vozpfUev1MyQ1jkjJmPmeLgi8ahPTi8/rDcFfLn6czypPaYfmPey1GMe9JOSpk4uuck40
XtWp4Pas8/dGYQyezD1kgY0zMygPd683T/Rzw2mtVoyux8p7oFp1S5/D+nGHBDp5GZ52nQl8W72C
yjds/chkRGNN++xa8gNZ3RKpkLSf45pKWyhuc0+T6h9E0RrVx6uH3mnGJzhs7Ir+n/p/sjkeZWFQ
hz86oxsDPyb1QaNBWl5kHDYgowr3SGyqWtVF767BaKVjIcJ+OIpc59v5x4a2rJK9VhNJVtl2hL9M
fZ9w9rOWlRldhXJ34w6FhsEYVPuVaCdqH7XIaz+bMslEhzwnVUmdXBvAB18rm4dpCnuA0jNvk1Ay
4R7peXwgr6iqXdu1hf3sEdv9kc8BwxpH2lOu792DKU2EfPy5t5sBo8TdQ67hzcHAwC4JxGPhF4hs
bhgGG4b/z/5V792f3h0ox/2rOmLyY63VO8KXncfAZhq1iAZickOnSP/pj6iUdO+9GATttiqEvFVC
52Zw4vo7OJSJx1bYvbllupCAqNIbW57OySi6looD3fSEDbE64iQiprghLGSPIDOm1zEa3F5qjAbu
+AZBbtewPiAqIkkTU6x3iQxC5HS0qqRsO3cHJDaZiuadTHkmDoVYSZBenIit2beQo2A7xDMb6kUO
xA8s9RlFooddHi4ykAJXCRXB14wSjC+NaPxwhpGeds0IRBXIjvHcZ1X3+gqslBmy2oBUz3wHVU8r
sNIgsdItLFCHNRFMHLFpf8XFNbgIxvX6IYcmjJPvRI29GAfn1HSQdcdM0JjJO3ZEqhJCHzqQWSaW
/6eQBRxd144lbXBKE/VZQIbve6mlGf8l7EoQ52QSb49ueGUPw2kQvMiliwv/U1C4Nfwgkrkr6T3r
7Y5aOIPsary/+Te7kPZSx0OattaT/+xGTGJide53L/ElY21whIazHetGHQjBPcfCkbkMwAfiKZ3G
waTcpo7HSR/DB9efjvKHuTH7EBJL0jgjl+MWU8aiTPu1blOa3tN+3sjDdYfnYgqH2xn2wYQv7QCX
uwTFgZ6hkg+s53uVYAt6mOOLE+ivPtJoyESDR9swyNBFIZg38qAnJ+QolXPsm2DPly+DWHqAW4Tu
7p5okbaYxeHJFhwelj77CmC4h4lSlwULbNfINH0+yvJTTBacvxdv1MuZMU2vbgctoQKuV62jNZPj
4ojiRMCZF5eQgQETf/Ftd4n9FAQPzak93EoJF8U6YA1sJo35UweUophBVhjCmoJzThcKe4ypVCHn
4wP73WGBKzVLPmkughaxv6Sl5h4kNxmHGoqCurQjVufLHUmesHPNeI9+5GZUnerNRbNPzJR6jBRR
GAFOPvLo9aSj5gQehbBhhHad7+ol9/SRSD+4r/nwHkWd1y47i0rpgcyR9GW5yz8lubyO1NTCgVfh
nNmgWXpESELVHhitJ96ZCIhG6z4ee9WRszPT9X8P49USY+CSF9uIO0xJCY5PEmV2saRhFr4NJ/i0
e32n6RVqJQfSNT5Hlsi3H6AhFgVzTsQ6VQQcUfRFFwUZ7UcXlMMtsTq0/WpEAZ3k/XKbrXlckYje
LebylJNikLZXrooiEi4k4NBAGIo3j3DT4J4LFlSP0cwwVPGD3+UdguJEsbl1Z7xYLym2CJroB9sT
W/hiaaenIj3JOouiI0qEEux3mWG0khE5FcIFNKHlXikDcBoXZRquyFtrDBlkqyc8NO+JlIVcO4Dd
vGd3xqkv8FqOREdPskeOAO4NcQvwEY/Zr8wJfNow2UFH5Sd3qfFP3o+WGKKuV4rrSWKnPPXPkiXk
YFrIKNycrsjljOv4JWsrKFu+SnkSnCiDrNOpwPtPUKc59erNupxKgV4a8HUhkSZOECS2B42V9BJM
EMpjz1NBzYMbN23+VGvOnspUtPgAZ8q8T3QtNuz5kfqHtAacXnmLCeD2gkU+qbkX/MctLKDk6ynE
0J5xwQM8BgUecizBo4TCO1MJRXNx6QmGvK3CtOhWVtQ1jydAbJJWGDAUKo0U0WQ8EsDkPF/AwLye
mHNBOcHfEv1C/e0J0R3PIJpL0/l4BE+bhg9yAGUYzIclAylDDhIIimUvvovjmtQO/1iKPCOFuRKh
27AYkgQPzg4B5BaHNFHRmtWB3SCMw+wTubrLTc8Kji/83fZVpD2zjVvmTvVOrYa/PZfaM+WV6oYK
kFSFIV1JW+KM/wg/2unAchSgWgRK/uqQWEWou/dsVqgSR5Os/ULl4TNId6xLZZCOUEpNHVdeborg
qyUTbC0Vq9t6CITnndg37FgDKDYdVRVZVFnitwx10cIhLG8/53LjxFhxz+9QDc2JeM7VTctLnSJz
fwGcripiT/Jwtgp/GIIWxW91/lYkdJ2kcMWCfMkbZkmkcSRkS1CAKNYNfQWnPaVUR8wLZThpl6uT
fD4VYx9zDzbTH7nINmA87YNYLf0pmRipPB6XBTjQgqqJpssigNCzadUgJTo709FKdGCZAlkGbhlD
5My48JJ1KtisvIMba+QdG8WptStni0Oczxcg53dt2P8ifXTfat/LouvCZ+uXPLcTyCPHZIkGNh6c
HR2GrienQP6M+/b2IOmEJIrICtQqCg6BxDchhaC7VjlRnlfN+z92XziNFvtREJJagIO17+pviqDE
bIqAaReTWwH3xzg4fcaduyO4Qfq9JUeKUgbGEM72eZg6PshdTRHEdXNR9MOKmXa1FKemQ0xY7rcP
RyjiTrc7g7foch1RzKfBY3EkuGj/cfUS9+JokqA3UPrRqK9MSYnk/2/nZI08ELIKNVdeQasLWlWt
fy8hzxCJysCjJdpUJMzabKm0awzZXF6c+7kcBlj/JSF0wLBd8MFERCyzj4PCl+tEw9aJWRX3jgLs
paN2+0ZWvfyQJXYVUxpaLlZ4SUk7TmayG3JS9QD4yJtiOky7n6kkVJxyWHEaegnTIBpycqn1UImb
kZzFC+B0riosrDExRIHZyhmSzzD9XyT1LXjvGhw7hbEgMK7W5JpUfFmSC052cPOgv4rVQm9B0vgS
QnPM+Bum/f5zJyDNjfEyBLIWnU7ABgUoi9xggUPXJDTYFYbEeKYqdeQdL5a2ZivnhOajhiX7DZvi
NazquSeC9I8gmHE7cdk2OipSg/Ok12vDSHCcPZ8NNNgIAZ/5fyG4vMGlCKv1smtYC6LNhbm5wYn0
T+/EQhKp8/yTSUEvnUEfyLJI9UeqMCAivxdOUxyVg1nu/6mRncAFB+XizHqzb8neNKYJtEL0d6LW
tBrVTXDzPtkkylYelLe1xYGKGJ9CG2pKNI9fLXhnAzzvW1XgThREhiUxO8i7LNTEqcDIstD0BWS4
1pIAxkXHm4o4VFSvJQlffbe9QoFNvZXe0cCYEEYNojFqkWWKZ8WR37/mQbdxs1/hHFPUsZuYiRoj
jdqUC2RTEpvM7VCaZx9r0KMUk+OTizGZfY9XSz8sDe+JiVq1Yzhx2uXkLbOQOrSIukGWZ5jDA1M7
y2lJVIRSiQLz5XIE7bUY6wvzmsLl8bx9DANKXM8QA24S7uaTOuTt1xIbxmAxurr+NEmYfv6sH/Pq
fWIxBr0dAG/LymhdzjbT145q+/USYKWyuoQ4IsyDoYChAL3hjF7Af6cFUxgVJ8JNm6hEtCEeVL+o
jI/31McnH3vubNQfjXF19WZ0/Ioi5Ndi2YHvfrau3cYYf7srfvqJnrBZkPEFvFWv29UuDW53Qcxa
G2SaGK/UHSY7tMAHknOQ0PUPLj7a64X4ScmnkoA3CDVbD2Ny7tgHPRzJxqgVgxv6JLdTM+PZTvYZ
T+A+aYRXz4yrLubf3/ZLvKn1FOq9ipIFjlYFw0qkwzofS/cGJhtG33ZFK2YPn4/fa3N+tnOwtJh6
pRvP6aucuuzgZPin0tGyjIjs9tatrcp4Os9f+C/tL7NiBfpGW1PgFAbjCvbbyG/bax1VbYldR4s3
Gc6sokfpNGzrhA5EyzhdhXn0n6PeAbD9DUcAiHc/+39X5nveGeGLpDSg5lUgg/Zoil82wRTlXKok
Yjq/5aErlNk73LG1RtStMTj7brKWjrTcMk6Zc7YibzoYuvLbCj9TTT283dl8uSpxcZJiVy9s23n6
D0NyBH1+Z78kfizDSIYPQlt6A9j18NQ3lA1hIIefkwuBYalIcwKvMzeP63/2/mqitvnybDtO5v9u
olescM7ZIP7PcLhDWUQlSxIcEColcHmJbR313uLtJPpqeUlmXEX1UCN5fIcXy13Zg1dT5coh9O13
X9tvcJbiSdj4SBj78/yxRa31lpzclu0xv7OV1AYpekJVIcOl/ND4FBN8ZxUxxvh7GBB3S8Oy2xFb
Q3UAO5PeKMBT5om3eDpKowtb5xSrs8n6dSp13k+pKxPVQ26eY4RzemoXtiYLke9Lmn8k9r/cGt+P
ozXYjjS2C0n6r7DDoci7FkiXV9dLMvev9tke75scUDU9g8p2x2Gkg9dJgMOAdF0xaz6MJQvM9NPm
kuazvBN5fmNJtg267Jfn0uqWHgtzT4dXLP9knnoDg7hX7BuPMzK950wzgPc9p4CvjtsM2FrtakFJ
UyaxrxbEuOSkMiefIwdZBmbSK2t0sUlKRus3I6J8n7VrtT6P/IbvvW2VePy0/YxbMvIVf4n/Wfb+
AtC7P9U2zkgkAPTHBt96Vqz0BqnlcdLU/15cCxp9+J6gSXn/cIuT7XebMVc99dEM7KR/Q+kivSWc
oU65WPn0XZYm7N2luTLayRduUJsoKGx4Jc8IYCzS/84hJ+asio7C99zNNknysLEnzSp25/tFEN/W
NHFjYrjgem+VX3aoe/7rW7QHFC+u6zIJnV2GxIQQQgWOpt00sUksnJ2i6Koz32P2llgJJwQ7LJEz
+3luRi4Ilu6G8VqY/0c85LRaVZKoh6i63bA6q+70lkUYgB84uBWiOsAVJTe7Mx64ueyqwG0/+i0U
3jek988aHwfZaqcBkXroaBAn6IHRRwrJUDFsmAJ3yWr1Rv629Ppb8A5rA/DA64hURGECELSLy1f1
/3c625veOnXT2VxzgOHjKz5uc689LX3sYjdlaVslDk4IoTkpIJAbWHM0boJmvCAY7GtwSy3HuTiH
aO4NOE4MIq6rCQEcfX1GfrDf2fuz3XbZsveKUJ2ViKxkRpRXpLugPLFAbzk5kuY/uda2nsMI6B/3
dakcnA1+d/FO3OIjj16vTnRRsbarsePhQiMYDPUvC744eRwsK3XtRDjzSKv7W+HrVTyCKHEAdlGU
qD2/O6cTjACiLheErYh51SWbVpwm8uZdSWXiaIsvmr5Vnp0HBNf+vlyoJLvx8sDezuR27f/lxV/R
pSfCURmRhzM3u0LBy8fA1uTVqnp1xEdSEccHfQwVfedsje9Wzwu9FqiKF7jY389rWF3FGVO1povg
dIMemfuAqJFNn1GkgOFlLnGlgco8ujYvI0oI4RUBsPxI61fz0BHloIxU3A5c0tgbl5uqAA3BTqie
YCoHSKAPLO0NzuE5lCUdmG/r5ppmWafWsDltgWZknu7KwNHhEg+6LffeLZoJ9jjbFmKBuH+pR1hW
AsmSr6Vi4c3xrp11h7o2paobpVUOHgBgOwtgaWQ6YFDsgzJUmm1IyJygShJborhFaMnByPDu7xcH
OpWrg/qcX5AnQ+v5018MUq0hJ0gqcS+GepRL2DgQ+GItvlBkLya8cEuwjhVFUa0qmJksxwPj/2xa
5fkkmzaMFDpNAeorRIGP4bXaDJkmtBfNrfFdi3sbiVbqXrqVvif9OE1/gdbTG1QraowUn96ePooD
lFE606cS5hvSWoJ9MOvl1DUC/mHbiVNytnltipmJJuhwrQIoUPDrzEGv/+IazYotwuqKel5TgnGM
QYxVQ3TK2K/S9Z9le1lm4j1PxpIrkLG8jWv+qRl7ibJBuTHTWiPGe9RHiW2l36lL3Qw+M0otxK5+
Tg08i9ppRJdkLjd+jrNpkVr814pD3GYEPzWyUS8QI+cSmBfS7UOSpe5ZzRTCr1fBfrX4KfvEtMsu
ktF76qhAl9kIPj8J1E3+XvQgVrEtLMijL5fdSrhKRS+4bfld9jW535G9A0WoQG/3vU4bXz0q1av7
4jhqy5ub9Qil+2n7zID37qtkTCZbPe3x5lwzVkXFXbbTc25VQcdellhBGZWhpoPqpI/g3SbKeYpN
47Yr2LR/S8MCHUekwEME6Kfn8Vejzg57v1UQn7pKPAC8wgV4oGWPtdC9x8qwNEO3j8cLjtwYISJH
VDHbJs5+ou8dFdG47FLasfFFHU6hoX3hAMVbWEIaSI8ewnGPK5BBqopupW/i6VhY1Nkcq2GWdm+e
Lw/saT4VQpU6ER7iZhvaMJRr3cb5nffjza33Jpzulyg9JtfcsZVhCs1p4qKuw9gQkpysSRO03UzM
BJEJMBIjcl8XWxGDNA9b5hde9j8PwrsbX06IOCH/5lQif1cnxq5lDPFe5a8IjnP1QTMGrYiVgwe1
b9RqqOWw79MMYbuwPZnUNhiCj6MQW6eB8IbhaekH/UAppkcWt/UZnGOKOLMmlQkzCiYmVQIqZeUi
PNZyCkXjBEwZ4SEZB2g5KN5AEl/k6QsyKHam1xYfPFZlPNnIxF6KqH2m1oIDJGzqVGWL0YNxCF07
yqK7AF8r0iyTnv7Z50ngrNEUfjfwdITNNky0GFkHk40uVRd6U8E7SMEnUd2IHNtynYdJNUvwWhmv
vHROYbgOvMjT9yflJ8dpBrVt+U6mP1S/OBctdMi44DQ9X52+QEFkre2pvdpuKzfZi85MPfXP7P2g
o4jtQ9vl/8vHchawrCXIgSAU50pqKVlEl5AqB6upyZQm8tnS+NkJ1i704azkntVw3ABHPvImqxrt
bSWOWYgtpIoAfjKgZjoX/vixYo4sgt7ZOB7a44jFkQcwWrI/e7s0eV5KOL33Ak97cb6BrmVCT+Ap
2QCWkAwSrkHdwAm3aXZvw8o49+hdo/JhT3zvNzvxnhMQf7K62w69aPlLwaBdwNxMNRofLL9Mj+4A
kx2XIFSFksfWwsgyZcHmIvemmoaukkqNGvlmNYZt/VFIH41Vd7BquhLMCXRM8lM2Lg2PMzxn0IDY
OuaLDrEfk+Rv8pcmIsdPJY3ZZwtkc0slogIlEl9FRFaARMZz0mpahypcDWBPctLDObtYORxzEBM8
V9LN1nnhnvsjUEHPO7MYVtIZdxG7OlYxDZLI4aj4ZnCVysQjn8e6TMgjQehq/IodWVx4j2tk451W
7jDF3E7ROIw0xSj1rh0dus2umDWo2Ne/30CSAqg1j0bIfDX/8fbcL0khYnnZXAibyTAg6JYPwHro
8BcsXIzDL12n8BM4ag8eftJaDyZnQNjBFEwWE0mWen0xBO5iy68lTm8zv+dyOwG7rHsN7EbXYa7V
gXloLsshM1gtXtFPoMmcc+EoEp22yJ23hm40z1Clt/WP7dIjDQJ7KosIjru/TlI41UBXpAeh+QCT
++vwmJCVHgOPLQWyJpOmnpHfsSAdXyujol0/hz3my18ETJFLPZfQ0Fbhlps7xLyGTmeBBelhRkZw
fWjZoObbo5j6INPmn9cBkj41ziQDEMHpZ1glJI0i5xJF15a1aUcJDQtp/Wn7x2nJ0d8xv5kUug1B
G6cjQztcweaGgNoos8tlQ4CybOVs4rMCBZr5aGofp1pdeiKZmIZ5FqtgdgUYCXuYIM1uKuQoAMqB
g9wndBbIGceliVSQ7k7+ujzW3/x5JdDUjd8dxHj7M8Mg+Us1ayS29F6tUOYe/GgytX0OvUvBWS2X
oGaiEMBatASXet/ugr25kAsdto+MZwGK/mXjhHrSE4RBvc3U3hwyIPQGRVy0rfbh/Jwz86G9MmlS
ncHw6elxGGeqvqHx6VskrVS+IDP4wFTPxP9mIoqnyYtLlcctAmpfZFB5zmFZD2TkA+GufJ1aEyKQ
kT5TWH1tBNASeyDqZMJk6EPbYbb5VhX2PniyFAiS8lMKZxNhWDTl+BfONMdukjhBkitDR9vuSTOF
DQjKbQKXuW5u6GCzMMaev1jr8ToHIpqy0J0PzXnUp6VsNArdlmhVg6QfCKBVRNF3bkf7wIHqtQGV
Cj01wEA5XgNE4ddNdpzem4ZP04XhUHm5pT31PPWjwa+ynrTHtdjlyZbytCstNKTK+V8cTOfzbCvU
Oem2HGv6qMCK8BMEYrUddIY7N3KMs705I1LBhmQMSnMprSFClp+W7tVyc84KXyo/us+cjGPrXBDG
lIqJ6TmbCnp7Bof2FFtNjiSQlGCe/VbuFDo6Tcv2YwpIBUYWJ0rkObjlLy72k85kJZzAjlhMhB3L
mlhdchZHmjKYEpq0fUHoYe8KFVeFDKQYOQ0AOt3v8d+Qj8yYp2Q3F7Ew30A/pl6G32IIGiG/VxvA
x1ImOYVYRt2+49I9Kt87ppJk9YlNw1f4+cxO6G3br/v/egKKB2cgJUu5c78UNeIpxOmu1OZrfcbj
xrDz6bYn+vJA+mOCZsG1T0WpavU560VcuFXwPrLT+EMPvaw3daSXT+KLWfWAUd7X5hfRs4R680tS
PAFe6GqEN+YI/70+JgC0jIeQQyo/my9tFlRoFPaIJXk/TRPzORddC0uOBTKa8gdXhIWeu6QYJrju
FP5RLWGczwd5uyxqjLwmARKi4HK8E33iY526924dCS1ORcFIv6DJLDVzH8dNy28Lq5h2DSPzHYSu
aO4NGsbhUGhm7xsk1usjX3tRkIwHvHtpI1TUVJusqXJz1z3WMPPbDiCELdRRvb5WKrU38/7mxZLE
6e7OEQf5jyLUmR1spkvFGM+WQmyf7dBFtOUhIemv0CsuqYYD8iQNthlvvjw1UmB5Ui/lefiiEH6u
q3qgpyoNTrK/Wwl0mcj89zYyQNZkQfxeN8gQvQaTlfewpsXPdflLL7dzzojf2dW5Fj/Xp+U9hxOn
GK+hlqtKiEzWfJ5+O0K4dghiKJkT146tDJGZkNThP8jjwU2Dag6YrqLZhTRR0sLwF32ct+Rx2JnR
Z2FqpQxWWaKUy67mFJLmd7rcFzKDk5nnQhYIMKn49CrJApuQwvwO8H0c2YFUk35w8yix0ieEWQmC
NmJ0uwcMoz4slb9O0qKJBGRLH0g+zpEFSyavO5CiCfm8MCsv5G0g3kOFcc0w7/spctOwLShsNqyU
jKIQJLShCUpBiK8QMry/GyrWqhNmszGfa4g3HPXqFsyfEJFvdlqIXT2Srm7dYDeAjshjH8pNPWyL
16p4V4b/qRj70Ar9RUqErqUGgQ7rvNd3mwPDtvi9fiZ/W+ONemIrtDVUMjwy9QSM+eASiDYD75wH
17u7luXovLhadrr887xMoCs4xoJ5ZlapJ9n6//Wffogc+IE/qasiTklD+6OHq76nT0OfgiX+FeUl
9PKWX+o+tzw/WtED/eukjypH1MSHxgqYGwwAlH8DerVwtn47idV/oQC+lb44drTaUfB3iS34e5hn
Mjk6lMUhHOv3uutnEIAGNNQA3hSZfnGSwT3l55/YnWsXAwFp7sOXfRiu/8S3wWzDWM89VrGrpaQ8
ScMpw4NTN9Loo9pF4mZZT13lRNpASWC/e31q+BuGVsVkorxfa3xA1NHWGTHri65uENJ+kt9ndA9O
jF9Y9sv/2+y/x0bHHNY1JSmYsRFoAXKao7k1K13k4NJ9cwRVB0djuDgapJHRi4jTRDucBSPie4bW
RPk69qkCr6o6w82szspNjP2R7SwarfQEHTfxL2shlQPYj3PS1B2PeuY0Bgi0O1zL/wBOoXnfhpQK
ZIubnWPS1x8tN2YheATnZjCydkX3/hhko+k8sB1hsuNNuuDAQjLZHPZmv+Mf1ALcZvAvy3cEEnjw
yKthmUHKCdea28J/AToJvxGHrBi/BP7hzEZ/NOhykMQ5x0gRg87wRIT55EarqYGVNbyhXedNJLYh
JvmypNjEh3uty7s12kLK68P7yq9l3Gai5xS+vLTu9nc4z5/54ndVPaB4bwPkqH+l8JzcRNRa7nZv
31MpAcebiy0bg/JqvEJDazOS0/wAcJ6Qy+46uofKIW1cuLtzP8Mbz0TJYWxeEO1IIVDzHJ+qUC0C
BF3KG6wwf4chDoG8ckNY+SmSe39evwM5hRnv36I7ujJ8hHPcqz3/4nBI44D1VBd9JJNhTxGOc0jl
1K6H4rwIyAf/bk2D/eJ+OCrj74EU/TrZzp99zq4egSb+MFHWJfiWz5H0m8B22sR/EC7Vs2kN+qSk
3+cuT+yJoifDKupaW5APnwFOGupCZyA1YwJTmVgZF1l+xMgJqXfLwuKRHejr17aa+GLd/7ZtYgku
6wtOZwaqdo34MINqcW5KcwPFFHDwvpWxPscb13hhXvSHV2vUhfElL2HXuB+mCzTKtqzPvkw0Mso3
kAHf3XfFeeoLqurJZZ6/vIChVR7WdKL0/QHNf86j58Qi1Ur1T+6phCKze63MGg5K7fQVUPyw/JYq
Up8yPoLuQFAu/EhZsYA6GRZ+v3VtIegLCrTaxN0YRmtauItMKjqRhhdZ/GEJWicETPrE3+Om2xby
LQ8K18uZ3IkAlwo5o605nw2ysDuqx5z/Mbe1H5QTYTF+HZj7tDoKgXZNU0G/6K5uPu63oUekKcj6
nxhglFASwZqXlv9QC9mMhXTym+RZEq9IKyERnVDx+p5CCd1Q/64Xq37dEPlgWi7+UVfUs1kWigBC
lRsVzbWo1WLdJsk/IGzDtuzyd9dZ+PrN/g+99hp8eueTou3s/OaKuQL7ru8HONPMkBksR8RzgFXC
7mcv0n2LGNQXl34CzsFlbMS250+j4rmvzAsZjsvA97Rk3xKcQjPt9XP89LKzPV9U2etEFgEOMsjx
eZ560IWNT4Sf3YXwzP5ur57zBOzMac4EeBAXqyP2daf40pjDHsMgfUrnvSjsbdflAH6/H+zqKhlu
MHETBEW8ylCLil3SWo3luSuM3CL1R2FmPRavm45H8sJd7xkIOVN8r/D1IE+kwvday0EkdWHd20mp
gal+Hn/AI5fHXJN9iRwM7K02qXeDyv9ayk60dzwPfYpnWhq8NDwZAKfR4k36X0sNKj35u9nO7plx
8LamdYMuEB4AZxsTDMT1SJOM4s4LdS/aA7iccHu5L1VI9cbI7OfSQK3reZAv3Z3px4MvUzc9X2Xq
lLVZqA381XBYtjliYldcy3cv0dFjgZNs6ceQou53niyLClIWiwj50gyI4TF055svX+RQFt7jFOwR
aY99IYT3Jma/K1MQRwFB9OeDeTiCja7BKDxglgzUpL/Untux5v177NI+3lI5J98JIJFc04ppBJvE
TootgQ4LsyAP45et6UlgTEfAdSvucmSiPYGlCZT/0fe7dP6vPX97bjtYtS7aWfbORSEnMyZyXlCO
7vfSII3hes/BV1V+FwBmvzcekSMFcPGXRYmEKTcGb4biHeJMVZ8C/4dg+dtHPxIbTT1txMpAVboc
aD8Ub0ci7EZJncXCntR4bYeKZvul3T5pHvBEn6SWd4iDso+9xCSDRt/0uob4tHeEry/6s+ZldGDL
HHVUUEamGoGERrS2032ByBQSQ76sqGTmXna9EOw97eWoOOmbiwYR9Nj19WzH0Inx8zjlyHH7vCKn
WmaisilDJjn0dWURXC41cptUd6/TpSlSP2vM5aVvvWNFRICXE3pZrV0oeC102GQrWS0m79vkjr33
orhHI3BtcgbG3ndkuBKL1tH6XEsdVybHi8Ti0HZGpK3gw7wGozMO3ycQL4EqlqcAxaS1c9dWLlcm
PkzzP1nQ/basNhG16OMFrxhz7+a1t4+p0ufCRYPCIYZ3lP4xziPFsAiGLJOcuCcLVK1uDdSwYZX8
q/hCnoOiXdu8lIz/VKOiTIk2m9E4wbGgrPsVU0czYiIOP3bR7T/S2+q+48ymesCWbyLPHz62iCqn
kwTks0HUagZp4I6aT0UfKx1UcSzoLrNMzhYYhkbQThavqTZEGaev/VWUoC7D/UzYGJ/0GFvX7hk7
ajAztXgpZmbYDx6O0w/4Tezmw29Kd7ThDeANRnljrRxZ7HeJEu3OPNbq60eNcZG6Zqq5o4cQlW+l
baOJz0opR3KMv3qMoX8syO8TKiQdq6ZeErsD6jqUAk4uQYN89w42xGagaSnLYn4UsmNPsoCA/r9e
UdxG0hTLrjggi+4eIZ0HpQi7dlTXN3+GzTmq87N3Fi7yvHkrB547o97pvcy77Z3TH6hgCZw0GUdJ
hGsFJLZMxCQHtiBe2H+xDx/VVsp3Kbhurc6Drsapaokz3QsQ8n1j4SW8vL7QJTepy+2U2fibgKFd
f46U0+cxaw+zE0n7GlsIT3rd2+BZa7EkEg/H2eDDdzx/K6lm9UiWmkJwp4Mz1MA6tGoQA0H0k/dm
VfmOHD19EUyQc4nkoyXbivtJkrBum+rC7NRPOFm58UwkmP78aGQnxGmqSw6NQnVkRI2v4LXnqy/p
MhWmZn6E4ImTLTBNarUYgwAP8VGRPzHkjznRPFL17EtZpSOw4LGpRprosUcyMCi18htPBYfvaRBe
NiBDSzIsDeB/1NCl3dGPQlEXw0SCv6ROhbmOi7oX6tAlQgyjL6OzpTPhKfHfr+SCDHRfYSAs4V5X
8c7tcNoHgVbMpyGr/+ULrBWMOpVwPbZiXaN+f7UNxYDklaYnvOlYLYOMaR59gLsQ3Np37+BhaZTK
L6PHDDf+uUhF1iRnj7hoqtSESgu8mYZO4MvTjGNnj0GhX5j8Fy2CsPhPnbpETeemmZIyhFXcadCs
jIHro377OuhXRk/z0MPposifvYIn4DBzptfEtofnmImA+I3slcisOMjQAosxZknd5u2gYlnukORE
YKJa7c+keFPLnPLKgdIUVQYQKKzquhfV+g34eF2kNSRELvz3eTPIEjN++U6hhX3yXF9vbXAq0+FD
LewYAgbbzsqAmPvtnanXMlUEwfyCcBi59br+qypAAUsRSdDKBw0ME2KtXwDfLtSen+CYx8TMssMk
R4KFxyjUWcholgtfpYw39KM39bz1paiw6ZA1fMGzjqUadwh2RcEMtbRatACqb/XK5ZmX26jhBmlk
txOc6/yul9cVzr2uJxayA/LxLaMpoWm+x6tKHBVYRsmXudC1K717iMa6pN5dnM/H/ONKIipFBd80
R5zLYaK/AynoEEhq4qBMZwe8vsn+Lxvj3GzR72fL9s2QvgXAvn4mueoL+5npnyqDeZrgdQw4sXvv
dYWkeRqzN4ifauhmZDICj9/Yi3fKFl5fS82BSUFowwpgZu0o6yzmWXVx9155UNUqqP9uhxx2L7lm
WOv/Ir7TU4EwEfH705FjFrsTlZUz7avvIcQgtjhBas8/bDm3KioIM3Is9oUtuwuslS9DtMDHDnHC
FxB81DBGugFwdeOtMkK5IUCWrIK+ZtgTjjg7JSmvs559x46liTuqBx8nu97VQqGgN1AQmRF2FxLD
s8RvSOlLpSrVfMZP8o2EshjPXFOYVRrBsJogeZXVT2eqeajUtA7gX4ayg/dqEIbXa8hLLKVZytLj
APnn1jHOfidfnB6/YzgoqH25bm0yhurqtetMY93oWDMPP8EwvRMitl9h35EB9M7zf3GVlSk0Xhzv
pazryOeJ0gLlxOY/dQ4fkBPpjTpe+0ZohkT08q8fQQk7Pbq4GyItORf6c74Lrr1tUgYVyqV7oAlY
qyvG/C+GZ78axaqy9gGRqloR9WGWclpAKKzJDIQ+35hYJjnoG49Vk5hykhO725OrFk5HRXAZvVq+
XPXF5JTP1gSMeedxOvRDngU5YKc5JtTzvFeJwD2BkyGX0cd2Z7qbIibCdTohhZC98VhirY7DyV/O
2BX3SOHuWLX6ZSw2psFb3NIC3UH9Fa+HDS+wMo+V2bkxfRY20vRsonl4Lw4fHEfHpamFE6JgoZwn
yviUoHtxR+7uyz0sbHD1D6xHndr6ylF3vrLLUj1Rwnxvasmd6zrcJMvDxV+dgAp6NsTwKQg3khN4
6yB9YdKyzrmWdEY+3LAwMetnxJdgozWkcOmftS89b5CerHF3CdexbQ83bROnH8VQiTqvdSUvyCeJ
HfLtMpv/n2caDknqBat2KIqIZIYsB1jP3o+L/aN6gA4eATcV7WW6EuRoA7cmVNGFaZtX2h68UDpb
hCsQpZd8klwj+MckflCRSS+QJWtYeIy+tHTtNjJ56bfAFz6CbdF6H9SPvxRO7QbKwu0VqRLlQU4X
16tZJh4veBRxtDibXpalHbP4a1j3O1CD9n2zvoqThsmKYcS7+/VujLtK7qmkbf/grbj9iEDuZySt
jNr028ndh6K8jFdXnVmOCZmoOE556SAjLenkFuHc7gq8IJFRPEWXJQ6b1ZgGE1YDc1VZ+BVVjlHo
TE/EKer/kCS1bQfSN0iZ3cDRyKYDFq1T3Eph4t43uip1PFUn6lE9kDCIjv0wQStyNNGGsCTcuOYI
/lMoOSiU2YdWUJIHClpSwR20JdmZ9N8qqpz6K+ME8VNODzaHTWkS24whFuGYJYmuUzSfApKPxHDH
7V/bmlbWcnUXgYD51wZSVeDtqyDU/EjccYIZ1qA1OdgsGvndhQONmU11+7RstATS/7iXOxv4qye/
Fr64OxlvE/9ZQKAe1XJ8d80M0XfSw3Ao0ummstSDOL8AIaqx61eDHyV1yMwbx2Z2ln56aU5zDP1n
03KwrTYgn2Vqgk+tnEBeyPm4UHMEF1he86bF1Ox24DER+QQaD/CXSlTTJx0JaSjTOaNxCyC6dOh9
oVQO1J/mFV0macMDGmeuoz5tsyI1zfti0d+j5VLTEe/o8UZy9gG3Qx0kjHo4+TlSSPda1QJSPC2R
TVoq43qk5m14UzAlPVJIccz1QvQKIQxXcaKYk/Mn8jaooad7pLej68BKD/WLtfW1jQsalOID7PVV
+emCb+X8AE5dGTW7TEp5sl6E37L/x7fYPohuIyMjaG4xsKMgaHvfM57yFva/76FseEEa0wuedWfR
BWOWCmTwCGAk8Zj057WBGUSpDNjsTljMosmz9S3PDgDcyYIXY6Ecbspm9OG4K0nNT3fmEmbssZtb
eJEcPOzDbvDI+LRoJWFaQ4WaeswnlipfOPkpD3fxGQ7iFVu/NY9aclhiLoZIH+bEhc8tz3rHB/Z8
1hvyRKw8JPntilJ3TMqmhxOsZ/eHnbbVyw5WjJgnXrqm1skr+9STJeGxBfGTfzor7wpEZPfgSTuw
keidEP0PFkExwrkB6Vr/1qioF0OdbDEW44c/fvbrfUJN5OYdyie5+TJzNf82Yb1IZ34VDiml/OsR
KEh76T/m2b6D/0E8s/5PEVdJuNJP1LEwJVbDgbierXcrpsACEOQvVYuoRfbxVIRVTr6rjjdAAcyJ
p409DhrKpDZ4BZrJhuW5EBfE74nKp8QOoDoWuRLnWaMU1suRNHxJ+hGNJWfgUH8PSYRqLJTXCf35
8v06n1ELkTFXprSif3fCcuaFYxvnkdG/oOMTz6DUyi4xvoI1w4hNKDdpiX58ac4rYPu1ooxWj8Bq
7DjHXaxOlpKo4Se6wH61hLxRJa59hTdgVtqGbPTHKuFPbIWsZJed+4oG7BzuVT02GzgOt4m1484I
tmjbcVqaP+M6TpumpnShpns/eHRfYAXPF+ayUKyj+hRvDWAKJaonVbNFB0EA0+T9AbW45gdxHFFt
FVL5Vf0lfBflWxYMm2Be/K67bFIptAfhv8MHflHJMKLz1uZRPvP6SUOgdRH0m2EsLJgNgTENFNxo
IJEVQvkPlx/RjcQbpKIy9BJp28y2U6EQBJ3G+cqqhXZeyEn00NJnCv29+DCIYnwCpoo9FH7hWEw8
Udaxzq7ly65WfIrryRYSFvR6yt581q/fMlok0G0vuj1g1hxadNe9lq/+fbh7R2dPwxdfrxGHQWX9
BABZucP4UfB2lhJfqdqkPt17Tz0GsBQpa7v1bez3IGiUAQV29t/iUK+Tk1P48Op171s2PhMNWeV6
G3F2tUl51GVtZaBh2Z8+FjufTK9FPBVaCyKC2OiuEuOLzslu89Uy3u6U+DZCLhXQyWYCs9pDfMqA
RxCpG/ViEg+H1+fDQ/BSTU1pwDxJfLO9MEWD7hkpJ3mt5YwrzfnVYcOSTl0wvjmLg1jeUPgOM3vL
+V9jbHmOv5sBwVRW77Vo/TdrLI+rNlG6W4qhF3irfrDZkBvyYTOlquXw52vmpMui9RuSAYpYNc9q
ePNza6eOLxbhoAAsZSS2I6oaprOBT7Sy+iNmQlSkHsnK8tRJdv6LpIqpLHUEXtN+D+MVLRlVsug4
o0t00QqM4cNuWpWkRnkpl8VCJnDzQy1m96IML9TU7NoN7VGcATbva4cE8SKcqMWXL0yDlJ4Ztscr
DSzzcduLlLO2w0UdCc/wcvejt1n1LkdmialRWqYS3jUDCIJEXoCn/aT12sibv/ivEuTs5VzVCKnq
RdbyUBHTC8JbslAMEWMlSlVMMufJ5Bmoo58bQV1gQSv5ul3tXda4mYTKucvcAN+3HAkqaUPV60hz
ecp/+C+lflxW71fxZFslHMWg196+NQwLbhDQ90Zt13fBOyejORjxI3LojdsXUiVZzoE6Vlgw7NPZ
vp5C9rWXS7aUSSGWISB/RdUlXaKyUn1Q323Ej1sY387so8pDlSAEV/xDUq9GDPh25w2CY+y5m3DA
khY1rD/suJuY7mzu+RFkALfr5fFYJuVsX2JoADv3gmPyYfvhg2Qz9ZMqCFeeMKCL3k4momk7U3+a
YhS4E8V6eOgD4qmVHNeDLLNJv75IG7TGIRw12ZbtNpH4J0XpFuNOYuK+Jb/EzASXkZRkgWKtCtVS
vA/KlpWMldKQFFQxmssgPLZW/DGjeukAVT1loTSFajT0+7R4CI/GU9eHYtz6+HrZgGXkBNWKTuPK
NdsoTRLkDeKaZLwSJ8oNhel0cXagfOjKq4fmyOja/SztUnRBpS0zPVbqxPJMLDM1VSKH2uLyZIbV
idNbTwrozr2eFTcxkKo83CF+qEClqqUfsyIIMYO0ac4SA8u004aTXrNiceSkBn3uj6Y6qlMjdSJJ
uYAOxRb45IcV7yGApPMBxG5bBKqBoXEhOKslvT2pvEBlFEjcW8Kl7pL3swWMItAFY1Uz0vtaa6ny
10oHYNxB7beo9wpPvG/VCyPOD0WWtjgNJ3tCQQKFPMvdHT1LsaS6bo7iVYb8/GzzOPSmb21h6V00
+Z0PSq4EP8TNGXg/CMb304MlWYIKSRqY7YQ9D44BVc0MARIJ3EvO53TPgd5S1agryqVg4kJN8M0F
N/IfKiyWj2GRAIqJ1IKCO0MGkixMheBoeL4nOEWtuomBqPQUoChNra+g8uYarneRiKJ08/B98cy2
L3NgaLdMjng029OaKh61kviJ1aX5ZlUy3zedsGMjqd0ncRTzteoQVXngKW3nsZqpCJRT6cJ4CA2q
BEQ5tKzEx6Qv0lkn7scI88V0cHosGafNY/qk8LKE2ggAJQVcDm/CSXqZPCL27QUGCTA7qG2C1s4p
KfGw/hgeMod25FQtS3fo1MNb+v26DwsvJ5LrnQUqDGlMEuXE+dFrUHbdAnLQHmtHEuonwT8s1/Aa
Z/aXXpr2npDh5SMwHwV3D616tb2CXMEhEtdU0LeQ+BKT/oCmdGqpVtdulTxz79/RljZ9q2P4m1jN
E0equXVXSZYwuKRGOV/N5prlabrPcVNIFLtBgkLEM9nrUSzSuvC2V1Qgm0dUwmFCYEY6jpQjzTbH
Pt61V5k2YB4JBi+VugoN3oRhXTpRzJkAgsky0OU/q/R4DIxaVfBkNr/zZxuY0iPZGtkefT9CkDEw
ufwyDq19J7OjDC5r1FfcoJARm/zb3Rw7RTdUg47HLcaGh8xu/24XJR5LEy8gTCMq8guedHeClOHa
sppbJEH7y9guBa95/l238pg9hO0hnyTHeVym5g5fjlOq1WNbqlJyo4JGQQoRJia2nQgAGmB61q3p
v3L2WGmYQIIgY+V9Mvwx1k5e/ya5rHJlrH09+hIebKsOgjyLqYu4XdWxRuejYZVjtX7dwUzSgjAH
9DTpbFMkdB4sCI50JMLZ51NUgtK6NhQvku9gl6PypVnuWZG0pAgUgvzEFDlDdOsn+marZZ7mRKaE
2vfsN62Be5YG2rn13eBKfp6+B1UMY0Ov8c9vf5tTqtizHma+/2nnKxS4ncetMZ4ar/hBO/pTGRXz
nINboIJto69orgW55pI2peIIRMzxaFLOPmkxVRYCwGaRTiYb/6MDllvvsJgTv86A7l9Ua2G5S5Ip
opDDRF4JN9ZcpFd77ZKYzIdaXh9PYLe8YGb6dtOd5OuyjDzg2XMRnYWyMa6DTZHV/MNylYVECftk
rwaaO26/MjyWJaZoQIP2zYnVnzDaDPs6bsIQJ/iJZgeRvwoPvC18FaeR0w9tsJBc2gBu3eozaDDo
jmpRdwhidxNVdvQF9YhlX5Qg2m+sv/O2vSLciNQVO6CVUdLu0QEP+xuKAM7r6ARJXgNQ/5Lju9AA
vfB8LjJAtY1Q2xEsMDRH/NPsICyUxNEr3gw3WnGQrFg6sgmyuofgGA7K+pRR6KaWnHUcavEe/auj
PduJbkUbsE2M8zHlw5nxQFA4NAZzv4qc4MVXZVslvPPKstARZdvr8FwUBB+lMR4jfgr1EStMB4ao
VYJZuwkd6VvBFYrMlO1ieFofOlUCx3btJ6/qNrqi/DK+94e2OUO/P4dQi/eqD14TT7B2ovGxRCsg
IfT61cWqxja8jm83XEKxXCI00NhCWETLPJyng++0aqvHqRezSOXxHGTtYToYh/hyPTlOqAAEGcRu
MAOpMDcn22Fiq7gqzhry4IOdjt8EpHAD5lriiAyO39W/wfusU/YKS5XXIAP2RqPXzWqblV39Ul2C
eTsGncBR+Qw9bKHW1pjZSC8lRK7iJTzGTFhuGCbqzLPniAJE+DgqpERapdwxEkdTk54fpxXSIch5
9hv9+Y+4PsEa1WeSoF3hdXVnT08rNCuIYg7t4R3XaZ46mOwB/GFcb1wan/ldRlheaPdwufiRp+6z
Es0tLxDLIKGPTUsuEv0YUxR8l3An4yidK6JQTdm5unH2jEl3ts8FPiChBx3tFkURfyjxzmueoSMd
Vk9n8ooPRs+BVfhdkz+eFAEJ+D/IIGWNLTPe1zLhQtMRAmzfRCz+Le9KzMPwCc0tTAbHNt0q1zSp
5zwI40Xyg2rIojF3m1ScF1xkUv27WcYDIxUL8i5M2Sk8AJ18bPdYPg/naWPXAFf5DUuaVvApkpAu
8CVX7HP8RRFWFWb+3M+X0Y4rRWeK8WF1K7L/PpDxTk7K2oHjBo9yFnM4rAdy+2Xz38TQto5J/+DL
HzRs0/8d+Uilm7N8lDPcKRcPMnxMFusPDgU10D/u+up4CkZSMEThhnVFllsuwMymTB0W6gFThtGy
KPdqns0EBfz3RRWMj9qZbGS++CK1nEDLagznK7xtN4XipIsgAXeUXfSsP9strmO3mqGtLZEKhsaG
kHJLzll2behIguoXgjfphNcZDwHbyi1qI8qR0S/wXHLISbMeUQca6gPTNJZ8Car+JrXGCtEDOKnk
eOUtSuC0hz+exk/GIAr9QK8R98yMe5rJDtnvgcSu8dYTMMQIfpoAXAb7AMED8tqNj6k0uR0a+vB+
rSLcgQSuSbUzsKdJU7tM33OK0uGWQckcIjTHhkNoEoiJUDmcJfJOANgT/p1Qylao8xSYUhEkKs7T
UKfg8H13tWQWG1F2OeiPvqYE/qGSBRo0Yt36hDwZKRW2obaNNli1a9w35sHLN2o8XUw+7k77w3qQ
6PuccSg/juz/zoY30najLL2m58g4VPYw5H0tugcKhhMu2bOho2xgyB81UYClGLv/GC7mZ5jOhAkd
5YRstQFKLIvknyov3fybBUoV0zeHHYixddTmVk0XlLV9TRR+jq71oOyH3fXJGUFdbL2T9MDbMyS9
z35IYpYnLI9F7i1VtzsLvHlID/OvSgKtWW7eMQJMLv6FMxS02kekUDbPJI6WZavSsMDtL2oOcmHG
LrqLMpqhm5unrS5n7p7KcRvh2M8qcWlwIJBMg8AVu7NKmmsutWZvWWt6wU0fU47cGO0ECkD2plOD
FNuSJp3T3yDWS/TSeSCqxywWqBBufoLEEkBrdMRIH62hzhHfRbeGUab9I1nX/5qdZK+9W2YOkA2J
VXFbeYiVupOJNrZsWjIRAKNXfeVGZBapMG4cnDt3nBihE1gW/D+fiU5qDnHvzTxtJBu1hu6lJyDz
yFb3iFv5wNNvkInTB0vPvvumF05/OkX50emf14et9y9NCzAGTRUYN/Z/LMjMI/4i8bTfNxZMUmV5
q3cXZaxmTC7pvoE+DKTa6e4vfWIplgqBTEhHvGhxBjtLBdo3itcyFwGC6X6cUFZCPTqskLLZNbu+
9AI9fTipdC9HnuIM6BRX4HtulfrqOjHg9ezxw7+2g+XPM1QIWLEvXYBl5MvlrUilrnrK3ZaxZRqC
v/YoGV0XEwm+PyIopyjT0faECWagn0gdk/0Id3pJpdbec2CwwmOw1GXGKqVgLg/ldpRGr3bLyF0S
CwzZSvQZeXbzhHBlpi2xCOgo3pMs5SH+2LmrVgHgtDloSseCpHWYNPseT7PhafmZYc/ch0f3C9pC
8Tv8O5xlk+R2vonutOdvb6c0yErNcHLTTZauWYo01iTeYIS2UcLYs4EjNKNeWQJgzKth4dGZdwNT
X5t94KFqd+lKstWuiBMzODFCv9+SajxfkhS3cU9A2hD4HiMF9s5Co1i5/mMP1lGeaRCeAgDPgT6n
FQ34NY5pIByG154WIV8sOGCuy7RFm/IDBgCMB8/VCh3GmgrxDOi2eG6b+uvRMV9jJ5O+z0WoSmN/
PVjWxi0bTaDJqZPmmymYBJ8iM0UdqVAfLfCK9uWenmd+ZBqgfDN9a0v4ncVUfFFCMpJIZlmKmr4z
fZqdDGH0JA8fNspfBNozQ6uzTBTFwHSLiE3VpxmrX3h3nLOhn9EHZeE/nde6fULtoG9rOJU6UryJ
sv87FSFxeU/h+Yx6+PerVQZijITtcRPUCX7E+7zlKWQfGXISXFnVri4lBpgomF7To5H2c59Fs517
zCj8ikQBJhyM4EOWTXOk59amhd7xN18mj7SwPhxZp3yuWKhUI1l2xElb8cjvw1MakWM4YAdEjDX4
EqTU2fi8ulSXIJ3fwoTsil0XohpsYxSOwmMauv3wRIR/6D7mn+TdRc51Kkr7UY9eZo0n9E9GyMf6
p7tMb9D8HwKIVxbiS365EdX5hmrcXkOOsqqkgYv8v2ZmEJY6mhJkazEZHqOfluL/413oHX8lbfCi
25cRMdG6p8OJAH6mBaDeHx5uHldjR9QxggXMPZrYpjeiFwYRflw0YssnoTzZIOiBNvNyQP27u8zU
OhW7kyi8zzqF53v1rYK92wG4l7W3LdDgDSE6elTbzBNcEKHwQRvZOJLzuOB8YOKhvnRC0LSyW1db
7+ipkxEENefHNxQMfqKIix8xiu+bo+Z/99OqC7YbfLJ4jcyV2R9AmTw0gXFbAd7sdlKq8JQ99L4o
d5f1BavWMChErXVBjeqgCRgMYr5oscPV3fXKe+BCW+79LJdojACxqyHxC1qt5ZgTrCs/n6+wZ7gs
yc12RQ8p9FcgjM4FXUXUjwq0b17PsVyUISci/eGwWL4StPbUZ+HiDf06d8pNX1r9jXtv0DjaT9Do
deOAyvwTWYxJU+jeUAkpT+KJHa8A6bmI+g/j9qFUz9IKW//Ppe5oT2m/42nWsf1ewLwK+CHwfhRK
JYokhxiWTNz7wIoW4RAaCmuRCNjIpbL/b8kgoOujKBMoXw25L0uIq4d8A5w5q8EZuDVbqkuyo9oh
kixpsOCJ6SsHFqsADECs2wYJSdUqTx6eAzMN125R3TBh1ex3Ddi1/8kEJ1cJTmRWwzz4qR2iYkNW
GNjifsYyeIM7fgKIFs3L/TNgsFGGX/b7fZrgkTvmJBMYUXMNv233YU1lJVBSuHpVfOjpv5SZzIzi
XUGqRekNwcdpp0FT3hQdhhcwJcUAotQpSdPkV9QT9PsvqErIdt4hNyi7LoRHfQMoBP3GQP8reDtt
ztld1vwJYJ00yBtA9B1dKNNnoqEhv0thrrd8ko9NnqYvddWEv7AKqmeAj+KfkwaCGRwBWfCTdYIN
JL3BqIp8n5s8oxkMp/qqiPz9jLwFvGfu1ueXBVYSflNo61OvJHzwCx09XIvzABE5wV4izWJWB2rA
ru/D/EvotEyu7dmQ3qr63mlj2Nb6xBb0OQ27UivBZ9/IH/ZVNgczzXedKt5+PTeniuZkKEUq5H9f
XDzB1bbrj1hDT4G9lNn+NdT52z9y02iI0MF5hWupLZqFICWzaVTgGelOy5CEUAyhpsmxzxEdyEfJ
XAT6hdnuQnTl55Ruy3gWINpW+icPTci28RnxbztlwdNyeHX1+teJy54/D+09rnUjaKrnu1BU4zP5
QnQxthzxzDrl1TsqrwcRdJvDpJpgSP3rJrpJCmFtLwQJ9ByiQMzyaStrpAs5CHhQRi3D4MdDCZ6S
V6n8pG/8ptg4fJIzPNsyNJCGq/v3iprxVRac0MZPjzi6vjZCd5HgbMLONdAD1b+R6Ee5XgT30jZm
2FdbrUBRpCOQPxFDsZqxzXGwfsBOPjzbPBh9ZxwF6uqQqXfPwyDWjkQxYFwTk0dE5fCG0kBQpgE8
T2ieYqBr6WjU6Xnk1ElYU3f7B4DoCCX+1K6e33que47L5+63SIJRKUuRnmSvacFHd3nb3guY+e4m
MuSwiBT95ykw21KU2Rf3zF2UHWMEubJdgqy2pqH+h5IqjNPcO7Q4yt8t6aDiotHb8wieVopf6gXs
KTvHzDKu/1VtlRoHsFbJTIeW4sfoyVyetxx/iqMtx1uV7lHAMfzrMQVayJomP8wQizSWbkSpvdI3
IRJAWJAk36/MrpPtewL2NSBoWq6BUpe4IM/fVSAG0R5LRzO7/brypFyZsenrZ1Pmqx+1po1Sq7to
aMDvZBJILFS3U9m6lzQYLc5vw1ZpyttQQ+tll2xql9TrqJtFa0JRqhZWdivbFeZ7Z9wlurdU3UjU
Dmo7Upnv2ur6efc0qlQapW6lSWQrwbb6nuoqiN/6KFjc6wiTk2wNBoIGW7hfywpy79jkXstLa3Vj
RJd8zb+tAr+Tac4csd3IPCRdxeHlIOIBhIKaENg7TAMNSSiwMRHbrUobNb74oGNCJK99EgnBjWkP
Ag8RExcj9txFwuQqEocg9+TK0A1RyDi7j3EoeizfXewZc7+mc0LT9d250b9+u8AZ45pzSHzYEPPZ
5fbxfp7y8IE6/XSO3cVLLtqYgqOeZUuERo7+4XPlnBUEIFXQTninQqaJ1hSZnrPC2q9uftciZm9W
KjaEclwoRpP85LVgah4eUTD+0pnblznqSXmD8MUW9b/8loTbo/Dyxgr7EJX7dvxnMkXHvQ5lRlbR
pgAxfcDYGD2oqmmBbsmDh1nFgREKo70yuHlFu7UKOg2ONAak3vaakaE95SAJlMIZQ81XkHfn1ezf
FMy6XYcXvKiUoZ1pZggGdpoEkP3fI03JwxQ5Zw0KO1PusJp5lGK4p9hsXaiDCYDng5P2a58tnMcU
omfiMgry0Bawue8W50s9famjwzoDkgfn3IdtBq1W6NwSQ71KmkjrDUSn3Vzq6zJWLgPLIA8HVfUv
mHyjaC0B3ulF3Ys5vX1XVYk2sYUt8dPZwT4FezBQW4A1g73bpasOT9ki8sbgaIe/NWxlPaBT8CIu
p6nJJMUoLkwe8GtbfpjXmnTahdrIfvHRN2AppLfUmdDrpG+dywQMfZZPdFA8FF3Z9ffiw0E+wqeh
XowLfdDe3ptSzTvKbQ9mvB/ggqQo791MKJz0fN2DXEQym29BPD+6Nzp+EpX9L697Mio3fgOYdN4b
cWt1BCwSEpYZNUkWddg3lYkq8xxvbmvJ0OtwmeuoimspHyeKXXGjLRBdgrANHy1SV6GhUggNMnEy
kgjAHaS6gsD2Zf03fC7LgEpaorJWFxjbYS02umRLl2IC9lVh5wzasjLz/sZ3MxFWZqz8xwF7ufeN
06szLlbtp8KXDe1dcHVhpDa0nd7+bC2Vl7BlPBq2se4/twrWXxWuRp1dM+nLzGmQM8CHiVvKFJR8
mhg4KBCQQVYCtkXxkvdmmaJy304Ryfg5Cu+60Fp952LeaDe4ByKxSQ+4wSEuRYOED8Wd/MIkdFaa
Zb2Yulr3abeB04g/gVLXw8otIReAxEBLlR0uaMKdtuIpjFISF50O9Wb+KzuQw8/JIh4LVyYQfnMr
Yeo5SRVmDdQe5Q1hMfn3CDjQFmxiS0DzjBtA2zQfAb4Fj8WnREmHmWiN21S99bQ1z7cK8d70b5zT
ZbYcey03ySmL+6C/46E1fuNobvPOlQs3pFQpDvuQLYlZ2SdAnCn8H3mp+pkudIQ34oWb+bZmjLgU
74V/Y+NQ0w62+h2ZWnhNPU7rUOx1weUhBIUhtRAK/KVcZMCXDaeu/ebEPpu5OcqEMFpvpR147f+w
5lgtVkG0xm1YY+1S6G9jIPRNnaBVOAXqgeTcEleaCcpKPd+EixDSHea2BVEmtw2SjlzM0+xTAwO2
1b+Wlj6ZB7eQDfUQPrM28zDRSFR/nLW1JfMm9SRGE8p18FZRvyRGoO6W2FrF/Pa/pBbFsdKbR+pR
2eKX06FVqQ9r1HI2huLAufxZFA3XNNBGI2Ke2iC2CXb9zagVQrJDi9I3KJSJWLdhCVqrUCXdLnYv
YUy+DF5rdExvZ/dajKBinAKUqCvi2SMiFv+PP8B5B/cFvy2qiC8EfS377DC99NK+zr7qWUGFfW5b
YfUtP0nsIXtb3O0lAAH5F+KAV3vUrSeHB9gncWcd2HqM+bTOrlm+YEwFo6xEv8J5ff9Z4dEvpzXm
hQXKsuYYFhXXELGBdOaZxAlXpFg0Xb2/4WokSyIA+pWNo3gUNfI35mysu91h419s/2aPjAAH8Dvn
EU4vcr7ZX+LkHpKZwBKsyxKf7NeruYDixqZOcNVmbwuV9JRnF/kcvnHWTkdTb9bkOVQTKlelHO+6
YXxI+MgzXRZLTEh+YRP4WyxZTlaJTY4yTb1FD1noG87J+oFGRzzlUJa1JyNEkBM6algsqj/239th
NQi2+sEn/TS56uZzYt/zY5Rl27CqBfinq8RAwqivqMv8T26pjEFksh3ccNmRpC7g+gCquBriWN0j
sgjLg2XFwoW2oLeLBZKs/EKF6A54oI/tssvNyYqHif1bMc8mR/3syMhFSxlsyGuwnOLWZGCub+FK
W2v6ZJEbvcD1sJu00Xlu5QMsZAMW89pS+RTSUHpzGkbYwVY4cvk70F4vAdDvxg7PqDb7zy2ckU0R
0672x0jZzQNq88Ee8ztCslm7nDR98nus2NZ8iqp+nOgS2uC5lWl+YuzyyAcCL9C5u3pS4WLMtdl0
2E4wQ7uOK4rQtXRduDDbpqG8ba2v9upK37YSX2MKAbyIwysv9qy1QcZIEvYFDEiEUDspE3ssWzB4
SIRbSm8oNgdx+/oulVf2PuS6Mmy2pmizchdanHVvx4Lf4isctWoyOYL5HZcKWu7HdVyDmQ2lrNH9
i0b1lknDAEoPfFVfDi7TJhPvngy4ql7MppRH4tcCybgAkeu53/5Xo1fvdua0lk70iQV5D/C/Q1qc
9/UJpONDzxzdkc3NW/u6+kleYet1+C1QSD5+G3ZXvtw2uwY/SWL98vRlf9D2W2lNrgLJv2srkzHa
TYpCxixHVB/2y+OLopXzsSdQwyOQicwH0CwWxgEfk7iE3uCPjPJwOe9H+UzZmK5gjj6a3XG8etmT
QUpEZDOVDRJAoGkBAHjdueSGLANuoFH79/GeqWBiP6vE608eE61/WaHNndWf/ahtlaLXslP6Ydq4
5DOohzepPbUltOlegSQtKDZvkGOCcEthEZlAOUMXtmI+ozRY63M7+YE8fLap9X/IZ0Rhii/wCRJO
wkyOpdh5Z4AKUGm/r1PhFwJQrkWKZtef+czI1BcOzp5MYTca2sJ+mzhne/zAw2urroxU8te2NJK/
f5kP+a87OoIIDshK4FnQ/+iaJ2mH+ECwDuBaVF9G9Dcoa3tm73G5N1dxnT4qFh1qYgAIAhXPAGI6
RlhKwzxKSXnKa5NVFOkQOMqH3t5qPQFftorDbVBlBs37baXVTE2rcUlTbZtyHkkUZTSv2q3EO1hQ
ztmc7l4wB+j7OO8U8ipaTrBZqDb9HOTO5CCuZBIN5gHraA306dyMWwPIW6lR/OR9cSQNJ1VYnF+r
9mcTdTIxGsDe+cpKG5b1C2zFUalV9jEOMV4XCrmADessS21F1JmENemXA57e5FjUtx6B7ZbZDN1+
pPY+oP0s8ZT20VTM9p8o3rtX4vIVV6BOeDX11CdsEKiOv2rZ4ru+bORtBayyA7S1q7MLf8/Ivq0R
U5bAcCas/F+dVgYpcNxhUIEk41hYmq9kE6X8mjDAXD1YuRLWg36YPYy2lnSEReXWJ6yeAp37AQ6W
wZWE9eGPnX9DH9ZzSdfW92polJRTMAp10jZFTYeInfBgMQaOge5rsI6GzMaZ2mZlI4La0eoQBmpx
wPBU6WGd/EtBSNWFDv/+olXNU1tl6Pt+FmliG2IQSjpAueC0QvcQPQloqQmaTkMh9TNECCaXhqV1
lWqTk9fIYakqHBP3oIJh37dxr6+qFY+c4aI1JMw/iVxMrgDQ598FaeElxIzBZyih+f/AjbJ5HwhE
CX82b4NiOA+/vJoPr0zdLXv6vHXgDFR/1gwEBQ+kB+9eOnw4taoAPyqX21bFHgHP+aL20m6jOrly
KR7pF1+g8xuWFtpn8IP++QeiqC2D2TpqQzllhz4IJ/vS7RhzQOenLee4gR+9V/N7FKnMNYmFog/P
Th8K1Z8M+ccWRSJcs0KdaKHRzobS6CtDbGgtjvgmvzblG6u2nQ3+Z9e4LqJAr/enIFYPet4JhuS0
gFKGx+bPyLERn75tEmJNGWLYpes7Ka6qkPBR2DhjVD8v2r0wBQG6Uc/nzgELdQl2iP2xflnR8cpE
wkqhVuNGI07cGDUqNlhv0uw5vN6wmJB+Xr2Lao6s88l7rOKHgiGtHOni5JqH2qJ4QmTuXdfbp8hw
8u7YmSSOEyJOQGmMZe3ehQZjZy9Gf5VnG6EZXaYcNeEhILnNziTUQvFicp+P39+Res7JiIuN9Yo0
xvo/+sO7HseaC6UWI4rq7viFtHjdp/KplDQ1hAIKzVgRvl3k1yHjAfWYoh0oNC2Erw6Twy73RrEp
eQVCrMbkgTCiFa8BqNyyKQaYJOGkOCK5MNXHIqh3hfhj+nVl/OuupHqDanI3hxcZX5SchrEFMgLd
IIAJkz4j57xbx7/Q+1GQNPleogFzyVF8WaBXK9RgveG5T0JLlvgngRubY3QYmiT+BfgRFkguKoQ6
CqOsUw9Zqv3E7Yd9AdS7PbXAkagnyvXJpgUZZNRXP6ae9U6UyzkxSfOJKhSsl1a86aY6p0w4B/Qg
xWjsnOQvibk2GIEj3yJ96HiovSPuOjJUg+MnRER8Yme85LP/c7TARasacL6x5+9F6CM9owQd83SP
fc3a29GBhvb/PHhF2Tu0jF7BA32doj5fBmv/zyPFel+CFaYS7lEDKUaQRZy5nk+KGgmosuI9sqoC
p7O2Kc5NeM1dHexH4b84Nzt7wG3Kx6y0Be8Hjn498olgJLNeoovRBopZb0ou8qVGH+iBWlaeVXV9
FCyw2tUvF1xizJiDB2YflCpzog7tnE/NC4gxsmG1Z+QCZy8gc3vW4LVh4yZRXZZrwRBNvl4jZbCT
ABOVk7MMx6vDbVRQATqsdDxwl6Oj+1GE0pzq+gu8QF2Q+eVZInGPhqeGLbI4dTpkOxfi/F0adJOv
31zPfGDwCamUKOfPJ4rB22SXdEZfuDApkfmRjuPLelJPO+6TwMqLvcdgHik7RCCiaS+3haf0uJ7E
3+51YlPNJnKekGaSFxEu1kjJqASsVsuAJiDjsdY72u0Pva1TeDW9NpHRBwMyGg2dZ2pxwlIs9+n3
1eqf6JktT8yFn8lwQ0gKpC4cEYmuy7NXi5BSP5nuSJWDcKULH5m/Pmls4h47K9lanpRNBckV1NFk
HXY9lez/phd1ggg71+Z0kk8IOZDh8Db9Uul9Ipp3Z6bTSid9U+r0WggLZ9DJz13w+BThq6HG6mYL
GjJoKeQtQ3RWeph8IYi2MOyfDoBBytY6L4fTxFT3Vf+VROyp06tgKU/nN9+Lm1BG2xVUSiLOTKfV
v3XQCSwQeP6W78Y6Rl80vlg9N7M2iksCkL8hpUw3t8skrzBbK3U5iJg/OaeoiPu362+wUcj0KUMf
+cGTUBFDbF+sHw10OcMF8M5WjW3F7FG1BUa1TWncej8E4w+1X4Gy8yayHRFc829j625GB6zGCuMF
U0txBCDNwhbBIA9GjnydIHTaXvk8GqD7eaxjD22dIKxOLEGLmw7s5cqOM/euxhXXoYhkonL0XcFO
mXZrNx+F4AXZMwc/4IfS+4b0OrslgM0+as7zHP5QnRO+Scdi+VeuG7yTIAtGf0u7b35/LBSSuhiv
Nkp1bxu8fN9/qb/rCmSX2SIbHi4av4iGo271KjD1j9cOFSPjfbc3/kVvoB9pLuoiCBkZOLhxt1ml
5raW5FTY0SxvAiTQbv0SGv/QSQNHPiG7qbZWD1TLNY9FqOjRUh26siLvx9yVccut4SrttS47h5o3
TesNDEbeJemhy6742TvIe5qDqc0ha6sSbQvF46rwmk+/BQlK1XE1SOHy1Cx+TXpVp9KKi0jWzIo3
DkPXiiK1FaNEUMS8gJ+JgG7vWHmyCgBhj1Sr0f08jxER5AqitUP+HHRY6Mzm8KiUr3TO8vXmajAw
lOhwklA95O9YwiBGKACzMO1ZUcVKa5yQ5mEXfa7RSpcDBX4YrQq/pfQoOQ5zMkQ18TjXegJzl+W5
9yTI410jaSACTaJfb+9q1S0A4PtLRRXRoyxyxFO5kw0TtwtFHWnPP4oAip742Ynfd7V2yr81JD0H
0K2VKyEEwSiYrB65iu6cG+z8odvl0Xczm3td74+UY+xuOf6u6o169YK3pyXpZkR/Dx8Ff2sgaFWZ
kx3439BojAdaWqceHVQn7gj+qJKwa5fAzoJ8OkOAty3xjEXFw+9qZ6VH9r4MwoUyhVk2s/dfBT5a
ozuC27ytIMAIAga1RF2m5hy4MDOBIGfJJvNko5goMbdFZ3IT3sPUyEcp4KjNA6T0FcTXf5BWEXTK
UqCPwIzX2O4lOcIuF8/4b6NCjWATUDARjMB/TH/La5u5XmbsldgkBiZx9QKmPOr9XzyGyTHayRTO
n0UtWpajZ9RN0ag5oZuqYD4tUwr6kZDAbxKF+ik2VgttZVkPf6pWKb4hwvb0KoJzVEY+nIZ7fIDI
c+YNo/x3t1NzUUvbSt9I9PENUQ99dMrFWQenhjlazQEEnO9pO/PD0JdvhafnTxdEFMpQv343EXrk
r2AQ/hv8Ehbgh+aBzxVgH+GL3PoHwNvAv+8vju9aaCCkze+k3M5Yh11/vsGW1tCqMeCvyJXUlnsg
Mca72FrfcnULcLz551McV1WflNSfYlY/mLaC5ofw1G6eUwKNDMR76zQ4m9RxfmE3IY7E3aBuZ3jO
naL1a6mkygXhpTDUrkmzmH7uDTFQHU8FvJ1JcHOEb1pAPvwUDbSjZyMcKRSNZKkJEGJwDShiV9OT
yL2OMYR3QWKzd/fgl6OInZi0YAjH1G2/ajiO4WbfofbpGxQTFx2mLd2ARCKsaY5it7mzbhBKWK+4
DcIYF4z2jrvW2PS1iUfPnlpDjPY0scL3KUmq4WNNYBF7x9Yoa3Wq7v5vKEM52Ljpxv/J3bA2l9xU
AyaE5Hxb6l7OU0wT+/J9kqnJOPZ4PHKDl16+K09YnGAs7OZujHIx8l7xQxmlxdHqPOkMZqY7NyJz
ZhksH4pP75hkmZzmtBLMm6nn5Mt2z0xav9Wky3aiff12NQP/ob4Gvtcwb6vzoo9SCvYsza09pj9x
j7JSLAtfGvQv+cMvpVJ59NzMz1q101L8TF/iJRHG4oUCZ6xFJFrhGs1w5fOyHzXwIy5cL1Qz5Abc
UWPBL4LfvmQkY4+/h3CxLBX6Pwpawfz52K6VogqBVscwMR/fEHLWi1A+k23/tn4t1mYCuu3aTMuL
u1M42ibMYsAIDbrpMMvlVjUaCAFqnffsBWnOKr2SKde+McDL21OHTfc/e2bU9fZgQxHGyli2R2lL
FPk5IZlJMkbDXza6UIt50HN6NxawcE87SHOuMf9MUY7nUHG0k1d9wm774OM0x+s6OKK/V2gvWoJk
T6IpuH1QJdwoz2wpBTiIkbDUrND0ra/jBBMDX8yhcPu/++6cOLrvst2No07S21bVZDlTMbrHwGyz
SRxOW//hhruUDd6moOcWiCP7ut5DBfgOknzCyum0O5Rc52afUB3qmU58Sla2WRwvaw9rg/bHnIGy
iSFYiXNFlzT7t5Cc6dU9qBAhTbOaUzAG0fWp2PJuPS0J1dSuwFwiqO9XZCGT2z6O9OTdbcRBYlJl
u0ihCUNc3lQs1N9feSff3P/+uQs6KBfAj8CVlTADw4yUvqfTA6CG9JUrXD2bqhaHN1/bH8ghwLJV
BHRUHpacRgmAvZeLHACnv73a5pMLTqNQUNs9QvcMvuAyiFz3rCW++qK/0Luw23kKqxXMWeu5oAlf
h3CZd7YwvNw345TAcwzpn/TAAsksVhUDsEHy1xa5V7648NrpkDU6uM87rCnwUtPcVdqC76VUGcCF
ML0zSwx7UZiiJ11imKoyKqDm2uh5U0qPATM3/fqWVPrnjs2Igkc2o4vPjyflw021hXcBIUw7K2xT
2wdLP/ubZ59BEyX5EpidU7GvBExHNq9UByl27F+Ic5Awx56kEbbppSHv+Ky67i7sRqBEZpsUuZOs
Db07H4vD7oNB2UhBAZ7j0G1eazhxIrdvVs/8vBi0yZ3HtdcSaHuxL97sx5GtYczvJj6/I6vzr+0P
nXOk+1QZEL3EwCeSSNgdSbEkFB0W0i6Id6zJvH4DbpSERMqfKVRrS/D1J3gPFfYbpSvV2AdQvcS7
UypYwAh8BwtQtTFbJ4wZfBpGScjSysN3gtVmbSlFghXHzbbDYIKqDyjtFJLqjf7H1bNJc6cztuVf
ARBl2cXNd99j5DH0E7FELMUSR902b2aZXPJXduwlXxuXRq7smnc1QPU+Zv4RXZyoi1D3q+Ymp+FS
xboh8wNkGzn+yB48Eu0+Hg1E9FlypwvoZB2QKWb2UccjtjsGakz/XXLSL2NScssgGbS4FNQKq94Z
stUU9urj6zj+TirxWjxcTto1qx9/wzZ5wzUvKHPIeG6WWbpAUlWQ8/GmKyqCPWbxiNsKBod4dF9A
v1dYGH5nU7rfm7ZEco6oeTkTunS7LzW0CGx8N2/Uafcf7FgMWFB5N/b7bsP9zr0IaawiFoNNpfRw
AlxwZztymb0QdaHHR8kKQH3Yje1SXCuxUlfMfFSvkoXCmGYAVNzblbGY3l5B2iWNUb5HoeqzbIQC
fFtcmpOd7VZYXSA9poyvb4zK2X38235YV5Ol7Z4PjNnae7nNQhbjtV56qysiV2hzaUVTI53HEd8T
Zrqb0aN9bdBj6sW+2E+fi4VUMX3fZW+e99GRwSicSsDfkfad+DiP6ty68FVntt2BqQfOVWGKIS48
yaz0xxllf/hmlF/Xu3jvhQyxu4zQcbdSz4l5NtwWjcAW9XZTuWAZxCcmj7CwcTcpd2CgAKrhLyWG
r48Y2QOejOrVI8OwlQvLIMLJtD3bX0FvzrIKJVehqz4Vxc+P+CfKK0+/cvUTuJdUVaoBW9TLnKZ1
8vNHF7LaiJGYGECPloc6btmNzLpZWTLCJd5ZmXD0afZTyHmM+xXaXY00bOrLufOyhI4Qp48eQzdQ
BGAijdfecDsZQ49yyhJ4NgOscpNdUHBL/F8kvCh7p7/zE5De8q2WqI+l+xGeAxpZzVleR0e+wMnb
KU8B69D5xS2qimczvxqPRczp1bEU9XGZ/xdRJIWyCTCxxJhBarOCiJTr4fCv0nsZYJU2fj7wWM1v
i+RHTiRGYWilwgDthAeJ+6S1GZDzWxX3pmQQHt3S0bxV6mRWg2sEU27qZsP3A3u3oMXIKTk3ME5z
QJzKimmGtza21mBU2lAd+3jV5bSEvt9Q5hEko/Pf0JfnEkjYVheVe4JBM/Dr9o63NEJ6UJ3vZCkL
rEUFUJ8xHWZRtNVFXh+DO8opbulkk8gD2Y6jCsnX35uPinwEtSf+5zo/ySDW+5o0q9YJwvs+vHa6
bmG8k7R9depbJsAIOk/MNB0zJX8QwqzuRRukUh5+ZqKR/6nII7gxUA3LFbZSnT4dCZrS8SzlyRTy
oe26C6UXbabGz4BfU9seRoO0SN3FlkpgjCOv5NjtdVhUFYIAnQoGWUx5ZNkqdKq7irnZlU60+e3Q
C4PBfaDwq2qFFg29PS6HH+LR+vi55ofqJqPHNHK8r4J7IX0QvewgoXppLgmuLB7SRE+IczBVidOW
fFL/sjoLLoFBAuYgCoS/NzMpb0c/N/BIapLayqdDra1siqD0BmL1Kxh2QblG3A/9thto7dYJJf+Z
e7s4fFGhvymx5PyeCDVL8Xv1ZGUY/80XqZDpAyzbb92HGwWj2pO+fzz3ksMmawl4X4m/JInQedsY
LCNbSjVIRCjcrVzrUWtJskZ46Xo9m3JeEOMNUyiQUeAB4hgc2MelTkFZ1TsdLVvKxJR+XjUT7KBr
tUeMzySx63Pa3BNSafODaUqk50+2iLmxKelwiioPPAodLBOGlqg4aFnRS8UjnODaJlu+mcN5Tdel
e6hEBD5Jqnu1rn5zQAnSZuCZGbn4vDV3+m5kZKzTl3/tVaeRmQdHvqUS2XsvHlGoFCO9AawHcvvP
7lcsKWR8/Pi8pFwgzawuYSbx5vj3OHRiBooPxJBHemuE6VXbHV+/HKGuvIkuGzPnHPB18cB5A0lb
c9tioaJBWu5GS13oI9DLWc3BJaQ4GdfhVm066UcZ5dE3Shxo2y2VHI9c11Ns3ajEn28lJjAi2rox
GpKG+zBRlnYxy4Mr3WHy8m1OCmfNNKxLIjyRfD0GKS4Kgfc9+2p8fHZac8TydLeLuZId57E7vOPZ
V021BuEn/ccTEyTFZp5czBQUKE1MiZ2f36bW8zAKkyQRiE5nZwgjEeGVvldbpkKsSlMISGOJ/Z6F
SoHldWPTVUrDNYjfyreO0zZ5xe8wCaN+iRzVYihXuNx4BhhbIIl72m171mi7fFdXLwCWOdC1gq4I
Y1G4/4O7sEIAijmVChQbmhrE9iDAbaHmRBUg88Di2L7jucZ0lulAsINL6xdM33xDAA+GkuBGsGoM
kiFV1uvocMQQI2BvWxV2/ImpPEQbXg3L6eFqeBftt4p9ZtFAzNH7muFek7M7DKfGhEFi+yhINXCn
cHhYQCS/dpnxrjLEYb7QaGfjJhRyeI1W5Cuuu80ZpByQNNdvmwWZZ8QmqPbr1R19rptwkGB1dd0f
XXKaUpgE4K5FKCvv0aqDJYPiiWoVLGLlRkQtCKkg8gDR8guldbkD6PPPPA9sJpHYFF2kSwZ++9MS
EdZBbke2Ema/vXa/27YhTuy0MzRcY9UFrWZYJ2lS2kJ8QKlCEhLt7pQAXTaQeGcJXekhPz7x5RW4
+tT670AQx3R3O4cpjw4Zmm3TVQ/AGYyNfuTOSSSrXCkdoDyEz+cXmObnvB3vVtJlqRAAv2cjdY8v
rcgwp/d2JwHU2JP5ggi1Exf8rpkVEOPZyd/8DmeIugiHYYqjXknPHNbK1DRTUoGXvWk3MWEfG6DL
2Y1W6V8r1Q8eOXymhmeOLGVALQoGLoDR/5xXwQp1UEtJHcN7+L6IVdtfkj9yGCHErcSCk2pm6Xj4
gLe5SArKly1J8jmLg6vPGvGrGq3rQ9skC9tydGVwWhO3P7BC8J1zYciJ/DY+vLkw1JF5E1RHX9li
GB63ri9bMcYgSOZFVM9In82ZJ6aLEl6PPSqGW8ewLgK0bVLmtOGFqoc1ID+vQpbyQDRWmOARk+cO
iUCMdvThK+arFRVkISLUPpabm3bIs3TFM0uUponB2Al6TVLVNuCELs1exoe7ISxw+bw81OeV8eVh
D5NTZNSfn79dMXgaARbqxs5rnzWO/HH+F1fZjjPLrNabLtNo7G5mgjF6lEhZTvb/9L9sEJsJSRki
qTmH+wRnKBXqTP+0dMGv9CO694HJVkgPrc+kewjw+I+F6GNTLBNqMQmiogojn4Y+/J0Hr4XfnG97
ZHvmhADX9U5QVpQFb+tTvZl3ayzP3vgHXR02BifEWbKxGgUkGgu0Jyiaho2l5TLigdH57w2RaCrz
p1erQUwbqkQp0OoEfwf8DBePWr0FkqWopRl/rjCJObsZ9XnbMaW6bEsEF70VIxVmCXi8rbiZrqJg
UtmWuF2fmKy70MLbyIoJeBsKnsIy5dAs2bklnuqGZB93vOuJl4/fw+rfNXhR9PhVbfwsySlg/DDs
KpPsAXd++mkdIgQX+4fslcRBXNyC0hqECOrIhH/sUO9PITlTidlAB+JaMCPs2AM8J8o+xi+4CWU3
QlDZJXDGC6hglddNFQU++arPCO/JAqf57QqSzTor5QPdBuxNd69rf3QkRjAvx7J9Qt4cEtVt3fFf
PPC3yunPplunVZbHdSTKVwuZ6uW7HqzH/F0wWZViY+UM9dzHypHPD1iXPsYX0EgZ23s8yGobg0vS
IQ83yWdwP5p5Gs9EthbNmi6I+81ZIZhNER/ocJ5iZxgzB2VVjs3PmqVWi/zWnAKi2VPw7CeSukkr
Rto75wvECi1o/fm3AZTAPLkqicdZniYVziwygZvrvM3tjc8ubAmgqFQthn5afwi2erA11NVL7LuY
iwYk/5zTfpXpiA4/ijgOwJXwJcWIs1DEJ3T4F/uFsHq5QZICORZ29f2sNnIhx/gEQQdFISNCmg8h
F9Olr96EQr+3b+5lW1sJPB04+XYei4UMcWNdt/HWejadgj5jRsfQ2tKJLqn+4Lt0BQQdFP424JIU
Th5770oFMyRy9Zh5fgO/v1t6QU3RjN5t2+nlEEUT0UOAYHCfdXgkTtAVJcqzP/gg749CZ9pijBUw
ZBRkEC+t1atmKB3I/j9ayNobfDCNaTYpQVRfPtAeCep2c9sOQMeQh17kkA0qBWlUTmYPZoV0Q8uq
fvINDj9faXflvp6L2IWp4DSm1R2e4aXjf+uwyF8iTss83DneQg11GfKLaVPFs6qu97ztBO6uVS9R
tiX1/jdoLf5QOokFAwev8HRDVhEDLFCjgpdJrOuX9NWZIVgiFrnFGGEqsxavL+nqeTa4rhLyjgRN
9QQVNx3RLc1TsrCv3tf/ddKth/V47WsKzKDuyrzXS+k4YlJP9bEaLoe96SVoTVaIRx/Jz4CrWiMk
ZhlNkfTeEeTbvchnB1mlxhjmQhUsq3zxwB+vglXbPWzW98O/mCm3A7xBTARxkaLLhRZjnGYRgfbr
kmQ7sM6kcXUE5/5bm5Eaf2fUxRaC7rWPYFRfsz6MYtZrBS0ilxSnPXewWLZdh4dTFfTu0vqWZQqc
Lhm/HPGYkYZOG0h02Rpu9gVi4Heimui60dZBDaQ6+Zy5QjmsPkuxrn8vHUBOWw398X3PBbzbKG3X
I+1yIJ8cbSMIJyL32LGYK2BT/AFDeAcQPRajboL5AzCH1EkeW7Gi6Zmn5GAhU/BRsTg2ZDW4IgeI
sK5hU3Fwt9LXuMIiD6YRLFDJs6FfuXcBVYfn6lU4qyJXri2WJ5cbsI/7gZkwu0m7N7Uq3708wMGn
rpnTHHl2ylZWOnA7iTxjwyRCmpDDFCTxGAD7kiashJyWnl9XfBlMVAVIcuEb9HfLz8XFC2O4NKYA
hvukDeum4ilRuzpenx5CWnfqY9tJYQH4TGOUCVeUK0pmnRREE42oZVskdmpthxBF1xwJ1erlxqAq
POevOcresT09i6Cr7hVm8lE7UgVVC7Y+kZqVNS/Ik/ZlcVxzB1wsBpJl+ixAtwYeWj33t445fIRE
TM08pFhrHrD1Uxlln93v3MxJMgmGzVqeMf5AJB+bLm911MTNlFFnKrTIdXKg6nldQxIL5a/RSfWP
KZ6vHxuT4ExBM9MYOUYm4X1oHiYVckVxM2qihPKhSAH5pqOdqHW24wX8QeP7Pmy3MoiP4vSnClLK
ftMnzK4YORAGhWrcMFQGh4uoFXJS6UzrpSyRaCTYudFnVbAmkpuo77YGdRIvcMXvedx4/6i42O/B
c86j526WOQGp+sU1sAiFzUU2l2YPfMl1UY9qIjBpJBuJ5fAqHWIkPRhJRmq1IXLwzL/jwMNrzJJn
GMGh7Ort/HYWm3qJcfK3x/F2yl6WQpMmgjHadQDS0rP1l0YErr3R+gASJVEdRE6MCd+pGjNZ2Qs6
D6yzHeHVekLge4xlOyXPdN2McqrK/jwxzdLUm1agoH88xQUD7UVCSqC24DNrClaBipWhk9gGW0kh
2kx3x0mJEiJqoLTMhVm6kUqoCQSInUlEqA5vNf2xxvEn/0ngKTvp7RfhJft2y5a2Fk7pJW+FCZSg
7fpS1zuQSef7GY4vhn+wmORPuH95hIhEaMXCx9PnGaWy52w4F55bdmQDF2OyEvHPP2TrdQHmeNb4
PTAiWwbyAIYssfpRWYVdAUs30zoP7t8ImAOv8MSyH9KNmYY2U2sAIs1XhgAuYui5FoQuzLAceNBQ
eh2DG5IYpb4lv/W6DhGe7kv5KhmkYRveF81j68/5JYb9PTSA74cz39OKLIqgftjlDFr3TpiyC8Ir
9PxoZbGrVpt8Tag4l7QNWvqSoZf0fp23ohO+pca7TdLTSF9Fu8trfAs85rmf1WNC7Uf45dOtge5T
6Po68GuSB+u9lY6XaSkU+SKfCd8FvFH4BiLLKS45I2ImuZ3DL9yGxV5tAgri2hJBP5zjrJLvBUAq
8sd2c9q2YFMeF++/I9P0vaR32DX5Rn40GmZxZhXe4gv09ngyK7mPH6FX7OMiuN2coZVibSGihLUA
k0dUMNT1BjNh4mf/MLNIn6J4Tqf0bUDvVoSG1FP08PKPo3hW7sFu1AjCgp5h13aJ6eTx3XNCytxB
EWVgh+dDrNkoH/j18V0QFLEPk8DBrOoHir76tTI/CxKMHWdwxJLjHLKir11Xp7V21SUid1BBZiJE
DpThCTiSb9pnKM7maynJnjxtERbQsN1B4lCjC8sVFe6G0Budf03F5t+fyog4KCa9VqVhncIuNhn6
NrHCmL9jE2dtpitO0GDCJUbF0aU+kZpfHU/IY+5rMBNMWSxzAMD16af0oOlM43193C9wzGprMDlW
DWqOlEbitDCfKX5CIWtA/cw7w9u/DIhVLkAb/AxDBzPWoqcJzlbyzRUJtSjNZy2Aqo7RslVESzdw
WjBXrGkRxKMgqYwQ9JpfdKsUdVO7lF2YKZ0ryYiWAzdFK0aPAxlGdPA0+xp2xDl97I5gaph4Gqcz
ReaHZfTMAkJ5KJkCRjZIlRHRLzYs0/JtjtADhzthUtxcyx0RKwKI9H+2M/QvoX6TcrOsaMqyBdSn
bQFD7qzU/uHz4LLo/yD17ZNdBu7FwCCP0lbvIeES5ic2BwWdWedaQCqx1D2k8KMLhDmDqoZxH4ix
OBlffx/Pi48A51CrLcCLYd+kzVE8d5sZjWgC1hB5ltWx3DtqgCZa4H9KwBGLhxOBXmXvcaO6lxLu
hEpGIXMmz/y//7Dum5r9LW4jTR4BhGq79DwTq6gvAb3Y1pXleSZyEZmmdJDs4LB88oGoASGjxu6Z
wQcszmF3z6aICLX7zdNziCcLWE86PfzO+4qurlwB7QbtzbhQRICOD72JVWH0FdHLn2ob3UZ/2nzf
8UnHEjCI7WOJJPn57yVJ2jXYhTw4H9wLalO/Baaq/Rp/T1cI0msn69XqB1uhD5TVf4F4V9nNjhrM
N+OGMecNpMdof0wfoDaqxbGOvUfWSzHbjtI8tIP2JPv/6IQ5pVvuiAAIVS1fswly/QR1mf8hiP1Q
cIyNR7pySAGvTRlZfbC650j6HLIv1SfAFQDc6+wG7EPal7wk10kxE4wGMJElf0f84e8RZNY6PsT1
kUogXhyfP6qzZAj+nrCHeD2zeM5T/ae7nWvkax2jncQQ0tJ4iMVlgySH0FaovpdY67xfjxG9WCe3
y3am4GJYRAotOZCDaNaPafhrwZG0lDjJ+J/GzE8AGXcaKiz8oBvj/usV4EjAqv6mechSPR3EY4is
3iGUotuRz36nr9QKkXqcr0u3UazeigIE3Abr4W+tCUeDOp9D2A/hpxbEclGdvonYsSrFDp33Kto/
cGwrWlwXkXTzDbMDU6ntyXjhSOB9PYW1dT4aVQKt6GTC5h3XFiDyuTbvSBZjAVauNCRvNWYW8mnh
ollcvLJpLYAntFgb46Kqw0xoL2gseefePyBOclcPpLLipkJgUG3/UGD2Trhl2ad0KQ9mvXN94ioz
RMx8YQ24akMMyARW1hU0Xe4D8Y1d3OxrG1pLwO+Qh5BqiJZypuVus1MPsdAOa8zZ/PQKpYy7x1pY
jXK4Uhvtd89puGsWbPUNQy+h49JVMTQXogdV+835e++TjgLZi/mcZYXDl/ib+FV4Rb9H9GFbd8cb
zv6mlHJUmOp9rFrIKP171yoMpgCFwuEo1rVJsjYGV4ZETjC3kRDLREJackV2HxOPKY3bODTiC7Sw
S6MVWFJNgFndFThfV3p1FXN/OYbGXUT63tck0tqP9JHI0X8+6rsrZJNfiO4NbOBtCO7/MIrpfoxc
H3ZeoJKqORmFP+cCnZ7gsbtYnIxmg11UpC5d9iMJTuKJlf7+s1T+X+5ntqh8Z7PmhJ8go+ZEQxhG
qlov0Fx1BJjoT+31vO6Z5oUvKQSrNDtGT0hjQ8RuTz24YsleZYsuOYbLOaRgBrCOel8lOuR1/9z6
yF3i7x68xAt9ukwUQ7rDWYZ8JhtetQTDV9iGEVGGkF1w/utZMIAugCZGvdr2bHlT1f/Fczn7AZkr
dU2wGkdcbr5UV3jsKREEr1ranhEQdliccc7EDxOk6I87RRTvbYOG8PjaZuRTiwFreCbO87pU7ef9
tMFBduQLhI4iVCcoJaSD5iLGZmEmujanwmvqQW6YyNUPeGsdf0Gh/kwotNHO8OhcyYGDdWeXfa6N
xTK4rv6xShtFKl0Vd9p5Fhm0wFOt5dm91MfQJBmAIk6AbSQJHG238si1+HKaFGPwoGS75/+qwswn
RL+mgREnpzrI3DYOsVl+ZyfbIhRJqqF47/384xYR36Dv+tXuqjt/iBtkkRPI4gzcNU97y5jadFUt
qWYGcRFhHQV2LPlPIipD22Dr9tH60zegPM/AVGC3OXsjUF33YsZQm/4g/GWjTiODfv7dXPQetA1z
6FJFvd4CDlPLYJj2Z4aurkqoLaQbDs32kCAC2uw9RBqltGVKChOJPY0J8g0u76qdd80fhQQYnp6i
6VJwXLrp2CWxtN+zcrojKwLunFfaMhzQVs4RJmlmBb5EkwQ3gfIHfKab+PYJxJKTo+SC7kZpc/fb
XKaL9cxxOlTha/lh3C7DuBM/FpoEe23jrgu6mbKaLZATDnKUiS3j9Bp3Dwccino0aOcRcM8Xyx0i
bXgQP9R5pnvoSZlKdwl/62Du9DEqCpUsORdyjJxJwD5VfvU7GzU/fcFWsMvLEgfEyar7BVbmLgpk
cYDUqDIM/0nsEZSiQQOTVDIktkWAyXswt+mbRKN/2pG65weLk63VuJaivqP/kw8BWkZWNcDvbDoT
IMYBQ5slMaU7wWmiQywwj6gjSRiJDOBe9Exyjr+7CJSUdSiRmQgLytbKfQnTKS9pNsaZodlarwcv
Te7oHLrXCHBEohzDS1DlGu6vlO4t3ugRwHxNpaPMR+Lo0RZH8xVQXSFN2yWcJe2F3VDdd3PleSeZ
ib0EHQJPGE3la2A64uhhJeCdFpmZdwimjssUTdyWkWGmi2zzqLG2+kayjyBAqTuK3dv3VSd8dOwy
kdoB1WUcoticlZeJ+2EqVPbexQ9LdK0HERmJOCO+AbatO7HJbJKxstHNHDoYcf5kheEhybQtco3j
3LIVoW+E3Xl/SzgTTjWB758MOhpgyF4XiNwKPfg/WPxKM2PZ6a3tTA+o8Isqk3OfXdt+xyDG0MTp
wvvsh/9p+EQ4H2AgPYEIhrCP7JqNAsf+utvBpCUK9pb8vSYRHBt5P4D8DnfQ+dmLdBGlY/ZjK6Cm
FN0p55HcRvSj08I7WlgqP2TJdWDBHGT1IT1edOSQ16zx/xYVBNFYpFhC5jBzYaqbLdPbjrsloLMF
a0N36Z+aoBW5kZCbcbpR0ns61ADT23af2jivYi0c3JSeJOn4f9NkdaT6jaP0yg8SUqeWLcFkwts0
lKWbqzCIDVRAcjrptoCJ2b04bATIrLia4kPwb9QBEx+wmox2H0IZxDQBgiEnGNP0hwa1hLo4jsOx
OH59Cq64fEMFSHiIoWanQvZctmbd8mrycQaNeAwHD1Cmb1xKjRAFSaiJR2+UCPsOAZseI4Mc3MZo
uPkfQII2s4JZWBz1wwruVJJPM6zSgwARvvhziIZv6S6GYBFOABfYmmSHw1Yu8n0t5TBghNVxdSPU
vf48eoU16CYbMudErASnPPF0/1KnAaiPRtmtGWDlyrGcyjVR7+VvwtlKY838f5CxpaDODVJIMWQp
yL84i8sg+l3kfSYLK3jgxlxU6aRASUWxsdkhllibR3GaNImJuZ3d1kGDMNsR942PpspgzpagfQS4
sNmA9XrjAYIMzZFztKiiBRqBAC3qx9g2y3KJk631453PyoVdaUkn3UD8Wws0Fcig9eXjZTDuxTiZ
XXpv2YLQdNy0QGcuUHFjg5qCWRD9pXKBWgCZl3qD3fIZAzKhIof1Qc/kxYDjGHwJzXp1mZKaNfwe
3iYnLq8FMS7atW62JlQz36850mn0a/anK2CEM8PJvxHwt4POXWye5z8atyxPUvnE+dEXFD5n2y+J
jmW0NfjDKzzjeZRWxODpIrGWna0rkt1AD1oCoL9Fo9qkjj1s5hxKuGqUHeXUNQsDM2fZen9IKyym
J3pIGNwFclpSu8BpQ5iNeqqeArFu80C7sqODJu5MFKwcv/bsJHyOjtywwSzE2dt5Wn+2zutyNYtL
d4la3jOwxnyIHJ4yizMZ18dkDf60z+IWAZ6fXTyUJOxyp/zKjpyZtsCiULuOOPNAy6gtIhsEvC+R
kLeTvuVmu+jdUOTiBgFz7fDkvtl43erV8T3o8UQYWF4n2FNRkrIl0oAVE3AK2/9eTtbq5Xv8uc0a
ZIC+qbaeAmP6a7MBEqDcN5Jq/ebjYM7uSPliDFRbpVUgH5EhrNioCLoMO8tZxJxdi8YZa5MxTnY+
ZL1vDS0qUbTNkrIdr77JHhScFA4QTUok5B6Zl7tDEqWjobBfvzbThg8iLevFIdCty00I7qsVRsn8
afu9eshPmRDN6+jqJRDhfvmFsDFIlEXld6qUJFvAigx1+dAMQ3BA+AgnpHyZY/woFbgbZFvj0fEP
Tdmxz0ySToU1S9+SfXtriQzdrBvkPhQw3jwrrmpO8DlR77/nBwng2o9d3SPkE+kZM1JFLSFWhxW6
S2Lzt4pjbSZAA3x4nvcQKm/C8O/NAh7cX2d2D0DXvDsQ3u1JsEBZdtV1FfykN4O6lgggvk1ZFU8u
5sH2EbipWtzypy58e0VDW0Q2Xu92lQFH+akBeIQWj49NsQ3RSa3UHfFtbDUMvejUYZKbVsI7vQVP
+6TgxqRynMoC5nsc9pk+UfZ1NmOseSylHQCWtMgz/DpcHkz6vV2UEFcgVgJVAoE71Wh2dxQ6ps2x
sOGySndsgkYY9xNbRMGe/C7/UMUtS0PZmEUTORYgp+++0VW6lrIG6aI3CGFBxvzKYr+0H/wPCs9E
3hqsSOggxHDjpbjCzcTC6kVrjNwnomq5msAwn4t8h1wtWmual4RD04uEe9gX0/ltBJrOKGJCflwC
pjXuAsB51sNtLAYw8Vu7PSy76Q5jWF3pWSVGUsV79ui2PXhse+7HLTEM7FEBmpkXylr5CsJu/Iq0
E461f0A4FnZKK4v0y+ZZIb18xwE+CSS+VO7gsazZi/MIgM5wszs2Gd8IOf9XfN0nrvc3H3Zeq10S
XGUJvKFOuMq2Vc9ZvHQhua+U4jPlxOmBVo+xiKTJBl5RX1DaZQ0hJ/8ZmiITRKwZ9s0+H2sG8iwJ
7FeTGcsRxjTLSoIkpbMOq/+/Vxuczj1OCYa2CLv0BC/OpFtnhyPdkLBlkTaejP/QBA43EfieZABu
rzdBIV0IqJmmqno3KceITAsnQ1QEx+heXzVvoXJu/7qg7nYgC4rXkHA3dgKAUR+Yugl33CqEqVtb
BZj2bp5dYiUVzvM6cs5Gp6NdBbud0Hh/Y8xvF3tWTV8V2AvJ1el6E6fe/A3LpUOu4CqvjNqou512
+7SCikjTahhV+XliOihNGnjIgSkhISDcLSXYDCJV/U+XmGVq9jDAUyuvHPFLRZnrGjfr0WxLo6VI
Yql1xSZALnNF3WEjgXdOxiP9sBN4JVFehsBNGhClmhkxm+eghW2FwrNRGmoL+MkqPysymn0K+vsV
kA6KwPaz1XvdyS+/IV9g65Vc2edDYOreWQbFN/lh8EpXH7XzoQNVIneKy0JdyFCvQTn6KaAsiPVX
CgV2ezXsFlUwz6yPZBqscKKN2Sjm1lP/7Lxk1iuCrI6lNyfVbPoiiBIUgemHlUoMAVhAze5EVYFH
bedNzoXAH2KhGRnWQdAz16oJIDIj5IL1IfcfyaHw8zSPiKcpV3Id5n/bNjRUzP1qkVwnLB8YV7Yk
mI7mbFMcpHY3ynwSezXSFxCf0CD1T7or/UfpieDwNdry7FwvQmerL+BRDy0a40TwFWWd1xGxNK5H
6VVl4p4sUorC6BlT43h/ri++6Bp51g46BALuM6VXABnhCP68UaxB6/AC57wzbxrxW/890J//2Z7D
3HqLanDl2TApgkgSn7uOpTm0yJeRwSNqf4SgqIMWVaROLLyAf2D+YKAsm/M1R9YklOGnTSgYqCDS
LznmAjzBsL33w+sm/KL64xPYiEOaU1kDAqCuCe5yUmhEfBPKWv2nTi9BeFHyNUeJ6CtASNLQr/zi
S9JHM5VHoBDJiZuHG55Ct21spl5Jbowos+OjVi8vF/zuq+nl/p2Rvw7m6T3/bhqs39UT2HPy12+Y
IgJnMs/cJypENH7GGm5aocfzGihYJakViNlg3yIKwjBMAHcklXBkiyfQszeM3PYSw38tTR4KlUBX
ph+v0pvQHUSyUSvtMja6mGKJWsYdKUK6elZiJRNKGI03VgIpFxzWFXHlDOIH0jh9oDBTbJ+ZhMwq
dJHBa66+W0fPzVwx+cGwO7jlDyt1RGdmlXaM61RmvgILavAopNiJldiKihQWmbRSI7Xgu9EtuYPs
niUuBl09yBDhX+PEBQfQjApDqmzqwNLg8GtB5OdMxGcAhZvaYB4rCXYL84cpQxOxK66i4OqoMiB/
Nst9ukW3dg2CWmqqaxDq7+E4K3ey9zCbBQ4wd0xkHE6f9a1tsWGpCPlqH/gWLxZq0aQ7d1sxlJvP
t6VnRBcBvYZVPh3CALYa0nuh6oDY2viaWu/IkjFF+BUpOZYmzxNdUtoxreJ+7COuU+KqhT+3AxPg
aLP+FzjV5gnQI6QsoOkw/hdiGiPBSykF9m6NlW5PD/Z+VSeDhiCKrXUS0DQ9axfCgD6ppI0EZe1O
oJ0NUshrPmjpC+akKIpbureIIDsDrd/3VBmjbcF77UIkZEgcT4xTH1DYth635WOSNBda4OXVQIOx
QEaZVhDH4myZS8OLOJjPdFwxou789XyOEhglaYdEvKg0vTVKUC4xBbAYpJwDk+kTS6iukCs89PYr
gCtxsla09tv/UY00wYf85vA7y2DOdtuSxdwPVvmzVdGUrgbMuW/HNYIwsYV8WaTIuY/dRd0TvX12
StdDTfWL4TdnQJgziMvud4/3x5bkGxSpwABVNK3Iy67w5antiCp2Nn3Y+Vbtw/wssQqipH6+zDGc
VTAptkkaAuAt9XFPRDAoFV+sC7PGWaVCQ6MM/BBHW6v08ntq4BF8FSq/6xDzwst5G1rFXquWsCam
gjz1kcVorK0spwzyI/jL/rATJjwqFyEUvqNSL2aGVKVNaTlJS4zHYJEo7dkAGmTmxcjwispbDN7Y
wfWY8FPA5JT/vDFhzDxiVhfuB52v4ZAW9uF2Ks/oHHa8YgqfC92vnWBgRBZS1gf8u8sceosgInxn
PK77mmvoy/XoUq8Mfkv1yx6z+S4sLQHQhrbf9D3OmgpfTMMQSiqItZ/qfG9GVWaTarIsuYERZIZ1
dU78J16ts82OBK56rzjBDFsVAkmcG0gsKTm7wQPL3QwRAY+MYSUI1zYqSpSkiHqIHFGAibOqKQwD
ciwLCT7HJFk4G3GUU4NP9cjvWGFoGDguOaMyjRVTKAB4vKAEuucCl27QAU9/jnQNKeAWP2S+7usZ
KQO0+18FoqLk6NIUBC7yq+Q6YbQVavH1RrufXookGt6HlN4H6/91mPKw2QaoONmcWbjejUFHKiNc
zOkhejJTE0jC/jPgiwKq1rBq9p3ztp0Q5sss1BXtqY7tZ32lq1GMq8tR4K6d3XNolzzXfwPszzhj
+tuOQvPoDQQ4oeuIRKSxt2QzjgxiurHgsyp9eFslzwAhMVhj60J8ygpRj25KsTW/e/l47xSlZQgA
Mwe5mgeRmvWNOJlaHKnupprcTu0YEz+ULWviJjaKBFdHYMCAkoXLOILvnNJQFo8I5Y+XGlXdQwaD
MHM7an4kro3f7+WX9Jtawf9FWaI64pCS9H8P87tE2fA9v3r5nEarVqlYokqKtAQ1+JSEFZSX9puS
8f4bbiWTX92ouxPYZlmSWF08hFs53X51GpBXw303fyb/CES+iI2jgaHzmDDW0UNkCPDhn+9w+H1U
FkvJhaGdFMK2o/44wa2t86XfILbCXIDRRNQcTSxy4upoTiSJ+de0uZpONNU7xYHWAUwauDTIQHi1
XWFa/oC37DGa8mFJfrfP7x5ZOpvs1+UhQzRYu+CYNPEjdnfkNtpHkdNmzUI1y5NZ0zpKqOyoSD7y
wgxwjJhGKyYUDu8lFrs/8K9ztOQXM0ZO0bQoepl6eLQ+3+z/UEVEBhFAA+INSQOAh/pkrOGBRNzn
FLwJW8SFyeGxKG4qEk7ak1HNmobVJZiA122QkSxde95jGbq6hq0bYuCEk9ZaNUv8h3XSA3VfJyBu
t59DambPY6+O9oD8amMUASzBQCrD2aBHrrgvy3ctUEeY66evu1CJgj7T3VGZo5qlFbrN5mf8ycEb
n3cTa2Eu/ez0xRvlDAQeTVdXvolZvkGL8LN2kHvVahpyqo65fyrjO5+KHVyelT73k3d0XwnLkc1b
NQl9NtwraNqNslVLeELAwojIkFqYbt3h6cAWAUkysRtaVZuBIbDCV2bZiEZPdciUpRG+t74c7HaA
GN/0bdR6xrwgHDCDhWb58Vp5afeSNL5L0kvGKbIV0xUbsGSgl2gyXNb4hybazc1IO4klNBD4H4v2
IHmA4CfL/3/ZZiqwo7hyionjYbo+FXaDXbydcesS/+l83MEc42GR35vrLrjAum1KWzfFsRT1tAdC
JKUa3SqI3C7FNEd32l9zXllHB0QG90qPlquQujSilzUS37hwq6H15Fg+NXtVmLRma+fQf8qc2x2i
xWzqSMy9LJ6s7d/Na05KaumgNAIieCm0YqLgByubla20Fitp1xyRDjOk+ETvZN5KZs/rwUX5Zj4V
W6H7Oq1jc24VinBzd07Kne6oyBy9NUVru4Wm5j2ASq9CMaYDrup0FSqXQz0zZC+cKrwmbSc6KAsr
BEkkYlZtdgo967TBhrQC/Km/+6e8C2zsowWpo1ViS3oO8pf37rvHnaV0WzwANn8OYo1MT9J87zRK
mtzVgizsTKD+LZLADsfMZCvCy6w8R/Fanjc8irN/OkBlDGN+7Q0AeFCvu1G8GO9hfKZyq4Ixxbk8
EwSAMpo1smF1XfB86v1mlxTkHQSRXsT5ks6ktuN+t013dxzJchuQ6RgoM/7tZSj3V+ELHFOmGKBZ
LGyQ/zNAC92nADIrU0zHm9bSBwaJQKcAEDqAczg+S9NES+DjCYl0zX5sqAdSslX/Z/vy4QXpRyTv
vceIPKEvDw0/kvuZk8rAs5PkBVbb1FveLxOlepKAYeRx6egikNvOo3J508vZO32wf1P0g3oTz2KJ
b+iqz7LABGty59NCEEmvQjZKbyzTlmCUzuqvEeSlL3bNpyw1v21uWBewIYt1TJyWRSXHhVb83UXN
NIsepxcfP5d1c24mpS2Jld111vyazeT/+lL992bbtUq76UnNXBvI9oSLYQ3iZxfw/o8zshIjC452
MGNF4Oj/ycvMdlYG3oBLHJTj+YMo5RkYPupahWdeVewJrgGbdZwHuR14dYxSMLSnvuWuSDGGZwxy
IGQNRacmk2oKdLWWUqKnkIDGqAyZqXJcWBgOgNfz1Z+bk4XGJ511D9GaJroPlic+phLj1YfMgmOT
ayIsq6rmOVXGH/L0tTk4b5Xf1RP6fiAY2A3peIR/V+fRCUYDJr7z+rWIBcRz/xPNyT4s8bT4QQIQ
9Op4EZQ8I8W5/TcYdTlYEUU5zcKbhHlRjKPlK0h5rKDqSygAstnUFGXZWXcjra2INYpPv8V3/xPK
ZyJKxdbKl9elfO7tXMG9ZgKK/OzBSj75XkESF6rLqQcOzPZBqIYvv0sBKMEMh0bbjuX/EsRxPHb0
5W6ECVXPBjcDHPjmFa/DKc8/nE7ylUsXCp6extChEM+t9H31uJCguwIBBioFE8NKHUtjPPrt21tW
xFtnB3KnaD4vnD48Mi3xvLP3Jvtcj0AVn5GXh/JgxEA3G18nSl8lO523AWNpnGFea3mIcqDrFOcy
bwB00VCEqHQ5MQPM6y0IyNR+/7k3q4X5qBTlSe+25LBxnl/xjjonuW6d61fYOpV9gCeNR6IM96+X
mOelpoD0ipptZLMP9RO6cnQbU8V+EXAMSl2cvRByUGEiSOtvQDNpHC+cvyS2PCc4+It09dW2rsQy
we0l47LTkkxw038I5MoeovMYk8VprXiwmaaWQBbUIyvMP7Wcr6e3djyOMb5HsOxURFf/hk5V/+bl
Vey9QKMz8tiPRd/W6emGwk8eWmlTBLSvxNUcSEs+HdWe7HBGdbN2FYMll+c2n5BTNwpPzDGyHvjH
8cLtsfqbpenq78zsicgY/22uM6yWvYO9pVPjFC7UAGtBAVl+thROLGu5CdgWgvk207v25TqHOn54
R/uThl+dLxpf9K1pNqJtC7ZPhMz3xxdCr4p3/uiqc3GY+PrH50A7nvSy2u38zym4lLX554jlqpSt
1Ejfw3in5JSd6a/dDolYeUQuLNVDZYwf0jNnaS422xshEV4ay9tOx90e0eblJqJ6TQO3HTuk7UjC
8GMaMPPVVR+d37Weesp+vCSSDN33L2R2QmEWYXRWqIwxkwWDGOHbgGZ+3pJowOYk7u2d+62malvB
4bG79ELRc5gKEAJggFwmZHHzUz9vqsauS9v+tJagPA/g0zwEr4x8Znx3i5QfQEtlIloQyEIt1dFQ
0erzCpcLulr0LN98/gVqwKHRTEKnwoLFtVpGm2+s2/g74Pt1rOjrzEbPx6abiRCYKpo4my6obzSI
ZNbm+p08h6TiTJPg3P0R9+SZqEX09Un3UmPTxsUTPLRXHV2I6apBj8/vv5Zg4huMVRnZ5J3XXl0q
vCffEJuCYy1SIJZTIJXEJiEMcu2FFLHF1pGZs3WZBE106fJzfeB/GnHilLGSiN5jYr1+8JbNhTP3
aWfDyiUWEXrLrqxqWXM1a9sOsG1K7JYzSkS7NVAxnYjaoHwW32wtPSmrXKClJnmngHBjSnIuIpBq
u44FlGNja9lijjhWN6eUwDGZ+tUVtf4ruWiuOt4boi8IGXfWW7lbo/14XbYjuZ+nO6s1FDPCsNf2
HBhU55CsPu+LzGUsZktX8BMnisK5F7tEMyIKZfs3+vJdhIAhjKBYAXYdnpwpcxYkoBW7tsJIHZf+
FHpzAFOW3zYaWHP6/wagmZQEPeNogZeEEjuUVFs/Tnggcc6pRr6KpBFFSe7ZlEK2NLl17jm43rdB
oadXLsuDCQ5h/+uaDlelSqdXMEp2sUv5yyvdj84jhknHGEM97fpCFhg5zRl7N+GuuiSv+24fH2Vd
1D/3hrCGx3Vf+G5GQywFgbzKm8ARxot37cpbQ+4UmMQxLKruq/60PKSMmCc1qhNYnre05UCR8lHr
OY3fdZHpXWwn7lm6vC6T/tMI0gRKK/7rTE8beA/R8OoWvrvpDE9mYe67pCJZaEvtTzkj+KBXLKSG
6UF+a1LmBrtorB0Zn5dgfgicv6UHO5jHY0M4eyM5LcIS4FOuEv8EVR8vEbN0wNe93wJZ9gXRSV6u
0UHrimJICC9cERTOwqP74hQgqqtnztPwg8bgcpr5bWv/aj+RuxGulgfmu7kSwZWnvmcMihu6i0Qs
jNdkWgC5YUk5PSpKugmnBjgpHNZpFaajwt9kJd0Kx0ZmgkeGaTyaZahqm3P8deeJ8EA7hfGUZorp
U+7ZKlVHpuLOhW9sRSmJnDxM2LIko+MrFQoC1uZNC23FX+Mncn2emwH6tvlB5ZRaLPahpKoxn+Bq
tNHZUf59xHQ5xfM3ObkZ5E3AoD+bn5jXcGQNDMHq9MxnLYdgrG+62rcHtDdrI739km0FjPFv0/Gu
/LKXgU+Tr7TVjQD9swyKDKUlfKnK14QinVXCbrW8WkfuY5WlNSGGQXTViMyobHuNRaPXl/AxOZ7b
Kfsjyr/6dOZ8PEjxER2rJzt+wFitiSJWHglmyX/AVXICuGACzmRr+AuNDoxAv+7RVMm0Aq06JNo/
Q5AcUtg8jsvMRjG1IMezHWO/d7l8XyDQbSfeSrtDF6is9Yt9HSGqvfGSGnUV8FTE9idhdN3o88xd
6HzGiQRn02B4adkpUdxQQFeJ8Pmx+vAlhLJdudubd6vqHOcnoxLaeotckIbMeEsSfd0iAA9XFgXo
VrwSFHCGcAfBhUFBCyxr7LXCrGQOjJczF/a603XqwHBjek3vE8c6PfKkOtYdPAV9d1ScgX7VIzrD
cmyvxAP46P3O8l9PDSuTjpe2gJ6NvzWVBCn5BLK16AB27lMHTZxJt85fA4y0yam6LxUkrWZMF/HK
nxQQlbviZKNKRsSlXs4LMJrOIepO6rw9xjBZ45/RBZeB+/MR0Co/PrQ+/BPcvzi33FNci3enR2io
I5ojW4+1FCxP8CMqhsoqrm9rth5zSfDPmrgeesFHuv+Wgz7gSJe3RnIE/i3oAxRWPY7SfzvjEhZs
gN/BcAzXLh9swYs7epdclLNytnhb14UGAg5+URAqL0dzsAVWMZWu5v3odWz9zqwS+I0NtXEvWhlp
w1zkyll49HjEw1WoKPMjsT2JFdxdal5uGj76NZCwiO0KaWPPVyavy1VjqTW5GrMQpbr3ZLEnLOx+
6JWIp1R4qowRIJ1KeWzpW9dLqFAdAQCh+SMCtDmo3+vcwRNfdHmAbR4A+VOyjyGdf+Ard7S93wG6
AoLpU8gjaXqShjQP7/knrvrBNO5K0buFplquE1NgFTRyPojDn/dXYKRcapfhGs7DwdejM+8RvpLu
/BknaOU7fzuPYY63DEsSrDfTAWxjUeQeczUazwPRl+/y5SmPY3hJs+Z4RYiG+kk9k2J8T9f0DMlh
htmEeBbf74K1RR2XerpwnV6LVoyZxCpF8vs7HtT4E7sxG1wUNbAL/AhgFhEKojvKcTVHef2C5DzZ
OTgK7lUG1OJYb/QE2BizShbTzduNCWVacWHTknp18U+JfBmehftzn4ryX4Z/jMl0S1hBkZSNJWJm
rGsvDQuopMtzdu5H41iF98Pm6BEbZF6oIkVhsiZCTGmGpSo1VyaGofMNlXIPBqdKh9sO5H7NbjKP
cYQ5kAQ5EKq/tHcWPwJLt8LDrlIF22bcTZT4JiJ/rLZZKy0x/Ryz6vkWsgPDXCscsz5LhUdh0UXq
dX5ciAh5Zcn577MNuHmt+nenV0gspO1JWxhknD/DJilBbnHGIVLjhiGFac+A+93X7Xl2cLOaEf6V
dRSEMHyWeZmQ0QKvK8NPVNEx5D9Vl4YhX8fg0ZN/Vw4ucwth39i3OvpEg3PE1vAmcFhFlkYzbvnz
jKNMWwkwvo/H9xuguYlBrowuSQeyUadYB3DGGahGlIbeDDcBtgUKoq54bGQtYI+rKMKU9CrDVDM1
ELu0MbHVMM6X9kokPyjuDmEB0x5qmwG1TcZhpLv35IV4QPRjJeEvIRlabrimxioF4+7FAOxVkgBp
j9c+dXVmeIQ9UF7sCU77tj2ew8mhkIm9S+scTw+ydgCJ8gjR9CnU66WTnVNSA49aZwcGVdKba2ii
5i25vI0g65sRIqbMhr1TH8jZUsBRdouYpiBrM1mGp23xgGdq3dLzyCY6DGqw0NhA4RKDJ/dS/Uxk
AAqRqnK3iGP/a/x0Xujf05O5dDUBEy3thOZ758w54npk3A5ylzJ4hjzStifV4d3A4d8kr5VXZd3t
bLO8PfiL28wv7AofxSEPAA5atpta+6VNqQ9XOVVqHlgJebiDCzwxm6/HWqh6PSO37qJMV3wjnOPr
2A7j3krbo/ZEikfjmUnjA22FJWbb63wbKPiEr8qn0/lGPQRlhco2gIl2I1VoY71MoFxKA5KZBdjt
XqQ531JCHr6c6cTwpGzMLCPQZGjdVHCcSv8cDa968MUfbxkX7OiGKL8nHpQJH1I/3QicZOsYBbOk
v0Q9X/cF5lzqGB7ZtYS0zPvdjDy23GlHad0JNJpwGoM+ion1Sz3ZgwsCkGngcWvEQ6nZn2rGy06t
uXLpcNhnxaOmq9/5qN3RDIiOHB3UbC507wENlKuH4l/hMdBpuGaiZ05wcbhG24526z0fhKTYR9o9
whAFVAMAfDv/MIC8tSMCi1dMLu/K+mZDTsddb91L9tNgddHIcscCJ7BA+RBnoiVZ8morbaOBo5V0
9NxEvEcOvcflht9boCUInbB47gnKBZ8OfRCiRMnRsSaNgO6t0ev/UuCxOf1l0+b+9KbgNkE/I5xp
KjWed5XABgeSQYV4rWCSF83tly150iQ4AuiHmX5d6yUVia8eqFuwKvj8yTh7wWP9yKKwXfHiXUdN
n33RCXJHoA63wW35PvoMm0pzvYnHZTAfpgxy9JkYYpStfYDWwH60meSV7npfJ93wEBaR611mhJu3
ZDsQdtRYUCU+btIWI9Lanjq8jHT+VbcuzRZHTAMEenYCd3A4jP9/E/qyf2OIkVgMWhzmBuyS5BDp
xPnuJo0nNTXvex98LXKMO0/K2nPBMdojclgqKbUhpxml9fpz2FRrphFDfVruH905XXOLyI4ejdlg
Gr3hAAGSg4Iywc39KxLx+e78t+Yozl/BEHHiPB518T3g//P5zu1V3vWcHP1cfWGfn7hxf64az9M9
AS6kEouBihGwz+HeU7litQ+FWefbS5tCscy79mlEgYGNHl/nv6F8YuW+k8JK9sGc65ORs6viFlxR
A1jgMW5cE1FYGXngwDNT2OVOX+/aH2WAv+WXc0HpKDP1Eu92KHOb00jg5gisjYynQtWFaG27LZgU
hDBPHel37RIQ5NOUXdpOknHOhltLNlqnt+lT37xgS2C0YjL0g+bwvgoTfALz6QYEC+/Ab/cV1BQw
yF4kZE7A/ScQ0xS95srRzhADgCHyP2Ahj00Gd/ZMMpjfTC7YhfqmmgvvTPgTI8vHm42yGR7TePEq
AOa2toJY/EPdgBiNIBgWucKXPqjka6YblrWvPacA+/8Q8gNz/cuG2MZikaymREdGzRV3BSAiqujJ
G6Botp9/Y8BkTGBEbvPnG/KIgnCSlrXpixLFonwF7BPTJKaIqZWLxTYO82v1XrVkbAF9INlyqWvH
4Bur1WA28AwcDTA5ghbMU4loYkyBd5qZ3ZR4QgcVZVO7TNvyVicaiVgdfBvlVbfqHhiUYY1Jo7mw
rXATgmBh35XNyCETVjKjPg3vhIa4sWtGgIQ3IYisJCiACP/AmLAADqglLksPvDjc4tTPvAFUklI1
/3fjIxuAp8oL+4CGVLK/pe8puq6OjOfmMy6tpvalBLbN4RQlFBZ0zj9o5jRhr3Y76z3LEZwSg/61
Y21nnYv9Pb1rZGaoS1/XnQJRqo3cHj3UILOQOAbgzQrMD7E0UaypU69eJejB+tckQoyn46kFwLph
QOIo/Sc3TGUPM9cgxgwsXXCgZAmADNUJUdEvVJr9T8ySMBmbiwBxZiiInRbp/6Rbvow0HAzN07u/
0WLeL5KtVc9BUF6tEm72OwOzUma5FIzYseaG2SvtifgAptydyWH46LpXR8tXsOqwnDoGnR6Pmoi+
JKuKjLW9rMPTNBSA5ujoVo1sbbZ6r0veaLPKh8bJXPiiZFxj5pq/rXvkfkdHuqxVW2WQ8c6AYexZ
GMfmrLz0zyV35RO7kF536GDbIiJKjFIOM+swLUuhZuTAYriTwWt4jaLe5pjvf6gxZeZcmH93zlku
9BffC6bZi7yVPDHFUcqaTSK3MxaRJkQpA7NO5L5rzgUo5PhJHA7Q/y7HYyLkZ8iYv9nJN8aNcBFF
1poriS/ur/+G0TNORJvAAR8vt3p23/x0NJSQcojODrAm/r+SFsgnT5SbxWSS7xOdL9PHgMVfPAqm
ELu5Bip5I/oWbjvFA90Pj73oCPUxFbEJa/EJmBficPmuaHLXX9nvlWIMyU8sQFWtAxvkj1mIXjyd
rK+2CNIcOdjadNz/stGeCsjyIeyPH3WGeT4QKTwkTyOz7Nfa6lGYT1/ksSS09AHtO5XhH70bph0g
roNiflJ1yrbzH/x427CCQPQUGrWtD15KL10WlUGv0LoGhdPMK52uNkUiTxlmxbNB+mw2xtJ71YoG
yZZc8p4HY1NmlHOeIm7OxXChurKlBO9PcfERaY4vkkSotEDeS92Ce16ZBIu7WvsCqjYEgzJbtiAt
N0OBh3QJAnrSaYnT5co7pk8kgbaBVmRKV/FRsiL8Sioe+GyGnDxT8W+7qPPl+965YtZ7wBLhRbAu
5NHwuO3ksC7gQIZRGYWWXTc4M+zTH1Wn5+j7R6DAuvBG4ffYTwDoCewoR2IlXoD75PavsUQw35yX
8KABcR9JwLYfPL22744F7r2ci1OrYU6N8b/+nLHabzxPUpLoEqIMysQdoa5kwOT6hqm9xr/XhmFS
1L+3jODhw+ch/3ejxz2tempMiXIp3Pk1jKjZ/W4J2eR11+t1GyC4iBHq7IYe/y1jD/u4SUK5I2jT
7TYW4WuU54Y0QcoIvDltbqCwm2mLDim7UvWRseWFdlplCVmSJryhNQHVeqzgKSTbU1exw9HU7hPO
+3sxny2H9PVcHuHAGDV6/jyZEpvI0fSna13j3fTo+R7/5IxcwGRg4JDDqZvQ+wb1HPF83SmJj7Ak
D7egNRqLe8c1852evFvWZnAxEcYD0mzvJBZKMBk4MLr0zUQWDJ1AD1IiGU0ti5RkpK6owYRcf3JG
g2FNHa+3tleoOWapzaKoGbtJthGzqhrLgNOqNNpAnAI+qaM0jbL5hd7p6bjPhIJFIBCbmoV1x9ny
hTEGmZyE1OIMc1WdjlPkrTyKILMZ3SDOMuupasNoazvkcG1P4zcXveDsacWz2s0CFH/sDWo3+yA3
SMtjHRQkoWnNHIMlMNoSGMJxoi0AiDahEjNnpG47AedGeJxUVT/Nw8ytu0AM5HqxSIQgyp2qIQrn
P2PobBzHtpxQekhbfswUkkmkbXboe1nejTginl1tyXEt66KMGwFHcig4UqGex5/bciPRd9EMpH8G
uulxhntMQnaL39RVZ+SK1rEZlB7Akjz/K62q4VP8fkC2qomPi5zED/H6+DZ2Zp+4RXnD15hvTdxO
/MQ/JsfwntDVDMqBE2ciPXG29w24S4j2cbC13lBd25sBHFkrhoPcnP8a2sChxCwjELYHw8qlgBHv
wCMxHRKTpEvJtLT/VBoYHBe6wlTGh+7G1hj5B5bxnKNeGHeLUwToi5uwn4Aw9lxJwh9/D3IKmHZg
9by1QvxIxmlMRIx9Bzlkn3JugmRAum35B+mk2f15pESxbt+sDF0NsURzzn4NwQRyP3SL/HDvGwl4
Jzj/7cgy1+ARVe14+aiOzsONgJpsE75uHVyjHIsyZt7sCsWPHD85KFeYo6tKPw3rtMyjFbyK8UvZ
lfnr0mPsMhuJsspjMqKYTjysmctOkXkOrknGalOp4F3o5UpvrRLV5Sk7biIsgTUP/f2e+40eG+1F
Ame0mazKnrKj5doVZTeBU9YaGgZ0hcNaadg9TGa5it26m9tihQY1AHx87MF3V1iFhao/PmcwrLe3
NrwUwEIi8PE0FcdC9RLfzGA46xAnTib/xMfuwHXffTYaBFvEuxZyfdyOVfwiV8zhxfj15DSKLdeQ
p/qZEoZ66NgD07w46KBro+YvlpQ9qtHeKAAtD+fn/EKQ+5+Bb2lMzGcnCON/Bk6hJtby2LWkRVel
4AMCZvsE8c02SPRTsomiWTLTM6bwW9NSyvuGEo08bi3coIRb90/kHxHZbgTuZsDBng6bCOJunVCA
5P30uZ8pxtXpzjur+tXz8kSZqNsQikYCXk4VgCa1FRpQ8yzyPAdprjORYdN6KuSN8Fye7Z5FVDiU
jtEj8o1sDpwlNYtlom2ZWhk/DffcNLengTRYNFI6o5yUjF7rTmdMIKaKIFxfG55cRQb/+xSWL0WD
H4328vu93APViTrbvSPcFM0fHqx0NwIVuon6t4wF5yte5sa51CvyYpEJjSNs7Xsgik0CzBnM+5ax
qXkdk52nLdP2BTLUL0u3ZBl3wysu4KR4J1dS5x+WfRDLOWkhswVwTu5woceT1+yhEI09QQS8S5KO
Tcu6eyVU9ZQfXqcETBSEGAWglowrR2Iuzz8oJ7z5LAW9CUxVFsznTf5WhujOah33RIrZ2sNGvM8p
aRTaGtZK+jyHgrLpUuBWtOJ9D5o8Kj3OsF02BLp1kS8XPwrGmLxJ6Khx6kot6D/qc2Gsjn9TrZ94
VHPOsdzLI0QSntnh6d4oNqHP2S/7Pb+WEnoYMeejCGfpQzFeasHSLzGHI4DFvWSlZK3JLZcTWG1s
V21IHyz3mbwt2+AFfdFXSHeRMOXodA3LFvD8tzbl56mm3AGQjOSdFUVTaIzgHzSaLOU9V2Nwz1aS
4d1/qLYcJY7SevK9/0GF18gogMxtE0rR1xynJCcNa/OKhPokzwBvi4RbXbHOXtAumb/BW/mRJ2oS
s4V/Ypn6Tyfjn4sKH2w1x+hTbe9rcBvA8ozgvAlM+7kZaxr9tGykl94rBiYsPmmhwJ77ZX1DIMEI
oqyPO2atrMGFWyaw9lg0UsYAeyauaxpLed6JcHhbdfrMulSSHlBSgTs0lMu9MJeX48ZyP9hdYlDa
mwOlzxyMx9B8C4csxo+a24o1QeCtjGbyFiNeDPhJ34QT8/qTD/igq2x2s5i0Revb0W+cdCd+AZBh
JhO2CGq3pHk/XLomFuC0ybQVgxkBGIRXi7v1ilCb58E97dyfeY1ip3/7Y0OlYtmef30SMUNiwvnn
5NU8Ol9CZ56eEK7mdT3BTpXUzpu0H/TgpC0c2VegJ5lVFudRY1Rf0CJZLl3av7r+g7jfVGcdrsJK
zZKBeQ6lblrGEe3Nq1XI2p815CHFZyeVutGhO2xTZ+o0vuXO68Yft8bcZLK0D+QrDjtWmyRZdaqF
g0AnfDCzlnR1xDESC3pPDdHNL9Bkujp7ml8MTt4goVte4G/qHEsI8nkwqzuLw/Qt2y4wTvCJSvyV
ZCvV7Ma2fpma8XypAI9fCKliy9sHls7VpGhK6wAZFhb4OmDTGumtzjKaaOG4PCE3or+p20uMkEOC
IPuDOvVCruUKJpV3uYIcgXuOUMDDmzesz93VaJVKxzoVIIvNSLPPwCGR961AWwuxZA/UStowY3Cs
SDc7/zqbHxzF+EUlB7kxAdkBD1qIRrfzWvqUeprnc9+eruVdUwOFGpGY03BVi5FgVorOwcxqUKym
UN3X3jN+7oMzPUl8VT1OtDYRgo6s0kq4R4YLOcAbEtC0V+bJJHJiRHmiNfTe2UZGoCppxHnBHWYd
7ZO99CLpwUtAu3VCDaJPe6D4eM9bDQwKAjf2aUUClhho6ACXCFXRA7WpCmJTzL++UqWLs787qefs
OV7aKQjWer89Vzz2r6Op/IB1VIng+cYCuNZSpZRddIllWm0D/3hMyYoS18k9Y1Lm3DcnjFxqHWxL
9q+pv0CguJGtlarM3pVa3iJGYwCMLht6DlCvrx1NtTRkWW8hGrMGNKoSWTmdzOnRW8ME1hoviGe0
tFd7clPza9YsryX2i/Rpz0e2nX4CZK8svwT8G0DAyai/fc89ROTZF3v/r3h8pLUAXQQ/4MGJgNWG
RNp62+jS1gb1sqWIqoFijt8sKgXFHyDoQ7rLNfdbdA3SkXXUP/0Ri05LYKnbHDcq09TrqkVZDwJu
ibQkS1WXBpzJcqjDgSPEaIeCfvsCNbVMkjkWDGCYyzc4XsT1UW8Y47OY2418WB4MimjpuN7LzQNY
vDvcV9AXkvG2E4DXYT4u13X9mUCBXx1TYptbXD/+QtFhkrL5TSXNyD/l+oPlu/UFb+dMGfEQ5ssZ
Ez5Yiwy03XKj1Zt/zMEpb96gnmemxv2FSzSrmJODUW2R1V2utyenV9dkRa8JpWYNe2VRKEPmvG90
CXh5KYTeP09IKdUstERCDjBOlw8A8ce4YfWrfosrblZgGeTpCy4qtKgRm87qjUywbyyMk5i7ESHn
R0CkjDhb/Qq84aqSnkSg9Ma6ifEI/1Hkb6PH3BBiDpqZCNmtGESoP50C+LaTUXPk1UAdzS7yFsJn
geZK/z5Q2qQGEH/xcMFc9QjxdipEnhuZc/oyxxj+QCVSSJQWV6XlwGLZNBpidF2iGC5xAPoL4D4r
testNh0qoZdEaaVyZnPn92nl00j7yf4LSbwb3OqVVhMwXG2j21Ec4bKMD06itZZomp1bSv6VzrE+
zmKWHQe6W6B0dW1QAuM16RiM+7dOVmBsN/pL5eIr34ArnZT5sMhRkde0m7Fg2j7YuVJXeJay2d9Q
6yfKfTp3Y91QF2r+94jSMQemA0fXfD5W7tzLOqkjKq4hxM5Mf4pJmufruWV2Nqx8YzpLVdfh65AT
6h79VBd5rIkw9wCF9M3ZU9ZW11zgDyntSVri75vrR2K7F+ZnDG9SInBHNpcFLCT/hcRVOKX4I0dP
rJm7Xkp9Y+yvEyglGFZRgQDBS4UwCGcdOSeyPyHLSgau/k9DwTwwU/5KHKzaxsrFt8G1m6LGCX4M
awrsQ5WkuqGz9ZrJF7oB6pL0valL7QBDn+rX5YT5kBJ18HH7zB4Sk4MGMtvrNm4ojDHxcrm0j2We
tDWFqGrMVaRjC3rwVhzeAZ50M11AINih4hbWK4MTYqSxN4hFShJVsQa2/Q18oRJInBL5oMOdbLBZ
1vN/Wszz3Ey20ak0TGhWxebpoNUx6+uASYXOnu++oCwRihf48DRWKV8dIYjMWjqWmFqpIKVkwojl
197vS/g9U/gQIPcPWN6lynboLXGHFCEuatULzQ8t+QeCwfP1ymjyMqZOXwJuJ3VAfVvDONddQkfj
B8U2S1McxQYLKKE4sHeP9nqzi25ZmNEmOgn6Nw+xohFbYK64BbTYYrMmPvwFNDTZq0FRiQPsi5cP
HGLvnuu1gse9KhT85syA8iygccvXj8DtYWrbNaE73zO+V4SNhC+LmJPESO+DV/ew/ciV54bgev5A
2Jmpo3+iChxR+39ckBvWhH+Bry3pZVt3YSbWaP8NA796l+RFcbkXdwLsCYIsXB+aUbg9zIUzCd03
+etyh4ELfztkvnGnNYcY62kTolwpzOh3b7qM6ggbL28VBfhF3rxDOGNXMk1ZYiGrp8eLkvSAJVj1
N9BuacmpqCEtAwcsK2Isc4Pg9aUcI2cB/pRx0ItgMRJCS4cB2GLhVhUHcLuV+wwhWYsDWZnhOp6c
n1I696yqKmEnrcHxLYQt4ZlG4xlh5e+SWTrVfD2Ly9hANtYcWReIALh7wOUtrRIohnX3dc72Zhd2
O6Kpn9pzvvo3OzfA2LRnXcHm1EMQMvVjdrXlOUFHJ70VbkMncaJv0z52DBPWZDw/leA5mYdNa6by
C06jcnY9hBjUCHHwbeH+1pO8nSgkg1XwGmMrLIXdwZjlKxQKd85FC4qsVzuz777XWmYHJggUXtAm
QHLt5uHaXfBT5Fuaen+0XXaqCpzfgKWDHTbzcGF9ueysQ7EVzYGlRny91FvNRBpEsbMelC9Yy5aE
LU+weuoUbFuA/9Tvhlf4Ux9WSAChdSBHCn8Ih/62ri1wpPmssZvKdEN3AGU9MCBhitAbx1iWf1iu
3wH9BmyVsYBmaQI9vIZx61f5YpEHW9ODVLOycTlIgmvK/E0T5CkGBQ7FHwibp3B25OypA58pFEFw
GT+CpErLYKN2Pw2WNsP8zENM+viW+EYNL+56yTE8bvrfByGyOP6laNYItZ0FqP7+1W4Vy0WOZiN4
IvOlk5G3Gb8DhnSnQOdUY/iRSw0KsAOMD5y1+ZZ3fZm+g3k4WAZBxNu4eXk6bohVOi4tJVb6/4sd
h5iDhiNdpxpKxprJCXint4cedwdZRXJbuKCw9RJ3xAlJ7x2j2n25KY6vEnIWBGuNtVAa80yLesU6
Bai6bcQXGAi49UEQody65Uk82Z7KMbmo/ld986Z6S43TVRTqwat8pYdG1a5pUF/L/vin+/Sk3aR3
8E76kyA9yZjvypoYlvp2QKBBrvCOvH4o0HQBHqQ1965NA4Q0XJ4Hu1Mffa8HDCK+of+ppKinXZob
eMOMzliXHZDJcaTPa18lVQq1G3fJ6r3mahL2BCSsnu3Oz0mIA84ofglfK2mzZkXH1rwvJHgRvO4j
niJsODk/e9tYT7TvBO9qyjsT8M8Dvtjpme7c415vIqRj1sNhQWi3SBwM6kT+tRvE/5uRnliUF7ku
wTIeWDFGGmHVx8nIc04Tcd/+T/bQ/tPun0pzScgpIjuRaZn3UoKAEnfpcFCYrXSMYJ6H30rous7r
I9imV/TDvQnAfswLcIpNtBQ4YAzMBIZtnKg8fh/6HyELJwjRJkodN7bd04WH3mbJNJR8nq8Jcd+Z
OjfDW/2jpHKYPeeeNm6/UuDc02kE2/oOloKwQGCQ3ZArPguMRR5A+LwoOCpwMwi8ZNJfIZq/8gbd
dX/Tuzm7uKfC3LQjX7U8v4/BCE8DHONnRfmjzA8u7qmSIbHzCEBPg+b/xyflUnim7b+XiAOjNMv3
XKcmzZEMAufjBL/IzkTLrXX1NPeGCaBKR8DzkWU1MSXs7yYBED/oIok7niKwzVorte5Q5zwaU3bJ
f/DK1eirewRNBMt6GohisVBqXNgVsInOC/Xxldusu+AaW11X+7r3Uy+xEfjj3SlWES6JqGQHPS/c
xDbUjpStr0ySGw3L3dZpOlvh7qWWDOmfvS96SnhVVV+bMXK3fOd+zYEJ1BZ6g4P+ZZ0A0w0TOula
bB9hLHei+2zJOSj8hawWPPZ0Mv4ueqfC7JhwFOnHGVpBsmbH/EIbgcfgMjYoGxItSFAiDQnVlyjD
7x0qqA2TowZ+j7pT535zOfxuLdiiSMTTXr0lSsNsQSQupB1EEnseCxvCzrJH05ojFHBAxEf/H62f
6juMDIh+x9QBUSrO6xhAMbzv1RbuGVmxF7zFUJoHSbN9nJJyp2uuoJGYf3OzCGaz42MF1KHrj/TO
ql7U24M4HE/hB21Wc6kmm/AbHaCrfo5U+vd2ncgV3VfCcHQc2lRkir8Df3t28wlnValNQqUTbsIh
ci0dVNxvdLX/5Dj9aCDhIg7576b5FulTaOFTj99NfGVoGW01dC7NAlzHcKySzxZ8c9Z55BjeYnrS
fdIaujNyF/j59ROv+uA4vmQBHJY1rByZ5JKzerUi6QwS79WTzCoijLcOfSRRgObeBNhluaOUuAhG
1eRiCRXkMm1aaodUWyLjvx6Uu8xroO9tH60rBfVEhqmhWI1SMnxEgUgTKMIzm23wyO3IL4gzDNBh
Wtk/nNigngxiRsAFN1yLeErNiQLvN2/TaMAwr7C/9nUXNTwgF943Df6Jwy/7TVN1l3t4NxAYu8ev
gcQImj2An72h/5y4PzXL+Lk9/7bC0qzff0C41buxYjNwes2ritJlWv1Ba4Zllx85vkTPhTcbtQhq
pMCeywcEE0US/6XAQZEgWC2tR/bSjPUK+iExSOXZGJRsEhbyVA1ehSXTC1abzCYas7W/PLfI8Z0Q
JuOxcBKdzXfc6Wedk9IKeChdxRDx+2TGPh5dOBkJo/j3ak2KJBsAKv1dMLcEBdId77zMoNvdR9ZI
I6sPgD2cqiH+OrolY4w/0XQTFvkVFUZusizm9ER4/3jxOhSLLlIFl1uBVKn0zA5VJyoJhEzvzuHS
QCIGHM8FIpr/pQtn8gE0ZVAnpeprIf1q5t4kpHXtHXyqv/bw9YdzN5gQjL+vl+wuvLUY2m3MrD66
4njf/iLseAR5HM7pEqmWO+/7qoJsDyBoKsitjZOvTD62wGA2YP93OFeh/sx1uGPIhb62X/sDbYGm
YGOXuHXCNQviOUCPisjJZSkqcgAcONz8kxRvAAndNL8qRtWfFTEBbMoZ8jBBYINfjtoma3cqfoI8
nad21YzkHmBpFZCQtNmRrHEcjwdzUgLpF5XbM+CFWYUbmHy5YRIrhd8UDd+JQNByVaOXnYCfvZln
ApWQh9WLNkjFcdVt1FyY8GwFum6Fsbtbn0VP04lHTwTa9GAWtP77Pps0k/qeJwC7Ew6JGhlbdQPk
zoqqzDIozLgZtbw+/V1jijc8jrr8yLjZWWT9h6sock1YXDoM8IWtSKZpVqY0jpMblzeJiL5xb7+d
MOYlgyEi2NQfj/lFyzByFKou8KHsi6C/uh60OwrOWQ4rYuhx5shoen+IJUA1CqeScoO6zktv+Fd3
OeM2vpfscaXAms9PrwuyESiXkZuWoBtBs5CTxCfncDts5ojoZs2H1s/I5fDlS0IISAmy2aR8fW72
KMQk8Ny2eZCjjBzU081AaVlD9gxCZdriv0cezQUkZWnJS61wY9wGUgcfdiaMz3N4OXxs9+IO+W8m
GSVoriq0wPXwr9dY1vZnvscIjcPaRC102NFC5yq9pMLJwIGQAPycqYBnV2DvgIH4LEA+lS0BNCfH
1JEP2inJwYmBt5s2N+Xe/L6pNI+9rE/h73bk+fh+tzMiZ+e75P1jlJqDCsDVs740IAwwbayoUejW
R9DLcEnny5Dvgj1PXkSKf+IBxEiaBQ6mWgi2r7bAEB4QFa5NFNFG7LAMkCvf14P6kjU5zAQ1Hjns
FogbHoJuqjaMKR/Fvezezzr7VHruaAIhRTyfgZo2wgd29rlCfYDLqjRznqkBk4IJei8sdP3Q5Jmg
PPgl24PKmqe6W0qXgGHihUPI9EZJBnn3mkXTiu404gAplln2FaUr11EoOf1w5RCQAOMuKCtbd6Fi
05oetmP2qAIrtSZzBZ6vGaC7d/97G25y+Hkb+sqMOfow3zMha1PIxmDRF/sad2ACinD0V3d2NN0T
xtq4ERHNPnP3bjSDpzjxfCAeqls2TfYTPwSPwaO6GGhZ2wWCyOcVyDl4gonthtf0RlWoi6kIehik
K28jnGsK0FpuZbFHAvZYRqX6pK2brg+C8kzGyg9lVPh3K8x4UZrqKLEsejjv3xCPLBjgUAz7841+
k/Pq1jKQ0xAe68eEU8cdbvXjD2/eVwuSplOESQ6bpetyFUMf2ev8fqGsg7sGxaaEtP01nqNGtz1k
MzwGP/qcqs0qeviXOCNlN2B//9Ogy/Sv5yKQocTLgVL1POB+sOLsCcGN5I65PdHbYEfRTTVF1QVQ
iW2rnsvk/bgvL+2MCU3nMFXXxqrEwJ0b3I0CB+XzqogAo4PrQOdiz+ME+INCYv8u/jQVVF1N2hUg
NQ4ZJfTjrUI7PoOsDlMOEROj6NvLFFQa3gGAIkaUMlC2B3Wt7oKvZ7j1L636yqpKz9bfYf7YYM6b
LZyf0kXviUrKO5Vg2Gvp7qatE9AFLXuCW4wvPi7HEPBXcDnIr+18ImSXefQdQYx3kx11ukegFG+e
Yh+N4XLWqvG2iRCrh3wUedAsqsFa98zG6AXcToCsPeQodR70tQMbYMQgRD97cWi0N4lmDABXMR5C
uNLnXygc7Bud7TjYNFUUFEuaAgZagkci9qm5bh4s1iylV8BYDps7EZv/gbrJjqEUZqZYNZeOMK8E
Ptb/i0wB4ic5AMVCp4cXmgn4UZ9NkZgQIW10a9+ArROQKDuHkuGXcwh+VVlI/HFjBfbBn4jxpJzu
FaO1OUVOm6J80d+4tL9cn5jsLCQDXFd6xc2Yc+riUfOYg52dLq9eJcGCixKIIP3nOVTNk1VtXdA+
+O17IUTrBlH4EArdT+B51/MSQtB54lotGC6FY2IoTg/kpbmhCOGBXvfLWUUS83i6y+qKhNZ0dfXO
shoipvv9KVkMaZv0FE3x8btj/D1Y5LFr355UrH0EQksqdtfW+ol8YCL/q27I4kAf/f0DNcoyZ3Hc
asujNEhaPS6yIa7BYJ5DH9uBbY2FNjNdUBP4cSmwE0Af/jFL44QfCSD3B6I7oHYQuojzMe0B2cUa
L89eb4jJXVno9LBhov8HK9a5uomO6zm2UsTdrOXZDad+hgdmuniH/VpE/iS4TGRS8F8naSCcZsXq
/ovdsRZMTnLYlJXSsCaaXrf3kiWNwMGD3+OnqEXi1R45bLxsW/d7EQ9nwNbU5FHgKS9yDimREYI/
SzdYkzNiBnFl2V2FsO2Ob10tgLnIwB8+U8yUwTcOeKiQx3NBEkm9jdtsPj2iMuQ/zrARJ2PuCMQm
QaW2j7jesleEgqJ1v7syJ0AD7O93eKPRSt308W+byg/n5sQsS5ffFAf5CKjbh8CjnAzxaCWJg57c
u7X2l33qViuc9IA+HxBVIlmkEYP2Y7bxy1cu8gvizMvAHjj4nMfbYzMZGPDjPYVbj6u9JlOvDCj2
etUiNijuqzCMLoqXzxmd/qtOIGmer/KpiUZq0JGecB07g56eL3LI6Zic88LOMsmcc0xMOkxlt2je
+B1Q0sMMy3667RvHgGWkWqaV4vFrBLq2ZR+JZ1gTj8mfN6+QVgh+CeyH9jXcvvrSSBGMB4+PKciX
1Cvep3ZGnkQY7CGHrwp9PYEuEbHoteqlI2RXXOVX/SdfER3YRbRU6Mkw0MNRmGQH34UFACOdw8Z/
4IgF2eT28cD/kr3BeEk9i9iZhlnd5LMU58CZIS+fsY6adNxk4QRmnUVUF7GjNDonu+JleQqGQFRx
3x9w2JPZnPG8203uZ50y2aKbHh8Qm1rGYaf5qUz50Dgcb7lEAFOLMfjK7NhNyqsKB03hsi80BKu3
GUBdnsy304t7dOOIsxdRWgBJbFO0n0L6yxMW9RMQzQoOvrQKk+tRBWDaRZatzZS3Lr6c2lifYH5e
BJJucRoUCYd0Yje613cMyrizjAH5bdqFPZcLZ3NeJf9Lmj/Nzp8gmFTzmQbwp3w9N/du7gJw0oOT
dn0v6BnGWeOLCW09NmlCFsUy9vePd3SQnEkHDFU2jzR+WBArh0kqntaytRzoPDQRoYaGLHhVmrlA
uCe0Oe/WaOE2+3ey4F5umRwEhRH/yR5c1FOApyPsaMSIAP+2FRZb5W7B18j066Gl3vBJYzw/HqJ6
C0VuGv1VkNc3UFdKKjWPB3rz/Egam431pvdII9Lh5zsOCgU62wopFe7/IFK0oldfPzGHqVbepMVU
tkAxuJOXUwTnCxhiDAii90CS5q0+KsMLi4YmvLpLfvFUyx36M1uBwSGERh312v3KNSseefWgeiRY
e3bqbf11ptlc8WqSbDgQy+Q/RVj16A9tMfaYbMcDh85nkf92GX830HCUEmxT6d37+qEsGznvtyIG
tdJbQL2n1RtysjUtMijhrjWH+GYCO4yp+GJ7kGNF+LGLKZrjiFYZv9W8zkRDnxINVo/t3CyD2Ckj
zlBQDmwR19ZYDg0DspLJ/zGdKd9aBNlJuKWyARiNSQSwoLxBrjolVm91o9XeD/8+W4IILzADCcN0
RVpWAblfI/3d7Hg+6seoL7kht8X9HmrwN5K9sJ7nc12+nvOSW4x2AXtGQIzWX7AN06aokkzG/qnN
u16CL2A8ItsjNgtMcD9WtpHyvJwjMBgeYBmw3x+KiOrwCRwiPHvi+XeUNS9s3sf34WtnRulvUgbc
ygTqVAy3ygxIJX42xtNDYIHwHrPVXGCbK091bX6ozcjlO1Iz8/RPWj+KuZfS76wqF9nEe71P92OE
a9hTG+xK/Ck8fZwZ5FxZFhTGB3UJLw6Qo7PKfcACcxquKtbLzYhjXBsmUT1w+SEXZwJOzwdJg0KI
j//A3rGzI17+EdwM5wGTFCwDwkjKfdA3MpPzQ4ATHPlAeIlaL1MFk9k15MrigX0bnzjWyJUsqBIz
4dTp+F4lT7ohGazVC2x0GQxX1aN9dXsWgFgN2MNeJu465ctX+pK1/6DRg7b1dHa/LBkPliv1DEnV
vkNCFeq2ZchOo9rbT/Wx1PlM/pU01k18KjKeBSVZfu83y5PS2uv/ja7aDKbR5KemBMxG4EOZUlQT
68/qvObLMhWDaMXhrQeoDB9aPZSwUgfAH1n3j5CeEWzS/l+Nq+FhIDkjplJF2R+wvaTuPMgSQN+G
Hc9sDaZb0YfhZvq5bxiVtd+9oBNnutEHrpxq/2yjfU0GY+kvcP7/6ITzF4m0xy+pU1tZQV0nSjGN
Xq32GLbkltu/ghoaOAO3hKgsOUmYvtQVf39RI6k1ogylujq57XmOBIcw37X5IgmYZaAs5va+yRYi
ACfWdeza/bKJ/lieLq93eQiqSC0hLhZANrERVa0IOkpX9Q6UaLKYjh/4fqM7uY0pEW1JXAFsETz3
/f8WDe/++9/IXwWzN/hXQ0juc+cl11cXGYfINYkLoHddi8bla9gD3RQSWo/3Exrt5X6YhuU7WOrM
coEXdsXO7QxuOp2ornek3Ad/ubjeKa9Yc1wFFYzbdPEVqYK6d5DQFidljjZrzwu5UeWtfpL36153
I+nPcssx2vxnretnNZuKo817cQuS03MNaVUpUYojXEYqE7AMTackb2a0JFas0OXnKAF47BloSBLu
tpIYHOspP1p22a+ExmIpWKB+ph4G5i0ptWy6VDu6ouq3rq+2f1h9gGI3A5h8wSiIzti+iFyZVgyd
RmZ0ZaGM8GZJfM8J77VQk1Cjxfhszfwud+il3mbvZCJOMzaXq65xfeIpDA5gN8dxVEtBV6sobDwQ
stOFo/bw17y2USWyPqZws1iUben0AZzk+Xb0ruidT44B4mgF12g4r+WcPc4/suP8R8VEFa5+PR2e
fFzpmzzXgI75gguQX6iEb9m8e9vGl5PuAk44MJQco8HbZnLVYPrSeGW3s6YqtdtApJhlbJ+CPrvk
7DKIL3+blwt3FWMpDg7pu/jo61hgTko+1v+ZljT2n66YvybU4UXQbknXGEDV96UcOo/9E0aQGZct
VYpKgXwz6JHCLAHuNXQfs0JeoHoGWPWtjRhoQQGoVKshUJva6WU++P+eFM13Md1hDxtHV5Fnso4u
W/ZQ3VerRfPp41b9/dyJjuRlR0ImMBMZvHRVbgsYX8s9w/npoZPbSyAR97Kdfig/dOR63eqqvi6B
3gGqyaQ2avfgbYaIvxzsNt0Q0Ya4cQdNn+QunyTFIBklqG1xUl6UYlQf9APJP466pkX5tKZ11eBE
1cypo3vSr+3NNQqvvHpZ5gx8w+B1ck+DPv6TBFYojJq6vHBNwYG4bJXfot2s43CAPc8A6jFahap2
oD/peM3z7GxwljylBzzYtYdNb4FgQT9G6ShVGthXg//ZDcoil5cvUPD+kWeiWiaa1k6YCb2qnQhB
Bm4w7K4zDDDrnmAIJwOjue7EsSUm6SaNDbxCBCtYj3RwWI161sUyN2hEZTgyLSB4eBz3NhnTno9f
ZQdpPDMQok6pIMANyUZOIVKYniOdUxYnqeNgjmARlMGOCsG/ryHXgCoOw9ukuL8/BDUNwdki58xw
0my/EYcYykdkwSAFeCHgjX+q1OXFzA4MCZYXvqiNO0FXwEezn2Qw72VwNnZ3XsaBw/Ezr7ZjtoNr
17tY2a1bfVPZdJyXvPRmU7xvZPm/ReAcMcaq+VfZnyEHuwoPkHXP5yo5Og8INpekPPRLmL1I56J6
QHPDVPlzp2R9t7SIiOT8zbaldAfHBEj8TkK5JnMqzEqe7p9P4VpJM14EymSXovAGAlYlcDLKqbfh
rHu5V+bd0pSB0kLnuxT2Tn0q/i9gXGC1ZbQo1iZ1kftwzLAyJ8NLfP2lx/GOyLmu4DbLJF5khdEz
eK3Te3scegq26cUQlPZhUNDKJX2JWtkWrR8NTlDjiFBQMDhVVMiuOBOYymQ1AEuEZmVEEwLDjySD
nguenUfX7H1MD8r9UBaaBdPnU32ev1LjXmk+oIzWVY3O92WixOU2sGj0Zu+lUPh8AgcAYzCl6zBW
NFew6jInls/ytLipJ1zFDVxqZkn8/oDNRuzAR0d6s/F/0qkl/yAWJv6QWP2gk8R7GvfIi9HSJzfy
ZEeU570MtoiVl6olVrgEX325I7OvKV4iRab5pq+b96ZGDMe57mjUwb1s5GfQT0HVKzvQ7NZtlJa9
5BGEI2rlpF+3PU5zBVycfO92IsPBfsuaLM59fmC7ASeBy9Wk6HGUs8WItDzhXXxvqZVB6QZyZCMe
+yiojNnMxbMLv4KO91jYb2kgehkaTMcNGu9mHl5v3ITaMracSjAl5YxiUw3Npk9lVm8HwOFq7QEx
E+ROp/DdJghb5Gq9AWUh/au2HE7QM6EKkRHfVjzXLuHAjJpA4Y2AucKerdClnzULpJ6Uy1MQiZsy
Gc+0UCkvtmPWna7IPcUNezp6bsJGIhpm4Oh4UnBPZaqN751wrC2a7KPj4mBweuj3iFxC0KdD703b
N8KNogWt3BnkFxKafA3tMgo+6dWLvY+jck44iPLXJUnrc9I2KFvsk8vnABVQgjmOxqD+CHbGRD7F
QEndI7W2GiHJEF45c+tnFFOmwLLirG5CiSlxGxhPyGI9vfZqVYvxyarTsu82KQlk9xMSt6WdGI/j
02FxzZrhtJN9DwUxEKr7R0tCPuOp2PoX+gq9zEdE8qsto9zJCA4aUsR3i1h0uPlq7Fq+XEwaUOX8
gt7QbU3+25hXVfRFBfIFrMXlE5+KrwzAwbpr8Q2tN5VvD3wPS1Q+X5MokszoVMClp20Hd2B3x1FE
4HN1oTL3HYb52HTs67BLFEG/BiPZj+D7G7OXwmACzwssR7C/QYxfm+vb5nZ3/l6jUPm4mQF6SCtn
+yPWyMCZCHFnwcijlkUwrX5WQ+VXHty5duZiFi92B3pS0qYBhltfk+NB/0LhYdwoj/a22LkbMqkz
AjscrmtP/TAXdX5hlVgKaNc/QQjQwPQorO0M06wykVDsy8+2GeTZjnmy6uybMf7KnWyS5V7HyLSO
/0lB/y2vkCCHy3mLwx7C2mm0NXsshlqQaw/Mz3zaCAx76e2IqIL4JySvQHTGSFlgH2DikMkdGjA3
inIfXa8wHMaahXx03axd0Tv0imcOdvzmGujoU47makNIx68967bfzWMTHrv74Cykx4y3cMOJGZNz
dQ+g/Zq0M1aJRZYAaHculllSQPJGpvYQ+eoh9bqAvLF5UI8xsu30Jy51MK+tA37KEXfhIuPaC4Gz
GRrsrkDIGSBDKepgV2xa50J+wTg6MahgZe3DzCLLPUizAM4apbRyze0OQJJGuUUe0Fyp65R4gLp8
vhpA2mMuHrQiPyIBKUoKuI6ByXyd19lFCG+ZUK24QgJ6MFYcSJBHtfIr2RcRr+9p75wskeCqY6TM
ic/YBifZgcg+HCQtLMzTIpLdAgv2maVpGU+SZKBWD4H5cejcgBnBY2xCUdD07eeDLhtAMrw7+u3/
wFPNKqW7CpEt6FTeUYJVVip/YzvO8BH514chZ3cDsvng9PFJh7YXZliBgSt4z7/34Ne9+TifdHDv
0gg2Oob2Ru554a5KIcYdeq0hC91cI+3MICuWs2I0QmJ9c//nPIwjM4/qrnQsKJHxM7EbGWhKh15S
naaiaG9EA0cmZxvff68qAGsJ84RchYpRR6W5vtLk8wKKzJc5iN+ti3WTXuhCElfJ1ayMaZEM7mVJ
b21ndpvdOBWUQatLAgyTdD9ISiPwDWSWQzgTP9h/oMpOoiVlDZjBq9H4scWIzZ1ZRRkO9BbfUP8f
KdQi74XeTr9Kd+igLEXImAG/CV1KkOVTjsOkCI1GtrfQjX2UQIpLXEmKyPPQJcfYxUlhuPfGlKnt
Y5O0/vqDXz1NGLXwKUG7GOR7O/tQhm6N3f0Z3lwRnsnkwr1bAAmSPQNkZUPDSQEmoLFEtMrpj7HR
emN9A7Wu+52REzWqtC/gWkJ26KH1qqbHb01Q6xJZVj9PiO5Xrw4H5zVdYk2/MVTqw2688pFz8zeX
ACAaYJZbZVcXLCng+FoBCgwEycOocDx0PxfoSQKO0VyPIDa2XKOtQsTMOM4nzlNkwhkh+Se1gv9e
4Xc2SHTCOPOVUuRmtV2gn1n6OcbQGD2VCc4lBT9mhf6vuAq7Aq5lhyl0MyyHgQa876Ffl1SjbP8q
8Ca8cXsvgzp8mLe3s3GEAwLM5++W49avM8dkkBAwuXEOWUyEy5Rj8W3UMvq/70Ez2UO8GrTTnA23
7OZwmNVAfidB0E0lvPZOJQ0AtKLIvp3Fe10WEjHOFHdJsqf/SfOhlysSyr8T/ThLR9kf0FUhoyi1
59rHbm/GT1T6Ylx7npUEAzFdgl/MnhpBGArZniUkqjzX7VkHaLDEaD2hlUwltMN7pq36v7XjB6DH
C/rNO0Xc1P77QchGpJ8ITMNd3rgN4PyLNFdM9+t1UncgV7h9JUT/IatIdk+OkklSFHMWp6Q27deF
j6VMfGdcyvcFbM2xcKXHoM/VwjiBrJ5PuzVd16DNVZQ3u9SwSbC7jHhODcMVEBpRaCnwfyxNYTFn
lcxt7/yd1iS0yIY4/wgKEW1Fu1OmJjCvgfnDhCH9cA2AiZ/LUm35Q5MXO6T2KdnbmyowmMh+gNze
ZSutHXg30npX2Yj4bnUknnrk8FPQ9uMwpcsE2+loExFz6NUyXg7gfev1R47WIzjF70D6QVRNV+pO
b3pV/3WufsISsTcqKeuD0ZcKS+rYQO+UzaFHKVKC0I2IVtevE6dapFnsVA3VomPDeoX3q6RmXiSg
N615GR8A5G0beTzSYrQlkihj1HAAcGjowlQcFfLSxRZ4RvWxdV3dHyc38zUDOEHFRIluGDIRSXer
9M4d7LtjNXL3gtKaHy0G1cMJ/nQBrUif3QKydyOyMZ/8VOk58Fq8+8ghu2jwJye9J8u35QGeeb/b
fFISjT9KmuSDV1yQ5sidlR5O4eKL/IZWLkgAvL2GhCdX4whULWKZTolmStzinQEJgn0WosppA4oF
ZwS0Q+zleN0J600ClP1rn6Gkv6nXyTGcEidMJyvc3gr5XlP2mte+d4YFRI9ILgmdGlovLxsnQsQY
n+6Dmea1diOxqxLDnrowFgy4js8hMDjlUzj3oTRJjAVxRHhXpxkwtclRe6T38DCFsclAyUu6f5d/
YicMWOG7cg9+VcheTijg/kL7O99W2A+Le/nmu38VwlBe8i6g7I9cgRpyFMzadBjgUEybeB1GIHgd
XDkVc+NA9Dp16/hR1a22Kh/qjaF/lUFaS/gi9Sx2L0YpAzgbLJZMNw/lsLSFwC3t/0HBiZ/bnLUz
R1hAm6ynWp27anMrNSZl+K3wSL3BA1OT++C2mg41bLvqaOWS89AY+UrXYSKV+C4qj/to/mHDhGwy
qHxFXg9D25vAGJeMDU4t+VDL/oI5o5pdoVEJ6CqL1sI1xN5guf9ry46XpvqO0YVxP7YhDX98xZaU
5OQqM9Pmu89HL51rjdMyfkY4q8M/ZCWOgLWZJBA02w7xARBNCqrOIm1EAWMJlRt6So6IxjOeY/GT
6/m64EFBxhKxBe4p0WzJCy22tyMBNGPaRA7UD2KC1Cl+1PgEyhC4uPu5rQIwgy9rFGjq/H7RhRQS
+Hbddmm2bvAFbGh36RfhK/oD+BF6rqWasByPzEcy8UzLHKEAYypVzmhmxFmcngWghozwz8ndf9ag
wHugEZF7TL/ouGHXwSBdMekvmpw62nFr4SIUyEfldU8CWuOUWNI167tin/vDTb3SUze5gftNEK4j
hZ/E3DnuYJ+idLVSrRQ6HgWg3UgmjWzai8CJGXj7aW3UMVfLuoLk8k9rqCHmSBjH41K4iGzuT/TP
6NL3QhnAi4m3NlRavFWno11OHaezIPaXgVBIksW+Q2ZjzIns7Q6D9Op7+XMtfK6rEFxlkOMlD1P3
Hu9MKuhDdINo2ZGQWT3pqDiRcoLDWJHcvCBs+dkExrPOg6r4EcQQJhbeDO4YLtN2x/ZeVPKFS8NZ
OO/p3kpRnofTrlr2DXG+GIep64ZEjgtU3qjYQy5ouiD8MPi6HlnqlRIDEac0VUqqv5EaxZyZJ4fg
eaMmVhHTRBWIeDzWHQLjRm/+1p2VeMyo22eVp1FZhANx6PHNmfID2iKtDt6qtBMXPNqllB70KDbd
e1u5eeSSgdWh/IzBAaxYVJ4JSxPxh5qusDRCvVn9OXIOHxxwf/s80NtLCcm4Fe6Gayvp5zIxWqZd
fhfDOVXDJpsLqIaY0P4dTnaekdMi0hazzTievFG6beGKOKCDXUfgh19alZ0GKVECSLjuCGeWxo3T
yjfgBw/3d1wKjkO2CahhpwtC0TasX3EwrFoun1b1CcMRxAsL51QYxmw2TFz6FkUpf+zf54k3sv6N
ya+IXu/3KbFm5HQkmMKUgC+pQPeIzLbhjzcY0aySakwi15syz3TLV5sOk5zJCFNOP/hJY5VXC95N
PiaR8Hfdos5c3XI0Bx1fie9xO397pDQzOuw+5DW+/12CAtVXhq/6xGDzz+WM2C71at5oYwC9Ovth
ItC73hj5alXgXCOvSGDiWiagMwaOS9CUjOnuUPoayeyBKgOi4Z+2fkiERm7CmiMnHUwp4G4u7/ax
KWoZIW2bii/23RcJzZSibUAvNEzVwbbaypRYCduGjeFhpKKbI1bFyKYRg5waVnI018q/vfe0qlZe
4+9lyXadXQkz1ItXSfJHr+T9uAyIYRVtF5w/R/UbwE/kczw123rHJ0vDsdwYfzceUCmCsKUneNRy
9Hv67qYe/Xxp6Pc97ZO3SdtdvYexMqrwenXaH2dAz60PUJL/Rq5ug4vLIlX3791EUHfFxD5tED5N
pp6teJl0TRFr1KlnoPXeT1mfhJn2ODU1xkcyGhdceJMk7lKxz7TkawloFcv1oL3C6C7tv1CLdNw9
eW52KBHfI70qHFnPz7XFz5N1dQNqI490MiPBgFHPLqhkIfeaZwJiuh8FdTTc+R8YrOLvscq1uRXr
Cwqp5REyh7dkODQVzrxu22ZL0Ld52LJ4yaqw20d//nLcNw1RHdYgbGSwfnXpgAxVh2rhLm0e9zpn
Eu1gzU9oRvPa1hreCPybVtFjuSZffYppYGPCLInjvL+/2dIhfRxi27131nT1nUgH3irIVSNkA5Nz
b0j6KlID6rESlo34gz/yuBQIz3ouYuMRVmSR+SqGXPlOpjKAjQs+INITdoFBc0f60ycRR58yv+MY
U6/cqAi6EYsCfi/+kxgo+vLVOtYgA9yUx9xBmNM7fstXdXkAARB3z86bsW5NKFh5iCxdbIYbFXvs
7Mo+Tj92Gt8e3OkKNehycje2B+dAe0zhJlwyxGFlEQKDc+DJP/VQDmADiUH7yDA6ncwQVkOq1Snt
YBT0uuyX0Lg/PdAShueK6HyHZEk6sGfui3+IskED7A52y+ZQQh4gjIRCjKcMGtI2z2AK8Gmlh715
KDpVX0uRgFDqyk/D2goDSoseQLy6N9nWoWte6RWupDDaEWnSF+inlgkW1VNrp0CZ+LbvCa4bVxqZ
t0Z0uxZQnQWs5xrwDX3Nh0MGN9OwEDfbU5r3O8Xq8Zw+OALuS7ohHJR8pHV8iEKR2g5cqx2uPpoW
IqkI4rN2jmiV4GoyMPfGVe05OiJUNxzVtjGCMD3GfbcYTvenbdWLEHFED4IiKMH130mnR6o9WLTM
CZ4LMlmMhA2DbZEmGJZjgnRo57PryfCtlpNxReFXy9xUkBhROiPvCGc3T4koAVlU5jWl/9fgXoHa
/2bf1QzH41otwRS68ZLrle8lMwSQtqOCij9UA32zOq8oni+ouk2NF4vkfmOFWA6gqM95BSFbfK4T
+TTYDeivNBxMrroEkN2fVWU4MKt/Kf04bkJzmCd72HLLezzDKmaEyjltYhb/BnaIW+GidAOLqKIM
cJWIFvozVornaBVxbgYHTdisYcn8Eii5iGKBf9GaXC7FBiwdY34uZqKu1bFZodYKe5i6Fjw6tl3+
F/LdSTfD8HNU86iEtLoBHG5akHnQyOtTg9Q+l2VdhD7ON4W/wo0wt53vzhHdEfa701bcpCJ2IqhB
m5IAsRdoprh+wBwBXd+440++KEIPv9ocTgPrV12LKLozk/RM7ovj6tacGCDv4ZwfhMxbV/H/3tZf
zL/AzRi1Kv+2qhoKUwXxI2+oTZc3olQk6yGDWc8nkfFxVvvuNbe2rnYBOwqlF4E10o87WJk1wPB7
wYYbLTmeYH6WH+pUBVDV7BtOOYIU7jwLfEnRP200WMbhrMV6GW3GkZI5YmuP/jLHTK9WedZvyQWr
M/4NrJxw+TnpsVFtiNuuHqN9GMfD/q6STHXtsH80ceyCGGwptqHVMdqdoKTuR69LdupJGu+A8xic
crGHIvDdGfT29IgzFVxZfyX238w4c50WfBlWicj2cYxED9Vz5fdq+OJrDMR5i1sZOfAgNE2QZgS3
EXsLMqsIuwya4b1ylvOOwIIwho7XoQXHtMHyTARsXWGqfqg73Y763UwhwMcmCJbAS5DLdmCZjX3M
Zq33w+TV7Uo2WXrCVj9OH6axnJxyXTr6ph4qloZJK60MPlQ8DWhUA+reIINWBjFP2y5cwjA+8Toh
whOjjW5wNU47n/KJUyFI9LzqfAnrYx82/JEApjjzdiPoZieARZ7K8KzKck1uLuMh4ab6D5ulh4Mb
RTfGSA0qxZTYXpLBHC7KHc6ZBt19PcfVdmxrON6Bm1d9fjkJoGLRFMXO48D3zzziWPZrz74NbGSM
sUF/sJS/Aledp1ZA+2WmKGXQJIqAjX54A3ANmQqttMMOry4bdTS9EWumGBuU6vRrDdu57EIXOazt
3AMtCKxa+fezbT2KvItzJuWIUee2d0IY17vpRaeLLg773aAI0OvxDMF0k1QsAR0ol+fKYSkvsv2u
G5lV0noOONlmw5tYAGctYuHL8LMY2MZYTociF7Qt8hRpRfX3aOX04CI8Jo120wYPNxxoR5cfLLj+
MtFQ4MF8AsIvMp+W0hkwm5xzv6it/S7YrcrY0FODCHc1sWcVLxU16Gr1Jis8d1wwqv7EXVYOjO4p
CS2ZWNT3R3hPUAXJ5M/OEwGJZjlX57ivT3ze+ZrX2IY5FUdvJtycmuvI2IlUPb685+JEa2qvRmEI
G2gSU1WwVTejMBKb4S3pHSYIwv84lz/TtMCktZELhgfSiPljgvP57YohLWoFq0DGaHggp/4SQnuG
lxkta7ZxT+AUivDyNWpLlhoy+Kf7M1rvgWjegQaPieWteNWMP01r3H5TKpEKbY8jOvBd/RP7sdqp
4NiJVROOh0fOiehJvXFSI9wutm5w10Q1DmKcOupU7pjRfiKSkFV2Jpd4GlHk2c4KLkPEsCvlMSCJ
X65GNoL3yDrQ3MWPXbQOsG4gkcI1G7xY4GTNmUDnDCB+Kr7+W+q2hMeX0haynJR5TO4F5BnGNZ+9
Ox2JVoS2+uu1pccaAyHQnTQkulreBDrUv0ehUXiTp8zw/S8I9fFiu7OmWhxbagCH+CP1cB3/nrJ9
u6l3YUma1aEUo7WYWb3xGjy4E7rdnIoUic9HKu+A5wxJz7SFjXCMcJ1m8kLlae1WVcdA9CVVWgW5
1IXMKekQk4quTQtSg66kjRkRQbFeCtrf1XxiSUPQ324dKOOyigB0cdBbsQeLEOhN/ehDjK2sdR9Z
Hs6umA1gKJ9lC4LxzSP5wi0jw0dUWpRPEIvB7pa4dGGNC3dyGQNHppVnmGhV5Ch/Ci4ZAQ0bKiK6
aCHo2ChvbXEE2Yc5BoPqQCxsKJkrsXCF3gX7PLXhx31t+ypdNL06tpfEsUaqoKest/Mrpdcw0Vb/
mtvvN/w+FSkhv9rvX6uEl2QCy74Xn11LBr+55ka/mFfTjllHKdK55IYPNLzrBY6o6AESudcBxpEI
r2gGDY7+R844Hp6T0h1W5WwHlPCfBVuWiuDY6G70inFnyNvkIK6PIWzwlTXNMkvnhXeceFqWJ8//
OzoLM/+47uFomxcmHKwxVTALs6eykolUdaaVqgG0ZLkARgKDZlJ4qU9LxbyFG0PzHbndseDI1BOa
VeA8rpJbF2g2RZP1ku3DnkRVYtak7zGpBc95m86IuiX8tQDgFzjEb8yCBWb2Ako2301VYXoIBt+L
uHumxHwuwtkCBZgiHt0e7QKeymmhvDilzqNoPXufieLEuFACZG1eKFsWCb3lK6x8rZhNs2lQnyxM
jA0ymz5/nGH3OIZ5oWiwtTMYlg5TBCn2fgvroHJ3hwmND35EXS24vJYSAfZBIn1hD0FgFo5g5Wfo
l1p8M3+bcho2Fr2IseKnAEfNySnw6xwNCX/P6p4XqU6m+ialSpU3ju4/NW+YBeBqbz4dgCNbl4/e
oSTHvSBRSAdcSloHp2OrcuJJdXiCInu0JLvvr6vcY4L1VKC2zeWt6H6UbQzdowWOZ5BRbmRRvjIc
rv/fy+JMk7wIylDtdlTz5B+8DWCBcuIgefGVaohfQ33yVqg9JEVRoRbKYZGDql9wsy+wGpL+W8a1
h3gl/+HLvxhGFmDf3P7TvQyYLBMIKKUBOitqI3NgOtVkGQGJHvW3OCwMh62BYlYO0bvYtlqSPO7G
ZCQwYWhP8qj+oqtKuP2rxuGDb+fP6yAWXIJYIOq4tXvpCua14r8jsVhr3uy4PY0U2tNHa18IFuY9
VaViuSAvv01R6Awmh4e/BkDAuIdzIT7v8lQBlOhyHTIpPPI1Joo66ikWvX6yVf0c7Lr7lLlgfYbZ
DfKeqt5AmV84NSmFLuUsLp6YAPZ9H9nntCarbDixLd4V2G7IpUmMlvcwsNCTvK7CzAgHFYSkECte
7GrICDbN2ua+tqT4dGJShtytshmjdbVbIES97zGFAnRrTPwSO/sjIk8mFiHuaQLMisWCaOAoaBm7
J32+aenIScvYvegqUAJPi9WAzpzLvYkh5RI5jbSbed6C/z6l+3uM3gd9+/XvE6rV0HTZnFiNCTQL
sv69Mm1capH+9jZjLf99YDNuydPziti9rXuq534G51lqWK2AsyVJVoD3LU1eUBF+SFTao58MLEhU
DQtKIlNWGKYfVV1mqf3KgmCGVKhY/+GsHulq8RfpT0cu+K4qljusxgvF2TEgbx57n0xfYDipiCzK
xabpHIQZHtCPMSJimXakiczptPbKaPgyyeywQnmAnKJTVrWeT/4Kn0dlNlEqkALp0El5XILNXN42
NPtvVQxmx/2AHdstLDzfSYZtDznRCO/uHBj1rGEbCEV5sv6GrO7izCBTzf5/sm8PLasIpWByYX70
llRWJuHHbmit9kjItuCntubrIxzy9CY43hnX9MseFB5E+R7y8ZgTOIg/1k2J/LYy6phXRm/kbraA
73XFZBZgHFtvJxt8398l50KAnTJHcfy2NY6wEyPjnkFFAaLQNJGgUkeo/IxSlO1/LhgraDgSnBn1
wzlqx9dZDR5oF5rjth6U+6ZY+HuYd9kCsRsQBhH40FhkyUVfHZPJCerYNM+uFirnDe/IIwyaM33l
9zv8BzyUdQG7dnb5HHH0LHIuX8pyvRsgUBxrBF5k9nmqacGW3pT7o86rstlgJRa04bydor9BCXiP
T1gM8hn1E6EpKIiprBZkPa0HEWQTBA8EgG7PSdLNeiS6K/Tdt8Bo/IDMQ51/eMfCZvPB39pEXVeO
R+g2UDITqxuPj+Gkzr64LlFrXbyEF36hUEDf5TerLJhD0c2uDq5vDWYSo/2e5Hw+O51pENTTJ8bX
IgE7cyxtrj9IXX2V+kFtXxO3rjA1rLolaRJ5n+0CW5qBbXqHqig0+td4dTsDQJ+mimwKiHbUMo+v
/yR4Ui65HVON1w+MPJbCnyi458R9kyiGxOmMj8s5PEXnlxIZMuXYRT8RfzXVwYz7G19RlJV7CJDu
GlLiUQijbpel6dQrfVvXu1jnHn5BGaPbXbsMCMnAvDzZDySGpJV/1DpayjQXrxcMLTDaRKo54JN5
xev6XNzBntNiGZfW+/kSz+SwBU8DCPEGwNucIPiuEN2xHtGc2RJV+vE648k3iIpNJVykYeXKmCWP
MV3oB5zvXId5iVGUfLpqxWKHBnC9nPGYx1iXOsYM7il4PcMVWIZX9V7VGd1mZb/nLymZbPULgor5
jVO7Yyl3DSv6w9ODKCjmoDGaS4n2v2Z4PIp31yWt7KCyZ3Sz+lIT8XvWDF1wevManL+s5QU39hPQ
JPOhR9k2dp/DvGvH/fG3Rl258e88YcxvoBaG6uPuPee1tjG98kgfJeTsRSQT8hvp3ha9egHBNiwA
7nHHeArz1GNWPwe7RqViXvQ26fc7QRh+55GRq6DjcZD5l2KammaiERB9sm1XC4FNYwDAmH7+GcTo
qLu/mctx6Tln9xRalsg4YHmRu2osBVJyJJOMTIAxUv0QmaTt4L4ZM8K5s2XOgc31hlpmQkVEhRHG
zQ/Gez871jtQZ3yTkFXH3qJXyZW+ntuvSyzIPVWvH+iHrkbXG55FmRucEbnpghwcCHRjeqg8L0gY
C5C/OLgi1NLdOD3/Cxe9DSbXpHC2cnYqPBbv9DquYZPn3+91Pg4DrMoAkYcFvkPMMofQlYYldzy1
3QfcliPTncZ6e72Ih7m0t2DU3asPkVlPR9lZMGjOMubgOcXFnEKIAv1MhG9tFFQyMXtUxV89xZaU
OjfWoe7Ak7bEWSz/S0b5U1oLvKqIWdT40udmF7nosDbeWfi1RA5WrjTckTykp78An4hSPW7YBRYh
U/6KL0HRqxy/4i6kjpJ4strBO7vkilzphlXsweSlQrS7ImfkzN7S2Ow59B4lJK+zZPN5xPj/o2xd
WAynI2k7afmNWNmuiRQI64yN0zI2hvp8drBXiSwdoy7DagMRcOGOTf9Uz7VVTgzfBeKQSc+Cgnbj
M3WS2LLO7Dn9L/jM/iFNHFbAhuKJT5VbV1svDVJAQTn+8gjwcTTFKGqDWRxEYha8iqNp1seW61mS
nNEWHvq2jGMNi7pUSgWgYvf6E03bCfUVTRIlvddHLxjh7zPQqR2Oe8HdiGZKBNUBcfRdIq8fZCXZ
jj2TVs5vNtirU/p2mctc44weORt1kkVF4lOejl6vMyIDkzsmoNGvbvY30qItnOuSowYvOE7zUwzc
i4KgBMHtMMgQ6aoe6ZVIVatTEcbd5oqPHfTocKo1pqSxHAWwPcTNzcCUGpDmPGe8qaKmDIM4O43r
xUUP5NLYHDZO4VsRxIWWOZOuXArMqoY1UvpTnG+1cc1cIH2Lq1fu8GJ0R8xhJuy3Y92RhPWgUOYN
9oz7GbRbU5hj+MlzBx6+VyDycUhVpDu2FC3bPwYO4LNdEfItXA3mkk0owy5NTJUFlnaYI3zk0yIm
inzT4DmB+iSpFq2fFa9yF4/fBIfBnlVDG+LFrRfxz8hh5aLuKevnMYXHtd7LCHhnbbneM8THAw6/
mMwH1QOPjCqccDDagrNhQ49CFFP9U/dfdhdgZ9fRjTIPKGIcsVB8UPuMh5zA193CMODgHSK2jMZ0
a4iBXiANE4XqX2OlqlUGD/NIUIx+oTI/Mt7+YICsvdAlOuS1fGZLLwGZM2a+1Rq0Y1FQ2YlJ6vA2
9XTrhJ9pjNuDr2ctsG67ZRZRM5Zv/qrlBAKiSvArvy20wE13l9U27URymmHmMwR//BlVTJ+w4APd
QnG7DNWJBk7Of4o6jG5UUko5Gx/CYJnAVcFqEdpGl0Bc9HqG3LVe/ApLeRt9lcw1j6NFQbWBHwxa
KoRHiD61BeKczxu31dVXBGYKYXDieTkdHcmekLhdKXPzigJ7WgwztD9e0On+SHeLfJGWZXXoL9LU
HolHOnKnI1wjCjug5mmR2a64nIKCogix7fuxsESbgbiQ3iE2v7Zda9er1FBE2FpjNYtftcnGcvq7
mhcTi2TS3bP7ZD7uzGLsSGj2hpsIEs9ktZftoWqkB+AQu2HBFi2C9US64st4QFkyqqe9JiD0xp1e
HsuZMB8ydUH2cA2JMXt/rVdj18bnxCppLP6SAtFDkH5vjPyj1yG1bcqNi+B/dFNXSSBycoTmgo3C
st2Wg1L1Gyjf7D68mx+LJyV3qtHES0ymWM9WMhd0LhqJPWErCZ1/q0yKeIeMUgeld5NzNJmZhNRA
JIaWdpdid3bf1n+Z1MfBDDw8QTMAN4OSIk8QxEmBJNW65oRdZzfbhlukwGhB51+2IkgjQRaBV71z
+ST3oSRm6nKQ5XZreEPgg2tLXd/AxIvkpKzj0skNTz6WszpU0y9ax+x1jmShDvAon7rSk/kGq7+I
z3TWgX391tTWQE2p04OGzbQX0Q6Gl1mWPkAS0f/DJg9QcH3wuEGpdmEY6+IQeJaGf6/FrJCV8NY0
4aN1PgbDlFUS0ceYq2qanEx2Y6Q2NAsfx1UgFmllH5OCIcRvGc7IXCpYiBnTA3yoOqyP1GgBI2p/
W9J4lBawIJgidoLwSTS4Yf4L8Y7UYS+wLa5NBpxlijp7pl8GWgUje5p0sOc01GL8uejLojUpoieh
trnxPHMEWLsuzTKvm/A5SoZsj1YIY9/XuRQedOQhCGW8nE+gNLagtBn+1baNl4Op02gH86bCoR5V
fxMDV+sirDuw92xTH/Tu4AD/99Rgod3HsaFaXaAC4wzOxrGS9xR4FShCkV2/qkixIhCCFoM11DM8
j2Wol9kcV8lYSOrVaMAtf2hwf8mexJB6Uf5wY1WhWlO2CXSX1aG2pjh4Jsaql57WggTqJZHhJR2u
TevRcPpBtWabqZvh/UMvfAH4la+AJeW4MY142iUAk2b+uOWHEJo17pLL/qURvaWk+nYivt3KNuxN
7iIrEKybT/Bm4pBtkRZg2Ua2fIespLkOI3lHb2tLGlzZMvpOJTN+6nwcHPy7VDgzJfxLWK0UfRpJ
PvVd/ry0Xa3nLCLwZKgpARWxoG5VeZJZGz70ajL8O39HYWxM9nu7FRyFsEQkSHeaIsK0U969/Kko
SD1EBgdBOJ0ZL4dlXJDXeUuJDEMzxejV10dgbhPLNy4J641IGbnGcvfrTJjbgb/VyoIZBIQZ7pBm
vMNw/PgIaHaHPKjaPDd32cipJNXb6zk7ya53DQ6RmMSdmUGytwU7THgU6TwEIh1a5FQYo9ZDGFsr
gnZ+qvHtbUgx9TIorFAeKDs1hnMe8UxMOKirTEgv7/5rAU6aqesIui1rn74swVGF2ZTVnjNB3V3G
eeoEZrkVwLN/lofQ/G4alBIAJhRPlDhTr0tPnwsd8y9sd6YoYwE2gG8EjeQDO2l2Y3qMVUsS4xEu
/5oQuylf1VyLLoxtqkjMi2v7sBqu+q43ulLvTcGLPnwJoFNHnX8O1KygR//8XNICxB1HZew2nAlg
Cca7vPJwH4BuwyaNnYwUbOuIWlcFEPybYZBBJHmiF929/se+c3Thg/HOjVlplgx28ErpHf7PV/dQ
sONySIGo8YZv9QIjeV/JagI664LRGah+udSUFGXabLNG55+ke5u3VJmMJNT0PCvCoPyEk4nF55sq
dDi4R1MX7qtGZlJbl81/fs7jkTnHlDK3tWNDo/QhqqTgUGtL6mjda3v39A3/AeapIFN2DdqCCpIj
CY4Tj9ZxH469zzKMRXaXt99sTcPzIcdzfqYAjrZb7/NzGCaVFMtkjAqNIIfrynlsz4vxW2LXLQy+
UrEOdFNjL+p32DYWaAPlxoy4U+jenvI9EnVxc670f7qh+R72e4NZ/eI5DzEc3Yj22dyxnlTymEk1
M5zU8AIANoimRQMQWx3rDrAkBqQ5ujqVLXCWS9m2Sb2xcN85LA9JJLCjOeSGuwb6bK/8clABsYdp
Y4NYNtKBCcaSbk8GoJGNEHn6DSy/pGsVcT3oSKW4WeXLEjO1UkeNmXnBxkBNX3/jP9ckPcbFffjp
xc8yHsxJlmG1pUDkn8Ezl8xiqlvDbirB9HvTl/ZtpByXM+prsmT7YmFiqsqoqK/jlOp38NcY7NjJ
0yb559LkaupXPp4u7SmbNft3ug4a6pt/inluK32iP/4qFT4RyRAsP+F/N9Nlm3n7rf4q6b/1j2qU
BLZuVyjL74h8WOqR/y1a3ApcDQGDXihgXA4pZWMKX7L4QAPhpTt5RI98+HbFDIHw9tl1AkSp1+YS
TOdn02hEpdmDur+G84P7yO2XDlT6H8z2ePnJSBvqkKZAdzZ4HUXvPzM3NKX8dJrnW78NODCEyEdw
kQR/7bFWsNN7ZKo7a0cFvLyQiuTeXwgrzmb4WDTCmfy59LRvBi/9BWu4zLu6hYgTPSXoEFhQHFHM
Z/zd5tB/8Qlv/I/AVLhwM/QrGGrneZEdiFjJpE3MaLYrVjeGUajwAActZ0mskP6N/eld9LzsibvH
darnEbJ8Mz1dNiMdlUys83xUb7C7IyRE3AeWV9wryUBa8eo/jBuHZ9dzGOnJOvkxSbsSY/9PckLw
rNkFuIipKfIKDAbK2aeM6erNozL0cs0lKMZT2+4HOOIPq8hx1YUhRqSLqvjhPhfBDOK0WvSttlHQ
9WVCKYPpxPDW80+z6h+bGiWDIdpQZ/FGfxTPXYcqkjVwakC9D0stgMo2iasp5v9TooAKYLweUk+P
PcLkTcDpT1xvwfP4C2Uvb1ldng2x6EIJsU2ujAZtOzfqj1iy8PQv5MsCbeP7m10jwjf2a0fg7VG+
/293Rr+W1w7KXfTeTuaPT/BiYu7ViZWKbMmAJeplkLPSf7Ajo1b8hnLmFdcklgic8HofT0o/UbN1
XhzcMovZT0i/CFu39uGWOlLF5cmkj2+viMPkNfwlFV/wj1oBf0hC9PUpVFOWZ/L/ml+1OciJGwpx
nRbmJhmjezSIim8CCXyMsuBomAkvNwWrQSa9BbOIhAJIxZrIcmN7fhyRDXbsD9iRV+2HaOeiQL3Y
58Yzi+SRo+ZJfki5mmcj7yq/tEPBeHL20/igdoIjjlOu+yj3VoEV4IL/28jEl46D5fgcar8tKBTt
JrD8A2eZ9CfcvCYZ/EIinMxTi4LTXiFjjiBooi6nIC3mbwWM+9VyBVDFaF9UlFZvlaW8ZMC152Mb
wTLa7WcBEhblM1XVyU/k82CVCndP6VTCymSO2sGbNBThW3HBRLqWbcvNUXAM699SMpZ7F4ZHUMAZ
txNxi4wq5CpVT0o3kBdGxPMXEm6Pzp7gqH0EPU5QlfJT1lOuUuLtsuChrsIQlaoC7LZVb104RWI4
hNXCbGXhCayAbJRfz/Cgz7ef9qqlTwI88bMt4qpbqxvcDw81VdcYYR+saoY5wY1kIyXuFW2AivUB
DyWwWjSXN0RJVQdxBDulTLFE7i0oZ4DBnOYnh3WbO1dC3jAePuz734GrDsPkcebqvMEEIAg6lNCU
TPSkn55s8YcBikvp68zongrfSBS7Fx2Avhwpxz5zO0RllS5fO+cECh25EMQOHo5H26b0dFMtTJRl
Rg8wtjy8a813Es7HDBIDnwx20Hsfkn4gbNKP9aE3h+z+b5lkmAlW6eyTFIBqaq4pyUJP6KL3T4pU
ReWy6WMR89BkRTGl90nfPgcD2SKpe15Hyk57c0qFGPogGP1+PYs2or4hueuzLnlJRVzebExs05jc
lXXVHOOgK+t83Nzp/v/+WTrrIRhVZyoRG2W84IRrJHVGwj36PNWO5/wZQaa8+/ByzLd7Vmw799vE
ot3mtzVjiurOb7QncptJiLM8LJbcto2+JxAdUHfLg4oG16jSXDgRC90s2Ym0Ea6VdONbT3q4tfm6
cgRCxgqvmcLSkRVCEN3KvRVJf2R9IeBFv3DYLs71CqedwkPsw269TIbwHoIHfPg/7IrbjLsLoapA
3a3g/3zVgKbcYFj/aoc1mZJ7CArqqPRtOeTDAfd0/Qe+7uhM9L9WAPRRMlUOoMbpSK1nKAlIQVOO
UYDw+Sm9j5DTsqiENaipGfp4zGFOiKaDghP7fL0OfVUJ2NdyF2/RYN3STEpU0Wm4SeB165mRrH//
Z5IXlH/hl6O+RRgMtigpcojOR4zpB6VSX10Xc/BJ/OdbTE5vB3q8PZRW8kdCFn+Y/QUnbzQIoOw5
HPQnWNUdcUAKgPDvy7nWNNtIcaZn/2B9+7QaJwAwGSNhnQdqqtlqwxqxNDbbtTNOP6gUlBJY1VVV
/y6KP5d8aSJ9RcwtiBp5jtB3foZ+NSUSnWb2vDKfn6QZQa49RC1SyWsuvTOT45MMzUaFCV8Z5pYl
7YijUWUDlprUq8GhmuDVLcBsAnMR2I2Vt7Y5PXdxaFkv1np9njbu0UL3qoJo2wvhCGFH+oX3Kjjn
nH/boHi1guYtRAPwwWs0VPYKUELY+G5R576DlFkrb2clY4Z1Zs/AYu3rhmhXqMsOn6WX2jWVPN0w
k1A3B87+Iw1vaF7FAZaw6A1ZWuQiVANFBpxhcjO+8Z/lyssAceTmm+TyNOS2CdOSzDZDT2YGHvgD
e9GzNcI9XXJ52OM/8oIHmHEintGt+QXZNEwPx5EHPeiNuWSkHNgo6BlrMEZh6dXZDZ1OEOfXPTEV
VF3lbFoZC1TAWKXhv4/OBxLjhKXju1f+QYcyED+CLvrKI3HaDZhNqcp8rUIhr0SPofglsaboouVH
eM9bxdVRAJtU/lEkk2NMP+yVt4h4Le3UlZ8OHvSORHhq5zKqhLntXbMh2wGzeFddQ8wfUsJrxC3k
9FdNNjiHlYq+tyjh5v1N0OmN0Tp9Ue2Mbx7Omhq9pb26Q2GFbuCB6UW2inPo5j6p/k+OZYA+oCnA
uthW4lbiNsjFwro4243tDHJtrgVpztwIDXDbgcCRw77LTTS9cXI3H1lWhVq7SyplmgnLjoi5rumb
DRJtMLqcauE1MWfcKI9xC7km2F8ghv2sMU6BxDSiUTkR8Vu7V75FGgnbXs1ojE3K7mN+94IPaEzV
x9J7++Wj8Fbaxonby+Yop7k/NSBhoRCM3YKl3EiXbDRXri4UEzF74Y9xMguFeN6SbS/Nc/fIXJE4
UP6mX25SePPG86r8n5HtALq3DbqoQgd6wiSDXifRUUeoAD1LaabXDoZU1lstPxxVuyuDrjJy332E
m8Dzp2Lyl8v3fmu5qDFxiFWKLIPqGHFJLwgDyFphZZRtQWG5FB17MPKl6RC8e6aUj2O+9/e1yVdK
zWxw3OQiWCTo4xDi+jRVkn7g7m/J0hz4OvDkCXMHsoirFIv0T7NKC45VDcX3HjWBzG6ZsYA61Lj3
KmLyRMGqvON5Fig8T0fv8P0YbZCk5ap48TI8jmx94pjRzWYoiiaL1EmTElBL9X8cjOXUYsC8kjB3
TUqfRc7mCwR1OvPMgRGaMclGWlqmUcTcs/NXPrkn0Og4bfHvu2QZj7IlOwWQWg9vZzWj7AS+FbHb
9W1hYihFESSge06z7cA3Fevah6ofsiebO35UUmsuvQF6aVL9cVw03c/krRfV+f1XH5jTDfPWwwQN
7QeBkbamEFZaRTV4rkeAbJ8mCSTYWmB3DumworSBwoGP/ZHYGrsTe3dNkOePbFMhgTKd1MnL1Z8n
vHp/5G+JLtG4cN0z3VPPE37UPoluLvokPkwk27VOoIb8VbGLB/QlWuDumSA1G2uEMeol4o6iBIrI
o6zw95PAEZr/27AwkHFvn6mORkvFYpjhyZVCt3+i7InB8scrOCa0jSow+D/cb4d1iyEechS4BWWM
rRuVTwb+R/O821lJyPjB+P+D/h480Fl2iv4DyBfTe4ZXzVj0AUefEj2jsFwKTf8491NMDhNIYe9A
pqOxWiDQ+34KWUWcq12I2nmRpZvVFpi/H9sfRevSinAtnxbHkNzd3e1VIEkLyJMtkt8h+qmsjpqe
1PsZ7eH9/Vnvl2egUjMlpYALaKQ6UKqpzhqmuoPCyKTSrWF0sulqxhRc9Um7UE6UgswPOapoa+2t
J6RRWAWg3MvXbKWlyykh/rqSkB191vT/SbB7uGt6m1VQaTY1nerb7cFha5KiVB+5MRGujq5clF5z
sx4x/0CBznMQIiGA6Yp5U3YQM2gewYYI9sl9L3SAFUpAbbe5N5/0ises7KGSXSPaG5IbOVxpvG3L
DR4R/ZVXvHWQeoOKYw9YkstAbhS4rHtP3bJXzy3MJUyLhOFSwCMywTAxgzQMrXPYCzvzFLnfNcKH
Bz2ygVlCjH/JXb1AneFElMxUBXp8E1D2fmuuchAMBFNTjqFrFswlVugpVnQKsMI0gutK+Z3fXjo3
rLl8ZmsoGCb/V+23zUOQQMAM7qxYeTUBoXmWt0RLR5m9UctiAtsdTg9UHGtDnmPbIiDeIs+9fr8U
x3byxDw+o8O/ivgpwa5w29vx++h0jY2/4XU4sFaUYv5DGQIm5ATkBKK5KmZULM0+65YAzaHkNT6G
4B6FhL7/bzjM2mNLcUXOaqPWrCpE2q6uftkXntDBnv6VxkgIgWZCETVdrtzTIdM0dkcMXaCySa9j
TiXvbAy+l4d6uC2GBxXvKOU85Bc7KDE5wAYWabqrYHC9wZmhR/GxZJP07qYY1hLdNN4ounehW0id
WXUxNzAAgL1KSvRxMEiEbshGEd73mqz6AIpKqAroKoF5jHGctOQqlA2WsmhPw5hAophWkjoSDheH
QcmTl6an+ByuFnq3BC3liD26qk9VVRTtEdCG7KOR06Oz/Ppej03/RRKZHUCFnos0vCvgcG7oadQG
PNv+9J1sGHoUM1WJ6ARIXJ8ZAGdRs7GBnK+Qaeiq5TEsbxdgQWixiusqZZ+PsG0/Sg0kfReCcNqE
d91gY3smvQMw5luMFtT9MdMp4wTPwupO/FIP2LvldC+fMe8EewcfjtcmJFRzX8/c5aBD+ScLywof
0Ojn9lmXe8tb3yhw2M1UE1LmrFYZ8ULcqV2zCXJDwsOG/Bnk16NNdDp6yyBzi9/D3+f0FaWw7uwg
IfYLJyp8mkG6oaycHQad2nZKoHIPMnFYmyoBa60Nd0x2xOUAssKcDhDMPTq/e+Pjbd2xo1fphctK
KVv3Z83CWTp8lO/+OnOJesfX38Y9EJx/8CjOP2wsJwz19LZuPdSRM5C/eo2V3lA04iJtzvkp89Kp
ZoXZz6RD9mCSPSXbT8QJDhSE6ogapwo47drVZsEvOsq0Xx40zEGkQwx6tO0A3c0CjtLcBC9/TxUg
65RKbyG7SPcf90HUxsoevYhi/Q2Vq1id6zYYnEgHW5FJlN6zyANS0qHzmHx6ys8UkYWAK3e2n7UE
nSV9p21bCK2zllO7fvBO1k/B55UaG7QSG+a2RUyxA2OJ5c2hsUjT/pkdU+wRu68N4uckstU9sO5K
whZsm10NwV4FIoAVKz/C2BtRshryiuD+Hj+W7xjmotVI6j95TQsbuxbQGllCOwnFilGEe9TCAx6o
HaToBXW2fFgfjFdbj2P0HhsVcdkAMiZkCf2x8S0K93izfOFiTWyIqjaF6rkOlXfpBvZTFimf2pvK
xT6GKwbyZehhW1ADDCl429p5PkOYPPUvXYYFYAwK7en5rQdT9uUUgprl1EhnUXlxeJ+VUm9XKl16
IN8tVtJ1uwkss8Uab5ZASPsEjXbjON5KVGDRYUXJM2/YbYi+nYJ9owAr3l+6hAZ0t9vNRloGjvzU
LZp+CMPhLfMjXxS+Hae0p8TgbQ15HyluV0AZAO8G4JgWLgwjTI7RQ1gM/sAmjL4rAjdqbVQ2jRkO
hmQxDmNs0vXUaovaY6JYV+1+26fcpyezI4Tiya7Qzzm1RJDrYXcfGyPiS8qr8VMSdNqC56tww7s1
Iy1pu5flIFeFP+xC1R43oMKHALxN332G/TwKYS/EQ8rQXa+GBo32P1IYP5RzgkadYYdjZaBnptVz
D+SLJb6SfF9nYrshQXHjq2euACVjpLkVTsN7Vz6TNj8hb4jl6LqCwyIEh+Q+YPebAjVdLLNLjmFc
VYyrtqbsUX0OjNXJDwSQtUFJUrU82jJikJoZry2lwzho/UKasWK8jSF3mC7lDgR112uIgzWx6Lxe
pNV8fXg7dqtgB2OVrsg/fe41Q/uZK5lt04RpUupyE6aLxOP6qr41aJw0XUW5oAeQASaQgx4mMv57
AWcdSOXW0wCF4E9BLH8IWyFe2R48I2wscBJ2la38Ffy//u+BNYQe1Yk95FQxTcTgmpIVTkwxMKWr
nRZVKVs/Y1nwn+Hjg5F5ob41P8Oe0VOaH/MdQ4P/9NoyamFSX9fJH2A1jxO1+Km9BW3RvYfnu3Y8
Wz9jhGqvtujdCBW8C9wAi/1LVWOMOXFPmMhmoMHVFTZqQFSgYa3NiAcimjfIZAEce0lxs8Syu6qU
THlDiTBacTBTa9T/qeDjDSznfuTIiXwJJHny9oEHsyVu/APFoas9ZuyuxGv4oE9co57t5eYwCSF1
Cz1FNQnCxAYpwhiXoiC8t32gAGpey3DBcs7gH4vv9vAnfY43eeBHPK1CNxJGJMNvzOiXHNNQsojJ
J47duNSbo2MgpFwAFE5L0FOJOAa8LN0ARBgn0Eu1dpA4ElWr/INJWJM3aiDrt4hxM/ynwS+0HyAO
cV8xv7vogHJ7oTuFQzpMsmhEJu+C0x8mA8dKcRQWLohBrB1qWcEgx2UY4EYPFBXXA10Ebxe+1wkw
NLDWlQ3k/1SMYoe+uS4jkBDD95bW2JXKGW+PF5Obvka34wQpklj31L9LHk0gXb6CpZ9jpRBdr4+8
RH8ycfp1N5P1E+JEbXwJZbm2yVX9LePN7Ocm+APe+0XHgTXjYdkClPygon0d5QNVmx9Dh+E+c2iq
70xgrEjxRFl8e7k98PqNNZZPEuf8nMm+W43wyVeps+355R0j4xoRxya+hPq4DW1hHbU9c16kUD1A
xe0RClul2nk8yrODu6n0OEzM00uySmeLJsEL4y3AWftvb0dxEM8ab2UMPZFWQi+HfYowwM0uJVwH
70mPXo8sShpsZqoEXDAVPEX7QXLNpTOykfpPQVL9fscb7X07NTi9GhSwo9+48CNhPkVIzPlw1VjJ
Hk9CXSN8JTnL0/8OgHmcFM24UJwOgqqgoVVQTQyeFmIp43PAVmnEiLCL+FmSL4b7Y4p03a4GqUGV
F0CziCz2FIgilgBKUF3w8T5cBsXEXXEDq7e3d3078hrwHQpwXfYRH62QKlyJzH9ka2z5w/Bj1mU7
qfL3iWSi8gGvqIAE7NieFQCkHSxEQpe3vBU5CS0AZuWOKlGtgymGWMCBF50BMSiesk4cQEidt8ha
kAtv8tLrpf0jYMTlP1RaU+AynSzTMAjRWonj3YFIzK07SFQJcLW+QF4i8rfnOs1SKEwj5ovGrGQo
euiLlyMeJuiXzaxGHdtYwU1IP+8yFQaS1+4lvJy6/HXe/MtUSRzirwdMwl+RS0M2Gc4TriRjGECk
iAKZnl1MZWUfjYrt5BRHxA0QFL9lE+JbbNf/mFSv2SMT5rbO3jsAlMTe3oBgIpoxMmc4uJvpsk5E
Vf8H6opDfH5A8CD31v+iLsHB/4JNkzoOrm5VlnoDdBr40dbbdIOe457G57jge6CnT8JAjBd/p7oT
tnzyPh/LTZ41wJIKwQqIitmHdyzO5kYryoLA9E/F//SqCvi/VjliO14S3ju0aRgSwK+ggsyvg9zx
fy9tEmmSSKYhRuO88gyEkr++W9TvTFtDMy0t/4Cz+t4RXrQH/u4V7Mau9I2NTSziyjQ9QceUsDA4
Jo7tPtHCaP4gC7s1zGU+AW6wll13WrsorSDFDcxaN0SWLLaLV88w9J7C2of29G2bkDt2MweTuyWj
a1brtG6CPaT9xeMraI6JF2Wq7FMzZEKVmvfyKjfxn8oPhO0w0DOa7dFFpCqGoPl8yCpzFQcHZzSM
Niu2jtNUXOh3GsEASfI/tZNp0CkSC77V2Dj2a8sqeiLl2HEtdkcdJ9GORVoK5NOTAOzmR/S4jTh0
Q9lD8xHAMuRjNjNZmiOb3K4FZUKzBgUPU8wHe5ywXEWIXCIOgfg3SMw8LkEpMiOfQ88dazFfeAVk
u6TFPgF81tXnMJFWKdiouWUmMMrpHcxQ55QfuWpXzEhPake4NKta5S0hoCMtNOZ6odyLlCIWrlWC
HAlmZkQF9nSnPf9ZZtKy1NdRSg85YcMT/Hu93dlDPfPN/pFHzu/ujV/48aVHlcP66pTjVukzYrWX
JhBX5dqxNK2ZvODpBq2fmYYHz2CMTuTE6CdJ6azZxxoL8lNwVl2iAGc1rXKkjQMG7KCfo5QooWkG
AdPpTgqvttSzW0URb3Epkei3AFyhQHge9w+MBOPLpyK0hxCjXOEJFGbskeMuW5vPxlxnMP3ihaYz
Qr4CZrItacyp0MY+FynEiUWLoC2ikD3mrKCd7wjROqDvdG/3vEyT1Mpkl23pQZL7K9rCHAH5VtYW
FV8ZXc9usXELF0CUzb5izMiiV0ZqgGR5kSsgD/lLRc1L1aNjTlZBuYUNudxzyBaCi7HHZxwdiPYY
QtU+tjTkBVtTj7X1LXyUvDntSVvBx83U1Gv6i+8SKZu/oGPpOyUGqX59uvDy0NJABLc9MCEKxqBs
a54HgyX7V8ii0m31d5TNG0/bomYZ3qa6wITQ1ca0TWbqGXtQTdI6DICCIw8sm3EJOQwM0/3l1xwg
2/MSwuk23y6Cmp9CZCnWENYpC9//S83F240XjAyyy0dw0HdxyA+5dMqSZ98GrzGYYc9+sXoq+xpT
jMAdNmYIPB7M9/GSYXAvbh9FcEsuavUx3OzsqURlSHbVTNO4egVCvlJ28oCPMw0vnp8fhyLhNfBA
SltIsE3D5Zg+L5pRDFSi6Zgg4IouDCtNvIcQxmaBcGhxNj5TnAvqrFdCqaMqyw0N7d+6grZR/7H7
HtPNhog2OwBbKz9NB7WNLLLmCcvYojErzF0kY1I8moknhTGEJ1dYjGje6teZf1/GxXMtYkPDNr7Y
MZYKxuQU5aNoSaCWp4lqK16Be7Upxo3pCPJDS21h3bReukp4B5fozmfgA2zeBs/FwTbyFl3n2D0j
4v9TDxWr+elzzUJkxn+s2zqDWDoQSMkwmkiD9mJK+kNOZuZR0nrWZsKT+PRMIRBWEGoVKMWNAdzV
DhDWO9wVjtMKBW6X5gOhqRkq+R1Fg0absWXaGtxDMAz3qcD0oqbhYMUZFcPUu9/erEXzp4WAI0Pa
qLUCou1ac/fA0s06tzAEsu65s13q+5j70lVbXQRqU0HXXTq76f/YH2pWeY233Kl4QfnxQ2adpRVi
IkWe+qtOotUP6+JZnQjbSA6F3ex69ej2RYkWzw28IPiDAjxw29zngmIIJxdulcqcl3hOgMRcx7k1
PuEDdi88w9LqN/otyP9FonspoON4BaFYXtqGCh9OEnMMPsCoZoedQF33FgTPc2rEb8LFbcHfOidH
8qVbhSvVWJUHEMe+6rPAd5mfWFo+qKOhilVtk2/4NylSHAGirjiGAIry40aFV4AByeoZSdD0QM8w
B+++mnj0evmuCo3Erm1D3giBk3VAF5hVu+EC0MDXFMc2J70uOaox6chB+YC0znB6YpmWooazFOyE
rjtbTRXw4wdiyVUEwEcQm3BectBeB/eIA0hgqYpVGwvL4HleRSVj0WCtznpGXypwzC4gHD/RveUT
TMzwPRSHXOkvjkxO13K5GXkeFDjwBs8K/VnrkuK2Cl1O4sknjRQlsFtbVHAodDdP6v/osxn6Zvnr
0MpWe7hqZrOn145meLVY83WfY164SISaFiA9LsVxd+tBUUBen9ELin3Of2F3YCMzxJhAxiZKSQwY
CwmF8b5NBWaQexGg2VaTw3cv+0aVysgoHPXEfwDyfx2rprTvribXv36j8y6wR6W1RT362ZljdsBa
YWdieTh8pnbvivqfoNrS+tjr3LdgglsdWQkk2w1RbxEa8rymfo4SoxItApjyjr1tz8MB5ZkJ5bfB
MN65RAHPMr1kWnzU/PcKeRPeJudvtVPVDJ+VAcrzgrE4xxI1IfOleYgW5yQsXwGTSp+SYdyB7XVB
z3D4miApeSsn5Rs6QhuMgIn7ZKX9Y2G3Gx0kcprc+/Z3JGyhFommw92K9w/YiYVB7OQb7YP67h1q
rv6hNrPeGVw8Xh8yUXwBr20HXN5HQfiLtZickXppKf+h1QyGgnsHTwbBVLzbvDycl0UFc2vEj23D
hvoB+QikiO89EARoiw/Cc0aFNMFLfdXwoZ/BROfZxu8sICOjiSCaF1ln+Uh2HX12ObIVxt08R2Ej
vew9RUE1rTJxx+C9JVAVmiwzknaRr2u+U5pMYEfEM7Y8R2/VOaBto/DuKMwgJ9RnyqcYcHz93sft
9An3feYqgjtICg6Ixl1Fgs57xPmBRBp0IkQ49jyU2BKw0Gzqm1OpWQuHs5q8qaJ16RZ5u5MCy9CL
EGNFQbsYKWj5Ik5wx0q9CD86xGI3fLh1QBodqZg57V3skB8v0mr1MZCRqXBBNVLAzLXwpiLKXldV
YZh6q3PMU8SnPHpCRgq3kQUVKkH2b2Jq1C86o401SCIeOZcnCmmEhCnv9JryFxpgqKqGyOIDdDrF
PBYVjOgnk1GNR/q9lk89Qh5CKkorP8+TeOKw9A7DHqQ0S1c/mUtAijN2rgUwzE47UQWgmVrb6BO/
XgLBBaXDJOECUiSGSiHayvTycF2oSV9hWP15UTA9x/XxUgIbUReqL1JG2xVnSnq1KfhVs80xzLxg
xdY718q4MdhQmLrPpmC+ZVdEpJfX90ziHxvy5lDJNrm24MXwV/p5kb64zdvJij0+Yqhr1eJzMheF
34wYaAvw+v++/Zgb2SOfctLbzQ0pV6KU/PtRfHsJsx0lg/qP7daEegQcO0m1N3TqhDBydqCidD32
om5Tu6EN2S5+m2lQXMKEwZDFWrxhQZSxNDloMyT82dfe7O2ZghS11UjHISuiL+b3kJLftM0z/+vy
k13YntChXMckxFM64KF0nFJS8UfgBeCqiSF6HFSPLHWb54yErzKT6JrZw4N1L2RH4l5iO5dlRCVK
4xpUHC0v7pLs2K1bWH6zHoClcdC32VsQoXSXD9auVs61bL/5DIw43YlMs2hnHBBdJOgf1rp7lv+i
yWjyOTp5Alfgp+/IMarlP9KA0XhGYCY3IhkSryKvnhIkfdZ7IvI4BoQMzvNG2go1BtWFSWMXhvwT
E5abS5lkQgaunayqpFiqqONynTShwTUdRUzJaLULGN6rqxYOoi2cDkPUGpFDOpMkrSMM8XFkCUhU
caexDMc2GYMaRJjOwEqBUdUpXpzPUQbk9j1K9Q6KSJgAiDMkYm8XB35TG54AQdRWznJ1E518osLf
jGYKcBGLz3WfPmHFDK8FrhWDuhScLXkdnoYjZP3vnrt7rfYiXg+J6k3SaXQUxsgfBwVJZzw3DSzJ
61Q9/EJ77UBspMTo8Aui3hLQ6A9IyIv2UkNavrFA+G+eXWv3klhAMVxROsS4S6AP+/BisSGOesi+
oBUnU1PG1t+PV5JKOhWssvSJFMlFMWwCGdN2ZjQ7hOzmJ0B0/BzKHxdmwJX1anqtj6jJrzmh7JFg
FiGLMGMSzK+6KHrSrgybao6qchFqLBVJ0ZD8xhqBPpNbnMR7lCyQS2AC8Yo80dv9OsGZgjzKmH5B
JSxekWsE+ye63NFG/8w0dRqyPx3plSvhVm0BtEg7PIpvipZglMrMr/HYnvVh/8168+qsOZbzKsg2
vgOINpiR7tR3SRP07BxROpAPRJ4g5cNl9LFOzpsN2qKY1+0JSeYzCmsExNRM2nwhqFmORIJ+F5rO
ZubinSXfYvQyAhUvwxsBYvwEbeOoOPGrZLIEGk70Ha8cRu2zBtwXcITDs9cJdsCnD9RKkY4V1gMD
G0G7ZNA8bMq+SicDo/hndssX/vERIQ2SSfqbtsdfyrCjPvH2JUiNixAmFyAr3nTXaQqY7pWXxEQt
63Qri9FOPKf3uqU8vjL7mpRD3VjdcrWcb+v+dm7WTG42a2B7NeFR51KejTg5hvzyqcT/o8oVeWTm
1ZoMzuL22AQHKyTgBP/YJpaekQVC6KrLv/Owe4y3l6AAjG5ZIzrAVHY3uotVZwwQtMJoFhObWRYU
NBJHkIDGBaeFYsklay7VdRvq9PRdn5E7ulyXfjVd7nelhhyKoaZzUch2Zh4sOXbyeSLVb6UBlH1v
ml0ed1kkv0sXEh5AUEaKSo36f4+JEWHUI4Mg71CAS/q6V1B/BORoJpOBdwSYAswMWHHOk4yKZXLn
AkOv2CljCZiX1jDSLm3QdHMJbUNEc4XPV361f3eciGkQAWTGA7X/Fgn635oBigCjdMcd4e6Hecw8
31r4dzOaWpOQbsgkBMmit5qUC2yLMXdtiwWan/R9e8516xScMYLU+3Hqh6Z3L8MjMDHrhINFwK5P
/HuqiMX69W9kXDMUIuys+lNZP/Of+0uo5XbS5rUZlD99Fia4qaCAcMMseIKs51uVr0MZYY02i+l4
C6LYBu5DSt9tZh4w59XBbd3R4EUvhwrBCGekcfIKmMtStsaxdIii6CuxcLUsOn5Bcr8y8ZF1tG5h
Ca/LfFU1dWIDax8qmjaP8agQwdPl79nRpABjCw0rxFF7eFTAe7j7o49HsrPYCd8e0spZUyrDirAZ
OLpax/emAGoYjY2t6YPYNVOMW5V1IfuLKyrmAqiCWZHfG+hzY091Ez7elG3AFrkQjFL0yprPJigR
FnuUMSh1G1B3bWWYVxZQO1FSb7AyBNBE2W9Z3C92ScHhcSi9Wp0TKewEQqAH43R5xWkK6REBrGmV
WgZEa9v4MerzpLjLbsAeT/fTjprsZjXu0geng81PojEzsGpV44L6fpc6Fzggi22UsojReJeoFW2F
SIQr+whLxsoeWm4/LMEFJyeSnduFc4LQaUYvNV3IX3Ah2sN+e19aalE8r7Eli3x41umxMsZB/EVn
po5HJgw3lAsHzYaAp1HRaqUqCXFLyubm0J7AclVMtCnIw9eS4JCpwYNeaiGgaINIqGVQeVqqZ6BO
iqyYND/wxhtMHqmg32oQOqO7Ocn3F7+SMrWtJ4zuwdbG2puFx0xW3U5wZaiR3JU9wyCxijs+lklc
6VSTQ7KayPyUr3U8pvR5P8PnwxZGoGkiG4uyDtqAZCDvYPhoGcKkqEgpxN1tbBcCAR/K5X4UZD/B
C42TPUojJCfEQjmo6NYlD+tQ9v8naq5+xxw8uZqF8n5sSSoO2o5ITTV0YNu2vRKbzD3ql9S1fhx6
XYLOWxXLhrDr4D5XwEygG+cJkcE7sDIwDm0SvnUDIUjU6Pp7plDbs1pW0ip4ORlN1CXo34y/XRIg
ISIAZmxMri5jpm2FiZWt1wseUcHWfE//P57WrYORYciAKyl+YpGGPckttuAmd115WV4CnDM4wWhs
56oF3BG6dwvHEzRO4IinVIUaa0TLwUOpEs8uCDpsfIUxyhZmls+pd7wKWPUvQpaOWuF3Q5EICCMh
J9NspMCBH6E+sNDgFKTfYZjuOtfXWHcVOwvpYRlt7Y73ZsbJkdn89rWxbNzKby6ZuS8U/1GdqLJK
xKThlwpolumvSoWMTzOORu8imycBHG3yDCQsg2O+6WrMWMHLtlYDQD/SJB9CT9e7VfoPQ5MqKIma
49FPMI0PlK66ejbAsrUWx0/jc0K12dMTVdwn/W0E5/iLuvyMtS+CIM7rseYLS7xQwuzbpW7REJcU
ruGjLFh7dBqoMNnyZtjRH6iI1ImQHLg/KcyYNdeHVPMmhuAO9nirwzVfHHQD7iUaAbujSIJubsmQ
ShRV565tlz36a2xcFtnPvbktfSxsD6Qym2pwp5zwtFPNLnjWW86YS+Ilp1g8/LCnACjkfVnHesD8
QeIg/g8iai1X6s5YqviIKXDWKJXvwkAWe+6imWYek6oJZ7LOIji2duKGmjnKAlWsbICsYKZOUqPz
wAAXig0Pk52luaX1G5giNa/0XeuVJoK/evfmTyh4nyBoL9FMBvdvjuO3VEqLVjKgfX+WPWIAmk3J
Z9BT2dIYSOb52RYmgQFire4GLNuj9kS5BOmATp0PqOnR9tpGFqiUo13mF741nCvG1OFPdNPR+RXH
5KJ33O/YDW/tZ6EoO3an5TxDOqhETlowg7q1rCoQswBIPTQUQRyTSZJyW46ympFCiIQ1j4FoM65N
8b8FsCOkZRSwo1qlSEGwRKFubxECVyjKdR/5gATUNzKBTj7On/0VSWHLHrUequWVtWXeGOtapI64
JQA8hlBd32IEz7TBAkuGBQQBk+WJhmYo2PT2BqkkSoRneddjArb3KGCmUnVS+DE2QFqyXRc+OE3d
00b1w/LrE/Ew1KKXf8dv6rYFAIZMiIkCWwy/IPlklOX7av433dK279eQIqowZm7Axxt1WeP4VieC
h0F9lBtO4fd/wXzULtRvXIMcrhcD5a9bjsApUbyRaOW2PYRSWPMAeXQRIqSPPfigGENvfYLIT/3k
TpagkZ/V3AwLWMaHljI2W8/iLnEjgR2tkJh1Z8TCA7kBBbdv4JVtzeEijOfH91nECQkK9W6r1FQl
vb2QipB1gYGFIRuNNEYhJOn8FQJeOKHSfzkzgBJfdEmSwblQhn1rTw0/tjpcSw1dTQkenxDd35xE
6Awev3F9x8RbP/1Tqk4VErEO1fRHWEXEydj0/r916Cts8uvy82+jZ9uOFSqRKBZ/tMcvS3l2KerR
o/oUQcL9piF11tNR4a7rzdH2Nb9blYiPgas50zGMSMm1trPZVnfjH+yeDAx0X/639f+qAVV8u7Sc
VPRYzwI1qQDN0cwLZEmcw3zPa34YhYekgBeLrA2Jk8iY0/MNfBjMuivDcVRnqgV/j9e53ZxkWkad
ulgADPoyRlB0hkK4w7s9RbCQD4KEXyasArvVAfXPDdvvA1apqp32NF3mr/TVZGZa3IkQ7QTVxkT+
w4D/Yp7Ww6KcngLVZivAPAqi/W5Aug1kfAd5FahgxpdGAIdhQcSJjHIwds9LoVyBZ1Za5Q3uMyul
RuWZmE56ZCyDJze1Hdn7/kL5AHjWJxxAYhM2d8D+7sDSlWUIgp3iTyS0XDJTLjYo3nldYLZYkW37
53K5pTYtrYjleSDiCfTbPeaA2giyUvUTtQeqgDXdQauzYe4XBnxpTJlQyL+q0BtyF2/GNGgQXo/0
llPxqNe857O+x4Z5RsGcW9HGbJWktotNZ1bmSTUgV+3IZKoaWJRHsSnVC0Znng7JDZR6gsD5XtT2
BsC6vYlsCyfn062wWGiE+R/YIVAElqJ0y4d6blkCRCJMBhs3B/mNDxVM6PVpZhJxHAQerom7kdoS
U1dMMNGkYx7JbqOib4l+i5ygf40+WS1p4yjJ6oANtjjqtZ5Pv6iMWN21OZHWuHj2IDQCzMNw7PBm
ha9fNczSDcm567Ucu4zD/nCRdTIRaXdQO7huXxp7MlN58pADgYJE148bbmjkPKvDSh4JM9J8usT8
+mm6xdj3cMx7S+2/IIdwWSBZAXYPT6I4tseVu4jtsgnUk+z0bhSspHeUZFFV8GJ0M9YzVlUGxDMk
RPd10XSYrjDvgTKvvbk0UuImOL+DwF2bZu0qCXchPeeaP4QdZ8r9QGWRKGdzOJLxR25aYHWJjczp
peKyjyDLtuGs14alygRTq/23kjeny/6V7bpKsVr1MHapzhPtuo2y4XHWKpJ5M3voP83Ocn2C6kKg
9Bgfz5y534NOlVqggu8dTJWiCbF4OI+oX2nMmyzC2hIpcOjOdWNDXsxCU1wKWWB8noM1BhD7SMDc
sQR3Uy1cLhZ0wa6u5FZrCWGNyzl0J5qPqMfRojy1Pp4/chpxRQ3fR2TWf+EpdCxQiWUStvGUhjaF
41s+b/Lxq5nOA1BHIwHXBlCYVIyDaM/gWOkt92e8UYd60oWsikQWWLDGQl9QYG+B0HsCgA0v4UIy
gT59OLTVx2CTmf3PolFixYQZSsMlJzcDb6sLlZkoHvglS13Mj16jMAvboalgNa41PXbWtUDxggcy
fR/MslTfLBy7aus+HOD0LDlPaJtT9hFFMa2BZd6nILquP+KWA81rqYryPx0uLZGcinaOL9MukocY
cEk5K+tgIDNgEKZyLRb84ZNeGnOhRcne/ZUWuHhcbviXZZ7gVn3qWwIenEqKQuvySqR/KpK7bl93
0Y91ig/d+F7qmmJR5K4/VvJFVXYK20PS9dtJKN5hU92jVqgBiBIKBUZGNg8nRE2eO8fwUNeebehE
oJWoFzFjHUwzgDy8p2+WsOxGT6ISOhjdqcw58ori1kYI2+UXX+ZwTt443fEYfEpPnqnK4f4/fHzA
lrgGHnsKPCpGXPBrMR47Of8J1hA2Sk4RjLEfBRfFsfd3Ppzdrc+tuRrw/15xMUbEmEPBjAmEOFVw
LqL1FpAv+3AilUYieiXwBOFq7QYopoVJz6o06+RLXSgjBaGz+DUNpvTbl052pURoL1ec0W+YEiKd
TNhr6hqpDlZpHKT8v0C34PH/g7U4Nvk1XiYPoe0ShmjEYn3T/kOXCS7v06Sl8WJ0U+ete5rmDEuB
egyYwd/ZZ2FW2SE8bL0ENCdEGdBroQAXAx6uUJPItTb4iB9gMjlGAlxYFg1qPuTy5efa6ymeBt2Y
ZTR4NJZrYsUk4QQaFQ+jH5PAPx7oSHv7hDMRdjO2NJM79BLjScj8IISRvnKWuzcZsVnpjXKXPL9a
M+13zvU+jAzN2xliZaJffz81oVIWOWEir3tPICksLX95tBAN9N0aIjAU3kdWNrk7s3QtZdcuCRcm
6pCRyZ7wyEdZxdkx5czvJ7HDwsHLKeIPLAEBppc4RRIZ9GMQvdbVl3HgJuJzS1mCz8gSe+A7IMTc
o5SSh97sAWdk6mpEdKssH9VrAAp1ffCO1J7i0V+pcW+R/DsqLgLPy36ToOGEXwbpZjF18DKUcZ1J
TbE0S89uMUGMaw/R4M37IOfT61yHX518hlb++pwzKleDQJe/Cf93ALUkJBGOsIUZac82GMPWJlFp
iKIZiq1CON3xwcWPt00R/qdhKpzvIM0pj30flHDTB93stYd46vh0UjK3i4PQ/0q46xMGfuphT1Zz
HROhEpGxp6f7ZP1wKVQWr0mglOJuxmY97EdvWO3Y3U1R53MroIqhxT3MMr9zhuMb2KNG41hrWqGq
o87QibVnxjuZcjisZSPY1/XBOv/KVgm0bME9TQm6JbB59Xi41AA2gihidC404tJ6mD6nOzrrDmmn
hxx/+8Mw7jmOKmqJuZfmVzmUpzoUfwIIwM08qN7RRggfRVPt97l5gH2mfUKgmpzXbC81GH8UXTp9
A3bBDx9lzwycuL5sHveiJHN63DVSi48InHxD5tewV2yaDyqwySgrjnhZBh2ccTJ06Js/r3TX9Hrc
//ONY6OaFD4ggKZqWkeOodNL9/Gs42I9vC2hPTrPl0zwCSNRnyxpxA+VNf2ao+8m02bcbbjBuT7/
Mzx/V4RUBTPVQPk6wpCQ5AHVaXOvSJEFpHoxpOcM4Ms0LzkuOL8YO+I6l2JWZjqk/f5CpNCZdN0O
uN1U+xvU+Oq3umFnXHqYp1QsdPE6FgVehZCqX6KydVTmabDMLLyI7x+2hLKIrNz1uz86l4ieEbaB
qpqs7bvHjs34bdyxBgVoCO36G6vqvsNH2P7zY4gNEOCSvaQpCzjvBgXZ1CglNa+CqK9i5iE+04Hu
CArK+AM3ERKCKM+T2gEK/g4cMae364+40b21alRVA/1sfPCzLnqIkKVpcNv/RWgZl3+Ipgn/qeMY
3GJLSVWDieKStBsxSa58o7MYPrJ7zLPvQTJQ1zjyQ5vPGRUvbjkmqLP9SRdnxYbYDyTjMLx1lUeu
KyLRJ/teonJAnmqdK37N0fGBE9TZKlbdbP+SkEbXf1pyj+IYkPc5+SehmLogkOIfahiZlrRgESaB
YgeXxlKYOm3s7RJBlye2fALlsEwRloQOmPsEtYY7bI9Hv/GbkTOP4hpnfpHkjIiqXybXyECzwRx8
ROGHGRiWhRpofFB2DFH/Cb4THt7UeqLzq+gvjMGpgBsuhm0DXV/OkCleoUMDYA8xFhoKQ3LFmsYD
P/dkWgXQ7efGKb+vAGZ71vKfb/M4TPRZvJLjpC9JgleKhW4+woIw/mmfO2V6QZ9OEI8PSXyR4nK8
XSVM+CuUtKolM3sW8rFiTzLAsFZR063ohHDFvJ8lazeCynMWzi4nHPAgvl8EGrdgziFnJHRS2mN6
A/EDzFL4YCz1/+BnMtROp5Tx5lE34t3osDndvgOXQQqZ+95M5IfGL1bJxiOw5apegDBv00DyCo1H
aCVabz2lm7O4a+ik966R/h8UnRjiunnO1O6sEBLNTQc4Qlkt5Sn3yN47Rq+kNKzyK/CfaLsf92YN
DMi6JUBkJQRRPYdVXFGjDv5MRCnfXY40HQQK+eUzJpFiE+tsHqMWYY/YqV7/4dhHXxRwQVisiOyz
q1dqzmPFEXKAGSN88Y9NVfwqNhzNZAZjxnL6MVvcLDYoOZxegCDM2C5gmv+OfUm4Vtu6ZpNqQgXI
aLzC+1CvBStIZ0Zrs70awQ46FrdXlJtGnJnJ1mNWb5meKfyxxx+CEoRM44WJBzaTg6xfU2AD5iQW
q8OYt1mgSUEVHXyCVLsFkTJnG/G28V9zlB5YI3xtCqXi8Be9cjaIkPaUbyKAUpjURuVfHFoug9hU
BWV2LtPZ/hrsRl2hieOcG3wnBYPWth3XnmLptNE/RxkN9InzxDJvEbY65aIan6JsIRJnprc84327
9tX5M3UWPi5BqeDRMAdglzGavSXvxr6uo2Ef8OSAhzx9Bcmck8ON7E972W8JSMpsA2gKHDZ+Ss4S
UnwKhZdOuXidAKxv1w2xgVP52ky1ZTSyfAyEZoho3AeEeBt9Q+y96BIo+GfS3DU9dUwHTaic6qdc
TS6H/nitbKUiZ1/4eF2JIcMgYzHQ9whhlEBIB3OGLIDh6SVhYxPOWFg1QX9QnI8TDAlqVIR+C9pQ
GEZyGJnioyp2YWDvxjN/XHmnx9sPQpHCZhKJUoKfMMDS/XjakG3uxHnwtX93QcoOrA6e4C4tAZpl
3xs1ZlWghw+bInCM47RqFvXDxIKIx0slovBol2Q1Jn9RoFuKyRqjWM+CfCSCRmW3hQvk1JH7Yzra
EqMTmR05eoSn2nCUzp65BbDW9pK7LQpwoG2YtutICFy8Rwi4KiAXU3hfhtfbaN1IQ2Rxuc4z1rvt
UCWyzNSjHD8G8RD2GVviut/SbF0Ir1MNC57E4rkAKiLirnwKkhikkOCT3qqYnyByZTdBpYm3RZrV
VHHRW/ye8U1PEjWwVCWbrQi4y+L/SxRp4IJNTJSqOrfNc4dEQR2IBJXejurDrlh01brwo2Tgkkac
uvybwzzaUhspf4hdYzSPk/Un2Bis7pD/NeH6kU6MTBzKQtoQm6RUl5esIKpYzzBmwAfyfshjeoo/
FPj1oIfqtCLcaEWVllRbxpvd8JTKFWlg4K9psTZhBuPlLzjR1tlbseXYjXQeo2iGFa9CIbBq3kzK
dDJW9l8qrt02wwysqeTaTv8i/1iiNGRcTTwXVguYzDd6djJwE5WPmEplfgZHOmjm3yEKjOvEQkhh
/G+49/1cuU8BPBLMUUR5SOZx63ZdZ5nKPVR89XQX2zwvGdZaH0Zw2TchVP0zXVAKDtQ24HDZOEl7
GwGEZxBZSLHEER4Gj6zrxfzkSHYSWzNWa/NzAas44SE/Txc2SAjsRZwNx5USC7+7gKJ9OgabYNy4
aY8/dmjce20+ZtbuNJAjh8I0SrQNVowKdLHset0jZD7HT3PqFBTTacYo0f332fyVBzRyQgFdOKXm
+fho7JKiG3ooDXhpbzU0IBfQDf2qB0tKqBLz5x6sLoeyrj+j3RpslStNUEyWWYoxbLj+htmjXVqR
eEWulGFt3IXcmP2R0ZMQGdKGoHGd8TpZVDkYhh4/I8Qf5rM1RhoE0rjhSFNO3bl0Ll2y+gDWuDfK
oNymStZZ3wjDcoHDUbYkvDusc/KoXqfoyCl56pkichVxTOCqL9jFPZ+Ywi+F7uK8Fer6A2F0Fy+n
kxcKkXu6H3dxBQ5Jf69ZhSTD7Pr9G9CRBuKcwHyJjZyINost9xGuKc7diA+Gj4AJweTMZaGVvQm/
12pz76iSzCOvqgMvpLSjNnK8ajjPQ92nskdkaLEw/2wjt36HxnXZ+krSy3SOgHo1uGBN/QjZU1RN
OAkpOGg8+TE4bLJa9ahS20pHn+wvY/VMSamWVXiR/fAoSWkvULx5YCUbzERXiLbPHeCTv1u23aik
pDdIsAieoXNkkgS3Hjl48QxM/Donp+yb22IL0dpAI6gszk4+jmzka158XARFY0UG175MRDbaRzFA
sMfZT6ncD1UJR9dkTunEEgyPm0U4akmJxQ09E4pQeGppRrIGlrRhy1Q6st9AmmJHPmc02to9VGkR
IXJr3sL2Bl/COqG6wMvrli22sYheylPinXWTy0ES1YLF/SM7UP7Igk2rxzmYDqR+j/FcbNy86tqL
vlvNEsNv1nbewKyYITfCXOYnSbP7ChdlgsY0iTEvT7xVTfVQNBgLtpT5ke4CzgnwkQ4Q2z3KEmU9
XZYlMOmpMPhphTdS0kYod1NVJCr1KsoCbsiI2b5hidWghsc2GCTV9DnpUCyd8ACvT05af0CQ8ph7
iMnasNsskZpoLkx2MapWPi2xFV2svb7+B1PVCRsiY76R9FUPvuHO4BLkZ55q56g13rEnEKvOWtMd
g7lZ2krM5xS4InnPjg/jpn8NEwI3VAIV1k307oFzqBTNERCU6y+aInLGnmtX+nQ3Or4/UJ7cmzdU
dc5wS7UsefLhDGvTSktTaDRkFboDQANwxIF24fGVyO9zymqzrqGsn84vgj6WfuuCYsdMRykkIg5+
vGmQAW+/zb9Cbd1wBIHpEiojvR4aO36NctKosWbv71lRgcwNkFfzTyBRWkjUvyayPWDvd+yxdGVG
G9yaON2182ZL0dKq0llnE2BD+Qko05a5PX2O2hfj59dd5bK6SqR4XvCwU9O0IuHI7OWd9Ax+ivV2
B8RmqroQpPVkv+/xX0O7ruo2sSGosXrBjTdIjirt/l0kyPimt3WHg0gLZie8xXakEQYmSMWk4r9t
L+9n4MbS00Xcp6OpAcG0mi1Aa962WLcCd3O0Kzr2iEbYJqQkYjWHmXFc7G8yvBWvS56lR2WKYsAz
BM0tZnWpWln8k2/mw12XzW5jeY1DHQjxNLL6k/E9HdBRANl2dhAQQnlf8GB4ozrfsvLjwQI4HzQ2
fzco4wT1GJrOGjBU/rLsj/5NF6ppNSg+YEObfxZjGkDSJLO+t0khZ3qpYdxu+hgjGpRLoXIJVri3
q+gPOp1SIpqJ6PP/uoVonBIiOs/8zKoNgRP/fL3T10b+/3JZEQ9cW5kkuiGGbb4NMH1PdX8KAi8v
qr1ocjJeTmciwlV+FoslBFfNWupTqf79LGAUDP2FuExk6Ea5Xihk540v9jD9RDrsDzRhYGkmfeyS
nWU5kpmLPr8NgurrgtehiMrOJId/5mzRP9Yd693xqBi8XJKxrZt3f7kFWB/mudWzEbtZYAkovWfs
aW7ImFbCwvK329Wq/j4FRZ3OxUQfBfGmnc/xa3dWtxNApsGiadaF1DZjGfSF5rqPTxGvgjfHV0wa
DesfiOs0BxGXa5kdygyw2QoSTJKO0fmVeO/BU6xcO3zEPwZhsk0JfWPwKXdK5fUkaCFtcd3ty0Z8
9FEkoiJPhXMSmPigDhTCnp/Eg7AXJ1IoyxgEQG2ha2xny3JQrHcpv0brfLr5q/W8CQLVJErZ8KPD
nwVLjKYiHiwa4YY2viY4kNt6/hJ5W89F7qzGcvdm5B7Hu7w+gzhqQczWSZjgRV5J+JboaLcYgQWE
34lFwXezGurMvAsPNOL5vxHiIcF4uFWAQQJXPCu8efXEXEmOOwMt1/uwAD9hFuSts1n7XqZTvckB
yjeEvrQhQjupA/9ZSavQe3CLnjzF7y6eZTliGf5NdMxWU5GZ3pvIQE3sUZmkzWrpyjwLf6fte+nr
6al+GQ1p1Yu/kWp5X0ZJS11jrgo9J7dypoqv52FcSVqg3kjjchpGc+hh5nFyTUOueuHdWNFy947N
58jXRPFkegJnIS91wyjbUzOLU8qWvx5iPjdA4mOf8BHveTMCkgBKkR/h6mQSdI8rcYoz657LPl9W
dDE9GB4auJNQfnIn5HRsvf9p+U4IcFFGYf30cVDZR42suB1kqKk4B5T7xuk88EvrH0cNmiogEU3U
xYAtfqsDfeYn5dMb/UoIue3YGkf4GYaDDLwmDiGk6Z8JEW2RdzoGoN0bG+5CzrR0fLCh8KwrvG9H
QtWIY/ZqiprGx3u2yz9QIYbJj3HpRY0M+SZZkUhY6rn+lkp3OF57KT/Nq/ayBKDkmMR36Dk5A3dt
ZOgRlI+RufzbuAxcV5dZlWrQh5oiqJS5c6n5ql6nalHdVvsV7e3END6QSlfVV2duQ7GVmOLWpZ0/
jApA+xUsxS4IQ+/DaQu+k7eYloLbQ6ff8juNRi8H+ldGsNd/aFukJm7F22fa1tbCdFYDRnRCrT6n
uKz+mSpyt9uGO8DS4nBogSTti4wssKfWwKZ/Ze8NnqcLy5lYvhzSuPR/4FEG0UlAsvrki9cIx9cH
BqpqZzStw/PjmuanuTA8+I7/rCFgyYdCzJViRDPRxYZDAB3gCkZKvhSzrGBJcqDIWFdqccaL4KRj
WEyXQP0lnK1uy6o2cXrnD7SvSamnJJdzU8QGRrnovSCHzc87tiS8u9QfDhHznbI7q4ORCteLSDYl
qHnm3leQO/jFKU+qt8ZL4OxE5H0TuRUygMyrk9TwfRsOvBVxx9mfA552L6lbOOC6flkCP2u/qoaG
B1leiqbKW+vAH5W3fBRUbkaoj1+fuuxVMDKEri9XpWZ84PB3EqeU17O6UGDV0ck/6D+uDxtq3c+A
4T7ItreIOHticdVfG5iOSe6Si6S8eJfDGnM06QDa3RexlatpJVydr8GXfJBl9ZWJpryfnzX/8yMg
vA1AFG5RsAY4404gx9LhmIThUu/f+lSxt+StYAOtGQpRy26kbcen+Y2DFMtcGq5v1zYa7URcAePu
2eecoI6w4OAqaghbjZhbgIadPyA5eyifxNuh5G+ZNkLU8zxpPYrEL7fOv7VVytpOw2y23i6cfXeZ
X76+b850O2yag+4MRq1Uq7GHW6Ji8WyFjbX0BBfFQdxFc6ygt4aZQ3AmxbZaGsikwkG1khHE2Ks0
Y1kCf52zdDcuFXRLY8V4e5u/z3n2cIwdz1xJX3wEnmFhxQrxz7D3o1UrtVlHu70J6ZSHWuf/GkRc
IdgeovBJmP98QwgKGttq5XJ0NJ1kiB3BRanvsFK6b7HydZXpRKC9DgwIPfuLGb3CfndZjZOcWK2y
dcy6kfMsu/IBM61wlMwYLyhOr8IrIPZwzrZpBas6hVqlhXzmHZ79vT+/+fLYP5i99bDyFvTnVwKl
RdiC8swUjoSw5rANPo9QFgd9wio5YfFo0QKUv6UK30gTIZixfRF7qdWkyC3LUA3YH7vPXKwHmmKU
XTmwxpvrTBbJN/IWiv3El6SY07d2tQr5VqALQTYU/6IB1eW5NcZu8pqwY/+2TjMNVFjwmwlVG9E8
6KYAMgsFPUIhgkmtxag6bGvdreyKc8vftLs3FyVuWGzrc2MXqbi1UMuXF+rSlffFuY1BTZfM1s+G
zl5TUlfgBRBBw9Kzkizw0FmQFE0gdpFfFwgsuuLLZp3BSn8RA/inkMkaicK98ZSN9juDfKJCDy+g
KbKQGEKMVU20D0v0NZ54c0dwZrkW4k5lbfzxhZYl/Ets27VJWYxlsd3vBGdGwyLMn7/3eaKyR9Ud
vUI8qezDi3SmhK+xFeF/z0faGaIMNFCeRtZ8cxYA7C2qEZOBjmBof477j/Q3B9J9EH/cDPgZtRnb
oo6ScUEJGQDvBl8HpwVcNdOBJlcxlcRcG7KpiF6VboTz90IDGbmKd2vkDMbuiEREqgi3S54FDl1Q
ImhYU8p2OSeVfIJVbMXvS/0WofpM6CA3dv5rYL08HgunfhCdi35/bEUFf9kOXdu1+NrmLUiHpkKi
3KRTHEo9XXMbS2l32DzO9jHSXscjA+QLq6YMa+gf0c17PpyjIhTQy2hNySzwPwqt6Orm0cTCd0Zn
CLvsMSgzCgxzq5bBxqQShbfTH0N/vdSdniFv20T2jwX4n0vKSivXOuyzbxQ9ca+i/WUg1Kb/HoWs
21mqbFN1vVfWvmQo5GTklN35ivnMpl5B9hx9XhoVWnLei4XbF2+LCdSssTMA2xusakCZBXUqa/rf
79wzMI5jfY3guhhJxMReUgcjUH3P+rHZcqSDEIJ5M8GO9JkOEiOzlyan/Eu1uYKpu2H+lyOJdBCb
iw8VpAFA5FADbpxZXyx9LDhCDD+gHKssWfM/5E2pvWDz1WtfA/IfIuefo3APzKLq4xlfpyWulDIm
Nw5jLu6WD7e3OJMVDvj9MgCMU24eXYWlPzk2/DQS5rZ5JbKlezpvqP+7pX41yD9N6LJDgkpIwkf6
ZARCbU8lqoL3TdA8ZA19AcBuo0cslWWUMfaQI6aITb3PdFbFM9rqrrsXfO1wjZZ1nKyFe6DUrpJF
5Hmmpzj+7x65tMx1YYTWKy2WlqP8bpMQ7Xn6h9b822reILLw2f8Vr5cPd188BryfWp82pIJbRgep
CyWJW1f4d/CPh8HTEXhim33U76wDJ8YmNwvcipzHZSKZjPoyQ/IXrBojJ9F4bvaN6NcQWesMsIyu
yjjEDG2H3WK8xF5FGaN2Dlh4RPB8vfnNccKJkhqLRLc7ZAqCycZE/DRCM+M87qqh2AyrrTuEUnVG
s+zaM1aFuEqykTFqnMhCqFCWIXfuNp5M6MaFFBz4aGfY3RBsb6THyB3DQmLUYEUtH3iwDdIOZGp0
obVqvw1otVY6eMN4NnnQfhYaZmz+l8w3BbhlxY+XD/EvgyULwj9ZLqYz5fdcw7iJIaAXStx8X3Dp
XL/f60NmYiaVs/BkPGfaDAt3DcJ61cjX8FHE453N6//Jzy5d0FRr25UFfYH3VV9tJ1Du26MPNS/S
VUuv7JyIHun1JhXiwj/kpgIoyGfrtI4BvEsM3jxgbdljd7deHqAdqb2DSvGIF5fschUnDFFgrQsl
KyZDE7ghggSM+nvAdTLtAWKHgmWzE8aTMo1B4srZ7Fld1rp6urL91QW3IzhRI6KzHMi8lXwGyUUD
9vpnVBYa8Bs+6HlrFADR7Ergy1SI4asEi3BcEzwSskHSwV/zzJ2xMVxK3Vph8T70GtC60g44tx/u
RI1PsLzTy3oBAXZA420zDS3bvavyH+g6WYkOkIyUaIP5jNTMUOKN6jPeK0AAJzaoNUvNRf8zG8ty
5YuULymiwxE6GVH67hQKyFaXcl9U+ClgHafOErW1hmCYnINP76943gxJRjXfVtu+AtEMiPtpeR0w
ToJSdFzJjvZ108Wydwo53X/JCW9Tt/GdgT5GYdSF8DGarvzL3Fpd/yJBVEqPrja/tlecYAXqwJBn
on4RIJSxW5qEyBxYPzLkl0f/8QJfAMvXNjz36kOj+o7nroVD0E14FhxpWYwHZ+qfE7/M6+PesIfk
0EH9+e9dYv9E0IyIOqIMZM4tn5OybMuid2AhubP1abe8RmNOU/sIdvNZtVZT9lgF1Xn1yrjyE4aV
OuO6m0+4VBZLTLCUVjuGbyVG5J0W8D+rzvCGIWs/AwtPo/9tv3aei07yHpkt2Xj3S2a5aVU09/BL
rC6Ql6QshMqkTvYHjVyacZOPrjekZW7zqusb+dU58DrU/9CEfbBqrVk54O5CVRJxFizRdvhASgEV
adukKzdlptZnNVmhiRFgvFbzLvafgsE6Jb8q1QqSkvyLM39QAv6XWG64cX2UCA3JhZ7+CRwHatbx
exdGVgZbLF/2OxEQ5tLiWl7JJPzs8oK8LIl6W8kcTv8V2vipC8E5entjTtEW5yVPuHnqJhDZtAtO
2PfQBJZu+Edpp+Pqt93bpdP40+VGpMGcmSH/FiHk6c5VsxZV1aDfUsIUTrFdRvKbM8A71+B8WVyk
ec21rffj9ZAXIUzYGPSSMmQUjdl/GGFKr42tL/cw5eHm814PW04gQg0uWyeR72Cs96bW8Jja5oSa
Jy2A2DxeYlvC31FTKMC9/QxJmZC4UVkJ4Q9tpKgOE1cEuiKucdtbmTRgYEZq7LtnF1/2M9MvrEI4
l0ggjSc9AO4YZqC4DKTPF9VfHhMqs435ZlF0enzWw2xJTTiKZHGdydewnXQOC8dmIB7e5m+9dJvX
3n9Y0owf+/tOTpqvUBSyO9JmNAyv5f6+m3H327F1chChSm/Ry99/taKsL0CrNSsX++grTBGdX0Gd
7hvYSOmjdQ13TOroJN9zaZWLtP67XH87H+g4+3hIYQeZnJitlv92Fv7QBTjBwt2LP98cPTajsZZi
AOCrJlWtEsscm9rIdfmwvN2w4TPXFpMSC/nQeisMToKZOgtLupVKUzSAix6UHvhfoG8a8BITEqqV
mjokhS+WmppGmKsUTlh1kwwpJ9HAt4WQ9v5G1V9ZLsR8dDPjrfKnoHIAqhFSRmhCFhcezxzlxv/H
XYI3WKtqs1MdZwihyZFo2gz9Msj8V3/wrEdnfu0nRDkrxwB5p1JZPNVSHmj3LylhsMg30CICDTBz
HmKuiAConIjcd1LrihRmja5BJQWS1cqEN47XVvTB7AIhE8IVFAorxmsuisUDMVqW3bun1yt6bCJF
J21du06miEyJ+J3tkG7zCjgDW+h5mAmCw666wesH9IfZlJQ0tK2wN6RXkU3dpXrkiHQYU1ISLjsn
1EQNxBdHDimgST2RpXlk/nBGJlBdxeX5eWS5LvsOGgDcoNNylKSAYV6lnrrbN/OXDzQXMfJ/ijXf
nJ35CVFdXX72ulHS98uUJ5epMsoU7VPyLhlHBLsES4XDYDCxkmfjCbxt/N3cQo81j8g4p/Lyx0c9
+LQ2nnddPms+iAgzdJN9zrXn5BHYoBk7pfNCCu5OIcYP81W/KrAcXQ8rHgy/Jht7PN2Imd5xwEIz
O7afchnK/YIvJrYTeU+2hzxZBBEIn3rZp91fS/yOi7JZ7BfNIKWO5SRkiy2myvgMDO0z78inBLjt
gaFauz6DAGxZSZCCjqNTvMjwN19i9OkLpVRSDngAsx+Mby07te4jA8f43DNNV9cIPGkn9uWPfiS5
dBBHPoAg+feWWmGMtG/F9rVm7f+PzpBmjh7LAuhF0lUX+9dslJENMwWvZuZBACmtrRvDeWGpKt3h
RItvJaucEVbNX5MhcZRUP+uOgWfpVULRFDFc/aMk4YZaSsZy3L5ALwGFlqd6aqIo4EFk3iKXgB+1
02Z5kmRx19hB69br69acq/pc3yZ2xKVCs4+c4Fr9cxbkr3BbBxkcQ9plv0OkBvoLv+AqVblyzyiY
cHvQjDpVrEcCNOXZcENho/jXDAIYs/kW09CPTzT0HnUEOnyGKgtk6TeGt8vuLTxBjReTDQyfYqO7
R+INO46zLwnulWedGcrqgizOJxIyEUbuUDKZWGPfsvqaouQQbKrNqRA0YPwGRz/P16D+SKq4ucX7
zPv4j3ic7TKaNetPULsJ+wLtRlw8yHuntdqrIw0Rz4jqlmjLMRwjdkB6W7QrnwUaHaWf3D+Vn2wd
cQFQlYYfv2px2wkpuk9zQ2o5znfSsRzDaiVVAw6d6xWxKYUf1UBVb2uOoGt7b7VwoU4rPzW/7ZWS
Xxk2F9UC3G8mbC8F8GQBSoQRrotIdKCmXT9iZwLnxo54PyZfNP3rhbX6uslCZ4QBzAsttjB/KSxz
JU6ULlDIHDO3bE0DqS2NfX22slL9f0lKIJqVMPxvBYgCcyw7nw/tyf+Mn5o4O1E/Xfy7VdQFNdm9
UURaYYUB6qmPHfPDZP/hvIjBMdsU1T/43xl46jESkBILDi5CZKFv9mVY1LjZvYKiePZ9KDS0BlyV
1Bw1Ru7WT1wgLt9OOgVK9/KqoEX1RC++OA5YKqsPoJU6xmOrn3pacgRyo74ZWVT7fWaHE3MSvwZk
AfmilWEpqEJpDgkc4wbY3XFqATgZkPkM/vwOjAylAtb9Onz97YcTN8371tbrKvdfwzk4c2JrCcsR
xPXZwwQEQI0+xbfMutO5Cu3a2yJqNMSA7xIlwrYEHS5RUEgHnyoxel/NyyP3h7+K4cCRN8jkV7uR
jsviHLYTbsRurUGwJ0kkSVhNZhkI2vRseb3JqVlFNe/+FKUlkhAMT3OnGXNpqYa4XdHCiIna/LRX
eVhBollWzbhxKPJk688OP5BAJG6tUA0Uv0yupD5hZtWcHFoecbzoIDFMcFWhNoWDEJOxrWpLlKmo
lvS37FrixCKejwzlktyZMU5g6xJ6SXt6kWzOJDJul1ScvQLY+zyMQsoT36XSistnpAOkZQEwOGLK
x0ZlKW29FExzIDoAYJYY+RSKR4OAG13D7/UXZwDm4K2y3zgH/FLCKRQnHBMFcoukBDhnb71x5cTF
e9K663WWSLxb9Agt0DJdQ6Q42pPEOLnkMgVXXqxEV1dgDuBQuZFu7mVb2VBZq/IwteuzXQYv4VD/
UP6tGf8n5IxocQt5pgQ4QOOUxJLlbHx/0Y3wsuTlJ6h5tMxt125P2kz5H6DbIfIc5kKfZ1K++iay
YOvaZl6ybghoP384SmK82u6kTw585laIjwqM0OSWhlztocXVuRhdaDGi9+wuQqcP3ahOXJeIz1f8
kINzVtggemya7P2iSRhJiLKzcwhbWx+hbRAUdo3KYdICe8LRe786rRE4oUmJptVxKY7dlX/ikiJh
/KH2QxokWsCBTpZnTDBblr917YAawG69nzDG69DOULGde/mBqCZ9nGVgacFf1+fpco0Tq49BcYD3
V8U1Wsexuj6PW0QDIr491AvUK7PkgS3jKq7SfaSKdexM+SaNIWSyYcOxoCGCajH5obq3gPCvbxx+
+XeMELbb+aeBYQINCDkAF+pgbYZJSLTYVvNDvj1+4CiXa+ExwQVzKqGa//RV8vFDuZ41iuwWb/0c
vY/GwPix4GQ+eUg3HwOMLpswEsfXJp5vujHtY8oT2CLnRq1tCCYbaX4cVHGMHqCahYgNhRW9G3fn
zbh/PdfSQSGWyn9R+DkICSgVQyWdo/O1WiBnlzZa0l8JJxAqBffaoDsw8tkUGURf/RDpgh4ZHIoV
hmQqi6tZqAQery8uk+ZdKIpsrmnYy76STTKFsCevmpY78hBLM5hNdIXOrjH3YZs44V8lCUcqWLF0
VKPvANmpoNRug0b+DAte/onfoDqpXiMaVhY0CXz1TKnMu4LH1A59efxGbOMtRUxGngJgCvIgoW2M
cTKfdNpK1a1IPLCJq2km13WATP/N01vwwuEd0UwQnIXYl6Kk6uKCNRBr9LBLuQjwoUTGQ6Od+/Gi
hWVHoWKwtdcbBV8Gn6fT3lYt9xtsQ5LcCEGMECw92TvbiCZsjsEQaTnH5UfeV1gCx0bbVCdB/ZOC
DHxXhSx35u2hWE+4y+kqwN7BEtXRuJZuJFs09mT3mKAlaqWwXbuGSSuwVNR5gJ5+4VOsqyf2Kbre
oY2DF1i6tv0tJT8MLJSQt8mtS1b6Kf3Lq+AYdn7uo4+/DINBPdb7pZFMNAnbfcAdVQJcpvIq3H74
ENEyZ4Owtiz/vtsF+y/gHtcZikIEUZWY2uChk9bxEjA50pOL4Qa5qbdPdGlh36dNDf3HU01DrsMG
qgMfa6x3+eJyIV/w9ypxersU6e+YRxcial/L+iBlla3BXY/TlULE5leAPt+ckVmBJ6HywPbAHYTl
y/64Iri5eFLuULnOPdk8QG9mfhJ81CFa8/XenyJI1AmgkzdVuQNXyYt7cg/YqLWCRxPT+8PxE7vh
qzW/YnzQqJpuzhUu+ZSsB5nS1eTP1iJ+zKG4UYuFcW+oIT3vC9ZCvF0g2aTMS61sckQYdYjyvYQn
e8i4WBFiWassyoMcHS+Ua57uce+tz1BSw2I+T7VhI7QZa9oPvXpx6HXK3LUFMyqUDO5/PsH7pzfq
PkJQvChJyAKCkATOWlTVvU4CB0kqvAkSGI9+wrU+/0AB4eTrj3kFx9P44l7IJj+EBlSfwZJ/yWmy
+JPPsrs/jcJ6ZDfibguKKH+0hLYySa6i7qGtUFjw9+V+i9k4SsZuQpylj0Enpu1g5PYAABJIeALk
WTk4yNTc3xiBbyrnF2PrTXRxrZeDXVWUz0Xpd8gZdIae6VMgdwrdfyQ7icvOjFqjwzMkHb/u/QZi
pL+MgzfZZ0H4UfqfL+v8chUEWjUmHQpE4Qf83dDPVGR7hO+q9QE1TWCKjO2cHs0GV2VNJrseWpMR
80hQkcYgAU3XZnQwtWsVUXZARjLLvBE2DxdHeuMfqzsiJdLl/46b+rnCuWHykuizQx8t0xWpsTsW
LntFiYNPwZHP/ul1llNYiFRe5ljpjTPN/Q70YaQyCaM2O4ev+go9I1qDAcX2kyBJdGtjbpqjVJO3
FEUk1BDH6/Z4WjvUQS2cTcZSdP1ly1DMduqC3lUeuiL0tqs0gdarRawJKHS57KCNSLclSVAGndpq
qv8xXnNEMXx5CpluNr/yKY+HfR4OnSecSw2FM+E18ZTbdM9kK3hSjiTQ9P7WPtHeqK+THSx3TcJm
C5qr4yj4l1R5XFaG5qxxHPM7qt74Op3O5/yt2reWYl/ujBDQ0brRODmg1NvQKLknX280EG99Liiy
20RAVLc7mlBFxMjxHFri0Zw6YpT9+IqktpxQNgEequJZh52E3ljhcBoeIfrekeEkbqRcqKnoqZfO
L446romcJY9DsSCaKWbBLHpP25naKlM4dx3RJWmrhtY+JBY9tAuTb6IhkzMucsbBWWO1zCleoTNa
iebhu7nRgHON4vOB+yWulO9+87SHK7SmPedy1dTbI3CQ3JYQTVAWFaq3XpUbZVEy64RP7ZOp9v0G
Fj19CWJyhkjkVxDzg527o0NMnbi0r0JOj6JNrn1bic9xC13La+oC/VRUvO5MhrTYDQaM2Nfv2s3b
JwCYnXCHf9ZVnNGphhR42HoE75qNzYiyaVh2QJNbAj4BEW0zvTlSTbusi3lzpF+mrG8Tli9oKgOz
AA1+Wa2zFNeskhgfrls+V6gcCwJs9yXl7I/uCevZsTSY/wSxHdtIMsoV/6W2t9JWahYFg8lAqJaM
uTASEX4Ia0kuY5cLudrqiHQ6bh7ipyySzWavZxcysJHu2MF6nGrBhMe/oDNQ5TKBemTDzAcjZ5HY
epZNJMYmeOWmLv40usgnCjv9iXtnmGnEoB6CbH5P4k+LaxwwVxcnutGp9kHAw3DC4r4rOLtjPoMV
jCBtjPve4jr9bGScJIgV0VnJx8B/fc8IQP/HXIigBh/aclmPWmLSggnX4R7orLlZEgMCMY2U/DuM
tOs46EFra+SShjcXqZSz4Sy5w1cexbl8gSRUx4X3Nwlo8hfXqnUhM74RPRIvZDqj6Iwaqw7S25/3
RpW8CEjZt/ae6225MAvUQ3NfcoYMihUlu/zker0+86tDDafQczNBK2PUz+SA1rSPoVvwrc8aptFm
OGKXqTPoA96KRplBonh4HDxWsDBoVi76BcvBy5JtT+DS8jLzQXi7c1+YR4xaufjLCg7NdcHKL33K
0hxMpCbBTFEj60FNpehfP/HOQdeqWanaHO9cqkAQ5ls7AW4QY0HOXDyAT56+fDOD+dLF5yKYn0l2
/ksNfP/cf8iOSsLYPu/HtO/c1uatBZe5V11asA1PCU7aHcodrzi8/DXQ5pXVXWY5g4vuUq9oEVXf
gA3xujYlN4QPm4TcqtUlFt2FB6NijrL7xnTZI4tL3H11lW0Ji5lbHkgCGvO+BbY582eAGrQEE3zh
EzdaTG60DXOdk/7Cq+GWMHMlb1po1QWKktCNPAfBMF0/uwUY57WtDfvCutLwzW2y6Rh/MWV4DrM6
MTH3hRZhOAy7AUR969EKJSTwMT8Dy97o/b7LVj4tlVnu3lCD+cZG5LVuWmChBPVqo7f5pemOh2fc
Nu29JYFZ9xa9P9gmvLoKwAs4WBPbGfHJ4XAqSNb+1gPzbvvvy9BfQVPqiY/jO/VcTdHzfrsapFpt
yeR3TZnfItFJmhKE9SHn8haS6hXXFHP5EL8Vrl+sy1gkG1qT4t3UnH16w5rsD8I+GSgzvq+degX8
5RUdxEx1sYYR+9sH2j7gf+llKlR8XnLZC/xinp0nULI4Q0fVksKQONvDGxg3mccZ5V5sJsOkXNUS
yhJIM+YsMlgh3F8AOTlUxRo/3/ZVM5NA97zUKUF2OW3FpvIgupc7fXE/2n8e/6cbzuLieZ8sJBX6
8cDmkFW0e9gVFVUejTd8XZdfRoL6u39awbrd7AteEcg+AxgCHV+jyd9bPlT2s/7e/bTh/v5mVeTf
mh5lpSuwWMU/K4h2SbinzY/SuBysmN5stnURuvY/nMbUx3f+4E5tLg3C4L0SzVGsJ38++rGGLc/c
fAdG2Iko2+WjoLIIc//V+Aw8cGQnY3cu8Me2wXW8f6EP5JEf7PVH/3u/1t3k3KakAHR9C+ESBiIZ
+LkqJwIJDRGkElGtnJFxa0xAR+daRrVqbxeHpVjoFvlu8SCzirYy7pd8NhqRuBAmE4Il7cEI4JEz
whWSb/xRhU3XAVfmSdVI/mi/WDSc7CldJ97v85a8HULOdGREBSH4/hXyr/veytBnu6j7D1ea3i29
08bgSVbIQbJQy2U/zIZMDP9VDcEfcgOiSOnQ1LIUEYEGSE2vC1EwmPaU2MzmmMjTBsTC2SpGPgA2
pgwa+3iX6LGutLFX40UzJBHreZkvLN1SztT2/RB++LlClMES7RY2wRA+Ypbmovc0gH2yCxrUIYmm
qopfPQJLrk8M3IU94ee6jXhdMj5DO0kn/mTgcI6Dy3gWD7IQTnYgU2S3P2yJ7AR8Uc3dg7GJkZX1
wXgOkjT9ZVUJiP/h5TgUHlZvUrKr2gnsO66/GIXIZvk7MU8PxNq7IN/unDBqHEwbJlF0ocMQb18b
rr+WMJ0L7dTWkjkqy5Z5spcJkUz/pC8K9Dhswcj+n83wYjVpPUQpz4K3uTLArqTQx8ZdQmp8dXr8
0q8O8XaSBegYP9H+giPZ+4IWa9iwtPO1/OhjrBCKognLeC7bHrZDCpcA1YGSnXWSrzhhvBitYLuC
aUPuwR7lcCsvH6zroMtLLjJcJb86vetAKO1O87EhAnqySq8FebZIVXvwSnbLXwTyWkP/v2KS89gu
sPLiPPeFfL9GIh4nvDQy8IDOr5P5GIRQhAA7gz0Oo2hKIWNpTNeXLq8Lwyxg34z+3WHLw7zP1+er
hoCJCupZG2LM02ugSteyZl4rk49laYX4LixDuJ5sVaoQXqvUGz36eBtUXeGYZ+EPfkMKEqh7KcB5
SRi8vjVPfuXj4Cv9x9cepubt2jg9szmbbywgk89tkT9XGs3paws4978Z256eXj+qGultCzzntVdm
dOFP8BAoTAm9LYGOMDKi1ovT7LKh78cHJbiLFosyzet7m/KGyrfvhxUbrxOoBGyXsDxEcUylfudC
oCH5xSa+eCfF1MZtnXHlZND+VYhdFf7bkPbEssAuXWIJHSgS+1YywyeQ/85KcmG2tVE2SXQHLhL4
0q8I41suIEzpZ7JSVdVLJPWdQ/3peXexuey5er4dbReR7KVnfhv7CTaYS540KkQDsN+bSeHkCIni
7fxjUrVpB/Y++pgcVsxu2trb8CsNKW/DqBIJ8VDl7TGkvkuQSREpaLU4nB6NZCLLXRd3ORz249u3
cfMWuh2OjAbOgy4TLO6T7eA6eBPW9CCTNzJsB0KmDerV9lsdbMKPczM/QogNy33WaLiljv9yte9b
Fo/tMjE56yNjOPirHO7nqh60I9AUlxUDPZhN4biLB7YeISZUTOPiAleUDf9Rv/3gDBvtihIWLX0e
KyrNYXfL8ADYLvYd8KVHvmdcqyjMSy2ZQkuhkoZNiIYzKzxMNP1pdnaND6hLAN1qWbVEBns2Fcvw
6/Vm39OM6wa6Ya+W0w+1WZqlZvAnQxWPjNCjqRpZJTbfeSns3jur/z3lX2UMu/jMVuORZuLZq+4k
TaH1Gx293qIO0Bw8U72Zqwq4VsLM3/vrJGoJOJJxXh8xHbzAztORgs9sszmzeaiNez+Y6b2igxnQ
y5aUAlWnxQNYWB4VEnrhUkx9bCEyTovGrX35AcdnP+7sLF5Hh7e/NYnWKecbiTD9/XA9Dxrs/CZ/
QbPhk9zkyXW9TPJm0hbdxJ7k/cH3D3mXJaa1fkdfqz8MkI1hHsEVqBbWntHULxSu7sfCjvBeyf8Y
25aOobr0TSYnndtNuUp/sbgj3BcbszKmbo0MRu/7xRaHZx9sTFt7VA8btN0hBVy5MJEmrQZeBmHH
tmle6SG1WQDRc+qv1vgTFev9W4GwnaWJe3N5IHLPq9Nt99WCycE1ZH5VKNFoxjjkr1B9d/Jnn+oC
31sl7A==
`protect end_protected
