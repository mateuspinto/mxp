XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ϓ��M�I� H5Z�j1-5�a��cꙈ�UI����)<gƲ��2�%S�(���mSi��^���d�v�c(�߮x�P7�_2�ಋ�Q��J�'�<QA���Ų*�� �]�U��Y���,VjF�Y\�~w3Z1SW"Փ�e�c!ͽڻ��P^v�2rnbxU���],�ή?E#��m}�C�bi7�^�5�(�7G�zRg�%ǭ<��k�' v�M��T�j�{LQܻ;A��<���l���n��V�������6g�=��s��I����6��g/�pf�r�,�Z�=N��{�FH��Bp`ߍ��6ҳ�z��`ݠ�_����h�>[�ֻa��������K����w�l�u�-pr?W:ĸ�Z�xZfQol�9�)�X�=�bS�\�������*�G�e�� ӽ?v5~�2\	�ISx=�Q	.Cu����ۤ�>*��i�\Կ�n�͐�!W�B9^T���R��O��� gF.�v�Kr�qHc�%$�:M���%��%���¨`���Q0$����������~uO^�aó�-�F�A�r�aI� p���b�N6�y��B�#%/����o{-���T��ͥ���O�?�S�0�-	�e���[������'�S��m-,��>�=�o!�ݣ��� ��zڪSɝtaO?����A�&"7>tJ.�K����i���Rw���b���_�@�|�>ڦJ|�|u�-�j���t�6��|X������t�y�匍0�;��aXlxVHYEB     400     1e0��<�j}��5c��٬��̀v� f��uu�Ql��]P8�0��>s���ׁ��B������N�'����f�_[���uO�ӭ SZ�^&���bڕ~�$��0�s�E}�4dJ)�����AN[�K��z�~�/�1��{��"cLx�L~U��uд)9�zx9���ei?�~f�=�R�����<$Ǘط{��x����p.w�2Ō7�����%��F�x���(ή�Ϣ'M�o��ޅ��6��&qC���D�� �T����R�Su�onBa�Nl.�`��/��ݱ�B�;��@I /��%����{���v`�k�� T
$D����QOF$7��ݯ��։�:ƫM�}.�H� U�d���yQ��F}�������dT�4��?�������9x��]�b_9���L�2ܿ���>�]��G���C�U�f^?�I7��_����"���b��Kb���"6Nkݳ�p۰�i[2XlxVHYEB     400     160��T:�Ή�F�,u12J���t'v�Ph����SHj���"���p�����rX	6���?R�й���)hq��_�M�o�������a�w�����)d�悟��7l <��Kk�uD�����P9,�����5�b������#���A��j�G��h�8�)���Q\�E'�J�z��_��_�$����dy�9�lX�bC3(��Q��y�|%�|��F41��n�,�e�� �y���j��uCկ�+|@6T�	1c��?�uj�3%z�(@���C'��Ԟ�|P���22ꦟ�z+n�]���c�bnU��>d�'_��%��6�b���{������:�����Qn�i���l,��XlxVHYEB      50      50�t�Ml�@'����j��~�HW���Aȿ.8n�k�"�]�W9���_�6A�U�?q�:�N��׀)�o�
1�z6���$�