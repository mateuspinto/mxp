XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3v!�{@~���6j}ի��-	с��i��1@YT���L�����/r�=�#5�h,���5������P�9p�W�n��Q+�Ƨ�o)uF�d�C����e^v���]��A��$��KBx2�I���NKi�����$<�����Kh@je�R�S�:�T�������8~g����'�}��d��t[0w��+/=�\�g|g[�*@��C�t"�����C�b�l����f,F�,B}t���"�K(�Q�r���q?���Ȼ�X~���3�?>�D���d��W���e5�W��\ܲ�����	�y��(V��S�/���o5�p��&'jd䵱&�5�����2x�}��W��`���5W��J`\7e`�-e��v���5"��8�ɀ��Bs�Bԃ����H�<Ce�%U"���DUc�4�ht��J� p��6� ��Ԫ��փ�ɇ�t��Z��vT4/+U��ܥ����a^�/>ٙ�t^n��1�Ls�^9��3<g};p�P�	Ad�~�m�ӌ0e�qEz�f������:;Q%���-�dr�1���@��4�vD�Wz��}���*��q�Eĕ�)�*�Oq��c��9�	k�n�d9�CU��d�%�Ze�P�4&���˛��	oNX���O�Qx,�5�J|���va&��B��,zD��a��
]���.�D&�r9�HԢ��;�&s�7�c��Q�R�O����
�|��2v7Ç�v��l��z6�� �T������vh��F�"	Ĩ�����ǽ��XlxVHYEB     400     1e0�7�?~����H|���$��*��г#�	�4y%�N����/���l�r :$��GN딽��3	�ʘ�%��@�T&z�Th�|1�ae%+�	M
><j�*p:&�[�+�͡���t��S�1NQĳa0��_��>��<�%F�P���J�II�H����hp��7�ɩ/�]�FYH�\U>R�#4?B$2����\��$Q$�~^ ��ܸ����bn�Oxʱ��)H��+|����[*,�1?<Ϗ��,<tP���]4m�@۷� ˆal������f��4�DL����l�i�ļLC6O���ef3�����o���^oC�#.�s�M���f2�}����3g)�+�t�Z�\��I��l��y��Wi��ꩆ�鰱�B�)M�F^����`��j��|H��AP�o�t�PWA}���c���H� �ˉ9�e��Ŋw �iN��X�w�i�d7���o�A#C�J'�j�B�XlxVHYEB     400     180[��Q��*�0˯��Մ��?:{��g	�t��5�6�����C7�ksc�T��BK/T���_{%�+��!}w7ӟ�i���;���\!���s��*c��rO�bf�U!ti\��Š<~��q��<7O*(H� o?�NqhJ�ii�n���2�W,��`9M_��-���>1I���n0���Ho����K��������8����K�����M�N�2�*�t���"Hc��/�}D߅������o|㤢_����<�р`V�i����I���9ֆ�3��F����2[z"���V�B�����`P�N��w�
�Spb&���3������~�Cݗڄ���J���v��P@�V���N�'�o4[���6�s�K
����T$XlxVHYEB     400     130ot�%��A����Ɗ$9���&���3�E;�����+������*d֠�s/��a�V$2�����!�D��ȃ��'��E��8��U|C�]������T\R\�QW�2�ڳ�=����,� ��[�q!u�~{?%_��=�5Jk^#8�u�O6��`�{���e�� �y�3�W��tvB�����q�g�E�M�>T
�F$gK��F�8�^2+2q�yDIMe�h�*��(�E|���6����h�i=�!;��v`N	C�ė�4��*ڗ�����S�!��D�%��H5_��#�X��E�XlxVHYEB     400     150Z�Lz�IF���Myn����k[Ֆ�	O�Y#�a�KH�\� ZI��ݤR4�r>0�J��5��}�=twRwg�5�i*�"��Hp���m@��%
�Kđ��Y�6�$.�hdL�=���`�j�N�ȢF�<���,	���������x��Ƶ�OB����V_߭��z0R�>9[jnڊ�uu�2�+_�MDض���R�p�I�����&]�Ǩ�i�䊿"��	Xc����6�Z4>�#1��h�غ��'����)��L��r�Z��nRk�ϧ���0. P���*���:_a�,j��mм)�|'�@�9M�v�'M^�������\Ďa�5�XlxVHYEB     400     1a0�?V'��������U)�ؼї��}��is���!��z���N��~M?�m��K��D�;�GH�j��:8a��sdϘ�#�7�� �0쩘)��B�������ʣ6��S>6w�j]��d(�F:��щ�zK3�'�S	��^U�H�%�܈-�!�J���muW�%C�dR�,�f�i��V^�
����;� ��p�����|L��g0t��-��Q��Z�`���k����v;58��˸9�r�s)?:��\��T<Z�5��e��W̢u1ൂ��h�wT���.ؿ���yA����C":&�|n�UȒ������#W��g�@��@�8���P7�ݕ���U��;o�Δ�#�B�")��𐪧�{����L������a��59�LL�A�����P�U����W�XlxVHYEB     400     160z��Ps)��M=����q̔�Zt�5��%V7+�g�.>ҟ���&�wK4���	}�|�B��,��2�H��製�F��+�ڳqZ+��5�A�њƉ�^�!t_.qC�m��1qX�s�X�n�K��2Ӌ"IK���p6��t�8i"�
g�T�1��|b��dk�=iVS�dt���a�A�9YK8/�`v��XtG�G�ϒL�e�k����D���tҼ� 0�T����c8��8u�5�w���4���w��qEپ���+y�0�x@���KX�C���^5楠���3^>z^,�7��Lm,���E����ݼ���� ԰��60��!�j��+��t���T�p�o[�&�e�DXlxVHYEB     400     180��	�K���a�<��GN��o��*|)#&�H��T�T�I��	f#Ī �3�1jP,G� gFB.'F�Ma�UL�����٬lњ�`������tO�JyX��ajJG�*W���D�<�_E1is�N��Hi|�S�j�Œ�!o.��f�2P�,΄��@��{��Hqj�	�d���`W�&��kt�h$��)�Zm�0W.<���u�'gh�4|\&P©1��*lx����L��\j��-�ஈ��o���j�j�!��^�:Oę؏s�:_ψ�oXh�<p9��m����<�P^3GJ/Me�9}��#*JF�_x.z6��&�����`8���]���b�<<�>hîI�j����l>�ĞÚ��O�XlxVHYEB      1b      30`��Ąź��T�����r��ZO	3�`��2P5ަ|�T3���_Q