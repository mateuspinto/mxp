XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���TP{�r���j�R^!D��Z�61��w�!�&{-�WUj	vQ��I�Ki�"��RO�#�|i���"ш��`�X#v��%��T������V�����}��&�gذ���b�HO���	{�@E���l�{y]|��~؀�v�Hb4��_��E�� ��7!=~+O�? �l~�_�]���G���8h�'��4f�n��N_S������i�Ə�cɾ�a@��ϳ�Y`U�v2w��s�)�w�7E@T������L�`��D� JBy���(��E���h�<sǲ(˸9�Vg6Y�<,}`Ք\��m~��3/Nrm/W��7�R���q<8�p�����ݕ:�i�����1��O�b�[�2��o�P�bEm��ad���I6r�:2
1Q=�4x�0Үʫ+�4ك�r�%��5��qW����MM;��/���{D�%�U,����'����Ͷ�h����p~���B��M+R���x~f�!��w����u��烢j��T��6�����)��gD;7��>6-����{
�#�vѱ��}L���C�,�:�UA����T�+�*)��GY�3��6�;��9����3w������O^���I�[�8	���A��l�,�'b�$i_�Q�����>mUx�z4ۨ*_����A�&�SZp��1�gDb��#:��N
�a�)��J 馁6|]�'�����ë���vl۟e��rG�r<`-f=��l���S|85�;�؟���[XlxVHYEB     400     1d0���c��z�ܣ�L�F߆�d�d�-��RaU�?��&l��|0
��&������[V������d��`e��ur�8�#ky���'M����y8�\ઌ�xt�E\�8����BM@]hk<.)�8慖�Qs��/�4ȶc�!���*jh��ټ�'��y�>^�z�a��խ�"�f�2�?�H{}��պ����~ �����Y`x,�q?
}Ȓ��Q~��\ѷ�Q���IݳsĞ!)*,�mPF��i�Z^P;��� �)F��}�t2�L���a�*-`�%k�w#�D��D��Ӆ!t[���������)��H� g�Sh�S�].��C���N@ݣ�8[6Q�KH��X��_��0xf���jI��M)��1��;�#����ۙ�o^�D �8w�5�%����d������v�*X��Ώ�xD��d�Itm��(�
!XlxVHYEB     400     140�+���)��wF��Ě��-��sτ��ˍI�l,���"�wK3� �Ps��q��N�1�r[0�X��6�?�Ҵ�@��.]�B�G��P!<��:&x��8�M���R�\3g7���~<o�d:��t�]��7�\R�!]WO=����3�H��W�_J��;fX�hG��e����g1�%Z�d��!��qsW1fi�����t�� k<�W�c�N޼����Fp_���.��էS@��j�ls���Q�A@)ʾ�J0�� ��//8f�<��u�E1�n��$&���ƃ�֙����Z���ܼa�MMXlxVHYEB     400     170d$�Z���2��׬XY%�P�m}c<Gk ܃�&����V�L�8����{��T&1��z��-4^��/6�o$�QM��ĭW1��⿂@�u?r`�4����saL��<:��u�^�=-$�])0��hr�[�0�O����uĄAL,a[_�.�w��L�$�����W�X�]`�b0@�,8U� �N��:曢�'2?k�X��V�AK�MM�[��[Ȅ:N1�����ҧ�}�@X��}
R��J�D�:�Y����������`�pk�!����0��>�H8���L��+�:�"W/�g�u�^�B��4M����ߵ x'��	��=�,��,��b�q�u����R�[x�L������r$��A��XlxVHYEB     400     140��Pyd������H���]���
��,��74�{�
8��:>]����c
t������~NUW���o�� �z��Ͷ���	.o����W��+`�.�q����e����Wo��y-S�0�T%CWJ,�c��C��WDYe��l�k�%���|h���7�bA9W��̩P�t[x�>zo�U!'FZ�7����8��D�*2+�JHй.����
]?J�OgCq	p�Ԅf�
|?7�7'3n��6�R|,i�蓐~�kzZ׼W!�=u��$�gkt����J�H�)>m2�n����T͌%�~XlxVHYEB     400     110��[jb����dW]�0��1g��8Ԏl��E��@Zr�)|'Z�5�L�О�L���q]�p���jbX�r�g�XBA�ހ�zj�,D�"r���&�����i���:޷A�Wf<�]� ��SN�O/&�$���)jy��)��s2�W�r���_bOM
i7xL��� ���M����g����.q�4V+	�d���U+0�g*_�Z�����l[Eq�fܾt(�x��2�4��2tg��J�8�r�ݛt��� ��q*M�r�]��aW{!8XlxVHYEB     400     120�Ђ1��P	�P$�4�K���ۥ#@�������OD���A��ܥ�n�JҧG[q1��*y��P`�k�T��
5c���3�ikv����ޓX@zk 4�*'��ѕYY�\�� �Lpr��eT���~V2:,���&T+ ��%��{�P�!�}_W���u����}���r����n���t���mʧbdbt@���#H4�V�e�8}?1��=��[��9e�{*Hv��pQ�>�&��n��NA5��yU��UR�I�c&/�;w��ߞv�',1�~:� 3TXlxVHYEB     400     140��HXk���wr�b����k��%�,��X/�0�M������fɟL<�gwFU^�B�^�3{Tz&2�w�+B��q��0)0Mԙu�����%U{L�)g����\����d���az�m�r�M�F���w�2�M@�kx+����zR4�|=x�قnѤɩ��v�&�Z��-��w
&u�G��H*��O�4�a�W��Ew�]�A�AU���G�3
w�r�����hl��I<���'��Pa�1Sp�0
���_e�8��G8��ur���wBĴRi������$<�f�|$��)�eH�</��Jo'm�XlxVHYEB     400     150�?���+�*1��fm6��3���[�*~ �m-�Ў���u��Y$�X�!Bk��%I��Ǚ�$=̃���*��};�4~W�	t<�!�͗��x����9�F�5}f*�3B-#N�T
f�[&6�g�Q�C�SYj\'�<������)����ͱ|�c��:n��#:"vrh�l�����a�_�i{�L3�x-'��u��?�G?o�	*W��@Oo�ʭ�lS��g�� 2be+ɇ��/�Q'�І�(!�)	��E7
�i�o^b�h�����vVV��$���	%��
���I~T��B�'8�u��^�����l�}���AAL���t@�}���nzDIJI�XlxVHYEB     400     140����<��R�Z�	�i =`%�0�����Z�bMV\�@�FM�@ls�Y�M��:�"xT+�J�N�y�UJ�`|T�I����0H�ә��6x?��m�W5�(zV��K$FM�:���>�n�9#z1�v�K����+t�����xpz"���dV
q�_yo��ˮ�\W�+��a���aȀV �~̏O�p������@�
~�|���D[+�'���eZ����K		]@*����{A��n�B���c����C�$nKJO_��Nc���a�b��!(h�rx+ 5��hHu�E�Ry�%!ūhXlxVHYEB     400     100`O�J���0�?@�v�5��3F���O3�^�SX�!��E�f��Y7�Iq�S���w쳾�w�*���2L�9�"��g�����Xr�S��	(s�:��}Q8�8�@ -~}����D�0�-�."����Om��X����6�����R�Ӊ����l��笑��+���c�������fે3�w�%��w���o�g�y����L (a��	�����_��H��!�6Ɖ�����Nf�YL��	$<�F^6���~q��XlxVHYEB     400      e0�b4C���Y�t����'�,G�[��:[< ���G��ц�����?��|j���)$i�Hq~J��	j��dX!�{回���޵T"䙦-��)�!Z�'���|����L�NI��tͩ+�#+F`����uc�j#7���j5h�V�����{�ro߹h�hv(��Y!�y���o�g�K�ÝBI��J��f�'�+b;\�N�a����s��VXlxVHYEB     400      e0-�����9�:�j�f/K���I��p�׸ ���C$�5�˲�A��cq9�<Zi(W��&2���#���۳�V�%j����hj�ͷ��K� ����^39'������*��]��v�m*�RY�|�*���]&_+�*RĒ�ܼ�RC <�
�N��#(���Y����bŜ&,%0և�e��W=�{��#���*��9����y�f4;%t����XlxVHYEB     400      e0l�+�.FmT�H��앣��;v�����'0�?��+�������1��w2���Մ.o��,���6(`����ΖӅ$���U�7m�ؔ���2��$�"��~t�{*�'��Vt'&�`"�;#��I!�Z�qݧ���n��ӯ��^ �e��Ș�0�Y\�7�H!5���A������CD��r%2|������<y2���x����a�L��H7�
��XlxVHYEB     400      e0�FRԞ8�Ź =��������������
��ɒY�<E��T0��ӥ�=�,��/!;v��-����� ��E5w=�5�ux��&� ҆�/�c,�
�M��2��L�������S$K0�F74Vp?s�J޹:F���Q#��s�hQ��X	?��K5$	��?FZ��8��iK4 �o�ķ��+Oa飪[��N�]VϨ%���~��Q��XlxVHYEB     400      e0�PqU��ݥִ�A����!j�r�_@����|�2-�1�|j�zw���I�M��VY�÷�%���{�^�OB�K������]ĨZ��x⛋��L\5���!Oҽ"f�U�� ��f1���p�~���#u�U��A�����K3?ysBd9:�0�Ӗ��K*N(�k��'�B�\+t��[y��ÚB�n�3V :�ji��C���05�N��QA�-�YA�|k���,#XlxVHYEB     400      e0�rYm<C}eh���lo{���~V �<��zE�s$��{yuv���XMa�&�g ��K`y0v�'�ɭ�sk����5�+0��!_
�!�2�����%��Y2.�Mu�QhC�f�\ɕ��w&�n�HZ6c�n3��Ҩ�0?Yb:�s���&2�D�k��X�^�� ���F��Z:"��i�&rk'u���)42v��l{;�)sy����.k�]ܟBۯ�_�hXlxVHYEB     400     1c0��Z)Հ�d$-�h�K�VA��\$���|�c��B��M�ڨ�Q�#���]]vaޡE�Z���P��w5�ގ�|3?Љ�ү�-/i�*���4���Ul��q΃�w�>�(+�����`������. J�:짪�̱e���nY�_bfpq�PY4���O.>P�@$��v���}��`�}ȹmv��p��+��x�����~� ��_!+��-vÈ����W	�O��^���b��bgS���Z����W�����������Y���a�%�~�L�{~р���{�e�l� m��SV1�`�r;���a˗T-�����`�?��4K����ĵ��h���F�^��w�w�܃a�9���8�M�ݎWm�\ټ��TY��a�b��RS�;|�Z
l��<����(�n^��E��F1uÉ�X70"�#w��fN����.{2cHXlxVHYEB     400     130���,zZ��i�H��#��S}z��QZ���X��BD�AjyB���K��X"vh�{��1�ѭ����#��ޚ9���d�F�/xk�S�HC�����_&�M�����YYJ�Ma�B��Z�3���52�����=\��B9���k�?Z�?u}[�F9�1�]4R�W��k�QRz�nUX�q`�	�Ih ��k ə�Mso�nB;S@4ah)}�>ύ���Yn�PW}�G;�
�jj�eժ��F�qWz��J�5��0Wٳ��J�%W�
��$�f_s�hϮP�r�58�h.Jp�~DXlxVHYEB     400     100�Y/�����}o-�r�H#�9B�atw��a.�F�����^/xs��bL�ZV@%�t���IVc���>��V�_��Rw���@����y�r�/!��ô�k�,���
 �;� � bl�M����������& �.B�H.� ��_+�x�x7��k�Iͩm�]+�5����NY����)sd�>kp��9�T<�t/3^��N�Y6X�bt�\���"�z�;_ڿT�TfPf�Bs�&��]̲���h�~h��d�XlxVHYEB     400      f0��Ϣ@6�ִ�b�W���Z~�:};����x���M���H%��&�/��@gf6pT#P]�a�x@V�b����´?G��t��i�>�-�#o,t�����{��B$=l(O�����/d�O#|��f_2�dB������:��|�&�xYl��7��S4�I�d%� �N�^A��a��].f��4g.�/�р���ĩ1['�Cq���|k,��1ܶn�XlxVHYEB     400     150�"h|LFu�\́+��:E`8��u��' 2(��aa��Լ+�7���s�W�,������63�EP�����a���ڌ\m(ĝf7h=���Ӛ�
GF]4�R����c,
�1E��9�w���cg��(�h��LR&��^�ԅG���S�IM��|7n�&4[�y-V���4���u�7�jU�Nd �*�}&|}���HU�ң3'��h��W"R�t�\3��j���T'Z�[�遧�����f���_�9��}���|Y$g�}�H+�u�蝬�9�:��ON
I"g�n��p���fD��-�/�@r���.���;��XlxVHYEB     400     160�㲈�Ǩ��0Q�o�ӑ�����,e,�H���񝵷lz�4�(�����?y/.x�$lF�O<�x��o�s��O�?�d�W��g��W��>8Sn$T�5S�C�x$
O�bA�P�(t0��|��CH��4aI2��*f^;�jz��Ӟ^�N*�T%o��T�S�rH,O��ϘK4��Z_=r���AߥX�4@h^:�2�@�K��noPl�,�n]��-���k�a��y
�Ԑ݋��]�`�Rm���{b=�Zl�䤣�ˑ{ڇb�'�Ɂ$��NHogsNS�
W�����W�O�,��,��r��Z3S�l�xm��d~��Ղ�!�æ�G������ee�}�D͢[GЩXlxVHYEB     400     140��)�R��eE���<��H�$h+�|Lw$�x�H�
I� .�*�_�� &�GlH�`z�tU'*^-�0S.���)tt���2pi���6�͞�MT8�D���A�h2$��DD1V�Z)���y�� )tߚ>�=��_f�@NБ�Z��үs���z��\�R�L�����E�T����ܨ�e`�It�oͽ!���N>�4��
��	�F�A7#�ـ&��,x�6V���$�ů��{>�:e,RVx�OB珜#c@[�j��t��ǐ�_�����p	��G��I	?�H�e!�i�鰛UR������^�XlxVHYEB     400     150[���bxuzM��7�����CLصt�<O�h��ݿB
�RgH@�W�����8�:̮���Й�Gm�� M'28x�9K5̪�<��e��x'
���cC��e��a�z��[�M�r��6v�4d��Ĥ+t�V�ϵ�KOmI��k�H_�fo�.�|�G~����!�t��_��*���&l#��7(.c�a��3�x��G�I@�_�ib~L�$#9��A*vn��̃;��凷�4;��7�=����9Ё�hGo�V�u�Rr�|����8�R���42u3K�@�hz�ݾg?�{,].ae��|�; �R���P�� �h XlxVHYEB     400     190dj���¥�(���Q��C�$M����ؑ��|�%��x����g�7`�1�}ab��4�=�ep[3P�;� �5�UYZ���^%��.� t���������v�OO���n��{E
d��U�u��i�W���/m������G���+�ڟ�t��ۓn�Lr$��.�& � ��6iy�|���&��I���9�PVn��]�C�N	jV8v�Z��
��F�nVYah;shlal��E�3��O�y�����Rd�U������>!�3��Ѵ��M��ޥ�ĺ�$xR.�)��H;�_�%v �߃Y8;�V۸B-K$M�B*4�����S;�y�5�O�����X��b^×��-R�M�tA��B'ue3���K*~��XlxVHYEB     400     120%\z��\�B��<A��?o�
��4���/o���$}*�ߌ��W5���C�-A$���m��i��3�-�u��܌w��;�a1�=������:��b������ �C�R5�q��}�J��9^��Ǵȴ2���:�N�,�y�Kp���
��1B#�A��C��E�f���x	}m1�dvJ0��q�������9;I~���ڸ�A7�B�Ċ	�9c�\���K�ޑ����S�;�����Eۮ+�&o�e%Xi� ���,�3+�Gk�XlxVHYEB     400     150Ǭx%��ͥ�@@�߲T�����Ǝs��p��>GW�E�A~q<�9�(t�����[?�"�?��2�έ;�H�ˋ;t�rV��A��:��C#��p-M���NY�C �7Ԡ�;{ Z�h�n_42�zC�y�C���=!�S�d9̈���_2���o?��`aEZ�[ٯϣU.0�R������t��焆��\W� (���dX��%�r���1{+�I�x��t�V�C
5`�����e@���(	�EwϏO���o�-`g�*&r�Mp��g,�����ck��#�J������z�+���d�9H�Cڋ4g��>�S
����Ѫ��1붷�,�9$��$	XlxVHYEB     400     160���`���U>s��n+9�Y>Y-<Ԣb�{�c���=���X��擢Av�bi�ÄK�!'N���FO>~)a�kW�*љt,��v�hq(��h�F\�E�4bp$���~����}躱�3�9�׹Z�&��l7:�J�6J4~������cm{ŝ����������q9�vp�6�jX۵;5��:���!���
PVeV�ʦa�r���~c't�
���Q$�$�,�-���| ������E��ͧ�T��y��f>��XZT]����I�Ô,����o��w>���n����
i�{pc�$�t)ȫ��0k5�7�M�e3�P��%�\��X�Xۙ�MXlxVHYEB     400     140�O�v��2�� �V�'i8�Q��6+�d�����e�5U��)��C���i���l� ��Yo,ڄ�&:��P���aqn�`1o�G��s��&�������3Hеl�*^�Zgh�xG�jo6��|'y ��-�ce3MJȥ��f(���ҵ�K�
������b>����l��h8q� BmE�z+�`��ٸ��\)����E�Y>�s�I�=8O�EW�r)c�!,ǵ1d���B?@��]�4D$
���㕶�p��� K����._LBEuol�����h`�B �+��T�6yc�@<T�[��G��I�����|U�!XlxVHYEB     400     180���'��` R��"���u��F��C�Q����+�(�~#�ڼV�6�)�����P0�hTHʩCu�B,֓�'-J�B/SQ�e*�� ��M�����u7�^����aN�3���� �ϡ�C�u��O�z�	)&�n�r�����<��O�D+.O���0.���bR��Cٽ�?��hb����)."�%p�:摨��1�;��O��N�~+)��[C�|�]�+��b�nQ4U2�a��i�>�uGh���U�`��6�=[l��<�w!LhSu�k�Vlշ��,W��g����ʅ�/:�-����욟K0i���`�z��9�?�H�X�b�����������մ����݃��<�	w:�o����XlxVHYEB     400     130m$���#�t�$RA
o@������&E�'�B��J��I��-K�5�\F��M2�F��u+a�Lj� %3%6� ]�x�̱�9�ݞ�n�jM���N���%IwV�
uW'�oba��hTl�#�G���:PiKv@��w��� 6�A?�?�f� �J���2����o����X\e�%5�Hڊ��3u�˩���$��Sン��*�%�9����ޤ�ג�����o*a�Q��&6u�ᨽ��N�6j����,��$���7o���bm_���WsO	}G}��FJ=����Z��p/���T��XlxVHYEB     400     100�K-�C�v�w^_@z�0�7�w /}l��~��
�o�3��z���>x|�VO��67{op�1��@tN\��*��F��G��ޒ��y�ۢ1�!�8\�t��.�	���+���pl'���XCp�a���F4�t�ǫ��^�N٫���v���[������W%�����$�XU#4<��0ܟ���j���g�`���N"p×;��Ҳ�~���ӵOVOs�qMp�`]m�_�/ 9j���ƍ���vM�䖏�XlxVHYEB     400     120V{�q�$�_�`���]�c�M�� 
\ϙ���Y
�.;���"�pj�Ё�����I��%�Ԇ��a�A]�H�hL�#�>!�Rh��|���6#FD!�5APZ/�֯�����~�d?��=c ���s���a}��l|�&<�������k#����X� ݵY��7�n�>��<�.����T�yab��fβ����{�`,�&�32ո�����a�ٝ-�`�hR\-��/�T��x,���y�C��%���������EBU: ��J�#��.���KRLXlxVHYEB     400     170��𮿋�oH,LJ3�`N9 7�ܗ��u�����d�����~K����8e�@�b(w$y�*} ,��+�����)%	+O��cLJG��ow�tP5�c7R7B�ф�<�;���@ʲ�]K�O��;�����(�9��㌣׮�W4�K����H4��M�U�y����rK�Z1Ly�Xؾ�����=�$�>u��^�%�asŴC_�L��c�	�Lsw@�  y54�~���񮰩wv�e�.b8���:l1{I\��,ܳ��#��\\Af��(�4	�#9�� I1	��Aoi�lZ�`�Ї[��pA��V�2(���S.�n
���(;��o:��E���xTFF���h�xM����^߂XlxVHYEB     400     170�wV�M���ɗ碎ѡ ��G�Bt�>�5�VKD-���t��=�h���i�͆��뜭'��Ri�<�P����x�V~�P-}%���#%ǃ������kX�D�
k�M.�o�jq��P���F(\�5(����8���k�4�ۧ>,�#�'6蒙�ߕ���Ěz�'�5�f@T�OY1�:�K{�D�����+7�J���&#����Z�xm�	��6�P2�c��E�}�����N�<�򖷜e��6�*�G�˴$�S�Jʊ�۝]�O4�S��w#�r�l�X�mdQӆ�\��nk����,�
������J'-�7"���ver{,o%}��B�	JS�l_��XlxVHYEB     400     190���n��B�4��9��nz&Վ	���D�C��/;��3��~�^Q��^o+_0�aY��E٣�L�m�zŉ�@�����$�X����F�+1|��,fg�����9A���FzkX�3d_\�=��rsL�����F���*f>K�8�ۚ�2��F↸M�]88Q{�a֗jˣ��H-����1dϋ�16�}�V�n
��������nXC�xE�⁄_c�����/؀c�gnD�Z����w����/\��j_��Ê���<_��ƭ�dy��Vו�v�F�7��H���}�Lhc}8ÿ{M3q���:E���#y��HvՎ�wd�o��!��>?O�t��`���L�߮���|-���/�٦\�����S�6=�4�5���g#�g[XlxVHYEB     400     170�K�g��c��Ѷ$YĎ�p�9� �������T�::Ta!͹��Gw��_��*ѻ�^�;_ؒ�g�N��!k]�t��H�(��Xy<�j���~����ݙ b��m-�1�fg
� a�RbaH}51*t�h��9�������5����C�����&�S7�Rf��v�+��h&5�8UVi�����J�G�d���_�jn����5s&k�����s�qT��E~߼�A��BB�9܀Z�1@ �szw��Y?Bvs5e�[���g����t�#�h��<?�/���(0����R����y�{�����f�	�d��l�f�\T�4sC��M�E�U¦����Ɖ{��'��Fs�Y���XlxVHYEB     400     150�<.u��		�C����}�q8�?�z������`	;� .�#�.e.PZimƞK�3��
�4Ժ�ҁ"��n_��;��RL�|ڷ��FƯ����������$ϭ���S��&��gD6�	�g[�_R��+ ��}�6�¯5*�[��?@Ȍ�	���?�,ӯ���aW����-ܓ�2qg��d�#_����#��0I��Z�J��o��x����v��ED��v�a8���B<_��<6�94VW~9W\��&bV}(�X�.b������Yfw-T��f�iR	�`t�'�kR+�5@Stm�w�%�h�\��,ڶ�@�?��L�XlxVHYEB     400     170�����!����H���	�P{��4g����OoXT;è�OV|�QeN��s���F�l\{z�('�-)'��x_��a'�~��$�X_�@�}A������_.��\�YC��ar}���zb%�%��-1R�QTN�Ư�k=�/���R���5��1F��5y%=BV�WK`pE��Iw��t	�O�*��p�0�Y�xt����O�����-����2f��h�ԅ\h�'c5�d�|�����l7����\�t
D��WWMg�6!�w�?�1�0���f�jZ�@�g��ˎJ�0�x�G�f$i՗�F�Cm�rv�ơ$l^�x���2sZ2�i.���W�ǜ��s�h���PEnXXlxVHYEB     400     130����Ǹ��
(�G��OǺ���戕�9��O�q�X���w�w��.E`߱�:���IrF����,�͟���~[+-̾�|Ve2���@rz`��Z�;��-pA���!������o���P��U���!'	Ԣ�cD��E��u�7�e]jq�:���ж��1<�����>�,<�Q@�AP� Z��g��G �{����0��0�j�|H9_]��2����K Ł�e�RIb*l�ϥDHYM���ԟ�=� ����"8��%����#�|l�l7n��*�=B�Lt���Hh�tP=���9> �����XlxVHYEB     400     180������LY�bvTx"����*�\����%c�+wh(�5o�8v?4��Wt�]�z4n:�W��Jd&�hu�{�L���^x�WxDE�{Y=�(O���0��'F����9~��a� ��J�k�I���_��naR@�w�F�d,Rp���ъ�%ؚlȖ�j���}��-�*N�F\�<I!�C�%L[o_�@?8&�dŀ{1p�k#<;�o�l�W�x��DJ��ޔ��u��_ЁO�(!���¢S~H�d���Ay;;�k�D1�e��@gZm���b�eg��~i�pu�jfv�A��r��ռ�P7jS�rz���H/� CP�t��G����$t��(׭吔�Et|�O�[P+hW���~��"��XlxVHYEB     400     120�5@�ϑbM�Ϲ$�VM����?�g����/~L5��gy�)�	 ����I��4b�� �>��B�3�j�JƮ��L�4h~�_�?L�z[��&Y���Z���������;�p[f.]�`u��%��ф�c�<�����Ru`5i����+Kx�$") �N��7l�@C�,lnY.�/`���|�(����4�%L�n��+��%�o���@��Xg��/��v.���e�%fC-�CgV2%�?��xT���m�6 ��'��/�z�G��i\�>�,r7H�Z�fXlxVHYEB     400     140`��+��v�e_00a����?oO>�勾l�i�?W���R
�S�\Yl�*���G-oV ��ı>���_S��V�\E/G�*�!A~�����V.�1W!�fz@>O���^��|�;/���Lj��S{Z級�5N�����=n��H¹�o�_�9�#�z��`,V��o��&b�-bj�u�\��{��X!��]�G�6�if���ÀIX���LX�z����=E���v=Ë���%8��ͧ5@5�G���Z��)�N&	�Ú=V�b�F�-7�>��u��b��]_m��1@9'v�v�zQ��Q�Hd����XlxVHYEB     400     140ʂ�³j��z�ǂ����B%A���yHo��'�$NQ�rY��^#�[�n��P��z��Ea��yL*��V�s���	6.Q�_p���Pur��0�/&}�wؠo��[4=k���W���xl n�f^�O��\�ŬG�<�--3���;��b7�G|a�S�k���wG��\	n*�������r+��[�����x��]��r5|�+��4���0m�����8�5�vjS��,qԈ}�r��ٺ�o���6^���`�#lpP.�`3�v�ӗ��']˨�5�Xt"3&$ �G{��?�L%�+�'� �<XlxVHYEB     400     1800r���L�{g��g��kK)���ߨ���aϲ��g��	�
7,å���A�C�B�y(��ˡ�y ��UW�6�W��cؗ����8,��϶���;BV7��xe��:q�{��x�Y��9;�7�ʥ�܆�~�7��3�Lޚe�fjߡ
��s��3/�iǣj
X��N�ަ�}�]ތ_�YrVg���:�$_�]p�Y�y����^#X�ݥq�����M������#!} ؎��P?�cO���=1叓���G�cGz[b{VV<��8���4Q�������q+�<�w��\�D�D@���.�����F��4}��|���L؂v��QD'@��-&�NK/���A=�k�v`J+,�׳��֜�-���� �XlxVHYEB     400     150�	��x�:��3�D# �~\==��q>&J��!��=F��^�!y��1�$yLV��q�
D<T���3��Zm�ntOU����d����V�!T8��	~xa��ؼ
�9��?�emZ �=p��n�/A��s�������5��8�7V��!��u�!�LY�&�w�������A�a7pŤ�����.�X��7S\Sn��}y��Yk�� ��yX�t���)�1X
�8Pvy\Es9��ܪ��Lr2����2τ����uin�=*~'��)�O��&��#���?v�1��*��Y�J�I��8'k<�}Դ-�O*hC��� -l�XlxVHYEB     400     120R��F��'��ޭPq�w���y����r��v��?"��
>*��~uQ�(U�3^`�b�A&�m�;�O�~3�V�s��i.��Xq�4?�3����=@�Ml �|�.�lcxqT�;["�ײ	><��
\>��Rr�R�e�d}iJ
:z�
��A�9��i������.�Pߡ\w�b���}�ٌ��p�Q�4�Q$L'zЬv���kM���2#��I��,+d
����RF��	 _�ՕdAK4?-��X���%dp��9�}P�Q�µ3굺�R�t�D��J�z���XlxVHYEB     400     180C??nj������a���H�E�:�Dd����um	�cCS6���{~�q9���}<=}`��\׺�'����q?{�+�:�^i��q�c2��B��4M��#��F��؛��ʗ�����ea.S�@���v(�����.���Uk��O����D�e @|��#qV?���4��n��!���� �8�*4��R���W��Tm/RO��ݚ���h��t�T���vI��]�:G�n�LS���[g\eow�i�P3��DeާƼoV����|~���މ���A)�}ZH�Vuv��8*Щ����e�`藫�ZZmqƣ�QY�ӀH3-d�Y�Q�R�a¨_O�y��{�^�����$��jfM0k%B��XlxVHYEB     400     150�����ś����jbE���G�x^vj��
Y�bH1q6�>�xGX�-�k7�U�8qp�G�e�a���&cX)k�>�zb��V��s�:C �zw>���K�p�eŪ�=�� �|��`�;Z�( ���S�R�]TL�k.�1>�_�y���<w4�{�+���~���r����u���d���n��.�D�Y/$�	3��5h�cD�Uô�˶�l!��-�T*a���h���O�>+륭))P���m-G�	�0mk�-H���q^����*��T� .Uk�]��@,%C&����M�-��5A�̾�F+���1��XlxVHYEB     2c3     120��s�7�dsyF�/Q��O�w��s;l��85�"�� �öL�wS>�%yY9.z���7�U{�o6� J�`u��nk�OF������QP��p�qU�=wã#"�s'n��6tg4���C㬝�܀��� ���fm����^���Y��(������H�\w�j�����F6�t掄�o�sm
�c9$5�A���E�������!��`�{w���T��|��b����(���[����s�{��~t�F#��\�\�-���K�px��CS��qk��<��$׊�_q���