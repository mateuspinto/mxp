��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{C�%�P�*�S��_7@8�Jٵ+��Y\������Ƭ7�)�Kfi���ރ��}��K�}��7ibb��.2��
�lR��G�}RӀ��5��.9@�$ަ.�?�T�� z�h�c�qy8�I$8ҍbH?a�9=ڻʰ`�A�-���:bi��-��3D�Iڔ9� ����3aL��[$��W䘗��Z�)(n��ڡ,,�Y�]t꧰߹����)]�h
Vo��5�<���H-�K�$v/F�0����]�B;cs�k���3�}S	�}���ꂺ��e+���m�����e�����|�`�W(�?T�L��k�O�;j�R�Ԃ��!�4�N(���
NYac��X|2
\����Tz�j�ԻZ]7�@�@l𣓜ǳ�+y�W4 ����:�rq#� :�ĳ&�{��Dp���܁`kq��둩�=��u-i�0[�4�N�o�
{��������ɀ����2{�����K�ƌb2?c��2��'Fj7<$0 J��1��n�5�8AD�L�m��0S-!f��q<*k�� k��j9UB�U��2�Q�r$@DJ]YG.s(=��Dy[�pü$��ڕ��s�S�>2n������K š��"���I��"�ק��bFJ�{OϬ8���7���7��!��BG3g���.��5�@�_Y��#�_�~�΋�Fݷ��0�;�j�K�jN�M`vmYEդ�A��W�s�|��u���^v�JI&�*w���/����7���ip{���X�#e��2)Q=%Kl��M�=�dM���i|}��ipٕ�h3��F���)���8G�|#��_&�.�s N+���ն��?<y)�ٯ� ��ߏzإdZ�Of7r��р�����ՠTv�&�k���X��R ����;2D.�N�Io����C�~�����7�䦸L��^�b�{H/�(��Ǝ:W8Ġ.��܁+�{6~��k��O�	�{E.�#2�S��Z�!�w���1<!�G�l��&>��W7����f���hP]�ei�d����p�yx^*K��4`��7B�G����K��;����[�%�rĂ�R���Ū"� �sҾQ!���㴍;�y ���۰\f!����½���W���8~����dh�K?�O��uS<C?v��SҦ�4 �u>�Q�0��g����X��S~V,�:�Y�ڡd���n܎�!.rsd��B���Kl�Q^��K�8��<Pz��OJ���0�� W*��������[FY�-��Gp}�vsc�|D��zӶ^��j�0Q��Z6�8�܆xPJ���� 0�����Z�@���Q�l��{�C���l�����? �o���)��m��P�b��l�?
c@Y���E�B�+���V]���t>=��1��q}��*�cQ�;gcͩΑ
5�W3n��eU�����q����	yva�+J;*����'�W74�UEv�4�igm�P�z�I�AӚ�,�����#��_p�$���}���W��/�>�.�}���E� s�1|0Xa�D�����-�y����ۀ(J��E���@o�,�ҾP���4)���lX�N����erK��j��e�E
�=~P��ֲ��G��V&��Entrs�!1��m���MCn�3n������
vӖ�yu=\0�(�ol}�!�����M�_�Xy���<%���i��F����Y����Uh�;&B�;�ZO[�D�� 5���������Tf·'O3�D���*��U���h��%�M�Y�Y�����@��w�縉T;;Y;���h��87n3�S~Ͽ������T�"�d:�
��\��33�h;�x���a��3-/b_�Fb}$�*��`F���7~�ze;�
[�u�0cZ0N2����0"�.7���d� ��x����4���B�诸�{d�>��O0G֯����S
D]7Br������c�o��-J�N@d ���Y0�M�Ў��i������X���sS�(�=GMA����s1UZ/!K�hG����k	�(��4NǍ�U�c�G���a�r�2�X�(�F�d��a���Ht��F�[�����<6�E�M)kc=�<�؆��9{�Hv��&Y|
�̐���F��2o]�OX�ÁO�Aj����'���@�ő}�ty����&&\S�*G#�*:y��e���9Í=p(���DX`Kb]���U��	ӻh�1��Q_ĥ�_~`L3:̶�!@�%�Awg��b��H�-�\?4�e3?~g�&:��z��K��3�����b�����.L��|��	"k���ũJ���������[ɸ��^[�j�n�Ei�3g dd����.Dd�kAÆ�SG����G�MTŽ�`F#%����,��z>�K�s�aY۪�k�u���m~�=s
�_�Xa0�aLasBgK�C�S���%�'�#!�m������r$(%C�s�,Hxyyg�a}}�
=l����9[�(�O�z�T���V���7�OF����(bbG�!��u��c�����h����1L�L��`쑪A�
�t���;=�/��P�\�2T��x��]S���n���F����5�c�)�H�����DR!W5�#7{Q{R]�K����טּ���l��$.�W�ŗ��,���A�$��C�硾zp���/�m"36t!�1�3�"��/���|�u�AGk~�S��u�4����N�Dh����t&m|��5���q?Ț@c�wjQj ��F���K�䔃.�x��.�(��S�\�W���;�`=�~~J�!�<�t�-������L�����_���a8r���N�q�bۥ�og�7
٩�x��9�p`��p�IoH�������b�	��v�#�����=������L��|�8�#|�Us���,�yo�����,Q��h~w C&&���p؏��T��r)�����9��Z�+�F?/�9�)��|΋����M���ry�e���M�`n>$���W~
Oxr�-���A�|���<h�h�y� e-+�էVǋf�� UE�D�wV2�3��g��i������G�}��Ė9���@0�$��FcM��.}��k���r�H�9��lO��s�"<�Pq *�{Q����5��G�������F|���7Еd�1����^�W	��/_B[�#`:[&�C��JϨ�&�-/%R_���d"�C���l�q�B��&�{3��t����P/�(�kRțna.���?˫~��"P�b�+����p��'~�(���Ϙb��P���h��IzEoR>�t���&��|P��ï���)�-�L`�zImi@���;�?�4ޭ��Tww���E�&&g}-���2[ݕ�M��47�1N�$��0�-�Pގ���Xhs�G�J�aHl�����R�1��p���1�c�u]�Hg�?��KfeJ��4��b{G�J5���͑;��)�"Ѝ��ީ�w�����2�Ԩ8�i	`�c�@�f�<l/L��.!ݩ:d[���W�o$y���c}���U��jӸM�	偁�0�wD �y-oDܟ5��5V
:e�|�x|ɷq�q���z1Oo�-��j!|T��վ!؉��2@�\�7����ZA����db+]�	�Y���F@��R��+*�\�����y���=�)�^�9���)�14%�B-r�!����_�T�E>Q/�Z%Y��h������K��>.��P�)�~���Q���YBp�����g����1�W��,�PPP<;t]opƉ�}�#��j{6�?X�
LC��N=���ϩ'�/����O��3���cXΫ�5�B{B,du��e=�*���1�dn[�R*n�)���i]�L��M�7���*2F���U�
���o+3�K/�ȵ���P��'XY���기����l�^��)F���ec߭R��[-�+p*�p~nc
�KE�Q&*���'��j}���{��$�.�:(�1zN�tJ'07KS�:r�L�YR�
ux+~�2���"nxO�T���N�����Z7mp��D$��7�����c����ѻ�##�e���G���p!� )ﴟ*�V�=��[�Q�P|CzN�o5~�L)�:�O��?��u�af�߸�B�k�����p�^n+B�!�S��
Zs����dO��S���j�hZ���QO� ��7_n$���WR�.J�k,aA��S��XwZ���ے^
ipf����������rua�c��N�G�3q'PwY�Gm�s!��-l��d�[���(j)��
���:��YPl�!Y��ْE������厥t��q"	��tj�&��%x��|�R�lLM�.Q
�Uz$0���>R�9�ܭ޼�9�� ��_�K��|o�yʸ1���%��,�k�B��P#n+����ў_[~��6Py¤ +���
zQ$t�w+�Qg�n��\�Dz���{^+����:f�z��RZ$?�em��_`�-�i��֥���9��;LWl��c̠�<��� SGQ�-hUoWC��:�P�Q�T�*@�w�=�I�#.L��|���jp�V���=R���J��i�������;�%y�j�Ȍ��lx7�y��Z��j��A��3b٠��ix����,�y@ܓ���	�S���	��a��.>�"jFAD0b�U�UCJ+��cK��t��9�Zl��kU-�w��7O�M�4�~�>(��\� ľ�k�9I"�f�;Ѐ�/� ̲<M�`\\���&��AXz*��_|A���r���dR�t��2��w�_�w�1C� �m$L���]�9SD�k�>�v�s������a��1#�Hb�Ae2���d4��.�ˌ�^�۵�OlD�Cf��F*HTQ���g�t3�&V9��lZ�c��	[1�9X�z�����~����'���w��.N%�Ѓ�(I�h�Z�^<&�G���S�ْxA/ȑ�1��c&���l�Z%5A��@N~R�弓�:��1;��RI�&� i���>qg���	��x i �V��3cd�&���"�(�U7�j�?~�d9�E����h��WL ��� �	��h�OL�����w��a��
��)�F��S�7�]���Lq�䬇|�^e�M����a]{|�ۢ���aK讫;�&���a�L��2:�l���J�qi3�0)O���a�&��25sv�����l`c�u��L%/&�'Y>�5y�'Z��V�*D*��x,R�0�c!ɸ^-�#���X%Zo0ɈA���,9Mh=��#Y0@�w��خTx�5T<uy��=:Z�h��0��
��i���#���;���h��\��`"[й��O���i�ĳ�.��S̖��@x��g'إA{����tw29Z��T���,�?V�Z֏M���T�R�x4��m��
��T�(FXl������I'U���5A���$d�֢�m#���fδ���}s��3��A���w�����
5�t�����W 5��*AB���,E�T�����{��<^r���~��X��b�ۢ�U5��{<~��G��ue�J��:Q1Veq�f����5�����<w�ؙ8�0E�oJ*��T�`^=ss�ӂ��Dpg��f��J����4cA� iYs%��"X��5���Iw_!u�S�Wɣ`��	��m����{�$�x�NaS��n1�+�� .}mr��.�e1�Λ{���>r
�E?���v�u��34�-���#jɾ�Bl�2�s� ���-�����J������ ���XTh�5�OY"��3?��_����X�}����7���Qx����D�`C����'A�J?�']J�g��B����+�C�� �_�	�<h����g�o.J��h�.$�7����}f+ ħ�ǅ��a��뻅Ṥ�H#;��\��䲇������ƀ�=L3��X�`T�RPb�w�7�+;��)�0=��ie{����G������Qk$�Bs�ǻ�2uJR@Z:�m���v����f�����\nO����+1z�����	-Y�Km�%n,b���I����N"﫳R>3ߔ��cmU9d��;[#�mT�����m�"|��� �
��A泖���0��a��.���B7U�&H����:��O��Vz�����&��"�2���}	��(�ЁT.�;�]5�vIlL+���v��Ui����)�M��*�8�zy2C�1[�?������C&��ܣbL�ZZ<�G4ť��m��0V\�.KC�ƞZ��q p����J�|���5X��O\ؙ2,; U����7�q�)�g\h�M4Q�лDQ��������ӅtML���X��>�oK�P�'{����s0��tx�<��~���2�����uM��h��yv�!�>�$����e�Hz}hD?�?u��޵8c2=1W�m�j�����я����bB1xZ���{���"l�$#_�JL���Ejp=�n߷�=�Ln@d��3"�w=�w�"H>�h���q|T��^k�9iw�Z�h;.~����d{V��i��2c�7�O�n�;�GwI/��0?��D��
�[�g��qݏ[�2^�B��D9J}j}]X�䈗��neb�?k��lG!����{�C+��R[j������Sa�Bj�����/m�2�u.���"Z�)�!�9�����ܿ,l15ȹO��)>G���d0PO���|M�2���R�b�w�	2N��$�>ݘ���K�#A���r���ɝ7��f��vpu������IB�
����V��a͵��e!.tn�Ǩ;�w!=�̝1}+������m�@6�9��+�y�E�i&nQtZ	�]Ǥ[��P]ǒض����	��S  QߣgU�W��¦�:׽x�_D!q�$�d��}g9q�ߡ��� �pp�3�%*k���f��*��ڐ?5��avw���;T*M���W���-ʔ�Ͱfk3S@C��AuC.i���@u��W��
����-�+`Vw=XK�x�{(l��5ͧO��=�LmY����PC�	�>�b-$�#����i�qgS �Ei��c정���t)e$Y1J%h�z2���LP�圕�j�N���t��~�S���H�8#��V�~C�_�.=9E�g�3�
��1fk�	>9
k9ˇ�ܫ$pX�t18�_���kLYm*C�h��]�Ր1��u�BD�η��|�C�4rF��h1822��~��SM6�*�<Q0�ގ(0���l~hN_[,����{��XАB��-��["�x��j��i�z���z!�Y�����>s33���ՠa��E��Sݍ�KeD�\��(@+pP6U8A=4
��Ь�v����J��p�z���Z��E����_)��yi�L�`J��:��W{�.d��v�X��x1F��\�����p2�v?�ˇ �R����ޡ�%�nU!ѿ��5{r@��TIA���[P-_�$fy�؛�g-h�Yo��@�F[A�8ݵ4
f��J��폗N��]ޮ�f�6��6�V�+�W)�xa���?.��C;�w���B`�����,^�{���'_V�LZ�ѿ�:��ҼjRܥ[�.8��~��y0��˽yX�-�^���@����Ok��Q콯@�g���R���Ф�1@�
�b���S�Cc����ﱯ�֘����R�&�6繉��J#z��,�4
���0�.�X��L�vF8� $��K��3m^.��X��,}n�e�ɿ���~X���O�(�o-7k�T�5qb�s	Y���@�ev����v�6՚c�{��ڢ���ǚCX����|JL�Q2�M-* _D"��Lyo:#f�4y����������[wql����.�ދ:�����}�I��+�'J����i$k�$�+��-�!iBo���=� Bp]ݵ�7�q�u����x�B�n�gU��a���6;�982Y�8��h�}XDE;�@�U#[@�0�%��muU_����J��뫵�����ZW{�	��<��$Vz]��+�$B��,�k�9T����
��1<�~�q���P@���/Q-WQ�+��/�0(�8H����Z�5_o�&em~ǸP�"hCةt+�s�-�:��0����KU���$����`��߭?�Tr߆e?
��[~��K���>ݠ�uI;<�ʭ�vy�&���S�.���� p���[�@ny8��E]��0�������K����^p���QRQD�kjb���s�����8��ѳ�X#�� ���ʐh���R�ڴ�����#c�����`|�� �� ����Ј��w�������dB��Y�"n|&��&pcl�у��Ą~�D5B��1�.�$���3rwl�6��<#�9}�U_E��8 Z�H{�+�gR�r����Zc�:��	�P�G�'��4<F��YMre��k׬�nbeN+�R���*x_�/�ڿ:VBV��R�-t��h�$!�œ�JY�b��g�:��7��U���BoKU��h�7"���@?�,�� %[s��]=�fb	�`��hۯ\�mf�hX��.��(��C�����:��n�0]�,����ޣ�]�����(�5�������fãҵ՛��1�q`0Jux	��M�e�c*=�󌧐`y)0o=��_=��d�a4�q_d-7.��=FlC�/(�sV%� ������U%�=<yϙ���:� ��h//�JA+���.%���_j  �0;{g!��dj9&�d]ɐ9�݇��%�8ˣ�2�T��B�e���~; ��c;�O�PK<j�s����"��G�ս�[#�����F��A5�d9�W-c�,�P�g�3gk?�� '��������gRv�� +脤�?���c�6\�O����9���I�R�&@뿒 ��u��J���7�3*]���`l���KDQly\����r�Iw�P��p�jm�]-�!F��C}D�_��S����2�'�u�7�p^���!�ʁ�K���� E gPqw����߆�\����n���b���5]�\"�_��wq�k����iW�Nv#�mo���ۀw�>*�����C���~gz�Q�	�f��
�zHjh�/;�M��ں������j��ʮ>߷����' Ǵt�А��%�T�t}�Si�������.3Rٷ��U>�����rRsU��^� ����|%�^�