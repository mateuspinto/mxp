`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
Yz2MQJITfrrXDMkqmlYANaVMpLQw4MSeQ0uqKdsYJu1T8QDl1SvqAl4T5N1USr2u1P4X01Epuxic
msbNzVAlSORSV5kCSicgiL/TNjRWqMV4+veFNSKU2TdiSoPNbTxFzjVtnufefQ4gID+XlXNZBhz/
uOxADD0DE5I38Ct1yvoP/fMofmDC65Yl1OOFPmWwi8RYNXJ2Dvr0SuDvj6sAkYTdYYmn4gadLVtC
LDXHq4Z0+KQZWZbssxOVWHiCkaV+7GGAx/G58myfFKJBQI5e4qkqR4phKXQ+keUxXrEOH5L4eygB
pWLxXM8opFrw4Fl97J6Oao32I5EbGIomr4Fbe95C3+M7JF68FITGjEEv8bcigcqQIQ3O5ogDFVLx
GZ1BbullU/Bwa4mgmF46EH8wMy+LDjLZf+jZkMXoKE01V+9WLtTO5MPV1BZbD8VNtb4szbLXNl+0
aBw4vi6VXMysPBu2fj89C+Jpx1qJmnIKgLEVSCSK6LGwNQLVEqSfbbf384OgEIa6j6+QgVY54GyJ
W3Mp0ecU9bpinrj2l7u+fopCgC2DXWh0sP6Ki+YXO1XuURQICfx9JvSvAmDyiUXBe2TJnXZ7uC1S
bJvzTWSYStm+zebvQyz2DHtYYqPCa9o+puNRqI7esqi+XmTq7mcJFqKmwEukSR7NDySpf/xvhp/i
39YPRFctw3fbPYDJJkjjFiV8idC31Hd8ajfMc73rQr2id0yVcfMNfjsw+Q99KkzhCiEigvrBRP7H
7RLh2EXZavmr2wnXeNVYztrLH4+NfA/8gTvbUJNtsawWBNcBPMP/GmHCgWI0AFqg3SCDdsyDuKR0
955DYPUA5eWqxtf2/IK7fn6jVLIbyibLeF7oHMvJJqdk+8xYkOcvX1MxqvvNLA/kddl8bW3ncvqh
G5at8TqigNXNFoPIIRzluRCRlRBmX2GJbD3X2Q9wgk4AXTuB9qe3jzmYStbfNwtmUdRds17D3TJI
6934ubRLubwXdorRh7UnSq41eaLsTAIBeO5SVHLGgTOcES8c9wSyiF2w7tsriygYOOQP2P2MZfiU
fsC+umHswUSzzHIrI8RA6KzWhX0vzVnRKjy/IEqiNoVlVmvakM/mHXkoJzRQQOCjuGYGr+O3r0Qs
5XMJ3UGFJbYgBymGBWFyiP5y07iHz3TV4CvJN+n27OAtyLtXQII9oS5aqXgz7b3vsRQMaCSCefVD
Nbr44PhGv8h0AikfK6H2wOxateQD59h2YZkglS2ifuL7u1ZZvJMtXSZ2a2LeJIrZUu7Zyk2TUThu
TgI3buOlXQSimY2ug7Y7w7/VqVGLgtx7bdVYrRG1Yk8Bun6F3wGePKummK78zAReHh2fIgf8BOaY
n3LHGtDZTlyGsRBtuASROF5nEoJKGJK1i8opmHeRHD0tllWP4BilmSio5Wa2WFc5Np+6PpQHfI4p
9BL0Kok/Um7sbCNXsDcrGDisEY1HjCr/92Vwu2XDAv88dsXT9soHqefLRhHyLtkyiJ8TeAGc2zQo
P6KVcOHT6xlAr6txkE4ddNXT21Td7VLtYxh/r3yJBliXjPYjL30LhdtZvBIrwv0JDW1n3re2yAHt
v0rvGEhPlP/4s/qu9PO092t0Oozkli30L+WgWO73fDYsEcmvvVdNLeemy+9P/mYgJuaZgWBrE9rf
B9ynCJrrO5dw/3sfBBPIpbFA+FY0L7oaiGMJyOdG3QMc+tOfOBwZluiOSKDEMYaXk8Xju8usUtWp
7ZsWYP6EdNZCp/8LWxgwWdT6K4rXoj4bXz2J0HXt5JQhGXsB4erPcja3kbcdtRhssbLmE2icE5gG
pF8D4E683bElvf/Thv04rfbovYyRbpNcWGdV/oBaaSH6eqG9Cuq2xXO+tgVqnVsTDbmaOF1CvLcW
UNwqCuYgAHE/jNlQuVGoVoXvH3n096Z2I24TkzNq2q9Yio2fVyXYGAhEkeHqRSMmFFudhV8Hj19l
/TMiVov8Urc0LqQdFsA5ZEzXfJEPblpNlRtAMGUhFKlPYpW8gRJkl74ZJ3vHuUtKC1OfVrEY8CUN
32U0pMmCkS4Jgky442GVJDVIVwm68OhS6C/bzA5GXjl02l3dwW+0vJcB/CAHw1vA7eF3790Y9YGi
s73QZekA8aNhQZDyhEjjqvf5vEKhsn0uxyzA50EITG22cxQhsU2XZY5JGBw0uFas3dpKSrygRBp/
l+IIdzvc5exUpcuA6Ze+6SIuM5MogmfpUr1+mgIaSUGvetHLGwlMr+YKoUW/JHwlMFBAcE9f6mH/
iSzktpmL1lVkvt0ttOxVwjlGbBr/0UiQyqkfc0RfQjk7T4LJgUneUoJWymSvaNDP8s7lHA1+TOPw
q/tv1sPmtT6DdsN8c4p91bmfpgQEjcUl4PMcypsAo26iBbWS0DuIT+Eq2KTjWosqgMRoXwq+rWhg
cHFFTKg0gZuv0nu4a3KCHctorilv5RbXx5fyghb91zaKURf0O2JzOsJP4hCqgKrzb0PtH4XhtrH+
b0liFWaQTDhILBVuqElMnLTnqngB3MZHFYgPOfCnAaSpGZ2J5BXwcqGimcL8EcatrOCtrmYslFFy
tQWgKpXdKzsm0XE1lHuls4er39m8vhCqZMQj7SzeNSvWifMtTxDEUrf1smFOoKQ+ztOvKOjZwF4t
zFlfxEF/EsB+i6utKDWtLQVTyDJjhL+TcxIS3+KyKO8yQoOJIkcAuhoWG6WT4xEkL/Rr26EFuUU4
yhoDd22Qfj7gBf58Z2tl8GvkM7BAb9U4LCWOLKS/WZoijXFXcaMssXmf+E8IiV8bFFs0mNmmRlvW
yt1z4ax7eJHXvOv/ZCnKlpMYmdTKhYuXE8aVeecqIon6qt5DviZd3Yorv/2uGcdX1Zl4RDGMI9KP
CF0whT6Xwz1EbQ+3Ty9pX4QKyoSY+uugvT1+Wqq9GRLsvckQLu0AMQngw4W8IhCX0ExYRxZz4Tbr
WzYjE0nwh10FmPybvhOtGcmpDZ/hAZ8SssVDBXHuovQjT0WOmywqZR42FwBm5DaiYP9c5bvLazOK
iMnGOh9OIKLGx6dpv9+WZyAM5bHUY3U5wC37+sMYUOdrvfUMP7gci8Rf/ralwlz9oGGqbsYhR5/j
A48uFhaTVVop3O68zboGTh6UfYXwMtxJgk2DcWgS3pMOpdkBTVjnpwXSYJxx71UAJW8vJQLvh2w6
RnsJwhIZ5c7aWhzqTgJwLK3iX75M05CMV/68/3cwrRahi7lZRX50ppb3tPrQEKpQknaPGvY1JPQ2
lWYOERyLwd0nsQc86lVIS/UwPB669OK+nxOdl6jrbdjy/pOMbMoLv++DbMjxl3NOpf7Y5UA6GREL
lmYp+Qm+F9QLu7YY2fSCYPxouExJErV3vBvkhHKUJYTSdMYCJO4qJByv2WZIbwdwa532tYwwuhiz
39Ko5kDUTcb+6hY6hyBx/ckH7t/8qapCiW/M5+txwQZ/3RWd5wHE9EumlllHhXM7YDkr66vZnYLS
yYJGGYh5LFxA41g44EcZb/xdW9zi5H4VGGwIhMxxYcB/NzBV2MrmnxmYpYio5GtCUjudIawEA4EM
Kp9rNbSlT/e1VHbzgACcanS4jNKWCuS0GWO5rHLkzMGwqjZo6sFRvWhlkc6NImvMYuYN/aMYNXKT
/DR3aUBOlZp4h2/CYs5Vx7MXrJQdufUe8Fd8pDTVSSdLGQHXgtTt9gxpqhcWSpC52cl+wHZMIUTJ
q9Ex9jTV44VaVJYRPU5TK+/SEvh6VHPdcA3zQGlnTex9RTB7QpCc/iKcawZwSeSL0MqGb2/CVwPC
6JhknO57rQHwMBhr4VmhITTi6iSCsBAHjr8BOtzHR1c//HwbTfez6hCG7Oc5vkIDm+iZqM6Ks8Bg
bi1AlWe23ohIsJSVeGFj+xQo39gqXNI6JwbiKKDPM2yDyOaV73Cf1kqy/fmDPxLIv+0yjp/Oghtc
TsSbFxV/AONmyRfTz2YtbFEYrBo6pO8JaG/rJDo4LC7q3WE4GWPFFJLwdDQfFRqsnuSZaic2tSo5
UDZac895Ze0Vy8O5HsKLaQa9OoPdCQTNOkCLuzBiUeQsDItUs02lMFIpJGx1OyhzcJkEWy9SxkHe
RW02dcWesa6WUInSFGDmAuvW9TVnRgYXssveV+1ZT/rkOJfsNil47gz+76fdwjTXKvdBWm3zaZwB
TM28R+iq7eWMDr4z8VLTclwXX3deVhcy3PfgM/JlfH5jP6VHvis3Bon/A+5CoCelpU/QSIBl/can
wjNJ+d+34R9iZw+KngvByn3VF2r3SSiJPUsgzWPfGrt3cxJaLfmahIWocxwLyz11AG5ZEKPOzlUj
C5SOExvfSy2e13sfc0WXYBCXI7j3TGg2zJVZHpXRn2A+LNpLDfj4kx1Csm8+9YvASSp9D44PZdM4
AClcn7a0UIpj51MbfkD4FdA0ySqPtXkWLFLrubjFSSb70VKZ0nRVszVxp4fO6ssZXAbxPCswi7hG
NPmIfkwa3AHpaSIWanXzoxQvs9GGeJ0QThJ0i2Qw97pjTJD3hBoxXvqRVXu+lbVqrXG46whFq4o2
Yi5bW565ZYHJghnq4SBLhBFPuB6Qyz1S2olOYrernhAIPY5jo954TKm031Gaq7DVv6LZDGKWP+33
CWB46B6rm5PFOKxhMvC2qLukSeO+aPD/IJ1eE7Wx3aZ7fJi8+Ijo2u3mM2nNULGNN9tBcwnNvFh+
8Y1dJ9PGWQkIxEVC6d6t5RjFZXWJiIM8PgErKxAXNPJR/0LEG0gRVG0uP3bP7EzbNFncRteXa4K0
AwiOnqU29Y4+aKzyM32WAJ3+jcYEa4SFg+Xj3apF6MX4UqS+OIcVqrTZytRMYYiJ5pXcmZ3vInzb
H3QMseiulB6JTNDRzIk+KX2wN0O5NiMEKb6va9gOIf6oxjHSXrKHsb9o7kN8btuKjKo+69v7fL+J
Xt/lSxn79FDyvE3iTE/9EWP9hNM3LBWgiL/bB2wvAeyd+ffXl3MeTFS/53M6sJtBx6WSY0kMGd2K
CBvomjEVgd26Uwq3QsxdRJEc+EpZmrucGFm0wbe1Fdoa1HIwGaDpnyAa/mVKLFSXs5hYEVP1xc8A
N2EkYooiZZQCxJcIpKmK4WUsodqhWF+30X03y0PluWNPkfAkgGJy99tLxJ74BlTC0/jinrt1aAjy
VqeR8rUgpJXjTAsfvuV7O+IxfGEQxJkSfrBMnDJAHsDmOxDy0feEwYy4PMXmxvY7pRBovsLnqQIP
NdOCQY7Dw6LfJZv1hNkoCQF04HSDmVYX1/6R0Y3QvTj7H/JQQDUXT7zilCLq5pGXpI0gbz0WUTOs
oSm6O8QAEd7pUFeRv+MymfOlvHN8MDTD1srpJ6HXZtUvAn4V8fCVnjwBiN18LLsoQVXWo9HoOB88
Q0NtfsIf63ydf5LoCvu30/TU1Fx3b4ep6SSBHmkN/vG/E034jg8iK7KfkXwIO4aOWxJ5YA3dHqch
vpLpMMfkQXz9q5kfUvyeLBP9eO7Lvfq/qhk6rU2IR3eMrs8pIG3a4a6I7Vl1AyDSOvFmQe+juOGY
rb980b2rMZ2wt7RNe9bTIaibOfFhr/I4alA7a34vHmu10c7STUgXv594QLYcw8i/U2ZwJpwAOsEM
FDrEKy3M8oAZU9m5tb1W2b+6U8NO+HhsgBl/WLK/EITDEQnR4DJ3Khju7leck/4BBI++j1oWUNUx
LTS/6XbDYN1XmzCulQq1nsxnOx66hCJVZImLI3qXo0watV8S8bZb8cuXMGDAYsjmzsgxMpMESDMN
vtkadbpFlJBsiVH2eW8IC6idf2U60XiP29fec3YW6ISgQELnwEu3QIzvNU1utT4YdsIRohxig0dL
lxEfFEn2fHsrSY/DbFd8GKt+YAn0iJhxXMc7eOkOeUp6pyX7U/ebOsE/R+Wy0gV4saEkEPpRrX5f
6/uQyFI1Vdx0Xx9p+y/K6fXbbGhMx1UMxIBF//qbqtD4rJUca3gQCSFwdKsUkic7rhQfsyzeI3YU
K56D/ELjh4ze6PK2Zdl504GynlIEnBh82zWet3iGiAQfk9JttjB9doGdatoygxZBz0WTtnNC0mpU
8H8YgNWouDlwmfa6UdRsfolysK91EaYKFkzX8Z3BMWyz0zIJ0cFbve4V3UrS33+qZ5a5dss83BTv
BJW2ujJrH0Bg/ZRZwkXjdsdYANCYWbYSWu50cBmLyZhuMBT3rrfkURsB2V8boFu28/9us158W48x
Vk014f58p5BgLEAgdRX40VCKKD/5RSpiLaLZPJsgL5D/EUyomL5AniMJQtwGiKUSAuzgl/w5vukC
6TUyvkqoijcBEqcRA9dmZORjO86ilPhpuS3Z94BgmUG4aeOhlvmknUznW4gJeEuTEU0qb1ftQdKx
2Uk0Bc12D/L+e+F2vkK01lXX/xy3SKZQEwS9ORD4cJdc0My6E/AI9ulwuYYuylw+5+JM3RiByyzI
DrlYcpJCdvQKYOiyIYHkhaW580Hryijprgjy9N9hWGWxvMnUudXAd1hSnL9QJfdwu1lrk9UnwEqQ
pLKsTcOQH1KtUaeea9TetGhbW1vy2HGd23ynBlP/VQAslk3QQXcuXdDnvNtY2a3TxGkQCzgJdOVN
CQIgbY0XAVhtroOJqgE/437BAXUSCCpyAJ0jS/wlc2MKPt02c/sjssULSVA4jlzL0PgPLrTYSQVZ
eA9ralC4hZCbYqqfZne7Yh2KPi9sLGrHJQ8vsWhAr+MTSB531+UczCqp4rUxwl6F2atODQ1AkTgv
lcASvzREAarZQ7BzRVN2Aze/0T824ii30T6ZJXJwE+MNG68lRjb2JeB8zumEUlwzNbGfd7jJ8e2a
MmQN+zn8ousYAx0b9f20jvwI184YnCG4931yq+SuH2wjlqyUXuo+E1agURGDNTZpOyv5drXo7/ld
rx+HvW1rZkk5Icohp7tJoY/hS9ZT2l/mXkBUFL0mDOKr8cHfTl4Wdj10dYX82hn5g7wvAwx0dSqX
/ConafFnBYBtVSM++VEqF/HFbpfjpa0koa+hIOnX6Q4vNs1+8/AJEz8HM+D1ofNAw2jkQfoUu4Ma
Xxn4vBGgWX9Ono67qXxIDE2Ckd1VGYuV/kSXTwor3XWbRfLodFQXhFY7me8xB3kM1afgAlSPuPTz
ZA3ZPcYjc4BaDhFFLFDkmJW/LHpMWp3vUlnWGgU+bupGvk1p9VDFSmOj9jnnrjopaQ0YvqVwuYhN
0TWd+hY1qkL01qMdnDgflQnR9rog+jjFDH0GBUUwwiQL0NBU0OYRUJi/tf4zFe+unHBh9y4ibdN7
C1M34AqkbHjsbxaTVdlUqcGCoGxH9lpUE2zmkweX4HvybAhrCeaLyTbzKrWqjh5dMq+kXztPwVJP
LfDcq2PfvcSt4QlO43tjCxUNtwv0pTpT/omiTRaMiAO4r/Tb7OrvoBMy25kcBTuIbZYF4LNT41yB
j5WbQ0tO4wecojoysslKFcm8HImfwv6l3ohfGy+TcwZarAKY41W8c/DavBfc7QWBjbNBwrJZXb66
bBGU+4EvGYdspVx/hOfds6uzRdMFVvqVKuEScyX2FecqWvcyKsAYIWCItl8DmluoTVa6YGW1ty1s
tcprjEVcdnKB398gy0EtNRn1iNMTjbrbkjDdpnwCGAT222ae5zINJpP+MVncQPxSx5uwWo7s4+6K
2QlgwCZUcrj6/LfUuTRicV6RvznCD667hZKbMHTZzFenvQWoOqHI+wqhClmRrsI2La/o0yYMMKEe
gPvg5uaJ9bAW/lP5nF5RJYaZntld99Sl6THSNKDQDDJh/G9OhkyA7OhbEfsTQ4hRB6MzxHAcw0Uo
sTDv284t/OnrYomvUrMUYkogd/x/pCFIeHNXA4kWkUssxfSexIAEcIGhfOCE5CP7O/Bfo+IlMudG
9o9YhFNaPMkoxhQd1UMtChFD1/ZFTuxg8iZN14fy1ru6aJ7dIe6Boi36YEnnL4SMY5Mt1rWNX2gB
k09gFqvnSbpyZFfySqeBu+M0/9MwnjPph9jUaM5iNbLy0Cj6gFQeU+2XatcbGGqrbcQx7UsS5/Ii
YO7aavLqFDpdZORxF05q9Vz7IIvXFYAmkl7ki9p8KTYJWI3DBU0jfrSYHODjOm3u21jTt28UkKuG
ZTAuwSIY/2eKcFVfSQP8EAzELUbWhNGW3mnyteX12qNTpgT1lgQ7ohgvDYA+VhXjd7AV+tnTgX6m
XxOC4HUJgp6y3+/eVOu26T5Uh/sSUYWxDI9fEJJWmhmPCPvZsWxnCQaq9614RLRClHqxXi+ct5H+
zvGTW/uptRbRcp+ldvX/ocSah8k+o+Zu5FBPagBB6NrOsPorXln/Ysizsg==
`protect end_protected
