XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��¡݅z2�&"Ո�^�ނ��9��$%���[GQ}�K��p{ �����t'X��������V���{�<;�wZ�M2a�AJ�%x�[s�ְ:�Ý�6e AF�.y�8�_1?��ʾ��g��V��/@��$���qpD�����Y�h�D<s,��0��IF�mu�7_o\X
l?�*`�jaҮ����e_!I^;�)�T��������we�bDwh�.+�	�6�Q&0���$�0Ut��7��� �����/4B$f�Su]�A���5<?1d�R~k��Ș����2<i�>�M�/)��j�2p���C/��C�Fu���I���o�\9Q��5��5�w��x��D-�d�W�[R� �Rf!����1{���[�.��aU���bDw�Ȥ����u�j|��d����
xrD��*��� ɾ}m�W@H.,��_���U���Q�2�t����$lB�G�0����H���cp����,(����iZ.�p!�v�I7�y.t���v8y)�=GU&L �i�sQ�z�
zҙ���,���������Q���j�^����eE�Nџ*djI_��o��\$�g�p@�����\�	������q"a������ք$��
9hSR����Wui����dno���BهU�j�'���#�`��D0:�˜�5ɱU�#P���C,�®QA�����2EaN�o�mx��F�|�$�ߎ�gI
K��{ޅ�S����:ԗv�u���>�	�G��gNt+kXlxVHYEB     400     1a0��M�rl�6j�JGu��y�Er>n��ͭ67����9(8��cY�ڪT�J �ա����$ў�	�N�>rsݭ�+�W�e*��)^���hkf۟�ñm�L6n�rPEY��)��$�،��4{��i�"J|�s|>�_l��ŐB�2�rP8�2���A
���S��3Ǚ��n��������UIB܂l�P������n��L���u��M������,U�J{5�3a�>'��~vN�NД���V%�qQÚ	����k�Fu�u:��FQm��x?�f�$�.h��hREd�i��෇�L���m5�:O;a�>�B��O�w�[���LW_v����F�����]��*��`��QLt;�UB�`W"�Z*�9�Y�fsc�X�����O��J��:l,a��O`������H�XlxVHYEB     400     150ȑ^�|lV ���G�ä�־n�Bd�˦�h��ݨ1`�����r���G%o�F�����0��i��C�ɀ������=tE���^HJ0�D�[�@��Mŷd�f�2~r^a�ƛR���m5���� �z�q{�?wb/v&�D��mf��q��F�;+�/kv>�ˑ�ڱu�=Z�ܭ8a��/�҆4��O�u�q<��S�-$Ҽp�{w�xoACŭdt�S�[W�
�FJ�u�-�%�]<OH�g
x����R����Ӌn�d�W�!֡��,�i���� -O���@��(&�|�e������b�OZ�H�z��.��]/�\Ț���KC/��nUXlxVHYEB     400     190Q'`!�z���`O]U�!ZHw�l���(��<\�Pw�.��-!�.�2 ���3��Y��w)��{)���f��N��(�	{�7(�]��5�: `őOL�:p���)������Ǝ�����m��јVxw�����}� ,�GI��γA�=XD�s#��-���/s��~������=a����d&�Y)��v/m��e&�Aھ�a�Gf�t\����#ǁ�'��~��Oyy�~P	�}R�y8�}��,�c��P'��	�\~��u�r�evC��x]uP�rz`��-v��&���?�SW���祜%�\�=_�����wmٽc����S�����l-� Ƀ]�<�T�2�z����S�wWN.�(���\(~|e�w��H����\���XlxVHYEB     400      f0s�L���Qy/��oP�:=$pB?�����~��b�_E�M$��*�P�����X�ŪH�H��Ϳ�N=]S�rH:����^�g�L�a�6�ko��~�xL�m$�o�ߨ���%�U�fE8�${�oA-�4\�f����.�RF`��p�	p)���;�<]�"-p/V�
K�Yu��˓�^8�˛X���������z���IR�3i�s�f����lZ�|_E:Q��/�FfN7XlxVHYEB     400     120=G�w2�*�&��aн��``ΉW�nU�`H/j�2���7mC� e�D��u��+.�c��iT�x!�1���m���������r�bS9���+%o�4ා[�PB�~2��{<�� ���z����e�r����"���ɬSX~L"��W�:�sqJ5%#�?��;�"g�iH��Z8�\�ka��L֭g1��J	�P��_�p>�~�t=��k�oc?�����ā�ʆY�u�ӿ>�z��o��J'5?�K�����?��w�T��H��9��`賭R�4XlxVHYEB     400     150n��ЉBk1Y5��A��j0�.������=0H%����+�b����g���?��h6��`�[�U�m�L��SP E���%Eg{2�mn���\��^3՘������g��տ������=�L�Z�}��3v}�I��q8+zG�����؛�:���r�T�����Ùņ�pkW���ݣ1���p�� �Ω)���@4�s����c(,Rl���Lg��}k��G|:_��F�Y?K˙L7랷&C�\hbl��Ϸ߯w��گG�����!����	SB�Jj��M�=�?yaJ��?�͵�O��䈛:�uXlxVHYEB      ee      70*��$;'���>V�J������{�@�a*��L�ֹO>�i����^O~���?F�)�4��5����Xb���.)�O���\���'�PGD+�7.qR���oe;��9�G��yB