`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
h2SaClnF7mJripMfda136Gh8dsWun/UUzVjlS9grcJbddijCQMTABO4YsqeubcTbLe2H1UyLLmEx
99DSSLtu7uZ5fqWtV5qPlirNfCsnMNvrm/A/e+i3BJ7jm3tfl6iTUYxetIe4Tjx62YDhwtJWCAkR
npHlMV7NToU7MuvUpeaZC8J+/SLoM6OfTVCeozePJv4Ki4ZeOMxACgvxW8oImgk7IvvRIg0DtOTx
s+zSc+m5jHwG5Hp/Dzh55aVkm+IDZicwVxwvkM/npFHSAE8xsyoEMhJHqKfJMbFeMHCbHVgGxWp7
QlD7Am1AIv8lXs6Xji2J3Z5lifzWdo7gTfsUjA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="TVS509JqUptsZgrb1OEDbyPKRtVfEj51k7a1lCYszrI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9456)
`protect data_block
ISFcW0BAkkkQtqfjDinG8ziQjT45AJ+fl9zVgvIqQj8y0TEzIY6E/xNZr98KV4nwK8R0NnHjAH6P
jo7tBBxR1z5dfKGPAw8K06z3LDXvrDhyIqe6/vcaGru/WcM8rThTGwtOs89duKDq1nZLE2u7b3SC
+QP2njVAJv1khgT0cjyBidllXIh0EgeGmoUXDoSiQ3gbBQS5Hbn08NOBJG9escSWh9hkQt8ig1ig
4ddxoRNN1O1u8RDL2sPvX5X5l/3j9qQRMOarNq8w6Uz9pPIyzXuuelT/1FP7CRhmgE/MMJ0WTUf6
7/uRdp4RlUCChO3O/B91OFL4bUqFZVsobSkXWq0OsuMcvGb5XEY+R73tQFFdmVlLkVarUtBQxZ9x
jJyhSVge8ni5KVrUOH4YlAHSVZVcbhQOrZSvGq3Uyjt5yRKue05WQQk+ltk4ZHPqDlmJ6wmllJnY
sjs7fUnm0oYUV1Cs/9p2IOIBO5mSt3bOYc8O+JjVYJPcuvDtFh8ToVJH6KgjT4GcQHgQ/VikuOdJ
aBBhErs8RZGPaJwF84Scymd23uFqUpnUQUNrTIwO43A+6CJy79P0Jn1g9sNJBYPHeTaX+YU4nyzn
al8ApbzmSCqWetxjJci1Vp/RL+Y/2EzyR9sLTtFuHJzV0T3oQLjJ0sqw4EeiBKq6RWbx7b/Tt2Z5
c7Z7ewqB1oyMr5gg2qY7Wad+3HpkMYKpHlofRsZSJDOf31C1tFvw7QHpgyvIAxz/6iMysQZAw7rx
3ieuuhfQditZb3TtXBj4vs/z5t2KR2kX38dKLgJahibLi6PB3yknTg7mIlYEwI7mOR6cI6GhNmVF
lO1/Oa4XzehZ8miVmnomQPdlUd9nN9IEUrUUjGtse+xI/sRVtd+pUa18Av/eqqg3sxORfSLO8NBk
XpfbxNNls3DWizdo5Ze4M9JaTD0fiDVsKuGJrIMW5iwLHJYQwHvCnmWAZjqnvfRp2mNb0uSiCFoj
j0FHwg/B6vO/pOqUoQasy1mnsCO1yO3RJUFf8Vqcy2CsRYM97H/7fXqN7lgwNLf12dGNO5aJUNCC
SP1OTXgh93/WF65olJWppx5FyagMaWczY+zX5CMAJEcD0f6dYXlGfWFEJAwuxIvirmA7VJ36Ew/a
2VTlD38NRI2MAP63D/jiKkrhfhJ8ZRwgzLHOph4cgs+qlhViL4QWUvWma0zgqE0FrKxCXYrIx0UV
5x9wlZ/1ffXYVkVSEWXHyMH7hpaQe3uq6UFrCnmLBhOdszndREUKgdV8eQofeB7ga9adFd8GFR4u
u/xYy2DeybhKnvW1eBAJMw0PwNh5rtUhKOknqhi60sFYTrvQdOg8oJIIwijAYr0A98uDfrVOYqYL
8eXxt0wfs80IrgIlsdDiCywnVtZx9dsDd6xBeQ6fX9Qx0ES/ZyGUhEszLqZ4o+tGQ2/bs6wJJFZe
Sk5JTxfHdgwI5QE4qE0Lub0e0jsr8rOLf7B830w4Hn2xT9sNR1S1yWrqnQcrtozX015xKrLmhtBM
lOdWN0Z+6UtKtBompCIEYGM0vNCGfSlqO6v37MnGIZ5XKASATLnL87p3AFPGk6IHnJjdW5F0gEkH
RcfY6MlfqiRzFyHhbqGMI/C6KMl2ZxDGDTENKUTa2sNsipFjFKYI4kAex6yfKQ73ETw6vvgvbHue
Y9UEZP/btRhvFobe8woB2gT9RGIvdj6n3chqCg8Sh7Mq7EKShkq32qsIKcHvOxHTYGCwhhCZhWpy
UOxvDV1fQk2Ru8F0VVJd9IaE7Cc98TjW+HAMjrZCeLxIyP9kSNVdNgrsnVxVTFbKaRBSkmulh5ld
dlW5yXZVLYaKf1p+hkvRXogO4Y8vS7byvqWnu6oMIbmAsnUNNyP3LHyFzt9XbJ+RYalt1tLhtkNI
5JkOLlyu7HukXfkFxXKR5GgjtZInWHKaZ4u4x3iUteAs893kLfs8Sfcw0TB18+ujrzbkMZ3d4PE0
LmpT7HrcLGuz/8/Rh3/3BoXnyvXJIIXFhwPfwclGplaVn/YlVHl6zE8we0dderPV6CZY7cnOHsH1
GKeU7j35Lsu+4RuwIgV5UZbap4atnYx8bUTAW8V/5vpWXoQmDqbxr+t9GH7zn5jQMHnadHIIQv15
nzdiv9YpIXKl96CGI8NsYP1BngK39eVKehhgvckkB67ydTOFQn9aMNM89/tTd4bycWJXQdzZLPh2
sYycuwm1ZtnbTiuFlNxy3viZsHk7sDmoFqb6ZCdVaY5YYdprcEM9C0WvAXjWL+kmCoWT+mPQc8jA
92m/nNJ12ymeTQcpycCoMkyFR+cz3paYcm0VDKErs+tRXJha8iiJIcFRYxAGZM5xaz9km22Db/rZ
/5F3pX3UkYSNRG4AlCjtoqOcAAP9b+mIfuwqQ+tmO8eygdtndmUmeDfNHNjoostTuC1bvk3GItd7
ZKra/o2xVaJfpkjpKaRTVVZU0n8Ww+OzBixLIkxnL0TxM51IigCci3BJAjuYZ2xsm5lZX0aCQxT0
nZf8zeCE9HO+4tEbQ8Zas6GKcERdDyKH/iqJOfH3D+mbdUgx8BJI1EmjnYP1yahgLmuga8PPGp20
k0FZ0OK7QL6X7ku6bf+ZnSDf33YbUyq+txdjflS4JbwG8kjqzu8m3skFpuDj4U1O4MgjmHq/dU7b
Eg4So/w7A+Iqy+eZZlxGWevsDDE6+nQ8pSrAkf2HVvs/NTEEVm2gUcdEkZKZOkp1fbyKFtXII98a
8v6PWtjasKs1hEdaJ4sIJtWgVBAIIrPbwLCCJlhDLtUWWBC+ij/MBz3PoTDjBbipVK8ax0roGX85
zZozoMq7ARsKzCb0kDI2DJlCWKsOX+V/KFKLeQ9ndL8ZOhXxovCmqqwmAzixivz4dy2J1ptyg5D1
H5RyxMSbyLmDerlm0iS9Do6Ipmk8eG+Se120caXZTLi6yII3If4eCeUEQlSSiKmwNy3Ai6PNEkot
7Mqc2L8Wa/xKJV2nyFe1dCFbDMPW8qJJ4xMczpeWUjkNYKY9e+8eIVH5dnWHo86QyAQ4vyphH+pp
+9tlG3IbZ6L8uQKTYtdheLVq2QmU9d+JKZfRf3jRhronpBvE+dMglFJRJpAmeEw4pfQwfhjI9xiZ
8/TPbGFGW2DwZLE4VbZesuh3Od3IIdaeIysfAvBGtoHPxg+OgsCMKPnuTz+WYeUZ/0mD+IyRnVDh
pXSeR08MeAMbUrQJOIlfwGD+/zfb1VBEHo6gD/M56o605BmpgLwfWwILjxk5yDrZLcJKQO8isRPf
d2GmOl0AAGNRgMCKxfEqRW8sV+L8rBJo2hRNkQBK0S/dMld5RG0U5oc+vmeCWyIRpsiVv03ebDKA
iyPMZASokriwO8NWrM05sIKZVdkrzFFBvq/6QJeQaY//e+g1/rQJSFN/V3Z/FH7u6jlasuDDBNn9
Q60Djz75lL+wvS14P9P7ff2E6WtgOiX2MsW3AIREeIAUonoBstnzepu/Z0ND9GgTNgL1iq5te0yV
S3BXQjrfWNb+gF9NaTxt5HWi0VdOS9IeSzrrxmkq1p9SiOTrDe1vxrEspm3NvPA9NMggaZNjTEuA
iwYF6HcKejiFJC8R9UlzI99fstkV5qQhOIP/gkCgPyHT8WBlBBhPIoUz56+peQ/phVQMYCkI2+Yo
sKE6UXl3hxij8tjs/McpK2XrKn5H7IIZtx33Z4s5fo37Gu+l8DIYO4PMG5enUVmDrvnxWbMz9nmV
xfqLd4mOhiPSxxMPWkwZc1mBXWoFUtCJAAlglcX2adaygVUqZO+ttb97ALEZEzH07eF6VbHr+rst
3mpwWGqjH7TbKfjLGzU7pwX5qojGeEN0OYZ3dp/s4y1YAoAoXub6pN0mBV2KCh5d4dxpabSTUn5C
GJKiKZR+g3nVSW9ORBbHsxa/Vsefcb80aGsZTP4mimvg8712C9Gyzcaw5JkAbRF+9sGcf1v++mE/
Hj97ZP2Nemao6MctSUYIarBLEMmz8qjubcf+XCu+O4pUWG5BZNEO9qm0mrajw/3/uAVees0XAeG7
EeT5KhtATGd+vkCwseIpeEo7AVx6Xy1yk/s3hFC7Cd//jL/X/6vg4D90xrODY/iJWVzHmWkZHJRc
YZHiFg2BQMDA26Pp5zBzacgfIi7r4Vh7LdgFdKvfcYWCU/0cRapOEvkbLBxj0X9FyYmaYxRZxbEN
7oBfSkTNKz+kG//hMoejToELb+FwfN+FXvLUf60ApyiaEoViOIpsggZSpIyZLxT5Oir1UnmaTPJ+
KTApfzR9nBsitxkwH6XhsXv/U/NfpJL4g+fnJ2C0UisGVnu9qEMd3rVIVhs4ox9QSMT2Vj2u1+8d
J09BkvLzL3uvScp+NSAuE+BB09UbAo/QI9f3W2KjkiANVIHgBa7wo5r9+CjcrZf/ahbzRcwlz5eK
oOeRuU+41mk/Q8k/pW7m7I+RVQzi8OvFJFEZQc+b6FIphhkdkf3bpqiYQ7pY7h0WVSVKpxiUuxNG
4qe2psBhVPrNofgB+ro1JCwfJ4tEYucAW7TNkOxblQkMb+Ybd500AmK0Th0wHtS04vpQ8lZypvna
KtDD8VtaDepzlzsyeyeXYBrvIif3T6HFM/h1nPSUeut8gk7b1TYB3XycWSXusdr2rFAGjhE8Es5R
Co+xREVfgd1c0Kk9MMyp0u8qxoBefimKP8nFf/kAb2MzXjjwVges3KumAmcrM2D0XUD8dJJGB9q9
7Lk8RCZeDilLAOfOfSaAH8V+Q0bXJvOurgva9MXIZEi4rIMYhEAWe5Cef9Sb43TNMM6/vwr7ZIBS
eXBgDPZzQjky/KB8/IYV/QRx04DVOPJqn9ZaHCdQ7Ug2clLoqzsl/UFCEDe2xjwrwpgc3Hd87rAc
gvAFr2x+iX108vr+vLuVIplTpEBqquHy5D672NnWqbbuXIi+Yx83jYJzel4q7xoldkWkzipTqMmW
qNUu6i7wU84OJS6DiFd/3aJCg6xNFNTjR5oMB1AKkeidMTJCDb6hphQZighDuyRLjG1jk6zZELTK
jv59Dk9KdUgqMLsVCapZKwUTuiJ47XAgkYF7KNWauCh6qRbeVLYLKxCLaBzIjNkkAL4Lw9ypZV4d
GcSn43YMCfEzewstt+7//47OR366y2YoPYuCFv84d389XyY8S6Pcj3U218U3ZnJn9kOyAuU7qXVN
9B99nSQjcpuHibznQCc0yj1y1SJkd4dgSBZj9qFWwdASnacIF6/Uk5J7CDXezBQrjMo0Xz3m5MmK
Ky6zMs41GAnXDwoSLb+qVcuPZ6tYpTyf2ORzf8tLWzYjzViglvZnYc3TeAiiapgBUU0qTWnzHB4M
fDWTkxVdpNqgnLsxysSKG0YeIK1gam/82G4PtyuKbe6Q1pdPYddp6U4c8/D0b1EgDLhOFWnxB4Kq
1Gy1LuT8zGeCk7byT+/TN2bEu7r1tgwGRpugIrvrMCUqwAYbUPr2mlnEK+5rCaCqglx9eECcLZKb
njEA7Es27CW6Dt5J+5KGD0Z90WUAxX0ed96BQP5oqB+HRmsWX2kOhEi/xyGxBgyoZOgjwYhW44h4
82aAEvasxrZJl8Zu3E5quQHHyj6y1NbvqFrz/a1FlyTi52IapSx6+5WExl/ZfS//3azpoiMY+eR0
3+9JRMLl3kiqVr1DWkpgn4Qk3GQYVMSEU6Vq7kMBVI7s97xUyC7qyHs/qwvMbSGuRqk38L/wiFdG
I1MwymcMJuPHkYECfB272QamrQbPZZoOekcWSJQRi1t+zBOKk5fh+xvTVvSvrGyybIFs+NvyILTc
z8kCIpRFqszYlcws0yCyS6uxezqsawLEKllH4PtK1FG0HMenURw4GeDWR0eK1H1nBOT0TF6KpCv8
F9PJc/jEkb4n6vvO3wUDih1Q9+l1I4sDYYHpxYid92KkNYsXJRabaGbCbEu0AbwjIT+tpuiHq8om
PLZw+EehucMafki1J8dA3moSf5xxtnbqgvYxef8c1ansrnWvDE4WSKfv9VU9k39oKtsE23sy28rT
twYifReOpeNOdIcyW1mlM9IDX2kiXE9DojXZ/uKZOL9Eza3f5Gkzod0y4fnXZUPLriyUdpvof50I
4GMKc9/rCiPhKuGOyrFCaQiJlb92TqAmaNPP/cm0LTd4aYKrW7pb13cR9CcwGBHzyNjjY1ipaJOc
MjnRecBnBOK/5yXSQiOixXQ9jkTxhlqD40qB3Hyg3scrryG9MqAQUnmtUQU3KIBYJMSmXophyIYe
428qIsHaaGaYI1+jxjaPtOe3q95ccfD6dFhap8Hms8UT15F5/MuHkHQn4U2iM4/kbFoWYxdVOyL1
flsww3AwGoYpvjI595sZsyD66gRU61iWplkQGz4RdHALGU2y3Y9nyfNEq3Wpv/3xaKudBr/ri0z1
3ipoexnoIs9epJVyfcbgS/wZpwMM8Es6jLe2Xe9IzrWCegMDC/3i8ddzo0ZtHiYZqkLLEIX0omOD
B+z7Cx2dYxvuf61aIzboCGMVhcEpld2bNP9Y7uKCyXswVNu0VuIXVlmwwIRm42JWQ1sj2ZvKFAPa
SR1dYsII9RoofPY4yUqu8LTLfoKWGaURrEfhIKj4UlQw3YQIGU8U5T2fanv67aJjUAaL2oj7ZMu/
G6Hhutj/S4+OqkPy74ufzZGbYJ9RliN6T46X1hRSk1EDULNSu8GFbVrG+oAscQigDtWWA7xMNC/m
LJnpXX3hwspqsdjuUtV5lLtjl0eftYTI//tmmAN84QZtsqvqXpeKsvaN0MrJhYc+2wSFDakA7k8x
iCvbGcY2OT4ZBhC1PspUwYnuAKgXV6ruu42goCv43JqVrf2lp+0Edh/Lt3a/fAYH/8GiLoV9gFTu
aXcjTpGwkspLEQbod8KssOqVX49PRTB8KeRW/jqiXR5rD8BQQFhafMEueq2f2C1VrHAhFRhecs77
WNGiPg2/kXtk8J/vFyzURkj5gM840R5nP+Y7L2Uamwtpsx7zAVvXypQJgBlg0tK7V+ZJ/SvnNvoB
pIDVki3BbuY9EwH77gCNcaH9e/8vqpcLc/0/knUWamvFFMMqIu2Y2ya+e9fUBP254lCK2pnA+y38
kyUcRb38h3ZBu8tJwgsvEvpscadqCfzrOrwS4ytBcNIgd+oa/oFRmTY6H3aGqs3iSG+O8JyaYSG9
8tGZ6sVoa5S4+nQgmLjoyOdSYKqWsDJv/QCGUXMPwZsr16eq0ebjb5e25txM8P6GUTZGXOF2VBht
53SGN6yfCNPBYwsANZSLqhXqE4pl0RupoKSWNe7rDN2bZSa9BNTbT6q2m2yVApR4qXAgUaetMyUm
fhAHk50qfKpqU11p6oUEX/cS6BvxXewuZdxzU+8ceS5SBMeiz6uFr2Qbsr6JsWsST4HBCgNjO4Hg
OLLn9UJfcJ8yPUVEKPlI7ZycCSwvzfxca+k2uqpW1ao/AkVAD+r9irBS2h4SUPkAGD2GN24ciM4o
CX8+PKyNs5oXnXtFpHbrXrDnY9S71iYY50/LVeQt7gVTTDR+LjcNIZFb1zxUnJmaHXxPhz4fu7Tj
S8vgo4uP1fQ9XTnfdWTi6IgEE2IVJ08TqOeF558JfDou1nQOy6l7JOdJehvnJzTywp1FOi0+vhej
VsKYw7B5MTHkXSQGVlu3lfyKi4D9M7UaHT35MJcAx11SCDXIlGV9uxJYwmGGIde8mbKhPB0OV6r9
y4934mvbC+TYqPGZhjWOrWOdQWTXJrWKxKt/p7v29R1iCTZCEt80hLL4YYLh65a4jS2a6roTIAsV
GSpJeYR+DpUd5u/igBTAJU3ukFT9OOrEmPO9dxxZTC7WmCKpSNHyGB0dDF7B4ueQCFpAxhTj054k
KB2NtjjTssLWtA694+abJi0tFF0cEdFd4+B4AL84U8XllbrOGnyUJHNZfZ5QnM60VAxGZkYDbztF
AXEwUJhahz/u4qJO2GbBYuZouPHU+KilggioItcSCxrLxbP5DMmgjZ3Nu79K9kXRuDL4C1CFExg4
NxsseV75uB2fs9bk7ohMtiE1pV8uOvcZ2oAwG8phAgiH41m7JcOFPgxxaM15Qa6QQOT67EQbb7XQ
M68iuRQcMXTKgGrrhr6oUvGtnXgEpmccxod7Z4sIj2P+P2xJ57GgL6DLcCoGt8r+pY1z+Aurs7nI
nek2TMhSa3p9u4d6Wm7Jsp++MMg3InacVc6tJEPiWaCzbpaMnZMy1OyThRq1GOLVLiA+N5bgkU4H
Xwz1OK6X8/ZH3zI9Po/vnmTsdWcmUbroy9qVDNkuQVrSwg4eqzzM+8wmmuW2m2Dvvi1zmVWqwEtP
2Yx0fuTluMB0ykaUc7ziCWpSWMqLiLH+0F8mZUeuThEogtzhcY6fM4+tcfzRbb/TTGG8lDA9/Q2I
mTFrG6qSoG4xJRWydm5jZ+s/N3+5Nv33evAf2CWgM4cq07azaACg4Z/MkLRtojtMivlkdtNxHizh
a4M5r2OkxWDpdfaHpxTjQ+MCSGgHe8tloREyGAzHRRkS0TLo4BPG1VhbzM8SZBnnhBlUebMyz6b4
+8tVSna5tATGP582J2iUWLd6w7mFcxhvc/iMqB2+BFTLVGFEotQYtA41mr7+gQz5dGAh9pv8XbhG
hEpFwxXMIBjsezm1w1FYwCi8gxK95TAE4edtnBLV53w+HD+zTn9Vx8/w89iyqIaGJ8S3rupUvApb
5lxpBHAGMgUNnTzQOALK37DBVNTq0RAg/rtxnMRU4+kdwbP+OCS8/jJZJork/302N8ELAOlMp8BF
cs6qyEoMhVaAw8J1RB3KQkFQzdQRdmt18RHviOb9H6glpFDCWLYVN0vWETGKUZJsTfkoYloZPN2t
wW1TV0eraEbDHVILCcb3BTltka377JY0xTrI7K5khgryPbOGj5tjZicsI01jM0srlWmglI01AkGA
dfiVkJ7JNdQsMqggogyo1shz5JVU0CDxDD3yacprSbG1LbrgjBdePsDQEG67xKbvj2I/zX9UrBBi
YDAHFeleY08bwVpNoFXyVrng9iOzSBHfgqm56/xB8b3zpaAx78E5sHULbzP2yqEAR2jTA7yUvLl+
YZdZDRW7aogesMC5vpLNrGQTUzKIwby/jj19ZL5njf7BcZ8JGYs+LDvDM4sKctY9SXiO0bSNVQMU
SVCov8anf5EODFpSym2LdA1mZLN7sLQLd7nJ5xP0NfYLKMdx3+d5Wv9mMTHMO+QvF4wWElH8htSl
XE26IwjOpbtis8VTf2GatNAHtBKPkK9hH3hqO+iHvST2uUnjP7isoPsIouMU56F9HA2Gyb5rV0d2
8y46wUumT5QB5kHMgwA8PaOkM8ufgCQrdNQCCu4loV9yRWQQ2y62uSzMH8Qx1hf+snEbmOtLO/rH
rfSx66876kh5drZqmln7Pana05Z+Hb47PMsxiJl6wX1r3cHmM7uqvNMPTn4cA1I7Mb8q6KfXF7/y
xEuw3IW2OcRKuqvTQjWJR+I4U0akyVarxOX0DifmipaSIHmcKRZxpdCHtxet7PHU4LD9dN8gzHIN
7BKQgpJIq5GTb9rOhOwEi72DO4QPmHNmFzfKbhZK4WiBr8ME5dD2Nrz5jXgUf5r8f0RxV0MAq54Q
F4rWvDQ1ageRwz96eEKEYU6FHIGmofVjXGefw1/NI16HHJbIgPRS4xi8AARNBGRlXp0Y7DuohtoZ
NB9Yy8XxqG0BcNn8VCpOQ/tZByMTphFdJ7e6MUhY+M89Sgjtbd/yCBDXX6eTwHUEt28+fo18/kZl
4m+ogTLOpawIt98rRfeOv7O26rvIxBuZRbtSq8ps9l/1+pkE/OE6XyghjyluXTY0fmO8AOuaUjY1
zg91ythpjE0MiKO2+C2OjajLeTb/1VdguB/qtUuxaVOplJsJvdypFipkpSS310M2qtBbu57MP0t8
6k24OeIjBVBdemshC+voatL7rlETLlRJAshfWGExfAbFaG5LjRU/5H4ti310Tbgay9B+/uYvnrAQ
+q/34UlUPW9pfHpSh+5YRdLsBwattoFOOt7/oXicNSU/ppUukCoZga1x7+ltoMjDqJ7lp7KorwSl
7HP72Xk8cz3Jg6GyA1cmmpMVyTJv7hjSXPSKbhNl8Q7t/g/3SsTm6yc0BfQQI5aX3mhbjmPmHBz1
aC0MxswCwuJJTj4gaHkQNdFj/v9mAqdT6lmWFvkHJlzxNBmy1toLx3NePDbQv8n/tkNNSXu2J5gq
z2q7CaN1CNfhqjvcfKgUcQqVxEj8o9tDLYtIctwASxdBiU2NnBhoyixNY+5gf4JmuTnZcTYj6wgA
9r143d/WeyIdqUdOdm6dFc9QllOT5siyLhtYgR9KEMa99MKAFGkUrms9AFkgIbjhvod5WdXXcT/o
EmNyAegeoEE5rYnJ30NmUrKs+iuE16eTGG1ADNRQ0G8lyeYvvPJWpKiJDk3rRx+EQJQCOQngEDp8
00JjQpw0esakZNmdawAE/qdjFg+cCLyy23/w5ZviATZ+HBD0yceBs8anfVSuQojTqz1DDJLn692T
Isk+pWuAtyXShrTta6/PHYjUN9leYLtGt/ILg+kg0ylLRGE3fgznikCsLHICSFRMnlQ3jhd5L9+H
yBG/NMg60XUqecOUbnqnM32RVBDyU2/vWABqZ/9BX5RXR/+EfDsyo9CidvvpB2TsiW2/b4atpZHU
qr5g0ZzdEBvS2c1e0grSeeuSG8vAjB4NffIHpCU6A4XzVD3Ew/w9wu0/n40Vgaqah6530uIVMvOL
QrQ4r/By17Dz/1Jh6xa6xVWW7D15mf8+l+hL5a8XqpzVHJqtiW9qt9pz1X4dbT3+XX/QFGTHlwv+
SdH3THjypbRXAsj1HdZqiCKZFKGQGUEckm7E1fmBXAW1mcZSzI/3f+RFTLycBPR9n8g1pv15BpZi
MRqcjzfExsW7TfFc6f1B4rqC58a+APA7sXth5NCKowAsArKsR1+7P2l+lutHIaPpqpCHun3Reauo
Q99jW6gKQK5ZSptPyW8uPlLtHaQexb/v66muDCQpdXcvv72WmU52+hCYDSvNQlv1FCHuBTG+ft7A
ujg75fK2Te017K9LfL28zxieNCDNmrJ1gu2l/TiQSnluxjo3p1FNiJcv3is521UdeRcrBBnAM/mB
XhfuOvpJNiZwelxlGTFh/zHIu3niiWER7wKq37t2P6tl9FCo8f2LLTsbAmNxrDr0wJW5OLs/UX3O
aY6jxwMNaW7hAkpTCnvEIcs8VE8YzL1ocNsmKkBJV7KBNWmdrkC3JAI7boYWqZPYgKLdq7MZhda4
JdMlRgD/0BdPlEpmBhTWEx+JwNlJarASsfSTZwcSPmd3LmDX7g+2je1zf4UyFRbTmzbYHQmNbkhr
pg+2T6itxI2BSRLNyKVkPyNl03z1qFdpWfDg8KR6InqFKNpUQvFQMKz8mXXgvKoVY4Jo2uTeQQxo
t4AOTrZIjJL8Y6RqfbSoPqCskv+xE7Dw2UlPpc94stBDaHhFWdBdIowGANqpkDASFWHUr63hTgwN
YLQF6RkQd3l1XoTIejddnMm9k6KaNdUBDF2nOSq/CGAD9aoLfplkNmt5ELdg/2N7NcUjq8okhD9B
PHEBUETX1GIj1UanxnSsYFjW7/MN6FHEpi2IKSS70/A6iZjnlfBNS2asnWuRP21GeHfE1NcXSVP2
Smj0SE2c2uN6rYhn+ZPCWuqRqO6nOw1wqhNMSbaOBsRZrKCGUGhMrtFJKdu/VjNk+YJAicFmEhT8
1dektFrLhjkRZ2dLlgngWQUw2VUJb/lwe+LNoiqLwEjrwedkW220g3g5mvSZurzSJaMn9wqvQ97S
P+ZRh0jKVSsCbHZew7Mppet/OIfVJl1y3YvSD/HyJ+e8m7CryRQPsObZ3LQnp5+GiU3GnhKE/msy
C6kwu6Re7UjKWolymNRyyuQtA0+pi2YA9q3pFo7CfvEgZj3cZTnsrdVwtBJrvbw/FSMj0B5voc9m
u5QzOLTaSjwztjjt3gRirNNhdQLE7jjbCxU3w1uKC4NG9MJS2oLFDaK4zHd7swKraEEWeS2Qb0hE
eqpn0FNZxC3C5EsXOri1lIcr5hw0tmj1DsrHjYVvbuvmdTriQ5tAEAqm0gnuLYKK06EaYnzZfW3p
VGastqlBsb0OVMvGnJGdxGMO9x3xF+MrxjFXfYVSV9EC0O3U8MIZubE0Ssp4jYw7MShddZbejJ38
NThklFi++YjTaY9fzztw2CQlhYg253nAPKnHQ+XO89MEO5viYV92kFfOcT9xqryJIPXftCa5ChjH
z0J5qUDJ/C4PJaXOOO8qLVwAPwazHIvtdwFxMktAg6hdS1/M4c+XwzHVfv+LMERPUsuJSgjvdXFe
WOBLOq6WM2vZ7abX344+KN2msQOsQ/H4oInDxbrKKoP/5NE7h2sAf5VM06QIZi4j8/jePcEVA8zG
sZco8GquYWN0rArpGJzdJe0E6U9THl0YwW8Rpo0O3afBJTSRAJbTloPSYWylKbYBe5EdrDSm76mT
2dTgryK8kAx+pLuhbUfKUhqi5Qy0CNhk0Njd/8doAeF5JjOE+2+wBeYO+vmY0VGG+S/hifqP6f9x
qSOW04m5WmvnnFXDUjy5sanGki+tmvm6feGm1wHadI8JROgOugm2eEMLMAXcKGM61ZXt
`protect end_protected
