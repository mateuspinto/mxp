��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{o�����u_���Y�:�_�� }
�5ݿ�u ����<�ha���m%����Oԍ;�{�ȭ�2{�Z&��U�1�X�z^�ŗ�!��E�e���T:����_tE�"�i����#�4��X����|�
C�ǀ��:�8\�����RZ��͓Ӥ#p6���e�0��F�!%>+�n q�����3�W]cX���Q^�J�2[�n�2���~�D��a|�3�J}R���׬'Qo&t�j��9>}wa��M�m�4��ǡ/�I�����%���*�VQ���z�LRM��f-X��oc�9����[���.���|e���ڻ��7S���|�0�#����!�-�_J��|Y1�?e�`@����/�nk�^����h�P���_ ��^|l�|��:�����/�*=I���p�)�?'���1t�&�	9��	WE4��6���)���aq�:�����Aߺ��W�Ħ�N���Os�#G�G���U�l�ݘ~�~��
#��)I�

�6���TWa��l(��(N�����y;����k�^[���o�G>�V��U�^�����j}X
t�!
N|0�q��Ew/$R��ES/�߻<t��3�\��OzK�Y�V�&E�7�=a�y@���=Mu�ȶ��jȲ�T��rtD%;7�?Ct[��k�kF�����E��0�,`��U�%���3���&���ua�x�+~�O�ꨆ��)�C���&E&39�����ZR�K���u`�c���k��;K���ySM�u!j-L��"�n����F��	���.�a ��f���#	Cϱ`�a�Q���q��:y�l;=c�U7Q{j�2�O �G��؂���ψ�7�_��7�<.�a��	�S���l
.16�h���7�'���(�ka�7�U��T#��dD_],yf�ð/t�����Y���7��~5�`4�8l�+���n�"�V�N�Gߩ@B �E�e�œ�Sw9C��j�nZp@j�}yQT8��0����e�V�>̋��C�%�f�7�Yfp�˞�	�c�q*����	
�TVS��_��)������<~�3���Ѓ����%�&���N��$�	�w����)�߮P�e��|�?ӆ
�ńǬm>�}�F�ޝ�2$[kƳ�Z2Т�3T��h�ˁ�wR� %��|c/�VI���)ە��$s|o�m�}ݸz)��˄祝�p^v�~n� 25����V����H�o�8�� �K�Ӑ)^8��K���N�8�v�H��է�O��#|��m��etw���]`{,��j��
�FY]ӡ&�����v8��͵.,0B���6��-."�@���a�j��c�I�Qz�P�}bt4�	�t<L�>�N�k],�GtA˱���Z�t��"�SsB�����JW�pڹ�>��z#ȡ�1Ğyc� ��-����z��zS����7�PtYHi8p�b��׌�QS�M3�S�]�qa���j��q �@���Y�Y��3(��T���D� ����,
����!��;D�nfA��f
u�X���!(-�/:[��*1��/.X���Ȉu���D��ꆻפ�%���)��vo���9	���"�b���KMKt�s�@i��4��=\�{�6� lEq�e�Q���EbA|�P�϶��>|�e0�>���������<Ž��������j�A��h�0��-P�Y�f#�L�!HHWtS�_�B����-�M�̱b��0;v�.���*H�^���y)�YIRj�o��� ,�c�9�ቄ��G*Tm����t�j��| 7� |�#���F�W�'	7�j�䒔��Tm��&��B��B�h�J	�c�&}�2<j�Cx)�#b�(HY|�8%�����q�TXI[ڱ�nXwGXN�X%����*��$�4���|����|h+�)��bm; ��� �b�_���s�O�����@�w�*t1t�x�W�Ttt4�eJ1�Au�,�N�>JgRP�I�zID-���_%�4�J���PJ��(�m��s#�bz*8�zvE��NZY����g�4�W�v���(=�ǜ���oP.0=diID�\�˧���)��-JJ8ǘ�B�)��