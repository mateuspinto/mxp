`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
XJmgH1KUv0F+J5PB7Lu5mdLdjFbRXe0k0jv6Clv5fMIoXc/5Z9KfzkTlfmpde1xJAmbr1pqdYac1
jtQgFB5NAWlTiSqdX4xOaIZ9S6aluGaB2Z/sQYbdTPbgxEY6Qnw/nRR80o+fdsReFa/13+lPlAmV
ugsbmtWJIpSSDd5fNu5mU7KBuicmHZvB9dRh3X5aTa81SJk2qttCr+oI2yEbTmQk5Lm36USuSxm+
x60UblCcGAqd4zUM4K8FzUGOZ5XF+n/7FzZfs6eE/pzrZNo4YAQ2oZE6lhj7h4C9mNtSC9sO8C8o
hUM+mNn+GPLgnOdMBrCRr0EqzIy4pLb2y3DEO+OcRNc/aQQWIhgUGR44+h6TT8CeeSa1LekF6y89
SYX3j2KVmW1eQMSjJprr67xfWTwLrrqT5BTBp64s98UoxZdeVpH4w/awO8BowGWcYoQQJ1o2rsuG
psX3Yrs+mnJqgF/Yze937FYZnITpYKnGDoMvmbVHkdChBLgPjGuQE2o5eXZB9TuTwfxQ6qk1Unv2
35BQBna/vENUotPJauFsd2bThDdZGlUrgAYqu5q+W0OXBAAmQrInd9ibCpIZtO9BcXBdAPeDil8F
IwBHEaeH2l9nJp/V5Wf8R6valX/aTHxkKpCg17w3aenKNy6Cq1SdMzw1mkNFEfhTTN4ZndTB7Qds
QfGjypVpCFFQ+2a9gogJwgFi8xqB6muIorSxzj4VgBYt8N91+ErrprbKHjoIEWS3BWwE1Nh1xdSQ
cdBHeWhpm06aOLig1pRSCYGHb7IUbwV9sRjjxhiCKDIFHDcr0IulNFCQjjqidd+m/c7BZsLPMqfO
OKSlN2wSi5Z7bgC53qABEeCDxV8CUjFKG4Q76wkyaeu3fd8EGSXIrX7dC01oVIJLnOMPe6xtzAOb
niyeYfKUokI4Y/TGzsGTuv4KjmCBlyl3F82koGFPpYJeB3zGoqgxzdb5FlcSMzS2IXa/5S4aFA61
5aXoCNkXvBeXwgnzttd9qsb+j8+chlE98Ke7NTLwppN0Fp0w7fgMSuIXrikLCMYfiTztdEYWKbeT
YYTGcXwxTTgs6CH953AeozoUVBW6mKZzrFr4y7ir7nqc7p1CoQznwbTJl0wRne4KUyxukycAU1Uy
QZhr8wswOXfmw59HWbliBfKcOihSeF/Bv8pk6kX4EydwnkVzuSEFas13r3kQpgIxwHpqpHPwdiYq
4QmN7WHBjMfUK4FnDHM5JYUwYD3/2imbIeeR7QpscSPl3JeOPjqv6G+ZeVzyuukPR+Ez29kUYuV4
JFir+Y0XVxd4dZImrqLjTclxHNM0xUbOgU8xVP1BfCoIE+KRUjcZpDswGTvN2hj2Cn7w/k52KqRc
qQAcMHa5Wp8fkFm+HSGowjNiKajpgC7sKYwV+VN4GzQWgasHfB9kfuAarXfUvZ9B62rxLmRuxsA1
Jt0J/tHFjZ8T3Aq5Dfit3WZkvKV4w25G67XCR4G3WSTJejIgWrROaWaPzG6mFERh5NhNeWPlmMrQ
txDM0SkqC9nbtdIGUUbpEQo9dPCp5cpb3pTZCr7Jd23nHa3p5rnBbwDCmW90/yPqVSEeBEaQEl33
QfcFRB+F7ROYujh/HmbxaTLV6+lL+eU7Mm5AW+Yu5XMs85Sz1dFLSXQ9D5kwtIhv5xKgLqP/KG+F
FO5kac+BMcxon8QHqDoZDMYTZH9nK/ERZjYnl52hCY979eqyIqRVSOc/BkrQYU8K42FWNURLyb9i
frQ+sXEz8ChHyLCysa755zFa2Ji0Jr52G1ubMVALpMJASIS8nUcDwrxy10nBCg3VcVVex9xf4jZK
MMjyBd3fezhMB3d2ruJXBXek0gzFaqsaozgHwykT88TivtBaK65rgULFKpV2KX4BhBV1OuzZWhLQ
LRRnVhXEyVIvVkghCIKdV5/F61kyMs1ru52kVfYwth4j1WoFrTDpTVsw13ZGKc41ONENEf92wIx5
MingRv56X75UZEZy8uewwcFQEPNeWi5pQlDvvGV7OazrX7EqQ/l65g8Umv/5XGeA2gOKfJaanvuW
cu4LatIpxvI+kkmd9PlBPGi5hbEdKEswOauWgrWQh7WSI7YFDI3k+iJNKpBlC/P9MfGbJB94IeNE
QmzDe4QI+h8ekH15SfJ8BocSQnVQkW+yAoPUTIY2C99xC5i+/Ir66bHrDQVVpnlVm6qTIvgGy3ng
kBnkVMmyJDOrcX64+/FodvFf7idut7jJAJu9lE3wfIJEDCKqtmk6dXPlixDARfLDnZh7fbk1E4wM
YnKnTBInTs3e0X4o++R1vGWp46oU1sCPOeQMhOdbf8Ax/X4zcNyz682NKJkusa1qduxIXKNLBGPW
8mXITUY80uAmlbCovl6JL38GyuwlqEFGYzb1lSgonlcI147sbrx29biV0AyGQSqI8P1wGeI0OoWW
TvUa+PxoTQhd4FbBfkERbCBdysA040fQNowerqT+39Rsrk18umSFrNs1OlzFq0IVLrwbZYzkld7L
nfTei5Kqq+laRLYll01TpdjLT57hp/zy9kPe090SS9QgYap/8M2JICHDANb8oBYu2QrOa9Y+Nw0r
/Cde355s7jDa16FtHSVyI9Z7NEHk+TpK5rZmhWc9QCanBKpoL84Uwuf9ms5Hp7ImxJKi5IPYtiuE
WNIqlInJtu2d4NHr3SpQpSbBDfEe/QSX9PsDGOs2++Fu2AE8eWF7luRwv+n16FFSczFSVUWaojPJ
GsMfoudvNKnm0XM79dGsfAW7ILfxWkaNxBW6cc+5j5QQB4UFVQH0/BwPxUiaYTJpbnGa1cXKsZEe
t6O9bxx7m/VAuGxUrd5UFy7IqPJVmQH2qYwKPUd6n1V2i5MPoVsA+g8iNPM8dJD8fHXobPHXNUx5
Z3nkaEUZtt7r73ZRJXeENQmhCSheqYW3W4C2+S9aktf+w4EAgSTLHwCLu0aEPa4/ozFvTppk6lxk
eVnIXdLOngSvGET943CApCGUfmqLO6zCxxjwWSaC+57MUndaWGRPTXAR6Z6JO/HaBqMCtclntajj
ATCeSznHBiIebfiuCFVjqo2F/x1jplKl/o66o7qHkfyYiz5nMNQkpBvpmsYUSnEU6PESShcys9rJ
eKtH9VRjz4iyqoOvAL4Db6O7Hc9sMhMncwblQnJHaDPWoEU5bcBKabORaA/ja1s57ZbajN/drZHU
NpDiR1tk83kc7ephZ2JaVs7q9W70oQxsMse1Rt7+MKlFY5tdNqaQFZTrgqTiaV/qZ8q/I2MF+CXV
4EaQsQAAZ8zqZ/ip7tf5X0VQJgc4lCQq4WEML157vy5yWnr4Df0z+AfZhCdpVx39kPUH/PH+MhH7
NPDrFSQbTdPg2D9xUgjxVW5TieRNAFGRJeGUvI407NatEmeJEJHaeNsvTFeyMZ5gnffWb5Q2hLU0
suKw5OxFCsUoGqNnByfzL/opA+cgA5f+RxqWy3wFo+2GECvloJBnD2cWrIwwv/DKoTAvqXjzfDKe
hMagOzSSnKU/voNEnYNc4v/PA5PFf6vXkyuTrcZsfuQCB9mZVvylfu8R6VEJSUVxN1c9SUqnxapF
QM3FjgyGBAFWLGA594TXw/tvNAJEF5GRbOxVGXPfwSagHtr8taABiRd6N1GOy5z9GrrWG7xd8jO2
a3HqKf5Qk61kpbN1q8ZLWHu2RLZNkuylYGuxofHuzorAe+sHDtXHnVVB/9Vbg9zxBmtI1olHPlVK
R0uUJgcIKdvHSr91U1COXUxHc67RsIAZO5VH/um2qygb/AYw/n8jBnPgNBT5vvEKkYZOdERtRIuA
u76hciZLQGzqV0EvcBWa9jJiwlqlucc9K+zBwqPNd/dbbxUPrBzvH2ktX2dkvBV3u6Hd2JxjvBWb
+aP62mrODy9f9GW0JU1rI8drfR3z80QEs7BPr3URvOekfu/cUlcZO9klPS1AXQzW56/Fg1e3JmAr
/WW43V8SdW8CL0iYToU2nGjr1zd6OHLMEVN3Elzr7oaQ6fjWYTs7Gyt6ZFTyUVz35XKDAymQhT4W
fdjXBmk2Ov1YVysNGxnrRSJaizn/YcBNkA4O8O7XwBoxBaj2+SaRYTPRS1IQQfEUry0b+IWKpR9f
MSTha6TlDV9UbAbwjAnRv9F4hTpJeTpv3rOlhi+GDZaby4OHvXiV9oNlDnAutpenssPNduTLbkOs
DqUk009H2q8rPzAW6NaU414Z7lCpicgZk6Dp4/JBOozQiq3ery1ZIf3K81POoOT+EV0ouhbPh3zP
if2+pfLbAmw5MbAOgCG27cEWIwS26Uwr7pMUjbFAMyHDWY84AHkFOmj5W4jLiZQmLH0YhvV8LzGd
fJZNcYVDevOQaFMPpqVRFwKc5eRsixMNZoJiAUv/sdXPhGnFUa6Eb7xImWAvDyYgdHx+g9ozvM+W
TC6dWfEKrembmGe2l/4z2gPRgNV0HtFhdUMyfQRgpkC/m1cwFCAO1f92GDmdXqVn9B0I6dmGJ8jZ
peoy9BiNBmu4WbUrmt4WRW5/bF+YYxoms6Q3RqMJYmIAKSTXHTlZFcu4Eo6uJofwblQvO1yb/Ruz
OV+nJdo+pjCPF8nsHWvOKOKgW2khH0P90lTfAaAzslMfK1uIbXPwVvcGX3JMCerZ5AfwzQcs7jC9
rt9De8pzjA+Jg0b3DvZ41Db2gOr7HN9JfluWs3dgwjWd3yZp4WMQ1GnhoCAh4PDl90JS3fLkXuDD
CTXnjj5h/j/v5fx7xk9Y4UMq5nZjTB1z5bVbjCPD6g/ZCOzpnbVAnlLvlHH0RzbpYk28C06HY5N0
zLx8yyePxEjQUBi8kyVUiczun9JYD1x+8g36pD5a96s4xoXsbFVtVhGAT5bs2a19x9PmxfJyXzJW
6AiKmG5yjwlhB0M3E16XnHqFrUJYLRAruJacG/8gu1wPW5/rxbA7RLRASFmD8Nh34Bg+CBcmxlXH
ADngXq6S3UMHv8rT4hCNpad12ChQv1DokYO5ZtV3na1tpieU5AfVq9HBh9NRMKzR8M3QeIq0rg1B
xXBBo9khe0ex3IAZZCTixScKQCpEcoRPSxag8NIuzVtOfWKNM43Qzzz3bIDFHYIcQJ2HXwXmpWP3
nHhxnl415Hw4V0dK4smOFLW6Sb4FNND/zyns4tkgI3OjxVSb+bL7aVbvnuBXrGl+OtxcWeAIfQ94
Ebafiaw7d5whXpmU2er1+QDXCPipM+V3368PMQENU48y0rFbeEqA121s016Jkiy5fGGPLR+ojoSi
MQZPOSxmJWdAL5/sgcaYoRcRz78hw/IMdfNErIkb7tSumrQ/gG03LFmr7B4PzV49Fzc71/FS2vCR
yD3TJsTUSkLrk+Num2h+c+Ai00fAbcUvV6kdOeyPFyDw9BRiy1LAGnDOT/JMejAcLCMQLrwUWlfD
j4pJyUGe00PY2ul4sWQuOybBm7jo+O96sesx3jbwPv66HGA+6FYT4lq5Y75X45V5m6YGIVn9riPQ
l1NzaWSpFpt2hAkIsb6v8CFyqx0gvT1tmpOJ8ThDhuc1f+hlsTJFuQCAWmKqtyoAUOu6vbWwzI0u
KFBJ1n57vLv5K5iouPZ2gntjHVmBPP1pER9IunbxDdW8PlsUrZCts90VTcDR9KlEHo2rYAmxcWWD
Uieda8UZzyuoSc8bm9ke5/+LrGph5QnDhe4AKIkkQYx5ydiEDGnTv35OLvJsOW0OMEWNdQKbm6Nk
hw8eoDbWXxNtG1sDT6zPT9b0yT7Ca9G1MRllyo9eDZmL5BEQMJq1rI91v6kQfbTmwPqCV/nzg9y9
70vvlmm0ZILmtgWHIyLZrUnc2xUbPetU2ailkj5DOki13bFCfMBm1ePQROjaNRkmE+Jqhpgxu59Y
YoiZdv5uehZ6JDpdz2i2ZJVUSrFDjo+HV82CZXhNAT0pEKYEXlLnSAMkdHz622YhaeI8iBd6Scj+
wH7ZG/vlV6+R84/J7oGf9L2YCKeVySMRsGLxZkbiCkn+XqbEyPVT96DC6r2SU1sMiKe4SGKYnwwx
JKZdLg31Xz+M09PZtTz7FPeWJr3alreNPrPr9pGOB0UIXepYzOeJmT5lolIIi9SApc2FbNNz+Rvv
iuTGCU1HoBFe0VjSI8gDd4l0aX8ngouUlE/0Zk5Zgd7mrnN1dAmkOdJDoAnynCalLgqoxKQNk4IM
Cfqh79BUWrHw74e8LY8p6FGsgKooQAg7fOHtnOXwb+90wvU7zJPsN/0qvttEWt5OkpakYEXMhUMK
xIvy0nawWD08D5taBnCSzdOeheAX+myuaFOgjI3Ax6OVQu9WVHo1YTSjgLFKyl2agVQ5PzWypZRf
lp1rfKon2Q++YlzNsuGuXfKOoRKYu4KVf6ZquwU+QphDbwrLobJYkrh2FDkmuX79TzerNqa1+dOq
QJh+bIXrOZvbi4A3Nzn0hn28M0tXo7VuQTNRovOitfRrvhaJfIw/QFWX6BlPsVST60HaUURTcC29
zQSVJwYtOtxu3g7TOyp9IdmkLrX3T6CU5IF0wEasqJeliSXLB860hSFaJUtY8YiBOODIb+W8wWr2
b2RJcmr4keulCM9VnfdAaBlNapiaQgx64/UYK1EsizDOB+w5JarQ/cX3TEPomlZpho2f8RrIym/i
xHRevgaXGgK7dL3+MESQUoxtWFoQ0DZITsJ6utJxWkUVOcdoZUXb9HYevA+5Lcr8Ql0oMOr/jngE
INvoEKQEwCAhQe1cVek2LltlqBmex9pEsebhqyvbYPCqwqHKvZwHG8UtVNcne0n5a/6wjgjR3IxC
hAQ+36KBxRXCtrmMxjV4of09jlsDte8B9uyWHiDz4IvCqnIo2RVgu8c9Nj3wcGcKDDaWU0/YYNAl
gZPIC8H7TSBhX1J5vWhigH1FF1D91KL+UpYI613ZF+1MhSnjlchCbpZ43W2O0yqR/358yCoydlit
m84S5Car8C2Zrf8smT3fLeuNSkl8gYComUqn504ffDQoLccBJWXK+/O/I8Y8my3kPpygVXoyD4CH
imppfJ1LHq0528HAHeoFOaKd6vqIJUWxelumIKl97g3qs92QT0a5fqgFGPOyCqdryDb2EPOcmBcf
uR+gg3R3PyrCW1QwICYGPr73a6iRMQeqN+/oi4S4GvHU93Uu1+JkGCKdZBX12NmaJtqF6bRABaUY
vZBgcLzY6sYfjhb9ya411HSDgAtz/psbH8ijxqdj+5r4Tl6QIPYeuDwwhHpqQAKRj+8MAL9+2bKn
Ura6YvfYopbu8AML4HKOgjO3X9qk5hYsL57UBQZ3zUirYIWdStYlRcGJqPnePONgLkxrl4XnRCbl
vGTkTWRyQY3AgxjY7QM9RZA1GPlDE4HCWqSNleyJPK/mt9bioV4amO3xoiiDaHaF8cS5+DVtrBC9
iNXLjy+Z3KgtMWZtZN6kzzj6m+93F+6d7PdlXxLRz/UVp+7BvrHsKVoIt/Z0aMh72v+JIWJ7iISX
+CsvQvOky0vATcOleaaJ8lOrGLNUtZeo8rKf5YdNGdJhRrxWCgLdcmAAI+zjXkxOHuctdSKLYcgq
GLPZmZhMGhyn/1KpDy7pMqpgw8XCa8N/pn9TI9fKl3N0aSM4u6ibh2x0272868h64Vku48AAKD68
oXRjpNolJ3cWjOozfMVjO5z7AClC7ba1k7ljDJnQUNCTEXmm8dtnpqXEruYoWOFA0EK/PIhBGsa1
rIWkc83vOTt1WCqy0aOafPnjERfoZWC7y4+wBHLrkBCR4ogK7Nzb+1xuLYLenwuJbBkaqgl0cfrC
UeshRFZShBwIekae+Cy9eFs0t5UTU+G+c/Ggm1YkoL03Mx99/ahIYnyAP83z8zYkKCWajACOMhRL
JDPeWV7AMqEUG3iK7wJoFiwi3EdHdVwDBzK0oDJT0/Xsiypv6KRn5nR2+w79rOX48FhCp2o5p4Zh
etJWjRnLzVPVdt8xFAiPpaLfzpAYpK+NOk4dIZAnOnFfUSdonHgQZmXSPPRzTpthBWq/6sqpcu2S
nY9eTNfVaNUDOolDxzZHpCO+env7+2JydnfQG2hK5Pf/yJ0FAwIed06Qyk6MCR+8+L+Lr/VioEiS
UgBV2DUBoVi3EoKaFMS+Az+T+t7ok58qQVS28+yXoyVX1GivhAzqQXYTfqCeNZwbEFGZvqLr6koN
AyDJOB13goA0cHpA7km0uti4qfsX4zrzACSPyw1r2rprJhxhy53QUPbUZ2qBUcKdvwQNKvEiV61u
YXadrEWtTxbsqFZKMQBVP6Do7u/ALXSJCTqETYJbHsWssA05Caq93ipNm0GDJeBRtbBv7dLq4/l8
x3VFM8Z0HBoQYWnSvazXI+xZKlyYYdQiDJKxbf3TZO7hGRG8d4vC7bf0K7FD1/TunF+Nxt8VMLVP
SsNiNPjpJkxcPzusj5fUs0xIysJUMBF0oWnbsx73IFqv/+wb25XGpBWxltWnc38z+Jm5qvT4nYxt
A6g3plV23TFAvafeHmvfqt3mKktBDN5CtHu/90bp+8XbPRgMQ6AgQB61mIzqdl2I++F/FIRum/40
lQAPPq+1eEzmgFN7OTnBGSye5m8ViMlL8FWU8L2uaPLt5/7rHMdlrEFm3XBe4PEo1+wdjqy92Xts
3u+hmdkROROi8HUNk7oqa95/R6dVdYwKeS50NXIm3Xxvo5KKJJPoTNCl/Jxc7SLw2XvKpVYpKeEG
rxtIqU2sBSAAoEqUQJmycWR0FaaWzHLhTTSrFky+zNeUSt+3FppMP28o352waUBKwgKeQwYqYhnl
pCBzrm8ItDlgQgB7InlX8JzihE1YLWxVEMEmGUF4yHe00irbbx2GxavvpMk4MAyjN5+Zg+P+66GO
otG6BdVFZNTM++nWom/DD/S7KSBd9PjLpTgdfqQSPxUEZsmTBtm/yXpiINqA0UD2m8i/0XJAGmWC
K2sDhzlZJAMXUUIsvKPhVFYJp9RNsNS2o/iM5fsQocis8bXFYDmVvjoYfw7S2G8FCW0YBtQLOqGM
z50t1/zSYbK3rBtpgvXUYDPwC8LsT1EYthkW1hQWVxMgeobr4auwWxoQAsHJWvjyhetMt7vytYt7
XmqpSL2tTze3C5QFpeKwMDBb3Hxsue4os0SJsM34syIMGm6l2b3hsT7tLzCxOqaXHaZUITue+0Bq
GQY4y1hvRRufgfzuOkBfHxaOTWIn7fQqhWRvPh0Zk8e3nBxYwjqkS8ARQr3C0mplddYyOUS2Q61Y
81+hbIcV1kSdmVgsrC0a8cREl6h/BFrhuoWpQhOIf6F0GNVL8x1rbJx5W0VPCG9Mxx88d57GTBUF
jJV4bSoGE7ZrZYrLwwp5VHaaj21v2lFDAetz9GeuAD05SEazbLOkOVCwaz1Da7JAffmGoS+0oBaq
cP3/5+6c14Hm8mAWRhNrffPQv3l8jeQO4k7TLAlZyHhCJhLE/VEcuWnXO1/l3L7mM7H+dcDa2QYc
kiaMCjBbXrLv1eDt0UsU0FlhnDXHMLFnzdOW7zD//CteK/HYqQTWJ1bdb4wj/vM/1gG/qHv+Ntk1
ZdNd14f0Jeik3HOKQ9wCIBIGZgk2qgFT8l862otimQZmdjh74z+6pZzTdoJEBNfXOCcIURvDU3wL
VJD7DE7R8CoxdZ63shK2v8w8HxvCDtIfRHmCswN1JJv6VaMXuacEu7Hz7srw+lKXR0mt2XOlRttF
lWjh8FiHoejgh6DEu9kKUuZq/O7vjNwBZkJAmJgzSMqmVTLRJSxiokF/Iij0xyvRKTl5Mpn5Srek
kNk9YMCOa2LOg+3zkXMEyouJIW7uv1dlG0UOcxZkMLz9E2MsCcuWCvWb/R4SSPCJf0+G6KB0QsiQ
z4PhAamvYds1V13urUeQWA16GSFKTiWcNP8uztGgejc7bkSFJFlZK+akKaky6xSxHMzPy+fBsqPe
jbfShPGbO7O+rycApH6mFGpmXfQN7IhaxbnKm+rcJn/O26nWC6EnCPL6Dj9qJwe+F4tyVUWq/APZ
mn4yFblCGpJTbV3RX8xWLuBX3HwOKQAsXOh/VvhvB3URDqIfAqcHTem7XAFtadzjjWMcv8lwqqA3
RGJvHvp/AcXC+SGUBNP3MUMQ8/DJVPNzipBFIKBBQu45lQDhNXhJL3ZoCY5uKLqJZzI/6n9ivGOY
MHMlzIud40EtuNcKCbdBCSjelXzYysnNp+Xg48v9EDSL9/OUmkz04wMaLpfYQUvhUAFTp8Hsaou9
Emkf5pZlO2KcB58jQuhMLKRcOKMXrCJdC9X4jmU+ZwHIMb0FJBMWu1JapQgAkpmw9bLCdjPV4X8w
N1GJXi3K2FnWF9fK/7QGWVZe7RGUMSHcVRgqtEEweIQa7EUCldBbKtW6d5CuOvZezLq5k7qrcbv3
IRQsxP/pavayf1oTpvjW2s0b3LekGoWxesypkaIx2A0K1dA4JrSp231/4S/CTR8Tl4DzD4dYRvfu
yloVq4kEDcJ/bx6G3EUt+gg9aJ/9qJve1ykBch/o95rJ8B5Bk0vBBx8E6EP1XqIjdyS0eHsAOMHW
tWdb3de4ME2EWVIhw/M38P6J0SxNx9ANrzMIYGy6ZUMAg0L1gJVv2+9+I0E7JObtKZqFa3IF3G2W
5hes1k8tQggjZ/ZnItC2wZ9IA3SUwgWy1Mm0h/9nluT9AUoKY2ak4q8ww17eXJna6lZT2CDLdZAD
SyGxXaypOdlDmio3A12EM2AnK67wnx/9kS5WvtW9dKVbesG4v3ePNhNt9SdyrccIJGWMknjwJZ6y
d1aYs02lnnrgbmX+JS7wX7HtZWpWJzsuiaaMr2F9jGej/LXzmayba369f4hVJtwv2+875rvresKH
2CVlxXIgvegtc9R52R9gOtFrkIv7x/s9hvAdZgzEtQmcVckGiImlBm3G24LObb2b/+IgeWYzP2Ha
N9qfEsOiLhkKGgUSVL8+OscAxWux2DBpImGSVnFLslnzg0Du98VsIVoNuNR2Ih8f/NiOWYs8Xnpt
FLYhQQBe8lG/FoMcfFrFTQGR8b9DkZR7AS8FMA99RbHOm/zx3hbfkHnESToHq4F+/kHi8gtcMGhn
b/dSZcatV6dAyHQGlhdH42XDbblWvJuzyi8Tz2/Grw9/O5LHvL8RCL7GtqaKmxa9UPazacjx+3cR
FRwn7x8H7+JWpEpPPc7vFhuS1XHYTA2keYqyH7g3d6nYm8t/cwbKuUk8xVX1u/cLSQdSHtMg8EG3
ihy6XcUWBd97mVLvR5TdyYUpZ7J53yCKr1VNv1Mf+F4tHowQoouR98CpSF9V35jSnTTjdeWHQ5MQ
c4wTXuVXKYOapnmET0cOuZMlzYBNDMh6IfO8D2jLqd7RqRX8FUJgZtENfxlsSyPfp+u7Ceg8yJJg
CNdetCtCQunvsWrbhPzEfUqeskif3aeE4cpPyzT/ymmetj8Wf2BnhQ08XC+DNGE6R5VQptlMEFFY
+U0KFTTyN6VCbYGWyZiXJ1uylAWxYgqCUDEdKG4Abmap3WWLedVMxselRfHkya1Jvlt3lKm/8OXx
pJ9InGA19wDw3duQi2YklARBhIwrPdYTYF5tZxsFYN/S8UgnVzvxnsrwUNiFQVEDtMSzq5N1gXaz
LLMjvIgvSP5cZMkUTkAvwIfWQKnTRxY/1r9bFXKGrRoC0UdU+VUqDQ0oPMZeItmcE8wBMxRPfThD
4YJh9Tcf2IxOIEsKQ+6vZvWG95cl44lb74NzOvdj3LT9fkV2czndUoOaXS81oMltHxu+GRqcN0Cy
YIiM2Rve18WaQCLNzUtdhQnPjIy+UG58QA4ihPm/thLzzzURsaZrafDK0RwVcvyQzDhL7yIkiSmg
IO2aoACFjwAsSggVD12jjbCPUbIAfA9SGf34LVnbISbY4Nvbnj6ww0RRvCpRovWKsMhKTpQkYdqR
TUAESROFiOzFn7LqfutLm45UwIu7Jz/wg/4WXNeramKFWITd3V+75WGgEYr8h5V7x9OohvIDYN6Z
3gGaa/I+YYfECXGoaB9eQurJe2v8ZQ+0/nwDJOVBNEcG3vJGvwgFu6XhoGM+6EbH4F92wuljiJwG
IbO+gApnOK+sseZP6YQoYv+96okqtl2OA9GioXT/KZzpkw3EWTEPU9sKoeSWbdfXoXx6rActc6Qi
eAegY2fLZukolgxh07VSdiSybBos0rs2ZnVUA7OkIQljXiEh88TCN/4zbqQO6THWabp0G+KSNcGb
2NRYMsuYqn9APrcgc0Abauma1Gw/BLQ8DWldAqHSKADeKZOaJHUzC/6zC6rx3u8BslLacQLUmcXw
jlwT+cyX1v98k2zpPv6aZGshlMVwxc/N6m3/pBgnSibxx2ABoLE0Aig37bUDZ0jNMMAyo88W7rrv
UBOHk+LgUpBenxYKuDTZnIVfG1npBNwOjfl8X3d04/sV4UlsiXcBV+X8jioLiMHHvZYWDWu5BPcz
X755ob0cGD4LcGIEso8mVVlrL7R5vM0rnOXolwHwYDhXTxXUTU/olUK7wZ5+4K2duzSLq8XZuvbC
CbAC/uJ0Hg8mUOn18AXg5SH5aXWbtmltjPkgkm340l6Zw82CKqG79zkzDJvgIfoF7Y99+IRhPBwB
w9lDtBLZelQjVrvnRlqLhQquwLlYWHFX/P5I8pJ6qkGWxzl5PdBctXLgyY8zA2GAib7cCaEKFR9A
0P8akddN2IIdh8N65HwdGo/aNzlrUF9y6pA+tq4Dis7TDuYZ0rK3RDH5e7igmmF/jindwfbz+CZl
uakyc712h9SFkqWzNgb+gXe6KopQNBFP4z0r4Fzn/VeeKuTw9dpF36eau07SB/sU8krqvEv7ti/i
GCE+sq5KhHC14METdHvSikYQ1j9EVsfbOIM2ZhW4iZTdnl/x7dQKV6P0r0eCQSsWBzO810Gfkt1Q
xw9L0G3q4+6R0DxT3dZuKIM54Mg7ZazerBP9HWCWWbwbMxPWhmU88AewlvADMCrnhSBIN58WtcTs
NbEflZr321TvS9o6xr+4w982x0xz7FU0CcqWe3Iv3R+ur+nnfiB1q7LagWa8nPP63BUjuRfhPISB
C1xF8J3CZNkhU4Tb++ly4Gb2Yel+wCiFNWj1V4+HrgyZnAYTQL/KIWWIfmZcQQReiQDv9Yx701wp
UTenkaLhraQdNBcbRYMKZL4RHe3KxCNui8dXoUsUvw8ThZYBp7XaHdGIqmPGidlCFLAsVDatNotE
01OXgxuavPtIs0+zaslD1d5ztJDfHKNTUyuKQZlnMy/Me195GtjIx0pPzH1T3PO7Jga6rs7nJQ+8
67f3MLdD/722h/8jXhdNXxZG/tRnugV0F38pGneh9R5Bnci20yywRDROUi6idj21x6mR4+0Uv9pc
o5C9/If7/nhAZHggDhwe7XaBQNa9i8hvX4YriEgUjCIdiQMP48dsI7GpV2Vj4QHd29c753Q2oB2v
JPqqWflcfRP0r2w9i7m05Ut/ycS6jWo0xbSPSHfJLXveUOnt0UXvry4Miw461lJQ9mXgHbpJv/LT
OcfOAB0HDyrt+VYpdzAqftP6Mc739rZpTxHmnIUDC10Kg3tV+E/Fo4CiFH4V4mHpsgARCUp3IopP
Xt3EwX6oc9LCuxyOh0FOvr43Z4AOfdBOX9XierEyEE0mgEN3Nj06dPAMpCHbqA3XAp0FyAH/Vwzd
HElwRMT34sAUDX84tF2dc67s20hmsML5JUhrfC46hshHrQHqEB8aBTRo7GBo1zSZy+GbZM8iODR5
OGyYc5KCjBMn+3Yp0/swxTXOnidf9dMWRMfXXOxOwHzQSPKoqWF/Z4krHb5M3Kj9q8ioF64lmNyW
4YXoRiCGNTriexl3z7ZMABqx0HHA9qEKIbRgkwZt1xVKstlAKFQ03SUDzsXY5GAZ16mNi+6/g/OW
K+CPkcnGdPChC7roivfPaMZd8Pewnx5RbVTYuu3+GeydPHw28q0dDijVbAcbjJdCVj8Q/a+GNtAf
mrVTEsmXKoIiS38aptFUYb+OctJ1RHDSgglBs1TYmoKG8QMN2eAmOsyqJOp97QXa44BxcYejCPcn
p71ELHFD1Ev1y58VNrGMf8SAprVyP2NdE5mlyKkjgXba6RwdVoL+zzld+gYxqFGT+8uZzFXXx0GL
Vr5JB4GOubf0sjpkw4+z+cjrODJxlNIbYSp7y06cYr9b6HAWjlwwVDI5LXi4GJ7+QrPrdY7zGrc5
6g3jWfCc8w+TWhupgu25NEPoXqpDPjw5G6PqUHPhjItiWjl/Lse5pPjT4duGcfZhOr/HaZM3g14i
EPLyywrOPkz0UNDbJAKiMmiwyTnJS7UfC0VP7+PdU3pPzxxoakbylcGYmGX5G9V9AB+RoOWG1aTw
jUnFhUckSFtcxIAz728O3sNIuT2Iggo1aznwEvgKdeLbTuf6Oeiw1qsSyBPNEBWMiewMI4p1Z5Yr
IbyOZ2jW+BiTpbLiuhin3HdQv2qwhIjbwNmbxlE/tGdpDUzEv6X9bLWYTX3Ksfm7c0M9x2eizcq2
qYPCGGairQeRqzjH0TPSBje8RLYExrmnEiaaKALmncUSooKzVemnBZ3aZ1Ri3Cafho44EroNAejV
HOp3zgUZsvcmJF0N+UZ4hju7BT7oxZyiVV0ehVqHqmIp9G5fo0zg6GPqlWmQ0J1bearEDl8wsMt2
2P+KJ7CChqdDPBDGcaveY4U/CdS9G/5/sZlJtra2UcIJdLqG2tfwpz6uDKEu6DAN0SWk+bW6oHxq
jY1Gqn2paH05uufCB04NEbW4cQb6TM3zuD+tRezMytlhIvj/h9W47bxbK0rb9GMbXaQtdxV1LDJw
0Z6dITIuGRkztbwn5PW9HRUh26+B5x5Xk/ASaYSvIi5ebvw/PJzsN2Qbx3/z/bN8dfLyfAPqOTRb
HKF0PRAfx131iT62PR9coe7tBoZ57oHXtKU/EfA9yyPj4WhpWdcKWuicZlc/yXG747s2PYkwoL/P
hYz9uPRz8xIutk3BuS9t3xEJOFMUNW8VovTAn79BfuoJ2OaEFBLPivP7nqTxnuFiwlTCR6K1nu9B
tmGUY2YZFtLsie1rrUgXuwD+w1IBESPjYT06bUjTWKzKyFRHlShNUiW/M+H9VNcwhu++jH0vKaor
AD6hrBDbUruYvn3it5c0TM6BoTlURpaixM8QP9iJvUDUGUU/OuyLXeTdYfOUrudl8CJWSq9mnciA
eEnYjiCVjKSZPMwtD+Y6XFoQMuF0IMbVx4Y8HCg1iT1ohyQPKLKmrul3GKIUCAQSwwOFMReSsOwy
wSo4PPIf7P2JCN5/H5mEyEW6UfLrHZnkXrBH4rG9CAmXQX5fjR7jW2u4m19HkcldmGz7XgrzPSqo
rGT67/OiTe88ygP6COLqqkYuAqsvQ8LHchqOu5izfxMDDeq68dxShNhsfuH6rxyu2WsLx+f5IVav
AMv6GPZ+w12dp9lS68UbDGoSvSznBD/j9QuxFKZkOmnadwiFjTsOtC2av9NCyRbEpqFrKCrVx9Ek
kuOXyci/kzw6zyIrD00TFcb0Oyua9CBF66iWACe/BPX/D1nNwuUzSbpTqyxKopI0C3Z2YuiBgkbV
Sqa48Uvt7w45y6FUA4coTNhnA/xPYxuTUv9CPWOtEJhUaI1Vtkmulw5cQkah4gqhnjdOkw9ECKZb
nWxzeu0NFnm2ejllj41GULBlIF/vD9Qfpa0BpaA167xaqfaZkeQMXCXPPH/VGRKsvH2Lg3N868s/
2GvnV9m1WCs1SWOp105UdqTTBPrq8AKMGvKeqeSN7Zq59HDy2A1okoMyvdTNCSLx1exiV8uAvhpB
rKqdUrBeSsetsW0UGj1h7vJLkNjEjFN31Wc9M75b1X/Ozp2VkWmmdOagEvvAweMo4yiDyQCgAyn/
CqRTZFRQqi2EjlUnnCVgTdGKTZp69XuLrGMossp4PB6TUnn2Y6QUxFP4klr75IbUjm+wTRgyXwdw
Cwut6BL3cL1cSyaf9N2cfcoZleEGKu4BBHf5dz7arWMmje1Wd7J1nfYPxjH4L0mhFqljkIfHcC8R
BdeKOqcuSgJBPXJeo6y4hGZLBAYkD9ulXD85xPzV432kC2/s5ZogkNEPxSomVA==
`protect end_protected
