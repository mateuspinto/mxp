`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
0USWSUGxovGsyBJteYpEodDHW+uAsXfzjLXhC1n6r3W0nWnqAuxw259tmAZEmL1q+eZ1EaZpb0Kt
fayPARvF4Amzg3E5JcB1nJrMz7DkVBQtykMT2hiUSR8iJs9XrglkQ2nMzKryHnoTzIba6VBV8EsU
8fgopKnrBqbWZiAejG9cmkeYJGTIOTIXVmsyajj3GnPt/XUsd/2xwUU9vDAqAAQw31ITEP5wQpGC
Axvj/SD07+BiLQl+qGRHKWnebL4QxoVqX5x/UQJaXM12DP8tKKqRWyuV/7jGlVI7fpQ08emSwc3o
MO5U2NODxjF0qdeH7q0h3CHinO1OhffBFxTrBUKq+49j6/QiQAo3QU0TpdB8z28vnmbTu9W1eWEK
ZXgg4pTbzPRGhcxzYUrYKvbWCSwv+SL7kUVdmIHre9UrU/tfTCtoldi1afhCOwgiv2w3fy4allP7
KDpJsa/qTK2MKyDMKQYycBr90Z5NHBTJ7+5f8HVn0OPuhuzbVfPe8mSzv1MfGc91YkrF1h21AfRf
ViKybIFaGccmgHA3b5Yl6T7mkbTupCU+Nv8eMTikSJ2CyCh9+zxuFYkAj9oLJeK7y4xmkQ1hxUvx
KElSNAoEH0l9RWpWlm/xH3P15hYxn8VSo7S+VVnX2NyrQhpk8DXey8ZTaqPNAquAOEoi0FwxsYQ9
NKn0ZvLaE8QfsSb9VHJhsV3/dUDDRQEzLkzE9hVVTy6g24hgEwnP26NgbiTo2kgmTRd5shAdgHO+
PCk9qYKNggihK1TnlAJ/f7UsDaUlXAlL+HrZF6t/Uq7HnyNGd5v8o73YZtlMhNoIlZPl22xWAqAo
m5w2ll6ai0rkW3wb/49R0P2iLFspq4HKQ2PIVm/cmyvJM5qdQtQ3IdMKVU8Ojt+QAeGmdQP4X+F8
sQ6tcNakSqHPWQ3zYxFx5uLTf+xuJJIO0DKPqaXOud4TymXzupqieOge6KK61CSdDgemc5kDiRaz
fgKwloPn81VrbcNFe/7iNnQUAk5zatLy+4IaQPtmSwN740fPYV+3TOB6xHJjve8U5x4vL1/zv729
CHJzFa+UgNDHAugyxxPAnXrLArOkekj+nnGSh3Rdo8995Rt1eHMlkOvo3WIkDz4U+VBm5c6arbBP
Mu3gaNt4y/e6LHLqhmlZHZtSQNUF2SA2Xtrzqz8I8gbHHTYIVEng6GVAtJ0EoJuNEA359z48G5oo
MLKg/0V8A7DWq9zycfmJAsV+ZBWaRpdYUMp3XNeqrm/VV6v7+bpJl4EX/R6Gj23fGHFTPAavKGgT
uNZm1R2VJsDhxt1mwG2W0J6i84/4RtnFQUOtQ25TUvNz/ZRmfqABIqjDo2JHS/JzxuHh2nhjqOTa
odYJfVvsaBiFFM/txPm0erUUf/gTNLJ3Mf0ooJRousUy4BGfN3++1Hr0ibtCvWov7RxJMy/7ghNL
+kHjbzYzBecsIm9ugSku9ZnwrOLNCAxqllq+L46am5z5NubtPcUh3hrG11NVMRHq7OZdGzjXrlUH
wxf9uz9RJrAPr5F4yxFCI7GJLTvmSOHsj79zDbYqid3YruLrcdy6wJqUxOqlwj8Mus6zv5CoTSvK
tsCC1PhD8UcQPVM4bjhKol8wvqiGdvchOp8lcni9/nW89yNJvzfQlUsmCzGedHsmUYZMOQI0aS8x
2k8iqMvJw8or9redwBJO+cW5dhdacKAUm41QSpJFB2t0hRLgVFPF8g4pZsJ+yCODBJ/RUl8ZQiVn
kZjMDxC29YwRCx5YXIQ5gdamzS+5JqP4DKKXdWKFc+zJKQhZDTc8MvloReY/YDEKOvrYqQ+zFIs3
fLCh4YwgCgqSKTiPimH9hizsZzYCYlp8hy89ZiOufEQ3+61O0M9omO9G+iZyYMbKlR7mPO37sI+u
i9qr/2qNznzCkgtgbKsn3kMa4fZcqPVpQkvo6Zvz6meOjdZxWJwgKTRWPFOOm+vM3QGJOXaBYmf2
p36kMSzd42ooJWblNK0RozjdnNbuIdVtUjA5xq86vKkFjHp2CQN9FqCu6pHuhKuXTzwGOE+fC4J7
NfXqSRfWffumxpHs7aOm/Wa4uo+0aFJpNdwIqI7rN575EZDnq0XmmwIyKbAerPmztsv0L0M+ih7k
76cl3aCGGysTOgntrHPzZpieWPJlk+VRbrD2IcVQvU+ryyjCX3kFV7khWjTmTdfGnDMHUJ3hsDyP
AMKfrjQl3iTc+6i6TOQyLF8hd848I5wQn4GMdF5W4yU2Eu2B9hhCP2fEV1387Z45nQ3y2yJiWvJA
fOKCP5fYlf4HOf02gF8tltZ6lfDQ//o2B6pnWH0g6QatagkTaNyH3XttqEssgFjjgZV5u60nu/OD
/cHRY5CZAYPxrDDibIKYZvG3srrnmZwNaLc0U7sHSoOUxs+3uYYT5voqy/GZkua1keqUxUqM1R8U
AUzLDQ9k+n9tg/0VU8icEo7vKle+7MSKbYd2W/qsqbMWlFqRab23/hBx91ZcLQq9KJU1FMUpX3bZ
dmy64H3RHY0NzaZwPG5toUQK1WtpBYgOFeHgam0ffHpMxvOTC+2qru9Vge3Q+ZkphW48pXNg5e+P
doafTuxknteVa2FP7QkNxHDVlvXnrc0YkradkhV58hHSsLTPdpm4xGhVJAaRwMcnSY7vmNYyhGGL
EKX/s5eTdx0pDBHy4fzZcZ4k0rqhe/7BZ4D/IqVpv//PHug1dcIGYK13ACSUoZP/arrIU3Myqaa9
lAYGdfoy0mrYK1xCsjuRXqTQUnKA/kKpFRV8YubQ/hvkszaEs2ssY4TOg0OmvHwgu7mYRIXoDB7z
h6S8x5afz/zZv1B4+BJ4xGTRz8x/qDkLdAd9Xcl7aDaCgyZwmyXzco5XynwqQ653dXSU
`protect end_protected
