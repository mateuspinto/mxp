XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ۤ8�ez���!PL�7�����[���ƅ�r>!<�C����RR����t���L�$����������EKw��#9A���,�D �y��j�3�}4j��8�y�g��V���.03q݅3��xfBD����Q�k��pv����u،͑��9��j]%�i�Z� ��i�|�y{�0d�(�:i;ֿa�%O��?q���y���U��^�G��c���m��`�e���Zhj�>(��1�]�LD�P��t�B��P���Κm�ʱ�l���r'�J@���J2\��Wk$3� �K���%��U��L�_���xᲞZo�K��nM�p�BbOX�#P�vY��獰o�F�0�e�/7�P��-_�z�Xf�9�w4 DF9�L�?��V@�SHa���捓�#���ʉC��T�Vα��^+�.��W��-�z�M~�<S�zx����p|۲�����t����|���E�����)#��K/z Ґ8Z���l�r�G�|�z|	P�k�#��I;Ҹ��;�~{�1iG;�Ra��
�7������P�}
v܀����ɉ�6����>FB]4C���*��ܼ����k��5`SBv�o�Z����߲WvV�h������u��]��e���d��'�y%�5rX/���/Ñ�w���Z<y=�Z`{v�7@0���A}��v��w�k��U@�l��,<�}��Ȥ��3%5I��7�TH&�V���W;�.�)�uu\
��XlxVHYEB     400     1e0҉���}�Q�d�H|ݓ���6&�_�3G�lmk��b��"��,WT]��DWT���J�A�ux�B2�~��Y-p�!��b�횁f��S�����Y1t���ca��Q��}�I��7��,_�����(�C�?��0NQ;��>�I=	�������
���_��z�7�Ѷ�e��N��eQ��Ib�M���r�o+1]��]$�蟦6q5F�bG��:��/�-��s��9~�o.�	�S~!w�R�.�*� gZ�4I�`Oi��eI^3(U3��~��� �/J>k�;۶�l�9қ)�]�8�gu:�0�������R��;a7^R��<�<hȞ��x�Bq4��:v�)z���[;�)�V����)�j+����X��%mųF�#u�B
,�2�Y�fJD�� �?���1���Em�r(=1�&�J�S4�����l�a�qu�@],��o!��xí}-�K�nqK��XlxVHYEB     400     1a0<��ix��=���=LA�L�hTG�mq�֖y�Y%�����k��t^��6W�8�y���3���g������;g{ڮ�#���6��b� �wp�h��䉯QV��Ѷ���K�[mEt	Ӎ�yw���m����r���k2m��%����÷����T��[7y��,�1�YD�F�1!B��NG$~�m&�q�ZL qZaTb]t��3Ͼ�u�����O�E��\�U������e�!D�oN;.Y܅]`1̵=�u&j�i��Tc��EM=���k��3*�1��Ȏ�:>���]�v��X)�VK Q<�����UՀq�(r�G�$�
��$�Mߵ�����A2҃�ukDM��p$���|��p���/�g%�s]^¿_�
-���I��8Q��2XlxVHYEB     400     130˟21�R�af�8����Y�+�T܂�������s��s�3hhR=�W��	��Ϸ4(�!�>�ė=aQ�Yq`��c_�FV�Tg�Ueu��($�X@���5���4�@��a&ݚ ?!��	0��z����^���,_�E��h���z����T�DKN�(s|��D��O8gT�����Ǚl�~u�DM��1�*�m�B@��^�4BW��oz�X�����cm�VH$+�Ѵ$崽_4���i�߱s�m�a�����=D�Q��S����-ĩJk2Pԩ�u~�>k7`!F��g�i�S��XlxVHYEB     400     150,tP0\���^#۪�Z�����:���R�lC�j��~�*h;�m'��]�dؒ;�v���Mc1�����:�M��{�dYX�	�f��1��~�@��h6�k�L�t$���� TaR�� k�t1����UoE�2.����6�� +.�o��'H�ۜc�Qr�j C�WY�25��8����{��	��+��o7��*�A*��߫.�3UI?��aYS���Q��+��+P��:���t�i.���QBq!|S#Wy ���%7�6�L���'�������tZ��hM��X.�Ŧ��%�p�tP0<���J��m:��Q$W��`�^�XlxVHYEB     400     1a0��H�����,	>���4��*D/!
��LX���0P!A5/����(�0T��.N
���紂�ݍ���#Y��ψ���!9������dH3ф����U����A�` �2�r�*��{�����Z�լw�����2�G��{�mS�����6r��D�	����ppE � �� �:���5
��_������v�WH�06$Hت��e "W'��d�L��G��~�%8� h@'�q5h���a�:���5"Q���ãN�}(N�A�ǖ�`_�J ��U�&����}>G��][��|����;��U�Ev$$���|�Z��k�R'k�a[;V��� f�K�7���$��c\�snn\tb�c�0�Q��6�&7o���Rۈ����t^���/�L`�|�by±�d�Sgl{XlxVHYEB     400     180�^y�$aE�MV��bl^LqI����a��/�F�ZO�;0먗j�h�:����Ϛ���9���3�U��D'��+�նG�e+4��4'A�U��r)Ga�������%R���*��#y/�z��6�{:��y�m�f4���,Ǜy��J)�N���LzZ�f{�'s�z'�w?z����Rbm��0;�P�-EXҙ��h�c��~���<u��vc�`�&/�N��F���ݷ������R�]�iM��!Rі��'�Oal�H�٭��S+$�p{��o�G���`l�X9%vK1�?b��\bY����Q4�m�v�G�_�hp�d��HJQ�`{mF���{�w��v�R�b&QE��S),�~`�m]�\��J�s�ӴmQ��kXlxVHYEB     3a0     170�jw�ΐ�M{��$�^q:�8S��h{�-�*��/�=@�_Pq8�ը����PX���!�1��Ȍ=n7���[���[]�z�4	歺��_I���3�.�@I��:��p$*�Bi#I�KrI�Sy���Z�-K�k�px׏��u6[��5?�K]��l�<�$��Š�A�G�c ��+D��BX~������um@����tޘS��qr�,��7�A�iHC�E��Y�ğ�>�֝�~>�i��6�G�kj�w�{�V��Z!����|qSݪ� �'�X�+�FPdN���"��lmBM��fUS��+ K�#e/���D/3#��N�����q�Ka�������mʅ�����F�j��N�m��r���2�