`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
kNdFPLzprnOffkMuiuw4xRvXLfVZNsmJDR9Su7l8sR7pvOVL9srMyYM20wYBSmobbV3wLoD2QbAi
ikzQMZPR5NWwxWLgsGItLLY6cttlLRqmHK0U3RV3cPrID9Qb6l3QPGHpm/MbAWxmwD2cwU8h8NU3
+pW+I9U0+GEAL/BM3WpeK/Z4OAbsQhHbkG+r9KW1pm4+wIASnZB2OtnmcYTLBNzX1O911SHF5OH0
czmtn3Myn81hT9XO2xg4/0kk6RkFdExctjuN0Oabfe4/XvrddfMpoYNtZrFyuIVF6S8z4I3k0vOT
WNrdzESaBQmeUkwd4AtivHeOqoPdyzSZolWLNccVJsyD0BXK7AHkSn8nGLDQOq55m/CJ+FnOwqB3
eW10PBmeyx9PAP3R5OaM5/B0MFQAwZhnmN8EcR6rxsclxYDsNC2wqtuS+JDkqBAmBknDykj0QJEN
APKQVO75l4yeToVqc7lZmD4SepKnzUQbm24RvvQUGvsIcorIp4eKN3lEyl00BrS8vueMLKK/tYcj
zadMUZGHPFNox+2Q4qxy0vq83a6KdFr8sRpzuzYecMh2ExiY93Og7NgiwLbJl8bzu6lk64QtRl17
rGoBKU7W/Nh5SPh+LbJbv72z1H2bHGbYqMk8HTuOtK1ayugqx5NGcFlec9iuXjM9caN0MdIP+I2R
TVyZZhofLFwW7y4HbpxE3hCvnCcxEUraJ26bIakekJitgM+5+xVNYJgjAj/GIjRW07SfQp/obhZP
OIHJ25UGr8ASkkNOBLuumE8KpRwhjzgFMXyWY8HpJUfK+cgA7Cy93XNnmBAkP0qscfXTWX11rYeK
IzC1ps8FyI0zuLnsShVm0l7fD7SbA8YK6dUhlntg0o8Fb0T0eHkaELHm4QdTRoyt2OzZKCGDoDbG
Zy0RqNg5sp3hXrHJ8MZanef/N8mvzv15j40Fei95JWkFfuXBNzJTIxEmGTCrZjqx8vlAG5TBigA0
MdBszQYQYR4ZLsbJu7Gn4j+6oPf0C1wGFZw41uNDyNLtUUz76/RCVubP+TKSUCkelSq+Q1ftmo53
KEyEH7Zs2F+ySjF7aMeD7wUMWYrSwEK7pqFaTiiauluOb59TE3r0oe0lpCO5EC9E0GvALYJRh6KP
/YYaL2vt56iGwYEQr5erUknzwhQHgO3doj6Bqf+MpERFrpTyPKJLvx6kE6+6PJJlPOWWQxgjfL6i
iWcEhIyMbq03606yufzpZ1/q/F3xmmUbO3kFGSrSc77CyAcfaxtuxQdZF7nUtrZkEY2uB/OoeRJr
m0owH3ZPH6i9xghWPP4pBV3GH164DWSMlrk1ct4GbrQHS2h22Dae6gci5G73oanFSlOlExb6gQG0
ebosrxtvz4+Z/mKSBmO7HMlil6onFrdhYfO+4ak97in+ztlJeUZ/yV6JKiBw5lSrRHQV2whOe/yV
QS6J8Vs0pO5Br5qouKOzPyK077z2CI23w588GYbCpJNjO7zBM7LnBes4yw7nNXma0g0BZlrM1Vqm
yRgfASeIJZgnmCUqP49MRW396rgFDCkE0olxfLAahe+w/FIdSvcz5NqvaycVxyAMGX5MfzaK0mJX
4y9rOdHF0J/ajwP/FJu+/EKQ2rn3UgVGJO2KMjLwPfYfHqUUoHMvZT3ijDLssfzmJA56i4BzTLno
D8AF6tSOQu3zwFYLI38gUNxXtRjnrPSFumIFdYzgXUn8EmuhW9iZbFEwQYgUKUbLCxmiVISjJiXx
Gyvd/5I1xJWTECs6K/An/Gm/0AIyPPB6qTrl4jKrokfVlhDgmKurkG0uvkZHCtER1plbhZRN1qrZ
GJ/5DNToz+96vcvNoHaOnaAE/wFoVpGn73s1chti/v/WevwQJROpzu2f9/eEmKdnbzGdR2VLEs0A
FWLXErDjhgTAiLO8QZZCvmbmtSQQZll4Tft/YWBxVaj6zc1oS8o8yHA12he9/msCKq+FdQDYTpAI
80x2ViPky1iWMFtj24+gduj4QaKCBP/egZJoyQWiX2pX9AJ2+XEeA9GIJG/ptik4x3m/PjGFCbRB
pX8eVWYiFWm5PZ7xLl3BjG2KFZJGsKjt3tUchkyPPE1w6eSMFmbM6Ont20k8LWvmud6eqyCV9PP4
nIqsKoz12uvnY19W5ez9Zm25IqSw1DL0g8dd5V/dUifsAF01CUqR+abAeuDPsbgvqY1v1scFox56
QDTa1D/4/tGUWzn6yo8ZLhbHyWlrR1t8pJRSnYjOhmL4TaKjjTVYl98xdUlmnlZ3Fm630atcbI4d
aSQFlMuccR7qtik3LGcEkM/aW10SOzljNt8Bp1LxA3Z1sq8NNOQs9q5V6nDFjMm8lr0S2JUcZ9Rb
WIDF6JC+GmfWYaTTZhBXglKjYhBDq0vKXuDw+Q9jMTJXzFrl/uoduteJp9fj9EzixFUb++Tr/Ukp
9RLC9XSn4QfMNNujlVsJQKKW+FfmSs5tq2pHv4geb/FFODqF+0/ailPVmaslSTkZjvhYw9bITPo8
nFUFcPjMQK4V82HsvRTmUtXq+Q4WpRtIP/uilW+AkQ0xUgiasEPo236l3MmjaWipUQ7XjnrtpSwD
SMwKFllE4WGkiKVDSdwDD7S1SFqx37rjYDHebStjOmq7La9JzF3au1UYu2tAiR3DTb0SFqJ79nZX
7fplLooXzgkMxSVfn+YhJJcp9DKYWGad3a4KWaS5hTHqyFPUDLmzQFPMRFoQkvxpTQAJSCJKwAA4
WgCctRBnqMFaGzezRsSwDyiG2tT2pQu3A6Ty0O6M4gm3NbgPEBLs2bzop9OKUHplxP6kvkeIkv97
e9pQNj7vbGWZX8B+xxC20Oubq2AxAN4H5HZIzMBL82IKQCNiGvnYEj5iknKtIwrdmIgiWyh6Z71F
AZ9T9cRTIWsXU7V2iwX+vTIzpk5dYJx9+426T6PuoJjz1Hc7J3DjhaFEzXsuXReiEovToHeyrsRZ
rst/p+BQOfS4/m4dzJSmcQOm3pYtEENyLXR0gHGNKGhaGuSgo0hhfxVV9jdF3LqcmrTrKxzD3j5P
vP23lGEvVBLNvGmTFPKxXkmhB1FBYrNFLX0TanizZu6cwAzWpwlv0NES3I7nq5BEmzLKQi7HD3Yd
JYjoWupD4TBVylEU+5wutVsaUSqedDJn5QoEjHMq5Y/JO5Z+tdBbk+jUSv6TaObiJGgXkc7lCV9A
UU/iz/qud7+NJJMX1vJw0N47tZi6Oun/rhc5VmHLF+/RuB2n2Wxaxhl7KILAwhAve9TvrnJA6Hmy
I1F6THuPUGbf3/FZutsshIeAU0hf6lUjyeAuRxXZM6thkCp/288yJTovlY/zSbuRXTJqD3uYwedq
rzqZFvPX3zfo44kbeD1SmHBFD/nd5+kkC2/7z9byTfJWDKnRvDAlTimZEJcsiX9herOidMAp5c7h
CwFHRqiGU0pvok0r4ZDf3hU90bqIei3sONsVco7f5w+RQHdlk+CsaMm4DnMfRcJT0eYeYD9o212F
JQkLEh0zFvMTPc4tsmYYuc3Px+9ThmbmKkVpbmrAXs00/1hOe84v4M34O5CZp8pVbyRhlxSdcqZb
A2ual2CMUX1GELuOW/1WZTGINNepk9+OdqUathry4/1w1pk75bmUQHmRGB14rilRCdMwpu6t5cTQ
I81fnIekg/yvZZIFyroip5wydJF9CIhAZgzIiAlV5xn8U7bNRj7eykuX6WtNA0QDD/VwzCXRCzD7
MeSEk4BNY4oNHj9Af9sKieLVlOup7LGb5wJqvk5YY8p0yktm8iR8HL+42HFkGINZiEK+lxJH7CnY
OsjKnLotMhGVHKxqyiqVV3r7ok8joL5oxPK6wggJXeNKz5OgahNHXQqLH+g6yilErgn2geyeBJZJ
t7vTeKT1UR6YBR0D9MWIDx3gbwdr+1zfVnwt1AHYnyso/vVgDPuNyan8nZQbbOvmW3Ukzlw3VIC3
8iv2AQQKfbW578YY48Tzt/aEmQpPzNJCVe0Uq2b61OQ5gZ7sN+6zeeXO7OzCmaScZ5rd9+4HI5M0
41yVya8IDQNokjKu9i6bdQGKclICUHhaLZCko3erJTCpCM9xCAVnKmo3cwAKzUW4OqOi3FY//wFu
23Q3nM4FlJ7Y5Q==
`protect end_protected
