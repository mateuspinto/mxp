XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E,;��G���L5a4�k��K���ȃ��Ѧ:sx���E��ĕ}�/��
7'Vt��I9ӝq������A��Ä�>�c��q)@1�v\�	��pJAL.�3tj���o!8$J �%��'��:ɹL��cr
 d�����P��I/s0MWC�0����q�s�ֆ��.j��~hun>Xfš���z7�τ��M��G�n�r�^��!���c�(d ��w��'NT���D���VPl#�UXR����#����p�D.�^#�b�߰j�`���er]�j]�1VP{)'"�E�e����v�e1`��%����S��/�^�mU�'}�O����Jp�9]�V[��$������ED��ryO��P�9�&���SO#kxo�l,*�e$Y%������ǌ.o1>�wֵ���)"aJE��o�����
����zG�8��*&����J��g:�P�z׋L��'�Xg��
r�p�e��6�,p�As#[e��)�Ò���H���8��-��C�0؟g��N��&4�*��v�Fk5���V��5��&+�L{�|�N8�����D�M�(�_�����y~oe<N��$�p�(�,_>����,�̵k���d���W'��ڣ����4�|���#�BYvF�=w���`䴾a��{M?�۳rF�_x����� �C<H��:���]�E�ݠ���yOڕݘ0 _�O�X@�ш^�~v)�耪ibﶳo�L3|]��<;�XlxVHYEB     400     1d0���e*�mVt_���@�ß��䁍�y�;-�>k���<~�goH�����PR�ը�
�>��D�6۸{�������V��q`�{�i���5#�K3�-�R���k6ao�:�����0m�סj�����
w�e�:`&�ꋦ�/:,�}��R�y\S�zk�c�!���g�Z�r�����XO;.$m�����	���^}i�t9Ӧ˗���3ɥ�H�? f"�? m�p^3�5l�S���#؀eC!~.�II���� �40��,��ɉГ1ۨ�@��#��h���Yc�%�(5���v����VB����������"��=A�:�>1���GW+�:���S�d`ւ6��L����}ȼ�dS��� �!�/Zi�s��7�>)�
���UjT��\|8%KJ�%>	=}�31��iT�+��M�]������`�f-��p�Ĳ��'O�X�F��QXlxVHYEB     400     160���W
�
�ߵ*o>�h�~�)��,$}���~߅d�S"@M}K��Z���U'��F�4ۂ~���=����џ{ɂ~�tQ��"o~��m�
M_����� ��"mڡ�*#	/���+���r*X��r��AfW��E�뜰5`!v��q9�O-�`�If�{�/���ۍbty���5l̈́��Osc2�zҴ��x�z^����U�n�dc|�!>Cr�e+����g]y�&m�б��-^�A>���W^Q<�s�S���h`��hDgn�^�WFU9�v/��[%do�+��b�+��E��M�<����}Sg�6~���	ҢOߛ6��l�$�T�s�,�,�.{ja���XlxVHYEB     400     110�3�9�\]��f���E��8����ۘ��1��+qsb��AX��y�H�:C������1'�!�"$��A�]������y5��6���Z&\jn+�`(+��Ӂ�U���h�[7�Q�	?wc���bT�WI�'�)�u��>CS#=�j��W��05���'UY�N�Fϝ��~����M��[�y���󳒍�/�9`H��5����y�Q��8eNA	�9@�y� u��	��Y�c<�0�;�y��c͢��r�*Jq�����;7'XlxVHYEB     400     110f$�DǛ��g��<1%\��9����N��w�r,<�)-�<n������
���o��J,��l[~��4�����/�w��4��;憚~n] �[s�K�E#S������wd��W �1�P�6�Y�ƨ=Z{�)���j�]�j�8�r
�g�>b�NC�:ex��������U�e(����g%�S㝰<�zs7
�JT �@E�r=&$NţL1��)�"��v��s4#x�����̎�����zΣWS;c��S�8EK:񖮛DP?�U�XlxVHYEB     400     150=��Ho,�4���G/�Fc~|R{3a[��8��O��z��	�/��ס���eH�ƀ�gf
���7	�<鄐m�`X��<{T���[ Ӳ��XP�K\�J|qX�B��ӒTl]���%|2�Fty���*�mAvp���ɰQj��}<aHI42��J����Z�־�w���I}�Q�ڪ+,�Ow9qו>��#�K�d���p�H��US_e�Z+�7W���mvf�R.�:�Le�w�=Ӄ���=e��QRo�����wg���ݧ�{Y/��*v "�+����*2aE��vr���>�৊�AaL	�4�!>��o@�h$��O�˒��ESXlxVHYEB     400     190�f�X�ns�hb�=W�Eށ�}��*���o���샟��z
,J�QP9��T	՟�f��9k�P1"��kxM�:t�%����5�Xg�%<�BX.�R1(�Z��MP(��`<�03V':x��V'�� �/�'�~�On@>���|�U,uL:��������&Ջ=z�l���1�f�8C�̗��Y��2�VQ.�a���`�8^G��k�7�8|�������'gof+#����Z�	��>�h���e��K�����BZ$J�S���3�U&IV����;	�+c��1A9r.�vHͤhă˴8K�}�QAO۲���� �eX��|N|�;�B����[�ݲN{U[��w�A%�\�U�l(�?�E��4fNDt���Y5��S��g��o�z�t�4XlxVHYEB     400     150�E�*��&f���C��7ið�4)�s��s;�f�|�
c����
V1 �F���^�9�7����E�*��@3��hK�Bu?KL� �iX$�7����4c9�@�+s�l#C^ըA�P3��G���b0I�t����d��@��h\Me#��j"�>�,��
�7��%!O�\����'_�؝�>�@�aY"����F(LUl"�a�v%���m��,cv�X�l��orL��ϧ_w���	W�w���E��\c`.��S�Ɲ6�U _�j9�!M��WƒJ�(�()&�.����S�(%��ʐd01�c6�Pq���3<y�9��W4�K��XlxVHYEB     400     160Mb���X�[w���2���Z#�/�2��m�)_RH�ǏKT�����v�o!��l��-�����gz�K���ʽ�c������d�S�zF�^q�Ґ�o�@���"L7@�G���N��J?������Sa�	�0���]D�C���x1wwm ���9Ad6Mo�p���cƇ�#ʀݙgkR낀�Ć6�vߢ�}�B�q�a��}c����'�\u7xH���Nޠ���m��$%ѶjZ�^ʞv�QM/����[J�	��?<@4Rd�9��7��Z)�	���!��b �n�Q�؀뉪�_0h��(��͡��`Ъ�Er�珻}&�b$��.��|�P��i/ƙ'��7U\�a`^ŲXlxVHYEB     400     120�td��+�v����f�/5E�B���fp>�"��Y���|!>P&��N���c��}����Q��u�r��K����d�-�<8�������T�宋k�ޘ R���6y�{7epvUv�����@n"<R�E����v��˩s)�����2KϲJ�&��kɈO�ku�_�C���<_�C�C+Y��D���5�����z�^
���بN�~p��=f����Y�q-�6�%�"��~5E�5A��/�㼠�w��]�(�eDP6kT+�lv�V�H�'��vVz�XlxVHYEB     400     1b0�.�nf�p�E]��:��|�d!?[2 �t=�K�y��ֹ��"�?�5�0�
O�d��9�]S	��H��7�{�\"G�G�æ��D-l��J�a�k$�r�%�ǁL��n����U�<��S�BkW׏x�� ݹ�Rж�k�y]*J��	G}�Wm%^wƒƿ,��f ��ؾ��ξm3���N�J�n���^Y��&ñޜ�v�t&F�VU�	�W"Rl�;ހ�|���s4����$��qZ��թ�R�8���b)#/5`zK���{H���9�!K�~��:�ܥ�9͖D��!q=mNh�V�+�Ɨ>�8�S�m�φ�� �+xa�d��W�w� і�4%����o0h:�]�Ps��dhQ�	�)�N�:�o=s�;ug�i?�*�j��P���yo��<-�@8ɔ�OSXlxVHYEB     400     1b0���]͝:�O�J瘛9��s~�*C'��dt��p.Ic�$�s�̕������8��Xmeje���H�����{�[�,
֗C�W�u�������e0ú3�������tr�.�+����f�DE�Xz����؆S�5u�a�k������]�~O���qV7��R�Q�Q-#&�$�h�A]S�_�~�&���VܵWRe��(W9[��7���Bǻp��^�Ѳ��iчtj�A)��\w�����Ve��9+ɦf/�e���߾�LF���.U��w�{�֕-���b��� [��äa<v!��SI|��k�3�#��o$p��:���P�/L�U��@rǞ�Ǝ��������ʧ2uO[)0gM�V�AEH��1EP qlVgj�v@�.<�����L���Z�'��:�?�] �����JYXlxVHYEB     400     1805^��C����G֗��sV�;o�(��,����B�M���ʝC��`�̿/��2����hY������W�ˋ_��@ņ
Ě�V��z�z��z��"�P�YM��\���ý�ϛ���u���6�Π*"���KP��a�q�wBy��9�f�$���p3o�F(O��}�È$�ݻ�+(ց��.�F�x>�p���T��5��D���$�����e�y�I�<�Q*Of�ڒn�0ճ���YB=.5E<̎��D<��V�ӝ?z�B��FBp�~wm\9_�~�0���c%q*<�c%S�'j����A���h�eE�r(�K�.�T�{���IhZ@��#I�O�����>s��`Z7X��s�=�Lq܅3��VXlxVHYEB     400     170�{�ߐl�ߧ ��`��I����h�y��~i����l鹢I,���+N36'�.X�j�;4F>����+C�i1�@��.�Ɉ��CMj==3��.ď`�j��]lх�cY�eg�d�>y�?�j՗v�!^�!JT �vx�����ia�a4���i��رR)}�!���ͩ�p~E1�ɝ���|�"fBƘХQ�ϔ~%�v$��! �vr�C�XG�:����ٷ�((����>�3��{�O�
i8ܗꨎB����o����:Z���1�qDIO�Rû&?�ӑ�9"�~RV�e��b����|���P$)N��\�R��F��|~���[S��8�W�$#�L|�29�y���XlxVHYEB     243     100�A i;�^�:Gĺ�y���i|���e6��Hⷘ}�O�*����i�v��㧞r����B���zjh�(d���'r�4e��~���܋�E�t06IǗ��PCjNds��(ĸ
}��x��Jc�d�R:�=��4	��`�m2�;�*u)�FrMw��[���T��Kɨ��s�q�p�!ѹ�70���T���vѧ��Xl4����R�T5����.�g�C���笗(Q�|.�)�z/�1�*�*�y�V���