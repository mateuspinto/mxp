`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
0USWSUGxovGsyBJteYpEoSgHX4IWV2mV+mtdsF+FsTV241EL0/CmWcunRsBCAfU7ZSBjjUq7nVyu
KiQSLd4mwJjJA1yrnQxAhdsh2yb9wnMvNWOrDIFtcfmy3Npi31DTWvDjieQINrEssNcPWhTReK2b
7I9y+1OiTDSnwt9gtOIlSQu8/2LdzB1TBBbUjMNSC4uw/t93lFFVQf+VkVUXnKy+3Tc1sEhnu3cS
xy2t9l+k1xHteJG6UR/vEtewA45nRIBMJj2dHcDlmJWc4kfuV3THB4h21OPUFEpOcOtRwgJwcqm6
yt9GI3g9IHsOdCGcNN6l252mXSIDx41+zEWStLPFTKWL6vBB3PRCoSReXOGGmL8s64nJ/I4iuiGb
cVv2U1MRLp0iEbzrlF/mjLicEb3yY+M4UNXuhfT470q3YLgWb2qfoPqe04gsD67HcyHhIRLpy7PI
hluNWYBkxczLKDjxJig+a3Us10LhXn4jxuaR5GeMw4syvnBz5hULpV3hvqrDfmpg/XGcIzbDZA9T
ARluzDaJjnS/7GxkDYSh9UeVo4UNXLZyy8flA+mk1eOEfbmoKhGR/3u9HbI5ZdaU6lgDMyI95HHI
4sXG9Pid8coxetHimSkdxOS+IDOY0TvuNiwyTKUApA9gGzXX4XAUKmg2McS8Sqn96sNhxM0z1+4X
gfeD1+UYsXWFXOdhOjK21ToH6YQzP5FlsEf7RMH7iL6hgLJ80omnHlzoXSIsNPCrU/0kn4feACau
SWoLtkvnKI0u74maJmzDyiRCsHuC+fTQ/t9a00iTWn3tmNbxNLvt4IKL8yCyN5nONWNZNLMyjTa9
3vI4QjOkEaN2FI1WbIjEviwwDoTcypjLSmySX2Boz49n842KIqXbxFtfTrM01vVxy73y6jY93V+k
CX5pHp/8lRvrJdIOXPHkmLZTKQtnNUq/4QpBrbkdPM2VTc6Ky4onRwjQF2fY8AgHhh9ZeurS9fkz
STnpcD48YBSPfT81CVPE/xi+vRSpqlKMIboDpjz6D27D6or6+aYcuIWz6zcpYa32w8uCke5exPx7
RJz0e4CJGpEEVCCfSAl6KpiWHRJDDvQFOl0ryDko8OXWHscr1MI2haJ98spqhT72v0sYrjRjkiau
Cp6rrx+dUByM18ZfTZHqi/7fb0viHt2Cwr8Wm0LgPOR+HZ7MEVvDqhTVmU/uNKU31Uo5aLP9z4GI
qq5J02g453OZtgvXxESbV82YDJp44IYPTxXgZFTDunGU/mjtg2uqH3BsgmYagNasGVAhUJi69bTG
YsM3hx85hqX6SckxmEYT+/y8EmyIN9i+r0ttufSqHgcv5btET9Z9bLQU/PgOQY/yNL0ENR8Kr3cN
cjawmc8JwGFLAyx7B97t0bC46Ex/rUGs1/OavN+oh39UxqeTl1nLuiUoMQf6Uz76kksAkp5DxsMD
suGDBjMNVQKnVGAgFX/u9Ac6zzAPmNi2v/lGo/KCM9EuHujly9sAoleh/hN7EAHFnpSMCnCSULYo
TJLo5RrmUWi6pc/4ceU0st+BouVd2Jrz7CfVpMA/kc5eEqb3ZK8U3sJ8JqWgSvbgglrj6JnV3X90
TiIlSoLmBh043AMa1oxNVGd+hgssn4tPvNL6+BMtnuWZnnYZKJMHvF4Mq0RkJ6GybXlqquiGFcEo
QNGTkIweiXHcSL7kuGUxzctYpHFH1GgN2CjCDNBdm7Z9woVN+Wxo6xL5U6AUmFjmwKm/eBE3BPQr
W/1YH8r96L8vewNZP0DYifbqjdatpJ3+wyCUc7j2GU9S9R8+swKBL/u+8VjbkIivEQ3k9D+WjLr4
l8Q9U2fWVXJ0ra7SnMvd3KYuPNr5nptjDPUO7cJUPbAPcpnegCNFlSnUxlCcq2vt3Crh1iFYISqi
DNM1s7CKJ1+1iqsqtlmikbguTMhlJAWTT6Q2EkoOMdiYnYCCGiwiRdEghoKUJGOPyYzsVBxqmsVp
T4bsyiV0gVQPyxpDD6EaUiaRhuobnwNjvcV8LpNScEy49+5436uSK9hNwDcMoY6Jsh+UHQU1On36
qXos/ObyBL6F3VWjsoOKspkP6thTdFrwkCnBue0hEaxMKFXhMD0+CbHX3rrZrHj8kdDCOC0r3hqs
s+GF5aCLe2kn8nsAZqTNHlhp0st9wnBNdrWhprZCmyno4U5c6D0aLOueBZsZ/hC45iDmbGBTLDCB
3tVay9coIBQayKH7sJpJM9c15I7uqrEG9zz3uCl6ZzOpcr52fweDEgRvzjMH6acRw77BKXyb82uk
FGxdF1LQSl+ijdDvQybYATSXYN2KCy5MbwbCbCsye45ivZulmvHKpHOyedlsLG/xVso62PNIkPe2
q9YnlP+/+Or0V1Ktn0xmtJi4YVQdV7m5Ij/qWTaJzc5tby+62dtuLJ4rZNWWA034Bfk8g9XcSuWj
qpumVGVlhYfG3/DkOW+SWE155cDndcf4qN/a4cRQikP1w1ckfy1x78Jtj5zjQ8TsSxfueN6yrxqw
L3ioFZC7wFNt037f9/+Q9FgyAAXpR+fsuwMqpSXJFiw8X2RAiiUp1/jRXG2plEEJn9VdWbYx+FRE
jkFv9ouIGko7Inu/E93SbjjRVMxSGctRwKuIp+Hb7KfIVLSrWils9gbV8gCIZ+wGjd81DUJczAjg
gGGGEmiJEVNf2jXnoubZoAvrRfc7RN2mFNNwBI4WJu+qlDCr7IxjyL+Y0ks19pABclyt3w+ze5KU
tTYMoWJVasuHVkvTs17hFJVhYORfnqHvmbPpECJH13k7yZKAw/AVKYYNo/xvoxtfg6ThBiV5/O28
xsLzbwmMx4TRdtWtoIswWiW8j7ma9OawauT7kEZKc2zfPh6O6FXX9MiqgutW/nB7o7R0FzBMfu7t
iD9DY2UoYjuRE9n46Lh0rgFq1yYJC22Frfwv0oBt+1FyjdBwPvKYkWTUGik9g6GCaGSFyX+wT/uC
7rg8PlEH2WDe/V0pV1RAUy+CuHwuPFYj1HWrA4b4/hh82slarq0DsLpknVLbglnSnTK0iEwTbrle
IGE+2srzH6Vl811S1+rZa9VCCyZv2oZZTqqNj9vVJUsz7lW8Ef7++DrJm8RrxgZ3YekxCHfYCVJA
KdyyKQNP/WKlHDzaFgRba5LDXz55zz0D+BmTe2ewabtlxIebsGlb4tUd1DH41Z5dPDv5/y53Zl+i
uvCui0Iv+jMIqxrw/jqb6ouXqN6eBpaKaXULI5Dyeh3bLRHNCZFvGodsTDQgavN/58g9mwsaxc5c
CK4w9Vs1ytxiDrGpDJqFM6mldvCvNx0Bd+gC4wo45G2UDG3ot19VrtOmVJ+OrQC7phq5X+Fwj0ob
W9GLqtgfB0TMjJ3ynz7cScy8lD94xZG0Anw2tqohYYj9GCnZSSVfIFNwaNuWvEBGfQft6b0PyA5T
1y0CWlu4vYDBVqKP5FWkCjleNFkUVcJ6xP8zYH18dils7haex0V3AGRWcCT17JvYrSmw3mzD39Gz
Dxgk7ZnRsOc69Z0xH4UDlyS2Q6Iu4hyEL9rYMOukBW1U1sIgn8JqOPGioLTpyfGbTSBTPlzvY0lZ
YqeZIpQag7yCShqS7pdCEShtg6dWO8/Xl0ur+liyDPSwZ+tX+MdQAoSnc0ivPG0Mvqy7HfYTsFGe
QhLi1vG6rwazQ6MmKC7fJsQ7JOmZv+QvFJlxMZJdblIM7za6slLP1XOoZvji6kY7C6+Kd9y+dldu
AEHyr/M5tkZ5gSeNF6rGvmofpCbb96aKtbfeX49J09TRWrT7oKVIHHwzmcHX+bTNacykKPonji3B
e47PxY+nWP9Ga8BwcYHdQrU8cdBCJsJL3kckLFZ7LM/3q8K7L54piLGIXJ1VwKlsRF3dQ3GRfFX0
jKdyk5hhTEJhsb08THrQ99oqQVgcKez6HqJS4e2BKuWnHJ4CCgkrRzj8zfdwRMXDYOQgkhRJgjaK
xE4uQChmYSd2xyizSzl3wtUPs2Ga6WNj+9ZLv/O0uJjen4rgkXmRvrpK357ffaZbFxE2tBF43eDp
ymGPwVrd+tsd+IC1NeZlIQSWC3/E2gbGPZLbw+1UePDAgSU+AnblolcxCEf5D43YrxUkC34/6nhE
UyqP3fUJ6N8vdWlMz/v7Cili6qNfc1YzI3FNyyKnz1osqotl7fzGGkk0VJhIy/07I1bVqzxLpPIt
Pq95jvBa5cc1V4nq9j1I6YLA8YdqWYlH0VpbRtbkx983rigZojJpvhrjn1Rr40c9vQKG+WCoQ8Cj
v0K6XYoofWMRxpmuEHj0udOX3o1g1ftqmAySJWG3TVQJlPP2WiikMg5aQu2qm61ZMzILBGG4n8Pz
iar1vifuIXEBG6I0tKfOZe3K0ricET+nTJIpbroO5iORViIKKyRd/RIbsFRpnq1cBVM5hGxnO3Yi
dJhxBgrrL1xL+itoo5WLKLK0rX5+u43NGkypUEuqMXmJweuT7TOUW/qhLUki3vsU1QPMINq3IySV
vnD6AVLSqwAtFh9+wmCZybrQAycUx97hlZWECjhuBffpcnQzlvwn3ijidsk/LahqjXydwvS4DtS2
UnPNcqBlIoHB4BXNGBumRspZIfqQJi5JQ+LsqCzSbWC1F7f95v2KaRw17qYkx+FsMnhOTAdcIqPE
63M9lwgau4u1HD3Pi3MedwTpZztGgnmhn4KiQ13vlPtziTaVRrhMMPkm+Cqvhso3Ju/TmqfLz6tm
3kjW7yROWzT1RfWFmO4HEBbK+VsnclQrjFxq79iVqNiltP98E2nK277sQPaYqVMkCcNieK/j0YlU
sXcXfABc5mpXa4BD1iu6B3lJaBKd2WySHTagabkfJoc4eJAzIDsnDzxIHJV0zztNNSzx7V1Wikwm
moYQ8uNKO/pkyANu+6sbovz9pLk6U3HNCyPogPUIqFYxhvaPPY2UN+CIe6ekNMO5NZ5q2plun038
ADFsJrl8Y8v1yzJZfZbAHpdWsldoljFqpAI9ZWQuhAW/1Gn3eQSjDD02GbjcotTxfGy+O2Vmauts
G0zBwaGS98oWGCmuYnVX6GLQQ42LT4OQ65Stj9tVtEV+6jkmQCTVMeni4h9DJFKuw7aoZezM13FY
v3H2EMFG9ccoTpuFaRbwUSqo3C5fEecNNaqyLc050qD9wbFfaFUUvZYV8vPB+raJ1T+b4k2+XHdV
tguPQKPruHpRDzRrvpJtra/wtyRp/gSkGf6wRPUgeqvvDCdHXdPjQlyqg7hDF4Kv/YlVSolHZm8b
jux4F/EgoFI9mZ8chrfjUp4V1HVguXxYw/CUzPqzreZULak9RPuJTnNR9LeIH7AbTq12ZoZvYjbs
h6ncEUlcGSc+z6zFC6DFpEbHCMQK1ZxuZgyJH2Bf01Gz5lB5XcbinxvhCv8pleuHPthxsMiWp27b
1OY8iSFQO9GH/uh95fj1oNhDbgzmiz3KBCMDGNXAgoHDTMqhk7coNaGCBSwI52xm0cIaaUDch1fU
MPm2Y0x7aD2wyGXU3a9RM8LvRmNG6RhTK9t9xvPOtaHRdt6xeHFKS1GEoDC9SwqEy5PGgT5r62GT
BAdj6k+UiYgaw9GxIC+ZkRjRcmAdPKn9aco/rlquLlP5gs/CB2HQRlHrqzNZGi61hRDm3ktnmHNd
/QhuH4Zirjj8Xquxctmds8QVcmQTo/E3m8WAI5odh8xn3tTnm3GAbj0A7SHUiZAeXN6otOXZoVdi
zZdw6JjinNo9wbfxUhXrmGIxI3rf3DY4EmpuydGeaSDbJWb4NOHgKPLB2gOoC2FHzjTCsaoHY7gr
ZJbi/llDOlmOwaaPUq67T46zRqbKbcTZLjQJwRADxZibYdMRnGLhycHXieaRRtC0Lnnn1DErAmCE
TmjNbGjBpL2Es5gB4p5Vd+hPfq1VYWwooXIi1xRpvZvDaftg+qZkhdI4wkhDHZkVUOM3FV3GzKNU
OGcaDvIDzA1Z50OI8r5P9W6XO5yCPtcGfrZoITZSIBr9tg5KndYabMA4PwNgXcBBzRfJqTfLCs6d
YXjVXD0bRN4Gh0BNdboiSqFT0cWAAFfXsKcvKZud5HVQayZDdPuPaiPXusNDynuZ4yanQ3B7hDOU
5r5qwOOeiOfVshkLVHU6uLdck+KSwgozjfJWKo5NuSCSNp1lDhRk1WVyVoKvgvXL3gsPTHqA+Xvu
qo7FrVcSgK8pU0xGpNaR3GJVVPUw7o/vcAYEqCOOaeHkSU8CMN/9E1qVb1mP22dWbqC82uDkbWxs
xxhrlydqJTYA+OgwPSLLde4BkRhTbHAh3mfsX7SvEUDYKxJUMp/YQHeLimEJVrz+Rix9uuBXn4/Q
gKtYclt9EW6DEMSjpSYlkLdogQ6vO+A0xSg1ztIPDxOvNcH1mZpuAN+eJO+LaandXOH/LYuOblvd
Ai6uJJE/8bc9cUxqDyBxOF9m8NDJcihtp7OaixtCoxbzjK4butRDjw7ZnOnZgLUjOLAAWAIRxUJU
5whTbYLi1P4T3IOJMWbFyO0GDDKUQ9/O8JyxdZP+Dar5SIJ6PprI2+gNxfDf6v6Dfecya93vC8Q2
xmGqZ9ec4s56X5KaWVkO8Mj6k6z4iY8sdI2xur0qcWHdAADQBA3ZwfZYDPDfEVXSkmfOEdTbib66
HTBMfAFkwqf/kMGDfwjyB7FpHB7HDjOZZj5P3LeCGPxm5SGkzHW96zdlHtstOoNu4rsCoZW4+PFf
Hmwi5CD6a4GZSWb2UetKVpHMcyHfPVLouCml8K4933zDwaSviH1KTcrzXv8HGYGuDkikseM9S4OM
0orQEja5EOTcK3S+XBJNTgeCNzxW8yQEQcSQNHYFS15B2syl/TvDAXYZlsJvNOLZouVSOV/Bf+uE
OhBJ7kEqNdbQ3aQn2ciyvamwbndnGne9ZSdVnOeXVR6Bw90vMHTRwf1S92xiD5I4+/XOguHVxwkA
8noa2WhsUXrvU2sqT1owbavzLF/kxBdXcPkuwWpWPqwuXuNc4ZiGb2jGs4jN/0LXqAfHKKvFJ4DO
KeGZmRfZKHD6bPkIxCgXSLyuHLiTSUoZupLXx120v5FK1ysloi2jOI8EHXVHBPv1Ph5z4gYPi0mC
VuJ36A208bxtCw8hrbAdEziUUOLvbpZ/BQ+t6IX1CqMt+f+BVNyQoi8TyaAMr4IJ/FB5ALLZsLhv
K4FHmaYdd3mo0iufKtTjw7sWYXqL88wXHbfG2Jp5W1zC3J0cRPZPlhUphm0IAr9IBliBoNEDDOYV
TFO4aY+kUS/FEtvdAI8XzE0VPyfpvTjp/4RmCixeM2EGOQHzx36NKk53rmvIKRdiiiVLwzEDifl6
yjf4itTqfjFtltkhuzgHGqu0nCP8LmQtlIbppFQgbZ2aGcYXEbb2IS4Q7+sF04mD2vdMsEOKarl5
mS5Pzqe95cZvmHHta5oeN1eC5nTicl7sT7eI6iRgzTl2ZCK4SPS6Z0Pf+YYgCq3y4usQ4lTiB3QD
uLsFKgHi7Rn4oInwmSSxyqoIQ5Kuxsszb9wLLPPCZ7YrUaui9F2dQ2lXQRdNdGy2gXuLzMaD28/V
pAokfPn8tabF8VHOUH/UjkJXe+r4wsO/rV7itgJipj/BQX/ugUQvAt6f5dWGyI3JdlJEgMWOKAAh
51hfveysLbcSo5qgDpZ2Lm9VzmZX217hqObP7EFDbAQ04+ZmwIwTLH9d7U0/nAMLLvtS8MNyOMQZ
D3a4pZ5L70RlrCqdJibhklrpLLX/GQATAk4LEQRyEko9iJ0KCYW5g15nNa6atgPQ+DdyXkJmHYue
c8MHRZlKBrLrYfDZUSh/f3vDu8uUJ8W50OK2o4tQG/MXhFzhPyFojCxT3YRENfk4FopbECRCp/S3
wJvnW0eJ9d+mrkC2qiA9RaKzKCk1S3wfAjAu4HiKDQaVU+j9xoXiKBa9V87GzHA/mpjGJO2rwbhl
cnFe+7fkKivQBEIw3YSsBZKmXfzmkb6p7MUkFOgD8rZLlWeu9jvHfqpOg4vhLGCBexqt8cVztMg7
JYSj5IZPA693/RcnF3CGQhu/Uxkmz38ah7FCCl55lppUiQ9q+YVhS8KYUjSnbzWf1/h7olNZ3EaG
2IEvdN5gXJXuFvQNr8oqDty6eH5zTfY2EC/5e2rNZdtGlTNWSSJj2obbR98aLdMDyfLc3Pr9hRRD
wnqCVIblsw/YUpODzEwmZzH6RI8rbMlUnnc4aOLLw1hqN5yMwSr1cJ1qFHc9p51Ps7jQ1rcoAdeI
o33R1yRgG79N1Qk0Cy0Qw7xSfhZcqOtGBIVRScYQMiCgDZ4BKQRnJ+0VesOtYM+2BZPsiXozwilx
fCa2TUNA1GE91AkqAHupEualS/dk9pUlaOuGljS27fF7XPkpIQQmLq0xHzjtB3d4byMR7D7f7g3w
Vbmh5OWPyIvBJaxTRg3NLaJ8ygiNOr2Q9MFO/P+3DhzLhXSaOI32FXfFLdKRt9onmxx51qRGmwOl
jszekdZk4tgBC79rVfapRhpMgZup/ndh2uuAMp0MzVmTJqQ765Gji35+xa0EYPEYOBcZv1lZYdFW
oibCrX23NJAuihwtuBdHQStL7eVW6thleNcPWCAU6t1429i/vubBA/1c3c6Ippp+nQTGMcJtUhHF
oMXNhG2BsiWwi3DwfOuOrH7eb4/AZZDTERkU6uGMioe2xLXGnjsVB1+TlueLEvykmDI6wuCWezdR
Od8zofpytOQ04UP+2y49coDIqvSb9eidHKOr3pTJPC/jvdpy114e890wZuwkeDKWMjL34OOiQp/M
NvTpkfkiq3z9gO4FfndR3j4Tcs6fcUmzQni1L5DYdfNy+D8DKJhY2JMaAseytNOSYIK7+qo5nvSC
xkW5GNqHobYRrj74S3zI1N3dDeW/jIg2K1u5KGK2+xiHLQgKpugRNwYE0ytnN1sox0B+qQIdNFg4
Ww7tY6kkAu0KLo3G3sjENe6I7RwmdO41J1+pRl+F7vWJbiEacXJfQ3Xz1qqwf8ZhUkOC+94v7ZMQ
1jiQ0HXeyr+SybqzToV5fbYpU5WMkUGpXqnRWFtyMLm51cbwqXey+ss/lK0LA0NqIaHwhL2I+irx
VlZbn3qj6+LCiZDabqtb6FfgJH/slFa3uG4MUaUBaF03vrzM5HCEO/+ZHCPOhrqijvOrnPG9zC2F
JhOapwM68bi4vOsXjVl2ZJF2u5xO1tLzgN4YNWN55Q4APbWv7YISFFCX0HKbsT+3lt6Q83MTedEW
k4geeIesWmVuP3jI8kLKvfnUkcAwvkt5X3N1SezWLbSvfSsfNYrrwvkbt9O9aT5HCaT0erQgKeoe
MDtW56kdIW8S6E/oZTDy2DJCxnvhNz5+LTNPbv4ZNqmMhUVFBuJ/RWmTSm80H+LBSzIxqCnlV5Bw
PG8EjLEZvj9sCCOu5UA5GgM2AHfYMCe0mt/3cyttuPybl+EMiZkTh730i+elWag5Y1tJ9y72Ai+j
rLI6Mnxo2nP1LqjPx/O0KNIuT5BAZ91+NJvq2U6SPZgz90E55wukYDRr/GmtrmpfYGvzAS5Y5vot
HLpfM2gHRHNHBqDiFn5NxFlrzdPkgEkC9LIfQ116+fAie3z9NfLPxQVeaivD9wJre4txu/Zv2MKZ
ZhpT5e/+uqY2VNFOyu2FvLEBAkhX520Aj+4qC4cw9X9UM2lyC6hz11juNCXAprqLMD0ZQ8fXPh9t
XTWYYNuWGlQNMfoO85gJG4vOEwiuZehJbpktWCgGBOQcTZHS5b5E4LgStiv3wKRP3z5NRpJ3W9N3
Lnp7hIP1uEUly0BnHxAwFMmom0Bg8O00GHB0SzQaQPlD95YzGa2+Da0hcSwWB/WBa8VGH0VYvm7b
6+oO4+UZW5NagcBqqPmAfzrij6RKDwTCHRyOJ/Up7Q70fxWr8Rfddfr4eZ4LhLTznEwZtOvu9pn4
EVLdKgAPNIZ6EvwLC9YbcKKFV04RiVP1y8DW6MwlRd30DtwmDxJ9vTC7oZ/BoZqBSk1qS8IoB4Ad
gAj5dU0JG//YLnx7XIbRJAq9GVV3/YjZST2/XzdvD7LRqky+Ve56ycR8Oe1SXeXLutLh8A0kgTKH
SZQAaPHhs/UW7yXihWM1wPLdVHbY3VZCg07lRv9btkpHqzuIdJa3Tgj84iwOYa5eUwPxHgcSCBKb
E5I4GBCxyeoOO2w1JS62loTP91wJDKOTvxJQynynC/MHE97QMm5BApdNc781Z7e7yXDxA6LJdFEG
i6A64LNhbbbdO6GgmTlL1lAfczTulryoX2IL8qFXHxxdaBxkIeoaZPDfLQWD/x7242NamaUX41l7
aKV8yUFqqQsmvIQ+ChC9RSu8A1r0j3Yh7NnOcGDgStR4tmaWeZuPfmSGgqA241oJgzgfDgYXSEHE
XzU/GjL4cccoimYvjuoxiZDWVv5PRfP94JCjddbsEH2nFxEfR8HqdUYSNlvYnD/2HMdkRO4v5hNs
Q4/ZQCoTl3qmWofS94Qc03xiGT7jUbF1CkAbXmurFx1prfLcmEgRFTolknHpEXOvLLeKqRfRUpCE
qOyLFk7NEAMGzuD2YEoiKEYgafO/gbg4HlmoYU0qBA2aI6BqC2vMTaGRGmmCOvmyA9ROQFXfvc2o
m/GNN276kTDQN8ZuGFezixe03qwpIxLm65woS+VbvnD3LR405vON/ifSAXqm1TCWWlPU8bxxsJ9h
vZOEYbefsf8a4NejIndufuGtKt2lIU9vZUXOvpXWV2EvqaXnWLREiFubBHH6HVD+AdKtm/XWxQ73
F41gRVSgCkzlgheIM0Yo3XqDsD+k1ST/ATUoDUwK+INW50xjFRI4MtWFhFPzUpCovBPN4LvjIZHa
NwWJq2HlmJhIktMU7HJ6p3IxKlQ841AOTohuwh2wqN3Tig3JeKNEEaBoX3te5Q7Xvd2+ZYI1Wi5r
HxMyPKlJnGMzDzORZxVYepv4YsWUroucqVJQEQAiRqx1IvQKQQe44xwem81U0fSjiOTSJpzuzQzn
IgGzEZPv4dzhb/eUEU3LAYJMpgBalYKmqgLRVC2feYGMDqVlmJSY4heU7DYLHFRw0iXhiNtljN+E
W0ZL269VYXJH4e7CderSOXrL1oKOyUBHIMGbgMwaAwifdh6COnXNVqB7ZG9pbhtyRWr8qUWsPUxM
Ms6VFLoWNFMayvMv/d+4F1MhJGnOarMUIm9PJxYw/eFZ3zCYRi8s6qPHrWtHB1rCPOWKYplAXPcS
uZZl0IhxMcWSLKO6+SyR758CKpW8
`protect end_protected
