`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
cHQK0/Tj0wkQ97FrrQnPq9xtT7/FnkGXkwBmHqIViywXnlcNA1kWr8bpbx5dWU7RHjyjpbVclCQY
FlAHSSn5UqEuKCL3aLRDgjefMWxMdqtA+6m95GA38KVY6SCnLefg2dn/ktaPC90GPcT7FehlbSbW
va5I9L2baz6UB75X0ztJ1QsxrijP/LrtEA2YuT/+QmSfghAarcJ3OUHO/SYlSA8Xjpg3Tx1aSYgY
bWy0NFg4RHlZluR77YbbKqzS8DR+wW/jtFPt/oE9dZwp5u8Nb5M0Q0/ZBThxvHSKovzyQnj/iZQU
MpXUYe0zcZO+2OyRVWnojVQxAMxiRVHPTjOGUQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="viuL6XdNgzN0m0fij9cRFr09IfEbdh53as+bK9iPRb0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16576)
`protect data_block
Sd/zIRldeDrXV9z146UJkSQj/0FA5y/X3Ij/52TpB3n8/OKEOzFmRx7S9H1/AVtCv7sTuqsBwVHu
X0lL62YzNsYMTtGsusi+f0rp6+Qgl9B9hMCuwFO/Xs5AKcgFcPRpOz1oExtCAta2q/sCPvC1UNjF
hCRK+XEhKtuBJ8ZbfvtNUXQBUXDEwDEozppfgCg7mYc9NPGxN6SuMx0XhMaXE8kPDPsPN1Pvj4Sb
uv60uvvSkM5LKCyHZTd4PFLyhETQuE54Rp6r16ksxZFAYsv7SfCbB4S2rENLfhCtl/cZxjFG33eh
CudQj4AxLQTU3b6DlMBMNMd9BH2F4iEFU3HFbL7tx6iRRUmynMDS3KpPoQ1he+jcEOroOymUT1Uc
FJMSpSd4YaD3ECQYZHO1uBexokR6EcAY8qCH4qEKA5yrwAQIPXfU3Tf3O4TpcFmYG3mesMdaKmaE
Wt2Ni1nVc99QgvIwC5Fv7NQo8wtWmO6Hkhlgblo4443YcpMJUJyd6AFh44njvP/VkFFIu/jo7toK
FZLDB5aeasPtlzfMMXXbDgydvtQOjke1H/zoWscaG9Ix0T9qThKvm+hMas1NtY472GYHFF8Y3PvH
HWfOc4a68UP1XW9aQ0w1Wmc2LvtkA6cma2Wf1vFjSmnQaMt4OzlhCLcEy4vuhO+KMfSrjIB1Y/Y7
I9848yBJ2zcyQ0nS1P2Rwc0RPIyHCi39Br/EX5g6aZC/wn331Zh9LdPU66XEQBlU3Di3p6c66NiN
2G1ALVrOj+geakYDKeFPl3mgseHFgA8h0GASV2+35aN+iA0rUKOumcVexHOXzK8mxNyQtxKHxTp3
s15EKW43fZGif4zHfH179lsaPq7C/hyZr1oqFjmUvhOhfw+BvUh5yFoAoJ9Fm+XQ8/e0BNCEvgH7
JvHOlvvnt9wFUfUUTzlieUs5wCzl2am77ModgPXAfrJ8/Ijjv5Nxr/A+rsBJ6qVnHCcCxytjzMWe
JA3Ak6hnqTV9IebW55i2Ik0TNlKlgzV05WZYnw7W1oNpl/Zpdjd00mTEIA0U1EBiW2NdWSFSjz0c
1itQ6mYpsPs+cF3sTc0NpgU6zEfVxobPzoybYODTnuedP40unvf/hWt70qB23j9FvO7L7PbxWOko
WbhIdKHREfaklo9K95hZYSYCP9vycMc7orbdRaMiT8oMUis7wsgR18xCNbF4InDuq9ckaTXf8Jqc
yleKG7KPC75fHexMuYUkOizcV4PD7765mNArUSgjTAE+ZKSOcwMAhK8b3nLotCcEUFa8j2PC+6tw
n6ltqcP+VdO03kMI3KAU/nPGbBKqoqIyciusA7BPFi2zvoSZfbMVIbCLuIKsU6di0o2EHLbgZ3ha
p4UlIK8gJfw+9q+S+q81Xel5fqW773bJanHX1/upmWHpxhGhz4XGy170XoCSwdsGOl+iljtOf3ov
hDGuTwVavYjUqmfniiuXbGiXwffNLeK0JV9T5HPm4RNVI+H/yy6y33RoZbAdk3wtQFJgSZAZlRfC
LZpoa2P5/XhU1tbrybDfXkizLDxCcHqlggGtw08+LpRulSjpVIVYBk4VfvqQVP38HS4MB7lc+v96
gsMwNbEUDjiKGm4rbV1ed99QwiaMtVKFufcj0gvSYZwraVgk+AkynXuAHR378zKGfhrGvNlSBywE
OMWyedC+iGb5KzL2Ym1+UjqlNsCYRwEh2RPjdAYdLQkTMTB7qclKxwU8oubCmSfOj7ct9j1wMnJ2
juYcdUaFM1VsTxSHle68xENNnOLjM5IUGQ89gpuMxiuHT84INKcXRI0RxeWh52tSGtiGXHM5A7JJ
Hh7u72E7xjLNYeUL91RhaYwlxBIx5S21jCiH+yOUCOD3oDtsl2qsnlg9HfkT9e+dINOP+XFzP+rn
EdjrxSa5kbGNZVgmmvPq9RTDvuZYSN4sQMWdzSeVB3k429r+gveSuT+qejipm0DX+0AVup+u6okH
3DMbipRN5NBLOyZQ9mcZkaLO+5XQAgZstDN1Ta4EpV7JYxWDf+vItHVUpyNW1fIVEJg0Sxu+f6wc
aH1OjXD6ZBs7BTNaOe7zdDDJBcHp8TDbZ5z1FF4e7UT7jjq8d0MfH3xVHZpnx4VoE0hZpVrxovGJ
UpVJPy29XhwY+HMcmtzhemSUOIssbU268e+O7U3TNk+FTwH26rKkmQ5K7Pi6WeK0/b5slX4j0tar
OjiXMTsQqxG6o0494hQ+OC4m7celePloPd64BrtKb1dRQM6deXmZb9Xo4PFBgPYhUhNssEqL9YSy
ZY09XrmXjkKIQycIt6h9KpTV6xidROKfBxxDDXiSXEKM6N68l/26ZEy9iiUVO/f4dVCyyK//JDXj
j0JmOl3XBiIvHl1N3Q9MX7K/DzMmI46cf/EjaP9nF37SwzovKNzNnPuM2RWpZcjgUZZvIbCl1wGx
VA+TNTmUZ9P+KX4i3VfWGVVQQOH9FW4F8Kutn7ijxi0+i7EIQ9AAwWeJOmTlZg1d3G5ni+fq3TxP
9B+W0zCl3mxdJq4mJVY/u4iZuijh++MAupV8g+z2Z3Srn/vybOlMeP193fVi6cnV8uP0vZmiDxOz
Fz8xsoGSKpR5dJcCxK3WKSV5JDy3d1EFiPmEIKlzpTIbBEyyuM79dB244TXqcba21MNn64pOYcUS
8lfrnMvIN+ybfUYqSB2UnjHixq/UHntv2a7fv0mO5VlbbrWxaXmqBPQUKY+17kbJ7BPio7SEIXrw
cp8g2iNDOR4KxZJQwM+IEUcQZANlY6uqKgPVvbT1F27PNWtcIdDlfoqCSgWpMQmWoVXFMIxC+wOi
dEOI+DJxUMPNKbeqLuSn7mGj5HuwlbcaaxmZwm+0Sth11i4a3A1h0fnarq18losRR7FBFypeAYOt
nzf0gesU8ExdvNbdXuLleHvh5IdPKMotDMl8GMtCVe4HuijTNa1Yaz3nZ0XvVOKVOSjMXcqbdnPL
7+VCF2RfvmxgvGl144SKz43a4Di1cQOxxzeF36jOWOK74c7I9T8BZjPr2WyslexCR9IPXTOApGbh
FpEZFbN9Hk8jRrMeS6TCm0OFIphs50ZeLQO2Kx1e2+bA8Akl94tBAFqF2ExL07mssvEjUzKltcmx
t5gCDJButcNpe/7LWEFi06jeqcP6sP8aWmQIYE+4amC38D0PQC1ScAyo603zJwOnVuvwcAYnDfW4
5OXYgNNls6ChXld0PVC3IcAjjmwa42bslOXKOUAbqcfVYJh9agEDbL1V9QIu8cM/BxkaVfbEVAUS
0VvBH+0qFJ3jXFQuvAOpzca4BVBD1McDVU899uiSlysd1SPFHrPX8DhGmyD7wXOEvKNRE8oGRvF2
5ulT9V9WclhX6WbcWIipMF8KlUiASoitoZfWQ1kciKVDd27vquGc6InvnW6vI7sOb8fDZE+WeS45
pkT+ZZEt6Je9ziR3EbMq8h9X47bf9DCw08GmhFFkJdnsHvhNpIfNpkb++fBmIjF7DoHZvCZk8gAo
2EBaDq0jtly/JPAcG7PX3O/tpLCxwwk/nhEYhU56QxQ/FuNxLCEKJhRT2i8bANGHvpM4DWiLMlXh
mKFFC7JtqD14dpx1uNk1Oazppf02i7OHgg/OXx2i3ZPBcHs2tjt6iAAcUGmTZIF4l/14zMzquyUj
dUGU5nZ7DtHmYtV1D2u1FaUyW6Ea+MsFgWqrjzdqonR6T+ZfzAoZ9G3OhgOQH1gy5ZFdSVrpMiY9
/5ESDiDxFi1rVre/uFibNy6ckfwIAIjQs1go92Dpf8Jx7FEvMB/A7Co/jrwStDAj9Pq+bpiIl9tQ
bt58yDksFP5ydZXk7BBDL3rXrhjIBzDfLUZwYt9a4NbYMy9cdIBP1q5GSaq+q4oWNI2/3FrBd//U
I/BzzRAa4f75pOTNobj/9igpInhJ+oNl6SREak5izhf5U/35bKwLvGki00xFO+Kt2f9qfVVrtXpr
NrMIrYS8Xo3Ie6v0fOIfCNREkMD6M7ZB7xcpqKGOjADsh1zwZS6kTg+B+ZBnCJaYlTyATd4RVD7T
hD4oKeimMe+Pi+gNS1CCDR96t7Gh1jQMRGwcPSgjgRO6ygcYtldodDyQ8rr+q6N5aTxaIXcfrZPC
t63CAgloUCiO2CvULRV/E4wjXE0+gTOjIc0WeKFoiQuo6qg9FloXPTufAI+ToPDtQ03TeaOh7nTB
U8BsARXh6ofz7ddPrYFNCGylncpqGK0OxJuprXvuQtAX09ZOOmiFzQez9wrzRYwfrBZYmf43C1u1
Q+cdX+y4xHq2fTbTzQDvItrLoYwZj1yp/W3d33UtE3YwwsZm/NRVdqK8HqRsX167WhH25gxY9K7v
zdzAOYnD42C1o200HcUmXF5TBAdTPzOhB9y/g4LbzEo4Pa1kTH36g1CgRUqUEc15/UYZZsh0oruj
JtXvcubwBrGhZRnFWe6LCaZex/Js/TfYHd4VKD0Ko+NxEkG73vDbHC2TIQtFC3tvAAUmcsGsDHCm
5es7WVoTMzBiA0F8E7uBLGVb3YzI1PMEJQTAsUO5nkc1Vz6RazLpyGZHm5BcdojwqJBps3ZZ4H69
vb6Ay3BZXG0nzptmHnfW69HDxF2db9eOvRd/WGJGysBeS4KqUUv2NVBpTNvz/+FKY7Pa1NF0buUv
vmWNKwdko99pKaLHu/OxsObHPXYKTBi+6dsZSkULndSuJtCgfiIs3ct7D0TAPoOgkoCdkotPPNGI
HHKCTK/1d0t65UYWsVR1jkhBVUFacInF4tUTebSpiIOdt3dPuD2OdioW8msYPublHrZVHc7NvrGp
9NrR7U+41OtWxVdzg1Fctp6kcgqdnZUqQGLyOsPug2MTRvaKMKiyX+htqADd22S45p6ECCUfsPdF
h8wbGo6P4Fe64YU8rAdxTv2RIwZJUTemqWCrifzu0R+n0LNEPIL/X9QX46fSFcym6Q6pspv+qpvZ
K9ZaO45fWdpre2c1LvUHudzu94FUw+y0lFqSlCAiFWnQODaR4UyA0FKf/9UeJ6A4dqGHqt6Xn6HH
dpM+HXzkuXtLy3vcj9a4NLL1G3RbYVg2eahsUIrOM/gff7DbSel9I/Rn3ZB2H9m5HWlWJwDqBSwz
JiSIv22a5rSoveBLeiLImg4qPaKFaxHcVhOBgBMU4xlI5nfKTV5YP76oVRTE39DlgEfvs1r0hSwB
Hc7BZLSTcpmID8QqcSfAZ6Jd04a929T1TEdQlFmanOTefbJjHvu3JysEgEZUqwHOQDJcWfw86sbq
0Efr4Jomq8euNtuQMf6S6RgdKc0JL2uB0IyInh/mipZwnFXADWCgr5LXk7+cD/OqZwZvMZ7a8NKt
Tej2/vt0NqF28CnMdRLm8rwvQVvcfrWUSVstRPW5/48k1MzhXSc/vqyAJkZZpJBp0Z9JNovHpcmA
3JOmtoJZnHXOu6DJyK5UsTkc33cWcgeJqQeSq69AZ4O7x2dtWXIvuoXQKSBH4xU5sT/9OtEYLgnh
i1ofuYNAFXv7xNBumPGomQkccqOaL3HO1bLMGvI/oZO9aFXzEwpe5YCwXGK9heqXacF4RfKnvzda
IoYgGML4IF0vr0t/COt33ZCess3P9FEVc0rJEnaO/6FgailH4ox+iG+ojwxCS40dcy8aNXgOSIaj
vRGUmscGFLxIKXgyNQiMFk1b17IoRqRUH6BUQVwuzWQZ5CHX68HE0ik+DVX1l0tEVSvpxvzYtJi+
TtJRIobACwa0O1IVOnqKsLlO/DAtjFZajgO7emiobLM/2spzipu9L8Db53AHR+zNg2fZWEGXB8t8
2ICQ34j827G/aMd88Wu0BBmiXarus1aaJVQJrt55wdgWSbH/Fs1TBzqvdk/Z+cP3VUNWJB6hq6+S
zmJ41mNSAxS0ImsuCdOlUansASCheyw1RZk5pEg0c9jgrmRFtS+lj5J8ypl6FP3wMAgo6Ah7qE/H
3zIfvcryDa3ykDIyM+Q8XpOSOU7tv88f1MJI4GAlf/+eKtx6LhV3tHw5MCJI2gyhSo6qXFmODHIt
KyVCbkvGNKNAJzTBPrLWbPKcI4NSJh0w48PnnTHKhztp1ul+0V6MhCirCaWqqpwmnfTXvtzJ5x3V
u0KJHTtA3ton7pOwPjXy6wcQZVmi4wHMAo48fspGE+koayfkhXYvV+KLXkVtWncHIXuvx3fDewkJ
tluWW86GzXLbYAdddtR8KjUf/vXkw5x5Z1YGo2UEon6WdRX2VWewOcbvm8WWgalc+vYryd7T4you
ywHon85ZjHn3sChldWQgW1RjORO4evnt5DtydueEUmsVceQ/LFFUZViUcCB+SwGMYj/3X3hmOy9m
qzAxQCmJt0aZjat308TnCcdsm9GI7TPpYOhqZHU7t1yVuYhRs7FAxNggfp14UQvF0K+XkHDdsyIb
DuDG/VLFgDH8r86rfV6tr5q1PJs8CfjWrRjb/weTJQonSzLYF2CwbxpHHXTwv5kaTdWaJgtOz6OY
2O9pTb6Sv6FjJIZGMpewoNHg3ukaDJ//xAHQ59vpdO0/4WK9vJTSG5z2qnK489KMKuiGdop6o4JV
BvDaeSFM/Dw+EXQwAIpx1RfcGkZFtIR6K25Fhkf6kj8Xvl5YTa49Hp8h2AuyOOMXZ37w+Y9Aoqvb
P1RW2O+ksAOMXlb2fDLjTY9U/LByIN5NWqMSvdYWjugcr/b8tESUzhJ0oh98pbjJjNoAni44vN5k
OQxGziISWlruolJVVMsmMn+i2kxZglpmjx6cIuIsFofPiyFjWDnFyZZoHUCJ5hogUdtOHBWZsBxv
aEAcM/FV0rtMn9mnWQJD+6Ru6MvzHeLTbR7D58Ogr7MoVtch2RuAeKGvnVUuDeLV9yZ6BqCp1Xm9
RMgu00PQRktsq7xwFtn+C153g1hX7biMTnRcWUfK66amYCGpkbc8X4VAb3QGhtTN/31/9h8wiez2
+1LqXDCG8NbW+FBcTZSbNFPLvKexzziuhxc75bkt3UfPrJ6StKR9cvGfIXoz83uT6cljBI4hnq7h
p6LSUGEc5exS+xd5nFCyzeEFzxAJEsFD//nkkp7iFRN3aiyIWEZINNqL5NYA2Ru8BW/LiIfGkfA4
KrMhoo1Q9ag9uRmikhjUMvfZpZBLc9qI2N7qD4sAbBgECrEga9+Ky8MW9McUUNAPBykW1N5dkPyU
EjaaZAsIuXm6/9/0f2vqspH/82rJeAfc6+5/66kvdW0l43rrIz6lrqwePnR5aKuTzbKjnAl/dpqZ
4Sq4XgRid2mUg/9+NG7ToHUf9QE2rwnO+GnX1viU17td1eykt4KQmJLpT8+9idLbe2X4XS+AQ9UK
49a2hBtCQwi5kgOcoPJdgR4d14IGBRGYrVjSF6N6FS/zkE1hA7ji1D85utmVOhui386ABr+I7FBz
WC2Ki9rfOQOTBzjKi3qtzSrnVzxFw6wO1W+jjVlDDy/i5spuZWWqO7z13YKgGEjfAL19QAdwLhlS
sCC6VLI/lvVdIsHC/DfNH9yHzAttjBSw9HmO/fxoqPS7RXNYNRyCZaBGWu4BoTHA5yO3q4UgxQbI
TYeWAlpzGlHvgqLDd5NNLctP3I/Tn6+0U5vCzrwPod1nmqrQLIt1k2DjLQaGh6ODf0uKhMVGgpPd
tQymBLMC8nauFDeX0wn4TL5udv1PE/wB34qWHGRkbNtCDgaJDvLydw5NmyYdye/z2rui0z6lZxsq
DSYJJBhgt4KvLgAQ7HqDfqljhvlu3EzjPQxCAs4qEe20K8l+c7UvFMa1pKdOPvGDLg204Moidr0J
kIj/JnYjl77Djm6iO832zp8oIdjPk65Ks+HF89vGo0GEJ2Ze3lrm6rXCDTALxJR0E8XovgT+frqt
IsK/3Pp5WkxBuK747rZJHWlpijHsHM0lsn5SoNoUen63sZyJL2WTDk6oYpvM+NpgHQP74lbZ5oZb
0ib4tljA6jPZyDzxXMcA4xvLCSbOO9PfpshIBbaeeHz+nqwOamNNE3zZd9lWM7TUjrRo9XtFg2AY
vKYn6hC/FwouxBPLfPvs+Q9SL6FGA8fyhHy+0KfNVs2uEU0lyEBl0BErQBrJr6sF0BVXZivf9jog
vfuP2mE5j0HTtc5tP9ePxJTJvZPqKS/Go+qWTyR5wOmr4nfboGkW46P/2mWjskko0Ul9AaPs4UtS
HsimhcFgmEuJIr0gxWSbvdm04yUqeg249X+rOB+6M9962KU+WFKpNh81dGR3bQdZ/EJYB/WpcTMx
0WbR7n331PaJvSksWkaVPzPJoCEIMqHQVGkFkHhgpbZ8QP8YUV/8etZtRYjN8EBr0+oVugrPO1Ey
0Syl5FXE72ysvcXIdGNja9hHSWeQPGlL6Ufw2VnptBpDpQgobVju9oFpCAYorQ6Hj+anKAjKcCQ6
CeuAw3klGR1E9PZ3Y8gX8o8wPN110UYRcUEAj+FKw2WxucVZ59hSrLFCdWOyfYC2wUqBrrZZFTBd
HZzNGxxsUqh/m3IAeLkXxwZ46Vjx4eXYBt4H7jAWssfvUrMCpQnslmQYKHrWb+su12RY7Zmj4fPW
5VsjhQ89BrwLImeMUSaveG6xwlgR6PI7tGzeZNPkRL1NpWutlKuOi1yL96CtZGCxxjMV4Pb0depa
q6zCarLJTbDTBT/ecGUzPXATh4PysWIior2IC6A54vxXsK+DYoArPyeaAq7x4Vv4mOQphoCWQKdp
F2hhfm0K8jkG/8/2vxY8Q2KTePoOIlozDYmogeQRHc6yMJYwNxpgKuErNLmLRJJ2mDEOy7pFI3MT
kHIUAG+10RiO1iyk4+KlBV5jQ7lt4LIHEkXDy3VfphLf2FbadHRtFc1EZ8f95jjL5BVmUjOboUEQ
3Z6v6SmGP1kgPuhYWett9+8intiTOJP4XeOA47ZDhRfqzNedVM/i6dymOMrsVl6Yo49jU0aRZXIP
Uat3j44MVyp19aT5Un1ZwiFIwk1Vr6eY7bHajTkY3tS6FwYzCGvT8F3nQKc+2c4rstx7IdPvf2Oh
HWt3oiRM7BxaXF+D/Xp1S3vJdXA2h5JrVLKz2B70c6et6vInEz3CX7mGqNEx3XjAZB4+2lUjmcnX
1UvBDZMVi28bseP/62YwOU80aLjnBAu+QIyrJBG9YaKHMt83JHjuhkOoHL+ZRxc5FeoyPtVR7EsL
zY+ya4xqtExxgJgsA5BG6lVpDFZkjTf+XlocwTGlBc4gDWllEgafh3oilDd4EjvBEM54HUS5JBBo
Gf++wPwj6bPX2dSNdbTqdFD0cLXLA+vkA0JOpKFrxpoJnuykps2C8X6mylMx8yeclEPNIhZCvayN
+RjbFnuRjLdEmgLSZ+GyI6yhHPgUrCzfCOPedBUQdUMExtFGmu0gTEv9EzIv/dV957HRpx5aGSxE
r0HSyXaDIxqXTNPYsVnUGHWNSx7Q2xO7N7gL1Q35dWssA/0WC+s8hJv2oy4yUnXfDMEub7ma7kIo
UvNIcbqvQOBYCIF6lcHrULmP00flIt5fN4iQo+rhOCMr7DEZvp8sk0LvUBNIc7Uh3LvLRLto3eWI
xPho3xI0ZHgiG5bAuQCN8YLLC5RaNxcBQQrNMsJ7/Y//ynSxVg2IRngArIutfv18ywUT6EKFLap3
202abf20dGF7FK622yWJs/3uvkkrU82kWXFtpYCNnVYx+29iuBpt7seFMnJQ1F/cg/1kjZO9YfCr
TZiVdLUaZqqX1S39d3s6cEgQlNJ9kBgUxSwLfbCfNnMhNm6BRhPshJbBON2aGZxYj+9FacoAaqib
YzvSWFjV55uqeBa1GQAZjDSImQG2L5jXwJrG6Vfuch/ZvNNs0U2oLpRauv2Zfox29J2oyjMlhJCR
uHkmsbubcYNawh+o/0+Krr+LWFlMMlEHymPb4L+s6bIAj3oIzQt6Na27m2ynR5q1FArOVhsIpeDi
pyOk29yhSxxPHtlHqDUUyJ+ta5RG2i68yZTqyEfW+ZPxf5fvmV0enBdRX7DJJBdULEs7x5WDgLqp
ar5CUKBPkms7PKTP2DOfOlv6rTj2+o27svAM4cw7/1QlBX4PFTMv5flsyJVZphAJVeQozuVzk86W
osXszNiAjV38M5K06nGXwvFLSyaLkRo9WSXy384kHy1HzTCq5DU8Z4ZTdn1uGyJ68C0BbgdOD13+
KAgUYZq2/+F98uiYodCf5QP8Heab5IyD1xCi7dVUH6mKWZjClTqWEprLK/afeFV3i3DO5OkFgDdj
xZTB2LqYW2BO1Vwg8e4VfMY86ou/DaZVwurPLA8q6x5iNigRcuoSF9qUMK8QUjRGEYQhnHyIbvJM
G5i3BEA0H48fDai8FsMidt5hjJGkGgL2tZpzgxwuJk28iVNG5I5Nqa+22ofaXJLEY69b5uK9la7A
8TXJHOm1MOvd94Ny4STGdj+dosxYna6LGssdvc2a3i+jLKqZQN6FhK+i5zpzDzmrq4oxRISPwjgJ
mmTCkANZloCsa9T29qt4TOk8QB7ECzpa/HnzZMgP8HGJXCBUA6bQZx5FLpPR7/H7mqOAc7yF6pEd
NQiSMSZsGjZ13NOQcrmhrO35zVF+mw7GhMvmMNq19HIGP2coFYh3vYGg2oxIcSXPW+gxkIZXce8D
RqyYWVWbZ22S8nLthvBy12uVupzFIejsZMVsFGyePMquoQuPSYZTGBifWpeLsdcy1xa7SlO+VFeq
15N7HdAypVMs9V78EFPRh4GLadVqhJFNVB42Z2UAgY1sfYgbjuWOCpjJI3qy6XiHs7RIY63kDRtt
+38rYyAdjk3Po4QYrk7oRX8amVR2+etSCryZbldT9PRncGNHtOmdeh3VzoSUlzxXoj0pgIjWYkaY
DQ/37NcIaYBD9ju342eOgdcYI9GxMbGGizSWrIwXc32Npb0Za7WBzonGjtazlKPlLdxg3CIRn7bo
Ks40+Fff5tuHL61BukcS6Sva4Ve4RCh7NeEIGZLl5NWkw311emaoHC0DnCXvgpzKQqbHo8s4ZlEF
oh6+0nc4JF7bFhe1mMowR9EWH38bzn3XNBNRNzodILKt+UgJxPrIrFTkiUtCY5YgFWIx1EsE4/w0
z5YHh6J2dvJvDMpp7xfFwaBAk2PZKAn4AnZ8h0km5p3VFAj2CttM1nDp1hdAxjaaPx0moBPt93KR
ivc1oL/xi1eV2sBQlvq5ajqlfhd/hnBgTt9paj5HZx4jpxFwBwhCNReyk4HhytfSIsnFoGea/yuc
FKvVGhHU0zP53sgAYL93UxS4WEGgp6EnBiF2vIkxU17QUjljErB7N37VEjswUT1dKOLxwjxUdcXO
TwP2cnvAr2pyvc7H7JoAHfZzCagcP/YyJtniyi29fiFeohtdFNDSsShRmEB1uwNLV0/w2j7ekOlX
eJfmrnEK+LinZcCTWo2v8kfmO90Nmh1wqI2qpl4TTuhzeHqNg0wvl97EoG1tZQCyWqUGQg+zrQDq
Jq84dmBP8ImWi4nzlAz2YTgi/k21IVYL6hIXMoeCDJ/VS3Ue1omyFiPIWIMKPl6r0sHxfnSjmAJs
DpI5QRplNxawF1UxCdEt+oUNQ5FU6/s2T+ofOrMOUzD5fw5wW9AwE59B1tGo6ILOtslbiuCiqlJM
g4gUgYL/fafDMqZNGP111+fJUGixVK12hiNiY70GpvB8OpXGS41Jz2jV1/nZJ5E8eDGAtFoi71+0
ugv5lDKmYXB0pZLJSDRps91Od20kfSK8WMRbykFi2PU2L8OxkNl82Y8drfe9B05OudpfdmDTqe9U
+ZndtJXx1ItIsNSJItL9pJyFBN4rvPEo0KQ1eHmRN3kemgPDSFe902eJCY9WFXF5+P1c477BwDc8
GMMLlaO19TkyiVhoYD7TmSknVHQ6VN+z0akl4XcsQ5wsO0/lK1YDIx8BRqKxe4UEVR+MWCc9bsU3
QCDsr6cnaE2/e/HYqAvOFF+bTlZMalXlcobARlSCZ/0FvEjm6N3EHjjB0T2hVX76ppVMgIzZxnUu
iw/h41rJPsUM1CzMTAaquUQ9OrLUHlufkaApu2XoK7YJxLRQS2wW6J1+WatdQCgzALXxvSFytxrP
52fJS9vv1TSJKzJoNSVyOR0WTnsFPNh46JcheDwWcRPfY6EuhkKqL0sm4mjjWEOXWnbZYQ2p2Bg/
VbyKUgjdpONVHtbF6oyjkXi6F1pJtRMSWrgA8DKoxDSV6fUqgYr0i5IiQvUjdms56kxYP3T6DJjc
AslM2dhC+vmhNbCHsl7k4v4FypTYuf1bkz/Ksseu+KhRnb/RcoK6XAvsbAfFDajGkudU7dIa+7fb
9oDBK+MwVs6Q2nwgLSEkqlAjOraK8rXIT0v65g1HMYOcuWpkyD4KpW2O6q9c2qo4j85s54vXVf9l
gMgbyoJgI4pOf77PmXPR0ao2Zs2QHs1JVFdJC16Mu4IBYM+s0LcyQNSUlE9G44fs1S9ThOGe1L/j
tjF+wdxlgqy3rNehZLWTJqBFZEl6dyQVmuLhq7lKOFfmg6A5DQKbE93e9R9hfvddBrZoIX09lcP3
jmPXpiRY8PZuBEEZV57/htlYFjp3ByDrxkHMZfiugylNvE1D1HJLd/yz6Am5t81N77uLi0ocRyeK
HDYNeanuRnt++r4oFYjX2qcnJOs2ZcPxCNVlGSEFLC1GtEYTFDAl+ivkY45Ikfxou4M5JJVlW8K7
Jn0V6gmJoTLkSwCc5fxzkB0KbhMtNJi9TuOjaIjYVIYCV3uH9PRCbl8YKY14bJyyrV32q1AaL/vP
J7N3CPuRmYBkrHncZu+yDYxB4lH1ApsXNJCs0oboHQFzABCA6hUdvuFgmHv0QE0PNKMKfDW+ktKX
13gKrrmL4gfTKwqzb2ibKQ0Qk+0uFdlAUlKyXuycstGIIzPU0iF+TC5KRx68PykzwaSnctDzwGST
AZB+4dt2rOSNnesIWISFD95sajVp2+r3ectDGxPLokIeRLniYep8iN8aQMBgXyaP+J5WwRBjA3Vw
QAEaqIIfy4HGaeCUGtipywSgNIgmGuZWOBamqddw4hWvTjUqFe5GeV2GfnZ+mcfes9u/66+5P8nD
FW9k5vW93Nj78YxG1ubXD7t98uz1ILcSBKJlXWmJULB5eMg8dtkTKEzTQegJuxl0RUFuGgtdxNyN
8w3fvTblrKyDgzBLKY7/gREjIA7lapvVf7Avlsl+hkWJI0Z/jCY9RLEHb7vFRJLf82gS0TJUrfF4
EwWCFgpYnkF+bjNVMKd6OEZSmdaXG8BO0rmlR5akTbirgpLolSDamCldIdPTQdZt6QaA5dXbWDnK
pvAwiux62QJ/pVnlDPAWA+AwDQtLS4f+vnpv7lxLyzKM+vdKvbKwARzgsV+9NyU8bVx1YrHqACsf
yI/7liiGdN1HItUXAYLwyPtWrJkb51/3J+JfWV9DsdZAHwH8WN0HtoVOXUXHpLqvhRFxaUSRToWI
U/frraZ7WyzgDCQuPSwp2JG38I4ehjOB2FjhrtYEIy9Qq2tcP2eriIMUZPNIgZ4WSuezchl6lCIg
IAAWwMFZ8W3C/uwp6/+EdZ7DIOtesAABTfgUgAEJ91GPf3zBwfGyK67kK9ODsdUlKvhdHhpF1UIN
2E/3koMXIXsWe3R+XHeL4/zXSH8IMF6LT5xxi0i8P+ijRBEOf+/F56FqniT3XIDJYtmedtc4QG7Y
kC9+bvylEA1qEASKmBmU5kOUexrmE6HlgC9OSTTQNTDxBts41ZzUj9xG9G629Re/NyHEuXZapbaP
ef7C2GLXxnzQPpMpJTVcJs3mnmzR3dz9C4a5+Dfk5IczfJNJlz9WveedEfJhHwkqgvfbaBRFW+Sh
ZWCBeoNsykjGpo416bvDN6uQutKbn23TFhoofO2uiLR3YWa0D02YpwRrW0QpXAsNcKFkbfSaRTZe
TCzukaEHLu2jFDCiKAoIwa64JhDrXrNDxUSYMTmxX/ccIzvT3cDvZlvhJxeOdYzn4ashdWFeJfI7
uZCMzdfYs5zUC73a2asgyhvrcj1L4H6YiD5SZ/xpAKmcONOZyluwhVVtoG7daQxI0nnzUDOBVVWR
97bAX6MUG4OVuHN/Nn5r2UYLU5X9h7rjkV2DCqsCEp5ui59rvRoiKcvPHi3+ZUTisxtN6mplRzG+
BAxgnNaAJv29KqT54DsgT6jbepYlzUr8Co0MpF2dlfCCI8nXoIK1xmE/EpnWpoHIVepRJTXBEqAp
vhqVQxheqxlA8571Eg8hinfupMIaHPJcD7B+OtUz2JjIIBZF1nXuINvAR0Ph9tM2odoNwdkRT8lk
fMQfmhp47/9RX2+qAm6oH92JGZrDtdVHS4EH2kyDu6kJ/YCZOEYd9pbsV5es5FGEbpCZ8KsahPiH
nSvKOvM8ojq36Dio5Z8rOjrmiMdDubXqR41qpknR8m0GJjAfTuGhi8Uscwbwv1piycrir+d5nM/F
ftFQ9cIZkPbeRYAm0hIA3vd0AEkYwujlg0dslszM6LvRHSarHyAxuQJZJJstaAgQ2guzBGL4UWth
q1XiIMUQvqivFnwSL+jdPQfMUMXsz1VU9jQBTYR+Y0SpP9vf8dvRB+gzAPmrxtH81AQq2OGFb5Km
S7BmcBZsTMD0onkdoKlXK8ddpk2AD5dh2UVY0WijoHIolBloLWXbvZDAiOk1KhdcrF/bR6ex/Gz0
jAKl/e1IHMIpS2yCrsT4u6NSuB2ivJ6Hus5YhU3ec0/vSvv72oZ/ODHWZ3Ga0KlDEoynx/53lWZe
to+VxQCjjh+3TSf6tv2B7Tc+Jbcl5TrbygOLkN174JrnvxcITTecmvV3eyfaYMwf0zD8UKWjDBdM
k/gvKV4+xZuQxSH1hurf4KlKzLl6drGI6CuVik8rQg1uKaxcdNkYJSc2wbHkLBBePtNO9wXUCQkm
t9XJSIsdQpt0O7s4hNnLqpT1uU+htCtQr2Z+fCW6b+O68P0Kx+O4NGJal97zm8XJVTmWXX1PY5/Z
r7gE9JZD4XbvbLNl0HB7npmBkrtJ5xA+MZgbHyke4s2TC2QB95f7UdrQPa0hA9m4PqMOzqjr3dlL
1Wdrlw+1CbV7Bqpf8oKc5FIygpFRqmaN0rmVUYhW0+3cTAsWqGDnLlHTXTBQISjU29DLesntRZPF
O7GxXSgrSwJJiVki9H5DIK2f/rQKhnr+KMrhmJQQajCzujdyt6o7qTrbiWSJbOEO68wy9wB6MU/a
w46SrL1LVsVScq8E8jQ0aBklZd/yBo1Uiu+p6DIXXJEjf/ROAxOoxrtMuapF+lat3NcgaiAszwe8
oAsRJJJBDcuFyquRaDrZJLy8WxY1ppryefF8DwlbWc0/ZhMrdcZKaQvaehrz06DKQ0nv+3f1AbZq
o+M3JiJ+6idkrhDG5HpQKR3BO58fivWhBkLa084MsLgXbeP8kjz2VfjOzWaqkRsQQi+kpGNooS0e
KJ8gwWqh46PjHNv3RtrdeRy1jl3rtiz6KMS2kvPK5Hw6rd2NCLJAj/gFrzq55mXmzKhbJqDA0s4t
9FlCiq4S/aDshQPYXuG8677ObzDfLF4H4OxqKVgD0HgopOnaXbdcP60Nf6uzZQqOcmN2cySZp8Vu
8hDFV1kwOWVcFBDUb4vkWyPdz/Ht5rRYTvQbCuXX/bSY0gcu6bAtzWIQP44wcTV+pKqZlz9FnaSl
G/6QM0AoUCBElLIyuQgX+ZAbpTPhDLj/e6YJ21LLWKABkCYYh4nfcMFbvoHF/VwKJI36VswpiJ/r
DsOeH0ReEq7ufQbQHvaFeerhWoXuq4NSPcAhgqsIzLWBYj/0T1Hx8vecVnQ2NVELxe0Zi0vf0knG
0XVQszQ1lGYyTOgBGo5BNxe16btyYyxdWj3dgyYhib6pGFhQ3kHdjviFwQ7BwkQ6lPFSRWH6vsQE
oAVNtqhioM2IFnj3edxzQuAKRk/W/SQKUYqwDstFPtY5ou1blMYyGhm23c9ZcPt9+f2DaZ0z9+wS
5yN155zR46B/pOZn3pkQQh6RfgD2BEEMVQ2E8WieelVvwcbLbimyQQNBJgermXMPaRuuhWoXuzaJ
33A2Sjs5Nw3hyuKA4MV3KCpNUuxY9ruGOwdOXXNy97o2HaTBl1hJRzHMggzlae7AqsZPEs/hN2rL
G9zqazDvk4HUjZTOSd2Ue7vzAf0CsVCr2oHrtqsgAWTLXTm3ptNu+2CWy0y+lVVud6Qp6XvrXdH4
ihb0UObFkpZkW4IVwpyWpkuI/EtG5EfUYbVTUeaH+jt1R9QfuocbK+cjJo79gPnpKE1ib0DyqkIi
ddQrgwHGe/IIJJFo3H6o7RE1X5LKH02zB8yx3DNjOEI340Q521dso83y49a+w+W86ytwJ2zT4Hdd
28QaPj3iP5nDMrN4iczixAyxIN5Re5EeC1fTw8rk9Dctv81okTEodlETz9Tju4LyMkQedFiS0wGt
E/uMQWtDJUcDVVO7vrECWtBUJTx7lFI5UQZKU6B4QEKMB4AGUyUn+qLETuMRXO5jbpAqmIvnUN7F
8iDQHp5oeBEVdlR7Fqtw+IaEeS1brlEJX3Ovpek617BEqbvoIIDeU5Fl93gldZUKysMNZOKRtY30
iWSNz3t7TgWwrJBSx7p20vcZ9FMc4MO8i+cLgoHpi+5nzJxcBhIdvMc4X3C7i43OV7Hd+dMiilpQ
lbs/CB/1LNn4vT+ulpsQvFts/b0xdLNgKXatxh/NXiaTjm6jwo4zUs9bEE4IdgY/Krc0sFKk1k9n
711oRXi7KYOcxcbb/yQ//PuSKWYknENe6/PxkmIu1kv9C11kAGm4agWZWC3wERfzEscHTUfBh22m
LMqzX7WnmxX6fOoLUY9501OKHTUyAOzSbDV+C5GmFN9NJTooLpxPgILBCH5GYqzuKWH+BLoL34Eg
qerHwJ+bi+Lc5SseX4vBdOPB5r4gjceD18ijwrvnmC6we6/enYdjLJg84D5Hg2i+bsxvKmKf1dUv
ZJH4dyzwwYlG/Rfqyv1jvQJD7mO0C3NNS06HaBIpcx0TZ7ntpcAcGnESJjgatGmil4/8IFRLkJM7
QhiPd2o9C2M15/BzMdK6ELS+l1xMUc+Cddo3//QBSN1sZLzL4gbn1EL3K7P5mJWFqQYAZ6pBuNk3
ob2euCgyRFXJa0dLtHR3wA98uYqXptBxHksxzA3GVXTZCUXRlwK6lUSJRqc7WdRMVhatpgL3Nuac
verNAaRcpvHAAG764qZP1zUUHl1wCShtRZ8WsqiCJ8nfoqozqN+DS51mvxbM9uLVBa3GjHToiGO5
WpEBbM6LUh62c73GYbDfNf3/oglzqjhxV5BPz2oLKValU1M7pXt+4ClF00Pvm5FgIN/3nXiWkpkR
LFXCcKlW5DRofZZFaB5a2DIfCh8p1objkolH4njfzgtV+JCURaiMgxpWJvXRzKAVjFmnLIsvVIcI
bBX/UO7B0GPFXyuatwnMSDP2RmqZk4YQhfT7mC2+r91LyntOh3jJDPUpDwTSxLfNbk21YY842xUl
9UWvra6vpa0zoICYooU7maDnKIzPtgrulgy6BKKKJx52PvjVPoGKIeD6Fqzjoj86SE2vYJUQBL9I
6BFdk9rAE+9FrFvI0c/G+P7FzWF4xl0u52nnM5KPacnN8YlyLQJdkc0b83m0K93TYWc7wLR9XWTm
tsGSZ+evoEBwOhQ24uILbH9TkxfgFUL5szvLTFIEcNa0M2FrMhba0xFYq0AnbpnC55Vt8e2MokOO
giJIX2Vcrm6nIywIURl/6v1ArwiD7fKnJlcmlED2205QScSg+mk5+f9qhxig6tc59Yo8TjMqynx7
giMjasYPu0yMrN0RplzQ4IoddOwdQkdUK/G4fvPleCWZYxMdTgL6XQCnJ8sz5b8tzBwWtsMzPEn6
nNd1ZCZ7tkV+RJwpUuJ9nwLOn/aGsRzXvAZyZRxE6QNuYbCP+NoZ7Wl397Fua4+0sZKGqKn39bV+
sSsLrJoubmtW+aqnblh6Flo7EA5QeVefArFRzWluTsFI5wFUYi8eyl1tR7u5hy0CvxQ3oyXX8ftq
miSYD0+E+YvUfYO3udOLIMqWPvTinzlFNEXiKIs6zB8LI+uAOTdS8D6tt22+e+YmUMLk9agXw84T
FY0WMtReYYZw555BLVbsT3UVJyP2g5m5JevIsotcgGeg9bSWYotpjrB4H2CJBFrEZIkXsjRrjNwF
tALdbNTtCGhQK3R2FLFfiDLFl4LE2ROEMsuHSrEecZF076Cmd3SaxOgYrOxHQ4bRgP4lzvTQdjP5
Yjcw2X70mtcZcR0ueH36IcjmcqUKbDBfpcWPVhO65GCwDMYpRPfJZyA186J5XioflqxSzMR4Tf+a
h4ejmh1fx9RRZKIs0Bpk84dEr8xsJjbY5uP/RvMx6ghQ+/HNDYQrjiCbzkO1SQYm7dzmTH0wWxdr
YmE7b16USTGMSvh1vLZa7ZAZLsZ0ji92x0vA5EAyQVof+Pkkt7Gkj/F1SsbkIE+DPLAP/48kJ8IB
rppYvhbfgWLaR/3R0xtzrmTUX5ANmmoM/h22P1tUHOaD86f8PsoSENb46zy7Qkyh9myysPf2XmpJ
J0Fgr9PBpzJdWMxFSc3wujHsgm3+Bm2hcDC6YBfk9v/5h8ZI8tgPKe+s+7PC7iGDi1JWrxu8Jpyb
7/7yphNqrXpeUJvhPdSRWfHJTwNu1yc944cnN+J5IiCNiubEwF++VTSfC27+Qhkxrgwxge0OH/pc
K/lFNEDWU2ZpQQf/BiPGA+gZk/y8GwCYNvR68L8vztRLuFSNz+QtWlIJj8AJN6KvRgy8MxNvHxfe
k3OGLPoqGTshq72AWawDi8x/X+r4MOT6765Hym+tiTxJe/kEbpSuQ2uD2UpXRIY/fyPrNgiaz7Mg
uLDONAbyccG/iDcp0w8pqMFpo27BQ3793i7WgRMdKJLUpA3FYtYYvq0jzS+I3qNz0G853H04T9Iq
Z2IIOaex2a2Dxe5aXoO0fX+dieFxV2ujKmraVKeZS41un7v6uoAEMEPdpASjLsgwwJJhOMZg/Hc8
hP+BrULnKiOcGa+LrMzjwaQZrMfpWnig6xdu9/sI0/8pkROrV+XTGOVdDf8/Fi2d1yKbop3RNBL5
VNvmUx2xUglQLhwqoPwUOFnC6qWEGmfEOEBvC8SkG0YiO/Oz0YGLKIbNTGkyd4C2lB4EOuM7foE4
yzUmHnCKEoUFyJEvJOVMQGqgSuOsPfrrbARV0gAWWhRufle+Q3kT/5mByH+ZBon1jCNraMxpQYoR
q+phNcMisnXNtFbCIfR5xfCVwFvYqbHOLfj2SO6FoZ3AFe1IaXL35vNJ0RQHQtf7gc/bycEWId6x
dr/3yKWMJuQc7mBkPuPTEy/4zaXFYTBoeCmKN8kILr5/cZwG6IeqBx4olra8xd0TCOd8olsCfdUD
K5/P8xcRjOk/3bHHl2u8MO7UfqJcb9BLIY41o7ZyZWbVm4DUQtQW8w/mpzNwvRY5mcdz3usbCm1N
1lfXgLvYMkv+20TrmtXuADTbS18qtpAM33h5hlisRu8D3ok4VjG/2uMcvL2mez92YFC/ju6Vazwj
xcywIvQmg0+HiOVNLFr71UQT8Br66IzkfUlFPAhuNCtkc3Vbxy0f90HQPhze6bBSzb3SbBXI/BQj
xIEk6Nv025H6EQu+eczTyLNHT/lSUhx/IPWeQ9DhGGydqOzF9Tcaadb4ca5BZBoT5fbS3QNXgHfK
7AyQR8QEYgcnqNZsKF/veyAMmP5kCPfahZ1NaC239gsq6tXI/JYGyXuuf6bBg2HfwNz+jQluqHth
C27fXJ+bJyEq4EzQaXquipE1PFa9IgOQy1e6xyoz5h+JjIpQfR6h/8f+UX5MqvShQV1/vRqXszxV
oPQ11usOZIKLxaJbBRhKZOl2GK/tEIq/SBh/i3DCcFOVCvOZqtg4BD0iQX206PGkPKRZB4QOZlEu
uMM70It9dpJDedQyRfA99rPu9k32A7/EfECO90h73s7XWcVLK3ETmNAHgvXgAEMAOjxGPo0Evg5n
4bEpUyrMhzZp2pQAom2WpBXowiAyB8BiFqHX0tXxZNFTJ0H2JVHW6Nmps+O2PiaRpkeY6k43QMeY
Vv77B9uk/UMX82Ee2F79ou7v/TNp6En2Q86LUgJaodW+6uF302pRY1EkC19+MGfN2FgpMjQyt6b6
9ao91fJzEOCvu+1b0mEiGg6eRbFTt5aMAGjEr72hH6UGDHXi+wobil8Cll3UA8Dy1IX1r9rbpYvR
f5wuzz0IQMU/gxzsIbNc1pgecG78LkMBvXrO+okNo7pHhRY/aWBqn2n0TtvKL9ImSqb2EhWOD5+2
mqG/DlVGpK347t0NGAO8EzpsUrxG6DBmxSezgiYcmuKIZmSTbK4BMG1hsvtnkoY7ifg800iS1hSZ
Gr2bHtQ0xUTogTiXUPBbtJJ8KT3teOcw2rXRPCVTPN+qG8STUR72KFQ9O9A/rO3wmosuBFt0oJyp
t9NYqcs5afd3YuMfIfHBrf63NDBveyx6TiVi/t0X+jZORZMxqq169hWfnjWGLoiiOsmk++wVSFeW
OvmFCI0ZiNh4lcVIlwJM5L209ltrt2SEkNzYPiw2tBYqcNW07noBx11BL0mS91iSqkUruJdi5aVy
33jalFTqgXjGSvdPYl/Z77P5Lag2PCk5p+IKzknX3pReVmq1N/6RMRwuiTyDtFvFMiNUawljaPyJ
wDMdCId0B/LzGW6CTGF+q7+GqrttrIZmzLJCdGuZmpxsw6RMmw9yP0gSt/WiCbopGpfzKTK/jphV
iwKY3REFMoebKyudhJUfX2RbWqzwfImK+wEjXPoFA3abMXemEeZBUQP4hNhTKIgGvxC55L9k5fAT
cZUzueBoEWPye8DAir6m1ulVO2REVSMsPJK+Jx2ejl3QYvDN1JOL4M/SkVHCm63rSm/ERpFBrZsj
JeL8/pdsYmvD76JFNV5HBJippx9mbtfMRNsYEz4wPey+giancuMOS7tiNj5i06e/0OtgvE5bPn+2
b4qj7joK0GMAjGNyK/yhzEefty/H78PEd+qfTjzAaoS+8UOYU2yOeCdi6bZ/+2uK/R2HKEWCi+fD
+8ilZFGrapFLqD9eef4LhwPGLSRgZ9mlMU9LrdAKi9NIbijZBKrQkCROiqR5k2ssmidmo2MBg3NY
wkUhm+kosA/Kk0K4DjkL5Syk+CjtTbdaZ2O35uFhjzFJ6aqOXnyWsNhu4S63aFzvOz3pDr9q6ogD
tft0Wdi+b954e1wyx+IZPybJQPzKrrmsspOo6Axftg2UCi8z3uzS1yh3pW3kwgJLh7Doi5Y2tT3t
zRdfP5kBsVUBJGZzTJPKiDjazMyTds2+Y7kdj8muQlR55I1w1QcDEGYWG1t3aUHzGfd1YgdsYWbU
UNgZmEwD0rG1SyyN7xq0YblxSOhGBrkrnSkiXzLkkC5C4pIiHs9uiCaRELNRcupmyLFIAToTk9/B
A5NonKvjbWaGvptFyiq0w6yQcl7toqkQRUpeTxt1zT8nQy6V2v3XhVheEEX0tEfmRZpHpLEomVC1
Oo1JFd9nn4MVTolRcCQ2V8SWBoO34vK7HR7Mxa35s3Fjk9yOX7JVfzMSIexdhcX0CwBOA2ObCRce
i9N4iedZRO9BSKz/Qd5B6MAxV3xXxU34hrpGVj9tVh9d1lSIVa6PbdxlD0k5uZy56nccC6KVu5aT
AZYySt9AdRNNN64BnEHStD23vGwnDF0hCP3NHz4jY+vunANdmwwvoYTaXcgboh2TlEneRqLGbwSE
EJeGgNKJ5ESkS+5EgIkUrMwFOM8IJWOiBIjs+R3V+Qlo1K3k76mxIBbJXxcWnE/xs7ds98Jp6tmh
YzT+OfAit9xvUkZg+Txu/CeCHn2xqcVtUCjtIf9cWn/MoGM9Zq5m7/CNa9zePzWC2w2sc6FeQhPk
jWeIBhf0V0faf2Yq4w1BKzN/Qzml08qrdT0FnK8uwTWYn1uUj9lD/LGZJsReJEBAsXe1A8WwpCM5
sVp9dvsCQno1L+o8ICCvTkJCgJe0mt+iyjeDIDwH9YNT2Yf1RAGxiqGsf1OlwxSqOwbprWdGDiuf
N64XAe1BQbodJr3jLfAggJnElthCIW2Ec2RJ4VlnCAlPnWA5V0ify7dWeYII4aCXWy65ZTIuwQvL
r9pwB5EYplDiDXdMl2UYL/m1DYYds1pU6zZxNrQDqi56hMkPBmy3cMm3UiMQWw==
`protect end_protected
