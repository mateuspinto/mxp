`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
hVaDHmomWbdDgy68IRYiY7NLSI+2MmGz0QwJvjpYA5Hu0u4nEDd0zB+XJWm8svbWqJhbR1ZynsWN
zcXb5PNStnPiMChL5AYGRUi/h9KMp0b1UO6+8mBuiIOngmcRJcdyBNCHpKqHhh+LoC0gz68CBt5g
LhAutshvKzeTaCW4um8q5aGkgGuGPuh3Y+nHEuGRrLoOFGu2ZSvbaZ+nyz3zxDmIHzNmlpeASKJW
A8thiJ1xGH1TjB3DwPbx4kmcDRzQ+0n4SymCARCGkzyLQyjCS3ShdUcHBcTOxCZ+FQS0lwFJ6FMF
ArxsVTyaioBHLt/tzds0GSv06vW0DXcMT37wUBHfLUlrA0yYWgUr7O+vrOCU5HD4RGfE19nbeKj3
5x49u/VDQP1bgYKnFrgosldEdC0z60aJwSpa65NXFtn74nAxpiKomI8ccPcfV8oeogMse0VNXTUd
mc3sGm5gn+mtWcgB40oOibnP+bQqYiSobPxGdvVt6ShuCwvsYEWvJ8mr0zCuh93dmfRgFufknRqA
llx+EDUVRRRlRZ4gJHARoFq+f1PZVhezPyD2gZJlA6aSmy/VtTlA92abwMTqzULP5HuPn6+vjBuk
DPXuWm7CO2ia6sW5K9Uhk05QuUK1R0ATjjPE2p4QQoI4Z4Yo1HpxE4QfAmYg7sJY0DCTS/2OgiLr
s5EntttTGFKz7/dxLzKeKBBbPcqi61JUwyxMenjnq2e7pB5wmkqmvDNDk8K/qGtP8dx2UxSFjkWA
Tc+/la8eC4ss9iyOSmwVDr97kFPD4jDw0kCqmSwwRl/coyw09bdJDstokL0ZfmB1hOz8hiGg53Hh
+uUCcTu481v672eFVEaNAKsyvesDZiGNWtR9ThgMpFUe/2R6OiEgtmsiX6yPoxZTG0n8O+Q4YVWw
vHZE4hgT0IE8HHqbARD+mqkmxGnVLQk/IGyMgtKBc3DyI6lD/mugjR4N+0TbqA1KOs0+FawKSyb6
tyF/3jId1M457mZQDcU6gzxtSRzAFrM2LGyrlCcI3LZyMeGpe9HyogonWiNPwT6xZfAlWlKBtkD2
zIIMw/l297PLiltrIbr4TLrAJ66qtHVeaPlJVlREg18q2KscszHr8bdUSPjipAld8jMNaIj+KyZI
Cwb7HH33+hsFwZydawokqDr0MnJY4Y0s3BBmJwdOAXGKB98yYUkrm96f56A6gz6MhiHAdanX/3CM
Qrvv4YmjmHcQxdfpjkIK37f39Q3tG5UpYZeWn2AIc/dDY6XeHbNeUY4d+OV/C09XMOHgP6BwTPuc
ju+xOTP+JgtXQJL2wUy6bPRwRquIWljDK27D7hwmFnGhRe66P7Xg0xaWL1dWi8ZSQk3GwBgoOkmw
OC9uCpe68BV1wdvLM6yKbD8yxxA9CVpdV4MHF0MgM7mm96oiFUT1Mv/ZCi/GT2CaaW2lZEKybE2R
QmE6hP4JMl8b83UwRok3PniZgnJj9iV7oMyz1Zdm6pjZyzeMVbTL4bHnc4hOHNr+rF09tRT2Zr8z
bf6i6ju393ptvyB2YsAOrPV24GaKKUMS8zRQEpQe4mSTPy/3q66V/N5FgxI0pU7cQgJSGa8sprXr
XfYY4cBWlUUZaILIfWGEuyS+jtdnCouBK144cVVvcK/LTnGs4X1t93EKgKXEbbDY8KF0hFh2XOQn
J77dkV//fDGHVHfyhrBDz2zfdeU3jzC16xpchi33cMJ0g0J0Bj+g7P+oa91hFMymsUE6UNkMR4hz
PDbRD06yvq/6Egc3PKzu4On53T26FH43THNjm3JKeDG9g62DqgvyeB5joasJwcaSFq5yTls40zPg
Ojketx8NNb798AuoLte2D3sbljo7Jyf67GHlLkuuy14urUqXED1OTvf1L5jidWEOWK4d5d7FFApx
QMNRLgPQNnLOY7zzMjnlJpQcKlVrcoX+n/sSqzy0B2MZ+pEmemxbjvFa6SG5sPGgKQQdPhY/iqKB
xU2F7yryC2yBZ15I/Kx8N2VEE9xx0QY3JyrLvQaQuNx2t1IHwwA1PmnQqyASpLrsBJ1TLHhHfhN0
D8Z1BIEoTP5hKra/CB86kk38eZiC3IMbiA3zRb/F5BYX2MJfldTRx7soGkGeQfufVY69rQHs0R+1
NmeR2yzlmeV7Kb7tvdkFGYwJIw3N/KPMrKxo71WfaxswNYCm2N5Awe6Jjyv58ggEPngz8WxWyRli
ZXXTjSvM0K8Fjc/vVmMWrSn3nyo1MtcVh1e8O5IvOnDQGWtYxo38Bc0TeOcUaKlTkcAjsp6qiGPn
eDte4KH9pWP3SdlwMH9Mitp4aPKpPszSnyZ0Ji1lOt1joCFaQtbh+MAh7I5LE9xOPnOasZgiQ/Z2
V0qSs3c5150ehbNo+eHPzjYhH4YvQ7Jw/UsSuFsd6NgblsOauAY4PbPR3r685ocA60LHZ8gv17sO
CNoOBm0It6kVgofk3T+8Y1Ny6PUVyDfWINjdO5hth5QdHqi602BOI9IMHlQLbNzua6TqJq45yEbm
Sly5xRiJsBiwBACSUNT0qrp2c2WIxf3E8R7EMfagoSP685TQ9yN+1NYSrQQ3nTwRJUBnlhuLbdAg
9h2RKb4EzQWOmZ6EjRCQkNuWvrWF3h4rNAbTMAekNNkjx+/3O21Chagb0mnw/Cd0uCAR5fjr2N2V
GyK+44Z040+CAt+vgHg2eO62wEr3rLQ+TZfl9rxEObkkGezGHNe+T/mphzM/Qj1nxwDmUpGwKWCF
aRd9bYJRb164Scm61uxPCg5jqa2a/8RZYbmOW5h4G1xmO/p+Gkl21aKh5+o7vljgiyF7jUsUrMbH
pxAC+sTaVtulGwzoq9PvKtERzbLsEwKoJqHQ+ZQNdjQTqUmuEqYde3HYDres1FEMvIRt6RGwBPPx
kjyvq/t+9InpZtiit963i4FN0m+uxjkjitfF27Hz1g3uIRj/WLzouLPDa7fmCu8Ee8UzG6h0PPIs
feUb2TWmSb3qdSJrca63hFZaGaKMX53bxZKldhhDUryqI+DR7xUovlEAfyIjncgpioLbO58HigQO
mode+/4DwnGnRL17LGEdLNrIBZWQ1XZ9DZA294PypbcIGAW/B5wF1YgEdtuLNIEoZuuMgk1iF41l
72ZCNMEURZAuAdh/AIM4377hrL27z+dSux0YHp6wEZercTkR2hyccoDU0Eo2CLZICeeu6g7IJAVL
EF8Mpp2IMXNWtLYC21uPgz9aPBbOKqAw/N4BdU8SC36M204BxLYwP2CyQsgFF9BsAR1FbvTY/Nqk
riIAk7Ebk1zNbO1MwlX5PTl5L/gcPhYhlDN5f963IyZGhU2uxm6FgxeYWoMHaDEpI6G19tPpJgPN
2XNDnj/KuTlR6N3FTUixWKs1KCu2FS16dhgWd9Xse06Jo1nZ7ExVimBXZufEHXZAkQrJTfqCPjco
fqNpPxructl8qABDmR958zKLub0WayBGt88zyn9K9xfhpJdLUyLMFDnwrCWnXH3rbeUs9/oeI20X
14BeG/gxHs7NkKghqWSdaATcd3FdFIUsuGJavt3gXWNxRF+bnPLApGAaxOFhMN3MvfRfer9FnCVz
reCX5EeJAdNKHkpmwKc08C5k3lALMovn3M/0GrNBOGbjpY7C4FDa+2Icp6Y1XR6THxMG7geNpjju
/wx3ASxqn30rr3vG4g6o/Hh29M2B6UlArJ35IxIHa6oQRB4Ygz+b3vqvdplCLp1FEWOUx/fC5tvT
gH+qh9DDsPCYPS9X3p3QcUvlGjqrnq4MBR7nr44FcNt0TfVwUqsp3NVE1KibETKLWXyNdzLEuUSJ
/rT25LMEenUw8ir2nYK63xKOtbCnGsJ1A1Pa2r6MueFrvPEX4HG6bVX/GxEJFA562A/vVnvhgunO
A/y4nomZas2IFuR8Py2BAocw1yfze1rzzT8UeU+e8lihlcJefR2xwePFZDDBhLeXIlj1mmSnB1oo
zIxu+CgBT60+YQDwaHBN764wtgiA/DNgShpTkyaNu344Dtf+ZVzdQeUnWDsc8USP2W+r7YfywTVc
ebXuJfOIXsYTCnqWAzgLf9FaMMTKm///67w41BFlX88rEmJJMOiQhi4DCNn7ZsCb8DoLG+EdLdjT
lKAqjMm23/Z7fmdKI3z3WsToeTLmmhUyNLxqOgrwwCTdvKEjc9FeJfHZ0TCnrSBZAmdCJFO/21HV
I3ZeXXPM1A292xBFTtjUtkyXvfsElfxIqelTGc+u46UQe6cbsYDhK5dQ8mSS+wl69vtqMHQauYo6
CBSUjJF6iQ7fTZ5xg4B1mdUA8JF/rtzm5qP9Xoq3AYtExl/LUmyhZS4Tres9LDmrqLRz+S1J1iL5
u9a490XUZb6k1zd7Zec/XVMuK94UiIK/tmzszA5iB0QciA8TQnlP+NFfUc0XbMTEsd+vliYXPneT
Tm6A8nVj4TA95v+7atLG8blUhkA7LmxpesPuU9adFtjYHihGSb7QegoIP4hOv63w64z88vAy7QpW
CjDkjJjzm4MMZtpPhUBpsj486qTffa5NqYTjxeQZmsePCPH6IsUL/QiD45atqI1jfAR9R/rZeOLt
QXFpiXCTqMrVZzIS1RFRfzDa15OJJqZebE6d81r2CRCJCBPYQa9z72zMyPaDBEKRAeJrnq/lwKB8
cO/cVMnCJzor/ZWQRccOfzlH3KDUfaNJ5qXaul0X+oexP9d897g7zyK8q0MqSW7s003464Ehr7Lv
wOkcMsRMpKApyysVVYS46vN6FWgVok0cUVi3mQLokKNFyKFummIXNomiD1UqBcvCLztmfTgUCT36
ymRxYuyTasJEJITL9+5V3f9ny3XosMyOBVlnh+uts3AP2KJijIG/FvJEO+rYrJyQU7IbK/hXjSPE
OaB2N1UiG1V16jnwwYVbuANnDHXNSp00bn7EJnAnyZDaR7XtCn+AX03tGa7HzO24U/PBZ0hguKvg
IpoNE4TIfFYj3P6spJ+LYOROAnavibdeigruyQx5S4thwrDt9D5kXCPPLaC9djXFdCRUB1mYSxID
pRRa/tpkN5/8OUgHmH7czOTO84lu3hLSAkKfQCfEdWLSCccAZtC8Zv05TWlTCPfS+OA86mt8rEaC
5HYbfVT8rSVZNLXsjRuL0BxXmSc0pBptkugRaEad20b3uHEujPDLcqd9iOGIyIebaH75srZaavCt
TU0JMEUjBfHjxbkLsFqIqmd42lD/EkHjubd83WxuUj8cL42nwwGgBGMftHLAlo8aFS77QhpX8CL6
+mCzOOPlzYIEJQy7stOviqjaYosH72tbCy0oXPmadu9yzeDi2F5mgjbqTol5zIsCOGEp2S2oRaCT
JBK3ztN5Jmft+L7DKyErkNniyhXTgsF9R4nIBrUg1sD6vUrnxL3WBfqzkZ3EqnfjKv7haN8vjnsA
FaqVpYpDFEHPCYBkci6clyQP+nc6I3Xr45fLynyW7UZQXBDFDuyBOWg6c4tocSQ/Wb3luBBmAOE3
PwRnlM6iX42EbDWy6DUNSOLZtO5jPebibxYcesF9NvdPT0QgYYb5LI+FhZYbAAWL3LAIRsmrMkX8
qEYgo0njSCxS2bP/pMWMaCGr7gVIJtOSMuh7eT/RhQ3oRP4RAwEw1B1+FRV/4n/WmVti7uFNlT3B
WaN2k+sC7c7DGRlSoajRDP/dTEo3hda0BUB0mQxYYEZSbsH4lWiGqRx6M2H2SOmXPFoTMEVHNzcx
3OqJuu2C/BadoetPBaRRDu4T4RmJ2e9Tim5JYEdbW4ZEN2Hn4y9lq95WYnK304js2Fa3M2Vwt0MM
CGEpNVA9+8Yn+XCu6eINClNR1dUHSWFua4Z5spaySWlIL1oDHo/MsGGfS3acsHZhR4VmPGTGm7hz
UHQoKrLOsYYuV3mbY8J/9BTS7OsB+ETjCfzVBJfRpqsOiJeJxkMYUBdTf+JErfi1bYR8qw6Cp+lg
rOotGwLZ5amPjQA2y/zjgY1V5aes5eDDY/dygnJBKQtVzPaEI13saIqJ+RqiLNKBk84m4HmxwUpG
KTfmB3aXKd1xXl7utsEZsRTK2BhdPtTfOWQJcUJWnLXQDB3570Ba1Nmq5gFprmEkILqo6arWmzY7
S5PBikV/I64JIzXERv1I8iIV+NnZKNX1mAgYfLSWLV1d8bw8bO9M6m0bnIJQbjaLtwEZlaf+U0e2
K7rkvczzFNWcMa/BgcM0Kx9Bbal+j28umsNqfcJowLvZtjuhdlQPOhO+1t04OuVMi/Vxe2uGGaht
IMg5kX1Djv74zDKoFEHb4c/wblao3sBzv1Nbg6fYDkPbg3guTRWV5fou4R0CFg00EbLSAnndKDSX
0i3edaM76AeP/p7x7NqojiZ11Q9DB0x7wwOzfLIEg10rYGjR4hl4VFq+KycxIrZ2LS0OYsbbxhu/
CaKiXPPeY3yUH88Bh+HdnuJC2+KsvFqEdjYSXsF6d+JRMQ+wDG40URVzxBgVdg6Vl3FeWYnbvY3f
OOPnNOPnaQ9W/EfWqgKcYiQ/KMT9iLw6fxENgobzXxDZYLTl2a5tl7n0WCvkYqJ06RHwU8OfsE9L
o6mghntl0N54hdHOTFKPiKTdbUj/fB9IQt/++U3oa7pYy3HlTCpmkySYjf2BBbZrXWUOSDNncd5v
cood0yJru4EtC49LoYv7luOSKET9Bsk9vfDEF4+5rGr76Q093xTiWONpYRhHaPQyWkfWX/3SXclF
SxK/sD/TKsrxXaOYTnU6M3ygKQazjyAHa5hGIToMmSgdT27oaJ/SuTvMZp7AS641c4bPA6yr2veL
1Kd/Uvac5H8r62jMRwIc5FzWc+8YrXgifgowgnjoPAYQJZ4H270K4hMqdZ/BCDsV+NBNp34AmEUu
tgK4lqYLQg6SJSeV9sCS5/Nksow8hfrPLnQZgI0rH8rcO+dcrKh3caupxseYSPe7uVHd0Ah4cLdR
58LQ2xOb4NrDDyOlLEmHOdW/6bTldYjfl6C5ortPVoIiy6vwzHozNFRZG9y4iT4xbxGXwIQlNSPq
kNtV+KXkFHH4Wc+biWWu4M/AnacUgnoYGUiHpJGzjb1UV6IDMrLGeJ8ZAEBcMDQ04cRaOIKq2jSq
+EnBbfuqORlhPqCpk2ATlixiKRxVAiS7ffSYgVpPUUstaBlQND2HwZ6PlNeid9ZdSBr9pno8BZFo
nBAB87pN2FRnNA2WC8034oQ/Lg93/7GWtCSbpAfxu6nFFSt+G5E2LtBWw/5l8HXaCi8BaHvhxnK6
yR2VAJ0c0J9DYF5Y7FspIcwhWIEJIl4fLpvWuV3sh3nccqHaizdUz0awZuHeGauZPVzY2TKo6RTu
TcjVgQXjGSvi2ZQHarru4r42tLGRYKgYHC2VrsmJqqUjDDYHVJPxsG4ebBjvvjVfTKhi8f2E57Kk
8Fiw2gLCQO0KN39LViIApB3AqRlL2Mvd6/rmJEgW5WEkTNWv/l6GY9nFFaGmnA9MdBCZ5H5+Q0NY
3KUtUEiERZ7FKXs5CmbM9T1BnU7cI6ct3CpvEHjqijc2wE8jG1jQDRQMGW3pT1wBI+lzmp1DKaZf
/SEDBKqr/bPwL+4509HJ+0HfOUgIEhFumV+HcbNlXbCJAxqpNcvMRdqlWhJ/UySGs+E1tEcxb3H1
2QbUOmYTS1szlp6Opp0BoTg4Z7M6ufvVdJOznSfuzSPNsJ4wQO8EcxKceJhO8zT4BFcB/5WEIEGs
/1w751n/WhuH0T9u2t4N2j7CrtRxDTV6oCg/GoOxxdb3e6H0jg/ParNtNVXmEyUDBre+EN5pDFqe
y4rmOXaCoZCmy5S2YSF+PjM3fUO/xu2YneLSkG6KA54ajowHWrKiIAecAGUyFQKViZDxb2+Dp51+
pMfQUc8n0YZTf5DQQX8uIsd8ODA5glryW9LJ95aFhlaqlh2FNMOsClnRwkDx2jwUTGljFGDwKgGH
q4IhdxHsxJ2/gTB2yN0Jm4AAyQNWp+s3fvGezUB5iTd3yYDdBLnHcrlxufITGTtQsvwLD6Gxaz41
K25NDbS52VVxTFuEDN0jhaE4YNdZPBE/SNFQkm2ZVtSRmL3p5Loe9/ZO5FdhSJ+lUY2mfKJYQVmR
RMil6cK1cEMR7k7jec0eW9LYeEQ1Vr5FCVB//7mXe8EPaFriRugBlgx6d8bzunX17laexyWS+4o3
Tdmzbdqfqg6MSbKLvOz6Wrffj0hJedvcdIV7iMCtDKpGVF4QH5l9X3oO6q0WuUUedv/scfdpwqFu
6q25+bkF0FlqEcJIujaB8GJzqhJKWGM1EA6u84V2HW9/AaryM1dyWM4PsgZO2uIqjw52/RHuZYEP
PBIyX0xST2sKswvF4kBj+M3JOEoirpIjL5cEL1ttohC3f9KYuKpJTCjwQZngzA2OKqB1YmrZzSES
BAbnDpmFoZ4o2FT+Si/4PWcO4NSyCqr5PqOrzyHSPJvuVOmhMRuiexFy0CnC0ZhflBfDcZlXrSe0
aiNeREuKS8JBLUFCR+euqeVWR8B7+lIeBIYjH3cRDdp6y7MfDGklRM/EQorf9oV6oS9RzE3GEa2f
NePxNAl9K73SJ+SxcNj2dA==
`protect end_protected
