`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
CtbiwgrpAs1rzDuF2zVn0Hxybx4efBT6MFXEOEA5c4Q3ts+UJYM5A7tz7FentjkCAISH4G2Vn9y0
RC2LXZgM5ONPHK2YmEQ7MkSBatyAukLvqpXN6P/TATeIVq/+KAky/MxvndSJe3xqMMDXbMnkYnBj
XOLAhVRSCfKA5XVVeL48Ay+ow02pnUhjpj+4GnACqAJD2CsJDe+a40s4LutTomdFzvNpCQMH6qPo
SWCRlYMBvqGemT0ALkdFUXtlQojq2Gi8YmbYRyA3vqiqXymia6/v1GqR2qJIV655I2Z94db6p0DW
cvPkqrSO8qS4B9bs13beuELZH3RBmVcatIaz/DBZNFVHUP+bmZgw4h/kZ3aAYAM8xtPb6upGd5Rn
RECX+0NTT41YCKqjvoOrL0lnQq3U7uS8FXMiLyWah6a/ahTW95MdTkTxKTkcIOib3NMxxkhV3Z1w
dHMYLN0koiUdQiYYp+g40NLBZ7ah53ZuDXvZ4K3wMY1luSsvAgvBDZrt7XmVsyGHQwew6XjEs0fE
HSj3oLkz4/t70J7F71VF71hwsSz6AVjxkTOgO2VxLz1ecUDWLBx/1Q2r5YrHl984egaTh6PxrEII
mff9tW7rBL2LVaKZyNJ+g0jVHvi5kzgrQTKlzIt2yt4shb3nOcqictX/bBJ1m+rbInSTd5HdxmmC
GeUgUjQM0lB1F1GhYNoec5x+0ZCLmTxuDlflG2uMygbJdKk4iboCa4Aywh4x5VUhGORXB5xAQo9p
GbYS1wZ13xPdKWO45+zQUnBRubgbghroHN56mfRCJT26RNDkk4UQ2NVGqfd9+iOuYVN6T5yp7Ju7
Ay1OhM541y0CUs+uYRAYDeRfKSuTydBag34/HIJuEdc/JRLoQmkUQ/V/vJA1zdwDs7VqMz97TSKj
7/6kshX0YYrIwDmPwEI0hT2Vy9cQey7wEt7oCsJsRff3zOQO6h1MVFhu2hCfwpj5ulW5XO2rIxhH
oZNiLLqaHwN6fBYr/cG2Uzckg4sjbkxlj9i+5ABgs10V0UPaamg9Xc6sxgTwiZVLKgTFpXu1Vguz
dOm5Dv0YrAwTqjPq6akLIcxe1hXQBWN7IuQTkSJPX//DPT6EBgc0poKG773Ez5voTlFq1OOS4pwQ
7zpxPGw+zof4Yh5VxQuR8lkt66iijl7QNbplRfJ5dJrAEKigZ4NQK7WfIZ8HNl71RdG+eykHHpgo
MMDqxSC8nbjLBxZWJwv4DeSV4ssa3Bfa0gXuYuToQHFLNcmc9GjmiYiGqNK58jPsADX2XLmoxU6y
OodmXezbYiw7Rrg9KBf6TZhOqlgFyKeqGpiiJGdy+A6Akyxy1A5jFdriVJv6bQcR9NSx6lIKgn24
2PR8PZD1tjCwQFbpoUnCDV8ITX9QeiurLnXk7rfbKACdC6/CiPB3KSCdG8hSbw6CskpQGAmkyXl0
DfkdfRC8+IF1tbLhIDMVXPkU0oOczC7OIZwcgz1qGi+icA3Mr0zDH/RVSm3p/OUhBk1Ku+6NpXi5
leS2wahce1HV506bjwgs2Mh+m2sr9ZWeSJ0T1KAwVk4o1mbprhUWYUfZoUYYMOh5U5RLX/ciulCY
PLCqp0uJz8GONsuQtbfN6+NLTDl5IpTe5LVr0vJE2KVAeZ02SEJjvpJCbJp+NbMF5paW+jyjuHB4
1mwwH3WZCwfId8CN5qidnL1vQHH/UdQWQYJlq+UxE6ec8AowYXY21qbv7ACJ741aKbTd4tgTsJ03
1jH65YGgBc9cVWzYAsm1Kv6hJ1w/uIG//KbEEovoKvW4yelQCiVVjzBK3AhcLnnYinZbjIkldduF
I5QEZCPaOhgestApyN0UdJSOVgyBa8BFRmONU6pBvsQfn/rubVUlrvDNqHARG5XNr06UKd84KiPj
0ofkzrgNqh2DAORrMxVFITfGtWhaNw8oi8harazmZIucK8lKqFp2L1U3MIvPQwRWwP7BD174CIdV
IAh/21K7hOlAKJQg1vqqLft/Q8Z3cBnnn960mcSEZ2fZzurIaP/a0/NVWnl0hiKckux6ewvIaC82
2zya68k2Tzg2aHgSEsTTwqRWfztsYEIYuRU4lhOd/e6RH8nB12Ey3isZs73ftVkA/6Adq0Dhl1W+
8nDNEtBiUIz5w5093NGW5tD6XM6VZKL99dlEa2BWbOskyFpOmKC1FEqDRg895cEHJXlyte8elV/Z
WHq7lQ6dMlP/vC866f7CNsOtbUsjz81gX51uH0uonJh2ytDAwqdFJawTkgPh94mtLS+3FDZfhb3i
LOt+Wz8TETTqFMVUEx2afuNJqQZJNsHE9nf97UC8wR1sc6dh639UooEKUctW6Pp5tOomCLjn8/pW
hjObKpQvO9TB23490C85hR8p/9jd9+dpe3RqfwfNLLrNFSNcaZYnVThIJZXAG+6nN6jEVBtikVBS
XahJ4/k0Nkxow4TmgrfDjmga+fT4J18J09nmRECzF8YvXpRkK2HRAip2JBjX4Y7Gh+yeMAxylYFP
CEfacBQbCNbd1+3p3NO3Gq9maeAqFA8ZYF+Cn3hCxqLqzolLcIgRv1qbV8ErCDj0aQAF3UNn6mDn
FKQiRV+k9zD4idtJB8HN1S6zTvF9TGfJJGjfxZKpO/eVN6N+mV6kswJGydxIuioMlLGj/ARodPTu
rjqdNb7cKXfsbj8aILLQu7c9mzr9v9ThGJ0Lg4bSAPXcKE42RtNmac4kCV1d1/ReIA9i9f/KotaD
SQl2yUlhA6gRHPCLKFxfA/9i9L6klUmvIFp1ackYtIAGedLVi0GieBIGmvt7+1yZDBBbbKjfSQ3k
i91ldPkkvU34uKYpVM/PXB0lpHORENYX4XsUgTxgce2IoQYtqKL5U2m2rTeDrEhQnFcEvKckRopz
9Z66F21eTbqRamx0deB62szQR2OH8/i46vla5Tn0OaflZjCq+ZOEZlT5i5/Uuuev+YN6JqlIEc0m
fp6Yu+4hW3zjBq+80sfd80VlddeizOqs3w1xpZrOJcWVOFkZSA/UIgisTEFpEjHKzrHSKV6XGoTG
LqlGCyJM9RTcUuQXvRIhwpwcbHx/zKOfvAmqnqflmO29iIv4Rzq6qdVVc1pZMnpyGa1X+9jnpp9p
cAKb7ApGzsbFNXFB+tx8BsYVjgh3vPK0ZyEGgwjpHm2/YU1oNupQWIHd8r0ox2Oeu6AUbX05ppi0
zV2f25WrtrC4j4TBq7mfi/n971cX78Yd0k2uNoFEQbVRtaJAI528eoI9o7RjmGZLW2V2PWcKEvlb
VAbJbj38VHP3JcVCb+mP8GvwYlLfQxoOFGDPl3bcpsZUT7wUqIAqzLkb9Uzvuk0OYZvmV+ICHwP5
luRHJ4UVYm1i/ki7VnL9HABOwtlTow71xtTSDGWDATw9NHvJFFx+71U7hcDMHiV7cLPPLbG8Zawp
CD7f4+E8tfHkiCticw7xHKJIBLCOP4qIxfXZza/2pMHMduLnNNQ0dv/hihM/gugs7U4vMOVEUwE5
WZSV/oZywyePvAqyEwsDeBQP/oc1mLMRA2S9O2PjxMccdbZbPQQDoLrZnvNEchpz8/qsUJWJ034D
0JAdaKUFAa4GtRIcss0mD//LRhq781ZLJIqqu2dhZqIaTJPSEZLsznafF/0Po9dsj5Mk6LQvucO+
y9SULlH8SbPN2NdnQ+KbBrd4Dm+fvZjuze+oiqM8ULtBYcbHcNmjypfp35panPYg2TyeL5CASQGC
Xszyb2riTUMj7Uw2SMwyveAwsjQ8leFq/tXpqznwFY53pTa8qoGsv8eyFHVPIC7+vhzL4cLirVbY
NKU+ZpHVjyMq08nNtfQtt3RFd1Gc2ylcM0UB8wt9zhxLEgUVWuo2cAv4VWQqlebMYAdzQ97SJ41P
RuJ8giGgAE0wxNyAnh7L+odG4kNDVJOPaSXLZYo64AETMQPeu6R7edkRUXv5DNJQ2fsj2uTPa6eE
itwkFdLHhlxPUMZsBvDBuzhf8FguI/5UkH0RLicGfCjxou7rk4Yj42w65IUKjQndjZ7i0iTKEUnS
7uah0XXMISFausxZSS0moBVOj6nN8+IwBGqbJfHr4hOUG1e6UT8x8sFpGvHGzIPsmjEBSFnDtvjs
fM0MrnzB6Zl+FjsTxD2zJxZ5AHk5oTkV02KfL1F0ajDV/CjXGpNKd2SP+77iJkjXtvu+YsRKz10r
dBciy93IiYfELFc36ilo/DZ1bWvexEUCK+H6giiJmlGE/WwYFFyxl6k93y/Ua2FRA9drDhMrB/ld
PHlqD5x+gXJZroGdWIOGS+w98Dpkcs6O6P9yRfKxF87TcjIY1fHvT1r0+M1h14GZIxgAlgKYXkX6
KwDgQqzLJfkD0Egzt1RNjOQuTbFPXEh2dlVHglo5rNerbtcCuq/oo4Py42VVSM8aKKqZ6a5GqI4N
um707jpvbbB9IX/qkoVRUACVLQdT7wdU+pbKjjI1oN42RwqPhtybS9K2hgddnouv1S0GypMMuM1B
9v2Ef37W+MOnTQlTVOGsFO63iLw1DSJ30eHiaYq2U/JS4Dpadzcs+VvhuTK6kehlCxfWl/uGoI6C
dssSulaTxTMf/4QH0pXZaiVI78U9HtA6m8IcYjiQUVL9rlQEewsBZghN8Zd0HW0ZUENwJRLw9w5X
Raajyue1I5sTzl3aUOAB25S07+P/72F9+SqJ7CWUJH3ULbKBPmclTgw4DC1Mp6Q33KYe+8G88585
nEvhaJHS15YS03zvcMotat3RNnGxxrassPBumFnTDQ55tzNWgV/2z0UfMunGuMg7UwEh3Bb1N8L9
DM5IJLOxAwWYbZG6zpFQAQ4I9NObM+WTwpORWt07DNfwokaDVdU2iUrBetnS6Bd81u3Z9wc9k6/7
DsZDWhoUNB1gmRC0JdDoWcglrMw7x4CWKKWgE6t4O+tTiPe2/uebZHzdUw4CVnNwwtHHMBrMY36Q
jjt9hFEC0G9wBEMnuh527M+CYt3FiPPrtKjeguhFqHhZcsjht+ve4mRRBaySV/I6pRdYw3ZM2nia
8ZbiKf8rII2s1gds70ihF53mduE/4g3JZM3hyX8cQV03SjO/dSOtgsX07uuUiaiQaFgwDj5nK1UA
g/2zekZo21Sexzr877zRtPb9nf6drItWJGxn0itkgyVof93O6yhQnwa9m/g90jq1EGsF2ST/KnxA
x0/ezsMTtartroslD0I7EeiCQQzB628wcmaivbWCkj39NdO36ZWoVeORez6iIiAjidxGfGEpbq6c
HhsZGVbmrVOmmBHjK66C6P/1Z4Uu3P526YuVHSCgISb30cVjtZDj6WviwDQPWTFnqVx2IDxl+EDt
Bm1RMLwcv0hvSCZ6Qsh2K0OuJNZtHUgASJn2XqD3mQMaqmqEkuXD/aZkqiNbuitbRSu6iciVU/Oj
ektRmluxDvlxcUFWOty14wa4HUwwgLukWMYm9VsIKKmRPSiNjLvd5/nI+EK3pq21u3tMR8w+OQjZ
oHjQN4maqQ47wCP/GA8j2g8Pi7z8jVq14+ibO580Hz2nnLZFn8q0fH7KjQfwd5ud4FXrrkbq9/oC
aHRgUyS6Cg21clsgYhWKEKRFkUQW4mtqYlUMzO0eI0nlsJC6WGaluQhG/UtBhzucORGd3fgre2LF
wHMgJOHEUh/8PK1qgrrNQcJUWD+DWm8GreH07/BwkBN2XJWxJH7S59KQE/E8K7i9DQxSTQajIwU7
BzwfapvG+HX9G5WD33yT5dt79mQQyuwQkRWlgRC0WKlmeQLMQRV1x9vWQkFyvUPm7HlBAoT9wims
mxJGVY0Cg9rWAmSd5XtyJsTBasvfbcu+t6c9xgys3/85kZ1HoZO0Ch/XlYfE8dTP7/J6/KL+JEfN
N0aZ79JuvfBePWIO00hPosKGNh36gmKev4H2Js4jQlW3vCFgd4yPlLOaC4yvZkGeGfmcT5PfR7u8
yjndH2xdpZt2yawZPHt0ukTLacjwHejm5BcBLk9IMcH4drzGDKhKmKHflM2GITP4ZTPN7ps47uj5
afFnHsVuhC54lRdxxK10+kwwB6D1bQV08POfTH40ZKubMpUgwjAByB3dXDI8OasO23m4/i3Id9Ma
LVd+fXJi72e2Hdw/1fc9XQhKS3bGJz806tLMFwUvrcw2YhnXirUpbU30burXbGjuZYc0tx14W1KC
9QOAxhKQPJA/AT2aIYqMCDhS094YnRTnjzkwAMGpzIovomv8Flov9Sju6I473pYUDE6UgjzyW5sW
XGCB7K1N2GZrRcRMNELBvwgyFJwpdaVzTSemIPPcXKOmnuvxQ0n0oWAN0vS6Zv6Ea7CDr8hSh81v
tGVDQa4eGYyxCXDe4ty0qCvIz0IukFANHfXd8r2QRQjEF5OG2+cdog8JtB/vR6QWfJz12IPLnicy
wMEa6JbE2Q7wnwRqvJWLkc41E4WGnyCrCrURcfYmhjzaZMtFAlWPG94751BqP7GPznEqbxnmpxEI
VAkj8H36DZ0LK9AR6nUMc/a+0G0OccUPKwb5Do5GY/7dxNc4MvktbDZqvmj942N7S0uClJEfoy8e
QdnAj2vhEXwgi/0XjCIyWkyBNEfVZSzIqHfLfQRMClXgJJbkmHki4yr7c332iD2EDEMmZ/4JV9Gi
XGHvlVRkywAGHH/Irg4tcrHgLz57B1AXOl8gKdy+A5/j1W47Z5TC3qELB5ZpCN4ZVqz231BNS1gj
59zNRbo1UUgTIzNBjeLVs/YXSTKJbMPEUJeFsy4hxKVXEKMRrMM1S+RsZgH886CZt6nhkFWWhkaO
X6xpTii2DBbrOfafdQPwRWzw2BPLn7aN2LqhQ7jqNroaKZqAta1XBTDy8gIGl92k7L+zbwp/EOQt
yGoF2E3oVzn6+srFbISKW0gW1PjEsp/zs5XcdNKM1K0pCGNHXv7Ivt2DuPRot0o+rdA8c+9c8iME
v3x627qG44b+ooYtr0p24AjnA8a9nax9HH0F/PwFkMKPvdHO8/dxp4hVrC/XHuzugtTbZmAQTJJZ
kCy5rERmb98P4vT/zyQwDZq/1GKaoKGRVIPyepq26Dt9Zre8bn7GbH9++5AuB7Z+5NGYPPeiEpTW
MaKaCWycm1CT3UeROiR4F+yRYECZLqj6lx349dfGirngjnAa6ITQ1o1iSBZQ/Gw7Ffz7csjHniCG
Dd2MCLgUczEvGNljlZVU03I5aKeujUr6KuEpVPqejwhRGJBxDjs+N3ZRaBhp1WnsaJwlvup99piz
rVWpQ066R8XgWCo0LuOgjtJIpB2d0VuYFb1uUuyeTKZVevk/oFGmqDsbezPRp9WtmVJrRhMLAO/k
W5dQUhrHYqb1v+I8/sBAuk2mr2RRPqwXOQboSBPboyek9pjA2lNHwjbGL6EYY7HAgcrinEBSrh4L
4YOO9qOZDH/yyQ0LlMfMIQ/ZLf6A4qGss7i8DszGYhG+OB/eXLikN13LWZAC6taxfXCQJ8kTutmK
mh6s9mGreV4IaoTA85B/6LydkBmT1tOdd4kDb3yblu5Dzus1T9/QeMybmd6TaRMtggZcIVoiL6F9
U7O4WKj7RT49jsHV/97eGvmXT+j/3nP25fk8JglhpxIgsT6A8plHDVZl43URQoCCkMszAd9Mhwy0
vsKE33YfM9Hn6y17NGEEnj015cU/AyZl4tSJWDkrXrEGHMDdnjH6/Vt515zmEst3u2ZSmNsYQ615
nRaUpnnZyzXBugrnA2ZMNiuzWYWxQisyoZtqqcGkrDjgChfufWp6mXP3IYC3RUzcjSyYxp8M90XA
FrWNnkugsbHR19CvOvPg+QtQIks7WzIvmKUA8dtxl+5vkLvlCH0wpU3bHZ3vCgtXBaZ3+EpZSYQH
F4A+fbNuEGSwIUuJr5qncwJk59IY8SDc1xo5tVQc7hmDOFxS1ppXu561RS4i/T8j1c7pyTbNrTME
WNV0Sty+BbDrCULwSumvA4Le9SmESp9XIHo9NTwA8NTM3FfrmJMyC9xTEtuQQoj1pct5iCL0Oj+0
9QySXgliax1dA50t2D1+2rHeUozdi1HcFgk3Dl+kqqCvHY+gD7pZEzNZUQuvdJBCqnYDYED3OGkT
/QvJx/nayn3b4UZyoLqIhUzWG4jOsimPDMzRvi6OHwsOu7bpj9+jD66ILayEBbTRmfjrDuOnxACZ
WudCUwVtxVnU/2SDX2T5H1RZLFpxQcghu0b7NlSteu0e+jNP9gBSEhDAkl1TMSxPUE2pUuVVQlfJ
kmRIRTMvOzy1A01NLLQcl5t1Lv+F3YgvXx6D0h5dHu43Sg0B4iRHUqUjJeehdX4xXHN+T1A0bBEs
WK9iOwhmn3eXTonUVXalGq8BApvvXbdA5PuvbyZDaNX/FOKYDJnnS3IFbe/E1nh9TViY9UhebbfK
nW1LdQhJ7EnWGZhg44mgnyOb7MTdxRhqlbWhQDHkyYIo2t9MR6CG2ucUzn7rP9Ba+kvKWteijkaq
EaN2Jwu0XbP5naKpq3WxBjGiA0KXJgw7lXyItjlBab2brQ6yWe/KxKyiz13B1Auvr3MXidy7KAI1
a3ozBIzjNKghPXpATc5LIgl7yDf1J3nrNhiQyQwEIF2oSdKEuh7YnTNIIhdlF2FHfdj8ihhPc8ax
nGEdwkd2hSgAXtyL2NZ5QCdxrAr4Ac01zQHyNSxvOj4OyYWIX8K2GIOHDhcSsbpz9fsx3xL0uIfk
VGcTZwJZcO0jmwKwIu/ZE9aB2Q7OmjALaY9bEW1/BBZXHz4nzwtTAWQkhxL+gcwC94HBR5cwJKqU
g+8FQ6Se8/rLHFtrZ4vzuQNEGAMHZusIoTsRj8lKcYZIg3VXWZ6WBqS0IV9u0lJ6aQKq1w+7NtOd
DvGf+ir0r5j4YOZrtxRYk8GVqwkXnP6ySdnqULUwU6QfMHqFMlf7lIKhnyO0I7tkoFMIV3XsHrJh
na1Hv0LtWw723n7iC8AZsQ6m8z2jYTp49sXxCOoDdkTaGwe4B882J8nR0FVm67vu9VirrED/y2MA
A0MC8nVEx9a4LvgTYZqzpViezpLi/DnjxRRhvTYKOD23XWUA4hf55EOb9BCq6FdNIu2LQw2I1wdj
TvhCYjOfOBh8op5/8PObSaHyx1ZhtvMZqUV6jDeoPKHyyRa4RVpCS1Ih0YFUbKUT06avvfJkXV7M
5qRbItrze5Se8JfFKFUAPYyu7IHS7Vm3b6e7xHMiN/e0hYq+9vV5ree7lN4lV8Z2M+2wwywiV8uZ
+JVmOPRvWhbUjCsH48ZkHW3HGzrtG6shXZefs1NGQ1rr7jCdfWvVLZ7AynaL0ZeIErrBp8DaPtDp
HUmV3jMch35wAKxgete4Tm8aGeYCw34DzxLNLMQHqsiDj9qyh63Jz9GduHdZ3hCoT4S0cpJAHnGC
Gv+DUz05/3+HAder5wbfcKRXX0ldlHUvo3qVN1hjn9azSeNQO4CbfeuKuL4hvq+ooAk34EimgmPx
ULVNJ/sagGEeLtf/aX9Ujk77ojuAfX9AvRfW+0oK+jkxGGU3PeEwq6ynldnOk40oSZ/EA2PgnjUh
3Iks+T0aMvJPVQxNxw6FaJdLHEL01V9IJnDSLuMIQwOM5VVP8cNpGuTEoA+sUbGGAKjq0tj4bJWw
2Oflv72bcwXIrm1qMiCC6099ZGoAfBT53ejNldEpYvnJjGRekal84F5zTJsBS5/U1hJ6Y3vvTBPE
uv9uy0pfA/v3ud3YmlnqRy4sT4fXs/6xjP0yzvRAMW+OP0IngwOwmN7gY/1MdFHF/3NmULj9GuUQ
UgM6ssZJNTLXq6kXxSvUVObKR06NXHR5bJO+zQd+ocdCtt4xWvkICjtIQXwBotn7V02iLr0g9Ykr
tl5OE/tDeHfjv+RMKnoGoRmgatvk0MBJz8o1ZdnWtD48+MXa78W2NRKZPVBDLobfr2ujQhVrj0Ou
uHCNTrIYlXECCTEhkWCQoGTJEdXMMQl4vRsYODhKLmUFvFk76K5O75SSU0RmiWwRtklds/v1mLkE
tgZccIgMu8EEGrPDJ1pIqISAO/Y9uTgCe1oBshA/Yj3/l9jSGOsPNkPrwnrGkdxaaSZZBBAoojBS
pDVaGrlEDVMZUUhn9etzhRZRmiiT88GbAhrzCdxCMkG7J3Fymn0Nk7bZON9Ne98Wkfn9OzP9p3JO
xoJhCCZbKrpY4shRspITDZnkSgAqhenX6L2/of6YtV2PSytvYcn3vfWbiBDQ9MeearQlhQV0L/FP
2EcFVJYRI4w8Z1Zpy+hTIHOlfz4HGzNC4ln5LVvM1PGR0gZ3j6jtyb1H5oIg5fNcEMsGXweIwXaP
mX/SiJRddwfPNI8J2/mHwwaYQ5atlgcXEwzkYXmmaTqNnGcH2qQxeLKrqci0recneJv5FRifLbBf
2pLAiGsKHbrECJ6F4C6V3XKC/8hhGl1JcB5kzjg34pJttB+v8D3BtAtRmQ37ctG0rjhHYOBEozmI
LgfN1MVPv+fmcH3KrEiiNd96ZExC8G4AL2o8Xnhaz8rrt8cp4d2UfbLPnfsdya7ga+dTWo1wQ/j7
oZhFBhuo8jqB1HN1DahQWz/lmdAs03HhSk34hEGOaHUb6wd4i0IoXtHr3a8SoUn3O6ySTdg946o3
gGWayHSk5zbMIsPox/3h766Qd+fr9J0uq33bqJpJi6Uxo9gabgsfOedieKm+KOcteNgTcLhK7jhS
KHkSQ65QjTCOJIpRTOpJIbc4B9BGKWvIcBpjQiJBRhii6BQtOvxUf+CQhyRgO1lLnuIryaSQ+fFd
rq03kiITD0+k4HllV4XvOAHwVsj5OcRF9mPVKWQ4qBpeG/OtXHEB6IDu7pEl9siDtbwIhuWG29h/
UEk7KMrfU29FpaZnLn1iDzl7DC/mFgSSTnwstls2Ikj29mqhUdP75z2a7rYIthDJjETnI1Ow12mb
A0xaoSTcRMBxcUpGj4P05pFtFjvTKWEkDauFUewFIYfHH/BpmZIx89Yh9ceOvziZ+ZsoIJydno4W
Qful8PuU0Ftc4kIVoYJ1zXl7ieGwlsnkAtt7SnLh+qgCpaHJsHoeQgB29qS09o5Dtn/oIFp26tO5
KJenchnU+G4Hy1r8QAVAEIebzeZudxs/FxYPtxAKgWiIT4b1Gp/JpaT8OdX2W0DWv4q8gT3lrNVE
4yGjGotW7+ok76g+LmXCZmpIzNhGseNHrzH3TMyAO8HkQHoCtW1TQew+gTWL0TIewl+GP7dmo1AU
K0ak1XHvNNAqq9/43NLEaz7a+N5wO5yVrKFl5r0uDJUiLXY9uGiqxFTf+9J49ZIwigOV6+DGukoJ
hK26+I7GpyuEMgUjAQJc+wtqM1cn9MRG6BwA1XeAlnrQycP0pHTl/D44X5VUevy4LL/MUQziSbRo
Wjy56he5yZuHSlqNMFr73Qx41Dn5LrJeOIWspDG/VZF1KzQ0DxyrUGdlGhnBe3uVaeGD9q/beyNy
EhAesFp8JtAbdcj3ak4dwpFgxq2/Ckl7CDY60f32qRKQmfQBNInhv4Tv2atEs+PzxLIY9Ek2Ikeb
acfAus1h+sxcw8v+nk1oiDoeEDuWf34AWemSTDSpJeZb1Uel41PAnxIZLrF1VVcwcyC49sB+sm6u
EWa+TmLAOpJy7d9aLMdYYYvf2m1gKYgaPVX/+/ueFhLDDm4WlkoUdoLbZOJOBOXZw3r24ZSVTLnN
aTdGRaHG3t4jQIRqXGP9hMmYZHKRLzGiPq4qbw/YTme+J0TMz5JwNuzTwGWwDIDvgx8x6Nd4kSSq
Ic9BFymM8v4iJv5bJtwEugoc3pKCvsofJzgtS9ya06L0vXTw4FBLBxeOzT3cVy87KPVBKuSfrkWs
coYT/pfNDqdmfPnUdabB+1d3bU7l9xjJY4I0fZiC3SzzqD4IIEE1xqltYQatsHrdGDvGdbhRWJuF
wntaAUwWEatL09nyLfXdyxbMs6aWhslj0IrE2rekfv80d1E9nBhZwhyVDahMacjtSdczqdCCUXon
qb1u8eQWdUljbr0IgkThceQu3ZX4cLzXxWekVnUYVE3VTXcZQxigWfeJn3QB8ifDzv/4oAQin/9P
05HCivZL8M9dD2mPsZ5ymG92Xit1DzEYhjH2+ZT6y6rkoQnGjV/VLIED1OIF6FDBz0BUxcUSNeYz
PqT4MbO3izlt5UNPX9iUrXtV1nG4ejMXPHZ/bSF3uLn870+TiKZURuSaNH/4wFVUdxZouhP2xzs1
AMS85EjnhIIZbgtq5ORpP2bFpGKoMgW78OAnMzwxQ8j6Yex2GahZNhJpxRAr3uVO16SoGCOXaU/f
rVI+JO0ujngeXuJ3s7q+JwwKTolldTJbv5irL/QSlSQL2QC2NGX6Hj5HcpEiryLy739+BGTG0UkS
8we9tZG7d6TzqZG5axknRvkzaHUv/yB5W8kbW0XDRJghlTBAzcs8XfgPrggV3jTK5YSRA0ecZfPw
Rj5KMk0OOnLAWTTs/9U4rAJCcuJMQ61pPqJCyglHdcBTve8ayJwEtkcKB0Sv+GUu6CJOAeEVsgpP
jbZ8i/p4andhJCeWmM9QDBcPuFmoK1+vBxFoNJeXGN1E4DBJ3c3NX+N7E9dsl0BA6w6QS5ck4Nzr
Tr4cJq9GuSVZkSfjzDR5pKZbsN0AtF9DEBcsUeyB0zYlvU6TFWfWQVo4FdNBhpWCtgvYQQoMKOAt
XEcYKjH3rZvZAQcd6oRJf671VDYGAZgV/iIdnkt4EQVik5i505l8FvBwi82X7v92OI5g9hvphg02
fEGijCGJxddo8XLVhm4p5Eo/GqOrRFioWm5gO+0TETs5XMFSJr9DdHPyknFLrA3JkLpkUxkJwwok
1PGjvBzb4IR2rUvOLrUbewCjuworx+xqW0dAe3A8CQoD+N4UK+TS7jvgHrxTFkmh6zj60lBCpqGe
p0NQ8EKm3vYH+t8gd6ZRPW4onXGJJxCTxiwtM//aU+3LRvHScU4SUFeDE0efpWCyXIfIesb9xy6C
Q1ChTFwun27LT0JOIE0oG0+c/ExADht53I4JETKk/qhOEMD9weDEJg3WzoUAZcT4Wslghn3X1yOf
BdSxwQjS7DaE8Mi7D+ucVaGDbcub7jiV333F/ou6eUAe6Sei724fiZkMifb3QZsEwrDaAVPAUFoi
T8U4ZNuGCHoWT1n/ify0QZ/nDF+WGxC6EUFZcql+ljaSUif7hgYbnqrqs1mN8XzlkTTpAqlZ02Xa
XTtKwcN0mgEoay5MW1oNcVdEMt/nNxcOW1MKmLIBo8kCdeTPE6X4Yg1BV4skaJGwCzKEu3QMZ/gn
MiJI+9AaeILV7vv8ogrmvqnabdXhyEP1eKT19mZHiG3TkGrufUXDbFRthmsdUMklM6rA7gRjN+r3
VSazH56ZfePBiFyFaV6YOHQ3pgh2/ONmuJ5rmDfbYX9oT2pwCJlm7wtBjfMoffLfk4LDylpAGkAe
Yvc8uj8eRUVqgKyxXrckcdl5YAy8j4Bo0Vt4th1wJU2tnkzleQqH/JJZD52COjGvQPQ+RfpjfT2g
aZA+jjMpJ3ap2PnTZHLOEngscPqYMTsvTgVOAJqdBo9ocJmTBohEQQZoBYQ3lxtGW48o0M4mcuNI
bZ729M1SwBxxkp2BRNdICOPzq5RmCw1dZAZngZ7e2FEULn37S8jQN7ydHAOLshBGpoXKIhXml9Uh
tf9vDHr7kjn2i3rBomqP/qCJIcTa0EykGCEZRH8pdOVLp1KksAek0BqtMGyc8c//OyqPLU5/66rW
ck4VmR+VvQCQtXVBOy63iRxwNba+1j1Zw7AFecxZZjho9gYYf0VcgE2CiFKHvQtGFDvZ+7hoWGME
LNyTcGumjH8MgukXjvNr4+fQLxg0NOrUhPwO7eOVb4G9K+/aQpo7Ck7UA84QxzUiaMlKn06lpBI8
444LzicgoCHBv2TFZTVJrKDM+OxJdMHvGLPj06nJjxUVpRhWq26RXX8kYxaOcDCdUMX0qQrZmzs4
tS14OgNw4ApJxXhVfL6omNazh5buiC0GwRWXKh6yq91O7BsdRwXD8JpCc4VH31kpKYaSgPyKaVsE
GfNiH2Lki5A5nAbDS2WM3rkObDf/9Hbl4O2ghpVbFvDtgyUd2FmUqkmt6YP4QXTHV7rb2HjDzwaH
76ZhGDAzQ72x0CZ8KP1GxL3sbCk1zOAjdov/u5xZQUdvZ16E2hZ5ozJOICmdmiljr77pJdAVKKD1
qKY7R73Lw5MXcrpLHJmD4citaKui7lVeo+20XUjIoGIWirs7doAdFt407bH1ZPSvzV9WAQPuklHm
YOil5QyN8WXJzwEsByy4nv76z7K7F3nhgjWk1BAzCaDTSpuuW8tpONLH2LNzYHexR8BvKQhhiWVH
1xIGh+9BT17K010IaMJsPbXlTjq7BVZ3BW5ZLwzYLMEII+X+Yn2UmuOlb1tRJlIG9R3Y2gMEkyti
zxNSvW/yfn/axcXELcaBKq1G8QS3K/S8rALI6PqkXQ3x2A5WoWOx2Y3dSgRwYlnEdBwxAlCwQEm8
8h7vnejXJyOUk53zsxVJKxBVfncmhz7SbsGU+jhYnAE/+lcOMyDGSE0HEVAacSvmkSnBEbD6YHE7
TF1OY+DX6yJCFKZ4oLKI61ee6PF1/xGw8Y2vLVYYJJ6v3kebT6MBq6Q43LSxM3x5maUByIYCj3VY
ubRM/DAHzzXMiwIGEu70zUnOAr9fxGCOBRnDcaqGByvmRF1m41UwhhwSJrCTStY9xnM/VgzZT5OT
KkoYG9y99xZRgOzcydNeUOYMuceuBaA0rcohIF6/BGpYV0S+CnlZsezEjEBxn8bTFxRYvmp1q4/X
rXkWzAGfrse7hK4qxWfnFA27EpiUAiqh3LcZumHPr8gfTCnqXQsCU17KShJDPi/DptfxeCAscJUN
3tNSOdtgm/7GoEB36QHUPgXr4ATEfKqDVq8ICdIjhV7Tsw7MJkWrLxXCWscyQOA1WZWPQ229EBEM
oGYeOAZEsjyksgD4twPZnrfO/l+dXU4X1sl2s4HTPe56y/Hy5A3RV1O8tcBr+aWHzLj455yplSFk
fa83p2f9O7a336PdZK9O0GzBHBCNmDUjUdoc1p30IxzMNd/VUM4UTu8Jh+16sZEGIvy6IACVizME
CidSzorwTRujWfFLoarJ7XK87z2jF2bgzEvuSHvLkKbl/WwmL4QXfvSr+C7x2cP3qzoebJsa+Vvi
cliwHP/BQ01Yy+d4aqx2E/Id+VwKTJqT95A1ndy39sLkytUmqr8BRKzMBY2zL0JbYAvyiz0yQEHa
ENLmZskxTl8BR4E6OZGxt4FAKUm54GFHtbYaSUJ14uGLKhZ39lR5EOHPOZPCRXnmol7hNkkzgcmY
qXOembEfXMkEq1OT8Wk7R6qxFl+KuT/Dvc4B5N31Wm9znwMlNiIMJ2Emwk3iwldHBg/KFqVgTUwo
HA1Vm17c81PrQttCZsgawQ6ZNjI6PpcsTrRWq9FMHDSDvO0ruUibr39ryiGO4kD29Polhr5ASWzL
ffF8pSLftigUTMjeZcS2NMoHUZ9LOMqiXtJ7eWfSLEhFgKmn47JTvsWeySxUvywVpLb6/pTWjBJJ
Wp1a+pyfES2el1XuQFzpa4nmMkOmRiJa4jKEING0Tx1wDK4o6mUJ+LHsUAmgxqk3qt+WvkFEfKSw
wtCgF66zOSb5on8F+l5JClPPeDVdRJCV3NjSrQVoG+LfSwSoXfzdL213Rv4GZvXplJ2YMUy749Kx
AfxbB0ASMTA/J0Tqnt/WK8/Rtcpwrh8buTl5Fwmf841pd8uG64Yl4eZWLTD/Mb2ajQYvdvC01+fa
InfccrKoRqFvmFDu0T/F8VTiNzNyb44KlqVuBMwlPQl8V1NX0IoZjPOcZ6EMkbmQ0iQQjP9dEKW8
tb8gBXvdAGLd/s1s/pc11Vy8dpo7mNDTPRHhSuxHWxDkd5vA553t4W8CtgMVhbFb9lm4Rb4ywNeN
k9Riy+bXnc5GXlBUAVReeaS/z15SNornGgNrDz7zzFJnoU22fQKJgxzOYjeuW5wlwJzPumf8NygF
PblkAMK2jAdWOL6rf31o50xTyEJfm/f7sZcz6B8daC6CB24i8sZAg0ddIHmEwbKeaaSOlt/U+7Su
R8Up7yWv8TQU9rXTzku6SC937Fe8m1xyI9EdC+y/HQxQKR1aHS3VQu13kz05T7PS2k7nvJPhCuMt
iY5Rw0R1FSfntENgb4fRTBjMLW/Mb9AN/UGklTUuSIMs/iMAkrH4OZoHHVaiPLtg6lmvcjsDPw0x
ynSTVeH3NZNuhz2v9R7x6NiKK5yz4tgONjw6LB32TvcHeNPOxRMweW5cnCrOYUR1XiXLF6TqiSfC
NbZJWzINTnN21aeYmF9kO+7v23ufoedRO2gySKqijvAwaY25kErgyeAm42kVA2BEZES/AmzMohDM
9WmUTmaD5BrP6QE5//jKpsfaywEnoo+jw/fe1a0vUAO7mmhe4nBBjV+iKZWxP6duUKHmDwNtiA5z
khoRSW68nkjvVIfGCvLY40hM7ftHLOplNtFH52KkCxN2Q1nd+kmDOxsWmfX4T1aZxNos7oMtKLR9
HiPsNnwBeU0RRlXBkNtu2gc5JrhvU4o1Z/6mo0PdUHH3n4mbdtGWC60/JTMxACUrgcCZ0e9e8AH4
yiRlRTLq8uJdpCxSb2j2rNvU9rch/x56CSm0iOGj69sujJOpqj9SsB2p3kXjRRKuk0diPJU1p/V6
puau1OIm0mEYNsIXC9oxwmfP6tNiMXnzROIszUo5HZ4OyCor+03DuME5j+rX2fNVsllPdvB+dirX
feX86K7BCvVyJmHxrkQy7+UsDvX9jig9Vu7qv1dUMsoNX756ShVh0qsQjy212sTelTRlsFRFlh0/
2A4Fj8SuKqbhVERjrUO/urgJeIPCuVb/Sw+Nql8ocMVgWDc/CUd/35srRmmsGNaoVuUIUz9oIv7p
BkuFdHiXNy4wvQAO0xRvMSztlNnuNUfpMAJKoDAAWMS/u0wrLkb2eqS1KHNJNgCjHFOHx6aos6KF
ui9BoYaGoLfd9cFK3wBA5FwNSh6vGgUFg2Cw5ay4GG11Jis9MdpbDVPfsiQmyVBOKY57Y5hTjJHU
ubkXm+k84rg9VnNayRIuwcAaaKNqvJ9/e9SaUT7s41mJYluGCr6xE/jJI9XWv1IcPnxFqq4ujOSS
cmkjRt45gaEYvN5ZbPRSBxBhbdekyb2krvtCJCOGJlOpR4+GhBkROQ89ew18YW3c3b8cY9lBkxjn
cBwF26Xl328CvDbMv8c5WvP2fyIiu779aAYeAqCdK73gwynUs4o1pzHTyF//EGFC8dmGpgR/kdz1
XP8JH1Cf6BoGEHTHuViCk74MBWD0+Yn7vbsnSFaL13xrUvXkrNiuWOt+iteruA5DNh9VNaE+dExY
OhyvuAGGGza57wDNSD4HizXO6Vobe86RL0ofY30aPpRVg4DTHRBItDnGFP3fMHeA9pwjZmuaXiwe
zPFJlDipJzGMPtfs42uiCTBLl1/LJSGXAakjjIT7HJp2JJUZr14KCAs9Z0BstEmAIBr5SVpYvkdE
XxHrHE8rSVgXv8b/dqE/T8G+gHQYKUIe5Kcy31cvcDt/IYzLCwVSR4nB1W0D+oDBD1vAz/H2BhEv
+WQUMthGqljTD6Dg+O0UA7v99xmYlCN9gYnDTyr5eq7TERAUBjckW3O9Sq1T8oHFmIsZqZITVIjV
RJbcJoZHVy9INJ51Kvml+VKxlwqcj6K03QtS+A43OMv+yxE/ALfQNd7O5yg3FowasErkdb7CLVRJ
0tQYnybKleNgKLdXxnUAAWSdFrdvAcvmigXZ/t+idGPaU9/PltS5hiUsWWG9FJg1LtIXo0HtDO+u
s0HIVxt3C7/SVrLIcyjLJ7HtyK8eAuY0IXUmWIUW4DyctXI6kukp04jjOlHTEQnUOX7WQtCZzPWz
oAqPb6Ez0g6xZZvQSGX9TZEDpmM29UWL7iGILtxrzj7oygblajAkLK6rSvcTTEwvezUvdxouygGa
KBZAwwLKbqxc92517up23aofGG/ssD8LyxyODzD0LmTjIkHQtB+tD07jY4rQFAdIOMYTtqRYt+vW
pHj3ySTHOLujAYU50LCT8tE+NxerMdGer7pSUi/4JrG0Bksz+vDsvpil5hOc6OpnS8YaQkbY5SZD
r5lcrvP4N2l7DDF/rTlOu5kzzlk2DMyNSRCs8jDmEiaPupIZzAMrLmGNlSfISvNdY10cB6mlax5r
Ye5Gr2Gj1HP3qyCykO+Jby0UKYXCQqTGOBTnqQMVvVV/twLY4bvjYWW/PdwZHugU9Sd1S8LYSVF6
SsPXYzZGpEgk2B+Y9NGCAuD7UTpU0MZJyghhRzkWhe6sbTVXRGKZpvb34/UKQ0Oxj1D8hu6jYuBH
3Y4RnstJ4lJJDDwNw9+c25ueYxTjBkyOfqlXWXH+pmZXfUhmMdz3PT/knmi8+DACRBgj0GDPMBNO
dQ0tLSztM21b/WbSVy+Zu/aOXnZFmilIg1Cg/ViS9UX3P2+IKPxOXfQKBJwB3+oVvECPXA5AwIpt
vZGCyRdk+g7n+bXpUiM2UrXGWA2M4Yg+dFPVXNvk1UCdPpmJ0CUzjiuTqn5a1y6xVepQqWDnmpyl
JJ1z/yYHxiBYuE3fuJHc6+4X+9jtHZXa+fOa8ZolSn3Y8SG7iYkfIlKRsojzlQwS4Wzan/NwWWKi
ZMBU19AM06B83H7fbZxKixblfg3LCHePCV9BKJi2vykcMYuQRYEbm2Bmbjq//iibyT0DVbbKRpEL
DzubR/lMTl5518McKlpckBdp/6nhbFlI99z5rq/XW88AM1UMOT2ddVFxXMjf8eopVquDo+cYRKb5
IOxcJbjV/jP0vfkGfJrupGr5jOWNv+47SUq/fnERBOvK1VQ93cinNai4XAbQbLgD7s49aOFO2vbk
/I9hizDFEpPQxSdB+YWFl4KJT+65sCmoLjXvBOuDgz9lbh04QOxgnTuA2x5dzLnPK9vJkpP9gvn3
7mz1PWxyzEmz5nq2sWR/xr4FQd8npfKFy9+H/YAyjpnaGsq8sn8fO88xK+cYLIcLe+XvjDeWHtHo
kGDyop3q882aO+48l+6fxV0ZepHfKUwWVrshq/2/NRYt7JZCW8eyRJgaOZMvjEwkM3VlhS5aqZiq
OoGh/lzcgvgXpiQNi3AxqrpEYdfBvrwT9ryJX1tSxCTHPez+Isz6PI7eeMfjOt+QZD68JP7L66Bo
WW6Vs55vLyykYyt8FshKM9TxBJoIMsNuMyvR3yCSK+MDFI9agMOyH7n19vHlb+ZB+HtqblgjDu0B
QOafPR7Fb4t63/+UTP5+ZAsSGdU9wA9MuZfKeo/MFvu3BqsHlaMq8Iz0PL/ueQ0qH1rSzJH4ULGZ
4iJ1D69wJrlXTUV2C242RT6T9lH28XYJagpURHoVu3lpRyTIxLB/eoMegzdx7Cvnd150FAQreEUg
PresKZOqlmiRcjBVkg5uctSsNZwzJaz7R/A4cm5H/hEpPcQ3/rYizFwgT+UybSUQGTGFfol4BXAc
OPV1KGwjBGpHpznPM/DIhvAhaGNX23rcdVeG4zOHXzqQAJ53+R88DJCdEh9hQsifTEdLrbUTH+B1
gDV7JVgH1OVzpqspevpMsYk3WnIvZq7FdVzrA3uqn9CEbXFrPhJr+oLl5olu1eB7O/shy0KscOJD
h8dXJau6K7eM3nn6xo2yA+ThAHJRHe7Jq8fj6zmqzJpSQHS/NJAK3ZFfC11EuVZ2vSmxhj1OsnSi
C2NR83+L2RuOzrhyKUQSoYDkPP8brrcO5IaG/Rma29/hekOYuLdvEECH3x78T/txqC0aIt7GjSeC
MTi1+Ei8JRIzByPDRzSDQ7ezmF2TiBzTwzoF06N4w5ufuBx2qqJGvf2gGY32oVwBkLaGN1G0rkRg
PRJ3xJDMMMAGKvUw+bN1tU1KHT45Jdx7Ujqb0hXx5mvbZsxP2nygiG9KZkIFoa42AsoebJOjrZ1+
7YbfoLhd5jMpQYa0YH4vvOf6e4qC3/Tyixqw/F9lVn6WX30DaVkkrROvibpOctLXdYQQCRvLQRdO
ltY2SStwhRtwEPeFPSPLDRqXL2TW5zZtXQ9I99845i1zEBJ9o5UCtdcHRubHfPtpQVlpYlcL5/lx
QW4LCGm6PxW3FwAciZsh3pThe+5PC/dlNbEQG4z6yDCZ8lTtQ+7XUE537G6YpqFlAYC7ZauSj4u+
/SoR95cn/HYyOTmTs73T7PknPGyx2crEzxMozM727/l7Dv5mRUzqhsYp7FkjjDlTOkEiR1lJ0TAI
xUgJqs71oW0URZtuyqP1EmK6Cqwb6qXJ93Dt47w5ad9C7A7rs/OoZX6RCpZG5kpx3Sch/bUiLFba
4k7Ui/9nrKSZ3UFxtKWpAVwe1QsgBNPMVIc6zI6D/Ai/mV+kBWVawEW+oCCJ+PsT7Rn5e2AbqX2k
hZiTPql7+vD10L0GlV509Tf7O7Pv3ZVbGqFhHw11qc45Jl3z65RgHuzX+cvvVb/vBZjEGftrCZVO
o/1T/TKFQb4wKwZV5wpQn7bD9dYLSS2zzErdn5DeMOVd6NqQ8lnZ5yfQ+u3ynTOG59y/8Vw1rwop
RvLoQHiV7AjqRxj438/I+xcKwRu8SELgjP8zE2fWP1JMRhaH8Ku64h854K7XI83viGDKBxJl8R4x
xSFC/3MmUU6HH+PpdRzOZ7bDq4So7VP6mCmfgM2qJdjXcSyBsSqiAKWtQVlrY8jZ8tRo2kVYGbHg
8SlIfcPt4sWct6VGBXwrHAWBSOp2YPg9JaGN51ehQ9hmoi4ZzNOpFMfP0WYZgyGqgVjQCBayGrig
Kn2ydqbNwox3E79dZ5Z+CBh/5laqwNSQJKQRds5pjA016xV3nP3WX5qtj0RyzvHSdedTa5sWEYFW
GwvVVtWATUdN3m89N/X1sa8/ZnZBC8/zFgrdnYjMX+2xtare4fIkbnjobVVImM0arIfoVZQcKX8I
OTnTPkfwv/e2zhAtIILeml0fOlHnEAMWc9xnzM1MzskvX84B90JENbfgY37qn8QQO/8t/BNlBfcL
frsBqAqs3N/rMVTKKBopyVEbLQ8Vciksvsotu0nrgxRkVfsaseK0uQ9NSTVyJovg/pnnJAb8w9Uo
UtNT7bHRYk2j8VgxG1UJ2Y7u5WJki8lWuafjLxOMxM/vfZ/zJ6sqn424DuMcnYVFVotwlPrmz+kT
hqUhJ8otFwFwFoz9nPekJ606JwYT5uqvG/4uXLt6grj9u+TdekiyrGq00M2Wb3mRGn5TGazSJKNn
tXVR9egi2VP7Igi1NlQMxHI03c/dOZWyOLoNdpaD/hqPEpooin1Rd/O+X7JCi3kiLlcBVy6X7wur
ewmvGufbng285wtKqESca00EHUJyRLCEY7c2lwSHK2XOGovxpuEuMU/qMjDnchvh6gaTdbIZ1PJj
I5wHyMX/gWK7WxzHR4eRlezvWHH5zfdctmRGWA82Vm3iK/IkYbgR5FEoxUGqydsgzNxi/btKH6zu
d18nfccyRL4I6V2BxVnT/FoXfJVpRmWHmzwh1UIbXC7SyMYz9IuSpoOSq4m0w2Ctj9VW70lbkI7m
7fOKFGYrD+yYfn43vnJUhFnjc3K4+ycVXq7mxVexikbVETfbD+NjVABrR0E4A/oze17sBjSoUvim
BjJdthvX6gYAK1tjaoMvdjoQ76bh02/DfJNzPlYELW8zjlpJDWQ98Wl25g72injPzixTT4XSZrRF
Y+WvzsnX0G2XsU/FrIjvU5cVrQuMDH1tahWCXrsbB34MvJLV3amGt4ncon4x7jeJyWBaYrnh+r6x
yylajDL8lh34FrFTC03EA48Gklq9LfakzLoS4EW6khBm5SCMebMywpvZZ6usCTHhxsVPmxmTYqUQ
4OBfD9Bqq+2LHkvonloMlHLAb18pU68XUqRKv94mnQk/Hs/9V5c/Do8BCYH8eDUT0KQxxRzJnitR
X8fTtP+EKW2mKsFKzKTgy+bUAEdyoOLIYStV7qdUDZQgddMUGrqaRfQOQadVZVw2JFhgk+QBRi/M
68Fn1z1yD9XlxbbxcWPkyb8JPj+nhdRXqnmH+uvW88ybcvFyJRgrxB7tsviunRNbVjkNLJQoqazc
v8xeZAa9RNPR5h+5Mqn1nWd5eekYI5bHAxfQC6Ne5BQQo7lz/gM9Apj5hwSqdx5n5+QluazMzLdM
hsb7Jcb6ybAAAFM8FjY8wYPlgoTIju1Mcg3B2UPj8VB1KM+IvxPR86CRGhaprGQN77/0W1JTNeQI
2/z9zD78urle13uxjUIRmBvggifXlo7jKsz7+2J7fUt1qWoZVuA7rmcOwRHqvrTdhCJifoLqU2NT
QK8Q+wOsCrWyXPz1IBcQF3DYBrb1Dm+Zx7r37mvTGF+0tlE7H1HqTxgRHjXdT6KNUfj6tcjEMrk7
Ei3SKHQWqmZMxnWrggR9qRLF3tEgrmV0niU7SQLkWQpw1KhWMEw9AFZ2qOLoeDcuIRkORMvyX4lB
0ifCqA8M4nyk66Ia9mwSX4Xt+jHD0hsVaR5XTxnQ5Dzpk05vRcKdX4Iis6SsMni6Y2Du/QLrUkIT
qEtMe7HHRO1bP4JH8LxY+erX3w+iDr4MAPPsKc7ohwGEDhLpPhKaEpSz1JrR4zWZMoUs4tk4YOtY
6u6kY9GQsAECHoge4hVI63mrhXW4qumx3beCM1qNsOoUJ5Xtveu9iPRPB0d6j+pNh8ty6LjQydO7
xZdadysSe4UuLOa3gdSIXu0XAuB0MaYbByo2k5oeXTfpcLXlrlB56DasrBjiXF53s/Uhj5KucnKr
Lf3nzEd9/iOF6j6fR5R8udZQPgc2VzWTHqKK1FUZTZn9npvqQfn4OsLbF+7LXuC7TgamOe3A48Kb
43afOM7CpPCIe/eXDYbJOacb+NDFxXv/kur0OJopWgUk2uxN5rELTRlVNTwaJVT5HhhaB1pzAzBO
QTydua3cP2k+aciTi51kJwF/neAt6apAurgn3SZRW2WklWtCV5d7UnkvPVXzrjWb3WWZB/Ievkqm
UD5CFDvmLIW6wNLPw9B/lrDAXCJCv4e9VzPPL4a1CX3bTZU8K0MfL/+69WcYK5wAAqIZZ0wf2gGA
hFv0aSuuyTveRXPwLIbRqFQfALXsoR71S7SYpmx6REtYXMQCDQix1yRIAX2IGMwFDV6L6unhNZfm
ovGlsjA9ueD7nSeduGzrddCiZ6gIeqkTMG0W9YUW3kwUkRdU1UsN0w76wxKxMF1ol3V2CuBrpRp5
ojLxDKNgyGCkhSF8jidbdtP7YJTw8+f5Z9y5z3sqhnpEG1n1+ieODMpX4j1cta2OtLZu+fMtXyHM
zNI0EeJqhJKzpjx2HWNw5DBBvvn25YEVZwYnkP6iv6V0XaQDYJfsoXr8+h+iBU+KpJJTXSWuUxuB
ktx9Oo2QSmPftlVd5el9q5NyCIU+XOSiyz4kbTVHcKGcpgkjdOBz8CymS1tPg0HynnLOwSmo80M7
w1kE59V8PPUhZyLjG+7b1pNVBfAbbPjY35xtoU8Dnz2BGCxck+HEv/EDPeitKUfW1Sx997mcheyf
YD2BwmlFddmXjk5/N5kAVWcc7TQh7gb7/EZzE1tRLJsMa1gpeJk6rwTwqEJOJKBYANFMapc8BXHh
BtOmrKcPsydmiAYoG5xOrgBX/EbbuIK4+BnbEiCnAaHNiDcr3lmNfq17gnxL0d12YJTvFBEZuPD7
1RwKCUXTHAUcnUNPPtTb6K/PouJtLEkVkUaR0ZnnZvdPlj14lCfJbZy4//9womsbBGydcWrCKnJW
V2qmlcS8zL9aCx7mrLUtcVQo8s8zOvwL2ToDFK8Xfp1UkTiWB32CHy+1IMyd3fMJb58ZWfC0RReP
0X+c4bIvuBRKf+5q4ZW4rI7jzCZinZkdRAYHYHf/E1xz52A2zmtqeeqy8f2aLv4LCRy9IfNndUx2
bib8IXfpVudGIvTEGClDxTzzeAM/cB/COCdCR6cQtom+QHPKafdY+ZENYqPPrBg7ZT/Ol5eFe2w7
iifflMOlRJZj7DSyKzdNeaYuNOl7ytcDF1XAQe6PNHXYMw87c3zqaHgyAhOnL8cVHnp9sE6wa7XG
MfwSRbg67N7uaCAfjHl1S5wYYvbC7jPDdsDiZzTw9H/lIkVNV68krKx4iY5031mIKjz/IrKDVGCq
InSHwF84kFRgxih/NFv9Ooalt/KOcCRdABvLFWltO6Atu7e37GKxZb423NYMn9ovtOBP0TLMvaqT
NDxXjh8d2hygyFbmfeBq7TSuB1z/Zhvs2+izBxzNyXc7TIBSRL93+Dpi6/DncleX2bZeKqjuKm0b
JInLhVUsG+nUipDsZm92lb2zPIinCTSf0LBxeU1LdrhdiFZ3SfS4rfcYiRShPOFPzo71cHpEtbQf
OJJKtx12RfaI3RqXijXlbu5Ff+Jq4wySrKjEdk68nVLdm2OA7dNc+awvZMHCwYzlqypYzFNLkkCT
8oI4TMUsOMGN+eiHbE/MY5UW2alS61cL2xSFRt6MMYJ5VhQYNvu6ynb4sm3K2kx4VFMgNrWh+zaj
ZaXdNc0VAds4+yia0lCFBFrQU+upgKIvkuwzVt2de4SzAJLWTcnko/r9Fft5Sv0LvBCrTOzSB0yP
+s7PGy5V6xMzht0en8d1P45sPxnYa9QtoqAk7ImgB4vAliTiHa2qnlsxNsqbkHswK4fXTMzcFjTv
inTvSfSqqUryNN2lQ5fL9iuoD8Vh4WBkiP9VXtKnIVbSs3IR73gypZVokL5YkCEGGl+S3/67egi+
YqHB+4y5UtDB/NHz+uDG5MCQCOfyV3UBsN3GTGz1VzF2wN4edSf1/VK16jRXp3lXSWUCKL+YLSYW
gVTuya41uUrQ+ZakA7r+QoM44XSpZ+vjpj+wd1vcq4DTSxEDPIrFBshQm6QBGD45rnzGPLdTqbQ7
CDFBnT1rxfqc0qxZ49749fWYcOpvvu9yBsy7OhbN5/I0jS0Idbe9n1aWiXe1oKyN6XaU3zVSsTj6
EHhrzoVc1o/+PK0m3ie36ZNUulOSwJNvEsZOfSIr+usZt/NSY0eSok/k+JsYlC2+PR33XOlOP1TK
EXCEio5WWv5siGTzr+UZCBwAt/xJuLPyiz+w8GYLw9mO5inYhF/XZ+zzLH5HYBp20LIN+Bu3Yx3l
RcOAVNuBSaLSpKWIeD0rvW+u3VvY093L3p35a2JQYxHKevm1A8CSSZBIsEK0M8/5N+Qs7DnNH/De
my4NKdAhbo1FTRon2vT+VmOJlczgr6aiC7F1i28ERF+6RSiG/vmi1RP6egePvgH6MVHV+VNtnrlE
gDgO5hkthEjhQY6RGXRVlDsygc7PFrQWng9OzSJqEp+L284kYYN+akfUHWycRK0s6pyD01YQNk+3
T09OJjJF3YyeoniDZAxrtOJkex3SyFuACB6tlUB9UKhUnV7mTnR+Btag2DtjizCslx3itsnh2QOX
D/WApzHkQth9hXaNE6J9Ecn7GKWo6L6koqd5h46HykxS8DQOincJE+h5bgbyeAl5HEOFyvlJdbdx
dfoQv5qNga6nm+HEAEvRpviRJNtsHclYcZfmBy0Zr3ojX7nUcNQsieyRFLPCGZBubs/SpZhzFTMF
CQpu/vFAyPKonNVZ5MicnufSWesQjiF+Gl0TnbVfwhy7V+jL8EIpWjqMHsLCLTKmvc8nABgDtwx4
KJ5wkp4UoRHHj+ex6nprG5LvxCn14LoNMYt0AmQD6JLVWtOtof1xNYulupH3qb3rTsH3SixjYzw4
pTbE7xqgCg77Ew4a2sJtOPVVmUXIsFp2p5DpJSAbrRzFtLczo/LZJ3tp9W3jHrGp+A5oeNfdSnZ1
7z+1TzhdbajRN/FnTo54smXadLSXAwJ7v6JUNgL0lQgh6Zb/aj/e3/TpPVzYCPmM4fP6HM/v/bQb
bmqwEyE18PstSdGm8inBQvGSftz3NGifc6V3TCDN+YZWb7bvXS+590MZEG8Gzy5kLX8LaYY35q7g
BRwGlnJcRuJR8WLedrxIUAHHtAluPLUP9lx/ikmk+AFmx5YBHlYUkL2MDq4FEWgMjEId+fbolCJp
9s8QS2q7QF1FhqrHYzPdNgLAI57MxYD9us9yF/FBDQJXrtTlaUflf9ZCB84MBzJ1Mh42zNfk3ynU
PhoekwhENH8oZvPjt42MPadKnSr31v7PHV4pd+IyultqKIF8qmSeZVKqjpmFdcnAAmXSGgmYr1mA
Qw3DQXwWHhXwYc5sGW3JsZXqx2rC28utwCOEX2kKp0xOX97yHkG29HKvE9dBCr88t3R75w4S1QNL
bnqIigBgVbl747FKI9bzdRkzlKOU/V7B9BkpjiTdY7wV8JHtoLhe+xPMYUksUP+2mJGdLdo4THJu
MGBXCDcxTmGrj7cJbsAH5NtK+yjNYob7Rti0xiYshLNQ2gd0ls0gZ5+w0aHTOlOVWSPjK1U5uZZ8
DLZ7kGHC/Qrqb6eEavAHGLqZ09Ekc+LAftGxOVTP1cu8Dc37ItYXUL2MUfBBd+vc7m3lmAaf/BSo
mERwhmhzZ9V0P/ypR3sAN+6p2ug9xMBwQPUhdSCaqARavR8RILiT3ZwhYXZBpqMnGS2Ho1Oz2ucr
mmAwb3YnBvt1mXxmu5wPGDF8y7dW0Gm6LpxyRC5tdvUXr1Rpm89utKeDBSRrvrZhyM4hwHmta6mw
SWygPT7yF2wiz9dSm30KThloJvIih9XRIVNRcSjrOFFZLvjisdO7A0jpo19gv3v6N5RZzmequgnw
rNpDerN9mfcAi7PV3aZvn0dywP/s1tp8yfrT7cb9BhRLfXsBNe2TIEv65l5Tc8DYlXa3K1GyqRCA
BxktaWfmZHkMnGVT+HfukpUITJnZ0z7dn6nJZhYb3sTToWdhKMLySr44ws75r9lkt4ND0l0PtYwM
St53uYzbW4eHo7ykbA0mawS7Pa/zw0WzAkh0dRs71woFXfKfpq4Chdl0a9cEN7sfMHnc5Kqsr6Gi
VkAMvEZ/D23ynW545eYNSfCXobHTOAnsOnB7ozYvBbPZ8zQh0g/NBjvucsG3xp/y/zdYpCJFK3bm
qlfkG7BiHgrcnkDYbM2s4CNtK7398qXezW6aUK3Q7miRZGe4x3UEC8J/U947m6ge3ZxojWBmqNVo
thUrbEUIHNwj1h6l2C3iVU33mCdwADuYveZoFMbGI1EtKHCEpQHhYG/w+kvv+rnufnzyo2xYRKHk
8rYBlw6Lr/JziHkVkJnibLT2w3Uxx+cBuRC0c9kcl7pb4nZgwPIfhUj+Bh7Wf4hMN1lZO+PhjV8H
3LFuwzX/DCL+G3qX5H66JyPgzCVLF2vYKUfMjVSmq0akkO//4vgbwXZCNm78Jq2yHS0S9ginCrBb
uYeVMZ5D2jeIzYbiehUgT4YUlsb9vpp6Ik0wbFdAyAs1a8VpDNeRSikgF2gL3hDibcEYOUJpz2Rt
X7A3sloMromZMzZLwshymem0j+6A3TPVkDSm124bDwz7q85my2YMKsfPhINE7WRJlOYwM6WsSJc7
pKzXOlSvfhdQFzFoqsfCfcPofXNKMsOogBu68v2w1hLXXUfP6dqF21p/52jp+rtCyEVeOC54Xg4X
+J63AjU06CElU5dnGi5EE+iA01HHy/+/xmy22HRNuRflk3vJQKWpa9ClEw41IZLCOZEMBxwqjcGN
yfdFtvNM3bOzX9nrmjJSGoeJC7GgDI0iYLgMIbHsd74rSyWwuMQ2c/31Tvo48nvgbDDRxhXhkBzS
d/D/CVnJqhLkgTNzI118v7i/EFEzvJTEYDmmwSulxB5zlYWlMJj1337Y+tVMkBAtxki0ReAU7MPs
+DqKJEKxrFHA9Kpa1P2OXU2tdDW0GZgn8afvb0slL6d1ylnpKjTDZyFXlSrugYEbEfP9gX5dAhGG
jDQ3YWr9tiwMnz8Rpkv9Ox1Ofl9JfBvJ8UGZ5YGksXykklBArykedMtTY+W0Z86mu8CpXzXvBQYe
rHFzrte+BE53FnHFekZPMZuMJevXaEFhANaCsdkzmcrCILuzb2++gnQGxMdLwXBOWf7d72anlWTc
+wbLLk50mpuHNczNTuQIW0P4TN/vSlh9vqP2d2KPKi0HpGtjJFJ2qUJLD1zMMJRRa4c/IxpKjEXh
RctTH9yIHze5DsoD4Ww8AN8QP6TbT4J8+r0GJ9joMXE9hx+JNimoGCsLNUAmNAucw/7rq/JS0jcw
WiE+VVnd3Bzg/ZyzgmghXJvCn55622kwFrRbqw/7ghR3xqF6kpf/ldTgpgUILHmyg88g/+0v9/8s
qFM6zOdhkX7eHe9KutOZdxIeF5pQ/QeHku9aWU+FCEaPsnUzH0hiISVnBmE9O9R1MlHg7Azvb6q/
fuYLpWK7Uy1S/2GH1g3oCYLeme3gb26nr2Ao/a5o3IT/GougKcmnlGYGgPBGzQjXLplvPAzA+o+b
ZJE6LKAfvV5NdpOZN6lvSveTZm2wwPrWL0Sz/Gj/3vrHi+PPZzvdR0Q2RkSkqfffEKKjVpne8vHX
BLduRAn2Ot6aWu9QYGlgcO6vCKRg9znAW4U5HNnOi21gqlcarLDjmyQp5uW3T7+gZrFmkfLbymLp
vos5iUpVo/inQyy6vVBN5L9XybMt5DMhCYFQKaX0dm0l0+5xH8rgrHkf8Jyie8UTa4UaICgd1G2h
71PNpsMDwyU2UY8gwdUmiecCg9Um6IoXgP9r9dPlJgcOVVQaSGTDAdrSg+fOADejpUfcj2qTlrPk
sd9lW2tdyW5UMTgEzYMS0eBvHLRy22InwXusIGL/odjlRTwBk2kTDYIUBUJUG6EfaHSMmD1sHfX3
UnUSjlkNj/QYP4LirNdD/Ji5fMl7sBkvUaNHRGOKOpwH6LNZOxtgMWy8mRZWK91ioCEAw1awQuJ4
ci/DcqY5Sa83Tv8Plf3UVes/R4uQvmghkMK1HewTacJNZE+tl5jVLeU0xORJiduu7GVKlb9pUFXn
8u3b//GDY+FCraeknIsYj3FatRMqhLt6V1W5uCO/ZSog7be1vLLXzEPhNKrpr3ZYQiw+Xmq5bf84
VgndSCXEszaNJQ9VAlk07eDFeGvJ8xRjyeBJJnGbV4yQoOWLlEKobAdF7MHrd/oMhmFhaL0YN2p6
TZHGH5iEoyCO7zxs5au5+mmMZaSd75E+7cwIll9lx/30EILBavS7j2IefJ26ZK1VtUQc1+cwRKpD
oSBfsZTYKYm6jjNdLCNASKZRXwEHoCME2g1ZiarVH4PYjwCeHVSYLJz2zGuzfUX5pwo/6if5+bBK
/nEWvghqI2xgFc8BDomcOJRXXY7uGqQC4dflMbN6pGW579QoNrW8sPQkjaaJ5yqctnzEPrYAvHXD
d/wzvxL68Js7ULk8MgdzVltoxhhWHoYwhuFDMIw5oSnre7a+S6UzcYYH1ode6TvciJ3IzM0H5Orh
yFCdl1ADDGG0FYON4GUGat1o233w1L5ZRv/tBd8ejgkTLefbD5Hq0BuUeEJzvpKIQG+TuvzQMCK/
xrjXoSbrqQFrWzgFHsGYTZtPQVMfY6P1gOcGNs4hbnoKZ5kAVhOYqrIrCD6HRBGJSPQikOKCzsjn
5SXtmQIKUTuAw2PlY+8bexOqLigamKFDBnTGdx5nQSdXHVKU/ps+VYCILsvEWaePQNIHYCA2KVoz
EiJLdSDlbfH+bBTgZrvPDMItelNxQXr7HQdJQudWNfBsKtxBoRR9BVv041LDkrSjsr7qFYcvqaDs
YkMoXTrPC8mYpplJk84eqimWxVpH84Ljd1BpHm38P81lymFHudxEryYQwe4v+p94jQqTsHv5p/8V
LY9X8gJJWhq0JmbGH+A/YRlJbiBLsBq3eYiSdPQQxQ1iLZ4NJbtsoIUusl8XYK3DQSEv/T/NzNYJ
cnSJl1YQ8y+DkEB84W6m0I894uotZJ3Hxoedx0Vba5sUqSG1vCVHQOZO8sGvvltZ9zcMrw6JfCMF
6O5q3AWag9HXbJCl+aED+khOmRBRV1LyNhLW7B8+mfhacapxLy8dcxMLeaEUsRexR6s4UDWeLQzF
40MyYJOqYJUax9Eu7FrJkiDLTMFgDIewUcY3G1hmbXPmPHMN0TtzIcwRY62GngiUq0LOtXhoigCa
vFZ+A242IH9j/+ItZ/bVTbT0KrER2pzyz+h/aHIj45A1Le1m/BVxxRtBP+e6LEvcUPBuMeIA5ezu
ZDUhMcflJqsi8UTXqMkSEnYGyYHmaY8c/GO8Qwlw1Jp30NnvHYFtGGvUXySJ3sE+HqYF6IMSbqiK
Lrh2cloZSleEQyQI3xbM+uu5dgTxVN0yFMv9qomUk3Px3SSqJ9BwiLk4w2zWdZkLEzYp/dEw3w52
/goMAWfZN5xEIyY/z+8vwS45I4K8puIE/uDL55Mnw7/ERWNJSpgXMIA1IkLH0Yys7BfId8hdj5B7
NON//5QcIN9bsszayB6sVJLofEOvAZPneLS1GLM7WBVkBEAxw5qDARqe2iViM7/w9GNwFcVcdYX0
5ZU0J+hJK36T64eWU3U2muCVQfAdgnodVhVs+ul4PfNbW623ZYSTsCt6dJHBKLnCe16mX9PhKVue
kiehnsD3qAlVQARmNp8Ad6iSYQP63TGJwX2YzhUHpuxJJANt4uxC5h2MZe4lr81VqVTHvL8PXy5L
7Kav9dRaOlkPHEcaaRlptbZ2/itO3oeaanCI9J+hgwnqD2ticDCyF5j1n/x8PsM0bCV58UZ/PSfE
MXQU1o8vBbn7L4XKofB2UVI4dmSccTc6++L35tyNxbTulLB3oUPZSRIVLWLdaI9+0mlVGUVT1S6J
s6h0V6L0QtxVW8DHJiJPTjjgonjm0ZNvJN11vNM5/lUXGy7Ql0NxvHdGBdy4bYGCornXPSVdUftq
Pe3BWpr+znSDFGRoWG0iWyNrVA2ojrH1wATMYyk8Oah/WBYLuwEbDR0yBMxWOOXqCMx90RsMH+ZP
NnbjuAQAvphm5v6zlVdCYJVnIH+ZshDWAHQKuX2v+f3tJrQoy8nSlJCQ5NpRD4vlRbHOgka8AkZf
vjjePVLUSxkDqfWwdys5Cb8eYOvy2wAGhgHiINKKLmFZOPDrfVjm9ThhAQSki00JCuti2gRAmHds
6yY3yJA/bs1vdpXaXED5BrsxPVM2KB3U/u5PvtL/CP6YXf/WKxepOr+bJcpnyVhoIR9A1QVXY/xJ
MCjqWRj/de5cyEHs6JoieD9oMNK4lrUpHP/wwfp1R40zChPsGd+nZJJplkU2RvRJeSWvgCHjMCW2
1Fp92HtYJ2mohfLao9BxVrRoxXgdKTntCL799jhtoRh2dsd5t3GI3xh4LY/gldZBt3GQaKYP6P9R
b4jkVcv7pCnQ2/qpAjB2/hn3UCaiAmX56/5W9TXuoEjYA97uhhwnBy5GwTSXC5HJGvOdpZTd0iON
rqRlK5GqVn0FS0OzmZ2VsRA6rupIoMhHhoSIO8wtYcE7ouFXx5PPw8NJBYUvNWsgqIJHOri5lAfv
OQ9Jju35NjgV3B4/sDCHrieHrSx9qli/yjETHzJBAR9WpIOrQkZTQb0ldxT27M8pPNB2QtKQyZg4
3kjHndayKJ3TlGL1S4XJLlng4dwmGphsWDUs1QGdM3VKnd5f3QGoYO4R2tTS8yCoEFhoBwF7aKo1
3Dnjj9cwKhGy5tbGkeZtvOnn7nSeVZu2O8QjqlF+6oqeItLbP2+8Bytc3tiCkmKbRF7qvoqhuuDL
7riKFB8OyIbn+LeesVwDBue5qZ/AL7pjAZaCSdegLARn9CSPKhGQBegYvC27gHH7jXngiqa50WYU
LIOsfB/bV3Kp6oclRyrxaKmJz8WrDDmNN0n9sZWaiU+uClfIQVnCtw0kqbl3DChNTdaD/Cw5Us5Q
O891sTkLrG3BvoLIH4SX20nGOQhPy0D6sFb65A0ZKxJM8vgjzk/SGeV4KXWj9DZynw+ZilEIk2RW
peR0XnnhaNzdIPIiy9h0DVhx/+Q5qiEWYfFPeJ5hYPvczdYrWQPOF+go76Ku3LAuwHeIWaxfo8c3
eihDFsFbHc+B9T2dSDGNPTPYH29qiMlm38K9SK4Am+awUyOl9kUJpiuDDDqndqqSJDUmaCuUIRd7
Shl+/RMQgdkDbpLhQ8x8IjcF7d8AyRIIFocok3hgPOUOi+CwZo4O01sGO3xR06MI3MNdUBdryQYR
m8flljo0hu2Zd7hZdnltBxABvdDFpEDl7LdwF0U3ka65BQkisULtZgglTE543ZKpm7ZDcjgeEQur
nAPyn85DHJo44SEQvPKo251eeYxp4d6eQsTA58wyQgxWgrDi7i9TK0n2w5xGNd7+AG7Er/0BSQEm
dQ4Xnkcs0zy9xD/BW4jtKbtymMDRKHb6lc4adq6cDlDkqQ7nMw0i7G/ACtR9vaO4hAMkJE5GR2A+
c+dJhbR95mzpa6vx9uW880FaXjbD0EovSGHXs7i6DT86fsPeoceQGTZUT+zdkMoaufWX8l5g6Dtl
6/hETknPx6SA+XVlKvnzpYkrmxNAzF/nokP3QqeCfi7OPiuy2QXfNJV17phoJ6JWx7l445RmhVzD
QmTlO5ya35cxnhn1+WNSXBDu7+RLUWgvM4e1PaSdTyPYP3TL2cbfVBBWvgcGOKfd/VUNXc4u5rzE
ElVXSA5LM7OkQVEHiVojc++Dj/Wl2BL1B9rOqoQk6X1OBkFqj9vUTO8/uySiwHAOUgKSZNu+Oiqf
5BfcSmZOHUf3MqsPpIBcRDfekP25bVawi7zTnvG+l0ywgYwcuy1qLMcR1SyQfdEkW7CmNkGmoCHN
E6w6UGmSpq8lThzRQdtE1Sdum7MAar2poA/WnkKFdggLvaaaE94VaolgeYuGRTGo7j/66DW2hi6o
+UOzm2s7ommrmZ/9AWdUi1HYTnNdtW4t2YL+p4wZ8Ku7PA7cVi2h1fRCvWTUr1qjVpDzKNE8L2Y7
snzSVU8a9+RTmTC5cEMlPt+SdayGnkqm2puiPUFAeNwbcVdMTAuSLJeXibCKd2uv9nJhmpUQ5jJE
yqWCbQqM6Hu/rAfeILt+7zFyV8++WoWbQChjT+MyAsw+/W/ekiPidBGXqBS45Si6EWhJ0cDLXkn5
I6fXDy2tm6L+J5sodYorQ59PsfbvAVuvrOb23LLv3Nv3IlyX/6jCec5SwJG6TwBDsNR4Ly7/KN0t
20vcz4fCah7VZZIUnnpKk5QjGWMC0sss/nRq6EE27GYlhoK9WLydzLweCPVpaK5uknsYtFNYmqcI
F6qCki9qV90ffnpi24/J3w8dKWB/Dg22GJQquPDMO1kpaS4rpI3d4PYgWZQRYQuAViYn+psj1XLm
MigPSQ4jpHSLq01FX2cDhj4vsjKMBByDkJz76Ht4tfnFnO1uLETGUkE0qDhI75ZEeLPSHLSEUL5O
ZPm5a+A3RMxs9syCm5IgapaR7M3L75Hr4+Vm2YdcyagwnD7mS+9M3N6Hu4LEZXIPViPnLk6c0VTk
iWLTHE/pRb/U+U027z5T1jQZKzfV5cubXayN8ebL3b+4Qz0+YpSnYDUeZk1KLSOLlfR7iy/3bUSy
5sdDZaRkoLOeG5oA7QNas4huNmX0Y+tAe2HkGvj/C8/d5Ao7sAtyVzp/uG2YOgeYNTwhd1K/XGqZ
6G5mwcz9st0uMuFZwRks7IzQe8zUXI1Y1h0emsIkQEeOOgCmK/WARM56oRqajJaXcD16Qj4dm67X
H6hjmVCXYN9bu+W2m1tRyxyRO7rlp9HL3HKVN7gbMLZJiXft4bBQ9XGANsVq3f/NaLr0WPKzOzsL
4hVG0h8hms2/ljF7PXayk//1+U1WTtAXcH/0nYwVUhc9nvZvANXv5F9+nABu6hPv6j4KlvVm5VIv
R0hJduHc5ANLJi65v7iLW9LgIxm/dVgIs7YaH0ME8imLIdqyu0ai2soqh4okUnscVYxOl3Yz+VeX
EosUvahTEar1fXTXI1XaLgLHezk5ev8h1L5ZIsLtL/PmGy4tBgXoEC4DOJ9wZg4/+Adt24t/pT/d
mYY4Bysp3W97KZM0X1xK8AK6EYpQWfKVS0YymTg7h+80i34CB16YrX9KKESfTzxV84dAKbfYaZkw
1FY/mPihWlqm+Guu6D9e4NargavKas3AMKCUWJzkqKtPRtB11+iNoeZPXTKMMAiBtuc1EfTtfB80
67XebUlHzzSKL1fIKhnINmRvFpHkuxj5Xz89gwHhgLBdgAsKQwVNnoS2/n9vWcp1llnPoIFyzta9
1TVvIkcsWL+iJrpht5+rV1Ecv5Mn3pV/YkIGYfwMZmG8JxkPXHX6U39AY4Ce46Z8X91Gq1sh95FN
JnE/dhyQhS6IGhmtW5Wn27NahpDEfUo6tNW5swg2f67CG8XLKkAzJzgryx+nfZP1uRwQCQYKVixM
ulflydnjGUjA2/L4+VduGCsCM0++cBe472b99ATuQ2Sk07QcEjFnd/3JUwtFIGmp19W98pMWiKBK
Ys7Fh2iEg8ZNmJagAjKLmnNzau/z8WKQHcNsv14ugx0eVku/rse0ojpldXCpvHvabzDRtoPNXN6X
zE5Qqsx5PSvNys2rN0FCX1vDRGjOMteZI5m0/aSjH4Hfu3ZBYxl/2stT9zD9f868nopFpILoqO9c
EnPOerADfI1oG4REmj76s3RuA9KFD0bbBsYh1nIRyTZiE2e2STwcLo65O+tk2lSTIO8NDmuN2Xoq
QxzrMxPeBsuHmO2jBbWsMyByvxvyHnaPKqQqbRsD2BPTEsiuUBZMpPgxQq+TZYce8ECWsF+P+Ndm
PqSOO9kr2crD0tGz+kWOlMpB0BE0rjvX8ixK1qhuV/V7+GT1Cvf2Mt7qHQuY5DDrFR2BVZ7zGkJI
sVspVrijGClo646FYwIt0+RUD7ZTU39TUo56p/S4jiQIHoiEYItva6iBvNyCPsqgZAHtQ3sKexIz
t83GPRZb/DGSxn9lnXExuXq33I7pb6/UZzFgC1RVUpbSA6HoFATUkA5zDPnTxbyQQALQH1ohANqs
t5l1vpc4sBSEIu0q1UfREwWWXxs4GGHHiMzHY6HXkvyw6T/+EfCeLO7jLuXZos4ARhO/zXFNfVpZ
VIxnT0rneCrORvxEbeL6jxMeC60XZwgfs5Yqh+bsciOJA6/mTH8wCb3DhvJhEGQkz9crcZyXaSMw
vCRcWRMd1WSRoztYrKNyJwe+UE37Nv4v/dSaC1yr5QoijqEINlwK5ERQQMKJ7HEfchLWAJuztCvk
MXCOud3P7yc/Y2fgdUljif4yq3tC3ZE7uA5HuA00TP8Xp2VEANfTicV0LbUptscTit/TgwBF1Fmo
0mDwTI2VwF9xyyY+xK1mBd4unAlkD4naUt+nAcjGyFQPqFamGaBNnpiP2b8qGsfzWT0JMqeXTAGG
1LlBrtMr+vLjplalt5pu5OdK9K7SVfSiZOU9k0MvUs7/AK0yAIozzlCuyGS0/m+Rasm4wEnauVYg
H8Ndda/aoUP/VAyYu531DjmTvZK8Yge0MBwJdK3a3ORnOTHukHjD7JSJW2lGCGKjVH+6kDPlNgsH
CJsCCz+9JO5jyyu1Hl6AJXK05RilbeuP4eUSKtAiFQeNt/U6p0BI33kOsE79zax5Iw9/Cn6988cA
rgrht2C8fwkZAPgq4DbyaT2Tn1wCIRu4gK8kfVCIT2y5hl6sIpIs05ilpIkQaBLEWLH8GGu1DnIC
Vd9218wvVny6CXjYMGZoLJn3x+/cJqDB/5HFz3cNsNnu55j/7PWULwbnm++mHneRumq9sfHbebFt
T38pnd4P3Stwh4KosxsxoZ1XodiKkdfZ/OfOVe4hb9NKLAdtJEYwwicueV8PqAOJOCDjSllfS+aO
FfU4WQEcbO/phw4rAeaaBGRt4YVRktpAqnx5aBIe7dck/ynAiFsbOPywTsRTJrTyIJJhImHEWY5P
4sxYEodrTBioo548gJnRPzIPMK6g2zA72gmlFAwjEkfzNE2FGn888LDcdsPfGohkhkyVGkwNLIPd
TwPB3YgJYpj85CDrHtI5f9XOhGsR0fIAoFFlbyj2gTugkudcpPdiu6cc2EXAhti+xzLU+veqFIBv
PtOKwkCaNybcoe8kSHb6wCw5L4trl6ORijaAkrbhxQ3v5xxAd8BLZYOLR0386PL1d1BWclLRNHAA
LfdPeLxKUXAhA0FTydzQsXwC8zp2uAcRcueqpHx+KGfb3RWqBX/AFaNALgDkSKA7VO4TzkT1doXS
LvWw6nbLqy8BwGWkl9sjtgH3S4+EogrmsAOLRwTBPcuPDG1+xF+IxH0mtwHuUl793ImOAI5nfTIg
M9rDJTlNraRTDRuB1aAulxr/Ou+ZRsnxrXs6cXsX9fxlSjPtzAsAeo4OR16LaZT808YKbaTuWUKM
tm+sHOm6wNkDdaF1+TxYM5seLHzeORSMQdRIGWA0TUCWMbjY6AjFgpPaDdcNlNxkDmL+NCCQcHFP
RiACXXF2l3P0Homu4hSrl8wl1N9LAyXGXfZPH7Xr0L6ji9zhdcW1Zk2rD6UOi05WDCtKsCJ9WBam
97piGbuRqYjlWHeSeTpvV7iDzDeshMqRcuNg6hahpqNXjVE85o1UKQVsw32YyTfmLxLVrBES0+EW
JKxhnrdE2Cju9kdm5AhrMOov+9mqknMIY+vTDlR+NHqt0TcE9COMpJPtou2qBOvEdbd7FsbK/F+q
3anbaaC2PJODcRmqwKmk/FMXdg2JdtlN33BTX5Kh22YbycXgTtsuRpX5qdnKSOyocsbGWhASFJQr
1HiBxyNCCnancNvCQ/rrNAtmrBQFDlOLUgLlU16stk7RZHeFSId4+CDCGWcq7uWN0FggesUbV5r5
X4uSNUUpqxZ8n7hnDnIuUzAGfoXLpG6JZ168df2rpoH24iwLxFmtm+cT6jG7CtozaMVt41PXYKnw
igWZwxOKxPhBTXhqLKJboLqE1yq2ga+jbGCeOvMnRAjgzMUht8CGwfdClP4ewtPCR84wy5cXIkO9
K66HdMuK6P7413yMzWzGIr55XUW+E8m0VUEnXXxSZoOpcF4ugxAFOOWLzT8TfZh+/I0/zw+qL7nF
YjFG3Ka4hreo6fFH8mVVrWzNPKGSfbaXte9vVKjxFFNcHLahKmZhCrRDNGqdVyYdsw2g1G6psx/u
P80Ikn+f1q2lqJULYDJHruwqjqqSxb+IgioD+WroQ8ey9tF5dHSDXtwieWK3Je+e3UVsmd390BYU
0ejcZRodx1zwQUA4N2SUrbg2Vuuuhp7d3K0B28VYgM4oYwYrmCMTduttf/2KbgUABPjXCjx/rhoW
gxo3FgQocO53Y7PkQ/c+aPncQEyf9jety2rDv9PrgqXiFT1xHiwvZo2ibkONkfVFktWWUPVmK9Q/
O/XorvfRuHJQ667BB6ipqHgLI9LVhiPky/cWZAhsz6fseK0IoSpC6m2GobuW2zNJQlcsyrwivk0q
vTsyJgA+htbsdbwj4+r1oMi5J2h4wo3/Grt6ugCo8rpxh8gD3UfbF2pScNO16Jy1obp5rQ9hBoVh
EueLnRYRLC2R5BoxnlI2Csbn6pBb67+IQt2Aq3hCxAkjaRIeTupQ3GJzqFk0bGG4bxxtCo+Ue1e0
GQSYsusTmbeDDMTODYvkcpz+BRbstvB/LpOzmFzyojXzco/PlgDcc+thXgnavId/cAg+3zlUXC5+
w8tcmA8FXY6owpSGApQbA85x63Z3FupXN5bHXwTFFlJvDLyX1QcPbsJ1f480AIY922BT94fwB3UZ
Sa0hww1qCGzU1edsRovHu4tTs4kc81NlfN/QnvlXCRGSyTZ3HQnSmt4iS6IBVEecR3pagmByBAnO
pwydnDH3E6HRnqxjOgLLnqPrha0ixsl/e/vHWyvEaRtMEYGWtYA1b16bNosGS0IDbVkMe90+INm7
ibzJpudpvwjTlxQTOXy7ueXcSg0maUvjC4RzBMCetVAf01SC2XaGuaTWpC7O8PObqZTQVW/oa2cF
J7rBDTs6UJ9VB9slKNPbcV9XxJCogV0s+3+uLiRGOMN/dn9NlyRsBWu31+U3oDjtq9Odh98GSnik
RPCAjYMrVwjTlmCkvBcCRXDFCUypyCqHBsVO7Dit6kAy/WJM6ryWYto0JWawpb9RU4/wMCDoEKpE
qKoN1UdJ5V+6kDi2uA7yJuvGESYpd3fRWfYG8ZGYgHNTozFV6RKqPomjOBPAtjfbtLidyV/y1u/7
kdDSjfVpZrKAT1uIf8MoiXoEo2J6NeBSqbQHFQc5XGP/jwXOiyZr+NlQcPoYiinVvAa3HZtLIqeB
2CzSepM7GJLNdfGZqAD805hqwPatDEz/tMB/X9meeQy00LZc2pt2/VXOGH9XInlzy7+NAZJk6PSk
miv4eMtWL+gjqQDTZHSg2h9ryuEodwzmC0Ld7Les7epc9nMPRGBS1NHl/d5NKIHggum0UrGPXb5H
+MDeoiBse6AITrJXQMx9vraTUdwMZbeyvkFdmn6tnFkezWFufzE9QGZ2lTIU0FvTUdS8lf5MejKc
g1PmHVR2xru/EymjVgWYPRSlDUoV9MtF17hm4KYARCq7EHJFypisWUFUPfh6NlHgaCHLU22iZwMa
alSUCBFyhCT/kU4WQ83FLNsmSNF1XukdoHiZYRv1kDJIXoQngzkdC2dFxLW6GlIWpvXBhq/6NEyH
H0JAix/zr3Fyt0h4SU/YqCb8WWyfSmWxY978N471FKYPwwRfRLVefnYOpc5wch4JQ5OChdkz49AI
HO7bALUWClK1RJudqNx0a964MkJ/duzCRqyOqbo3Pgr3QrAZF6tojou6WJ/239AnwrONIurwHPPy
5Zm+B6Iotd2rWBzuNvPPk2AgIQDPIEXb4MX9YGde+kxgSBaiEW9VWzaQg8arb0Qdx6sResbD2Srt
r1CU5jYxwNzLAVmLrq+VdxIkGXBGSIGMASIFo985Ir7yDiX2QPwodGU6s4oQsDdhZ808Nf5IILvw
h9EMBq5hwkVzvD5prSOsyx6B33VcVzX+jup+aDplSVezzN5gGASMjaMqUy5BPyt+DEjrkjBbhRvR
51GJDra+hsZwWG4/cpdivn35knwIiejeAh9tWnX3iPWGHv4uTDn+sl1NDvELjYbNQhcUNNLP/jfG
8EHGDtd6wveT3Wd43jaXei4OyunpMYEzcxPdlX6EqOPalOxXMXbvKbFH4GlwKo0FUr1MwxlU5kd7
a6I/VBd10NhisKZru2eEwToRKoohk+sEWkwAIf8uy9FNghFE6RnTYG4/TvwtcFMEQEfBec8hK+Ht
xKZQ5/YFx8AgWMfNf06NNZ9HYeKhqXswkugdm7e1apcOsfaGPbecMsH2E6SIShmo1owVJ/yiaXWV
wcVnIbYayxQ2Xt3B4jI9QmyJZgd3dPKUflSaGbR59kQ1tGt8G6lcpp02UsMLnTRsAWRVbeuI1b24
t2pXaiObst89IeMNTTwVYoZeTP3ATkTZyIR29b6lp+5ck+WLKg4ypsFSECHDakeAZmc+r7G4MP89
0de/Qj9Z9wnC/bAYLb8ucCOiIgZ2a6b07FfJIA1MOpoFKGqhZNmP/4QLdBVJveTrXeGaE6He9AGQ
NfRd7KfHs1Q593xx/Knty7+O+XRbAYvRO5VoDAsCXkG1ce4RNyEP9CLThJc6p386XPlPOWG/XDfn
hSECH04ge+aWr4bn8rBpR0UC4GGJnEOy9iuRoKZcMcwdF3vx+2NKSaakZVJWS+dtOrPeeCT2gag6
dhn9eCnfurfdHGUpcp4E114vCmIfQyMoG0IkqCgLgbS2mIKE2ujYeXFa64KeT+IssfZ7gfW8A0iL
pY8JI/hPBkyPOdCblIf53UxAzEy1FS6zsCTs0hATQP1ONe1gZhihufCbcLvAEsmIwuIFz+/SOIf2
anNW9qfv3EKsuhoFo0vZipZ5jsKmFDlwJ8GjFDTLFrjCuMSJN1hy3yaAmOn6y+mszQLgQzyliXm3
24HR+t1YVZnuD9FHisQsNFHgjlg0B7ktgft4d51IRFmPOzoECs5cafDQigPDsVqDf16ivRUJNRYZ
QHw6K6LIF9lKBwKMxQwVvaKpU8mwfr7mJff/d2N/LYJulcusgnFD3RC6mtHnMBZi6Jkrd09ANmMu
dJpxilwQlDvzKIUspb5tW3yX+/ZGRRLdskSt765KABqcH98Rs/wNmYlhDPnYZuKLxqjUUCypF7+M
wWS4tfXuuCGvl7oH0bozu/z0OPVfWEGu2jMMVv+E7tZ7L9vIxK92WqoCL9tCeckaPgfxkSDSWLBy
5yd+16kd7C6rA9f+IBuAzINmWMUJHyDNxudRL8JHgMVENAjtWyNuzI6WXHjGWmfo8FXItZf957G+
3wRi9NrK01iPVLBfDn3mo5MUIOf8TWkPRtCLHe3Lf3EtdtndFc6DBxyYHT9Rye36MbDx1I1MK2wb
qJ5PDhsyroL5UkpRLvrWsJeXQ3rS+4tr7zGrMIZT2IehLdyZJuL41J2R6th/G5Td7NupazRaZEv+
hMRIsFwOpljUQ5ttWogjDyW5NgxG4+bz56o2TXIF6ay2qwWbUGmk6YuZm1fuit9QVnsd9hPMFpk3
xvcnrO2fjqM73M1a+fuf01nsc0+ZRekR1nV7KYL0JRQnujl9QCSbsL5psLKXgfMV83RjR4mrtJUb
/0vHY3HFgKiWYz/PB89nPOzSYbgRg2/PgpcBnkMOSu693Vf7ThuYeC63J7E1UO6iDm9UVM784Elw
RtzfCim6cBPJjTq78S93ZnXpWjxSojJqBxTYMZvHRKPcZRjw5B+TKjIHh92NbCJsA+JjfQGKo0Wn
rCbI63RUl5ZENXvysF/1k4PFQRXSGPb+iBaHGISGeBZf0WiyM+8rESutHiPxcAhTKbfxKruwxk9F
vd5ME89TIN0x8h7EH3GYka1FRVS/8Vdgeez9Cartf0d8BInGcOaM18TeiNTeqWA+3fuMbw1cxxLi
roCgy6xamTkUVIH16xAyf5RnLbTV8exvmrrrvPciWOxa/dqKRxYEHeHKRUitMo64XD5kEslpz/J9
GZk0pEYAKYBLhSDfi0Ll6p9M8CvP2ToLYpo2F9cWKHRCJ0HSf+CJ5nJv5I1HMU2WC11g4wcSL2uF
Od9h3TRJAeaWvT/YjYUDWc6N17v3kuS+CAQWL9xHazvZitiphyFTacJ7hhrBGPGR1xI5lB9xWqGe
kwyzA1gMpoYyrNAe2pIc/KGGv6jrMqyqMEg3cjcA9vUrDpVoiGvyAevS/kPu1OxnT+35dDE+Xrxg
BZ/o+1o8fhulvYEZiOZJ29q4mLBAq52D6uif71emOyThHwLXgs1R21omXdf7kOxMaljqbVlozL8+
izrGyDQJ7/B0Q5xh5VdN7jOg3BtKWtLRNMxG4qNnMcoWmDHEoWLbcSCgUT/qRUZ+qsGOZYFxpAVF
0UGvHSMhwijM+to5SFVVNPOSOh9/D9/T4NxqwzEKU98arZTMsXCYReKWZHdhcVR+vgI0IyUEYAeU
QjYhXgZMhHB5z0nkrcc51QdmnC7H+iH8/Coi5JRKVWaMTUjPDDq7G12xCcYiugr65LEG5POvAn74
LLVD+5pn0ibXXxDeLMRtefiMfKldJHEtLYl0PMU+kQgQ0gQwQ2I6UeR5eMTqAHftaYcaPjGR8P3V
4PIjNWW9unPAk2DQnNi7nYUFKiDATn3bshBHkhrQpwB21Zh19JU8FOKfVFa8ZUqBgozQO60UNO1R
cxgim8+5xi9RjAtKwAV0ZuMsuLwiEZx6ohIuO7ADJDZJqE7ENa3eFBtyzXsQuLsNKQs2A69YVMew
CC3KI5B8CzeYC9NpkSQNjkD50J913tSeDYDRSee1Lwyc/bQWprIbVG7bolCRI+52q7uUY1XX6BoX
4arqFpTypZu/N+wJ6YxSMENOyKDP/38npAWK846UV7gquLU0Ld002ZUfH40+l/xWspZIXQlamFJX
n0SMWhJ/2foWGRqq/QcH7It9KfdRMdeOKN0PoeNFJlPYLyIL7+e2gpC+zaepsbqr77PN6R5IkmvS
F7uYGpayV0eLJ/ZRwkh5sinzOnxmSFhDGxwYUKkw72ZvRW6LRZ+LLU2ITP/T+XU1/7n/QPTcH0FA
GF0S7HlBd7eXW7hdOhnJhRuF/LZsIn3HFX2F9D350he0yYKri0t3PnLFs0gOfutwblm/BS48KZck
nVou0rk3AiP4UocZyCYV9TfGtm3WPkb7EKw7H7xVyOFyvD0EW3A1B56FhaJInXusgX1FkaYoA5nB
kFU/qrDAly4RuOClam+1NK48YzOyKH0kXNqAE+EAp9VVeygX6raI59VWZX6a8Ho9Lorp2j9FITV9
Rnju/M7Y5T0OXMp+cnM26VKAfAmyrGliuewCUo6Zebho9v3lJDKsbFnWOGyMpiPk/I/HSynpKiCQ
e1c9BMZFZ0opTzzQEmBBoNKhNyj+l/qNhmKCV/8qV4b7OmqmGfvDRpePsOS3C8jsa7FNnuAyxQb2
+LuaMX50uAB1Uoor893q9Ddmwc43HaPh+1KRM8zWLaQ0hyvwkvgWKqLSv6jzut5GBYC+Bn6igmiF
va9lsJEr5oDcwf8TOvPuyByV44+lgMtOztN2fMmQBCpSXEFLYMnSUJiTIaS5rcMWE/EQ9WoG3AaQ
FPxAd004sLZ6waOrE8ZI7dU2MAbuc9wFi2p0hFP0ky/ZkwLZFjj4n7jnglAHzLLXfIC+nHnIqsNT
ybrbS8BIZC4ByoA32ppuKu0SXchSkbLxSeS+8a1UuelLMvQplvjziBRqgJIrcglnRg4dqEVFMwZM
F7V8OjlMsaCGKIxETQ9CTbrSBU1LV2EinRgQFp+Cy9nJD83Lglcbx3SBntSApS7/Q1RvHYxCfBSe
ouqdCzHRwNYJPXLUNOwKol2DuTD3M1jM7UODNDl/S1xJ5TsqRHTG2lA9KanjBym869gLbOpTv8Mv
MtXhio7UzcbPu01Fis0bPa9/pkfhROJoEtBr3Zs3eypxniJx4ulwulrE5HGJ7oiSg0rR1sh2tFEs
siCn3hCvptbYai/QGhmt8dIREa3eW+b5rfDJ9NybAQN2/oatOeDSV75Bvh9kL+b6tx9VTKpp0cTi
MKQ1zOzwexK3tSwzVpNKPl9teoL1C+zMoxtHuukNhrzJfnBBqbKH6q9ZWLbV7Mj6Wfx8jxAhOjQt
OP5dpQolbftahAlJMY7wqiB0c1/9+SrC3QbqhNb8JiETor6+9UuFzkjw+tceR2y8Wvygjzm0Wr2e
W6P0aMxfqD7ZI/hCZzbX0fUwIH/mQAhrKat9lesdwJm+6pPpRzeM2wtKHivW3o9FMvfA1QZNr1RL
n0GZaSeWVZpja2QWzsSUsBaUTH74uoKDokDUl8jLH1IX0/1V2VIFLuwRxQx6yqon+vVBQLL+99No
t1O262NZYknA9zYpdAnsHStLj3XuL7l1P4MFFpHf7fDeQD6WYcyvNRe1jI8hQffzVTU2dWVB7hfh
ktXlOc6wsBDd2IG2ZXjOr41vJAntKaSI1yjzoZiHwlJX4Vy2dhjVwARBpBCfWEvn33n7Q+YVOOT7
T+YJnh9b1DDabFoCNzYVnIOk33isf07NX7k0YM+LMNboEiib+zRCzXo9WkXfARMm4i2nHdtt8jVR
QTRjnm2ZQ0z2SNOs3EmzOYn8CHt9slTfIGEuko/NwP4C4BTcgwg6rTRNgKodKnlL9NKqsebvPtMf
UoU1lwKq4Pu2aGrwfFgsbr2IeAvuIFopIq1njVG9739EMx82u/yz3N5u+jt1aXZwOLMmFncEoh6b
pzh1biTz1m1CCX+SltLZv08hx/E/uf0dc8gLW+MSsFYRFsF/xL47zc7ispLOYNHPNfoSMUesU99U
xTZwlbodbHOq6QWtg0BbhIs/3gWsVgXYiN4oKlvWbdd8Nt7roj7tp+5Z54uF/F9E9EVJJJblBZHQ
iFJxponRHMpqU/gXve7JEbBMopEnuzQ8hf5qcoxorYXbEUPMAnlm4n7GarlosUD6AvmAEUAwMCxJ
MUg5qXTLiLz0HvaFP6WHNjipkZFNCD2swGAebPVxt/q2tKs9f1O5vxX0MQIGu9a/C93rZ/AHZ2Tm
73BcYVQUSNjtpSX4SVSCfId5ojT7Qu7s6sO4LkQCbOA1zZujlpS0GkvTAa8ert1zwup/NuzXVrjc
dQV9PWGRCDOCK1VdCkigo/q64OZNnWus0hVOT/Stmqq+2mgHp6RuULAVHkjd69vY3ITX5IzCtSu2
CCjwHhjD5RITrMpoOpMWnsIXpcXLaZyvs7cfxhmy8Wi23ayTUemaVZgHSl/wTRFP2iDx8E7U1Ach
iiEisAcc31LtQ5r+4ErQXtR3WjrYrc/ASWIjc1sUrioFy8g9ElfyaQqMO25lbwrdU38fpLt1L9ae
oADxiYE27tm5Y0zh4JUTgVnI62u9Da+zxsLbv0NyYtz3cIcSzNnU3VXAoEFFxODjpa45TOS92Br2
yR/rtfYH5aJyZOnaFoQTCKpr/21vosUQcIuxS5MQ21mTqsXPRptI5eMEVKb+cpENpVC0j9eLSDRw
1E7tj9yoQnLXerfjIcJJY+0Mh/eDuvaRn5Mb14PuuAI+g1nRpyZe1AvcH/ZaP37LnWFoIo9SMt+5
ucma+GaurTHnXM76fiZRDuzlbaYpmo+ERjlVgiRnzKD8gad0SpOStVIKiynBsfXp3uqFmnju4YG5
Jd5g/RSkmy4LmL2m+6keCIweIBkG4/NHz1JlBuvu6KgDQvkFcQvwnn5vGayzb+K+3BxpIoRYeqrZ
rIK8z3kVEFxb9l8sFE6c5aKfaR+D+ixHeNUFyJwnn2F9Nw/9VQHCh7wcC5skwPaODxuuv7c73dGF
BFXwsKelGOOK4soAYL2IJ7KToep4AwV+nYFF/NZOmFVDOcIWBYi0K5g3zXc7MQ2xeMSBREYkQUnm
RR6Rtnuk+H4qAiW11UYhVAE8Lm6+6EhscsPc7tYwRu81tKe25t1pZ4ebL0nx1ubd9PIvDmmx9/hI
gsZba6SOeVWx3+uAqk28ZYL2n4QDg6rHvnv+Bbzxi/bu0m+0B+fNHJsTIrQNGlxnZGDtxaBFULQB
5JJiF3D+RLcAmsM+Ij6RXlDZxfNwcr6EemKwsD3c6o95Tsylg84wc4IbNNp40wHbvrAwA3zx+TDq
7GJrAJfgiklrzFC4ytm2a7k1J+8LM6CnyRDa0wzqOgPyrGHeWBvgGYTDukvP6K8McWXmHpAf8iDK
R45g/WM9g5o8kO6WtQlhDPpV1lcO/S/IxhavZJwkRVwRKzniFpOjqGwDxJDxM1jFMyUxwdTZS489
NEjgpSMt85XWr6rLU6ct/oUKfvCKsHmvGLe/tvpmeQgbq7pn2+kvldjxUXxHHhw9/Ep3e2lF/49W
JVUsMqjMjnQo/6HtzbwtQznlNeTOWqoFn3L2MA+NNENhhbX6oIzC//1HJ+sMl0C+AbPBdoY10rmA
LfM8UJTIfFvdt2QGSz4UKz2Kb561PZghxVb6MvQmh4DkWaltGJrKTUfIgd4VJHoVcJvWxVGhKPto
fQgnIstzrD335bM3uafnrdMdiswmG+4km+YUJnFcKQlDiBK6B3dIsbizzOjuB3F95YpUgUNb18QK
5SxmN6py+edk1gPNLMsmsk3GQq6TLnRoFiaYRcFZ0mFPr0ZvR0aC7L+QlaE3tsKVkC/sWXg+Pdsx
V7aBnaVaRPUOk4UsV7+a5zekNUsS3lQ4+jE+Ibt7rEfRuG1pT0eT2gboaqpD7l8gTnxB16deMR49
xf7duQal0eY544s8nmu6hRU/JYRuwJaF4dEKpgUQPfcKadKBFDjUbtT4d74ZV5nBfywABeqllBEi
MxZ2Nhz0+izF7tl9TWZxJ0CQQEnuOfYqkm6xXnha+UjO69CII/SntMgBzuz7I88z/iqUOEoEAbv0
olrXmP/gdkxifF4JNSNXIgimw0qRQcret/fLH5vcTdE4c6iMUmdypQtlHa1OZhkysc8NnVE+pD3i
WfVFKhyNUPAEzG9rH+0Tz/ROvH1/kfDWGQ6wSbsJ/FZmJ/snkLtglLUZPUDWdALjAqxN7xUrpKlb
fHw+u/7xwF1Aw3Qm5GroUprlXun06S/IUOpL8HjNshzYlgJzTkjI0Tm1sOEKhQNVJNudbScgN8sL
gbLoW1IpqFqD1NVrC7042WkOkiovzjD4u61oWy7eLCMvLd8wFe4VVd69hrI3rkr2+7bpQTCHmmol
dd6dTnJXcTBvxPxIzLh/MghcHA381puLGA52sYTeboIz8VHaZo7iB8dR4a9mS/+tvmEqfVp557sX
W1vEGsaDq2exc4OUzTgB+iyOXgIuv5asHmroinHQgjJVOfKR4QjB7EYp6qmT1wO97KFPhvsRZtHL
zb4sADN4mw5yBJEusJOWurLEh+FKkfxJG3e6/L7mqL6YMNz6VQvTWHwyqr8MO4z/QCUqQ9O0X5ut
Q4FfkoHy8ysUSSzicfcD1XwAC3SpCs+Ua8BeuGw48qcylSXTRV7wLRpqP4LrSANshl3rVSSh2YAB
44HOdKFtauD/N3FbWTNlc5oAs2B7tTygvmyru0D4ERhgfLVt/fljZSWBfsqI73Zd4HNHApnI+npe
1M0uMKk3KIuj3Y8T5OagFktG7KXMlofHjxrZ65cH4Q9InahxLqWEdCYpGMjRVWR6syrCOBl5vUG4
ACFBfaguKndYhfdBF+pEwIkpBrVu0BaaeMd7Rjr9legvFAf46qyE4QLyJfwXNk6myXY0+7D5ZqN9
V92zbcALZKaYMyZ2r6Cy6IAbkYa8HffG+DwL4ioWSeU0klg+p6edwaf4lNNXBejihSNHcUHAO/5s
LTvI8Ey37x56dddnulcqvQUywxhftWR0mKTss94BGvCgl4rBJM++8FsBfrOYUzcCxW0CSC39RuVk
cUgL6KzorR2HcVHkqtq76yxznwdhe8gdVrijKSdkhrQha1aB2TURDGKyJiZW/0OaBiGAmN7HVo20
ga/rDyMoqMQi4ItFVkWTMWSzNJ6mBdffa8tEwvZI/tZ/7dKkZl/y7BzdAa/QLyn1urt5DZmIKQ0J
MA9COmhycTedFijllIX4BkYp0UjcPxn0Q1zbUh6GOAlsV9BZ/UEE4RU2FgNMfJyfB39MvTeW/jKp
rHQMs3BUpb5CFw/rsQYZGHuBGcKQI6nvS+HJGJFjLeGI7sOCcc4ymj/ydV+Q3UG0HO0MDWn0Dr0L
NDbBseuUMMrYsHoZpKfV0CEqVlQlWIVPNwxQk2igmqERemCXw8JUif4FEaeIhqW9ZHJiARThujDU
D28qo+T/WEF6UlHix7/uEf2KGIBilYgT8At0QfNvEzeeVRYuP+4Pm1bJXs1LFXSlAKlF4xUQ10PF
GYWvZcsXeYw+7s9yGWcJY0je0n0kkehkUB+Y1BCEmySz+/p42zIM2VH7Plem8+vbcPJRXR8/HIyl
WLTfjggH/psKoQRA3MxhBEIUdLklDeJ9B9Xg9WtZrQL5yfaA9nAvzxSOtt0vluWOxYK69XNC76nS
vUDUS0FV5GHDN1pBlZV/8axRgnUFLzMtkIVZFqub1ni/OBYzST0ttCCIRx88ARKK+Mqhr5ogVx+c
444DOTIFY+YUYiZD5U6dby0w0ZZftYsyQp00mvt4zQm2nH5ZEs1ctyi3kAz+as6Ph9ao3Ot5We8F
VwlD/reJyEt157a+TLpm6aJL/I2G5k5uLK8l0YlLHV4PjyQutZLtXI/Cb42CYTBrjakKaxYIpvo9
VsZicZ3g4Ud8TY4BI3SuO7U4hrzXm0bQ034pfzcl8oiGuL1aG+dXuuNvPNeQI06cIcRtK/tcTYNv
n9W819CjzC9MG2VdfNSS33fUlDVBdKf3fBhxnkis+WR/uULvXRyGWSAOg6fr+VvnBTvQZcz4PztK
dutYm3blod229bSHBT0ONeBYBv7QOP4tUfE0I5cBgqOYllg4DfMyMp4e7UZsre+OAUbQNzdUf9OH
bX4leVxkiwyMk0+tNsIHcXDu9nCj0/4MG2XlI0QhcZAgNMMNildLMxXnWzmwf4yD/TD1G6hOOMmM
jiXveZlamye4KGMp7G0IN63sVfpsnwQcX1juAwuIRAPB6NDw0yXiCkAiZtiN6kQKMnruW7ERXAov
61gR4QMzixVQfPgrgYOxSJqLKBjw9F1+lQaFm35FtQLS3f+zR4RMZsTluEWhzfem9/no3Idz4llu
5J4FfWF1ikZEPi3RCUgPeVcs/gYGNFl45bcwCBp5Sq1qE5mcgw5Uv51xByT66XtQfxBa7slDrKcv
XSYsRy1J9DuTBgys2klV95B5i1nPpJ5XFDhQbhMS1VhCB4TD+FJbZksnCnYg8aLbFxnnheMz4YGh
V53HndXV5E+h992iaClhNfW/497mFAq44M+qOK/VKoiKoFCCIRwynDZBKMZaUglFqM/pKCX5eagk
WfKLIcUeQ3sFHZ8CjzhaXne+uJBsODMVpKUHevrr2JSCeNAinVENN+9rwphh5CRiyng+cz4lBOm6
CaoRFwtdy7TBKIBjhNOUxboqQgeB+gnFJxNYYXzDzkgpRkjlnx4zCcunyuBr7v4YnFWou9knf7PS
XRfWLaM/CEBCEx/vWVM3NkLp6VaOysQnhO77Ky4HCI8QTWE10GnBVQSIujx5x1DAK+eqzciFTuYt
eT6FJByKZacWcomkCoDkaH5sbINp7ATTi8w6O6gVr+dMnEgDIuqsw8RaHI1bLmjz87fAhTqc/EyZ
3V87Rz2wobC9ptOIkX88dPMx+JLriNSSFHwPM0ki7c3DSMvq2gCZIvW4MOov3DmEFu09rwKlX8Ro
ZiM0s8ys+BnkfR9y0y3p31gDZ4/FjkZuWAJ+NxcowW6sGok/z6e5zsT5qRU8q7FhBxYSQgAEqpmn
kVcMHG3EnkXiQBSTNj7lv2lYbchaC+PUty0YHteEpaTTDbGKmI7OBWy2PyI3v0n8rLvF+AhkdNhr
skY40vXqKJ6uxz6i5e8Gyp1WabxhCZQkoV6DS+xqv5mPxLUlnDPMOtTtavV6+P8CxPCX0iJjFDa2
iH3gCfVvJM4xSXrShhOn/VGFRvt8g5Jd/+9I+cFpUAe4JcSwxnZQbYfolvFqlHb4AyWbv+dcytSX
H+BqmeEqhunTIkorwhMYfDDLWW7P/hFb2O7C4IPmIn/1OkFOWad8xcCxuW3Bu758bepzLx4kgC9F
vx/13JSioJK1orUkDG3YFApxvXvUhvGG0nhSot+qQk7DfltxPto4xZkT3pF+/JFsl/HPRkWR4pyg
6hENsv0dXvP5PaPLnJ6oLwJqdBVqSTDOEGu2shThQcBH3HT1dnyGDmcIZfL2pjlaBdlllBbYYNHG
06DtwO4GD4ACc/o2abyVxF7lJyAZWaAbphA/StVy8YCLkjjelqRCNCDmutmaGdFoQR609yQNLDHj
QfKFAF/jLyJIrdApSveGN8b+h154dmM+oOg0EXm7L8LRoSXpM6pyWuinGOwma0mLZXTbfQDzPjTn
FyXsirhC6PHVtaHeKD8/C/2ctrwIDtXC8CVYCQCsOnEaYV/pTgra3lcc9A9e41V7SHZ8VJPRZGyo
cgD/wH/wseKt2jn2a5ZaypjgoVu9d1wBn7cLhPf0FIywiutxaUqUdWAonpl0tPM72A8BDLpt+EqS
3K+u83dguhw/T7/57DGYGExlegWEZOefREQFElibvPxS+jGxeai/hlsncrS8Qj2p3bhLX+nQjFnS
UqUG/qoL9qPsYDBYj/jsUcueOwqJDLfYJlEcHGyThkcpEhvxg2MHJ1qEY6A0cUzX+XlbKIw0sZCh
1faPmbmumXARojew+pzweIkCa80xvgxLcesoeupqeNpKI6PWMiswgswY9s526aPZQnO1RRhrN+Xy
LV1ITc4P9ErB3w6iu+I/+2Z9Jm+6bDNRLWrsO2EaoutwUY4Jo5qCchUweZoUvlg3PHVLdo4dERYv
uBQHkGXCqoxgHrQ5Kw7DPjDmqGYF5pDOZ2rwQh4SwU5Z4l8jOS2W9tm90tJv4tHhrmy+FcIofOEJ
x/fsS79nxFJ4AcrtUjWfactwU1RskggmYoj5EJd9WTtNh3Ja6H59vEL8+/ofUQwUkbrerWJYivlU
rX8rcHo/UEkjEvIIAqmcygwH4FcGc69j9W2QjuPsxR86Bj6Aypq+JqeDopzQDmqvwvdTzIhPni1P
st7B7Qw5es5AM89qWoNIXX17vkVvnTYtxfkhBEsZriWjk+TFKFo/TjtZTCJIFIvwoqSqOC2oPsPX
c4KVDJJ+Fd+cYYivT0BNv5v2R9A15Mrcjn798XFm+jmQmm0JpkGlvipyv8eyY/yucvTmVMRpqf7O
yv6WmckZ3dBXvRLhyW1MC8PntiN3uxmR3u3NGYmPRUA+uzgbeiOx7Tw81mD/x28+JL5UODN+A78L
lQ2+gPTKAEir9U95twF/KSipmVf+/kAzzeT2e9bOwMgI0PlxZEfQUQGEhIjWkvAAs+rJFFyVKOhW
aLBtEh4tJBMveZM96aHY0SPyev+gp1ZITl6CSu0knWksYzs6HFPUzU2r93uiGDkx0gmV+LA4InAZ
o3xr/UkwBNRBfgt/l+LFiseVoKRfHeAqohx1TidMDtoRbSHlRrpCzR9DJC1kNJsw5w5tZyi0b+gQ
m4ydtMO6Nqfd0pMyh7Mkccgaovo03g1lw2YcQFesc0M+LEszoJ+vDbtimpyo7XGEXLp+wT4pr5pl
5X5qJkgRL62TWlwh5wtYWFNWLXr5YxI53CQM+0ZyePybv1Du4xw7c7ksJ8xCRacNywWy3Uwk4I08
nGBQZE+qw3bKKVPIMUEdYPcMssZOMs6kmWpKqxG1Q9dydrI1lNeMDJRddycjW+qk9SFKIgmOdDtG
d6fG25DB2/rKD/QRoxWlyOaBL4PPLJFfXSjHUEJ8nJWh+ATawha5RJj5Av68lFwDAlmzBxVM1XHY
czvFBOUl8nBe/O3Fgbbmn68HZUnBuUbHMIip7rNMoJKwVc+IoWPIs/dzbVZLPwMUUc4LD2TSsdpZ
t83rjtf5rTSkIPsQ+SuywMmuuNn0/gedA7xpn7ztdOaYKePkn0H0d40XEXuOG6VjTIbWfedfufNV
7csvFFTLIFoZi9tzlZ/k7Jtp8ZGeyaoF1YM1DbvmMGl5WdAW2pLdMQLsrpwS8/1rZ+hyNruz/POz
OJQ87ZiX3ic4grW7s7i5WznjDoxKBNdZO8Ygjf6mV57G6mXu6cQIInbYpRBggjenOd1cDr0ajlyp
A22JyUhZ9n8DMo9DbI/tB05H2cGWVpCEtTlpgQnPi0+EENTE0rc+uZ/gCv917EuF9iqg5wpi+zqF
kfihaQsyaUqFXZAsOVri9E0nPPmu2fJz6Ea1j8eCg7oUcIHnxrDCRfRdQcgCtxOsghopb35jF638
kRCssKo7pThBogtzy9EgE/Cbo76bD7R1Gl7G1SUJQKN+y2ZQRMdx+YFFN4P34ia6nsi7OV3IO4wY
VNPhlTg3zBOX12bba7nMyxlz5WMDy/mOf5fvGJSh3z57wllXzYDwGyIIQ8KP9/3ALl8im6OIMbAH
cAkQPsHh3GXjcju41PBLE7UKAp3DP74/YAJ8YGicmXDo6KRdXzZlyP4P5y4tph8CaPghXSM83e0R
LyCXjCEAcHvKFe4IKdYND3bH8NRyLKSySO1zZsGn8lvjdtMeYSDu1NbRb0J3gyh7ToXAxDfk/ERY
OaTSSObiNT480PsrxRe3z2ZWxuksIadgNYKFVJwEAP3HXA5xP05kW/ESsDZmhk1p5ERH9uvnVyQ+
1Bs26tCRQFyDMEiRwSbaQlK4nUmldBSf2BM3nWr+meej8JOQ4RAt9nrqgGdbmZkVlUcW6fc2SP/Z
8XSrmLkVd++V/UPXynOUR9cmGW+uiWe8fDavSkM25+fIzrE9REF57Yg01gyIG+Ba1ECIF55W+4ZD
hffaN9HJwcxoj6b/vQL9r/yEdwLYQPHw8DDyKv4r444QCHHMztRjNRF045RVLvz0zCtSABUvMvv/
+F8C0P7KD4abVuBguWv+3vSeVpWf1W/QUgeGqBUdqIyWAMfeTaWGQSLoKA/X4B5pTDBW3hMYxNVp
MZ70qbau+bSIh8E6YlMnAH9bMsTrlZb6xC8eRMXPf7p5hNcs0NLyk3FwClSjHBpfySxnQB9qGtcR
B3BH6q8NisfvZQWBt5iXf2fMx2IbGxOxn+P/3PrqY1KRj+z2i2bOWAAA3uzq2V/bdIPdPT2Z+Pe2
kn+72khp8jsDkzilIBpdFT5C5FAM9OAKVq0Ewghi6nScre7b2e7gLbTodoeo/TTRHUlMqwsbc59I
1KDKPFBgij/6RGFtZV0GIJ3xxNM0OvCwhm14S7ur61pkK32qdsnw1wR4GCJlrPGMQarUd3ASVLTS
4NCYyjtocgrcMhRLOmbUUtOBCdlJRX4WnXZFBNZeXe5sikgnJ7YlHEemhhonLNbJjzGQWRCaVEjo
7L/BKdvk4o7k8x4D2mQPGTs/LL/7N6uh4UA1vHP7zoOd/fOOpfWbKGnZj598tZaSORrMSPIKsGAa
QyFHD+82HNF0PqO0uKGHefDSp/MLNEygID0LlRuaw/r6za96A7WPXKrwE8gcQL4syTWVb6Zhlewr
kynV2IPfdfNsdAAQQZ0dgyn762djJK7OgdYkyY8p4TA6YWAvUm0hxtU1RwsV4Tp/OHDfjr22/AVR
38gQM2iM0XeTqJv1GAKQLuZyCMI6TvDOSuRrUMdw2IcOLrsCJUcuHs8GxL6Tu44GjuYUjL55MfEY
H4bxFQPQHxCwH/Na+Emf/dBW/4mzxfS6Ipc9a3w9nxr2lAyAgErqqukecr6Fnd2fq7Bt0FjJVCh2
qJY36eLRBAgMf0C8c63gdWvl/baMtDrCm6fNiwRpUllfV/hTaJa8WsjcnJR0qzJBeVYA8L+fvUIe
OhwQP+0pbR/IZ91Gje1FtT+1S5NAfwg1gpZGS6ZZ/0TH+VN0AY7DUGeRA1+ggbIFWWgCg9URhq8i
5TMk/zPUkK2aysIRfc9qLJSu6Bm/q7f5p2SbSAJWbsysPpUWDGTtOdAVoJ5tow56T4UJVHiIznoO
T7d4rdBXshAElEyzTftUfA2fonOFk7zmtI1b2HYGeLB/KOi2fJXCLuKJCLZLIMEA0302Yj29XS0X
ZIiyxsu2GzECoXIJRBwZNzB7VfRZYUJkym+R/9t+w4w91QbCOBAnF5oM3YRV4OR5j1H96RYtvsCk
GwZsdtDBQFn9Zk5ppM4m+3hT7RIo5aCtbShGOTE6c1Pg4hVqT74wHbI0UjmmGeCUOZ+Jb533A9Ou
h+uGY0r3GkuNhHVnksC6RCZMGmp7lPsk/M0417ucsVymgAmgcffOPjugXzqJlbGLNpJx4SJGaBs7
o4etsHLXxOBNQiN6ycZLMgKN9a2HtBz25McPKEwD0l/SunEnJvXsPzpSzjA9SlqYBW20oaoDSUxv
UOz4bnOEbReikV41oKGHCA8URTctQp+DNsMkf5Jl3dMF0798MaI+F9r6GpreuLdQUpOc63kTz4DD
Qkxs/hGM5eHqLJxgtUU66tQvtWhde5jy6BZUOmMxyfcahdFGzAcu133YsNUCNy0in/FZGnFo5NfW
Sk4ScdJXxj99QwAsrZWGdEnIXyyPB1o3NVG8/W6jtFDfWERu7iukqnYQ7p5s/S/I0hdZXgVsHkNV
HATxPoVawNJ/ldLbBkaBBQ6HmPx0malMCC3EGBQa1/3x4NoXOZ6f0wWtSe+5pqIymS7bojvkmR77
vvdLIjw63+OwoLrmt1587CLJktQMb3wdFaA2njZ6VvaevxozoZkRQ583M/7EY70urUJgK5Spv0E/
8K5v7h6wFw1p51tnR1lKdHnhmd1Er1X4zCV1p9fW5f/Dg+upEZJFB5I+IlGVqqJf4+YD1b4lEJxa
p2YdwIfyGWCv3U4tGW09PocKfwjn5x9VsREqAHtT4Tpja2iDZNr/uhZ9XGvHx2G1uMtiD6fyc0F9
jF6d0UTRMk57pHc5L9EY17BqD+MMN+Tj8w1EwkC1x0i1Nvtky4zYgrb2BLzgTa6/M31FiMXyfij1
j9hFoqU1Bx6cCpPWX5EV8lZFxELl0d0jSFmYWBga87dPBmkVGUlsD6KfGLjOweb09pqyVyqdND1U
tj65giz7TIgnT4qzUtTMGBgtXGLl9gAkb0qf/znoj+Hx7MyMb6o//5Ht+9Pc4Ytlcu+bnAI6afFB
cL+S7BZPqc5uTgX+rvLWQfevNTjb/357ShZzML1UbQtB9+px7uS23TI0kdNrgzbalFaOl4/qpba2
LcDEwUqu3qz/aaL1FmsHa1giUybygIinmHMlpBsI3XG0epb/DBuTNUi+JiJp4+oo9rD1XW0WxtB6
ql1/HPWwatXOMgUu6fi6NRADU63I7ewdw9hq1tkxY/+RqcWScN1OUFcPbZ8hqHzmqr84HMQPxU2W
Pgpj1N6/qm8eClR6UF5BGWJgJCgqBj+OyGWbBevG5NF1/xMeyGcrGCvVAB0OEUDvg8FcwHli/sak
JVgkltQRXYgHaNFOddMpvdrg5AuTpSGsGLiyDRlgNnXTl4OPUH0j/csoXjNUuw5Eh+kbsY0XoHrr
ZzgVbuxgKs+bV4GMqYQi7e1uix48obm/QI531RAa5YUABx7FSXxhtvn2JVhgdv0rMFJpCeZvjPTR
ugz85Z/lu0dciVPBTVR6GOigb+z8OZbvbZrQl6vXSkyKKweB5oT8kZTZRteteB9Sc1njmyZ+gqY3
OtmI8DyokkNImL15Jf7DZWr/JxSbd9PKYivk9eWy6AXPeMNtlUsXKB7KTE5F0OVTJu0aL2KDryEj
mJ2ApNO13/RvuFiXy/yBXY4/3mj+eCfdUQ9FrYPXV2qTlLy56qNOwTVkdLZdylI+olpUgBBHFjI7
Ncnbyy5bsThE7MGcaxlHZ52OwfObLq4gddoqtgFyF+9Sc2+3vkjwuGuUO04YAD6bxQMmCKpBBM2m
VC8AjyGGUHFDqmZKVWckYadpHQEAOaN1cx93FDpDDVvSFldZiZ1c3s56NyspwuloCqIQLU5p9qxk
PAPEmbg4gDY5Rgqidik6YTN71T3V5X9h5gS1iJfvTwQIgUwVOZB6iR3hOxQvA4O6WL66taaKGBnx
iE9aLZNDB4yiObO1MyPzwxq8ziWLrOiB/H+QWU2AHPbP//bG2sOa2WejV0LI8XbQuVk/mosINxjq
deq3f7YV3VidUATZijwoo/2Y26zj5YKR4Z+BM1RXklZY896pkbyNTCRRmGpxSYJv8wdAn9KMmMOG
qWDI56TlpyjFDB+gn4siWOQE+4xAGtWXJ+8UWy15oPPvRF4/35JoSpd/dSxaYUhLpS+d8VEQ90RN
NbpLoFwQbjh+y/snH/eE3YifAIIDu8gGpP7AxCggVeS62crO5M07gG1rAwllqM8nuRG0HMehrkTU
oeV6/+i78QoWHAfWtOqDpLU6YybP6+f47ghi/69XhQftIFF0L7fJv8VaUTr9AKkAsYaqzmvyL3rX
xqxPbQYcIHHmEDQcdw9ARhlPOiVo6wXZCou/Qh4uEKQIEPDBtBb4p9j7munNa+BKxLz5WCvNownR
MtCJzHdJU/Abkcuke2ZyLyWedaPjDZ6h7Yg/pBLByAM+8PRNtIvx8kAW6l9+yZLfqK71SMynN8S8
WUHkKXiC8vg83k86pq+V+TfjOGvbVnth91bxGqMdEEBH7spyMjpkH/lqSMy5+aY0JoaKlVsH8xoL
IgORM4WooWnJTITFWvNhqFOPwWd/ItqAPYMG/61pc6DbSwRTXKfgQSAbah4x1WwOptvcq+LC2oNh
CCg2YWnm6uZB83AmNyHjDHtnCW0NDROBojj38ih8kig5Rby4ETsdFIRIpZmQZGR6g2qcyHFUR5Aw
bjRW7+JDNXzQC/W7bxvIS77FUupV4u4IJlFdHEqNzWTyV3fI1UWT5nMxrZmQUeYxEXTcTqPHOJHA
ZzXEeUVCQFmJbHYudGxmfwXqGo6/D5eL2xs3fwj0PGVV2HSAN+cei2j27ddERQ/dqjNRz1X0jFSQ
EAuREQqCS2N5mLfIO7LX1DnIBZ7wXixv8U22ETXDjP5YEPoYE6G2jai1KptgTvU7NC0VAdhVF8J7
IPom1fzLkzVDDj1QM4MD1Gcdz1CHEZihV7SgTBoCe9mgHYRW7DKolWmRlwks0jfuH7Py+YWzJzW/
gMoEipjY8aCfdxPJZ9XtQGGyZEf/TlZm9d8h3yz1fMrwwPKOo76wiS6Ujw3NW1ya2Hqfts7iSg0q
2odrBFHegUUUjlJv0ibrKA83/uf8PIHtkN7h7ZwNHmlC2/ylIB1cwZq1FSJ4zLN8MzErG0kcHRGn
EAu8lWAdDYHlwzRDVt57KcbCEezJ7qKbGHt8UxIumWgSS+gwtBtVi0LxCu/KvXiyWq0eyHVzJ8WS
X6065OoH3BA3PyFjWViFaW5oF9kjmB6nWzN5NvupEvG6nNx0UTtscO+w1SqZksFsN3y+u9N2oZ9J
wmii7HclWqT7984zx0irjYBQetiLMndJD47X/+W6gJNCJ+nLhgQTpUbZHHunYznY+YFnc6hcFTmD
OkKEpjEW4Tq7YGUuCTuLMhzoMK6qGBGUIzsIcUAkuD9yq8SnAahNRhojbm8NCc3UUwHEU+lvlMRr
FoGl9R9L3ueh/5cBCPVMetFjG3yfGAfiHZdGu4dOVikZ5dM8ottuyKsETfLIb2PcPeU0IlIxpjeO
bqH0Dh68s1c7NEU9D4ApewEi7x7jN4YqgTC7gC++Z/MAoMWWOD6n4hxKgdeTWJmIlo1Zj5aGchm0
SRQuj2YMlaMuNxZvW9yPnLbflqA59Og9OWya9M9tfeiVXztd03Jin1FEkZDvnmW7+Egh9VR0HtLb
ih3SF1SlADjpPnjuwdSc3JFuVtNEpfuMdFJo+tlgOkTxmUhP+jeIAylxQZNVmYfp4X9FcTvzHH6a
yDX444JAqFNyvA9+z26d13zXq6ZJnx4ooZXRM9mnCqOjBad8aV1wGBu6C/ku8EeNFm02EvaqOAOc
ugtGwlJ+ipFiInJ1CKiTkXT6k2V9/Pe77s50Zdz0kFOjeHHrlvYxZwLUXwCBemXBGUs/kiIIDLW5
GRAmu2UJ5b0wMk0Uww9kdQOoKKlMi9/MkOZ0hiC1aljcXHTuNCxGf7BT0Ah913+6llseuY937dav
0uFiSsI7Wo0CAnu1qsfLOvpmCHGA9IZaRNf5R5vud/SHRxVCqjuszPUZ+2PgZAqzE9PacCmloTNf
6YcLJI2oqpqqJwnjrrC3lZ/bDmEH+vUdVMvv0Qagp1Rl2s0pFe6gzwq+5INcHtARc2OZvyKEl/NS
41EKMTAi5icJ+j7nSDAH+dIYGFe6UbKypZWq06qQgBZcmnLDMEyyd9AqTpitmFpiB782UIXX6m8e
REMZDc6QrMhsykKWDow8h18VAFrkwpekiYPNTVEdCFi2IRDks1b6SJqSbFK+OGOBYgqPkFnhBIbf
PZlAWIVVQuEJwOwFjXWimWGpxOHDmKCAtK94DYUAq8E0CBBRQXrf7Z28GyBqyXSaVnnJg2DuOrrX
30DRnE8OYweiSztQYGZ5i7embMZWdYZzHXHhNPiLv2wfQmdcKnYsuQhYs6i/OwhVvLnEbh9RKU79
ogyylKB7OH3Ma6TKPSqgqifuBoRASoM3alyxYCUx5X0aQ3kvuv8iLaWSUmxsc37f/5XaGKt7akOv
B7/HieNAcivNZl9+/mnHngqI4dYT4NslRcoDOrt+WK37siCU881nlluK02DD+/Pv2nNEoRr3olc0
r7xk8E3KE/TZp39P28elxxWAr3aM0QTk9vV0JRyaKLH9szbZRaWKDSNOqF6Ku/IHr1l5T1r0zIk7
5xtPfdCRZ3mQWxZu24uQ0//rmy5XwPzBxjxMIJrBEfZZQdrZ2czHny3ezdXNuC8x4wuotxQuJ+A/
57nGcfgh9oiCgYjm/EG71wWTdGzEmzvmbX9Fiiim7VJodvDW3nMznkfhEMOVHSQF9eeYy88QJMsH
2698cmFzW/RJ/7ZPp3pIYlHNy4zmtaLqc10/lc0su7s++a942dleTmrIHXJ0SgJMJqw78FzjBFKE
LJRdnJZLVyFiZndww6/DBGE9hZQG59QVPCyE0rt4FQbBtntTXVN3eeTFMj7BHv8cYdcHUx/yEbXF
DNzz1uC27g1J5j8WX8tiJ/oeR8PVMK7AwzcqcoRwBTsGAXNNKdehZwWamYDzshxANDWmFDMqgzZU
A7k5T3Rbaa9atVHQHWLNEiJ5VU2lgmdlDi3/2y6k5oXXLao765oF/FIskspO3420uggWqHmOXHjZ
+OHmGF2wU7eB+/oDaXP6OajhTZOYd5kfhA+qefiUo2sPrEBaP1nt5KD7Lkx5nYFrqDPDleeL79r0
d0ULjzoT1io8rfPIEPw7HmHABORO0OiPh7wQYTSZlzbk9J9fR6Zk/iXf3WwCYuaZNkGwfUOipQjU
dKRdE576SR68Rv6TQVUnKy8UhZbMu9Xnun7nHTV/9NRCFI4vHjRKIEioC2Q6lE/rHdJxYRhQl9pz
Hr0+pKAYuj/2o/eHUU3UvcVMrsAcDWmY6NoVNWLVL+j23mGz7Pmm5NnYqJWvI50PEKr0yhOt6Q8D
+jeF1CscWPv7oZDZxP35ezaf+6LcmDh6rnzXsK1I+d6BMhqBqe/9LjR0tbCwK4eyiRI3oDkPC/y7
l7tw4cSdbv6NYGJZdlM6j3n6MmDZPqTBXmynse/qZoXyx3bzQW7nipjhwHNb4eGaHdycJpSlwPaj
C/mR2DDcR8gcGlGQJuXclzIRoyvCipj5t8lKw80bHOXIsUXfio79OtCZc5Va6z2Hsjy2V/dqF2vO
wSLwuTmLitOM57B8tbzE0Ha5IyXkNcY1urXbx7ZjcmBok+32oKybASoDYugT4k5x43MkLNJCWQn/
Lb8FPA3Dm432YNirlvtNDAkO+H7Myk8sBKYTHjT0aiYpFt5Otwczaj61Bji0fGV8DJxx0mZHMxHY
2f2bx3lgQHLM3kUc7LbFeOVJnVLugkPSnuat4RIkYpW6ByezC7kwJTjJKrzGLfTeYUfmFgjz1kxl
t5lmgHhrLDMV+/NPpw9EZaxBHiz7vlM0Pljv2/zxyk24jG9vrmeyTcOBEzHebkvAt2TURrzleGq9
XJMswmRIv7vgkNbg12gUnX8qQE5uTRsYNyEACBCH12VeuInMrLLPbnstLnZ8krS3pipcQEaJN9Dw
+sylLa8ho9QIlpD5U2Sy/gCGRs5P4adhVSKcfWsWHgGCtgok2F2JoKQnum4lSbJfEFL6pib7oJyf
QM4CdFxJLp73LY/MSerd4pXfyA+RxKXU6v5eIsWeoRzuA3oBiHXhYI4zb+p8ewjOR53grFSgxk/A
K1bU2ubVCHIN7yZc97jO/WfkeN3wI6vIZ3+HIvDFyU6SxFcY5otzkqWHLT4nLfCSCTgv/rErorao
qz/yCxY3BPhxRJzEC5DXMZqA3auToL0nOi02I2dK8zxqM1eJHaoUw6o/nLTlsn8EnhOIGFOvAfcZ
nikUzycx+8+NZn+FLN7qUnMzuJlcp8fyS5Gjc4qwbeCfPaW1tmXEwEQv/q6fOrE+LA4QmaVzs6g+
Cph0byw33YU6esEh3349DB9OeHGD/3Itpcz3zazboOC6T+X5FECUodyIUUxyogjdPV+t7+RfNIR2
AFVi9+EsLnfmKOvl0DymGbEqS3+sU3VkoKW10Gu9BCm3zW5PvL2HNXXP8Aa7wKdLVCl6bmQ+TjTz
AUsoihgZuwq/3HyYtFhNnGCuK8vKOmjcHCb9asnMr3z3hJERqSXQwMlLHbjw8PWKZkup473EkuyF
+gdA2Mamwp7f0Pw7/cb0dN5GYSduHlUT0BM+CSNDXHYXAqrCyQkg27983Jw1WCOPTxi6qqZzPDZX
p3qhg4yB+2Scb8zUAjjazBOz3PERLQ1zDUmqqKVPFiEnvE68YYW8C/C8ApYnHFS5e+szmH2uRkki
ld3nRrcFmYAAoOlvH9aaZNRGZvSJslVcAFGRPHTqU5+uktfwtnDKSTTSF38Ezg+DuZVTEm5pRqT7
0N0Jm6Mu2FnVcBrMTyyvJSEp3xvhYfaEydzdMXzIT1i86ur3F5y5JjtKudUzT8lcKFYDzJ22DTrL
pc77ELhxFvzrPKXhn+B/8p2LZgw475elMngJxGj2HOaA5/TNtX8a2EDvgQ4T6fu/Ez+MkW6ta2ir
hp8+LThqQ/8MPiFVL86hVV6nPlEfTLLtexCnRtTAAaOLy8uFYNpcA5lEKgYjd0CeKbCRSYljGcfA
oLiz076A1Uaf67pDMBwOMD7+YYtlmbZ36wMXbbJEhQnqQv6Uq8o7ScPgSTIc6VMGPXoUuh90FBhc
ryhDpnLcw6lKG8s+g5FOMAeU+nMovKLrtsV64XOdzxWyynU4ESh5fl4SIUJO+20rJyokJIUdHvDR
EjKUx52y7r74maL2+3I/W9EYLwV0eqjKzxvWgWQWIqZ06+Ds+49yGHyecUip8r/QUJdq3O7axXWl
paw/yMFad2Ad9etKT7IK2D/qmaGpgzN0x4WtPZ3OVji1LqbtA0v3rhFnVfSL/jfByUmzc1hlPz2U
ItF/9s+YGmXCbGjEKsZkMQKv6W7Sjlj7gHd66XEB8OIvZc69/ltn7OrUkkJALWGYBdPsWES5Kpxi
Hvs+nA7Zn8QUIOt5xi1WXwPfIjeBRhLbEQItpXjpp0R+Afu+TI5L8mc4SgWNu1LmdBFgNUChTz3D
Ppd+IlxfexUXUhXFUq7A4nIKprmehg2Be6oOQXyZKUEpo9i0KS1Xtr2g0T89KRVAKMlHVq79aMw1
7yL1HFq/NDB16Mz3a6eMrFnTWipwcWgc5V7A+sebYo989j4sCmdO7P99esMYSfV441QONTFsXQuR
yVi6p5PIxLk0IlTAfEd7E6xpm8H2nuSGjhLhdOp+yY4hzAVQq6QZcVZRbfGq8Al8bx1uboVlQhvv
xaBylUmg3xPALjDd/RiUB5TGUIewkR2aZjYQDtTdYaFFm3A4y9i0+wxnXOorsJXVKR9M9ytBax1c
gsE8XaQ7Rrh5c1Y3PPlq/ODdEMMF+IdsO9ZoT2EzeBSNE08VsZ/3Cwp9ii+XXDsTG1TUBjb0U8Dm
LLGgFWAeBTv8rsJUifwYUU+WoTXeKBmc+LRfW/bsrtzoRBRsa2a39fLMpzGDu97EzXOBReDEOQeG
j9HjghPAk7xfUk6h/2xgzLkiXQfqHjnyCvg1u7jdQHiOu7r+3GjOTaSMWuS5satuDb8TLt5FOc8y
BaJvAUby74aWKX6bXTkLsssJb1bRmeDmQAMdUki4MNBs8uNfOvu+OrqsKvbwZm8aIernJXZIb/6O
oATJRl4kjRZbrDUaqm83E7cgpnW3VGmyjBX7rWM00M6Cf+5Ypz11d6IkquoQVMTW7gVkGMKm2qD0
6Hi+poCnbZzWDNRi9sQryjAWV7gxe5/WB1/7rz535USF7qBis3SWpYH8A2aQPXTW2M3qKrsglbuO
ajDgxAmR2WImhuuRkDwYGk6CLuIXRTRZuvk27hjNXhtfGO23JgWnza2OPx5g7Xn6JlDJmOXR7e8F
GsUylz3LBnSQesjzfqNScAxuoCaJMTejid+mwNR9lqLCrpP5S3h8oI0/WEltPzV6fFfMv7QTYuHx
bEBpXnLjUGxUMkOrCJ/qdyn0mCGTeW4kQeFBJA+9k6q/s2BTAUxMnZBHjS+MXfM3fpeyX0mKih55
hmGNcLysHT5ivlj7NBMgWiju7ivXpTiZR4HU0RCNqwrOLXkqOAfz2ZCPPH82mHvBkmiaNaZ9jHoL
xeM5I49XZUS2a8OBjH0Mwn7nsL3J6kIfYfkAtNTjxBTNgQ8iqXRscikR31FiPV1nmfgjvWBsvg2B
xNFxHxblcyJPO0a5j2N6nWrP0u6YHtOJhJEuyR42wep4VVDIg+osp+Prlo3YpDJ3gDqMJRF2wHIL
sg6bV9IHDWTqIdZebpBNfFxg2QHzmONdADVObhy7XCC3igynYIoWuSGj1lc9hdtL4X2NTNEuSDUM
bH6/K/ePMXRqo8sKijcczlxaFcZ71PWb0W+FtfhwfgmqWtyrxcgmVbRg4XDlx506cDAjoWEJGYC2
ohBhVeDl8Dt8CmMyvf5GE/zdIK4JTVAdhwgxktZHOchFMLyWZEsKok+azhDa/gToPzP4MQKhdSUc
IJ1r0ZMHJfhRQuU6RWqnOj8kelzoHdcLvnnET4FEBANyLxp1fyosi2aKRHxuJxVQVOBfgd6Eke3f
dMsCFACBT4qJk3/hMmsBY/juBsKkD7zqPNN0E9eQxucMbTuxceaFW1PNYba8GFBf/ZPpnSv6ygZz
ThMUFKbLAD0o99ratk/OX7amsKdAd/SgEhhBziADiZl13TkEA5jQGy660xK9H28fKyVESUQT55Hw
G5NFxAWD8cvfFTQLuyp4Kep0ILAp3GvVHVr5nSK0cAU8A03douRmKuo0K15iP8EKxojy/MeB8Xq9
a6tO4iR0m4C9MmvlJl9M8qj59mFhVZY/LNMzvOxS2jSpOnfuxXyQWYhb3XKrhDZX6ZwZAAKAf8Cq
pncK/0OfzxdTrHbbhsRXdOZOsjT3qG6VMDoiiR/Y7Q7+4wF4hzdFpdwT+oTzraJH18VEGpYeN8xw
VS0i74vno3fyn6e8tfNDQ4nDoAlumgfAbLy1L3jkpwQPfLwepzJu/7/p75sTsFrfQPzTKpzxkKHb
iHBXTrLzqCiqFrBCbB64ifHpAZOgAHX8+ont1GCA/TJUFQLKFzQ7Kgm9kit+3wMmIhvnQZl6KzTC
dg0HwYSDkwRET7y6Yv52kbeYyuM3Yqr8oYIECQxtoG6/CXC4KKkaA530N/rJwOvaBJozdxTjkvLQ
CdD+XBlyLu6YQntzV7r+j1uRWLxDv0hKwvJl86PzE2k8cUGmpYYeY85z+dmQwca0mHCvmwtej2bL
lEWzfK0y+lpF+9R3LfuVmL82Palz5QnG0aOHvqZkMiCOkgGwAhxQ4ZOxlIZcwgYEa21bsLcgHeda
b92u5XxuLpJ2iAEdt6Hj7inDBZjFnOEkER9KOKMwnaePuRTaEvid1WbsW+jCWXBDGFzjVL0KO53F
81qeIgoJOQ3RUFirwdxX9b1C/oJ0YuTD3IpZ6oq3rcKwDbvrU1j5Ee2NeM4AlO7Uo/y4rEvnWNEw
KdzwCkOgh241xm+2Hk/+BkVcCEc6iOLzbVclifngPxFJecxS6td2JIR22EMipWdmi1YZAAXVEOHO
Fn3qsjR67HZLbkcYVQ5XTKkZ24sP3LdlAN4x3Pm6JG9BVfMuyqMhct7DX9Gs5otAm4d4xas2Nm0/
VcqQBVQAeXwNjB2JxYuqU434QqwTLstAKYdKanUV5w4aosXz50qH+QuI0VxPlJmQXd0YHX7ESvP7
f2CefVSCeEOXdM9w2rDXWhg8tf1FLWssGKr0ozwBxKnjIvsUe9KPHuACoupH7nnF0eE779W3Keyk
HrU+5Uz+QLKQdul0kKZNyWM+4hp0+SwGL6NuI3LfFeIDmmjgdmR54uSiZ+ZtYNOajVaPE8xR0GnG
462KL/2ofaAIcq5lPK23TbKc+UiDrmrHrlTLYzrlLjMK5FNCmh2Gn8ye+lKbECeNugqq5X3cDa7l
wXuI31RjhFD0X9mJVL+/biTYvbRnIVGl/KUGjj65nZ55l3dEKhPvqOCheE9Q0qYstwgyTQVTGYvJ
6tXA2yW8pcQz4KahmzL+DmMH9mvnknD/G5EkRUv3r06XLekWzBjbobK+2Y0A24CeilUYuiqysknx
RfTp55LwmoHoQW7pQptM3pHccB8JC1Vy78v7dUvLDBc3sFPnF1XPYerHwKu5FlRghgT/FUE/0LyI
TRKNtB7L2YsabL1TxAzo9WnR3dUqgFoPC1hqz2tPsLrkitm2tp53n3/w4TOCgM9uyjkuOc58MpIo
4Bdj2jqgDwuz1KxuoBjYUw1WStqio73LqyvBBnR8jDmqeWMjHiRJku1DfRe/6LWK0IYBgIVmmE0w
wk96Wtm6ZquZ5RhQ0SzSoENUIE6uATZc2Jk4JeqMTojn2m2/6KQY7F2uk+AbJk16XbBGYIvVSB+M
+CkexU9R9qIe3NFhVUS/rzkQe0ZvYSUDw2AmAxxx/ciar296HIJ8O1GhRXhxQziKR6EzEBqMI8OT
Zebd59XG+Z2SmHOJ1cqc3KjAqYewmLuEU0fY9cURhlZ0ik/vQxCRqQcGhZhOfe2m/pLwSAI1sGD1
XYtQdeoZT156LJY+pe9K/Z+lEYK5Qn8QEtgbCWnzxIZTj0godZWLi/sfBeTFLIgDbXD6fosPVkxR
Eg8ZWNr0hHtdvne4vfwjLpuOaGc2yuwljQq+cLTBKGLeuqgNzfvqL79f5RDnU0gAA8gHER+SQIZU
t/LJcU8nbaXT81ZAa0XUwdP4fn70KLHdgqT6X2AIa/PvJGqn2YW7XgGs7jvcVxvT6bFGgVZktoYj
iPWXwbkD9IqD3Ad9762x9TzhjGtmvENDCdzGjkejQI+dHcILPPjbeuTIfaau6TnxyZU3cFbXEhsR
/zcI04rZaibfeWQtsrxpvuZgMUlA3nGQ7M35D2eJXfuT0VFvo1Z1NV0/tncvHAp7Bnic3vbC+DIv
0oKpkPlqJlgCk86B0fyRw+0xODFceJwd+cu56Vy/EW5DrmUs3gRCcVVtrziKlzdSSWzePlRHzXeL
jTC/G+Zx8/sXh/xELcc/pGFE6oebsHCwqWkfEgDPWlE+kR81A7LLJ8T2gMbJhDPZ6rAuB9hpw5KS
Miu571TGVWpOuG5N2EwxmuIvlQC8ytv7NFLrNFM6HUrkgXVqw/M18e1+mO0PdfB2rZTcyyak+R7w
v8UmuaVfCAEQEZWmhcbUry4eCemCCLk28kb8ScGifQZHCYF14n8ehRBd1ytPbYnLciNSOB0IFY9C
pckL5l0bNYgELYRPMfoneodOHBvAo7DaKxrRDVXL1CZhDplgEEC5XHGA7DPlmb/SzT61KuSQXHdz
DtGQ8sK4142x4r69jr1R4gfcrVOhgqBhAlagbTHxnQZnxTE+iUn/Pkvbv6C0M3lECKg6ijgilltW
zankxZ80svoBw7odp7fIlXjqIR0oyTLMkOg/ZysxxHsG5k/FnHDzRQ7Go347yhNhHncamJWOjHAi
HdKXm5KQFcSeipDj8hf0QQYs8Np721Sqq6IZ5qjGfirT+z9wzCP+8MSLVbGNtTuat26RpdbB09LK
Lkmt38n2J0qaXOZ4EgPiftOhtcyMJncBOfoWijzgBAN92vCcV+pp1NrGkeEJKIlk2X9HkiMZuKPj
7YzPORAwyHJSWzKeUE/NpO8RuGptREEXXV/4Y5yJeFGd2t+1EcJI00jQZuUnrZpgEtxJREc5+doB
4PrP38NPc6rLAnRx7vNISHh6WCedF+DWwC0/obdaD1b31P0hgixJ/YIVtKfuben+DWA4BiVv6Nqt
g0a9zq9MVhUsKXhHSJxpQRr6UvoQXPwoRhrB4gVlRqy64+zSHucSO8gGPRuQW3LyGHucU11JD7sp
ox20ACdSfVokjcKx1cI8sxrBirNOAg34DP2Cf/2SXVIuD/QibOoLUe7Ji/eEVgdvhbgdYOB7lgZ0
2oOThBBjGgD8FtfSc3u6e3Plu8YSayKwjPXvlo9okQLDoE/zkuk+dHOEAHOcv3oVrnDO3dwk8M+d
rq8OtdXj8ockgKlp9vUkk+o12dXTFCv9MisDJ+oSF2LgVzW4t/Hs7XE/L+/WKLPU9l6LRYh5cffI
Y3ByKqkq+j6pXVDI3DXvEZYEqvT6VOIK5CkmTdMMloO4ygFtvLIxg2e4fcCG8MPW4XE7oeKHqP8c
yOmMA9I6mxWpL4nXuol+X+Jry3SkI3HMsS3ryE1w5g+9icUoObxr+gZkIfTIJoXuM+qXOs1aiBFN
hw3BIfJMB2iGJ0mlmeHEXA7Hk6wA5eaVBYct3wtA+dV+BzAf9I7yGVauy+LzMQ9xzsYVvNNOTjfV
7U3AYs6IYBd7/W8lf+NaeUbjGhQLTuFVHcTmHn+4e3PDNBRA6jDNYGCrX2RVtnbbUO83wDpVBuxy
m67Vix/yrw1w1GAHO9wXWoIlhKpOaRTSWBzhQSkS9jv4SCwh2oUceWuRyq9HYhTkc6RyRCOz+HDl
wS/JPFytr3t+445TMjOZo6K/OxIPuMdShuntgw1rTDn0fNRjxzWYNIl68uJ/dDkmLiFiCPd8apLd
6ImLOskItau/eKuPOt4RIrX7I7dVycNoD18Bzbm+qJA/GplfuZJb01G9/iRuRUymYNQOUSk40pLh
sItxL6a1gO8bylwC5M1sxyDAYr78Y2d4qLmXdjxlkIZWhH47aAHwZP/JGWo8WniM0sCrrkug9Pgd
nwu4dq+SRRlY4mCJlWZWteAXJ241/1WE5mrPNtuAZ+ltYEiFzofiODACtI7fWkKp7aGX7jKV+I1b
L2+Yyyeu4uAywHcYqdodYOvtKobKEFpyelOQMf6H3F3axw/bjeK4K4Y28wM2UKJq74Ra8yJT35qX
A8pmuyfMgNdgkBNDoffC2LeBYthFpk/3xc0/zYavUHKrGwMYw3IblD9vLrcwE6ruCoTQPQCT/scc
Gl9/F8y939j7beH16yOPWNGTMecQ2e0AuZOK598GLIe93mFQ96t0Yp5ZNu0AZCB98Nt/axN24ZmT
cv/I6tLufJq0xVB+zV9VlrRASXOG2ycz4xxgbrePnbymZbMTCk8wb8ALkkKMMz9tzlKejJBIU1c2
RNzP7fMJ2JnGQDBDGlm/MHrhvf/DkqeoPWJIHGW7il0IBJ3Tb9LL51j41b2ts5B4Ks/Sj2ilKB7g
BE5eFL8pqbr5gcwS5tnRJnVw7FRPqemanZ6zPlbT9GM//uCKzgS9Wx2DQgdx6qt0u0EKpStqeeIz
WZGVWkKCFjNB3/wYCpu/PhgPvNpSjy5NusuPVh4miWm2nX1KlpX9+QMT5my1tcpS19SSDewYdMKJ
t4bUTREHY5tpu9vtytjpYpcvmPtkfCLBBHdqjiyS9VAqJAD5ChuBPc0oq6Zm6hLq0vawYK9ofULe
JLYWCq+gBTzgYta657F1GzYz6raCm8uaL5QujEHQonw2izori/dD14E3vp228gPVlwRzzuBi4zq8
g8oGIN2RT6h6qff9XbNY2vI3/rJLVt57W6hskkulAPF73ze+xzoVw9H5sAk0S+/yQCWNVgXjRACX
XUx3pnRqRX7Qt8EGOUlXzJh7QAN0GWZ7jkjqeUBgXsBWnhefs6GayqNTIrMK7vnTqn96OXRhJDz7
ifFSpP0Hkd71hcUb3GVUQWorUvizx+bPlbJ9xAPrCoxbLivKSLQhoabPjYw6nqma+XLoKhQJsWdJ
Ceo/ojYcjRZRnr/ZE+LFYChGTBrnJ7MBqUaicT4zJAkfIDZ2clVKCp/NXNyBHLCNJZLtXiHKm66q
OoUJLckhdkQM4dEH5rSQhn5L1nizcHDwCh9GAIEdc6TW2xOcbgdeO59JZ2L8jasWZRPlgfFkZt/J
dGy5W5ZwAgunDVNbcFLS2b+DRZoWkCYYp49wq7pgEBcft8imx8xIExi3BRxQNYz8/Wqb4ZTE3iWI
/LCemH99NAgvUjY49NeWiWCanix1W3Xv/+y55M3HeO0xytTYUtOi1UCnv/jQdVJsE0FaDAh088Lm
AbwBeWQdzbwU6Od31RN893kMgv/27SKMIe8Y3WnlGRzc5vlp+48bQ7dVX/+uqReWli5I2/PhDyus
+IBsmslvIP7/r3bjfI6WqlpBFl64UvWlUMsyXqOPxO5x6cVexEdD0WIDP3nuNU1iSbl1SCFtU0tw
JrEzn44UeFcJUC3YX6PsU944KHVdrvZhXdXE1O7kIF2PJgdpkTl6s3yyywrvOQaGXGxhaVNiBL5W
KqJ2Sq3N9aYdgSJdpwrRdry8YvBvznf0iiXVD60yv0YAt9QIf6vxOw+4Lm0k7LhAcpN4leQuEVww
bhJEhPmdkrDgzytP4M+biyIQlGgKPiLlJae702V9FSfjKJ1RmuAxGNwMfFrMX8O2VDwdyjXxgKSP
8GxtgtrTUJmvFZ7GsZ3IPzvlrNOeWD8GCuScMgfOv5EYB6cEkUD8kgO9BsImU4u6NgpMr2xk9OmR
Iwgpf/lJtq4bg/5cKZLTVSY91DvnHLLEu8zZws3iIDOPMkmWUWCqX0GpCm70c3P6EYy6lFbDDqvN
hyzg9Rr6Zj1amtAoDpNvR35LitbPAtCu2QmMYEY7DicWaiOt0k7+3oGnxg+fFaTm8WRknEpfXtfV
uYfXf7b6KwwBTPO6LvoLNgC2cWlJoj8jIrLepe8ZHnzc1LKXGVXGH/R2obNtPEeUdxJMK1Sg5bmm
S0uIbnz6DFQXdVgFnBqSz71xpV6dTNQej4XU44Wmy0istI+B7/GEjdlcpju0nssME15sZY/M89eh
ZiJdJie2qBsVZe8XS19PfeYUYqHxGsoZ/z07FY5FbtbmA/iNifeWaAQBjcd9PhcDScbGFiEpH1ld
I0wIuYT5Ptbma2oBFzLT6Q+hL8R8++yH1mX+MFurxToMCUk7UJII7d+QufejqNY5ufKC/AQwMNIK
s6TkxKOxN1smjVozo+WREwYo3UamlKQ06L4Gsk4Pk5TE2S8HWwMGRRT10XMobRtUajGtFDKVbVXU
jvbxAXqYEVkLSWGsOHNvL+xYsKGiaDpdoON/D4GwytIUyygwKEpz0+KB+xIr31A9UKewCtPbRQUr
VEyzmqlnVYCzdiDjWkfgTKWnhj4HP6FhE4Ki+/zXtwv+5t5yZssSq4upWQ6t0qlTLvHOw+0tusPF
jCepbi1hwXP3tGUI7EOQ0BoQbLbqpRgQH/p6rbCJodzt8VVVp7j5IRrDsoSP/OgjghjyclDZ2faX
8W8gRukqQ/tVqQMTdWaDr/wPEBym7RfdlXs6iV7rRU+wLypQlX23WinF+kJzyRoTzhP9x8wJTRGc
7hN24mePythNBYiKxFPX2bVNXlh2vkr06Gb4KaSB084LJXc5ubN7hFNKalBBktCoQ5Kt7cgDDM4Z
AC6nzrBhY+d32y22waXJ54gPVQnW+6e+2eyXqJLF8bLPJzofSb2Ob18f4+BTzXcg6L48KA0K9BDx
rlHVvA4qwo8kWHTjtCIWGJivZ22mf0Dlgp8m/q3kGcmVEu9XhnTiSvyh6NpvaCFsGxPZlWAI5NGr
JRPaxPIytf8df7XUCgVWfGDpBKIgCluuOOHMEj4JOZafVvQhSLPmxqfI4kJjvwoT7/nr53tetqkn
avJDYIfuSSHkxa8TS2wBY+vb5PiKYZ2IZNQFc8nJFBNfC5jZAcObWqd8vhz7jPHAPMOIqnmGjUe2
ilELdJ/5sq894+0eKFL16FoPecAVQe00QfyYJ/C+gjjB6me1JVrwgQvtsSJinbIin5C123YxTFmE
wC28RXoGpVSKZz2oa2pHAnli44KVJQtNaeFGlgA4TVMF+XRxpDNIoQmgdM/EU3g8spRVpCu9elyE
K8mVAQeX44/QrntyxrUmqqPQsl0Jr4RziFbBnrQjbqJcTDdFi/lN8n8PI9rzV8vQsujI4Lq+7STk
tEVkG52s2gW/tdJoWCNGia1droRzta+j1xpQQVnNJ8QyHp0DlT/00vaXgDokSbb7TgJ4Gas7g23Z
jWlIMhk48GqgC48Lii+qEo4JNEZJjPIY8ZdvNKIvWfSCXSqV2K6Rq+ZskPBnKvWauZS1L3ZlvfG8
fqi3nfJJZp1UadzH825ctzFnox3yOqugJD5cNlRJD6QwPFeyvg1XAqM5Ld0J6voRgZ8jWzMcQYHZ
vOore2vs+DQRST0j9sS9PQrdrpDOqJoHiYgxI91DXLy7QNr4ZwwGKlrMN4keErM3A6+O+bq6AP+R
xtdBfp6vCaHKc8pkQQvT0rPU1zvt9Wr9Pi5B7966w+XwIbhtJwiUaUBsWNJLheK4ppEl80ngvffM
4mKhC8tvM2NRShDmEkFcV6PdhXWNflBLotXHt7xNe3BfFyXLaQOTlhOveCPRgS3UUOAHqeB2y5JO
a8/nwoaZf7SCpFZd5RkCMVw8QRQ9U3uKFbt0RfWSn6xbVeNWvwkCjugFbQEeiLzI9LNGfPi9azHm
x6dJCw0qkUqFRU7UArwvBddKID3weGguH/FysZoCWSV4PmAMs1+FB02Nx7sVLdMqjnGwjknAAVZQ
WD1wjdtJ0neN0Bf9Ghhj/SR8elkXfmw1JB7iJ86mclOCw0WpZadUSieB/zXGkOY3QPkgNoKZkAm9
+Vkx3rMTHDI5P7nA/pVb49m6bBYc/Svr5oSe9W8rlVkmbNdDsQQ0h/zlYAr/VLTxSvpaGeqsuk/Y
Oq7/DX0lZsgxj81dllBAlDWQOQ/ZXAgZ/VmUrc2FxUas9q5SDRv1Yom9E6Hx8mDycg6lQ+YPtlCy
LetARId/0HYkAp+uQEHdVCEPfxjqUf/c7b2AEBlcWyy4XOffQ9fDdXfiVs6CZ9mh8xYSx//HY2t0
E+FTwrRewPBYf6mTLXuzoTppUq/5H+NgZQZEvaBIzQV7p0/6DHOLfIUklx3TIWHhgrcRUazVf1eA
kurxi8bk5jjpZrANtfupCbP9sZIAR7iPZLKH6nJ9QmKrpaS410480UEsUfxrYpnCoVA4t2c4VHxe
GpEZyMUv188ZvxGLIUsn63CSbRNv+0YDFVayp8sv6XrrDfbdaF2b2tycdppuQnd3oeOvZ/VkpaZI
HDHmCDPo0DA5hksoNnu9vQu6UwOVPa1cXzH/GoOSNrARZPGsOFdUl6DOu2/Jgf68xaX/bfkbA+fz
nZCggyP7ccaf76uUQyL/gFfva+G0qKdGA9PLjY/wIhYJE9U7HZCZxVRa1si4upIsVmUv2zFveWUi
/Ee+n2cXHJ87+y6XtsGOH+drybgrC9gnl46hOXJcpk7ZwxLjiy3BHUCbYb9chaWUlT/dITlwB+vm
Xc/s2qXDsTrJ4OcLGYcUmKXClnkEVBw5iPbEpjO1AIHljrm7+LhbEBkr0yBsvFAX9FP2mUWfhmyx
VyxRM2lE4izyPAZOvyujwiwR5/FijaEJelfLt+X+IFx60X82D4wcERsMq6LnRPVWCq/qGsPgG3nj
XsdWa+z/qxVo/6ubasrW5y8VjUcvK+gzpE6mokAKRSbQZfUYQ3oiJLThu+c5ZaAB9KaxOmQhRF1Y
8ur6RStGmp+HeXpfKO1cYsvs8lHa/OqHwsrWLWtpot1pHjYfINoLR2W1mdo9E645SQrgE+HWyH9i
zO+XiS9praPgNS2ghcLH+t/geJb+Fl9dbAfkgsb5ABg7FmxK/BagfwasvgxvMrHAkjLsX8xBJdHP
iXCRz53deNh6lf06rc2ZtPrXjMOwkPd4ar+z41yc+Gk2YlM1CHgHIWE+nVqOua2DlJhRcu8SrGXp
UByGlwYZucVhllSWB2Yxcxm3M2wjaJuIVBTlVM/FyacreIJu9VRs+y4kfdaa3GeIbY2OgXcJ39wO
U2S48/e3YGnEOizOUazJ00UdrctnOK3rfu/V0s3xRD9rPeQ5iXAUWS8tzrr/+wGzXODzotUZiQmW
/hC8ToBloF52tW+zqYemQE8K3QMiyYFtT/XYzp+968W5JESyntHCrpN2y0MhLbPSoJO5yRfBYYK5
0CCvggWLnG6jmDE/Le47KNRLJzHPxb9h+GVlJCGt5H84QB2+D2riNErUiEzShwSb7BmTbNgku/EJ
6LIHHC2h8e3MqyBdq7MwHUxAIEHTfqPEMTaapOAWPCwTqIetgBFvXmHdHLck4b3xq5cp/3917PMi
UBe/5qYdUYm5MtwZjyuGnMrYFFrYKuloLjtHfECeO1P9+Ury/Nln0g8zuPUBQQQaTK7j1YJRnmMy
SStMAmaDIA1ag+/M4rnfkEDAqJQ09SmK/U1yGGbFR8w84wo+y3aPt60Qsl+cxCbatg1t1ZxGd5jd
0pbcz5Um/m37VQRHM449EfBnuL46TCF5FqpgpAKoecoKH1p5dK3t4k1SAgJHmAWEVCbWMnpYSxJW
qIoVsf3f5Kd3C7ybjxFDgWo66c2eYw4F4B7tIUY7YQBz/lYbz42TMQ6tL0xz0M3ITtlYRSKFU9wo
3QgUVUrXBzr68qmQZxXR3F5Ju61nTQemJgBi6FgbZNmemCHeRS0sbxFlgCblloU6lmHQQdjDqw98
/YITcCyMFI7JLMvkCfafTMgNxURBQPWQpZWx3JWDD6zEvbv/uPLttSZqUyUx1qVLmZRfW7hj8a2j
X9PRzBjuncvnYJTup65bTG+7QQdHW+yhOJD6WHTNTZg1y6quaYqxpE/fWGraw/gmlr7t6c2Oq6+T
9Ymr/FtDpcunencnN86fdHhBY+52UpFCnn1UrCM4HkazqLiiOeT1JjJIFGsCMhO0z0EAPN4ors34
AwSkcEe9UmehPhBnXYosFK5RJck46qI2FbG9WP1tD9s6geuyytbbpe6eulrRnqKFn/AHKt9n4RRO
hQzPKSI43AwJuDjZACNcON6Rlcr4d3V0NxUAkuUj5c24MO06v1Iqe3vZLFbVJcV+YHMq2JHOcdMx
ypk+gDUP19Vsk+LUuXcGFmfR/Ub5j/2qCd1xFZJ0hBeJk8RAYmHKX6z01cmPFtoD1BBpPip2LCAX
pShisDFtlqZIGW5ad/+2dc+QmGoxsajXDeyjcPBdgdGqXq9+FvIlOuQUU941rBuKetZejxsPMxZT
DhB/PE1kjnTZGF4YlN7cqv2nh94msTlZqBteyjyE9o18SRfJh5j+hojkuBXevHIQOpicaiQKj0ko
gQ/3gFXnbI4y8qBn00dvdmmqEHU2M/K5bb78eQCH3N0n9i/Qy2ArhL4D52ed9rlvBmmEN96Oadf8
Z1j2W45dO7Y1H0yOFtTCy2P16YI64QIyfg1Z52bXBGhKC1p2+eIeqq1ymDfMdga/1IjuCtExp0V3
psx6iRK1DQiAlL0kGQC8eVyUzYE1KSOLuUitxglsEpgEzOQUeF5Rtvvqw7F/qvECN7Da+yQ1WUWm
pB9zKpoEM+atd6oHDTGjBEYBtjdhlmJ+VaT9EhTtJLEJ2wFkkthTNBYnzD9+gA0IoonNot+HIeQ2
mT3PNbHTZi7Z1riWw8YAGYF4kMpoEuhdVHG3JZwC6FsdZSZjy35CuFTN2Kq9vcSx11hYP3gXVCOt
Z5G1Y3B6X6PuZbZBrn9FldRW87E08zQvcVlFzlY8YAUScoGJrT2C5xArxacV9Ah0bGks176Fp/e8
w/9BYh85z86NBaJ2hQXSA0kNJ15h8RmZ+vzPP1CKOUE8qMGk/J+ScxQCEHDOhjImgYfLKWIRHN2J
GZqH09b2OLa8eAF+1UH3bPssWQClCVWf3tTc8cd6Ia7NN2ULOfr3RLHYqEoJFjQNw3Ua765hDjnR
T2yrY/TnKzoVEbjffQtkTPFO042keFUeYoLWA7U2QxLHgan/oavO6XeThtx6FTbypWpl/Dcx6U/T
ShFUFV4aAkqzAtZvdzRxOxZaBHyWuDnMk4MZvlq6pgqxGODKjQRmAgal1iCJdQmz3tpL/JJu4IiY
SKidIyGzLOflwmjvVrL0C9MiWgd572Ui3HCDSXlVfLDinih3/UIA4GlkeEeXflFxk9VFoGEerzkU
PbDWFxXjly47mudgP9vDcFZejFTjXWdKEP7JZuXUmRcN7ycD24IxVyr6Q7M6xFlTy2IpJ7Y3TDl5
zu+QPWw9PSfBkfTElyPGb5EhUI7GT3RB8lyOmeEXB71QNEZEjyrorB8/4YQeCHy06iWgvTvX0cfq
5dzpq3qNhcZSVKhhw5Th7ij/xJi1dRcQI9tl72AjbONPtVoWZxs/WggY//9lBbiqjB7ALYMMehkT
b/jTEt8Dy8JZtx0/ZNWQeSf+yriEuyKi1cqDOP2pnrZhMMgSaxadIoj0M0XxyoWYY8WSBcSYtwIA
yvV7x7qhLYEJ3T1fZGLEKbYcE7eRheuFueUNBlw8mdMLJ7GG37bWNpctVCE9FCCmI5zvAzAdibtj
uFwHWe27UHV+ChAURnl2oFKVHkHfSVpUeLJvlDde2n95OIXyqWEozsXFzC3JV2KDaZRWppH8TiEJ
Havf1v0pWXVJtvG39T8n3HRZ5tuZ4ZtfzV2uQclUmDEPVLNf10Ov3oy2aJ535EHTjbjw66LHltJ6
+jxs3W6C6OO2wRkbgznwhrxkZfgtFl0ucqlyHtQqf9slNU2jF00HnWqhjInI6W3BbeEZKBjbS96O
ZSX6v/IT/EjJch6ZBvpJlRGMSJK1Az/vkWHamJUc4A4iT0C9N0qntqA3sdXL5E15Mh7fi0D4eBD9
wLmL9y2713MbqXF8FHeP9mHWXvaonL+0JxTuFeNg143fyXRo/82z8utBkofDZ4IxnQqU24ML5YuD
Y1VFwu/jo+SDx1HXX8uESF92EkZr1xgCOOXnhhIEQI/oi9vmWmoM9rqqETM7tcoflkdgrXfpMCSp
D6f3mM8EBUryTN+oqLDQlvCHN6EYpM6lUDG9/1pSGw63JLwD8UDzNuYAZy+H13N8daWeWRjprJPR
drU9/dkB7+9+oHB7Rd0Btjzls/jWztV29ByOY8Xx2otzFg1HCe9xjWa/ncJ/4OrtJzOf1qNh1/hu
TfICyQ0FI2R4YfUZN5dcighhkQonjfIjFy1fsXyrI9tTaQ3CA+h8shY/V4ZJWy09WYaz2JbJvQ4X
qNFfb5QmP5PRCF5816uVlGtlqrRdtABMVRLIgsdjwTq66oHS63Eh66TsLfdHmKgLGH0iek2f//tv
HO9LOYuJQDGWcKcJAHP0s1laTaMJu7lwJkslwDBYaAQn7xYUisUy9F0FJDGKeH8VkQ9qGOwpf4ra
g08x2I/m5WLd+ksoZfmuZenU4Mk2nTGJMh/UBnrKfoxsP5ozsJOVefD7lmXdUc6N3U1ZNT0gf+GE
njwiu6QHe8fJTbogrkRxeb4yoQdVl9PJgqGi/IuO1EcZozrjGkLIa4FhTJQ/c1jE/SKRkE0Yyfia
14yAEAWk+ZaaQ3tW8yaMo4F2zoSJ0kWKU+fuXnWf9D8lHmArqS3cdvQHtjllS00rjEfi8NxzjL7g
3kBjT3yn4GscBMT173OeWRKqDAQmEeuyRaC4x2p6Dmdf2KIrzZphGWFiJcZ7tHo2GcRcVoCB0+mb
7rn7n9M5dkNQkxPLGr0xG1N9evwwjKV97crJsMZsaZGgP9buYfgIFx9a9c7NN3tqRC1M8aID9k0j
M+eQURIqSqPo3e95QZq70KD4pYnANHEvLzZHXpDJ3Krzl2TYDAod7B8fWHpuC7aSUgFpPwhBpdSZ
H8oyGXsYMfskwGRBhFlsfGxF0pDHeMpHedCLaJ75EETh6xcn6kLVHfCUggStpRwRnvfEhJ0AJWa8
moaXvtP78kYf10ODmcuLh7meRlHlHZKcn1wT5Zjl56IjpcjKDRZhU25Or6QU8gCkBD3s4a4aBiug
mLPyfWOsfnPfq5yO6MVSlIkzjH3LALdavokywj6MFgyBUkjGNVjWwnPHcsryoZHIUd629hmXEfyA
J8Wz/7e7Ki5+D2iDw5g8XS67UlvL+5heZeZQc/KPOXPENeScPE4FS7Lu3N8Jurvtx+rhpq2iyXsM
fD0QikqjW062kBfMZ6PrhdC8nC1AaKiGhSUQvWlS0dxPelDqgyTv/+AjD0xesNciZhdIeGvr/7WJ
fxr0QpKYOh6c0LBoqRa91PrFgeH7d0Yfo2YClVHsuIrwPg2T+HCW6d/VtoG7oZKc+V+qcjR9fMTx
eLFO8m2AbSe3Wp+kpqAxnO38dHpWea62gLqnDW/U86tBy2V/01rUxFNH4cniV81IgbVMqGr1Hxhp
op2HXRSVRYLQ6TOYVwTRC1rRbt2F9fKdFOIbmBKatDXq2SKFOql6/sVc731O3Lwve4rsikwDsrDh
3Ro5dbZkwDqZq2GcxbyebtdyzNT3qUWnCUEulA+EbmMST9N7NY74lDqJm73B7frJVjcVtwdNPksA
fwpRGL6bVNwNpqycBWqcPM5W03hQtvN8iGqWM3sprsA98lvtK9u+KAAwGRCgm7ZUGboIL0sc0XMh
0dYzp+1P3OV1BeNcIv0FwyoLWmfzid5dWkEtsro+N0Q+5PshRGRH+rI+TAvpOVCCu1safqbUqHQZ
pjGkfyhyOBDPnFzNpdaDiWuvswAM1LV1oPLSWfg5891o48xdSfiyL4Gvc5Pj2gQZo0B5BgexVMUV
yVCqN0ZapqDbZ062AiDR5DQ1y4/34vsSBbAV/p77+jkf5oz2tGnYJkpByv3iRybX/+qPdR2duHIb
Z1OmUXhQOMq+8btp+fiFplFngN2/usUKex2aKTl4244cVHerXkVaEBC9nA7+/O1mqijzWaY3XT8A
6suxmYN+7XWrtTJY4tu7+Rbl0J7ik273fuMApLD9fnXPWIm4ZO0yU81EHWLAKkw0nxQjUoWJxxOB
R/PAkbyIZ0LhxNOCrN0lTqq34w9KDSL3J//VUeyXbVda44XOS3jJzIocuyoFdbO1ssFH7wD7tZvV
afb2bgzbnWzWLSW3ZNqBqZWKWEkMINbZ4BuFx+HAIpwEt9DNnrpr6VYpPBc66nOcH+0AkkSMQ2ih
DGL9u/h3oaXnnvr0HJAOfJyczQU8db7aXSzHGHzXPwF0HrvPrX8usHJ1D+eN6BRlNcQ9HBhpDwXK
7TUOUaXMUj9ciKAu3rb+RvPs/zmnW13ffvDbpFW69/it+rPDdiD6IGuBn1YLpbrVzzAatim6H8WY
VevAZmuX8Mr6JrRR0L+JGAa1r2u2RXZmxYE7XiqMXJ7w5fveCBivbwWKD3jTVMhY4OE5llM5TZkW
YQ7F012g9Cp/pnFtCaJpiQZDegPzI50FejrF7xOyFtFrO+zB1EaOcjjrSyk+qULD+IzCAOnAN9OD
CE2zcNlUIzdbGKzul3/tTL4km/PDVckLTsM+MJpeVXv1Ts2yS9gtz7oiDKz/4nrYjUkCqebdt1r7
ZWfaFlmpizvQdrFLIwDf1VTEXJ+8JLXk8priQKClOXG8ZLHE7yaXCV5CmyEcgfNFxPmoG3chUEmR
FHesp9bO3vtkn3mb2ZG7e3yRDoGEsOMdd1aQcWBLU4ltLL5LxmWB5YuDvcD1VcifMKkLoM6trPFY
yuAR37lE81TgDvlA58pxfgdWt9CSzjf/zgknndFaPsjVr/7NATgvDNFc+ekQzBZ1Xza+bOgHhVVX
V/UP8jYrDrAyPzCZEw7uLXpoBtlnVfa/cuySRk6z9pDJ0Uz2PhaaIdobjXB1+UPvwcVnh1+E25Zw
wtgm5g96TYvQJCw6XvBrf3PrCGz7K0Th4f2AgzBEzAt0z6p8vBDBu18BgPGxlrajWmYNfSyRmBdv
H4tvbsQMuuLs1Rhe6eALVfevL0hY0l3ibASU1Yj4e/Ju0JGTmPO9y6h3mHKPWlJSHVGpKuwZSXWr
s6ZZxA8xqAwD8BCovV3ImItvngjcKYnunQbOVf4AISj310gYoL4sOLVAlWp9sywOebmhs2UTWk5w
0xeKoyfCQ9RKskP8QlN3XImDGp7qTV+ewDSnfK2Z2JotlyviwGdInrT7rRNdwVmti+yBhv87CtBz
LWF1fh8uD7H4PbLf5Wmj88UOh/NKheQg6yMRUaFpzGwJADPBxShS6edu8E9zRZ8BKYu8ApmrIANM
OVb6IsTUXIH1OCkXb/FXoUXZVmjTfPw5TOnKFE37dEvIjkNeCo7Gu6ZnTVecdCf7g3aiV46Z4N3y
0JR03d/Uvba/0eN/5hYiLSExp++o++gvvJvqbo5+lQ3Ku5XCAEd8jE0G3EBZ4A8XF5QgJzND0pEo
FzF8NFV1wuu+W2HvQo1sVZeJU7X6DrfBYbaGVZ78Cth8LyWfpsA8CGldMqS+0Gr2lc7Ljfk6HDNr
KYki9Grao/kj15VLQFsA9b7qZqlHbGL9eh3wSoC7tQgvJpAaRByQQx4kr4SbwoWQK56O7xivjgHQ
r/DstcVfR9tZ2kpgpfe0LBW5Q7kyi20OVrO/5r9ngt3gVMzhMLJvKRg8O/YVociVFkMGzb1H3YPO
w2HyshGLb/GeZszBmWYbSRiJSMYPD5MInmwkndUBKF3I0kaNqHGOIVCY7Q+eqeIMIRciLmowmDya
eKFgbiOJFIeAWsrkXJ/tQR54Z+lxkjOEHPwQK8gwQvYoOEszk0Izz9Kq/UaAgCSoegQDgYMVP34i
wGGcR5YhnqxdEak8lFWiNYbhuphGAZDfnF6wVKWzvWGGsf8/iEEHvlPE6ggBMF8wLTKVfmbfhCcu
Lc10BZf/6wSyipZiUYLtkPAu0gCMdwNaox0UPVsLuEX4IohE7Yv+2FYZ7Y7O/e8Xndx3YV0cOiBc
5mmFt2OtrABysVpPdIKnKyEDmOGcfmqOCWz/hhcuikiTCXsz0MwAIROWtb25xXs1Q1zSB6WE89V6
9MPJg8v7twsfLVHBPDLBdbVbdF6doZn3qGfkgKePq6QtR3RQPsSC2dGvihKD1DD4JBfDlI4WF1jJ
gku6BColbgjRQGC0DxPhjhws0rLpHKGh8gUVMcwNfKM76IGddCOq2P1uZC7/Ml9ZOUWb6jfXrUI4
y2PXTWnqOMqBkS2SsYbI2dbilyb40+X0GrtJfAJx75YR0OvOGw+pF142gOOUbiGyY3sKiKyaegx/
82rzj0dqBeMZ2K2x6y7bqpv3g1DIeJu5EE8tQgF90Xl9K0H8tr5XC3Y9p+/cMJB9DnBTuDvQSAYC
kYyjIC7RlgSBcdJV9Rle4iPHdyYMRhwa2cGEJkrHfAZ5qaKiH7w3QfRGz+X1dbWdPDA/ZKE9DnU4
ryyogYausBwsskmwJEyekcTwk1Iz4Sso+J6nSbRUTOMLbYBIVEF+eneEvvvGiNP8sN+lMBvOooIc
lO3dd2FbcA06CKdIlneBbRRU50heHqt0bVDE6EGitA8h5xlzd/UzHWLpKeKYf9NXLp8pNiLzOq/g
66pbnz5WIN44e3F9D0Xrsxp/IIO4paoFtgeF52wHLYlDc/j7CuA4AZG5fnCcMCVoVcGxVijvoRo3
Ipn1zQgORW7l7wha+1CZCJZ/or6ssfPcjN19b3T2QqiQtHNkPgUH7HO2DNbk7H4HovUZICuKeo92
AbCP0sy4VJfOmJv/vw5xRQAvZw6HN1tAQ9rMbs+agZUEViD8Xup93sNzPZLDVxkRjTZYU1Wxtu3v
n100d5/y1kRxOza1bcdcb2VlY5/6LdRFieRsDQWRspsbBsNjn3eUFlLA4HWGGM/4ipc0eAK3G2WX
Byy57IFnFjwe0S+9nMD/n77wCXJGeA9X3meuvTupuT2gGVhVIpG1Ziby4olpT/gYoCFMdvg5sHpP
lrixGJg7x6+rfnaRCFPTthHx0udtoAUA7CU53jU3ApiKiq383SZ13uaP8pPT3p7u9CVwTWuGpxdJ
aJQ66Dq0j/A+TJQ35KyWRzEopWyFu/Tj/8rqiopkmqfsNZax3CYVJpPbkaG+jvYYV96VN6czyeKv
nx2fmryCg8xzmiHEe8y6dOp1Kw98CMt9z/xlbKoS+otOVf4uvZxrclq6DMF7wXWObRyKVI+g/1vs
XNaolSbDV+RbrfC3bswZCaxG9jtEiGUht++W2kSbaMopRKSOpN1ta05QKChoslf7jTWAEaEH1zgi
Acrxss8NkLy5UwOD6uVBkdaDKtwNi7Stfkr4qKFPyjOSVfdF3VoBlZWnnLuJ+HgZtF2vKn+7DFnM
AvBhmkukGhg64+Iu4Gz+umQb2tjE8PwR75lvqUgn7xOXF5t55oob2cxXWxSNCOeEva16fJNIKZg0
dJPIEAswqXpI0y6nCT97EiGZWLR7zs1a3+SZLSABH2BqWV8YTseIx6TDQr7oruIm1c06QHbNfpMO
vysSgt0Lea8ffzr0KRvFqa4Hoi//srA/mPhxbtr3W/ITWdPEO9RBqxcpL01GXFjaGPBiXShJjK/V
Dj0lKRoQdlqdbO9LkSHHxKrQA/Mm2axTOGlzBiH4c4qKRbPXPWWrpiof6SrZikGK6pWaMRr3zfDV
rO2jr/nPPSeynWshsc6FoRNpMSiVrWz7MkgW6u2nN2RbPfrAaAGE4dg41zfCxz59CkQ0VcOBhBHY
1AGiVksjYdBPDpNN/Ttklhl2KwEswezZGrxNZBRGc0LA6+/NEQVPKoPrPSsHv/gWSXG7yU0iavSj
fxzdtZOY24Y1a3DjxXCODro2oQCp9nnhv1qQeXTkBLeZt5F/Ykbi+JML+SIZwFIKJTAscNgam8JZ
EZKl0JoR3pShXcPIIPLOheiyo652NOhZ3FnaCBnJAlxUAXAx3P15WA7fRU2l9CK6Fsy5lxT/I3m3
Zzd88JlmGckthb9RNRxK5GG62/o59whIXy7q6akvdQCM7PYGkrVF+l82HCi2yREsctqNFkhz7CB3
l6rUCcYT4akspCO6p16UkicLzzzqKufH7c6KVzugt8rX3zPzFtoiwo1BNQorlz6kXH3wgrH8LQ4E
TEiW30esw+zSDtAzDh6SjwPtM+FpaqYOgffyWDZIsFDingOR+cFykf6xm8DCrSGXwlJ78UFxZMXa
hEcd2nX7DglEJ6+FZ69kUGcVLsV8HqLmRzfPx6RVmx3PvGPLOEU52pdzlEjqPtg5t6OiPYVPGUde
DFOmG6XS+JDP2qlRJgmy1G1zTIdrUu9oEkWSzDnVDFBCheb1voynb/GwDyOw+eUyahWO/DaAQrbd
iNnv9ss+syZp+MkbqswHXlst773cMh0s3N70Fxf2HMEOswZhfbpdVa7NZU4ZfJfi7h6MzHnqqIOE
/1i9Myuz8ymgASQpMFKs6GAbvC+TW8GeXq7y6iHMf09vftzGRTBnlaEq7hX1mBSwvIggnzqezdze
tK/3t0BkoRFTX81xYMqzz9O5uRxnFqoinLZYJcIZkEBG5B4AZaRx+/IfhTLN7p/JROWumG/W6FmN
yFbTHiEs6SrjID9XIjMbyE/xwnioEnsrXpXhn48I9OZU/ArU8nkAhgf8qQ6DEC31YIVT/D/QiAro
+4XTufNAe3ZaX196s6ME1txijO9jlbvsKKkmVlZDPbR0O+ww28yVkt/MgrWfzsyHcrIhCW+WhF54
Kwi/FOh0XJ/CEv4NyXWH7L6/aM/lODZP0jvQTYo0ZN+r0oaJf419rMGrQ5mXHoIlrdWVKTAXKcBB
JkyLA6+Gy1YoEycl+CuIkeNdlVSjbtZTCSZzvU1dISBkbiRQdBFVRI/1Wx2a9BQHZ6FrNF1FLTG+
9WessruIKtT3SKC8J5pHVNSs+CkVdtPkqKIgA4iA6IrbEXr0XGo9mvVbY3MGJZt5+5+JD5UjEoYX
Mp1UB4ke2maEb1BpoO77HCtYWtq03oNyesItlH/o71brm35DDNOANT8jMb0LEfMXFTkEbHvyP004
VGpxoKvZyPW8xC9J36T4M9lWzjy+hA0D434Nx0N3mtm6G9nNzhkDqbVghEG4GAT9Y9G3wb6aDd4W
/OS2Gz89nf2oI9yVVRsNC6qIKj5slz8/3AfpH+Jnw3WJCHOt1yjvc71QV1KyqnOUZZVTy+3uNSiy
AJmCOw1pJgIPPTZnD5/kvOUf9j6Ssr2YGR7WYBLm6717CcknJzabeuPB1JoqAskAW3ikXZ+qJqE2
h/kIUE8zo3W74utkVXBrE7ZWs1AgyVP5soVUqJC4+ECbW0ET7UC2qRX+kPwCGeFqFN35K9tMaaWX
zv9fBfYWmbi9SzzIwB+5fpqChddTTyUczkmHcf7dAspzVH/au/C1fbDok4k/w9LAmUlKGwIFEsN+
8YbqNOODNtGUF//fNEr+zPhk9gfO3lQ7Z5BouUNIqAA1QNH8M990yoKC61nMnTPu8VSDwxWWtrev
HOk2WHcPJcGYWiJBCTvtwMOA66fGdkx9+8Ben41VXc5MtssblgXOPectpkoOLTm1yf4LdWAOoQj2
ZqiPrfdvRWOEG6UVOfqdHN1bGFEGvC++F/f6qgDmqxTiQD03BEtdPg7vm6HXIc0B7cWbfHXS4Eu4
lBVuuTpg4uPKrL4U1EQ6NvMK/8rPPVkSOwtX3FnE3smBjz3C8z1HBDYMTDQjGGjOa6ZjbN6E/y6p
crlDL0bfNH/Ep7L2v70pB8iZK8/AfngmZmVLg+gIExnHTzpp8v/TwEjkU88ioTjzdLgrzFoNjhuJ
yvaQSWevBfAmrGt9rio3hXkFJbRQuKnQg6zJKIpPNczWqicINhNZMDYbaPPAUWwXFZUarY9mv2PE
jbd3eoRkwu85tfmeskvqcLXKCyOojfrtRCTcgTO/BBoDWZSKmVqnx7C5JVw2OSnAKq1ldAftwh1S
rCn1aTj/adomNoPdcZYRpWyPGhflkCJClURvLikrhlhYZWHLXwMb7+EFjBruN2PicOB8ummAb61n
RchV4rikx1SYU2Qna8mYgSW6CL4ZDt76XfAqXWqb+xLtK3OVs+vKPLd46N1tQ4sMG6Nb1LyEZSxo
t6X1Wpkj3ToTD7h+CYur0zFKueN5fDj4erzpyjG01u1tj2DCNB6joo33HiNa7XJfdSqGka2gxCb6
kZziEpy5aI3XQ8iWE3ejBKUweG/wM/Eh3oSCpJ8SHLa803UPZZNEZrlNWluzHHhqJ0+4Uo3gWMXa
EDTrdNydv4dtShcg6CEMXSh7nQ4tUvAst1gOXsdRyB6a42mDvrtkYTeQlaakWXjV708OPmxLH6j9
Z0QavKGxV1h4XT7KtZK3dhMKx3x8PekE9YmC/Gof0AAu/aqSyQWIJNFE3VuIohZXYxp//uMc5MSo
6dqffl6rNOaeteLbACb654GgdPCLcpPqWT+Mekd4N6+LmSJBmCf3OfvFwHD1vBVnFTIoDAjxq874
uk5jQmj7nb+Q1bfqsxVmQFkza2tC57UutB/BJiRgc6nrujpOzW7muTZCAD49KiO+1O9tdYrPDZgJ
mLfpkI0wEhN15znUJBZ4bCkwzHZON6u6Am8gYCZvwC2GzKsL78/4xey2cccHwZm9718bxI0E4URm
233QyP7sC8jnDc1KOj7b3oSxJG2KEihphzRz+xPa1QicUSA6QYEmbIQHi9rIJJwbpGgVByLqmeCb
/Ld+FbBhjrh55akr4hONkMFoX6Rt6kJ537M5Eg+RwFH9v7fqe0oHDHtSa5+HGhOlPwmMQ2+MHzxd
MXhGHsOfeXAWMnQRPAPoMAs0mb3Tp7B7a0fznfPz+8pgh7snkKcOO6q0sfK7ljN7wOC0wZqn/mkP
0jhTh14jDa4luJoiFsHZqqT8Ix3ACEU4BQPfXXIM8eGUwldS/+EVPyPyKeKxlMdjvIGxBH+MOo0a
lN7AEYvA+aWBJhyod15zE7WthGpOyF/IpMgObI0JHOxmdfdfcr5e/G0OvVDqehhVaReLLiun8mt2
OF96GS4xCFy63dEzCKCxG/IJ69X98E7Zr5UdbfngbXzhSclzGea7gsmmOWuVZQJWU94xSer5x5J8
/MXP/pj+v32SWo7J15ETxeLPnwvWM7mQHsHLKDQmHzAEdplNZblIej0W/ZWpjEpL8lJU0+K9QbAX
UnneJC1TuFj5Rk7z4EOW+t0thGFnCcuxg9KPXm1G3UWJFwADXuQDi6e7OHBD0ogRv2LpFltyz5mx
KDxzNejEFXJFmrabDSzxIfuoz+EE31FFmmXUMSqEorbL/a7BeZCgzgRdmKsuDrsEogMH3znxmAGq
l+YchdKEKZ/ZBnLCXgXD5ZJWwad2/Z+nbBWcRqAFGZOAsHi04db8nJiMbZr7Lc2DKLqW6KmfO9xD
bzYKU2VqU8Sz6ciad/ViD9BJqycuy1NoWqQGBzz3KPWpekoUhIeJ7G15B4zXc9C/nXj0Km00FmS4
u28pig+OsyaEIBLItZYfzykJYK2i1sD4Wk06ZcdoOBlRmHwlx4Q5Mc/ItKSCuQdJ/ivaVvFQSYb6
pzag9JKimxyB4POxM2a3ndHeGmmkOAmFokXuSt+dtTo0++5a5kl2rPz+DNyUe7LoQTWbwCMf9JnC
50Jguuh4JUhSxiYixwGud8d2x/4Yms3Uexx8GfLX2bZlH7jKxz+kyCXbNYsjMPOQSfFyoBT9dLqx
hfC6/nO5D0aAo5gxbYGD5khC2QmoBHssBsU4klzAYYSedvjBu6jfODgqHVaOABmHuTjkUghgcxUV
ihk1+OVsDWP69om6BnMTJPxj9PfOHzIEN8tcfGApxcecnsLD73l35NDGY56G2wY5YcU+wvLCxmJ2
QUdbbcEsdxPFUQQLgmmNSSCnyzsMCoHR+X5guYSpRTMu9RO4UBPsJ6FOJYqjrpv/7F7BHkXiy4l2
13CPiictqn3EkGUBtpCq8TKRBaVP8c8QYVM3u8pX9XEZHA1+GS6g+xhQUuztfJLD8GZeryY2Y1sP
YiGxc57CRSgjhHvm/ax2vAZp8Gu/u1TbC1CWUnMgQHgp75FCbkSHFoQWJ0+xrYXYcn4d8nL0r9Mt
89Q0tQGwOS4HyiZzjoCO7jaUjexcT6PuR0fR8PRfxO+AeNdky2NukspKo+6Yfo0AWCXomzKgyZwh
/u/gnG8AVBiVgudxwCn1PF49smTQbxidiAlLxuOAZi1LW5m8mqHdY7fkJLR+sv8X6OjFk+8sz2u3
z+ODMxS9dt3sUfoe49Ql8i7H/JMYm0im7PXRiWtZxu/Uu4lMZqlryJibfylQsfjT5zvbolROpt61
OWKYbaEXIr3O07iXcj9h6n/i8N07y4pzDBGO3VD1xTKbQ/LdCOHvzItl8m8zI2K2SQ7OB+M/XPi1
5zSLoQy/u6Xvtv2HooY6jFuskxXX6i2j/0t91KC2x0JT4fgCpB8S5TR1KalrhG69kWT3vpAfDreI
gjtTozi6YbvxC1sz3sk5y7npBAHjTM765Gtuku4DW0c9lotf+42CaMNCVw/d4kPtFeIgp8NI5Czi
EjVLhSW+7uMk1oJStxrC6doBFF7RiY8ZmAxkGQJK2khgKtwOTADT0Q2ubxI4OwT4jAHrl6G/cWxa
WwpWaAnpLBb+ZVAdlMG31WTQNWkK0ueNnYEoCjna1vkYjxVGMRjbBTqG1yD+EAMemZIYj+5GpAb3
g4CRQwBYgMAeAEoQUlK1PQN8qxcBlift49PXkz2usTbgQ5A9Ohd3i+wqNOgNO+VgnvPPSCHfYN23
zoUZS2uK31hIKp4As2JvA1KI4VgqdPH2SFRQPU07vWcs/Qa5kYeKp/SznEGvbyWyIiuvGdZBHO9B
WUnx/tMYxkpg5f5JWgRFMha6701rI+b2/yeC9AYwfpP8rQhWqXPK68cmZvOD1/kTy7JHZBHnt0zM
DJQ5YmVxE0VIFPByOo2cS7av8P39KvEWZO9B/zUFLqHwwe99B23EYzrzVr0m792tb9VTxMOyhHMr
7WnqpC3oYyOARYtzpCE3Md7wbQPXIT/FXDnmxKeMlYlsw7pdw1QFnyzsvQS1ahgpochaZ5PMPMvJ
nZpHpPgyEpybnN8CHYVa6X/i3BTVwshh89BQbF/dqX+7YhrGNITpfDyT4xV7RTJCZuhcrHGyALL/
kqMBjtyJfkdJe3iX075Z/lbG5Mj4wtJwn7DMB33Quv/qARyv91YBGoGLV12Bcs1wRs3MGiNt3MtB
/7Q0CigSXCnlO3tspyMan3eHW1O0eZNVWdJFbBd4HJtsDQPsjZ6NsSnqpMTOIaLYoFQNq3yIF0gx
9kO7Mq/Ax/R2dL6hor3h/OQ9Unz8/msk7bJsnPW3H9PLE037FHy93x3GIjNIGmAJnMyGU6mpGd3K
B2GHTx1LeTW/EE8t1e3k7qw+QONQb23Ehnf7mDZKFUi2q0KDRP1qH0aNZeVPxVdtIGBTD0iR1JJ+
aUwbdAkZaGJo+105pgwAvZgSO5SAnyV0fK+12IZDKq35JiQpllhjIum+RtzwLIIGmdmqMiLF68DI
wiz2Zyp4fIUIr5aV+ga3deNM2oiY1SsJi449zRK2mJyjsAwtLWVf+Qga6NFheV2UvnvZSzMMELUO
f+G7w6LuIRbLVXxLUxFJysedJU93AhHZekomi74rS6qpa53upLPZGMiGI+wQCreFJ2ySooEhkeJL
J8WzvjWmSnLSUiPrLpD9K4Qb5DRzERYFg5xgefMN83TXSVBVjFH8g1/tnMUnBp2INQXJYcOuYDuZ
dmM0UqI+IfqtLce/Nx+XXHbpBy15CUIn6/nsUvCREIrK7eB+hf0FuXaFixnH/ecEZDLrg+GYGU5f
ASHDTbBvdaV9iuZbEtAFgJHs/2XX6wzubO8E44w2RNLoABrtkWfvmv/Ib3Rr/nk9w8w75Pf4P4cc
XZ493/OFE00hjTE1Af1ok8SgMKK4PCm+6tHb5V2T4jy9Kno13KHHdxu5loZ5eFvbYcsUqfIEhYuf
ASOxIm7grBE+ANcJ7ems9XHIzzQw0pNDdlRCPFUJ6+Mu7We4p3a5ekQ+Kx4mmWq3MEPlYr5WqCwH
w7+HyF9sDEpbwbOGCJeF/NvFCiitRHxiNC/ADvuA2RWS9sw7Er2R7iuXvt5mir2J0WTxi7OFkA0a
udORd6T1i9znCHZ3s0NJO9r0m4+D5DbY3r1PqYzpPFZM+4nEkt+8cC+Yy8XAk3lh8e/NPvC1EBYL
pgX2ITiPdAOL8c88HAkvIKybkn5n/pMpz74MMXnWqn8vHmpLJoUg4XHTPkcSZYcvVjUwL07tds5A
Bq/W4Y99avy4rNKBBCSIFdol7MMF9opqgOxXlmfXIZccSf+ZahJQi9ZJzoCZ8ucw06bB69qizpI9
0VW2SMHNY8iAIrmMK7foE1n6QpEsKxIrxs9afvpHFJ2G/MQ29lzKfqJegL9xFXrnMWeyLx/0V35O
kgRTPNOrglvk+gcjPPj1T1myw9sbFCabofiEZeopnyIZhI5VMdEExJPdTerU21JX71vstpeKzgED
Ag8pN7zSQnQHJ5njVcnBy46TicOrsxJeo7uiPbamM+lEwK2uirJiLcpAYhUqH5PHUDQjHylnNJ4I
VXkXU20XvmhVhw0o+aC5a9cuW34Kft+G/l0CuPiZ0TyJehVcZxTlLdRQHLDh09s4ujat0TTSTAV0
8Mtkf3WyiNdAV8xsiqmGk5crpgRy0dkWP9u3GuvPTvfqZc8zCGvwcqduhSIzWIzAWg2/m9aB76dp
3riz6t1AZDf67I17EhDKtocWfpWKo81Hvy5CS8YtBaWa0ShWzttSmDU/6MB7Wr06chfsqpMYHM0b
fg+azJIKRy3p5XCaykAVjAZnNKceyKuNmhBgGXlSakL+u1k82OP+V3C/7RuJuqwkCvlHA9KggA28
iZnUxXGQTTSESlmEdxMI4xQ5r4JBPTuNcqMUD5Ul+RD4gcYtb3pCR8tMAN9BvR5phLVOZL5sDK8x
1eIRzJra92TICgxPz2X92vv6UgviMHuWJBhpcBof+r2Ty+PAaTpWH+Fr9kLgnIuBQHd/ydtJuV3w
65vGR2vlfi30XFj6A9sbib6mGiYeeHpmxh4l403RfL4mFK+IHSQ21Hb5q1FAC9NmQ+672dH0v4ha
thG6uxUAHScXGocedlCr6pWjiA7pNwDJ+cYYr8n1LB0zQw7ICxW97l8uFAfqj6esEkfQpQ204/3o
A1E2zYO6mnb68zx5eSAAk4QhfpkyFOx9YLg3iIMidMd9CGv//JinU5Vn3/HtbmY4/m+lJEGNjSng
zlbgQopFFmrM0icQXLecjsbIaK7pFrxZp0+gnzNAlAW4wcLhnzZf+Pz5olxjFYoLQ9V19vGVw7Bx
Do5RlbBequxjaYkR3CT0f8/fCf4RpciFPwAvbQdsv0TRz6dVO1sUaXucbxocIiXIEo8ZOXSbxLQK
1m7oDiv45eCU2ctJR9CR+JmJckDd6/b+FQk38uSmDvUCdU8M3O6slChP4fyHkXaLTH7KvsbfCY8t
7ASQbVX7cXU0jP0loUMqlQj5OISglIRqbwheYv2KRLKzzJRrwzT+ZYK0oJNhMyxUEaTCHtLD94rA
Ky4UY7AujAmCcg4pPd4jyzK1OJ4zcArdlAGyUsCDrGGKyFUnAHddK82efDxboIxn5lqk25nlq4DN
UbgsyiIMjR5QBalWXXN2IRsPSYM9QWo50osSoW8m0N5afsIz09GJdaPSUerXQLa8RrHRRy3zMVjI
ZzHmv6CyV5vm+wrKIhRq+kb/QBR+9/CnbkA/EjvmveWuK7kpXPJbrvBbPAGlOPhpjUQewMh5hRmh
Cz7seDNRoN5lmQe9VZiCmJNyn58GmpfcW6RsdIM+aOITXdJPtEx5Foswnczuu7WCrTT78yeAfnVo
FuFtlqdyW7slA8JnyMtg+BPeHg7hnX2j9EyfS8rkYqzCQDjzk+n9mWeTC94EzPQbnVS9vwzcH0VZ
Co0RCAzm62M++6Btxg7Y3TqiIv3vGTCwolhqoMM8PbFsPnkELYoCR/gPycKHuXHF+ecoP6tB9Zna
ky08w87mlp/zChL045G1vib2jhN21ctmBQhYbDy5iYOkjWbD2zh5OquLr3EooBYehgiixb7QFglm
NU2sMFjgZs8fAN2Vksbrx+uTj9np3TN9Qkp/Aprf7j5Hvsw6elb6LHC50VloiuZVkOYrSHe+LV7+
kk5IfB1y3At54chjIRwdwuhh0VWUh1WXp9Hm8g6tn+4yxvJn3RFhkMWQyA+Nj63um6lN6Gm5U3SE
ZBuTQI4QMkMu8CGspZABlHUE4p80goWn7j4CllFF3pq2Ui1r6ZBdMywPKB6F8nrgQu4oMdRe/+us
brzAVI0wnUgCGDDyqGs2q2Z65fIooc5VWudh4MVF/FBPKp4lVcI8gCPMiL/0EE30zvYSL+OXPWdN
+MTtkUypyRyEQVUCbuS+ZJ/RDgU/UHFK+Vv5lMfg4Bmk5TmHNVYdHto0iNhPhJfRrmv2jBmGE9pT
Quy0FL8xM9bWLttS0idI0+KjKTfzSrxp+uvTFT1AIdilqzidBalmGPNm7AVHhewVEI5HLeq+dNC6
weNRMiC1yyJv+/fn30+uvbYi5IpmKxQJmJSOh0ij2RTartCOI0fbiYvhU533x17ATYDD/6WEK0BB
HCLl5Rx5H4A/1cEFMkSdHjS/WxpwsCE9rL632ms1kiV2wX9kOytYB4O0KShuWw4dQlTtx7PqE9PD
ng5v2GIjDXMez4fCXf6QTdWxF5cdfPYn6K/ituTDC60aa/9quyomeCPvhPXgYVD4mOwliSyVYBMa
FTNKwUSSmXIIU3z0ztjwhzgD7hEIWE3IQmKAM6KUVKxUQMD7G0rtQmwyOptAzK6uPCL2bxUijmlD
pQ35vy5RkfUU6TfPF2kBwJZM7ZcwZutijgcr0gCQv7SwIb6mLc0lBnGObd57d/5ljX+xtjmEdmaE
wyoc04ZOR/t5xquLwKSmILyx+nhvXXhN78CbmsJDYi7WlBt7XkifHW59m9dGB1tpQVKkGaTzlSw+
u+IwZ7yo1xMSG5y/HlsC94kxLJ8zdaZBXG96txNFx6fjgrKJELIjZ6sBIR2dZbl/NpW9Xkn7oDeR
fWalVxU8kNq/SpsBb63IePUQx7sTFtrJY0TpTjdqc9p4uKP1GhRVGnzOFzITSIpFeTPO9X59ZmhA
NzZYfjpjYEUCppHi6a07UdLDVi/0YOhCgYWg4ONI8p6ni00RvmbaCRSoDk4wUoofrGAE0SLlqlV4
UZa0npPTUk1JoFPMRqMrHDhid/g0+EspyZ9BoN3U/5oGyP3V37hz99VathWif//oyOa3JVIxZTCO
Ey1AhWnVfUzJp+N0g0pM0GAzerbwHeTLNIgH21LNOHbpe6WcLMLyEgDTaPZGLIcN7mFaJ1ojWo43
xQBkupWkv1A+yarZoKkuWmmRnVuL5SBQnZVQ1Qw5CHmBgBRKDEoVC9VLNcst1zShw1xgq8S84Y2A
dlnIpPobPky6CVY4VqN3RuZQwUDXqIWEKQ0IR2Mb+z74MvUzAXnk3RCSJ35bLKpX42+z71lIyjVh
Tid2QtsjUvvaus9mvQ1tHhPpEpQsKFEe5FFjY7MpSv6zeU5y0C66KLQGIkidOLRbVxEQNNAGCD+L
UQ6Pa1MVTIvPiz3LGbBJRWNgVM/Z9d60krdYbx0pQaC9SP7Ok8BAidImTekI5gr22Cf3wPGrWkTx
caSaATqCeuo9ex3XT6qEMu7/Lo2VOiZd5texkwBbpVz7mtfftZTrQYZ6p6CkYRO4SXGowyCvHifT
dfQr8z3CA4ojrhgDAAbiaUbUd83L6h2MZqCmIy9Uga6CMu8CH+I12HCdDYH77jiXH16SfFKSZ+xu
DOvDfECPlSWzfcCHM/CncM3/CtAzS/2RWop6Dt4HlKKALxlGRYzJ+t3ZjgdTqiekBMfb7hbQy3ne
Dd+m/jrqWuvdufFgUyaNUr1q2kPb6IkFeP36XXE9CP7cFs0vulmBFtzGq23Y6X/GveakW1SxC0o0
odh+JTzsC+VhOjgC2fXgu1mwDlz6FgiN8uhBL0PVRR/al7mr+pDvslJGVE/6DSPZk7HUtxHnPeis
s81lUfKSx4jFejjB5cwH4ERDF/8TF1kxBOseKJoDzigSm2PPLn6Nm0TwuXGowWwV8NKcieq/tfyp
4coT6pAs+6sZcVyGlDo31R2GHmVGQsyc2Cp/E7AmUB/ucRveawYpGNbP10VR9KKvD9P0jl1SKF5v
MO+E0d5dJBZv/P1nNUY+aRZNhe0cyB4wP99TjIZbxQ1i0qAKbNDmhNeMxQygY7QSk7BuffGoNkah
8t00RoAt1PPU65o85ytPr5KPUurnmz9QRCaLy1jKgy3m9gnQgMrYrOHxcyU+3YfhlUHmMdix/pa8
8Sx2SHeWlbbu6uFgmvtoi9RS703zfBM8HXRk07MD4qI4n220W9uvRM8KSIUbuBY/zXnHKK688p8/
PSW/AK1y66H60qAcXdFfd5iRZOI8TP5xsgD5vnFHevYWC/DJlT2ib7Xb5r0u35UH4FtBcSGWA12+
YH34mFqldJuVquyqI1X+MfWN0fH8/miSpDxUatDcigrpuyI/yjVdbf9B0UfL8ZB6ovifqy+qT5yh
fg+vZkmDAaA2RdKwyeustrHf/wQda2Z4obvUoHY7szJLGcedWdZRnaXJTL4BvJdn1LFDR2xdQIQI
Fcq/IXbxNNvviJS0mt01ovL0fw+VAamuwdnjzyXoImYkrYTZhigTDi3VU6igSJNuIeVr4IBFJSpf
Me1PndAwsbC7QfIUppHtyQhLq3usIBJcy3SOgm4EFQtYfE2zs0viRSuSUyb35pvLUQ3Th5nN/jKU
tx69oN3VUSmX2JJEEgp4ULWe0B7HL1MerKZhyGV+if56R0jYhUHh8fZ4jfN76B5z9N15oyK8yVJ8
u+MrTHrWGBZQUUtwndyhCLq4CU8OLKC1fWgJQh4zF4Om6XmmcmCN83YgEirON2PdzV5QMB3w0kqx
Ezx6j7BIOOVSw5O4BGe89FBxRjXWKeSPOlPSqGmf1tJOD12of5Dez0Mx4SYZNDXhtjhyC1ec8IM5
QogLmTeB8BsOqpiekvWjiKOBY5bvtSJhBgw6voZmgMdxGszc0QMpXJHds3u3w6iKSi6LT3vVOybZ
WzTzX7eMswiKAmOPMNNXiqR/SCj5SC8E8hfe0RzkS4VCqQvJnPkSvCzmZQzajawJGx+2CGhaaHhi
RvBDPytJpCPc4byepnIqwUszi3XKyw13WKSghY7aZXB+p5knFzu+tGy1iIXJq/clAah/G/2UKYgL
n0zV2R5fSFwLgI4ZIxC8Bvsq1F6lgLvndPLYUxPKtnok9lSKPddvyIePz65IPPXI1E4oEXlD+Sk4
9SApZpwjms+UBIbRfl0PS/KR2CtV00FKsMMbnDw62ol3uTYSaBtwkeDvFbA83q3E5Z/puw0Cy2tN
Y4Br3ZYItpVkNDm4AiOIa9d2vTvHSZWgSkSeSAyjVhgRLffftEFnjqP/EAeJROhGRVrUKtKjcQl/
MlcoRAJqofzbVQj15c6ibXxi5UOH91S0HAorCp4XmYuPtqpCvCpylXEjOwt2qGuhQqqYWPf8N82C
pAheX8Pi67i9KMF5dFKlOgdBpu6u6qF6r9bmCQHa31MCN6nXHenYk73X3/fB2KWeg80ps7qLhIPj
stYrt4KNiH0NyJgWTtEf5YDUmnpflshArdj677JIkSnnn7a9WSWT3Yh4XB+r81XSTUnj1g4PmnYZ
CUT5ks11zpTj04OQtGbfQBFAG9VfmCx2bETiLPPONxJsmQEKQt7jIj7EXmULTgCkXerqX9xu99Ua
9SkWRRBEp75DMeE5IZV7MMOslxyj0SDOSwfhGzXMaObcyra5KLxtzrr7VUBt81r2AQnFE7jVhzNL
3L+DcDhoh+UEGsMCj30Ulm/BV4IG/cHDkH5CzSecSgxVIN6jRyFyT1jr5WpBAV5192xsTbB0L85z
r5ILoVFX6lxGomqzW44UlMVUSDjyWPz5qT6Q/HO7Z3cOlkP2i8GM1QedMJ0E0apRis0aHYXTF3Ck
ES3nLt6WGFRRVHSD7cW/8ULM/quGlixocSz8LC3nxfJ8tuPoCxPkG6HpjinaphffvdiY8H09WubE
BF2WvbEV5l7pei2q/bE3IdLLoy3/mWm/i1J5WbfJ9Dic81l5h+TCeR2E+cOlPou5VZxOICaIAPEl
aOJmlInPjBohMa6hfb4F2NWOvrcSkcRLmA524QE0BKY/3qtq50q6k7cvG+w/PwiALJVFLIvZPmsF
XYDSJrGmWsBv/LR1BoNKVgOA+h8+ChPpS+DUmdDV2r1HV4IN+c3h5TC3hAMAlCrYpMVUc1gO08pV
LOBi53c/G2m0aWWtIVb5TTbamIsfm04OyExLD0K8NUxdGZRzW6GyqIZH2KTBnyrkPldxqvWY0sCy
b/RldPudWyFuHL++FByUGuaW/u5AmObuUi+mr5m04OQBSNBOUfJwGy1xGicmkszhBcPDI9XoAo7J
ReMuzJQS+Wb8msdMjGIvODM4lBifuttagIhhTqRZxselAClX+M6NdJrrk9SO5aHYDfTVZ50uhgrw
rfMaZtg/9laO87bHTbrica2kje09VlYgSYcI6iwxQ+SCOHQ4phcRTEHcXaAC/nMTMlkZ7/ZN1DZp
Qzh5K9EhLnQZb7rQDyTw6GbSC0fxsC3GZm09gCWgfXZUY8AcjpLf0y0WArF2uY3oyIQNW0KIpjA2
fWF3H07laBVv22tDj86Sq+VyqeFQgtoW9y2KWxjTf8DGx/aXsAJxvNJc2rIm9t56f0w30K3VVTUT
aMiDMyXHYafDThS8VJ90fArg8/lgK6tsC9hUytSjdFAwFBo3pudr0uRCOt3qDn3u66CILUxjdWd3
xFJD4VeEki2qZ6ebEDqlt6tSUFoebdHiE+EEHtcDqwAKho+YGMxkzVDS4k2BjdAwSgpJHZ218k5N
PaECXqUcBvjACEGYWp3hYYOhwdwtujHmSadrW7a59l8eZvGVIP23ZOGPHNFEpBZ1YPdLagBICl8l
pkZx7ZUFBcsiODkW4X0Sso4sPWa85rc489ZENOQxPGgfsYuTyTxtb5EwA5A2lSFqiFomynP9q0AX
U54kfMDCr32yR8S5ld5JfLjUCmBNXZLakdyK/As9zIrrSp8XGmYqr9vyhSX7hGjC2SlLrQOris3K
3GTCIhw9Rx2b4CdyFp7RG69a49idvxUIp1oyNR3zG5Sbn4eWeER02frduSXjfG/nUYN2raETqy2Y
FIq7TfX+r8+X6ii+J98oo04C/FJfufldkfuKG5KH5zvp5JpZcsll87BerJh00OYCx3hB1gfEj/GL
M81XlOittv966HhWUPXbHQyU17evc75zpbtrVoA4MtyxZ2sONs3/GOXClpg/ibqDsztBP2y81IYM
qTLzXAkdpNTRJW5W2+sFfO/cMShQwgNY0zcS8BrTXdvwrBvvgbBC1iWn+U0VhCijtXGYug8gjuB2
8/iMEt2VslD4xJE+tEryCppJI5+QK9XmRxlFGrsY8tqdQ3YUzk2E0mpshMnxb3x04d6wIFid06rK
ZaOWSwt/JfR1dUX3vC8glIDU3aw1v0ixKd3Mm+RJF9XkifnDIisBDaUAGBJxsiB042Y/FaZHcocw
KSLNGjxR64aU9fsAvTrt1y1xJwy+pPV0ys7FShqd4VhQ5GUXkZ//yERGYYumlIGEBjW+pOA5AS4y
h54hyPlpTEWzx081VQiKLLoAEb3+AB9E+thRfGhxuxAQdAx0gCzCa+21aEHdRqGIQUbL95XHPWjM
+OoL7rkx6pFM+2FDlfJ+RrMpSyqmokshi0YSX5joee1vyBnjV8N+OuZ0qxoGwqjiEApv5oAh3vpj
w3PMmqjFwq4ugEj+ykecspbgqM3Atfft8MVt0I7bGA/i716oJ3ZxGIVlv2C9XlnBKwJKH/JNrbLb
24J9rD89zaSvHdfIAk7zLxDUh3TR9iqVisnBQfPWb/7qgKcZwqz8HkCSQJpUN4/Iu3wW+wc4sbm5
3SlPFZ+QlsQVG8K8HP69JCW6S92tmyC30UWJcc46Dt59wrcyg+2bZvt7NtrLia1im0afrhLObCyr
yB8LfcbpnKa/UFoAB3CAnsCkm9jnSRKhvND/1HM/z0lJEy6Ea+fouyqd5VMOLsKvJhhDDObTRBB/
NFRW4Vl/5EFgCp/7VaqhxQ13cegESNN1Egbn7pFitEynsKztorE6ZzM+ESVpfzoq40VR8lmQL3I+
W4K6+k3zcuTHtwp3FYdDNBL1vBkHmr0llEFHXfjQc12K1HlUZG2oF0qoz3XlSU5Ux2R8PDYJql6h
H/KQ3JF+2y6wC4WW233sdPsSfGazuv5rmuEWDtFmPWoNLCCjFZRu4PDhLmforAM+RUld+2FrBOPG
moyUwnuulhqBuIQP5ZY3rrOJZrk4YKwYa/UHQkcM7k4yV6ySvRiVHvclWnh18vpOf/mivhqkSQD6
1CWsTo+PZPbFTcxTGfv9LGuqOAI0C8JbirXEkIHUNOSp5poqOz17ZjUNDLAdYdpqmztqsdjpU3yF
vX7eY2VwZv2TYwhCYsFO7O3XSNpyBtIHsjGI77DPvF1MGZSD8LUZjD/h5xavckB/KCkEPt/vB0WQ
0JnYbbhRGt5fxu0OniicWCMnFOBJXJ2tfFP9WMH/29BPfJ9JewtoxkWdh7dlQu3W0sP5TlGg08T1
G95PqiALOvb7x/z+5lu7ka8GWEXs1HCls08Havme286oz9uXT3JOKhf+A9L2usrcUO8Ji9nKun+B
zlVEt3qhrc73ADKURTCbxbdxrCPgexK9ePYYAmE/tWmz3f/sPlcBwntaJxr5TSK78/1mvC3Sh56w
gicwRoyUAuOxLMUr6YZT8Tef2DvAUmF07qhADGha80AhncUWc9yUTHBnfRIwcjGikW/JmkSRh00H
XsWB9MjLGTUUHpZ7G3HfKTZ0JqNVyd06ECZq1lkY+AkvTpjmEQhDrf5r8eULGBGX4a/7Z/AHT6YY
WnxxjWrWb6uPonor6zHptGxCVrPJhJPyxQ11WKdVLeu7AHLMxqmwu01meaZyD8GQ+hxYTjKnDr2j
FE5mq4XGMf52TU8UOQ2RYSnsQOxADsHmuL9mJE54DsfodGCBhxaiKzYZVkFjPpVaVs0YaQ7JmvuY
QDhRbj6Ur5xdtgmXf94m4ZPN9AB8WyikQ/E1upNZpe6mB8D4YpKdFNUGQt3cVQ6xUEY/f+0ht/7J
zkQbv0I/B/wFin1qaOm37B0XCNNkgkq1AM04z5NOYv7EZpWEku+NKhWBB40FHr3TrxTa4R1G3yY4
HNBZJ3IcZax0ZJXq9JHk9RUfJbMpB3/NBQA+WjmHkY0rqjzwaOpcE8/1ZlIEyzD3+g2OMbo+VdAl
51pZ2zf56/akEiL3r4VL0YDSVHFpvlvkR4y/J6DwM3qBQPVkccnsvy6JjaewalzZlLmAaE3ZqIBg
WXa/yZz9QJuR0L3TRbdOfl3ikaswRFrBK1TTTN5DrGmk2Uas+EV9arM8kzg3KuiQO1NhthOqtult
5myjSlF+rQjnKFKukKEpblOutGEj6ecpXdp4+nANRbVB8uP6rcKvLGVlGNOFU4uXByvmmKFCsyx7
ziBtEk+PzbNsqv5nC/w0MGWiPaC1UO7Z4gv+NfPE3bjgXD53gqlmmcJ63SOaBBbooymNhmrrMd+W
Lhfc0OSyKYExIOmrT2qgcNg5V+KEshAVrODP6GcTmaDvBXDqwWdQuLbl6nOxdZxni4VgAF7EItnA
ZkBolQnNzqy1n6pNTvhZ9DM7u+9hkeQ5g1cIh2fpKHBiDuOu7U9a109yPyY++liFrSNzRl/WKrQG
xrj0X9JNZm0U3/++fnLBZUcScpAb+5aC55WQSqk8OtFiKS4x0+uSKRHgnkH1vb21SyN8RmbDw9J/
cAcLMtH/6PoL7wTwCgxlk1UegjFRucITFmX+JbElQfBIeiVzcXJmmhLS2sEmAmFyirGcUr0ErL5f
0t8HY/BAddXjQJgp7eG1/g+SnsjbLMgHvMirclaysVWzNp5Dv/9BH0cZvJz85243lfIRevn/JlV7
NaEg7imYA4eMekVy1Gk6biKTzDeS/XZdA65ivd2zomBgYeNdN5uqcRMVU0k7YePf2dEvdZk2oN1m
TWBqNRg2cm7c1NGzp9io7gn6gMKvGoz45/3z+4Wm1szgZi/lJtST66LAhmiMYhoG2NUuTPAlUCnl
zUTna7w+XhvR+aKyx4XC4Ex28vFkFcrkz7p5WbCdd6GxwSrb9R5pBi7f9NC3iOTsSXMr38yfNmKA
0ISAy7qj0yMy5EXLAC0UwRSALPnFm4ZuCSbzcGpcq4h/NYpqvGSHBbSiBsuj8dfnhfAUi9vouNTL
c1w9fjSyRNKMZ/oAwkuZTkBxzw2gqgSH/HsjprV8tyVLXKT+lZjrunmeUvSYtShEudCdrtCKLzC2
JXJXJs64l/iwLGYTe3LcBFSOCQ6lwF0xd4ib0r8tOHD2npHkFwTsVW4FI6WM0ASCcnby00y7JE/1
9HkCkdklpxtBrLh04sEmqsK2U548Ab1OPGZiWyNGBGRDpb5cr5V504cG2cyZFoGs5AzlT+ykKlSt
M+qtq4Maxz0k/l7zHrzFF5MSQgHrHgdzH/HFWtJm+iq2i2U3+IUc4755rMWatBl0prGFSOe7ijLN
6M/5gHiNTDAbVBhbkOnRJiTjWWQb69Hi2ntEdowKS8SsDImlJNkvwh3rULdTUfogWMqsteYsLe7I
2Ydi63sdoCJviloSp7Qdf8GEaNTFsXOu5SSnRLazQIrelHs2dLWUV1AkaDT4sQWhR/I/ogGQXOR9
xdRyvj14vkbVRJJVT9ZaDoHtx2dtsBXxJ8wbf10K+F8LRYERVaASKqfib2oZsqHall2a9Pt4G9DH
fTzwltnneXmknn02vncWIuIfVoqoy2pGXhnh1h2aFFRT2ufR2wGiJCawC3LYvyo2o4VF3S0Y+AhL
jqaIe406abDFAUF21gg7ucoxi+Cmbx1mIurOJNdj3U0/W4NQY0gCY8hdDlf0XXqEpcb+T39YQymW
o2sXDtUwFYQv/eHm2jfB3acQnzKb3YgiRznIasq8EN3JZJFyeMrkQ4oenrBk9z6Agmg5TDft8E6H
7ohCmOBPTrW6SU4nbBr7KBBLsfhssxPJeRW04HlZdazcVjv+S8B5uIM7R1fG16Q8p2QiqXvniSmz
J9ETDNIDIaep/WhuUR7/+QqKUhHZPKWL6vAzOKe7js6KMizF0hKwk73KNOp96Vbh/hnw72bCdSVx
yMkqfOvOFp4VMtHkIo+c7bz6T+NxDkZwqyrIesenSdOtRkdt+wswno3HodwlAsXjbdrHNbJbiycp
51H1eY0sHlqndl15NhliTGjmmPQa39aTheYtyPLIWoYdCPA0b4snOjIGKCmlWKwJtxq0RfJdwwmb
dnLF9+WARy6DdlgYQbrVGaLLHc7CbKzY+zyI8wJqzt1JFqA6hTvmygpU7p62EZ69FboJ0EqJbhh1
4n+KYQ7NvhmNGJ8Jeh4gdNU1QXvDlr5WKtgGYXBW6YyyZdhvoMU7NjPa8b3LjEDnUTJSpSDLARqu
JzM4skaZz6Y0ma0PPLoWe5Y2TKEcRIQSRieS/JYGz6OGdwgAc9IjvOOyVw9CiqzojEJ6GsaZujia
u7LqrTLtOaU/MRyiNEwmDN/5v+vXcmAvxgLrCW5iLbPpNskKVjH7lOid0N6ZgFNPgvjS1Ov4oyf0
E4mcvWoQLdD8grnPOKNaYgDMunnWFakddN+I30t4fWjbQq4k2gJLxZ1h7w8JXPuZm5WbC4gqI1Xr
ZeqDwx7AkLGaGOuWibd/CTghEt9Le73+jrrVlqW+dZznXb38+9hfhBEzwZ4HKkw7OC+qw69vTQ5k
efOmKEGALnagebHogsuFHWOTe1cE2EBN/VnVXMUWHAj5lmsW69BYEWl36yzdW13Ujg91NbHXcFg2
jrbd2YLWVrULNLrzANxYnlRCftzSv3PBeBi2z5RcoiHkYrBFmwqyYLDt90eRGH8Wo5F4NFaG1inG
W82cFTfYSG6g7PuGbLB8MuyfdJ2RIGZMWu1PKcR0OlJRuMqI5V9vAyJ//OphH6SC2zLrIqDhwzr1
TInJgBRbbhkL3FyacVmOsAvr+srMnMuljVlZOtB+xFBbnoNfQS62BktMwV211nQrRSC2nfJDE8L+
SMu84EQbpbvPpH3dAOfKAGqC1xpdF7VJCx+/JeFjRzmV22QHGH2CsEe/AlwlAcYihggcJEoRc5EC
IgV/nEbPlVHEr6pnLDnCqoYzAC1J2NksSHy9OKLEzX9CZurUvZuugnzjIdlxIr7dAzqGC9faqisB
b7O6PEynutTBX8mzY6J9eumLM/Bi6Xo07CYUsbqI7GshfR5L5rqJdhIlq/YkGt4YtdTvZG4m6EAG
2rqdxgWXIIOIRaexc4TVZuN1oiFgc8VPeH00e88ngGiRn3pZRosrmlD+LH0dPOwWG3rvCwzmw49V
uMko/UVePWjZ2lhk1fR9uE4fbboX0pDK/HHK4x4bB3sksuvURv59X0oDf//sIsp6u4PDRnzDoNs6
fHz/2R2O1FioA2AhPICPVpz82wS/FzHyb43dEx7q+yVTyyFTbsAhJuTWFHYOPNb7n0lQfl4WR4+x
QRzGArWabGDLa9PY6w9wQBNHdDc/a/MbFpdj6f3OS5Q3d5ZfBhALSM3R8B4bkqxxxyUd/pVfh20v
cX+tY1P3qvB7wW6CSR5ihT8uBA1YARa2CzpITDNALVirN8R5Yp4OFsZ4lpD+ckm52Qy+FXJ3+t86
ZU5vwzKzr/SrLTzP5p8jRjsDkIENcjQVPPDuE5PMSZO2z03ojKehp9KcCTiBJWGE0zYDKNUIACO1
KZger1xiT5UhkAI9f7qk4i6f87W6tAy9CpyJwkBpr14T
`protect end_protected
