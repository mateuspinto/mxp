XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c�]9��~�WO�(�(����������@{axx��tαrO�֝ Q�ԧXO�Oow�:rO�wkq�Qq��ea����"���|��>R�@'X��D"CH���$�T�@L��w��L����
��x���!5���[˙�4��|�NZ�ANy*S\ĿE���#|�aa��ajQ0t,ć8M����h�G���x�r�l.��trƭs��sb�"H�F��vjv�;ژ;��L�q]�ML�{1a�%�>ٓ�(��&k�>FP�)�}�
ɝ��Ĩ��ݺ3�]+�l+��+$�vQ����d�����7�9�w8��t��)vi?y6���|�r�K���(,�=wa>�;��=Gξ-k��6I���D6̶4�'ǀ0�z�j�����v���ۋ��/�h�Ta[�ٔ�3?��*����qV�i��wng���t�"�s�B��ʶM�(�kߥӹP��E�5�=�ņđw<�?4j�PYD�	���H�0K�n`��sM�7T����?hcK���mbOS'����n�=)�n�k����i�<אx�Щo���I��_ˣv3^�F� ��!}����HUz�����i[�G��\ ��A���{L��Ԕ'���zj����Q� �{��kVC��>����cW���/�˕ft��m��
5h�:�
�����#;�D9�-$��#�	>O+��6��'��m	� �"`��i ��'m������qd�,�a�0����7�=a�to��	��{XlxVHYEB     400     1e0mXgt�����,�{��i�(�<X��c��yf�1�|�&�W�H}�Z	�H̘�Vk??�����X�kJ�R��h.G����4�i�l1�^̑������*�7}�<��$LRn�Sؠ6�HUz�r�.�
jt;L�`=�1<�jP,KJ%P�n��x�;��@3��S����S�]7��=��<�aRJ,�<�i��ٟ?�j���~�@ew�+r>���g߉�ilз&(t��������[�}�Q�:��������C9 �=G�312W�:�ٳ�eʗ[&��o�h�m'kͼ���E����_�|�P]0�oy�هP���y�2�uǴ������:����OZ�����"M�ƽƎ*�Y���ݧ"�+�4�!,0��)`�?&�Wp�߫���y!�Q�įB���ٻ0�A{����F�l�޼�����R�qd]�&6I�[q�F1 �~��%����p�M�B�� C�(|�Xs�uz��XlxVHYEB     400     160�;q;�+���?5$>�+�ɑ�?���"�����YW�t9�/�-Ð�;>�'!媮1�]�q���eT�S�x
+Ԣ�������o+t� ��Z�ӂ��[�S�ͩG� ~��T��O�7����KZ?h�{(��F����Q�:΢�wBG��/$�ԐY�����164Z���V�l�&��%	��dF�:,�nJy�
fQ��
n���_e><�Lڣ����-����p��Y��Qw�.�[��_�QJ�ӜK��qj[��.�<[��B6�d��g����"T\��sk�@ ۂ9��W����X�nY˻�8!�)���0}Qu@�|S�?G���y��)�Gx�UT7���XlxVHYEB      50      50D�;6�Ĝ�|9��E��mm�<2�6٧��3%�-�Y�ܐ�ԋ�vGS3��p�e�Q��m��J�@�`^;C����