XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ib��8������E��қ������������ ���?_s�E��4�4$�����%5�?��TLt�;kv���[o�T��Ĳp�22��E�ΑAh��/L9`��l�Td�n�c�.5���7D��Xmr+bs2?d<�s�{��Q��@͋�PS�| ��Zr><���#��g5q/N���^�nSenK;��ǄY���E����.�z�c{�����yvR��Z ,Դ3�#������!�!���Ի&f��u� N�l�Ֆt�f1Y���h����;�N-�H��y3��J���������ڭ�=���P��v=F���?�#����� *}2�F'^�V�KRdl��D�&��*�'(1I�8YC�D�<�+�>�⺙�[���2퀖�,�Fx��w	L��-�/�tj���4����j<�,d8ѽe"8�;��q)�$��P���(���(�#18>b��4�v����-�*`pr��/�A�&�VB�L���˫�F��Uz��U����y4�Q/i[96��&���Y"?�)�v<�9�5�����xS�|]�X�y�M���#�~�wf��|��цz�V}΄� �B�B���!�-h�p�]�1���흕��^�pS=��@�Yw�l��	�m���B���d5����Y���5!���S�~�i��ft�h���J���t���N�qp�������kz�ysb�3ש˅�X�Sb?�pm�!j��Fr�F����3/GQ�eO�ʠ�P�?�-{��I�h�XlxVHYEB     400     1c0�u�#J6��B�77r��e�a�cSy��5a%��.t�D���z&����;ޱ25��ų��3��,���wa��S?K�􎵏@u�V������뤃GK��Ǐ��ȏ�f����������e��ZJ�6U'��L�P*D�M:
:�����+;&�5l���:���$L���Ԯ7���9R��f��E������t0r� �N�l��WZ��B�	&�15Q�������Kw����oi����ھL�(82�'r���F�>�4z��b��Eg�8H��v�x2��TX��R��Vw(���'3bV#�z����{���W^�/PMR�(����漢~�n%"�Ml	�~D��e��ӊ	VG����v���|%�:]o ����	�!<�H��`85G�^/Nը@���H�yV��/3Y�PNt&�^פ>��6G>eT�XlxVHYEB     400     160E����f��OS�_"9f)���vy�+|њM�`���?��6��C4QN|�����\���^��c������kh����Q�.�B�tC��}��u��=}��?v�5F�#<��o8�������M�]�o�!"O-w�u;�v�^AO
��v��}���.(�	����O����Pt�k��	��߿��O�U��ޗ;�������F�2�q�a��l�9Y����+PE.���V��@�� ��=��e�(+��C��|s�o��l��.-�4�����^��~�;���(��,��Z	2[<]�є@Ѕ��
/��
�ّ�\Ip�*�,$��:�@��pN.jg�l�.IXlxVHYEB     400     160����T�s"����9���#�j��t�Cl�F��9o����S�����]"���^�9g�L@20���#���M��k��ol��q�F"`�"�:�`��^�L�W)��,�H��Z% ��P��>}�<��$� �Ֆ�p�|���1�H)�C�%ܑ��\M�D��?{����<;%$��z�8�'u.�'��nP�U�F�ػ���!2���oF�$&�0x��F@�/)�U]O0�z���������[.���0Z���]�ٲt/i��"�\���"M�hPr��)X�7쀺�G8�Lⷅ��~�俘H*ِ���g�K_���k�e��G2��a�WұcB3�D�	��_��2XlxVHYEB     400     1006�C�Z�ܝ�g��'u�b��l*���u;�y�����'Ɯө��~�m�B!֢Q&5�7����U�.����qj.�M9H�+X�Q���\�b]��(���yo<]�C֏�R�tg0��ZCӴ�$�wx��d��|waVQ;d�{�T�g
��y�!�`#NLv�<4�Ic��N@ַ���`��>qD�q/�wYS�'���ɫ�����$�%)~Y�;��Io���B��'���{'�]XlxVHYEB     400     1a0N���G%6��E.y��z>�����Q��K4]&�0��h�c���1������?��#�������#�\�xb�8�C�� D�/&�f~���5ؖa<	��I��O>��w
קˡ����a	2�'� �5�����\S�t�HƆ`�-�霔����1�x���w>w-�(I�E�챺�����"���3�q �c��e\���<�p�v_�`��}�����}�HhBaP�U�U�V�0�7k\��!�����e�Rh]���d;s��І��������w�P��\�����|1=�k(�����Q^��"�%�6��`�vK�a���Y������јgc�3O��7����C��l:���j���`rw�A��x�����+d���z��n�oÕ?$pphI�¬di����)�mXlxVHYEB     400     140���~>����d؟}����n*޹�������%鬓튘Ԛ&7���7���X������j���q^+�n�fa��B�

�~�L(|i�T_��]����+Hi.<xl�ə.d�k��B
(�cP� ��'����g�9��D�.P9�a7ZE���5i�Пm��v�.
9�I~+��v�ݹ�������螧%�o�V;FS��������أ�?Drp=�*=a������C@&�)�������1d�����*[�V�W�S��)���({��=G#�n�w㔤�fszj�,h��d���k�u�����XlxVHYEB     400     120]/Yg�w��-�o����`*��,`"n������1�����%#}:���7�^��%.k�G/�
�)�,���D�#�E��ɋ�ee!�����U���R���ӆ���4�$8�wm�f�,�P+ϭxjȤ����+m.��O��Tl"�0�R � V�x���Lx��E{Ș5d�����p�L�������4�j����� ����Q�����]�����ʻ���<iw���ذ��H�?�=��I�3c �8�������`��݀�t��Y}���xg����XlxVHYEB     400     130�$����c
�Q���±c<�}�<�c2}7ʢ�w
��S�����SA�!�p�ȴ�Z�)Ό�t�|*Z��UGQb��2�a��jb˄n{=wh#��	BFr㯬uu��37��+5�6H�3�ʐ%��ȍ������X��a�|���}�P+����m����~�4I�|5���������=H�	��OR�,r��=��
vrq ��y2�<O��hꀍ92���e1�4̜ (�� h��~���syY���ڿ�A�K��`�>���Ii�tH�}��Ev�m�Ev
n\
�W�r;~U�XlxVHYEB     400     1c0,��qu���Y��pu9�V5�|!]���F�ې�0���U��t����1;?�Ż%r,KAH��£Z֘������(���N
���R\k��c��mg�9��c&���S�2�ӊv��ڋc%؜<����P%�UKl���I��Ch8w|��^2��h�k�9s�d��b�VtX���p�;�I����l̚}N��X�q�S���E��� �W��Z1?�?������@f	���0Pwę�)��3	��˄jZ�+�vrCu��!4��Y\lxE��k�2����tUJ��5�o�-/�E�-���*����(���s�]��קO?�uHZfZo{��V�Y��R(���0��k�D_"0T���jvsĽ}� M�4piiӸq�aU�Q�������P:X��5��1��R�_�}\[��0M�?%"��� ���-���tXlxVHYEB     400     1a0�NI�r��DP��`Z�|hlM�ZL[�5��+*+��*�����[���Û��TD��N]�L��V�m���{^#e�u=S����9���AVk��I��(3I�)�iC䉦�C1�U+S��w������V7���CNp����d�� 7މ�F?b\���%���CN�M��8�R�R���0d.����������R�����Y�{5nhF��:(lx�0wQc$ܐ|͒7����U�!����	�)\�S���@�p�SN\�u��	�?2���j�"�ء����"*i�M5S���Lg�2���D���}4�)o6c�eǀ����q<�;��6�62�Q8�%Vq#-�0��|A��4�|�uQ��v��蘿�M���P\+FÄ�u0~�e�"�x�l���X5�?��XlxVHYEB     400     1a0|�Y8��Zg�e>���)4!Ƨ�T�����r��K��0A_�.F�l��?*a�4&tɓ�v,�@��C?��s"N�F��ݼ��5�Zȣt����Z�"�@�|���m<^�x6�2&�]j�`Zt;@����>3-I�+i���sR"?ەz��_2�1��{Ë�1{'��#&n�w8�烉(ψ��-ɻO����ug������3����,���Ap��Xn�}ް���,��}����3� �d�9 �{��/9[?����k��:�N�XPg�ncn�ᑩ6{Y&����=Z�u��0���{��Al�md��g�l�l��s'-���;�T��c_
hX>qA��ЪN�\����i%��T�i�n�W͇g��2n��&��bN)�p���p��� ���Y�����K<MXlxVHYEB     2d9      e0��m�*۱S�/��W*`��|�,{�6d-���_�]nS:j��r�v�L�E��.}v5��Ly�I\2����R޸��X��-`��nƍH����3v���|x���3� UT��<��=�kqG�U�������2�v&�S�;]g�HX�ZX�?��+ c,0\��h��7�5㖯�i���ΆW�p�@W�A�S�5Hc���(����_�"�6�Skb�8�Yԅl�>�8