`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
cGldVO/G4klFWHnV5a6XSx2sZjiTWGQUaLHltGO4wj7tCSOvuH7JL/cayLHTNDTQFczqFjOY6tST
gaxX0SwlTVIfWMqngR/X4TjD6AZkG4xMoVK4tRB/9GsjuCYy2hEgpaCM3UhrrjFjk+WNa/crG18x
Ej5OyYGlIdovUKv4J6lMhDE+17jFlcysauMhYwWzperoqLE54cG7YFN+Dp19ER5e6MqeTRE0FUj+
1vHCywvaOq/8cIP5rKMmJB2PBHeMqMYapPIxAscgEJWu9KhJRmYoDUfEBNnQX1bwjE8nE82qv5lq
xFFGSoeYFNaOHaYziiM0Guz4Ye5MRIF25O+53A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="H/Jyjca7iGzASkkM7Ici6wnXqN7Dgf6MMmQGeyqCqDs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11648)
`protect data_block
j1F785Le6X1LKkYLuBLPuDjLK7dToo9M6QvBsNAMSpPBkEXp0tHGQb4bcfw4l+/bge3jauQi9PI3
rSQtljgiGiEm4UMyZw88lkavY8pgyzPnN5NbFBuJQMRJKfCgMOg7jugjipSJxf4D2hqTxt2ZwAxF
hOGVT6j3q0yzivi7SjoYkReNuxYfH1aT/TdLoP4hKLfQcnwFn8XF/Z9OqjFT2LdYkcJ0vRdls6//
XqRETvIHcgJDiaaPHkgd4QyfP3Y1LMDxUtidiqnEwBGj92MBjgW6UkkkBYut9mPfoXE6FTlB8ujp
GMwA+At6N+FFpdW87fKQ+ACLlBZW4rKpOu6RQJSdfCc7OE5F/NWT9h5AKKWEjcYV4wICQZcOJhwg
jp9bsXwiAzJfukALlCtIbrZLfRX9dD6oXubyLAWhvqPFKHrpnSoutzNquE3ExamieRkkG8VD03So
bKFSZZ2+AiwdTOKr3gHh+ff2SqZ/0vHaEnMJB3u2MypdzmppBJAWjUNIfN5VxcRfphel5XXMj3xu
CIz/2Uu2tF9S2OtoVhFvqJfn/+EArzuD0s9W09L5VmNQ26XIn2NoGh/maDjId4OwXoGKEWyIORoa
4EPmUlXPO+C+4XCRkiQkcNNiHbQqpFcEYnBVzxZxQzVIkA1XaWpl8lVlWBnMen6jQLlG3jVc1JXr
0+RYYRT4GyZr/ySG5hazbun492hViN6/bwbCzayhGCSEBBaOeUJzQ5xufSPR6bn4KruzCXbZJ2Tj
7erEPIsuevRbq59L4fi8cHWrlMyFlst72NfFW4yj+hgxKxJlwxQi2P0VPOayMfgZA8qka6nDd+L7
7kd66sNrTvUDdvgF880aiGji8dUiEUiLyAdbUSiU69IaSkRa77NI5/hglm5sX9zpBH3Lv4gniTEu
oFA20GgMxKOPBKug0FZSp9mj7UoOdoOh0FPGZ78fJ7i55MhcWsbMFymyNok8pPhxjU7sxzq68V57
E2izMEG/e2JDb5Bb/usnxREEMUtYrHbbrZTDNUSp2twG6dxqHUwHrYgcez2rvkT8jtvwONTZLF2Z
5uLb/5Xx0WSSqfIAo5KgCiSggLjLRqxHKxdwrpk+3rjIab4M/Dd7ko5XjIpvZyRhwkw8Pttua+yq
HTRxU6xuq9NgeF2gSDyor45x+uwWQ7dxUdvwzkGDmoOHmvTuvWPL/wzqyyV1e3OzatRhOpZNzXdw
0zpLuHhUfzy8F9o8tZ2hSuwEhvHihTNHpiV23bHAIfW1PtsuIhZK44OP4LRPHtCVJM3ZZmdGOWCJ
mOlBKUmEApbaF7QE7LTHQoFZKFBxp3MugaUcA+NJC5l46WEUnCC1LzGNA4h9nOLqepfpEeMZ4ncL
A19PwYZyaKK1EQBElZYH55IsCdj4BjXvU7AxxbK2PhextFfNgCve3jTun3XPv8R5gvkyoRwSMcy9
EOV99LbgLDq48etSjpebxUDZ+wFGIkrCJtbqRn/2CBK8JhjRxi9Xh6w/QD2/unBk2vKa/JXh3w3d
yOLF+C1OXR9wYr25zMk+JIKLVV0k9Bm2D+VrRpuJ6av68WXbaahAOq+VwVXhCBvHKdX1FXlnSnPE
ijNXlAlfOzRSpm83I2y6R4HUe5Sd5Ctfj1b1hxBiVzD9CvIZI6tSWW/5gG0LoXTKR1uBm8eUHgEe
DjwB8q7mTaYfk6eXzvHwNiFW1qOKarZMnNIZ3WkRmPPFN9JyeeqG63tEporOWng921N43+R92ioJ
jt1dOhOkUa4GyhGIaazumKJblOldS4uIr8QtLujcLsJXPo8zf2JPMd8gvHDttpauyBCAbSY9T2kV
MPan0VJB++T5DlkZVRGLg4nFL0p0hDNkYim46lFVj7ytF0Tsf4oO2QUiJmrFbdiGRtqv9EjYc1If
NKgI+lJWrEl8Stthq5fLtmJI6oOzpAtFUTDlq77+/CvLaA1WeLzoPN3ydarME8VkawGCD8mF/jo0
92cagElW9fkP+h4SiyAZlA9UuOE4z00xHJjt2zHbF5NgxoUUIvpNQB9B8nA+3CyNYsatrvoegCDi
6nCiTxZpwjXL1Q43bEC9CagJdJYoh+ohJxV8FY7zeD9zklxvwLi8v5Tfjt40WFk2CLGKrX/PK4pN
Nr5vdSu6OY28ciF2krkPZUyb8VyK3DI8T0/O6ciKiJTyGWVWSut8ZC4x8p2BiCCr83X+nKu/hE2i
t96UFI1+fv1U6k53Odl03cKfYEdXMEQ2NbeYpi8XD016Y/U5WkPHCB67JEASKWjpK05+FYY+jPBB
no5aGKCPX/ytlnQYy1Sr6SkCB6XTMZZgiOorj7f26VpMXGONDYHtVwv4dsqGHus12J5TslKT4r6l
FW6GjELWHpsMb73doJVUbxdXxWXibCRyDkUh53kZ+oXO1wJ5ByLZNX1EM+LRMEht7sPdW5DfWYI1
EvL/vKPQTHuU8vInvgmbPvLNVdqo/DVjQaZ0hxMGElz11MoQoBMKqoVLkrOsXfvKyX+M1qX5rJh2
gsaPi7ZXXU9YXgtneaZLdZw2DmwU4SiHfvt4QHRypt6LdemFAL4YrBA3R3IqT95DEvh9m9xbY5pR
7hP/eWXFGIC1PqvMmhFMGUNaaszh8oLwIp8HJZevLh7PQiAeGpVeVUXipEaX7ABHd7eqWbEfj5fo
oiXbZvVpRw0x8FkdkslwPSyfPdxZvsQJnbGAldKPtKxcxykOy2YchBrRpmQlcADpbNihk6cKm9BC
697gjI0B9wY5Xg0XL6xQb1aCenzQ7VeyjxQZa79dQd6TmRqMVvA48nFKZbN8WghR6IukkB6L7OjH
pnohsQciE28pzrF2bvwDQG5pfFxNVbtpBQHtcQhRZWmbj+xAgkzDM7FE1hkAJBvpkS6Jb07FboNk
pj0lRjr9tbSo+scEgJYVLAiY1etRJpnD6rVY1nQZr3GINqA/wnsB1+eoZZdGyBI4wo719o7YAZ/2
NSVUFh7Hdv09UqtKo6clhSptUuB9mR7rKqRMuxtGKJrN1DqlVtqeO9cegzZPYABaDClVy8shir46
TuhWFJQ+S72z4ie+SEVx/aN+YzDNK9VyzrY8bl1jY5pDmOGY/Px26y5TzeXxm0MtZGnLxIlbxBpw
KQ/TprLzitOSeg/c2YIi1vXGKRzP4ESaQzZt304vMt5FB2/0famIrLEOGEspmoGIT5e8rwVgTzAy
MEyRDtPEDozRfHGkczoYxuOusaibDWR2X4/m/+aMzb7+FdEv5adUAPEBKEumWOjk0EnUrPlXmqLd
kVuEvmPdSTn2R2dG+sO2iVMi2dGGLN9pV8QGtUS/FkzZF0L27j59yxlc6NQLWRWIr5rR0Cr0Vc/0
H0oyhlAImcPX6cG9phJEbubum74nyw3Y26k54YP68X+tDNkN4RUh8JuvMZGOwIS25Hg8Qt/RgEpX
3CmNcn33k/jKebRkf/7hWDUawXkY0gF6bCOe29OhMe5v0+AUmW+rUS0PDqmG3WM9On3FhnGy7sAR
G1xnftmn2n58JGN7n9XwPqPqFs44TYmiNBEjv57nD9J5m3Q7NUqB9q0kgaUu+YOfsN9SbUX7ARIq
S3CVbZatmVPtkTddsMic/MBGqkUY5H3IxCjq3OkPRpL81lDYGujCWXqtp0IVlVwkZCBpOahZfY6F
ccmin5jovILM/kQRdy0Wvegqij0VRuG+6wEp5ok2kjOsw8MGWzJVFG7rmiLQJdcr7TZ8dEu9FtUN
V4k+e66PWg3gfHKWr6kIxobC5zML72JkD0DQCZ2QU7hG0UtudGHwfbcpcqvjiiYoXKo+a8HijbL9
35Xc2mCn3zHDG7k4rRXrn8wEBsP5HkFV7Uy4rM1I4ifJT0lmWRjX77iS4514bbuwd7/A1a/Um3OF
Ojqv4hJmH/eg1M6Xkd+f5Pd7kCKuSwSRCMbMqJXajH+CESVbv6Tf/3+3mq3W+JxFrC5N2e127ziA
Z13iU5Lk25C5pbvFUjRk0lcQu78rPNXwqMTkLzmFSzURVfI4WOmznUuIxCmngRrDPeDHom5VE6ed
K2oKY7UnKY/FFRAoWG8/SDo6HkJXnIGQxoBxpRE+1KKdDhpcyQqnqT97CL1Hz89IM6lbUZArHrmX
Vu3tediHwoeFicnZHzWnmYpaTqZivrXzvOU1xkN0KNUZslTLxmTCHgEoqCzT3Al/HTBLhZipWemu
j8lyZc/a6T3rdD1hLR84L4gWzgu3AjOS63m1hCHjVp3LbUMCA8gl1HSQrBth8c8vDuDV4vZ5fVoO
y26OoFSrbNKSAJGByTHJ1CTzcfKzNuNshXkdWfkNByylB5BOUWPLHBjEwlp4s3Y31iKbPRFhEq4c
160J2l7G0T6IBOINosPTeoVDvhPhJqg54gkFaKkd9mv4QZHTj4W4bcuZHNMNu48dHMSmU/JsQiRr
ddrxgTqdM/63E/RhrC6QnQ4EQI5BRmETEW35pwsY5vthDgx1C5pLyLPOnIU1viiiLzqdixjkXs7o
zY8nYoIwhHdkjpS1HLVOX9CvjcD7iNCOfbN+dghG1Rikd3A7JrCHR1vGhkExCBOYhIeIG9puU7Re
fhrUyWyt24tyahPJtlmvQP7vHYMewmSgh2I79LWMAjcsohlIOsj0nxJO3ESvfFs03Q4Y0g5lVJWc
NWS2hkP47RRnMelBf1qr9WoNCQ+H4+7fKlRfqAl6dWUFssBXpMclwDMMJJjqAvRRmkMll/IOTcc9
ezAznX0d6put1HvP428oAM4mCOuR1mBd/CFkC0gK+BPrZC3LxPG3XQD21zS7bv/4JA9DAsR8uRLP
DEGOuO8noAF34kEskE1mBsBXiTmHbkPy+iSjGHleOVFtzHi1LzpbtH5xzRRX1SSA/xzAa+gajf05
dnlhkLTGBg1geq3Y1T+xKAhQAjD3J5IX6afhHW0AQGzLDgv+0i0yBka3rnLR7V61Gxo55XoTSBEh
brP/eD+LvEXlySmkTte/ok0+RTRT6J03yKEgGs/smrbQoNOjTOJ1IVcXfpu1WipepShd/gl4lhr2
zUgF89T3YEI9y8i23NiHdD3/URzSE1k21rNr8GBdwUBekmsWoKC10dVOV5de8JE6vbjLlzQI8PsH
FdBgcBf4NRvWHbt+1kKsPrdIyzVOVhfQVddOg6igQeqBOlnwrHleeFsZ3uJcOrgf+QLIFaQKA5Sr
oq4Wrj2ZuwWwu95kG6Dtt+4lOXaTsORrux07shAkmCz6OqcfUWhKad7Ym2GYW1X+aHKTj/JGB/er
iJpQqfWdMVs75FraufI1XCkqrLr+2VVd9/tdnfA3d2N+ttp9me15m5gJoJQ7YSoXW+9ZxIVVzG4F
0X4c4/AesXTHRSJfdnKuBfh54EMpZNgV0puotUPOSnvzbIyMQNVhoEBfmaRUNZe0dn3qQHt0L26S
lkuEOuUgzynb6Vc2Hw7S1w88HNcoEdKiBLGi0lfC5WTBvwyOihvZaaYmgplYhxAbLjUw5SJSyqgU
9O/NoC01ZZsb7SBBGIldvgddVjgzmmY6SicP79tiqR1UBdf1uD2F9pwVQg9Z0EJvYaU1tV2cWD8x
fNhT4op5fHUgV+gJtKxJvYGsHo+AoftIUSFl5LUfK+OmKrZPPePtxyZln7LpPXk0aYqQLmyLx5yu
xAMUJdAPWMlVDM8nl5PUWwwwLsFACQMWr6+VXy+v9KA5NDwcIBqhf9UMBnYY6mAyghuCV2ss6+uL
Fbe9zY3vFU+07sSntXKEWMNgvQo1SByR2TyEOmUaAzJDrskJFpyPp7lhuJwNqQVeiQ1VJKhHt5wM
VYnwEV6Og4T0CNicsX5EJ0SDUDfjP+YQ7u5/hRMiS5wp0srglH1/6FG60ah6Pd4VjY8IeEgrgBLR
liF8eXh0+x1DmcJrvHtlUIhT3hyRAO9LrTb+fwo/Pj0vOR9cuAvDrcE+wVRBHtycEinSsBx4Z133
PNOnlUzb/kiH7UgSczZ+8gowyPczGLIB+BltbDYWYd8mhYuLcLQqObnrKhhzTSkolnv28kBq9ECc
L7Ip/YYnnZcqTXdRfpcefOXRyZnb/2A0B/1Y7S7dxbLfUiI+l/u/pAaLUo+CoMeVAd2SvpxN6gZp
7mBYI6fFKYkz94LyWZKCT7Djfh2mh8SFq6o05dP96s7w+A0lGfpnUVZ6sOMV5XV8A0s/4pfjk3v+
3wcHEbgntDyMHQLC31HN8zVvyL8giDg/pk2ivtf2YkKoehtCuyHxIamayOGJ/xAVH7qPrBNVbIhD
Y3kpxJG2HQldlNF1B3v44PgoLlzS2+/pRQHonNW5KH+RwXR2Pu7GBj487gzPInWzfXeZhMjsPIpm
nmz4uA+8K52H8HcHYvuBCCdNSOhMwXifIXLLaWd1DjlCzrzLqCQA9xPniMOQcS2Kz1DQ9l1J8j6L
kHuraiimPE0hevX+S5W9oi2eLnrMwhnrAGUmascGTXlFoZrg6uMhXWbAPXiEX0eUvk+tgcA0sulE
TMHNkqtAX0BROMO+ZsqH+DDh27rZI7akMVTa/qj8aQcOoKiweoGyoC5HxtKXxrmpooBUyC1yl3vq
XDmHLvF/UQ/solE35Wj5C0WkwRYBkPDktz26fCIbjhxY8eM7XzTyUllk/BzRZgQGOQhxbwHIOD6Q
cyOOeKGjpxhOKwVl2Sodc6Bmxn8NI124aZX/X9Ns1g4zx4RKMzT2/1kP/AI8qxARfr9YntNFki/e
+1CH+qOdsNt937gD5d5zOVb2cdVGKm25tfWBccve71jA5QwZCJvbEHHygJs2FWSTzSY44wQ40wLW
aqB3iBDmTPkjwqrzX8vcSXLU8XLfJT4HjX9ZC2NE7vPvjA/HoCf5SHk9Dj0pEOkCjz7MvQmhhC8m
amDnFyhYRvm1zdH5G2FUNqHvQQ01Nw8G/aASrHtsE4ajGXluIw64H+QvSY2HdemPvz1oBC6HW1Dv
zdPY1/W3VrFkkkobdxp8HYaoKFU0x/R85FPYicNeQ70//cls0LeBjwApZ7iGsfK2AN9m+HdBRGFz
TIBmAGef5WFXYqAVqL5kOE1nldo5WlnjjjjyCzv9B10zr5sPtOPOSwkztxB9J3h/MvSw5vfM/RWL
BCywNuKZBC+g+Sd3IEGImgTG8d+uxQlaFXvWXfq2tn3HQqBNwTzk/6J/JN18jv5dmAGVE/HY5fvT
wflknr2GpIySFnVUPhdlPwfyF9k8SdNEugQC9AoPOwroq/aluZAecJkgIqaUYWKQSeFLeL1jYWck
ZruCHOQ6y5TsjgPOvJSvzD+rR6n0WNy536x3h2QPtiEbUL7Ehtz15VhyKIAjjivBtXwUEUfDN7MJ
FwEY6dPa3qrpQxzIciNrPtMPNPh4cv8fu/Fgm09yGuZ+fuwGfw9UGw5MqyrNPDK2hBsdbnrqMh+q
qSq23agJjuFBnTPikt21rYKo6TnYjntHstWM4ChafCCHL6fYTmtw6oQNXKMCnDuzU1rG8b9ZLZnT
JjVNp7sxtZiHLB6C+rlzsIchev4/7TxL1zr9xqpHUGcAqGi4Ef7lBJRobT1WsnxPR/9kGIDNbUgy
yWWGwaWKpviOg3YKEq9xUjQQk3b2tI5WpKxj07M1J47RJxdUV70X1I51PaVJ40sEtbONuHETNR/i
6v5gLJAmA/4L9x+m71mnSv/48APxCnlhjfGJpw4Cvan2Kl0Niep+iYXKeQF+72tJoco9nxInESsP
a0nSdrHW6inodexmsYOLr4puNZK+Ke8T8+ZXoIGfu0kYUbG3YDg/vxMJqAHW4UTcvZdxADjg9s9T
jXKa+cxjBx6A5dhFp8LJTpOG8KzfAz74QWiwQ5+7OZPmoppV4G9TOcD80SdRHfCJa+XI4+jqrXqj
HJQ2qnxts7sbmP3YkAYmM4/zEJsjxJ/cxHNoWhWSAVZovArtmK9feODcaAwKSL2UypZS5GiP1WpL
P2vtk8WDDSBqvDHdl6DiMNkHY/v2U+fpD8lqvkKVoQxt1t+pzoHhbLthuobIGtg7Gsk2lU3IjCJO
CAzWZvSiDVRY2W6U0hJ6AzofW5ADRMs28RdupnO9cWB6xlkzHpUZiYnsvviqKzbv/cYBicvIjDjZ
AQfLuKMWR9TN4VhXMtWJI4bMfLmrz+d2njNwKpmGcHTwKH029B+L+iGJ3QKSOz5SZnjQ+lOETnwF
3osKMuU5kRgei35zBswab0AIERhu0j9mxzR2JAdclvimncO9P8oDlXTUFIy9kFAZmKbAq0Vsi/QL
agpUnYkZWmaGBAr+FBQq1R1NzVVwCLwOK9yRrW8GwsKGyJmLRyLMmaD2QcpeFtT2xmIRiGXHBtOD
UtfjCz7e2L3a9wJFKDraehkl4nGYucH6Bz1buth6l7PIoCMwwJaD3zdKL/wBrzSohSDdo4hA/BdZ
e09OCli+qtfEAT408zSVOtafA8r+6NgYiy/e/qhplGyItE2F339iV8Z0wVuWcHL7o2nHBQ5+S0yu
sICN53aneWAI5CId9hb9UZ/foDo1usDswQ9p1Ri6WTqyL2RQaD72z/BmYw2SJGx7Qs/xoiWnpGO3
Jdt5jq/WHZi5SU+PONJvje/JfB3bJfG9vTjocipiKxH0KqHh0VxSeuc4kWYkaW/wLFx7T5eWLNcz
egTsP/sM1oH3HcOmmLNtSkJFfJg+QdN+IidgzfMBsYOn3r5ysnJYK3SBagOOqYrRIvybXJe6Tc8q
JzsTvGR9XDnPkWk1dq+B8Pg1eBTSGL9a938/fXmihW12hBGFZ61uGA6xMJAU7si17tsMDy4gBTad
XnQ2nOuo+JJPShtfcIptmWwYlIFP8TwfnafIHi9lsUF9g4ZPGkygQc4Vtr6COMNvSOt8SYDqGLPP
m257OOYP0n+yHIrpzhifU6BU2899xY8OwQ/u3TvDwm+g2Zni48/boQ++bYhWirqfJOvonQwKGz2f
6tWgRMRwS3rP8je3fVSXhYnZ8GmwKXZrjvZ69zA7rPyXZhWDVDHiv6iAFN4OqfbOJY7Yn2dpu2Fx
wLroSrg1RfmVKLpMkhzXD4APW2Yxflg4P+u1eUItyrEgkzjSjj+C3KvXHA+KWkUjN+HJ7zYBxMk+
5HMVGEli1C+x+gTAb5RJKaWDrXw0Dz0lBEa+K+fIuLWZv5CPFoTQtpV088+JtRGVSCP+UPyKLEeL
Z9aa+Mjg3lOrXkrXdw3se42G8mdXKeT/3cZg2Cy9Ey7JvwP4BqqshmDaNTKqlXz3c3Aq95X89Lu2
MgaySadzfb9OBNQgZ0SdLhaWWZdsKvWqdXjytH08xulW7zB22Ap8PdYRC73RERQd2UAAT3XHqT1W
9sTFA4T8nMSHvp3VKSaauTv9nAL6wRoHuA4DVkrANS00nlsiREgGV/QlpG+f0I+AS/cPpZwVrBJg
nvXtBN9tYjpPOJB3tPkcWtW363k4szMV6/9jdPvP6m9RdzxBHE1Gb7GpWKW/dI4ezVL6ZEZ0UfZo
AgfYS+RtjjJHHQi1YH50D43qf+cKWJ3cJ/cRWQ8ux5jMYx6CeO7PKvKUebDe+Cos7B3Jg2O7mudk
ZGdBYoT3jJ/NaGtNEz3rnXs2RWm55yoaDP9e29gRTx5hgz9nGinORgApBit/Ooho8fpsU+dCQ6+U
Cb1obJHODtEOrpBzqOu7gVq52kDKZ5fjtQvIiAGE2DusdFVgtegFKQC5VOy72fS7n4JnDmw2N0XE
sIUrqLuAADmjrioOZvBGohwwWoQmYcFApkWEliPigdu9MUb9QjWxgE6W/tvJ6CzwZoV4WXIxibH+
I3C2H4Ty+YuRcrj+dpGI4JJTMAK2UArhrQc9IUNDS4mo8+68RJKuuPb7OWxsnw1v8GcLq7zBbwNQ
XTkEXEgksUVEHaRtXcKZV1P8YGF8e2qgBnIolWws0mJDml8s17rLurrjBRiRjnkF+HJ3cOqGmALM
QXthpiJyj53vw0pqoCcPl/62ou5KJWAVLrVham/XlI0iSOX/SIc9PAn/k/+egZL6D2BEOWMxXEVK
LCTVFeAqUYPZCicTEHWhVTCD95RoD1/IWRwK0AEO5LuyAlEjVgh4FF/rmHVPCI1DdHs4lt419N0p
eEVv0kZdYurMY4jh0sbwnmztmK5ujx1AI0WK7v5u6KwtvnJ0sUfG7Uoee8URQylT5TO2nTY6mxgX
ztmjzI4hTLPHWUUfgZh9eLoFxydUBwotZHMnvih/k4YU1aPjZrOzXA1oGRAJbqyLtrHVEUwI5t58
kKzKKvTKIrt24C+KenEQk8VXqG8tzwTUNW7XCapBk9K4GcpQuTaw+fjZclytpeKhQXApYXz7hclW
Dz89gn9EkDD9UFzta3gxaZ+ZLua/sxlyT0ReVuKM8O2zsqJQdBH6C695lrqdib9cguxbu3SnN5WY
CuSHASBMzzKU+eRv/0IhtxqofKPV08Jwd7VM/JjbQwhelDp31gs8smmJcuUSOYSrIcn038f+xV/0
2ImiS1HlW05i88bfk9iVBkj4CC+wRN9w/aEkol/L6z1GfW00D9dFS28YsznYxotpcfiMEU5b4y/9
yRlJ9QQ+Yd3t3gP6RPMUEzp2AdcXXPx+r2OPHwjt5iqSgFOeCYX/rnFmMQHCtwlk1YNmKnSG1uXR
JxYsXGATK+4JmG3sssgjE90iuerO719wEl44hVRCa8REfQhRn2CwjxeAQgDW63+bSelfq3QFmkuz
YfTDDT7P35V6YMuW7N8++/D3rbjJ1LZg9FnE0npWKxsTqjtnIpCYqqbV24S6facII1kG1Xd2MvAh
Uw1Tibwc+QdJyC6WMtkxDN5EEakhlnKpOBrw0CP+ge/QO+GEgNHnIPCe2gLLexm5XbfS3hEGS63v
Mi+eZLydWJMOX0JprgQTX/WQvcOGfVAnlPzqUNq8fhHSq4wBfVtXr/TdvrTKobg7F8nhzuoo0El3
MFppVPoSrt2q1iL+kIwykcCTlfIC9UOFOWNUH8rjrVl0OGwkbeOriMVc3qFj64cGq4iy33vEMkZC
xjuOJPDVp2m2NW9BPumn0kDB4HZYgjqUIz3+hQmmNA5aqXAQXCEbm3SnDEkUrxtlFiwzGyFtlh0U
LKW1hREcLOHYSl7wkU3g2cIsfwXW2et8e4T7bANkbdKCotlvTe2AbOpJ2kP2xESVv3t0Jv+jeX4A
9OA58nXuMAdeBn9nbF4pJ1XtbECL3R2A8u520Zg1HmSi3gpzwCicuzYdYEXKSrv8eP15/kpSG9jH
obXH4cMbvB3C2156FlyTlJoiuMepzGbvdkwWnIjrZAHVsUVdxxTSLZdorfGrCv02fErU0oEWic2d
xGET+GImAUpb9Q0C0kD/Ji2D4lr+obsFSyOQJIwgQo0f+apiaGfmR18wxe+EKyS6Dey+4uIsHoO5
0xrg67oHqvpljI0u35dGetZK2p9KM7f1tcztJTH8+0+Mf+SfbrYwqtsYL1Q2IhFbvJdURUbgCnqx
zSAO/MROZa/zBo/WnaffxAg7KJzjAI/lViaTq5Ky0Ii5nLujWVijyMXcWUK5wZcBKepZ5iD8izUd
4sn2+2mtc9aKhSe+tJJOiMyMf1PNOWs1HCPN3SjAooeyMML5qP7wv+F1l3Rqzc/LmEt8J/nzoirD
55vclEDnVTI1aLN7+Ohgji80p0ZjQb4dK1R0V86vF3Nsmn/5Gdt7QAkfLrRYenvGCmIoGQI8oIdh
C0ZvBbm7BL+wKyUZ/gKtDMNkS1CwgMM1jrTJ3cD8ot+chXemDE2d/Gy2hUAeP46SD0P0GdM5Z/KV
CmpsQZ8FxZl9owhkW8bZzsrMBuUsyQW0eCPAaBPWDYfD0mtKk9UWly6vD2jPEL4STxeDyDD9nald
KflJpPtxFpHTlKZR4MkOxbGvCPP+8R6fa5PtI0sRhzYFV4Via4bmsxV08uT75k+5PElkGVAwk525
jBiI/LLHXIi6g1aWUgWK1jsQspaTdgs+9N1CyOoqfXO7Lbw/foCBsbSSxkYkjtdZDI0phcR2ekUb
ZlzqJXXot3W62kEFPjerCnjPA6iQHyEsR422wWVSe/DFaZkEsXXMYxacxm6gzKCZUz0gGubUWGxK
2+jdnq5rhP2Jr4fSJ9NPeXguPMnBNQ13cs/1X1D75OlwL0IiodTZ+A9C2qghl3wYLQvdkYnb0Z9d
yy1V2V+hRhTpdgrJCF3neDRjyAcE9aerz4Ven2C9bV7U61kCCmoR5H1A6C86reL4TtJ/5N/y3AHb
pBKrQ/OBEV0tQXVczZ4jGoYKq+Tm3E21k0cZFTcen4SQS1OL+s/yNLEm5Yh/CHAgkCqTC4I4xCn2
cFzH34ux1A8xdQcM2hcCzXUkqtXyzqiLjQ37gdDWY3x5gQGV3bFGgS6OzOtV5ZOhEFOyuZ3yDLNj
EgAYVZotcBQaeejnBz/2Wix1zM5vVgfFQc+2Zw0QTFAX5D0RZHzFTxBVno1sCEWOMyBRE+9HDzx+
QSYDQlnKRM1OiqcPDMDZon7Z1l0thww8MhWtzA4lq8Pz/7F6cM0oTgqXp0IBn4XJjKiRxtBDiOkG
qujWXYhFKUzPq+ZNKe1eYu0so7k2Pto3FQhv80Gw85YBuWSF6ucPK8aDXURFuBMPWPn0kDs9OCG1
2ukUcPcbCkUo6DmLXOKE8ZzztYTncAW4FT2JUVfHkBsp10DaQnn5rEOokKLNGBqKSrr8SnaizOUn
uCpZYDzx8mo7BItqID8WMa0zBP1hGJHPxW7/BVOIb1oIc2BJHelmwFXouGotx9j5NU2nEqO8dx/s
PoOBvEStbRexcmv/LF3sKLc2xBlJ1sqGNHiMpNC5BP1260pMchFyq2NtDdgG19TRJmPJULP6AhsL
oZNE7/CuVP6izjhXLDDxjmkmRanUOAO5Mlo1duISsz5YY3jma6sJFoUWz2vrV8A3PqsK33dqEsQm
MTj5xWrbYU2YyQxUzNZVR70CN4D8eFLix9+G3vPm7U+Yj4PBLfdqJsSEfqBLTTYUIkB0DwhpZDgR
DPIGiz62naLyfpHICCCsYYG5jkTbr1kgGczjXhClTnpxoapqs46XxBBeBSi6lUs/53tpCxnx1jCL
SnsG+BtaEbrBc6e5I1lot5af01bVEC8h3haGBpKEHofD1c8GXpZ1Wot/Usil4j1Cer1wj2p6tbfF
hZwgrV45adcnyq1Z0qmyfWwu5jeTowUDEBaHJLJ2t+r/RrWoHtsP8Uho9BZY4rX8MVLf/+Qe3K6d
//i1J6aqTVBNPTFdjBL7Uvgk+gGsMDikcllIOGgNVdsmAAIGbk9SbfNcLjGuuXlQ46IBmekBmSfX
yZiGFlSYtJVekR6GDC8/icpqJjGUMOWDNXlg0Me1HWA7fyErn6xaZWxZxzHyMNG9tUsS6h6orm4h
A8iCCxjbLxuodXwD2kjpi+AVhD/IRnZamxlLQ6kKY1wKTFteD+E27vqmH2YLLGndN8Q1Nk9i708Y
s3Znjt414PykuGKwHt1fR3ZNUCdawkEwXUhxsEuo2XyFM7SIdGh27hrFNzXWGcec8lpnJtBVMvR9
c85FUNbxGcY/OaTosfCPiPA/m6Qvm1azyH2j5mUkQG0HM5nTBLvj9ShMSlEicS9aeN8lkIqs4QeZ
hTlsN9T1Hc7DwU72sFX0UWHrwmS/J2+QL8j74ml3V/Uf/2cSRABx4PPMNUj8BlOGRdi6vSG8Z9IR
zDXRAayuQ43wMNn3V0jWyPpPTHp+lxH8lUExGbdYGLg1zscz8aBuBtUnyAofKM0yRzsHk7MdOr2j
kXlNgr7+Ik6lo/IS2g0vlQgJwzC7fKYFM/IPdUDCZsL+mipVOkwtGSnfdU7PfaQpolUpqWsO9uqG
fCHIHMoimPxhOzl7jP+3tR4x+N5Ow9HOxV2Dg6T8i7ENyxR1X6qSFfOknKQrjbUpTiUqqP3FbxE4
04yk2nOnEy2NiBlZ7DXvi2jLMZznq7axWjGCBxLLhBzULRiUZT73zWtXIXs+D69MfZp6UsEuZmLU
/+K2ZM1VkZk5SHtIG42Ltjq1L+mYLvW7qEDLbXrgJxBiLJBl8C3KToYEwnGDXDn2X5EJQHsPGCbH
hLPGbWZqp0FpZZwQ/dsDvNeTXadrcPrfL052p5pNFobzKkyQMPXab/BV+K2BAYjKXPdSve0kAX2+
UaKtRUhbBWofVJQyfQjjhpSnQL4YaYoZHQaNsOOQkuu/DBFuBTeR3RQiMGS7SuQChGgi6/Cm7Qlk
ZSFPPBj5S8RRKj+clO5NIKcEEjN/Llc8kRVII+MPXoiXk4wxf8v7tlLVr7aTbpYI1bmeRKSlKzFm
Z8rjOR4EUB6kx8rKv3rlnrBsZPeySzghOPiSLzj+SSPLl2A+6/DGWPSqRdyMLXZv6rJKxTnd3/Nx
3umhqeXWzVc2HTD5D0Gr66ccseB8n2OfwawuhgyBdL9ufw0xTgbwDGc6K9MWrff9z5wfXo03qqbe
0yJ0M8HhwpE0kkPE0gmXq+kJBzzVK37idGLXKrAp3HI5lzJMPkaws6qzGoZfvF0Nn3RQzl3umdH3
OqOcXCXUJTuXBI/yr6z9bwbPp998/VUQBJVCIuYgk9R5k75KWmSmahvi0zHfmKi5VsnN+O23Wudo
/F0/tNkWDUpDyxAL8dvp2syBGG0U9wP7P53T0dDGlTU4lRhQ0N+ILl1CorWI3QTxi9uIE6hVm/il
Jx1uilASRHNmRA3nvj5+9aBQfkPPjzfR5YsD+wB8jnmaQYvsiDeVy7xjFQw+2JUVplScY9rjnJGp
upwd/Ln04NIRU3tVK3IearAWrsgF+fYvtqim8mjh74pUJxksETEBJaHbR9YTxkgkvi6j50KG/vwL
iJ9abOKyYwN93jsCmdmtpjW4aHUDs3T4Gd5LlloE8L47OI5Wksftiq2kPZ/fZr47P7Yeto+aSorM
O1AQRvWph8oWGvFXrRUjucz7oLWzNaKhwCC7RedfnVnfzIJ8OHz7KbexYpc3i0QeU3V7jIA8XYKh
zo5/oW3Fy255RtLV/68H/yx4yQ5GJDrywYZGEp+F4ZYhhR9xWKDWrqeehpI16EipzX0dHFyuL+bE
6W2NGYEz3EGtl7VFrQCV3SSA/NBlrPQjZ9C1AfklDPxRBvlMxnZdwpc0ejLLYrghu/t/Wskt6ozu
4ahT2czMQJxWmUzWL8EgPpk/TaNE+y6yIEYh0DIMuRMsPN12a/MiJSnL1+e3/hxE3adnIMyZOFO9
GvyZ6/hh9oYTE0ZpbazxsUeDZurZA7zWO61b3q0XbdkVQ/nngd2wlYpgl64mM62iz/TXuGgAsc8O
1ykseM6KFABj0bnsO4ytqjViLnAWxRJCCjTe6Vn2CylCU1eL5J9vLW00y/MB6G/jI1JCybq10F5H
3lUWM8chUBFj08Wr5RYAt7Ro8EzPbY2hdKMXbpP48LSfs22W/f2+VGikEc78o2USZPLVo3Ueq0Cx
lNg6H9aLO3CnV6DBLUcDMNpNO700RrheFe3jjqfjO17zPEHRJPdCI+9+rxnXhZm6ZokGQfywjFOG
ly9KV0+xVRmBN9ybzfYteC7Hle7tEHNkGL3R4jAc8ed++ru5GpMEOJSagCBJF25cD2AXaJEe+KX3
NJXHIU7GtF7WYpWwgJIPtvYLJHg=
`protect end_protected
