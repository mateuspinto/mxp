`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
j4l2GClVhK00lZSFbmDsRJyb4mTIS7wLXWTWlvFLwLQ8TbYCPYmoonMIktF57eWAI276i1Mcweus
CyvtckvRfLgnWrjBQT8wWxBMU66P5eM17Jpk61MzmP6wz5nNq4YPczViEADv/iSWomhW50pzHlVZ
oLOj7ScqQ8/nHxmX1yGAw7/rni0g9BRbXF64wuhHQbxC+2AA2Oee/KBa7/G4KBEQRn1sma1DpWzS
H3WtDiWWbYE85D0Lai5XfvrM8SiMBtaEu7sq8hz7ocUXW1mZ1zh8I+yqJKVni5q23pXM44PJb7cL
MehbkV2WVmYHRIdnj2Atu5+SdUgnBI5RB8D6yQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="vcIrgpjHFSOcvWodsepFCLf2yiKooGYdwgBKXVatU04="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`protect data_block
c916P8eoeybwaqt0oKvCzvnwnvbTLZasMrjWeIu9VZqcB4T4wysSco+vVmdlvGZsw0o8nETp6bNo
rfv2+jWg7uYj5EayxXviSg1AwU28M4iVBTPSDcp3gZ6gmVZGwTd0PCIs0GTqrU2GgfX7FJHSAAwX
3a6R8ZcdslbIeWWLUtLxYyPGb2p7wc1+5E+QUSN0TJW8lOpBGMEQwlYg9vcx2TMtyU1INv4vyU7V
iLhtnlEdHS8Q2Ff7iqO2+dw9KvVRt4iJS8HAAdDLFIC9DNGg7sTRTGrzzVN0CPOmoXSp+M8IMIuC
8fR5u79LEo2pt1E1UKXyORKUPlkvDrf1HF02B8Qg4gieTYzgVCMiS3JbPMnoXXVVfwZyaJ+5u60a
adosaKxI1dqkhZHDyByG2RDA4bVHO/mG/BUbcKSxEs20sJviLbN78+EpojLDHgugH2p8SYQz5s43
p0T9nBnSkmrJRQy2UroSWuUjEssKkPL7QXl/Wu8xzbht8yunhnnSatWe1Dn7l9BHEolsOjnFfJre
Nr40/4zS3ByIXa3nmalgE/8H378cMc7tHlmSIcJEfDXYa7wW7321Ai3A2I662GVUP9ToprUW7ek4
rJ5X+Jlo+OJm6sIAwaAGGjp/S5OptrHUYSg26K6tKTcMtyirIC2nS8ntscNKMzjNRciPQLVv5cBW
7VHdazFssTqYwMe7X9RnoG1lXjnOVWlTWCXTCo3i/hhFQxHlywUa4/XskJINsD5OlJLUafuftJKz
STT5p11T0Muy7BOQ2EwlwXdiVbbVJf5uc6Bd0E1DLLe6+OW0sCiBqNTUEalfIrrAGqIOvO9Y0E7d
E+HJ0Ubxk6xHbEY6IhOfFFyinaf4KhcB0k81lT0xeF4K9S32UmSkSpWdgAfVbfv1/IT93OnOlxvp
TEx4gH2uYdKTPWiQ9MIwAfGf8cbcG1BM+q8l/iJ9viEJUPSFeMgeX36l0uVAPoVr/zIhJEeG6pYs
xs48FsSnSBQeabm/sAaEijkP2gepfyjpUiaCfZvr3uxm5nlctO4lJNWiQRs6Bks4ezEnWgaaFeYl
Pc/9OfYTf5Y3wBKFdxYEvlAZJV4fcp20YdDxOYo2mx0Si07HXXPk3kOSEIPyFbuykn8fJztqdFbv
usGufaNkO9tZi0ycU0PC9MEU+b1BXYxDjZ6xteDjAjEEWnx1CqIP6TsY04HMy5z9ctPzrMmm/ojC
WvuYB3Er1j/XCIEYM3/jbqfk38tykwFE2tB2cQAb5d7pYqCfGqKJmGsQLMQjUtJ9kddJ8CmBnrWZ
rtTNwlYaM0HTFyOxcX1BnFbucZ30W1PdOOAciJudx2P3xi+DxFyjlw7nmZyIA17ziFIR9CwDZy9C
nbGoMGG5Y4NajsThmR6FtomJNJjSwXwIIcYwO5QIqD326K86pPo7kgafPIaOWLvznDbh8ea3St9/
1xNQNmQv7LrbywToBAJ9NFU0bE8aliDkCkaadJuSSGTNFKwobh+qYXJSZEbYip1QqFawURW68nCJ
MbXuQx7iDKh2K+rg7lCQvE0gkdpNEk5EJ0mzh1ckDSs+XXq7qT7kc3e40J2Chh9TLYMFzycuTCQJ
zDcbZJ61wkcX/egZG7AjodFlR3c0jFSVrsgv6l8zZEmV3f1ktz5U0s3GOLmO1cUlVlqgSpDIRgYj
NpC1oBbC3HPLsD9lEfXZaEBGJdZvqdzPunEaPXQdJlkn8Q3JcZ/Qlxuv8pOKWsPiW+mUIvC/RQQ3
wzRk73/7wzzF9QJH84+5C5cWNVNGXgtWfSql2W6hAtfa+Gtyk7lbYmdahmRX4GfJr6cD2/woC4cl
LNKMr1eJc83nJWcdE1j3q6gQW1Wxh+gm5wHTQKaXpldZirPIkEHqJz7igpG9I+TvmaMFgNQX94rP
pBB5f7RMsokHYSf9s3x0H/tyPwiOZtyLiy5M7B8kEHC+cQY6EmHgHS0+IjI52jdGZheq92hJ2CRf
bfC600+ja/l4NXMJwpjdFiBdORyHC+bq1j7j3XouTTlJI1ZwY2rWQEXXVUL8ACmt8hU6oMRO0I9U
967VI299FA1hFxYpukP3U6Yt6mFoOwCLHvT7bmrEBsplnR9/lRvjhpwgrNNQ73KsDlX9O0bqr25U
uSA/MQeDPwPuR9NEGNKGL5FTb/QfPuW/vM878q7ZiK5AQ57P3nNzUynWI1/GYTgYQ6RiAbyeU6Bb
kAGhW/3vf1DU+oLPVs8p3kd9zhsk34gGffUQvWoQCYGmnRZXqN2Ll/d0Kpa1sauRCjMn8Bw0oUdM
/h4hLS7KNdCgAJJduKYqvZ3QGGiZAnzT49oXPkjZVtUmYmdFRDlYKlhEScTp6sUYhJiMifsx3CS3
8voP4Nx51COK3BGqCX9N5nz81vlW+qjGCfAO8bp+h7HvvUNr4cYmxswI6mUSNjtDkbfo+n693SEg
WtixaEGu+G+7PyKGe2Ozm64IyTKuZmXHJC8WMTCIqEkLy6+i4ihai3+AapB/WQcxLV7Sji+kC+Fn
8sebC3pyEFnaaZQsbf9qtoeqUY6EsGcngmGo3Dqoi87YBaTLiS1r5PeCUK8AuM1/FYMPuePVJpNr
siCCmKvfIjJzeq/Qa6IUhBuFnh1U6JN62GvKxjtC6yRC02Ia/c1ag+s5xrUZZNvqS/iebHJfD8Et
8MidCTxjlwOzQhrA4Mz1gI4cgKJcfKnjbyGUztg6pn94R8wRFIspuRWPoIR4w4vf+ToiBoVjbJOt
ORa9PmzC+EJ9UhKoj53MDT2JJh3K8+hxuChjoz9b835Gk6grJbkA4ReEmt6xSMnk68uvemyyGNnT
fcRSuJmcLbGjRdvoARd9+WJPLIanMEpT0F0XX/aOkoQXbfRvsDP+/eSHySy6CzpK48vHp4ZrRQJe
OU4bZUrAyHs3mEOmlF3zUkZVlAERSmLApZWIEvhZXfKpPmAlFdXzj39BKo1odkpXW2wUrh22bU54
k0aoSqJk94cKJ9ETNDDc3VoUXHrlE9vSxMiwYZcXZdZFjlUJD5og12zt56b7Xre+GLCd3u7/9sSR
5cefbdfyijczAEuxKHakPXRimmlgjCEM9rWXLLKaFHfemiQ4wjkG899gzWnjPBOrV8MrRbY+edPj
AMINqllDz1SEpmc5oao184y+MNuyk3rk5XUP25vWQkHZhhauSIvbMP2avY6AY521qKmH7CYr88Rd
chzCjATqa+1JVC+YzqE0T/8TegGE1Ec0rlRfO4HL+9+pd6+YAALPMjSPRmYrS9va2iOLu2hwVU87
Ip/oDpylMBSg4kcrqV28Jx7U0WHFhPfrtt0EzqddyNLDxz98omnkD2iPBFcpw1gHzvkLeTQNj0bH
5e2lOKbeJFVfFbMeea+R521l6/pLP1tZNW1BNHa34z0CoLk+q7urez1pKrIYFLeu/pJwh8oNICCX
xrn1CNNK1LvyoGMoK/Pld8xICqhigugwNdknjLmzVcSrMs2UxpbnzkNZ7LPVYZP8Wmc5HE0DdCkP
uSmeXfmQawUbyJ+5elLJnrAA7xSs2AjlBjTua6U7oaXFkOQe9Hw3TzTm4U7CwZsRBCwCM7IJPZjA
N/xNEDpPvTmZylLugevjcj+u7mKVruzbElr16PYde11z7OyI1vaxx7pqEIgAWmeNWzrNkd1lQYpA
8yNe9GmwQnA5Tsj50VTNi/kaYO+PjQKUKqtzAvwJOFJbJHuAV1eQv06e824dHOGaCB3SyGXYVxwQ
0enhWBlLq1jB0osMekJBOosBmRpKTV4wTD8Yz8SLa0t+H1t+rXTG+OGTqg7nA+CVNFdWc06Xc3Uw
xzL2RqELH5xBU+e6kn4O+mANBRt04oqxblIULWVP1QvABy0QMTJLaQtR9id51Qxc69k/hmpiHSV4
wawjlvcjlBbEP3itEEvEw1TEdKELlLu0+wnMqSVBZhms60J8w5KwclxCvUTwI8DQ97p0g+DMJ7iE
03wd8PNsNwKmVR6PGcoYeW1thYPN/SHInV7hj0fy/FZykm46tl1pI0CM0hIm8UPnNPApJvxxKRfs
DvZRPblMwbRmkuLB7zLs9MNzwYTRzaz8meLqet13tFtWqBEYd53z4pJ7OqoXinZ3eGIFq3wHH52o
fXJZO3Eqzjqng7hQW5weQzs85T5uNi5KkILxdo17LsPnVtJsry+Zm0UIDGgLu/bCc2/3lwz4k+6Y
Ok1qy3RI52XGYtLppC6xWLQdXI7ZGo+ZmfjLM8d+bHD75a+CJbLq8bgQP73sMPqkl3tikQBIQ2LS
jHIE1kQMGZZ9uIV3EAx2NMlfgedE+d6ky4XkTLDeYFOGhQMtjGUze6nNLszT8Zei3hKzWnGP4u6+
dJzHyquH75ltcIGuvniNtPW8aqYj5F62ylUAnKkTLRSx1n40N1JJ3ki1efXJC+ykIg6l4enn3WwU
nNkwHRD2Y1qNFWh+ZH+Pg23a1QnKGYZOhn877u3bsTI8yrasQlPJuvvqhYzk+0eMvk9k0PNyWi2j
jvNxAoZq15MWauVmDbyyRu0+F0SQji4nWJ0sFxN/Y8WXifjqmrNErswXi1E9IQ4S3lBP8Y8rlznx
MwzMUMPbuWzTyOQkB/GpnemvUhO9Abdx65ksQlvD7UZJsMb15qotsjEmcRWikF4fZukDpTluX7Yk
xc86l5czBYAlxhPjE6/Zgb3bB9JaRBNz33ft5tkUU4PDRyBEa/Z5+saf1tzmb3lnwVnQDuzFWKEd
EVOpe2Z8XqrOqEljk8xknpjXyIwCJm5rEi8pF0Jtm/3M9US0rxRSTAdq1loUMJlY6qiaAgBzEtYG
zD7GdQytjhl6gqWuLuYc6XyX7B3lAy52m1tPg3iy5kjmtA3dKW1VR4vd0b/rOwKqZJXHP+leYf71
DYo5Hd1iBLQiFJq51SnWjnJq5X0XYNWccdecbEycqU9rc9IUxL2Q+pAIdNltrgSr409iQlzhbePX
d0ryLDkz8jjYT2VSrxfXr3au1PEkr57I5Io0AXcRSwZRkfoDzxVadTI6IGpY3HnZ83BjJYBIUBWQ
blLICLff1vhgcYObiJqotyRGby8UeN5U1w2fOkwLjEivDfoWvtFsM5/ZfBscdq81D2q5rBVDA70y
Sxx20j9lm6F8lpC7yoHvRdyl835B56XZ1HbFPZoeQ0Ti5LSqJ15/vfazslqE2MQtlAdc7ix+siEA
54Up/4czARL+YLCZDFPynHCV86TZKRcCpwKONlCY3a0hgohlgh8GwiMRk3I42cU7fWb1BZoJBPwC
teMhh4Xy5H/dHqcKvVMsQFS0zi8bYnJw/f/kvDIyKLzC2BALzpdd5R6lIcPTv2ouBUZ/CaEAiyKS
VuqIE7d4ZjU9/5TXw6a2XCGtLa/w1evoRp3OMLIiR3iPBQbCylmnZAW4uXOTJUTQz9MQQC/Z2svX
FcAIsbX4ITHD9z5UeCvthMUjivcVjV9tI9nLNLZ7tZ2VtXFT/sm+WYpc1NHfsqmDe0FNVm+Cemx0
AzJdiqp0oftiwaEn6YRVuNGjhi+0hpM0T4G85OJ7G2Z9Dd9JTrlFzxPEDf1TdqmXvjTn4x+cAT95
o3O23yEc1+2C48u0CRZbwXIdnVj6RX8TVU4yw67j7hJl3pqMw11oQY3NopM9g972uRw3ogMTSAPh
OGSukVpymFXCig7lOU1fKQwlKA86qG+7NhwIZ1j/BvgAiFUU+aNZcVDV8rJc5HdEIbnFdOqHe8Fg
sF8z4NFPuWhEbLHopMEeAkf1aiA/TRJS9vnYCsdejUoP+MHBYV7GUCu4wz6j/e8itkR2xF+e6fE7
ptXHH4q+UkerXidxxk6dR/sYwTMqbdtGxugEgVrNfZpoVM5UWeIMnkZZwhSFWg/01wg/w7y+v8M/
53kkLXjvVpyeq1FCiMREMtWZkjvLjha8vUuWBBzvFCJy5LflqRM6/n65YgG4lPq2IUwzKrBwsVb6
QIhl6QK7YkyFoMFJlfEWkS4UmZzJDiSorJPxXCvyW0yI/Ckvswyy/5G0Ekf6m5VLMymRJfkObXP1
IMb64f4OLeaZrc7znaBCdF8GrT0jEEOwQDzTurTunMjBykZlbf07yZC5EYb54m306jjtPeKI653k
+d7uI04tPBZ945UTR/+w9x8GcRKbZu9p+/pOUXhu8MUvCqIRO72hwrWXSWYi+gUqh8CkGBNdktSB
48V7+Whvqj+FAtg9fNv0cZlPFkv/m1ZjbDZnYSGuTjJayNl1U6c03uVvK0sBEYJn1v4DY2pBCEa1
hwxdTFnZpc9ETAhy54nptkYwosj1TmmEpT2bvftQhHwiFkRMYdXszqethhWrhGBybnBk1oUkpnSg
8vKxXjszUcP40VFLmyXV1s7OUMTfDzl6jXYntKe+1rpXXZldZ2bkiyuFMAiQi+AnxrCO/k9Au/4M
vE0xLGf0hUKOt8EgM9n6rDbDRptEu1hy+XdfDSCb1MLIJZ470vDjFTXqnXoOuuv5Dn6dNhpViv54
qU2hwGf4u7OaSansD2L9g7MITXnIk0W2f7GmNztWsKGfFpiCMwzjhyOtHJgZULarEf0pBa/bh7bF
K6J+ip+JqWWqUMFVQnqPd22Iha6XefBTTQ2V1pO8DalNIdLT81roeCQUkKQOCplvb+eclsI/aZ4a
FOHYiTDvt4wWYw9XagH7ZQ/uJpQoEHR7zvfCxquu8JvyEsn8zGfV2x5hdQJSvk7Pay5l0CQcSbgY
EmzJjiW1obLJW4s5N+4QhuHQj/JWMtY8ttaXGjbH/2nNNtVqbYKCgfN7nXTdfz2a3AFj+8MxeYpy
jRAVvQu7W4eoylt4ie3Q9rwZw7yput34aK5D4hgWldMW8OlbzwSuohoDHXsa5U+lSUfR9Y50alCJ
XsHJ1zjfmr+piLKvX1kqVEdhjzTo1b2nVdQCAwFhwj9jrhEEhFcNuhrtf+h6FdSWSlO8O3n46hiL
Tj2cxx2gCrTnA2yKbw0f5PhgrFQx0ulPaAfDPV/twrfPfMYgB+6sU52qTYPV77JzotbpKbcCnBmd
sWdFRXBHxqe/kMUY84w+Lu606CwH2cuoADaXeCzTS7Nl/fikRuKNNpEfDYFFv1eI9J+rR/jDUBBn
mT4oygDNx2QCVWtAZr0bSE5O347YqdTIaiXqkY3ag2f+oNXP8aPCOLlZ1nJN9iKcirdoZNwVCVfz
MQkJOr6VKnHCnQ9A0SvKv06cYVYC2PosqM6zqO0Ft9yrkewVj915TpRnUY184ktoAL+BbICNVc5X
QTOhVR3zDNSIZk5lAqnZpqN56+t2i8KqYBgJDQJZ3amL6s/FSayvYdtXwOrCUOONodBf8igBy/au
9T7bLqghJ2ncYqxiVqL183HxVH5roTRX7XPaQlNrRG8/kEpuh3k5LqjaPY5FmR0E7gM8nheyQ98a
l3mdxi6GzwO/Js5CsXIcOe6Rl+fqQscX96a696UZyYSH9I5JzUZDElieVfbSTRdJ++0gMKuXbWcN
no3uc2YwBUUjhQVGRhYSuqW4zV70MQGh7YAy3aPM40dC19WPeC3WB+qndd9LczJHTyirDT27PslM
21l7lB7qfEbNIXPzuI49PC+Vrk3J4nth3g1FDY/AuA/adK7gJ816wU7LufbfzGY0lv4rwZYvXgNF
f/Mh6Yn0vSxqb/xmUfFOJHo9xMZZaO7shLqp540IOu0CYNOcpSju30kwxnHc/gPX90qq37S0JjCG
c9VNh23+im19nVULG+7taf0UA8V/8wk/TY9qtKR9t4CCP6KmBFPZAiw8BxUoqilXzx0/Jd/ZQZPf
R6yx0Gf5rB0ocVhj70qfHuYP7It57wzvkE+bMpmpv3nlwvFwhoQkyiAQK5Tk7/eONQ8hHdRpFe4r
2PSk3wisizDcaGkIXFlh7WopQRYorCQjZnUQLxvPtB4w6l9ViPmSCB9eifmMVnNVDM3XuTKs/udQ
6hDtWViBhtcOtSJH+ajXyRe8NQJE1aXbmYYAlI/bomYEa92us9X3ZKrQkGor/MyRKaEe8f8rOLal
Qw6Gjo91tiltlRy0RMkUoqOqrbZ7//1d0xUB6y/MLoBUYIBPjQsx2+KZ8oTE5+nG65tif4K+Kihs
PrAze7HEpUAXieZuu+o7kn8Gy3DmLialCt1kETiQVWtGrk2RMT2daWCZmdT/4GLhoM/J7WTPi3wa
6ksYxMrcFIjwER+IC4k6OxeEkInHHOYxcjHZgjXkOHqIMfMkF62aeny1TVZ+nsFrBeAMMusWKRaP
JNOqW359iH+jIjyVwD1KF0h6QsdMwrfkHeLlzFM4LiqpdS63gw+ZNeHBLQgpGXWv6CscCazBAAJ8
scB/8e9vJqxPAY8f9IyckIs+fBjiKY+CtV2u6OevCsk302nEV1FbOSnLQpmKg5JPKYWzFSbd1piv
n20bjctdYZue9/Nc+5iNEuk3+Lf7XScaI7d52B6fT7bhcC/x+UU8YtBFMW6nuBjvcHZwTXNXuCfz
PKkAgNZpQhCzjb80xjZCqCQOgxkFK3C1OYYgmTi+E5hMdRBTVlHge2CZBThaHMGcxn3VqNL7jCMq
iZpQcYdWUEtXwcvD6dJJe+6ZcNh4HtvybNecqtLHhf6e8neN+UbO/HIpsCcOrnOgggmJiWWiL+t8
msq13FbNty9Ig6XP4gkTIxl0KbOhSZSe2OFjKxqzium0WG6T2mIXxeOIm4nzomoDAxhLzAzaTnYg
oh5NEklKA4QUMXO90bPIBcVHOd8h/9LVOMDjYHnZP6flqe0AtHPs+qWApDHb6u27/1tATUKsmECN
Sy/fA8XBVubDJwAOzrHVlG1KlKpDo820Bt1Dl7MBqNX02PuUQUNHDNO/LbOgXwYk7MstShU9PUZj
8JhOjBn9UOc+jJUDwc6lihj/L/aOyf3hBhDm8TIWQrfbBIm/8FoYbjKppUQr1p0E6JwUIJvPzw27
wOggtQpzPWjR6LpVdREPtxJlwRv6kfv49P1L/kCcFO8Xb4tqVKxK6kqSOACZFQx/4wdZjeeVlFYO
7w2JUdxTxLBX7tcSFgUtRHe3UazRelVhJDBNUflSjHZfMLdptmsiZfHQ7yknFux5iHgxUjveRujf
jMyM8/106TynzGFenIMvH9XOKUOREJEhGWr2s2VbggAY4Q3uaDBc63aQBg8k+4LWHYJR53rWbVZ+
XNltKFpDshlYLb3QicRpS+18djVgtXpcImb8wEv3sk5nHjGujnqZgDWG6nGW9c0KmKSQF1FVpLW8
uUlWtumEFIx2/0R/GtS3VCV9rmYTU9QTHLHapH6R4Beq15A1lUtKh1Lk37L0TZa7lbdLr9mvrvJO
H0vG6M+vZ92TrYGssXXxVgUwh8s+ZxlNzfzGvQpc+MTftbEx2f2Z2arwGeN85COEPNguTphhS2yc
SZp56hKQ5mCmYsqUWXnEP72c5O+HgwikwdRW0iJUoFnPjZh+LxudBYEhHf3OT0Jvdp6gezCS4zn7
e+oc/juOMpsBwFHALHDJoCksz6j3OzmQgbl1+1X29pXjCsv/JNbVZ4hWkX1MbUo4eHhY1TQ8HQyC
fu8GmIfHiEAi36tgGjpdFcdXdvA3Uk+UANS/u8IcmGIZMFjbD0aDRQVDUu9XueGgmReMXvNMgaNe
63Zw/xZufdkOCCn051c0pplj6xK1eoiCxAQnIEjRHhnCMkQYmFvpE20Di0LEoRmXnQQCpE5161M5
P6plFZG532/h6V+xW/C4c1kVwCZ08WZKGDK1dFx01W7buyTcDP1n1NMlX29ytlrVZb8+yJbRI/T0
DZuJi5txVE5gnY3VyqZXXrydETNIkZaXionJJzO1VQp7GP2rFF/2hH9gUl92M88wkMFKYxoxGK9X
/UqY1TnXHNfizKSsAwhamFZMhlC+MOljRuBp6kzd1/iduhQN1/aTs/0bKXhh4shD0DU0i+fnBgCX
ETew+vZCd2GCZrGOrRy45Q27KlZ6/Va+6xLeCWneaIqcOe4m3Dq+42fQbKCJG0EsWIBjO/hvLmOm
DIu+dPnzAMOCv5yT5weVISWgYCLjWM2USdclfxTJhw8Lrczme0lilrDwapVucvwe6m8bMKOB/tki
m7HrRzIuffhK7p/BBleVLMT9CkW75Bk6wqTlMZYIcRtHIkBiKiQEz0DBS0mv7wbk6RtawlumLtwh
7aKjFr5FQLmiX+PeCA6UyV64C5GQ6iAT2qdStGa4kN/DFVu7TzQNR7WW00dmF8ETxPEAl6i24iSo
0M9MGu7d7VtllTTlO196yn90cc/cCZbnm2+jyL0dporeI2ZjOYdSThSFY6gebSWKpQvsB1Ao4OAe
mnIOqA+dUkbEKLxRJYU84g8WTtZOi5WuccFTOut3Kb1A47caW+Xi2ITsctOBsIMK6J+TPvKx5Dh7
sTingZcezJ3TlHhykjHvuWb9CRQlfo9rF/+xTuqG69afvKMHq9zbUNOZ7mMtNN68L9bTdwnfuZhj
qTCwCdfpx2gs5IrG51uiAK2S/BUE64h8niwfuP1jyAylr6Gz1DSxGjih0b+lWBKhi3tConVihizF
2/n0KAWUloWnm9wtKcu5ZThxTltoTZtQ0IcLf/75I6tlM6cshhkxqxMC+hikJTjk8rTt3qFcLc3+
3oLoTLr2KqL510PaXKlFFB0+m+U9LJh/OufqOlfJmJxyJJ6HFLN+Yfzt8TWJC1FzS2OyPh45gRi0
4K2Ehdrt1WFiPA+kmUarOcD/t9HKJNCQZJb40H9AqTNyBeHaDodSkKJ5iSFKsGW/aPtUXTUS0yJO
RwVFoJ2ea/zAjKeZT4XiIWM1anSIy/4YCNoncP7gae7fMu58nXfkJkS2NmuIPJZKWKYwWKuIphGJ
SgfIqqUZtceFKRKQiU4h4mgsaTBUsJSuL63ZSeZFZbl05uky8200AXtnQSSNJa76tMynt6l9Q1e7
D9Y808TA2dYB30aAUowYyEKhBMTw0AITF/EiTI9uBS9M22r6V1mg3+cK6JlAXjpn8Hu8eYhW2hPe
AiQ8Mzhu19nPq9f3VPuuWK4rKZuA6weGKHqI04WomgF1sdLHpdlo9ru741Lm7hT1QpaTFFQWm6JS
5R2YjhVivwrNQKzB89iydp0xlTLmKeltFhej+oHTsmiFCN+a7aAb2Sb8hb74mDE1dxn733I2OjN6
ipe+HrceXyAad5XPVAJv6HT89uWBN77B3DRbKb/XkJaoASGWyUUnyLM3nu+pSVQqosPR3g1Lcgvx
LG/j9sYs9HPfzRybSbQORy0IIxZYwf7KPUoZBTv5G6HJWtfZZjx1sh1jB72gJC7ZHusfsV6ycSIp
uS2vlE91Tc817q59JABKhFElaDDfXxNKjBXeUbX2hCRRGSKMaJJ7nXnU+WmRNSEaBz96k0AqnrH6
W+TgkZrsLACyclShABkFjS0/Q0TLossBNnhlnEHoP8Iy7Bb92HsZt7H6yhVDR5VUSApo1jScfW8d
K00iLc3QMDHLRuJEbfoT4vc4E01suTlK1KPOfuEwUebsGsQLlvlk/4QttkX2OUNSnUlN+pYK21wA
NsyxipmItAkd1rnhLZZoamlkrjvaGI1f5LkfBA2j/6z+TYnzCBcWITe23a/sC/ov93d7evleUWgQ
1VIatwkPw4PfeWiF0Fjxtxm86lfaWeS5UFRW09qZEcig7uuHzzWRdK5W1aPZLpc5C9/PufeYoBT/
GoZSUp5xPt7Io/jy4LBzU9bFP4wMaXKA7ANacQV/giV9G3YQcrVD60mCSPfankmvamheCMDKh3Cg
o5U04jHrx3AFcPw6TOySjeHwsxWv+H+C1DRreYNzkfT+DqvIEBUSxZ8bBHm4MloelPlHtQY3uJuK
xu8INHb8hJkviLFxk80zNDGr5bwLaFwMsNKsZOR3AK9+hXjMZR6QWBeSifnHwn/WUEHliN2JatkA
fkyXU17nbc1YCQJ9hjadHMCjqHVA5CO0kepLYa3bBjG59waOasIFFTNwQ7llVj5OEd74h6EXJZOI
ZIjd9l0OO3aHVKZf92Jh5YQOffBoIZhCVQvtcY/2F4WTBu7NLVGD+Ee0vSrpcNgitPR67WmbAHf3
Aj5sTAvdgWYaQLt/QTPmqE/hOz95sUpSa3zOc+1OEB694VKCXNqVVpclrO9xhASDf7w9YQCNEy+7
ZhH87274jntTeQsoyJz/I+nNC2uPfx6GHbx7eDquvxPtpfe/b0RVjHEd9MAQDzDcb/4ynl7nJtOQ
Oo71jnnCMgdVp6FwBtUUwaznvzRhu8/BrGHqngM74Ry3ML+MeFSqDnTLJmDuMsBBZ1jfMgssnQ9O
T+nrf+Bn2hwI1hIygJZRtKDBmGcoogvm8zZU8RBvCpfcTe2rcDidA74xRo4oRsUDVD9qZA29/gwo
TxgJTItXSMtBr8IU2ryUQWZtaTS6JqFPwaUdHtV43oZOmMs2BQIOV/rfnKeAjYrJ4p/j5Yu5yaSf
SkZ9DWc9e4HVGPWbyNkr7yyXci3V8phmR8NosIB5UKy+AVZkwutPbnK44pdQMpUqvrKBvhY8m7Ic
uhdxjQj23TSuO4C32hrjm9GG7wU+xt+hZTQrocRN7Z4uv637LEmokxh+oV6Kzx1vYgKRuGQmENEc
cKzKvylbmoKqPQRK3YA4u26h2rssZQBy427a4dlXfMQ0ApYkd2dQ3eSx7mGPKphIGocAkd/gqhra
BsL0QgRQsooPGmIP46WPwZWeqFzgj4YhHzwd7TtykpR75Pb9sTGP+JAVYlZ/OBkcrESStbBrM8Td
6QlhIBMsRZOsQfI7vnDrHzbGW/X9m698wJidIR4ey1pm3m1u69au77/1f9QDrWRd5ytJ/5V8ttPE
a/OI5b7StI4qNrkXuyA30atFRSABD0Tudc4i3woBZoohqQ3oQD3RVtRuYfk9rWMAhtx5PCdnJMsi
e7VcOAe5Oh1C+w5Sdq/tSRk19tvpn0PFgD6zH6lXkAiUfG56EtHZf3otXG1VO4RwuuaAGO+AVGmh
cZzpZP59SXlHkIMo8WR8mbtjtzMapA4z+EGoGY/KcCHxyRS99uNDM0auhNQiQ+p6BgkYuxqtHgYV
w5dWJrSRypgaQUHShRdKsZSgxPwNuGLgraw30Ibo5fz24J5h/tAEsz2kvOzQan5Ho411GFkJldsE
VKBFBqtulOaATnUIs1Q1CmEWV/ZRb9sP3LJRqyi/4H1JC+2YlTkG6fJZx5GICFxvvvGxk0LHAUDw
Tuo09w46tKoze3yr7W6AOGbIrYEF135T8ULItGMRRNFYW6kPAZd5+wy7RTeV/rBKGy0gEbBXceLE
VhhsJKdo1oaqnXClEacmphgC2Hj7ZL+u/KLCnbBfbkNkjHN+d7G0sWY83oeXCuMNV1z6YX5by3RE
Cvzmaj+1/XQHoq5uozw+KDIUL3OJ5Wbb0HUD5cW1wchQU2eAfpekpRiT8mwacY8xLDdVn4fQqni7
ElHryjAB05zqsp0bq+/fBMtXPHkb0igCehwBb1yMRGgzzxybG1cs7fCCVgST6X5fJYDcxrtZw6lL
+phHIcPKo/PFEIIPNVnoNubxpWmrx2AOJ2RPJXUCkGmLqTnaZ1nmBVHF9vFTcsVLzYFU0mcZoCCd
xADHFchPpCcmDszbi0oSMdW6lOO+7znLGO5M3W11rjs/GCj9jjwfMitw1SCDdGIi/dAUiowYTt7s
3sMpfgsYXRNxh8ZTewd3ed3euQdMKm+lr092UeBmlTyCpGCmYENg9f5cDB3gvUiXFizgiZ3AQgap
WAAlkL4PydoY5lJtWAklOBaogNHQvzm+zIJtshEfJQkzj1Oh2n6vT3fmjRZ2CkR+H3eRSMZT+WSF
2W0Xy45LbvkZAHAUmXEhSoGhT9VIQrqC89VXb9pE7Xi1oJ7bOrtH13p/f2udrrVtJ+sBB32PMhy6
832YWsm0xRcoWhJGkAQctkG2RDC6fgS1AtEQoR1TIWZ5zrOJWecuTVcrf56ns+k0fAFRjvJ0iIjW
w6PKv7XmxJoAXgHIwCrCjIHyMD1m+zII+aT4FM4F51obQRsyTBJUCLNp+YwhCOMjNxVfoGYT2fjn
Cj5WBTJ9a4g/ASPNOYq38aSxvNopPEWcOcTxQxYYC+J487/TfI36YaTDXsmkMr6K4PB0AoH1cVRb
MQwUCWSZPzBbh+5wetMCYMaxpshatiQw6VSAVoTYj7FkdNniIiZHAk4WjP9v7966wA5jL3/qIgPG
xee64F3rQj9CdejFVIDpvu1ZRRypDeC0VdmqRG9UjMNPUDEHEAqGvodbBvBnnOcTv6KHJXceacvE
WOKhQdzsa3b8NNfEV6ah51dpZ4Fe7i8Qv7Kso/3EHrTvoSgcbe3hUgy42omfPSvKybcgOY8wF6LH
YyOdmlkrnnNUP0Me4fFCuIk5XbGU1E0EOA9UzAxIEadZ/UIzKJXe1K81MKHChrH3dA9dLq94qAGs
r+pqdmkGABZ/2ZzFeMsbKJEyEgCnGUBdHGPG6oG/NKJTd+FGqzibiIxgrow9ZUcDPDfoQCV1VjwS
RTAxK+4aYJ+iBmMDSEQvo2g8XiMXNxKk2HJli4WnUh2ofKVlBcgWjWE8BPIUpwti2p7gDm8xwbWS
mAqDcGOXULV7FUZhXztOnTzopmZP80Aautk/Cd18JKO04H/DcGz60sshq9FbsfAcFvId+1ceNZeU
ZkCiPV0pANRfnGqbbu+pgDFkGs/z6HFVG0P1GejuklNIHraMcjVMJE+uRkVfdGLfXkEmtxb2+14d
xEiL0gREoesaxe93TLkeRBYqAO5+xyBLDYmi7Jw2Qd1r6hzOiDrH5V1Hl11t0jq+kRFEyM1Mr+Qr
KKWnw74wVE1+boJSl5K1Lb9IcibmGtkBSWXLzHigEOYf5AHZiADHRuYlrd6of64FWoUf2SciHOB1
eNWrlYf9SJuPc58y5FNgCATK6XenEFWD9wjDSrrYk6zngdjdNQdUVCW2+D8dK3JzoYNUseaDxqkD
C2h9cTP8zXi87WHQL7tnJMC527Ye1fCorwjDR/JFAfeOm+pkspHqd2bniWZ5Pia9xRkiv7EQUJnG
Nvwdgn5D9649bZ9qzKmKzJj3/WQ2XfnHngvBTgHno/OzUNXiV4v7jPHY16auCSJmiGDksHCKuUAg
hAEOSMG0y2bMobjeTWgRC2QVDi652GFc7oZR9oPpv+65sI6EKJ0XNY1i3RHdmfhnEyaPby9ABzA9
X/C5lZVvhWljEwWakfDA9VgV8Cxvxmf69xPw5UyhHs1TwhriktQQlQ6joeycj0fUcSKBYM61Eloo
oDNwPKlLa2IYlIV0DRlKg/IqYiulslICfEyai9rtmZ/B9+uYLewMedLzMKpQpr4mCuil5WZlAGlE
x9X8so2TlymNIppTabO1AjS1aKoXQqZAHJ4Lhcfl1z3Ol0XL6r3UZHq9/pUORDTFbLqf4Y+Yxhep
ZFuWRnvTFgbzN0NEzfpc7sfuh6HkQJTUIr2D5G6AZNq96AGyioF/rhW6SzvNkKAb3o27+YiI1mGY
1xP2Xj5o0PwcNrwuoaLkpKjsZCrVEK9F7tjD49na1oZHM9WJXtMdJEYu2sE53pK+9tLStHgLgiQj
swADRjglJbCncO2ZqqlZ8lPs2w7X/9ov6DVrbPGO3pfmuhZgyUNyrvd+EARtn5uQ6aa7wq1ADzhQ
8VUMkIKxo63Uz71D8O1wdpCXT8JUEDP9MUigF0p4exmPE49dhmw/goj+DwbFTIIfiksroBe87Q9Y
LuG0Kwq6KabWEhY1vAch29dPWh8cirGszermNOq08mz2uI3C2TSZ3MsKpOIF6aZ+idQtEpl8NNya
NlGy4FpHTb+peKVvlgnVpiWd8Wn9SQ2oDLCQ4rOFcUwnwpjkVCiPaiSznlLffVbFH9BAMfYrKo9U
vnBPpcZYepwK1E8uGW7MqlHftdWaHntE3tJjRF8qBq7Dny+4VuS9VwDlwDkI/5wa+72JRy0B1pDs
NG7mzpTtzKlRb9NnLiWtfACnvybHPQ3GMJlAjsinnTqNAvceveNFKD7sdVpYdOB/0Z2EddGfi7IK
gzqm3gwC4812cQFWImo=
`protect end_protected
