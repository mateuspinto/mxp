��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{o�����u_���Y�:�_�� }
�5ݿ�u ����<�h��4�o8k�W�d����8�ӕn� i�����"�G���Y�a���!R��a@�4ŢM�p���ߞ�suN��H�H�!s��L�i	[��.�1Tk�E	�����rL��O�tLu�b��:Zz��i�-��	��������S�4C�HZ.�L{�B��`Q��M� ��D|8)� �S�Y�8�m��r����d!�:��S_6�k�9{'`u���Q�=6���0aT��mWZ)׼�^�r:uV�����_璴���I�U'
eʤq��`��%/Z@+��&�K�F+���9I��)�՟���&ʌ�œ�O��O�*Jio8D��)8V����
�����k(u7�����7q?�'x�?�`��e��{k�26tY�|�2�e�l�/'ԣ�"�>A�d3�K����'���=T����$,�bDxۊ!-�L14���Ws��nd(cm4uE���W�k'T�⚭)J�@�v�jT�g�N�����x/��_���Z�=�ǋ�B�Q}�*� ��g[9y���h�T��l�''�=߄��3*Ű"��^��ԱM.��q��0]�����`����'?Ek5�y���y��TY��=����#����3�x���F�x�c}�`����5u%F�Y%��6�J��5zR��l�2JΤ�*6*p֦t��#�o���q�{�חY�%-Hރj��G�X}|F�I����ڌpyDkO�֘z�o���n�~�������1`=2�L�	��C.ƥ� ��x�i%���ڈ?p��|Q���;����R�xo��mpi�]�ct���������tupK$��{����B�g�B�C��?���B�<gz�9 P/e�m�*~�2��t�6Wp@>��"G��q/�9ܘ�����=��:$�x� S�?�$��f���	�Sph3V��X~z�[Ht9-/��"rſ�^�БQ8CZN�̾R_Pf�A��/�����ތh����pq��g��D��7��4����f<,[������>8?���Yl�_y�ǆ�e�*�\�r4��u@�NR�JP����?��AӰ���x^2����M���ԟǪ�%rf�᣽R�%�iqɚ��u�{i��!�Z'��P����fsm޸ua�$��8�OAeC��Z˿�sB��Bb^xi{� �hbˊ��+قX�3�UG;�zQ*�y�ݚ+Q�	̿��	��t$��g�f��}o[���Ħ��]J=	_U�O{o|��x�,���{��$\fSȢ>�|7���~�Q2�!�U+���Mĥ�m����r�Ǜ
�$��Z���H�To��J��Э�׳�l���r���hϪ8!zx��~���;�%Č�����gw��f�j�V���`�B�1�:���iB4d�A�����<O+
p�*�k��!s-��@5�L�{=oʢ]�?	���� s�=,��Þ"]����5lNKZx�}���t��^ǻB1�$ ���)�N·� C
͔div�E�&�&��̩��ϼ�N����҉ܘ�=n�s�����SaQ��'H?�� 'F� ӂ㹚�,���q5Ơܑ�#	�	����xA��ջ�����0] @iڛ��_1��tx�ҀL�t�٬N�yʲ=ɢ?�Y-2����jG@�;&��p��D�����9c�Yp)�����&U_3>zD�c\/�S���g�<v�K}�V5�26��k*����KF].��S���Oy[6���`�0c��� �I�R7F*/��:r�)��P%1ɨ���P�½2Scu�눽�a`�}����ýE%ߨn��D�{�P%զ	���+�*����ω��]�Z�G��k�D���r  �;�᪭�{ϸٹ������?��Z��]��z���ф#z]�el}�2"���0�QO��B��EĨI�D�Z��kA��w�����VL�Ro�I� ���\V�)���\S>��/�u��>Q��Rr>ze�G㠾Z�!��jP*�v}%����񈸑�*�b	��
ף�S��'q6�T����3Q�K�X�e�R;�g�k9��ߓ�P� �LRdH��