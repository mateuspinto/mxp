`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
pK2KSQA2DPANt1RB+kdDNVTyJEPKsFe1ebtnI+WCsfgSKaM85F1gYcdC1d7him65iiGmyVXZWycC
tW/NQHmDU8kQqgbZJ3xPqJXtJnH10+NSSnDLeJFtgeja1INJ3fPwuf3ftn9yKWMjnkHixbd5ZGar
efbEvfqAt993uNjiSWoY5SN30vAdQ1mp7BfUgAhWatFgeUIndP9JcTNJkhAXdIgB1Xh39q8QIdeC
E4cdl1//PuUovcuEJQP+5aruAYR78RxndWaLXLQTnMW5ocDmfLI6DQlLu6vvXc/pjjJU1WpLgRtx
KWMUljyGig6T7L/6XT8tsubZQpSit9lrnLjS9zVQ0TF6hqv//hR6g3HCoiUdxv5YjluYIJhLJRKq
cZuAKuYeaqfZhfSyX+lpdfYoWFL08vHrXfW1RWaZXgXEqZiUDz9oFzOiSZA5QvbA3rz8HvzWN/HY
+kYcdQTRvFqY4Z0pbS9pxZeYz0z1sTrbQJGXXOxHN0OyrlwDKci/NN63YBVsnD75E8HEzSzhj2zE
6LBYwz51Jt5DTXoP9nY6hxovSzvlAZ67eTxPkcCBTLw5A9BuA/IK2kj8nhPTTaJmJBm05yi90Kyn
575eX71s+fAqhEw5mc4F9XBTQ9Tt0OOL4jmIzWBNMbpK/TZEIkS7/nlJU5mYvmHOmrpI/VzZqImk
3f2AQblcnXPS9DAX2RkiNDpZt/qYNe4II3FWq/ccnmo7Ckx6WOnPLEE4NKQYurROeyxlIxmeem64
JEOUhd8TvKk+SfzHLXurFjt/Dk95pcUAB6KJs2zC9ll/MlV5fyMGjOGT51WL8ju/TklYeMIhD4t2
IswtJkVs4uO1w7lTh2EXrb5sL4WUIa1QigMKrszTbX4w2gnc5TnlydwfFludg0l7R0MYRu9RUZgW
HJqsWi2vrOtp6SL88okbs9yuR5PfJ6tCRU2IkjBoVbA2ykrth6oDT0U2MmhqQdZEISTHJF7k7Cw+
/RBecTGoAL5sXV0/JO9UMVAT/+J7Qdge3auRzVG2TO0n6xsoyFt1u6ox0y+WYEhgXvTn3mv32llJ
79UUZOoxSr/0WFT2DT0/4GJ2aUF+LSDnmrWkfBoYCs+dHibXzzVKScr+EWeE6skveBKejEae8wiK
3euryeiDdejYR1RU/TKY+OmjBUGdpf/B/VZOjqvxqmpZbwrpOsNy/JFkkBGXWAnZ6ae+v6VzTDtk
DpC01PZccyNxoeBmd2LxD4+yT9wJeEvGnbAE2OtqYO4frIJjJ+RDnVFktrOwutTLUS4uYRgp5wyY
t8Iye416yLpki+cCk1/Vfbsye9dOcK8FlB8hlnKa2Yr7ii5RFAGrpmYvYHGwYqNml3uk/khB/qM1
138Yfx2vowZFODoAhP+b+h0trJbyR33BpYxXHTFPcdq/JikmEHgWelfD0OOh2AMa3tjHwIoIcU8t
m+k4dC9WrsInKTURnigAtzZF5iLTlLR3CrOg3SrQb2JnVscYFePLEhpXF4bdOp+hUhulKbElzgim
zF63XM6Hq/sh6SY0lCk5tMJt4gau3A1hNid45tqkhW2cWvNmgw61ebysuJH0HKOEfBwqN4mHj/2h
7E0tTwCoT8fHXivD2OV5x6uRqUIKl3FQ2Ck4vRM+IYF6gP/xsGw7ESqK0Zj6NNApqR9SJ5jPInsO
WOQZ1v+Xb3bANqMOY/mCGLc6nNXlrs2qoJnO0LxVmvb4uVN7hBPbkxAAsJPkiEw4n+o9U+h71bnQ
a9Hb6KGzPpajMloXd8fFIvygFKHXM8D5kBRQ4ILzGBpXCG9B4EFbdS8VMHuJOjK/UANcxS8q2ode
yyF//0WQNXvLl+Y8MjPTj9wBqYNmKzR266BomNMA8/OKkyC1uI/oqc8Qrwa9UIWgXnNMZiIkfc31
2kPDmLxZBuJRy4En8BCs01Y+MBxawfXy4XpDFdCOXL/nin4LgXgsxEgXxyHroWeKr89x9+nGSiIc
JP0arE2JZbHnaspe1zZEdKjjl+qaRxI55jVgFJ27pKvY2xYDTkv++VAtZL58ZlE0QwDrBJ+599qR
cj67y4iKGPAqIuKhJUc2B6RWiLwACIXyg4I9dEvGXhwCaeGA+ZKYQqWQuRDrxMumDP3s18YGjwkh
TAEltYKX5QnySzLeacJFaQCDhWQBlFVM+BNYjHEgwkgTqRP/VRRSV3jIp2XHaKrIQubAjlrgKGiV
E3Zvfu/sTzdysXAdGN5yQAXkP8E8FjBIIZMcoY1UQT7TW6YbNImt7nlWErDNJbyfJo0v7w0K9RIl
NAChnI2nYs/YRvN+dmnqMREtp/MLLuDmR5OrLVYiGOTrjc2XuT66Gz0YCMvE7qwDGVu9fqEEb2j2
YU0/0WHuC85jwdDPrqZuwLqtelyrKQ9QF5qvKYsaKWFf4VqJ37K4bn9Ajbw8cCAw5yzLTSnwci1t
j7Nc4NzFxI50NSG+V02oRxIJYWemGrjBRzZL39X1YQZa4KfQcGV1OIkEmH1jLp7gp7+saIafa0r0
K+ewj4nlI4mcjO4OCGysbsk/Q7NhNZd4UGuMEN1gd1oNfazBxvUuomWkfBbr1O+Ea1QY6vMbSoNa
LrIaQmj14Yl9ys2O1Ap3j0XqTwCik7aOZFEW+v/Pfa6gA5M7WkHpl3KmT3BtrNWYzwj54kPh7fbn
HTph7RVAsLb/nQ3t/sV9Z6njacccmI0QNW/+YuWP+Eslz+icF9QUa39CFCAGXNwJrbNO18U8oFYQ
Nqn6Tl/FlAAu8Yym8by8DE+a5TSSwl/4Lj1qDkhzSs9c9toYIWx6DLhWzwnbOPtfrvO9ScYBX3ES
RKfmmgCL3GEm1T1dLLAaFQjJf96YzIi7vU4Viw1N+TDSIqsutDuni5w80cInl5WM3ci9zMkYBDLZ
kV42gnJpbOwpaxRrTkBGCNtaCxOiUkXY7q4Sxyp3nOqhF4WZhwGwewXFV7IMcHKHt8lJofYhaERs
yKO5Q7pqdbomyASjXNcRFTlJ0qa7PVm/0Kt8JoZU39sOOZcC7k6NCd4R5NQ8BZSdibiweCNbI3ui
7qvNGKbtt/ImB9spaMvYt3obfHuW6h0aWfCtXYIoOK+S4dCNckG2Ql3MvUJMxk8fTP4jrXM8c3rx
CtgBIp+R2jYDaHQgoN/hyyczoC0okePs2PFcMRv9je277ehoNme+9wPUwjm204mvoBM1/pPI4F1q
0dKiFZXj5500YnshfyaINyDc6FqFXw0wkPvJ/Tgl1GVLm5WN5i60wzVSTzx4Xz7JaqB8g1x6bc4d
7cFcTtFQtNhQ6NGshnE7MknIRSBXEQ/VWomdp8TQvP84mPjyYrq31CDXNRaUcbfdSWHZtbSOWOqL
FXtAuhGHhoOR13XI5hYbKT0Vj+s+XbnrKaCKywOa2PgJ0lEYkz2YMJyHyLE1R6bMZJhZaxro5vRR
tcHJX6qX/fcS3S2jTinHI97e4TMWNEgHEKKWi3DdALiE23es0WUI1jpiEvrFPK1jx8KS/oSuY9G0
Zdjl353sgIt8xtLBzJJPOSOEyTWJlBNBK85sWekwE4jtqk+uPpwH8g2yFULWyskMvh5QMfx4Ymx8
tuDNG/kvA2S+Z6TzSihVU7Zp056a2MLawYykJV7RI8cB2tilXI3cqi925dGwcP7oMH4xjWmi8c9Z
VbziaITAVgd+GKevsF7F1jRr97aEDxfL8RYBhIY+cZPx1m2UysiFFnzZvvsJyfYdUZ5Ju5jP02Hv
pLu9W8hBLJXvtxj6Ynu1zXfwQtCwQS+81W9ZbdCAF8+BQPp5v9bGgvLtZUY+k+f8JJ6MDrR6UyXs
LKM12UdlXsEsB6y5TXlQZbXX59NmLPtNagpM7gPqSKxCqVKIQ2CwUCc3FjMZSZn0pZujqIrpk5mr
jKR676HuTefpkhK7LwMtIH3HsvOoifweNK5I96b34qXd77HJRMWqB+xqvudSGryK6zO2sZSyQuJi
EuLlUMU0eogGVKi3qrOFl2NE2NG6y4oCnbwBoGsOfCj7oLg8qHasHn0mZPOosMDQja8YYYAj9WFX
dpYACufAcSWLv+u7lNNNAm8W5MUazdY1BzCIADr4/YRV6DZPKTj6oq2S1iGZD7XbfEwneH2QWi/9
lOBYRxUz2Xyh/0x1giM2c1cEdX/J8IRRMCUWU5ri9fO35N4zRWTP2qDdiBjDl2srBpQW+kD8/YrB
B+ZoXdIVKTuTD0JXLAMXwO6B0vvrcv6ZdgFWnvl4IuRBJJvbLfqp2ZbLT1y9fE4+XJim2H585QMK
AFznX+fw5lxrhSZ+N9hRtAyXyZSYtL0cwNOlYgkw5b75TN+STpgMGrZNmThEVk5+7udZivLVVozN
cV1okAhq6Wn4L8pTnE+q56VJLXBd0IIspl8UGkprnboMKDcJq1QNAmZlzybwJK5Fh3JgmofysZy7
/xpMLHEYyD2ImL0QWRoRzCTpNYuPYowRim8uBAiXXTbsKioUXcQ1I53rNS5+c3xBLoTG3s/tPJ3g
DWlVzItsmAamigMMbujuI6f9twbOzDm8FxkDjSIGja7qN0kEJfZTgXNqdNG7CL4ZtM8u/Hfnv1OP
3ktYJAEXwp/XTcelKjqNyzkWk1u6GQ24dq/5DGrCozhfEnOFgLmFuBEQN1vTFFNgcLsVzofLawWd
JLLIrfBrZ9xmsj0v4yQ/ZvBFPSJqgDbsfJM0LvANBJxlSQH/3QG/xOOUPo4nHEkdlZxw2M4k3MZT
hpvB3jFKrMMG2QwDbkQjxgH4QMZQ7f8W6/BK/MIHDrnj7WIaSo5IXY+SsQIkY0gJZScr2XkNEZDJ
bIQE1A5aXDAVO0iVJfF5vat5O93USEgy97qOoAFFGvA+e1YWY9EahOE4x19b7r1cDKfIFLL0VEbv
3RzOhOyGk2GYTGdVuSBhXyJNqEkHC2/QWGtH+we8ph3nnzjuCaiwDFX/JrDKDy7p/eU7yKoJ7AaW
fAO3u7HkaDG8rxoSKliU8FeilZdrb3P+Q3A2scntu/PjkXGupqq4V7sasyBqhYe+GFFUiO4bkIAE
zXGAprdE3SV+uODPc1aFzOl0XaYPFPLw3NHuvba1hAUP/2MBsolmRYDlptXi7N4EqWbbd/WKfVlh
5/iA12jkfxeDn5NW4IciHq97HyjVh6rb/UJrai+D2K7+iFUOoFtCn7VPECz0EPsJ65Lb+pMKa+6+
f/uI12ZdHNI+baXLNN0ot3tu8EQ0aT/iSoGaPCKR5SwNbf+IN+4GXl9uzvGFF+AWNMayTh1rLDyw
BIN6gdSiD3A6bj+t5JLhPRqMSwi9pFlT+Mw3RBBqkYVn/NuZ6xDeqkpMWcI/9YEDgbIF3YGfNHMk
HDd+q3xzmHDrTFMuKOfdIcHFpWHYi7bFUFmdeGACcJE50DXnKsmL403OCDwaghpo4Xzs3khIyh0A
yalIFeD9bCo617DFQF5UbSYNddpmLiEuSrM1IO+2S8808eUuKHu2kw9EZR1ETVUgC+KSYVqX+rUQ
U36HWlZZmTCWO/AJfjP+nVGq49Py7qI4Rr7s787kV+04RCggspiQy3dcEdobGnJXls6/ZECF0QF7
MkfWodXG1ZhbJ8eD7Nlk
`protect end_protected
