`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
0USWSUGxovGsyBJteYpEofJpODTfrn5rcRKpdfedhoYWyWArL3Ro+rr0dvYJQRSgX6pLxuVeeG1s
4gSvG86qhzvGkQ43ylKgoJVreJFZQvYYpfEVShnKGJJa2QXh7QGFe7XtSvXv5hQZ+xFJ9RKLYZ7a
cTarv+LaCasVJAijqzVf+eLA2Wz8L3i2USeCrjje+qDrg2QZgVel8lqj4QpjHrNyqOB+fsR4eLOH
CQuq5SunXYLW+nUz9r7l0ivF/AkDmDZNmxrnRdoJDhWcc4U9OIydJADIFqUQz5ZIq+F5R6ZUOznp
wCN9eUihGD/TBbvYk/EOdN2RsUpAGWMXl3x5It2oFvGD6VrudnxdT2G8oOCOmHN6ftwYwmiBT45T
4BfSKMD7pXXJ4IhhlWCetkArlGvFSs9dqcpPj9mHsYvtMYUPQvME/GyoGpds7Semlhkyr+VnAxPM
/5bxRrYSfcVtG70FcriDUob4gA22I//p3fIdrHBsa1n0nnI+TO9NXgL7QR5+DjU+potC9V6Cfy7J
3AqOvlYtuSaN6YlsCRXjRLODlmfCAGwNsruCWwqXCK0zEdWHKE6ii9D5yWBHuzvnVca+XB7q6V+7
Ak3EvCY1Mb0XH+dkIANLeA+NCNL2XRUouIHk+bwgQHxeYwr25e+TNNIiwZCt1ATQdqtCJbpTd2eb
zquK6Vp3H5tljiFAIZ9QwrU1kEiq67SwRQACOTitQgCb/0eHfWxVZqzUZGYObHwuXe/RyvU9+dx3
wvIoEMHCRVPHoT2Fi4iMnB0PzBLPs1vGqrrEuvoB71Mdg/prWmAJ396QP8TYHyS1qihkczoimfIb
N27RdL1cdjt9DZmyfdwkPsf+nJQ9DQI6aBnq0hT6t5IJdfEwvRmRjh5AAY7vRr3JD1KWSUkpiUdU
TqAlx2MJqRK23B5n5ncGDdDgY9y5slULYfGGvwi5/+6kDjQdVtzkgOWNXGxhxu9E71MA0KYrkhY6
CWCkSeg/n5VYtg/x8lpv+M6EVsGSipeSiz4t0mvEx6FlwUDbR1vkZPkk08daqgsITIkeuUlEyo2n
nAy1Ow4N+F9xOVt2OSohgph+BEh05SARMSw4I0SpysyJT8QbV3vz8T4+bHh9m1ru6zwO68Nh8x95
+AmRfWXtlDmjPcHGK7Ip7VARanOUCVk5qLQ9Fq0708QGg84FRztVGgELDDqUdAu7QWIIRVIyUL81
YbNxLYBiGuGHzn4lznnPniZDKr8YHXdT0zQHIkX4BS31dlAPNqd+h+NxeUk+NLWQlvAST/mjJR1i
EzJry8iQoX86gdpAyDTsktgY67OQRCw+lrvPj1vKu/xaDtzJSRA5DSVGAROUynWTAc6bbQdVhLA8
+VWaTsTlUvGReAhgTNTiQ8k/Ct3pfHQCGQb19zOp66OOjDuug24jHuZly6pdHBC6++Ix78wB/l2m
OuoA8/Jq8nNFpumSkq1xJyd1FnkLJdicwILcknOakyeJvahlJw7gLE6HG1HhN0O6vdV+z1oOVquo
wN/XE7vQeIx6EOWqzlbJJAdLs+ii0RNRTtHBg7Bta6cwCy4je9j6aXBsowRQe5xDwBIZ3Fgj8veu
a3Ak/390k8JxU8oVeDPvRnABng1+9ke32Tj09rrqrl1qsKYbF8TBlOek6ccMXEl3ianjmYa19HC2
9sz0883uXz2q/iI/ffbBT4c982AXLLZV+49nqciJ+FB84+QxY/oXOefrTlfmo2kMbJyU4TjvLdWq
DrhCKaBKRJQMDePzlut52u72cgvWHe6rN1d1pv5lpAOFE4x2tSgS8gmVPJw7HOVmu/6sOnmfTHqy
h7czLxwHvLapD6N6FIGGH/f/fMHXPtQCrUAsokLyLVL5D3qh6vQed8PnQNOvkVjaEc0r5R8tZ3UR
bDgYFBczGA6p6Pn1nngRP44w5bsxtiCPIAiC4SM9ZDxNlO+nTNq/dV2aXnAg/kaLsy727KV4nNmo
gILctDWsg4HAxQjvCic0gnqWGrJCZJAEe/gyhLCoNlW4h0LJd1jFlbuNfna9vDHyqjquo+agofU+
FajmNizT91RY/YrhKJBG11GXLFrpIsVmFYKa1JpSCHDPQEV+MlucdO+erPQVCtuwQaTlnTZ2sxi9
WkfDepeHZ5YTTCuugxJSUk8aa66qoyaSULw1mjAjKlYHryKwAq+vKhVckyHqIT4po0kDZ+jN2ayq
ici/aiK0vfMsYab5y/eP0jZfk6ZpCY3m4zrq1MQnQ0on+stZT019aMKMVEVlwkq1xJTo3yMFWSZd
9+P7UraikCWEAHpNFRsNO0j9H8JZXpzD8P2ZmHCUbRgOQtaLvVeAke/5OLhKXX7u3nr2wEGVkSFt
mN3Y6J1kb3k1rQqeetELVJSb7VI3y0iqNK6Iv4qlq0mlPAPU/lObNXGop9YAQxkTUr2i+BaJUw98
AbGMRUq/pJ2Xk+9j032K6N0Svs7PR9VZc0lcUqli6VsOOkspItU/qHRD0DhkWeJpSKB1wQYjvG+Y
7sMh9jWhrcbDDF0P6IKd9YCro2ABd9mVq+evYwIpWQd7y3mfqt4fM1ilumnE4+M8LzRAXUYsFWFQ
oWNnI93inejoq0vKVO39DN4YAwyRGymR5i55CQcQ1moKng1Au5AtnFYrOOCshkOYWqsrNWI4n3cc
4hQrNS9V0fmUZ7rRyMuMeAYm7FcfE4pPqKx6XTFmA+vfQkttMTqxRczKi1HQDGxUwL8qJ6NO4spz
uLWtpiCVRjnkiUFiTfQ+033od9A9p/1XKCIl/S1WB+R98p9z3WqRVosSyuk38F2pfXSy3BWxeLpt
bmgjxD5QhTOujGD0PI31jBBfiiMUa3kL4rHuN6wMkL2i33Vk/8FMWAR62tXBABoCJszHGeeTZnXQ
1Kn4tPgiONyFbR54rhYVOvvxtkis7DlAzsMRFhx5813rfVs4ED49BNqWmDcPrhjDEvfGT+4GiZrG
gh+PkjxSNnEk7tdMj818R+eHz4cKmKR6+U1TJOOwrZI8laO9hKXld8TDE/DU2524O2YCJLoqsFha
aVg4jXQ1Y+hZ6ANQSHnCv10aAOs2CjbMUpy5tk3hjlzHZfVQmovKUGpMniMwLnvqmbabwU4YdS5+
gfBmOUfUCBkneI2uraaZLBRmEV6JEzKlvmJh1QwrAg1s0qVF0ZpKETLYyyuiw2mq4JaGIDZQqvE/
agKPEbeF135ockA9sYNugSd5ppTO8UTyasvaZjGTfgXPP1H37DDqd4Vn7IgtGI4jyci7hCPVtJ30
KBZo+sSelLxbgopdeF1AEwrCmZbXTi/ajAFztA7PBI+0t6XSoECD1lNoq+cuUyQgi4hh4omqRanh
sanVDgvCdec7qJxL4T1V3EuFy9qB9MS4WNt6M7jI8RoQ3H8VnlWprukcl/icykDc2eXsKTEMlh8E
slNtonkSRkGVEitJhUvRqLXgnT67NcmwOHeTWhXMlfeDaESsHkcaufoZ8jeUWRB90MwqPOWNrObE
8gvsaca85nnAoeMTgICzydpQW08tgP2iELFyCoQLbGc2vGX1HaCCx41SSlmGWy25/HN4J9DU8XED
qwFRhnTrUCR3e4taQEGScMF3vZSE10QCxatlSST7gyZYLDtX9w50igtbPvxRqfkkNqptEJzty6pu
78VSGoguBDrTIwB+f1wcap+Jbc8IY21wXu3nO8ePmVmI7M152GApOK0rb3HNzV5Uijpk0i7/Imd+
4iSIgp0HKlllU88fre35KxnuMfBSJ4AGupzTNodzVEZ81TChGMf56Z8I9zC5McFSgHxfrFUfxYdD
O1cCoLXlY+aOUGA2IEVSs2p8cK9QLuYW67E3UuG9dhmcIk6wmpYVhgTY8Z9e8oF7AdVCg3P2zMdd
ABYiGBXExQ0hdsZUAFp5ZjerScW8o+QXBIqWh0iU+1NcNdBSMvUnM1ZOWTSXkW91Nqcj+wuIB7R6
Fz+T6Xq99Go8KbWO3jpr299N/+/mO76zMbaildZJ13tx9JgCsZCbX7T0XerfoxCSr1R3oPf9PE3C
PgpDVBHa+8tpFUj/6/miiWDKKGaf57bAO1GE81CvPMJ42hNeW+p/q5uRXi24zQrec/hK8xBb1EC1
0/jXdI+mh7m2IQdZjYBWXo585bZJrCZ8BiysQQFHMaHXU7z6IBsa+V5Vk6Xnk1tKSEdC6DU6OEpd
QUXeC1mk8oevLB26jTE9tq5wRr0FQYiZwdV5yqjUH6QDXOIj+eApJDmVJr7Ipa2WVA74E8dJPJTC
kwZ05iDU30IrDgzNY/ACGJcLIFT3t7JJjsNudLaHLC+fsGJc6sls/CQolFlhMknuCdW9L8+5kU7e
7V5Z413bS1xpAIY1kVBKxryhXXVYa3PHyNLcTtFPJO+WPOHV2FFCjfZS+Q7ZWnRITnnqHV3emhPL
J0TKtHD9/xJ6MmIs1+/NhhYXDGrCw+Cho3wwSRf+H71kVMjVajkVNVpWXTtVK5wpTC9W6mTQCpiP
IPftrJwvYNtWs3JovKGufvA8BeXGLWvz2UVdSObN1usk4LBiHTLT21dJVo5UWoWIpWu3lB7eBuJS
nB+Aom8jNpoldhohhawjijPH/3kTWq6/1yeEeKXyLhV7i3Y2jdCDOp9FnePHVruyumZ0bankt/5r
zjdl12LzLubVVDxYWNY80sdipv9AGS1Zy9v7KnkxFuQCSqAc7NfcK160QsoFEA2jCWsnmcITw1Zj
bnyBDLzxAxDZavivZrfPh3YVskre8HNmidgNg+6f2jSK8qwp0vBEYK0MoHvod2V3nXwbN5sE4qtG
vKIVUw0jxgd+BeyA1owkjAhrnusjqHVIY+JDtLMy+/0Fqzkw/HUeTaX4WrKo4V9EER5pTEP2tlUJ
JI6S4BNvVuLov4QfqHuH+MOqPFak1hGYl9PZvrrHmpxXGIMJ+MrQmyHZ5oU4t1X3sYyVqFMdnDJl
DK+nYU9ZLeqpOmGkxRImeaN3REBW8NsykQ+/Wjp6fgY4rTj3ALUFoEFKqbk+SjtvrcO78q4OWrGm
NduratecLG92K9+KrLj3SCzfWbml6K4s/5eQQ/JtA5rzRh120QTIskh6aJ/Foq8V9mdFoH9BWbLr
sUl9ddf6H8yxWi8QlAAmJ/ibZxqta47k0CnsX4obgKagdpz4Oxh9zUA9NhrEHghmsxM0sLNqQAQZ
Uo2TXxZvnoBt7I98rNIt8RamSY7aDNa8A1bshF4alff12nOQRde++CssktCu6syTOYKHn9LlJV4s
DJDQj73qG/0ipW1ONmF3uTS7F039H5ozt53feZmQVYAnat2PRkZ8OQnFpofJufkowzCpm8BK4Fin
3IKN53RDyUekKtgPO93JxIOwbAyepaYo0IfXRMqXa7I5rOZHe/AdRbcIuklifEdvFOdc7imIpvsy
k7i2QBxn5sE9j3qEnc4h8W7dUpPcPKQoS9XN/kbryeK7oX/qmPYW0UpPkc3QAIEiEojXR6B240mF
khoxv2NNwqfwM9unnydUMlGiF+BOlVps3hNz5Rc45/jD9XD3i1y/rPqlB48EHR9XLdPCRZVl4+rp
f6Em8SlRUCEBh9RbFtCkFiGWcKbVbI/jgypz/pyCMCombWCBJiVKgF4QoAQeI4TbLtro0piPMPnq
cQ1xtQXQ5KIpxDsIAu3Be/5XLcCmNfsjbLi5cHsyB7H+SNXFY5yUQp5vOd8m1gxFhYKXvBxUpjo8
hP+9sK29SWm6qdghdHxxBc3xj94tPktOOh5QlJO7FElSAKSWeIVPNPYoavfBR7GlaBUt4DKMu+Yq
MZHtXrvLf9aUARFQCuFRDouF1dRglmC/IkEyhFLaV6Y3bUEF413iOIJIRb652zCX1m3HYn8ytddU
IjH9CTlJpLFz0SufWsktV5z48CCHI52i3wFnhGoQt6+jVzDfd2HmjxTDa/I8Zterg2ey5T2qlRBc
dsKloutodjhKqH/qg6pdK5TY1/Xwh2O8kLra31WsuJMpYodfLpJfKMtpEBwLzlK0vqTvTbBujDjT
QVOWk48imBE92gB138IBSxOzBzJm+UL/ZeZCWDPB1Wy3kUM3YcBbAZgvCl9lhPG9hujuDu1BxeCH
lXhk2JbS1MwaY/sG3bvo01gONH2JB2p/wPF8zgHfopeajeNRbhp+Nwambr3zNo4JZ/2fw5XOk/jg
shCLhAiWE2o5uECjRRLEQRJjve2/JxZN7p/cegZNeBU7AMlg/FYkvRLNLg3u+Wz4SKs0SWKFhyAW
CdsLNBWdLWzD6ZnFuVtJMf3ftSF2fkMQb2HvQellAUuJym0F6Hq4x+QLT6Qsnvrg3skeJj2hzG7e
GQpmxwkitvs/tifYMIN+ngtXhpdQrrVLAgyscBIICnNWoHb/1l7GPT5zcwqGq7LV7XntpGM9i9IH
HxZJ9qK3BCdjvSvSTZmh+2DH0sL/BYzbYNBxT8+eA16STqJ2NjHrkNd0hlqy9eHdHJEgzQVvL4WB
pRBtRRABDyygXV8TTeALCo3213fzzaEyjC8k2yiiY+X0qH0tmTkmJRCUKnusJqghdNb4ZjcB2HND
gbuVbG4L60V9Svk2OMMNS+Mlue+uqgvbdrNJgNpKlACyiyZkZvu+Rt3ZU6Gv5C2LTRnS9SFEOo0q
TCj1JUCSqBZdD2q4yYTLLVAL/VCbl9ht3KJeYdt/GvglQjwpBCNUX+to3kmXKJ0pENh9GPgWjrRV
fg1nEvzMcKYcShwxdnRERe6I5SFMnO5N8gDLfopcs5z8GcrdXgeBslHVkGs6exDfL9q7ENBIbShb
5g5mCi21/hUmpf+8TBryMHDb1N9qSgGB4xYmqcFUmyU3zxbz5/uKLKdmip6YgFoMnf4XbUdIjPJ5
lwnF3peyWI8AYeESUqli6t+9jpmgJdch2v7vEhdpyEuTIaByHa3fYcf3UudBXB/960BD7bhQqEyG
JveMUzbc2plOZCGcQhBznXqnicPyuNTOw/cp7OWxkfLwpQEbw4KqmgzZELHczMkti/ROwwCgWDOD
i6OQYDtdyjFOTPWJTWduXFmVZStjxlD94UIbEM2fzm4ESyl1w43a3HfBsz/S8YH6P1CvfyP8r4U5
2Q+1qz67k+Q0ufRgTh8hS8piPAVD/CWPuwx099nlOX0hl1LFtaxEeGzRqn6o6ErZkt4TSn2QWY+u
aA3fqkiDcS8VaU0X54JTUwVVCg3eyKmLO+4DBJu4BpaGDc1jBAX0/uWPShMzFll3cvGekZyoY+0W
AG2d2OdNoh/C6Oa2vEHvjFQU4112dAwuJCvojdVKSEA7DrjnpbWBWsXa7F8prE0GAtMHQlCzlhI2
OKAIkxP6RzfTDKoEb3DsBhUsk8gfuMTD0iak9Cza5W8xk60Vum37CONu1ZEiaR0GlQ+bS4l14VA1
NfiEnAEEaTfhH+553au8iKOPypJbIVWnJ4JV8P4RWmW0dB85a7TVHECUi11Xo3f5IwnlKbyq+5KZ
H5UrzTMVpnSX/Sel9ABkCFYxx1Z4QQyXMaGOoQLwhFFcp9vHzzhHfEqBGsGFd4+XC/G/3uk2sy09
V9d0gDckAEdrlABpzFdBqguIp32+n8lEvl6lvOZuN1NnGpMeV5l0BTW8NpPZDnHlP4dWP5Qsbq1E
B5fUwe5KvJrxXUi0MIqZuUkey0C17cWdf1d2nBLutVnZhT71fPGyBespfIhKRV4W/cVVh1UOLnak
Cv9IfmDZLNxkaTI9HKMrUvYAoa0kJ1hC5NHsv17JzYhXV3rSf3nA6gDcYtmapzxJsO4wccIsO/pW
LWSrhKWLP0HuAgBKHl8cF5xMxQauW2CqzUrxpqvWayDjwiKOrhlGglbgHPAgKFWWrIdxiUvm0Rhq
DiyO1uMm4ARZVWTrJsyXVsN5Hzb14WtzRCxYOzN6vb2cNzALKDEUgpnpjBvC/VvTfjUu7wvcsDzh
1Jc8MNVuZVJTuOUQWK+dwzHJZ88xaoMEG/dUhnuUoJ2UlJr7pJol2Y7nxijE/QWjI7nL50A0kI/b
hfIxhcfdgHsUHYztk81M1LO88wyeql7AIxCf7S69eDnxz+HZfuL098BCBSsoG20gOAkULWprHGXy
z/ofZVM1glMD2VgZWicnooDAS7cvqoIT37oo4Ld0mTswj+SVcMwcDeNz5vyF5DhriXscSIUupSKv
dKosMtGxeQtEupPpmaMkG64MnTk8vDUdjLe2FMExC0DlnBKDKGUGRJ2hPZROHK9Z5JA0FPoQ+gVl
Mvt6p9ALwHrwqLCOLcBvryw2cJ+QUGdDLy3UzBSD7ltpQJJqxEY6SbSXZVnYlPUyU9jRCi7iaOOa
+kMmagIJwJA9He861UswujMppd/NkD3RUKRyDyW7o9TrjyM1+8YeC5MJFSUDkF0hmBUIWCdpIh5L
TmtNb/XkZX7A0h26O67KzqQnR+U9l/CYV1JkxaT8CeMGKdnOx2RcryDq0ltU8iUyZJw6iPdsPkEm
fGZ0HZ2jOPjqdSPCq45GpxVDNk862IpTXs2wvA+3yr+p1BbsXULQnhaS54EgPf0vYfexpjXjS6Eo
VbIlyliKR15BdDqwrZytu6n9TYxsbz47ivt6VNG5SYs8qrwmnN6aeL3U8T/vzw+biF3eaqaxSfjl
vVzGEBO4m3p1j7YV7q8oI+XE8+DBfWxZHvJSkDIyxWY8TNP+/bOA8wpXOsQhA+jhab16NrAAUGS0
q9YRWuqztzDZXA/f1X2qQXEZowFNjBse6j2MOFnxJypn5ElB6MUubXFCQEMwjUwxuDY2abtDxtdA
GqWKRCMR70xbqYXECxRpnVLMQV2Rb9rPczLas3046z5SU4zUFvTjLxdQ6P+tP+NqDQRFYOdvUPqZ
HQhkAHW+VCpa2RFKICqWtl1oEyxo1o9gWV7UDfQGQlcNh1onlo3dG85gUSwFEKWFuajlRY6sV5pd
bDe66/YEZff7SCkopnO9ZzdHXL1vR9QD56F9cXNxuCCf6UXiXVe6KFPhKZCWI5eYVQE/NRYYITk/
FeGZidBEL30P9PJbPRUgcccoSsvgi0F2ISUMJP5wnuLwbCMgJaGGZYEIrKS9OShwOSfwqZ+PUQm1
PKFlNLEOjq5eBd2W1UpbYfEby/jxDMyCttFVuN2NY9BZ39piB1z6kTRtwNKc591/b8jZnt8hb0PO
whE5hm7vPcTz0YuWzBg1t6dgk5nxzg/jTYHRSUNt3a/xwVDMfAO2aAycvSHuTOacmX0Raj5/TcGZ
jj3ZLLkGiD/XgXQEimHyXWKou/w2fK/EiFzlcvOcfXGDMWRq4hnZ9lR7doYGJtuGqjNWW5sR6i3P
FdpKWFvErfmzqjoSPQqa06imagipVRtbW976DZWuGyfK4r1cKjAu2Bl9SsVOStevHgOvbAkQ+GsI
KSrnkwADZla4R1pMusr6LfZKm1s4dqqLwbPelM1iJxzdDlNblC7YDUjN7c5gX63o1/PxRVZaLvdX
sGLKHoUfRjKMlUGwSHxJ930CMgIo7UfWxqpY42fmkV5J2PcQWkCxNAXvpwVrkd/TtM2I3YG4VZJa
1bYN5bJZaSUhhPcFUtk88XH1iopn3AT0lkSUWeDjIPhKdRjYeChuOKN7v9dg6TkzM7c+9gGPO7Fd
K4/aIQaRQbop1u8A19B8rswdaSh5xFt+0+V4XMNnrRLQGlhvS1l3wl0dC0cO3CmuJY84QexiOe4l
VrRxAoIYcARKXxE1gtipzTHW9AQXTk2i0svzicjna7vsKHA1BvyAdd6KpOlbclf2aEgZJcxsxlX3
oZy8GEDbKgDS4ioZ5lamU2DDWNuIEQbO4Xkw1OyePvpvEXHs6l1XmatS8va9q27EOvrSR6nh199M
+Ki0VGUd9+nqEXNsGm7CNjZemNhrbxpuM1T7+gERhM1y6Z6kTKDtrLGQ9vMz6D4oSFfS2kareqOK
VjGK951koiPXke1KybKrfocsAabCReHW3m1pSMQ6fmThC6cY/3Bvr1UuxWfdfQi2jpl61wYxkLW4
LTHZainPAfj4KCXChyWO24h+Mm263lvVZ09uvod1YOW4ZnWV0CwYHyBZocBDxEABHIIcSocMtFmB
2nErlwqulh/+x4G5yFAG2kyQIkPpxwo5NkwdYxWWR59G8OFmfo9s2JSW2eQHI4gGQVm0RLo6hF7z
Y42nOjRZgf13ZtvIKcztJ009tDur+9q+AWcVtMMOwFaeZzveQ280/llTII3Bqoyym7TPwU96AGp6
T7ldbxwmMq+9YrxbZScy7coMtDHgouKCHw2T7D0pIpqG66Blue9jJ1Ez8Llv8UDM20L4wpWIQxVp
hZV6iHn8QSfQxwUFEB7kFjjOdWsucf8CGWB8hvLx4c2W5yLhaGQzIYwFhluCHRLwGAS9iK08YNqd
0Glnj3lKzk2EDmIweJd68aGokP9k0hyATn6fQCKpzR5kNxr3+s+EeTJVvIS+N0pBPUkSZCMICU0b
wDIEZs1mTPkzyfKbAhsBb9VZ0Wca2gQZiCM8wPJnSf4dVEKaaQoDiBPe3468zomNaUna62wKlxKW
9129fPeDbbYMDqo4yQcOuyyBEaMdmdS32nue+iIyv3tT5lhJR9OKIccRAaEa1xXNM/Xp7yPcUcD2
V1DKqBfA8eMZi4jNB/j+F9C3fnXsJW2fm03LQdRNQgCXtAx3cSh4Qpq2zIHdIoK3JzRg11VwwlqA
fx6C52pap/jKl9w5NL9if/iyjhJ4MPKssadQrI4i420UidL1mpMMRehYt1+bDK1gX1WAckfhhODp
1Yg1+1hmLhSQ7k/ZUA6pht2SM6XVmJRBla++mna75IBk5DoSluhmtLY0sarg2LT4hlkO5eredEUH
WMuvUkPXehFeOcuHLYJ/XOszaUfMqVWd01RxOJrLZ2ND3wOyb0mWrarWw3hw1iihxFoTssgQmm1F
j8tbivIyr6Nyy4Rtqu1jQt1wLqnahnckI5arVN9qZLu1nknhebGKOSrotN1sEs+8PfEcj1NIOxJE
BaqY8J0hXMzz5NNHGXp3IS2KCb4uNLmPN7MjW6UlWVH+tg7BTnjuhOrTFImq7N1FjiULRCDtCr27
enEutAtFv0maVNPX3NDbE7+gnnw21T6vy+uMLe9D78DzUFpJwhQ7AqVxKtBINZM+hoR0WgrjuIpT
aV+In/uxK1I2CbRTcJubJ9gOsFoANIANR0F4GCX2NavCUsgXHAJyciZFQzJAl3JjPEQALR429Man
0hUy9Mtuz3x3goa8CPu5Sz8vsWaV/wiYdj/w7PcEofcGAsm6E94PzVdUZNmlyfJCJM2WRmnGD4fK
mRJJBMB/O9i/uby+8fE2UW3JwBPwd09lLDb3kt/pUWMKWuMZx2QJk2U392mcJx0JDxizQgY5PmFj
st8g40ifMb3P1H0f8JmL2rc7xPQdYy2+Ly5a6ilDs5KMmyBB7tAwo8GSoZVedJe3Dyfd6e0QSsZP
Sja0FSca5Z8cTH+eAnP9Ydbg1pM4MusYZaArnM7YaYUx2xX5QDYVI79gZKk6ZgsSZFdZfj3oc90o
iFKA+4e6tjiT4HySrlEsj1cmg4vmstPnqAINGU40TiI2rQclQto0ttxA3JoijdaOMO9h3AkDKu3w
nAwzNRmEeAL6iL3YbXME/u2fTKbinETXCs0k1jxkaAyzrsoCU3jEzonIJBn95WIeuJj6WdxN2ma1
obE+zrWtsUiv/H+d1Qo9nyzkdEeJG2TjrPwMVSdtjsGCESaaY4mHXffRlNSwtc+mTPH1j09dnpbO
fCdKOhW88jweEkV7xg0PMwjsMGLXqLSJN3n/LBgn4XLuCGdk3yOwnw/vs93prxd517Y1cYI+c0nK
jHWg09jUEIaGocwU+iQw/tnvjxUcKfosdDbsXRl+yYtQXhz0gZ57jn0tfYxcOwkh4p/Q2PgXjHtC
30By996yRY/zaSrwIFcD+afnAokXGIv/1GXl0QnOAsdEiR+FSG1cUsKSlULaiYNp0K05PPOxvE/h
iCE+ByC80Cyp9DOPJtF6Xgff0t4Kvh+kREKYJAZr8b5VrLOIDbmGkIMBcf5EEOv+CMJtfxLqQVSu
F1M884kplJ6TuA2IVwXrXU96AUA9nEtuyzG/1LJtDIPBxUZEwjJJqgP6+zXZYs9rUOSL+LZjYkph
WyRSZFO8Uoi/HsK9ETg+sstJYdYQNAQ4iu1W3Hu0qGnrvJvgbJHX9FnCySSvD+Nex3UG3SZth3XG
Q4jA6qr/4qlgK1b9n4QN5oynmNQR1I0zObTUyLzsLZJTAZ0KgCLFmy3TrblRwvLWvctPMr9if0nS
tJrp/DMzqp4K7XAr9lJ0YpJ9umKoV3iCFFtu5P0o82cjqNGZJGzjRGz3LbIZAe2oRscBempjC1o/
B2VknFR7OgOJrIKTzu2YN5zcYRMwV+654fcWh4GRKSsQoxQJztduNgOoWdyC2rMhF0Qmc9FH4Qoj
JwqaDMfVE4rjOYvnjamQHvTiJmo4kAYrGRqf9SQqICjVpPDYPMVHXgaZKJ6Ib8I41VyacjbQBV+z
36Oha4McL/BFtpYwgTE8JfLnEVc4IuqvH7lbEZbBThIGLORfrf8hwZOHMDg5lI2I2lO/xE5nIsdT
uihBJji5xymUg81HfPEtcz/yhPLW6IhZnce5mWhIZded/Lur16/RdkgwJgxdS5EDBPET3rBmJas3
bcrwO0eESVArhUGv+yOYfq7umQTupSNPSLbeWq7DGaHGiFBUAkF1Yy/LzBCJmVFcOt/x79/58Wjn
7Tz/vl7zj8JTrzZI2jsDgopBXWz3pqaSP706BG5ACJraUTASar/0VUjkwEX77FsMBteCL260dSrO
WkOPh/NaCPuMYBtiBmsuAi/v0nl5G1EHlSIiXeGyPUapjoTS+I2hy2JILHTvbcWv4Yz9/T3cEJ2+
htAdShtQlZdGUCLPf/7JY8n0QJvT7fhKbLbCzLSRbozZ5Loi+oyd/2D+IM70QczudNq5i+0C3/sO
icOjBqWQDvvwn/arAl88232B8iETG/i1ZRpIVXIOdeKlWHw7x1O5QMlgHEY7fWN+4C+icHLDFXBm
mc24bdcs6V3hLmLwbov7jW/W4kuW8u/hmGiSeUzzKC2rMh2oEo+4nZxrkpLzBKiityNFhhTnx6MP
dwm0eNV0UGuZjzUudBBjWRDbIGoAwD4D8KOyfNqbddm1vP1B7r2ibXw0UQE5UXL7Z8IgoBv6cSx+
0It0JalM+7aYVGyZ4TugMCpkEzBYQf3kKqhSHL5A+62XuxUL3SFALGPsTuH0R6VllRA7gQPAWdrD
RPleanbWp//+IwXqMx0I+3bTY50sx9tHjlsQLVQKWh3J5GdV2rnQCIElJddulTtHazJebm1XOBVY
eqqMnCLL7fSnvACSfO7UGJtbZrX6kRvM/MjgPN9b0xM5xOTuAS9k0V0KIZuUEPDR4OaOu0zp7H7I
5M3PzDzHCdCMpoN/amarzFzuGn917l7tm8AJ2xiKaRMkEG8rCEcyFhPjJYKMSnIjf96RgexpdMQ4
F6elcLQDeBDoHnMKDSSIQtX5kgyDgx2ReYRNFkSUo/6dItezKpylabUxq1RCTXojWDFfu+omd9sM
dEEd846wAtbyPdalfB72GZDqXXT1YKJmvSlbfupoRaoml1QV3j5xLEeFzpcvdAoAsbCYnS58wYAI
YGm3gJA1eaZqMRKaZL9I6n6+WlZAck9gIz2sDq16RNAKZ8Y/mfp5tdFGvBgHjs8hswfvrJA75bm4
kuTVpI5ImPUm1EHBqiwM5AIOeh8Mt148iEVBaU8sIbJr5fpM1ojcRalc2YdJ87vLSEuJyNVe+1ME
BbcY161EtuikAs8bNPkxaTq9qmuSQvZdCSvsiOmQ3jZq0dGZ9ss4z+1WKCv2p09XZmSLR6ob6KNV
4NCwZ+9Zh+PfyyJG7GrPC7tuKMKjr5j/RyqUQRZrSZg6+iGa/z/05nD0cFW1UdpLOM7GCsfuSG/i
K8JZ5dSUrOxbCC4LZS9mg3YABqhVdqR1K18nfr9VlsPvqVSWegvx/hLUqHVBBijHd18pkWWVzn8J
+DZlaaoxXEaWIF2stjKkhsiZdJQT+Kd4iGQ5XVuG7K1iJqOMI94HV8Kq90+x/qrHf8QIgqgNGL5J
1dpzHUU1p0eVbWNnFYNVuRq5haC2aIjyi+D7Fn55zF3IP3ip4Pc8sWCFIXNjnV9/zWNpoMtiWvB8
2guBuMo2LOnUCedpm3VKFh3wJzoE3z3MFlPl/v8PHYddWqHUi4oEYOW/aXmLDRb6nmyhW9nu/D5J
mcAez3vnfySYOyKQn9C8/3sM6gaVJzARfuTrs5SuVUxw31noLNzqNNygQpCo2zlRGAfHQgri30n5
Me+WteVLupfCQVL5F230PwcUdfSEZ/gigITYdSyF/BOnS3rj/GYAgZ+iylMxtlPi0Z6JSGataMoB
jFWGGyeEqxTgNz23gTTApvDkW9dDsCte/SGvrfRTQKVY0bRW+CQ9NuRW7aMiugEjOnzujLiHdFxi
ttzBeB2vTwjqeKfFJ68Gdd0kCrgNQrmJAt4xPJ/frktCeTDMwLOWihmhN1onxY00Qq3vgHB02H58
H+0vUjxcc206bP0f7cFgV6tRIWFUEvnk/C2UpV0no4+xjaimXWNXEF38aZPrEcvKZfSIisBaaLyw
YR6qjnFKTXK3YnykqxmtzyQhdJ7qHglVzIr8pib1u69fiss7+kcFObDBjloh13lgYIRLQWMt5yVE
66t2HUv7UZZuTX5HJ5fziQIKGIHH5u8YDzJ45+B1p9dLwkol5bj6KOMB4YvUUNhvPrZQcJwhC9ab
P0YXe6y1BO/zPvD7GFkvRJsV5vnpkRSpWaFfhQfOD15yGA0BKDmG67rDaHh4GsmA7DrOQZjewWj+
JDCyYMycyCx+R4+g/8FWB9ChyrLNpARzFTj5uxC5VVgNOsUlAZdbZ4U6i4uP0n2hupClgwYDnX3J
C+whJPx/sm2jjwwFUC45pdU6X9+/R2Y3kwg7VtCoHXDSu1SUrNM6yDdnoCaiNuZ+kLMkeJ0bl2eF
5CRHYozz04SILsWzBJb2Ue8HNWl6ELm7jyhJB2SqWWy8Ilvw+qPsNA2blyUtqXFY7nECmet5mwIe
okM3LrJmp1s0Fqz/QjPAJ3ZGyhisYH6EaZH/EtyrFVEp2aP6+FDBe/wvHSA1/ktO0Sv1DOVEOyy7
JmigI09wcIj1GZhMmySdZldOJ9SWYzTtsRZU638LeWFaw0JG4IPIE9K7k14rtLvXxdKZsqBPLFba
8dOAl6/HD+vf9VpFTADK/UpEfSnDy/oISVrMrVksEPdThqKiRwP3Q/PDkPPXGuAOnCnVVF3a9xOG
a7xAAVkwulg4chciv1B4y/4kCN/ozGH3AoooipWG7EyjClfrQJlkwX2LN+55hWxlmJP8a6Er78XB
LoI/nGaeRbo3u447FR+UuDXIP15XEN+dVa+MBUOy97XAOV7mv7RuLlzku7AooZu4AaqYFzU2OrfB
aTaSOj1A1a4I6YLpYIJn+ad23KaCzNWgPTvvm+4zmWNBSB9jYINyzBKCWBGM3Xa1uMCaqzy76t5S
tPKa4DEcJom3hcY9yLyT2JfywOcOp4058iJiFnvPLpWwGh5xtTQBI0tamwEL09iDP4yba2F1h2ef
0m11Rvkfn32h2Tnlr/JVMWHfglYLEK8/m+8uxK1tEnNdhp+58rRBsx5i2IdlqcJbqr0Dx9O8YYHh
TVOdu3Ln3Uht+izlEIdFxZBpOZKydLHoX/rxUcMH+O9JG/fiRyrR2rzu8Y5kLFQFssK8rzIVGRez
EOAkPIMvyqFNsjMdSnZOjGrsiMDOj00PA0N070BIBq/ckz8S8Uqczl00yVQuwwnVMDKwyN6TDhCC
U7k2cLcqE+2yh+w1oGgGwErXpeTWrTgkkX5rpPpg1HX3KTYTPdcOIfUZ6+N5ks+KizeG3bCZy6Bh
j4+pm/3h/OKKGLNtTzRROVp9p11PTB8d3EUHO5LEVHn5QNO11NkVUBZWGHjzSmC3a300C0TloJVI
2UrWNUPoBvLaB4Ro7rBNz8GCO8xxTYTFli21YG3WnJBBvAVC3rqU2SsiDqxQUvcwp1PTH4dDEq2F
Y+knov71HK5LNQvkjiXjFPY9rN/s917RwDeXM1xu93LcQ4QNN3S+rEvkufHePYc9eeD3ATFl/BsH
3kJRXom0qMopz1nvGJ0nsBBQZkkCJe8aX11f3WIFfuMgEE+7e8pnbdJ63NjWz69mG4+T1qi7NDcw
C6owz/aNu5Tgn+sloKVah83iIs2PeD9mzs0fm7OEt3M9PZyjgYjCpyJK8FGQpVQ0O4UEdwNli9Ux
NxR6K+gHi/7pw/NE/lwjt4tVUwk++1YWgmk8Ugy3qfN5EXitUOz89TU3dmjmcGSZcw8OAPLhN3qv
7Nt9oLdmUwDz6eeXQjLaAZ0ZN4CEpJSpvjfiDUXNGIAdf5MoZUBDKeee7sa4om39B2zHbwPe8BlM
/Nt4Qv3AajBkKppX0niBbJXQXiEaYto77hgYX+pvNCAUdqJpjcQR2I/x+CVNBH+bWo++njzCpSE/
jjmvFssBnEVd+Yv6sUWqBX0qtjjLFeAVAdxOGhkyzIlDBSW61CKpVyFhvKeQQ4jMBddaSA1wH+23
aVXq16hGLhUPiqNzFB6rflVG/d9kwo5yJGvFJ3zDzt+dSrnA5wQXZNuvQOiUekocwKEIuMubgL/R
vKijA/FCJC3KMpznFyUZ52+ZjIyzDuxjIJW+lvT+XDH7EM+icCkWkxrOUiRCMUKYarzreh4T0SAT
oSui9jBi95pds3JdLszBXQj2yhCmAm904zEBxOEIM50SoFPE1Eeo5l44oYd7OCTF26ZoVsYXVhL2
GDMDZNkX0y5+IqR9V5U5xUV0GwwYaTMKmGCWvnq9gTpv6ytfuCYzZhSJVdH4fjKAPHznOp2BDSo7
n+9FGn7dhEoFE6UoU6F/I4X5tSRHrUwbMA5uOrssVDlGzugf5c82x5nPK21+nxIiNFYHuzCdXf3k
YqWWztNo11LdKBtpuifLeOmeG69RcJc0A1ZBD2Y9611j+xzXOHjdRObyHvm2EFXB6QnZMhGxwm/w
sEsG98PbY/32vhALIBwnOj6V0JazKqg0yTbBQJsvEotJBpHdaa/0Vp6L4EpQkoPAtFUuQplWye3F
2Xh+bKyCebMbUJYHrFqVMusH61iuiiddFu4Zd5zLjlK2vgYwf29R/57NRCBzWjAIcq2EYzaMSL5i
vDobyK5oeM2RIjZymiyKlIceqGEHLg7PPa2mQzQ2pN8qRTjErpegOxfs5a7Srrct6Ig3N1eNgm2C
66rulD1cq+qkQOsayHQ63SnDcXs+Wpn6Itq7VI26CFwt+lCiWGCv0G0M67DfC0Yvg49WZNuHxMje
9ykzuk5n4yH+8UVk9b+e/hMdbtm+MMp5CaQnjDP8BIWQECjRWHT/Z3R5XQsHHYH8ertD0djhLxfu
NtjDRdd5UOCNl3xvd1/i0/DcIzF2gZv5RsWSK813/PSBnzJFMZfLtJX7dIvMKBTmsqftBqyOcb9n
nLEdsVPUgFfiXQ0VZQSjzUJqfLvS8IAMihKj1NkD8wvL9QoIGgnECH0yBRaqYO523p1ipqY2+TiO
BwSq+2dwcqDhom3GinbsY5ZCI8Z6yHLbd2H6vftRMHQFY3ecZjKewCBt3lC0iVK9x2A+MbQw6b2I
vUcUbOng6S9Ve7UCmVMM13f8MUc25ybmBK+fG9CQ05cl6nERle2nJH8Vn/jp2Uq45LtXZv3TFY4c
K94IEauR8YdmseCFU+KMYzLbyVQr3/s8b8O0bmGJZhanHnn+uvQvxF/uA4TFVnpILM4cLDvGOOwL
cNXEdjj/0PHMBwbLOGrh6dzvOjnQd6d/eMQ6MP+Etid9zGctQY9k/UbNOx1MQt0q9tzFJpO8/6ZI
v+mXstPU7dNQjmWO488EKA3qzoy/qiSFzn4jlmnaPvk4mzv0jZfbeFV1w332VXYBk12aoYCD1Khe
dgnWeYURSHJaoNK5IA8F3AU5eB5eu7/TQ2r5BTyjysVAX6bAGdk8m6BQqQUSXTx/OejA4Cjo/6ji
/lxbLEM0SuKmdu53GKxdrgk8Nozdncx7Jr8x5Un5TIGX4PHqdUVch+bkC3xYZnhr4rejLtm3KNvp
YauL5svigA4c31gNo1o0+prxV0ML6euj89NrBn5Xv6yyGY1cuTERfdJjafZ9SCvLbBAlZyyqALt8
XeBX16Xx1G6mColzp6Ztiqefcuj0m7DTZXTZQPKJuvnSkF8f6u9fZJdiP2/GSorFC0eZHqtnMr84
uYVEFoSHIwvE7SHLNRwiixEOMFMuimlDxleWCClYtj86cGJPZFLVDjI9q7l/9qoMbeUiKIzrcRtJ
US0C4MTvGVOTGrPgyfnCUQVr+xnDfb/I60gsTyvvCWLR4gdQg98plFpTxhDiYer0rMITQxv5Yep/
1xMnobx1PhS0i6KQycLQZeiGBD/GdL0PlTWDde6ThKapwKUlxsWJC3CRM6VEtAHjbms9NKtywKQR
z8mtKWFPU5sXou9hlWKsUYhnbltbdbq3Nzacv0K8SyePnqyYP3NL3aQLTdd7s6IzKH4NyYmnG1gs
ilyktzO4I6UuGBRFa3ZNZS2yW7CCHTg9D5TXTLD719N0GzgztG+Z0jds5gL6dzqO0dQXt6ALqQX9
gsGhENC/kP/QHcXxOumCmZ1/FqQJ3qBybD2qkBiqceRNT2EWG0gBLyv7FQCcyuSlEOcVg7ON9GAm
aq2U8o/+kEco2+v5eBZTFOjcBkz11PTzC5qL19xn1zJL/UY6zyrVwNl/VCSjHIaAUthpAyIixBz1
HToc6fGjW4G/zLWf0r4NU4AcvG2alFKJixWeeG8aEgMKM2yFjSlp5KWTxCRr14NmQ8MvvxiEM3H8
4vderdizD92KAB9fjFpDaXgNpZGItE1Y7juLcS28ZnEbF7aaQWHhp5/PoCdbJ50Dxdq47AaHRCRL
0ux5bFVXElgz+qE9qeZosd7xAQjFQoyv5bvWWDRgCuKImXT/gUHEt7Tr5hTJY2xHhisV9tpdayxD
kGaXU8F66C5OjADwhv+UdDX8sbpXZleUb7u4JGD2JM8o7Vt9dMpZzep5t1njXYWYNYYbM3/2dGlk
IU0fyWyJKwRVHZ6GbMqhZVpLliFY8zYy68vJ5fTlJRur+UI6D5zp3rQb8T26Z5ouKCcE4jg5uI26
PAtN0oozfQq91YN+wZGKiXAWEHhkCm7sWeK6yBULMDf8sp9jZMHyW8O1d+GRyBni0Y/zj2o95Lkv
WVS1XDdK3EsVb1DYERsJNoPJIlFEA2uIJKW8Oi0GFV1PEnpeoO2p7Q+A2wLpcW2G3m/5mMIXr++q
F2fY1hIGLCNPeQ2kR1lz1DSh/iXBxi+QIBQl0fZt+YFR8xfVP73tVaUUvWG70w9mG+/kv0CO/zKX
QHAVSADk0XSHh+hDGMRW1B5DHheAm+9xqQWh2FeZ65IBN8Y2MhKoy04Hlk8v3qM/puxjJ9C/aBhq
lIYUVAFoVU8L3RawCH6NP5wY8YDFf6s/r9m/9seqL2OKzkl28gMscM5ho9t3d8vq4PxIXQfkiTXW
yq+DJ5OzoM7rgdKBqUBRyjk1WGl6EFGxvV6i5p4tpm5vCDzZNu4zKYXHXPU74YBqA0C0eXRK2idH
SYFhDss7SO9JWa30tQ/wqN4XhGTHSpb+rPRaLAapBJyuydcbPrFp5o+rGrUYCxjyRzB0HunbT2IH
3W02kIPozXo4rmmErxZBquvoODQDkXfDwOnM+PHl2bdzEOvAfbkn7dB2U4MVjnZuzhJb+ztJmdws
TDUTEhqA0lVHx7ZkhfD9SMr7XWZzEpBd1aavMW9AjL4E9e1d0R2ePMZsbQloob3O2q742771m8yE
1uA8J+sb1MXn+9q1vMeQUeCFiFZq/vkIyY7ehn8WN8KOr29dQSDT7O5iGHApf6dnRhmKESdyHher
7hVWi4Cbj6wEuyyEqXmbLV5JvDsE4gbGACfiFRGzWUGLO8zHOnVkpSbHKthjPWdemP/ex21hnER+
gsZyYqvOrChHVF3WElu1nOGMHRJOUmRVHxSUAoNY7JZi7UwN3cZRZqOYK7jEoCjqJoGKNrvbbA7O
uq/RQRBd5iraGI82EmIdJpauPkOsCiue/qeU5b26YeJx7gfoDOwe/JbyrCS+qGYkXpgIq/yahWVJ
QuozkvwmmMmezPwaiHgq5IMVoQnmM/Uq2yP9hkrz463nSnHfemoGeJQyWbKv2oX/BSTVYPfg3Y99
IqXF0nmGq7qj9MuQeoGdmkdix5kEv+zKNa8SBhMFJ91Y/UmdBUf9tanHn64D2JIFkqTY1MtXvfx9
xt/kwFp32R9Tru+TDt38jnCwQxD3SvNBMhEPTBDBHv9qiJs2/3cpJkOwIWHckHJSFHlIAej44k6U
OzISzWKor8LDmGn6NfvAg5W34aM/Tge4lh9Mojuh2h9xzWfiWQKL2u/T3DCR+VlLGmKBizYQnnKH
LOMj9egy3uRf2G5qXA4m8nbc74Pd8ARFeuAvb707ua67ogqVYG/O2f/ijpQjIekmU3SiGtB65NJx
T0r+m9fmPO7WkiGhd6iVa4Hd1KMUShdN8XoP4cgBIWTRxZiCOp4wLZIZKXxbPpssK0poYLCVdofh
C2USpUaUh2HkuZ+SpMTbuQFabS6Mc00hxw6pl4HZZ5MqIqyA5WoiwuYce44bCjX/SihfFuxJTOry
kCPbBo2LNNeG/7i4G4tQfCBnSlqU8gjWIDMZttkP649ybDu0eHqg/Zv7zFW0En8HmldA3xumKUn/
jvgMdq7bJQ9M6nrxUhXPyKcDgM05YGa2atIG1/CShvMJGicdI4s5S+PTryo9RK11IalaPgDdgYI4
Z3E1KW4V8MEE+DSZxL2WLicr/6uc3qBlwCoBejOFqGWIr1kX0Wd9Kfg6i/J5dxrluDa+W+hyRRJa
x9WowqpS3T0cQwoMd4ok4hzihxTf/9WMZ3r+FKDRfr8j1RIAhyFJMIdBSEj8hm3NcOR9BFoerA8M
qdGDAp52hjZBRzjEUjOwvLdSs0YIy2whKIs0vbLX7IvG0QNoNl6FGEebBzTlb/aadwWl84N2DkF0
VCC5JEqCmvoOQcXD1IbflPZswNMJY0zEIrm5L5VyG2jnHzLnB1Bg3K02EW6csHZabNqCks5esTG1
qnyGgz0CPCbxoOiwEOu25oIbrO8Evxhvf1roNnLnCsFoviJjJKOdfnGHabLyFifmiH9iZyGf2lcB
a6HLgPRmrEZkG2r0+11l65uNCQgEvpulg6wgsbeZUvnmi/xXkwNIpKskNy4+OAzDD4/bYu9nvHzr
FeTBscDKTWSne4VdDBsZc1O3i+jJbiTxgMAEWsYBCSeThFyQRXJhhTzNJ7AK68q+IsrlKmJMJraR
r6vw5573gRhD8/Kxm6TK5hzK2IMJYICF7UAmkZ1V9aWLhzIowjQ92/vZKC5eINtmRps4a+7mDo1d
Z/ZyMUShuBOV+HqY4MEkBSQO5gya18CANzy1Hon87scsqB0ezLLyA8kEylvOT0uruzzlHeAT1sYq
0sOOJzaaIqv5bajAz3qCzHo20bAzUMmizuWStQfDdMGVv7OjhTcllzPkY4uSKZE0Hrm1VIO0RlMY
7AdeS6DKlAvF6Ld1RUYoiVXoAJnIdHuuRb6SqwYXCbAa9Jj4BN/Jb0HgGDpYiqRMo0P9Xsb4E2Is
oeU2gTHyAH7mINnzNp+2F2CGuUp5m1986ZW0P4xNVWuTTyZRyMDh4Hw72wXpSTD49VrzRW/4bYwD
I9edHSy9zuA68u2aBFm7RWMpZOgE7H8BMvr5g/zesQV+8VfQ78kyhiyaytKom/yOe2GoQqxmd9XK
3Y+HToy4xaKgJ0rbnLNtggycFyTe/XmOEz81tMN+vLNwOFwULx99fKvZwo3DOlRCZzdlgiPqBPof
MvzRpNuZ0BBSzRTiQbhd3mF2KrGH2aUUQosmYNSVanbcO0N1GQ6WRw105p/HQcegkMgsub2MwYUx
oS29/Nyq3A3H706IZDGaY8r/vWm4yHzhEicGUkK6SkxPwM5lZOPvuxjoXn4vH7NzA5jVATiMBl6l
EkuZyP3ZRK+GeUxx7PFlOEnre3OfDDTdetJHd/5s/BzFrd/kQn5ZvAKaQQxCEoTkCnS1KVOd1KjY
xbUybzubx+1z8hn9bg6aFNnTf1nv48yFWU/i7h3pGNk7vyEjNwnUZ2ZG98hMXWSnIHDZn8NKih6g
FtLqz8lWYeg/Y7h1IzS/LvUhRvNrzY0vfOIplh8vUKDKTNZ1AgFEO4dvHasUVrawJUNrWaWtCsAY
MBJ+nxReg81lXxBkJjYe+wY0jS9lVM/+Bp3S1+e1k0RiwusEEUEfikbKlpXcemGBnoFq0TIWOLW0
rnS/cY/T1allIFUAMfcUcc23PJl6V2SRScB+BGsD+1s9lbLBKqokwSj3oNkSK95khsRgWJlMgNZL
zVG27RiIyWe9TNTMIQZE7H4YX/ZV269h6Z9/tQQX7TkfQX8Q5e6aJuopxv2/eoC0owcDZ/oBeM9q
V1RsOIm8DA0DdUIMas2Dr8towCAzLB0jlwmiLTQCjV0RYXkVypSq5dM/5RRvhvJa2Es8YIjvcvSo
sb11A/YgzkeZ3dUsdIjslZLhTFCYUAVvqDa0LDM21/g35C3WL+LeS4nkq+aHS2Fr1TIPCtFK6JEE
IglbRGVAZkL6XfUKyEa9C0s6B80G0/WCnp/QTDrOFIHvW5jVD/blJl8eI/Pn3/KLK3nmczrzFLIc
Po1q2wG3wzhR4nNyp8umK4KQXAlyZYMQmmISChHGwYLjCfiqKvWGkg0B4b5V7jTdrt6UDYb6p1ga
09BC9kHziLc0xphI8s+AusHqd+bVb4f1y9HssBXNGEQdxgijaFy1BoadpH64VnDgCjqd9jIHWfHA
yb2wZutwu/QMBgACNxBLumXueP708xD+2CP/iK2WB0P73Cu3PGAXIzjMvH2LjjPUY7BAPPldokse
yHxPc2ZCJGRGbbFdmZ1It/BAWW1kgwTjn9F099HIGO48rx3izqIk2EZIDFywWIu/aW8YPaOZVH2w
aF150sk7hDMPDbb+vZPTfahmvFXtFb/HI9dfNpOmBJQTh+AAUbChh7HErxdgm+9vRwUJFV5+Tzaf
sDpVQ7ssNPYtyeqYahivrPYvdeGK2uL9S2BqTjcClZxK4U2MiARz27Fg/vDSn+etgTxoF9CpFWRH
Ynw8lqaCtaIugdxQRbPyZVW6MPuZ3y2s4o+YV8wi2Vn1ayYjT4OaTSyVfVaKQucb0rHxNBP4N9PI
lJ96t86Hed/JWMHrd6Q55LmioLnXv2ThePG97xrrQI/HBwRxMx/AqwpFnpbKk1JtSENVdiI9miHN
rLZWsmJ1uvhqy27EMDp4hpjqyqnAHAkBazeOZMg2Rxpu0tCNvX3Q8EhBCXDrwX1haKPuNaFYN38r
OWHved0QGM5NAVPTR8UlvL5N5QsZnkIdpPveMopdPAapEmA4sLDCOf7Un6D8sjmPjtnEs43JqtaJ
lSZSCykNzVjFctiSoeWutoUmSbMYdGe8x9pT76wfHMR1ifwpEy+yH4VDFCIXcn/7FJA70YTXraAL
EPm8/podMlc3srLl3iPsLj+T8TVbkogdif8L0nspgnhFfm9oz4xYxxAZ+1pQR84Qg7Nzf4vKBggJ
Cwjq2ryz1Y5MX6UFIRQj1WWKdlOkCSDmwGjj9mhYO5dRn3k21sCxCOsA027X2XDg7h/z59UBBtk0
ka5C11yLOjflZRFy4c2NCvW6sU5kNzPzdDmilLHo8kPo5+MKaaSj5s3P9R46q6zrW5AAuV9BI8K9
CHW+S2Fpst1vLdI7PYr/3LMHlWq+bXJos0XYwPsN5q+51IH1f45x3hw1+YkkjkIYqev5QyroxQXX
mEaNNQYwzny95K0fbS7SVqO0gITX0UMJ0rUTvyOF00WmI6u9dtZ0a+D8jHStI8YGu2JjqOVmVbMa
Ze0GwEkY47L/WYwQ2r+SVrmNTW6KaY05usEnMSxx8tJTUK8C1DLvbv7IxtCPo7ofY9/tGyxPOHpy
TH/T4AtfzTVcJBLFaO4MshXh05VrOEZRZXAUTEpHfo7Oh15BDPADsFmt3uRMrsIRXs51kt2E7lbc
TAaLzBCSGdWXmPHu7DmHHzZJ9wOIMFOqxgPLVSOJv9YpgbEYmvlHRaLwYokCJCcSF7yvcmT7Tf60
64zQSUCecU+BI4F69uBpThozWVY7qf8vlek7qGP/W2jvdIg8WrThKnzzGX5nJ+4M7vTCp4KUmhRx
zvduIRggKwH68JwHq68NpIMyxUlCNF/5MeisGKtYXE4K21v50Deq/ARNgzb9Z109Bc33PSLlMthD
HQBEi6R0qi0AKyQ2jreRe4qzR+ER2Vjl1g46TUJ+4V0Ebk4LKPYsRkXhlM/7GrNgjz+Dt4GB1aTv
9N63LLJqW7WgEr+bObOt8RwjoBrUjyv44BVb5Kd4J1duoUfPTsQWZ47o5XD0L+ZNy8MBNCSESNBR
nWsWWVrCTPqK5+PPuFRceSKZjOJvrJHIKb8bGn9NK3M1rRIrsuvclx72NdvIBd2+GFF0HUYCgsbH
+yMNJuZMXXGSPJJWZ5sH5iPGDSeFO0q3lcyOINhbK2KJuugo+DCNSKzx5Lh6q3EuMRrBx5ghrhLS
K8PFk285qe7zDAvqv+hduSR19lFLetdcWbZKZ/dqdrCDEDxbB0sqcr29Eo6bzW6o2RGvrWd42H9S
uQzkb9Hn2ZdMfI6NINyalD5wDlAPy4FyPY6OZf6N7RtrQ8GS8p9oBSrUmhdPk8Lhu/78ZicBgVdk
r0QyjWlZK2B65yxVKGZKque6rgzg3EOJGB7k8hrFRbhc/z1JCPS1SllzHGVzqPmJuM1di5r8oI5j
tZ4dnjmmcxNHlOtqIiPWnn/yMUQVgr0jSitT49pyeC5y+yu35o/p9xaR2qs4+8HP8HIvwN1emxXt
94efPJK3xpTBF/GR7JCJQJPLj3P8SlD9dZu1lwgQ+IfPWQlIt0wEierNXvyNQeT+JjpKZjEccK0X
wdxyW+VuVHGquZ+/uxwrAcEWAilN520Rni9ErNQr1nQZaeobrhC/e4pSyNRYzJ2E/gqkSNUuqmDS
Kfq6PUU07V4tjxgUy80YbqhncYp5CQJou6P20aB+LuWYIpLtUPs/iubl4bg7hUB66s922SmPuAXJ
1jECx/GfvdMlIm4+geq+NoDGNKbY6d6Dup5Vozk4SXOj1Wnk0xrpCgluWxlxEmRMs/CiVPvZgwhH
ngiCKOeDqfp1FwQufEndF+USuIhTy9kWRIpNQ0SerwgJ4XKnMuqhSRVIZ85qhAsNsA5TClN118qh
+yzcKkJbyJpL5vp5vmZXL9JsoKIJoIQiJj3oQJLmwTsIKcL20st3gwLas9HNloEt4tyOiKWwyTzx
u0eDreOJm4UdmLImlnrxpYemsYpROPbsMTLQVBOegUPopF70LAgdZfYudbyaWZmDxXoPOC+MuzJK
QDBJI/X8TFDXUZlowQYcg7dFYXfejGSkfVKQQWLsvsXXvpJsnREzJC521W2tTuTG7JXS5QhDYrWB
5FfOvVjOrd80ElRaAjQo8qYKbgE9d0tut1Me3TvEvpGuqy4It8LhEhBVZYQFl9G/FWEiS/8FfqOs
cPbCKaNDCyw1TucKF2Kyni9yR9opBXAw1k+56uQUKyc+Lzp02SBivJoSLc8kd1VdPHpoB285ikAk
Ynq2CdxtFU+tIN0I14jRP1aJn3yDxTesGOlqAmnXQ/LmLfVHcoMvwbaJEWoEJ1aqLnCTr6nYUxZ+
FGkWw1DDAMuJmR2jHLbJVfcMcyh5oQcaUWRL5Z6vtPcZxOlM83aE/+Nh72d6jq7dUS/yEmLFWAU2
LrnOAbUUxUGKQth90k1eaAuP5gUDDGONgoGFdtVXr+nHldDUOx4lzHXbqi4SFr795Ih/yGL65EdY
Cg51IazCn0sjB2RpkBQUCXvedqSbcUXhbay1Vvz19wnWuYUIntDG/LhJAAo+1g2lJ9JEJm/132gt
+2+7rCh4UkqWFtUee8jYBm0B6RThj7WgoYKi9djJS5Dy1GAUPGNwO5/5TzhHwIDgNEJ1gjqMxS8E
EerE054X1U7pPKiDWv9mojlA7MlGnK24UiXu6XEWF0Ibwmq2uhamR7q/2eYDbvvvYlhcWfNBxJeS
K3chu1VlKONAsbzXQK6rCX5Aj1AuZRMygWIb9smgsnSJeQNEfsuH1ZfzrcMv4Xd3kwyXopylBXZt
k0XptyUOFAhS0XIGWBd5d06fjKxwSxmfQtYmZZF0Wo6HoofYBBl7KZW3t4QY6W5DDxskFqkqDC4k
cjglqdb/yjF0KGA98ywiQXZAB9uoVAceIY1FGtZUjDRGzM5VAy0k3MwWXDMXIGrBaEVHjgR4M6WS
iOxmdlt1p02la8cKFzDEdz6SwAekfPO7VV4BhqGdaeACEK0ke5H+ZuTuJFwJs+f/LQZlaAJ/dTMu
GJJQ8CaUUuh9FxqqNdOwuhN7V5HzMdPB+ykASS35KCmVBWrvsAVPbBcUx71N1SnvcA5SO/bZMaTR
ZK+aBV6/OTCi1Uk04Q6DnOrVwxN3KsEg9xDMP9PzYTXybgitw9YdG8clm3sevdzCqUsZczgAaFPt
PJMkWt75pNz/Ijwws57oHncau4Eor5rFU5dB6ICho5Qv0ONHTrVUGwjZ3OTYPQmdHF5DId9u0Ktn
LwzvoR5YYNf5FmQLu7PtaPqACr4s2CVTTfW9WWUAFlZ9p68CWCh8wHlCTYIStNRwnyIdKsr7VBaJ
U2JFBRCzhO/4AxtdnLdL1L8G4vOXT3Xpmux9kf2OO+uOYLrI7YK0Tc8quuSzlgVYGAOrdLl9BXl+
VbOpBCYMOUKxPKB+k18A1lVV8d1wuyyCOBHcIYEpnbvUoIr6VcJv3+pOGQnS7SBRXSro63LZreIz
QJ9PXE9oiQRgE/f3FgQtrBHQpYzshpYhjsrMTEdH65SkAyUlnlFgazzDQbBBe7pxMA0Vaxw6biNt
Tg9tvXo6fbW9ORM9J977SO9YLRcW9Or+Nm1Hg5tJw0nP7vMF+iunscGfeyLoEiWoDh9HqbpG9dkb
5y/phhAPvlcEzheqT3Z1nu94dzZ/OjC32px+/dP8Gphgay58CfazQvUTDPTAFmBTWddj6AdEB9oV
OEVZaLQFAKu6ZSmowEZJs/3AP9Ny8NldSgGLeWtQar/1DpK2PfRQ+bu3z0Ik95Ztc0Lqb+/Bp1uY
kBLKne2wLvTRoM4QO4OdTGgYGBD+J1xHf5nUCKVFGcpG+yKAxR/RQLykEbdSqyX9OeNrFqVD8ROH
uSQi8XIyfY4h5KIaYPLs5+4FraHg+jFZHO8jDXaN01XbyaamtdZ+1bU3/1gtrtUZfxK3h9hWcrEH
5w4jTjRd8plLptd/zZLmk2CLidvPWm+Lah1CpXptNvBATeaPc+rI69xEiTO9mm2jIabf2Ibkww3f
gTd01W/4CwBD05aMpq/8fxLnGil2V+YnV7vWtKh261ddAwzS0pOBs7JXAYrwwv/BqKQLc97t7yhz
7fJQ2a5p9hjUGe+cug8KS6a1q7d4bSdNbr32ho8iVtWirhCvQoCs62eBjgFwQf9d/gQQwnDGrk7E
yRKnsoO+j0OiBCb9KCd8r/tmUhnhqjVAGAQkzNsl5QPb1ot/LgeOpRIKh5w7iAcFOVcPGohhkKZt
F/4PYjm8o+iwyWlC4pxGylVTdhtLNKrrVM44wkSDR52zxnD+GZnXmmLYFvJHuzyu212b80xPRpZ3
IhNb67miyxpmHnTT8+EarF4a4kEuvN96iIeMoeAgWrrKn/i6EM74yJf8cR6AbfF2Cx5aNvkCZhOS
msu3x7JzgpimLI5TdabSLUwd7Ta/QRG7t+SEWGZkXQgV45SzuXy0gBbXq5u/5SjTJ3PnVutdiFa4
ZjbFYCMcpLe/rNzFIU0chwIWM+U32kc0QLPiGXdpMJ97iAAKWourn7WkLHUD4QVTx4/Nw3SA3rDw
Ohs5VZXXQ8QiAZuMIIJ/I7qtIt2/ga0YkIt3/pnhuePNiX6mpoj7iLLBQ8CfYJOls2Z0FZhIAEOz
c8CKS4/YDVUI8IMP2upzE8xqQ+NAMOjsUXH5Yd8blO8z7OU/S4Q2G/pzT2PP/e5IQZJjmFfE3uhZ
A13dW9my3bYYh9T6JZL+Qdgirq3ZS+I1tILahlXyQZ3SVFOagrrxxefZ7KAdCTemKCU+1gwZ982y
Zmqtc08nXdt6m4CarOKLlxmt1s7007t3w3XvrR01tAVsyPYps85FhqBjFQaZj1tw8F6eAtcQzj+y
dB2koX1LRoFIEb8dzfHL8d62I5Y1Cd2P3iIqOQaTJW8thF1YrgixrTex3vgza69Mp+RCigb5Q0bD
xfiedRN/t9+9FJwyjEFO1c4iCyLDwRY9fm/787u1Fp4q/mzoxRdOX+tHKYmDbqQj+i9PlUT10Dbj
ohrNtCwLrTwbHTLtRk3jX9+z75+KVWfa740W3i9xrcPrxrrtl92lOGkHpqfM2j+VRAzVbqwT87mf
2isGX4n3p7UVJ3DeLnVaRdtIYjBzCKbHWldZKBOrHksi5o50sapHq9kc+AtzOMFumdlCgewxfnTa
iylE6Dvk/2kCRNhVD71Sd+vorVdll7S1t4sWT13gVAaeqycEq0bGQs9gqGnTCOHDWuXUBhIx2wiO
oXtPzWo4r1IgIokS/MEyWdLWvVWrlKFfBpy4PcaeNNA8rLar0Fco7HDEXiDf3zOze0f7uDvPheAk
EiboYjQHwz5XERkyMbHEG40BTJoykrb9Hf2OoSdgvYXGtHMXGHABQA7rbmH5x6rP0YEuyfEV2lhU
4ElAckmIb5yOSyJyS/y0YsGWvbPCnVHzfPGWqem+6lhmXEIY/bcdy5LICca6Hg/oVW8aHL4jwqGV
5aIfN1M43csSTQrejzcYivdHd847TZtv+RP/F02VkYw6vylrbeoJ447tmZYxCP/+LK05uDLJ46ci
9ATdV6Ji0kq6FHgN5NO4ertfxz6dM1enh5+72M56rtSfI7O91yZrAl0hPCgePWQ5peplrbvVb81c
Udr49OHulda50pW3b8TeKREa6kIb+Jea+kGE5ZsduiR+I16BxqLvriQ3DeyDntABsb4lpwUbOzgo
hKykrCLSKt0PcyBDIhLMc9o61Gg/zQ9GL0aQT9Onll/i5jqfES9F7BHXdgXlB9RUntA7ZdhGMhrM
0UNgdR1GrM+9/8jMuT5JyI6nn1X+xQnuaEe0lc9HILUgFNTpSH7Djg3BC/JspUOniUXOw0gXvE8/
kjDRBYsQ4Rotn9anxPfqrGeNDklz8zV8EexR9LkAfUm1WC5q2yVKdhRqvVS9oaYsgBotapuac4F+
a7r908cCovNXRoSobkz6zaJSxW9Ycgda7BGQAP1aYXdo6UDXsb40W4tanmad6EioQWEjFdbe7k7q
ajIKUj58Wr3QrYvN4Y1Amc8ahyrwClKYHhaFRJ2PQkidHcS1gVbfqfak+2GmWpgt+PqdG8h+GV2K
N99E6Bhf8SH92ORCH5PLoAUds3dlheU3HKzQSGIhkzp065JED3q9t3sisvEIzc7qCj+B90rLm3Es
5zk+Ha8XFtoPic71uPiOEEt/nOe7+tNUfnYUjcbtoPkheGbnV1Tn7y6k+dqKnvBnJqvbYULMQfQG
7KMZhMDtDG+kBSuik3RwFj7lS3+zzdQ5fblu5iM64NSBrxwlHUXZ4jGhhMPX1scyNirAZ4DhddVK
U+eOUdTaqMyppbXx0mXTmooRfHkiwxgEmtW14WhLyKPjtbbaEi57bUUEP5ogyZtGLJdlnH9hgLf6
XSqlTQH/c9873Vy69UcXMrxaKBpd3Pm5RBM0MOOFPOOOZ4SfxK/hwbZVhHNwXnUnL+lmO1tjC5hb
p36+1gRtxNNGexjZjiOZUFchoFRNCjowv1iXGIohhdqCksga+4+h1XbE3TveBgdB90WTtLFTVTeV
6JyfcsowLjnFrRoQEw7FmbkwzC3OpxbvVTSg/iWTR7HEKEtp3ZtlMiaqQO2HQgAe3d938x9z8nSH
AWH6K0NX2uayhc6e0OvThRi6/T6qmwrORNqep36hWz1mY/VY4qE2PCopjkK+v3YIqAshDDmdYE5J
nHOhkxeejTGmHXIHji6cNYSnGmqxCgXU6Ur3FJfdTVywGPWsd/hdsdQiUfGoPbJS+ozgq2klaXqH
uvXYPS/uihs33C1xzGCoLu1h8RI5UB5zGZH0XC105Fan+LqPww3YMQO3DuzxD5CK/JZ7veUgWaha
KfBh6VT9ipoT3UvOwRZu7Q7sn3UeDlEVsNdbg8BBfNaUhF3xKuM3Zsnk4LEk+wf5jweIihplMPmv
GKZZyyGZ695LD3IK2QsoxXjzetu9Ah0WsJdgEoyD8njNEQWIiDOfhQNLVlFdyH9fZ1IsbqwYg67O
1xdlIKRSPv2nFr4v0OM6U+7M3u1Dp8A2wdkUoHeUjjnyWP1AOkItRigr1H87JX6Do6WXCPyg9wYp
Zc8CZmr+4cwhhcIolaARKWRwG1xuHUsO9swCD+2ODGAB9xv+6DZ0y1Kd4UtPef7kwjPBcEDehvQY
UuTw4Ww6C+El8xohJL9R7MChPbTHAYv+u5daUITIKDvfqzPQMb7q4GToK2IQkX+9DQkoRwjehn/5
2+G6Fu4PMCc1Y5EDRlyMJFOdeI+f/d/9z6iqunHLdb+N6gqLVtr91R6ItYrCG//zMXKI3JYm+W4k
07Y0kvUnNd8AGWYVHJDcmic74Jt/WY+pBoYF6qsZ5OecjMpdqf+tLJthEyPXEBzxE5XSMxQdKMbq
tH5nvabmUcFtS6uled2Eaf5mXcbGUO7iWDx4HAfs2c/snHTMB83tKlAawcgennwVjhty5zsC0I+J
iSfX3cmBzmZtl/Ph31L5rzGvfxgxCyUbTKt1Xh/CnMLzShkVv5lg+wlDZGozQNreDYQWw3RZNVHW
mg1vcjbooN4G+yDOFqn+1xLZNX21TofEEJFBE6ofsclyHop44lHTj2IA2IxtVZUmIcu61xXpqjGR
9fcCV+deXWRmH+7l/QYsOqYdmTLlw1f+0AMhi47176gD3N5NWFTmxQOLfgmsBmNFEuCqooFzQaHY
K3jE8Awx1cUPz58CzVx1PDat6UEcI3AZw9PpDqlmTNXo1fD4LQ5tYWJcWDhSffbMdjcOxgelIdCV
AURDWb88wZ/BYmYyhL+I4+Lb19lcV62sC8UE/8oUlBvZxJIhMH6J+bVQqd7dDZez/HyvjaGLgh+5
hdfzxQIrYnutvpj1SraFUcnqTLKIVnPLobqFkiwbyT19I7sD4cUcc2uCDop9k7CSfmO3EzWL/wCh
l3K/5MQdrStnPpb2nnJdB5nfITqb6wkC37D3Bouc30/fiLAvN7yExdVMJ85vLFISsjIFI5zn9r3T
EQ0p0OdzPEir4ZDiYX6qPpkhEFmgDZVeMF4jqDvvkPjmgjQTkcscotzhkuYPX93SWVKEbQkTPiOF
OOeTXBuv+yOVQKVJc0y+qzLQxXj+hxHxPIhUWeChrI2IAyVM59CdnNgnKJUODHoxYMjmJlv3VVVI
YnScP+eHumto6X9GCH5iXn/XMNpQSLPxxFq4U9gXUuadqG/nWQMzMS8p4+4Woaa9EvAEjrwcQBIm
gQXl4HYBMRdacshE0/3Do+j41Leu35q51lj0gyrzZptpAHo7CC7dbALdTE9PRpZ0HUEaMosyoqcT
Wq1h9XbTHsdzZDTRUDcneOuoiaqth0EZgsW3E0iF+yW0ubpWkTIGeiXIygbqbwqdYOp1elMzlwXN
BfIhcxiJXhUfsxZeh3nXe9lCPuaDfDQqZRDNDVnRNWOs23UASQgZawWtyMc7uR6SQBE2jwiZeLi3
HQ9w+5hxLsheTikBzh12Mj5K7cPbOIp6dTKnDl0IQ4+yOxtk0zkCBzSCMOcWeLyglTnnfib0L5Kw
ixuQi17yxc7YhMZQVeiMWGUrfdV5e/VVJbg+MgtTmJXt5Z29RALaUQxrjOilF/4hz1Y2M4uv4/DK
rpAB5yIBQW9Xap62YQisQ1gbPfIQOx84RpxwaDztBvW4OFEMlEOahAcGtQs5acKe8L4RBr7gOijK
G4joptMWRNs6Hv8GcCt8ONWQkXfsoJ6JctdjoICzB5tdhUt9v9EfqaYhqMMKfun3OMvdwFq7ZbpX
lMpVZUfO9/pO1AdCv8QgEnNpi7YSgrO08EKjpsGMZDsggDfiHi/XYGTbT4bNkR1m1hETifr7k1ko
jNGoRrQ9FfbUB1mUWGLCfoBHk/vHtlN3eEizTTV3Ezsgi5nk9KSgXvUmOPFxWwqnbhkGBw37UAf3
tVplm883SF2tiqTO3L4z6qTb0/bqvzSInGYgiR4+oqJt3a2Vzp9OXL9tQ8mOMU17toex09S0/BrV
sSbRafymxRVi65Q8wN3VkbdxR1yZkiyBVSXyT9vTmI3NqaViSQZWoiYHj4ZrsH+eOzxHsgNHWNQb
6X6yMT9FJJO5s2P+7WiW9VoB7Yt+vHcD/cv/L0yT9Flz26v2G+HbYoOXb1mDKdzkT1Kk4n1v7KCh
BgUwgMQaDRMIuSr7EtRIw7OU8/a5En6WeqQvQwFDoDWZNe7UA2Rxr04NiiSvlGL6sy7jQdgYdZiO
xZXF8qSflk8SU3mhtXjhdw/oonjfW0AIMTSp5JepVdS80CuNQsPuwLXTC27OOrkNHivhn1tXCurp
cz6mIRJLDN0JBMioW7FEWI/tdHoB2wPe80wDGzTPJmiPkKqwzEwjseBosgMowy1613cHf4Z10AtM
Py3oyfvCqOfaDm6+Ot3VCMGSHPLeJY4hQsmZhL430tUNWLf7zyR5Q+aWkTQrbZfKXYShU7cHYRta
7JbohbyVaGpGnpptb6SZQhex1qoHiCuskyYEmzGdoLEVr6bcryH8pRL8INT07K3xKOVqSX0TZiA7
zCZMNZmS7PCPyyxeg6lmisERuxJwh3qbCAQTyFOSf9A2jILrOgHr0AWHymXXoauRZOUhzCZKjI7w
gHKFkgF83v8P/FP7jyNjRytVmqXBUNnQNH56+Iuqszl7+/9zknXMLNUYOawowAHX3MaYSQdxK+73
x1t7K/pXqBesuyGQdtAo9Bl+ujZdY9yZcBmEwg7umcRV3mKa8mjbfXAT2tdVs+3GqSiAVbTuRs11
5PRvhpbOBNrfPSJFgmp+2p/EJFsyM0tz1fpm3doIcVX+CFeWJ6QrMDQ8D1+QbLefgU1W8Bi5fyNk
rKZ9AYCmXdRGFBHv3WtAk5uqnNGeEPJnjHLLu/2Q7DeVSnQFF0d9NBBgSaxFxd/pixwpNMFtwAsC
ZLhMwZFacdUpolaZT6sC1B+yh4/rpvGjH1rS3vvePwKpzga6PB4c7J/HDBRUDuY5am9ifCRe7kx5
0Rik0sLgLJ+bla7F6Wkmkuv4t0K0ArCqB7PBIxYU95CRwuqCfE6g96tlt11qMT/ggwlsBqqbfvmM
GPv9KyoShCfotCbqJ2kKiR8fHFZ19VOcSgMhZmGfVslRCNUACckzakL4X5Cynysuuft25MJvFNol
xAtU96ns05s6ZcXwYJUJdDm1zbCWO0BmngWadU3sx2ZfALCqirBRtjBrmTK6zeGYiqd/PY1JK0xk
LcXV0Sg9NL8tm+VZ+koVVYmSXPECU0AEg8VPzRDgnzMDt38Ssz5ZlP9mha3/pj5kT5dqAcJ/RTmp
uSvDDUyqww8aA5iXRI696ccwhXOSN5kaYAI74Yn2HvJDMsgyS3jt2+lclAYKuQpRZcjloy8KbrHV
p7FpIJ3NGJWiMhXEKYVtyNNQZoRbdfaF1ky01mXxu7h+uaec0YTBD7C0/wtkMToMhSxvsBF6q1mY
vcnll093lWiP+76vi2cRIk28foNjkw2r1RkPaQ33ANCeUiZGmvpbrIDgQyJjUZMzpirdk6OTMLtT
YkN9LC9gZPtnCj2CjTdfDWAPNNTI6WLHL3rPh7BB+rcMPQgfeArFcobvKLV1JS1nBO3kiG3wGsfs
ufAfc8WHR7kLDQ6deGQeeM5/Qgeo1Lf/gJHB+ZkAUTGGwwYwYGovOsbdA72R7NXViuh+UhixFwIU
Vj98+/qUhgFuVgTcRNWVjZFnBzmwwezdlb8K82MJC6dav+nhNZe3c3bVM3Cc767bGzC5tC/ue9Ze
yxcVSyHQP5mI4L/5r79TDMi53Pz3ZMN6uhgGoMDfXiywrd5YF8UjKu7+aY2hsZO+RrrjIzSCwr9y
ih0y0/c/AnYM810OmXrslAwLgkm3Y8iCuW5+su8j7//fh0OyuWJkFaRMrNjN62PYHNe/t7h6Tzni
lA3M6XAQSljNK1BuP3n4tm5X/wXIjogR+rQ9F4k1KWpe61agcBnJe7x2PaX8F1jn4JwsrkgCvgoY
B9vo6tU9LfPLH5hLPGhxaXoFC5IvkPYcXoFD3B47ycEv4e9Vkfabr1FUgL/jT6WA2FBJH7g8CxyJ
B2ZkQsrHXmlsGSywk3qH0ITZvRxyxqBVi4Wtkdps1tG/dXIUoH28TNY5p5WEnBSayO8JM9C7Px+j
cb1KiBOrcVOwjyUnckKWxpMmIh9uzeA43XrbUiTUikhLZw3jk4XERFWMJJVAAqWxVypdHfg0m4O1
7RtxpqU3QNusizhuBJ0ILHsywSsj+6c5wmzazCKmhQYI/x8RLgbyCKuHeCwHMeND/OoE6XxKa7gr
1z5yr3VJKJekiGOrzQv7aBEYEmneCixCmwKeR/VY0u+dpIbXWakmPK7LtwIO6XRvYGDVL+mpIu1j
IYMhVVRJpaSKjcTCDZmu2QihScHPp0sjE0n3Gh0rwNoyawQmNxSeGjg1ecuwhaQU6GQ3XUYZOpcy
EgkTsl6t6sIxx5DBlT/jA+z/DOvQqMU5Z+1i5zdEzvrV/JwsxuUlUBgxFvGGlgU4aLqAjOdzqun/
xPzFUwNlrKaarzSeoVA/JqaE/lRzNoLEUibKhWGJrHJt+sAAkW6VfLv2NCesHzuCYBhUrojZykbH
kVCxy0NOR/uTw9wga7RiOcqeXWD9chBqHVyPkoCXP3GVoZaVG7tjDO81yNDTlVqOA/6gnWt2ZVSd
seGf8E6nLPJPNaFRF3hv2ISbZgH0FrkQJW8FbdZALP/EDI0BVnpWoXCyLkfRb/KoY4C5EoOisseb
sddbSrRxHNSl45Zwit8rDu4hejeDSsJ5Q/zx9FLqMKmgfQBxurqy3xqduS9dBkN0rTkEY2K3oR/M
qw9IMU7EpVyMKjzvvsgn0JqkErLIhUYaUlo6V8TRgVNHs2wcv6MRiNd23bducS7il1829/gVg7BO
XCoTk4BbjpS0YfR5gMOWaTM1PrOIPgEMpoDftuVn7tryUPlfzqI+3IL0OybSBmENVBnkZR7Fm95K
9dN0hizia8Kfkq2f6LHMa4hRtbvY1GViBle8ZqMf3wMyoOwoW4WWijeDJU/6pOFb3l3ThBlEMDAi
I+R9rNOW2JnCV5YNdXv0gs7fmikSMoR+4m5+T2lKQWEdNfIBClXVGtlYU+DyKkFocoVJXlYhUR5d
kcCAqdKby2WnjFIWZQYiK9rTxdcJLhQ0SgzKOLc2OAuvwqXT9crEJekaVr06cOC7hn+7lMb1h8+z
F5ExfEClID/V+uYLgq2DTiOGiajZg65JkSUYMa1r5wYhi7ZckWxidu0tHwXjB+wo75wAbnRaESem
GRbUYdokap4Z9ctGopSg5RlBOiy1WSTX7dbNGB/R/BpwbNe+M4KFTpuc7Wb++FNbcHhlIEG0edJe
sSkWZH4FKNVnltxDVcX4buje3esjdXy57aQvSRaFXDVNZgDd3CK9LfFHeuoxDX10xYARJvPjbhWs
AkZKZu4Ldf0ooZZ4IwFL9XD/N5/fhxSiH7hYKoOYyU1z1dtedsNQ7TjLabhq8ITYPIJ/MeajNSh3
sV3vbxYJPWn21nmNo0cmDowJrY1UiEO649ZCPdlsC0opu35vwGLkWPsBkssRSqBB6K0mSmGjN15b
dYvNK7I4s4zCIEeWf+zhod05iId0tmgY7SpILCAWWLI0/6rWVNPB4wLnbCKTGLwiTPEwwMjZ52ec
EOmN/T7QIGG4xiWWYm80eZ7sMAEayirhvoqUUGMCqW3gxufYWWlxG/zVAbmzwH3veVSpbe3GCI29
bQTTkKDAWzVQpTgiV3A3aBXuFVAtpMP7mWNo9bqJb16UBl8jEozQgp5jfRD4qqycmZ0BsjDj1XwX
kOxUjtXhE8YkgHV1Y7QmVYLkS3KfEzc0WmDLs0gMtVL4JL6mS5i8Ao2Ar5vIquZQB/OFoY4zZEcr
jG4L99QHe0fSoQKxAW+die/3tENgKAZy5oJ8+m4lKOB1YMq1tcqcyIFJY+Xi5vto5zKqL1MkR7Bh
OAt3pM43F9Y5af/MzuT6mLS1J1yGMjwHDRYXPEAO3qGKmBETKHsJ70go1zdRQ5diPN8UUS5pFf0Q
98rC8+askpBDBSGmIIONGBLFf2yRxFKoprReb/ixDzOT+Tz+DT9rLlJg+/lnNE9kH/qplXj8Yzhb
2siYDwmKM3aVuz2amhIH1hV8y3jPSClJnCDwAccyTU2DAenCMFIRVd4X1qyHIOoN3koeZpDDUMhW
QzsI6pTXVgpYyrlPpndhYMPQ6VKLKiEUlHmEk2EWszYXoo+YfSDMhFWSl4A5hwauWY/949IlWI/e
pxR7CRMGqSHJGYao84ffOMdii5tJ1bbWfjVKYCgXpJMywBpUxahKp0bEZp8hBAHNfUDl/XbGYCWE
sZbc59QU2h6rQuKVZrKRshDpd/RE8SSW2qiLUepv3rDWu0dS0JbUsGIyQdXMU7J4vPfcrnfVECdr
pjcic8kttaUShtJTYBCa/xMxhk/t5qgUgeWOfBaYuzHpnD86UqcnZcg4/eEoZEPuXatPurDn9eYk
fNDQP+M9LF43VdJmOEJn4wsSWN68sizOl755GT9vv7s9KBrKz3/bs+6cD51FGqF808wXEz+kgVcv
LSByNhwaQR0wP80eQiMeHgEz6bj5KEf99wPv6UzF43888VvQR4ZdvU4qNrUv/WdThe+1uZj/5OaG
Yvg3LYpCqcIrlxBpsFerlP4o0lm4izY7Z4Z+eTmnZ138wvWjPYET7bW43J8P0plQ52gJ9XGV6GrN
KhiUpB8kPr2v2J7CPnVDbo83vYBSIh5QlByNcJWFp+9ux791nLcsufDg5Ku4iuafv4u63N+dvdru
e2kmF85qZUz2w+4UL64VDOEZmkdpEGkxVc8EI0aXhf+ceExw+Dz0nPxUWc6v613rc2/A4kPS6nK4
ZcMKk0cc3hN/AmBbvwbNz27RFcSidAvl8VocyqxEdFf9ctxWYJ2yKQvxFiOESJWyhkdy8fDerMjx
vFsbNmAyPRO1oZq/mxX/V0qbsSrIV/fetTiocMo0ijRFmwYUDbOJrwyxYbvz7rHLvV/sa4uFQUEb
+X7nN4wp2LiVLi0ml8hmcIj/x8jVE/HmnLEJJfTZRWk6V33D83V8jE1ObzjIGr+nlzg6A6+xyCpk
5TpJCml3Mqhsn0neBJs6+4+rOy2NZecBfJ+vplWtnc9t3LhfhPgTPdxV4uN1Vx4d2l5YArzsB9sk
ep2hkJUNQ5L900C0esE7CwccfuCxyvvy0ooxF+g3mLVWOMAA/zZPhz/CzN/sJPEJqP9NGjrMnWNk
TuuX9oYC1RPeo9ctxy8V5b/Fq8n12H751na6w4qkUdCQNDCgXgHLcZZoJxZ+v69StV+pPXHzP251
br68GuOxmI5etuO9sgjLoavI2te4HND72kCihI2p/wXNpRHYyyqRU75K4jOM8g8xDrK6jcJif8cu
8ddgh3EUybO6lAkbF2P1/8Sae8QahTEh2qb1AlQX2Bbrbwvyhzizgj70+1Gml+UJ0cAMAhEgbGtt
2QotkwRi7ttLExIH7g5YZRoT9SSwYcbqZ7ng4Nn4vqaxBBQw9vDw9DduyrCTL0XOANw3yMF+wH8X
9yMpoSINQWDd0tNSnnwW/h2FhJEz4BwRplzWfy21vSJwyThtxw8Dws6HE+6rWo+FioOo9yJzBUCx
x7lEoC7YVgn7Iv7CdFBoBb4xVoWUllCVqRjmXdVg1yQ35+JJvZT1ce/Imd+3IE/j9888WNjRwVVT
4b62oewfCjKOXeqcxcVx51Uj6LZ4iCYcLItj7TDWv9er3zaAwXAChzI8P9ilfmWF9piZCOG+F8QO
I/VMR1BLhuu3H2hB4TUH8QKTwcFJWLaobQKFTVRBSOHOFJRajb90dLMOLDn16B8BTGL3seUdjlUM
PEbXs2x47E5hNVk1AGpCkBIintyhAy/a0l09JG2Yj4AakBVYTTmlHZzx7i8tsUtcuFI/pK3z8apI
JstlVVibLaC9vO5fnY3vJWl+jGQ94SN8CDev9iaQQ/pxK308dhdNSQTJ6LJhCVT4DQZKF/Qe6bZC
vmTeRXw+d0+TBqCZfdgrxabeK1PmoQtq10LMhb2syi4+xnyyKZwGDqe9L+tr+kHqh8mpil4SSIAp
e11KSQNn5+dqfI6WKy6gTHfQGhV36r9zIu3hTNMI85+qa08D477TG8xOGtEukJ1HqqvsItThsC0/
yNUU09LxYkx1ysG6T5uezTSW5ylzlNniFvgPFeL68+mEwDBOSKSHTRMX4FLEpo7xjv2feF6cwcwp
jVIgTV68y9Jwf5utcL+AEMdENHNIX3pSIiLuvYWFWH8eIR7/6RFDxAWlkxfcugZ02Otlv1YilkwQ
F7MiP3TC+fEUsd1BOFGtmW4IrGieYtNqdUalIgxjZKmUkS55+kxt2cJG1Jdt8jidC2+MynXb4IJp
yDExpE+q5Z/z6FZfxy4BDNc5SyoSaPKOdl9NY2ZGWfeF9tDLPYUlEv//YBmkoG6mlkYXFk3ABgM9
s+3c46y5yNd9bdkItuHzfZZr4oAVMS8KhGbh+PK505Z6BpZpxGvjfivyk3vwzl2e6JF0fh9LKJs7
lqaeWPXnTrQOkJ733OUq86BTU6FFh8MqTSG4th6FVJv5xCxLclnAgrVdvtcz3/+zkpyQLpTKWAxu
E9bmMUex7oZ56RwqMPqwi+ecfNMsDVAX4SWiQsp23dM+sxmumE6cZoEK6SpwoqV6/sJtLv/GNg/C
iLyiX67oGrr78rwUlh/Fe1BOyYO3JxJgey2i40Vv62H1413pDPHPvdzkZhavzInsU+mv71fhm8nv
cGEN5dSQvaYlWCXlxQTlkHmXDxtp3z1FhTFb486dydZFuvX7bwSbQrvDI0DYJ6+xI80daVKK/tst
S2co19qk8Sc6kooe1HSRfhzuNb1E2YGi52LnzJvJlD1FIHKr4j/wuWYlVExGeqsBvDP5RQFDHTrs
NlvE0cohFYKe8d2v0AOqlWGiriFGx1aJ81Afg1DDxYCn9f0zumkUJAGxMqOwWBDfCWkjBv8mO00P
3AG1xWyGYaeU+jM7qbpq7xq2G8gjb11J9AdDxNdY7a0FjYev5bX3Zx8lSrHhplJJPmU0IpoKu8Ec
ZaWBnWDDLpZfGmtDAvDoXQkawVNUJTKS1ncITcD3N9RWLP1eF8IhqS/3OehVe8pzsNV37Go8g+xr
Y9H2nxB0b3jx8hQzJlwri2eYo1osi9mINMm0Jp6Ioi0/G0v87PTsFcR6FaQZ/vctvKFbfR4HAFRs
nnJILktqIledEt/zAGkXS8Vh0dNMMG+R0ojUTWswpp0ra4LruAMUEnybwN+Nfjuj4FSRvyTE6IiL
IEZ2Vd1EXNoO9e05aqHLVc6sSD+8Ev7uPdwPGqpST37Z/EucaJ6Rgqaw6BNi6Ot3hDAfFyupHZ2H
Pxs0TFHFxfDp6dh6zWv0qxy74D83AtInJP4l6U4vJLSfhFUxY8A1Nza/YZsc1zN0Zj/KtfZoX/Cq
f/QXQSSfm4yOju8qdg4m4wpgEwUriv/wYMWo/+BU2ed7OaCDTEA+8bf97Ts8KT2wxi/aFafmOCdO
6mRLVL543mAp2CYPORCvdniFhKjTPu0iOG55G7c6IWOIHxwx//nYRtytncS31uGRtv922e9ZTQ8f
vYYMcnkV/FUDnh0GaHs8xkJ47h3OML6rGCYJNiSCw9RnHbOfxOodSH3vH9P4cZWqrH5jxTwuoUQA
JXEcMdMoXBhPyVbPLo4iZz2OwYN8/eWBROeUlnhJKb6Ei3ATPjpgQQ0yQ+Y5aYRy8BS8RIKFOJ59
6KXAqEW9Y1f2A1ZejcwYVO5FqCqXO61RGlATYbUrPO8vYz1ZG++WvZS+fUg1Obngn2tYsKxnXktO
lJqfUoAp5zv2dVHPYYRZEGo9sL3XLZs94ImBqyEvIBwwpdap/ZuwMSBqtktSa8SRC787Im+nRa2i
UE0TnT+B/ei8LQuWlHQ3k1NMnMe3lO8ndBprBlehgDhbFS6pHfrMNicSjntPfh4uP6AmYFLKRifQ
yzd8xwnCETEuwUSTxDH/g+38ZXfHWZ4Vh2nwtZlDYknvzyW5n+V896Jeu9R+QEiZc1UzbWiiD9D/
bQQ2PdbtDWQy6wCK4T6LSdSULFMwItKwF2bOSsUpBcAJ3payWO0YUHDGjCG+UdB9Dj3SN0AZxo1G
YE5FOjGZ91qnr7ULWRHQbYLmf/4FFy2XG9XGG1eTipNrmvqnZhqE3nwWVioS+lUqOCrUB2LtWHVX
tNmzKoUcdn8d8LNN25tdUfoiw5B6olhUPVvi3rC5oifvsLNOrz2QDcazOp8naMrOJXugZHk9ck0E
ekPlC5j9QUbfGHxmlPJtvl444YN8RtqAcEnYuolPwcnQFGP4xHF2Z7rO6GIwx3M7UHlTBzt05WnF
KQeBzAp8mJAjU2Hz1ANGRl31cDV98ky0HsqTN/ZF3lsj3DkfXpyJGATz10zmp2FbwgQeX01F1MNh
8CYgTTDxvrudUZ3qEBzjxCPji15uhksGfsTy2jAg6zJ11osFp5RFz7FFW5BUkbQ11EMFb55zzKEr
JcU45z+w/13c4TMaR1CgALLuPaf28d1zIJ1AV0ArjJL7o7C3xJ99TgG4vKuKbx4kIdvUBh0CGoRD
TZAH9H9/wnXrhGIPC7HbIvq2ZwUVtb0t3E1Ifmovs8g6BLyVHL0iqmgf0VQc3xsykME7BY53h8DG
9pSS0MKEXkBiExiO760i9HP68gI1kz+91O5inTd9FChhQU3gjTGf2bIWxHaVj0t2Qci0hemCQgRZ
/VfRhHs5xMKJnm+VTShTwU2CJMM50LBin+7ETvoHJoaFiZoz/LonmcggBpGWsk8J1aiUsckag4Dx
kSxsAaPsEt4nxxyJBqrM8y5Fx0nwZ6jneLkTKfZ13RXhk+jBYPH1T1qfI8UVkHXInSwi8KyU2ARO
Z8NEn7Xva0q+sWHozMOs7DiMjoxlvp3E8TB0o1yuuDjkDlc5Oaa5Oxd0m5JvY4DQPCB9Ecv1luOi
Y/iecXg/jEagogxFGH11UAZnJ/P7rIEjrrsZuGmlQTv+90OdFVyrnuqDCGCKPxdqyQg0tgoLo4uu
noocAshupqfX7UOA1og9ZxRLoI2eiAAjY3v7SXSh3H3HG8Wa9Z2uOjwXbmU5JmzE9DOzU5jlzDy2
1Pgo/bZjVDiamemXQ1nuGfGkmkER78Nlxk6+HCryMLpIVuw31uE0qnQY3GqJzdtbdUHnpl4gqR1L
KRZJd17by08VtgIfAaKj9QksL1rluim+8ujy7Mzb6nn3kUlbYdOeXSp462FHn53VgRxsoKAy7l3D
5iODG9CCNrOuUOPoHpiSHSAPhLNtVxBekhslOiML9KVgc/ZoAXKL5Ibt5b4nPR0yHhmWi3gzmymG
V64K3pGBpNCWr7ArwG2QKTI2DAatfklQke7kXwH+nkZpmHLrk+faP7j5ex0SJLoa0cI0zZG38F/2
4uTruJ+buS8noY6D5sLPut3DHcxU06LPglJ8/k3PndyOb5cRQxcwiasDVk4+VRMTNon5Ex6WEw6h
gC7FzPqCmcbsP0Bnf09HQ1rABELZjTMD5zza1sEyz3IzZYUoBfuInh8IpQUpsNyT1wxpg6v3sf9L
2hw5v0QSuDD6RZ8yA2Hog+GIarPw4Y/wqRNWWoVfXSZ9gq6AkrjFPxAOnb7ee4u+u2//vlu2m91f
yPCyk8hpAxPtvyVvrEGopQCzuzPlNfWiw89xlIdbnU9OD1GTqk5bq6AW3oMXdHR+4ToZyT8p9FOG
J4aWwIBlaJYRnypUrMZizgtkWTiz5WLpGfPRNcrAtC3VlHMlnJXemK+OTkT5VjLDPxBqNHA02GjI
oMW6RKbO77S++yFXrrHCyChdI2tZe6HwdocEY6cKCWCXbBhGvD1bMd6DrybQuk3nczE/AU2eNtCj
PWcVj/salCKF+JhTZb0VPKFFB4/8mNXSruBM1iu0+bU+rwkm2isVrKW29svQU5ThONJngbSYMEPq
Y13Akk3e0JBg3JknHl2fFR+LuNNatLk6SahVnP9WHQi2fNJwTXsCG6q6Ei/D3d3jD5tGEq3/D/UA
bCgSDFMzrWYyD4p0NVeXTr86i+bI3msq1PR2+J9f51ik33cUG2c9CUfV8d7masjt7m5ZHg5/k5IL
rRbxvrp7urhVuhSHMo7WXze1by9v07vsS0QZiiWSEKxzWdvGdUq3wjj6NaOCq7X7zvuguturUuVP
LYccxTEj9vGbAoqhVn8jvGXXq8v1vSTvLlOK8oSF7h4nZFAo9Sxo/mPhK1jt2qE7CF8NZGDKTcHI
yNjnSfczfHUXXv5yCK4XYqCviVKVebBJiakBU3BeY1tVRUr/5hgwIzhSun7afQqKHjwZy1Yj34xP
Vx17GWBWnEgPX63IRFS3wr5TIyvpfmZWeMRlxcWtmtVgOkovyMd/Efohau35SxN4bwpB4y3KH0Vc
P+o8wktSgfTlg9nhyTT3XyFMWN/kuTbWKJHVuNsurnanPDX63OoC35ymHKHNSJqla2TunnA6vcaT
AyGvVBnsQ31Sf4Z5UltnWZeNk0yz2mBreuaHdX0/a6o+/fuvXFqsk5Iwc1erYkf2a+wwDrk75S5Z
4hAt4SYOauCC+RCbX21KfcibS4i96Qkx+NO+gw2TvCAGfpQlY3GeA5k59jEZS/lIhgixReN5Xp+S
MomhTtfsLdwEI4WGLCIBk6W/qJPc4EJ6TIx3dF+TKbuEbvx8zgSln5USe197yBYTb4WURfbuMLbh
OhdhfPvhoTfQguuGRvAH/th/kXJqCoFuwr3zcnXaMPYcmHi/gIKsEYhhgEXYvofTVgHsbi5C1ulo
KdXPpmFu8Cc9NiROztVE4plygPZsfjnwE87ajsuvmWrxiktO3KrkVdYriVjGqEJcYOWc4yWjKdZ7
76CPH63NX/cVcs+gCI5Ab/ZPvbBC8Gstxmqb1ORa01/wqPLAUpobjiKwX3gNVutobMvcBzzEW7Bh
LuXfvrlcXIe1fSTwvm3MLWwQAYNakjIJqEkPb92cB5WQsSzatye2ZIBVmZ7VSVTiXMjnXNUgxGSg
/Lhr9YsfCGtbQE5hkf7q5i3GCrOGvvqKK0zz81h81IbDqMp/nmfGaUN2XTF6BK7GVWHOXV1xB1ZX
IrSNVP+uh7ln+A+2z9vNH7KGCZfI221kEFiK41g54hVCCnqbgxDJeVNMPA1dM8Rmkhq21nDDastf
HvvzyS1+pkEpPCP/Olm8dHUTDPaV9LgwnPAIFeqxPf2vWTbB6TPtHuvqq9auMOPE/H2+RdX0eCMR
iPh4lP2E9Snu22jnLvo4N6wNCY2ig8J+woUibdA46l1RTgOhOoei1Fy9lCBsIzBJC9S8G2c71JHI
MgwUCkxellaXMBNn7cPvPBgcjPSh/FrZuubwlv/VnE3gXIACeOYK5GoAHjzNTInGCfnoAQYObOJH
VMtzYZj9+4f4Hmzhzw9ZkLRBWfcEg/MzTtv1pzWdqn4xKK3ATlOg1WDrDuh2l1lF5tGDYl8mIECn
ukqOpDuY3V8BEdSx8pM22urFwVxitFakC1gXDmQ7ivw0xl+OBtt1laNkhpTsJ0rAXtVZxyuNAEKE
nzA2h4j4H59GG9WlOE6hm3KgfcVcyL+W1uFo8W42vfHrCuYntuJ93jOcEfWgqSt6FquINY1sE1qK
5IDGSL/VzLtE0ISKCfSJTNqaZCoeRN7sh7pZaBjtKzzJrtDYzY/3+d4C0Jj08m+qa6ChpNmimH68
DRdr2rcrtLLW+nQOSIpCkIoIizz1SzlaY3kSbKqwcKSod6vDZVyaR8PE6KGTg1lQhWEMnPFEjnuy
upAoKvkLmkJ/u8hw/aFjRx2arxe7FkkrezOzB2TlP8UuP4M0UV8zPUyjN2b69gUwN2DVGIikfnHs
gET2fdKjsJWig406WVtzFSiAidZbSh8D7yCIVJchaOgC1K2G3m/38M3VRlA+BjF2dg8eSpvSdMvy
c75n9ZNaBuUtJn+wlpwGiDwRO81Bf3JFJvi1AhwWD4/aiFmvoCrpb9NtvcTJlOMpO7Rf+MG2mc0R
L7aQODBCfrXK/HxZGUnr008AiJ1X87F4zfJI9P+CBVDDZuOtylZhH1ewpqUmdCFYk7vbJhWgvNLX
kQW7O9KZzke1C+hP9JxGqVUoXdw6IRzaVwobERFoZec+T8Ubk4lr0EaCAJnyV+TPbXK5EWFeDPuA
ISAuUeV8Yn5yMDG10+t7Tw78wCuR2q6Wf1edoW56FMBVMhvVWulvzoeRDQ2bqauHhLRFClmMEIMj
jdMagx/TZZYAuQhLIUM5Ri2ieiZtv4ZsIBwzHh5qNJoDyCwO5A1x0TJqRnFpHizK51LZQlSXNaDQ
FYdnEFUnx68cpYSMsGTSCIXpKlf5fQAtkwYuMSdvA9eL4A7fGJZuOjA1Z4AEJwfIss18FcJsNq8Z
TgQz0vDY7XuyaiT9ZNuG3r5MjJMUT6Rjq+7kuaiCHgiIr4A6m7bo/SDhCPlYFla78vfg+gBgy6oX
aO+8Lt2zPGngxRIkUwCO4F5WEizrprpOUfPMn+bWFOM43HkZupPyvYQbc92++rkcZ0umUhllGgsd
joXUhKwE2gFN5VZQZ887VvQseisCytpREodx5cE520OdYOfgAfef4OM7hvmfzp8wG2gId1iAcARk
QLxVbqbV73Q/GsnQxJeyeBQk4NEcleIFUxgsjvY27wxvyeBcumq/T/QQep0esmwp1Po9B2C6gBmw
SczrQZFRJzh2daItk/mskCOYXL44fYS1FbsD/m5u/JvXWlTXBkh9cKDdbz2AWfHTs2FQRaPADV+T
jfUqDYFSnzBmZt/bMbHxFPgNuAWoG59htxoCkrkxnJrPoW5UE4b7eMZg6NVhhrH0aZXXmonXTGMt
jQcbE9KTAaZGoAjpvSxCf3DWe5Re8R6PfwuDOGqaaeyhiVuD3rptxxQwVH1l64UV6GxZGEN/ByVS
aK+3kbuplnzFrZwuXgqd9xsivHR7Vbgj++IpweqQ77bYSBdyAbdczznXE9FBnM8aQafX3QDbwrer
8dDJRD0lzZLascD1QTVDmwWAoF1cXehUQMegdi1JqfQC4STWYLlcasuiCUXQjg0UXfufktJvcnHK
hfvKHD+vHXf9GtOKImW21GrQjGMQ3rKNB8586vVdFqERpPcZZ/AIGI2EeS8s6EEAPcYff9tt3EsM
ws2OXaqXScsFc+r70oi2eB08dx5/sqtWTToI75oN685e6XHxNxlVpyOEIVKXilISLpZNYajmd6Oi
jhc9KBe87XT8ge5mOcczQDROIH5uHThC4mFan66zV89sNTwOdMoAk3KVxPhr9RADTKatqTCIOjgV
V6z0Iws4lM6qqiOjrEFlzOIPMJsUqPFMceCYm3Dyudq5txXLZIZyREiV/DuU/l74K3CpFKwOnkaE
pkTjQg9TpsEbT9qgh8HRNXdRs9lGEOCKcxGkjBAuFKKAiZXACGfqx9toR2oRtxpamTmSQXBbvIM+
+EOiMIGM4UmIL/4HMgxtQgnL4tOqbfSbOlGS8Ec4yMlqHV+2XyN7bdmiGyPIFgAmEZxtrfAu05w8
ChijzSoPBWaleWx/cPq/SSmyB6S+h7OlMtl/uOeokY+Xoageg7mxQq/8+b2OzKUIwMOTELJqIIzH
okx3eNoN4Cys4+J6w1i287KRLYXBB29Wk6bOBCS2wVvh8aKXjPZfqRtr5AQg35QF8fpYELOl5gfl
crkVz8BI1Z7FRnJtKAiJ6+fweLr1s6HEPSC1alh0Eg62PEweb/yBiPKDOPd6nOzHIsSWKjlnPyUv
1g2XNTV2vKmliXWPB1DCDJ5JKvJg2pjXBbtyYalEa8elu/y4AFwYW4XCDguhuk4b7FXdYcpMfZMd
pQfPHO1vQfBX4KLO5Seo3DdCKeNb9lmCBOWAZO8hA1ix/BfuUgf9dlo+VmHIjNgWVXsn/V9R+g8h
U5oavaPvBojnl7ZhN9uOm5pVpM929Gig4YzZNgIPlMS7b4Ana2QPwXxfEA6EyKKwx9XJVMTVDdz5
smgD2Q75q2jMyCljHEvgiswvNj8Sa+zAev2thZcQVF8K04qxQcr6I8otK/0e/TmRw542TfPvRy6L
1B9M7oZLWVliDIkvf4b1sqDDJRZcYDNGFUVfMCe8caujPFa+C/atb9qXa7nxIu/FRiefAdqs/DIG
RM+JxDYOcc0+BZNPd1rDzvmWE/pSLrGE4lQohB10yTUMVq5oH9YyML/6c5hoY5lIF5havKAq7twk
V02y9t2qVH0SSen1k86yBfcxV19kqFQBMmO+5/eHigiX0iBBDG5q+VwoKxZqiFbtLjpXRbHTZ+A4
Y+6zgG6ILzEDeFUqqae6hu34pfoDbODPzZp4KtiTENioPr9y10UVSh9Fwt2/Obnzi9Wm/NkaoBYX
UaFuOuDs92mKvJiQti0d3aOoeFHOljtI8ufAcEKyxt5oMuoe/ZOqlsMWr6IEN9BdxfkdmU8KPNDn
9uTAo02TUSoIbsaIKCnJ1w2BJNzTlF4nrHFvrSv1Kd+t7afnbulWJrtUdPB4fUfHRHnNnOmz+1Xw
cWlwp4JZRFt67F3fI3BJ8w3x7WWVaOh+qSjSGBpulygQQm94j+wb2j7yfuHYg1Z6jnZsDucu9kfL
mr/eX8ITVLvCOKzP8fapZ1xYglYkdJE+g9Ax/Id6JoJvsxcSgE/4EV5NyjmbwoW8R+oIGFx1K9t5
HVzFYbrseAfk2HEadwrrNZLb1I1Yt9fRi71o228rRVJX99kI2zg16RRR4wAyGfnTi08yjShvs50c
OM/jsZRWUEUg65FwzKHEyIys9MgVlqJxAHizcJnxYPJd3Gnpb7P9vsEy8/LZv78isAiBMDF0G/mX
Qmw3fKO8VFjCbhmhp25SLIKNPvZxk0FZ2ubqOJ8N6iOF2pXQFuPjGrdz/uyf7PAtBL8fV1NGA+Pc
7kaDVtcHfIQOsDki72BWs4pLNBhHOyrmd2Vsxz5VMBsi2kpxSqklZtVV5DckcR+MLvbwyI49B/8e
jK13mqfMGTz57GnVGtTBtrpT6rPwcoAx+Bq+bPG8d0To28VMNUSY8P0yqr5GNgEyuW1CxK7FYUZr
ZNCFD0q+HAbvunMz9AZOmr//ykY+fHZOcbffDNAES8GRJ9KcqtpSrZFCLWcNnzm85NlYCjoTWiI5
0AaAuzRRkh1V8nWrzTnMlgtaCy8yMnZJfp5nuzDRDITp0MZuuIL21fUGll/J6yHORGFolWVziKCy
sToTgjKKb43y7WOkvNGhTb4tkAkFkCJHSmlxJFimqL/YVWTc5ehkmUoJ9EFFichnr3fEhVqeh0l3
BgSZaf9WLFYABkrX6Mjfwm6kx4sIWahT8szZJloslidgqIVv+1tUF5JKNrSWbwz2N7nPId+nwIgJ
fLBuyVw6UMy/ti8Q2zoPA/lXbOsVtOPGWC/mv1pyGqENybO7b7vKCplzcetMwPuW5POYuOdYbV7G
tAxKpkIA3uhTx1a3hOeqL/D901xK/dSY/L3iaATkzPOqzuR7sbLqdVgrV6cvauRKZv4wzHeIaiDl
LT/fRmps5DXFpU1EMP293+omUGMZeThmzTc0yo2hxycFOi37xCQTHMk2u5xY4ImkXeJPfMqLyFII
DbPOhury/jPKUIvJ/ShE1wfB/p4SDd6FAcRl2OeQO7UB5zezE7pHqfDyuepBftN6ewpho0Qg1acV
b2LXYH2192Ej2s+01tKw3hjhc9GFUcHdeD58JHvlPZHDggm/FDcVm/KdHwobI76e3GRI//c3aaIm
1eFqXxfZ7FjhNd+J4+sk8S1e3wKYAWPxxdDPTSUnFuvsaeXzrCjqrdBI2KDd9KzDXsI5xMjYcFqM
1J5bpWzAkL/N8d7g9J42W4RW7g0ByNKmoAX66iXgcCsqO4V+UJP2uHf937SfhoWLFnU+Biey8nyp
oVfaYMWXPuJmvhJvvzjI2NQLWrXF60+xDCNRXkEbSOE/if38zpwVSVFLSOH9xAXIix34n5vXSkGX
6P7WkDKWU5VG7iwpynlpw1idEqc56vNHevsBYlJi8t325xBu7ShlS8/7IXrIetONxYHVZKTEklCn
pYJKM4PTUceW7mNXxSMHTF3Oc8pjeiW5qw+AQXnx6+CuaRFl3iPa59TRMtOgNSKPwvhT+MhsLUd5
NF5rmJx5cUAfRMb0U16Z0siV9YapfZceqM8IGDq9UVbaW20Mv5r0T0NEYugiEdddS/o5UtOWBRiI
ufz3SokA6md4OYq5stCTMosdlHwlBHEuDFtQInwgzkj5kUhGNYzB0KwK7yECepBU3SNQRSXbuhGB
PLy/EI04KSB986taxFLbDSeDt/e8AcmoSgd09ysGb50chIfLPjFkAVRMkpeXVRNmgKQDEuEvnwPN
q+zzUOMnJGZZ2Dr1M9we2yg4p9zi+JIRmhqKd+DeWaeXARmJ+lzO5FqEwdLCsa4kZDfqozOvOsWg
HwRHTaDvq8QHKY1P3PQZz40PFA/IvK0N35D/qkllUAXxHWQks+04gXh/qceBNn5evq3QXD/WGE0J
IjIPXVc3Pg0TEvihGjWVu1W4+VccnZdULwum+z4gnCG+HTP/p+HZ+dPmKkC8nXeuY0pf163kjPUh
RZRBDSvcHVDJFLFZucc5DHAyXbjNPCVNqj8VVHzfNADAdEFA5U08/JbmbWz+QdxOzf0eOlEd9c0B
f3RXr+KNcHgTvgFgkglj6Qa75IuPp95/3d5belctwVjc/AQObJrkLGan/MY5881qb8OSQOBNHiwu
XENd8EvMphaY/2K+h7lyPDSHvJgHsnDsZFvwdZWx8wJeFwLbY28TarTmP0ogU0ZRvWxlmciqU/0A
QfR823wsi8oIAVbkFI42XlTJHE3mIMHpoikzb1i2bDQpfmESY3n3fyQnKQauig2E8gD/Ii4Dns9Q
CU0Bdp0SP6KbkelZDLNyq0jzK9hcLdxylvxtxIwcVzbXvAYA9Wy6KJqUu2zcqzlXI3pSdT0FKNd3
dfLEmfbuKfv3Y4dR/JJn2RISX+ROFN5FnmloZ29LwVVWplv5fVytaKCyzKO8s9+GGRgRPpj8cP29
5q2Bnu23ApA3HXVg/lBNEHPpdamsgn6FuMrprfZQnpuaQldNoUf0dH6Fi3J2aFpqsethMZHKSiiN
xjrjeqFSiWm6FvJT1LnACiKlyX3kZYtU+JgErQdgFH4MA9vwDqb7vY7WNNSCGie64+24bDg9eRz/
EY3GoDvHM0OYTC/BbNoulvWoeHQMtdC3kZld+4wJokp+5SM+p7hIlawts1okpwEh7LvS9o0gd6Qj
FHmLzZiZddO9iWHrtlwQ5L10Mp75WzjDZHrj+DM0DaPaQ0iSBPLYe8GnnXfLyAmR7QUBFRN8wh4a
U44fxgO6ViYZGmvm3lBTmVGNUr88oAZAVh7UDeXDvqioQB+BQ09w1CWw6DUsiwUHkhp0yf5IXdb/
k/wYr4sBnRixrpCaey/PV4d0HuxUbxyW5S0KV+8guaquCDHnP/iYc6Gz1v5DIlEl308VtohN4Nyr
a78kyzaFO8hb+5TkDFuI3VCK+gHPUAfnSR5NW1V3sVfeRmWSh4u5+GJI3pXEUlUPM+zSyXJK14JB
6IGj7rJvuZ8wKZSWNxR5GwuSFAvJI/fEsKdmFZf1KygdeKnJPMS5AfQ9P4j0O4crxeBeWMrleLUA
yhA3fk7droUIqdKsvKy9Gf/IHwIKnIcEs7+42747onBX3vhlHxIXYPMZvp4Dr40nQ4RgGJrQiVrQ
VnQQ3YjgdOoUKtRtZbbANlIEQDbzhdj1JdyQZu+j5YIhDRjsGf6IB3emx9AB83KuhJ3nqsJLeiF2
d0cP5z0bdP/+QWwl724WIVo5vS8qDZoBaEvXUf6o+/9M5HsXJEWsUYv7wLgWuHp8U+0A0vqBOyZ6
RtKARPHesKNuL1r5PNL2ZKiEAOwsCmLUho/dEKtL7HcuV/W1Mw0mGssmj2xmCheoFNFjdePa/TDT
aI5fMN1FTSGqtuItnuXo26ZtTB6pmacB3r1NaZC+OCCL9OBi+4umAFNLydP5ROZq4l9lyAwn47dA
/zAL+BmfPqdiuhKCwM08YumdFGehHH8vTGipia5aInxpqzH60gp3vHvNIXFAjpNpkqA0N2plRHDx
8OO+ZMWLpjU1ZY2GY6qt75dFBW+NkpiATR9QoRg9LizhOOWCRyVIo0Zh9prYx13dKhu3llQddk4l
9FOcXrTzuwHBbeTr6C2x2VyvChfs5EZTgPxYLNVr+LOlLHoCdTjKf4iucW5Y2x+uyDgp1u/YVDfc
+0rRXh7XU3UjteHEtCSFPVawqggc85YZ/2tEE3OnwWL5dn9RacRd32r6ach2tHu9ZCa1C2mqKCah
23fYBfFVC9cIibZh6nW7vqjC76kz/AQ0syMt6EN8F8GzeMQq8BTKur12OltNRDZV4h8nOy5+rKDF
spYJPwO2Y3UH5Tn9jglPi/a2vXXDLTxERnntwYnhNyXI7p2Vm/7CkdLkQ+yuqcBr46UaAT3XoxIt
VAIRFJkZYX5ItqLl204sGS4m8trJFFcvoHVvcRVbIOTsqds7oJdZmu/iraCGJ0eFmelyqMoNKKjX
QjCREhqsPZwfkrXi6bowg3ju3tbqNy1FOEFiy0Yh0u8/08/uWt5gaqqgyYlvAd+O9IT/4qv5su6t
tFT+mrmanPsvfjVa2SC4E9L24ed4+RwX/hKGG0o7xnvO77QOwz9C42DYuBVJLW7Djt0qwyE6QRPE
68Rxcb6K/NgMK87qPWD5t7CecMiGCmt+9BvFFqHrHp2wjZssfn/jflXIkOj1TRnfBMZdcgnXgGKD
Ok8zxTfSH42yFg4fWzu673qttQTs1+lZ0Atqug2ad5DW6ZHHUn9WZpORJ7MoNQuAIaPo1q67WaJO
Bz9eezstT48zW8taOlsVpENopKnCJ+05i3z33hfhGFTVyiBCtzApc+TGcv+mvuGCiRoM0OSFE2RY
Vj9K8iZl36Er2Pq3mRIowRZD0D8dliKD+slTzUv4UYs49uI7ensdxEdxNV3vJZXBo/GF8Ir/F+fK
2kTKJT8c86BMTtr2/o9HbVn2z7gNO7iVUlv+C90MtvQNW/Gp4vPrx8yg3QcXLaWMiHTeQEcZGSRG
2mql5MzrxERcCc8iKkemq20wJwa3O98DMylD5rlj4GYcEPd/Qy0R0P7Ed50lOPnww8XyZWR/Ix9Y
cQJKSQeQewMxfBi2OpsIQorL5SMwQow3AtuxemxMwRrC2PRnjrXR/YWDpBr3XTibKO6KBI1EtNiv
9ro6kGj7s/k0hJMOIDjf9qrBFvN041dBb/dExJr0HRJhgfVnwOhfL0o6D3N4kFnQSpj5WxIHmXfV
as7duK+kCIV7avS/tXq4ex+NW2DcDFvWThCxOob90SBy4FF+nIuyQhtAivhIb9yGzjsBu47MrQZw
7JB0TRWD+vCyFedb4z78cyN2A3qbCsTRjMIS1NO1vfgafRCEVR0TWM7Ya262emaJtQSAuBWPspA2
OOB64SvJVgh2o5mTJpMgHicfCAgtiW49gNfuk2DFjLWzVHO1JDPhmZ/OB+OmtnnMPh8Yf0qgNfhs
cG4R1kZfon2OS9m6yeyx2VuY8tfEhWQkjZS0G0RUeEEKGsQAvg9yE0VRVinvwa0r31vfAq+a1Hfk
LTrwOMwegF6iAqo5x3J7VhAYTgd5wPwoR4KfXe1CHts+a1Gu2yszFmaRPRa8mnT1DCJUJaxrpoLr
LVXGFdPQCTeuVWUEhpy8La5/35SstdG/XHMzwVqqKqzitji/rybfwu7oJeGiAVyqPjpaR6XUo3ya
8M8wUJUiPKsaHbpCZAtpRHw2e62GKfzTZIOQHfH6vwYLT34kUsBQkspS0vcE3cv1sbheFMYggu9k
IusQ1IGAXMmCcpLXuUZ2A25FrGOy1AE9B1Q4ylnvIHJhrUHnEuK+jh0vnVPSTaCS3dPCtaYrFU7B
47dScXtwQJkafFg6NVw7cWZ/0onVV5R5GuBtmCFdbwTcXG689H12ckEm9qVPEbJakSAPj16cN5WV
+hEaykfcm5qSDrw8kMMDyyLb8MMhthc+Sgq1Qjbcw6j/g/sXNCSA8O1iaf2MlxakC3q7j+Cwf/+4
e/SXEXaCfZS5mGYSu3J7ChGLHJuyKYiweQzokKNILDaWEjQ5jczVcSxo8P5Eoz0SAeUcpQdXqTIv
R1xf+q05qxpop6s+QIZBvlQO85KBfjI0wWmWksSiEVU+ZNdzvPHxgk3G7i2ndVl7zO6EsIW2e1vo
/HnJHkBopK2Iyb1bpv5C0APS76W4CpgZ1wh7wMPVpuMVb/WbxZtl/8Uz/16vxqPpjcIDW3i/6Ea9
as9QQcp1TfPNBf66TPq6FsVv7ozLYJa26BEnUozEGYKHlH/QmWyU3HZ/2729O8Zf3mMxeKPpUMF6
iEYyzCYP7uVnAeD3ap2F9xd0f61HXwhVz8tll62p70UfZiIJLL4PxcRChfYn33o69rm+SojHv2JW
l1CQXCkfv0OWjMd0rn5I81iu4tpChYO8qoQy11oQZ+YpohR5bOmMwdOBxxcgaaLzY5nyfyIJK5J7
nuLUy6LOhc5OnZ1TmtIt062QutBvNYgez3EfoN/wddIYiJ0teQEsNmXPjjpNilVBIzDEN1z2x3P4
3PtCvfffvOdGXy+DGGXW7D+1SFbPGTrQzQWsKBz/5O5KY9M6jM8inzdf8q9qzMNvfTrE+fA1t2xI
OBVKVV2xzERMDqBjIMspsemcSuP+8KNPy8UWcezJR9LAcrgAQNYgJzHPLQzVTTVP9fX43Mc/Pow0
xVByDgy6arcz2+hYrhRWif3/gfeNwmfTU+dwb91voIZ4bCdSbUrIXdQv2gVWLlkXQlOdx0Tn4CrO
9JS8jstD3PAe7HBg/DFBc5li0XMW8/2Cmq3kKZfLF37NX7qlBWaaNzPOniaSgxNjWIvlGHNT7H6C
AioV8UQAH9eyaUvJ2w8ateUOCL8APhSvuyurQ1o61Y9/le+FxTr08sGX5JQ9bbks25E8Sv9Lzozb
ljUQwD3FXRyoMZeQmhChucDbIWKZr3P/BqTVzj10d4PJ4kWajad94AI7R78OKsHmIn/m3k8e0mH5
QfpnFpHrh1Y92AereYYJcyw/bor14XZnidSkkHpZ8ATIEoFmuELvfYcqJyvNT9g4t1FFlDhRNeZX
r5MyrG0ZHe6a3dAXIdONWntLs1QXXo9nSF3Qt00J/t352XAN2IKhOOzB0NAoH/xJCqo3IIP4GxJi
X9Kb81D0ZJilTCLlECNy1OkH9tv+ZVM5vk8R4Qg4qxBFyaOHV7yIPcdThcqU4lieclaHgAmNpwpP
mfpz25gxQrhzDtE8+7gPnXVxat87+4ifEaiYoueCGhWVuevJeKiLx/v8wODpUAjXxxNVJtfk+2G4
FyB9GN1YAOxCF2y5dYPDB0mAe1dZ6miVnL7J0u00crhZiAvBYUgOFJ4tFXbXj925DjOvg/tNWd37
wPX+QpnBmbBZzZcqokIKFxt2QxHTHnqviuFi+dGBTC3B6dCLGI26RMeub64GQo6gjeNpr3a8Ryps
lLzxlSMvmCRu5LtEsK2Oo9YxP5hwid6enW6GfgZ8KTqmbzydkuWl7opaEB+cgpPW5Lzo/Ls+EKrL
fwkkIro8I8OYZi1yChYuOrNvPcUm9nIldTbuLqGKE4He35nuEtiBi/DYaiuL+GdsmRBS1jspzS3k
ItiZ7xvPks/X3uVdBi/+KIgiMZIY3v/RKf3Q/tvXlVX4pkCNlWHIv71J9XuSpDkbFWe2ZxJX/tPt
H+JdZfRsbYLAYTHvKEtHyoUuMXY08rGwNiDPPkvf/+JSrhcKX7tgwRl46+ux7IWYKu9/cZC0i+r1
BMSoxP7d8LvnXuUGEW0QoEH+eipoCZ4KY/HtV8cDSwCbIOs2ohliFHErm4GWrarxkMSMM5oG5x+4
vQUrWp/J1qGTNc7legV6Q47uVC4YQr50gktndF2pf4ADlx/zOW5J05Y113robmWLqBKCBTn/mT5c
CyoWRpaq5H7Gag5wATvPoM3vj4bHE6xR5tiQDlJ9/HbUG8428bqVtwB1hg9ETQr4ClHG6Zq3yPxO
578SS87b9156bVXF3CjezSvk5F1TTSf9W/Zj21J2frEUTs3xnw6M3BONY8IhB6CI8PRvaIzvzjk0
5fbKJOVnwiJN6O7fHYpZ6FjusYJ5+Dl3turKb0JaLPRPH/v3KD+mQ86huVLo9Vj0O3zmu3fGoupU
GUj48Fx2V6l5QxMKKTlayhEf2A10vSFrfMTlA92w89QPm2JMeDYM8pq6Bzf5E+kzj+x6cAfvBGyo
KD+7cDJLLtBEn5inK+14jbt3LyqtvrDCoxRKbEvWpJpdbRBxALQUADfWaeIttiwtiSB2ltfoKv0g
3JpeW/OsGZkAI2nPyNFTKUe5mqLDNtAcrAnKfcCt2QdyooL81kE+w6r3pk91UjqJ4uwRioh8oSSR
LDxsys362ufwXjtpxLyc1xfeGb7zGEHX+YJNq3BaKpR+9G3DAErDI2bpvSsHv8qQJITO2VZPsP0U
5MAuekGAGJBe3vYTAlT2uCL4zVxyPUquUfU1IM5OQ0HOK2g5p0ZbU2szYlh1Q29nyzRqFqye3SLG
7mlF+svviS/t8SbYP75vt2gdjsaPQH9ZawoClVuosfiGU2svvhKrj7kSsWVWa9kKrksIviAMZEeu
o2KElEM6vr91FgsPotj/ayPFj/KI63CF3SsTyVq/zwyeE12XHYDNc6DZhyYWF3aeVIj4bc+6T4M9
ZwAviZfoO0fOyA5IwBnrMI5CcHTftukcRs4IyBt3BCZRChKP7m883cUnuH3WpMhMqPYQipjeUIT0
S7SSrez75eF4E4jqQcNSqYkLI5YC6SyiyENiBU10vz7ok+Koq1v8bVJBmJk1bhxyvVp4mm9yky4l
0JxZLw6dz680dnTtXOYjqFU2QHUkv9A/8zsc7PYCa7FWzJad5tGUIRDS/wq3yNrfbIiBdg6x7Un3
OmUTFrWQmrfr9lWI6wJflu3TUsjIx47sJeoHvmnO0ZYfNdBChIZqAPPbxYom4kV/3heJxgssVDmM
5rmrj+o7E2sR3NexsGApT6RXel9YLjCR9k2kIbDjNOttvAOuTnhMgCvom7YgG5an+tkWg/fCMbfR
GkaI68uuizSRANZgy7EJImK5UWXHvXkcPY/cjv0gbifYpf8ntVfhzWcmbfR61oda5opD/0xoxmxw
yZVEx9mZP+lvo28C2uqzkhMWbGQ1mPjfizz1XE22VnlJ2kuEDGCc/tskZPMu3eK6UA6df0XLq4Tr
077U7FXKomilvNDmoZi9kC9zI+EFWC+/5bNCmIjuiU9cCift6jDu8T4BQBVYs9LaMhxgWJdMJEkI
nBlfO5CIs2CL+6iz09nw+4TypGS4fy7ifhENM3JspF0mSKrPwlKIGgLB6BmFEcv81Oy5syjPm4N7
8D5e0SkbiaYHIKLAB6Rkh33x4DX8hM3IRuMX1Qvpe+6wMP8ihlw+XPa/gqASYaeUIp6AbdUi8Gkf
sHnWigbTGErLshW37H3VU+vKizqVizwu5s1kp8vSmMpyLQgoVahml1/OBFMYZjPwIW+ezjFOTXpk
wr3qvJ780SSbvEmjjX0v0YTihQlrDq0EDRaihySgY58ioZK9JiOdeAdudd/JgxwqPXo9xd5HdXpZ
pIbAg0lWZsH4JEurp5ZgONpGSiAegGEIBxtkhKJn+hz5tGdJVIgKv78nVYGIV7Xj+0U3iSE7HVRM
pqf05MKb+8EheDdHfaChVgZBe7BtDg/PKF+rRjxvsKXe1EcEeB3YkLuBwMT1qY1nptAUZdG0KVo3
sUviAfHvkDRzT9G+tCPlKya9kKn9/0lQkdGHauNUekbvgM2n4/0j9F0MifG4mNv5NjU5SiAmtXGf
t8r6IJmxHzC74YsmA/6SM1YXj4J5dueLszTnhLgBvulJoySoKFg1tI/k17/hZsogwc8c/cW+k8o8
9S8cbbEiXEYBGbebuOuBUAJwTgmi3/GJcECpMfTBGUPuaudEOrFNd/0175JWDpTi1Ks0XnOdjGBL
fpIM6MKcLha2csYdObsYT3aeDQJNxxN2/CpmHLJzA2lkcjPWvdrFOoNVHzxSF5FLd8/RsMV89N66
aMSpxmJhPg6S/0CzpL9Br3ahQWtfxr2x2dxM/pHcsJXMug31Ao13vTt/pCasHVyRv9a+HJzMPGmE
4BdSj3nIwQvdkLjnjRV9xUhtM1PT/DXT8SbhqIqbJuq8C0XcsEkvfuKVrxhk4I6dTa+PE4XvZrW4
o1cGr1bGB3OVUFJGRTpvs+i0JA5P1vf4j13G955JFUd5GjDlQODZNfZGHoItT3RM1kZuT8uQKljR
NzbjgAN6b/qaXg/ETP1Pzq9YR/P1Ewuzhbtw8CmDs8vwBPQhSHUZVOEa7w2k0rYG5FO8VdN+HROK
+vqg/yVEoIGuWE7c5aUNa969yYrOqKPCWZZWq4ly3rSFOGJ8mDMRUSXb0SvP83ABQjebzk0jdXI0
kXP+gXs5e8L7nL5wHpPnoDm9K8/95HjSIRJJwOy3DxzSLkPgQ+HqWs9nOxYWz9jDeSpWHDRwYAv6
pcKgp0iSIIHvOO+CHeX7LAXEsri2ZyVz/q02aoUhmhcagelogcDiZHw3roHqaivx/QEl/XdsEuxV
nkOQscSSt/AGaORDbCeq1hPGqan1MMXSmj/15jldlNj+HR5NkTcx/xz0DYoe4UxTtTRqJkOF+yOb
/5fQBSl/sptCiW8PgOF1cXi6ztJkc0tu5+tv9EPUP9MopZR7zF37F4rnREyYxEnnfhlJDm7F+7kH
OtG9JvhNyP9srlpJ12nJoeMIscQ/jaweC/r3a9WSB9FISQb8e8x1KivQymBDcu9Cg3GgKzgIJiGx
VPYENasmZBtHEe0c8/SPawI7wPN5rF3qPgXgu817EpNnwlrZLNiV8VWgKUPWYylL+LVQmHIlix5l
gKhTvALPxa/4E5SIngb5PekQkOS47vzF05P0IOLMZPWEkWR3cMFJ+V1oRWUz1c+/p5g85e8bdcLk
57zq2mah9EIGDoRfvStz84FnXOezAw2trEH9o/uVen5FKZDIaVmHGXWe3Dzr5CnrsuQZqFHys5Ws
WPCshXSUbNqTwydz1+YNAKGrQ9ikfTQE7hrMyJ9bS+45exXxzylojkK/VZG/LPs0oZCPvKeNOpRu
qxpIYj9zP+oJcySyuUOKUEhjyKc4EHzxGe9gS1Jn9c5izo6jahrF8YliB+IUvhyshlRYVq1TjJO4
z/1n9XikQ8G2aCg0WRgYJeDuKlmkwClW18ZeDULpYJ1j7WXt7Ik2xHfhNZdFBMEeFwjugrFrFfvK
0H0AXl/Yp/H2Dmnz8nDkMW0ezC1zraA8twsE4/RiW7Kctp0VPsCbmIGJulG0CH/K4gARpULPFOUw
QacXyeWcsyYWzdGfTc0UsXRDsbXeqDUtzRob/X5f+WQzhAbeA4wC16/uGq+Zml7bhdLSXdyZmhEp
ilIch3DcuAjaoG2H+0MKuAzcKldY+dLUxIKRraKFQhZ2lM0kqV6hBji/EMDDQiKLGobvigRw2BeP
JwoUK6HsPRGn6nxb0/ba+oM3Bmvc7KQQHVCfJxfR9J9wVKjVSyyilHnG7OMq4NCNxss7SKXiG/nK
XXCN6NC5mM5nZ+Ny8p/S4AIRz7BGmVultXmf49TtOXqN+BKGtLXFJp+DdA7AGSN/vvzJe8jGzwtv
G8ZrU41jEtsmLzjppNTWBfccsxCAVCJIVT2WIAn+9FCEGxVefUxsP6+mi4yD1sAs3dxvynqbaxww
yC2TfdKCSo0kxEljdyVswSJc5sU1ph8hXEbVjiOBXObjdzWDnzLxnKOgNMqAnTiQf7Ecgjc4y9fz
OR3J1il/VDaRpMSHqLm8h7M9FkU4h1iotTPiSdf/JBiliqrJiFtP9YdFS6Tu6pySwwRnyoWoR6OA
bw2qXbh7V8JTn03WVffDgKUuY+nQap2ffVVzbbWecc0lEFulMBGHxNvUM+eTlXBHAsXh8kMal1q8
P/J/0L08vZu3sVwY8RibINRSqQ74r9e33IGSdxqIAj8m/usQz/F8g3NiHAXzv6u+SNuu/a9kRVra
X4djzEeWpQcVr9+BweofgEftW88VnSYOH0wLlycymzNcUphOQCAyhWY+gdJF3eYze8nRpObtdGsD
ZSJ05yQgDV9GpTAGhNby4TIpHMfb0JT15elmBE0sD1drACZvCrFWGvXWyAt1u2Zw2S+1cgZK48Py
tStZDiV0iRRLMb5l6GlXwFHdBqZ9v+XmTi72MWd/Tb1mmzRTnd1pzQx0uMFfFZxHxqGVxOeJWP9R
Evv9C08rXDW2v4gmQcxwjRdq+4CMh2NlP/KXoT3MmmxnnopZ5RZR1d3CY9WB/jqiWOd4fpx6yrgo
Oe6NzotSa39Qy9wUAdnVky29+i86LLnbNorjNJXilPv1P/wFWfLLR4iV27ROoLRoRJ+wM5UX1BUL
bHJQw7OUhMpcKQmw7A+ENSSwI92XWOENDio2YG+GU+BgDKbZjd1HmbYUN29yphNKq7nd8huqEgQc
Z0Jfir8HJkN/ue7K/9FBqGh/8GAUc2P+wEt4PCpOSJ0psu5+jOK05tnzAnGthUY9BISBozY1W8/A
6amoSYEDA8RCK+SVLTCd1pI+Z8wJaptxUHDlad2tNuctEqMGzFp6qynhZ00bUtFyY69GSoHwRFqU
wJ+wGKx9cZM9mepC1hdHXYKp1dfqHEk2xg0ja66Qw1EMEZSIhHXNfiKrCJoZ+GnU0GaJ6Cq1cV2J
PkE/LNMOI955R/xerGxXK5WYUKi4q74uEpPdyCw4GT1/tI1xdfrbClN1tybKgamTuUdPX8Vyadff
IngHggNfoQj2a9v8oHW2EiBrh64MM+p+ZEMENKzmY7/pJE0qqgm1jss6rMK+FsOvKDTFN6ZdJxgH
6bSHuDKucj9UlEoDkgntTFBs/v1DiJf3LdQJJsilJwuApTr69pkuB1LZf5feI9SRhuXwN/x7E0Ap
6TX+3NRUJMllggUVn98m/zSG4F4h4qJAFFE3fgRujcQkpXA+vHfOpLKXJmROEuQX/3mlyx7j2thC
kis1Q7F/63e7SkrdTN8I5UmVwxMqHpbyoItbIJOosrpZ4OtuXFEwktLO2P4m4/2SR3KYcE3yiF5K
R/0DUp60W1wqYWB0u5TELlBaenC5oCjdv1bvUOITDylyLulAx17W58IgfrPbQYq6NGXRadtefrVs
5xEX67bDdMcmN/H/jwKZEFH7zsCPKSUfYcsGJufZkj2L2hwx2q8+ENScHk9Z1Wqa5D5/5FyZ4wGN
I13Ajm6QzdhTCe91zMhAoIPmh7TMqEf9VJB2B7fFg3nxrTle3DKQ3l5b9nt8bIQcaaE6mseLnSMo
98/kx4O46OUQJNqRAy8m4g1SWYmyyXj7lNFWq3VSl7JVI6rbJZjWeP9GWdRfF22K/Ss0xsOPMSxZ
OkiY2DhT1MaSzuiTJ+8bNcaAbmQYxyk4z3yw/d27XOr/5w5OcyZL8KOQaiYz0UtMWNyrHM5z8MBk
P5Rlu9iMhs9fh/dYVjsG5Sc7+ixywOvk5GvFicVESt8vUPkOdWx4YUeyO6X2wITytv2RQ8tZV1vw
6t7dXeGY9AevYROMZoanPjTpNlwE99dR5RfpJbC0bD+f/zzyquYpjT4VsDOqfyVJQwMzUhS6BEmt
Ux3jQwBi5JGUSP+bAPZBP9lyhhz0Fvud/KBMASZYtcuUKxni5uw1xe3SP9qaSF/kSBhDNKO88Mhu
teucmDPP7HvljqqKo0DkfMG5dNEzaE9Y1yDWEvn25nGZN9SiL5h8uVDi4c685R/VGKBcBjMuiN2O
uyf04WuHd9yNJZZ4FmfJBMo4+1KQsKy931OhoXSuvd9MgJEspgf7gt+QARA79mvCGrUpcymD+6MK
7sYMCP3KcCKPC15faCQTi7+KXnZ0CcjvXN7FvGJSbJx67sDAJmt7YhMvbJR7TpX4Mj/9OxmqZAmb
bhraoYlerZITcl7YvjKcx5BsGm2qey7CwHh8+FC92wwzG8FdAkDVE4D9kmJ2SqYF+9nwQugWPxHQ
wts5I1B6rAJNUcRurvXea9DvLglICqg/Yg7OciUg+c2qqWXGFNBIZLRy4qhSjnQKFVVa2qi5abxI
sSemM+JjWkeTbm3Vyb7hl1O0AYdNc6ZZuVNpOs34iPcBy/9GAU7sgNj8Huc5RjyLzjrUSrKPjqnK
fXzr6GH61PBEYKbA2Wl+HAjaDuoZzcaH3bSJwfvq9me10TSCdaMDnBBSMQiqn2maS3vLwudzkKO0
Pf/G+xHL+mQAmd6ufCln2swJ6BPuekbAEfCWyClIyoWH/dmnVU6lmnIDmV9pXk7TxMqh5V+wlE60
sI50P2NY5+sMqIwkgEHTipS1GobnWCxFy+U3dNdQXvEoK08S3EITcb+ogjHnnym8SZI496bJaXFN
z5//yO/d9sjePbrpHMO4usJiZLppR1mrwYtZHS7kPeiQ/jZAYzGL8ZsSIFnnnG1UuEnGufsQg4Pw
ZcNia8k8U5hrf+bSYdWzpt1Sorh7YAakRQ4iWWFK7uwFxEca2HK1SH03EUUyijsSrdlRBnMBUNkR
TOzibMdOnUAeQQ0IXbgeIibyj9N6hDzP0NtlX2MyNflIdEyA2znN2NR1HlkihMsPfNQozQJVZrau
BdbxHKKEMni/ZvEszYYpPbWlZnhgAJzTRg5lb25UdJWsjV0B/Ej0hcOEsGPLGCzPd9WP3MKr6QDi
iTinqOjrXTJhyMUKnMaqYhsp2pEJ8vO9r6DbuCm6fnocgBIiYCVjVWKhY9P+ddIkEPp3yKZthhBn
bcHK37UYjdONTKXjcu64DUaTnnR5YK16aTXOx9SnfUSOxw5rpHvWdd9crJ9JfU9SPys99ylcoti+
6iNx4PKgHoT3v7b2YLqNYHixoBLRHnmXSzkONcVIaVjGciYp760Hm4KD6BTVf69QFfEKJPxJJ+dq
GVxIoPUZbjYUlqSIjh9tb9ghrxanLZ+xxt1e3DoSJ9OgHgvL0dfDiKfqaDphO1WBtMXrwCQ2wTPd
kAGc9JOgCZnCS+jWNSlSZ8rPnOT2cXgiw2BsCiSw7GY/ovZmdizXKBhvvL29oFXwGv2Dy11olN/R
vrE1dG9sXZjOmy4Aw7XbsAcNULBUzaxZ9yPKRfVzcJaNNzNBX8D2Dk0NBfKyU9Mw4x3hj/+KlG81
PHxM6TtB+YOnTYTqUsFCyIqCuy4jzA50miUVi+ro3NDnVKavL42xRQ/iH/SFpLZ4SrD4vZZXLAvB
k7KNYu4G/on8FTbil3muRC79LjkIOFn0/lWvyGFyMTuyyBk/mKwiAacUIfiSS9ufBAE4+dQ97bBd
CzMcql0Z295SMMO2hArisWpKr3I3STwuhn4IHrP0Exy8DrsM3DXAWv+wqj7FL9KxQMzkP649ra/n
RafsmJS0lVZz/UHvHRFDWlMGof94mUaDmPUkXaqRsE6gvEtQnEYnc/2wjDYM2jUjQ5rDamVv35/D
SoWmPgS1Sf7oCcmFMXrn5fIkcREP1OZZVZo9kA13tFMQtfj55Jg278//yY9l+Yx4Okk4xq00t9CT
ax0zaqdKqS3OCvkFztUtAVdMya92GgJUzaI4knBlGg0MIxK2IDmKEsaFQM+rNdFZyEKQF6BU4QOz
/5tSyz08p1Q6nJEs6d55XqrFjs/yCM8nm/GC4l7jqFwFqCwyqJFRtjDqy61bYLES4WmUNSO5oHhV
ivMpC5qTFO06E5CXavHlrTCfD8fsvoglg1S4xRe9s7Y9bMFu2VwiYaRlrC7UxEJqPkdMNhe21okQ
4nQq1CV7fuv1RRjC6XF7akAdXNyz+PtsmkI/6MKZFfBjqypd/P0nwVCExnBk2AjwmuDz3OmTL7Ho
TYP31BN0ITzcdF3/0YrhFYWg7VX1Otn9RG2XigB9BZ85UzZ7EUmQy3ZfLpDvRItraOqxeS51b8Ue
uT/8K9ygZfDTxlGTJXZOa6LxOkxNEB7jVREhCGhA3ipmlODhzhyKt02YltXfLK5RqApfnxOpK8zh
QwH7P0zcwB/8uMBHmKd7lUu1JmZld3jE06cJN3csNxDBgIrteO6KGVEMN1wiG9OYmiLWL/3HGdnI
dqJsGcFEiJmhPZJVUQwgwPM4qrBZyMhzZJBLeziy2uOOHW9ja2t68cNd3/gWdaRWFeeUpkVFt9wl
jXVkcImgcsOJbq+QuVaMIGB5gVH+V+zo63UVlgYG/Kwh9FTlRqFxMnhOsQAknJI6hbrwpUgoZTNf
KYYfaI0/duWrOXO26un9BBqY/ThL+jjKi+Y3HUrVjIBctI+DvGz9m4x1h0W9+83D1yntQN65Htc1
zhIEqUSGYOcjhQ/c4RFP5onBnVI3Ubbdz0H8MjYhI4OmNKJsJdqaRqodHQCmTAU68U531UkhgP9U
AiVmgmxQCvAR+S9SRlT/ySMEI80sbhOmLCDGtFDr1QRDZ+Od/MFmUd9bwIpxOBhpU6CKHORBkMQa
tZTWS/zdL7PtUzCwuaWBwnF3wVpmI7sZhXN8mT/rX3Ilz4OwOM7PePRwG2zHlhWL/fQTohUv1ons
fvoMAxoFgaFciBr/aBxPb6wZQkYFQsZr/2BU+x7IF12qHb5IvZxD8xllzalVHVLtehvsF1JKIMei
oSS/hv6GFpawaPeFF2qQ8ISZoLDpdduBD6t2V8+ZRVNiednBADj3Nte2F+vV9ZVXQV8ptCV+WyCk
MXDvGtkWSFgmtMWW8vZAZdm6djYrf+dnaNn+q9gf8Xih5OW1Kd4yETP0+dx7J2rA4uLffBlaklW1
V/oJMlwrsne19g+zLqdEcujEi9AgnMvbGj3m9JViIil7g9LLOsy8h750PNH+wWfKYFzxDc92ln/1
9L37RrqCgcaA8VpjM5lt5bOwyecga+fucizEIMX83c9alSLYK4UhpOG9aem43D/kzV3vCj1c0hiP
7DHkr/PFPM1JpYyDadG94mcaPHbtiPOBVADYaQ4mUbiSuKxeZWUVc1xLk5sjOMFOjWIUtUVzeZlc
wcOJvA7fzRj0pk0y10qcLEQ5uVVzXiEph6UAbSZtdiy0MyyTFCmX26utjqSJV7jIgq7EPiyTSVsK
ht6J5TwuaZhXCQAmfCfLwcRV2Zss8hT5J3tkO6SYDYr+6zKfQrg54D633JRQJkjk4rJ+QSaLrh4O
EKFQNlSEGPMjowLgzOcnnKKc5pVXyAyHatJBnFXr0D1KPmB7N5CikNZV3p9O2G4CnfHfzv2wGKQZ
TrWLav/qdVCoZdWgPxMYIEzpkpF0uhG3JiTS2G1arOrV5x3tMpsh/ITDudpB43aHrZtYh6SEXRA9
hAIHauu7hyHdB6lTKYKWrO8vA5WZBMu6PH5akAG3tBop7DKcXRdDld0qjQUvAKDlrhxcphYraIwG
bKb6C4fInp4YWNyZFcPVt4Gml/uGaY4BsAJ7B3nLNro8IzOBlioRXhGlH//Yt/6RJ5MchR4hy3C+
lcXAosHw4TJNG4m6uCPfhKWz9twopeuVw0ud6AiFB3rYDNohNzIt/yFJxmpFD2NtuJ/4ijtax5Gg
tXf/omDOV37BrUTpUzj+9HoF0ORLol/doE36lclqnJ+BM/fe+3N2/SilV9i24wteo/6OR+3Mbijm
hwVNVVpOHaZE6r9nGn63Mujp3+P/IIBB92x8KhPcrMmgqG7De6gaEh1Ym98Uj/+Y84slPqX57Bd9
eURDc6SCC1hoQE4IsRkengKMR9s9t/b6tRziVxHV0814hbS3slPvDwjle3hlCfX02+QmAsdGYzSI
9NOnZp0pQCbxWcpEuHIUzjD8nwOZahPa9fWa/qSo9xiYTEZBhbyDS9Ko+GbKBENNt5G9KNIctnhI
ZFeb+aMNPaNbXhO0I9mNmryYRg7hDsFh4EsYWeRwVW03bPeBjJ74j2JyBotcNAIqY7adllW3b/tJ
VM4OdAoMhLEQSbWf9K6LT4g4LiZXNSYmISWAA8eVg8c58OSon6szFDSeuEHUdHskg1acw+QYJ6fd
sUcZuGZKEoL4AwwX11I14g1sVU0CIbDUyTgVt5T1XVDJRNHEYOCQw85zDiRQWMujR4RjLzJWecns
HqQhkrv0u7jZ9mlQuMGh9qH6PBA3jXvUjISWiUEeBJrP5C7/znbV1tOg63XgbvCXy+wSI7KDw94v
nmsvdbOfWVQEKQzqVGKaLxiprzlqACys31y5xKYvr0x47SzjDrYmAuz2dnUYtiRzHY3C6SWF9m/h
Nw/VKiRjd9dk6ureqplKm9k5uak7az5mafhhi9coXWPffmCmPhjH1AZBntsJ/a6HHZN7Xgy3xRQ3
fasrowvWUo/Fk4mbysvTMX4sXCkYa4DxYYTFIvNFajA8EiJah8r72Pjgum6pqGgED3BDjpGyRV8A
P48N5uedoHkDKrh9q9gCY5UWHfxj6RmdhMjZ08hObIXLH9ZiW5SX7CvQmHWBsmrNFObXja5n/BSr
798/IelYmc9r0SsrqCAdcXTYxeP6+SseWZnIPYVbOe8471DLBmk52Bh0HY0O4V7jqQmfAJY+IknF
s8cFeXd+apuDrJtU0OZr/0xVo8VPB9hjV0knZXeeC7Pa2DYYEzyaJwl3TSQTjhD9s+eeN7VryEsX
GyBp4LL1oJ8FopN86My3TYkOI2I2AxbCdtwW2IuUsZe48lJOw7ihYUl160b8TwIHx6JG/foIWlcz
Tsf5d77izzWiRLuNKgwacqqUKOnnUOG+qbyeiLt7RtfE0Xwn/rOtnftdlyIi9JS+ZEhwW09VdyQL
X57kx+dtOoWoSD0F5YQ7ieL8mEVLNaObJgpZRxkrJ+Xq3p+13/o73Y+tozNlWgc37N7mUi7zuQc7
4ytmzwvrTgeSWbjAX0GYWDvjbFStTfpEdo8RJyrXB+M5kd4F/d+F8EjKrlwFEp03ywlNeQEoK4aV
EIJg73bQvjGu/ZkCb6IOzpJ0l4orE6aagyBZTjJzKcose8Tu22V+vSnp01iImB59zlAGXEqxJ9s3
DgE5s/B1Rn93Ugai1h19PrEWCqq5gsEfHeUsV2tBmE1iFLIOR0tyirr5Fu/yEqj+6pDKiQF7FXGO
phls65yxtNNmjgsNWl8+o1K9GHEf1HRoKVgeo6nkN+PolQg3drRwRXVSM9vRIWJ3FpojYgL2tmO5
9HuPKJP14jlSQ91TVBBbfPhK8qvQleW0QuQM238lkOFb3PEWgOofl0a/X3nFkUDWN3x0zkMOUkY1
7h4jwC8MYJ8sDfR+fNp4fC8xuyte5pGphKu4hk9yXVNu8OePD5+qlcFBbQQwrbEBdrI2Vap0pOVg
RWo2yIByfNCxxKLmVBHzYoNIdLDUR4Byf6W/alEpuWq/xJregLGqAVvkojxka6dnZArgMU1JchOQ
qgaWS8iViyMdLxA/3M0cYaQJV5ZP+DuT6Vly8YceS0Kpx/hl/35ZH43ryxa4MUJ9WE+2E3tMI0S9
HNXNiN7O/+BEZhLB1BuQB6B/u0t21IUxodbomh4p8nwBH+UhpKCKU5sjA7emEhxGsE0hFWBEQg9v
t9U7zOvE3cVovVboR+WSvlaHBI2hqFPD4PHvBaIplGs6KCLbuC6EqJxUOKuPtmGSbD+zQuIqu7oC
UMbrLXhdlsI53A8shLg17XAAKDFzu9hbD7WcLyIl+/xBXrSqIP5OaGb3FKyu7gkwX8LyrYzpomz8
RHut94eYrwa1bKhpFSa1QwYXJgxpqUbV/LmF9Ggt/QHtlUQK3OL+yfhYZizApixYlJPDwQps2W66
2LaH9rRf2hp7jebZyy66+6Sf6fBFAJAloTw1iR2h9pqkB6JMjpWgl882mSSAAnkPT1sPt5LgB01p
+1dx04ZFA7NzbwA/eHLUoUmvgLfUj7fhhmLWOa1cQZyow6yVQaZLk2bJDRFWys9etUweVhP44vLx
Col9nZmaxtfRuIug3XKCn6tgHVy9eNwxi1tRUkDsF+t0nOvi3oFGCMhxewLctGExwXNvzpjUj5wH
9dXqVEBbhr6VsAanKGJCdvqVzo7b8XrWlbF/kGDicD29X/NGU1UKAfzAxBlI9pZV40h4p9jYiSBH
0kiet95w/v+2M5QIvN0V51wk9HB31nfVlpeg5YsJRv+9u1ONssJFJ+TijFbrQMiV8eDR6V2lgYZc
5hMovbKB+MHrDG/fqrLOM2TvviLVNLSbpp9A7SGf7wfAHPJTYKXk9Wr+KpDwUnAgoGJCoLGRfshJ
CYJD1y8YbA8thEa4TIn+ZKlgtf0n7WQ539KZLcS4NICbwyTqdlRmTuk6ADy9FqadGrpv/imfl/0A
XNFRjIA0qVxGzPE6SU3WDLVXFgHQ2I49TJypyRrccRu2h52nadVQkmTt0+OKRZXZZbpmBAUO7Spy
ngCJubiXUkESzy7pJ4PgcugDlZKhT49naPlTmYbgg0XERPrjdvgeqE19xAbM0EP8aDdQycqiQ9Pn
anHMawu/iPGpgsGfRaJoTYJIwICQsQ6uEsPBy6LUpsIsIaG7lO0VRxLUVk4m/KGoI0YY2FAxV5AM
l4AbjeZ9qAzd5+NHvzMZYWCRYUsprXhF0dLzUCIK/Dytgsem8W4iqp+6L1HZZ/ex8aL188XBUJcF
uq1z8VEEFu35NB9j80W68lQt59ObsjSO1tl3CrOb3j32rjCDqjTyUQh2uK+D0/iuWa2pi2SgZZsp
7oXnfnBSRyyNoLVRtj/3rzTnEkqn6D6O5jis3mvCJNHQ+1kIjNPcXLyoZ9zv31vZZDPAtb7VlXlJ
kScoT+q0bSspm1sXnyN33AOzxUSuDjmOfPHwac3/CM2CrtXnJv2T/5qkfYVZet9ht7F5Co4TKA2W
6txTwtEpY0zH8CsvfSxE655l7FoQC1JTkqlczU86DnfX/BK2cH0tmv6Pn7fTMRMiKKrmt8lqgT7W
3BSXX3BYe+03AHRzSUkF7cucjzDXKfcUWykHrCaMq+VnOqxIYwUmQK5OBSwg+Fdto93leOw79CAz
s5ZHldm1Mwaj5lLnGAGNV5+14E2lpN1VIIQZ8jIFxPOCEmxgxGMHFs3EFA6IGqdmYmZmjgRMkbwJ
a9b31JBC5UzGkKo6/N6kJ/7VwilsQ+LACP+BXQntOOS8gjOF20VPqyhTD7bLdSlyWusvONO/jgSW
A+QS/xTwxt/KAHau8RZjzWKAzvbyJRUOWkFkgO4j87djcBsh1D6pOVWGK/hj142THHA7D9vnsY3m
vkf7Qx+Xpn/ALOJX5VTDgk9pcMtyUDpQFwk4Fv5P8f2KiorhGV5PzSS1OciGQ7SUFUoFkrAafgUC
qQuQK9PKVR5x2yltc4cY/f4f5awx7To9CcVfXupsZ+dNsYyUiUU5NvG7bd3SuGOaIYQRa9xwr7FW
Aoosp2hqrhy7QIIRQpi+tmdn3cDI8TXYjeBHGqf5EHyGFZ6xRDVIyyxYFSD0DyAgvyNbi262cTmm
ih7eYuqkeZfvK1nIcnylA2E3STZ5NKCyLFGPaQ4BwkoD4dT3qWMn6n2rSFO5lvd9ctc93Zj2mN+1
O1SedIBQeNQrNmvK5+yN1SA+GBdv+Rom0YxXtboA7kVWa8tmft4jtTCznIXtAs0T81OBeEVP2WB1
XMG1GKdBfw9aSm/nQtutlakC6KNnqQDCP6Ro05RBAWk7dty1bH7/lpY/Ad7mXP/h4jq4JGSLVt/o
ynA/pGqcTfZqIw5qRznjqCeg6qaYIRimtTmWD4lV94h8jPCkNZNvICLDpzn7PFvhkmnryT/nGDEx
75H5c4MhSIaEqxZHq5SP7ueS6O7V+PZcsYbBG0aQE1qR20NyTiarMnDJ1WWO70N8edy+getmOS5k
VIMdMqqrJyMHG8kvx3gGoYfWK1MdvdxI3w8M77LKkMWELZZnDzNtuz7CyFaxH7p5ZWZJhfR9N19J
AzG2a748K/RZ2AYAGbGRdJ66OxGNuD7HO3oRK5v/jLT7iRL/c6uK/m5V0MknuERt10C2S4H8iw0h
3xsVtpnH8f/JLQBu6MfpWwz2FSXe+L8Dc2KBnKTtwaMf6ZKL9DePF3/tD7BDVr62Unl+fUyEXJoX
BmZrhIP5PFxSGzUEVRMP9C1Ny379Kp4OBkRNncKj4e77R5h7XX8OlgEXG2cdr6O3VLEXO1PenHrV
xFOOTn0Z2apLzHjENU4m1FEKK4ua8s//tpvYluRj/0E7CmL5RzYwl7F7JKtd1VQ7KXKpFM1csJWV
JAyifG+qhSRhOzYxFsCixHu8KPSmvKZW96njHdI7ncsE/ltHuvpSIbdHBtuqASHMTAyAegStgL3D
dSPxgwvt1XqeXXwMPn3awPVFBbsOubOUsJ3Ld/poYgyWoOM4/G7a6MFNIVdd1aV8Vs2tjMb2uqC4
UQshvG1ezotddOaB3whVJ/OKBStrfhw8XfcXWZ0Rf+XK7npz12/I79AnPgfRVu+3IAQwHRvc7qnk
8TkgSG7BxYRaB9TK7tBZdSqI6s5f1ujirtbg/3x+5DyF+qAzxSVlct22Xh/ZewZ3fIkN2b6uq/xo
PCPOHBGk6h/YD9Von9lULAtv+IP4yS7JqTIGScR5mlFo1ARiYYmo0pGrSMyIhuql1/F1jkGP69Ez
xnMQWAuTUwIH2z2RG8t3b+gq6dTEA9W/FGB/mOzcVnCCPT7jD5jkVNYie8dVCkFeBuguqkc+OBgP
11WkzX1vRQwgfqT+/cvkUEqCljbJRPnsT0bpgchgMvpOVwjs5F08178pVVb8lx7+dmzzl9VMaIwI
8a383Fn9mcaY2rEErQb1n3N/wD1OAITAlUAeiX+sXlY3fQik6l9kCWKn0p2FFrZzmDE5+k8BIwb+
lS03SiXDJSthwEwvabATY3Ze/U6Ci/IZ5I7a8JZTKeADmCR4RA+tljm550zVFZI9FWHBbWACHu/L
acayWdAt3zkAZhn8OXoBJaKIqKqHi3DPXAMZc7iQjjx16Xw4d47Qc5EKu7SltVQnRsvLO4wMImuw
PEVJ1SKl8RvBBDccD3ipWLqU/wnal//Pcf7md7kr0fnU9otf6xprYn7hQG0v6Mzrr6bexB38Rr8+
Zgk+BdlLHN/9eC2rqGBpW4q1ao0jF+/wkPaouMCLwzPo/UPBLotWoTauVa1yq6BV+1EHk3aXj3Qh
sNIglz/O/3yuqCGkLzQIv8e3XycL92Hj4rOaXlOf/ZMErwhvI/nHE1DF/JgxxTNHs087lau9GUom
7CTda1N6XPZasWHofKe8JAhLeFKGJnT34aQQO/Q7v9ZYa09x1AzAKB9eBVqw22VmluJbQXBytV8/
cmnqR/1lLFJRkkO8mAsIG54JEYmww5cJZIeG+Hp7GKvgK4WP0t01PFIXhjYnEWfaNZtllcy1y9jz
xIUKpi6F9H3Hb0QV8YQZ0Nu4M0FQxNyZvvW8wZhLerTa/QlkJhj1CIYpm0X71NxGgGdRno2JlCFY
wlGwn+M9R2WcO6UJP8RxMORkhLJDmAdtx8N1AxT7pXFEkQfK7lWK14FMyveZWkj69cE0zDA1lxia
s3+Sa+6qN29HqizVLn5zlYp3yJU/f4T3Tyg+r52m1G3lkXGlrIFmqAb8jKexzEwfLDUz3NFjUiYT
uMVA8UTdnO1YQuUpSxU3UHYhl0U8VwT7tMauhx5dsxcGE3Zn+J4KHG2aNVDjYOp3YGuyQrqQkTx0
ZvYyuvyFpW4EK9onZgTMdqFro6K+EHdzYciNuHU3MOXYd4OIWEqWExjIYvjTEHkgbqQIRywlzNLb
ovCSQU9jEIUaAoeLq6Inxn+9tHlFCUB+OosajS7W6q6MGK7eXx2S2y8jc1LWJRcK7OkoN9RACLi1
7dUpIiQ3N53HLKTCgxZM53XlTkR5XQguRfV0qAvl2997I/BJ5X+I1CqGmRFWx7AjUpdutUEtJnyq
VuQL7LMpADDKWKrXFVmMwcELmSvmR6WbEt2X0Kj2SDaI+abFPofQdJFel1uIHu8NDGj+XZzoVeV4
sT9+VOy99JauFCp+RK4rr5V7vE+WgSh4Cp2C12swYeMnpmkiTP4UtWJoRVHjKKHivNsi7DUM9LJM
gHL/0kXeL8glXgLQu53w6z8hhg7vedix+kMGUMT7BNzh0Zg6O0aii8mJHdEqQPj2QfKTVq6t0iwY
gr6wimjp5/g4KALopWdXA/wQp/UVvVWX13bRxYMRFP1wiegJOPFqLWwpeWTRhWSitXxfxpKmzei9
0M7iYEr7JsRaOIXcq+F6ijSj9sgOCtRukMwm/C6WuWH+mN9EPEVkUOANA266eNBAbxxuaw7f183C
pQs2P/B+ORUeNWzrz05cLQSxdYhKwo7xFDcDmdW8nCytIbeC0WwShS6WbGd0/RT0dItobyyNtlqA
yI0QCVzLVxwH00EAn8kDyPxwR2iJu2qjzd7mhZTVaYIq0mUfsPviJ/5JhnLu4Cdoe6N2ojCas1pg
D8tEYsls7XJ66Afi5VLaSatw9PNN+nfkAZEXo34XndcUr9OnLC5AGiIqxdwgd/ytoH0cku9Me8vz
bV66apVizIPsww/mqqUcS7dD0oa8MRLwuNByFZwRp9cYOkas5Yz3F70JU1kLFg+Na4vESiZKuhXo
Ek4TG+TMy1xAJHPXwPHvnho41ycTHPDD8kMDy1dQ6D4cF+cGQFGsjNAAnq8vSXiowWi6p7+UJIyI
/rRTGQFKTF2t8aH/vsfto9KGTCB1Z1sIuda/SFM4mL9LhDqsKCQTxoAr65uyHeqR+UWAkIPSx9Y7
hN6e889mvlGm8srqo0dyg0/jYjr3hkCvEr3xJRayzY8mnJix6TJDcYbAHgagxCB8JCWoxGaTyCbJ
fKkSPAhaKmKcehLE5ZjoivKJyOiRB5ODjWPoOsSDd4FI8G4eKdLAM5HKQunmxjvF29qawHyZBVhy
daiqQr/dcm4QnFQ/pJDrYyhp9mB0bO+NCbrnbZcb8DMzk7LilTtVWxnne/rpXOA1SuxW52erGj//
7lPn5ME5PpxIldXDTqFgOGMxHkAwY0IgpUAv7pHAvDZnX5WxrlxVPjWMEKZKkaLDvTFrqH10sUOS
j3733CchvW+0zSn9mNBmKEt7V6kXRnaUBxkqG0FeTadR64mOeiFYZtFm/xvjz7RzFrvGNZdYc2OO
Gt+2DJ1qKG/r5whBvdKfMuHL+yOzOxEumY5UABnMwRZ+FQJ8J14Uzm668q7UHYpvmRHXn8OEco+Q
dsw8NsDHLC5+4q7QrHge57toJ13GsnerRIZznxm5l69b+E4yi3IttUapDRvqxrBAXEDOGul+v3fH
1r6i6DkIngxbBYsuY3jk0AE/iuRIsk2EM0TqSDuFsANg525/PUEhrkCq6vTTnHQAiMQFVwOqNaA9
5ZeneitDvKrw5Inl53aYVe1p6HznC7nXznQ2JMW9H2yyLBM9+CfOzLMVoZGZWfN42EpysKBUzkNy
6FrU9pM8VL73OOsWfRDIA1fOI8HWoIT6Dih7gKAKLocjjegpjFE+r0veqxsA9gxGq++mx+MpNzy1
4kVo1cWw6XfII4J9dmvwqoYd+aTDyKZZNOe88eosN7ZqYuHf4BztH5qnauQB+4lJ3V5F36/NJfou
kuyfFcDeGtAqhHzR4vSHBEy4eu+QL/7hJmKQrrQNVumMQcgIpr8/v16QDmy3eDD0UudqI+vPim/8
zdMfEHxLqD4dmz4KaSv1bG2d5+ykyWhtOrcUBTBOtNi540Wrm9920aSCyuVu1vWvVzzqMkP91ahd
04MC5Q69XCg41RHiAIQcHBK32CQ/j0W8heJToV0z/BPihY5imJnmPGrMddPf+NBZyl8yB8dO0w2+
wt+gE+RIHEvz+51D2+Wgf7EErsEaDbZRIvsOdErFz5MWz1mYoRvdV36sgNo0THdHgUHwdwgfrd+y
/U0uiID+q+xaROk0Y1pMboGdKeByiox9thwKGN2sl6TFyhsXfqHyevEIZVxB3+Ev0MUUO0VJNBKX
NAh62AH6qMUNXqmAVglkyTN8uIwV7ciGzSvx5WRMjHMz6YxrAsXEAfC/hVvLzIanJwnvMISc5BMQ
o8xB7uwp4rJ6/yvAjT5sVwXkhpYbZYjeTQJN2sKz+kA8heCiiIN1SetDBbVbuSS+Cthe5J23E2sf
jXSPUWvTyAWr5v/483HKkx6VLrkQVjl7abtvksaIsD0Jv0zY3b9iZhttS6aGr7jXQpyrPaWQSyZM
MF4WZ3O6AOi2Iu6QS6GsMVXBHoH9cXckZ7xs6Q41NdVBsL4bPfGEaZxUDrLenJ7BT+05RIsyRSvv
MP5kKoqavX251gvSP4cxrFrkBWzPmS3ZlVFhsQZ8iX0EcyOh2D+D1UrgghgxG7qMIU9wmyKmn3g5
GxHCFIN5LDcdHtJMwX5Kr2W7D9RdjWrQsXfmrL+Dt7+H3U2VPsb9jEkIIpEwZq2Ap0AEvCnsfgD5
6kG3CoV0fCGf2EIXTQKiCItf5UMcvm6sHkkVIng0pi3X+gV8wIDKxLbeHjaTB57QKluufQz83no5
LIOBVeJ/+oqBQNw2IMIAn3IqFvur5eZvw/ZFN8efujYRvsBy1PsPkiZZVUKP5FlwjneTgAaVZHfm
lHonPzfc5gE8r7R4mFThNoZJaWw8Dym5wzRYHrr9EKHu8QP5clJMyRfVHrOzYghJrWe50aDCb10T
t5fTMWA38/QrsjcLSDqgG04ujMpJFw4NEWY1mdMWClP/0lPWHuyIvvJ2tSFJjuQTKRcHSaB397hT
ztIAYx/nIZxBxpoMf/GLBcOzUnmJNuR7YWArGpl3fsVuEdBDjSgph2tx8ZnvCLwmx9+siGl5sysV
z3NCCeI4JKJYuAnBwHVCUoIoi9TXMmNdh+4lpdt7nYLxfAHihMuoPfw2juXBAr+qnzeYsyS3xsfT
ORTVPy11ZeHlhzDRMa5/dW0OLT8XHAfuc6mYFXTcWDwrFHP25R9ZNJ2lEqUABqDI+XgnILBSvA5I
Yd/bk95RHgLdK36BTgxLzwggeyBMTidhxYMuw6z2GK/aA6plm2GJJ8V8aCt3LcrK7DzXTmk7mupz
gzDGo6t1rdbiDBdzPdvue8usHZH89HPnIu+K69UU1Azp772zD17s5WoY6tTN0WjX7iHcyqjaskXc
WYvw3UWw4myRMY8vn26qKCV47IEJC53eTaEL32nNqS4HUaJFUw26mnTXiyQzLMHxjVIdFHxGgoWQ
qxhbUDE3lgx0djFcuFrg6LlaMy0XBwtbnh8EsLamCJ5VwFv1qEDsv6pt+l190Ihul/5teMITbqmP
BkxVhz60piy51QwX62gR82pRUEFGMRg5g40Cowx8EX4dDR4QCLjklFE2SpJyX1POlyAn+s7E0L6y
lQA0b0wRIflMd3tHo3kJSY+Aoryv5u3T+1YVDgU3duCS/Jn1QX6aDnfIKKLS7SOFvOoT4gPftrmE
2KZ6FR8/lsSeZzSvP/Da8ClN4eVjHws95R4C1nPhhNrwj4PLjG8+Kj2nlwkkxoaTYBY2FzExibwj
3aEDjrGxZB273JoERWLDBjyGvT7JNdUvG7t39denHvxrzu+TNS+ifZMugTQIN08EknIrkc9iRkON
KWA1wv7+lGvawKL+oVmTTRdTb5eWOoXkTogngs7HA4oA5lw9SaKPJfuEv2QnywThpi5XGQFn2/7L
5ZPMmJgYpJ4yAcehCmLrv0dzZZJHIoKRQN6MNo2N0sndFeGHOeektWr68UQYasgw66WLoc70q3rH
h/nreVgArKwRmQ1bmqGJOEN6BVU4fPHFb+a97Y8ZMV1+yzkByNNjCDrKqDzLLYA/WbbduvblxK9f
FU5LZJ3qcbUdvTUE8vJ6chdU1gWdCPYkYgNvg9E/y0rdqHfNQddZbvlXiZN1CxBtmA1VrOccteMn
eDH1b/8CI28k+lduAlDLEtCPhuYQfjZhpD5DoRXpfPfwL5vL/XuKWGtD+A1BaSI0t7z6NxXiNSvs
jKXvCzGb8x3wPJJ3d0UYOlSxSrm+jMwwJOwODjVg7Gqa617LogMnT0WtKGma5V5RRY1c0HEQL+lT
fDgl2w8ShigiNt6EgvUB/PzYCY9oFu5nrOoINfTszwjEoGtg1t9zMtb1pOrf58ZINxufBOubdU3L
KI0PlKwS6hGfH7lv8AMu6jAsE2wLCA5O2XPmSuWvjB3eNmTK7UvUKrLHn5HVwbJeKp23lABCzNIX
y1UY6KTN+RsFPnxxukkhRkXEewtAggIq/nr+GVGNKhZIo/UxRDAcDBVvzpdsohX9OjwnPwnKW8o8
Yd7jHwEpbTups/AyhGsfCZryKUIuKDIHzr/U+5sQ014mPt+04YI78GXO/Kvr5Tzju6JOrIAofN+G
IIc3RdIFRulhA8rmDbEosrZmfkGQRkf8wia3fblL207zznFYN73T+mBk8zdy8UbSeDrAfsFSblJW
rgg/iEVytoZ7m9mcvv1stbOVyXnCwv/UaYiJkrkMT3hW87cmAOxEGiFJKQoQC8yeBuUpbbwBSSNW
FHd/yXJJWekJnMMmiIKzJu2EPy3H/x13GBasHTOYLfU91GrSxuARwPA7Hb5KtLaviGTgINHuXDdQ
qEEjEA2HINT3RdSYqs4bgZv481ziPvv77U69Tejc1BDy5kjZ7ih/ZQYrOloG48sSG630Zgsuz4pP
QG7E0A+zhmrbnwA1/4EYmp2Ep3w3Hhb9UihdbloKlIoOdsAQrRNWbZ5Wdk6YifWCBRtfA/f03wJR
biDtpBSzG79IdhvR+40xa5aHiB6dXcGtwg4OfpGN3sicb2W18ZkCMPZQM5GYCUOXAsJtuadfCbt4
+rLGwZj43vKnFMqsha7MLjKL5pTstvgaK/2fnTu6AuLX1h6yvkyXhn7y7B025rXDHWEpdPQ1TfXo
2cKjySLxhrk9V1xitiZC2iTvisoi/c5KH5/tFn5nqxMXpAl/VCXK1TagnG1fnNakO6gVM3u3BDoa
T5dTTc0hh62hotPQDG0O1wgeKcVWPTEbghJ/CpsbhXPW5i5IjZ/pwos92TcL3twY4g6oMCnKHn6W
H4ctettpQ0KkH0voTrEZyRg0SGGeESHG/GT/2ruKXQcLCtEFyO+L/3cWIbEwOS0NpCze9B+Mj3i9
abXn7C8gi9cO0W4u8fJSrBq4seUJp7iokT1MBLlmCzxpiArXVte1LXVy13+2gsBZMr7T/lO3lPum
r8mHKOrO9A/V+3RnmTOv6T+8zrF3e3rp1xArvgl+NRs8082Q8Tvg4ck/G8MXDP0FWM0nH0c6cWI+
KTGwaTLknyEUmXzt8AFQlDU470Z3O5s9h/SJLOkNsBtNTxuJ6cJnUCBKUptJIjIk30B8/i/Dqs3+
Pd8kUpsqwkDMmpX9zIV0vf55lBAurgFt7YtUA8NOH77naphk5kmsVyoiC4bpI7QAvk3v2nNSWJ5b
DnaAQVJExnHY6jJc7AEtNe+84LOr1qIiI/50PMCc3UUh7m+9bMG0E3i0X8xljW7Z6UqP8DV8WFEp
XWMSeClGSvL0abS6srhHIiNw4fxzh0wKTsb4vhQMeV15DPawGdSc15R0ijBDkK/cdK8qRJtj7IZA
76ITNbhBlquSJlq++LdBkIlIgu+kKWTBKtb+d6BwXV1+39d14b/faQYv5OIU9lxmMLsSKgv0irPi
SO8WKbGAyKQgPRnNQLD2tzFdm/TltARqwM3TnhNGPCyuTE30NlImR5nbbmIGn1DOYIUV5j0IzMI8
LvCBqb4+cN2U4c1YpWgb4FWtbXvYo4G8BNNhqcZpNJYRFekShNNbVprJj4owK/DIHWGPbBiOXBHe
CGAuGEsmesANv3CdHEeNMIYLp6/vBK0356v9CTGN5HZjilIX3Expdu8WTTCP4c+qNYXnIf+wqMt3
4q36rb24vAfcN8vlCIZbZEVb9q7eKocOFkErRlhxzFJ7cgKwXeDWuj7aCA4RAA7r5fAmKZosU/LK
QswL/vWmJ5WMVS7rOB0GdiaXlM1WlKEFc5rcAElrXN2Y1dpCby2nP/qWlrHMuV26Da5ecgn84hG2
VQQd2+FdbMCuUjkZZyhbBsl034HkYviaItaA/gcB9HeAvvwKnHr/h6geCR/0I1CECqrquV9WEBSM
jxJI9Bz6ECYNirIVHQUTgDkGJQpzbs1KTH/VFD3tMEUp/+yLFiR+cP+3NCXXhpNrBjeOzabUzYvr
WpLkgMGW4QGpMMQhipjgItYzMYdNOOYjfiSnfsehDinIxdHdOA9IWCRgxvzcdFrAc3wyAongX8BH
mUMi3lVTlngNb3h5TeI3s5TwPglZZMsowKgC84q7ZSKspREDfRSHxi2DethLbbFdVEKr4WnkvdsR
eJrvI1ovX0bhpWmdnJZpNFFIk8W56xX0NPExCRMjga83fuPP5WuY2+3HBVvmiYDJ5+tP6CZ3Hghd
Mo1CmzhDrUR9B9XX25umhV6pJ79S/M1t7nUVpJ6qMVVravLtM9HWg1cy+X2nBbw/ao24No3nSwwo
MDyWgbLvjwnpsmVyxPTaApjCDWhn5UP2I95lA8gLTURGuWc4tvatQaQWsVodlJsdMwDZsKciat3b
pYDduRTn/d90p0SBDeGGsJHrtbDQvmlvH4Jgid9EufcpGLOI4dmeNn8ZxWbehC/2Hem8emMsVzh3
bpKtEvMXEXr8wqOKFFG6VsFE0RqjOvn31QMSpJ0Kyec9Ns3BYWypb20fDZcdQ7BPwld7DY7Wrj5t
oFAjY87/jZVmCzFwIfWXuppI/m+2Aunze5apHO0FhCPqUwM+BJROu3W5v2FtCai+CN6jMIlbMJxx
eVLuvFAtA1BSFLhN7SPrlo0hRQbeFSONa67ikEWM7FlubofOZWIUE1ONQZkcnQTH01OrnbZRGMBi
KJWEVmV6Nf0o3TPF0+zTgE223NYEtuW+diVB7e0iAsPBt8JF7G7XN32lnODwBU4KpDxaR5XAQIi7
ylx67ViHhcoVkI8KlzFydWZYAV4nl4AKNXHQFevWDzIPrKmXFOdZRe0W5kLkT2kgpxfHHGzbswzN
c1zUxv2FftteMeYCEotZTcHsJhd+xv8GiFweQwPRfthfMFHsmc53oAsEmHoughV4+HpsJ/7svjx4
EXzAKVYdutNm5RHBuPmelMv71eIGQAYdH+6aZkXGpXa3K6nE+rPp7qhmQziZxGpxtjekdbT6IA5G
xniLmb5HUlg13PxBu57UZ7Cv8d2CD0RpPjqX5ybdkoqGbfs1Bih4OTTTgVMDA/ipLrFhlkNapGSb
h0n2yM5JMTdQvVwgnBSPv7XjKPDEsjz1xzNBUiG/urD2IXcqQO9ut8M1Od4XVJHZ7tKyvHwNvPqU
XzIomYDmknoYjyIm6Upo0tMjWBanQHzdDNkUJKysHh0RI6L+5il9EkaONaftEM2Gq9v8ZM5mRrP2
OgBssha1yGZWLls6snWj+jJ6AawdaWnOV9iGQcd/GLKZP2NREgy6sbgFRs1Pdc9KzbZbhXYlVpZ5
kNtsJYHY4lLKtCLMpK4NKbCg/wLusI4pcekYmF1SlR/ArP+dbTpYvYAJVUp29+xwWtmTcW7kWZNU
BAvx4k6NKIWTqInTM45io+Jm7oOjhwXidozfNbWEdHENnngBVWC3CY50ConuJN1J5DbmCRQaxZle
FkD/wXHHY8plVa9Z51t4QMDajVvwI2V5BagLbJMqPAu06X8cDuqa57KdIybfd+ZQudewYgjFsKP4
vBriacBa/7txFDDc/sr6HLBQfypJtjbSJokca9DZZcxJ78xEoTsjm7QI02GvegvLgkKbb00j8V01
jEi7a+IP5QZ1hxe+81YDl0EDTdkl2SbiyxMdN42OGw/apkfzU1Fc97QuKyTCVGKrvwLVqzYar54j
KQ5r0Xvbb6VzSpS71TmdEwMwh2jKpQxrjGROtFGt+VFUfQhm3ass5tQOMGFV9UlN1Exqj/JyLfMG
A06fV79ZoSN4eDO7dJNZT73AoMVFGCEDQhDA7DBJie7avuNiLDurKxV0ShU0Mvz5BT8DxcJEeuPo
u6mr2BjnjuOlsnpv7IPQOCIg2Y2EkMMFl4D251Bu3uvSKjSsFPXVUXzyId7oVGu6xKUOdt/nNC1s
hRDQdmKWGUrgiccYD2K66cZoXGX50wdphmcsaWn+6NQyM+612B3Bbpjdg+dkHDWD7rC2P6T9W9OK
GStVX5hsvsC1OInSj+o5YOcn5D6oQLMn1io/+xOsYg6a9LE3IuaFrjfVIMTBfFEU4PROE/5tK50U
FBVet2TjNNjIKEg6QIaYSmER/6vA/BoYtXrRNJCucUNalFvNDIpdrC+ICFa732ijhQOzVXvEf5VW
P5bahp8TlcppR5Cjot5fpizWVp3SqBp287RbH+f1YvILLilugXJLJn/Bfet1PflDlYK3kFURofac
o1qk4HjEMrGwOH7jHPOQ108LHBPcpW9j4CjFIRLbu+SF5lATDOu3LVzSoU7hTJHjLw50ye/nL9Io
jDo3QKZtLrgZl20DT+KCzmhfXqI8EB80/PeNOMJ83I6XsGxi7kxfGxJYnAIL/0lkypcHA0a/ZAz5
1qz8FJEnCWPwmebEjfxohD+6+9DuQa//4r2fsCVE3X7lM5vyQtk7do/BhY0eF7pZHX9Op7rwGBmY
ig54oeVnx64Hdk1fDmrGLZGIOYL4+GOIy0MoLtvAoHzBDkJesTX4nATRlhenmqWL4aJ2BgQstrF2
FeD5Ul6N7zmliuz7vOgIRvY4Qv9um+gnMZSKPvqQma1afiBtXhV8FC4mqStNqnuOxAruByhGhCrV
sc4ANF6EldPS/1C0TbGueB5uISrjLWsdTD+WJIXp7cX4h6PutRIaTxq/5t0OSuSPX8Co4Ps5Nzi0
RTsciPVFRPuU4qjK3dGfKlzZIyKMppwzQLm1eTcLS4wyxWgM5/878feSwL3Pyij12pwTFpxzPDEs
8Wx0osBiisT2LqSL5UzR6YftkhyY0G+e9gg6HjOPG+TAZ1iM1ER3LEQY/YvgdC82rcrZT2LdSIJu
Yvec7QU4kqN7FAb/AyPT9Kd8pylUTPwH0Cm1FPtd4XbuyAwqJrQqB9Sxi647A807RZl9Xn9A+mYr
ODyf8HmwlG7vm+aUNBR9B8hRXU2Khln+skFsJma7RNxJuqJxVDWWA9ZEUt2YPHorlNOLc9qVEN8Y
aycYxpRyWoD+WV2uolQJGBlhw1emHz7CedLIGgL+cx9DAhIlDFWJriayIfbxJzqj+Gvi4ZzjX8ye
PEtmei7Je9q28AJbkPTpi3RRqZBu/h/eoGOSLl27e2bFg8/SFBak7fuEPE0WI99eIo/ysx9Ypd6h
06H8mpRAjyVc/eszbaJQWneZz6nxa4ouhovi9dziS/ecfoXAkE5PL5haT6PfgWb1MatTOBrELhZe
ZiTdGCciXF1Gkt22FmSJxRDsUrsiXMPpCzlBiwWP78vTOqp+UbJbsWcQMEOyO9Ht7VBcPSFnF02b
NKMArOuIKbeF4G+RKftWqb66o1oU0mBRymwVKS0rdFjnM1iy51s/78tHfxo73EelosdNABi+0UUc
JmyYIa+bvMGlIJKhzJhzV+PXdx5dTrYyF6XS0eb2Ycr+SADu+hCybhLfSI/HYRW3kp3g9icHLC9c
Gg5vEIWwXMQnGcuGtCBaPO+xdNqsk5dYpXi/1iGhkD/R9apQ5T0M6eQAVGl3S8RB63zXyje+FYkP
fgyrmSovAXYL/cObmHMuNg048pU3ZAwOI4sgs50w2paaF0xuLZTfNJa7rivZ+tyjcyAr/01q5avr
FZIwuK3D4TgfbdgdkepVhaO2izRD6iOydvgfrKiJbujPULoqDiZ9ZB2eqW6F3vP8rrFRm8pQtr1F
h0kOH24R/Lpt2J6P4/U6xXTcQ6Iose4ePRNrQjbfltBnIdYjLbouSTIrjpVqrwOtqEZ4t73r9RTm
0l5BplTvI2HN4SIdMpyoE96V7cMtJbz7mREdWrWMl4YjpaDTRabkjKFSb81+GMo0SSo4X5AM6YU4
aFXiGm1V8ynBvXY0CrcXUPTODsxw00B7fjlxQ6BGXP4JI9HuQ7GbY1emkl1wtdIHYhNVo84xLfqh
SRsG04FctQrBYjqrYQZHVTBoowWZAfbTFr0T6ja3KsLFbHiIPlco+fJsmxw82+4SkxHu9hC0VVAS
L/lCVqbrMMa+jaAdIykS4dLJ7zpO+2jhXky8FD7djFwx+NPkU3Ftk+otWCxkXPX0GNPTVZBaUStg
eDeZkofzMbEujOsPHBeh3nDUtSxT/K4QW2A9RH4wuOCMmJ4jiIgIzfBMjdMHvX6qa+pTKGh0u7+m
cIH5KBgXsX/jF4lvfM6Ky8imaeBlTVlcOi9XRexqRDHvhneUCjf5tVzOBE8Jf57Yfm9ZXBm5ISCB
nr4tTLmHONiyNv32xsXavoZmWQ01o7qoQvvkrQt6gDsHRz3UppqDYLwy/2epZtG5pUDX/IeFB2RK
bdE8gvm/2BIxFVs7l9VIBUy7g0NGG4GjPDzyYmJfFuA88ncWxN3A9SbzlcQSQ4ppdJwfY5GFtPWd
6FTC0F6OmBXYJJ7XKR+J0A+OQiqhHq2diyRIP10Gd0B5EiLRIZ7iorrvcoXXD+jjdqXL82Q/gBW4
aU1Db9BSdExTqv5hq1Sg3Ad9YLh5+PQOCJJ2WtQe0pN0BSoXRGotHAX/hcUSFIQ6lYDOyQx9R7O8
rrtcsTgowd6o70fflLhz/fl98sDX/7UNS4bLVEDD17NTrIKIR92rWnShrDfOlehpoENnjO3ablQR
DVCBc0jTxFP+INfR5MUwA6afDrc40LTQSK5xC9UFeBfePjWojjwPpQFtYGl4chvN8fxTlrvLjHxr
qxRk0QhLOzHG5u8QjNITexyW+Eq7n3RIzJUSElnV5vc0wC3jmetrpaopueSFseTryE1c9unvj2yk
tm0IGie6b4l5X1X6GOQBLw6h0sznI/IP5gdCRow+HJGpbJVobt4JdUNjPtB+f5EiFJ+J9BCzPReQ
5CpunbFxoPQ48jTgCvZvKlLN88EVMLyBl45lXjUoJxM0P+Up8jP2l0VBT8ij/KGKudTS6O3/snP3
NeGdBudFZMg7cR9zs78H0G/T7EBoqZB8kSBBRZ8Aq009L69ZGXXmkqTX5EbLgkaLYtY5aId5TDBE
WSfFBj6aQgSW6yNkp45S6jR53/7bN2tq3xHOderKoCUCtwfpYuzBmoFwRc3vivROJmDdI4gCfZCr
REG3KCd7v9fAZ2O1S4SgPnP/RaacoQj7ZmfbkDpHs2+pM7IqTk5hPMKCcwNZtw86a9dg4PB6GCaW
T+n5ZRO44FJjT4XOnvUC855asYp9gFpeQhMaDGKB4HDFT/Whfwj1n1DxANvH7T0ZSuS+0nRsiAL9
2uXsGOaKUCi5pbE7huP31LNZzFBIp8fwyL0wnt+dKwBdIJB2qGFluuQXpdRyKWuUmHY77VgODOIP
4TgQpLfnajObpsf0aLetGMqio5vbkioxY5p8K1Z/0JTHbo2WJydSsnsYLv6ioGPMxugDYtcRiwqP
nVyHxEWYAONLrMZKrI3WUkgCPeTZl1sOB0K0yu94mW2Z5/CLYGMyHLWKd/uu9dx8iWrgCjMRxWfK
7GegyZIWEmn2rygDOe16/0c8cGy1EPRE+ptiszzqGiMXsSD6mrr7D2iBqCe2POjjbc/2z80W/PXx
+ovk2nOPAuGstFkmJ5oz0YX94I8hlLdkMbkr6TkGebHBZptYMMUa8tLHn08qdQU71QL1ZwByQcmj
IhnTQUuOgqmh8DaJ8ov10vhb7/ClPLRwfG879XV39QI1ed30fh/7kIecWxerXurmlRCdk17TcB/V
DBVwtGnQNUD4wP0DvtYvYn4sG4vmRpAeBonRXecsbAAPn+FyeIRkGPvSP+//W+lxD+LI2hFTIvgv
UtV/0H2JpBs9jSBR/aa6OJhOh/JWaYg0gmLtU9+3RVhapZXWnDK+kCsOMoXohYpSaeHNcxAL0glW
/HpOo/NIqCgYz5AckJvFfj7nWp0m3Lk8tz0bS77rcQqWR8QhUzvAojFed7MQE7A5ozX8HdJ1GKWM
SYu6ckBvk7r5jdAuUE9VX10Iw2lT4RW2dcAMkCeyVbehrOEQ2jTf150kK/cuOuYMlLB9o8XmQbpp
YqfJFKiFgJ8bVj90UnIplMT8qtQyHdwBBebE7tmv4sSbs8Dk6NVnx3FALr6jrbyQm7yMF3K8qXF7
7r5JK1azfUJ4LB15u8K5is2TzXTzmfDFYEZLHvDzYOVU/7ZNW42RU+MpHs1ju56Et2UtgT3nMMT0
gAgntY4/hwEaoUOKquCpKUerJmK9U+xIy4E28oMUEl/AeRp+IQJyRDj5wdYa7MpSPdwzGJ2RZDAG
NIv/u69gAqKGlE0yCD+5Vc+b3J7h/XjpenqjDdcvTwQTL4cG8lLGlBAdqBwh2PZJc8l0LLY2lUcr
H8k+6xMUmGVsKkBzR9bbT5jhPXu5ly5nt4txQtFo2yCAPvSz2JpajKXCaSwt17QwJGn1sstumoaS
/F+gxUF/IoqA+hXF9fSmY71eSB6V72CYXXSUrxZZEprLx2qt7mEvARD2nTXMcY5pMRu00Gacz9aK
g6K1hgML8q8IEZpUd7f6r440RIuWvVPIdqEEWkSu+DtuWO9k7+DiJZzSCj323Agw6neu51Fqmv1F
zSxC1qHvwpUuviTRM2TDFzirpTqCtjO+TKpXMylTkznnkK25y4duzWlVye+uKIJHda+4F4TaMNBs
I9bLjG4TBNl7m8qpK5jKLkxi38Xm2yZFyxOO15cM22O7tNf/NkG4frDk3pn7Uw3+CJ9z8dFJ0Qqw
cs90eteS0g2pE4ptIC9R20L/rPxDiMvzNo/VZloToYGG8TkovnDI7TA0eb5vVIQsDRqcV52T7Otk
v7Y9Q38+veGS3TKsTpsUZQiRb4x6cTcrE9l6mWwcwHBl7g4ML+54Q+WeAPRSLXnM9ViQRt0NX37w
F1K0y6UxADTkxuCnD9EqEO96YfYOueGyeMNcANAKpke4NinOLojXiop+4JppAQ0R5nBsVuKq4ikN
PsDMoW0Y+3oPSXtFMcnXy9UptA2V9pq0ZkrT/Qal0LiAigwrjwr5JVEY7gQEOKCtGGcDPImd87io
LjyMXTQBioC5EFpfjEBg0nVtbcKIG7Ipld4Zo1RfKNXWEVPZGJwis5vSM4PiVHC7gZtagBJ5dufx
E4jfKLEBkRQ+thgPW/515Hy6+SdyIii1b7lS4EOuESBnOC2Ba0dPR6XjuGlrFIEIdrMncDzx/W6V
C7k1K1qfFyg80cgzN3uXnno9+bc/iydms9VAQuGotIK43eKv9rS6cp8/8lc/vSDZARWzZciePKg6
gll9MeafW5oeueg4NBgsyNKinogpa4q5sBSdAbQidNUgrZr7Kn/Ir99K5zhrcKsf3OXvjfavAqoX
YCj+dPle7LqtDNebLlI/7P8CDp/t2kt+slVahQFEvE3In4HdYJxUAUTYgkwcq5x74h8N439nd6qs
SKg1qbkR4xaZPXo8qegB2Ee822eNPH3XcUP55qHLwiQnLfBJPD+r1FkbtSt2EAlWmsT4W7ImWjCH
Ru5EHEo/K/NMXiRkDPrrQ7F6cK8z0evoeWO3V6AOxFI5obHlx4VkXqLQGvDlKxi183H2VSl7c33X
KZP2hnKf/Dtv1cK6SXKh+twxZEU/+ELPnrqM5n9T9KUwBKwTBo6rxO9yRaWpqlMvcbujKxQikEYa
XuDK97+0acBijCkfWkl7TRwbC/O7psJSw4z7N/ML5MD1e6w0zJYNaw/xsiRo+Vu0wlO4bOQSlV2v
DAuynSNMARUjzDpHeyyoGC96EJDhVAdLzIBrrZ2VCkoIITRzwT+JWp0baxpZTWSqzqpbPl21E/aw
zw2l39uxzqJ+iJB/hZoUhnXYhNiIHgs2r+LPoWej6WlKBz7GuUX8jpMpAPXVDZH9DpA6TVB53wv4
hkCSTaSZVf9UkTTJutmCAi7XLTUqZzehntVmr4gMv20dRYam+6y4Vo0ffpqtrfNsYTPnbVqEHBdj
xspo3yTgZhMIG3DsvHnqX1dyvRphPYJr08TySQSi32sRAKdO6MFGnLCyzAAqnb8RRNl8KJbXzDs3
p0QIEIJWjSsT5PfM3nwMK3lkPyJJ0+ZK6c87nCu7EUqsQcO4xKiD5u5b9S6dVIZ79oxaPrGEV0ff
75FRisXC0BIT0QWQroZQdM41n0Qz7Umxx45HFS+vXvptguvmZzFPFJhunm4q+F6L72UQTnODp1Wo
Ub/IQnkJn7jy3QLfToiu6egu671PVn7k4uI66+DecFUj3Buuc06Mcl5Xj123cdB6TNc8rxvwfyKU
Hd40ma+TxfZUev9JCjO2Q6ONvPn3BJz8iGfi+Ilt5BSH3wlOmGNH1YuNNzzj0ZZqKuGQ937asXC8
VtI8/XLZPW92XxwIzVFxDu80VSuIJTjr1MuEigVCk7Ag1MIh9Ct8Qg0IrI4uX2qecqB7z4uPaUcP
gg8bR3ciRXpxvqBBHD3+h1yYsLAJw4giXk2CPpiL+20XC5bpvr8I409ouoJkmlBWnk5/LyKlX+Bh
7DtDn7pHLzPGd/iBm6LJ3fKYp/yQK7mvu53v5OCdjkTDWQuflCKq9MbOv3xM1ppTEUduKZWxCbyb
0oV4PoEo3z322DMKhIGDxzILGUlmITuXnRS0G7wYFG/AkqUtlaDP7p/LzLxJHVzgnLHuCq80mzLg
nDqHnrGnGJtnJyvs3fIzOw0k/65siYF5G6YJKiAbQfna3KMcxLclkUs5/cbxtbLNjQwiumTVf7sa
nLKp0c7WVXltulYthG7u3XtNfqP2bvbTgKtEW471T1b+DFA23P3njaAUEh4kkRU3SgyDUwFXvQDp
bTvRWvPs5kZZxmL5+AaDMgzfUtmthc6kWlFkHvhgedfZjD3JobU6xnISGVd7Gepf8qLw5Gl+doVw
bmD5hGC2FiemY4oNa70QyIDw3A0SV60A9eQ+ofJ7Y6bD9AeOkQ2PENSjyNqQDYL8WAFC5DzoXnFj
I+v32hUYXc3XR6cdl7VLDDe7N2WWUjbcRgnfXHQssTibLy10yy/CsXVD7zPF0nrRVGlvYKiojPaq
/Ll95RVsoFUpkhKlbmZuYmxveOCyn+pwXfd2+1kj8NGMlDcfla7p0vCHq6KYlcKTMILJHFMOFu4g
6ndtug0HlwYzFJDRUjvBQ8AjcRntFleAoc5Fv3Cmd9x5PEBnKg1ubwdff0OxbtqCqFHtZ7Lg4Hmp
4rFMFVJG4wUZu8EXkxHK6DEPJ0ipJesNJHQRgM2KmVsCxBP81xBqir1hNBjiqApo4yZwnSncniVN
vUiY8MmMSwVTP9lU7lt2w3xfwH1MIWBDMVccpf2q632eBPOEnuqyVuyNKhEDB3wZNanAlW6Z1qjm
iWAfcrJurcKN5RRRXgqtwAJddLg5ZpkwMcYjRDekyd8VWBuSmNnjC1AUMkwhvn5xsEDU4ZC70fgp
AJR0a+F0V8e5uwoiYPsy11L2HNGlHdxqAUqU6BeZTGk3KVZHAHj30n20hYl/pJINFVPQCcYNG4UM
nU9o++IIKBHZMReo/lLKf0jebPU4znmFvAzFvQun4yODsPX4mmObSKi/s6Fqy1BsBCSM8dzlrJIJ
/NMX3GUJXpyjG/WWVT+rn+NCt115ryqOz538AwYF9TCpRQrogQ6xSyKeWC0E8dSMJ7mmPJuX8OCI
U/nXClwhIg3tsf3AQwdiWlGufveqFbGBYbY8qlSQzp8sbq5uoitWISzACRPHFFzZnRDjHoKgZKJg
e6MK0DyYJf90hrO0DaDW4XI2Gci9O9/4PRr/82iVdwpoihpMkyKlH2WUAQdUPTgD+G46EyTkX6e+
DmcFV6veATcFRlZfsR4Js4ct8sArEF+AxAlMFEuABHLkbcSzx0gpKY/fNF/frEh4w9fSUNiZbmVq
ppFeKpiUSOt56x+EW2jagMtnfWDOKsRuOfLM6ELrAOaOjsKgEYFqRRyYcAyeOz2pCuYAvtoJZLd+
28evCT80NOpmjj4zN5Xeg8qilz7wsNXkuxL8T/0c94nO3c4bzePeo5W77ZnOIR4dQlXJDUwMdGYg
rVClQihjabj6lDQRK/Nob82sfc0fgIu2I8WTQ+zlzObw9oEfRiVIEfm5x+wZr5F7tUw+VErcsNlB
6wvrnMgvQnejMVAtFSWtf2bCs/jmb31MiON9fzZnAt+kEpI3yWWeRXGNs9+nATHUzh6mxeNAE2eN
0qoLYu1WDYiksZxpHcIJ+DlYu8SmHYzvDkdD6PYxO2rZsaQayAVeCm4O10QGOPpTTCkZMHppV2sD
8ruBOP/VzeAeLevdnkTZuZ9rIDj2owB3zms7VI3wkOeIB5ZerPFQ+ACJ4HBwnCuwepp8X+WZXFHp
2L0QNOtHhB5cTmA+U3mtv83WUrdCvvB2s8ufYMW2z3Jn2W0fkEDDe6Vr3jqCUye+MBNbmC7FYtYJ
zNKRIHYS0UK5mmpe5XH5zHkJzVx9oJ/I7C9ZEUN/1UTRCJU0eoyLG8BMWz4ZNuikwuuZC0TPPiMK
Alv63kB2pPh8bEBbnriB/03edOTwsLD6wl5xnnMYo+eC55FJsSqktqchJ12oUQYWgD+iMXhFXKm7
Yk2Bwb9Sxga6SMlW1v99WTvBbHckWnW1URRrV7ODWx6MHN5vbybVXaC/zjeXmXr78ub3ZrXg5Qym
9XZk0OIBOP8MUPadgyKVr+hBulCUR3jR2GBJi+ELkX5J1RyWmN3206eDqkcP+pOlJclYHND0khQe
xGlVw9PjLAys6TNvbZ6sLyjmEYwAEYvV+9Kb8QIz4BB8G1KgzhlyZbHU0qeo4NQ1lIUslSHBHn0s
LXZjc/12y2nGAvUr9yvHcBM4vnYXoHp77ra1SuF68tMp/aLmub5cYfA0m8gYIaOM/MKgscuNLTY7
UQuX1tUlHdNDShMeRZffe0zEUnQjo94mFrzVscUFv0deTtH4W7j4zkYFKpvc+qnmVl02tCPmTbCI
/Y3D6pDjag9mc7pzybvkI2UKn507JwfUnuMPsIGv0scZYv54DOQtMIK51+fzA1QPSUcdRT9MJ+61
HXK80Ii48xy9pIh+d1+XTeUqkMbb4WzH6iig+t6/G3xZqZK0hQZMgz1Ws9kkFXQ+cErwpT7eX5S2
E1pvT5bnMRxV/mFXu/GFpo4TGKlfsXf0hn1oILRhrz2y4GMxCbBfTGVwCg+ft2r85h8hqUF6v15D
WUVaCsOs/fovk9bsam+z33HeVFIwEih9/Y8kXeW/DuJjPPhRdechOQ9Qy9jf2mZK2uTztct22hk7
7YzTqMXoucDNvKzz0r6qYA/2I9ABuKHQCAtxcUJ6fvLdPyrz9gMbD655YtYA8nbwlQgzLp59N6QQ
Kt8Vy3dBnAdttNzSR7tfJZqHJK+PRQvs1UbZF4E0bZrBBkUPWJUs/OLC9H3w37Lpod4CYkjXHgVz
rTBtqBxv4KwFij+X7PoxW7uYGyZXJfhQSqCDCkU9WmEuFw+v6fqmO4rrXl8b0YpofVArvIjKZCCx
+dZUA5npa3VuO6XVwPIO/RjhNTznmCvdJpY1xB2XS5/RuSHCG3YluTY4Gb6RCWi2SKZTr5qZt0Ss
Hl0FBXQZM+PrJl2m09EM2H7dtpy4+lYMSfasft5R44zO74jTnWouZpPMJbHnJi9Rwrd2gk/VBfcg
gQsmOURcCCA26rj5FbIVK5pozOqhHpHEp995B5ziesjiz1QeRNvS/lw7qdIeEB+KxXKfZTseqqk8
1Za1DTB2QNmajSEqeCqV4ydU02xzL1kDPql1iPX2ix9vRlqpnI8Sb2quAxMGCUOqxilksqaXOgZ7
258bkCaWip7TdoaMTCCDvJkKpdMdRLWRhnD4E/AtXU5H2jF3VzhvrfnNyfuTkAKWsF2ByKPYGiUN
nQzhF2RbMDtsxYxMxiLSYRdB8w0f/9yOSkkO2JoNapEhKpnhH2e9tLRxaftyU/e/G9pD1pytoWhC
9ikzSqWH0YD3Drr0mNGoIPUYrwO5ToN6Mw/7qcq+8l8nDrYJykMsEQiPSADy68MsNCds8mJqPedC
PvrOUXwu8e6BUsYn1rdVy3H5j4E9d/DaOkGr+FKYGFpussczVNcW+2zwPUMSj11nWgOrThvq/x2k
63gPMdPwUmkt5NrxXDt3WYq+EhBNk5EFhtFF8ao2M69vZd9YDztSqc6l/coUcFE7bd8uO1zfoZzd
FekcbVoOIoD16UwbMJh9W2KhzQW35U4KVWR79XDY9D1JZIT+vHoDEzKmcEXrwW3kuVOFCCrFuUGy
N3zJWAVWWvtN+wdDcNffJr/FAFrfeUEMMEXVGTrbovN4SzC80kXBRtCXpZC8P4JJl1pRIiYEjrSe
pmrKhmD3yd8JgvfrpFsBikkV3VW3t37uo8NmNHxIJqa0PYfG9GmX5MM5yeqgL7GhEvLQBKtll7al
sJL/TEh48B26h1PgTzUC9azqc1Fc9xumlEISZhK/UG6AQ0kFr8ZzwaN4PWzfLMFNlU6skmFGbOMQ
SCBgbc9SWFpZKRMlHS49ZXsW2R8LgPYIKkMdmexKJemrR8UITW11f3hccqdb4M6tDOvsAc+aQS9I
yFeyyxNpfdP19VwuF9kqkxa6ztqP/mbjb4ql6BQq0bET9eKP9WW6zUaLQrAj1+LTsqr/6TJHqW6X
Ef7G9Lb+eQQb6SS3zyDyR22mOnZcJiKy7dmFuDfyo+0GhplIQgKZt/Hpo+gdGS48KQWky8lrsiA1
myqtEqWIGA+3/P1BzIqc/Z6I9lKEjpW+BVvXx6kQIJ8iMVQMwyyB9A1xvmo/zW8fSzJ7w1yrPhWn
H1R3H0FaIijYIY+fB1dsmB/JBMq7Fhftnw2qUZtCH56QX9KMW2pSqf2QlzTfwJTeZnSTeYoiGpz0
EXIZNg/T12u5AGt7cPRVy/sv/uoYfaAEra/dmS6KxaL8XX1PpqIddv+mdD8WBH/ld/wHdX55rjEs
H5b0KyHNmFgfAFRSGiII3lvk7Uwn9r05v2U5x8OwZ0Xgw3XVofyGRONbbtOrsmv20uWMwVL+U5hP
EXSHtjPWGDQwECmnvl7FehFuviET2nOpWcCGVzbrm8ByjGEH0DiqkFxGOFDeTFG9wJIC42yKH6BZ
hoEsSBmBX8/N4zjFs4W5HdxsHkhD8gSs9qIe1DHTI1tkcprY4GuisbvFNvTXtRsG6GpvXwQ+JtBh
/QOAnOPc8A96G5iG4BJ7Dg4smWnN2pGOaLv5ekQEAtOfyMn2XdfnhpEu0c1jIl0RR+70SPbccis2
AjuuA6j3tKW/kGc0Ij/c+THskCdVhT0myyhZpVopdoE1ywjg6EiOjYmlhJDFSyYcIPtDWLCznOxz
5Q3SfCkQrIOSC1sYudMjO+tKkSpSGqavughzb9gahZyj+U8HqsmXB7QIy4UxvyQC4+YH8B77ijF5
tLu9ETiVLE87Kl9LiSdA0Efp50ppe9jjCUyZeEGYoXAziqpU/ghab7IeVKrmfjdsE/dFbK/j/3HI
PP95GULEJz+dRxUmh5FEwhpHVFOo64/OfAtVxwvSiqvX140wlgKWyfcI3Kmnm6yUmSy69L1RdCAg
9MkyspgYp51td8+T62Ub9d6fj3SLBNT/SdYcbZ2I04bI0wZoDwzD+qbspyJg7uvhV6/nLBicCg1i
mKW9af0ruelGs+raRfoqMyzmmZfOwFPC0kE1nTUHVBNX/koD5baqOMADsaXPlQ1Hf6SZZBkGckSn
AA43xCCQf5RRkWwpt6+5qLz8Rml2tYiOJD2hvELe0WfmKcQhspiPW8hz+ccMdR2E5vPZmaUOD2wK
rnuWc9X47aIG3JqoCbOp4SdXb0cZaBWhNm7mP7ond5DYKxDt6Rx+8EA/dS3ULC15AFJP2fb4T1Hb
nCCV2DHlYUGuZSj3URwW6SEj2LEOiECLM96nnWI8P8PWARbyVttr/U1uyaMw4pg1PS6CpUeRHs+G
FrWsIdrs0ynMepMOucMChPPdR2DNZn7FqQVr07FoecgZkPrhhfU4Ys8x/IVl1tguBYAgO1Xcybdp
dNfZeoNXz/O28rXLx1dXhATKqqPtIFb/W4od4w1NfEPJjAqxk0cXSLQ6vIRy1PSmtI8U5OuozpZm
GG2FY1GPwQlACr4EhmVxmxJ5wkxr+DSo03F091qVo++lXVRTe5E7Tddyq98bjxQu+2lMdEsxcBLO
7Wc5EjW+ZGlbRcTYUPNvFDtD4gSVfNEFTIl1zhT9b8cONZkAtSQD37LEW7Y9gbhi/B9TWNOY34GL
V1Wfn0xF1/3HT24GRzTpPCXtB9WlZtcjXLp/9vjNhIGMwUGMNkBp9XYdPNDyjhRgpsXFSNXQB2jz
1QvH2vzxY9HgLwKvvlh8JVHCu6jgPoGRAc4m+Lmpmfep2XSzLmqKGOV2BY8WfJ/ENfrjaTqYl7EU
Sqp3Iwggz5EtQtclbB+z/O0PWOz0274hEl2fwlOr99XXYIk8BeZ0AxDzJBBWAK5oPG0mDrBgHZQa
WtDDMN+Ar12QMgscXfnprtH3gNYxiRYqsR/qYz5W1rjt8ackeDh8EAlIDmKgRf0x35raAadm8l6E
CHiu21J7P0YnKDHukiF9cflQCBuf3LG0Khqo3zX8iuGBN+B7AWpjoMwNqNFFRgY4vTgyh9DDrgqg
UflY5z1lqJLZR72nGiTqs0qugabS8fN0rrWj1lr2YiX4dAByyf4kEqGqeogylTUQ5TyFWSPRybbl
R0bF8UAPUBw/WmMimYg8rKrNDF3YzVPfO24+fZFIcn19q4jQyPkN2n4Obamxlp0GVLO7teMEQVjI
ElZ0yxdeal5D22ZmiyM0D/DHAsZcOxBXNoXHASwJLx5FFwbZfbZzz6uYZlznmztfB8qfG2D39BYs
oHr8Lr72SXZcXwsJ8UBRIG1SQ1X9kFaIkD6V1p2xJfji8jFSUzjhYq2V4Q5Y1RY08JJw7XLrEusO
t17i7SYYyCBBa/piq53Y8iBInMkktqG+dEZImB3Z/WyPSMmSGr0PHYYME0Xtjcy28WQuxk88W1GT
3UXIw4V4gri5mAvvhlXt1WRjOYbGhstOp0zjtd220eNbqLTr5zCbHuC2gVA1tjRjL60oaT+hRO6x
vKJelopee+IZHeqcJps38LY13y9+ZIbqVXNp0ydX8KYpcF7h71f8d2TwMdgyQ0y5rwjuN8OxB6/x
oaFc51j2fOsPMoI1ud8GBrwZMvorbTIWbjOKNXKvM2MYfZFjDq95/Qh181F8aBjl4qBkoT46BpOa
M173bwP27h/Pg5llA1AYLAIf9rWAKOD3R3YgLIADWeZKJcPH4JRYvG+xIeFjDW65ZGJK3lM18bo0
4iRGj/CdM2Z3t/2B4T3vgl6uvkkbXD2VMqzCXu2nt5bGuJm2Wtb+sUwnFDo1NCv/NzKvj2eMTFSN
i6Iz49UHCtqB4pISTa7zKaKkbbs/x3IcErZ/S2SDmp8aaYAmh1Jyhz8mRaYHFLdqtTPtOUcgSewJ
0jK6bnHlwtwkZBgItj+YVpkhK+sG8rlmDqBVGSrn5tufLjFEb+XYyJ+TLbjJA0Uz/0iNG+BLI3LP
7jd1XTpOd1CR/4rJzOgSMcO8urh72w8+Wudf0/kXIvXlVSJStOduuWbtImsP6qzz3o92aad+U4jN
0n3VRuSI57or5ymzk4azwTaLav9oNFIs9cb85WnRkLBteE8qalOj3ymfaZqjYBM5haxjqFBTS0T4
ICZT4WP+NcHriu5YeFiJhDJKTuzHeaBs71SFr37PbleWRUV8jJMlEqU7sJ3ggsImrJ3eK7LAgscM
hU2XoCVYJEcfhk0JDyU4X/VeEkZp7u2j1ZZwrEgalIplL+Yqda5Pyd1tvcfQSDW6cvt3CyW0Eulw
ub+hautB2Z+hzDxHaYYQhC6I6dAHEX4alo1EtloG03GoCQ9q6oos2wjaNWnBAJQ/uCYp4XHWRWFk
qFSnSt8u6hLAwZUfluSxTKNP9bkXU76UWTpSQlRWATgBz8oDV4QqwW/j8Y9PDVLSeWBugNyGIprH
zSnHypLU3cpTtVjB3mcM5owsAEkReSNx+75QtattX7wdVRs3+SfU7Tq7h1DvK1Ab7evhRVVdbNrL
b5x+uXZQroCXgW/w0khIV4pYoue72XYjFUVJOwgsZQkYFtrpQd5zZbJgt5PwIn2QeA/0xopYuEnU
o3L865uBnuM1IfZ3k+rZWchHplH+3F2wU/e7iTKpPjDj/RRPm4mjulRVjvNSn6xho9P9U5iCh1lW
sIxeYt2GYFSW7VqX5bPAkdw9CUh6WYHpxh3Qj8NDjgFnU0sGPqnIR1e1X+ooXl30kyCokYGpGjDu
/J6QNPnMW+5kskOenQjVjH5EiVFmN7REg3K3mu2KHBAE+WwvvkvD1ZJHuAK4inl3Bla0t5Bj8asa
B07akKnqOuFhW7WIvvsu6dIy6cq2VY/nNk+zDVuPZbmRgEEYgGSpfpCKSG9hH9H0fq0cj33x1h6P
apsvjfiiRVq8fL2UfVNruh5Mhb1hQ+WysLrWN/SiD8JsV2W3Bsl9Fv2bKZ8jEKE3DVwbIr4CD0Vh
f9+wuOpoCNwzKvytEzP88Dx1dMHJoxgDXqJvkBkxvlBZjt/Lw1gpv2gjbtVFFc4SiubyX9NKfVEs
jskFWGz7hxZ7hWptbwJdxTuR+UWCg3kRAauKgiII9M8zNbtE+RVCuEv+YaXpkYvA42ygDPpY716N
dCmpYlGf5GLeVnwrYPxnf5L62sV5YTcWKxv8B49KGLSdTvJQnqLbqmb/IRkQNeJky/ZH1ISffO65
cpbjX82MMaYsDSokaeuCLCMHRPkIkryd0jE8upxt/gvHUWgdBZCWIUqKuLp9BywYSQgcF40mAedc
hfhfQIoUG8FrNmT5LH7r0nTfVrpc8OpfkyS0znmSqZttyJavap+BgMNFbFiaRg9nzfzhP0eVKIeG
RjVtFjNsf8XZB8Kre6GBgi3wrrydrk0AkqCNF7Ix0FB54vxMqjf6FwHBB7LPN/2Nxe2AQE5vNA3A
crgJ5L5fsz/2+eYfoHANly5UKvELkYE5JfsZeYXiCa1M6N4/DQJhgUFVPafdej4HhtIBiIsySM1o
dFgFxHPBv68qtgmf2nlRchZvDSGS3IF4gg9/VTkRH5T9ncr/XpjGn/WmCWD/x8ESC0bw7NWYw0tl
9HCRH3mJhWzypzv1Ibu+EW49spbhQ6s07X9spXMBdvxdjSFSaNU/daN+rh1gELZhgYg18u4+jiBf
Wl2dX8SxNjTmdaq346pklyPDuENmsK/L6YPftXa5ZuinEZbftKTCHa79efmsj2K+QERqAfQUJt43
2bPEWwgmpY2cD0UIT7kraxeNxR17B0097p0SnfoIcpx1vsGfEmDO9+zeCnYcfoelcH0/rM6ChDZU
NOGGvSROfzfNWIWZem7QYTHF/7G4kEshzAfwjN4Cq+qdASmnCSu+67KR6Q0NzPCHsJT0h+et39cI
hHsZs6WzhXOILAh68xBZ7pQse6M+oaqNk1a1dYjLIPLa/Z00IpWTGqikxZW+poJodkza7fPjmfdz
lvxDxDVzm1RfU5g4E9pmUj0D/A4Kpt7Sf1PMsOfZhdDydFXFLtTtjNBo/5Dew9aIIwXSAciyhO/w
8yfenPWWWMZumJxAQrmeT4P9qD3/LcAc0jKqsMjAQr3bA36bHNMaKVnUSZZiG1zOQBo7KTD8Gg/k
aB/q0AreRAwuRlM71Eo4+V7jhhbZSIJ29B4Rls8NTAbwu0Pqdo+KSaFP5mVkmGV1nSrjUCI3qRjF
zY7Y1fnnBhaiCCIsLpsOshK0x+p8Pl8rC7Pvmv1sdVxhLCM5FHqbbydFhyt5AbKUlrAI+oSzhNzE
Di3aD2JDx9RNxQE/wgROVIQpc20hW6Pl0gso/1H5LkaDiItPqVsLX2awCo4fxFSlcdCfZEOdD3XY
luvjESECToW2zxPNgZCvhGIIps6KzpKaISG57f9wzqjVrjntTGI5yD080jCzFX/7+4xyLn9ihbjU
Vtw8pINbrnriw9AN2Zb+HMz6iQppuwYISgj2dKTbPYsWQzmGDf0XeBrmlXzVPVZSwF/fh7OBnRJJ
dETSPBAcWnvb9CRfmfVfmmWc1VCUeCKrAYX5/Jr68o15TxZpsjyyKl9i4I9P23nLDJUurUEXo+tI
+aZrrpA0QtHKIg/LS7tZ/TaAR1kaNQnzefEW3YuBZq3zxp/EL0MGYIMvVIluNrUAOKwE9ODcgvPa
opaLrlPlkRrNLGwwLxmSc/JC1Eih8mMju5eXS64ex84ruBQ5Ioi9LoZAugwh2H7IA7WkACR/4fph
wsZvaNHgVGUrokJMpfyGKLH74jrieHmWMRQCBFw0vNOaPJIBX7c5AcuF8dmQCtDHpnyvq3IF4n/d
Z2F8ijxfPDtRsVxM+4F5xyk2h+p5HZ/smXTiEhIBv10/ayocM8YWHDFjZdLWkdOsDSeEFa/YdQlz
Yry756ULJSXDghFXxvUR39gDr4qo0GB9m6lntwoz8Gmp3uzTIf2C4DN3EsK58iGtB30Nwv7xiLKF
cwUuG4cbGtIiATnS2IY9LzoH5kHXR2Javi1bDlM1zdFZoELFM3uUtjbDLTiDs2Qs9fNRu3baosDC
0gxGOH1qX098dbhELNlUpHY31xto2P6K7Df/2Wl3IUre9NNT9aYTPVrpgETVJ4KKN0aC2EEowwtf
RAq07iHZ+SmpBAbP0dBwzz/p7F8G5vNr0FtEkI8NmdAPb11PthNM6vb5VI82i2XVp7Inp/2zN7kz
yOV25CsK8cQvjdjp5gtbTUdq0F57PRx8o2wDA2M6oAPYsDkL1zTIdVtz/ErkJF4naDwcvG5PeXym
+lOQzH2AlAIEfJ6K6lxaI9SdY6GcLvTQzMj+EHzmeeCg5NfsoBCp8u3/+ZGsyFH2JguAPlyMiMpl
lw3LFCD5Axrvep3s9O0s+dQI5wjy6DPnrkeIqCIkuf+pPD31OsjnwOGU6PGqmw/iQ6/urD/ynF6C
UWLaMI2eIAXI4uR+UXdIzERGgkBpHB/IzxGLboZd5wK3+cFxUXV08NCYNU9yanJCYhiZDHnXtJqk
kca2UN38fWEaBQnYEcbgekNJ0z7Z4lsclkuoLRWvJExZdsnoSfMkeZ9aIM318n3HSzYNA949TuJ+
QRyHC+K9AtPsSMIczr/7OZOUG/9pZqbWMVXdr8gMLRMo7P4J2gwbQEp1tFb0WgArxTBt07QTnNIE
laiqH2vuZiGqVZg9eBOSYMrhbyvIouFZV/QmW6ke3c5VvQ4ydXqunqPO0rhL1+nSCE7PSwuggqG9
Wk5PyJPGOaoVkaltz8f9YRTzl5LoBI+QNbTImO1/jsf8o6x+Z6owd49gSnFe54L4tqSbeSkpQmDC
BQSWHoOuPs1z6GFDwUwb+msI3Bv+IGdX6XEEeZwggdMVxb/CF1Q6vx8W6Rd1JE4MBNlItN6bwSQI
exPcSuUsevMZzOf4zBCqyZqJMbqzr79KtbO0sknvZwSOcnRGez95IUO9fLjb5phX6wWROHv7wzoG
PkKLeyq5xe/teTZw1CP9VA36UUTNMsxg3kvuNLKZpUR9Mh9w1UAisINOHAFgFxcZ+hS7pczYF0UL
LZYhd0duqY57nJiOanTXEswIQnWtFJfpizPfTB9krO6/oum//RUYLA4DUqlXCCtqKT/qaNXYmd1C
2xFl9pn6MKAtvBgyDB3TNPue6VQvec4gdjaUXF615wFUsPfzyhEKHRHq3R0VoSPem0a/SrAHYxFA
G9NNU5kfEzd+kD0DVMhH/MQZgVoTn8WMGi4C+xHtHSnaIjZWJojM7RvZYLruBc8rQwKQ89M5DEzj
nN8uATCUHwKJJwnjiFtPNaFDOJOkDzdSL77XlP/V2mRowHGQIiQGCnlyFGUyM3yH11lKCPWdbp6M
BCaUqad7A2aVqtcRzLah/qG5RqNKOS4Y78ev7KQKLEH9ZWRoqkw5ykB8CjAwzghzgH/THD0RL20O
9SV4+ziQThZLkX59R76PHUEB1VwQy/5ZNn3SJ0qtUu/VPj5tZUwJIFMjFT1cDpA6CFNxuXo9lbHC
RtFMNSUikYnyPEBDa7iqMWtHY8dUBUb7kCOOpK4RgAfAWU87sNIatTGrTPXUWrCE245zbCQafzKG
panx0pat+Y3ebJwwRpvPUD315NsuFjRC0VopAuZyVK9B1Amjuxh5A3MhhZAtlqMVG3i4BlBU+gAz
2YiXPOc0h17UzjXttO05Um4tabfebl1uF4gCWE52RhNkCtc6mwCnxnLstte84i6kCR5bCMDB5wzp
V0ROc4MSAi4Mwbgswhvgrsc5Fcd4DHCMphKH1XwqTk8goqL0pOoJ5049/wtwxe5M9kORbrEc1JKO
OIwG70TtwGPBSBMsPa0IMY9Q89rkGZa8gQTpC391GYoOMVHgcw724+6oEh3J6sqrhG/9PLUF+WzN
1fo6hw/XkUnKVJF0S0OGJKehFHgtVpIMqj6jXus5j8+2NjGB6F1uQAECOcNkNVpuTOwedZbxkm48
ClJbmCAjrZ2mCg1DvwrmhSj8li7IfVYB+J+5nSZ9cBibzhf3TRe8tWdGC6LRuaeUJx847oOcMtkR
9eVSiUM5OzN6N6F/XVqG/IDQJMgdHQviT2TfDEu22n39B7RqYyiodrQJqStsUtkldc+R7zdLNggh
0XE2GLwiTd+JgA6ABNR/WucbGAnXuhjfxyXBCPZ5LFiDXV15wwXGbLkLiC1YfWSjLlB36NJWLGV2
UQVSUmzjIu2MFRW/sNxwCjya1syAaQ7Ww/3GdnhvsaV99WRB64WKBf+3kyRwhpnwehmpbdWRhagS
juS4E1Q7dmt52Jo+BF7B5qAUxUqX6DHK/e1ESBUlPZNkt5erFmI2Ta3Ro24/GDBJ2JS8q0d+pxKp
Q3f2i6cN8f9e0EEnPfHTsVmbW+O4mOxVMcOpuFKvBRG13mq4ZpkaytXVLCO6ISEgpYpKpv/XzfW8
zxci9M0bOHf3768gldg4QR8Eb7a0uO/cv3Ev6NQ5W/LNyok/z848vzJsJjjUo1LcEv3GIgf4XgC2
L1p4iBLt64FRsTEOOkPBOwuVbyRqYjPqys+nE3raHbZVphDJ7xl4JmEL1w5nMKZhqFRNmuVhOmD6
R7CyLJCf2YwbJLH3O1p/7mI+4/AC0ojBbuy7Lasju7L0CUQhs8gDOMR1j38s1r/AYlPCEisSitDC
9Fjmp+j+vpjsmoSmaV1RSb5OO3HXuJZT+RXGb1gBo96sbJsq9zhZcIbmx1HiBejTFMLSZmkQzJ8w
2+UmzUqQEdFgVojf2vCekM3MrSXjZDPdt3ivDMox7lINUF1gbXaYWFrL6gnd1SHeuRKxGSDtZxdC
yYv84xZNABHcXO2+MPZB1I3+5bssqrMPhOvWW6yt1hL4vZq32+Cuo+Uez5RSTAiwFdP43HKzGVC4
VeCOgOXGlgGXdDB/KR/WvE8TfZD4jomlB9ImQDhHcrFSRioE5FIJCZXdgNCSKC2JHu9BP9EIJNKR
RftqAKnFQFKsbGVXXB/Lc7ZUnN/NGUgY9rvjyUQ30hhaSOC1P96C7z1Asvq+Nz2wvRbvAwCtC6gT
ATivjcQ0AYayz8IYt9gDZAFxbcZRAz0SQJMrFsz4x+dwpyDZiEDRSzHhMYPOTBqMFb+LqBB+QvTk
0L9WF/BHBEdEEXUBJtRn02espFCVQLUtWMGDKOqfJMWIcSkpumxHiR9m7y03xUDA2XR3y+bAmw2w
ae3sAqNJF7Z8U7WzxoB2ZtfdPq0jUt4n+jWRT4nlVYc2SzM+xn0hNovoUo0Fw9pmZBwxZtmXj1iv
s7vvNAucNZQAjc09zvQ7PwLf7Hy/RmId+DKVq0QiB+PTny9Af7l5C1hsI3PU0EK4TI6S8sy+4v/S
C+4HOWtdJQBCSOd6uw/eoYBzUXIStYKKV4kZ2G8JDXRV0V1mOALo9bLduYyrSsUwfiWofN05Rpv3
YfeHth6dAE0CQzKGbTY8GyplXf54HrK6w2cQa1Z1uc3dCRd1gpZGei9/WnuuMb683qOx6SP1H+5z
lsKU7GlGNGMjTGESaCO2tJhTUbfXN3s7M0Mfbd5zpHYjxN2pVkduE+lsPDMKAvEIrZaMTmCwlLIt
/XIsB4/zRqCzNOKJyGU/ALb1FdVpYuGLNkOxe/m5WD49VHCdW/qKyY9mR74XD6rpPnv54/axCoyj
tRj74x60IjrfGUZupiPFiwI0gFPVIDdVZw329dzt19CkN7uCXM1ikOs3TQRE1GaTEU2SJ5qyz7PI
r8PXq3TKhUwHNbX7jd2ovYV3k5SURVnXgyp2Zkbxuqw=
`protect end_protected
