`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
KTNs5rYcDOiviP87YnqKWxkkIbQ9e+LvP7vW2C5y86dmrQTbQGQMfvomRC40QDX27WKpTLb/smFj
n2XXMNinvV+oEdZ2ZODpVLG9LN91tfBeW5vizfdwzkC8i5OAeRHp6eHv/t7/2VEgMiBA/EIuYMEo
UjWkDC+k3y13eU+V6l78DFst5TBurLiLEoFZEU8CsMOKkzXLwYIwYjUWMsnUofMNaiG4w5LWShZO
gB7zakFplbpgjF8VDgQYzUVQlqhdlZ4vKZsAjL8UPZI2hQhdo85zJISgnVU1FF70S4SfAbgvDwEQ
F3lE913eLMmBvRO9K8Ihen0c6pZlUxET1tFKh5GrUhOtEjia2yZjJiSvwP6qZy0arWLEo8s3AX4n
pi1kQyiprh6jkkzU3zwlPRQBkEVhHBIIp+pGZi8ZAbH0nkJAWTEHLXi0DQ4YjuXeraWmiQjxp/8j
iO1Bxdi7QV6Rf6CAzk1WXl9D5232yX+nDIWL4MGH5huqqDs7/7ukqH/mMuTZsBzyJhoURTeZxSEp
fMoLCJk1Cwu1Ej545/AGDe3+8cef/CbcHEMPgC/S+PsFpSJ625cizODBjumAnG6IetKGNq43aGdp
Ce1IjyO/5/tw9mw9xvrYaqitVwuYNKOfLyNkSCDx2LvZbd8Mz6d34Yxh0CWY+M7dV9/Ba7s8QYdL
DP5I/W1HidMkpB9801PXIr1vsS2sGzlOJq9+VTMpM9NReakbyqBLSAF2SfOCWlgUjUO3iUgr/aAQ
AUzfemfhzVTRbwMEUBfXh5vtnG+Lw4X5XFlMQ8QDzepmphLbwnCGaqib5nQvFrkSUVDsuba3ElJQ
P+Lp7hXy31bYgKK5/ftJ/enI8lACvt+g0mSGixTPXjkL9fVeTr4fuKj/MFMbQ3z0EdV14z08ciWz
ePrrckxd/av/H1KbicAvNSnXdxT2OoQOY9yeQHIIIGjGwPDJNUJMMb2dim27cJxi1SKDqBvS5mVP
vA/zAXckDPw/CH4HrUHFPLf6RuMci3m9nA3Q+6U1Skz00o5Gsrd7oHVcp0n6DDsEnOCTfVYmP4BI
VSxDAG7x6S75Edd4pBH5dD9xcgblXZLqpnQrdnYP4jTx1lEx9Mr3+I6xmQ4/vYL+/J7mpkJQ0nAi
wmEFpvSHL8Fre8q4dIoobX6x/lEzbLQk74cC03vQ7lv0lg/dp3qQP/7BjedY2bGjfGwsgzD0GuuC
KTaFiLPKDsW6BNMRoUBFfMejiUmF7w3JK3kGvzyfDYI19wtdim7jj+rktoRfI1FFMZeQ3d92ikuQ
jXZULna+TNFnMrSOf0MwSp9LPWIb6hj4G29k4w+D8jl0k2a/qJ85t6uXqR9pu3DOOFprch7rD2rb
xq86QKQR7lnzjhYu9eQ6V/LaFAX6MhygAtV9+HKIkgTFAxIkkCOcuOPZ1zzKWPxGj/qzfWOGlfDz
YZ5FRstEIEdH/dD+vrpnegIMB3oWWlWroD+uk9NetvOmD4P+1v7/GYMTqiuSpphpACx+9arDdOOv
e281IpevwQv9lMlh8gw02Cx68EbwBwsOeSLGYKg8ReneTUsrbJEvo/0QfRKXmxAuRygJGKoWtRjp
IAoLb77IwS/42c5E3pYPmYXNz9rYfutKRARY7n0j/aNtTtYDomds+2bcBz9o+l6i/nR6IFxx5pW6
BcGuH13D2N97JbiZHVQHBRaoVxOsVx5xxjgLdsGABD9MQd+RkhGrWh7nRWekrZQaCk3+rEH7Y3dm
jKu43Pa++hQ8OJGoJUEaiqW1sCovGGiDlCscfiFdD/yXmPmGS2S2Vync17MutZXNSot6l4R0KmH5
of3Pwl6UxzvxIPEOk3lhiU4GPmvrxcwhzvH0NfLWfcv45PiOmtNw8nt4xsS7DE6TQJ9xzLdD4TzQ
slxHmxVOraLQ7utAd9dzWYkQ0HQ9btzNhnyZqi+YJhBW2s3u83MlHdy3tif8lF5D3pKk25LFn0nc
tcITzZfMbBRsFFKNgADoa1ULI91zJHVWIrZJY5Vf7yD3eBXoXiQx4RJf6Sm+rAlagskmxYhnBRR4
gOucIPCyvda+347x/nib96+sB1P0s2PgOFBldHS4s/IIwMTlGYnL41Hb9qtwRrY9m4B+xvKANE7l
2AS+HsX1o3lRnopLEf2d791JtQwJUqrI61aLETd2+6NeMyzFRwzIolFq1Mzoy5mwddZ+B6J4jo/5
WN0Dria1r1VIAlL+581sdn7tPKF3NGRwTQocVRrZnzKnWfmmNRK6Dwz75YCs3jbsoSgbQAsbtMuG
DfbL01zCll9vr3arHYXEuK959ZR7+X/Y9oeJjvx6L8ruG2Kw2V0XBJA+Twg6xA4cJxpec5galulW
Lgfo0LiMHdI4OaQfJzKHjBqV77+P0H4XFvnsXJ+H+le98MkWwZIkHNegDPvrCaurq/qaf+Li0GRl
BcH9NeywuALEXEwEgKEwz/QODHZw3H72griTjNYhKyLxIUEWbLD3e7dEKcwsa5Ldb+j8PNtgK49N
1OfwgGvGjJYI8+VafMQXEZY2QO0W1i9Cb7lXDBJ7YNKeH1wUNv9DzvY/Vgbdh6gMvX9YyURooUw0
GdtnzymKNGkXi5DmpB9SBvHltR1G8AUEASCjE76QM/0Vo9TUlmDRBxYj0QTdYVWrHfOSAb9RVJa8
AM9AocvAaHB5gj3j7EliWp8iLg4cgojjWh7l7h0/avSns7E32BQFqltxtTkdSG0yNoEVc8E3MrPn
Ywx9QRyybyietqn0CVhR9OAvV3V9cv3Q+kx6V+neKf/QAZeJzlGypf4+yukVNL5sd9ziMVhYP+z0
/O8Zfkjw9L8eT/xaSFmNpscQ/H0x0ulV2dfrIO/+XRE8yf7aq3paB1M66Vq8lvmBSnEW7cp66+3G
Ci+ffllwdTPjKkUiRmIwrsucBME4M6TVdA0iNxGeLUFi6WDV4kVSGf638qhIh1P4RtV3R+FCccOE
k2b3rRgdInP3Kr/8VjQuc+d/oM1Wtw3MIz+tU8y1xadFBQEPoLdBLY9P25N4kEXxMfVj9bwJ2ZPn
vYz5FPxDlz/0O6wAtwgUD6wd78sFDmRJY/gt//0+LMlwS5kxPu+e/UUIMMpmLaQOTbxve22Fth2O
+ekv4hAwRX550Z/DJd3RmEweuwrLi3UhWkDkQVhNpw==
`protect end_protected
