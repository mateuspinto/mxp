XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��鸯��B��_�I�L���u��Lأ���&S1��D50���X�z��y�!�"�G�G14f�(�՞�6L��=�]�.H$WUU-1O��$�7����#�J�<����A��jA���%������Cxvouz���J3��F-r�i�������&�hޛҀ>�="�oge�g���P8E��4���c2㕠��5Z�_F?p�[#�����_�\6.�l�:����G4�P(�/d�/�q�և7���ޔ츚*n���%�	#���J霖w�,㙞�D��0�r�-@ a����!�a�8�F��QH��ZM6��-�_��"�Pի�������C�L������BF�BC��k<to�t�p;2��)�'�ԝ�,�i�¥�mN@ �a��<���,Q&+�|f���L��.Vx�٠�0��J�q\9�3�\78�L�<i"�_)�#�eGԞZ�T^J�.�kn=�ӻ��&�&�����.�O�$��k���MO�܋�kX�9�O�����}dv�?���:����n$r�P0��QeP9��'�ΏD�;��-1oJ��ws���3@��gh���B[��{(d���\�M�{�mFj��ݍ�^E��z��N蔯�-�~7yo����.�ɰq�5)�/�����cLnZ���D�=��+����������	^�:�&�a�[3xz֎?��:1�;'drx|���WN��� �R4;�{�/�U:��6ukP(Y�h��V!�(��-�3�)?��G�lXlxVHYEB     400     1c0�ej�}�N�
t�����]�zta��O��%ȟ�TiN@��|f"˽���M4�(/8F�H�+�Q		1�h]�-j�?�Hбz	5~:�J׈��m~��@M��?& _L�C��������e���J4=Yۿ�W}�t+̯:e�K�N�:�kb�]q���k��������U����DW#�v� |bơ�j-V��6���)Y/IKЬBȬ�:�[`pRZ��8&V��Qm��ܫQ^��k��"��O��ĭ�@�8iqµbaG��G���[aU�kWo!_�o�18'=����)�B��V
���~U��c�W
��{n���	�ΐ�DK*��3ԌۖU�;:Lކ�C��71�S1W�|�� 3���W�&/=J6���J��1�Fh�jdBs�m۸�~���E�L­����Mj{y���8���q���|;~�l�XlxVHYEB     400     160:���{�wH��X�_aL����iOu��]J 3���h�J����	Kv�{�U�<\S]�4�	F|��t�O��01�#x�'ӎ\�
��g�P��;2������IU�p8g�P��Bq�.����N�$w_xA�j��� ;<iT�Έ�|o���l1�l�u���}o�è7 �El��xk�F���$��>d�3��7/���3P��2�n2�q�w)�tW\��Jӝ�s� +g�)���~.�x��z��=UG}��Ts7�Db�v:G۞?ւ�������d�u��]bI��P�^�7w�I��7�0בּZ�x2�7�k6�����&����1�O�E��a�<N6O���I�0XlxVHYEB     400     160�����~�z��k-�&����C���=O�3Q
t�U�����缵8�`�R�.�;э,Eh���NI�&m.��'#�d�@��l�FP�NT����JG#c��9N=�����6y����t����|�mf�e��к|�l��O0�P��1�j��f�ۯ�Aγ�dO��<��DH�I���f�ZI�����.���� ;�nW�wA��D� �����g�J���N䉡�"� ��e�8�I
�ÖT>�Fh����EFk��7��y��g�:��H�8n�/=����/.��R]�Rc���2�h>�͈��A�*�s䵅�[W�u�-�>^61��,��XlxVHYEB     400     100�\?aI`�u$�ɥ�l��Ý�|��AJ���U<���j\�5)m�D��o8�Ӧ�h��ѡ�߀����۴"�T�݆[ql��W-������^�����ae׎ʖc<��q$�hn_��ǀ���(6���_t�"�\�	 Մ.l��B��d��zj��/N ��y�|)���k��񱤟g��v�qN�Wͻ;�����r�9-�=�v�KO2���������w0�����W��d� ܵH���7���;�	2�zXlxVHYEB     400     1a0ve�k�b3��}1���Dr-{��w�!��2#N��t��@d׃Ғ�Bؒ��eI��}����fB�8�\�'�!���ԙ�t;~��% �^s��?6�\��H	�-��.`.�����:����p�]@��V�F�.s�\�7�;w�_����'O��;vQ$j:���;E.q����e��l��.�
�(�Z�Y3�+�@\ ��V�ʙqϷ��J��X���_�dC½C��( �`6��Ӟi^O馐W����������$}��o��(lrA�[ ��e%#�@�A������`�¶B
�uh-"-7�+X\fb�	6'��r��7x�r/K���a�19��O(�H%"��͉\t}_����v�ǻ\�Y�Ԫ=����McA-�rVd�6)��I8\�?z|�q�8*k�0[XlxVHYEB     400     140>A�Ć����I���=#R� z	��K&���`zy4c�M��ǁ�{�搱�-<���"oxS? ^�/D��X����1!ց\����G��z�G�WP�b�WЧ�1�5u���*+����zP�'�u霅��?
bf�;N�ˌe��3{YK{�_��@���E��1��l�
��ٲ�s�*S݇�bD��w�c6�eg�����.<<�B�9a2!X�7n��x���;��vr��p	1OeX�zR�0��O❻�n�f	���J�7�y����c��~-{�Ck����\��5X0�4?q��n��$Ti�Yg�XlxVHYEB     400     120��U޼����WB��}MG�%�8[�Sc�������@�0�z�k��.*��PI�K%("��lS��������+�O��DpQ4��C�6��[������r��Z�г|a
Uq@�(8IO�v]I;�N��z]�4�S�gKpz��=R3 ��)���X�i�ȁ�e�IEbz�+� �O�nJ�Q4�[n�̾�ႊ꽘��s��W�XYEF�"߂ʅ�� �hB-/'l��e�,f�d��jCU�|=^�Oπ�:qs�y
���g)�9�]�u�.��_XlxVHYEB     400     130�3������J�R�~�����Y��XHcP�ߖ5+��2��J����>b�K譆��^a1�]m���2A\�>�Z�4��S�w����ĠjG�v�(�������zi���I=��[��e�oz��˴��P'�:���˼ڲ����m�n�̺��Z���w�-�f�\�N�t��ץh�ds���4XG�7j���lg����ڒ��Ȯ�G�\k�����yЛ�+�m#�-��� Y���ѳ����D����1Y>F�n���q�>˗vL�9�e���~\6;��3��e��v-��XlxVHYEB     400     1c0������V�M	�u��f1>�m�gPyK��s;Ex%_��nTS���Ͳ�e���J߻P��Զ<����HCn(�cK��	�k]>?>d�qs:�X�V�f��ه:�Z��Ku<F�H��ld����F�h[|��@��;�w��B`��c
�ES$q�5	��Ȼ}]�D���m��*	��^�8�����=u���E���5yF��bR
_@Ş��Xl�&Q~��G�fg
���A�t�9�n�_��G���6����Z�u�
���B��h
�U�uR�D=ܩ�E��X�wԦu��h�Q�Vo&�Z�n���*��o>]p�h���P?_ՠ���J�-���	�9�c���c5��)�D�}5�ѩ0��ASOH���\���<�`�'��f#C)�v�*��K�I%�ԯ~Ò�!#D="��K6F��q,�IHr�T�XlxVHYEB     400     1a0v�[-d$'$�S�_�k��:)�ٝ53��=���7g~z	��f��ڛu��&5xͤ�%S!X�s1�y+�� �%�|b����|����ZԾg�E�������m�۝l��z{`
Qt�ʕ���4#|�1h�;���Zx!���x����樗� yf�|�V�_L& �s ��A�Hh�,��G鼲��@%��?�<΀���т��v�/������uFd������zb��Y"�- /&�;�q�':k@��p�Ң=qB1_�lZr�ַ���~:�F2�F���t�����=��r$�'�-���˺��T�<$j'�\���+Xd�/����f��#�S��%�����k��%��$X�����,��>����~�B_�o�f]�0�r��.#���S-�;�XlxVHYEB     400     1a0��n�:i�c���r0n�t��}� �-�~D=�k尧�JףV'�yo�R�����ɿ:m�b���՜ztbO��W.!��WW��#>���#���hf�KH��1^0��0L��I#�p�����e��p�zO�:�n�Im���h�B��V1ث~u�sk\fSdi��˷d��"��ߣڲ�f��������az��7�t#1RR��մhx�r	0�>���c*�ѥ�e9*UI���B��]l��Ԭ�Js�(��E�7z�4�U����4����H��	�7��гL��=�|���Mz�B$qdmc���[@ �r�6g	��'vlRR	�d�piv��[�u>"[���R���:L�<t�.)��k̕yN���2�!�M7_5w�L;>JuYWG���1��XlxVHYEB     2d9      e0����.e�e!��V�%�2�����<��2�=S]�dJGD]|<;z�.b'��h5���5X�$3�T������G�bO@ȕ�b�s4Tf��f"�/3eQ#@i�"ǚq��*�~�g��u��O!'9����U�_�NQWT`p�צrH�V���%s��ـ ��d�'k8͊P� R+�A�r`Nc�&:�J@'��(t����J��16ڙ�4��x�(�!(��