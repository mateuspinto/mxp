`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
tj4qxJILTJntTHr8W6aQS1/nxrtr9O1qC8B9yw0TI+27SVyez+LI+wElieujRCfvSg+SkOOj9DEo
vmntF7g5wRkwMSMCZHQs5tyeWAWvZ+nCbdgx+v5JdjJyamKgRLNJSp9MJ9CzF2UfBiForLgygVn2
a0zoMKPqiHuNFYazAhY44xf551CcDh9fJWCd9VqvhMdJSIivpfnAkHOZ8F35NY7Ixaw2FkncmE5L
yNd7eHFdZhFEd4TYtfLvXGb6K3wfrFRzq7sD7UWov17F8CatwGPDpcAbwbkRNmCyet0tmpFjZYLy
/8Y1A3InKYuh/fmyVhC0+9auC43H4nAzuaMdSrnexPRaCOdNWfXR8+e6seZGOJlsny8voeciGoOA
4NBEtTJyEZDXI0VBWQnbMhjxaQIrr4GeeNrA2H41L1xiahKDiMjuz2QFe+Y2I2KUv9syDJam9Lsj
NjAkEio9XEThUqvwpxPMkkX2jTb8zKG7/It7skYqbPpbZCQtJ3J5UBBDjSwowLCUQjoU66gOwpqc
RtnvWu3zyQnMbpJFysr3wbbGyyk+8BnGOSELmleMifI4JlyPpk7CJ7rqhC1/ofI2SIXC8BOrH6n0
vDgnVmsmu8f3cUnmhW7Pvppkspp40fiNvEphX/ki+vIJQRtYGPZlHeThdYPKU5JXVZBdnxyxRQDi
Gsbdvdlajt762WnEnzhN/4pY7i5+302LUGzgt8Gz0qm+aT62YSMu/auLrvoQLksTZg2KbGN4qTPM
xYhHat0TbUv+F2Y3A3cFDneB1+Q5HLXRro4D6B418uZeod6jWMJqq8HPw149nK0l/jdg6ds6jmcE
QGRGsaiOxWAAz/pKH53FnIR75mTKDkuGFKrOkjJZtuoNYLe5Llq4Dt2kV/BcI/Zl6mg6OyE4hRDK
RXZOeUqj+0D7uTBF2h5I4bZ8g6cbz8nc2rWYRQOKHFT9HVaPR5C0nly/yj8Uoe/Vdpubx4TtDj8o
PSPi6vnlfT6imspOLOmlNYdfg5kYjCMXG02b8PxSlZjiPB30mK1bQy6qXjdaQZtLLM4sTuN8zEU7
+sXe2JeBm8r9MNo6xsudsAyw5f6wIGZQpp2jPy1ATPdj0TNmIgKV0YnXl2t1ME+zMAtAVDksBEgY
AOB4fEDyztZUT7TTvMD+tDdotzQnv8neeWVfIxx2mkeJlkv6MKhFRj4F1gMMdPkM2/+l45/xrBpd
mnR+ZxUqgH31R4RGgl3EWJKSn/pazEUlCUJoGqQJMt7H0ANKSeyDz3Zb51T208pBmx4zfAovTqSV
ehXPfyV93dt+PMPql/K+JX6acgzVwVML+wUFIPM7iV/Jf8In7IEiXhYojVS8/vEBxpcCpAXn5mtr
VblEif/vdlQE7gS3V6cwKY0UUGIbVGxuzbkZe8ZVJAOD3/xd/nAIRwsbmte/v0RTavnWxtTE5GAM
yK2dEB9SE7/ZmrMbEVh5cjtOs3K/jLscftp7+ytFqIObkd/5/48+hLqp743cAR3/V39MJ7FcZYRS
ibbo33n0LeRH9BV+a9wMBM9wLVAlQQg/mYzJgLHfi5ohb9D7SXLZLYiMA4+3Q9OahD+362FC/u4z
1hNiG5si2jHLJH82s5/s7+mNzcB3MXw628vBxXdOtAl6xIAtose3lCodaDvJJV7XQs4OqPA94zZn
rBlljUJbxqTcqpngBplSV5kHupzyJ5l0lwalgz6pkLLCGiVAIfOdM3NahHKAi86gpDxtPuU4MjYq
DzcmhN+rw+Tn6ssJ5INbJj554tGt/OasMLgAKZy0G6zMJeoUumjHr5YQnMAwMe0MfJftGXnvqcgF
33eLlz0LjlD0pSpTZKm6yQ5Iea7Z2bQBmGu8Wm3I97fJ8cyug0RC3jLu8iVvLbtQptW39oVCXeYV
yHx9Q1WD423omQDOsFdmn0Y4zszEEO42hp6dxaYeRuZucTPF7hLsguPUpm5WiaMkiPsvOIjLTafp
45jHlRleWqT5KXxh6guBRsW/C1kxpJGBXpe0gIvo7Vp2cb19laa4eAkr3YoZnrXVr/5qtXE8sKzj
J9ixdbE9+xHsQsWbT2Qum5kyTkkPZXVdsb3jr6/aXSQy0ox27YGJBYULCQPC2xaTbP8vFEqUvfE+
MrXFMRFC8JUZa7/9Ga5kr4/JFuAA6QVGug6iqyR/fjEOs1Jcx4yJHsvmmHyJreYObPvCvoP/5mjo
jNhngXIaY890bz4ECIuKFa5ZoQdsrfuB8g/KYL2Q1Ulg3qiXuvegBW+TqDC4CVR+60vGBDA0TWUA
4H09UCiHNV5xcwN78Ia/Ud7yLY9+hFowxC877E0QmbmjqzEnLL5J8qKnvZJ2Ar+M2EREkOH6aUuS
+yqKwGqt1UKaA1hk+7kHFPTKmkaBNq6ExsZCF29qLymhW7XDR5vfkhZTGlfLdpi7+UaUJBbltK+z
1SJJTGsgfxUL17CA5X0nU6jk+rLpzJ9t8JUZ3etl6Q1LsM3PQkvbXM0cnsG1TJ4gsQlxuZRWOKRH
zsYO/Zdw8e1SZRmRoERhSqXgzVspmeVpZLs2hgNkF2K4LYnEcQ7YGFAFDpW4NbAaZva1Bu4S0WtP
AUM8Epi0UfqT5B76InAHVAYZWI2CZEYJiham+kpYLU4P1NhYbyTDDGWHMDkwzdcqXaHEtmXm96/O
YikuIdnO8UFtv6/CNziTair/ChCfl0t4UxNkSYhzsfaBIIzCbpukYAoNuBS9rNsfG5TY3Fh27zj0
J3Bi5m7jVBbumhxwlwwqwsgbSeWBVzHq7IJGLhZL9DrUUMllE45THAXIaRRsx/06VKM3eb9AQCm9
2PcVQnjtuqGSC5t5lmSO205mzrAeBF/il5Fsm1fFD2JilRf8bxockk/7XecWkVhUmO05DJl/Awr/
vGiF2s+8yKgmaUEo5G54KcMW6sCjlmPctMFN/eF4roazsUR36WueeEEqtt5cANJaAFPmxeFOSUX5
dY3b9HqpTmci4I118r60mB6vtJGca2XOzM/5JbYwEwNizIqVfZLBbhcWtadDlGCuhCEsEY6ohXOK
/qCPSQK8UhrpJNSFxeq0p2D3Pwhqu/W66YRuYOAvAuGEh2SGIgkt7k+dKO2kc8sr8EJRqjxwEbFn
catv6CLxROv+/+OffnZRamXImqlIf9UNGNBPIAoCzuR69MN+xsyKWMivsSIYcNMLzLvh9QIxteSA
6+JzoK52WgkPY9VkQdpSqnMhYitZ5iMd1CxPyMC3fc1Ax0WJqlTU0+HFXRXcIZ7k4WUE+nmUGlnt
24wQw9wbu3tEwuoj5rbtNmTnYYSbk1Vxge1vAX0SnC+09uhMj6HJTfJ5NuEDII7EcY9H+fapNvkX
/j/SYFhg+3aGLUpq5Slw2VX9BdrEyjcKx7P7BaretYcaSJt8jSOYe+7YJgKWLr+bQXkub+ZJA5WR
UUjNOrz4olTevKih2BIvtp4rW1ZijTZj3hI/DISMzcahS/UwHNkwRWk2FF1KBIOHLNf8S89OeuRP
zbyGPFcZhBmtCBod6nfFLs6TKo9XJVEUN+0FjzXUqZsza0qFmJ8sN+xDB86x/+LQamOjTX8aFLc8
ngEovbV6QDcaEYYsTKaZZAx37br7luCpHftso/ZIIc3jD+2nmQWBvt7+caDrsHMu1hyC64g/hf+T
P2lqDL/sF2VXX5JVshmoY9APiJlWgtrF/yVogvbkQfGJwohdnbic/J5Ob7xONJ9jVertGlcM44ml
64HtLouHgshiztRfNdyhy4XDworOaeaYvMKmNx+XdZV6IPlbmnq1MStsH/7ml/NS/Bvh1QTqMMin
hEDIBuMjLRAkB7MF6EyeMFd8r/4Ez8QbY2bAYXHQ6Q2ZYKrEWxOvHLaer0M3aXU8sE5DCzEXdMBi
QcxTAXqYwTE24J9L/s3ZfDFgttb2U5q2bCT9RXbr/ahW2rGSa3OjZrjK66skcsheY0OCBcqWtIJS
OjPVN2SJdpEtGAGdJOMsDl4/HMZxmFyULDxRT+EJUnWjCari0nfZzvu4n15Z2OSka09FuHBSxXBY
v704d1yJfBBCkWpAktAPNFDK5R7woB5EjxgpEW4IqQv1o4Z6w+BdBGIh/aULYeR8wS7uE+LFKVjn
QX9e2QbWCBdWOwtTbJ8LFiYrRg0Mb3PtPT5SinqGXLRFbkmh/e09+jgSF+3QGEKjJl3RalJfZTAW
ZgACIKAADAyAlO/3h9gsBmrIGiOLPHAHwGaCdkDzIAOK/OH7MFxElXFUdyKqZreYAhS+AdEEcdzi
wRGu6obg2q8N+eECnHudFN5kstTXJAltOV/o+e5XYlpbMW4AdYREkPwrrZC4cx4Jtyu7E+SAzFHg
MSYfDhGhqbBbbZma+9WT318Jb7G1lMNR+/VPDo39uJpwe2krHxcGikQCEK7MXhgztvBNWvNwH5ex
M60l+76TnsCkvzn+GU+Mx0TSpCWj2ky+GHI2QEWuiZhDF0SklUYVf6U4iba2FP56UR4JGRrfA1Uu
ckNECzJW5+h3bnfdsjAPDkEvUg6c5VwbkT2Llz8bxgrgu/oJFWeOCq8mfOeUsW2B+wxbPGNtBIIx
deYL42yem3n9oM11Zr+atYzFgmZk1Vo8A+UvtCMy00gcHeeHW3dL1jhmpRz94j6LZ6htikjT1qbR
jO4nz5YtRa8k777pPYjewL+0um6DtAJgCXABaK2H0vuaaQzf5kiZJsOJ1vRoM4GOgNND+53f1Ca4
/lvIHavoqZ2bgFsZdzqDhDoBcGoOAwh6DVrT5JAp1d9L1MmP9kIjR9wzoQF4C0alFVB+mY9jttmQ
OtconrmWDTnBlgNbRzE2nctWPRmPR5acTkBJdaHtrYlso2oAJLeotwHIGtOY1BQWdA+xXsdpge6O
AawqcHAdM7rmM5to4i1yVS/UCMBj4F2t5bKecZ5ysL33TEvnj/Y1suTNIfxItlXbL4BZDHtq+ScZ
USaIBAhc3a8dbXXxz0LMrhJdscoxJx8TTDTmEK9alvMlnf69N0tAK4lgY9o46GAxLIBIuB2OREXE
snPO38ssgYd2JNIB1MZzCMopCddBZtJFgSA2Yewfb6tlQtc974iQKt4OLQBzlelPvGf1H3ExQn2y
El90mFi+dzjB3uDz6yzo6JyUWPjTrNmSU7zsYRoIlyT5ZuwWdwd0f2fLwIF8SIx1JGXyJahEmgO7
UOGQ42JOlqdjrUhvcZGxpvA1qsfb6ZNBNgDQIKvq5PCjfHGONcWokClTo4z7BbKCyQe/8itwUx9o
QB/vjeMrBDu4VU0aSYAKw7VgHryMpr4dMC85+Zde/dPAPDifwRyJb52ZIk9Az38hX14kySQIcM34
PtJ1XfkTYaxnF7bqC1VSAyQZCqbtWgq7FbIg+m7k0wwkLGrHSwO1atpNLQlMamczVAoSx7XHAya+
3HlW1jEqGJySvn6+/bkHX+jnap7m8Jcj7PXjZS0kfGGp/R0xCYhbPyS787dMXiFB+qTuESWkGHpC
RBSCxhX9+kzopWrVqLWdWqY4m+4IUcZpQ+uEaIIHZcaRJXDTCxr65kRDB9LX3bru2CPOtheB2Vpq
tzlbtKX2OU1wO0pgG6+CEojDwlNthCGG2LtS6vC5DN1BvLJCe3q6ouhidX5GNkF3erjlkxl2AV0Y
jLsX8Pa5mWMiqP0gJACSMqonmIaUQ0xDpL0591YkcUVFU5gt/VqKbIXHxMDQEN08jyOjuEQEbTX6
yASHHIGsUh7DWU1NkcvjXbJI3Hscvj5tOiB4ucg+gAHeP+9qTHo5BtraHXnB752jjlqmbCNo6zKr
KUbCRy0abmOTxv1JQqYZrF36+5Sfnpim1QJ3sLenMR8rAJKSrSyzd/GK1NLHhs4Pe42wbsexblzl
ZpBfZwsMO+yb/zGPfb/Z20kO5u8rjMZiNhoWO4qxmh81AYV3bKAmmqEUZJ6x+DY7dVPe/KymP9eT
nuT7Lo+/+IK3rBdft56mMpCyWbWNrm/D8G1uSgLl3P6oawQ5QQpLMSHmEOKq047iIgar+ryzZANE
XGkWD5sYTh+7TLVksw3JIr99Gg6DWxRUDfs5nWRzfK3z/cloMDTJgp71yiagJ7/MZ/3tbZTtFNNG
CVwRYtGM+jJH8JPc1iGYmJeGikgS/9vSt5vEu5wij6lPuUaW7uIkuLm/IBAJH4TSVKkn8BQnXorK
K0G+l+8QQQdX5Ey/hEsQpEkYK8HozxNFqetD/sKT+EFzhvKvtaRINgCfyjv3PT1S7XGUhp8F18Qu
fSYXNZoagxjBO7s2gjVaO7OqqiY8BJUnPjqwR9kzp4TRwijiN3J9yw0m5oS/kMEbvtBdFSBe9nvM
7vWhq/m8fxnowk5e9CbfD9eZNxpUYevzKdczZ0AXyhYRqlErVwiMc3F3LJcSAOT+7C5RX0jrQdHY
zZFArVN+oGesm818E/4qhzYDV/tMhbUee6JoWAWK81WWPu6hLi1qETkekE/UPHZElm8VGhzgBa2e
MFnnwmoFFlXd7gg38ttiszEnmoN8P2R/OLXPRK1KMq2BuMDXU0bNEF/xCu65WnsgBxVxoAB1EQAL
LhZ/Ud1VpN5/0Ij7BvzivIHrp1khG46VYdvDpI9LbnVBzytd9ztGNL1KD0HCeER2iiBmFEnK2sf3
7bwDqI0yKUkzMm5M+JehVRawVE3b+cvDnfMnPZq9WxAIV5DJM0jJ2xV6NKRHvfLgRKk7Mr9dViCl
1+Ru77qc86eFVkImV1yaFDatjdZyc82arnp4kSsM6jsblzyg1v3QuSgESoT6RSPa4aRhvKgYyK9S
PGrSNXHqC88/MpomB0j9m1PjWbL4SzsJYYkze6IIgvbgOYJkxawVAxfw3SmvZGgpWHSmHxzEufFj
FTHb8NXdPhlghIcnaFLkvW9X3rVPT63uZoTn4QmptzzinX7MbIJJp0AuUUw7tf3bWfpIMJ9kl+kZ
88EHMmZmZw95NXqZCdKCeojX/VmYL7+aJ6UFqNP/+H6X3mxHXy+nLft1PePq3iWHzKDWADzFLqTe
H63OzaEcT2Q/UDcNbMfBpSAHL72jeVWH/xK/AJTj1S8JAHcIDeiPQFWbvh454S0e7DJa5pWUdpce
SdqJ7pejo6wanYvbw//K2Q4cpUHIQskSJx3P1Z8ePp3u/fEqZxVGuw03f5HSlY4gFjiBkzNKw+49
mWcQoP5ekshT1oEjxyDmJWV/ntjy2dFov1KitfpE9MZ4YnpW97Yz95pn8FnrnvG1N14TDO24Qz/c
NWj3QSlIRy7i+nFC2s+dJNQye/v+2Gn70s+hkvKlz6VYcjKJOyxYl1JNasMuZ9ulj0TF8Gj95dkV
H4h9Mv8wYR0suLtTmJxp9dKo6SN2YbXxc2APWYBVNLHnA8avujD5WsTukhiwh2AbDCWTGg1dZR8u
XYOpJGA7TiaANRJ/p2iXgrxhqgXXMzb70lRpKDK8Tkfvu0cCD4CtgcHyJGqRi/RJr+DTdKdkwMQ0
sZFvEnzkLMCrxDf3/S2GaTBHi5EY1EEMCL30DGKrkvrHdLohZYJSBoTG1+xMIw2eZfbmSu88rd9u
FgLg7+sfjUuNvXto55zci5OJGoOH0AdEcdqFpbBYUp+YYTzyMECRI5Lyn+bn0vOpg3KzZGLMwTIZ
QAPDpSOX5a9RfzPjzb6StZP59pP1N75VR97YuGQGWON0pKtWhxHcV6hNmG+/kQpR5EpnwH8ifLYG
dVWJam7MptfaCqguV7zCU76jNAgVDzWW8SFT0ZCdKYoxKUQ4JLIqW2Otzp45B06BudztMPQ/zEhN
PvSmojzGh+bRXJoaMhcDHl328qWB8G+cuBd76Dge0ZTJ+ZXbKvOlBOKcupeeGgp69Ps6QFYf3Tjh
guTqx7rrDVX2FwgYDQOf1hwMIsk7EO2g7D1dThTDs4tsUarLtD1Md1K4uRgzonpnUSJ+05xXSOx5
/Wd7eFpcHLAxM7i4QnL/5QKYFo483OMRgsKitDxlqMYu7nO8S9oqXZfpoJyMqXOg5UX46ZhL3ufj
va9oEZ6TM8T4zNJCSIXeyLVr/5EePBZOW9ACUwYrhtCpVJban2V9lHKLSpNQE3vwuHGaFuFczM+A
F8PaAVii53VAGnzU7M/u18HrrofQbIx0/6azqLbOn4rlWY1qDfs6jIH/sbcNIhSXY047AiXgYL0u
lJvTq+mCxhpCL+9krceq9y02t1DvMJdPTmRXS9IVlh1KsHhQwCOE6hl0xSfG8r2KEkoDgoC3C9DW
KBKq2aXPKZztQvVtCtQhSc8ro96exv0aNn7lZspucXLdYCZ9u/0WLUTe+DhN76hFwfijE5xjMGOg
FM6eHtleRTFE+KV0nCxN++iJ4zmXIO9Q/e9eKntQCLyTu2Y23frv+l0S2DYaUatH/jq3h0vTU8lR
mm2maUsMHqC2wog3zkrK1X3XJjfJY/ct1Ynw03tqc/Y4efms34sa9D0A3gKLyK9pfHgxSuUkxZ6o
s6E3AyNuvvNPVGWrBA6/+lGfnQKjhN1yjBnSjRNX/Th7Utr7dg414hs//yxntBe44Qbme/0wa83V
xHaLPsBflJXppbqGB0U+ZWWs1kd9v+aEnyVqoKePZbd3LL30paVlPTvgN3DejuT4pmmdMGvzpNbc
vYSaNzL5H5DVieivZ8f0XhVBwLPeFZQL5u4JsdumJ/QEWXAnY7L4BMWYVMXXzYEWkHsQD59ZxEAn
x88hGDoXYDmOsUoRTeuOS7pykL2mhoj0Vb3aHwVak11tLlgOO67sSQ79liicCQQRno8CU2MtuNXb
t2Fz9UGnjdjdj9gD/6W5i27Bw4/UggkFyUgB8CDQ9b6F2GbNwKccBhivqqDLReBgdXuTmK1E6ZnI
AZpwv1U66f8Is5CSBSCZcHjT2F5rOETyP4cetyMiv4fF/P6lpcEMulkKAgVwCVDpMgRd78WhwaKq
oLZHSTXeVz0Nk83x9zbBCQC2mk64zdFL0yGzPTp+hjv2vPa0uuxlvnB72kpVw+1uJUh5f0wwRNXe
4eLbvp4sM408ysGTIjNk0i75eGATTevj770tyiCyu1mj9jcGG7tSYNlyk4paX3sixTaH/KhNL93A
iw3BaNSgXMChLGtBCZTLg/KeaG0PasZlcVXON+swXDcdcQs1woWLwcvh+CZg4WTDTVu8Jzi4TOD3
KCO2IIkRVyl94jv5rIB9RMy2TcqUpplqPowKYOBMuZ3lpYlMB1VKZAKs8ANWGky9/pqGpDHVNRb1
mA7nWJG1eidKW58Ut+u2biCbDZ+Vo2Q8LSy7pmzMRMl+jZLNLaRocIjSZ8Sv2W5TI3AUIrsd7Oyx
9UhKQQHo3IHMIiEG3zZAT/X3rpvWEZKMVi8geJ9h7QioZo/2SJsm/8F25mqYnNAl4Ams7HK+zCAG
M0/fd1MTHmCWGSSz7jLDoTuu7HY+2XaVUa9LyJLsIG5T5Q2/DBue2Rfk/dVeJlsP32AEFATHZmvR
znfiHPM4Ka6mvNe84Fpk7N9az1pP0eZIoB1WEa6s/RXP+XQ+lkf2PTEf+T642/VnhmdZemg3Yvey
qi4Rs+pFZtN1GK3SfA91MECUlrrorKFI/rj+sZ/llUsDHKomyOFmcXbP3nxdg2nTU8kjyrWZUK+g
x66srt2Cc4JWGaBft5zhDIAgQ1n5sYTWu4yC2EBUN9QRU3KRvL3z8gaErdZD2c/aH31ME/Q7mv7o
lSUBTII4JZKw4nycCosTYEEdoYLzwRI44KeEXJIEyPndT50/S45KWeVPm/NhrGBFUcI2vff/lTqx
9cYNyFOdB0VqiP7sHTt9UmOz+5Yt474foZTsKa/bxY9H6vG34lGtfyuTP5o6oczmR56zDId8rK+M
vbFia+AX6AN/lulDcj3ZIw/Y3borthV0IzRWeniERSMJ5AFkDww3rPYnLlB7uW7bxKy1yu6iOhp0
9KE+rQ1OXIxbadwqv4zyCtWb8qFaChBz8ai2wx36i3LTz57go/RFoFObzdKEfCqz7apF9GE7UuND
xSXyCaz4stTdRqAjMzKXxpA/s/tR4GgLw1ax4W/QjgD9xppRjCmZdMtNe1N3O+TK7QK5TnJ7KW7v
8SXqcWCgu840LpYP5hKncTLvu+CaxNXinpes1qiv6es05F7JuJeEwS6No3f7VUAWBz16yuISE76S
CoC94F+6p+vqodDU12dXxQcV7AdZF/+fEDfiTZuqsb3WcdA/+cAUJOzvMu1K2gvRWH3JJ3NcMZAD
3yUR2h9gWAcXcr8IQBXoEJ58SJprh0yztjRPab0Gx9HIrrPbERQ/cAL15lnvigbgEkNqCqxJdKON
oopf0i/9qJ+ua6fSGKmqBRw8fIUfiNdmu3s4ZgJr+zF+WpTjTj7DlsiQHfgVqPc5oryRaoz+vdMk
r11YUULtkjrp9sddhQYl/Kq9/Ztk9c7rNm72dkyuhFHGuYzz9Yn8i/dAXmn7MAIzvcXx07MezBkN
MLVXoZm5X6GnC8kyFX/3BUmbIZpxEH4ghIURDCYAgsBYmY6nlmrFDXtRTM1w80yex2En0BFb7KaE
epwdUuQ9VXMVLPph9/WoABXVgFdzPUL0vnbGSFnUVmPSVf/inVPDT5ahflLqbjEBuAShgk45rkoW
dmm2ymEmmFzmqbpGjqwQh7d6ON/ze8tGeeZG0Pvk/Uq2ZL3vV0xpGBMihqIBxSfAyHIKZJ5ulAnI
6T9BuMuCcaJfvbDwmrKoZLCVeTQYn5P8Lz92SRmpA3rJ2tN61y0gFh3Z8jfE1XwzzrJjiVYH1aLG
rPvhniIsiZBheLC//kTnEZ5Fqmg+EsuOitIiJjkRfbfQgXFn4or/aWkHoRgAnpyQDPlwTcHY46Z6
CoGC9HxiCZeJEPOy+QlH5rWN7CoGxqHON0VD8iUOwBmT0P8iaB//bCvTLaifNTIqclMkunsP4Yq8
qpQF7GPCScTH6ZGhh2Qe3LEVZgSX+Hc2Tp4fQnF+U3qhWEJA1LTGuw2B7G4bI2Jdqys9yi5sdiEq
HJvT/15zS9+MTPePIsIHLKPaQspxlr2j1dOUFEx0d3WCMfSev+kseYX5YAwi2BJhhrc1PdtIhiqk
ckxYBW1ObaMj94A+ld6I5bVTH7UeSW9oI2r/uX8SatvI4eS+tuWmYr2Pdup4AsyLQBzl8U5yULo+
b3ItkH9uZ2bNlcoUEM/BwXdZvzhR9xDvnP8CKN5Xp5LiHO1xINGbLqCS8TDwz2BhmMVZxWrvfqOb
wa7eNVAgQf2iR9QDL4mK/JuQFFmms5gPnrsixJA7ubuPPnnq35Rjef/209CENqMy4WZaFxqbK3o2
H25Osc6cljChEUYqelc/VqDvpQ/ksDLIA9+FddW1CiAIeLdoa5kSit/glqE212A2yqB/uJ2WLZR7
hdt8EVP25bG2oQyoDvPr5qu8WaexUz1urFxpR3BzquuLz4dBA2hSH/yPx6VlIh4Yc2rS2lnfMmdN
LcJHN+u14LVOaxkRAZaHMeHYn2FaJQwKWc5NbDMjtIyrOmf4dAzSWA/lk6I/M54vrT3ALCCsSKeo
dZ3ZNwCwrVCEbiE6p4aitfh0e4MoUVmx0REn9ZNtH1+Lqm29R/gqhoFeWdrDOUAfq1TYy9x6E2QS
GLjfdvx+x/HYK9CdrkXDwDkvPP0QkI92GJjLnQg+J3HxcgUdJgHzJuAwQkMl5tKfoNJQRqTwgMlD
TNzbx1yMPi5t46xvzgvc1DdFzkosQ+ifrOeSFrdobM63OTuLbZC6LD0WbINZ8JguzXThq0Vv4F2t
NySrQGC8du9aG+AciJ+NnDA2LAOU3vTKusSM9vsth5tqMDlRFVD4oYbWjFskKRlofP+pdRjiipQD
e9bvB8PlQEw/YARNOcKzxYwJntZ9lAXJLd0rnPGQFWOABT8wj/00WcQd+MqdcRNDCvIulrMnkAha
gTTLh/Umb7uY/+RD/DQ/4ID5LbdtnYPPqmvq7msqNCo0IWaza+D2zPN3KBSiDe9R9nXNzjoq0JWI
k/DcQ09+gCSthj4WBsFLRDxSIxlX0ix77E9YbXYI2WDzsr97wAGGt9Tm/gBHD9abOHcrlNSUNbMq
q55ULDwWFhsE0yXkJlmWpF5Ms8M4m5p6+CT7BKkl1VzZWEQ6PwyvDUvAiJCDz2TlwYEyt/el+YJH
pWbQid+SYt6CHzSl9NnCh4QqG4CG1l+grUPLdVYolQJxcZaUuCwkqrIMoyAwAJBlvefZDDtGn8Jk
C7d0UYV+cATNXR6b9rjqC2wY6p7n0KFPDD1G89pLkqVf0MOy53C2U/6KojaXDv4o7O1Edb24cYvb
LrAqDa3slhs63IemoVcMLH9PlMcoq4pR1/EZuh1iH3CYD6CBsUIdFGvTOlDJiW3tVc9dYwKlTRuR
giGj/vhj1kQKj4bua0gn5dJY0smljyBlkdy8zGS85n9NA0LawK2fq4xHTKbxs76Y4LMUYLvUxLjb
I8ymSAcoGvdNZsP9XFcWjmg7XgIRvN8XFxq8jKtmS+wK5IVOlgFRDAv3Kw4yUEMNrqeeCYZDSuJF
PgsgmMaen/i1PatfesJ4wmV4cGxNNWicqxzimfZRUbQkvLctQy2GZ0D7Ed/E3Iqre7dfopzzht+p
2aj1tK/KfZI7AN5VLOpzregeCpQRAC1NLTFgArZfU0UKm2gkDp8w8BMEodGCTfXp5bC7sen7hKVH
4mg7T8a/sanzlN2B+wg7UVKLGwO0L4RPMktMG+P7aOqiH9dWsrjfPFPlTDQJdzZ8Acbmo0o45Wj6
6m2SB1pytt8rt/swvVkpIhPFdjeE9yj2EVUPr8opOR96dDQBVZUhPMjNng58BDqTn5pYKim99pjD
4dzKGKzpfUvE8qmnYKmJ8hkO9vfbYgwyFLfWr0cJ9GAkIglRSiZtwnoTTNmmfdHV7Q/pbiOH9x8X
TNR8P4xMZh8jvel8ZxKT7gCtLGdFF3vjL3J8zCX6ELlp6xDjt3J+idvWC77TE5GX0PN3GSfoaoj3
t9UfUImF8NKSbrU3twyZ3B2gKqXs9/IoSgL/0Y4O6+9QItKts9aofgr2hylZr8T6AlINTgJz4mca
mv6ivfJXI7wYQ7+MPqm4CWfrov+F5MpQ1nMQcJMLA5ttn1s/5gQamIt6UgsJtymtZEmk0ymxePle
EuchJfd7AdkJ4mwKMqFG2845xVVyOc4XFvOFpMN2477MUKehhbBYhqUQiGgx5tL7dIT5t/bHz1ps
NTUHFUSfo+L7d8cwKTmos3Ym5Rahhq/a3oMpCalN56VQdG9Vi4on+oLC8LOE56l32c1Z0jqxkKdu
Kgd6/VRqBzETrtYiYzLZo0u0E7M2T/jJfuCksbE8ssHoGIpdyUShYxMWr/pKmyf4KdCq4UHQsajf
1EYirI0lEcOrO8+SqtOeMwXS5dG3xcfrU+ogCeFDYAOMSuDakW8TCAO3ObkcNUY7UOFZy64U3a9Z
s/m+10yLpLNW4bKlJ9np/wjU/U/sF7x9KbnyfI1xpDiS/fWniRlHxWuY6RojLR/yWFJ1wgEb2yjR
1fjjvw/pZkJT5AgUU3sl6OGnZwR9qItJwdejApiXbW3/HjH/Bb2WNRH/QFHim9sI3sZFE4u/NZAQ
FGjY3GYMrxp2wzN4R45IeZ+hGw9qOdne9AolI7ydlZRXuGbrbJG+4ZMONFpqBLaGyWAxL5snfbI7
ThuN8xd7fhhnefmQYiKSmDmfpJK/twpm7N84I7Is2ZOV2HIx0xPhXDkjSs9+K9QDUy8Tl9UB9tQd
yBA++ds3zgpGO/zzHctNT6jWalVNC+PHiHLKk+2u4dYcJr3picIYHYf8WI0t3fgn1abNt9HvH70F
LX3R/B4fihbHpLyqOkzXlTV6lAdRwl85cmldg7hlaAF2Dn7XFgpA0uDJxEoAsLFQUJzOW466bO3W
ZkRrvm+UnsjkvxiOe2+a5lnRoY6pAcL7KsIYgIdNf2IEr7IUiaU4OfpWyVwiNSxpouhd/GB6JfI/
WistBN0NzQvCGoqMnDDtIjqEtcPi6fHMANU5Oo2UUi4LXPc2u4pP1pABHtfyeCxNTJgsuwB08tL8
UfQHQA981N5/FuekSCavXtNi3FIWiY31irSfgUFsnGmc6X3ow7eMU1hc4bXgk/g1zQf4/1nOpAUz
HXGMmMWqopz5V/EW2Tv5M/iU4FTWv+HUgkDXMZHlPBIDMBIXYYHNPVZ1mHD7qCbucpROEuH3+vO1
63u+xYy78qGkvzHyHyVm9HhSQqAf0OHxBXRW1t+3d2saph9qaNm024DggtCWUl+7LOp4uAOIEArw
mjOinqbisNeAeG2VsVzHsv95xf0/71g2x8u9OP0qPeoNFuqeTMohmhRjmqbIOxD09CJRInfWGNNw
cwM46srOMrkSKIheQfimK9bB/UGHMgF2Svs22d2sZcM2V1QU0tgdRK2RgwPKG0HXExOUZAL5AJtK
b9zCPIr3NyGPFAyWSFLkNiKqrxZoSzxsc1Wg6wDCvACgwiE96VD8/cLc1PAgzjfSJGmt97/OsnWB
LYrThEiAesk5SqMijO3bBFJ3d7iu3fBW4fLC9qihs9C0qlGJmh1q5/27nEg79Hu9mEDw0YHGESka
xmNpioxqLbbDIXjk91oHnwX9JQKZeifl718EB2WaIBgTvmmxkpBGm5VuuWhpYe4OW9XW12vrb0k3
PO2piehbM90YZQENW+SNXALarviCVIixQfIcy61/lzC5cmM//6CjfphgnRLvKeB1gh9HJTwipvSL
8EqRtmIhq54ee2uXPerzxEBeArS0PHe4LIp/RVwfzULcwv5qaM6HoC02ii9evRMi2WvETF5vt17U
oQYqFCgtpZG9DGyvmPIN5vPPRUhsphZ7J2CF4HfPZLV2wRXSJF7WfZ5nJNHyWCVQOIBAf4GWrt8T
HRI8Tfl9kvYWjHjsJavCp5V48O9pUBgvfj0wBTYJomiszgXCSDKB1r1wuPRYdPYzw8aOO0arSFkW
bfE/pimNWoXGGR38P3ejSrmR8HoaKApy+Jr8Xu+YZHDvKchlio9RKRjV5ydUJZNuZULWI6A+3Tis
PVLAubZUSB6PKBAImzMqqpeLQTeAKYMFu0Ihc1ui0FQqWgplfjstO9EsdxjgrBQV1cJCCNnx/sjh
zF9cf/9uIILDQiEXvB9uC22fGxwr6QQdBMmzC+Nifw4WF8ai34kNWUGBW1ZRVx/KDeCkjymBuUya
YX6Xds1TnOea9jw3UTkiybgAzH8iQvlOZIYdFjKwmdipS259dyuNxfpfNe38ZSn/RQAWlyZtZL91
LAirH+Cd3ZPHnYVIYkPypxyATuYMi2CeAL4aGCfoznR2mHMI5i9ohBg0qchuUC4258ibfb5Fs8K5
mibYIhTNMo6TBjw4kIOfftj3z+Msiy9z93Bt2FwrKrwcHZYuKoeqmbMfZs4/kDJ80YM+LtpMKhzI
tr+db43CFTr8T72iIzv4IFBHkS9e1jb5OJSTA5/NhlEA0Y233cIkF1B5zn8r1AG7TKe0LFM6zS5V
kpDwqYvTuAL0rR2czMY/YizxAZQqzv+mXfoluDVq+WIRYuTV0nQkzhybRdnFch7329VG1/ETPVxq
59VH+ZTHwvyx174BAOE2zz3veorse+lvmg5I55LLB4qrghY/qtItRKDTWBYAdNK/oO43fqbgL3/3
ewEmJ7pi4gGsO/tNfPNgY16fHP5z8RHSBAqwLboVCg2rnYSDiTmC4qm8rA5Vg2637wkGZdqRRCdg
mS+6mD6c8eIcH1Q5iPrHZMJbMgiJBDFutN9XFJoStnJ6YCZ29zR+3AiA78oAaJuUGSorz+OL+lAm
+LHwZfFiwQuJQO8SbWJ5Jv5K9P6Kbd9G5Uf16pY2bR58TuJt/zCQKmchH6UKAnxr84DlvkTNQx2O
aK2sa587ja/u3kh16PMMS4dqBtayz4LbmZ58PMYjMSmTCAvg6WuKexYYHJWIPSUfKszQe3RSeRVZ
327yzaSx3+ueAVhsIHnLFabY8ojm9cVMY6bCd4v7HjEeEgSKK60b+MTuOgbHdsqiWoYDeTXZMXAV
ixQp7Euo2BP7msozJdZeimwz6zRC0NSbeNBWFcMHDX/cF2PD/BBWMoBCjkIedLPVUfLR9u7GxCiu
PzNqdHPGZn/9ykQeu+6BVSKYSKPa1UZmqycMHCksS4ZMCYC9fudxGldy8G+Iu4fz+AfvDTKpOWXW
kKyNW8Ho6Uue5Jd5Ws+QgfsYR2+x9x5YfhKTSOL467aXyBattkLNrGydsI4XDAuQoe3gLGEpkcuL
/68P2VyD6WkLn7hnCUsNMW8XG/xvoKbLe9+i8pW6GWKBrvdBWCDOsTsL0Uw7TAqIKuke7qDUlYt8
1HtdawEM/jC/M0iU2XDGJGDkJrcQfExpQnxyBVDb9r/Q8bX1gfohAQf+whHjyXTRzXaJjse2xDg4
Naf30eruXckl7obQJzAAc/9YxKGJF7RxLrMul8cFF6vVc+KHsMSmU8MXc1f+6/Tlxw+e0SCEiSCw
w6SZ1MYnJk9naBOcnJ51yDmc7f/+c5t59Vl5Vzx5EgTTvWhOWP2U/WRCXvntCP9XK242wEytcZcJ
RtnM8M2MkSFErfsSoKLZkfofvsEgkTSx4CeOWJL4RLYdlRRceuZ7a2rPp22m0A/Tm9hgi8/WImYl
mxR/Z1+rRM1P9hDrPWINNcEKUVnmhNWI3cDXFMD7GLVgRJaR/iGU8uMUjqJorN4rgwLhD94owLru
QqkrJYdR+zrEZNlxmfL6Snc7Qsle6FHMcziBtOq9cWbiOpvMfTXqvp4Kc6htdNUJZUOLwdXnfoaM
cu66dmaihzMAapzZ8bgSWkTMCDcks6zPapV+mCl9kvSuzbAO2Zvy+FhDQRGwkmbfpaXEReCCXmit
pTWgukFfAAJTeY2XW+DTrI5DYDdOaT1qiMoRCUHvG323qamGlTgNz8sfjxGvHexsAUSP9r8lIB1b
N4re/MxsxMqhVajtVNYokuI8TLH1uvMNYwCOT0uyf0MZAISv0h1ycMQ9JB+EF1pBtQPoAMvR19ah
KeE01Amkozb437AhwfHMYyQnYLPBkGVlDz43bG684reMgJz46ndhZG4tVCJiSLqt+PGqMJMj8YK8
+fcbOhZzh/UoOtFWJDx3kzgXy3Ei81fPISSxg5VzVb3+epzzEvvFHQwLvR1hkuxPadbRVtiHncyt
C33etGOARdz4J7O/++MVbqeI/3kIrh9an9cQQ+oAno3dmVG85dIiks5PEsoSAbExUSmxjhCt9pwl
KsaLHoEK5Wy7ElACstULCSnGXfTPn102pnTprOkrFs/Hxyen9TtX88QKPLQ9OmForQtLvWdCFzbN
uqb3nKu66D+S4CgcvGe22dCe0np6GP1QL6qWFy1IvRhlZt0+odBlogAkfbwrViua+SW/5C922MlL
lSQVboFIml9fw6u4gHjawtu7OxTRcURbBzJqPt701NxYOoblRisbdATczO1lLsrqREq9PS0iwlOP
AKePod6XtC2ke+3eBul32VYF0+/TF+p8KPSM6fxmQKfV1loX+R2eHQ2Pkmpiyr7ccBbmUvFBU8Kg
/LObIMxO6Zdz2t1pLa727aO6ewFvZKxeBSmIsEnATvOC1cSfgT//8NToRJ314dTrzXwsy4hE6WSZ
wyiE/o6Pznv/CfLUZCLRzh1bG8yhYxFBokmAAsxB5/133zZegFNwXKHCjT1jwM4rD2OwoT/RnrGh
uZe6J0V3T2Inp9FCffXM+IfjyHXlgdoZp8m7LljF5+2pDktVTyPWyKPMFDCnThPVKGGCsVgC7M9W
23hpi+cc9zt/hmpc2ujyTEr0K2OLTu3XvNltNtYz6oE7MSp0wxSxsZHJRtLnIFL2XfxB8/23vzmL
YFVJGvs+CYP3txOQi6NMgz7SR4xM4SkykDBiQOGOHTj4O8JSGAoO3SG4Sv8Z7HA918vP0FSv47/Z
ntCZlGPLAvqGIqRC5TjzEW9muifRiUvjVwxvUiQs7VVc+h/XOm8YFjpn82Ca8Bk6yk13b6zepOZ5
napLnSOua4ezZ+boUXwsnWSj9L+h+9cqcm6Qbr8V2MnPL9RR8ty8xHekIal04JJSJT5acPdggQZI
8/Sup/HcGfOG6ZEINUI/Gf2/nxEGoxF61fftIfrpu0c2Z71COQEQu7jqz4r7FFmdAuO4BEhe9qvL
QlAbDi63AKFuPgt3M5R0yaSwYNva35VaNsnPpv+3Ye0Pz1+k+cZMr+YbnZ+rGCNmNR1VqNtyGkAi
+wwsGcPoAlkhGoujBBDzFuxHfU1MKdenzLHYKXde/d6U08obrrWFagMEKROIVdCJQ2PLRtPtcFoS
mC/nxCwnDr3LGiD3GutyRwXIFFKSuuAdzBbqIeNqagoQ7bJUFzo9Mpwoz2RIfgudvvvFftqE7EAZ
ZDzdZJT4YhCuHGDBZ+4oxe3oXJNWU3Wk0p4eYep945Vz5J9fA7iprey71TXGXJyzTR/ZhvGa+3rs
lln/qkFOuiTu2F4BCkNTqYwDz52xJnVspSfNBPlSa2ov0VFafUaP2lZd4aL1Hn1ntb3SSF6MUXM/
gOEdX600iFsrvV9iSpLvl8Md8oeEVWJueg54MWmwKgPVZDydyl5DjSOp0yoLDBJVjX7h8QsB5HUk
JGOBOB5YQe2LMpRrmzL10lxtPLMCzHfbfxtDdKX9+VU7dtOvrG29L60X+4qALIs4bfJTgkYsEOgr
kSP8QlMcQUEaTh/af8AZyHsH1ZMjV+hdQHxpl1hVKQ4WcFwkpQDeomwRWfP3Ht1G14XAIwx0OSnR
kQTeM2FjmvLIslpDXV0aXYc0e3OGjVe5apbsnUxkomH8KZs6YFPFXkttvKjDQgYEnURV07tX4d/F
B9kIfstltgPPZ1YoIEUh4pQzbDgOyLzNRMvj4WB+S/vz1+palWAD2zDlSYvlG2IH7brd1bmZmrzY
r5kMOUCVw8B8IUpXhFkA7MaAiWjKehk+Bk94vGKVN9csjxUfNUgC8q3Qf7QzTrGCb0WsYxiCQUEY
PvbTG2wbVyb31MqavIQJ+/TuAC9GgDSNOsPp8+H9HbIl3g80LaW5UsjQ4aXTD7tqFjinlKPebTvB
SFZGfDXEfc4iVV9rge1NBGQfGV177HruoO+yMPsKWoPpav5762JAHlpAdmZxEavJ9ddzVHOSchKS
raYiG8E9MnIjTIYV4kxezudc4MH8HR4kgqyBvYe4U78gVf0mj81k+0a7mvWSPBM91xoonkmX0Bno
oNoti/4anaS3exaGxgNezlvd2M7d/vCEmGN3wzQNWlWUJWLBz8VCxyApLxFoT3CDck71J+eGR2e5
nFl550LwCduQKZQuPGIgjWOaVYmhSKkH+cDeD2cG3YyqRc1esYmOLwa2oX3JaoVpy6UTSi5H0nVg
3DJI44izUWwnYZDoCIq5YDs3Juro7C+r+u+sCyhc6VtENUnukKpBUewGbeTLfKDg70ZNd7WT9iJW
Yy8NLegcFEQyKTJ+xnQVTKwZ28ek8AvkPvM5vGNvQwQ3HVkGkg3WmnT5EfpQ55Z1WG08x9ImWbaM
rPw68kGkIhytUWSlfWetxWdn4ON9LSZeOVC7ski/ybgH2Ij/+2Clkfy27cX2HU1C0vpPtbCYj9a3
erDBvXBA3vWHjEpjvwA/ti9pO/vL8AqXKP+Z/QEIYpsJdfMHacPFhlxkIc5PaWwvKg1BKYU5cdnL
rvkCYaxqcJCEkwswiEVRMG0nlge6JQut3cp2gYxum5kGe9lkCVukyVbbDHULkxAuxFJFw1mVyFOB
XRMOmLGtbkcqWLDfY8biq5lf0PmhbKid3keZWqad+QfHcAA9Ci13qIgl6meK49PYIolkLRQNmrGO
tYO+EV91Oo4Ckb0kBRUFIOy4Mf2mk9irQpiAd8Kn/bvfjgIRHzl6Rzs4tSS83ga30SVKt23Y3J19
VATTNOJz+1wi1UpjZ75h9t/uoRxWDpu/g5hg7FwQiRVlCtuoFiedsjQt4tLsAr68FGZfPI3bBwyP
HP/KuFqX3dWn/wlxetcIbaexwECc4Qkev1hDactoxddagNbSDkw3oumCJmA+vuqKlVcRnuu3qnbO
mtFMHYheaY0aEyHxEnXWqReg50YMx6Tx9nVI0/pLQnDvUNjnLjIFIkOg//dhE4QXWaSfdGLVLxBW
MbCobNAY6PeoBOt4OBsqmltwX8ZzNlpHE2tJszuzVxbi2I1h8SFcgddrXMTD8l37GjbTYjmGqQJ3
0y/VAc8ckgmkCZZFmsQWwrFxyYqASHggCmp7ubRkY2zOcS2YFami08y9zg1yWE1EcL34qsgwO8AA
2tOrzyYB0jkqkDWu0KGkrH2AupTWoZXhMKFKS4gmnwOJmJFoM6OgTsj/lEXyIf2YuIUHzNWVByzU
bmQkQ1FjZ5+7OVdgr7HRhCBvHXid7rxwnTRDGpoWDxkZpocmIqabK/406hm8KUoi4CNdLV6EhjNR
Bp9ONrXvl3EXibdkcwEv2wlWti3atCvsC2Q5N4Q0BxVJfCY+a2nGPWGZqLNTsEqqNlLWI/DJDL85
SNcwRJM+0u99gRpzGT4sGzmAdRI8Tw6o9CEUin2xWiBeigVJXbA2iPgO5Bn6G1hDSWDUoexRGxDj
0f49LJi9PxpGoHU64mrCVNZkDvlN4CXdCRiVcKB+4GprZxieTWVtC74isRI9IR6/RcpDvEqX2Dzm
tlpIVFdqIsDl0hztaQbNI4Y2PzsHF6Iex/SjXtYmVLtxvCOIFH7xQJxfaU8dVUQftcr/NQTbWxQk
zEcsqrWQY5hH/DMuJcw23QnNdCrpBtFIrTcqeTIbeZxvDxUwqd7aR72WXobqw2flTR8lZXdwQxE8
+LXkFhwuPFeps/QGaqyP+Zp8gXtfmJi4hdNSpI0MCwCnxymIR2MHHblZgq9jjXv6KTGc7L6VrG54
hDlI0gifqLRXQ8bMpMLKHGGwQxEkvdkpKwNTIJeF52qRFRp5AsUbAJxGn1q7IblywvOEpFgFmMcw
5jDzdruv6y8OfFjOUFP103k4n2Wlvn7DyM61Lmg99tAuAANsg8Tm6Ibr9wh1D5fRu9MlnufBUEY3
IJNtJ0ngAzh1mWsgLawdmOd2184qksEaFPoFd2a9/wwkVpIjjIL/GbQdfvbJt3gEJwM3tdkOiC1V
OrUJLv58VHraXV2rgkBRIrRzKFxvEasls2w5Niech4OSWOn10ASbkmJPK2oUK3vyiAnU2sS9VHKy
xIg//Y7JO5dfOtj4/w7l7WS7h3+9meeP0vcil+N9fSn85X/sgUbGRQJp5ju8pU7ybLhWspBkEoA9
D591eEY4dsurVdSvZ5qkywtjwB3zZCGpt1kOqRhQxTK+YqFnkTH5eocoPg6daPfts21y9wgwWCoF
oacafSVO89/KEkBy3wRwSs5l+3Y5vA0o6rKfMNe4xOJDMjk73v8sSldvznszhwpTAC/kWUpXalwH
fiFz4zU7LVmqPKH4f18pQWHKyr7EfDUsGAZ6BCf390/xoWw6Sw4Rxg+AnYrek3OrqQeGo+HbvGAD
Eu4x5GXw4IDvkiVvxdhYupcyAl6kor0rPFeRr/aQqkdO1Lt5KYZp44BI2pa6xZsIls+SeEsxvr+0
fXU1PnpibCZJeQkLmKOQ9dGa+DAh1PXxPv2+Rixj06fn/Mf3YX/txlUcPmXG7VQGvSsBnVHnDVzi
DM7F4eQS8yd3YaRd0vgQb6YJtBK6Wfn4f87cOEYod19in0xrxxYQhU5PbkzdFHBWzWR5Ujb0dy5M
gJpnEgf02sh86ZpneCE1NeO8nV+FRrhRqlQTJ1iWNBZnpNx+856aYen5s5sMii8vElwqE2FkoXRB
3SLDq87rh2k8TS76hfN5I8PJ18Rou1R/B+YxWEHQ83ZlJ2PxcSg0IT3y28L3++i2fggngnQbFGbg
AkVkZIdl0pY5WgX0OWQoAXXP60QaKrPLIvwwgXeDp2gUhy6zyCB7ZLQp9enlUnGgEsa1g74GC/2I
jHnlPDoOQ1WWfCeYH66ZdET+/rl+ffBdN3vP86lOr0Bm2M4xnS4WcyyLQhOB1YEOcQ7PMIlW/mI9
FcInHH0BaLkBUtXXO/BZuNp9iVyLA3rIWdkLK/hH8sy7z5JEfWF3DYlT/zHyvhmNSFFeaCmdcF+8
Npv15yNDxlwYfWG3mBSuT7onNazsKSl+rYs9YMt1NQIB3exPVrdyPGSEiRGAwpb/P1toZUHMlr86
Bt4ZII46BWlnJOENBQOqkDj9BcspemolvCRsrhSUJOAF6fZLJvpEJTlUjWcdmbEHA65vx+VykOVW
FWrCUK18hWV6K+gGzKmfU+WrVZRwwoX3tdkVRWm1AwwyjXTowMzxB3shE4OL5om+3I4PQEL2sXb2
p5U3gWD3I/nza5iri2K2BYhwdx4ZzGParvkZ+7YI9YTc6eHe0QRnhhwgfmO7mHkXBcYTxRKD2Dcq
OyLyOKdkaWVmtjveRjwANrmiwtcsoJtzg8dlySonqtO3uUzZMkuQ/V6ramzJKfu8KDni7S2W5CuC
rqvqVoPHp6z1CiGAa9wVEEu8j9v1YWJRRILFBTlyv4IeKcKgbsd4r8hYGJwNm+w9q/jHVcee+zvz
dhQFav8xsG/P0gU+l2pX1O/0pwppmSnmG4B40oJEVHPjLSU8nc779Nxka9iJhRLcrxVR9UTwYhYV
lT795vlWvuZpUHV1kX557nPGzfnLIkSzjqds6hSujsU2Z8L6jaN3n9UoJWvoYS4GEPZSn8V0R0oQ
NkOrFgoEII2zjAO7U+ocVHP7WIDP5p00jv2xqkg/+tSX1dpVJUwLfhZlP/ep1B7TKewGpuifxh2W
vTj5mjyaled4Sz3q0rBEgUR0tJo8wb/M570WJu4ShZzTepBQTYyqRUGNpR46bNXpXN29Pyxm3Blw
xI7WhJSjC/Fv+j13JxQl7KrKil+uyFYII8o/TwGYKEOBHUdGkDb2sqX62kuA17c6tlsZVlO5+C0c
NZAFgAweaTtQjqjrbPJilAUn7QYyoglgykmS8DIpS5M2wlXXbieEYBOVvWB7GFm5pqtTIo+Qra6G
SBWJjpnbL2AjI7BSleZk9OouydwZE7XXI0++0QPWqjYjauiKJ0x6DzmyXmKi0tZ/njEMkmKA/1LB
1n8stAeY3t0i1aCpv6s6noqF0oUF+0TiRwY6h9m+HZPpQ7HIYtsjf+EtBXmyRLCM8ICG0bPFtjoD
8yb3BuVuQ4zDdlJnn5PGUf/kIt5qXZxicbiy+369kyxcYDV1CYBhSrsh+4v2CDtXDGYY9sQuxIXX
MLqnQinRjKA9yUy/F7FdYB4zsQMcX4AnHUy7Fs7V+bJ5CnUoAinbn6mJOI816NwsQvp9mdykocjA
wieU57B8U05fA+FpnDexV9orWjSOzDSsBynK8cXgwLfYiK3lG0/5mQqZ5cUjuclpq+nXbOM7Yu5S
sLA5kqV+0mowrJxPzEt7fynYFn99xek/SIXDd3/Mra11mGMVN95Hc/GrEGtURRl6zkyJQcpqpem4
0bQJqM3SBnuClAjsMAigeP170Melzg9CKCKOlBkOoB6hJkbkLHQhu68A/aRp5xoNNfp1NdV4kYsc
iOgykFPvpwPvzYFtwNggi7c3xHtXWptLWWExqlENZHWtzLIEekFOrg+oGM2mVNLhiJ4qyNgDb6bp
0KqMnGdVDH/0aXTQwud1NWnPPyJyMZcdOCaSkou04lDv6rv8jawP8xJ5mtnYqys7d0RlkeMAstfU
pSybynrkJS2iS/LAoDkvxAgyaz0KHPcYKKfFxa6EyphfmCJI3KMADB1WgVz9Dn3CceUK+JoYd11x
5u1QWfzHHEYs7EhoZebOrIhWQJN0ftKlMVKokfhAbf6iX3KIKaw3e58lgJGRhDZdj17l6zYOLvZd
wcpimIkly5QYe3w6EVomcTLfYMw/Hx5CZyMNFC+jSQZqVtU6+hMDMBhSAXZRLLYPLE8/qOuJLjlY
i0P03j8iExu1H3g64OJQ9dXQ9cL3HqOx/0dKYOyIetSAatDqychBaelPOpeP/Y1JqWs/gx9uSNeO
/HvF8bH9FkCc6Uu/YFmGIYo0Ls5A9MqvWOZvHh2G7FxELxMeH9NPk58yWwe+eDm7XfKJe7bL4mnn
mPl7EMqRpqyrtLArSUaa8jePiF6Jz9up/wX0KSfNK60t24U1bul/jtZ9PXCABRHGU7L7kxLULEDs
2lC4jrC4ooUWViX1DuilpKP9A8bkVqsQHzKvz3OT18XvHG+Y0n9ONlxuW8SlRcBqlFbepPokbBqQ
P5PFwy8OfWLPjO7oylG+2uJ809T+ctnHhjYhCxvnPpZL3XAknhU+JZgpxDA9+SVrytiCSpzdbvA6
l6iB2j0lZQzClhQQfOQ+0tf+DV0ofVzL65lUKM1wySwf6CB8+lL9izDCoSq2rYIRbEgrlMzhlwpa
U4CYnho3Ujh/a5lUGmKfqwxcvYdBmJEE4pgPMdWgSIycRlVTTH/cE2oxjlGSZrynTyKOgWLOWNn/
hFGHC7IuIuGOA3KcThDEBtiPfKkJp9w2l9Qaz2ICf/m1Mpp6T6DxcBAcacaYR/JNCy8dhqaTI+3m
QJM7MEHcT5Z326DaPzdnl1NrE3Cp89qv4ZmOktKMYHyEi+o9uG0PwyRn26350DeJHn4lfUAql/Zw
hp/ULEDzKgcA58sfzM0NJUSdlUIu22R+k6zBXMOzubQuW4Dq++ixabcLN+e0yEasiJdBZoMglSnX
nY79BVQi0Gs1QeNB23chJj1HT8+Ny0PNZ05gn3kGBpY0brocscB1CKQDEsCcpNVZiqB+aW882Hyi
YMVa7ZbzQvBW/pEHYex38KFD8nShuieLqx3PcWCzYnUtpceplu+56u05TBO+7fBWYTi25xP8VexH
mxawSOYGddggSlB6h0hcPz6NGUnHNRZzuMWnaX6ylOwziW7buPXUjpWYNj52c4OWQCj/P5t3r7hW
ZXu2ySVRCa3/D4s1kpOyol0Q6Y1TGUHwoGzVK3+fH+QjdlZsJsb3sKshWewwS2byhVXAGDXd/NTK
6OPQdEHyJtdUiky90ce7sIW4rFIDNrv9EXcXD2ax+vjLFJWMD5AQhqzzcUVQvRGk9MLhLJqBV1Dg
/eO1p9AULg2XVPgS11ynnh/hL+j0PPBUgXheBAzbymLahQ5eOoc6KB+IZa+evpy9x3HQTUWEg+QA
WilQII9j6hDaIeLoiGRUpLogwkzR+K0qni5fo+xum54T4tFANSsr+nOPYiLTOXEsiVLlRIls4U6n
WFgQYCU7eEOWKoZHHk4bNvukrko7wTawnw2N68gfgLUb1bM6xTKtXc6gH3uOa0XicP/a4VNoFd9w
qpaqHvIjkg/2zekeeW/Jj1dpbOZwMsUNGqOmXDQUeFpHlzz0fKtNJAwFwSzagS/VWy+4+rx2xkJY
l8gwwb+QMCcoaSL0AF94IyyhFN0F2gExvTvS848zJpyBhpUbAwiJvUQE5KoiiaMnMClzHv9+Gr97
1RwUC+8kYJnw7SDhOW0kYe418Jlqit4t7kGE9uHG07p5HouL0Grq5ofJBUnJ9KrTUQEPMai1TAnW
6mX0LPTxxT2qOGMZXsvbzPieYXCUhso7ol8d4u1KT6ExMzJxQuysfu49M6bsp0ZxzQTm3GYh08zT
CriSSchD5kPc0SzDC35xz4yXMfKo3xO14SCHwXUUHa3Bhf0mbWpvEEOtS4nEKgBOlTUKunkCPkaQ
pbrtRUXzZc93D+JcLQ0OVqLSigljOJgvzv+d2ePkuTyKDbvqi6pIGvx+A9rAfoc9DixHqDV0ORNn
zAiE0UZVlrvyVRtzReKK1jU65WIsD1evzvv4TEXwN5EI+yXByDTNv7mg6bx2GW2A150mrNpGNcGK
EMWuAGr4h3Yg6fQ9BY6uQp9RzLYv595EfcxDKYei36gnVXUr2aZpWf2V2siuiNfeywGFRnYWG8TR
M7zuWuApPGxteUkZvkFxfXvAkg8+YrmuQ4gxX/11HWbnOg39eJJ8516QZuGd4ZAx5SInv2TdUtA+
cSp+G0glh83UsSmjNVCrarEQVeWBVEZaFGTZ9shOeppYe82DRd4eCcuc4sfFXTWmEXk/wFA2Tu2B
PCH3EWMIG/aAYIIdc2B8Ov2mgvKUQDK4iC1E7DoTxO6P4lguHj1xXG42+d3NkRJT4ujC608pYQH+
ORzuDuImj93G4IlxYpKtzWpPVkyGnCZ34NJXGY1P8yhYSeRc6C1T/j4LMUPuT89UP0qGmjknHbr5
srMugbdVhJF9qLTk7csCmQ8DKsT0DsBUXuVi8y4Q0NXcOPUUyRHmV69rSXgQyyRrVTQbCLE7Rpod
EcDYv5M2xqWAPUkifQU8bI5NWqFF1VSkBjRyrIgwTN4IMO784baKKbKXWtaDmBI6tXJ09lwUxrD2
m93Qe0M+fWmW4huyEAhWM6VepTPmCVcrk9hYuUT985FDc2agOF4wZh4zlevoiVhVUp9c4QcFXEXI
NInw7z9aJFmMOQgccNNFAAByQMeKc40cxyZwYfWJ+/4922KQ3wa/cmHchgSM0n6REX2RGLKi0hMq
XW6uaIqTMxpDfw9CHfgI2rZldd1XzUZsj26jx1m/0+Gd+4fWHm+1CILI711Fn/uULt18pwq3qdnv
KL+myv1DOWCTa4R8e07WfFDyCrKWCw01fV0gg5GUNsU2hhmHLbmtDzoZ1z9AmKH3jz06TVZjSJes
g6cOV4yHJMHFFqPb5VQGjnmh7Pk6jZz/7BbWYf5TWHAd7AsdLgx1Sd22/MH+91wv+kYy1Egnn1Ih
JZ8B6XspVMIVmeAWzrRaT5AcjWpew+OddZ6C7q/GUw6S0Gelm5N2jLTY8Dp0URarJ3slXXyIBpfy
0zlLxKB9PxXO9QQ+fflC3Kg1/M0n5uCJnEeVEYB7Gya0FvtaM1qFDwdJB8SNYnNCtCnEF6sTko2p
3eJu0rRKNb/lJ6V/3qR5lw1+cCNISRpZsd4WHeD5r9QOGDCwRO43D1auYeyrbJGrseWR5tvoKHHq
PvGX7pVSUnzlhZIs9blY+UUSuT5EpbPZUGjWRDOaiwifsizUbAHrdaMa4Enw5dPph/JgLjN8kNke
eR8UtvmtHQzyuagcO154tBVIPQbIV0uNf9MDO1PoE5oYjGfRtQW4M9lxR6495ZfkWvPPG9hxgWcb
HD4bFtrOtMvxrsV0HmlSXyV2vsiMLCzTgb3HiPRj9C2JVOc54GGOf2i04rhcH2+BWF2c0a7PcUdF
IqvW+DcmSAToJQfSWovY/I2FJOtzZuuywNqOReBgaepJlRH7B0/jd6C1oIdm3yKryhZACVsGAHps
YyJFY7uGlB5eu3HgrkKssqDucTqsqDR6zQRPH/LdDjIbsi/DNyvtMZe+KHeUmixrRSWrU8Qe5V/r
yCEo04gTPBcTkUzzr7TYvIAjEvSOPfZq88KO2C5Ma1+oB75mgnVj7t4k61S48ik/0LWm/CzDzebX
dPk59i9bWy92DvOyljRuPuuG5xFl0/XRNhyAqUV9eZlAQowT+yTwbIKB30PNwqEbTR2V5PYJLP88
qjN2GS9Tn1IwbSO/wpVW48ET4CV3rs8QqQyxAo5GKB7AxTcXVA5EAWjXSRuDhwg2d8H1oBv8vfV8
H+4GrUS/67KH91s9Ahibpu4cEDsdObNN/y8U5IpUrhfxCcS2SRRExxDXnkfMle48+pIS+U+suoll
5qVwHcTbYauXV8t9Sd8zkNNN803r1qQ7AXXLBNQRpDvrX0TXiwleG3cCx3kBXUsTO3rk7uumQjgE
2Ao0YMqbqavguFp0D/1y+EcXgXms3qgOqA1+HJ39dN/dk2CsYTGzjGokE4BPM+TmMCEHTWC+vuTW
/uvqFcEAqqKWRsYDzhenstsLa8Rlu507PCAeQaDZnGEkywg0FNjD2G6uXQ/d1lb3smtMokLFB+BF
JAq+wGhcG1qdjyA6c22f7Se7iFSVj3X3l493PI6J7l3IGxlAEJ58SwIkoRIxJJU56MXGYByYQz9v
JZv6GV8ncbYqWNhN3FOXTXPUGylR1jyemWH8dzZQGi4eofakt/jAG3HNjuym1w9rDr3xb1BhsEfY
cVPXck4hBhWh6QTKril9S5VbUaO3//j8pKuShkN6Vz+jDi8fmvRstFqJws76peU1RIegs8CqrA46
NXUso4f9IcvZk/hYPrnuU2GS+hN2RIcyKPAD28acp3+F+xw1Pc0aezbi3H9aW5ttR0C19J8rgPbq
LY57ySAe4UuQLpWXnjWBjix6IjZwc5PB4iBTvRCO/bOiUNPVgoFphCsQY4nesYQPyTt71gr6WAjo
38nul7LhM9uEYwN2m8AsJqODcHxIQfCmE21MTBHwddQSLFfsNOpSsLksmqQu1aUJNSYqZoMriLGc
+iH7UWkmqSNm1t4XKwC0vELabiXz8+9Stixnqi/IqlFyBHMO2REx0aN+Z9aJUa0juF7Af7eH/xh7
oIT4Z7l4ysZ63qnS4rmP8RXI4hgidU0mhJ27onrMn1VzEkLvyfZyeV0IfJHL11NPcSeGb53oLv6y
rvjt5XXY8hcciP1dtQd08cRJkkX8eUS8gwdGqyTbICsWvPSu8Nr+kWF+rfTlpaAMvFJK16wy5w+t
u7SYqKHty7q587hkXDq+EISMEqWuvROHT+ZKtllGWKMXYCsSRdfRfbD9obstm9OHH2i1bp3hotia
zjyVLFZQ5z41kj1kXnAvlqtd2UsG+YW+EhXr282sKA2s9v+GEB64jluWfkO6hsGCkJwiGNdAU99X
5bIVUqGS4OT2Ifk4HuM6nQ0S2ij8LjP6sIM0lDPp3izMH03Oir4U/fv8vrXuzTRUzf3c8q3ysEPc
FR0zkC6oBc3QRmCvyX2ANRDcpoKqZECPzYAdClX9MR3LSjvEh+FTPSkj9SoPdpx0wlsisr88uGR1
W6D9ijCS5SPYe8hNes5Zy0RD8loBvPBCs7Rh4emBTz1uqcQzieBrB6ICa+vxz2Plw25+Vb859h1l
aEZovdDToolJrLc+4+ECT+OLeCnfsoQCyWc+8PP3R8m/Zmot5MKsZy1zuDEr3rXXbBulHq06fyi4
J9DUZVvPg8POa4C8Yu7cR5vbF/kWbJggf/ECK7779O2iRfvQtYzqpM0tl8HbveD4P3To1yicRINF
OgLTnIWahZhaV2Fs8obHrteUa0fWH8QWntcJLyYSMCpsAyLrWw/3H1NTgEKHJIDWFOJ7nJIXCJBA
78kUkSZSxupZvB1qp/94G1ACLhpkRhkcBH6rknQfaQtYTCq+Poai7jG9w2cBc6/ndXKiObZPKw6f
o/YIc4y4Ho6+O++Z8rRDrdVhqNWHQcedlUhlxQuRME3isyqWcBDfHwTuCuviw5kVkIs32iiOFj8x
2ojaCPzzWXjt9sDEE05JqNB/NNZPBSs3/DlEEsctDFM7rJtGsVeDRyPMKSuKQ+oY2KAoXwZhfjcZ
XNPp1y1pgEDofXQwIstoz/Lla8IQVfJ4iWHDeMcAp7bI2cK8gedge5FczOctp2AuvTlnKvWZQPfw
0VWwd3PMJ3BWSTTq45rdsKqWZw4jF/NQP+1o2DUTIblnx3VjEtT3ecyUhmgMbaxMMR7a/onPwTZ2
redxVPKym3fClXIrC03E4BbJBfAcTF3k9RixvzNNV0ANEYigkI/ODFxmmnO11fFeGDegItRy7npm
r6v9uxpsbZNwW/j/kRjqIFVMFvnSU5vj2WkFceGCHrfIqAVolKB8K0wC9jOydB7aE9tZuwjsXegU
/d3JNcwjRHsyM86AiWLHUIpnhJt2pPDDUINq9jH5xoePr+Sj6SNQCRipCMpP8ASm015wP7oK529U
dTuBauqS2xgQ9lhRYA3SIp/nRjeX1LHkhPzV15wGWjPujDW4U6iZcViW6tkIiGRIT83ksgBVSwUo
VycTTtd2OA1KqlEi5DtNt5wtiuaQgL4Aefuy9OqlxgMtjf0CPF0P8ZjUS+j2D3wxgktyjYzdWdbz
TMwlrHj5PLGP3gSz+1KzOSZECO244TIW+bBv7gxMBGG5+XItnprRV2KWuI5eO++S6ebHww6TNluw
9iPiBAxO3dosy/KiIKHB/rtMVGD++iOAduQsn1z2Yowh8CNwP7ADuxCBX0HZq1raksWVRt0V/DIO
9v8LjpnIyQULZoQ2oXmDtR+caftsddGqkKdU8jQlHmEnQg1NCmc9kuiMclWb5h19mNE4NZe9ND35
FlL9rDrxiW+p/B/S9ndJCyXxCewacPPRYOHYl+iOkySBdZkZpsLyHs0IQzQqtrGwUlKzIJkvKLgG
dg5+C/qdQbFh3Mz/A2OCirhzLNQ0zex/QspF6pYNM9aTSzQ8Ok1yHPw9d71Ql+vxQY2wWeNda2zb
kk6FJPHhcSm+7bWAs3MgA50fd56+uB9aR2c3XBm55wCkgy5Yl2kKVMSeaLgbcrF4DbdL7tJzvP8l
3+5ma9n6+/jn15sH4PDV2QCtTBpG/8q0IDgbmPhG7g4Osma7QhQt0wKxCyCYi79Ex4tbOOPVzK7j
qKbtMDYPv1dhfdvm93e7eZr8zRj+Kugg/+ZlNrlFZFkW1uw5UVwWM4R4zaLdmdR6xwZUxvJFEqRU
H5exzi777KqcqFipb9Mgcir2h0EgFDR7Rfem+XWkxJkVo6LW3fqBwrNhoAI7nuJEZcnazbTVnrdw
HxfYocvIIOMUWQWyfIpmW8GXX/06Eq5bB197SX/VSv2V0EHyIx3Qs9jNvpM9AVer0QNyNhA56dfF
NOioFy8B49Lfy6MD9Pu0z4N4ACexouIhrtzko0R7K4RdIw3PKiuOspAK9MiYqiRCe4jkTzOi072x
IpRxDEfVhjZOojQl7IZz/86E8piSOe4kL3D1nH/Spi6B8tRC89/11Ku/DCaOwKocd0y2Ft+UNOBw
igv/I11VAiJt8bA6CSjDCpkQW8RkICmULUr5WQhEtzqn011AfpSiZbrqQP7E5BzJhDNgzdDahNhV
8vN2ut+k8VuWsDwgJhZXb9jN4v3HsnsvG0LvtLM5FlnAO6XXm/5mxvDQbaRa5hU2vexStopvqHuo
R9QTFY9QX9KJLH1RdPmyQJ1Fhgnjq5C+qIC6IITsTEmqWb+RDvYbUM9BIokPuR4FRzjVq+DYBJy7
qDgLM/+fvyIws6DgLKsJ1iqsQ2zBzcqZ8ilnLJ8wh1CDRF3V9JY5YrkYYdNuDFNnkA7VPzxXV0Sy
K9pfPZLnd1ddndUfJywWO5AJ74I882Hfh86MB+Lirs6mW75lYQ1I9Z1oLgPhE2ylQH3BVEZ45gG6
g/b/uL0/WyHxDwdWMqBM+MLtaqHK8sTYbRgA1FsuvmPA5RNxR4hv9qoYRq7/AbNQ4t9casUidJfG
4J9OYXrKCSgO2xyP2FDfSHbYhJSA3dfJwiyv+lV18Gns3lgF6cvu8U5Pf5ozVlnaerRs37lqa9+2
OsfcMORihXi3BLrWG4hFKpJOtSLS7Kyx1L0FuuyiB3bBY8C9gyTvV05xHMtUa5V/rMM3LmUGVPTZ
+dvHNut5K3Gv9XlMupAJgTPclDKZHYDi4ydYZkyX4q/A8t2ytz8lmr9s79agocA9cAaI4/jZn07u
5WSwoOBwQy6gEWa/mvsmWPB8hKjcElX8cATl11jzdm3/IPIykLGahurcZHpHpN5LbTbfbpbwU/Dr
3l5ajfDWqVY1hsH50FPRtVP3sULXr8wgPJBOvTGrw4Hr1Ux1cGekj1RaRAiPDiA4/A810dTIFAkD
H8KmhpaoyPBCBXkRNX9jyfPD9i4eMsdIMCUMTo15UdhESx/FhwPM/ubRiM0eOqnhLUEVU7qle5GW
4aiHHi7SU96ANHR6AKG0lwrtUsP3enLzOsRQLXwDNfIlRihcBRfdpaZLGwi7V0cd0y6/VhqdwX/g
klCu3aWbmmqfv9eaTlAFIWv1Hp/9y1xo0OTBhI4KJs95roMZVMI+FbQG5LOJYbeBu3+p6RdeNRKc
XS5R3Pk8kOURMWcu7XGgtpv736mKCs3wI7Tc+/9psqKJNIQS5pWzE5rxIgK1rI4fznOYUTjJzu/g
OOioiRn6qP1GNv+P2pJINY3Yxf6zMk+Bq7b74AVNDRIvwUALcGTaDvJcHxcvEc96wbw93F5Mi/xZ
HpLu2Hsx7FmeayfR/xcRuCj6fG07asvcOb1iSSz703o4p2oP+nOd5iZb0Ghvxz1hwksvDiBda0io
ULDUBgKIoUjBPian3TIDlMaAXQTSRySX5OP49K7db3WMEMPUiSoIlgFqyrenWbg6aVQy31DP6mDW
/3xaDk3O5iJuyD/oABmL+MCWEXx/+pSaEDFogb4StRGQCcM6ZoYuhqXBnbBlANVZEN0FiGG84BMu
R97O4QGeNzmk5kTWJeL8VfkDwgBUIo974qbfX6rM2T+0U+cftOSVwrTWdDpRXNdcjxeouTrs4HRA
OdPcksx+FOraDbX7YNK6zsuhCDi3cl9WC114V931u0ZKU+vcR0ROQY/RM5qz6ZpoRyh6KkfW01ir
GH/Z79uNWIRdsUzkhXHoBX9ZU0OvPPsfI0p6y9EW/KoB7h7uFVBVIX64h/EVPPAjOn9FHKTkSDg2
xbzcrSSuHksGiKxwr3SOpcLb31TbQKVGx7Pcg/yb+smRhRHB4ZL+p6vvNYaaCaiJRyOazIOMFCiK
g7KDiEKh+SrBeyiY73VdSqcA4kG7dP007jZ7niUrxp+sTDthjNqPSzY6jruMNdAWTZ+mJ9EsBAVh
H/RWO4iSh2/p+XMet3F0SoEDFkfJ/a/XPzC0fIprTh3tqyYqrzFKZBMc9A/KOox9dUSfmoLww7aQ
Gnd4pJislI+zOQHnFjWcxi3QnrE+nt9lkax0Hxf0aGicaNAaLGlS4W0wuX6lvuNWfpR78qHqq19o
HZsgCp4JLMFjZtXDINFU/pxf8ClVhHlpXDrCJ4FwkmWiwdahuJWJmTKeSQJUcAyPpYb9HpkGiA7J
1xJwWu2Iyfpf4xynEHEuRfRrN6MMgqvhDr5VUaM6OgkfXRi3BHS68o5a4ORwoUYXxVI2QqQWN3V2
20qMbCzH9Mf4bJ3zksaK4yNuXOWGGv0IdWAGWF4f7QysnAQc2zC188gMa8yeeSQuFHWNpgtly3e+
nEitZpSzn7rnhOOuBZ95N1YlmJuDeNa/b2xm8tOm4GSr9wZApCAgJmE9cUo9np/tdaEKQkjxbxvG
44Ef8ZFOtQYaQBFP0hkJqtCVPf9RnJYuBM1CgpiSEgcgP9WQt/GSyc8mbOygJu6uEYw+jk0aPxcW
7eSMgNDAapxH7l0ALGXaP+HTOgAJDC+EIh+F7hTrNsLZQyeZ7g+7KC0neDvCGAv4g106sl9p1dMD
SGqhF3Q3rMPGSd4x6lHFu4CjOBkWtYkRbcQ413Kx2Dbj0klzoT5zpg6/0HDCJzrN5pPOo4cv1UWd
ryGxMbhMCLVZXrLU7Lxc9D383UQ/tKfPJxqyDw2Cv8nhVYEwFMsIMspWV9pbGFiXkwbQP9raI7Q5
fLi+Wpv1Eqc6KRjqwPrMyqaJQYRtHx38P1eC21MZE+ipZx/GTpMadWxn1x3rVbGjU0DRWnpGv8aN
Bek9epg0refXAKmhIlFvTsw5p3TReY3J9iHEuFj1x9MYm8cIoCoVrAr/4AYJBJl/4NYkUW8KnGUd
ic0b2hY6lKayDJnNsE56UldP1ubOz7vwFPmhChzSyENu3FnSiLAJSvZ3blnsSOPrVx8EpYCKGKq/
FNfSZnbw/rt6sFASEBfTr4pyG4ONejNu/+QWVkt3JAfmjTMkkaKc8D8ctKEbSBUmpGvHl/0fB4qQ
kzgURL+K+ilLACXh4/QqdipKQGMLA9+dD8Kvpr6lNMK0tTJjDEDIbu/SGcCOoaEUkkURVSt4KYAo
rxmhtlKtl/nYiY9l42CaivY7B7/1DJWsivl3Le7saqXmjbVtFSRdOzQgqEv2pGPw7VtI9Mi7cx6V
G5Ly5kVEo1qL+lpEWO6FH8GQ3T9OauTrnEzZoWtc+3osHNt/wI4+Od/NEWVObY5KtymWUYIOSvIi
YNJr7VQEhFiXvxvWa+3v/ZgCL2S8/rSyGAi4ggs0Qji2Pjh9fYrr79ajR0Ctgha9aE9g1hGUakI+
DilU9gmZdy4Xrzu54zD8cdm+D+2M6gcMGUe/zBZqZuvzvsvZlKXajNpjjhQ2bfxgumNvqwdspn7E
vw0QKy5R7UR/6M9nC5TBMKqf/jzqtACV0srw4Fu4nBweLKLCbS1P0BQBhEHs0sz95NpBO5FGmPj7
sOPPn8lWbcLopORe6f6kSH9PC2tnmuBrW2spdpBU60YLO6ykr8V1ylM7FCUfWv5caVARIBQCgE8I
v8EFAPjsVMMg6opazLrNtq7QTE5vuCFN+QGyHX9v/l6LTDw/9IkQ/o/NeMvgkCeuZxR4+DgUHOhg
/s6f5VQnV6KZFz6QmdhJzM5ugQd05nM2Zu3jD4a+ciujvjU/VOBvmVJI5kXAS0sj6il21eH3LEEM
7US0pcQt27SEf/eIblWecM0gMIt3ry2sSkiP4L6HjObONsCdL14ceLwGaEaP+x4KBIUz2MAL8peW
TdpwRcJp9gaNSv+HT+8eEzBEx3MxQfsbj1W4xtxsvi0ruzN4iGcPnUg8nG4si+zKXBZEkvBPpLY2
ZpAj3bKh8yCPN1oaC9nKE0tOdpHGKHw5wGqMRaEkg2tsQAocQsrfY5MIa2kQO14cZVJQVpw6ox+d
QW2KoZTY24OdoY3tgsW5EPvViSUkVdN3Sn9tV5fqz8hrEtaZnkVIFb9mjvgw7rDPfbepuP0671Hv
rk8QEfcFtNNdfrOjZaLLYQMq1ta9z1n+eB13WO1IJDkIxnVdUcXzFNCGlP2YKE8q0G1BUbJ4CBOF
3oAg5NDpwASy1XwIrk8GMw6wPHXjspv7a+J7h9vUmR4PJk9MY4aPYMqrydf/JYhUpfIC+mCBjQWW
prawgjB3atYe4bHh+A6tfv2a3DoOSn5jPrkZLVWGC5eLo7vrstGEggRHMgDINRlSloYyKwlPvzgu
h6QVUk41ouPbXpCzpaPSBgqnDHrJTD6WcIJH1ZN+YwHvZEIv4/v9JgDWPJhHslqGGjGAMbJNoY1C
cQJtbTTPOT3UEnGsIPrqhfy2ZRgG0FX8zDG/qyEpJsnk1LyLKtDZwCjex4RTPyGxpLDCLJ1zhYMw
Op0UrmOd0pRY2o2nnwAQPLmP1MQyx+x7WAezIyJTuCZ0CpBfAsn6+mjnA08/wrCYnmGBBnCYbqmP
8KzHxLv8xFWmUJXDqdWqJhhH8vfjF3P0qlTa1wqmPhl703PynMUVBOXrXS9RboniddX+gF4CiMZ8
zwO1jBc4IYAAG0Tn5l0aCErqwz/UbNsO3AQd3Bp3GNozMaycIOYKEBeZqubLmgc1bIKsibGy7zpt
PK5hYsqODCOBw9kXECFyVLLz8jTvG/3dl+gA28syMg6Q5ESLBeWD4S7QEqYOr1UqwofApelh32RA
Wb/cHcEqWYPRJUzyuDbAhr7J4XcXFQiX63weT43aL5yE+laBjjGtzOEc7+fNOIKWdtp5rH8MfWc3
H2McVKmg8j5X4+PlLojBjr6wBepEIxgzNW6A4Dt0ls4CmHLXdD23cwQhPjv5LcMukJw8X9n5Pzdu
UjrHxO9LB3zuBReebahqa9vXHkfaw7SoqLw93psFXgu/D9F9xfmqJDY15rPwT/Nwxc+qn2pvLEI7
oZj9oRSauxBF6EpHTDiciFlcp+IidrsKHYRgvGQ99F4sVD7pbfq+sxKvEJBnh8Qzxrm+Ur3tmoyT
YKZEti/0YZPD3UDM4qtGaD3cquUwzNrvpeWG3/xfweQIyTy+qGp6yrZ0x84GyHJB01hde15YbKS/
OcaIEkWBEx7TkQD0YaitaqGnJPJR6jPKYta/hJOejWM1UOuD+MhS0zClBHeeuqRIhZTVY2U37d4Y
cW5esgbSx/LGmj2gwoBJ8yqd7TUSZsg5W7Q7fWHuTx328nyybrKkeOitvCZMIQhqtIl8H3hmjVQR
ncJrBcbMDUt/gHKUrLrgDPey/kU+n+mj9Q3T2Rcnp6GEpYFM5/xZ0k+Qw+OVGhhNJGNCBp9qmegb
l2/QJCjmjDHXGCzuX/earRqQxKmVR9xDWoQrd6OP4Oi663ngVBSNivWcVEvSPqVt+D4t8Suym/3M
ISQl3fL+Z0moWxG5E1qwMIDFJqoz4C2YVwo8gdfdFUxNcHYyHeh+whbqeraQ6K7oXUsrZWfKW2s4
eIGE09yR3wcm3mfc+SdHYR8IVO7c0NtNLblsutmwRtJZOLilrIWy64T686/9sfWj0gUyQxOvq5HN
rALpGCSMNUQn5it2I1HVswIapK3yjsMbUmQIEiiMyRt8Te/LuS8JY7yCbP8ZIvL4iQ/26pv/mC2R
2q5LJe6KvjELi2S+FxBiAxP80Uu0XL/lJlRrb+sV+Lay25SIA32TKRyEOeqamm1u+jwD//M+G4j9
8D20eH+hOkZt0Uuhw5oQV4V2I5C2rgVwoZiWPMphvrpd7auVnqrj3cyua+lxsyrffxKiZdfhE8dB
1ZNAw1fL2yGgybD/k0fbMNJjG0DzveKWXWK/sJRuOFJBiwIuxcaBRcvJ3G9ko6t/oNr51Ffxwl99
YU5N4N4Qm09s3c/WNn8oW++tm6U16Ct2Q1yrxJ1QgliopuqQdg6CxaI7FsjxZJRjFn/dFnnNr/EE
z491NgAyG+9bNl87hGAhtWUiUe/gofQXtZxRK+NZmvs+FeEdqfSw5gJ1e7UkY1UThfWRA7GFeXTA
VeyOFXEMDbR3jbOwYD/nrbN4Excvi1HH5IPycGpwXqEno/MTXzK18VOOw4GDzSXSsR1cQOBsZpdU
dQfUPwodflfggX8CPsDwR1cps0Q50Y47+iWnxo18F4M8RdQi0wksmSBDIpk1L9doEvAkx+02G+Pp
hrizjLx1cCdWTJJyA7c8P341zlU5hOANtScr2aN6ONUfoCRyyAZLcAPHUbTa1/OdnVD7FJfZ3ApG
Y6W1Ibbx2iDdWr/fiVQe31bdW1J+fCsqaDiYen137EmwtzFk6ajaxAxJefarCDhRhoAKNO8uL2YY
mnTm9+sou/GpQUGAKExAxrUISGRcim8CmV/RtdQBmmFmn12z0xVRxwiJQxcVp7eLmk5XUKMmzGQP
zeX74VKdWY/GqdkyE16bRcZkegC3WOJ2piTGYe7rf2u63drap0MTBEz6tfteoRecx5PWL8bYRwih
BKOzkWJ4MYviTDWcT79Kyu/lYWVPE+ihxIM3sXhbuymTsthtM7RZsmm0bCyfXt5HU3KKfSsbq7wL
KtOyf4QQ0kF72gePGCpJU+knSemB19+BpHPFLEzHaBEWtqwVUWCVRdaDP6RvptpwKURiqC33kq60
Dzwo1/R19/tQQzz9ieHLY2QsrfN6WeqypI44GtF6ciI1FjP+QopwgS3Yley7RVNUWmvgKkywcHgh
TnhcMRTMPgZCcCWoRntiBz8mUIgs5qulJAf/u3/AqchWDn9EKee8yPTNm2BZuBldMyVxLsGn5rF/
JN1rgrqfZWN0sEzKc88QDhPv4moOnNl6R5YhaNA+gz2yy5tBnGLNJMjEaWm9wMN0zgWML6LVToMk
Ps3uc0bK1b1JXdtCQnn/n7aEg4iHlyyM5xa8c5O56MzRJ8rvK69kK0YjEwe0JZDoV60s4cwZ10pH
gGw4C/BcnyfuXBeaxOhLYrs8oEZtLgnSaEyYCfcck6ntc+IA6Dwp3WgArbc1anazTDJAOKxXkt1O
MfKu63pfApJNAczT/0iJXYpWvGSSfj6qiHiGexzPGTUQp5w7hxrjSfzPc6C1T5hG/T3TnwztxAd7
RgaZP+ArcLv8TzOIGSO0f0tbikSpnFVQb/3G5KNezCJppVwPVYp9lvssHBpevU5Bl1ZFFdvoOXX/
vDm9b4KtslXnUphxgqqdIsf+T38vEkORpZ6Vj8PB5ro1lxtJFDtAojmQ8ixbxKL83UwqBEdEJYSE
gVem1itEFBPbWBGqMulvANClvoRQRm/GvHhtBlkzIpQeaN9cK9vR+61V2oQ801/qkESgt33nxEjA
2AIM0MbGuhOLsTNK5iGTmTmcjZmdAPDUwlUEAWMwXsqn5h9DB6MxJm35075ilurJXPj95YxM7V4X
whY8qcXFzlD5CjmLgP3BCBQu0qwetlhAhCKmCC+oO+eEM/NwAtZMicD7iKR8dbL2UoQOrF/UvT2v
IOiD3zngyCDl4cRg6mztNiTP/saOoKjqV0OG5TqBMQuJCUOtTZIq4oszbtjQ06tY5iz1eLu9JCv6
k1QMS5MGqiPsoqbuy4uhoawXNayaqm3DtKVoBc7OQzehsJHGB+MKC1Dp9KykkbGeeS1LQ8ZhR5ch
k/x+7tk4WZGJRyJ6nFzH1RxGWDBxdxv3pDCssqrNKC+uN77Xyg0M6H8ursu1sP1wEMj973KVWhSJ
58qOAqVrweGWrNwBZ+cEVApa/lrzaKrawxxpEDTW2cnZ55ol+D2rmG/7d2tA27pOrxk9YL3VOQih
loTY41XdRjbg1hqITg/Y0rLeWGANAhEUOZIZW6wzOrUsEXHcRbsr8DPQw8QXjwzTj82BYUa+x1yd
fk9FMgTZHWedumaSMUagOv7+tGI3GqwYsURtKt7f7AkdA3sEAIVmnshTKWoQgDQQAN0BUO3sPGrL
+zdV43BGJh4BAwgjDwByzUxeY5tLManutsKq1IecbAerMdI6Y/iYIpRtfQrb7SRkjVU7tih36hU6
1lQSUyqvlFh0fSbKw1fZwZja7h1AHfwMq9/GJPmyQXxpBieBaTrZY4EAT4rFxbLyQKbBUobzRPP5
B94QGfPS/s6wiwC9qkcEPBXBe4T8/fHFUINZmcQD+nmrIDC1ff0uMiVeY6RMrA4evwoLePAmu7Cc
n27/6k7V3M4ixJj7yHNiXAdxy/XWwwMQbNJlByGY3GfTp79S/PSjXyrfz96Go5XVb7Do9AMasoPY
F5SLInrG+3oXOxhUth/Nn8ChGEWH1U1Lb+zdjSfRhxyw8RHbjToC56sUJihvkLm/kFPQt+2fMyMJ
W3z+DeNnDzWm80qJ8I8YfNOnbXT0maFhioV8RWM8DNfcGkyAgwQ3qvK0Ag/6TsL7/zuVwXz1oNuK
sZ0J2Pyr36D0OEEvsTdw6bPR4dePKveM7ylkSqlQjpUabJM+i+bXhrZTm2s9x0T/a7gjJecAyS9L
ecqYE5BP3YIFuKKmZE0jmagkZV+zxhoOaRoQ2g9L6D5OKtagiSj63YKtkYHf3cKgIyNMnJWdvcnI
c9pMCBNArDGi+Qpm/QefzVjue4aYt3+oT1O/Bl5isCgetE0Xn+nbDrBpXHlaE153o6xklKVHUoQI
ruWMWswcDmBBaW/kUOP6lFXsOUuJDI9rPVRLhUSkTfoO3CthqLxhd0840pClJ4HW1gseEMKEBCyK
BTE0lK2EKMInde211966FeiVx+I9v4YRWLi26nuUB+Rm6FFfnlIpZ1gxNDJzzMaq6UGEgm5r1Rnn
QpK3RBGBB9xu8Y3gyQBQ4VL7E5B3MMVJ2YQUBSf5qD3kh9Db7hDeyP4E3SaoLXDQ3K+im/iQyPRX
XO4KbMOD94X2ec2LFWl8SPct0i878bEXLlh26PMYxmwmCcbewJqdnTlryrnrGCvUI+CnQ1u/blj3
BPC4lN+qID7OhzLNIahK7Nb4aIAxIoee1m014RLWsPRkkQx/R8BQzLPKlVCI75nBzzYprQlLB+6d
Isnr9Y5rnAebAKCKWeJOMKzRpoi3EGVEEdLhTaIarCDOJGv57kQTSXROtQxNULjjAjq0g1e+vtzx
qLiK05meOn0EJhNNJVsuuFpwgd6gv9CFgWQITf004YllL8yu0oRVeHSgevhyZyHX67/yb+8Mq+B6
1sQfXD3hBPLzzvRbx67T6ybGbi2622AKdf9SwIKwuf8bkIgkrC25MqHFHkPr8W/HgCjxZjzCyRf+
O1ZogKNNYRg37htqB296mwfAX6YYtz3HYSRm3D03fR79junb4Net/lARAMB/6IHHh+ev9TThXG7i
KdtC7qYffb415YnKwylIO506LRarTJgc0xA4K/MEph/V5FuE8gH7bLEiNIWt/yAaAdEQME4LaAlm
OfmxP3HDJCcC0mCuC+3gYcGNOje1tlgZI/ggoVYxpy6E1uOhEMTDd//GCplKNYv969eFa8wGfKO1
dXALitgwlRgOFFKK68IQ3XWBOE6cMoco7hKTWDjxzcXaTBF4bcWWVO36hGRISCBkhgi8k+u96AVB
4qS/50LWaQIH2Y9foig+Lpz5Be5m3tMkBKdGhTH9I3P6KGB5cxa/eu4WyS5SP7apvMhXqhDBu/S9
i8M1FcqIPMLYH9QflifyL8k/9zY/eD2wi7A2txKlk9pvgsE2Fv5hFDnJx1G6+b6gdZcJM05Gwvwe
pm5ZIhUltxRrzxcxc4B67rBu1xkZCWZ722eYFxvqKwh5wJkEUgIx7Gxt/LBaZ5iVhYphb8thjYaj
wgD332BNbx4xn2nvyhBWI8YEuD6VgCj5gAlzMFQJqPM1yAj8J/bwwvtxck7EDZ0lMom+AiPUxPgP
k2fMNV+rHTxMT49e8vstKAOzTjekX8GrcSDZ3ZoVdy0VKi/xndxxYd65CoCNqhW9gjKJ4WoFZIl7
eHMUcsmAJqoHnZVOob7SukKcHHgwuGDpo8tQZHWc2mJ2Xf8zek230/B+353fJ1JR7JQILqFC5W5K
P5BBgf+KrJ+3nFPDnk/SN3Fex5Q4foRKtxmJvxKTaiPFg4qa0Q5XuCPSv/aU10nHTIRUS8XUzRkH
iGLbmgxtd9ZQcFq7k4aOZ/4TTJbJVkV6VJ3Vfpdbpx7o81HNNSVsxkgQDNYPi33y9gGS82ZRjNf+
aIcJ8uZ4ZO6fTiRXPLiZOgq75U32J5H0UmZSU1hADLUSBWUqcdUrBYvM7Oj4CU1tmfNFjue56yKs
x+u9cELzfoR6jE0vpkRGThfO6b01cTW2DQQMinJLHIcSJu9kKslT+hbXdafFyK9gZjBpXmSBItzb
KHse6vIxazDgCmbdYjMNRjnXl882HvRLUnvZC3bxpxqSY7SBWOUQ8dBVnQe042K0NO1QU387EyC8
GTrVCe7uuYbWHixZ83BaLxaqNvqKilNG/9/c8VYfgXYB5wkh5uQLj6UN4bchd0iSVlwvxD/b+22e
mZAQuId7vBSJDVhVC73qfuz8OnjQSIubZr73piT9ENYojSC2Wvb+tT/0CNPjaHoBnRrvRCq131cD
JbsRSp/rxsQD53Cy6PoFXUE+fX7TaXYwhm6kpQSKo3sKa7o5TopVonfkHKGhFv+fpb2FdUQrhWj/
Nkjy5hgNl24EmDbqfXocvCySHy0M6PirDi1nutVRWGQ5E6hbL2PhGFMRwB6NTf9pkTMBoQ2m+HGH
auEPzme+EC924X8OTXp6gDc312jHSO/IMHFdNKyriD/JrGozkKh8VLaPp52886gJ8EwcTa6sts+S
q0HWIlubyBLMwnS4+hcxhYN8EFp4LUBfbYUL4jKOtt/Fnwk3TzHO5BXwgPpSG8f83cGE5QyroAes
lHU7HaYEED9MGY1UyqgRUG4nzkOhBN5zhDxHqvGwmwnNwGuFksXHE6Yh6fH1Co6YWEAVpc+5s32V
aOe+/N44n0mdX8D9KCl2EEH6WTsuXmzxskaHF9j/uykl54yGv1dK/g6N05DQDdJNAfR6XVZArxAo
8HZeZMpfpUDTj5ddRSxwltQ95NSSy5S64w4Zm9JxZYlfVA1waUWitS2dCXBAZMJIJBFPuGb52x39
yubOupKYBs+aYCFhBAiln2S+0QkHmMQ7jlYuhA71AiCreu38oPMawrxLd41Her/fQULVn2yhRS2L
+9L8puPxapBMLbxCIIm0KS50VusE5jNG4wyx/4/kVhReI9BF+yJhZIOIXlAJ/YjxraOaAAn894Hy
oCln0KxY6nan5b738ISe0H/hz0vErhXWl8UuGSQS2jgs/N/r7cu1gEIjIT0hsW62ZUt065y+X/jQ
nAdvBPUk878B/fCgwRH1JR5T9YScRlwiidxISr0/IKBGEO7LHp9tQnvF8Os0ANR3hpjhZscIG3J0
7Y2Z5xZoDiNH0dAzZKU4x9mKfhHMCQRZ0R9D6pKSN/asZccmRIiGeeeN31wUdXeCpxNvF2BFChbC
lduG9ZmS1f0oPyztXDERe3WzIOXYX8Re8Oml6kWEVNfrwCZa7HK/k5f/nDe8+i2MJoURo7RvVh1Z
0bJ6vlwMlJ875TAemIdHne48X41cHJZTQf5fVBbMRhWk80dHlbuB1yKtttWvt4zjI+2niznrrqur
y1VnLx6h1WQtZtoYBSx2+ERfHEQ0VvmlH6DsCoiia1RkN+5XxMYc61BN8qHsKosfUL9+0LNh7ud6
+UvZy2xXQfMOPjMk1D8CPSlRH/0jixvfpvheIulH9VK/IgQMQ9PsZ59cpz4qKU1GGcq49KQM0+MP
5ctS9j6AX30onlOxw7pGlg77Ule/RyCeJyYySxSSK3Ca523BLefdJmaR2XqFkdE9gPFMjn3OvqLT
w7RukBPbWoe7GJyyfnav/4krILnyVhADbFnpD5E0xxBr7s8k7uL3sOt80ndf/1/aWA2WUM80SkLk
yS9hvyOnq9RgIt+hz7t9ehb3Y9S8nFub7WqsFDuiyKUjON0TLJ8zM8Ta/XNDdLP3QXsS28UWEOG3
Y23su197AgYsV2YbV3EG3pi011WxXkQwE9qAGdr9ugQ5P1srIYu0QsCW7dA1KULLqdnsUagg0V6y
NGHKuJFGVIbyOwSgqOICpeEI54ijq20a7oKApCeWq0Pws2mixA+2HVWUvJkRCfkJ2aRCfm2NrSZk
tzFP7foxC55ZI8uxgU08kE0y1nf+rA/drSs75y1aKnM+Wb7wwo7vsAPYwvP4IW2IbTn9uU+xc8Zg
GfZlUtiDzmAlKnykKLsnp8mSddlLBbP72WG5DuFkaO5vesz4Dt0f3POAfEzWVeEyCkDzq1bdSIqL
uLUSadVzKcroTmRP9Gvm2BkvxKayJmKyNDAW/rFSun2m1v8uL/Pfq5x+LbUXSX6fwF/ZdzryZWas
98CTkSn/PoctT8gdHyN2Fa5vSttL31qbQ8OaCG7+q9H8ewhAZ5V/FhhBz7jwWzW4hJqxp52HG81V
8a4h93CGirNein7bXbyuEcx35XRmPdHDDzqUTmQiqk6v3IQ6tlU7ZNQbpb74oHYAAU6mAplzEkGN
Jflv7UjsrS7fMUEhOU4UYYXQ643oF0H2KFBtDixqd3lB2oW5ledtehlGfrbNITbeIZ82P7Ppa5gf
IJiVyHsN608p1ziKoX+nyedWokJfDvqoYJmn92DwlrvkUUOLkwJsI2FBr31El0IHIQVE5dPXWOTD
/mMvw6fgPyr9UZY5jt+vtNKt9S4uWQ6Zsd5mNZaoMr9eoD5sJbsYYhCR/u1GcvdBaX+ZH2zTQ5dL
RJ3PQKNQLotU04wh1e7BSs2WOFZMA8tntfdGWt5iqQrB1fVyo+3grs8VScpTNmNXCUWZaRVNBZOU
+/oKpZPuKCz+FI+r7BMejW7U+7lfruz8ZMTESfy2YV2+OWIka6vIzV6sVGY1cs7hbqoKil+f/mKM
Ki32mioijde8wZZ4QCdurbyTrLVUyd2bmav9wSyO6dPscLJUzK6cmxKjuVE9FreuaQNiY+zP0Ck1
WaYcMHLmr5Nsul0tW/N+TFdHhP+mSA2hMCA46A5OQtlYNz2a16Sao8FAH8pp/CkpLb4tmJCq9gRp
IlWh4iWt66p7OpPU/zxl+ZaSWasRoP4hazcDLYaoXU3ojynRc7RuLEfY+OMr0xwTQfUdE+TSq34R
JPs2z1y+vE1bv3giLyvJ3uUFGWGOu7XYaNkKkoga2Bw4cbmucFRQmnYvqN1Eaomb2ZdLLNHgOSqg
bRi6D4RAJYgOPDexct+IwA4BluHZAG30/YIiBi0S+1o1Meho2gLXFlkian9gaH549t9OchtSWVqm
vBQl1HFGiRaNtXwiGEeWbqt5UzPGIuMBV67maYCBLxVUzCop7Nkat/+R3pasmag7zq1C1m1kuszv
qnR4S9awvraHEgunheikMAnRrg4nLGe2O0W+n1oAGQGZJ0q8+esCwvGPfq00KSjBsUcaPgniTAr1
GBNp7InoyPKQxNli/1aAbrog/GKYJM6VStwVbp7qdDcWgxJ3d1s7vy5tXK1Jy3BH2x/mUv5z2Icn
0NxaDie9SZVIvJMbOfkElAsK2fFYNbJu11mnEzy8khF17SzUnLJPIXg1FYxxvC44NTa2GM1utGHV
aFr3AmDd3jrLal9zcKfRCr6D5xadssVpEJ7DO8PJ5HtFlzicUq8a+o1WrdJcUcrmpQFAN0/lIuos
RPEPyvYWvUHH4ip3xJwqvV6R51/HkzrH0x5J0UlOYGQit3jL9UF0IoYqSFpOEvy/HA68MqsADCpe
NweQ3R9V0Jc4VjdPhKjLVd6gOnxyuXkTGjbNNQwI55NV+Ua88HUZJenjyp7K/39UjygCOEyd3jAG
rwi+5ddGmR8SykRf4/xdDVGRwnmv/w880+/JALM1n5XWzdqf1W46nY2HiX5kFp+lR8OpHJehdH4Q
2LQhefRlPIrMbwZt9yqlb/H7vBp37emXuawIGfR7cf+23l6ITW8nSCOzAVl8nu+knLsBY9QelOUK
8C0wl3u9w1qs32yd9u+O7tiy+CSAJqFbJDOn5iAh286KuhkwenbdDya/bAAC+lfxXlYmDDc6dQCx
2nF0SNw4uj4zrvCUJcpNkGCJ9whKZOKcXgfwC+0khLBkEkFG6brVfGnR1PkYrtzpuoI6NMU21LoK
KBUY+6AVcPb5Z3OemdFZyvtMQ9DMB8IK3V+NOkQUuRaehMmvHRx6h96fVsaY8A3cCiS1/HqGRYWY
/hoZxmSfiyXh6sFAgs4fXohs+i92APaP97uDHp4ohML8KJeuhWUUesHH/h7y9h2dECVVuStVL+mM
b0oSWNyVyMmzkbK3I/I6kU+/meTR3ukFzACR+MEXkCKaRJ7ZqeiUPMOOPX26GXZB+57rE4wtjYt3
8D8SWW1aXVT62mNey8BfP75W7cZQ05gkxibwDmJloqkorDv9DNyVOhb8G+/Z46Mpy6xk3dqBqg8a
+KOtHLptQEiOpAMAQ3yaLGySz2FyGqMnNSphLL5csKzfQlBveG7YhEBpBdcEcSZ0L84olYM/tkwQ
cScKGmcmgzN3hyybeyy/PY6gdQZI/9YeATdeOfsm7+LM2hskOg9S+8iqdKIXsamSOskFLT4r1JQl
r/0Wngiesg6JlULV4Xa0zZdZxHPVwNDde/ciADvqYZlSTly9PZT5yViob1OJJC4GVC/E8qCp8tSg
65yXrsEy0i6oufUYqxGUubIvfURtrd8CfvFQYGs7ntM96df/1t36RTQH0L+0rpY/plcNErVu/RnH
md4oWKaM56iHKKLoHV52ebRoZI7pPLse0E7v1/zJqgZUJPMfvW+/RtLvrAlkgD7QY10GMmsY5h45
dsc3YcHaVGvHZeUY+OUIXv6nmT0HZBJRuRVRo5VuDI0e+RPeUiN8cpgL/6cnMQCREMz1McVEnqD7
r9F95bvQpVZ+LPvTH590r9riXlvei0dcGgJ26FGf60/DR9hN/c6a7OJ2Jdl7oKSwkqwNVf6ITQts
Knl87PSSQ8m/fqsR0aN6mRcNbcCH3aqrPzudVGwR8f/X3Bhhxi3nlpKJskpRxehICt1RtyJJSQaU
q9IqNxNwR+nOtgfY6l5214efsW2ZExgK8eZaf/d11FHRUKiqhwzDTs/v78P2VmBPNOagVHyS8B5O
vRxU77imnyPD9K88AyimWTr0ciuCceDcE1N1nu+7TLNwGRk0xt4oSr0lW6nSmybaKw3NRzdsw5/y
j0mCmtx/Fj+lg6k1nRpBqM+Iu7BG+rOaJsnqdlz6lJ0AIU0d17FbVY1DFit1Mlja/tfaQQ3kDR5h
ocTCyKboTa8YReMCclDTIWr+PBhFImbZsk0mYgEG3KJDQrZgXO/HCNKiciSnJNlUdiv+4GGz6D4+
lQtztvG/mL18oWroFnWbxNsbJ3l0gVtFv+AsnRpWoSwEJE2L/rrCDG7LwsWvhFArVlJjmt50ke4h
w9RT6ThHMJOmSzCwDvEV2Xgh7kdFHR6pXDzIzzM1YcelgHuZVoh6HsiU3VdHMHx5SyhjPHJT+G8M
pywn482btIl4c8pF965Eqxxsr1w4oiTThy7KeNuBLc2rP4X21Su5KLwxhZ1DwEcsG4R60/mkApcu
QKNx5hb+ixNX1lKYYlK5/L0LVwlmpIXYkuDMgqfpLUDI3Kg0JbjEvYEFcIgmk/M6OJmIL25ieWeK
x5KFSdMvpMrOrRsXLZnmaJuKbmX5tAyklJNGqQsoLDyfIE7aVaxKUmZS2hcPIbifhnPhYv0P0Fvp
3uHZSex2rQ2/P1kWRKg1SdguAt6d1yFx8GXc7smoiokLXqgMmy7SCHnvF/Zp6smP4U0Uy5XA3FiT
niiPK/tVfWdpVL3PouDgM36Tuyv2rPnSiQAR/i8Dw3Q4IAI6/6nrJrxlMiTWAzFTy1G9WSrgqRdk
Q5NFE1UJRExUzK06/UoqqXfu0htAXoGKjNFuUmnbZ42ySHlbXjrvP9VZQ21rjxkO9/bevoiJFqL9
bhvEk5jttsWyhbvBPxdNePUJ0y45NNaVl48f9/YMR6iQRJrLCKtQjNjDQ39WAtu3yVwhx6xo4uBH
ynBC/e72L6oza/II3fdTRT4c1XvpigPhIsIn9GvlHugvpsJ0C+O+I2PwE4yyIDuEFuKJrvMQmwOf
SAU1yYu1i5bF+4kXLMTnYrynsP1V0mcCBg/uNs2d2+OXEzVzMMbvzAhjqDKHxlGVdgE1uMZ2GORl
rHLqFhK9MOHW8cXKRJzejBEP7m0DY1MNvU5QCxlTwDioVJqIQtxA5JEuhVuZYFntpSmEqoyeJU07
/Pt8sNQnE7LAuaoVoEJUI+UXQW2lRrKk1HFTZDdNDUeJOV6/axg5pAm3mGPd380EPMDjIZhbnvsz
dis7ms/bWOLuW9Zr7e2KDVAGSJGjAzaHo6cmYSL349azcjIORsvz5UEL0KoUrsaciM3WfrKhA+Lh
XYLFwDn8gU/wns3A3feK8HlH8TU5mYPPFiWodjOCO3Uj0HFngnjsLLXrAFVbju93sCDay8wnjqV6
j4aumR/rmL8Tz7hRXc4/rFwvcX8/LOZ70i7vEyknWEaesBgST+oLRzBurPUjJBoTixYEa1hTuAoq
FGdawJT2Y4AqsIt+HWo8YE0a752bMw1/XkSa4h2rFflzzfXAFH+MErhks1et6SrT+lReCEfsfYji
B81LmFqIh2lFFXXRkfviKMKP58Zoy/BOitNbpjuSL/v7dSiClT/1krCYBHCWVzTkvcKunEQQeZk5
hK5bCbMtRbZBh1u6Mt7ayxvoKWBAogD5WgQosRN0I0MWcNlRI6TNqIG6BsIwHUSI6CeCgYPNdFHW
bY2wlI7+ToEXDgowK5pehZa0ysUTspW/AP7MAC8fvcq+tweEimE6NedVB38kR/+PLxATBqgwAqaw
cOJ33+DfpOw5Tt0IRP3uJca9BbqA3jb1KLYfuPjK9MgaEIgD6sOComqgGPjMnyqVYI/1PpfjKDRf
o+RXQo7aFlCzNStIoMkrALGgbAYUiCwttM6JTBF3WF59GT3Myo+NfOQbOLHe29cpgHvdxnxrT/kJ
IPGVxvfF1B+KoTIGMK6Q4K8zb/BjfnJY7EhXdQGYx3OT8CqdxtuD2EO1DtniWhp1coO8i6Z9rdHE
g9c1+mO09r1CxH8s3tM07ln2C6KcDXvIb1rCoB03nH8aErb91qnvH2dYFuIytuucEMElT+mhVFiU
pHBVxndA6LOwx8AmaC/iI0g2+Mb9oVeHc93nQqRAaRixKqb5k+ZZ2td3ay1jmEVIYdZZVImj83L/
cuw5ZNk5sLJqFpK5faMsW+DVthwFWcrpKrrpus0re6gcbUAoYFjmQ4r1RxOFqZYPQ6Bqa8cD1FMs
j+N+EH/I81n179t6A321Osb4x5xxPo3RwM049aHSbTr64g/RFJMkySb/VXi6c6D89Q+AhJeR8fe2
z+lVQBxyzlrLHJEeELfosOCunuq5KoxdWxKDxLuVBNm2hSA1jHjtGIvbtuPzgz3G4BIpApbRvI+6
AK2ST9RqUNZodij/XOO//vuXeL9jvPWpE4usP6lB1rkVSOlI1JKVm1zMIUOwx48lHROXQxSb8t8h
HPIOb7SxeTZtgt52KPAcvSYIfQD8qHMG2Kszr7iFZjDwz/NUeawTGgrx40mPcJSNKN9q/HPUXm6X
qoAJrAnpXx0bGb8wU2QkeG7hYPFWFpBodD1IZsBfzY4c11jFensNkV2zupXFMgLnDIhFf21Jz+ig
WOpKteycJmehs876mJy2PTiDPZ79YeAD8C96jMnCG2A5kCns/HVoRPbJRrIlbKGCB6kiiBT5fouZ
vcwv1pY7i85QaLbJz30QSCyCEY4nbUQvfMgMjUsAm4GXn8+ghTluVkeogzO0egkw/M5HsW3Gw/nD
2yvXAsi4fbCPFPAGyZgXyHwCUaYaFDZySAcazPvdgrloITQWXLfAw97m3sJLzDp+DWwkjYjA2XgH
xcHntrhlFCI6tDvAdyR9pboAjzrEl1Xd97zxfkPcoiI9Wz5mqMK3lvOa1GwNMQ9j/evRq8aTL8v0
QXD5ciJW3sIDT4al8ifp0KVIR1ZkriC/+UMbD9O6Emgs7u/5o3i+76HCygpZWQyB1XnyW93SxMpR
EZPqvO8uN30O+8lIL7J2JrPB77eZffd+/E5qVsdp8sHzlIy+iaiKDmICGJeYhV4dlClY3Zasfd7f
YZB9SBBhw802iRiqcUHlJtBeUysEKj93co7kg1Rd0ljrPBMXtZTA2Vycse9D5I88W16zkkiI0a+1
Uqk+CHUlNUT+zB+Iaf2DIULQdU31Gs88lgUsUVPZ0d5Uai7Vpb1nZitP5nA205hzZ+kIjt83j2q6
Uq+Foq5kfJ9k9SVgxs77iJmDjB4tpBbKj13RWv0djffmK2nPE86oiiRfbI5SNM86uEeUIfZTEm2k
dwHfRMasRnTwNDAZ3BRx/c7onQc0G63QkOP95ddgoIje22KvA6uKNo9MiBo2qUyLuQNk1zid7fYC
noqljHwv/aJpn9/886QM0eXsIJylzRcxaMEakRAyM/ZBv4Y5uxAS0g6ozPUt8J8w5mV2MS6qKAvI
qpxPCfBcJd8YvjIrNQ4YKJmoJlAAVLIkkUUvFRDVqqdO+pkk0364jnLQqXfFwbajdag9h7HekswC
H8xZmYR/u2olRsEtXVaEgJYetqD8bdun+557fuj4xvgq2BWsuc67kL1W9DFJ9jJxPuyAm6LmGeyZ
fykAukIF5ZjxM9A+pqFhRcCQ2EddDwrxigTRWQR+hF9HKb2HdLHKEfvg2arqGAOG5scTm+JE+OPo
kZDvfJk08wh0Slla0LE/b9xMiajuaRnXWvKt58xRoaBgN/1rn7jvXYVh1bogc64Bh4dhiUz+1uRy
8eFwMIZj/+Dkw2OA08fazrsLX2+FfHeG7Q2KWb1dRxlMtB/KI0y25zslqx2wcokFUytkd14zCUQi
SNHqh0MwJqamqDVp0pDiJOR/V6edrKLOFsP/ba3QRUMcP+1qMaqXRiPWh/q4odYHqdS2ag7fdC6t
ng5e/v1l/C7ebcs9f2a9U2Qeb/rv1+sZ/27W1M9RAv9dyMvoptS4b7+geRmSua4XmjfBzLdywz3b
oEBtIeP+x5iSwsr4PS6Y3stRkS8LuQyK5PKW64H6QXzwpoIoeEmsSS48QlyqN7hVFCOE42xhVWtv
/aWm+zQ1CYFQk6O1xH50j9t8QzcgLLJZCFekvK2ZFgL4zjx9+tspOyjyWzLjoHMgYDnDT/jYJZZa
h5I1GbEsWp9HPlUBwvLPdfnWmWFN4oJfwDk4W7VYJNZvDP/+fNeo/zznKPRdOAJl0WOcHt1LxBEB
jaIOpIIoDhcASMMwKkTm0+k9QiUihPq8NX/bnkGriqdeQZnaSct3j274CI8eVIun7uLN84U8gsvU
lYyKllY675vuFJ/i6jWptAsYZqrWbJ6sU3Sea3SqqEF4byOODLHzpHEsSmC2OlPDTBLQ0n9X3hAR
m2uWkZNSEVGrjpRz9Wxl6UK7oNI+xODnLJZMwgVrutZmH+xsF3yZZ/MXhefLEPnqgiYoEqH1xOUl
3SnLpkNgUgvhCdmhQ5HH3Ahaz+HA8kWWTk/dVLtwKvirZHoljNjePABxKPn2fo63SB3K7jf/LWIm
9Z7kNFA0RqTca+8wOX4CuxnSR0/kri/bFphcd3RYIu1Dbmj526krNtfMUdIwJfBgMSIOWfDDeXkS
ylAxyinPmk0Bpro1+jSreYPq9SXIpiplbAZ1+5zzeO6DGlM9Uvjv6WPAvONerRcQoDBK9ST5VM5k
lfCU3qABarp2QaDR1ZhZ4pDLqI84wmKlrCf8r71Z9Q51otxKtolTWBmk3SFjpaPS23v/yGp5NHbc
kY4iFXbyUQ29skvhkki3sCgZCnt8UuLbCam05EGZP+r4gMScprA+zXKdujV59gmv/1CZtMv+O57f
dfU0Uj0bszg6NtxAE/fYgIO10O7oAM/FLcMxDQYE9j0RzJQBRZXVYvZ4za7GqYJJaxfqBML/pDRd
yTd8I7Tz9MX9l70R9BP/EEhxRKEUe0BBFiV+DmYpV77COqORdl00+DToG9YDZtSNMw6Eo/zKmGqF
2S4acYqxPZxh1T4EGBTKeHwm8j8IGOTohVK8QeGf/yOfkkvX1IByGaf9kFQlyWalIuRXVG8UORPp
ofXYNTMVl/LifQd21sq8rB7PFn25XMEzzlwN0bMTkGwpDLkTT29+9cH50DZUmbwYYzs1P6mA62Y/
44WG/KYcAwrSOjG9cz2zCAevWgyQJEUhh+qZHpU1i/EnegIhFwrF6SGs1H+vre1RI1677jVRf5BL
AypNwYT+BnPZG8Ak4IbQztUQmRCkvcC1eUG7lHW7Url/TaJyaDRSb6DafPF+ZcrS9BWvAxtm8dJd
5M0Wg0zAtXtzy3QhceXHpogKXg25cS2IUzVtz61vVghahYMIBt32I2QjvUARdyLFrCHuci9YyQ+/
ZVE0YG5TzibM/XkFlp2tTB9H6MJCZEURF/YgcRHXbtBse8UhNDznDwImzXssIDbwgWbbY3jmwl+7
04nWtejpAIFgOdGZKu5QJE0ksPcKMKEiQIHBWmRGCVmjyH2RwY3/jcmO/goAdv7OEprj2WuxYWB2
1tfZAXJgrhDIcUxFuX6n8hvdScJ7bJAw+NwiP/ztMsN5Xm0q3HwJ3rmfxr8h2oE93Y5i4hoEUtyp
hO6fWiLBhhU4vSMsdNeUb3MKxcAOItrvuDJqasZAK5JKR5A0/Ff81yvWOO1Wu8mxu2ST+CAAbu4y
Hhcxqjhpgx8GmBv4hJXw6odKeZMdcCQIgy9sdqws1zngAv9y2mSqtY30PF6NzBJfVrzktMqMfJuv
xyAzzhh9VdUVyzwi26dLHrepJDaBUtzo7qUOm6GqsCR5POHQc3nrOecZuCGbre5DH7tYfjgrrW+l
avocXz0kA2GrgDWhPAHa+/2AJdkufn9owWE2gVY1GF4Gp+qgcdL9sFUM7/4vI3wvXSOsk0+cs8kS
IrpdbcUL452oASNSll6O+Z31Z7zliQTuF89fNE6Q8uwz3p79fAMSAtyIOeNdvLJevrd48hISp2do
ea4P1N3g385IgT9xNyimi+chEbSokvFmdCiwj2vDgBKp6XZo1k4wbdDcxloCJE1LDbK3hA4tdHB+
kxEtsgTD0jlmAMAIeMoVxQURqsCrUcmlD37DmE6Lg4OkGqGGvR2KFyHMLDgAOQFLnK21t9r6kwez
2dBQSTu/rRZ4XD3TPY9bVoXVLgLnlIasDiB8dRFNT5IbYsyTn0ayPCcmGTaA/4TRDwTRx6CBGz1A
Ff8nSrpSvC6ftcwoVZ8PrhjJJNJKFGi3siEFnWsEjE6qrkjcFF5j/vQsCGUPsW3/r7mNZb+CQTuw
Nv+jr+l4SfObx4bhax7sKy2y68GfgaRk5Y717AwXaOYTllIt9hY72gphL8D7pcH5mXVs+kbj+3nQ
Qees3S5lVqYVEot3sysmpOhiuebBsuQwwLemm3RqawVyeaF1W+Mdu7cWsbZOOJXW6YcVyVn5g0fE
c6tGJMXkPolaIlkuoNj9kApD6G2APgRO5VF4HX3hIm6gkr4opbT90/1dPxvM04g+2b2fpEPrL/NY
cLFzupbRMb/Yk8mmXEQTwzNpYnvULAHthwKHQpn9kiAM5OGBGCE4K7nhASjOnGC1LvKj72xqnLt5
Kb6gvDoRohJ2xYTOjIa8C9y1fCfP9vwEx2U2XPTDcwTU3qKr7USap/Mrxp5rfK745xH+ndsmnC1U
A0QcuxH/1NzMfqTcU8P1B9FH43o6pUQakNmcPQT58QDr6V446y1NjUVo24T+oUclrnyZUjgAmDLf
ArIUEz1Xh6Z0pPXU8GTsFWDxXUxIY6UvpqFxN9T5/9iRwcZWG4vAaDeNm5/ODUEBp7BJIAPPS3TE
lrvfxlDSrXWvMQ2iaKyrXO+VQeOvc0LFX0uEgifFLhTbUX9FGHQQ1vK0+iiY5dpG30GXLrNuYbaZ
1I+B/as1XU00TSDMZefDsg+koEASMhCk+pIPTpDOe+KVn/z1tPiobu/ixluQM+KiRFwjtwno9pq+
KVAPM+ZDb1hawm95G95Sa4EPP7zkxee22r/9ki5Rn/8u2CmsyJIsdiv302ILEFPYSfBBoRjdR4QQ
3MpQegJjvZbZxGyHN00j4vYJ7u67/3C+o//HnAnbHlnYQZ1RHAT0PQ9Sve3jMLBjbTjoQns4AGd3
H6tsP1eGqomZEkDKGXQPnaWsyMKsS1cxgltMyvslGkdJH5A+SvhuoLYZECuNsVT5jvZcgoOs9eJT
V59704NmRCKeiioeNtM3eY2ZPED2iRgtRr7tekrqjAHL76yQjm1o7LZfNG4UHD6XvLjpolT/GKRL
8ong8PWDudrRk5dvbx3tcO3zHyTUvdf63hvyCi4er/Hau+fCHXmyiH+ITdp2hw1V4tCtGUMX0cPj
C6OtvYvMFYoIQ9+hkgk7cdkOjh8TIoVlVLmTeUYY3z6cs8MQng7I1GNJn74WBe4Oy0sJjtz144Zl
Qz2DnYLiyVsgRW27YkAbcZMJd6Zy73tk3kIm8Qiw7Ouw75usyDdXbOwgLVH/sNXc9FOVUPpImjpp
TGpbVOFYlA5G2sID5Y1cfCHYoPNodyEfyfjs+NQWE9uilNl8/NrMNKvwERXZinL4P00Mjr8XfVYm
dymsi5e8Lb/uIq3QGD2NaXyJIoa6u9UbA3dRgz+lWcRDit0gr98wBJRHyKtGnjggAw6xBmLWlp78
BHEgy7QZOk3QzO39ieDLlcdGd9zm4ZOpGleG0qN+ka2E5k9F0HZxzwxQ34Lf6FwH6S8qtq+9bp16
wZYEKpQrlJLzalIrd+rdivfJDbPy7yLPS8on68xrdm1N/1CovBhFP2AK8GXvzL6NKzwLGfOtbIcQ
ce9tAwFendIMqZSsFrFHCr/U17lJWvn3gjOwgcfWwLfNtVC7Q1Wzdn6ycJMg1tMEESXQuFiREDxN
WjvUdKRW8LepIWqGqUwN9vS978l47oe4YTWu81W9GIB5XzrOzELREEHB2awIwQz1XDz9URzBS48c
U8QNKAN1f+1RkYVZBhuzAmvF4LxIZgrZa5gr/VeHYRCWFUMryxNzuRAy4A5AZPtLLpjQb2Wqc1DR
GSeXIgfByPAXRTt+m8q3u3at0Xnl+3EvBTYmuZNkb9Tml5u97t/tYCJi4SHzM39RtJVihdsUsmBf
rkJXC56aaycKCXvx2I8ORz79ObtXYT6nCT8K8E1htu0p9RIxV4PLuCID/zjwDL1bEVrTEBaTTLsT
PqeLuby3MYb79uvhkHS4pzu2r/eKgDgFRO1KfuVJ2qgD6Rm1GBrrh7W9Bw/aEE3IDa2E7TkeI56Z
ONsdPU2FsisMkJkxdy/ui+/XaTOa4qC0ya76Feyu0PWapZiFB7HqIDxkxOmI5JnROegcoP6DC19n
XKGBqn4M1/Y3m7LKGtu01Wfm4uelvHd3cijIQ13MWyx6lIyaGRwc6IjZ2AUl19Ua/cIH3TuhfWS+
AbY1sK0cJZDLb71aFn/tP8L1FXiNnA8x78n7AZ1P3eKc6UItTPhsO4X98VZB2FwHQZ6Ig2IG/yNr
KL6lb3X5eutHlYquH8TZCcmzBhNXNdkOwWg4nmZfm/wijtxwgiHPHU8Q7kb1UTc6W8Krt2UEVEyK
osEdpK5J7c9T6fInW1LjyK/esKo7sgRar07a/JS5YnFLqAg8AQO01TWfbybYy1JNkdZVw4Nn9JvZ
Kl7VH/YgB3nNvGx/orWAkw4P4cdjHNOF2LQFRexcCVvy1J+xJ87us5UbIokGAUergioST0FnArYA
0qZA27Hp4XcwAaPTIymYhS5QrVvi1ihtsbyVlzmzMCpwFvEcBuH+1gFFoqiwYLnMf52PP5x9Et0l
e1IzUcnd5vnvrUCEpCqdbzzV0bvP2dB6xri6Ew9DgDC62KKb5QYxaOWGrdEWyTm81Z+2axGzsbhn
kRCOaZXf792SqvcuLzsm60G7S99OPVUdkEZafjJUlr8HnEYRaZLAZEICJx3TIuoFdo00pRsKnvGu
gqEsN4q2ly2LxRYU/PztlrL5+sr0GG0gHJwWTRZuIHQCWh5+LTh3fuBwwl1zixd+rPvn5Kkmfii7
nHKnESqyHLO0byPweU+rQOOOp1omdc0AEWt3iYu+umSkTVPHnEewU4VWMtpXEegeQUVDtrbfCSib
IvTc3ZreMS45RM847UVQm16f/wiRQe2j1jPy4GjRFGN+haCBDH+IwC0V3NQLCMFD2Q9N85DdfNGk
gGXBItSlaXmWEJbo4EDvTZZOGtGQdQZ7b/2Qd4ueNyL1OovS5p9hs5zGZkMlrTvEzB2f1xFF24F9
xZKd7s6OIkrCwZ8p+0RKFIxkDqDoV3xImKRJIV4OGqrPmS8ImA3tqZcmsQYjQSL/YZYt1kR1TuV4
Pjuhsvl6uiSbH2uIN1HtEiWbqaC7042W+rKkP9eAWh9qvzOVBMC04kWaqtakAE3Nbxkda2SewF/i
9h1vuf3hnzXWuljn9dHTotPA/pTMo0SDQ5T2A6IUPfAqZrBzX5nqtQFxASJVslSKhsvnqw3Xc4Ld
uT/SpAORPv6VXyvJg9dVpuqmIV3euNLY8Uy2PQaW2Kg+N1ns5ZUKXyypnzXRV6fi479woKUM/WZ3
ewzMkoH4f5xHvGj2QjWOBW5TZT3pUXwZlTKvM0c3URCY+drzJ/M8QV7DHNfhKilOM4N58tGTUqyo
t7pHLTZrWi6kzPHYNCrQYom6a/PDV7WodBhTCwbqVArGQ0QVGhY3/XPbHbiEKwtlUtmgVApEdgxf
3M2jh7XXQkeB9jHBdv9mhWihQQbE203ZTOifA9b4IvAPaNXc1DoYlDZF02Zs+gJ7nQ0OvqxS08ND
QdREN+0uMoookTv96ftjrWVw9fgmpLAnhQj2tFrx2lc0f8RoPiVg0Ljm3fD87fAh1fEwy81yXER5
PURBp48Is+jHrttGvmmhRcyZN2naI6xIHz+fbJePb+8qnOouSHDj1Z5WkIViznwy6iQ4Odp6yeS7
AX1a1IH3J4zjboePvpsHGw0xwxXaxcJsqnJh7ucGwzdUnUxz0dhbhKMJy77f8dVPRhMSwYkt/HEj
eVicM6TeVWmI+EldvZb9WBuUYJ8uBoB2eQGSTTFnKJ7J0GNdznLH34de8boQhODl+PVQthjLYUIp
qS1lngKl29oTo5T4ne+FUpqvREokxVgdYW8KSTF2wBCDokvFiDfcUEn1zckP3PIzURAmiY+omvG7
U4p7T0EA2PmSHZuE1MLsBc8PWrh4mV8ps6edlyLe6cFymqi3kY2z5mYZcjJAYfMISfzRRnbzPFs4
5X4Iu80h8bglLUazg3bMRgHUCaHaOHsB6NhOKciHyYByV5FjuYIce7BtMY0s/rwulAEEPPm+AxoE
Mf5VYiIcUsDO4FgbcJBPnPYP/61KaqyoS9Me6wYo2wbzIkuVEnbilNDp+6ayF3E7deksZ+Ff5jQc
p3ZOe2Zub3CRqrM8DDdg2OiVTIAZKvTrxeI/v1NW8QfENrShWZVvi1KJdsr5qGGo2ikavfcqIGiF
HMo0IGsNyqp2McxXq2Cmj871fOXJ9Dv0mq7P3aSfjTtWgaxQyWrRd0w0VbxewwSbG/WaUPnG0Oo1
OdPBjDTcuDz2iFRKCamJi+v3n1s9wggWXGpVmzTKLW/A0LWXQ/YsU3VeLjoHoG+HDoP/NCxCmeH0
plEaDwBjIfEXi1xgW0n9Bgk2C4sXjLNvzaXN4BQ8gP9TtgZqIu6yu+diZBZmRyT517f561zWrGM4
45EsnRB/wm0UkASHdFVNMkkQCn4UhWzzFbH7dYMadncMdyl4SP4Ke5tX9uJ0g92oNvb6qQMyslJC
rqHzq88w5XUWNuWqWCInY8Gt1vO8EbkbFZbeYPalhZ7IsB3iRoSVKKf75pH953TE8y8zndLI2brA
ZCe8LiZ/zWt3xuFfkQKTaUIMfvhUO7YgMbLsX3INpWz8AMfB3CXLsh6w9asyvgHwTezsH3jiwtrK
mhjk87MsG+xGeH8VNc97BIZVvbUtDx0g2sRBiTzep+V8WSemwrm/9wWbqvroe3s08QNubOmAJZOA
Pl01lAcTQQ8hReAryuGpP5wrS4mmhyKex3Xx4WQaUM36R4UwClw+ZN6LzW1fWOI3IXAZb0IExlVy
SaWX91ijlHCaiApw10okL2HOFIa1ZFV3yoz7g1JIJnzFSfMblZj0q/80oyS4GaUrQRywFkxAKbi2
KZl31xnj/PeZCco9UiVdTf6bcIIaDfcxdl34zecxEFIV+0L7I5I9JAbe9PBodnvYFy4u8PP+xKYO
Zl9oskSpqDlufINgZyX9qhkboLy+upx48/mp7ScxilMaIs6T+155CfVQ5nxDt+Jd3/XdXWrkmJlh
q4UwZ/KhsLPJdachIXrQqozpmarlk+2LS7AVZamJffLaOruVQoaPqeeE0dMhDt54sA84+FMjCP9Y
UDK6le3gmsEBCcjhYY9+nNDF8WfBoyBo5OrnVuBpGv2RebC2rEMyg113ZG010R/oEAlBS/FcEFyI
YAEpTX/eIFZqG134s55kdUB9tVwMcbWcAxxOfFiP5d2NtQbfCmJHzqGdEYM0Chnfjh/q69elpFrv
GT4snS/4o/A5tZj+g5krtenO405MVqlIi7rlIUzs0V9lMUb4PfbV8hAcdBrY9nopmK4dcsrwXkW1
vca7woHwlU7L38XeXO7RK/eqNkxrf8GjWe/R+otSdfvHGS6QuSb3gM9Ktfm1tNKy+XpoQ+K8qaGP
82wEbSeotcnh20eul0wCNk2EkBg8xs7SHQnqR/MjbArYKBqwViN1zgqMWItbRoICr8PJXbW5eZ+t
nqCs3zrwPB+ryIz9b+If0ZJyYAs0loCkpfNyf5STMJ+zIyoMGO+j0H/FcGkM8HqQ2gnPT642S/mz
+y7eS01V9UVhNhg/Wpv9pGIP45+HWOfmSEYWtiv2IMKMd1yOJ+phvTm0719tb2IdMZOoF+7zCSRh
G45v+eCnethpLmQXLuVPkwl3DlJlj/JCHGTa1zbNpiQ+vGtcIlOw7zkP1hjC999yrH7xkzr1Gw2y
K+mZaupS4mD1rIdvx+QDzX5zqZZqQ/4X7C5meAo8dB9JkWvtl4B/sZBmnk1J9JixvqqPJ326TkdL
gpkvlOaJnNOC0wjrahLL4F9pY24or2XEjmXpDbISRhZ0ULHHWbNhnVnwwdmhSkSdMbguWWrL5nFe
5IZFZ1C/lb+hegHJx/N6r6Uusq3nAMKiAH8mPoFgOhbZFgGxnjWdwErwtZshfq0lf1fFQJjAv7P2
CSy3RQh65O+buX7qyxJlPfTTQvpcpX30EncmjaClFRiCqYoYNRLmL/km7GCjVxITLbnEUvAwZn7O
8eyjVGFmg6Q8CLs+7JiIlZwtTfgppDnedwYQn7i0g+YwnAnpEDu9Y3BV6aOOFj/bmVbNAEC8hE5g
Mz4hEigH36VfgVNn2B/WifYTAqC7cl+N1U+fHtCGvdu/k2l5qGmfuXL01szIXSc7GKWP3gCCSku0
c5Z3BLGeLwfwekcTnnK0nDStFAKC9Mm1Ew+xvlzQTB+lFAuQRlYctSdFJ0HCHgwxSwtyBji8PdJq
oFFUHoLripSWpw/JsHemP31Wwv8rH6pIVmFu7eWgBUPw+fw1mmFoYaNeJhOBhhV8kMM8/xEqnt65
KoUfvl2APrgpmSTsXPmLgDSOf4eFAEYPNXvXdrYqucLKNhru3+y+Kbxm+pPTQn/GmfuSTtrKMOwe
hWi00GFWohmf33xv9I0lLnCfltOr+5kwzuPo8GERPsno1mSnbaZ3vm3zgpyPIwx/FELhopmnQI2X
dTH6R3h1PBr5Wzd0Mr1Nlqd/HV6aYVkH7BIEuGdPE/EKOTlGTCtCYovs+R8nC7JjO/S/LXlFUZIB
7Is1NlH9xvB2UxXrDSFF9abttodgXXVNO8l6cRypyi4QcUge1VaFGZOPdJYj5eU0bB2b4jSsDfgA
KrwDgrZpnnZGkwGpHacSDPi13+BsqCI1DsB/M7eji0UMkUcrF1uwOUgqfTf4BuKaqwF56UDb2R/U
OofGV5lzcOfM+42uK+EF0Cr9BiT8lgAZ5bEttD+9nrynX/5mMYNRWZ0ZLLEUs3wqgcbUo6Pw+4io
JhoXiqWJpQRz1DvOcSB7GEUDRXFcT5+B4hJRRv5BnECxOzxfekGRA2fbTNxhLL3wy0eFkqQWVXoP
JZal+nSIm5GcH1gCfqUy86Nayv+5f5iu64ncLEM8EIsP9lSo2P85ZfbNSMEK3jxeE/Kk7bBLflDF
3tYfysKWt7eFV19OnrdezsYYw1bivEoREqUWaaEHifuqfSe3E48H6kdKnR3dj083ZXpfAQ/4Xam3
NPnPWiINBltvpQ6a1ckKPTVEsPT8ttqOZ8WcJt55HACGBD0l9/MFv3AFMXu6MV/S3l8TAovzGBO4
U+b4MjbBZNz/fdQl3OQDvJX/3K0p91sLrBCacdjLxxeOdy1ALqWNscx6/ijUyo+Y7cl2oKyVYf/S
Qlo+XfHygBxorXXEZ2MTg3j8e48777JJevGZjhok8l8RPw8ExFDPpHdA39v4BfX7gIcKT2viedE4
D+vj9STTvCtr+OsMvLP8Uy65iXtXKirjRF1gX6EmuG5Aop4FuEUgqnyYpyzCjwdLI9NqwdmAMtEs
Nk+RKIH4lx52fEXU1Adc33JN3V38pvfrZl61R7mVaa7G9oIsGUiwTnnL8ElcVMdJ9GMa0DGYjw+R
13ThAhc5vvnJTe4jIw2hvqpzwK9wq7yFh8bsbNdDEPvwfAuLBrrFaTwr9fzz2y7ag7Qt8nNPULth
Dv5GdG6eVguR6DcsNtWWuT6kF0+08pPbhp6kH8XFgKOFroMjlyT25IsQGySt7Qv/hs/qAbxA3sKb
VagaO6vGFw99d2iJGdbc3FBOC3AhaKCcg6JI3bxLIX1kJRemBBJqw0hZ4UWZYGLocM5pP2iTyObf
w1T7ajVWrCOVo5t/PxgnEZ8RY31mAcxQ64WFnO8/ZK+kCcHQKm8++do9Jvmd2U9DwnQ36KfgCRSM
EQwqanEs9zKETvbpxhvAG5aTLbcjL1GUffPgx5sdaPpC7EjAtQ5srnBGWSCcIINOGHxPli2/Os87
9lk4PvxJuTClcnZuSEH9THdV9rJZa4CL9jIOD8WFNqtHCAUWTsajuYbPtCed1glD//QZNQeHc/76
EgVmiM3HsWurPsieggW+/8cJKaTXxnN/bt+K+4SBPR2q1ZYlLah3bs6qc30NsBm3BzO7W2ijcZWx
pYB6/2GbCn00CSZ2uCocI68cAe5cXxHHxhuvBFOXJjUfc0BpxU5Tsz/45yim4odSO8OREsf9QVY4
52GHHTy23rgQ8c2VeW8+rf2FHfmLZoGo03hd0eqBtZP/cmSMerBB/Y5MbJ+9Ld+Cd1Su+mv74ojD
QmtwVy8CKLzpYa/KRcPDWQeBYh8DCgX6aPwijyraF5o/syD56VTBijb0n5WcaciaQ7G4DvAYNrIP
Lv0iLm9emRmhvtUxblYGwKYzDGgLwvwE885i7dPkE9vqCKLRKbC+P/sbquOsERtjxdGn6QZtFPiF
8GBbyekeh2Jk0VElxmERKt34ic4zXaH3T4cctfOzjupO1bA9R0sEYy2bqos0jW5w63bujmECB8Sk
2CTwclSfSGDJM85i9dtZCN4h0smwMwraPi4qg/iXQubwbBialhuUotddAnqZaoPdBeItwGTuYdEO
gZYE5UOFazRY8IGtTtcVm7mPhA1vyQOMoFtB6Y/6Eo5NHZ8ha3FE35fF5rcRv359LqJWBDfKIIZE
oAJAa2hQCI/jCOMq8weslkxDlvFSjIYZ8wnZBy+z6BJTjOSwx0SEiRqY5zS5qs0aBqsXN6uR2ovR
GBv7Z4l8oUDR8nCjXDNDZtW8HZ7i44AkbABQ+7vwH3rhJ8LQwc2UwAuEhrJizUjJ+cBj9Mo4O0e+
a5zYh9SXuMxsOfX7oFI7MT2awfskop0GsypvT1+zO+StwmLErVdM1OdSwp7PiTOiIy8SADgdRtuB
gCQvwCE2nBq2aq71D6mE+JyYvKCSXG60DCqCAO038sUU1P3Se0ef7I3MyXxG9z7NHdYhZEz44pUC
7XNveUW5P15A6V1+N5KON/hiKHQ5UEv6A2WT0HhrjSGmoIo4/yiUoOb49X8hF09CMMiCYRZ/CzOO
kPP1pwDfInYQnNFEWx27zFAuHLK4M8arSIjXbZFTei+MYhg7ImqLXA5EB4Cltj/FESBcAdQRabHC
fFs0/CgD4k6wLHJU3b0XxTlxCfAUCMjYWsClWtfvfC/YmvpJxRQQvH02bjlmAwN3FLnHeHxPMee8
2BzUxH+iLdZTqoNGcbZjQZJt9NCKRDFwetXl+YiZnimPq6jQUxw2FfRtpoPquUrbfaV5ZupPoSyU
/fVv4GY6W1b9WaMke6I6hmFaB4riPG88bCJhC39fTt0aO2SLGN6Umh26nvE00DNBziWym+qZOCeT
vgspa9UTIXiXWwbYY0x8GY2NAx1Wew9akHZ8uFSbqVXmV7Ci5WjAZQafBxQ3YYADW/tZyIpLNzNv
kdvPiXhKuT9Ep6VKX8qMLbImHoCemSC5Xd51anjOWNhedQmeiQdCueiZehJYwmSAAKZz1Q25c9xz
DQKO8lxuZNEvPE1MD4EbOGvrF+doEkisRNJp+3kYQ5n1dnoAkQByygDrWHcYGZ1O1oYVSRJu7FeG
PTn+k7+mbyO/SIC1S+8YdctE90/7iq0powWwc6vKYxs+GRCsXZXKA86jYnvX8zBJWmh+Z/JHjnDG
KnFYApVEqUvozH5C6F+ICmE7Q+7RBYEAiSOFTd9Cxoc5OlvQTMzGbilNccJHRRw3bdLM0TFFZXEj
ol/Lak21rDj0SP5djDGQ7QKvUz6F6l8EQuBrui2EEYEmEHBWIf6zs8hAhqJnbejfgc2MnYRD8rWE
8RyQEEgn9p7r9AshW5fjcYEBrEHxIBdJLW3ZoxmOatodt8fn6mNF/dkzvQibqUw9DWAJ67DA3pN8
o0zfIxTS4Hmh9lUK25mb783p9hf21p69QPhq74BCrUawMCSgs2ca6vpYbnBI0oSovfMpJ/T1WUY+
4SsxdFgJGmom6QHQrgZ8U/fZwrDR2pPU364AgfK4UKRRpWz4w+td3koBJ5RCH1Kui3upWTSgxuGu
hIpAExW+MPDPKOe/4mj6X4nRM1qAorvXLnsCxJaJjmxHE/DB5MAZSOABV2HjsVjwzhXB6NphFT5C
+1NwwImDKRzfOjKplbDN/+NPGInxCGS7ORj6hcWSpcXM+0WVMJ4M3t/0IwsRXDVcs5wkdd2+mX5J
23V9m/8sB+HQaR4DmfrRc2Q/dIXg1UZ1EqCqjJMljvFcmLCzyLclEXOWBd8pje0E5sBwUY67wPXE
zMQ1F7qfhXLkpUqr6SQAq5nvIniVQhWITDV3HbZ0fPWp/Bn6nIfls4PpEAj/rqXpSjq3o3MKGX9T
QkG82M9gLYdwGhb6nhU1tqUwcYhXkG4FMp9U9CjVrw2GKOwm+aZyHs8X0Qed3kmFNFcsDXoattLy
JCGldF86i3TsA9G9tubj8KVLmTKEcYilFcyO5/0oiQFajp34hpRZ3SEn48ob7UCoJtTjau5EPdNA
5DgH9wRyIjJjiir5iQh12u605o78IYRy+xWacL4pnR+xfoSZde7R63SSsOHWELZqJMaHqaF7i69e
1gilQn18W/bfu1bFHkHshKck4UBd10fYrc1WESPO3TE2yGXU9j8ozMfz+E47IzLVMfqoECtPE3V5
WNBM+y1ZFFkK7bTAjXTjpL8AfTay+xRzkJ59S/GRoF5cYgB0/jN63OFLWYFlJIraIbKqsdNO+xtx
k7cBikQwFJnYmd18YVO8dvE2SjX0qwzuUOLhquCyGMylgHV0M0OCqFax1WbldumCuDcfFFicGcFb
lTZkQSBGjQMIKsJeQUI001alhGqfPCrEFXvA9nvjMoiQsr4z9iGsqmGqaktm9I+VoTFBSozp3Q7s
Vf+FOCgVmJX406VcygeMcciYXMlYgSkyRTSlh7M4sCjCy+bw3e6+vG6Y70db7N78bvTTieUoJvGE
1UL3UQTPbhYDqyhmnKxEWYCvA9AUDrfIKbgEPQ+tblYjBKIoFoNwDoxa60k55RQDz+UiYOyTwRt+
HnXdcRMYQdrafA7lslrHpFaKnqdw1tXom2kwfBSyxXd6ey4cVarGLe9Z909xiZHZoB0l/ZhnLUKo
hQWjX3lufbH9eJ20FEtF5GCxmYGCptD7GmVj1DTmT8y9Ibl3svz1EMnXfjt2fe6+sCSRVEZavM44
O9wNmPbBhp5Rx52mZLtxd3ZKfPdXzHW0KhjiJPyu86zK6bbd/2fXT8Q7CiQUqDedkm1p9M6KYPNe
cJCpxXoiuOiohsKmjhUBAmZgEpv+WmVRF61GxIJ5FxJriUlzgUcJkKgiM9FnOQDINz4AK6nwubh+
6f4bkFce+E4Gz260F0SHS5HmL5Af+jjkYLHM1dU8APmHAP/ow1/Qf412Aymq//zfjGeElhh804EN
0CpEOrXG6XUZLgzoS+Vzvyemhcu6UhkS5eccTStEVxz+iKvouE2mkIIFWfwkLq+fXIrbBxlxkIcL
wnQgzyz3eMnnyBUoPLVBJi475TwqJS+m0dO5wKQYbSNSraJmWwuIMs8xPfelxVvYdD0qL14i84yY
ZuFsrQlRTwdkKbgnZWda6yTdvTOx75NfUIXgPvD9a27kntVea5G9WG5US52jGfp7SsyqfVXCLC2D
GMHAgRj9OPpwqANgANQJLpGcy4WYL79v1bejJbs6Mp7Ow6gaY7rSm2wqjOOfjBgSpMrr3iZ+b5xE
pon61DzF2uXDWE8g3JNKF8ParzcMVEyODQKWHO+JXFXzO44JG7k+q1xEeowpydRTwD4VWjhRe67m
YCHWk3pXFanczlC78CUzAOEwFfyrMtM7PbM3Bl49UUCruthMLFfn2jUdF7vVvMkwXO3GMjKLOhS+
rWW67CpHv3q9TrlOcOCpTO6laYCixVA8n+EA/K8Vy2pyoHdSEQyYwdjQGUFI57cnZqPwbH9fgaO1
YCXHxwTrHjoetL6VMLt/fD5+HweXxeilPncOM4jfeZbkSBt69lp0ypfijd2VoM+IgxElc5nNqTao
vyrv74o8LMlOSbi3w/2ipDCTBjpIXshvVwmsCXe1dFOOLPe+CsWqxs7j9PhPh2uzQ/kPDCItIcrV
tFAzxYXsH/2py09X971Cc9XNpgHQumI+R+xggVF7+vRGVtEie7hx4fXd7NMxFgthZQ1dKJPrSQb1
govHxwBUUaW4BnNvb6sFrOmusfnQRSrqYe/0qsuknPP0BFEejdVQQ/CHlkVOVe2oK9cJzOx3s/56
1rHdI7fgLyivKckmDZ9vnkw8aiBngyv/MHCtp1zPyOmIOip8MT1u2AtbCelUwfYd1viuM0FWGtfx
Jb7xNVsFn7biSNe1nWmSjejI0Bz+U4R8rAA3mpZPkV0c0pAAE8KzwT7AuWK1Dkky/E+jzhj5wbkV
0JUvnzHw0TkUcz4/TBrbDTlZcOMfgij2UT7QFtHabv3afsTa+hQBxJcZagkATeAu/eB+PjxnEPjq
hmWdmtjK7JQKdue/RsjTTDpBPr5Xw6K8Q/orhws0aAydYEx8/YEjV5VRmmLFIAhrCkFqijeYCEn4
8tLbQ9rFpRMZBVeVAitVAQHQGdDsOl35FfSHZhPFJygF6z+GcQy2nDRQwViucNCFc2Gr31RJKLpR
NR686il/gkJzTiuhWOSCzWSP3pOEes0N4U52cioAJ1V8zKsPWJ+4cmzQlp9wgtTIw7myVMP1DEbV
wv4CB3uSGvMk4Ohyud7UNpJ9eQckChq4IGoYGaCnAGLyq7zhDfn9NPzwe3SF8ndE1InW4k7ntNCM
R/qp0ZxuAPAAdqu98teCVPBGvFgnz8kdeCklbKrTRIgkDeXQryQKtGmM3sIWykMAVKWV0ZXM4D84
4zyWt28EJjuQOpglUY9iWbxKX6d2or+s2P5Vo0tKiVAu2KRZmZkqAQrYzmk2tJzHbCcjcUqdQKIy
XTJ85NIgYwxBLQJ2JRWXO41Ei3r9UjP1TCMC7YsYaqCDbJSZeSQeXhRIwBVQ8aHQzJst+t/T7YeQ
FsJic1ayz+2laZQw+mRGCK8kfhRSnDZepxPyNNxYlBbMf+/Ecsv7serKYsbXW8HL4cQoPDrIBGYO
4LeuBowgoojfGmmGPg6Cf850Ndg8Cur5sCcQ0KMFFKjbYUw8euVUnJKvsbWaPjRnehwJLjkU6uEy
o7nlXXP1cP75hkljn6lWrMm9K7Eevt3xifn8lawVTH/2jd6Cvzlwexk3v1bKZYpYrAdEkoOYH6Cx
5zBh6u8/oErZthfT0uPK9o7E4TVlHBHsSQ+eao3k9wPgWuFkiVVPTkk9CSwV99m/HTwLdxtsZTt4
vaSrcXdIIVLNe1QQJggLUPR0TM48NibNGIxqMVeuD9o+UXZnMtX6mCIk71L90NYmHiTgpCQefBNg
wjBBLo0mdvTSvW9oyBtKBtjGvr5JMyvLWr1PpaT0Ff3ShnMnkIvwtsTvB9xWQvVDhzHlmqH8pFNh
GW3hnY3SdxMDrpXtIY+l1EAmB5ndxP5YS7ct3F7X8U5iHiTmBe31S7T3dcEPXGKgzhtwjzcyIVY8
GVqoFH13btvNb8+vYUt6D3pNgUFHHMXHSKoPkU13NwBNbKr2yOb9pjHjwOozddM/4RL1GDbcZEDe
KV9Bcnwkz06rhctYLrGUTCdadSukBlRRhVKnxs7krC0kc6bOiTMzEmYp6OKeD67Koc0cy1GAu2T7
BshNjMnF1ioHGOO9JinhezGXgS0XrOGSHQOrhULks4l9fCjR514ggt4ZvGwmrlGo+pGe+xO65UqB
LcRmFdHB/eXZjW9DGgGFkit5s4+gaBZN35XuuKzfUkAr1VHQHk23HIu/U50hiIkVNEpXly7cLxmN
rKx2g0bLoMrE6GNNRXca3HNgWasCA0iUyGmV7qnSCEtZOfA7DcDW7u+0wKmEsoFyIPOzMJvVpEe3
A0tbpxi7bol1GsYHxBj0LpExuij+oiGvS3TouGcfMDd0eABJL/4fujZN5NVPeD2zULtFP/kn1J+V
eZHL+FzLkAWnOSRgGugh+gm12pKX4TjssYg+nR1j7bOLOxCf5LkpwvQUB8QRbNx4801/azE7qrYp
FzrC6XChU63xt6L0gF6UnZYjmehWZUS3bdSUna/3dHf2r/IVi893FZKwx4QxGhwYb/aiuSZHGq4C
CWljhuSKzpmyms4lMF01ucomkllDDCzrA9LTQ1Cijkm0/wgYNF8beaKagA21LZpvKErgfelGJ6gv
XxveOJMXEolqje0R5MvtTNGAy8WwjUogZSjJ7SK20L2+PUFisXLX7saF6zWCZll38z9CmfjrZvWt
pXgn+7l0jo4DBGDrEPL9c3YTuG13NKVrr3N0aKYqe5CjzjOFppu68K26X34zleu8s3BQGjDTLBwP
Wk3FoM1SStVFIiw64dl2RTw5kecDWnRR4iE8TTkp7DtGzwBpAhDTzObh1fsb1qSN5Nti1LYHH/wP
m0oPSeCA0V4a390hBNXhNd1nyznIYeJGdwrYZPwu7tQv3Mq1+OCTK86E3o+ApbJBKz0jrzlN+YYa
GavWiDD0F0NY7Q+s/eH8ciTcnstoAaBmQMHLGu+Y5n002XZAgm7SFy1dUBWSVELyw1D3Wgiq0N8O
UB5NTumZmm0AbgF6iSKegt34hPrzwASQ8Wgm+B6qi4kJnzztWsQHVmemmZWvS4rtsmh5+Wo6GOa6
IRQCM2c7U4XIY2nxPdfQww5hxMbLPhB9FLcrtt/AMUYYXqzkQN/HkEIi53+kEG9od4rnrZNwEAkY
folAIoQjQ6Sj6vxQgQojNlU4LUB5JZgoUbJ8rpP9NL7gk5IxH60Vhn1bFDPUqBE57inDScZsS1W7
KstQCe3if90Qr4zOtUDEh07V56kRi3vchJM9RX64ACuS6Udzn051agoTF0l4MpR4GqCctjkI9hpf
VNS8ukcPovxYLLiUl/Z8cjCPEPz2SvwNQgMDu2jkZGHNCN2lOu463mFBVm/XpkOdmGTTB+YRUfRn
XOSoKS8dDoeCfZM3a7ABBxVRv4KzP53hGF6Yp7FX3HQ7V0Oc4Q7sF/uhHKKm8JlRktTrqU/VjWVV
4Fgo2Id2iRw/UadKW1EdqOouZVmRHFQmHrjGlREgIxdfgJ5jAQoQLyrKbzgy3lhw+cq3Q7vxMEze
rLvvGPK7L/a3noGj4Lf2Or2Ufb13Mz2B/vWYFZHNlISUlWQBOXPKc0mBMNFBbHCtu2AMdgY24jL+
hLIcu3fAXn9tYE934QbP8Ia7x2fixOHTqIAU8ts5fWWqFeK1+kS7aIjY1DYD8EymMs3DFj4WWD4E
9Ec9cwun3eVKK+GrD/8OwVReEALZ1vV/ISUDmHLqrjrDJOHwLhRbf8BlZIgMV4wVe7FgMBLZce+W
laqaiUq6AKLbZHUOtZIola0R443qW90/CHkB0TwA9nD0vp7IV2NLae94MUZODgHmJBDZq+cZSrJA
D3P6qrW7GOExayMwusiVzuPo0hqF5SxXJ8bS/6N3jj3P7Fhpzdym3ZrC18Fvc9v4aDEldBgGd9+v
IcpJTCb1OP5deypk9Zw2+Q97kNFK4/fqITdKcNWmWz+p3VOh4cePuWNVn+L+Ksd+RxR/Z1QiTIqq
ja+q52U3ceStddqcqN5fu/lYmcAp5x4bZHC05uXsjCXpywtwWjdBwIyNflky3uCI6DI3tKbvg02e
Zw7uiLRy/POZfGUm0RVCEqgVvn4buXuLOQphjQCMNizogpcwRoW0xSIDInViCdsWRV75YH8mFl0M
Y5hVwUxzqJMRyNXF5mIhLcdFBJbF9VKqIyJ27jz88m6DpCWN1sfPd8PAlzrlY9LAviZ+8w6eYaqC
ryDR+FcYotHTjTRGH6Md2K2XmX0+8/8JuPp428Kg5olfQGmJzShI7ro4Px6wbR//ZiS3ARIuFjk5
2vkNPLwrMmi12o2W9aW21vN/WTQGKWaVOtoP+8X03FzQaV1JQhiwQbhXVoLFtMpj72flU9aTZurC
OrBiyrTNbPAIFSXNufmSoX5yuJn02Bow4j8JCGaXC1OdYMbeVbSgJejxQPsW1U9vzzPFWMBIelmE
EOF+SgakzDAYrLE6MKy/mhtJpNI/rwgfUy4BifU+tUC22rAj1YGmBT1XcmqeKn0vILt6c3gnmj6T
neZSdLI1M6g8OC8qQ574O9Y12WQXe86OwQ0bj8tg9+7okMzW5+UbTinq7Jt2YZG03MpUzc4/BPYL
chr9Nna/ER7QyfZGkcHjGHSSw6qCvi3rDZ3SxTqoU+BsKzXvehCMF40hkCvlK+S14XNFpoxjzojX
SWSigBntdVJkHnLjec4664wpy0airD8zs/TlvMCUummA6/sgz6KVR4V/FnYc102pOxHtOl1dYi/z
lHEcPn8zd4yKdWbG/OaQKfb/GDbdDc3A144dEVcMWLykOnHwnhpuQyk8umHoLFIJR5Nsa0lo7otT
XbLBPxfUD82Sf/Y46MmWPfPyZ4hbJDpXg3R6yhZx68qirBubUI3dJSLlDvW4xmKjHklNeF9E7L8Z
wA05vomX3LY5pud+trsEI/HW2ct55f+4jzn+G/Fzg1LnnsXwjiG4hWYWskBOoyZF+v0nsnmbPiPx
WfSGO8A1du32tKI0Xy70i0K9VYJH3aT/TbG0N0pXVuYkxmwiBcO207lZE1wfi94YfI6rH1UB/rQp
QPQazA7fAHaBijbpLLioWg5p+GJ+80VNNlexfC+iNifKSw1TfL1lioUtBDRDqt3vQUH1hce+pE4f
R3drKuzO8rIhWRZXTChLU+pyVsdbKK99wBK4v847kmg3rtZadL6aKphGpzoZSb5HWVaCEyRFpKuu
eLuzfAoKA8S6cLuYSaOl0YctqvtYjRU4xusKvzK6sw569FGu2NEm7Tz+EcBXVY0Rmw3/LKZNuzeb
SzhOYoHcDxqFgUL3i8jwZzlrp6hPAzT8nLpwSgqhu51TIEhNdOAA9R4jIeQfj/vGsJnfgLXC8nn/
fgg+z3J7dl5yLyHAkgGdFD1rfk14AWG4/PJ1Sr+gSMNo6IDd9EUBckMw1j4E/1V7yf4wItY77Erx
sbL7ewUgI4rn2tRmMkO6+fCZ5C49Mx9dGjtd5Xov2717CDOy1A/vSjiwcToP4AyjkgXZlHVWUvaD
6mHJr0WwGomP6qgomcjMtWMkFoF/Ph0j4/WQW/77HGWZYpcksOR8aX4Oi+cNS7FPH0Gc6kd82W0L
mnOK1jIrpKr+5SevaQpMXJLrCLS3PHuwVWR83+/X9uJUcALGorezK9bVlcNWYQ2uNX4H++HKryQl
PQgOyffsIeh3Smt2/r5xNZmf4f1tyDWWp24227/ShnWeuJC0YalkhNyVSuuODHeWG7UL8YqweQs1
DudEIHaUCEQlGrZT/JOYwQ3lr1xdvXrIuY+KLAzizME/pfs9HLsJExOPQKDyoV8Y50ugz3NKUA0v
aQxfvx/pTsf9RXVP0bItZ7wJnx9lfv36nrSeZ2cPNDHsFTsrF6nq3qNYvRRrXzqgNPpbWlU4naXy
3nIR9IvJdoHhRdpOfaoDPUBBc5MaerqcKF6615f4+mcT6qxdqyoequXl/kzfcVr7hyp6bhcuGRyv
EOOuUMfww6Mxrk23AI43AUltPFX7xeznpxgN5CgtG98AWaT93VqqwpIDU4V444srLLJ9SO4fOyMw
D2ZRJLTHs/wdWYanrnzv0H7y/s9LqNGeqPcVfhPfUvs/+yjKJLmbUloTCXaphKkr0BgxlXsY8zkD
mfKmOkhuG8iymFUmwQ2/b6MZEVujF/dBS/FTxeydAG6ilCQmatWSycE0Re+xxrqyBSJQdR593G+X
flGWG2YTX8EHy90L5c0Q5ZUWJZgpcGojShUKv9buAVlu8fX9XNxKMd6mgDXOsIPH2xCdLpWIrU06
k2Ms9UDdPZGaLEeqj2eHlPqCA6/sQIRR7CYPXMQ1rNXSK4fAtJ+Oehuhj5hdpqyvTvtFgMnbDSsU
kYDSh/MfJ/tT36F/srb9ivp7e/i/QC1q4zSTgnUi3CXliF6ZV1b4XAMPymPfiEUg8eSJqEZELurU
T6ZPQUfQxQN+kRVcFDnJkvUvEEhDTDnafduMmvmDVPGQcMxGr0b7N27uv5w6cLInMaBX74ocnX7X
+bbvUKUdw2Wy0m2W7zUbxZHLB3CRaEWq8qRK2l3RyuzGf8TGoOqmFZST1ETEdiwxT4Vy6fSzi8kK
J9/ISxY3Nf9mRyuDgBssYT57asITX2f2QVvRzzHzE7/Sq+U7y6EC9jGgZCEIV4JlSplRIOJCJZdv
BZXNIGFsNzmePxzN6qMVLO+k3hwRMayXJXctubuDtVr7MrLgRl/eZf/Wv1sxuICQIONIk8XHzwkz
/8ztGNDxf3/A13aKqHh34YtC5nYVcXmbxJ6oouwI8lcXUCdoPldaKlhBPPOLj0PRlPMrpEtXtjL0
9wRFtnq8XuRR5LWIEm3I5hzw3/XCY6nbRlc47e3Q3csgPgw/5R1G3+5JIf8oRNJ/vltlh0fHjKtS
0gPEel6sGvgPQGVeyC5mXIPxkal2b9jViHVcABSZdHQA+akpuE9LpgCVf/IL98w8ugvGozf0RGoZ
VoAjqKK722KBnTf2MtmGh1QUOXfCX2Xy6eqU0GtdpahMKm8EIO4jqj35FUphL0QCQ2stgvY5EUof
MWOSuz0dxZ9F72Ih2VTjptIv1sBRUXsX4h2wW/O2sTxciVgKXRHNMl0fF9xk8aMhRUO9svY9nbon
VwMVSkwxOygK1nFxhXB9G1lPiGQbx7Wqi4SeQi26hdvF+jSKDtgqDZDPtosQ+AW79y/QJs9III6x
ygE0raPdE8+4qME2C3Mnx9UGNsnE5tOVZdVmDHfRNYa6RUHP3ltL2oEd/zQ/syW82rrAXjpEup9J
ZAriKLZLn6cO1Rzyl0cUc7FEV+2ptysjUknz4gX+FiRKbFBO/Cb/Xv5jVQczTP6R1wxxF3RbpZAw
yE+UdynvDsbGT7aE4b97L9fSPvMw1LC4J5A0hUEvGwBAXbMU3WyYgnrmImtfv0QsNRHYNrDH6bb0
CfqWjUm3TsvMd0otixzqeJVybvrNAdjbAYM20cVVSrisppJhHV4QTTXShJw4EjJa7IOWCuLwjiwM
MYjFre1B61OLeOOOFVC8YLvIQWgo7V4urgaGRsfQb6MeJT1pL6RGwRdSelDOCsY1i8OcP2zRfjdq
z4F2KeIpe9ivzN87Y+bwDME4WMhyM+Na6Clggb0R+YJ1/kO08bA1euFNHXoTaR0OGwfY1QxIMfQS
1wDM1KYLpfbnz5wRdhfR/M4bnvwWrvg/K6DtyU79ZgeY39amh7dTBqe+cvL56GZmug4X+fQbnfZB
1scRVSFr2v22i9IKQsUstSXwQI6CrAyt6Ins5yXZ11LEWg4iXF1+FUsd+OIqYr60z3IoEqkmJ6s5
OYVsEBlW/6RI1qrQHPPTZW3r+hzujJSxk8+gobHytr2PU+xtXuKNRRV8vNzq4aMUwMjoHgjZhzvb
NPybWXutF1gfY7X2HKLtJESOgUkwWCWY7Mf3+OFNlLq6+AupLgsLiirSsUtiPJbxfK8VsUtvzXDd
1snJVn8QW7oYB6aj7lrJ2uU9QWK+XQSQUIvXaHukUr7GB2hrGuojegIGh+Jf+ONxMWYZ3IjYcwzf
+Wgq7EEQjNROjAigY0bgfIIDP+sCAo1rwJKC62BiKSaxCnm2OypAvz6V9T0weImT6pSvwiLLOrdG
3jqlMwL6QTptepRVU/l46oylZRGlSXHxcQ/BAbGrydjcgQFpneMN22CjHFayLFJEOWAhW4Se3dDw
Ix82CCis47uwhj+ZktPWoqzfG+FfUuGbpVHq7UujJ13j5sWt30bYCUjj/XFkSfhbD+GJukZFxw4K
q/OI5tHYUmFLbTdI/1u6hFVSxBydJu9ynyj8gqkxQ6YrEqTRuyLqN/fPHGFuvlzd9qAkIWtwm8F5
5zLbSzGVh4fTfzWHsWwNp8x4iIBCnNSHH5ncYI0TZC/2oWQLwhZV/hW56p5PDQ6X7kHyXg/XWt11
3RrNthOzS2jE6o9HvK2jpAxNtwEaWNtcwK9ryfOd3PARXZ33WRai03+KTmatKW7IIOjyxuN0mxoA
9KbmNhYGk/q6WLblXz57NJqdp4QAPB5ACEI0xZXFu5gJ5rv+NSItjfVhQbyPDsfAnVM9Cb0Oym4a
hJmTNIFQ4W3t3o8F/XIDbL04+61aSvnS7cxnAZnBsR8u0a3IpxGamHHi8LeFSLbdr3WCyPxoNXlP
xn4GSvFI7fz3NpECDCwhBtngBSKOz2M3S8yNfhcvBFdaEqenxEfh2XOZnhOiDGtHxKpeONyxMiHx
d+syP58RJq03NSd1vRcVBX8GKYnAQITxNtq7nA8fhq6yiefDwYt7NNd8nLmLCt2CzUuTLppfl7Hx
6XXs1VQ2D5cMmO6LM/Q7PZZFDK+lpABV9F0fdD72zz+8fUHnERmQbI9WnA3OPsruzU4jxDzvr/+D
/zobJ/G79qTC+4xulKIyb8nGb92dfA1IfnIPRP0aeqncrZLXQocI80Ivqj3lbC0jAaQHveMNR762
P77ut25x8m8JAjrYukm33L1zMrX2Hnu8T/9CZ3oCmw55IE3wBpA7Yr77dBqUa9pMmW8ymLFGq+pr
yJb32FKmrZ8k/VaD6EOgb+DISUahz/1lz5NxloWdxEGfb07nw4mmBmqmC++yrBRiHttnm22OCiLu
n85T88izxbJNhFvhDBkp79uRvTwowMjWDiXmc+5E5lBC4KFLaVLpixLhLquL8UZ2tnknBxThEBgz
z2fIG9pc1+lGDto7LWr//sg2JaxBmoqgzHo7EJeCVlV3qnEfTQA7s1xvItxaKpxpvksBbdyFTajA
5D0JtE0rMiylfOlGVq7LWi8e4Gv8F/wMMSaOMpxWcQV7vrTf7GJEjXeUqJne71x2si1s+eOmygl8
lxjF76ghR/i09MI0pGPif0efGPhopZwWjbNAVq9fUUSpxIFJUvWiPbsZ6JaenvFDgL3zhv9NAMQP
twAvtKch5ceE+7WVp/n450c1Mt1lkw8wpYihe7vXAJqrmL9kSf2RbAnyk219CzK2UcGRWcobNLgq
mlLSZieHukR3/3u+XGHj83Kk8B9g0x819ulmiGKNAAz36iwkRLzRtRvZ1eVwLIub11kbWIUzOqf/
HtpP46ok4jkMmHu8vRB23WWQjK6utLyzYav9dojs5hLhlRrDb4xqH83pEbREoNuvjK9vybKjQlsU
yEiolMp8e3YNk32bUNw7jYXt9LqS40XGFlXVGj7N9xEjE46lVc+J7ecrMIqtuDoXW4vJNOMKO9+P
iHn2RDvPauG8qR+0r1c7nyYffNwLSPHRZGov5zM1YDVjPvmprG6nn6UQ435K9Nm1vWqe0PEeAg3Y
cQPUvpHVMang0es+E8dW4cmW5csN3bnqOOWK3V/t+eBsOvglKChrYtW4/9yTHV+z31OnSO1uKUrm
kSNGMUWUJzTIc/PFWqtjK+SWK0vZLo28rpKxvdHIMLHYT9kErQDvqpP3SSRXaYbI0zJTLlOABYvU
q/1j+Rits3UyoeIVpMhUkJyxDdZqg+rzdvDsppiaZi7TNjF8vVgwJnmByhnxbg2NTK5GFz7AQdUM
V5jOt0LWv4Cx8mcadNtNaQcAVt9W14sUvwPJWY5L3zq7RBhTFAPRDZVYxRrtMXVSjhaZ3yAAsoQ0
Mw98LnMBvX9bp/6KGiPcqi8H4tamFOZXOqdBYDd6nVlpC2VbDsdDbcS6y1po22JB34eLBcixVzLW
gnELOXDGG3vtPqlYcyB1BPnRBK6uYmP8eAs/HX9xhMmp75XaOFO5EFGHftnJ57nXzi2ZAj6LaBQ1
ckHHB+R/cw1FjtLKXH5evbVkzMo0oCNZWuHvSZGApfm4ze/woC7SGwM0KrlgmLAQqtbH4rSVgbrv
5HaxJ8XxpwIRqMGVkKDyNUApYx+lHlaXF679sCmO2tuuOBGUQFf5vluLXYbjT733PCxv8u2I7sUr
2YvRVYpm9XSzlXIfsZBc2bq5nsV+yejHzp0ax/iStyav7UOSH4T/hHT1wCPN1E9IWQ+5dzdG9anB
vN0eF2flApCjUwSBn+g8zcezxKvfJvPyESmlJwwEc3Fw7K6a8qRlKU08CTG4HcEBaqvfHiRWEDgu
7yWeE9OhtGZ/hKyNNwFI6LSb2/flBqdVaqlVjsOnoHwUM7EsrVVs7nloJpBtoP0lF2IXTHu0t2DA
li5sshA3O0j3E/+Ab7QU+cVal1K0FsUuq9KRDkI2dnMYmWwv2zRlNLqlGwnFP7kIQ9lQ3RDVK/oN
y5jU0VpM4/EA/UKOXeIFfN+KN6rNCHKrLrNVABdBHYKLebKwib1QjizPxCk4i9BAmIN5/1oOn1bL
fWmpOXnoWu1IzXHxia24DQYTbJ7cOXf3Cbo6IDuJ8raGdNot73LFaHu5TQDvIS8j2NfZsNPNsqLn
YHm1u6LjfLZgZiY6IRvIIXzSLcYzpkqQ+Wn3RLExAUva5q8W+6aNyYH7MhUi7i+PxC0COrNHI3yp
10TRYBEOSp0YJRe5Gj5QrfGqcbL2VBbW1jakKtQztFBkLXTxMim8i8IFxQDoMxicUDCXRF6Fs78A
JJ2Lado37NsVaqVX7I2GDdDxemrf2PptxeNstC4oQrQUi3fBDnnSmKkfle1/EG4XOjfgLxlsPpjY
9MP8l2Ydb7iktznzTqBcMpCz8xWgTBi1WCOzKnnViP6nnbN0giJE4ZNoIDcGYU0q8GSp18Bw/Ye6
hBApaQo6gwZIHmTN/kTQzEFUuRd8pdOkEBPlzNGawEY+Eqnjg4mXq8xrUTZHs3uU+s/kJ7VEbdYF
duNOUNv3oWcIsCAPbggwqzbfCWNW+Czh30hy18LH9DlIqfouCORK8cAhr8P1O7QmfmCsVAY5t5Cz
hJV45HpcuNTqS41br072Ym2BL1LxvM+wn7C80VQxKRP4h+tTSKO3gO9J6uyLgEH2EA+TkHaT5ot3
c/Ei/4TPypsCmpc2Kuz52Z/+R03+SFh/HovTVeHvj0vuYzGk6UzJInMECq+sFr1ReW+XUT2wsDPL
lGXzXy5Tk6EOKxt2ntR1aqq5rkQZ0hoIh9Z9SspF5Y0u2oncjsJmej7UuAxxEVlUm6GCD07qIS/e
tLqLyvOmjeUp3VbREsPb6oSJsZZG8m9pmtRc0kPge33xEaLXOjR7SBoNz27vPP0DMW5S+m+n2FpJ
Li1sMb3lNN95y5JNVYucNbAEQEOaz+stMq1a6G8nbyuGthzEYMfhVazPyOtOJ8+RzzJqOc1+IZlQ
B0wsze/111iWZ8L7GYvixyivloYEycLe2ElixXEI2Plb0k6o/ZuUkfVsEGjCDuyiooJH90NDDDMY
GkiybJIzUMlIJSU5UrX9p3M+Z0GBZogS3HXKWCKy0unaVUeb2VaH1JCdl14484vHiSxDzCf4FviH
rIohKvbIhj8Ihm3rBXUy2BIRMcj0JE0SXjmZNHV58A2/YS49kR1BVW1dcgu4Dte47DU2vQS71zvN
nNCBvm9TRFuFj4bzQft2+hsMa4KFyllb0BKYOe3KbfZ72mN0gBGuPK6PGv3eS0JFAZkChr25HPRq
2RLiQXHGcOOyDUF38r5Rf+KK+MH6JKcaP2F/+oM8k0sYdmNBBEXvxwGgqxm7fimAZyzAzLpXRKQN
APvZtBP39XrwIOH1/Dx50CVu5tl4p6SIpMsjfPhkDmi1xwVNmxNhERH2yoGhkbc8AV77So/rHEpU
LXDslsOG17xFBFHoJrTbB0TPAF08UFdRQEk0vHeuFKnsQ38b8ru7JREw2wB0/axFE54beoGwdrGG
5wbyrmBPOMbFvC7gfGowxgDefDUUcNiGKg3IweelRR+Y7enrTycAPznPWEC/JQbew6dGerRNHz24
XpX6ETE8yOydwbywTeJO5Ba4c6V8+t2J/fVBI82fh86Jm83K5AMIj7RlONj4+OlQR8tyCTyiIGYa
KgRiwcNoqVUOqn6g7ga8lxGC1iULgg0I8coCWBTbv31th8mQCqts9RqMR0JhKqAayxnB8mcL3msd
ghTZgAmVBMmRh9jidnZKx14dWdHHuRF1TbesPoiYhLyL1Mu6rhpfMZQK/5ZCEF419czk1fKTPk0S
c9aq2BBUldYj17LykiyB4rO3tqv1MsnzKB69O/O0Y09bD/Hil4oa9SbBw5F2659ZJDUdobTWIjTN
eMbNbQFNVqbXILxAqdbOya7esbGLwWIabFYgu+TUOEQDD9ze/bYg8DbG+zPxeLx+hHZdiAQYRfPP
kdGNzQ3D5Lzx1XmDigCmxNJKygUSv2maYWbZDUgdNBao4J48UqRu4DqMuDC0GHeWlUsXS9Der4dc
Z7Y+E6UlUv08CJY1CP0zcO5I+kNkCahTJqMILYcxzGgzOPQFqe0VYoG2c/XDbXgeDgPqtgNNHAQ2
3+N0a1BYaVpBsIneXcdmipIMeHCfOR//83/yGXn7nDyk/xmfpQryhJW39ft1QqjSiVGwDk9IMGnL
t9KmKXfsOq2mn1mpeCLI7TRzhV9JM8j0oOskhEDnpj+F6vTn+7ubTJJ3TKTSoL9OtIZarbXnemt6
YXtEuH47OffoaiybQXBykKmR6UaWrpHI5W3sde60njhGyVPeXop8sQHgk09dvyigFE8yTRUrH986
28zsD+1tZLslsKNauKIbElpA7RUXw5U6Vm7wx7caZGno5kRn2DhUlRpntzMaDaSTD2PLH7prSilu
ZgwqREiPSFaP9WcAnDqNiazNN4M/65sVA9wFyAM5ZQAe7U1Ii1DKWKwh4giYBJpJzqccLwzJ+9QU
EZSTPBQIwzLZp+AX1NOd5UK89spMIZ4ovFmhqDQ0k5q/ZMSYMGy2DIL8DXQ2Zj9/Cae5Vm820PrL
4mB9iow4hSPRAYEBy2XeMhhX/ESlOh0InBL2jUy8RxpuRxaLBMc6zYG+29ewmCMxO7cTuz18KTkX
4OQ/D8maOss/xIQBslLYLonm0tmwese6RCgCutswvAEOLQB+9/vLy1yD8JKCU6izhlAPRAfaVGH8
Fqn/KkBjvmya74XjK8Ejx69jEQnY/Ujs/geIMe8GAFQZfLsodfsI1RtJSmusaBqZ0CMMb7atqPjG
EFcPi4pvzyeIaxnIrpvoJsZ+INqgJSqxMhgj10AvH85uDP/jMDIRl5vbVVMWdtkwJHoZWOP8j9WH
kXe4M41nvqyV17fgz8UNP3PX1vcvI+OBSKskyyEWB/4fUiwHTCw0st4uGKWm6vPhFPbUNz5U6uaV
rmJM4zraxDXcaEn1TwvJJfzQyArqlwQ6sud9mKf0f6BedbJudvWGNl77PjAC0hAqGDIM26SSu7zj
ifRW6jhOuqg2utkRf+N6+u1i5BM6oRL44fCha+iaQh+ADociJtBQd8N6MI0ZzpjGr1T8r4R3Tevq
IrUbFrVouknB3CXOxZPTN5LdoAsxcacUhRTQ4ebYWJKGd/lXHDvJHWU+qyghL67dXM1aPzXgTmpA
A+JTezkfnjAeGSHikC0vpQeoNYOIhjsoKWa168otFimSB6SeFRn2hP9wdw5+o7Us1n1Y2G2WJWvs
j4YtM6952CzOBs58J4v6wccJPrW2kerk6MZDDNevfP5eqBeQYZbtU3AzAx/X4ozl1dz3PB70DKDB
UplVhFYm3Cm4ALFwuOZzLtMZTYe6pLhWgHXVYf6/cOka93PgWXjt9xfEVyKKDz8Q0d9pzMHmAMp2
ZGtXnIPv6x6L/S+hPkUPLHd/QTbXfiHQ1INCPIonkLYF/c1jOZT9KNWj2oRdwUuHJJIqnfDcbiQE
wGuNGX+j1gk0BeDw+bvdg8hHFLp7UeyHrXHRGBRip3RfTZSngHgfOvzPtfRTSTIL6PMwEttj5pu9
mia0QASuHISLXnId4Vuw+w/Cb8kUVe1Du8H3nK4wT+Dp4VC15eOtwWijxmxjSduXJphiP99iZ4uG
Cl6wrx1e4rly9fAShVkdOzZvRVD0mbUHGlT2L279ds7O7MC0nd63IQm0AKuU26VLIxlWTa5bEUs/
t2NsrcEDZCqv+3yNlVca+ZlXPBWT6JW+esWvCiHJlXSrjdOtbJoQWPX52LdDxMd+ZRlInqqjS9Ug
D2DE2DuW8blIjiq7eQdVnzEtx0cqLFc3G8CeKwBM3PFtzSAcGJMPyU2I1XKvahseHaTlf+B8JEQh
tzIYFnzApWUVvcfLmUMWY/gApz3Q2LZV8U9jtHFh4vhoi9NLqHoFKs5SijN2TJobNwW8rpS2Mcmb
Dw5xz2uC9Zf9G7mAxvBhGU+Fqm3Z+mkyxUe2Iu7RSyE1S14WvrWKVUGEMEx+GDtM5NKk7fguvl+x
MKWCoFosIFzQwRyH2iaGzecETevdGUu4h7ATPjaAiMOzKtc1lToAa6JtiN2z+v+jQJ1+pQ2nWayc
UH2/GkpApUUfnCy8hUAsHr0Sno6pq1DZ/2aGyVd9p2FU0P8qED/EQGSnJLW86dfnmfYppI8eOYkA
F39zsYcilluemtf3OWJlr5oy3//tYlRheID+81a5MMh8RgmB9CnNkWtKUt3SC8SguIH/UCtWd8/6
MXoQnrmoAzOcnRDKao/uSfTDmisRXK3NFm7c0jM1Bwov/3GtlDGTyK+9TUMsjT4mgXTOSO8UhmKA
KpoIQj/Wn/vF8+Ett55vA1F6Fs3rkVy4UC6ZwW1jpWMhTxhTWwW9lnGYeRxrzwdjbHsk6kr8VWEq
yI3E+jWX+4e0aa7JEcWaWsgM0BcEGY8U46kdxydWzJ5GSjhNsZHPrlddXoUsgJnGoxGDiBzS1FXg
WYKskjbf7nuSZVBeSB5gTZO02HAKYCyN5DZHFZkh2LNystvL+QPXhcawwgui7tEZ3bLXUhbICr8t
iOan8grKEZ7qp5F0MoGzN/A0hYbN1TzzMqNw29Z0mAZFAiLyCXIFGOd01V9mo6i07ajMpHPcQJ+H
yQ+DlwS7ENs1fbOS5YVbGJZvVqcYiSEjotn7dVgxmJPmeFEWpfS+vvNzC86/+NQY6cS5U/d1RS8n
W9LIbZ3mJLE/lByLIO1SpadhYTAcRnaS43PzMSZu/nIfiaxaeK5Zfu2DZpf+OnqexcwpNJCoj13f
yKW5KmEdhnCkPqn2WoKpCFLVwlYkeAwR1P3csATNFqrwh1tznMZJaRysGejEKD659Y/jMGtdNBlN
7eCO2jZ+5bNmHzlDIVqgXVyyiSwLli1EfnrxoMSqttaNS5s5ilJY7vgjhlSdk8+taRMju15pkCUz
aRhr+KkySN37lv3ndglHgls2VX/JVeImTJhkFCm8ZN4DyTUd7Wxb/V/1yx7uPmSICoyMbJYRYahS
NTSpMq48Ys/tVGMF7KyJNixQYI3qZpoCqYJvYPSTFj1pWZtIGVmKd8l/Nc3c5/HYh2m1CYDxjX1u
3OvYAZD9zFagoFIKFg1O5kChN6VTgNO/7UOLv5firyRHEvLNmaZN/Z91GOipQgoz0oISiyvXC4/X
WjMfr+3oha7A5xY1O0OJy/nOFLNc+/rrB4G9P+0BUUuglbSLp/wObBR/oynQT9GtCY6ZqyDjxxea
NiFNSUktIGlAoHJKgYgL5xuagMyQq2H0AqG8ii8CH7/yVO7Fzix9FpYBoiS90NroH3Ghp37FDac9
muDDi66aSUTC75iK9giETSG0unq75EM2uI6tEIU6qAgfjLnNWuKaf+WPhkbwhRClL+cY5QQJ1hy9
dUks+2eJ1RJ6HMw3Miba0y0iRyEbRUpG9f9Vn/b/ejMdpqHRhXr5sPpRMPRFAqPN5Zilk3EFd7MI
k7vPZ5DF7yGibt2nnRToDv/hJXqnNHNQfb13E2kLcSx9VKqs+hD+03Q0AWNf/706I9Gsz2bS1ef9
/QGGU8xMqBaFQ1txkMbAgqRQzlNlLQlBhEBO6lqc9wqJLeXzwj9wQVQ2HvFBBCxV+kxMjfBnpAit
BSVS3lkmwVPPeYkVDLNRG+Q7mfnsnXEYF7Q/mjsASzkVQNJvrYA+Na2vnIrFabEybfa136dqW61Z
3SMtNyGASv3QByKrkqzBUuhyO8de7SyBdwREx0/qt+RrQe0RMQN7aa/W/nbdLfP6Y5HZLiDgIunI
sXexE0pAPxVA92e+dzbRh1jVxcmTCJdtmb84EKE3EiZGT2eC5yKVsbWcCUxHsqqmkb/pWJuPAIiE
23xexhqTSh7LFhppLnqgTc3Ix1V2/GOmQfBhRZx8Ookxj5exaetYrvv82eWOB1y4r4dyn1aTN8Jn
p7pCsvPPFtQ5YdauDBRvr/lKNkfXHaIs/9tTxY5OmpTJsffnZKmK2Yz4eI+dKVIqbFcXC2a+T1cr
z9mZvAegVEYERjTdMR5WhQJuFY+kMZbpkNN7ajY4+GviZocFAVTDyfQqMMDfD8NrrxB6YqOdRSl5
FOu7oXvdtAe18qLqo9ozuqhaVw1nQe7BE11Dhh5oFBa/0Jbhi/HBMgboQoxtVzlQM11ijpW61KD+
cr3jlPkch1Bvf26BlHm8bEYwKnzJJERvdy3GssBL5SqBSDN7soVgklPK8VHZ9MPTmzwFQs6UHoLA
wS5gqziFp6RJ/3pZ0wYRJb3Ak5jpHmYEC0BYQ/i7LjMfGjWmu1QUg+EuF8UW/zE7zBlfLUEh6hCI
uBozn4GE6TWkDRsrRZocUPlTFtD/1q7sodT4nyq/8+n4sHN0K/LO+46Cg1ax3BSRlJMSuYVN2hVP
5lvjBL7QwtOlRg2GF2oa47Dt76JUuw1KHIV0q92Pkvg5PPoi2sMPrj0xejO+d8FrKaqBmJV+pxgU
InuPN9ieO5VETGZ/JTxn8KVXPEZHN3sXPhKzsOV4/U0RpBsuSrH6Uwyt4zhqk0B9H4tAEKYKWAeX
ClKQsUT9laNTxoxIYwEsj6mgr/CakzeCLlRtU52DQeGjjDZs0PXhmaijQQ3CX4V+8V1Q+uMwnCZz
LAblx+AIuakVb/SMzV0AGr6QS1rphE0tzc9rRqABk/RcKeXWrH91LTuO5udwpp52Ulovz5BsOzgJ
ymapat+7vDaiMWQupuMtkUvADTezO9efc1Swo/9oceJ+HRJaKy0dQDY+8tv9Ch/43PshL47zkDuQ
jcOYSjlqBaORolKzEnQX/ywv3v/YxODkvzt92LWd9F9qtWR9hZxAppjxg7DN4ITjWs9ZUo5dYVxD
aq59DrNwg8EsLLuFL5STodX9IKyqgP1C+a1PEHH4QIBC0qIoqQ58KKHAuQObsb2+4fZ4nklPubI8
6kW8nqYmFt99kNA8K6qhZi2o9IbBTDMNWcrmL1N2To136UsUu42Voc1yfv+0OUIam+OZczc8BRtc
xo1Hn1fkrNo3wC5SFVWfuonhN0rTwwsizpnfAP9qKlCJQ97tEn2Fj8k70OZ74LZb3HEZF2x0Q+7X
WcsLPdM20Oz25yYhFVo6Jh2WvOAJnl1t/sxh+qsb8v0yUIpTu4uFcT725tk2IoCpgdzpv204wMHf
hf7GHj9ptmCwnXZ25LhVf3LCBPIcovtrMIG8b7i21dic8WoAeI6CQS929xoz1vV8KiXlyFrz+BVA
M+7OSQ4jk03e7rYpx1t1H6AbeNXVMurHGdRqB5GA7yCAIWUfEnspSIs/Biyy0DB9exC6PSINSo0D
raxB/hGQDFW3ThOgYGpIHfLR4AkWM3JmpxIIvjiNibRJpwW7ewGGoLJRPjzoSDDE56HaMwwP0I27
OjT33dC9pgMBzBdiT6nj/dS2CvFe7iu2vYipNkkhoXvsJnkbhgIIr/s0m4GZB8bC/CTeCRc17DTQ
PW/NayABwTxlV350kmpc7Rra4ndFf9mRJfPOuj8b7QjnW0722bCzLHEbloEZCIAu3DgdZN+ZTRkg
iUSTFPrd0PoisNGOHN/Wtsp8QysXCFaGmsnPjBuyEUp6dBnfMX1RBFdT/PGhEpzkjWkCcj9wihDM
8ELA8bFGv9Oa6ZGvS8SzagwCvvNSb6Y1p8AXRyyCM6wfb18c+8ugJEV5qiWEQHvX0fJdVpAMHlK2
v1lJhAFkeJLhSZGOTn6ozyTTu/hHOiZPMqLdj/Ek8kr/im/Bazi0aV0ru8MqoGkNDTKTOueNCgPG
26AXvXj/YAzbqkyZxCJgNsxPzLbNOxXeZu4Dxv6djoUJ9MDmRunfr+V8eF0DXXRPK7fIIBgpIsfh
r+SbZoeMwESkvkARQQr8mGLEt3AC6nqDjVLhzkjFQ4YMWPKMUBiNhkUDZumxDzj3mLtyCCjv6I06
+HnBWW4smywWg9mB7udlPoX48FgQTEiKcHnWtWtshSlsympkAbvGmPQvpoBANbizqsVqGyPhv/kE
sAbAIjnc1KalUTRqa+NaJURVGzbfsNBbEPg4DvEcRZayJDayknobJazVSG3SjM+P+VOtnStATuMo
HOZfVD5L6Oq/TAPePpz7qc1+40S91re+/joicUkUFqW0lRLNVuVz6C1get9loLSoe3UWCGgfWXxf
2Vr2V55+bRE3y3DesR3i5iCUznlDIX9iNtevuxac0KMacPzUG76Nqd4Y51QIW8yDkeWTcsDgs8i4
p3ygxdAC3hmtJICDuTu1QJ0HIO6Z/37ECd3BuBWHES9DFVqx+lDOGxsnpILKGS7imfk0d+P5j1W+
Isv3xTiUSXW+vYMpWZQ4mMgz+8kXtAjt2SJKCSYMZg3A+nProaZDZXt5lWniW28G+XJwVi8dpEfg
ZPN8nd6lTe9/v4WyuWcvLzliBxZyh72Z8K+sScbhAW8o0EpFk9MOhT71C6BhZUiMr4G7768cDC8q
lTucr8OrUstrIMVQY97wGsuTWRuhYQb74OK79AOm5UUHfBlLWIMA8h5TuDSSRkqbMQ6VI8Ik4tU2
qhFEByKBlRzvPhV18Rr3VCQyJvvLhAddYjoOc61DqaukX7sllurh3OX8WoD2LIXOXnxvq6TyFXQy
HLuI4WUTXThJyY+DpjSn6hWyIcneonAXeGVzOS+OpqTMY7QA/zGE3coh1kK3CAFWcJ0/exPLRclk
saSa+6P7mfwC3opI1hawhxdPjk4M6hBID0xowW7C68jp0UiIaJYk/r1mE6hy4jgTRVBkChq5iIGF
FgAm0ENdf6XiJ6gAhHYvzmnPDK0+fZnIz0ulyWz8GY5sWT/8kO4NO6/LtB5s19g+ToPbNw08R5O2
ZAh2befSfkyK0jyfVkndQDRFLchGyV23hVwGnVAT7/UhJkInFxulOtZNe6GIgV8300L/8NFS0IyN
cnE0R71HcY5xERYHk23rs0k6zaiHHwDgPRr/T+2u0BeEb4bQWFHRALU8pidfte2HhbCOA2padfeY
AtkcpYLPu2RSogFR2E7yCkc47wAODLGPiAImhpdCSrCBeJuGg9gJRt1p7zHtNOJP/ZHHFfW7DDTn
8nnQo9EPj/33q5vPU+G8w+YuTraT5ZrFtMnMWEM6h1GYIQ7M8oyhNgW2YNlt7b405ufO6GNFIA6Y
JOkaj1hLfVebFNLQ2jeDS85Ar6EXR6vY4bHjfcZIuEU924qRMxS3EUCZFuu2lTWcInfRJhY+7zD1
uo0eE207NKrowLMStp5GFCIgnAcxldQpQu+fU/nvgSr72Mg/aP15BBiAIqzD2BtxsrPSghnVrc9S
bRW8arcoT4g7M2A7oHQO5vbhdXFKw8R3YfFLQ0hjXDA1BuaGH/ChrS3btKhitt6DaGH2GAF97lKI
lKgbvsNZY2z/6Dfm4eXMgotNzLpUrbyygSc4uiQw+TZ4qqxAgwrjsoDjXUfCFSs3ev1adCFaPK5q
a9xkL+INrnhtYyIWdhsh4vAEIWwWb+1aoFufDXZsEbK84LxjdlHDdIAR5IO4rtIu6VOnGv/wOId9
/EEjYx24OHWJgGgzRo6B8XJ9ktYnhAU6sXtIfix4PewVNGkBlXK0wIkA1rzLHmrjQ3uyAqvO0W1d
wdGAdzaE2Ay39SSbjZXf95g4aKToUOCXL91/LciDLBxFj/tJuFEXvHr8p85lSHyRe33pXgpbSf9+
Th/c6SnJC2jnFg+U+mWd5rgBDb7LN/PJxa4Rn9Xliyzpw1c3Osq5Ad9Neht3KMKdGysNUn4V32iq
5PQFhwSmQHI2Glh0WGCakscIG+/7hqsXLDKzdXDyp1FRzMS6S107jV8/CctX/XL22fFAVIPrgwNt
yoqh84D7Hu97gCyuRqhGZJw5f88NdJUGcLAHxovR8oEEb3FFdWz0euLL6ED48HQpBrCxQkYNigE5
BsQ1jyx0IBf9AfX1bzBcf5JAjghWY7zVnd1WBMTCD3Qdu4KWdGg9ZJKgmdBzGYYF7i76/XNzguFt
G1aalgC/un2gj89rQ5eZM+VzBGzwDO3gmLqYT3UIAsUE/xC6empm3bp/FXNgy4pXEAG4BD9E0Cg2
JNdE/fn5o+63PC82IG0grs2H4ICqkduZ0qEgqldv162q45np2GIiUR8Q+hpRKQHA1waS+5+EK887
JeoKEmFnsXRWM9W4MAkwxp/ZCe+hirvPndTJCl3yd5jQrHLuUB04+iCNxHnc/BQzYnIzAXCrGOkV
N+k+I43ItJ4GVvuFgKZhj4mO6xTSjHeCUrnpOQDAosGwpnmWjYrlE0ptJut1KQ+10FKPEtlQMaJs
9Trul/ub7x+DiL64zc7a71hQc8muOiJUoYS991WIa9j7WJYCThmWyqwAfgNIiM11SEo9963TqIq5
rKktPf2MaEr8CblOvsbnf32CtsJZk1cyaGqEPHhUooJMChJBvznCBokl7jeFIU2zmp5zUK81LbCr
7whSLxMe9gwXhdnM7dCzKpZSBzuIo43kCMDNHexu49LRGcvCo1WPI9AkJWvWa4Ds8eIa/bHluO/d
sUxNXVGVkfxJW03XNAqvfoaIbdPjBwnzQEyeyzbqult0SFi7Oh6PMSvAbwUcUz6HS6A5TqwXkqpf
gNR3gUz91A04GB/3AQjWoHOW5bunvO3IiIAV1rRj8W3npRe3/rgUPsi5Wyn4qGXUGutTXi/OFnHE
kUMLSnbm6HGVx36NyCkc16zV++XU0ZM0RWmFk3HE7noTeXfN1KtDB+Sd6ixIfMwy0M9U4r4nS4jO
DVi7MPB9JBkf9AHi11QPc25mFwA700P2tNmZvwAyFankDr6X5iMBmFE5fDki+yOSXP6PEEh+QBrP
OMC4mgBmtByCLZLrSeiioIHoNW+frAAZobn6gK0HRaJ23jph76+SKLtqOMIQ9ZdrRMgvmjb58rug
k56t2LQ8gVeEOOFrd7j+0VESLkdm7n6s8YaddK+553HR6hNC8w9Uj8jap5RNmo+oEJxaBJwhddZG
rTkmeTKVwll65IflWqoGfM9W+/K5pVbm0S/tt/Dz5WMl7Lfw9yS6gCrFY0bLaZd6AhUnpxrgj4fM
KAJA6lS7z3j547ZPwdWzI4eEZx7SoFxYzJmHEXnS6r9NR3Kw5+RwzuyIhNW/0wKoIkYAUa+DTQ5d
B87b+VKIdTwhX5YlxtTMXSMNnbdaGVymGmj8oFfZV3pJA2XTNp1I+ugg2Ahp8GBU14T5UnQffI5/
IK6xCoeXMnMpopyeguzMcoKIE2ZqsGbTw3PL/nf/gfNgcDlKPJ3CP4KpKfURPIgT5OgyMCPP6UbT
KM8p+nEoBTAiPnBftP6pq4+JKQXaSnmmqV2FoP2yMGWN427R6J8k7qUGMnFw4SMc8o93BWiQEDBJ
XJbwacENtahRcrQxo7BzQ8/EhSbt4ZpTEJLC+lRhmhFPYpAl7JpBt3qL9M/MrGyurOoQ88q5W9pu
VkjSBKAUNlg+sI89UcHscCFHFynCwPx+lkJBk9EsKcFktJi2oYaGiblrz/TUajmgS+m4ckFFu2Qs
JUtfIZQybIqgIGhqQL/bc8y11+YxpL28wZo9yq3A3mofPPIpm8Olt07fx9UvD7RFK1EwY/fO/eOL
MwkXkdYjJKj1DO+O+vCauDo1RYk4wCgMuyyQYOSIpsfVAplLUod9iyqeXScjJ21/N+joh3pvuE3J
69+7shGyoxUQOj0fgz+JxS7VfjHOHehSx4q6Tp72K5I+W5I/FxR7bBDp+pfME/ede3SpwbqUkj1p
4sbrVieaHa2i3HLPy9TULs126ELk2Py0b8md03qy/eSa+wNqWr3+7Mq8xW+B0nKbEmeojXIGF1FT
0LpLgr8bUYNgBM/RWv/qblAodZXY5V+1s14o+PFP0ixL8gcd4n9rua5q6DdNk5QI0XAj2sXj6yPd
ZYXSTAqT6ODrkOsbctEYRQMVEbej0kF5Hq4Kr5LbeRYxhGMHBg67tDQgfgLpmCWtQXJVd4MyQZGz
2w0Ka+uIoSzLaUCDXZ9rscgH8WoFX50iwSguppfZcObrQKI4/BYlMNZAuMoQQv7xtq8xulMBXExA
S+kpNwP1oLuPsY/xScGAv4VviTkKPyvA0J0kTwesELopDnDbZbiabhl9snXx4iiEw9Z2tx9hATTv
1BVRayUw5/kaAEaz2/iXkI8burzQeYMBAXZaz+1nVmB+WCgGyCpYCAPYijxjSZgWQ/V3issymiGT
I+7ESa/1+8ZjiX8UHJ7JBhrFBaoZYJQ8GRnYhZPpizrwv+Z3W7YQwlA+w8G30R7AkhHQbKAHrl6F
8s2UT18nu5X7d+ALZyao1hrrKpPCdSVw60mTEAvA2LU4XBdTtfF414L4O0KBVz/lqIGk4tavIIEg
p/JyT3jqzadTSQ6br5JWBEIv9/Hq/qOf5GKtVnOqw4oq+wuMGz849+SlXB0oLPxSmA+3knop7FOx
6yKE72DkEYfhzs8XHfJEt48du7WIKBGc35t5WEQn33/wgCo2iV9KTkxVizG4gNx6R/WUbkbCB+bL
m+9YLzFjWDtOJ5SnE2qSbRaqtE4Kk8VAHrR1UE1iufoFXjCmV8JRos7TPvAm5dbe8ZOmOEdTylnd
tgl5xiK3aq+3crzt1QsuEkVqo66Dsxv6EL84OXbX9cGFS0X7Kofl+N8gzbpfjUjN/ACpQ5BzkP2K
RzES9MWfsC3TLWP8w+k4sb1iA9f758URua0HDYulNwk5VfsknxflLaYSw9cQRXNGKSjy2Cye/xe/
9axCT75+JKg7wXW5mDRR/u5nCVX7mzejH4fqz+pVeDecs89TFNmx11ex5czFAAr6BSksxoMzAANx
HAvHQeZIpAAB+QBxVSNMvNQp8nq+9wx7Bp9YXjrR07bK9EY27OWLL36umsIsWCNPBd/D0iWdwnqZ
oSAf3y6ScMuHvRhfcGsiDcgfYcUMW/H45nmGlwpDkujPR2QYcRY7wFxl5eMsmpJ6hJlyrI9tbbtQ
mLdKkuQAouonpS9mHEyNzuc4+FgAbB3YuaVZyeiBssa9Z6FuvgVDtsblYZFvB89my7iJkA3Ng258
khWj8qU3fLyNozWD9DXZlEfiOvMpjs69KknCCRsby1dQkgNqbWjmhud2V7IWO44IzB5VOV0DNfEw
3pFOdgmdgBv0Lx6kEE/Tmhd4GBPSt0JtmRcJuFxBHA2geS3VRjyHsqhEv/N9WUmF+VDx37z6fzwM
GxubKGTupNn/AjCo9483cganog4Rms6fYlR+BNwZGe4rr4vQZQLkdWVmteSgN+Mc0qJwyJm7Nc2f
QLE2KfNcmKhvhNDHFOPyRLw/zFEhWjPQdLyjFzevLTC2hMt8tFDzCs19aS0CFFjXlKlP2qVe9x9D
Jrj1slG/qPFIx3NMUgJ/0HnF6vbuibh+t+x4SfyW6/RAvb71ZrXapeyUK1hw/yBeluMZvABOmcqJ
otrDgSG51thjEG5u/29G7Vk+raw2YmyZZp1JYxiLxzcKIl4B04hQKh4+EO7P6ByLXAK0KWu1CyCL
5/G2xL+eBCSWpdJFq+o4irkRU5qkHowdgU/F4gp0x9M9YrIaLJx4yDUpH+QdDY9z01V1Sr61+/L8
ffPYwfGwVjuaC+YpRxWvse7MDbx/6bbGjxunXA4QISaVi16u9JKW2wTWUXzzx9ylS0lmDk8DhZYh
QLojARak1jbocuVfD+hmFreY7sq2EZIWyF7+QeNugX8ptGloBXE0VwaisRNCxDf5xaADaemtHBv+
p5clg5GwWqqB7aJa6rHRdJT0Gbaif2YpyVtfrw3FeQXYM+vCnPfNIh+weZjXzkq7MzvYV3LTIVU5
0keiq8z2eDIhtyc3u1VcQLBvbScUIAV4E0OpSk3MHFsUNeLZ69PLW1jRzuMlAGA5R1LFl+EbVtrB
292lNKH3ddFg7QkvqbMl3IpWJPGgCLFY88f9QGGwUhYNso5IdAYqC6N8Grh4WuzUVtrsUwuIGyX5
XVO5FhqVpuLXwAHTzaJyj4Nq0TvEMdm8pClwZ1GYiDmUKemMGqO4z3pHP0l2Nbt/bDPO/4cd+iQ3
c4z/tumD3efFivAWC/eaVrPlVXaEzuP7BUkF0+mq/IFiJvzQRnPEN0Vhh7qYXOvZXEVBASFzKdZ7
2fL28EPOYBnVsMfPuKBw6DZg9bz95q7UGbb2f/QRIU4o5KHj+k2VFVLn9fPFWP4wI/xdGciQO9LM
Td7L3LYbHT4403++/8jwiN/nVB1Rnkc2SJGGXawbb9gxQVDlAyy3lQ+vdOWJyGgvLzWSKem7HR2U
hSx0q8j07nY2+7OTFXM5tUQZ60KbleezVj7zAKBxpjTzReFb9uSiUdcNzpYY/M4ImQe4pkZZJ+PO
xuWwwKgJZoO9uxBbvxL34d4QX9TidUnlSdEkDpT3wsS5dbCUfhTzJK9uEXsEdTxqtuM2GxDVrEV8
SqdRN26ihY2gZ0jrSE+ZIw2HC3JVfnur8jHMp8D+gnlnFhgle383+tYsOgrbSDpg9LRwJSN634cv
0s9SOfWWnTskI1hSebEMrzhySe7GByCJBZFBrAVDZvEE2FEpXQCPJyaHFD4/8Gk4O7/VKkYnJNua
TuC3a++CBTtQIph/+KeUGUnfmfVfcexsI+hLHO6X3TrCU3Z9Jmng1dGt5FLnrpr9QW0r0cP+9yuA
Xoo0IuZ1tKyCpc2WYkKHVL2+Hl69KSzzK3PDodTsRgXwo+OijX3+2z1jTqs3auZw47g2/LxeOYHJ
fdP/++3iabsq9GMTxUkVHP4cqBFvL/uTjnF3TvggYVzzDGXC/jPh+Mab6o+RFBNjrXaThA1DmZwj
rWLvDIdVHOHCR5XVRd2e6GApCJ1b6d4+exu88Oj3ohwspQHqTOPA0G82A1ZY8A/99Y0bjjE+wPqM
FF3fki18APpgUg8sBFb9Y+clcrgAJzimtfHDpTDk+vFACFiCFzb9/bYz0RpxMVZoksAdilOf/Ht9
BIsqIKbFSTIz2KVTXI1IVhINXC2/mO6HZnujuunHfYIj1FfrrLN/o9Tcsu3QdVNkYVhHC9+aIXGd
VJRbQ1/IYFhbXHBEp+mvvfJub9EMCdOe5hnWrHuAEMqp7eBlw9nQr6E2d/nTZRfDrUseE2vsKuKT
psnVm15e/HlkSWQGzJ5kW6sK58GZyefuiWxttPPupwV4PPqFjzp5khfSOt2MZZ75c/AD2IVeRWso
KCCmrmUH9yewhayyQxxehXVG+Lewuwkd8wFdEFmgxxShNIbzI27xRJMbwWVMrCP/Cfc0sYh9R3tc
vsnYdfGjrT/L+CXMLHAN1FdSgTeKrHMmYARHa/eZVhZKmaiPc80VO+rlU9YpEIuNT9zJT3UOl2An
+ZD3XkgAsK+Gvkmh4BRAKjRtlL5/qBz9m6hLict6qLZtAZ2PSVYEzc9yNfE0HCvxP2nTHVu+iTy2
fzVj0ksnho5/YQyTzhC27GvtLep7MRYKVPD0F5u7wcHB2BW273JGw1eGPcIhKUo6Qq39iJ1ZkJPH
yAjTftO/VzeBHBt0z2hrdqoQVwJ1wOATCzQGl22W1pEKqTXobT8svjYA0n2wcVPMM2ngRZe3BoBJ
48bKFGncvL9PjlmmgKcFOZrXxV37WsD64kx+cnDa22Cd/KphDLwMWybcAO8oe3nsgcWpKOs876Lh
e5CfLg2WEaRiq7T9fduzBA87YqkVjkRsMNFr5lDWBCZnODgePjiQyXfY53ODX+Ax5r+IFi4V8tho
pCAvA5QPlVcsYi6uis4qRdQgFmmyu3GuFU3U7uiqUxMOuyhCy+cejj3nKkPAfr740yijEwzX2TBj
H4PdQZUrqj68wuM6LeJ1gEAj0MTCQidh3kY54CzxC/eXJENgN0cmMRoAuUvFAgPBg+zzQeCowoBh
dRryw4bUMkHuNUUS5wpLws56GwetZ0Ogd4EhJas7p92xBjEZQbrZISFOpL8qTDbnZoDK9wAN5q9q
cmGqAWIXHcXV0N8gnARsKkhlxMsSESWb9AO0aM7X/BvFZti9JiV0JWiPeCp6TdtuGxkbdcETmis5
54NKJJrtVDI+7PGd58KzmniRhp0od3FnMBTBaDtuQ84UacxW8iOVOxNs7egRJSnCO56TsWszUDH5
IbAEvLiBv25htYz8Dw3NQYLAMNUZ61ZbKDV7LgKH11U+cshdSWAh8yDF8BrRBkYSh0T8x8IYOHhw
kp6R/UoZ7XdLYauxxfa9l9JMzV3LMKWl5mwcfaaGX+huJyQaFaA6LH8/PzNxU113H/LlRF12XYVF
5Q1r5gHxBMVi4DcNyUEa+uLWhge0oigMKONFu09+VeJgaGwNFsnzoX6HkFJzQvmQlP84TRPTB0fD
AraifQAARIWASKi2gbCG1FZU70T0JTnc1esBfyuF3xGKV7VNPwPlCFIFsKPTfTfT3rkFrhDcjmjq
aH2QY5uHQj3Qx7gfF5ZTB4mFXZAok0XF0T2gOvTnEZKxhV9FC5icwYbISfxBIGclTO16V7tvAJNw
FHwAzaz67ypcNIFzojMcY/zqeYS5bIQWxLcfVMk5RNV91dNXY6FUC+s/maQ+aTSzXOHHS8/9DMK5
v7kAiSDhsEpkrojlnQMqhSBdI26IlrZV993lr5swAQclr1bxM06QFJ30/faF8mDtDRL5PzlbC2X1
xnvTaWml1urRVxvxzg24fX7APSPTNrRAngaeR2fSq4+Sw1o4/B8McmqcQUmRCe7qJTWce6Xl10m+
Nqtpa2u1kDYJa6Ll8XkYNTkHCIt3IU6scujEG+qDSaI7txGsuJXfASEnPT2hJEEJJ4WU+mqN5Oub
DMxLZLwFmxG3e2EjEI0mPFBBV9HcpzrvkeM/AuRaJHc1OUEn6e5mP2Z2FGID8z9vi3HQiufUDrdu
/LrrDKJqHxEScAkbMnynhuLEVPVwWiWzygHyavtyQVXa8C4hDY3AsQu25OMHakc3oKWpBPSux7VH
bUWvgeNVQemI17JLItd7Cn42dunkCUg0gKdWpJbCIA3JdZJi9K2H+2h70QNkSONNuQaxjQTZdVtA
uLX9pfMVtHx0Dn4EyEmoVEpJNYBs2WclrOyX8ii/JMWarBxy7lj0TbY1XJW6vGC1YN6Y8arjgBqZ
tUltBtXnw7XluvRyuoqsETwZZdAPr27TOe3cuodvEjykWEZ9Lr89hNYfxkuPqfwyYshJ501eIw5L
RVzrKEWCZUmz2ioGvLpDIgJg/PrTG3Jl2U8IfWxKjWV9L1xMhvsNFsCTYEvwuyXUbGTdexAkR3QY
7wfqgnZS4VE9qsaUmMjJOKAqPsiKkRvayHjnLRPVXBPurLDq291mGlXT1x8hUCdwk1U9l/lCdOsT
U2EcOYxjyOA6CjgYPSEqz3Lx3U7IlymyA/1tb9tIrF7Zxyq58uH4H8Q5xpssRyVIbeAxE99XAUwW
Zq9UO2ao1547STzuIfXM1XuUpqmYy792gftPeRahCojh+VyvvGi1mMetihyWTSoaY0ei5+iUldXw
/Ff1TfTIN/jdmpnts5ha5MyyrqX6q/gjYWrjBwXu7CQfCAX3lRJV3hqzaYcdRVGVvWI2ttpQFlFf
MWfcjsPt3kArX9Uc+tEKZM65P5isU1Se+nVIve9ZhhinDncFzWph/YVqJSyKeYJuCmBoZ/FKq0uK
rR4O3xCjqHGFEhpwel9OaS7tBGCCsCgLijxzcXClg5OUrn42CgcvLeG2jFc/rBltJI1/GaCqpIKH
VLxKWpYlc7+bISDptTxFZVGOBK1n2222y9oNPDJhc+PGJp0J/CEQIhsONOYgmotANnr4B4CJYyfo
GtV0hKLoxOild2bX3gK1ptWPTYR7j1tlI156tRSJTW0RMuTg+i3/17KD6dKCk+j+O6es2Wej/Z2K
PhcX0DNvr3YyFIuyaZPb544KxFIzqmCT8NnpNC/iLMmC2r5Yjczlu8JapfeHM1N4HrzAQjn4KwFD
2Dx4NTHGQU/y25DzmT3POwkOtyNLSb3A1niiLnvJt/2PM1jD7X675kCEdv16EVgzMpqrExcywjCf
hWuH5KXZJIWJCGr1bzN0C+0O6KtOXgn2PzkTp36+HWHASrzojJEgq9m6fqUvR/so8WLMTXIvAjxy
ry6XXlKWUt2t+pvvf8W+7Xvdd01opxELWSyQnX0SFAkGyqbdgDgGVO+wCQ/U0Cryz9G+ibKZoF7U
oZpk3etvmoNeiiMoZiDwQ9SSDQcGtrDhUnz89+TYFUw3T9innoaiwJZFxAHn
`protect end_protected
