��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���w��Œ󓔼�sA�e���atC���1��Z+H ����|�O	�@R���usE�n�u�ѩ�c)��>r�ID�2't���(h
�S��ɿ�T&���Du<����X�(l�L�b��穕]��ǹ��	���Z�tf�eסN�"����ڛ�3="5����[�oE�id]�A�)��*�Y�Hg[#\~��^����B\b�?v�7|8{A,�{}ͤV��m���"Q� "�w&+F���7����YȨ-s���~RŤ���4buH��D���ve��B��U��?�C�>�0����^�6��=����F7���K�lx~D���a���"�̪��{r5[|�K�(�V{��@6O���)�\3��AO\����d�Ys,�q�� ����Uc�B��%�R�B½��&��O��g�ƃ)��������ċ?ϣ������f�>��5����*@�S���>{��9�-����ˬ�9���3�����/�Z��?ꓭ����#5�y���q_Э�w�����Tz�O��!��Jgml~�jN/��n���w��z��ࡦ��6��h4r�2w5���3���kIi�ek�$�]�nY9��U;�L�"(P����N0���a�2NR��)j�Ц�ͺ��':
��2�����߭�d���)0�y�`������o����
�L����7ll~�Yl�}�4x�'Gm��{�51�~����(=O%�07D>n.����-r��86���`,:G�F|}I��-9��<�CT�?�>��%���3i���!EZ-f��?�?^��78�P�gHZ��	�yPg
�P����`������#'�W7QGg>d�P/��V�.|���FX����#g��Wk��k��de��4}Lu�P�15|�A8�\I����X@@>�a���;Ȏ�&MS��G��{�Ae��P��܅-����#��(WZ����6�)��Y}	P2r������
V�d�/�V(�0%�.z�-GH=|D�F/���/z�V>����^�h��k +)"lp\7r����7�*��U��:�S�A���=��j��"�vwhO��&�bF�5���q���_#�	";�����/�ج9I�b'm���K��s�&UmɍW����<,��7[��X[��<ѣm����m��\)��j`k>�@����R�0WH�d|�#��D��Ry&��i�F��L��U�-�oaj�<cg�]�F�/���2����f�M%?vr��9C�7�%W�1�^U(�����I�-�4+�֮��V�ٗ@��XY���K�!:����Q������"��/`���o󣈽"_#��E=�8��r���ǡ�nx\���9��y6UpN��ג�>F��*Ľ�U�m�Q��_wq6��s�7g ��)v�d�T��ߥ�W��D*���*����Mu)�z�3��r�NnBd5AI�,��j���ˁ���+D�W#؍�����4�v�_�`���S�y��焮P+�y�U���P,J�7Qܼ��!�q�2 b��,�`�҄ܮ�>