`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
IEzqR/+bOpbRQyuvzU3bmLkHu4flbmWDhphUB21xsKPeNxoPE+QV/f7FqDcwaDrZHm08j64dnE+/
U15bZavC/kg5sGChZ5h9H7AKBt+9Xkx3vGBiaGpLnjorkRFlJWXYB/vrjl0dgI71XPJQgo1nmkeu
HL8seC2RydEt3ATvmmBi38XcJvLUuqdevzFlQ6Z3au6DzXRK6i2b4QpyL/oVMM9/T/nZkpsXMb9O
p3Oyj3qqb3GEDOBrexj2XWR2hS9A3XbRaZCDjZauCFBY5Ae1N9f72ZAb/AGEQKuXiImNopvgtMlh
5pR+R3YHDtYi5BiKz58d/Z3n4B7IIuOcQVAsmw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="zrZqUC1zlEGxlBhbBM9aY1EqtFsVcyKPaGuGMxi3cFs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3600)
`protect data_block
oCxbrclmCQO1xEqB+gkye4i8tPFNQZfeuwKbLmyoRw0Uet6pZq9Ge8vTGdZxJjma0lbmSjaVIYYm
ISc3bOfZfVhXuebouSedQ508RwBHABbco5prKQP3Dn98UmVX+a9CMZV4gku8pkiUYQgIxd97r0gY
9Iwe2roOFkreqtWY2rToMBfWMY9+h6sa3pTAEe1wWbhQ+1MVcjIE769g2cPbLCHIHwV/JiQK25d5
m/e3xcMIzBAFhNuIcMjOw8L9o7tww1ngoOlf2bwtxBXvNF9/adD59vm+3rXAtlkLj7/AU/3btDnu
jEqGFGi5s7zdfKdHuHt+NJmMyyXS7tQaWbYFmNdfJyi1VSik3C0QtDaNn4vJ25m+j4yL5NoWxivn
IBDKWO779veA5HGRmM89TZH1jC3yd7euw/cx1uQ80dxLrASzFpTe+jIx5pwLbuzb/P+axiXjlDvH
LFxP3pahfKbhfJdX3ywzIX6ekgWwoGuQS/W2vM2S2h6TUTaV4lZ2nyqW4Fv50WtrkWW0tHPQivPe
i8z6slB+wEhTqyJHqK5O3/N/c4IlVLpYDyFL4t8WLZwIKNSluuRY7GiFjGCljgHI4OCNSucy2A1N
xm3CKn9BaPPt/lINqdbGKjwGPoA9r2VVmkG+KRkCFC78vP7m9WCD8Dn8iIOzN08jjJ+115aHw1Ra
USkx10DXgj3hVJT4YCRgQuDxvX2NXoVJrBk0wfSjQ27XQ+HSsDHuzXyDDwxE7Fr9KbGu9Ix4QzSn
cnQmZe9RwHA31P7u2uHHLytB+euX0UhpmUo9vOH09pJHedgz/LsI38M+WAebb0AICOVUdC/Ib4dh
/dolnce3RQmKXavfn1VS5NvgQTjkzQ6IajNCRF7NOYkZPBPJ7Gn6As+FsFiWw7fFo/lhggUdWIY0
O3QJhToruOfRU+pEjAcFwrvuCO2ya0sAz3AIkGVSZtbwnn4xy/TON/NLrwW4s+3K3E/VAcRyXCGT
5FhtvolIk2WLa2ztZLtAIa9kZelggSsrkgWE4GwvyKtWuI+wLz/SUPUvMThFl9d1ZSsWH3qkI1gO
jKODAJpzFW0mvIzTYRWmRSoj8wks9TNtLPaKO6xmwpFzTaFC/8oIu10QD6ChlsLLsQafqi1U8wkp
VPQQrj5U775rpwmVdrUh/qbhFOtqPPxkPrNdxZ2ZYE+POMqacaDuIzYdXFdT3RqWpZ+KBxPVgCZo
vxpPDtfXE63seTqlM9HoKLywdnuVdrPwQCz76HuD/BUtjYwkeZTXnkeeatA+pqCTL+Wnq9n/mVV6
eMgh9HGhbmPMBTgIQC0zhWqgPM/qeo2kEoBBRzla6+hgWO49tH4wM6Y9dNQ0LoZ/2v84tuZDufSc
sty5mfxYDqi9Nln3egwCYUL8tGudcZ7mFpr3EtN5u9yml5qcAkhY5Jc7N5cCG/b4969rVu02wiXC
i6Wv67HAv0wFvHcHUnifJQbAiKvBgzHzjxshtEERsYbfrN3oceOXCW0MoAFLejfzQcYCBrZSb+Ui
GDxXTkTwWDyhrNYwQuQsw4iZJnIHLa4zE2zXWqi4uepa6+KI8myq1Yb/1I64AYFT++yKg0//VIf9
zYZytCOkRWTvbLekq8xg0ot2esd8+5MrGqZoMQZvim0XNRdQnpoSYS7VIOzR/xYDPrbMiNFzR7sz
oqRZo7Iwqarq2qGXfbp2rc/BG7SnzPz+QKJ49cXvQH+MU3rnwkupYO86VvZ8+JujqDI5BpxN0mos
GsqBbEYowZ6F3xBjQiithB0Fa9xMQrvOL+QsIYxzji9nTVAozSPtyHWyE4Px/2vSGVDHPVkX1jbq
c60jJgofU7R9GwA0YYKRmu6vFdSfqEpYYoFywVFK0y8ey/m83SYCXhHGTpFVsJv+2KQiLFW3ykFL
IqAz9LdGqrQQriRhcvGH6kZnFzz7zZ61emt9lerhanhyffzl7ZZE0FfkAt1NULCilV9juJw9FVkY
Vwcp/1u3LHzVzq1MnxFUS6u8QwhxUiVwxzfJKI+6Qp8qaG0A5Vv/zNYOCp0tNVc13gUo+BDSOGEf
yDqQgYi3/dySranQxiAUknQ30H1Dx246of4bdpVzTOCHyL+bnKeQib+90FS4QZ6o6kTKWJkrcc+j
3yvFbC02x+SK8S6SiT6iO3uD0KOLqXfvgnfsbccI2EE8VTjxtHkKLyfOIjz3eDKzBJcjluU4v217
S5UMVaSrrH0Mwfzz1Ce2F3QHPJ7Dnw5OnH61CzRazSh17kGnDKINLln4a+tX0enbnP6e2Q7P2HWT
M4ttO8QZRPjJo28f4HYdUJlY18wFW0T6UZMK3Zf0mwP57XjkHr0ABjnn58/iVSK3uicSd4dYqViM
JTpo05GbKDMqnVhVy6QPbfIeyVteBOW+Sr/Cl26KFvCaeHFVo4Ic1yGsUsUhg7ogbnQpOHZKTGk+
aRrW/q0uZz88GBm2+GIQo7P0HMR2Ul4OOQsHlkX3Zm0h06vg5ol/k0CJl4rxxS5Vfj75MhV10GkW
65TK/Je6pWBLLcDsUIwXZiUHZTlcnCfylfSKOlSUKYgBdTBJPZrJrB8K5Ou/xEjZFbfaCOCUQkMr
86ifdDUERBncFSXtaf+QqPp9556dUrrYENj5D1hN18E06VWTPlWpjMMRuwOqIWrVfq13BoHp9hgn
QqKQn/xE86/wmpmSFOopC4BtjcIHIqPXfYZxsy0rY1U+33XHb39ugkUllIXV1pkF/BvOW5iWCsxI
1//yXlpFML1cArkU2HghCtYPPGCq8Svgoc+2At6qCeR1a5n2rGMeedscuu79q4ST2uA6pf1voTKc
8aTr21qHr2OGKBy54KoGsLPhIDmflp++09ZA/hACVdIwA9QAMswZag7I5OXwD9GI8VShIuGh/wQi
bC0qkgDTRxJCAm1CqdCfPoehmSZfxuzQSWbv+yd+AYAGQMIHuyKdamY0j8XvZTPaHWPXBuUbIhvN
cDZsdpzK07MJsc5qRfOvSfMd6RdAGUscyuYRaeuHGmx2aOnCJbTKR+ioMvJeMGkhGOtXqt57wxN0
Gf7X9RVPSlgca+SOsGMeKAhyOcO2aK0J4QSh9JCFS04hl3eZhcFnLRQfyRDH5ctArM1azW73OBC1
kplhVin/DUIocHBDpuYwKG7IGJ6YAZ0BGbihXuLSqEyp44A8Hc1sh12+X58TXLxLlYhliC6DQVrg
hcHDg5HJgc13qvKBiwDrXOe2XgC80iZLo5gL9jfuxT09468bJOjgRP50tCtwAlQyhikIWcZFn1tq
Mu3NDGDgXxqtQuw/rmqrhNN3UuLASrJ06sbLcsvcuGmRW+uJ1z87meox8Yy+OWNlYy6h8p108182
PyyGlo/E+scL6mSwlo6bwKIzAcCfM3IE/5ExrJsIx44sV18mbzBAxhOeiicEWT74XMTB9o3r6EsG
rabUI8Ag3gVSGZjEyiNrL6rIHltGtbRomnmTSV5TugbPBbrMWVeuup4RWXmrH1yG01irdkEecD+t
+7/Rj9AbBFe7Uvbhx2kEDE/cewr306F5fMZ8VYXtMtzz0F3mFajXHouJwWW7bCIakK4NlDsX9Wmf
YbEqAMWq5zl0uLtFPnVVls9Lz8yLQRR/PW3pS/1l6yCZCXz8OJvmG1n7M3bN2ouUPcVruRwaGcil
edCytrSCcLdIpTkzjb0lIR6WeLBhjf9Y30nBr+3obB9XCUsWql/sz867pTuA19tKs6sHonlNmqwK
on1bOGuzwwNpZj1oO+py4GF+r6idrDOiF4BSC+rF7kMAQMnGpsPZYTLUSX9LamWFCggK6MRum91b
1HE9Akl3fhPw677nXP/HWKhwwZPO8uJOvh3U+9aPumCY4cPxP1h/30EtQ0lvACv5f8d82ktFG22Z
tIXkM8zFUvSCKowHF8AkZAm90BA6pXGTljPX/najrXUyTDJo4hxgseAodubpUacHZvVMZrvMD34B
AvNupuZYOn+QZybtGcW3tdbW+M01glvuS8svz0LHd+UqzweOzk3PMRBpVctfXHlw2RkD9UXUqkw9
xnNNwSeryHTnhaqqBCoOTRlScsj2oOtZsdNww2zRZoXJsmEZ32bVQHGS8IczzrhvC1J1o7SU2HSY
8eBMF/7xI5lU0sPMbwV8MdAD5qXqczK0Iqp4+PD81WdVgbryOKpzU+ERON9R2SQ8ba4OzDtSbTZ5
4xKSjwjx4dp2/g6Tk9tUyQ5GrK63sxT63eUydlqx5m57wJOVS7j9ZTb34LcQACgmFrtPKDza+7jP
WNcKw0tPCDmGooceBHl6oncFuWCBn8ZCcudGUfI66wEewayFnj1sv5wYSIyZGsGwaoV8/G/37A/C
9c2DK2dmkg5Yy21/fUvOmLsd5I5/Bu8Rbgrj3uC7MaX3AwlOeRipmZGUAJvC7cmAnGDM3Y1ZYN8A
vAx3DbWIIybCFHXWb+PT1t4RKfFsXGDQ2stpHHIJj4MWWNakWbOh9jRm/pE2WpX01Tp4yPzKkrtp
pKDvjepQp8pxlUmBK5J/h+SCi4g8gNCTq42sqJqPGeHebYQISoUUj3A9XCgPezLqiSUARAOrShtp
7Djq/Z7bURPg6m/HyHd4rxwslndLIMVVXoV3Mggql1vgICDhnKxtayOog7uXbVhO0r3TiTlNoI7j
PdCEr4KLH+zhecKrrWrgTB8qAp/nx/aFW9ZA+NeD0W1zEQRehqaLA66x4gcyKbvopxHa234+1D9C
9u2eloiKsypo01wE8LN3R13MTf2CYAfiZ0MdNiXXr6A55MZBGJyauRVKS7bl0vsH4AirTBFd9ldt
ZvSKRaVOhe2T
`protect end_protected
