XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S��X�$Y-�����4ߥ���X����2�LT�Y�ĂOr�DkՌ�~�鬹똞\H�d��Dz�B2���!-�0�ݥuN8�k�>RU?�韤��慶�W(��}�[�����B>�H��l��s5ŹN;wyj�6� ��^7���;���q��AIT)�w����7~)-C'��'��>0!7�s��u<�k��a	KN�J��E�� **���N6�,�%�?|�"���Z%F��S�V����w|�X��nY�=��,oQ���	^ձ�D!}��+��2l���l$yy������V&��/lӣ}��;W��  #%��S����G ��H|c�r ��RT��ۤ +$���@�7\����尺tity�'Z@�&�lj���ھV�B{J��PHd�/��;��R���9�J}�S�@\kR��o���Wդ�Jn0�-�E �gup�`���>4��J#�3s���c\-A3?bmW���e�d�}�`�x��1]�]�`jrhO�D8�R�Z`�rc��� �\)�ۅ�(�Ը����5��@[Z��L�� ��iО{W��}lTY����;�I�kA'%�c���vKi�C?�?y#Opg�we)t��Z��b{��q�}�R�p���Y�l���� ކ�8kP/���!�[v�!ƪ����3�� ��b�"
0�QK�5[�M�j��!J����BeJ���VRq��G綿lU� c;�pgl��i	[c�(y���V����t�7�5��K��oXlxVHYEB     400     1c0^ͥ�t�t+1WB���a��G}?�/0���/�+܀Ў˩3c��,{��O>n�%�e�PE������&\�:�C"���H���M�|�wV�M.�ǃ���5�3���\bq �40�pSj�ns���Wtา:!�2����Э����JA��ް,�0y7���<y �%�Y9q�ь�Z���6ۘ�$�`����������(5(�2���9��c���X�ۢO?�{e2r9N�+�2��p��a4��_+֖7�O��p�O�m��>�}NM��1�cl�|�r�
㧐"�4Hs;D�:�Xe&ۑ9�x�ff�i���X�S�iQnr�r[�!K�`��<�E{��^4����w����ZP��wQ���
��������l=1�deڐ�
 ��?����٥L@w2V7忇l�t����ɝ��&Pp
��P�d`>A�n�nXlxVHYEB     400     160�b�ᑃy�߯�Vf}R���2��y�	�B2������,��4Ptgf��9� �����j������1��+ ��/�3�=W�65��d������:p�T���tG8r΢(�`KO)�%���]&9�q��YR��w���[d�r�':��6_k�?��,ܱ5Bя��@���؃J\gV9��&�ѝ�D�+^�m��/Tm7Y���V��YW.� ��i,V��N�5��I(���!��* d���R�yY�%h�@�Ia���<�3Aa8�B�;(�cϔ@=�.Xg�*���z,y����W��)�2�S���f�H����(�L�'�FD��&_��XlxVHYEB     400     160�~r�L��+߱%���щ�a�M��@�b[\}����Ώ������L�0�7��k{��u����z�vx��3�)o�	�����1����Pۙ�bG�;���~�R˞(��S��+1'a]�e�oE�\!1��$ �6z"����5���6+?~w�qUI�YxX�ӛ�U]�})��#A¤f��hY���/^3YPM��\NҤɿ#h���r'�����B�MN^a:���EQ�-	οwژ1Q�$ӡ �6K��HXO���ٵ=1r��gF�rMpӑq=����������C:틤U:�r�>�C� U
v�#��@�RլL,g�}A rU�XlxVHYEB     400     100nւ|lߗm\�U���Q�A���	��r�5���g}L���fû+�Z�����j�X�J�8~��8��2��7��S�� ���vW0E�!��{�1�u��"ס�L|SJHo�F���&ض�Ǫ.�̊��8ئ���w�eΝx��}��+EF(��[D�Lk����?���P�⨂��cNP��ܙ�Ԋ�}��^	�C��w�>����t��UW�VZ��YQ�ily��r� t�<P$	s>n�E0�ÝiGNXlxVHYEB     400     1a06�/j���u�i��Qy,�92q��0�'?�~7H�@�X�~3�jW�4��d��܏xb�(�
����flڐ��	���ׂ˄럗o<��!�Xs���8��,���� ��-M������'�>ϥ˧��J	}����5)����6I��G)Ȁ��u�����d%�~@'�X�BԄ�9���M1ia���Tq�4�d�s������֊$��
�#xp�1�������)4�Tn@w�Fm�'J�
hk[T��\������V�����6���D��M���8�He'L���D��A���4d;q�i�`��]J>�EN60J�2=��^��W�u��Cy&p}��e�=��$[ͮ��/���SB�!iGnb:0=���H��.H)��Ȟ!����.�ij��5��?�����XlxVHYEB     400     140�H��?L%�k�}��ei�`�C��@;g���_7��� Ovƍs*�f�.�X�[�)u_녺��6{��	\�	�4����d�*~1B�L�(KT������iM|P�DyG�k۳?����|�{5�R�j�Hä�C]�:_��7e�u��f��2R#��a<��u�oE-a��M�-�U�	y�KhD�
�zx�،R\$7 ��t�S�<��k]��#˕}�rs}^���Z���Աz�\�#X��'��������[H�CM߃N����߿���i:���%�f�+h-��+��<Й1.
ԠY�@XlxVHYEB     400     1203�u@Ն�T�6�/��59l�
uݤ�'a���|����͜!������׃�mڤ ~*� g�3*(u�k��.�4�^�pIL�j�&D��<��o���4ȿ�
@w��#�w��5�v�����I���ꪘ�����A�)y���x�%��7�4E�1��6�����?���%�.W�)����Ә�X�BG+�5�n�p�5n�ߥ(�xN�ȑ(�f������ �
0�.�dsYj��E��/D�ӆ���D��TkoU$/���4�Ԉ��Yީ�%��XlxVHYEB     400     1301��N<SY60�-s��tDM����=p��˛�����!�,�xQ䃃Y�b��'[�0��lf�n�:�=�,aws?�\��r���BUz"bn�y��u(EVSr��Eה��q�Ex���m��I]�HX���zu��eֳN,y��墆׭r"�
�>���B�uH~k�����3�ER\��� ;���ŋY�*9���T6�G�a���-"�,ҥ*'Tg����H�i��+C,�lW|�oM��`i���)Ǫ��|Q�j�T��M�#JR_�9Vr��a4A*q����ι����K�p���XlxVHYEB     400     1c0���pn;N�tf�.�#�
K-��ԻJ�����f��q���a��j��׶��W��U.�[����"Rs����[�5{GG��S� �㆐���}��;�n�"�
D'l�|��9�R��Е2<��@��`c��1�ͮ��	퓖����_��d��z|�����.v4 ۽�a8p0E1���'�FU�?U�E8�g��</I�K�Z��P6�n��9��]��E�h�/s�61��զq�~���p���Hg~w� d�z�ڄ�U�f%�}�ҧn�6� ��h|A�.�L�­�!N���|�~����0��O����v8>��Tԥ=�&k�KrtZbv�n~1� �"FK�?5��M��e
[w�'�lb�i�Ǩ��֯��%���C,�TL��t���R�xX����!Ӑ�S�H���q���H}3D�m��f唙�K�XlxVHYEB     400     1a0PVi�+�O��N�E1�����`�3W_�Ow^gwJ4�U����i6��u� ޼�m`�4���S�ܐn@r؁��Ӏ��w0"���E����_v pRi�܊	���� �F�j�"R�
M7G�'�?Cl��ad���
E���}�z�<3�y�ߖ-���Kw}��t�Q��{a�h�*i�>L���r�~:B�x���o�g?.��v�׏�5���ہ
�Xʱ �'�pݙ#����R���c7�KK]�;�ϲ�#(�.}I�CO���(�udWx�SM'��_znb�Ƌ��
M�~�ًy~�7��L�3�a�E�[��(�3�V�qJ?�_F0Hl�V�9珛�-������Ӌ�Zb�#�) �&��8�,.#��1_�젯��V�8�]}�1G�G������le��d�ޡ�XlxVHYEB     400     1a0� -^*�?,r��R��T�s��1�n�9H���%�g���W�s��PL����s���w1�Zu"g��Y��xY"�ڼ�u�Ѣ�����;53���u�`#PK!�鬤ջS��-\s�d�B��y�n�#�x � ���K�N=;e�����f��z���R�Ql��>{YmK4G��T��l�<O�֠�;�5v�Q��0ypގ"D2S�	m�F.t�#��{����m�_�Q5��=2Y+����w*�<'���-�`��VQ��Vz�/�����ʷ^_�+>o��s��o��fH�W?��c\RBj��5G
ݭ�KL����_�����m^�`x���̽;��J��)(��wmXGIo\�Y�O���o��V=6�
�g�g�d�?�4�����B5��ݥj��`h��f1c4�;xO�XlxVHYEB     2d9      e0� 6�}�a���Y���2c+�A��z3ax|�=]�]	n���S����)o�뻩�qd�Î�{��xual�U�¶{"�Z�T�6���ϸ��H V��Q�Z���-5���: �7��N�A^|�^;�'7�ϛ���<!����&8II9��:E�:�.h�~t�j[���(%� �����0�R=���S���5:W���~Mi��`a�?����L[�|M���2\c�