`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
sAGce/auatifVUBSRB72aCLMiNNsExuaADDAPQYUHdTcu0Qyham95KY/VyzZ546yhFcuRsXMR6b2
ePjXyz98QTGd3D+YhB9V9b1wi8NMCdLlsIWUQWHw6hr4F3T59Pr7PaXguNqLEyeg7KTbOk4N6kJA
+fVVEZrqjMwR/fLqBtPtAXX8QzqlepXBk8GDuRgcJFYwInCZrshMVwUblDjbbmy5ZAQQ4HZR3VLl
Tm/Zk6V8QDxk/YBElHe/ra2kYNxfVE2K0ZgUILAQgcpuLSU4xa3eLqw1OfmcTPb87Xast5Pe7ajz
vbPap7rpCkTxvt53WQfxoC77gz5BSEhHSji75Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="eYdAxExifUYAagPhZpIFEkG3EIwW45ycyfgp4EEzD3M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 46704)
`protect data_block
7nI/XpXwhRzg4WAK8Q6v31B7lxWK6syiJktKAjASUCEsW7HAJWVN/Ky32vvE/0mwB+K91oE+whuH
B9+1iAbW21NMmh/ceB8aCBly/1tyMpHTR//qsD/nTabViVrH3gd+IAg4PWLGFa7lhfOgwl7+Z8WZ
u44ZjSGLr2HCa1WUTpCudE0SRGXzsf5rb/eOceyjlAgrcf2b/zGoJXphSzsNKJEQP+Lu4Rhl4Apo
tPxNIUrDPex+oQlAymQdb3UVj8kJ78PvgDTBJ1amH/aGGiHwfkpc7czIiXrk7JpRH1QkcjG0wuWV
PzO+qqApOwg+01Nf4o/WDIEA9y8gRr4tNYFCnzcsqglAbC/8YS5LpASRLzKtAkcVojxlMRXwNUn0
Qy5szezv5iciK7/SsvvtWSPW/dyjHjypTI8mDXhyg/OiuNuV2SvpIByc9gdqKH8a+lm6uJ6RtWah
+zsELxGTsStbxbmKlRDQNDRBwLkRadDaAeZITcosImgE4mgC5l6EPdNPoFte7ve/czvZTPUogn8V
Rk39dnHcGsSY5XjZHhTlOQF7b3UlvTbrj853DcjZk+BiEV1EUCQTXnC9D5u/MJTMJcqv/dYtqcmJ
bpQYu2Ekh2oXXguEycPXHad1hRYUx3QB+notVhuYhWW4f3eChWs5S9eISMKA78H+oTDyU1oCYzkh
Fpq6prC2zLVdgt1NXaUMcjRXIgK8HCjkwANbSi3mRTM6cvZDlQxlP4VFocNibedX8AEYrsUoqQIA
EIKS34NqnpDxPwq/cgDX9eb3rUEBU87AWp4sX6wZ4vwJvuceXApaNmWkQtpWxLU+p6+t5L9LpOwM
t4ENx2ODdQsQ+zqW9AMdwQ8YNRaRJNFuTDn1rhbzEhD9AgrAeuK3mjWBrmSyXYeqExLxNV911Wop
Tsvgc7VbCA1s7jpn/lUdm3bmn49k+rKOkrLyYEiJAEAJMEXYBjEndXlsm+J0vltWfgnqQrgvV2S3
LN2bPHNQqqL2n6J3a6VwRSXxRwBDpS0soKQ4cAkU/7lZUE/c75whp8vIjVbtVFdCbZMpxSXpJscB
js0VJ6KFPOuskotXMe/mz8opvP3fRglJS4KMUDK4g8IVgF526axklJl6KAgdsMGVRbxCdD+ZpMTl
0vs6lFSFpjKL9/Ge5IU2LTZkMR50kM2VAF4PGY3/ktbJV5/NVDsTBjaiqllUJ2na7std/bs0MoFO
jwW6Wn4/rYGkt0Kk9vTDqhP2+AnbzwEg6txQ1aUkIT3R66PwC1gWxw3PdhvT8jZY7axt1YVVPc8u
leadj0OoBcDV6PeZIf91TE5wyIPuGBYwDCF/IPD7pjLCFeHsrCXPiOUcUpWS2bYlkpPT5M+JTvyN
1dUVqAJ2ZaC+3BYCkP24u+9ouFk/1zdSEBWxRzIMr+y+lsTcc9c/Nm+XygcExSSpV/Cy8PUOXvjN
LNfxB0YR5Npb/eck0/vxpqAQBbloJVIj9sMu2AYAzRu31zlyUoT2hAdWAH21k3bsXAmxAoCW+u2e
KiI7VQ6ptCWshS3I05La4St/XNJYEmjiabH9p3I8wQJsRneaaY0ClO+DM2NKFJkiCBtROv95HF14
jT3AqRgLg5P/OnMhxtipmgACz/+nPcssiiUF8Ca9K0TawPqDUzFT/CYIrTATHUIO6wQbk39u1SQ+
i1Y9hoCMti2oDTfqLxsocyTALgMkE/wxX078UlxcEUogagLrifLPTM0na7HDycBrFkdJeOU045dl
MbpNhlOH5W1P5AcRx16HGe76UXBBEbTsYpWmH2oRvx2Ui3A4HhXD5sKF2FOoBWg5XfVkh420FI7z
FsbqZOt8aFsioq/fKQxa2U5a0P5Jf6MDDaz5OYRXgdp1Fu54RPZhUgVVDSOp8Xa88nVdJAgbrLVo
vx7oG/K4EUlq4GM2tLuqGo6zB9e4+E9dhGQfrs5CEnkiZ5KN6iV9a/opioduwBmFlJATQNzNJgZb
D6cDRIgsFdi7F0OVeFVS+CrOoDqhoq2OCJeRfpXPuDeT3u6+ynlFvJQeJWzQJP3IgVx8nvvHg5IW
sMc7Qge1wntxnzSdqUZu0LEtOrehjgEeJW3pBwXEvMV0OD5dTjLudqtX/mKaemEhX92YZxGfrkTa
1olkJGbKbRgPRFiYXU/r+/AeJDL7pAmJ1z6JXiDC4Y041Tvd8ZukJ5AVSQnVFxWXVkoEEYmd5r5R
NxN8Ldd9IxuXij1GsdXzzkAhD1oOyYXHwOHrxrWffMw9SYpLgE1cVnKe4dcdznaKlDZXajJeEP4z
ufFKWAnOOk2Oh46WGsztJRKMpQ7Cll4XElL+tNGGeAKixkpinjj9bfrmfHB4DTLRzJr4jKKogp3b
RsU7+80fWXixz6n9xlmmdamEU66wqPW8nNvpDM/zf8mCSk+LAbDz15ibyA8Yf36r/ELkBDL4VB5R
TAUc5Gl1KWSa/232RPu1CuyaEtsQLEWTxY7B1kERAI/8t2pq1Mt0WMWhsH+gjeG3SUtvuQgcn3XW
2iph8Mv6HIscrCZdC5zzg2FCQg2yqw1frvP2NQg0W2v3YKZMMQSKIg2Z0m1wH07aoWCT/xQioXlL
m+INtaL6+e0ct666o/s/KSZh0r5f35SmD+4Dii2X7x62b18NCz3qMYGjc+Af73jrFRNxMtzqitqR
//6NyDUDMRTOUEuZtJtW+4p0rr8+igHOsDXSbEOl5R4nxkFCVNFMQKO9VEYy0HRKnsp8LUIIYlOO
2ZgPxEokkF896OhCXUm4roOmyNJI7pTSBEqKvlwq0ErfEX50hkgEnibTMm6fJ/gdBey4JOgTNX88
mIIzI3SDiyD1E5fWawrKLy/S4EktMANHsatfyNJTIN+IJ/ck/rgEwGa1yXb6RLCKnI6iKb7FFlSa
kFV87MG33p72iopHp+I2NvR2XOgDIDttoTvyG+NpGc/BdCWIsgbJYTUmKGjaWF1/JKOJNf6Ym7Pe
4fyK6T2KGiezAchT8EUMZjNPliPCZ3LrSuK4hRFktRl2fXb/39Vn3VIB0ly75EXsKpRtO9BuZeoQ
ZsjqK/Hh3/+K7cpLe9u0pozOTrWv/vO+uR58fmt8dyICwABTYShKCLPVPzb0GcvaDH2w5LCjmDsd
COfSjLbxknKc7TxbOz8NQ7/N7CS/RL3WTmpe8qN1Gy4RtSfudi3MDufePXWURt/dJlpOdQz5eXNV
kHVojX+t9YnxcwHrUnAu30hL6az0b5KeERZDJ4RpfwmdjeLDrguNZLpdYKVZNV7ACevnl0Rc3cec
w5SGaeLuNAgRN3yWDUOM/VIW1MqWMe8IlZ6n7qvA1+t8bfx38zKLVcnoIn28DO7Thd/NxI45DYDN
Yd5hINaDGps65kwAmdD+Pf23qlnlwHftCxFpNxYwySW1TOPOsdvBEmCcl2sdiMqaG6KRY+TcQaBZ
npivHXZ9EoD+0/PWhHsRAneSJT470WSWZlB+twTaxv5SYbhIXMJVs3bCd6wbyTltNeupGE97UFTB
wkG6JbewMc88YNIYspXcQQNdpMns+ssnXzAa9dsrYSqj6GDaYKNyYt6szzRpOpx/VLebBnYeulZt
7BdfDrR4tSlO6dC3+TMVo/NxtNEMoeS4HYwG+cHjOVIIE09XOcdgo6KYsIevrGy6CNfOHlYcgjEA
N2Fvn7Lmdj7yia/Kdffwn9UsZwJ17zKCr2TJa13Pa4Hu/Bdg+FnoPW+DjgZ2G3Umwczr4EkVQBdy
CUB+AuF/tqlYa6qHAFH3xOgr07aXeqe6SgZunWmKSHaN16YBnfILCXCwy98UMM+Ww3jkoGc1YM9e
92FvsQrYHtK8ySOX8TCKJ2gsU50M04UkDlyNMGhaUFQPRXqboEUT9PcNoBr4SrdT2Si3jHn7EYF5
u0zUirouXb4WjSjLUkSJfDqROKQiSW3oRFTqq0E5RwQDIqJCsqV9h8mUhBzxN+YOIw/21QcxtZMW
HITZwNSQo4/pYyl2PUxTT9SBV5r1SSGorZBA97JlyQ6glNBc/r7OOOZ32WNLGaj/NMYNLBVhndY+
+fSarKDF3dUEyHfdQ47bGB9s26l21OTXKb0IMrgDW+S5LlN0tjGv/FJDPWpJfo8KJe2Ew9J+0Cfa
Ov6e5b6uOSaCNJcOk3Zuc/MgoQuFsCzzyWm24vbUOE2H78maMXqiVGlcNLcSG3vPPiuG6CFxZbZI
UXDVRfYPYHVwbly2L/AQrNIdPJmmucX0wocnXx0oClVSQtqqQfpHkzGQjJqIV8WlpD323snyhYXO
8oMYivAEc3cmvvFEVFFpWMlSCwEe31ujk5iVdFyzmUwRTxMfg8F6DRMhfhASS0M2xEsrxA1a48q1
v/6vwPm42b+i9tsCLicZVRwlUBlboxlf1lfH9V2UaFhOQIsjdqKl6U9dC4upQ1L9C6UY23m3aiCd
aOC+IDD8GYjlKuOAWNl0Qpn0ET5h1qXjwPy+bp3gP/q4YikCRXId1WJlyfJZ8915IdpSdGzbkShm
Gzdo9jbqiteGZw6Ez2cWL4v5/eDs8nn5f685xkbrlZXKX7GPTFnDQLQnphDQEYsC7szfSu6k7JGA
X2YFfEw8ZBv+ikIGMn8GgLiJpL8YRoOuHJyMG3tXdAODfTbUkPBLDhtUs8zdn9zVGOa72ltdQLmT
iRaBLKDsCSqAgLE4FnUsUF0IfyeWmB/7BbRdVV8UW9zkKuHyS8TwyunOoYWZWSFePVS+NpEyj/Pu
kHz323PEKi0ncmBUr6t+oCAPeVJWcxl8e2elMZnBu32X1hXnB0MMj/+lLRYgYINmzYpdhmJeHU7E
OoX8aOAgzZSjN2gwa532idTlu+Vq7OmyfX8Gc0BQmCZ2oy+HmErwvZ+nc1rlFiP7/X+nc1UNKr1c
rvVCczhWfrQmLbNx+6CcoBrIW+6lvT8HiYvsVUoJBvgl3nEhXs6uYLE5UwPoG53j104PWqtbsFZQ
Cfutq3NVmFG6/jcliXHFcy/kGakNQgDHtuRBVOia+qHa3JDfImdd0V69xnBg1cDnxQbIFfKgDbCD
SUei3VhIT7UAZ5puFd8+/Y4xasUXTA70G6H47ob8fIZfyfqjGjBwVoun1UVucwRo3ZkYOe1RHeKl
zhuOaJxeFuHeZeGff36ThkQqPDuypC3EI8EZyNjDB4KN9mfOTJIvlHynRDWTEHJCelB95Nmj++ms
xJgGA3/eImeUouwvCI6UcBARABlxs2IOlNSAZWewV+tQDIGkkESNHaZ/tF6LoM6D4XIxKqlK53TC
kWZGq9K6Fe7AVY/btEpGmSqIK4mj71eItHTaBtuPEbSJesPzdcoZ7wu7ofrKM+2gzB9qWMxnx5H6
bhjpKx8dDAhHI+PYTjzLgwQbXEnUT6i6GDczKMOJJ9WFTVkbk0JXjWMJLY64+2oG6yBxUYBJ0WO0
8reUE7cGKqSh/ywUC1dBnO7QHL3ydtreBI8U6jvHFpWqO0zFTxbHj4NurRJnYuZmFe/up4YgQ5is
Emm9qSfQrTm+uv9MOZmRTFFE6RST6OC82J1kjrfOMVcxu+rc1xPipMbvhMJILtWNT+ISudJz0WCQ
S3y1xkQUs/mzn6IpyLx9zhTqhTbMkYESTSG6TnOhBbJI1pepW8lgEj9bPe+Q0K2XcMA7JlEFPWzT
pHeRIhaQRqLNm9I0B1AF3oUEQX40m8N/nTgRT5MRJ/+gjgE//yJDUOPNrT+7utV+QSr83OmZJ8oS
eWvImS1U22uvGz5zKxKlL27BwHBtwx80EjJALk4urNWrcj4Yajvm6jQG6BbKlgMuZSARuYpJ2dYD
xh0jT1/SpohQ5MguoVMtNobNA+r33nI69R0lyL3CiYV3fZmMNbdHk7XWrb97w8f9BP6FuDfF5xNc
loet0fT1KVebbFUtr+GaDCWdf5KDjLw/4qNUkzs3y6+GdU+i6jxZvIOnsQNUEzBLQMNXroTytVmd
yJJZMPbQchbCKxv25iedTjY7wSlEhx7sqaAgZDdtuiwaYB6wPzSg39gzYoRMatGvUnN9RdL8dGMx
dAO9Kqlfv3Gys4/TPYsDtzRwqBIuoMqg0eaW8AJEKrNNiPjsHdXuSknsoLREUGChKKcIekqAjONP
t+nb73nBhst7t8opc7yeRbLdi6ORfPEv/nsuc4hKuqkdq+ksA3ZuIQM2AfsVzOxd1uXm9ClcQMXJ
CREC7SirFP4OIsdKUby+4Mb8hOjvCVBAJwqOVXOgpdxkszpTmp2maSMmasf/XxziVwKpsUCctqY9
17Qbec+Yc9pgcXl6e8CHBAjA3XYPXFDCs0cLMjRaaQ2zUIC0X9sWqpk3lEYC/J9myUNaU7AEOxF2
k9xqUx8SLaG3zgG5aLkHu+Z4XVdDdbx2QFIOz/GmOtcLKMkHxEJ7W6vErVwOkudYHmJ7FAw5mWWG
ulqMHMpnlQSiEJNYB7OYtqZSaTBB5bcGOMdrc5aO5Ylii+ixwVccjU1k6eB+GGMoX06pj48HuOGL
kcxn8867twMURVkUe/P9MeJjupPX3LPQwreWWgen7HBMobd16a5yF/hfojk4RpMYjVAVXjfc2gMW
ppjzMIXGJyoJ65Ml+YPrvrL6NaUPmVGCOoJdgGN7qTqKfJdscBQcgMoEL2mqDZoNhgeYUhPfowex
dnflIbPN3L2Xao6RYKQjxiZcDgkjq3ODpHzLnO7UoRwFN//Rz7kfW0NX9JsAi3CJ5efd43cUEETU
6FH+scKQLwoVuoaxzV75ZlwRYfiZdvY4oOiEVXKlUM/VOmZ9uyGGTfr8iSC2GgaP7TrUemtBPkPu
0KkVa0f9B3xDpshvgcEwmVzEsf2tGmIKhxo/qaYmCV2Ccg63EO/AweA2B+kYy6iXkmVq4o1k/IrY
eRcytUoMnxs6KK+pLswCaPiZyY0Hc6mavklwJfyckh3WSV+Ox7977sRHGLiu/L+Xcd5l6DjTQYk3
2aV7rwz3wZVtiTyeLKY4uLgjuOA1/xIDkHPtayG5V/ykntNfJhhoGwK4BtEbm8jPVJL0rgHE/477
Il2wbOR74ee1OMFx3vfvnXcG63sJLubE/2IvrCo4XevNpNebMywPheljO5sgbQI9PHBry1J5nx53
Q1+lZAhpKXbbM2CbHnJCCws816YT8J93t30n4k61ckC4DRAgxYFNNNzn7FV98/N3wgwXLQWXNYKq
yFD7qK4uPG/GnC0RggN2IHCmXOu/u6koA6HkMYlgRGzNWVR6R/mD6OAqUEoWXNC8+gFv5NC3lrU2
vQszOS+S145rl1OG1suL0e59MWMNjpqqaVrPARZXvyoMgb1AvCQDgMHhIJhBDtQGCwOC0TAIOPRB
AFsrNENqMs6A9eZ+2w/5M/H21mFn9qyhiP/0pwB8GIrIIi081cjRVdrldUF5wgYwZD1B1tsDDlMs
BUPYPBLjzJo8r8F8qVH98SSHbq1uUUdXSzfAW2dRtabFdBClR3CCm9RS2Ex+METL/qF+AuHYh7SH
S0j/AoPpVcpEiYFgaCSa+sPQ6EGdULvxaFqZdAdBpiQ0KDOTLcwg6zB651PaL1Rld4+pAP1PivFW
jBuPYHfsxDv0RparCzVGlH1r9CE+kto8zs9RQ/hZyjwl/1gQpE2m2Vkym1gg6ltt4fMYDrNUmHy8
n+ZNi7g8kKyfe0w+6Hwa3OtAZbtprVRKxakK0V779VfwGP6SelRvirEkN0zRLRaH4ZysIP6Nar8B
uJTuo9gG6a2SacUmvpBslK2d93lAbpNDBpb9rymBpjj/X0v8K1VNy5nqAI5nkyt3Nh8+nipG8cFY
2LcC2K+hxlJolAZ/Q7Ubk4Vpl45rs3Pmo2kB3yMKehWWlI1+gSR9x8+n26gzlTH8dubr/74bIvE+
VpXhg92YCekeKaHcS7lQoikt074z/k3HrpfgWW6CGfoSR5e6caywa8uceAu+jn0KX6WrHvCZzW92
HFehE7zr2cs4JTThkcc4DfZmiW6mMhPLdEHJ+eGtXiN0/0S2UTgpYNCaugYxoRN4Ho6MIHXTlkEN
cj9F9adtdH5V6Jhj+y0kNd9kJ0E3rzmbYgN6oac5MtSDdazJEuaD7bQNnVa/uJZsr1frdgeEYOVW
PGEf304g2Jj0gyrL8gZ85c9ZVx+pxUzaExE2rpI3NS60ccVIdkKSktQ7arYRqsI2N14bEeEuNwcP
YrXOTyiusieT9CfqXLO/bNM/spv/4rllErIRWXKVap4yw/X/fZ7Yi+U5cehnnAAbFguuCG67WDc+
F8WN/jcRhF3b/NFKJ2zVMsWmGXmDMN3AhwA5MtxyuzSuvJjVxCzvJwtWxcqyp1V3K/NCexfj9N4Q
6OoPU2GGDDUPQhFn0/X4oM02MGrRfvXmt6A/Is0zFFpPngT75n8tH6BUXjlmI7IQ07gykudXo/To
pXKDzMnE5suDmbvZMkH5BPwsx+5X/ucsapPtImGXtimZWEAKUSt/AfR38s1kAXNnSc8QAlLbMQ1D
VbCbM28CZNgfJXJbMkHFXAlnW9A6Y8w3AnxoRVuav8bZc/5oHQEubj+VO1L9AuWOzfCFU+Zix8n0
mFlqTvQKinhMuiIinlG07v2ARrjJhpnp1MxyrQusLwhDy8Eb1t+U4w2zvKhBb62Up2WVxFom4hgh
wwOyBhLk5oOawkOcS9Y4HUeOssr8N6W5qvpP4idDXtsuOUO4S0ovRwVR5LMJz1D7GvCDwaxSHqTq
KQXJVkTlmYD00xmaC7yv+C6Lauj0RBH1mfIeIWGv6RgpZphdbhDX/SFxGwx7Gd4XB3jTXrw4YLPD
/rXFRBwLiuXff1nMvKHvRhafvyTZYhDohaGyVltOcRm8sG1TlDoQSbTi3wMZFqc0sMJ4TJn22I8J
fLuUTK8L7ZCmgocnLO388IUvp118Pi+fJwhkfpmMm3Syhk1hBoVr/9nusWvGIEyjrVnZigNtTdGm
pQRLzIXbmW+OJBXZyrh01XXJ1onzwqWReW1mn+Zo/lnlD8XXgpKMjtOgNfwLHtFq3MCKrM0h1dH+
ztTKTKppytFKRTTYmL9mmsTGHjxWbJGjgPS4/oMRTnFalxPdD01bRjSNp4JwKbpjrckg9y/IJC8y
4mFVH83LQqHCLDG1XVWsDNfinv9jpumfWfjcDxqwrvWKl8jFSYtyfK3XO+e8ofFBj8RZi2IeHuvM
qkfssivHXn6UXeiecqQA4L7v4KnhUBl9Aw85mrC+NrFE9LK/Aho30qc7R7Xrqr3cFbe1Cd6aC2J7
Y9Wx11eHqrGCsq1oIUuNCMh9tGQEaRfb2SVYiOT9bW+yitYpjFhc4ciwFO5xERuAGpcm/AI5T6Nr
5/VaCnDvIhSa6py5o51bHvcpHvGtOBk0InYq/FqJXhpH9Y8YJVPPPjXYfnNPrqEbZzXClIp4BdM8
747Z/xSDG904IXXyKRiAlMpJpR0aEVmNCtwkQmcnzUolrsjMgONd0h9v6lMe6PZVFun8WJeFtjPM
kfx6ZBPfG152mTxy94xfKdJufKPuRymHSbBdizBhozhkwsnSWlGusL9bbwOwF3pVvNJHkiSCKInK
uYwSzPqKPGtBrXnpgEKmJFvJ9q+rzu9S7SlCwk1kN7MBAYTYOd7SLQT7swpg3xYo6AKaBtB/VnUp
FGY43vycSYDCi9exs4yVYiThPa128bn8MMi7hX2CBpd8OYy7Nc0kUqQmjJZiM25n1rjRQG2dMCpF
DzZHtF41zS+tpHG28UPiRLkrpGuY9DMJCmEWrTOjI6ZrsAxlqaQU7eRyf274ctl0DxK4H1WzA9dA
pruBFDpXuW6SbrGr2komphwODXQW/1sSLri732vXznIYmF5lEqJIm41HeEnWCVLDkbcbfjUycNkE
bSamwuFV17oIDCRo3yImWVXzYwTofoK+WhSzwjLsPUfh6OCsfbyLH/hVgyyRVEEvo8h7edUgGml7
KjwYw5c9z5ZIfIRaJc8VbDufP4DVsG+EvmgvP0rXVbAAbzLf1FQqz/vhl3SpM1jdb9YNpGfyuj32
tHaytVlMgw+kUjiYUJiSD7PuV1Ekxf8RGBNvHaSDXTgYH+WTsK7qYTHije0xksg9C1rOC5X6y/pR
8aOfVZcmLd3j5RI4cV7Km21ueJoEjybe/cgC7zoexSRt7ZazWgkBz/SE4cjDZhh/NeJHpsHfsFLY
/q5+FwTRu7gxPkcJJ1EUfUH23fb9eKi/yBViNgN4ToEIIrMEd9zvd1+4c5ZOHFAIRSQLgN/E/f2e
cz3tv8uuChmFmSpawG1Tqazt2IgtAKH5Wj6sD6ONUgg7NDwyDo0kQIL7FjwhXOY5iK9lZGt/3Q3j
bQfVRKlvlnmb/CnLbO5JCDJL1mu7cBH4thzlojJDp8FMKCIwpnvw9jUMZESVgiVzxwo+DSVzoN/o
Fxt7ezz32OT3/ohmEHbMrSMo7MBOlGaCew9lXFU0B5FHyWLGB2F5gGKdUdZX6y9CSlmYW5z3uEVD
TZaUFJ6tH5U97paZxPn9m03FmDsSeogH2ML9ePw5EbJoeW3VRkGZM/vRsJDqfWbPAU62GKXwnpJL
uUTiVeJoqq85QtnSpeBQ330pLsJTObZXrhe03MBEqW06IpWMMc9eaxp3S9HfU6n0q68cQWAywrbS
+ORmwJ4lip2ZPF/AeMaOis5JRLxWd76EFZLSCgQxehAb33D1iBopLeogKcyNOLJbbSQrMCk/CJXz
RiMbOXiE7Mx0LcV2W5dKOTe4wqNWcI10zAO0/7jtkzk8srsXe7Mkb/aB1r0ObYptScg+4yhc35ON
Hm+b9cqoxgvbARkJ+wThNlIcyIpDebn1MqDVAKYgt/oDSYwC7CU1h3VcTmNkbTJ36SyyOpYfyOhV
7Sy4fweobKiXys9bA8Fkj2LHoTc8nZRVj6zndDL1XM9YVwtdhI3oJc6BH3Hz3IEfxO3HFUWhRLUN
HUgd/dMwPGxHRRK8MLHY5g1A32GrBiO/dDTmJ+wYggaShBeYoaB0r1W9B6W8Ifr+dDqwF9ikHq3N
7NXcj1M2vDYVtzCuVSh9RGiJOtb6qZAmYCZM67D7sKY0qoMNx3c999gG0jIr6ruGh02x6U5d2rns
Sz/2r6Wt/C34C359r5Tv/fFf7H6dFyP9ghlmj0L95T/U1G+jt2MH4Gjo2PgYA2T5bf8u1dNXDl9b
npuLUmPGDPfS54pdL20/psc1m4Ur2HbVx2boNoElt0l7OLexQytUtbUMCuzZp3eEWgAedoPojh53
tZyLOVYPZA7uFcGo1AnQ0l07dscQiiACcOqU3joGwjqZWTUucxgH7pRFA70ZDBfjOJT4EyyRVeGT
0J6YgQYcEr31WIgwu9ciphmBxmIdfUbVeQTaFMiUoDYL7grW53L4kdn/gnvPbHnn3LCdAZ8JKF/c
jasOYVyto7v8ay3n+qBycG1+r38GEELMjRdhYNbpqZnwRx8Fhj2CwfI3iL2szS0m72uNiQZaCfrj
Utz4YUidIPC0LqXw08+jRjAhFBBhhMKUJFms63IrHjA6hl6gn69kUMwC3MSUNuYOagsc+kRqCkbb
aUIlVtHnqrKsOmqebUp6Yg/F1jpRlAzbASAmw37T+mdKEKNrBNIoM3YgUrRqt9jCRjRkyTet+tc3
9WWjiVTnR8Oc2cbrun4ldvJH8gwCXHWyRom6ISSrDJl4yXFKz/hrGuw1kqCU/wKfVvoOpRD4CZ9p
bqX5JLwkn5kyT7bChijkGJDXbLdJ5B2CgfdrnhSvDo1f9KrO7QXV+APlLzj7jP9pGR6BVUC3B3Rc
ap55Qc2HmqQ8w45Uk3/oelDXunyBX6SVVg/NqnQ0jY9e1Ob4VbO++HBF5BuEKt5xp5SRAAdZ9c/H
Cwi7Du9SEBi14UCqrRqd8qvTQrT7zD/ICTdCQm3KMG+mspkoXlwLHxmChkUwZ5bX2eNFQO47KDmz
ltYVWiUIT/V1xHyVpWY2GnF4RwX4domNnqjpuRDwXyZBLLqtl0L58mAqhBuG9pt1eFDe/KZN8ofI
povEDbz1PFiVGHPcyDCh4yrHe7/pk8M0gySLS4nD9p4k1383hj+3kjRFsp5lr/c15u/LKZVIZBUT
0uknlstt4/bp7qryj2gs6Cgm81UfDyl0TVMybpYm9jbS43+7IE18TG1ZY8hQltms8E3o7KNb0Aw1
I680CaSNK6S7w6lwvunlr2wcCjkpFxOTgyoc0tBmmuU9qKAFVkGxpROL9vSVBaBwJGtI2a5O1us8
jwE99i7EieELkEh6lSZABEyzcvRq+x4JC9ctxk2v/ESWEA3oEvAF0QowMwNGA8I3DrjEBHJ5i/fI
3eDJ66eIPxtltwuo6Pm2d0oCGbQ3NTjTn1sUbGJJFG3Cub9D0NHcfmMvJc+4gSNyEFuGqpzaQUqL
DhRnir7he4vtAyiVt5k+X+hJbJXmE1zP+XJoKKCNFqE1gBCu7bZAP84O+3L3TGn5jXl5Z3kTONxw
OZrPu0CpeO7J/X9QzXJMXwEXUv4T5ntnuw4UGfzFLohV2bYiKcw0226GWwPcRkyKO6YSo+jdpDg6
6+AQQyobJRCZnPFqKYcENMVfl8S61neZqd4ZblNSRDzdUFyvcHI3h3JuiDfOHHbYybKrbnAJDrlx
VKLIJYv0YnrGGV4O2NsPLMi8q5XOlBrmZSLSxZhHbqieaBxAmnmvZz1wCXjPoxlLrdKOuMah+FWG
rTYM47CPuctkR7wV1FsvNCm7e0L72tO7XOvl1BG55HoK1J8M0XXJuomdZ2uVRRihQbBCE0RG1c0u
gB5Zd2BORtFViQKKSTPILpc30R/i81ghXD18onTbyul53FT4gg05fiVoaGjMJ02Hb9D41oCoEdEh
Hwlvj3mrQaPP90pzCs/Xgf3lcMduzrA+Vu2WibcFHgSF8WTFlbWday/123ZWAqIiBylMxvRK1QWC
qTJYvOo+ayTEHKIIIb01QvqAK0B3QfSK/MIP6Am/ZNsk+z/bkdlSXQeYwD0/QENtis5QYdSB2VqZ
g4KOOYmzBonDAbuQlbyPW/1sPvqnoAZ+NPFTyWKgENsuubpkfI6SI+ns/NgBPumlTyU0l9HrXVkB
6vkscMK4SLJa1ioMpwg8g506sm6/vbM92appotAwGl/mSb4ytfH6SkHDt7M7Vc1jFp2aPUONDKhm
QX+II5Sie0Fg8++eZ/qOzNvRDnZX60ddvIroA7Jbn7lLustchlDWUzdBWaQetgI6HvRimwudILvZ
/KARW9lI8EBxIuPzMsiJ1+lcmZEQogJzK/LRKSD0CI70Rt9PH7LL/8KF8DqjwkBwc+9fCKbO2uRc
DQ36JFT2fVJTpYQa880A8jGXxPrZKfyHcvi2BjHl84JsxbLrAGbCAj8P524Bi+jG3TOQAQDNRMko
eskj9ZC04uItrDYyaCGBhDGzYsEYtavPdkgba9unRde4Ij2iPKY2O783sxe1t90kNr1vQQo0LC+j
6DDF4PDbA2iQu+9VK8fCh17mVowvQM4w9NshgAi5TBFDMz0OASkAa/AdR6zi6G4Y0xkqrJWChpx7
YMFnh8yqbAL82W0xI4Up5G1nw6Gucyhu/wV9md3HHQRMDfCz+lVfpysCTaZufGd2d+9MTW57rIL6
8oL+BlRXswpM03UhZ8hSBrFvD3gmCJEfZnnR0AvbTat/5ULyqrj1YtRcjtCZSV4sFOpXQ6zMcpZH
VjYQoZNig87VbBhWfKaAxkyL/gtmLndB9NKZchnakwVc2t0s+DbLifpp+s4m/ixqdJzJqTd6jUZp
MkKxab/0A5JC43CqJOElnvczXQg6KHbbjVnXSHjhfQobjHBskdfnsPpqGirL+0bTmVZL2Lds5GN8
Ic6Q4TwUZqNQ1DHnUHdC7gjilYKrLBExOK+sRmikOh4tvcSvjxEwea53r8EwXQk+jPW7yDv2Z0kj
pDhgmieoFwiDlt0GWlCeHM20TehJLu9EEj1MMaZkVQyYOqHM1BPRRV0X1/lB8zmOW0WP2adWaK03
Wc3OFYGZXWYaVYN2lhDSupGa3/984hrD+UzKIcWBseYO1UYWP5Wwr8STq1DVGBv1QZpRcnmHdR4+
tr/+N2Sf2WO2GE9tm1O2p/zgH6fkYH3LPr29g1RziPHIzDzuN8EmLyWqGR2f7BCb0keQp9v94B5d
tylh2Lx7k9sADtjVjdVWuQxkzPw9vzTcz+VItZUx4q9z8Q6B3lVqAsP9mh6uHCR4/DVYghxw9xJN
7Ag9GBywPDQfLJPw69Kx7oXntxNLp7TmA8Z3aeB8vGEmRNUgcCtE8MxdREMUkJczvlynwu8m4LQ5
zB4ZRDTGP5iak5hNN/G6ztisKY/PHApxO/U2AE9cTmiKq1uPqWVFdIqw4eqiXtqfm5shVeeSujEZ
rjKO0U44ck8qH7ZodIfOKCbMmhauIQi15tzZe1L6qil0gHSv85blOXFuzS6/XxuU77l2q1V1DUAx
e2CuxUOL6IEqutJ5OWuWtg7/lDqQGh1k9knN22ZWsbVtpddY2D+UfI9TSkUKGS2poy30QkDjIxr9
xj+dDgJJ1Otn9/AErlT6PfKDnc8ds4J0S74+2kVw0x0FQ7hUIAGmNMcM3+P9bAN71lBUThaP1uCk
vrmWIXpk/2Qt+WgWajKXhnGxJvThXdrObwZakTtmN8JxOLxRCX/S/Ue4lHss6axlZppeR4ZOBSqD
+b0ojtTr9D2ch5yV9UWozDmbB10nuu5j5TicFLbeBzguFF6d5VGIgqFHrdObRpwgYDp14c9bV84r
hW9HPEFVHvyAMpTDefYFA4LjjPA9qAGLb/w3BS1uWNbaraujMTdI6u7+0UGEmk7+4gGLzDrBJOFP
V+Fhj/Qm/4PtuVQ7u2r2sSCK6wJH0IbtO3yaivGUWyINbDtULZLE9Y3FkWhFJOVdYusAni9nHLNQ
TvLHlcQpC85TxXIZIuvc6WM1nJRUSyOictbh+NK9IGPjfqu3yaPWdEwz42wrQINRPkHcugJhls1e
UMGrCZOBPtRZ42a7tpJyKXlLCWsEpo9mun5IAwrQ3RNCYMmQ5QgggozwBAhiw4smaFpJFdQXrSXC
qYDVEa+DEGv1MWhPJE4FAcDtt9l3B0kyCS1nP5zRYr/hAvaclL9hG0h4ww8SVR3RKxP/dhtSkKt5
sRCyfE8d0IKL21BCXW1ObiJJX4qdIKn8WpmnQ0ROHqqVztxebZsM3kJfB6nYQ4eBjPq7LJpyeWpL
KWNRS/WJJBfMjzKXL43UAycJlKuxKCrCkgUPdwcLwmzjSGC7bKpcS8sNv/zE2xgb8DXmfuZE29w4
3ARCUEvCAygi30AkvQxM7Fj1PmbR1tsynuC0y70Y1IUMPNMC2Q18BtRG9QlR07JUZKIKDN20/DvB
xRltSWbC5tlIiYo1xwYDVPJUiCr7xSK7x5DZy5FiMGTJ75YM9hVnupnCMwRodlNxkQF7OkHpm510
byE2rVhW1/48VszVkPGDgXeDsvFoPmYZIMlsmYP+Nb/ewfEPQ7O/AXX/cBtaepOKk4JLxwBb8wy2
zgogDObx7vmpQEc5nTdhavDFzyHSKbAi2IjLHxsYfprbdGOrO29Ltw2MQJlJeAQlh5NCHKLow9EW
xEOWj/4xTwtH5RjchEObF/nxIV7DfPpsNj/UN/GN6pwAJ2jwt2i/uZDL/rJFO7zpXw9gTHFzeaxY
q82RdZ5jZIK9wLlk+ja8hR85gcHRy+Twb6VJJA8JfPcSlV4a9j8seL2RiTgcn1vICwf3l9kD0K6L
52hRfpv3mqu47vOk/tRhrrxwTPmyoJOmDsznM+KmH5C1ob6qGXbBuJgITpZZiYL2j3jxpRFVBMEY
Lcl75/n8to8eGhgrz65IgxPnFN5VglO9TQL8T2UpZ2OWRAA/3SY7EuDcTBVoxlCwIVzRKBbixHtG
D76ug/Qg3Z1go+PRQ/xhCf8CuQ8PQVgVUD40c8dEhL+TBBeNxQH8GzUlKABAqJr+89TEZqXBrW2v
BnvzKs+3KBmJkL38dcik7V8UPoX3/pXaKAkLnUpb2nSguWeCATIfriIlMWEv+0J1MK3uARzJf0v2
PaUnL5FWF1YPeaid3Pb8S2LqGjyvPV+SKVHwFnxhfl0UcerKSLkhz/1EV84oK0f0C7IAVnbRsFhl
FbWiu124GyL9evTUYD9/bTiIJDLhvMYsrW2aRZF7nn0r+yir+XK5Yn84F+Yfn0fZKKU++MWlEhfd
8oUqVu7FxYPJLSwRVcpkgULqFr6t31IkxpW4kWhzS8D8UfWQ3WISmH4vj07D4a7CroS67750NW8u
/mn3xEDFz7IF4I14LKc3GRPdbT2clSPgB823JTTNM2pzqUetNcEMectmKePraGfmZAKll7fyh53b
4sefotViobGrs72KKH1jZJf5LY9AYlxYQ1iyA8A0/nRgTmxCol22lSXrHIcTbbmcAADXxP1P21AV
ERRKzUubtlMqKLNfV3CSMBwIPsBYdUqsbqme1OrzBVpD+jNqOVA8BmcEnV6EodMzbrmxtWuj4Yuv
IlS98RR4JXBM3rIB2ERQ3uqM8hHPmFsVOzISf7U9vsKus2cb7i0brqgm6MwuGdaQeVIwHyooiSzm
sIlAzUY2pnuraDP6q0MzrIzgjEtXJFeQIbWE8N4u1f8bYK9jEZPy6Nu7Y2Bv8zKmJP5QI4eCubgi
qO4XOlIPpuFRz0fQnEuNSGctDupWo24qNc8NZxGI3rOySQrJR1W5fNNico870nvkCBUs7IiNnVnv
S0ApwdXIH/qQszNQOl37iZGWjmHLbthbB8/ti7oeVtVoeq9RXcSvA4k2/TKk/w1lnXIZJYFKXRBO
L6bj4oJWT0nusaxo///pfuESt8/XdkU5gd5ECmW5GBnR91c3uPPo5nc0rRIyA3RIMHNOfuekKI5p
zOBEfZeI2IbjQ0d90/uEGUhMDfIl7gOBYDo2TeitpvLGejyiHGhlq26EqK628kNK6t1h84hWmBXp
9ahcbd5WHVGBxv+zB69GyDkzz+rJaa/aWlKIvvld9wl2sUpXnh43ZalZ+6cY5xiRndBQQ+9vS+8p
O1BcL+oX25Grw28xWZhAG3G0zCDZaGKJoQp/iHigN34mHVYdJrOpK/p8G+rjjztcUZio47l/Z/y6
4LLsmtjR9VhlqWdJ8ZGXAgsLA2yKbnBolutjWyv02UfPise7ZZzIkmvyet3uPFcIK/7WovW+sS0E
7z21DbMxTcGiM8W68gN+9IFhb4L7xPxkdoHzhhr8QoywF0Eed8cMCWgsJ6sA0h5PfUG7Q4EVcTit
YWDxDFl78zr/y6A1BHIhZpMdzz7Ed2wwkp3hwZtahnIPtIMN1JGrgy4SQUS+VcipjlrgjezNyfCQ
WFSt26sRRJ+q1LkAw0PQc9f/GjaSySWaTRP6+4dFkA4DNJmb0Du9QRLgcMDBVhGglnyiIteAsAFO
CplFwJt24F+/Wktlg1INKgZ1Jq4+aCDjFzwt8zYur6AvQe5YZphDqn8FRBXhmKAUYWaFieU13PZJ
5kVmb2qaJQ/VxUVGVWpdj22BJJe/+Qvt4z/jjFhH1gP/n2SLo4OPro/YX/Wa2EHQ9v/3iegk8KpO
rw+0abrxv9FWhN6ffu0fuWqKIySHL3K6+f5QRrf9PT3f1iwJ3kd2W7jjaBMW36NvkCeVPsAjGQOR
mYN7cWZWf6zRxdUZ5dh+nOiAGC9w7P9j0km0VADCcfXxZkMWT24vMTn/D1Ak0iT2aIyRV7swpieV
LGDF3i7v+pYzUqH7Gp3TIVFx+XgISwaU/E/8XUN5TSp8BgYs1lqsikL1RTRCbrJG1EWnhNgYCuaB
q73SBjkx2W2fpMKnlTs0Jj76Yx/ARe+ohvbaY34Pa0NUcJQqTwo0ecxzgAll4I3UhsS6WuU1Oril
tnpEmZ4INW0Oz8BmmpmT2GeeCX0aWi8zwxL/B1V813ExtvfPdKazG0w7pvJsaSgD24b4cNG2zkCL
FBBtNwqlwc8zxIf8azsfa5oyHnzstWMSaawiT6VKV0A1RzAug8W4qxeFZCFmm3+aRsKwY02N9y27
A4JVysBICp7BWIbLm3GwuD11fUnd0wk8K0AJi5lzo544U+jQhy2CJHF836NlUXdN0jOEGIE6y285
XmSPLbFimjOdmj1x0jgoqSJt0Txc+/U4K5z8b6nI/6RpBrYJcIPE5GY6Dlza2MW0mpybYgnA0mcX
sYBWrQCxGSPzVwIDc4RpDCDAPbtue6KEp76f3J4r4f8Gg98HNvKWT+TT9qOQkOmp95sIa1Z0+2pU
5M0/27DevH10jqzyUI5+K49WYHP+oqcN44CyAszwVAobRm1Dg/0kJhAXJEGhk9wm3c+l+boLACkY
GNH10ZmQ11QX4+iL8xSrwFL17xLjMNyZoe2IJlDlmfJ2Cc4zvXeqghgjoV9Uo8oLWO3MM/2Ej43Y
hM78u6eQxzaI12sSWhGxjqN9AALIRpkG9GDaO5TSTNSZobRoGclqpcJf63YoFHAcBJn9ACsypKkq
WwYNsArTTgrCaSmZ86WYJL2G/l37s1fCK6FB3SqSL/oa7TcFzHMcdpuHaE/RyfWmiqq4aejsFauL
J0wCsbnDYsviN7HuTxMhfwMOuCN7GFpWcXtNK/odBHo2LpcNhffn5jXAs1ljESZeRnt1rUVYlHhC
zaGf+yDNVxry2/q+3rq/GVdiLe1emYDnOfm9mzfJeaCNgEjNnIbUHuPF11aAsb5scyqNMx9qpLv0
CFrmGjW2pqOllv+B+reWy5iYD30mVNL9Y3VuSKKzrgHYc/bLYOAwKnfvcqVOAVfgjLMjnaAueSYt
H9WzgQZOdenGT7gtHEYEGJKAwyTRP3rrBAbzGaCaFrafxhHwx6FNQMuC8VFetmW7QBNNIaCK8+Hj
OMV4BaCCrrvwTmPVZlK3tFnnIPTQz1toP//4AHcl9mBpjbN3apZqRPnnqRGBgo3rwgtbXoey2cci
cSR/PJPKxvyPbS8OEuS/ibdQ4RgUfu+b0HNWJ8eDj/2O63xQl7u8rG9goGLxWyAF1e8XHBK5+YQ4
I1Ff1TrOhQvo+JYDm1hkO/SqpTRodTTSdi7wLtiJxyDtL/pEURA9v2KAlDT2dLkhQkyN74KHP4nR
UzNevSNZrU/EPmLSLUECuv4RrFztClqRJjLqQ9eNzjWuPt/oGV7u0aLbZksAxnO9ZrydBPNUB85n
O4kmQuIsFIrHWBhslEzRlzKWdnHHr2fhmA0quwyR5z5OG95uJQKnwGAENqusrQLo9mehIw0KkE5u
ViZo+QXL13jJT2rxkQnpxMeJ4mA++HnmMU1V/IEF5TebJwfIC8h/nAMY1FKqb319kPNh0n2Hj6ER
4VRwjUnbC2ODqdK4x0fs63Z4afq0DIVXax2apU4vjmp0PJ0eWG0FN1b9HJbIc8y0nOy1qIg88dBY
oxXWWcDY1H6IwLybrV0ymuP7TXJg/d1eF/UY9dpLoVR+WygL+g0n2u2RzSo+wcLXtAiEFdE4qwSK
+35HCJn28BGNC1/T7s1sp99Uqbcw09zXJPfUotIjqdwbYJEKVDPEgXPgjSzxo7rjoiygHSNlKpvI
ejoJeEX5n660nBMZYUQJsi3cBRIl1CkJ3fGog9dtCueGnFt0TLGPyo4bzyWbY5GrfQKYMEuN9iVK
zGL5QpEF2FwC4+TXTcTOvswwVVP5n+mCOvYqW8RcWF+zp//HHNAFxJFZKSO/tX2qxxlM3Rz6GNme
eM4yLN+Zz7u0joPQ6zryCQ7TysL5fu1IdIa5MdLhfyh3cga31RES2mqAziCQX7NOx8XULQga6TQN
o8RP6b/E5IudXuhuD2Ij0DcCOcVuYNLteHDHLX7b6zcixlcv+jmA5dvwooIRG37AqonF7xCMvRI0
90F24pRJrJiQB7NEx3Bt5cYf+oxQi3m57su4GaXVfPwhiY7F6nZBF0sUfAP9yGUqTJ2xxXI4ZsiO
Kh1oWSrwDCE/AJrcAA+4EiGoQ/H5x2K23iHkOZMJRtwn1TgEljWd5pJs7r83j/ruxT6WRGhxX4op
Kf3KEZ5lnJktghKjA0lNC8Gccz9DH0Hj2AFjx4nMyzKSkNPcTm0o6M4z+peqfhUUOt7LkIHa8zSm
tjPFwaL17sxPvBxxQDdwesExEVvJ3hht3hA2jjfzS240IyfgM0atg/zvAn8suoSGYKssQdmsktLl
5w/xQfnyKCwX2i+yuRP/dSCp5bMQ8zKLnV/PToRNuCwWsWS1ICpk6c+zIOCfyLi4HKdLpsIiS6Vc
YHbQgJI3IBewJbiKh+eh6y4ep5jz9meCKD+0EDZ/TGf7XRq/vULnjq8l5Y440B2TYIsVNZEoBjah
TBYf8AtB9UyWVA8kZ6GlGgRgJrYE9eFIKIyawXoiWxh8+H6xOe1Tv2Ixmcx+fWR5AMH7N0IPQ4Y6
nQThEqwj7eBuJ8fbo17nj8fUikIeA+mLODT+hBTQ9O9JD0LJJS0xFcimgpEPXzpsZselhRhLkEsY
Sna8ir/97muiJ3hzoOs8jAJm83Aens/kkI8k2CRsygcnl9dwFRBBy4THXfXMWQewG4kNYdFDJ0KA
dyQEr272Tj9M/5LJKhYWyhwOEZXH+UKfzGLruDRV9LAYAtOx/TpIObRdgOkRFyemphBlE9pY6QDw
6zs6LIXAH6HM1sRhf3LkuABy5Bk0BliQ5gmpIWQCWBD9IPfSET7dKZjmxkwISRB5azsevx8waJTf
SRHhgG2ryoVbSOI3xdc9nnSzxKPJfubzIOIsjSqPGYgGDR/47gP7P9EYGQlrOUPn9YyAGLSiRZ/t
3a4+VAkeHxtdaNJiOsEXmPZWxM6jbRm3jqEmFSTsRgGMwFhSVHFcqeN52uddKmqS5cnEX/3smsPK
gAMz6GZ3ZeDToZozRbT51RwVCzHW8rDLO+zB5r6AwOmtHIp56+lg/DvonKVQ2j6a1uZWl1ebe9n9
YTygUdro08n+tqz541qInXvrwEAgVCX0wyWLD810APlVpyagRp97O6Q7zsNVvBOwpBvgeY8Ty/d1
lIeE90PwAYA+b0nU4lMLJvJb5enX+mzn8mUpNq7IpBjSdrZkmvooi1tYx2KVm43VAgZEBBpbJt4+
ADcxa9cBk+Vu167xjpZsttp8H44HurlQFfvojteOFZ91g5Qcap7a9bY2YySLs0vf0+YPdbr76fHn
a3Yjr1qbyvUzTB8QKx2nUByOJsuGkT6ZnsxhLODtcY5abKc3Wp2uU0/kmKFqeYPcWxwqzR0QMTFA
Mqk5Ux9lPdCFNiEWBL6UKY2l/VqjnKIvIjn7tu8P9NxjjZ59XlFVxCGreGLCNosNlv/s46c32kWc
F0Ee37mJaeQpJKCUxdCN0n6rFb7krB5ET5ncFE96OUmUV76MvZF0M0foWNfUZeA94bgbYbbi3rMn
AAGkv1XNsePY5s4veAZ9ipbK+YDAfi3jkCn1NIsSXEf9C6zJZ1Wg49sZRuw87ETJWlLtQzxNR5fE
OZUrEax6+bedsJm9i/bJmRBV2nx3xn/ST0KiH38XYzwt84UIu5hhscPaeO27fsG+CJzXd/UiWXFh
aUXdHaJEVQKPvDszP07Qcvy6tktE49rGqfJtWdbB/srGzYbN1oL3b5/xm2ud3Tq0YcAHFiIGEJ6Y
g5RZImahM95j1Li/mCLNoGQ6sdllhKdRhw5gcZcZkev6GGj2d2OJ15eayZeUr6raKc5Kcu6UYD+t
Yl+nyq5JARsQT3mkfAaqfRY8wdEAhcinf3XrUJwBtyfeL0o6sKzCzNbA573k+00jbQxkDtbbStnc
Jv0t8J3R1u/RawM5MYjx7GadP8EwkHQSkGM/1vLK1s5bPmhfmbGwVTMxLR4+NeG7gSmvVaYXPWRU
bmHrhpOKz7dI7UsBUnqpGb89+3VPCIHJkijjpN92a9z5fV+cztwdQLymFkSgusFhBDOzFUCMrNJJ
XQZKp6eHSUXUgKA8HzcIGludUlx45iu1ewWFesND9WGyG3EglfyRJV8At7jkcXRLFpteMF39i0yq
3pFnT9OqIoEPGVhshB7FHuRNhw0FOv0iJNu9VwawIF0FaX6POHNE940qntOt4tTHTtLZCu3bFA6O
n21PgW626nBoAlWVn+6B5wjTQztQr1rw9vWT/ELUrNLR10ParS7xM0mp5BSEiYW3AvBddXaoemlF
fxtBUwub2GWLpl/clm5S8dhLS/Phh2CLNJN5xYPr4P6/wC5x6dDDTT6CBGr4uk6Ra2BlG939bxHU
v0WLnnAK08FSm11p5znleHKLx/Yju+kL9/0FyP0N22Xbd0kuBDSOhLJiJq8hxFJfSzTmyuh0TPgh
coEA2/4BFK/1frgcTFRZ5CyfazYA6/r5CI4RfUx6u7XDp5mmJQYwVzzL/2MaMdicEDLIioWEO6eG
h4AbRnjD55C2DEFe/+4xEW5ODRd/15YN71+tw14xb2sThmGIj0Qcb25lCMaOykwXvJ0U/rGvqbwd
FRLJq+qoohSfUxIEWti6u2zZE+SQdAAk2BKkmqJ/I4tQB7X27YCof5BPHI/JJXwwL3pV31t8gN7G
6d1DBMaDxFWoU6qkioyJWsvp18CA5leWr88LrXNZPWcKEDGE8AXlPIff6QbGpaOhFjXTZF/y2ADH
KyAHVun2kbyE4jhhbrWdh95Ej/EU7JMDxt/HzJy38VFmRIWphqsSHcKPKbZwopAtl4BpcYYVEAN/
w7rN2Cmi0h/OrrJrk+H+r/LnogbQ7nTK7WVsjxmLZZy5mfMy7WVWvFir/NB1/t1h234ddTUgRi3K
5jlyzhDykdFaYXrZbaZxcKMMg1As5SA3iwb6TUb5InqMBGce/fDMJQ7pbEVSpk72NuyBOxyV267O
Lvrt8mVqnZsYQhh5wrvnc9MNg30Uni+2dd1sbvmgiUiUtM9ZLAX8+2slnXSI3P7FgXZTs7fFrhng
PxN86efRz9H1OU/zUMczxYx8tr7TcXXFU9uH4QSweqe8OoeBHci0YSS21k2rXM2t2KdZkGy5c6Ce
28YgqS8eGK1HIU6fxPJmC0AFzGfD/9q7moczXxnhJMiTxPT6ODmx1a8We4O4LxOxG3EQaX4JjYI+
10UQdrFHoxAzjT3INZ4JWpjG6aGi4yBIpDq4+j0wFgJ+ARNoaOMK08QW7xD9Cmlix5H8i7JjcNkj
E6kLyy/XBxzT0FAiyo2cOZi00s3Eq6YVjkxFwmWcI77dmDA1ws7o12EHxHIurMlTJfSQBAiizRaC
TLn1QbBygDpbA/66lsCcdVeYENp75FwqyqpWBQOKT59MQHbTd4hmPuO+yZnTuXaM8lkD+GzFaAbX
4ZF1HLmem7qrSQXNO+vjAAgRQOxgbFb/GZJ6+89ziHuY87Ab2xLr6lhNPAZNxVUSJblNHLcYLE/K
HlCoYYzMGyJ9Y5kXQfBhn8c0dS/omUIJAF25QSYk8fpcRV77pk9iozWPf8+WaseudeXDztePABrh
cjz+WdMdcf253jbHcLJhmp+CLVWB15H1eAlVFhkJEuiSdm/ouz8uvlea7O0PmAsj5Cy5xSXcK+wB
zRHBdRnZp4mh4wKrjo9PvkQ3dsgKlD2Jw6emoU2kg84975K2aflKNS5ISO7datt76g12WQJoWym+
gVcaci7K90wWdL1x77Cght9W0TPEpwml6CBe1d/ZPqnIvf6bWEqXp9tJlh7zV/GxWSH06WnWfh4K
0N24Gu4kwH20yOKB2o0cASEOAo1TEjg28DHtvkHWqjKc5G6AaJZ+YIuOkIRU5qogA5NXsqD97izl
+Hph1Oxjik3uI3Bu3InLNnsulpA9/+HJ/isezmqXveyAnF2m0jn0/mQARCfy1lkqIzxSXfWwM4s2
5rUk59Avg2y44tL1LdnsXmS54Fp0BZN1mZOZn/XqBA0rgUUzCdk+tHQonXgyl77TIa2FtwpYHHPb
Ngw469Im3DN5nMW+ED8MztCD8SkZB/07WhKIOGj5Ev0p34V3cgbT+XXC2e6/l06Z4D8VWqfOoIQN
Fn+16tz+GAIp/LxDQVAKiZpY3QWwKFBEbHBh/Qba+HXVxO/6rfefDjfPkFocLjKbGGP3blg8+2Jz
7K+aAekIglo96UtvWqiJxDy+LT1+FiTcMZQkF0JrsOWA2op3jUBzr8lfJIL1kmgUdIAsVR8LLdbq
spabyrAqMHmSSL5o2AbLK9rPBkAyy1ZFjaGoDHu5A7iaCp8zoyAOhrmAPElJQBr+X4S1uDQ+0tHJ
Y4s3ND5PMdUdRG52lQijQ4rqbkNZDeZLX2PMhVUP1jyHyCsoDG0qUhFqFwOBDweV1nn7xV/fNUl8
OZ/XmWgxmT8oFp3g+EYzdCXraK/4o2yfe5SX8ax37QgyfT1Jon8y6EJsiNbTX2m6AtSQd71zbfbZ
SyxIZsuHJ4zsJAvcJMq4+iuTnHXqCUiU2bIY8TGEN+nVwm2TovHZbG7Kn+TJ4OS9l8P5xGhHJgma
QKCbfyzbDtyojyVFgxsjXn3+Y6kENesiU3CaHFNzIo9X/lxIi7skcaOJ5oGpKDH/iKnMRNQpobNS
XN6vzRDJCqJtATpJYqgouHNma1XJ4hf3vwuZ2fuUgcz5LLDUth20qkNDTW1zfXFYkAV77TmBgP5B
AV65Cu/cF1ewEjJ4ggvu2n3ylUi1yo9V2cX5rve8ktNw+HEnPiRCk3dbuCnRKbueqqGQlIyNk++x
is1LJDgJcbCcwyAM0WTTevXiHIHRwNZtacDfiw1f9emohKm8iCJw+pJwmdzE7Aikkyo+6vNcnnCn
gmMLv3o93Vr0jY9SKgnXYP7NA4j3lhpn7VhQ75UsUQdBs9tCZUoZqEknSMLVd706g0xJdHx8fRTd
TjgmD5ilYPJTA2cZgAPzW2x1FKVksLDJgzjmFMQUpdm2ktv1xbFlMQDhV2AMOE5VRZA71DYhq40F
JjnggxPoXBvVJt8I2nPqx06/47sc74DtPg+ZMONVu0CG5jagfVRIxXXqU7nWyZV1iy7y1J3gyr0H
c8TZ2H+B8Nu0jmYSrVGymcSuG8r/Ean+ri8oajlNzM6qWyuyEjlyjXYLXdbXxyIkCGcDkm10vkxG
qniNwafEkG953resAQloi/cMNOzYFrZ3K+P07lRsyJ8G7+M9TKxYNEBU/c0bNefDUJlV9EIHbW/t
zSW6KQ+btViwc0dMHnrsBJiuceikNRDydm+xShm4pymFgzo73I86fKbF2+FkfUPEFVp+eV5vjniP
BAYjqivBO5N+c6ZNh3N1n31oaglaU0LW/fPEcEqTtUPgK0kX/JuII9WKc28EHUVuPjNTdp0UCII4
bDwJqMxsFcrsPPudaORT7/cWubuE9AQ7H9KN1LzJIPWwWpKQzKBmAQ0lMLdH0wCaemjkBrtT7C2S
ppw05Lp0wvQEGocUkEE25sTNG58VwrQ9hVahpycyadFeKGjTRCjNNWGNX5zaDBKAM74Fer0dwGz8
lCMMgKSgyBPCy/FkLIyTTdrHnkbhiKDTe9FhDPPh8OJJqjTKD+Y1COSWtzHMjYgQOw9SSsReYIdD
4FqzGYix9MbY64PloetvLJ4Fg2Ehzh6A65LWf2Znj0L0+7ola/KwlNoXLMqfyykgar6qowIyyGsN
Q0pFC/yKLpyKPRVFHDgxHMzkKPFhhn83zQDnr3mbPMRnUyC9Esnqe67wVnEhv38QKGb9C+T/4FXx
kSekSTwMiMSDRrGv8slddjSMC+L7a7Qf4kOiAGjuhomiwaIgnuOF4s2fyx0YaWbKTfye7bvn7GFw
ESxAPV2HOy7lt1boQa/AN1nKFezK4+yclxUCO5px+cf86VYCL7OiH4zuL7aEIGJr5Uivohk6lUvt
WEHrbWuTQXX+oO0AuVn8ArqcsZS8fmN1bP9d0THpMyYVj+laMyvhIEU9kZdb2B9IB0BVSJlDDDaM
2krdL4FqjddCLXPNKsWBpN8IXXUO1ABWc1ewyn1k+x4lGAAeB96grbn2phLPVUFsUHHZowkDqoTK
MwcuHApNO0zIjANIdgGqy2GybmpgjxHCqzX+qN+Rz2nSz6ASymLDor0uImJYuKKs1P8cCD2e12vx
xrtuxbUd4c5n5PFZzM303DOBpm9mU2aWblzhjvUQE3h8RCSlUK3ouQP1G3nJZKE7FWFRohy9tiMv
Hu7Z9i9o45MkVbBPA8mi77ZLF6Rp2pUc5H0NKx+mVEzI2nyEquo1u/5u9OFw62thqpPR+L54Ae+V
/sYzUGd8u3WcIqMQ6Ff1rrQvZ3fhnnmZCfqAYaEPG6G5AKdDmWUOqeTP4cJfigQBdXG/ZpjAJoCp
khLKPy5fVsTja3QkznBfsSGVrjxROGIYgRCErgEPrlttxVKdIwiZr4LIL8PaMgbCr/MESHGvCDrK
AdlIJAnhx3pfuWlTQnyZDnYnQhUHMlD2RnXzRyQvf6Ri91M9emTnn2u262WjXv3c3CFFndNsoS1A
4xWeC5lGpZOab8iW4Cr69axkONopq8wrPFo1QIOTDwy7Wng+xcR2MmvjENxcPq5pM730n3fKkmyn
W6seyOwedZrKbUhZ87HmyiPYkqLe0PgNJR1z8rqdeweBxoDtml/ryBTTheoIml+7LllxN/WPqHy+
9DyykBoNWHnq2wFup63YODqzIYjh5hv0OPMmhmudx+6EQ7xAjytVTRkezxLmOr1lEi4FEzbstYGu
rA1S79XeM3IgR1SMZ1u4Tkkq507C03aaffcS7+tKk5ApdE64uOZZ5ObTB/ePY/86bVbGaC8F77Ph
B2dIttIoiiuBnn6kSXv2O1BhQXhBTGXZmy6uRgCks+oG3CcdkKk9Wm1m4h4F0Wimc4nq17eF3pRx
xSaETdmlBGAqG7urKewk1z7hYCZUssUsbuz8prjSfOY02O7ARs6QR571AMYE/lwL6uKyf9hHijkM
K2cwUcMdP0KhnXTgyTzxypIzV7gtQ3OKQw6H2+wzPTrhOSKE67mHetee+Tr3U+sy1/Er+c6fRTbr
/HFqwbHfkFs+BN3Fhmlj1dvTNw+fW+Uz4Z2hAy6eqlwt3H8xV+5TD8mx2EY6Tzy2OYXtsyO3ln7s
NSxEG7GJ/2XSDP1qCZYjMwbey3Zz6nVZqljqZgYskKJCy+plam85MW4p9B82IHEJ3u2vYO2baIdf
UwBaoYrd+MrHY7Gwzb3eeavJpUEAkca6mQUi40f7J+u+GbM3ehrUKGlir8DxOzb2xlPbgLaUGD0W
QnSvorV2sJEmFhE3qDi8V8O9RMWU8SxAwVwuY+0Ew7KHwk6xQxuGhMlM9oVw0ad8Of2miAVnDxEo
uhTfDThp8ya31hLInsn30Im4fpUxelsLxrSrYqHrYZwIHrp61JWXunNCBnGW+J5Zgedxo7PEwhtF
ZSHRw8eVZmUodKIZBdctM0UBMuw7bqHiYvTp8lBNPN+oYIv4qE1p9AyWlSWA+T/RETrspOYUt0Yw
lo7QoQFE5id0v4KB3wt/BVWgpWNexjtlSh3vrXq1OsW0fmz2regHR0m4jkO0U9aZgsMMTDihUBQt
fxG8XFx465KzGkGCL4gwtjbgG0aCTueQjIYNQL0BHu8nVZWfsmZKfK0i0sXxMTQN3C/Vg9LgpfqJ
1NF8vzM5Y4Hg9P6nF8fqfWI8RV062xZ18xEEt8szSO2DN2bAxwuV32eW9gwia9vpW4qgqW/9PURz
XqOQv/3Zj/3PUo1Dg4fteZqGWlQrmbGrEpNbYeI48Kn9vE+yJZp8+HPVcOrVrayRpKjGUsiYJb4j
Z7z0zCZbatqBTGuJ0i6JGbkZb2NPDHWfE+dpXi9HuO1yVWlmlYP51VygTxbBSDFj74M1oNr2o98A
If8qmIsnN7idkfg0HYFHTe9JQzV94FKqT41rCsq0gvdAZ/+Cni9SR92/Se534wLM+guD+LhpIV1S
WABKVuqCcyzCvukEN5zEW4D6qOELF/Sr1W95/VtU1GLmMdX/AFOEhmxaJbxrhY8FuSvxAhzDWUwQ
CkodEelp8a0YwBikIuExOln4kmh1P48W1eCLP+bb0/9OwhvaeSuB3o5bZPnWsY2Y2YfxHl1ACBs0
cAtbv0tiM1+Hn8FfLXTjo9pAIHkWnpDuJL/OREyLEB6Po8zcTkxtMtQnfhq9Zewm5cUee5qksEMI
zucRohqzSqdrcp7Ttk60nEZ8/vVAwPzbHQdM1Pm9faCQXTnWyaRYvkjhwdi04T9MZAu97ZdQLMTF
79IWsduYKGuAVd3SfMv3vnPCyfI3gOULwB+YYriPiMVHx6iz9CW8zNOnj7bQ7KEPh7vi43Ry/Bkk
pS8HJNhjso2ed+3K9K8R97NcWqvJMgx33Op8086Eqkol/ACrKVbWCqVgHe7lXSk+1b+fh1/owXWz
3hNeOpokWBlpFSs1CFyX6A1I90YxItmacVp4V64N49SdfacHweT569fRCzNpY5fS5FjSTWqOQY//
W51kmilbXqNAMytrWJZmnINSFTtABUzw4GwN1NtRdYUgIfJLQXAjNJOon8L03+Exls834zicxlhp
vnVzt/te68FED4jtFQma5usSx+JRqBr+4gnfSTKK+ZFKdz32t3D3J1s46EYYw5TNTDDmyBvacXLB
PQIWm3571Yqoge5ZNwtpj9c2bNO7tc/ZPIRs7M+bgHojQNSyI9RyYTFzue+FOnlZN2u6Vne97nBO
hnujMKG9Dxw/V7AUXdLDSbBOMksN6uSvZoZqu+xdiPQ3zqkRwAH9dpHFSHRHWmA6nscX7AsPflVQ
PO9C+AXzwYEB5Mx42MX259t0LOr2LuJrNSZ1gjFZ+mhT8LJOY57JBlgr8y8Yfqi/ESEmfUOv2eIv
BB8Nkdfhxend4ezNG5hyz3JNHbDJ+TgKxyxWGkqv+sMPr6qXu+CJ9Xft9PcgFMZZ0kwpP1qnqfJ2
AMRfXQSTAiFF7piNqNpYM49gBPS4by6umhFXO7zji2g0uxuws+YZ9WCZPWSpoFLFG02NJoRShhYQ
t1wKig8kbLCNCrLcczCD4rcydKXo5P5pyZYU3/CcP4PJyzY/6UhWVdgLgI/ngOcjou/RlRKHq8Ai
dQnZj1sNfjNHjLw4hYk7rIA1HDR5bRPIFc6924GsXy+0buL7VmCbJBmyhvaUkajKQ4nE0D65XLNL
w+vBZRJ4O1EnyBSEFws5ez9RyaE+UXyqQ94tRPbLsVnb5Fddo9p/biQMBd+weznseD2KcJJZGJMn
zcOuQzhS0AwZkGA6v17lHe4SXt4z+S1rH3PlY0M1usrXMdqu1Q2UTRPIf/oP5jnYSsuz2VbKZwYZ
xDCXTgHJ2VKRE3nncRBSnQjpC4HVKh6Ulp00VZlZXDxu9a3bE71j56VtMhWb88siEMfatdZlA+kQ
a6+8EvCkJINRHIALeJmUN/NM1uZInsFMKG1cxmZZnc75IcF0CLp18+Z5l1s8PonsPlFLTV46t56+
pwxr+cTPz7f+AhlN+8l/PhecHCEfocAwqB29IgJRwCiMNgNt4l6KLWw4nyvTLCDJ8DXROSYzRNCU
WYFT4DxZWo0+jDdHJhLPySpMwom8Ic3QaNpNpEPn7nRdi+JIMHBxrxT6AWo/Simw9Zbcs0lJP5q/
h4XxkI9xZek6hayQkPQthRDwqrlvP4nA0gfayU+HkrVYNUb1p9RICRtsKRHa/a8x/7un77nLy8O5
E2OzzlpWuOHgCn41/bxk6OTRatCh46EKmrsBvWkQJHPu6HJ5HDHXKIF7EHiI6Q5CSioj/g6VH2EV
EnuKK0SW/9vn+YeQqGWSdqmA2T+23mcPQ6SEFKNqxGdTWf+pRjHMZ/hwvwyZ9SBJyCDiivqoLEwO
KTGKyQnqcEXQcO1A9V7Re3ZUc8OzedzUWWSSOTCA0ubRU10ZsFGWuAeUsjL9H9djH3vTvJRhDNd/
p8lU2T44XEqg505onILjS+MF//AImXhTNhbGBwce1Z2Ihk4aIaQyvt+iUOooNxFOChysDvvNqWHd
AHYZifnwc7SLELKy/H9r5FNAIGiJq62Trtk9Oj6X+NC+rxf97pfpL8jThr2CfMpkh5PK/O7cHmY6
D40tg6T883xs0rKe2C6M4o0cpTnUYINPCWm4QLIsgwoZEghUaROszo7mQdVGyDdgItPuDYWusjv2
PbevA17WcyWg914I6H+BI8C29ttUWls0DhGccEdXfxKFxyg0EGlI+9qU6a/9D6HhOOFo0FPwam6G
h6Qh8rQsFTWlWB2XjqvCfkOD/zX3JNqbxGg30y4EcIiEp2u00wol1+kwi8Iz4C51YefPKLMjTWrS
m/F0s7Ll0+1JQbcSZQEpgdNaCcygcbAGghtfLbmby4DxgSQA31Pb1uqL51/3dJ5OxBSj1dzSoW4o
MGMSWfDPKlyumWSZwMaHeiiASAm4CBs26DoWswCca4lFyRp9IuTi7M3RSUSIQHgbrl2p1lhDX3T3
KNy8ZjRfYVmHo/GuXQxS1tGmd2PesLuuBPGSeZTqPXd5CHrEEZx5RbrG2I0/G9vmbEW0w6bTwUsD
XZHfSswablnuQpFjEnvPaDzBMMiY56gNKhgLqhG+LAYhyiq25HCO9Bjt2nxZisQpRGJg1OWprpqG
hQtzXeVH3RBFa/wI1Axid4AJ30kWDnoyAseIOK/o9tNk92yOENPbC40IPr5RTAb5YRXX+o3q2QOc
ndXJ+YuBizBWVEoNu/P4ztjBzJVmVvkzE+ZA3v+L55oBbo3jfu/xHRixa8iRhGSbhqN3d452kdUQ
xN+H7mqgcVJX1eL+LmhtUXSLdyd+982+tk1vGN1TZZ3jBjsb6oTQy6YV6K4u3p+V7UeaueNpT11W
ZLy00DxilgEP//c0JMCO4+oJEGMZJTA+HNW/luRRJEdL5QXBB6wZovE9VoXI8g9OrXUrYmgNQsO2
wTz9SV+Jhy/cC3e0pdn6w7RT8t/8dNQyXtoSEtZGG6ZSK/A4niCnSW7jSOigMd/8DYmZRk0YFI44
FeH7wILZmLX8F/k5QUi6HpQ/aYLcdd8ZIp4Mnf4OEsULLUWJZj2CfRE8q5BdTEMy3nRdIL6xO4Mg
SDJJ0M2q7tBeihdzRWLHPTgOBfvMTAC2c5KAJoKWWAUjR6U1UvUicMvwqJNig8CU/+pUgXrzp/lE
ZpDVDvaw1wp2vrcAfNSQgxIW4I+SsqVFysPWUZ1wyjvMnNqtApCCqxSVqJgFpmDErQX5TOyqCFdW
YU7UCHmuMPTFUg+fB2nGi3b92JVBhGoejPYB464IPDjE+v1J/Iaq5CqFGPwhLapcAV2cLVEBwRfG
kec+0gKnOuOYalV6Q4OvfvRmqDwUI2hz8jt78gZ//O4nrtdpZYRcqShVZGj6qxZF83AJZqlpwfCc
g4zmJLe4eM+KzMVzHhPl4Uan/vkBcWkA//nWwd0I6fVZ1sgcNte/cITrW/ZK048Bv3YWKFOa0mr5
99tKKcpjbHStfk+CPsD3egT00bHkib+aYYMpNmQLqQ2fSZJpMzqxAXdSlogqIcDv1YJqI785OAK7
g7aag0qZYpoUqjuWuHjon6A55dVee/KMfDEyWXBE/4b9BzTfUbuYqo3lS+kwR1rbnkvg8UrZZlTZ
x4XFqVF2pvRKYS6xuVIG/E5nQmtKGIl/B/AtIugxcv7LDP6lRwW+FFrDEwJt7pPfyzP/xnMg0an4
Vr7nFz1BitVbVaTPB8sUA5nGhdJdVVDhLYScUrVyncG8UNC1C2c7z2BjNFuJLSm2u349vxSet1D4
AmJ6740B4HswaXRVG2kk9DrjFwUG2CtuG6Nssj+q/BL2f7YBqNYGHqkeVbpKL/sglQag01N3nIx8
l5FJGr2K/1RUCgDOKY/cusJTY8ilnPCQByC4pnznrGYgtaXRuO2yBOC0c8eZQu+ObwE2DJrnqHX5
xGmAi8GFYpo9FzDIAL91u9LYIwGVOaDR4ztOVqmjjkpgV5BYM0gT8ozBm94MwbbMVZkShBvTnLTk
Ta2xs/js+22gv+2/fakPQzG5p/yKwDDJ5W2Ljn8v26CcFdQsU6Xp6NMNvPYxyc5K9MdF2YxIDB65
wxi6ez9FIS9uIorVmpqBZ+vwA06EvPy1FlxjJVyF0uzxtUm3mT+u3LyzxZc/OxbHE2ZRpMLNp+2M
Xl0lbOl6JD6gQUY315y6YNTGCIvpeinyYP9WoLO5NdA+k8wcmufb1y89W1LMjUySJkkp/0dp6EUC
EASH8wt9xeTLnRYK/SxZnx4qA+u7kZPe7zOdFxhPiYxEHqujIKOiBmZWCmdJeu/wX3A50I4Bn7wH
l13Oq0pALbuIR5g4xWRyCoYpfCxkDL0xlOQ5Bwh56p40WcG5swqx13gHldtYHagbtIIyfUsQSk2e
YfYUjabw4RXeFyc6RIyviThbpWCs9MY6IvVKfJiYhF0ZmvK5XXFD8ngEvrjidmP9FjekOC/Ihbt6
8xLrNvxEdSAzRduBtn0ZsIG9fLK2wSU3OEd0cZ//Z3jw9ovt4XdGi9RXTpz+bZu8k4efpZnUcgCi
HMoQnhN/PDeQMptA6Q61dip3IHXoLo2Q9+O5RoJXBtqXS1i4KzLVpSwsZfWwgNJU9ItZSAa3a0sD
rMpYJlHaJYQ4tNl1Vn+b7efpltT8Sc8bmGy9fVEIgzda1HFpvoVDmANpRkrvj+FYJ+J7HSzdffEQ
bplknCsB0yE4LLBq4z6cqz2RWsnBTdIiT3SAwzTZA4JTWQ+TMTEqDT8nusjxCs2U0ABnWiV8UJcG
YlFPfRTinN9CxntNO2tBdNIqEDZwDgxAKxBkB0ngNDlAYO96b4mn9fDhpUPleA+9FS5VZfKaK21p
an9/NG23IgPiDzfV15nTCbwXa58la3xhWk7gAMrCoaHC8egMbMgqyuGUTmrgDjbyrfjbPwElEt4z
+3ZgJ8V5PM8YvQtnPMVGqUZTJCRgrcJ4UmpQZFQA+MPYe0ks9DKmGmJILy+y78ERO7vK1Nmh/3jx
Pr3kKaSqwVjFmW4UlQmgvxaI1eAqw8RZyTVIbRlvZZVfmVLCeC5ERYOCpj/qR7LmSZAswgcd9fvk
rGF42jA4LVlMqJiiz+yRQKwaJDBL3EQAcV9/GzfJFst/3DShJIIoHDajeKteoPtFHQzIZ25SUx6G
Q5tvscHtDtD/LAfhmcYebDf9LchL4LZe+ip1Ddr1BhNArFCFt3zdSaZmfWgvIo/tISrdLuSsZ/kL
6iyNYbBFi1Q9IVFSa2vAXHQIFTcsKe+FQGet4O7A9S1K2dta30ac0mRhD4F/AwlY160QX50wG6I3
1GMnq6T0SsgsVj32+bfaFS6311kpkM/KjVttq7evlaeY3J9D59YRh7lUpMK7iyjENaKMx9nq2lCA
q2o8sWbeiHsZdFxK/wgJeCdfpbjgaAfDcUVhiEdt6NdjEWRXvdaOdRsQOZVnr05dBOF9skvCfOe0
ysXx/qPRIZIatoULcbtedkpOd3hF6ErWhY7lYUIypZLhiMZRpCpBjHwkJ/2dhsnseX+2QHvKoOD8
Sba+vTCN31iiLeHemobZUrxk7oE+46mlqc5+d+kccgAWBIziNrTnmTq2v6K1AMyQryQlONf0wPOH
YL9AOKKlxLxreaJsduPzhDNHV+YHfBz+Q/YUIjl6TQoI61Y8DAUzQztDlP+62w8Cdqz+WRfDiguq
V5tpom9Q0J3zaIH63MpZrcdHz5vDuGjcB6PB8shNm6t+5Or1hJvJiA3FwWrn3CnlMTmBA39VpBxL
EvR5Sn3EBls/5zbEDnldKX+KwFdYjJ+yWvyYgFPPAiI8Vg7hIKkw0Nng0J6g9me5qMh+54egUROn
YYOqCq8l2nmhkVsuHAsysyL12N8kLfPwJ/ssJpbcch4J0yPX0gxLEO6gxMlC5gpIHkCrWfrdX2jl
esz71Is1Vq4MEwP1Yzx3OQMm8M/+3PQzTmHEH0M4K/Qd8ebp1gELkbq/Mw662uF/sf0d/ApPvz42
sGg2DCzsHP3mmDU037W/KTApXH6jDzZ2QvIE6jbOnoJ/bucGJtKzvutod4Dupi/LxPn4xxGlaVVp
puoAx9NstvIxIg8XE/tj/Usxw8l6y3/AhakF8ru3RCB8SPzgsWKSCspgJEdu8cnv6tVJjbwmRj0P
8C0ZVgDh02FicjCdqjahGfPmMEBXMb7EjAo+doyvb5BTP6pjde/xeKFyCJlKooSofRDBuSyczN+C
PiOJlul2vmG6/hDXLiNCcI9OK5FjCQn8sg+g2PP5grB2hKFUg3BdIksvIwe2afJAf29wqv6caZc8
nSThGqfZj0cKo+OXTalbT/aWRyQ91fP/IJl7ttTHgXTryKNTu32MEO/SDqfiigK9feSF6qiP6bVB
EMURyJfQJ0NxhZTHCLK+cPwCboJ/OYQNaJViy9Ss/ClgIr5x1TcZL9YrXEOtrQc9r4oaJkqZa2mD
Jdxr3pym3Km0e1nFyfyNIS33mSThWfMoD35IkIkKf3+fvl+q6SQ4eH4U6zYzUbdpfZNo8c1gRRhm
Z2ECJWF31UMfAibvLGz+ymcVr0t5AZe4C3E1eqChCz37jNUWvv3scAvPcFp6dkwRAKxy9MO4NFUC
izQd4nFKDbj7Qlb3hsTfYGaQn91TX7wuoBHySbT20h/ipO/NpcDVwphIjSF/+Rm0m7B6uAYW1YYQ
TPqG53a9oobdBsPCCohA1SZZVWEOnBzupIgBYx+1K1ytu91FnY1UDnqLRbPit96M6neUwu52w/KW
6QXelqtt/KYjGFztGXpigTeVhZJa3dL1ixX/gPZGPcJhjSlXDzmhkwWx0Y1mJ/OOXnBt8G2UM2Cu
XZGFhhvZv/TQzvUzKCfLrUS2DIgmp5Ye69yBNAI9rwdpCZ4POoCaSQwv8UekTrJ5h1TksAHeSl3d
6mDL8cwnfvK/94uo4ZSWk/PP7Ry2YX7W3Au9tfpwH8N2pv4kHmgjYnt5bf9hpVA1+zxUGSqdhe6S
czjMbTjvhRtfEUBUTZSd3/vPQLrzwBneGna1UXtjqawOeMrRMlMpjPmWErbNdljxlIYF0x+O8IZo
mu9kaGEpXPLPpYZDgROOwDcBKxxmYCk1OF7uPbqaQ+RunNqYXAcu7I+vd81T5GdmubKUTnVVMAe+
PL2uk3EDQAUuIwYMHIurEfSuricfY9iDIpFtZ4Bbjrkts1HWM95gEYSPQmfPQnHhQAltJI/K8YTB
lIiuWz7tQQu/aHLjyofWP7dFelCUcKfz1jv/53H+/vLdNqJx8S9pAopeenkFnFM3ZREYFrfKg5Oy
cWUl87OYdLZknHuX0ttJXdl5SQl+gP3BxwS4Naj/GIML3K1o+ZEx+lBEjggVPlo6bPNOJ6Zait1H
CX24IsF+IqvS/mc72pHU+AjO5ZULeWg3cJgPylUBfLj7z4q2qWKa0wNLd6q7np1rmSp6w4YyIviW
Y6klly4Vg2QS80mu6trIuoEi8JN2CaTUvue5ov52uU4GrpZPtJfEuJCLMu/wTKPq8C/73kGnoEbj
qAxYQvTFxGrp152EZjZ4Sgh6LJjT4W6Qb5zhymVPHRgNvwBbXyXbcpDWWBFoqLdlTTMJtv45U/HA
gu/V2UHA3Pfn13xjezOmLIcKrfz2QoTrAwoaTrxUMZ8WwOC+CARWc4adFQ0LblsHp0fUC9tE7Poq
kkMiDy4EubI/16hdPRt2oGpLJWg2IXUBBqhM7QuYZ2qbYUqdt9vLmdPhp0M696twRC0B0YNzX1fK
okIh8XAYIPGKNhElIMXX8sdDa6X25dsYfu5NY0wCu4SL2NScsI50x3KdvxORnG73K51vCLdMa10F
MjcKaAsD9lM1w+LSthZTh/OkuQ0J0ZHPFb6YeDxIHvwOS0uG7F0vILRNufboKrer7oUx8VaDkPz0
C0bdut3anr79HdErcjgQk9YuHHOcIQGe/4PYVubI8bNBS8+syTdJHvhFLKm6Mfcgb3YijbNgy7nr
6chs7iWyTnt5LnJBic/LYhau/Fc0gyvfkxdePyXF87BAOQmH6uIRMQ7C7tBxglVU0KKrexiG3ZHH
S2ni7OYZfRDKTTi7fsLC2AHzgZQJhHIzvUtsZLVuXyfDe7zJLgY6ih4YTgL7XAEpCf4hhZc+1kS5
iByIBnEKYSXNgIE5h7G2U6YbZdygANpsvI6PHXgXvR7SVlqg90ZfEbXjWUR2jTWxZa+6dO1ugxzy
/poUBnewbRYg1ZYkW5kJkWWAsPQ3a86yvphvHaXvaYvV0+v93fxkzJ5d526L3rpaHjckzmtZPz9J
nh/rch3uhKkKf8SzuIZ0HXlxNwAH49azjz+bT04BO4nu3HQREZ7xsZYZwGZ0w9tJTO0R9ZKis97A
yeQ95rZoWo9oy1GqMpI0AiAEz0HeuzIq4OxHY3kf14DDlp16eTBJOxJCD1Hf+LOHDqR7AaXNg2mv
4mEefC0JqYRM/OEYp1A+V6cVXV8gSgK+3qSiksoTHh9gtUx2AcrpURyP6pt6tCXHgwzJnIUSq/+p
ZYMlnaT3zRop8ye9ZWAAUcPUnW1NeKH2+HOtqhCP1iSJ5Qp8ivpHKyiapy8YSz5ynzCsugz7N1Vc
MPY6btWzACBMzFFwjYp2eMJFOzVu8+krDQ96++CdLJbvy52T117Eu6olF/D7xONmxrMpD1aeSDQu
LFE/0xviG6xqpX5aI5ADDLquK1eGd8qyOM4pi2gg4rFOwvgg2xY2hzjq70l9GAnvBi8IamSptDH8
k6Mv3EPjNdz74d0cLzMBMZSmyVFsTkK/Bm/Urnn6uyK90IGtmwJ34++6nA3hqnCyAzArd7HvJpxe
pblnLxEnDPUhkUuyTw4vpCOQXZMaIMEMUWNUMv4PkRey9HOtiggM5onCtCRjXk9TgPQErWihsEND
4xzSwVOL/NFdjyYGGsATe4bqKavUmoDBsrAjITpUmHBIwEa8zLdxRT9FCICSdXFg0GANWcYwI0e6
8aB+almSUO4z0jwJOidqcPSsW1EMbMtpfNIfSq3qUVJTciod32tq5arf1Kdg8ME39g6zh2LNcVV0
z7ziDQ9Vu1MKHlw5N0e0ZsTmEdCOeSC0udfisaEA5UM3KdS08XVLqVTwZce6uEn0AKLXTnxYYia9
ja69dpj77wc9Ui5KUVaya/knCOUke/Ju67rlMMFR1dnJmMKgVC1j8p0WcF0SfGQYb2cCFTZRbYq7
u7PEPdHrzLICS/iuzk/clN4GTg0yrf1u7F8YIbykN9EXDr50X1YVXRl8Yd58xHyM4sl3uU1MoWML
rMVtrLvxalTPc+AXlQEZv9f4gZN4Jd79RLAAhyX4NHmgKwHBQiAu9+JRm2DLQBZ88WZ8ttpUPe+q
zNO2jlHNV/Q7URGa0jC2XxCtAyR9Mc7BQzBR4ng2AtKgym8ChKEtgagrwwoAaVToQnZvvTROWl4Y
Siw3aXJ7TPB+nkxLnIfgHk1T+4PhvIYmsGcaeAjBGw0DcomlcLgcOjzEMyUU2kzFum3HpCbhoHth
yifG3U7WUGtSsKokbDQ6fyf7Lm14+Fepk2notrr+YPkK9E8/TmP0ClqNbl4Nub+aNzlGmZqXLd6U
Mzp2IRn4O+l8hogpW0lQ0cX7iB9u9RvBawA1B9FISpybNd1Y4pdAjWc5sQkR1CCtHAf5fWaFF7v9
RGu7IUU1JY8B/oIYxiLj0qCi/sjlMlsU31F4esLA3a9hFcFH7W9+iYshfEA2azApMtYcVtw6+0zB
rTDKzTNjb5pAv1weigPs8+wEgxjAVq56RlwMTM4gDyVODbyVQVDooAMWINuWyA9kH2+rrzxyqS9/
xecQtzCHcxowzY2WoMPk2FpEW6wb2Scgo6SHLzBR9IHbHMUFP//fzZ9JmogUNvqwkqeh9+YRWXMe
0VuqBgqSBUNLr+8dNrVMcyLcxddkgq8MYCbtD1NMRXcOefyI+u2hwcglJ5gKdhVG+9BCo6s6HW2g
FLDKiqX+AaaXkkT5B+Pc+fi1dYvvubdZYQfIllPZUa4GW34CzBLbbpUo0seRKav2s3NY8DnP9FN9
g1Fi9eFNap8caf9dy8mb5uOU1dQTDdHEW3OFwmjG3oeVD6YpHbDI87lmeuMhl64q7SC+S9BhmUnS
Rfn3wV7HQKha0ZKySmTqEgbTkSQXoSvAiumz42Qh2LXM0M778IDSBhHOxkTvHU3iQr1A3x6JLn+6
tC21RzxCrMnJ0rrr4QEuTuwXklIdWEhcKR6plx3/Jz419cyRd1HVRJ6ZTFCvksoQO2p3jS3K8RlZ
I1EDYQq06QCv+5z0a/oiDXq1f8LtehwDZcvVDKq4paBitt62cEtuGEEpr6OcG5TIuV143fiQZVZ/
VdC1cP1QB/vDV/n9IJic9FkyZYvvMPW2EcIRAPzo2G6OogR66TE3ALkDWYVWEWQCLRHHzL+SmsAJ
J6C79ISCNEph0a7EFWLFJdVaGRlR+YOm+2oRjGo55BbD82yypvDhIN9l3Wqq74co9W55XCzmVjqq
bhm4OZd+TWgEELfhUnUqVkwWzjQ9Udh9eBb3a++y8bt0jqMUE3vOE/qesROl6t8HxVoEKkhxvDRg
h2C7LQSNzvkQhochEFWrtVXZCWLfa81D86pdwCk27STP3XvLH12EEoXlK0LiNaWVgzjAZfG8oCh/
GVTVnlM5GcoQvUWjLN3KAJWw0wuJRZOOXY04Q2vwfPpGZF7+RfCMLpnwnN9PPWGaQOjhc1A6vSwC
xpG8lgJIPmNxauGkqVWu0ilHzOSwQoGYiucYHVCFAqRaDio+/Sp+WgG6f9/bTsrKWwnyZlf1sOdu
kTgZ3mFntlMI1cWHWq4lw+95L9o5CaoTnqOTOmViN77IIRbcn7CBrpaDCy7w7oeJVb4zXQ3J6qrZ
g2HGCbE8WU/OudxekpCkjxShgDnxAk1SqaOo4+e9qCTmyYws7DQsO7C9uOo63pudDTrSm/SGf9An
K6NstfkUBTv+vXOwLPBojjJGLPrTjHaAmtgVh80LtNkyHsuksVfPcgFGLiYv7jNVnPZDqv257IaU
Bm9O5VNPvphNNESPP8yBmM9u/pAxqioTxdP6Kgk/JRKWgokEHsexSc5AmIU/wtN/QXohwRumB5oT
ucLWKWlJT8TwUwWy/ubS/zqZpe/x0Ko3a87KE3zoRiTU2zfsHZ3ctpUvA/CsK/FKiGrg5QvwXMwJ
TOEZzCX6IWIq0IQA0vsKvduXjOx1jpqJAQRtuEVdRk9Qjqw5fkQylTCnQJkwppznJ+ge0bXvKg41
RfjRNC1v69j9hrWkisBRTVBQJe44vVP/yGQtuCPOKYQVW8jJLQvkUMvPTimmcmxjPil3W3kfrjrY
zCkLBQwJ0Wkl4GqAxaODvY5kRo839rHG0cWX3xZvGbWIW/YW8PBPNEXGE6+GLq2IV71lz1t/Ew4k
WE7z1NfQj/glFh7YJSfsldh4Oej7xDNIlXIl8qi7PwKELq+zJiCJxm0xsyi7Hp5UAWjEhrNo4sda
d7HKhTOgkbAMbh+YLIA9tz2jAJcuVtPVbH9l/8Pjp9TNlXsXdIrTTx1qaEOlN8K13UxPK947TuKQ
ZuGgfq7h7sLwBbaOLiRSLOWbyGJifo8JOb+z/lyOPgLpItc8OnHqlQTfcXenB7ZrZvW6/m9Ee7vR
bjdK+NV5urn4sLR4Gm683zri5mNr7867N0xYhkk5nT3MsoyV3UTtbSRdN4XUFeKlEqOXjBU4w1uK
Lh+te2TELlUuDU/T8ZmBOljtGG9WXdb/mCYZy79/cmVP/BWqrCDwIFX3aruaS5jNCm36++aI0Fod
rw8F2piyIO/MA6ZwqRLHLpyyH/XcxDG9FZOGqe7b3YU5LS6XRvWG/K0YFArDjzJN9J2/VE7caVY+
zIPwEuU7yHzDfgO92QMIwTISzB49mlMaUYQIl7+RBpj43qAv4Na/a+wX7T9AsDvDiGZ0QdfRdgdt
4SDnYD00+/kTIISf+MPCKioi1z+cAJUDIO11jPJbau5RgXZzqMuwgUn/TrBgPi7mIAAekFFsFeFb
UZFG6kaJ+pAyG9NjwTOLUIdOzh8e6zeJIe/EN5dWAVX+ItfKb5N08n7JGcCwqIMX/edmI3Pw9hfk
7Q4UIWzlzFK3Tm6nDBaBs+ZOXV4s+/yTmKzYRMQrTHtwLEKKLui5Qje6hmWeEZ4PZEKaeiwd630N
tlu08CYgZl13vD3uhegMwuqwNW3c2h+u7JZ5/Cyy0Us1n43kxpHVS7G4s8MAygtpFhkoeBlSG6Ya
tA9ssvi5guzHvt2xYKRO2jJASlE7XGi4Cn1ww8RnlwopB/nZ2XoVg6qVcKl2f8Y2dHiuMaPL1bz9
7pZ7rzJi6t+AOI34t1+E1S9SXmHqWt6Z0BRlla5edgq2Ne9ELhCLId31ULVTJBVHXWdBUL7xVF+M
gjpm75G8aZXocA+1UJcmGddqeGT5+MWS1dV+9H2dJ1Ix1vH761zTRA/RPPTM3oo3sgidG8yUqy+N
E8quer/RGn+JBZEG9OkPA41KxcpTb+VHY0RRe7vZ5Yswc/HFFNaldcV+/6eIY6nMyc7wU3oRpZit
18yQOF9DRc/UwoLm5OwnnCoh91tvaB3GBFFDbhO0xTQ+imalQOH15I3RGlojnIjB4oz+QZmS8LJB
iBf6YmYcJ9lpmooHmQS2r2T68wXI71J59QS0TlGH9BB+AFxaRv89TSIIoTvFVLbS/qss5gbaUu64
KrVI++w4ej/nC854FLe42zmwXB6OPsqee4a9cW8JhuVm6yUOoDurXERcEBEJKPsuFshrFKi3qfsB
52u1UUUE/wxlUlY4IAYu9X1Lu7dnm1GagPT5M8WRdL0gJ9M8jXmERyssz7qw8sNq6lnnrFZVDHYX
pG855JY6MH5rws/XlBal7ChvF9R48wlL+89eUJcgq//xVYInwddbTXiNLjIJjyieP61RHDwR1Zij
JFggWjTJTCv1NKKuChdnxAmyozMC0FGMtqLK93CPlWf2jZE63gccq6ufBcGzHGh5cT8130MfmPwW
WItswSBT5ohJwPMfNn8V7pa2h8uqTu3vglpZVd8ZIcL2k+gncbV2cTpPZ6ASEaO/IJuYtYjeNNb7
2LCLlsnZKkC272F+sDFJF0L7/VKZBkiM9i3MZL4DBtzYDRc4PUKnLOz228EJo/xi0a4ASXZiDpia
VXYLNwyER4BjuP/UZ5CfIdsY/X6ZSopYMY/YNu2nTJBuubG2Ds58G/e16moALqmrIBnBhLYHGd73
bia/FWaDObQHEAgD0OoMEeqTMucTkvJltUvYpLyMPCAb4v8gJ3DVhjSYnb0XMRmw7ptIQ705wRHJ
LJOBdK3zKc72OsK3FouYUiYxNEfkylz8TpVYbixoTii6XywDMVwO76vw4JjLNOY2fZoXmM8yrn2A
J31EWmYPSA9pBwSO62PwAouX9zqq5DhK884TLZb47+2wHF2Mul2Hf2vN04daNdv+Ux0w67ARsBCw
k1olJfwuHQiJwyDMRvPkp5roxv9XkU80qf7uWuWxBrTzeIHZ1rFhmlV1oHWJywH/oQ96wriqpBlQ
wzyw+3mcxL+6Z/8OQQsoyugI4ZLmx+yfdsbfTq2W3MrhtiQolNkR/kK2GUxZqugCwrqPNBulxdYO
YeLp0UjAQQNofqNBaz4XU/MEzJO0CGQ9Oc1+8ZfRg0R1DUezPvoRTAqH+NCaM3l81V7JoIGV2wwv
beQGnaGgitBxyiNtvhzuEoio9Lqp4/PTfhbBnttdkntS4d5MY9B/uo2eVBZYaJhGhjR7T2GCTfyb
EKMBcfq0oyP7F7qHjNSsGQDN8WwZSae0JgQ+jkJLFm5IkYTTcpgOofXcOxtqsVTdFaJRjEUrmQtU
lWUkeKpL4Q+b/+3PObXCYjlZrX8LLTTklOaeJkWGBh7gne1G7849hbuKMT6ip16LXE3czlSXFPOM
F0ol04kuSm8nbWzfan5oOS/mE5hJ4YMQBdoq3Ox8ZgrYgg8tUuC6rstVlOG7IYmXOPmvDXAw1PnR
GvtmTfQr1WtgcZ4RDseazc4eteFOfa+Squ4nNCxqN+1NMDafu8uyYrOuOjFO9mKHpUriA1VTZ2FP
BHcIm1OTQnw2W4g6KLoY6/mRhKpVN8XYOwf/wTtTHmWiinMAOAlGkLQ393pjRLwrRxJ0qZQKaX32
2XqyZK+Df9ivp1PZHm/jqNUSDHUzNIWqTnyMdoHz5u34BWlmml8EZUodeOik69zFoiW1U7btcJ6h
zUvPsm4zAbT/54N0btVf7jejlUPeow3DqJ33VjJQlApyLt0bbhtY8be67UNwueFX4fcc1SAmppjQ
MICMzWjFfi4lo0pHmewkAVUfdWlqorHpYvFcUV4HxHyoEJhAb5ddNJNRgffL1nKrIp6jCpTQAyGq
Kq6ut7xY9ZFlN65BB+k3KDl0emKQNlMbKAOQewdHwNUjTDtJ+Aeo6Tz9b4BAxCuZt5mzyQm5EIMB
a42VEvlqOCwhsF8Z6sW6yFLBqJRXk07gi8nPEjt/q0Q2eN7/fj27h7ykuo8wyH8SbmXakD7rGBrY
fR/VarjdiwwYjtAn4vWarjH3h+bILZY77VdRCJ6s9u8B0dpjVP7me5gk9piT8lFhZMLVsRAiVVPw
uS25ChoYFN/Lnpypj3gmv+YzoVvd2TblXtpzfWSVgh955kMJhUIFnLg94Rpxp7jWIgVvxwUxzcoX
paY0iVu4MdPCqsJGiVF/7Im0UCaWVlzjAalKttArfWgjY0hW3zXXvt2WXI/HHvs9h623y5SEbCiu
KxpmVRq2YbUOmXED1tFgvQMh+rIpQKEeSW11BA11CLPV+DiA8/psfe3LEXBQRldM8bqNIIxlhYgG
B5kpM0QFGp4qY4y/h9HwJtSLVtiHOubVVZ7yrmr0kjkf5OhDBmJMg4N+yUQD0PNohnLQzQ4xIoTC
iYsqCXvaWX8HfhxGOa7VJ7lvv/V9/KmnTGZaAS8tJ4auVcmRJcu9STsEM7Bp13G7WsnpJJbTV58d
ZaXE+BKHLDvNHp167IpftrR1x7qaM4BuqfcoJfufHejAEOPbDXvt/9DWiT2SP/zHD3JGlzBn/iQy
W7y6ISMgcCEadrbSApdM1lPa+jnBjtzt7+jCjqNtdeixSXnw7pGUQlM0SvmD2YQauymHOpSyOrPt
G4AMrx2zntGEnpPQha+QwocmFv+NeENNGj1DpCVBHjJzgDgpEq43WqEWG4uho2s58rrkwD01Dv0U
eRoLw7elnoMQohrBwFwa7ZV1SCT0ZIykj8QFlW4KZtr90LwXzMvjZU+Ti7fMDxoauvS3hl59jS6B
XDPdDpVjms9ZNBpd2rQLjGM0WO+N37zMzruVMyVEar5zeqqv2gidjJ7iNk45qBD+7WXXu2fHfxZT
JkVdb869c9Zq2e8e1P69U/ls+xAyV8q5DuE+0Ctw6bS5Bh3VO9kPShU3u/NJyH0hLaGeDrs2UBB+
P5sKzEXdLPfjZd6Eqo7T2UdI401a/CcT53ggcaxjbQZ9OUdX8uPjGm3v6hMfqeyv1L5Ms5nxXFbM
l7xmTtRjvD/PO9G9qPgUnWVcY+cpe/LXleLaQfrIHznN7HGmg/JddTH4PqmAuQGG/3vqrwc6EzKg
i20UTKcEmkLwiBLJq9P6cyWmgp2+CfNsTZu+oEawZ4JgY5Ql1TSr+yu6vlMOpAQcb/3WnryTLe1L
Sjn2KUQG+LsWQx69QzzDGxtC+DraacJ5emn/y8q8oMdlZLMX4nzxrp64fjID7nP2W+zK/XzTuoyH
GNev9kfIi5ynOACq9fzgGLrDAPPLChmZRW/YCRyV295AFo9zuoqIdlL91Vt40WGwzSio+p3VWAPN
kmLqdnqsYdDllcWiCqXSM9rC4j1tyBu9Kd+xIyzvGMq7RXOgspfNs7rH26Y3+RPB51rtXXpuOZtn
1nev2RT/S5dCixUUagvuI+/3HYeZL317I/gVe5yGU1U5wOC3LVL8lr7wFNmhdfohMhTPIotEvspb
Dz73MTmt7JTST2DfTnCEN6+7sGuSBIg6Z75BteOnPvh4jAyDUlgnmnOm7ld2frEiJkXhaaK6tKk3
40DR+oZrTZamFz7iploL2Yk2aBd6ACd3GPRruU2/qQ8d0KB8g4CkoQe+vQ/689AB46hksK1xhD+N
F4gM7iZ8NFGgM+RhAmJDkXwcm7W/Zotgq6ZlMXGf9zB0idhbseyDp+W74rd2nMBIMpHfY9lk77/f
NCxB8aZ6Svw0ama/TTQvPR9hPW/+VvZw2S48H+LJPuhgWtJIwyj29IIoCKQJhrgcf1pWGUYah1tM
Z0K6M3k2ar+B0g5q7K6TW2WnrebokHkQhOnrdNrqB/QTlUwRYPw9KHfGVywWn6fOLR/DgdL2zp2O
UKsNElJIDGtoxQo/3oQ0IFtfFz4ypWQ64v7WXM4ctrtZfbNIPlO0Rkq50La9hHJHvCq53SpLXay0
A16xVKNd64H/7GvF7BIKkuEAG2NDdrTlAs1hN1GOov/SVP1E8DFtns+tad944TRSFJv6RiRHkwMy
tsf61jnMW1cXudqTJdytlwqJRArPagbrjD/fIvabzEBToJM0d5EXeaJXRylMLt9d7PdO7l475dKP
qx87fkUeRvY5Ah04ln2jz0MDtuTd70iB9Xy7fXOaVHxXcvSWPQE9WAniUSdzUwHXiIR8roZnijSe
C71zHhEs5f1tYHrpHIqb60yn6kGxHtA4xe9Wv3gFldahFY4F2H9XsRJ4yPm2YsOkIueZq9yGEc99
5rr/RHb1fDFOHXm4ICjIXjiBXZsKBCdZmglGgoCOrFnIsCIwWG31s5kBBiXtV+FjcEzVgYLA/UYK
ByPl8CO3BowLmDUIoXaY0KnEpWjP4W9m00StshDk0jaHpkffJ+a/SGuh/5UfkQJHE7yiaJllk1zl
Oeqa9YVIeYcqjyggNbztfUhtaKKL8cmOJvR6wJc7VfpCmMTLUfV2EbBm6UlDumS5gyaV1Ptc81sQ
lgzTmZd3cepVCHjEz6P3yj0rA+eKrls1hKEkkFq00lyaNUTcJIXhk0cbLsbdqSwMcS1zAUJkbayi
TpLyH+W4nPwObRgEBZB9uyo8Ak780KlOU+w9PORrKNUkzVTGxhkrci4JZewv8vG3rbhuQskZxdzg
Ut+yIoTzJhvjL/OClqJcScnxoXURC4rCEarBtYnenlYTP9/ML3f4Ax3HPxnFpxptyhXfud067jwb
NpdMlrtFuGGdSszNEc7CpWXFvW2vq9bgpqwxIgaERDZQZDtgrQTARxJRw46CNk8XX+krRTIwN1BV
zmO3+W5Gv24LoWkzjuQaPWzpdpou0sP/VEytmnGOucCCTqbxN3VIQk1vxQbsZcEYjZyHjBq3Mavi
FU6bUsT19IWOosSgl2LIKa09Oxq3TlJsn/Mw6Ovi7CVYiz0OgZh77dHbRRa5IkjIL+xi+MIAKG7I
vQ0etyN0oY6U3rp5TQ/TLsqFHonA6VPajt3PNDPt/3shLgNnXexKWYYhgQn0VIOJAgtX3NGGwvmy
fN+yW95MU3omF66kQj/v7PmtzP11mrvk4TRqyTKA85XWTJYq583lnExNArN0ftj7t4D+P82EYvKH
/hWANdd0S2qnIjEcqH3lx3XeWs4CK5MbCqnfymsTkZzgwfiKjb/fHwAG2Ru6xK3Ya8OBlotMWr4r
BEL+yHTMKhvHdxczLF8LmP9Q2Hc9s3Cwq25k3j40CjfOEaX+QyfOCUkUnGZflsOOWEITpLDh8vSR
gTUyshayvAXv2Z6YNhqeckNROZsKrf0TjjEC+tHr4m5Y9xRoHg9yWWju3dtHrOoQWwf97+noh2Y7
nQ3b02/l9MleOAXw4xK4w8E74Xb9lBk5LLfjkqOu3Os6iuo4UvU81aXhjOZ6ol67xNK5BGtgJ/nK
kqJtJp+xj3uo9x3fMe1e9DE3sOs6QpD6B0+NluSe0d9aquW1p5S8f37HQterSarVEtUHrLyzp5c0
3tBBiLMJo8I55H6CFPzy57MrfNqzlQog0XnmsdIZrG96W8EDIlft4GYlMbrNibZ1JCfLG68pt3Gv
n8UJTn0nEbfVTxtf4oXYVgC6H3cujiuJv/VRMfZrSkwY3ggmxwdLcyOByAdjP2r8bSGUvUrG47Kv
kc3tUtZuu9TJd5W8HEN3q9ZqsX+TTetLtCPGL5vVgDkmlaJT+21YFME5EHwLt7VmkdZp/8Cw55lh
CR8ZPW0yXnjkQSMXPkoF4magI9xtwPh0LPiaoK8UXXb7aac+RcMUINLTgRe3fl0gkUVrrHYeK9Mk
o62tvTkhBtjJhpz5ONAeAH5/HK8sAy8K18qViPngQhjbGNi0QFf9zmAhpfVLtLOn+yrAFEpmDRtT
E0G7KTkfXbF/+jT1qp+9poN30m6IbGxxm2tMYI7h78LkeVmsfrjS2ZfG2qm+V4bGwHEtD56LjFyF
C/yMQC06nJTdvllgHr1ENd4Owvvz0Ws+LSxPoAOPoNO5CequDMpLsgw4ZaOqiE/tdggaShan9v8P
S0en3xAgcVAc+G+KRUCaNVMCJ42VPXXWIjacHVZKSY57fLttcYsjGirouhAp8S89lPKzZgKnbyDB
9Tyfyg3Oq45G8Q5IMDE75UH3cHS4z5XvgOU8rGy5JbJ6qbCMMWxL/8KZ+Z0zm7emNp0/9C9rQot0
ihOTbXbnk2oHAYL8ZFWpDcxeC8ei1W6NEZ8kadXsnFfkPcA35gdW3A21HM9TmVAPf1jE87YAVfWv
bfDX+SAI+b/RmHPim5i5BwLUVIQ1OHMZCh7lcY/dxaqUH9Nm3/Eb8ouEsE9f3pD6ga+hratO1mTT
4GEN5ZdZhP/AelARPVUs/mAlvd0nXjR7RFGhMONhbGwbl6T4S0PdyQSGKcGLnJYJlrqdp16xxMrQ
7X5p9zYXgHkEwqNHqWCgtSIA5tJAzXU7IL3Hn5gMdo6+7+jCNyQ5GWroWevJzM5heQUF/tvHZSey
LVOVD9lWpNBYz9TdDmQsMfYajQCtnX5voC4OlQJG8jfZl+0MJbc0KF0QAbNSiYq2xo72SaRodV+4
79kdT6MND2jAsKPpoUBF07sO6MiVCPDLM2AZ62Vx2wHoqfs9qFsFMDsqhahj2ImTHy5CzKHMx08a
QcFaNHMu6hThV7vtschQd0qP1rtfTgIJ+KE1iYTPlf5CevKDOE+ivKm6M9gySiYy9rfX0Pqr1TNF
PqUuZbrAyInsi+w194kNUQHImmXd0WHesDmLnpbXpjq3ImzQmcEmDgsDQ1PclglX+WN7hloy9ptF
pnfb6GVVBpLFQR5wS3CRxaSVuhgqWia0Jr8cRTnB+UACRLjoh4/ON0UoRWHGGzgFw1Bc/pmpRZgm
RhLCF/mijRtivQ6VjQxgPXJSYQ5VEpKydDQZZ1k/3pkcc7ZIFuurmm5ea4W7b4z1yfSQ7k9xRKZ9
guAk+5sbyBuc7Xj2CgdfZoJxWKN/Fs/fBsoC9WMaptE12AjnHKJwAzJuRNmONNSlBGduXBzbybbc
fuE+7M5eFravqwIoptlMKGRLUIxqlEhaz7t2XV4B90a4f0AN940zRyAG2XUHYAE8iyx9UBhpG8nF
NO6tn0wCyDpFK1LkSGuH9uYBlNgRcsM1CRnB3WTPuobxmRgAJA0Gos3pGJqxVDQ+gNtfhiIWUVER
v1lp7rvW0w1/UfH6e5VOkCKvWykoOOIpNvB6WNwzlC82Xc4iq6ukj6i3CVzivkNgZHEpljP5WR4Y
oWLapCFB3wHJvdcQAWNrgAmuMxpgOdnctFvzorGQbzvJcO9QNUVlpvEvjj3URSewIABY3WoGQI1x
BmAfuSJxMGaDdl0bPvJKgkH2NsYxgntwVDVjUdXiFuIL8OXYBKifNj7nhCA+kerX66V9sji9dYsC
aZh9y24VT7mfd0Req2oMjFnsiVwdhzu1TOn/d4auS0R16p1wI0+dKLyyhtXk1b0Da13xGw9rBlir
YB+gJ8Nc6qt/dQ0cmAOuPNK/c0khzyDaqVtbbwcdxy15IsA8ME6oOP4rVFkAPE4FmJpsqWaKZFaR
70evSpWTaRR7D6ykq/VO+98WyO75cbH2hdfJdpTdThcgQGexR72WY9ohKrnimNek1xdExlwvZFoQ
dHJOxGd+h38B/1nOF/LmtEmykfDKT51HM8n8wEqTkjXdDH+StxtzgMlvx/zoTRlw4MObqjsqk2DW
7TrgCTuQThUUbGSKBUE491L1uttGavQEFKx/YzHR8f8uXqItpo4RtCZpyDK6Wkxm1eOBv88CeFca
LGVsSgEmMiIU1f6l02cUU4iWIvIRvV0iUj1ETMwx0E99FPX155YyZ1/ulWtlokz+wGI5Y+IUPT+z
SM7/+DHRSv5upSkPz8vkn/1BaW5Xz1u/wsA/gT2+ZMi3IL4QoARFwONhij4MicFvvSqhHPucsvpP
o/8UoXoGNYTnd5XsCDxfXBuUMBiUykUZAOrybOFwZVpqbNNhNELH9AHbfDSSyU4tqlDgodSMosmt
f7XsqEzlTus8bPvmBuUlhJNRG9XTW62gYLZyba6diyc2pVoFZhMKNzSa6HdwgX8Amtxjf+FAOnR2
Bh6p7NAtYz3A5qNdnOS9x3Mwr+q6g/3AE9AK2ftlbm06hX0ADhZXYRo+1WTZV9Kv0gHQObanH+Bn
59XGIhnbr3sJFRfvFiVR0DWE/ea3ArJLKlksSE7/wv2SPpiBCx3ymcDriYcL6LqUVVYY3tXOnmnQ
iWsQoASu9+CVPp/G+iAQAaK7pcn+IlzLk0a2NLoiI6QkvoU6DcBspM/L+sjJl8HzqcyZ8LwJwBni
sj0NHWFCegSTF4/7ZUUNRBrvohN4EuZCk4joIIpykb84a++MpYq8y/8lWIAJ1sR35DL/z8OPqWu7
qy4pCC50MdatoKFwL0WpSv99nQlxLeJ0P/NrFyyGZqksgBuNgVrQBIL9md37Duqr9b2y8CZAC7l3
7xb1g23A4JS9gZqYSNQE1+LQDGjH3qaCNE1jhzGovkEeCCPR8MSeqMwq2dc1w4GJXiy04jBGi6uD
9V6L1rFlQybnhVUvEjn0gw5fNZto+oVbg8kVuC70E3i+Ujx4RCcMmc3bRGJC4Gdt628KIpSUxwJr
G8sWrFO8TQTNe0GL8x5FskdJuEBbwwliLuqwQoSv+bfeozaDLmS9ph7dffnioJXa3IumuaQYcX30
qJD69u504sgY0N+DrPb2uUzI6/1Mr3yDg4bB+2DnkSUgH3r72Tmh7RpGhKQmvR0PNt6uzo8acear
zXpODLN974dhfsXRllB1noToZeri438Xc2ozgNJMs4XqbJjc1X+vr2KI6E8stkgamHWZAXj76RhB
5lWd08XTOFClri8a12CX9TpeOuHNHG+lOQ/EN302yG1s4V51WWR75AQOJTFeyEZCIeJjKEG/zwha
un/o1GhSshU9FMegWK3ZwZmjvu36WWvuMpAkrbS8hbRFh/kkuOjJ2EyNFdYXN/X2Wu2hHTbtWdFi
GIjN+XQ3BBHjk2wVXDA0oK2rU4gJIqE5mBIDXPJgHyVWZIxDimWZk7dQa0tc7YaXsDJ85jeIvCS4
pWMK1woRW3GLPxGRVHxXrXeibzwwjwG8SnvTJW06YEjvkwlGJgNGsS0kzuMVGsp28uijeCcpM9tJ
ygFBNZfqiwWCrf5HfjKcimq3xVqaaVH6KBD1OJcn3StpB0DYGeH5mHWGZ5dNgo5YTnJMrwA6CZWw
wEQbh9DS32j5co9o+cFVP7E7+hLLEcGIkCCkk+HexZ0ya60jnGjWyQ2WxxhZgak+KKMDb7kzT4m6
TdbWbMByLH21rCPUXBIEwTi+dPZ+fVushY8gXiuX+pNEFx4Bs56Ds93zeSyQN9X25B0iwwoH6eip
w23KK8wCDlhJkIGOOaMn49GTeLHm3lN7H6VjvWL77MhCbzY0ox+2sQEoDJEv+A90zH6gtjo40R59
irc4Yv0kxcNG5jrWivmijirTB5AX6ws97GG1WbANzH60neqkVbKPErpoH3dwCsUI9hcZ1O7DL7KH
ziVCb7iBLzbK4GwH05HCli0gAZKyQt+EalJjJKFoWNORPu4AVtkyqjKz/zEIf1vom7Np3ISxL1x+
rbjdyLYtDboDT6WhoXGP6Xc8GKRR4I546Z8gMWfCNu7poCsqYVTop/kJW88rJjHHNH1qkpEVovyn
KBw10wrPZzoLvGYsWActW6JUgC7cU9pUhtLJaVZWu/NXLjjLG19blDNPJ67tIylOmwirt9MHBUqb
i3XfTFjCRqnTh3BMhyK+A3PbrD76yQu362oetgCuLPER+T2vGaRkdOdQJDjsUuIzKIHChXmvUkuP
qoyiivCb7NXhTrkKTwmQZhdhxgXxdzf1lwqN1LyfkoqORUbpxSmpG1qfcFRi4qLAGCtna/0aLmxI
JqrRsQBI7CC3GyMmBFcliiJynhKk5t5YlBCzsyhuPCK0whceAe+TaXRoBRggsngojZUuFfPu0sE8
P1uxYdhnXGM7id59tjyfyFz9E+8TO66ByuoFUfFmtQ1Vsfsn7JzeW6AFO2uK8IRd8NlF+Wdk8Npo
CyRPe3rkQP3gp/5nMjqEt0Rx/Usl1SgT30XkYEvqC6FqoVrXkJFIE39QN7ZUSMUVhJKjAMR27D1N
0ScDkFgkUR8L5SnxCCLqD0r3uxFiw1GRfz/v7xR10f5IWAmJ8tyD+C8Gz7iTg4PyicV0bSD7Loi7
ZMOWcKWDKhhgXrNAL2+JTae/78BhWFxFq/2rZZj7f5mmUV4abgDEdg9KYrGrvIEngd2iuUFS90XF
JeZwkemNgfvubgT1QWZBBCCgf6DhELkER8b+i21IyYPAv89IZBnUQFsCtHTOYXCOgupwVApZoVS/
FQCR1cYJkzCe49xh6GaAUdX2TsYRBn2RpRGRX8r54wnkMJC8AK/mnQliI8yvY1Iz5WGnPHKin8+i
S0GpyWuLqO8o8P0WJ6UkLXkcBcKmhO9VP416YXTd5V1/NI+bHB3d7R+UyRZuCNjNpXTZGs/SmCwp
qF82TK8CMwqPhSpSOQtIKkwQHBKgN5715PQ/kGNljTPzfmLqX5cVqcM4yI5Jyc8uVzX3kSXtjHwX
d0Ktkw5bi0QbQJECKx+C3o7RSFEIYftQpMzTK2Oz8Zxldi/Y3LDWZ3rRMqUofcuYu5mDRVF7/ezf
b0T9DZCy2VYSHUKLlrMRmudSRk3An/XLOsDWy4fRjmzVycRuoOJtlbvPQBNiVgg3wlY8myuyWipn
JfP80wiIGSu5hTia4fd6jWj2gjOWQ1Gfa53C0YwGNEkZ+061xUSNaECBItrX8KNszcMG6JpmTCWj
8EfQ443TjXRDs41uBS+jfn1FP2YyEwDBaGL+PZCb53FQVonFCWDIZX1+OSa3zKQZnn/stYIWWAfZ
BvD/p+xtINkYu7EEYE+1v2Xsm2MDJ7TuCK2t2PBdcJV4Lw07GvGgdYJmGaaQEatzrOxQYJ9wRkuN
K4hsDLNZOx87eC1H90BcYIkBWJhwx+ZQuNWq9qiA8Agvq2+TUCUh9xHKsM+Jaay0MbwjohPb3pFj
jHLivnuxNB+vgp+Hsoy63t1JDfG1t56KmD5DGUAkqj+/Nu1o0DW4eLOUIZ9IRm5AExuPIVEaTzXJ
sFxdaHi16AUmziF2z6uo4yv7VMUHDb2ZTdTNJ2ut5Y/8ue5lI6/8o5AS+Zuj/Y3Lp792lZ+Fal5G
v7jtBNYnGg8latwnV/zgsQIgQpn10EqyB5Hw5aVXspI50TWmri3Pm4SVjXEeKDU4mCLBWvGug1kg
7hDPa75c6y32XRM2gfaok4Z9xv42TKWkt7tlOLJGdA3aghjxspQFx9IGm+H0NerGWYXlgOCrc/Rt
CwytTcBxJ6V332fG/ILSXuMlN8lLByAx9iCHPkzJKZ3GSQtbjklHK+77mFEVC9Ct0L7Rrh8qyb7g
FmKRg9NQXNzbw47IW7+5OJjquQZDUhyYkpU3jJgiS0XvDOeUOW6VEgIdGnTgVsZDYHD55kOXoQbP
Drg64hUF2H+m/s1IEgNbbZtTDK9IbLfPCLqA516nNjgHy3vBdJ/6z1Dr7T8jpxVIaFNFT03gaYIc
j/HpVPCbAemFoNbHmUMNKrRhxSBv+O5NnZ+ZCEHJuOkGfkwa9kKn39T9y0qjkwDzr62mAE9+WAGG
qFZdKB4dufnuF3wlqx/Z53RZfJdQVKSgi3rhLtluE0GbgN+sIHxu8iN+xr2VabtYZm/xPrkFtI/Y
V96XbyikpZYzjaPbnlxZGQMrqUE3Irh+M26vv7lRzudMs2omHjU8AaLu2I33tdagaa2VZvVGEKti
0xOmhn58a1BG7MiEgtaFCaZVwt22d4mGpOQIWvmG22g6S0ZeMJqhIuizjBhvOGY5v9yZiN8kJErm
UgEVL3eSushP3CqZZACBilaXbsqTec+tR+htwdijIBfo5Xj98A+0TVoFcjBPvcVX4mITeQ91gNL1
N6ENHOUrMeWLQayDjRMhn23W7d6KhIjVaEQOUISq006NxsPMU6WrJQHgtqPgTlfislBtlQrslcv6
OMKfwfZ4gaOQcNFO3zKay6hSBqn0SyHgYpICr6eB1jFFFY+COGQhx2F+DQSZj0jB3vspq12sisgR
3p3sPC9vj/Wvbh/T5fRSbHI5b2mbkFvMEciIgNgFFUpWU6rPbRTXQFmartVy5vFCD43b6uIUtsIO
kovf18E6yqzxQjKO8/eF2dbZHghNz6zd1NEwNeRT916Vicq+Cqah8vzSi688n7+hWuCNFWbVwhrt
cwlTkJw04lbJmkCdklocWT+hEuB3Ay00wfQFU8gs8d+muXOn7N8CTgcFPMbGCAbhxMIPNrXWSKYI
o82TXRUmk3xovaiSYB9kwn3hOI2jezyCwEzq9YoJvs7gWtZdTb2ZDT0XXQQ6HcCLdtD77TEUk+97
IFIo5f+uNkUAHxmgLzuKonw0qgJYZTJfDJYbarp1dV8YfdZYvcOuvFs01Mg0+PiKa516+HuO1cFT
SCdMaC8d3jJ5hsg+72a+bbFuDpAvAJ8dM5Tje6Q+a1yjA4vAbw4ohrqbFqBjgZXsiz8ZFjuOm6A8
5ZuL6pD7w/y9LBaHhRMIO/G0O3Fc9mFC+ksc8FIyvX6VvTjwX6tgMUObmJkNmkUKrrjUwAFwfEhv
+h/sUd3QoitpYMXvTPWp4iWPUAjWAhBRHvm4jD+uNtcTK3N0uJEM/gGQc1ZJGQqD3ygLa4ekL9/A
0ChyVUsaO4iUa8Kv3ogkzRapFrVFIB+x3vcpcOSX7zIHMGncpRR+veXS7xFv3jYzHDXV0fcIe0l4
wAnguKPZI/Es1jKioui/qbD7k1SOvpwL//qU7FsoCMTVMtfu5Jn9lrjgAWX//tQHGqYDc8iConBi
ewHf5dSbYyTi3b3+zocrbf3fZGIZrOpjTt3zE49N/r5VSMqRq+TYfITd75d7NcVUHPGUmZnfPnHm
pHyNORW8F52KD5HyyNzbeoKB9w/K9gnddH+BmOECgCEzD8WNeh3JwNYuKF6pW9WgFclo9kTfuE/2
Xci1hqX6Qg4SBt3zO2Mo2V62DOZc4HZkte3WvwuB31/qvSV3QPHg/XkufD4ykimizsMMxaT+RAm8
HleE1oE/aLEwuquji3faoHD0mA+2URxmyIGWC3hcdemOfRGoNONzrGK2zua6zgHX4i1o5EODpX+u
7BTx6EruDbl9FXZ4Vc/Xr7Uvt1Q5QY0gsYzTWjlC2TfMPLZAPl09A6/k1HVDNFI+PVdyHgl2ku/1
xtuwLWpc7bwMgXw+yJCcVa71Zx9S8aKN13FeC8uZt1Z4CiErYYj8ayuuQUofj33zmHyfRAg6b2EB
6yBfSEyeZ6YAPRawmRqcvm1M/EgYhumedK/PVRkDNvUy4XJRYIRhGkcPUxu/KEQ9BSXZGXEYEidP
9uu4/QpHkrafz/8uWfB28cIL+rlO4NBxbNMPEx6BBepRoHzNR+e8G6smYCi+ulLRrk8e82apFZno
YMpD0jNBUIRzQnFoasqwzLLqYY1+F8ih/j7m0jRSx53aFIERUp1axgC0ub+obRaQ1qiGatr8qcII
rosIebZfzoI0gj+ZFGsH32f6MV7D3RTnEo78Ge9ObTE0hSLdKMUcLvDcCTQ1mVNhSk5Y71/4yB7n
DI0qs5gWGZN/aLv1lGNiZzjG3eQSNwUmQA/wPhSAoQOAX3bA5HgZ9xIHMSwD+5tbw4By26O44IGb
9eTb6W0TVK7v0aYDrvWdBx3rorz/az0Y5QMudli5BYrZcomMn/+Bc75BYSeYaMU0Gfj0AbH61UHI
B8AXbyJ/tHuBP4lvZBqsdhPpNd7yz0jA7lUaqJ1RQ+ZoUPdQ3c5TP84mZCRKfdPd5jaY6+JqY2Ng
ey7eYqsO8Tcsf+soctqxRqdodPdgCFaJ8HMPbdujGo+pkPRxRMKT2EAWas3VEtp1gNwBHGPJb+rl
GveFU6J1nwKyakA/ZUAWFSJZiVpsfkKbYQwfH4vDBOZfKm7ehCOOXBNkH4rspMSiZRVhzTYbPVNY
Z33znQ1Tmxso2JCHW86VmJRkJLT1X0osRTN7JrMXqN8jp14b/VzM0sDy4pULHdg96tZTxBUA8jxJ
jt/fwMgCT7hoPK3GVuLwX+/oZdHPDImzPUTeZD6waV1cU/nWLyhrHsBCPMN8exn7QObyTu/ZTPJy
jVeLzqSBodPo2haKRTqacpg3wcfzEy3s+X0UJFkVkZcELPvikw2c+UZq0oRe5ZIZBV2ZmFz5hmdJ
FAxk82n7EtnCSBC89G0f0sDd+APpYgKk1vLkK5vlRuoFWcbY4d7zKk/XB1yPGHEucdNMOR2FY/Xt
b0d5RsogJrQk3NK339ouo8ofwhjx9KPz2VUVxDBqCexj2ptzPkqEcmOp8r91Aie0Ss6m0M+5MqxH
2XOo26rXidXsDE6twzdINu4FGa3CQAsSbXR4fKamRuyQ5tPY6hZ1A02pMwVi/Yj/olqgH9t1t/dD
7LywDPQC3MA/oyT2pJjtR7VXvRyoRz1zoXBoML9MkVZJC5ixaZKny+6Jl9WcqrRoqoQiBsR/6koI
RtQfTGcn8Yz0zspOH0PUx7vUDlOHmip3m6SCAazn+0L4NKS0uL6i3tzwHWfafyB3K2/qx/7ggKaQ
XMg7VMxavIcioHmWhemNUjj2OiQek9qrkVp25uzfGVO16Vn9twu0lvvGcjHKJMZMKkD019+mkTd7
jy2HNcpxlhIZrfm/viyqB4Blg4nU2E3cCBhz61XKHQrHPWE/ImoSgeWn+jgUKy4QXG6CpEVZz+xa
86vRA6ye+yUH9bknHCL0w0JYled7/6Kt8jcHjb7gQcIR25zX6Ls+fKTI0UUn7mTfywLzIxjEsbcD
fzb15po9kwpKhLntYT+2AY054nltoSU4zcKyel8HthXRxKe4F5SFT3yqdEHMV9V+Ks/ugxUXOass
tGhgShOVtyOkg8ONaUYk8HmO/RRfPZ6J/jE9VfCqewjizK4VIg2zeFx/zieVZQeLBvl8A6tVKlB8
Cv/nUb83QCQJuIr21s3V/oQu4g1tqoLDYXVxTtQLs13tMI2nV3uKdYVlnQuzZPQeINgaxsIFqIjk
2Y/OzTh0whBoowR9A51MwStngVY+7UTN/TGTW9gCRHH4EyJc9E2yd8yjpvmD7HwVWQ+vF48aJKTl
urHKWQdGaXipjGbOLJlrPyiXjLhbAE4CJlfC06Wm6FYMSAC/xoHvta21WYDNvao5s96gCu9N+H0e
Y11PMxr+BBG0RCn+GnWM/IRoJqCEX4YPRvrgicrYqI5SOVPs5PMa/AzOFmQJUxsK+Pf6HIjyHWfE
Ef5sZrcPFMFTn2QF80+JtnCSIGGn34OHyuZImCSoau7B4UGUugp6WQlaXA0QCcrkmNz/4IkDpDBX
2odtrepBSP4VqkE74O+aEyoGQuzSDbTBrxDiiNuXyhhnXazMCULN2JlhIZMWeDIhJ4aR/0a26+FR
t3GYbZunitLZ9sOD3bVBay7uBaV/YJN+gcICQOpUOCacNpJ1DkZgWTohrb+h5F4SaLl0uhl0pB48
CPVUrONdpkll/BuZVeoVtK7pcs7tIuBelpena2jW70wXD/G1pncgaG2IMhJGSYHEwrz8KkmzAFws
KR1Z9TNsuSWHdPA/kSKLjwWOWYOaxgjUwdUVU76pWMpdEyz0f7s2Y4UkU9igVqPezV4iBGrm6ifD
dVEggfAvzHEqeTQo0jtJjWf3jihwEkpiYpFZGAYd7IfCnw4WsVLi3h8Nczw4fxw7dsUGWRfkQ3qS
Yka0tPfeqtSdEt8FcEroBAHNsqDAti1hQPhP3+9uuc4FNFfJpAZvmrbNQozgIhH76IQIq2qNdOvs
Ed6THPhLtOuZ/NiA1tpz6b5X2QG3xqFPOY6Ma5cAUcVhVo+QJiyZWC+H0GPuqMUlkANTuL6UmjOH
Nicr0dLSq95dHjcWEQDVP+CuwMMoOmGQtDanaGXb95qk89xG0GhscpfjBjVr5/vnza7SWIi6f5tJ
TSyQG7qjZlKA+hLiaNXZ6ghfq3azEzVfQ1eIs20Uh4vltPpeHVBcQk0k2X0lPgLgj15M2WeqZTzi
bSZZcr2v4tKX7ObCg1d5qFRs8CM57F/CaXOlL0/X1WjIucxOCUAyK8ObJUecm3ljHx8sdJoh6Asm
aFbd2uKURdYHiwaL8YNFTmbiPmy1oA6IDnH6xcmRPdF2A/6OiROEia0ljqurGZYxdTSYDc9PXcdP
V0ejcXPS45s2RqPlwV6eRtmRorkTzM48cpqc/WRWRi/TF4z7KpxWPSflztHjYqviJX+8jfwUz/5L
XhMFn7fGqp2JP5zwxO6XrZEgXc18H83UuMo4Ot+bCEgNoEl2lZGV08rm8tMpx8rgyiEwEYpD1whU
IbsxJ1u6TWOZqlfESIHZZJJHyC+2S/bmtwOM819RPkZZpVZmPgwK+NvH/CD/7b8e2fp8srVtAFI5
DPjUNeIywZaAmhXOtkQHNiqyTpiRPKkcUjsyvWdz6C7enLznpX9KibKfIW5lUVymhmEVvjCquSsi
fwg0NWjtyTugknUes3AEWKAuoc8wPr7K6SwaWhpiM29zAf39yR23TxGN5K76uR/eqOS5OFOK191B
BU3dWjYPWRa92UGd71/w5RJFZDVLD0dnl45l85ANjOoTPbEm7oHJsbEkIdaV7rqrsjORw97A9tYL
ROH5w6lehBvbVGvxe4+nAl8Groh//MPSHRNaQwJ+34vIHnQ5JlOzzUJBdtXD4uqxKYUDvK0BTgJC
H9UU6nqhF67irYcrhK4gFyEW6e1hLu2TUCuCnNN4Mly+gRNCxOCU7DXPZ3hU47RxG/THilrPSAo9
PpE5i3m43OL4cW1crW4JCZXZrgtZS4T8vDrvRzvN9HegJ1ofti5iyqKGP+qAI0YoTBKXMvtqgOt+
IJ9Y6EPbtPquUfL1BcFBFw9QJW/s/Op71mjqLVsMEru5EoE29kV6arZ4wuPDtMbjXnm7BKVQ2UdC
uOe/YIcCeCXzGf5sa10YsLMDbbIMAhFXk6prhZBSzeqKIvoZ1V8vTdLbVBptgGmG+UlxK+EeTSae
conPzMPRXyISd4fRNSx1OQB8EnrKQ4t8Pea05xg2AnHR8l+SDLn3nLQIpKjEsyRFuFONgYtDSm+w
go/033LN6kN6L8G/0ln3cOVaH690K/P2PQbXJKfXo9TDxrxYNegEJgOPHqZfBcy38FB4P+iylrNK
uGh2QPYxmAGzlcwTprfROaZitf4vF3d1TSBKcyHCFdR4gaoiH45AK2q/h9ZuQZtqDJSQJ/bzeCLu
9OBAN4A1KUgsPbffohxhYTl/f2af4l/OvXnxN13wvdiWD/44QQvaGFQ7/3zap9BX6kWcno8ibguB
DNRJc8v/EgkBWcTaAngGE4GjNGzeK5o1ORXT/uOHOD21AavvEIH66LZwXoH2K2iUGAIn0o1uWYFU
Dv8YZd+tXDfpSvZ9puuWMyAOrKvgSx6Sx7w+aGfDf3SYicwr5IuUbnLKPuNKBomGfAe5MRridght
/zR99DZCv9E61qXlF9oy+ob3CdBuCYfF5FsB0/w9Yg7J4melNs9DWpq2HuDFGO5xm0Tdg+m0T7pD
TxdmI1xZcUf/kedutaridFzR0SeHrJnGp9d7nNV55T7Bzoieh8dXzuZhV+VbQsi+3T2Pr4qIYzh4
bqxMsiXJ7e2nw/aJGN5O0P+b2quPH/vskTWfPRuShh6pJVCo2Uxx6HeNwZHWrTsuIHv1mz2gEqx1
7jQwaaRamRGFr9BDHXw9I4597clGy/bKOxsRKyqrwHoZYVBXfu5TUySLZi/xcGRPJI+aRzngmUqG
ONMxSn9GmOGGDAespxwPqwK9OvEV4DLC67eDMceXZNCmNtZRf3LgigIeOX9ID+bYgOxFImYV2Ge1
5A3fWQSPhk+AcRbR1bLhacpQKo4nxxKD2o2kJgvLyE0ef7Yj6fZlMrW1GfRf0TSgPWp4E1TK69B5
QUaJjJzsu1Lp97NZGzjpRK3CTni/Q54BFxpIft/K0Xz7v4YIGlxmOdO3GuxJ2X048hMqrn9iKdgi
krGPriCV3lgf4gjcXajCTKVrf2d6yjpOhWnKNWbTBaJcUZiTmnNHCVYWOJ9+aYgeGcq5LsVoxYYZ
glMspF7reLzw3aq1XR0onCJHMYKCA0h6UfCK0XWAg4ApyJZAee4NY1FfTvyRje2sKrmAk0Xtdw6g
trkMQrKbz/h4lONS4Oi/CI7HEVgrNi5HXY7hZGCB/WQCR1Zw6+KBrwqEK93Z5hEUMU0OY4ui9l0r
DF5WrDJqPDqTGewbO5hwertNCHQ7KuGxwVZnCtOuHtlO+HY4lYrhXrVVAhnIMLNXsAR5R4QuHrlg
junEqWYlzQsjHsSCiPCicOWYadPZfmDjbF9lwyakM7PMKUbZfF1kZ2oJc0KYNy+fiNRPmhG64Fw9
ckYzIsNSQg8WuVe1XC+vb6TwsnqyUCEH+AN+O+XIGp+0jqqywm5Y5cEu5F7NkhajvMunsPLifqz5
7gjg0pqhJbZ4ijcYs4cTr+bhdU7yURY21wjgNbSOBiIzFkcgaHdG3yoP/CKBeLEpnv1WKOmeDUTZ
m0xt8snFbCDhVbDKIViDX+gdRGWzOY8CUQLGM83qVKH9rd8GzGzbQYQu9fQuj0CoKS8ARMDuRuP3
oyYSS5Z42TdpBRek2ppr4d/XT25dFi8Gh+qUwC/aPZzKZ+kDfsbNVyXxveFTSOUfbKy7S4i30lEy
323HN7Gcpf74ZX4k86mF1Vs7Rbj6aRsmBD6HQCkOxcjCPBJc4XYEK3CdEupGPLuo3SxYvTL+svfB
rE+3pEpP+eu/zK2zbfgj1sWZRvo8o/YeV1R/SLDGn9ytrT8+XW5yotsH84ufPIdBSxMd4gSj/4Rs
9j8YLTDTbLKyXhCmn4xJcSyVJquHUIahbgLkG09lDiupubEBt4IfVQu1p9RAvdewbMBKwGGycgRn
lpJf7toYUUbKOlSqcOexAPuMtoh35nR6MGOsSjqSDYBePchnLmliW4MyfV+DPAE3uIYuQnjFvTjC
yf9FZTtwDcH7XaOnzy0nTOWSkQz98G4nQIiIF0yHcN7R3G4adDbHf1ODwWmKUHkAmAWtZy6d74fa
sAR2pFD/39t3RmcxL6qil8gHzbUF7zQdfIMS3onTHM/lh6Ue72KJ+iYZsKGwrQJiD9LUPAhFF/6c
Ovs9puhHKoAbVhsGqPPybod0I1pObgblUnsNbhPN64MExNGKW3Qe1sZgga2qAQutctJQZr+6PZze
yh+cXE80QKKuYvS6GAmJ4TvWbhgyqFfi0CwxCXSpbfJ08YlsYRyBbGspnCAk9UTjCokG3XHCuE/L
JTAwfZ9PatuBGuazoBqRmeKIv8KpWxcM3fbsf2EOpwj9ZvudTNaEmwq/nmeV32TP/JdFP8pWRlIJ
04xxJpWEXNojGRpJr93yT8g49PyK9trquhdGFRh4EYIigMg+rlrXyOwhQOrwTJBlaSIK55nPuCqg
JLobB1beWdnMdcUm/B5NjMXJ49Wj57GtKdsVeXuNYMkQsv1DBlEcsRICtdIquYmeScaFTnObmuoS
fgln3ocp2bmfbQThpPVO6rPw5u8GR8vQ/9LHstmNkQOZJaGwtTlY9EsoBIlyrltjj1CX1cU075Ko
ll4vL30CnoIQSkn01TBOywqpuvdSAvlTXRhFE4TNm/yzNVFZ7PPiGhQ3+lYudgR2fhYC3tyA0xn0
OJ4oVQaBAOmKvnroqo+XLNdZT209i8Ey/0g+xtLzb9Oxt0vcYF7N4WMnmZjaBDdj8KY2tZC31tDA
1dNM6Fiu2ByqMdvU7wY3Oncga9J7Inz90IoqeWhROI/ZwJteiH5K6H+3a/TO6HzO4DSdixR/1KDL
Q86cXKnd0efhnacEKnCW1LaK+XexxxBoV5bIGKkL+TXQewRCH0V25iA/DsO/n2eKOrcVTH1MXERH
dys8zFe85uLkooepTkyl5bMQzZw2dXLG0fKAR5V1/CitvwddX8tQUzHbvmZCBBO74bx+6u4f+pe1
8OEFqKYngwL6GSUEyLmo0aXM9MYAChtsRZVipL7c7Y7NG5f2kOMG/BtNDTed1QZ2J6m1BAv3Fi/F
8cOMk2YnMGg1t4RgxiVSp8sJbt3Zw0rywA+9VeuG2HZMNaHZxpZvmMwpjC7obWOEpXE/hSB0HMtt
o/EywyaKX/CTABhBUDnpZn1/v5ZBuEoUSCXnJL4NCTzOHqzN8WfqKBvX130S8l80HcDeK+/FQqSg
ODXnKLiTLqIw9ifV5M9zBmRbRUzgFQqnL69D7tx+bFsDUCwGD9KtixZ92lqAdQ7EP5SuKFSrLoel
8xEE8Ck52PYBoT2mV+W3dlYB7Wq/m6fMfbanLpl+a2IyHI4v4y232m35m1RY5Qah6kKnW9mBMbdD
azr4W6U1UcUhXwt1uChiuU4jwZSoA/U8zz7ME72nBByEskkovGtoBQIktUdXOzl2q3LzErY9eRZE
K/0WlWYVB8N57dNaOMQDZc0mw1pT7L3oROyipTEqPtTBFDu39lYIIWNN284QLS1NddwaMtDDVsUR
c9aBfSA7bBgVCmm5WQV4DFRPrxRQT3+zCp0GOHyDIvVGimHAPQ/xEDQqONmYSgAu5ouurthjBzK2
FitVrnmEz+UkfoNF2jvrWtwMldbiliZ3nNrM8o3m0MULtfxVjJYWpOM6YVDOdE5IOd0FBCI1UQPG
T+g94aWLpoHDuSgk1ZMo0Lq1GcOSeYR1OWtcpNzQTc5tZNoC4dT9Qqz8+cawEgD34td4VWVTgaxV
K7PZZiYMfxrSFuaPG9dwbJw8B6MWBSRUwXGLZm5FRurbjCrjUDIqV8hH5qnTwPqSGxvsHJB1LdTF
gEwfrYMsRMu5bitj69jYD0Ng1DQZtvHtC/nfGLd5PNhSdHfnNoFRStW1CcmAhmGft39Py7T/09Yo
N3m/hZsosGtAlFoQtqeVyTz0N3U+JHY1ROMTwxr09elUggrYQkzqvsvn/3ThEpHyacBSmTapK7Ij
5/BCMIMyV5pS39RXNH3/2WfBjqlkcn+mJza8tTN4p0dYEasn4OlznG3ESGqNLIlHB1ZzXz+crSDz
AU4b5gaTiTwveLfhLGMYkkTRK421Xs9L2xvROHbMpY045ugBbypcnEpsGfk9nrJ9XFLvY2dJUh9R
HEoAm17fVb9oBS45lA1Iwb/UdEotNcDPU2Hp9uFGt8nPDDhP5K2xnd2JUmOz/eq71o7hPVJXToJy
EoZxOsc69xzmWAoOiDLcYzSu3+i7/yZ++9EMmxxVhCIR2OSuAJvjhoK6XRC5Rk9hFUULA+y0ZLtb
VpiAvisI1fF+25O32e/bemBbJuu/pfw3bgRpf7jq16oMigcBnSSyVlY8xO3Uw4QfR1q1nW+xnMHL
ROwqw3+0DZKlyuF1eFBQzrSZM8HeNmv0fI/WBcFtpYlY2rsVl1EeVRL7yk/2bGQwgd12yxtoB/TV
7LMN8zmZNhWbV2jLmhhjrIzxlZMZTbB138PICUEux6R3qHhIxGcvj1zgsDk5ak2NykvZgFtLNy8n
XukPDmM8ba9ODLH5swTxz9rzIrK+xwW5G96wvU1nJyYVIszimv80wkfIPGP37DyVcN839Lv4yCa8
1w/q4/Zzv2OkDsIDBaH2b386n0Zb5v2jZCTGfsuK7jXgefCq3u3MvI/NRwSxIBadkXjxXW1HSXo2
llD+bAhykK7oZCw7aHMWqKSzAfv6eOfpNYtAAf3j5kk48KVsg4X/0KAYUjn+M7niboPiUuAo+2lt
QrbarCr3MuMO1E1y/1+JCJELrTA9Lq+2zlttyoTDafpK65ZYzUWsXCA070wPeNy8un1viLvH5JcD
Qf72ztHufl4v4SOrm8lvw2A7JMNHYGU9vul8GtWIHPfbqONZbpUq/vxGkSozWtOX9Td5pDKwj7jV
aHHf4IiFAdNMTxcsNGYkBuoYAxxcUuFYtlvIHaXBujT0Do/rOeDfwM1Uo21+5jAG7MlmzK3fPYvQ
72+KyXlgLXxpbxpvcYfk7chdeUOReqvWIAYYbLHEimM+bCygu+xSmKet4D5JaBWRUmss9jf8SKof
r01bpflbWTmeabky1qJgO+Pjf0PB
`protect end_protected
