`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
R7maltAT+EIitkxYKhWLItgO7D9YVmKtur8NRR/3FO8Jcbgn8jKuhuylHx+EBWlT/xkflRos3hbu
fEhGekaB+ZoreKIAILBXzi+NO7IIVRrNYd+9Q+sdIBadN7XBw2r0ZIzHWRbKrBhikMLD2Cyddp/u
T+oxQKrDIUiOHML4Zq0KIpHrU+He6PS3MKKNk573X53BqLBorCl75wJnyz1IH+cNlI5UIRMZ7q4v
d9c4Og5/LAluO294/KWySJCY2caaCQRI53YONI3g3MUPNEWKm/PnLXOOzvuIYxikBcetuFaUQg0e
NgaIpR0l6ChnKJCr9I/xT8vMJeVX2UqKbc0OHg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="W10Mi2Gun0eedIR7FI3t7zxOIPY9LIvUeH5yD5qa3ak="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23040)
`protect data_block
bxo1zeeixeEaLtDzMg3So52S+ObUNlYSPe+vcjJZFHb7sno5IFQzX+3OGG+NmuYgmXCVw0THMMc/
WSFyRU+GfEFFcxEhVLTbyYfqmKE0mRj6ad2Po/zFFAQQUkeu3q0fkDLY7VuULUiklqaggnY+VxVM
ca84pdkl40xFmUbRhp59ja94wc1snwnOT/ySNgLi2+TBvxa+t+capq7D8ZfEwWI9HWUibB5cqQIo
aNKba2RA9AAnvMuGWOf97BshjcuoRYHLraiHBNWbmB6aMg8Dl7VsFHNSIq1253JEocfLKhuve6LV
w1SGr5EFVUtiQxKtfk1HbKwtgw+L/fkiskWaZbaCpeEmcTWQ2Xfy7M4oppBYacGS3F/XrlI8LgJb
rzHOUZkoouLxni1xZiMsdQqnHIYWDck/HhmMMIKkRdxqZXOR5Btah+qv2JgIM/+uAxXvUps+txyO
ZJxrLeYK0yGWzCGXf4S7+sMSVRs18bzpGkLGLUJwdpTGsrBdm38maabHIibXDKVTfo43x7Rj4He/
mmHsNKUZ47XwqVanQ9P7pBRymCoZCAcNWFPPQyChdNH9FaQD9W/260my6jpYvEYT4Xgfe3Z07dtK
OQuyGXE1ueHIzJwqkTRrkju43Q7vtY5JgwKTlVF52AL5gneABtBwmTft2MdJ794lBS6JUcqnjtii
yXW3az6bMIQK4yUMndhjr/elnhS2wqyXLkq+Udd5VWH8dLAYuDIVnYIR6U0RC2DnS1zoEeqNqU7n
gIM8VPg/VVHXDZUCSD/dSt53wBm9uuU/sfwjJDssniFW3lM3sEpm3nhX2T2KqvjCjOn2Z12s+IfG
3KUzZPpk+wwjicz3rJQVfgRUesA+Y0qvhKZY0yCM0/uqi5lpP+zAOaMt37Y3a9pcbNlpDdmRQY+w
35+lZrTdpIWdX3Al2b/pIc3IZ95OL7dSqBSie1I1DzwQYRbFZzba0f6cUEogvD1NCS9SLiK254WD
r1nyBPYm4YMahaONPKMk0tmDXo3ZQI5qZcU9LkXZFVw741s0tRxMcytPx2omTROp+ZMUSOU5xRbk
gazfgWnyoX2EKVI9/79c0+08dpO1sv/rqqNYfzhW9Ufo6frkS87omJ8u/HT9oylEGDOrMbUlhw0q
OMYzsCS98moMk+E+r0x8K1MVmOBODOj3KTDXkmOWdYq84Mm9eKe1LzRPrT+ybyjkZJhROepQ9OQU
B2XXtmzTc+tdYFVxz0FgccZmICzs+MrmMY9uRz0l+R/i5ONwel5uRqPbjYUKAyByCga6ELT4bker
ihSMc/3pA1K8uI2ovZJ6VMxl9Y7LESb82BZ//xs6XZVHWmTxli+tTRdbGcRBdkRkDCsuJwE6Qsz5
xCbdcvOswT3lURCI3vWRayAxtc2cyrE4L2O6VHFsZPZhGPiRTbhfwRXkUSeSfkYJM+iTXtKLW3dJ
skzifqcGlxtlB+Ikx8PgbkhZ2UZjIIDa/8InE6lxb86hfY6CY2HpfFq1pqv9Y/trSi0rY7GAeOy6
pt1Bnv8DT1WZiI3cad4KwdHtKkVdPX79B9UkWyIonEnR/1/2dYqvBCH4beOwDufl4BJ4Nc+y78al
NjwlN/jK+zZ2DvlGCknQM547rx3cwxfM7wiDOq7ShVx+sQ6Zou70pQN5/HJ79+0301pdC1G1z/1u
5iHlMIrUGNJLS/13etwlRFjdVSdHV/hK75G5P97DUhEEE6wE4I3iXgk0kIiHZF1GJRgt/9e0VgAC
uYVJDly9pl2wR3a6E+oeVkwa1iB6q8T9Gt4MFMfqVtSqy6CnzNxUW/XXGCw6WOcr/P6HA0RmCW9t
G2O9Gkfgdp8yUApgyWyCPMCZp0sct8ElWIARu6K4ZNmAsYUNadGd3YOoiV3kC1MdnZ8NkaG7aYRL
jtU+4fEN/j92I0n/mte8ftGVL1hiB2zCXooyIEh2+WdsnP6pJx3z+Ry5uON5XwkaZk5VuZeDc6KK
lvLsM/KcOxBJc9nUfXE+psZ7jZjK7/qa++m2NAvQIoQdlzBXkyKwZeOVaxYVSUI2Bmb54P1vIUcg
j7W0N8GbctTm0PLyLWHnURrB04EqXdMqL5KM8ncofl1GxZ/YScBeQayuhruBpjaMv0gipZtubZli
DWC3p3gglA5MIiKAyxINhRUNeUJqqHiD04CXtHKQ4vhrlj3fWLtPd8siiDYRKdO+QDXJ1ALi4Js1
6oci5uCaLbkcOZQnhPz0ln00FTCZ9JCkZZTo2PHlouuorJ2GduKktYT2jguLohJNWVqMLIQJ/wNs
SLS2kbIheGvrIhCA4SEtVhzkF2rNhcFGh6g6QCmKXoRKONFt8WM17KxeZ3kMJbiCIDzkO20zcjuz
oWvd2+GlP3R66rsKvTzUXOV2uUPNrU3ZC8u7tdUCcRGSK8apMFaerCd5oLhw0daN1WKjeRL3TN/b
SDHGAVyxSDH88HYnMbcHGTQ4Y/XQ63PQ68Uljyq11IGYT4QEb4HNnAJ0ymWsPczQAPxSUBLcYqAq
CdUjj5U8HNVzw9FDR5IfBo5FGD/dpssKl388JOIDwZEwFwTw7Fjl6JbQJrYGuxw/pcvLwqy9PDgN
VYsKfbbRFyLksKbpa8g5fK1YCbOWFYvUrVHRUalw/xv9meFxpcKLhSPN+kMQ0svZCXsXMUH2HBAI
sqyr6pAgtUGKcnfXnteQRAcalx+jDwcWMX3AprH+zrrLDojWNNsyKeoOFxe2i0vyBgczomiKyTrD
p+1fPb46TA8YEbbmHwpKIXM8bym32nvLa+uefjMfvVYnj/k1RZKBWVHKyP8vz4lEycAxovrsLdeV
HI1sXaT3jG4sUmP7j2kvKcAWLmOcHIfOsiSbHadbrIy6UAXeUd9yKgGAjr03u2XfEqv8HYSfxxaz
zi6Seu/Falt3ZHAr/xOAD6kCSYw0rz++9tYo17MQtnbMF9k0lDVy+IJUZ5a0Tx30pfGnIlZR0sDL
C71ltXET5yFLwZZy36HM2UxQc446S8MlD44aXqoY1l9m3lHhiY8onXQoYzZsh31heKTFDgvyfZmb
CkZZuaUCFUOehjGC3fkWnhGEYChA/dV5XXa8wL9scc6gLFNcqdyGm3Z/53kaIm6TARIf4jXan9gv
EHwLamKSRSFcKEn6owqXIYefn4r9Mn1uHdDw8M4eqSclWNaB9snChU5hhDMKMVuN8wdwHtyS2Exz
7XckwRfNaXwTyxFiuUz9oeXuP/r2dSUi+vd091d2XnAQPflO5cn7ozoBrVglLUPAJhlsDBI8J+MA
N/ynWR+mAmwUMqZIfezAPK45dAGm0XB35GY1n8llSV/C5UPx6vyChGJnGhuFEyHpAYJhqCqLFYHD
Z7ByfmnCtJkRFrDzZ6RxHC/8LgkjB2iMpzOa0ulMBEsMsMUgGnEsDjaFyU8K0u4O6HyeTXBP0Gxr
iz9GOApF1rG8v416MS7WQcfJy2ynjOdEaOLEyy1HeIbB/wn89GJD0vtBKyU+v0uDyxsbakOaakTY
VSbJBHu0YrRcuxIO7wfCYhDG26tT+I0HRBbZoIOdPVACHykqDccOclw26bBdAyvLtgOIrwE7CvGT
RTSCYAtAf+VCD/mUCJV4UJTvFtRrfGicO8MSP65t0GiEMWQX97+qTFbdK4belSJoMKN5WwCCZCAP
be6125hlwjSlfqyoGp1H58lOE8/+cRyEUCiiG6fm9HKDiRPGT9inlTIVjMqhjk60N0NH9gakzMXg
GEqi8c83gi4mc1AzYNjcenLvXEqq8+KZDPu6ZIoYPgCmWxBHnm5BLwkewch2r3XCVAZMJF30/McS
HHQkfi1s90fHdlaSxkOp0NG6MjtmavcINE4YDh6UbJ5hDIqbV6IRhvB7Rw0TsLClg1ZbYUE8zYYR
RnfDFf1J41/YRPHxcE4RcbjgrCbymAl43Kez3wRi8JoxEtYD1nhbNrRPMWb4B2bSwupm3qn6rZ/6
oWFDIEKyHjNznVQXz6BJP9fPMpuM3KE2R7KyOLVLoIrdgrKK65zcCV3skpRYQQMpVrQEHUEHuxdo
ZH5d0xoiWJu43vlvn+bL5sDOrnfVAYvjEuzFTzNtG94L7gWZUKVO44XhNUkJzQoQvS8nfmVTcZEI
BwNKIKVtUp+z8PXyUBFcOUQSclDdotGJK64YUCCgwACHBpCDKFF7q8UbgjWAKSvYVOLyqwhWckru
NsLIw4sDtptzXby+FPfwQBPaCacdYsBiU0iqm8X5FocU9XDEf4GpnFBMF2n8Vq3guv1+ukN1UVTG
HxqiGpP4FOqX+BhEPa+4SJ0iPyxh2HChqqeTREThOFSXbdUk+sLMF9aBkpWC/6S6Aii5HieC6uSX
8IxeyB7PR7E3Me/DalXX4byWfqx0t5TkNl9zk+hAW7ImaLg/jpKdcJsZpoaXSFz9mnieJlZV+NcM
tWw8SS1iOYyk6PIv1fu2ZZSmtwvUjaP3bJC4s5npDCamdzf/Dzr3WFBk8W+13gv1TSneMEn82T+2
wcfReM0j7TPXMWo0s8gwUOqW74HA8keKgHBhdZ93CJFdit0jSyRueiSdBRBFa19g9W858TALofPm
YK56eppN+gOQg9sXIGmw4zfhvX3ZlTocHL/CdkHts9sI+ExVeIMGNvbuZNLgz44yvo81pAgnu0yV
3U5KRqBYsTNyxT/6hf9SNlHvyhZ9d4MPDq9WGWpQMCNaSXK7epoIOGjt9WuIpq0II0qL32PK9XEX
NC3Y7XcZp6j36VwAgBDnD2XQj3vZszcIHU542P/b+Im+NYKXNXiN3BGcyc86ycRogPBVCkUwedoM
tF3KOjf0WZ4+UIMRWAMbsR1sfY2gwZFA4913+a20wODvqNKVX1flVFGxyxHNXeQK4LA5mDOfOCCw
lHlxUjZGwTIK64Cx8Wa8cGEkgxI1g9Qt/d83KrrvnUkhFJuOzZsXbkcVVbHT2GFRsk+3JKgzqNQV
XRFaYDEaTTJCuMEHEHQG9MgBKsccrTa27hSub5EBl0ZURqydLFtUNiCmBACXGFAf+C80tz9HQz3z
HY0oZ2GEmUbvmIdggl1W3pjg/I56zs6asLE4la3VeRZSUXFVOw8J7gnDum7XE4nItAiXmrRq8tnS
j5AwikLKuy5j74/WpJj0qoXiPwUZio5aN55iLJhSCAJX3Aado58CcGtgIs9d9Hkg6VTM6/Tdw1IJ
WdK4Had9/3Lt1OmflizMwKSwaDIcSclovphj2B+xEmTEl6t82TppuVHnEc3MDW5phmJy51tYimDF
kbEGQqt3cG360JUMrA5Zc/Tv1mLyuAPNn6VgF3ckhmBswtO/jDaYRHa32YW1jx1ljRAz5E91o4IW
cYSiTfihDN+HNH+39eNCHRSJS5OfmsYKRhxrX9I8V7GdTVTl7rIyEus+phsJlOdf0mnmdnJ+hF7D
BylKoKTemgok+T1hs4RRVeWNI2jhNZNpp+yz+NHm19D5GOYg95M+G/UvIFtjbmhkSDPhJkt05y2r
msuOKG+E2H1p3cYXy/l0JZjjL4v0lfMEzvH4LSs4jyad6r6jjdzhydSKpeDnC6dLVVpSf9KZzWVc
VEgxd9BxVHlnuNwCbs63xwdpRreYiHPRyScG3AAyVbIVzurX2TpSY3YDUaOX5uwhll4K/Y/k9mx4
Hmukml/ZItWLUp/0jHj9EPnfMFL2MQKzUMza9r00dgaaC3wVnId8UTu3O4/7guEFacW4/B4BIh1E
Bc10t5SHrjxxqaOPp6I11TzsqSuWXmycH/1UJCm5QKjwTRVW+zmXn1M+z7IWBdPOlGS+pLsVOuJN
9T3dPMddspJVAxYpZFLN3K7jzBn4E8cxGsfQOffmkPwdGcuvXZncGHux8T97DtDDpgKY/f1MiCRU
6RxOICbAH4fAL2saaiQttkO+798OccAtNytT5AQ/lrmjCzlbYTlwdoozDZEE/M1ma1IUZBR/2EEZ
HIhTDfIf8tgVDVPjb4W6LNF3WFBYqAfaPe3mxI88jwVb7zOicQbN5AX452m51P/K+lGvDOkN1eNV
tDAQoxIBSsYG72eEQem+SaRV3ndFAKMZcswxhTX6JADUkibiGvlOKrMChU9jLIAcEbc5eAWvoMyB
7Vc1z9qWOxW6lTHifZhW+b206aACYNrMmVHRwHwoDod7tuNobPDiwJQdhqmySRl/+BgGPDI58I2R
evUZSawtxp4MOjbd0COl1b1P+P2198Ckj2CLP6QXq60Gqjyrgq2Rb/egrCJDYSYcAjSAfe35wrxn
i1ESTvNNHix8IMV9ISdbjvFZb+yFjqNho+LfXLa7ZkX1bUr+qa+TGRWU3U4uS7s6dSwSNPS6Qox1
nzdLwbOf83lsPouU6qqVxNn07UL/THH2s2C6/qk4BSdd70qCuWF6bQztEE+98jvRlo/MgIoigWLL
hAJynoj7ducgRFMF7PmdYd340l5RPI8I4nSL/nUb6ocrhdi/WYbHjTazy3HTo+FJP6NL6+8kntf2
PT+XO5r+lo328O8EM2YiK4Qf1UyCjmSLOnyvIds+jCmxhLNdQPyczgHKFuA/RFX1y1l+tPMhTo3c
afA5BGgoa1DIbWjOqM9gl/o0I9hyggCqhViDWqi1iLXUpgdnhzktxPd4I3r3AUp4OmuDt05hM+XF
LN2s1wpXV6VivhdSaIMUoxlrtn48mRq9HCgrDxl3APJwoILztgZevBqbRprPhLma8FACa2C931E8
dxmMSL+vf96+4/x/zTTQLCELGtvNzBCmqvN13MGmgmbKtFir8JblbR2iZ0/fPTv/9C/51oTkFi8S
0mp63cK+gTI2DHm4zTR5trbDjgLB9miGOoS8wb5zsXAws3Y3GrAT+BhLWO3Quw+SfFxcUlZiiFJ4
jspOswj9AAFkPRej37tbSaevNBLZXFpvaAdHaLYTgZSO3cw71lT0XD5laPqsyPqC3CA/D1jdvxm4
F/hEtWE4y2t5Kw/IaE15ECZg57SS0oTER8V6TA28ni/R4AAUNK97CtgXGCwZd2wn9nNcUZbFuzD8
XulZdPILYTvPE06TE3ITd3qROLUTExt8Bq2JeoACB67LxN7RcVvgISsZZ1WsWMmI6PnSp/+qzvBL
JjQc0usvZU3WVvaKZr+wNq3yqjADqtMfEWaZ6FqIQtBhVDKlX6+tkHrKy+GWhAlzTPVlr085Okwr
rKTFbEXhAynoisSA+x1WCV8xLO5OwFmjLyqNbn7RbtlBNE3nOuMJ0NLYcqRXFU/lKglpKNMnZNfU
X4PuVcFtEWN7ERMRmcJMAJ3rCB7S6+xH4GGJoQ/8d+W+430FqnqjdMDRSq8uv5huIkx2QTpG7pfG
4ktFssi3Dn1LmE1wwpdwF/6MpW8Uvp8MGwwqLnbGFfIIUJWrficN7Do3hrkLl498VAL4eKGPao0S
0kLwwYtRnz8tcufLV0S3Vc2L85waW3ZKWL4GErVR2xnw6+w9gpZD8V8lCOjim538xaRzE597mYII
8wudPFvDCcAAndOb6KpVSOczpNXRl+fa8YzHuVSgQWyKITBGS3w1VEmYSQKlpJe2WaND4APuloPA
Hv7nTomykxaD02NIwGgAwdgJN7wzJ/FT7Qqq5ELijd72RQaYdJ9S6gHjzjLbcvGSCBpCjcaxkAa+
zlNpWp9OoXC+/CkxCbyE36GM90xNg6jsdX8fJkEXy5jBZNuDXaGufFSY46zYLq+9EwhyiUEz1hSv
raECpoUI1rD6hkE9hgwB+NKDD/DW+MbmP8K4PJZw7XYogwoXpcM39SUlxPEkgntpBWwlxW07W8gX
2yBA6ap5A0JcuZ5KjhqR7C9L60zaNS1G80iocJTD8dKjnPVMMe+Vn4FsisQQqs9aniSdeRSr2emA
kq5HuIzIpMZo5y3vqKJ0FhbNYBSlI0wj3JoXCwZr/uAJnJWW1LOfBy76hIaiyTBchLllqOr7Ww0x
JQ0j2RrQptaF9znYDV+CGdD4eX0BQdDlwOk2U2TvDucXRzMit/u3xTjx6MrdGNbATK4snONAnWk/
/jpf6bo7kwidVA89+Xjopa0XQLZC+FDW+qRokYkTnI/0p0CqBsotsJPnHlTTQot6kAMKD1IrpoCF
OXXgm+oBm92SlYbDqVBQ+4A4kpt+y5M0fdICcF1TG9a2dQmHdVFC+SgscSxycRV3EF4xOaUpSo+X
1KGHrNQK7VyI/yGxjObcFwTsa+yV5XBdr3irJvvPRukAKup/1JLxquP0rQuGau4BwpEwcEHP39IY
UT9YbXIdq7jadsAmR5VzNs+cxnDPYgswtsYWvkRu/aspQNG5IubH3U7l1NN8kma6YHVTKSHQ68mD
BM+hIXx/rTyYbxEFD7qVe3G8VCMt4DP43GQUjJ0Rw+KbejJs+l/q7GgYgbWbeNox0QWtCVIBYGAn
MW+drO2A4rH/seOYRL2EwELf+Xto24ZncUxzmsZ8lmkK7gHsDj6HHIJw6Vk/GIKA/5G/3DIiEsXN
WaW7y6jXRmRXMBjfw48KEoe3OWB3w+YvdFCMAK8wZSyD5bgJUhPj2RJFTtmlA2sF/RuHtcQmeH0H
7oIyvWWkJbEcvqZrmp1j6OiUiw0xerKrHvGl3R5SZd41UW3aqJrTbSRMCYmSmLebloHJiNCWvDxf
eSJdxBzshVxJ5M4XnkB+EJyGQlnFS0yQYuNnB1puapmqHCxEQMPcvlxblymdrtAvSDaIut2Z3BxZ
2M2PbidkDPuEAFF/5WkPcFeMBFLv9aqFUMd+C0dLUgcwN89Ismlb5yte1iQd4fxG3rG+JBB+WAq5
t+bu8fEFsFAbcDcbdTEmpbvgg713m/XXQByu6V837UBQastFRUMhHchDkQISSF+nX61fXaxT5/6T
QeQbxTerOaIdsdE9VCHU2LpReqwcQ2mMCag+kxP8VCUq4SX5Xs9ik2WfvRQdIW+1vtyHwrmlAoyh
D8c2Mp47ojPq+/mLDkF+Go1ir7enZSW8QbXBO/1d/68ZrFXEEXYy1V1qMfh0AuJcDPlVpSXdAxqE
rMlZdoG5pMn8NkN3M+BfWIwHG1s9hr2cBSfHuqIE9bzAuecyss/iI0VIXd0dfZvU0CYQvQ2iiATp
97MLQtfHE7xO4oZBbPdwJNPngK3Qb/liiRwjmNNXTrbzHT1Ih0hDpM7oE/LhZHacgxjfKumI+eZl
nIXBI3zesvdLhoQTO/nil8zW1P1GS6H6xxTOWuoeOZTKo395tugbVtgCgnzVKxGBq2eVI4Ymn/is
xf2Qqoer4lO2fUVUXuahD7VFtGqW6gLbaWjWPCWi2hvqC4kPZ477FOFy1IC1JMnB2N2zUdP87etM
PVzFz+BPxeAOVSpJUyh1lifF25wYP3XZJXSwjFxu+YaA2LyZcYh8xrlTK3USvNIarS+ZrtwvxUoj
QtqD27noHtU11stebRSu2X3qQqMw1YGWjcftVF43uv3fz44cmTh+oFfOH9upiX5GfG/vGCTCV3oV
+fE/+5KEX7QCdfZlE5uHIgK/XEaynwoAWW69tv6/4jAhSGpPNSXbd8HeIeOR85mdHriKZeKxTtw1
xE92PkxS5xeEmbKAEADZBWXxjgN9upmpCR8d4vO3ZNXBA91g8a+q/YlAkpa9d4Xxqb4yTZ593LdK
dSMNEV3ZdLwCxf2a2R50GsQ94zEE6WrLvBX0J6N7u6wPXqqr3mJCv1BCeYo3dJsTXxXEUiFlzR0C
Vgszg+jyug2TcZCSDzduGaqNRULz9cc+KiqrWYrjWk5cwzA9LbmB8RuDJ0whLfUSremJ8uLG8UB5
jwoDtRk3jyeSgrJsNoBwEsWX6zjCSLsqY3IRMUm2pXRNrc3hItftVkSpukstco605bSGczR2alhm
n54N+a08MTmXI1MSoqLwmpQUCSwAlE3IQ54MWVSvuJbBEZfRyaxyMpEcN4yX+umE/KGuZwZXG4sg
aWUIrVpSgcrNFmuxnziv0fIiIuCsH/gJ+/JR9f8BLwhplJkYo1OpA5iUTIWWUOhUr4226RLLTUZ7
hNxYavSpQLqNkpPCJohb8LD5TdKUSccc60H9XyyKXb+nstmWUPJoxu1QFQGjbp1TMxZfZXcogPkx
MOMid785W3hGTvA6QGCHTek9AoBokj7alVW3SEU7GToITvfR7dtokj3E06qy4PWHsuFq1s0pzvx6
yBDlTLmFGA3yRpGjte9ygoJd0eVvlp2T3ovRt4HYIoA/b10h1/JfU0T9NwLzLG3bfuLRmP+fYXah
MynZHydgbCORy5rjXdeF2KTROCBiS7olv+BFOnGTIhwjv+wnnQSXBWE70aATj2D0wy1f2tJ/jR87
HrakC6ZwurQeN8c7lCAhBCtyCqNasJ9iCOSGKra1vcqbJqJxxrOauayXvKHHOAHjoVOmTBdmK1XV
Qm49hM+vnrDwsPWNoBSFPOOBX60xrpPixfpFlSur5r1Ssh87D7WJXvqrIbN1kzBoj3EfcjzUPDow
xJ2q0yvND+fXvxu1TxlXvUkQeU22C/EQFQA22OrPyAiNS79G9bMpFFGM7Si9h2wFZ33lJoMh0efc
KBYl9Jtfxmwv2Bv/oMy+lnOtI5w2NuEIaXtaMukCtcD330xg0KNZxpXw5c8u66PQKTVHQdMZWrft
yMU0nk6G46d/VdeNTDSKFfCBiY4Mv1xJVQfA3/hLwEBq7zGWlF8P8Hldvx73zVJPWbgE/KGL63YH
LZs3tFdNJuuFHMyY3T0ufpe9LbG2qYY4j3rnLDp8/MO1b7m594+XqTgigFpNWrfYtNhHp4IuCvGZ
GL5kpbvVkDsexUTayoFxvRSCj0rTLKemoClR8/4HB8m2mpPIBJNWet+VIZ/qEzLhbm/480pD8g89
m5UIBB06tdcIr5FTfBtrxZ6Qph8WNJACG6N9OlvT3E6HDuMwW+bayhK3Xajcwqfd/JlZWVi9wb8m
DuHyWzrlMUXb5qfGAiOvlVyudkM3S9ZVPbwPpatYTgpfd8ikd8HfM6SY4/pkMbpjKpV8nc+CZSRg
4PoQcd3v9tAAu38+z8CJp4kpEk8xw94jOrjWy18/nzUAJVwnLsAhSer1n94uTt1kGVkKcncMiwM1
yrtKL9LQuM1mFS/SBgCOne4zaa9NqkcvqrEX8FN+pYcHQ0UVH80kOBjPJcjt5dkoYCy6M9GXhCIN
KW7lwXfFfW2cbsbXQ4gL1tfw3k1/yzDXtGBt4NcwH5bcMRhQWBPNgb8mRw9ER5cO4Q29nTqTiv40
H/bOTZ4kPpAC6GCC2rjLr+vGbb+6nna8Lz0MKEFmbsts3pC/6VBm9qPoaA7qZNS1cJrv3CEzYPPV
mRl6BLZtQacBLbQ17MkjHbRXY8mEjFZ2QN1+gVED5fx7sP9puCVoHYTHiNmTq13DXojrFU8CH4qA
MnMMfQm407omWLEYB8L6agN5CVd30TzFden8AEyIHWQSPZgBIggq4E3RwOWD8d3f8/LahAA5S29A
xpt4S9v789Zh59b9xDlaIvZ6CSfCEoFwzwJiSViwheXaHYeKpJ4rBTi5QNb5ttZgR+APvxVIZFCc
pQWyqlYNrwt+sOOfmZ7YJWKZhkZA1Au67XUtnVhfonusZ6/smTw7pp14010RaHvo2o7jq9hxC1k2
qnz+v6u1XUL4fLPG3gMDK+n8j3Y4esuvrnUORGDg0DAYdv0TgAHXD9JsKy7lzD0wbXR31bGPCe2g
T3kxETVJW4+2aLxoyFrUAAZmkKE3l46uQtDgaI4oyJTlBfYsCcMRdksNTzZ560J6y714XTNIAwJz
OR5g0m2jLHm418h3KAHIEZmXGARBVcDWCtM8Zd06TgyPzuEYdnnYqSaI/cLU/ldYDFFUrSVCxRYZ
w/ic8Q+1YpSLvnEi10pR6lvQFG7UDk8Y1IyBltYoRIChDntP0Xu6rQEVy9iGRTLYlIX+68ienOiw
pUzp4BqUSC57rWfc5EyYMe0mS4V+2AXckMq3pRjuMOh8XdAui3C9ymqVsfKwutxumTh9Ut5rud2F
7q0L/FIQ5Q6hx5jnWANJ6PHg69p9ShxYHY6wXeHROpqWAg6qIkzBD/UC1/vi6U2uKk3jyhOtLpaX
2j3ow3qxXWzTV1G7NpBZgdtG7qC4qhGsinmTuxMhBhWT/MOr/n+gU0amlqGlQyauFOSL7D9manJm
93JXAm7GicyRhq4+B6s7Dhyz5K2sznGQ9JPtFEKymFl4Svp91U6WZlKvc3uCatWoznZmS/74sBtx
Ybwo/RUa6Ubzt3YKD9qe1y1fPkPKCuwlTOUkpDjkTR5O0zDXj1Y0vstOJHVyzVeFPfdyTwPDimUY
Yad10nrTyN4CIly3TG9bmR40URrKGC1F/CXtgyDri5nKJwqPO7oOra00BYdgu1yAQ8dBW9ozm/4m
JrAn6hYeEGT/ZZJeZUPfaYFQIlS2D2X+0tbPMzL2KejWssdWSYIL/RQPgfXecGP4VHzqpzVnLFUM
0dAG1lmbKM/C/JU8IvH8a6eGoZYCNMbmtDmnl+aD7ewEBKwrYsOqcmHXHCJIxEXAoYiuUGwR9N2o
OcreT4ryIWgbFoBeLDpCD8BiSWriqMMD9Z+bzroGd0k+KGUaOkQ+P/s02AEla511LKP3u7ZS9uUC
vKZmoprUxEAOWe2O4F85W+AFmyaAWnnJ99dzHBOlfejkIsSh0SFvmtIu9nz8+UhvLI3f1LyLFOjK
o6tsLUdzPZtOG+XiLb89dyhGgWlrBPa1m3uzauAe7hJ3t8XQdOnJbAGErhGncCB1Erj7T5cQG+f7
qDi+HOOIOsbQjZSP8TCbW4JwemIgihtoyxb0bzRkEIxE1gknJQdcGL9omO1M39BNMpIdI5OqLozR
Fjs/RoZIAKaud3v2c7LiRtQH15R3WhMztUiitBX13L7EXhNSt59vMizPtf7WGDTSqO1YUSR1upmQ
+lo/QAYIlHvGjs/xLraZuWcHGcXkflC4EzCqaUPBVEUYkCuDktL5S+mq1M/0YVqami1w4A/4W8Vw
Yg1sDhTsgb0efSAg0+CfdTTj7U7waStsfydxwCTbyFnTno2L6IIQA6Lbd7AKrm8hP7a0hPUFVL5r
vXK2w0iQSQr9uVguOE62Jf0JxgUdIGzY50aLKQQuZRirEUusXY2KCjizB6BDOhdeNddKZcRZK/tK
5ycEQw+Gk4obUKog6ALol2Id5JcTXrslVLJo8WjiQZ93LPOVKm+4iK6zaIfPN4ce3XkiJZoqex1b
hRPG8mb0imMHw7oYgZxCJeGYkwsHZLVpa+EE3mj1Dhrz3Rm2LPIqIgwBL3RobPuqCB2oTbDetLgE
G543wnooyuY5qQB5/UQrIde1mKRbzQ5m/UEt/3Yokz0fkq2XaB85sXRVZ29oBaNmr6rgCvjTbv3x
5sf0UkQQj4gHY040SvvbFZFKL4ONo5cfN8YTSWoZtiNDL1g3o2lGBuv9hALFvMRj4TNVo4bPSF1q
8i29lGWHJ5s54GXYCpfvHXZQ8rkvJ5wPBzbHWIpw5dshc/QpTAKXI0ThlZdWfrv4h12+cl9ZhUB1
UlhdbGwIUj/bOq1IMmdk986kfC2WClTpgvJV+WRZrvf+0yzLp0lsQ0EQAysFVdxMVWJCxLz+VW0b
yxHnuHuZIvzv5FqXNSd9DQqpbJd8LesSYwMedGNZJz/I8BbrviTVrpuKqpEv5eKDCv3sd1gpCkp1
NPjx56ERV1Y6JbdxnH6IS0hVf22nsJb966ll3DhzvkwYPQ1jttEmeNi3WEqv+LiUNQyyU0/pKxCh
OoiPEBzsMU7azEJc2IPUMHbP8+GWpFfkJvQaAY4MSyMNI0kzc1s4OzDK0MKSB29mRGAyLjYr7NHR
bBlGM+e9oGHlyPyBn9w4774SYK6RwIbFLA9HOaDxkiiZDzNRmZtmBDYHjdHhRYwFB43h8958NFUo
cHqiL6fW0QODsSd/uqlBoTN45V3fhcLTR5td25R/FGl8neWUa/Nq3dunFk2pC4ignMbMlIOihhZV
zF1kjyVk+v+Vy2POEFlvAeQCcHm/hYjwo7QuQwT5gNQpg537TehR66Q0MdXA/KcxyjJSvKzm5Lvv
ClBXVflcombK4Iv0LWkH6g/aRYZOtJbCzTjXBGtqPqS9AFBosBbRBZcCftPupWdvfbRUnG2Ej37p
nFdoOsWbxskWACLWOvSgw2oby5MdN4U8breELZBozyV9KXvtlY0uHwe/NqPSLC0xBGORRhn+aTMP
Es8Irj9opaJ58CynJOv0RZlxxegjABQ/a1niH34wgMUI1Umjh31mDoRbtPqWPZLbTm+cBZrfoyC5
ErVBvhIU7GOAxlsu65tuEmZreuKnpIKhNqiA1tfjbuJ0Xek2ye1qkA1MesX3aD97TXN4M/DGCUpn
/qXeyEfdP38qK83FmIEvz3UXu02piEu+dhXD634RLoEPVkyWAr/XJdaPDZJvBrUBXevuZ/4BgN35
85ZcUhX3zSTTe21w6AajVg4Xgddas/3z6EkVYnIspo78fkwP+UAC4GrBka5ZYWqu6/9tWbUpAG2c
xOsTgmobHUgScE1r8u3BJW63DZCwrhWLGDNHeyyYLyoiL2TwAZ2USejJg/QgnltewnIz0e0fZqqo
7dRbS+xuKYoyncR8FTM9beEbiA35XNv+cwuEUS2xUwbFpdLHgQfnD/MODwiS/+UstcUGy/RG0vMC
tSyPGdjRLMKeJf77eWeIWB6+fXLkOgmxZDiIGGqE+xzKv36lcwv9pNQqI3wg0MjX7Mngy/gZxxqQ
rPVk7+npcoWr7V6FJ1R0n9EGxj4NOFoxLCjKiQsPIWBYK61+DBO6pQTO+e+C6LaO3IDGZD4o86L7
mZYAQZaTAO5oX6jXo73WGVyZYwCDFFpbFeO2fbBu/mwApxMVMvmeNZ+8PIqXXC5/v72i62oSXcNi
JrRdcWh5PGzZCXMeLLuIWzjmg0sgnbv7t4DjK25tPawZnKn5NcN+e70vqxV1auuEV8hjlpNC+r8E
gDwN7kKuBY/hvhuL3aanccd6a+B2mXaJ7+e4vXnV6HrM84sWCxXd2BugFJarjqxSWCSjQGHc798O
oYjdMO1d8k2QmoIaDqEBZ4+neGhza4abBkV/5HlPv6Dl2c0WSAWe6kKGZz+cJqK/CBICCc3GYmfK
1QllTVbtCWBvH/i5iwwUejNVW6krpAMta6uWQOKiGJRAmh85M1E8Fz1GIoklbVHi6uwHdQCFk0NB
3V1L4GsX6JGhNBBcmtARY67eR5TtZ0Cs026Os7SvLo9MuPQQ29odmU4zq9TWRAULMwVyPRrnvabB
OlfLktOddAd1YtTxf9QA3s5xUiLUDjxSUyUNYM8ZXi2kiRpAI+6qaZKZDWNz6/vebFZGBrYQaub9
z5BvL4dU75MLt54kG9NOdDtTLnbOBWppNR2f6FodUTojwKiQPmBvz6K64TYsu8bpvmdnjDN3ivAU
01C+wSwixmErL6quD9wL7hPoDBWliQkIRSmGdzhO1m6Tjb/yY2MKmTDz2BDDSXphtYv0sTZR/tjO
AfjUmyjNcv8N6lrHVzjIoNsKBSlaJ5AFlcwiumIW5ZB449nUlOuA/IeGfXBrs6VqP3F6hJxGe6pf
Xc0A0yHEs4ULaz4/MoZsRyrqq6Pg3FkdjzeTONrhDnssouRvG6j9YaFtjwQjhQhkxp7dTLQcDVK4
c3M9F1fjI5zVgzXABrRWJ08Isy9jK1RScL3MP5DAM5+Gr3PXrwqzQY+luU4Z85boPNMDMzsANvPu
Fak41B7NunBJnkKma7b9k+pbrnN83Noav+9qiOn0Dw4sWntAAOglKhnnnt0GuiBCZjRUQXp9WigV
uAUQu7cpfcMdqHo2WaNnsq3zKbUIlL+aan1wEbVZuA3H8fF3Jczu6MlclMjAcohmWxTwACBP4puF
l/mvL4D7yzHQkhiLXmK1WT+p29Bj9MCjnb8f3P3Cya5qYzXhbcnDmkbS/1Y+qSUpar9jaljGxPuM
NWlnCKYkGHdbw6mP6a6YLI9xzlHGXJia03JLLrlIVNbfkuV+RP9oCB5ViMRGytPpZZh3JrEeJZVA
nirdGSwrG3YpO09blIWu17RCivTpUpLjGja/xUMHNZhoX4Iq7J9Wdw9cibXM3EV21xJ/O/i71p0i
9uAYn18rrjqIS2AjZKcLSzMr+WEjeCWDPPHtcdYCsoopHFV9EG2yASC6oQ12S657auDBRXWucquD
+/FURKZYjKPmZUVKHPu4rQbjjwO336VAhwy+ZOCmWaJWHBG4tBAdnpgFmnD6tdRRAr0vk1ZLMjkp
ssxwZLt7nkNArL01XvvhEasaG3tkJFKKNz7mLbeqBtSf8i/nI5D5V7DjIW9PvVO7N1HbzZ+WPvPr
uDZsz69u4cHZnHX5vnfykrWEwrLeaBoPn9gft/HshrQr70xaVl7qSIC1NN4R76IvjYSu+kx5OA+6
+Zg0y/B53PP5upGq7zVWBk9kb6AEZoGR+ATvzzme84bGf394k7ViI8bNq95p7ORX4jiVY0V33NrZ
NqjLPMMbD2PPFbQcDQUfq8vRzG/v4Ra0MNHC2SlwPWCH8n0XJdP+rW8oLR75palKgAxXi/8AC4uO
W5TUlO2mlXnK0bBkJY1CyPHnGs4uRBEu1g+wYjj+ZMdHCyUk7QtwWHENXgxj8uUkaovRQtXK2a/e
f+Kui6i1qICdBytlDI7PLHWRFnN5ozLn7YRRE/1UGfbkc9dAUL+A8q6NvrjUfTZ3gzNOay6Wz2dd
fPMa/AmfzowGg304IAaAwF0pts9dMf8w0W9zupRR3gs/RNzp6D+E97lnG5mj6Yl5DUyJLYrFH9me
5Q9kjnUsTfkAMA5821cmNkiRrAf8FTc7Jb5IjMhksrfiSsVnDoUG4LuC/4K4QIS/Gt7ppqoa49vF
dCYWBFE+bkBZg9u6hfB0nNf+RA/9VJhDI0e1WKp9FIainhjNHIZoLv/cJ0ObgUAKsDaqzUBe0i6J
Z9GD38rI/lI18AydBM0ovxCG5VRN2Fj02UKAOxYme/U5gesCByuJv93PgTK9ZxkQfgNTjUYI3xgx
rF0aNoojFn+oMKBnZQEFJxjZK6cgbaaiRZeDXeLpRYtRPMFJuwb3laeLGuY9jccsvh7mG9xrL7SF
jL7dD/0cIEpBVfUaKaHvtfljuM1MnLkdoV19tQp/GuutIYmocjPbrZkpnmzF6MNVay2MQoUzlkKy
UHo5yH46iYdcoEuPaxXTiWYKUPmEsCPKXV4tII5n/+VNqk8r9aq0iX+42zfHRo0thMCOaggApcbu
pp0NR/WGCRTMJaD5/5Rcx76rhvd9jN+b42c2+ZG+0CsgAPYAp4GKTS7SY1z/5TB+ilwn2fs8Q9Ep
CRg56GmfdOWvuiHMoUJ9amNJ5HU9KNeJBJFSIh4AXbIgx0fval/hPuTX2KwU+XQAKqZHLEx46IQA
650C72nqTWIoIoa5Lmi8V02Tap+TUX+OLp5Pn+9CIzZ9g9GP5xWuwnebl8iyv1jAnj2tW7Fw9F2Y
aoBc1MzHgX4ERHL5UT44LmGQjTVU1IiZQRkMJBFwo3xjNIoxnEfZgO9wjFTuG9MOeRhYWdxlLE2+
lMlB8+od+Zy8YOm5ir7jm+sQ5vx1Qi/a+ZhbIA6f6Rgq9yAkYwz+blFOlOiXCC7RdJ5eM6/MCKRe
woLSv+raC3RBvR2y8Nlh9dNRtkDS6BCjduPriKXAcrV9xoTIuqHB3prJo17btBLpontUCiyyD9/s
/AiPOAXEDQcDtQ8Uz9S5ci2czqN9SXSlMtHlEKk0ILX0nxJuEu8+2XT5nP9czjLL7Ai7HvE8P/9q
RJu5QKFvfIs067f/oWNK9n2u0NUxSd1nhG+b6iPwA1JlNI5OgSxbknwSI//ye9MDfx5caTmrOI5s
NngG1vWpdYdTG35LHvGz4PUJhG3a683FX0eZzg19sDhg4vfxW8k3nj07Zb7LnBfCq2s0gEByBxet
KsWZ044d2DR1bIciNnjpQUfjPjbI9xZko5n65aFXhwXmMaqUn+JE3f/mCLCCToxgjW6EA71DLWAD
USQ/wM1LjNn+TYdGN02/A6AfQzFNvCg1da+lwrzREce38qk/4p5KkUsiG08HfWqwBCQONwEPQws8
bfoviM96J9hSbLY/EcSVFTOUx9Z5h4jlBzdwrDduBlKw+CyA1f2hqJD2uEadhHBsW8XAbhlQFpuR
YbTP8cXSX5sUvc5lVXrFa4sbswKzoT7EIENYxO47vmmniDk1fFyqCei4xzs96i8EdLKPEpJAjpF0
kuNj+6b4HIRqEoqJb4z9EJk8SOSRp1YcQ7ylWtoULkgavVeA5nXDUHxmqEStCoZnDM9lMEe/4lzk
93HDosszaHRk6xNowAgZSnglWRmDf5MHL/+aJPRfw9+hHzQEQBXmt1uCZA1IxRopInfdOeRoDlzk
eiJ2Da629I5YQP09plsKg4syV+rTk7GI2c2Jm+YE0ESbAsNdR6xd/mAv8WMgB1sTtEKZt7AAd3xw
ypx/dOBsf5I4GWILE0IYvLREZpkrwzHd3YEaltP3Z0c4VdownN0t/tdIIqB0TY7CD4sos7LYLkbH
ffOgKU4hzlzApR4//zwAv+3JzrB3ppDVFlOovxurlvNXFqNnucXK4g6JW7FgeJVdw4yrbXBcQYTp
rR+8CAq5C8JLsu+ol4tXm7FPZBSzMOtDgrhiXN6dA3r2oIMAiviRiTLAyaIUzz/ni8PyIg63+ADb
exTPEkkvrdbtfG1TcGUhzKc2OcoSQATk2ffe2CAVjLcqtJW6oAcb+h0Ip72jwzT9o8IwrXZbrMdh
d9R4cH8jqYOtTJazgvcmWKH1/BNOtLOVGW/eTeQqPf46WR++3IHGb0xS6j9+k4HeZm2DjoA7tQP0
zWDVORlmajRPxvKqgkBW4pWs5vOPz5UYlUQwHHR3PCeAHZ4HjcWNZhvkgNCv45ABBoV5MQ2+lXZI
lecitmYmnCJ1DvoyFbP47b7AyDZbTMsGrxERMV7uJMDhNWk97Gvy7L2YN0+ZDChIyNCRaU9C9NeO
318NA1H7h9cpMmxtW2nCoPYFz/PNk/M4HtHPyeiI2DgBq1CkLUxvfxGYHGdmgzlLNR6nkQZMx+jN
5DDyCKCTjmFvOUvXlGUCc3SjXpeDmnkUefOVAZqEx2uB2aTAHrhvXvkULZ3TBfxGHjQNgB935L6d
bVvcg7JcS+gx+za0asgu1jfl/q4Gj/Pf7fWl2WT+7oE24iEbzGaAaRaar5fbqo/eHAC7BKCt+q5z
DCIyFcXlWdumnBjSbGhUAi6l5B7ETgXN6+LETMI1A983j9tTWqdc6n6lXBOqtmUhi5T5gZA7X9hQ
HkRq+5FuvS1Seq9tAsjlM1TlQq3J/zaas/PP8NhUFRByu6dHHYuXR5qL77lu3ZoPoOuzzTScBCPu
Aj6Be3vYuF60ZIbS01fxJeHzEtSVIYn3+vKfhRQmurTKS5X1KlhQzgWhlELJK30bl+6Y0KVO/hbf
GzfucBkNZ0SAI8Vq9K8cQQ+wDbuGgxI7Vm4AnWpvL75xfhqVqnkyo+U73HwH0SPR2MTdMZRSNQR9
9taGHonhMAB0fLkphs73EJZQKXCMbw6lYmpnyhjzjC5beoxGoGKaZyT59i5XIJaA2w7lK/VN80BH
E8aIygnxD5EN+DKmwcI0+rzr8N7aXR+WsYqp/8HhSuyQ9to6aUP0dmPOCkXZR+ZptuSY1AHHgRuW
x85uOorZCZKeqftQwYyfMijU0Q9oRUEzAeJUdw4vd/C+Qxvz0W1HIy0BFX7ZFDJ/AZiQjOOqT+Wu
TgPjCe8FTFOuhs1e4A1aSNaxx1ZQqbZZ/+RdBqZElMxCtWrorBVc8OP9w3Lt/UlKhQ7GTiwsWziM
jWecGfbV6/3gfPjOYgPg08PJuoT1Ur1iq9TTGOWTB3ls5E99Qs9QO6HEnOTygDklxe1zRrChhIyW
uxZwqVhvUeQr2xromxIuPPYrckNhEx6hKHm6iJPgS6um9sLJUNl5MsUzzdHd3FuNeblHLLGxx+8I
8Ph0MuYnUo/WDR1dpZ4r35DrRgOtF+sCBBQiVFmwp2OG9potrjS4qiyMXcd8hMga0eh8on0hhuSM
mPdKPLRJLJO/0lFzD5nwG2vsnuNd/manNDG0wf3l7vI9focYq4kJjfGXUYTgZLJgY7UsaWsBrnvD
yW6N1gEpoJZux6GUNPrHHaCnc2WPOpNKzDoDeOAKmLkP2ehwixOs3/+2cggpq5j6nOI8hlczQ4qq
aSAi42UJKlgDk8BEWcgKtH3h/FWEnJ1ULzkyP6JAVOUuSWbFMTEcfMaqNAKuvXtoXmKPUuXLXile
CLTgXNodihv6i8Ge487YVsmXF35fd4gh6fvhIsHdMeJZT4kCwENi0cu7tpz7C02CGOnITtLsX9fk
SbhuKXjYXOOTGX6Hl356LNMOphmHLa9zVo5g0cjyLrP7DnNTov+Un3IRou9pUQv2HJ/cwiWnQ9i8
O1RSiyM29q179fjyIPipts73W/DHC6DnjiWJ5+P7xFHMdkbYDZOsXIAupTIGI9H0hSNgA4VOHwGo
6Yo9Vl9mobgfsXPFTBY/3WaGpMHUB2vTf4J9KuDfSMgOaASCPpz0dAUzNCzH5ubSm0a3GwfgOWqs
BBbo62SbUa7pYUX0ujNiC08a4w9nztVn9fkv6lv+E674bVhtctwLIw5lrDfzRK89Zn6XAh9ydct4
lq8YBC4OBGLQEdk5gTLdwLFoII22xIfh4z5XythJexA2nlX5JBrVV1c0bPjLjt/bZ1AJ9kAaBRnm
Wp/Vy+VQ3EWRAQ9/5X0mhde5Xs+VHuuyrZ4pGQdZtQ4NEQFPNQsWAdM9sFVn9JUJaB3gkh2OOp8f
7EX0ulJcAU3guYGsnfQr94Q6C6w+L3IFdSRCeia2MYzTCY0z5tSiLQrz8RfJ6DpUMTeyn6bmi7t9
ieo0+sTa3OpBelUTu2HM59DBzzNX24mT7p9nlnCVm+MHVkQsxycRvSNnNJA+Tgc5xvibteJkbz68
CreL/tnBSybWb6QaZlrm01mp2oSPasli2d1h0KK849UwGqqSm3ioc0a7AckFyqXjSptHdOYEEJ6R
WmSvPFGq9jmEkYw8Lnt/LVxWKWueVZrfub3YLC+9gqUbBXh6HKor9rYC0Kj5S3urNmD/jhL/1U7F
BpP846HCoJNTc2uYMwYlrh5aAQeToRGjBndnfpvGL8wq90Zpt9n2EGK7XxCfURlfaf3+uhIflSfE
w959tCzXAA2NBnM6eIM6XTHLyf0WhpU7JmgogxDYBKqpcdIPlfgVjIevwoK4MBfHWJNEvXZR5j4/
VK7+sm6s3wXI+7mO5Oz5u0oyo+Sb8sCtWwMqitPL5gtsvgpaNq6gPXJTGrZEIQwJUCqBsni8ovW3
FPeZC4cw4DjqKLRYFr5qVc7Jwg0t3P1r2ZS2bGEy7syBZj/WFxIhTg4RFdMk0hJo9Pg+rvdmR/KR
MwX4/BdVkVLXmGMq2beDT24pVn/WADDwOPcRBd6DhkzI0L9x7gCM0s7HG1mYmnzScA/FOflda3Ii
y8SiF3G7L4UoZ/dH69u0YpZA60T/9a11+iNrpLUc5Mv7fHz2w2wSL9Aml+aDvzy8ARS206Rhpw4D
yskTNvCxOCwPwLfWIRv8E1OXTpevYuAanjULaDr2UA+gU6yOGv66yXyhMvuWDcWtlK8L5GNqDatd
CW2ymUsZu/R3QQp1c2LL/BqzmovaTiKI1o02JVNG2qBZFgVOTINxr7w9kEyRQghlw6JeuP8YOcgu
HQDa4y0UcTZBr+it/gOOi/yj3sljfcrdnlG3aZSHDqJoSmbffhwEmkPqev3iy577QppvW6u+yMJR
p4Sqtu3gjZS7+UMr0PioNXPunujy+yBnm/T6Jj0bqacyA4htUat/5+oSYKxIDBhWzh4EZmGVVVul
Duqwbrm1EtRef4yQaMmy9D5+3fe/kpFiftXOXULHgnGGF9dSmjZkuUGJeOfRLhp0ajmaETUP4xC4
P6zgrYHzAkaaqC/Ypo6ELDespU3XkPeL0c2qwiXNMZ3C5uD6e2q/KsdWqoyVy1UaDJ0YAT8r5tRn
Yokj+jqEyPVYnB/Ium0CGX8pGvBBEteMl7pQHrJjUBC7u5kTE4kP1Wv5M1FuSKnmNYcnORDeLut0
9rZf/yC14Qj+eJ6fp01uydAu6HMs6dMVueIAGYGkteHwwmdEdmyfYYhCXqySXYtgmD6Q7Ih70hq8
IDA/rdcBP02b8tEZRpe3SOTMbB26DIyA6e6+ppcebbX45KcRCZf+NhMoqENE5bk8rMoneqjaWVcO
PTgfSxyh2arpCICx7my18gOWaUKZsdJhfRwLijypdI1Xrxnco97It4lQeyuhzUbw3KXorMJge6pS
2eON/A5rWVopJVMrjF+VZRBNZXV/l4UuzltR00OaAjKL3nyfh6Kw3rqB4hGFuOHxh2CIi0eT4M25
FtSpStjHDU8ATShK84gXEPBHDVLj63YlXnbaaWWgFrg/XGPgOurk+KAHgCBLswcMCaiclrjE2PFq
6GQpT3PYf06jxfGfd50I+y4ChtY48wDQFNwkXFU9/7opTiLIrFmVDg7J2ZKS3srijZEKz0IrXpW6
ar+5ZW1ypLV5DtvM4nI1nsrHzbFaiQWSBRtexY35E41iJuJzoKWpjjpAu4/WBUWOVeVa4Id5gO4c
ebmN4dNaXq95LpQT/3JoPES5Z6evm8DkOsCCIDjQr6ugoGcV+a7mXVbwuklaLBcVpfaqHnQgPRiy
vchUPhGOSxwpmgOY4mZFDlIrh8SlxS1ASLhuXNNsx3kZ8MP4iGAcIXHmOokcqSpu741D0TnBAyzK
IkUY83q2GkrsYSJMB123A4NyUsLssp7hRpPzRtWLUtP0ihA6VAm0cg6CEC8aVfG4XQWkIbTm0HKR
liFbTVMiRx0o7ohIwGXclG4Q6xnPKimm35asgtfU2JriTn4y6JhTc2kZXlbHSJYCCdpcvpBIJrnr
EUAOVWhiPvn6GQ4H5aMhnQqvRKpdjHoasDN6mKt3IJmx/0lqRzwopgW6nhkvnHcx6fPZ1eL/U3Iy
0d+LQyjCkhezWO8S4Y/Q7t29pyAMRVDsyBeDdSJTKdkmEyhqjA+I90YisDOH3ECjSioi2nMCovYO
YY9Lk9fkGRrJYdqJBe6vW3xkN27/8Wge7Hww3x++W3E+VzJMdu/Rb2bdb0zZve1bWJqEJxw/ImTO
wBtvSZTvWDo7yhw7SSfF4wO+fXSlfSq9rgDprHtds7kMHh5kCV4esKK2PJ7PXIScLRZVKGMx/Zqb
1zReXgASX9yl84uV1FoGaNskj3m+FzKtIdkB59EBiyvBaZZD3xqSt625wtDSAIPl9fc0OkY+GDW8
Nt2CYeq7flDbZgr9O7vDRNUWad9tJI0eZl6hQHaGtV74vKWcATpH4Q0Ry/Gd09kGgaAVVFIK9HAS
kb7Tcyx5SyYA1aLHEElt/pfSkzOy0Ar00eh6v2NCFqCStCWfzdrBwgtG33cDDzFYNk/xihstTb87
SojQLuF5zbL8QCD6e7Mer3RHvbV7OEdgCgYX2B8CEpZLDSpD+Cl9j1WDc498MJT8UcLK4zN18Yc+
x5uXR63PGapg+Y6PKdEya2OUbLt6cbKKd51MnC7dDKYR1iL3o+VdXs8Nts4MMmHbKGYrVZgE+vjL
STT49e7coy1+PxuXej2RGk8xiExANXZT2jn8fxnxSOXiSMJ1Nefl9nlXkPVAc44TDE5OxPApSNoO
fdf7HKxY+chf7zydNYt2STAG59ZVxhZhCr3TPWQiLcfth1TFIn9JQDa5ITMB6+o9rfs7jPtNSkZV
apLycttxX8CcO/J8xf1sk+Vv81u+/1VKzZ+Gl66KCLTdG7EvDrRkozOytfPVVq9+TzdWYXGczcdc
IXRzt12fbFlQOkCNJNsFTgry8DXzz82vqZbucTTS96hCl/bVdnPPYDAWuEo33VZl9smDUuBz68r1
lSmq8sohUR1ByYD9dQXRkOYoYsuQpwh/ib9jCIiVasL98vSewTg3eOYp1qRIjDwR9QwQQzaxwxdG
APZ3Qyl/SJ0UEqH/0AlqdUmsY5ALOfpMDRQVEAAob28c9GBI84NfbPs2sfH5bbeVM0TYZVXje/wQ
3k3CDyHyGYof4ZfhK2l4HYTQI3Rve2CIDsc+SWJ47b6kwUCwHTp9PsiB7jCTRXMLsgk+0orvFTHy
FSaHnAjVGa7oSrZ0FYPR5xI07NkX3GOv3YR10RfkzM9ud+1wSxWZEWJkbO7AfU0IKIdfLCsF0MO6
JAyi9MninGoh5VJHbrwhCXdSc81CjPObT9eojETfLAmFMtLJmZ9zSZGtW9khtOEJoJgdXpZyN/bI
x6wjxmHB6byT3DUL4hF+r1ok9pbU05WDRYKBnBo4K8OhsHO7El+DTvcuvPjmNcbkhzLheUi938le
ZywOZkmnfDP27JrQDnFfyoFGsqQj6TYtHAJH0f+UwAbAh/TeU42IFDdJqwC0MK55b2fo48VximR9
bHOrqn5X8bbgPtp0JPomOuFX7UeOHbs1zmLv+iBCoyWM0uVurLs5MGOFf4fAA5+O5ReYhs7B+ZuZ
GqYWpf55fcVT4wIeFbvvzyRwRBpshmsx4ndhzqHAK3AE9LexYuQ46psS5S5bCeEG+FVn5+ZLXJRG
fnpEu/BENhjfhV5pmqDvq3sZy/rISwgJ8gEtvwBGIqxtimLX3l55NeS0TTLmSmGM9CgbRFpj+gYp
F4HY6ni8x3qPi5aHFKFns0/lTAotd1s6LaXUVO/7ibwA+TEY0sIUVI9yJY5fR0jMk2E3WKSA86Le
utZx46CipVr0AEJ9b/DPr5fc48QPqMHSxbVDJu6w5c3v8IOUhTnZD5I4+BddR1lTHW3OSJUNcods
NSG/zbHwsoZ4ZaqLV8f0kl71pc8MA70l8g3CNrt/LJF//Jm/68PqOvRbEIPj5bNHxjJOnpfW+z1X
UUtJDVpdPC+nPSTG0tbdCEfpA63RlT9E7KbW0Wtu7ucH4ayLM/xtDEe8SHo9P9xfCv6np3QfWpso
7AuNw4g37CXfCfqRkCU7VCO9i+xmZCAxz4+lc4ILt9oH4lXgCfm7e1CQVFxIRCxxeDJAeDXbsWuZ
ipjf0wGv78Z8tKKWddEOtioI4Wq1YNS1lm1Wr9ejecO1lbJfxFvn1wing9K/P/aapCf5KInUdaxg
wr4g5/NRRAQ1s5GHJeHw9EzqfssmXPfv25VkhXGJJvLjwjNFhMZxiu73V0ZXmSlrGVxuiJW8VA+H
4GC3+fy5xUUaD2qh51s4VzWLWEBTJRNabvDdZKbcEbRoqS2ChZt5U7/ZL1xsRVw4bM+nZyl9UBYP
2sEntmd+1w9rIxJ2ph0dlaHuOmtvuBEfmASmv2ayjUZA2rbiSDt6lpmxclpo05iG0NMPvue+xIq9
b70NUdNdwg7qeNTMHTvECEzHWHafg43drvEdUmxgWQjOhTRk8Yh+dM/OTeEkn4xHbj4FxrF0qsrq
msYuZ93pUWk8wikAZGvmXTuw0lFF5QNhgKjUdRiF996yLt1uz9JRscF0DgEM7jUMkESEyp3UpOtH
sniGmEaStzFPZZIpYkeAZeCJmL3AMbcA6i8uuV77TTIANL7zeyLZDOI11/pFGAVJJZuet2xTLKu2
qpRzbcy4b81rQwoMa71Lf8fD7UHdcFAz+nUEIXg9HPohSostB+2voA02AR/iJqlbav33Q8lrS4Z+
ww9Bv4j0lmhbCgc9u1v+vAOuiPO2iLkcbNmag068QyWxEvZDcG1EiJs7UeKDWU7uTGUwHwnX15xF
JyI+ZJ9H8BeNAQO7AkfTNs5GlujO5fdUABoGqGWyo/iOaG0XhXi9WDbZSz9y6wZtU1Qlj0hz1BUK
9YtuxiURRcmjmw0/JA3BRt74SmfgbJuvKkUwPKyXP3zkFPK6BANb1zwquOL6n+BFnj4ak2oFfyxT
/kEbFWrXJY1ZprHjQGlSbQHfkC4Iu85E4ZOvwRxTRip/69ncdfU61DuWKr2sQ2il53KLnMlyJhYB
e5aCmfLS2/6S3ftG5gd4pozOWtCBMccLehXbze0b3u9ysNaux/lKpUGZ48OEWuNktc9dfxDaw8Oh
As/7sVimck7ewdJXWTuFnvCYhzUCEWbDJfEQ211Je3PuxHg/QX7jem/ShQr9m0ycwl0GaSxpJ6aw
96xzhvq3WHR3R6ywTXiyVLuoPnc6L4TrKdR0Izl1ppp7CO1uOBD53ucJ47WNlssdid/xTnOkxnfD
sP0ajowJ91ohlpCXNwUFYkHcZhJvTKGOnHRkKrOFwQHGb/qmsncDc1n0SZAkjkPnvotfYM29AXUN
+3h1oHBrN6YcziE9eADmfHj/2XfE5o6Lbmv08tU9rlcGywzfZWtYyE+BII5hjND6J5TUtPrIIhij
52kemEUzKrhqy6Z5/3/oADYLgIwrMwrkOhrAKOgcbV3v6ZR4ipOjWKShvegjFFc85msAGX0DaJK+
y2Stdmr/yRH605P6qUtN65/noET5cvG0bnBYQeJA0Gm2D7mJ0LPn1YhIJcRyyr9HfB+gLUiCsDbd
Og7kXVUnY89tn48v+R83hYnkNvonKieTs52hk0tX1R7DcVTAb53HsL4CvhA+dzy25qMmMFyWjHiE
azzZOF2ofEt4bWAPv20Ruqd2faSikKICGcSSySpuSheDri9nf3JI4i4cwzNPCs1TdDJDLbqjQMjr
pMxbPfh4DVoPXEaJ6XgCYA8XRVZ2bkNAELWz7XLkd4dYVagc2O4JVluzaD64jebrwFruLIm12qF5
OnyDZfG54+tYxLkosKGMkzPhx9dfdWVM9yk70IRUp149j8ftYXUSg93afhKvvmriUfNEzJ0ZaYAo
/tmYG4QDpFAP8llY1lvI9KaKppyFDKzHnS/YHjA3lxa/9bowVtcYYA++UTNT8FMOvBOTTuOXufoX
6c63g42ce/hhLg5a/yl8ecgun3b9dQexH5i1RtCMCmOAscjcm/3uRjE2cs8LoeB10bdT8E5Hr3CP
tu/qrfMMMYjnJxyo1SCMoGy6fwQgwosLok0TUZ6PqrAQEkOG+uCTOhouI+1fzp91AjcKv61duNt4
QBshF0DNsdrmrBIajSzsR2nRdQ+o+iX3560foxKgfz2bs55AsQrEWrzWRzWpSrvWbgxUY7GHBwuY
9/9IJdKNb9cX4iIO+zNj1VbPU1YiQbuiX92vEdnnIaTQZW4Osl4Y/QaFdaJMDrxZALVYCQSh9T4C
4n7kqjCKeTUa1PMdi7wnHsbheQTZganACLj0v97Cxv1cj63m0IavIjV9+rQlVx03ZLtpWKZ7U/cn
ShbLb3RR6Jk09qs4bUSf4FBVYDso3JHume71+z9x2AyhiED1N7ZIMhMfwUGS7UbJ69QEwoQ2D9Jd
rccpC3vdWkV9JnmtyWj8v4pFoWZC/oqK3ghZeVnRg79GcMMIdTQgWMweF1WPwVqP16qDWdE08s83
mrmf9JmGapYL+ELnC+LaLShKJNsNw6ZXlNQbvRBb+eC8ui4MfrUdfJGKSmiSN2VeOu2WDTA44Cvb
FpMerohoqlDcqhhwCAPC8N3Z+DTP9+LO+uHBpt/t2XZn9h7olRbETB6T+egGz0iRARNQbfbA3boN
LHGSC/l7VDz5b3Y7Q2CQ8D0sYB5RjEswaTVVCxPgYVnD+fFKL6getosn/lH5GTpcLWqp2/r2YaeT
wOo0FQ5I+rWhvSHM92SebmQ9NTvRHeF/WWfZCn9qoEiUwWvxQtPwwHJuj9w9A2dJmbt35YYpfM9I
yKGK5Hjv28xTeVt4t0uJGoezl1rl775MsKX+2H810bvSqY4BQqbENXuTOfRQMh5xdP99QfU0ICsu
qdHa5KnZI2VAMns6wAP3ePlzqt0CykGZx83v3QU0Q3PpowwlYm256F7lAswx7oaJJL0h7a11vZc+
Ex7UTXyeSFhlMmXmgBLvUm35sOyazLK2B00/BiWidYJPxk6MkRg9oYQyY/3jHzFJfzc8qvJjWluR
rEid1XPT2KraufDOOc0O87JVIZiY0KaLLwRvE6WKXpR6Z82bTo+3QpoH8fYjc9WEv46G9Isu7yoB
/xaANJBJGaW4h6L4xFWRw+oLMlXSUPVlMLYPYJ/7MYlVlYz3uwIXmciie/qEXlBKZKtalg11UVyH
tF9BGmmu2+Px3yiJpD8qyo0fBecVmImWxrMOvHtBW8BIP5UBObjxcR3R/7CUzOwXlD+Q3AUDVnuw
BmcVXjf3M3wx+3OTUUqBVW7tMdyyhyWuotKlbfje/w6nnvntFPHXx/qJ03y41Baf7YpPtq4Hxaa2
W71BziQykPKXd6533Vj4fXBnpvVC2eZ/VgKXWBxVkWF233xIct8l2L7ungTH+pg7QsFYOWrtunUM
qELI5ncSs+pQGV7HQQCK1UAvAey5G090e5kkMqETrklOrVAx/qlkbVJpMnu4yRFnM6k3xLnza1Hv
XzQxAN0dPGZDezjPv70lGwlZeadVNfSUYv+2qtIHDYMn76itQPUFhvjfWyk195wdYK8PFwi1vkHM
RGDqewZGqgPdYg2tX+qTF/XD+hCOJdpS6DXDk/ETmR3dJ9Pei9zkTjyQJdBbOQs7UyInQ2o90LaO
OTGOF6UH/wA2egEHJIYCPgGIRdKkwBmcnqyKLqye/1AVmrQtYhF+nMWpupSbKjz8lcoLOrGm9EhL
kQN2C1ebuDGrkdZRsJcH4xNkabMzhd+PkRJeIpZjuW3BkHhSP3HT922BH9wWmvKQUTjw43Ic8LDo
P3sBd14UoROABJzDwJDZSYUTOvnDlgswJbwsG7art+YoHIRUpTjdclDker8wuGZGLsMiZyvjtF7o
GrmIl8Xu1Xr0bzUuNgW2DHB/LRG8M7DRFaEkIxUfQ/qd2OdqwwEHNMfN62wbFoE3R8m5IwIW4E6U
MWOjaBLhop9+EU8nw0LgYbkRvBctYTsUuEt+cMFOskeZyLT+1mHq2ou5kCTZrZgKJ39UUL6vpFsT
0E3s4RMJ3eEXjnWuIYNsPSYSD7+TrcK6tdJj4c8Awk5Z+FPWbsmvHIdI+8l/FwqQ6m4/0M7/JCAE
bL+YLpq7P+tUoJd3F3g21XISNI8Bcs2A5JUn/0jb22cam5c45V1IiUKnaEcfa53rJcHVYp9tDfqB
cjwCNsz6O+EsifWVAcikn0JXjelNP7SuxBU/QUqVDBn+OIhGbbBSj4FmJunITsA/cn1rcYpbttJN
MqmdfcSwU/rpsm5Fx+fEV8mEqxzpD15HvMHjhIfnbT37PPbbca3DfVD4lzQPR3PDkkvoXM3+ywfo
7vRHJ4qCbz4SvP8/80aRFL5AE+Q4XI4Z7XmaKBdna/vn5u2aH7EcrA5Ev8QV8Ce25GiEDZanWs2g
eq68dmMcMrN5QpNecQGvuMfsSboVyhDivwNVbpfyKT99XgbEOjMxRbkZoVD+IcCfXxbyZsq602UM
CherF1IaEWPIBkz1bAKBm55rJBumL0dilbKlU52vNYVUb0ua8SYgjk2hZDadFFtarTCaI3Q5CKr7
DL2yKOH21bwZFBRKrINhgSKDQD2xWUkYk+9xE9bHO0h6NSFugec3Z3832tokwqfzLDhUSFEo3uI9
3lxMk8FHv1a4U/G3O5+2406dWq50v1T9KafHwa+70syrwbu5tbmS78TIwUNoxUWniUbLtrxXbvT5
v2VaXAxSJ8wyRuUwBLgx5eaW6bCbJpncnAaCAfl2geyLyDngARvP1mOe03k55nyFMTPk0W+/F7V5
wTXntxTEgzF8hhLDdIuDPvJPtIaZapU1QRC4fYQl1KA+okBVGFc195d4xp+P7EpFVZW21K8wkNFt
MbQSIHfInDCtmapG/8qxN97vCwovID6MaXqivf43+KJzumTScOOeHGQlS41e4MAItG6xHJWMt5wZ
qSKAOuCTq3FDFx6uw6lifaN6V3JN0Ya+5qzbqhofRWt6vjBSeGr8U6A6UCuXrLpqDDwUsl/ZlrxA
S3Bvj7ApnikfmyrCv8ilfBXJ5F9q1IpdWJ90qzpDLVkimhuR9zo3I7dT0ClWrQgKdqrmW/qCcwgp
bAUJhVWxGhjz2G2n4Tu4EUJvUUQOseAqxbmgjlCRQuiZ+LB/1Wx7LeKKMj2nKioRKiV51SR8g72E
8uq4KQiYxhPqwj+J7S5HnNRvmRXsWArlLyt3qBm6/S9V34PU3BIqkkdlU1V6yMBVHfBBoHO18Cob
DXaitz1SePCqixSxw19HS7FLeSUiJ7Tg/YERCnxyaWK0dFciRCk9bc9I6FoxyrXtCcs24tsJLUT0
ZKrGRn/Cc8emrX/cYSGqWzzbvkGDDd/HqBBlJtBSaRO2avDusvelEDnIqr9edUdVis+O3BLHIzmj
s3xny9mFtmKfFVCrKOcnVkZ+u7NOUo1nAlf97FlyzEd7nMuMIjVqTBrKZobnbln4PgGx19qQzluU
ofEP8QW29AiQ60xtjw56cJawDy5a9RhA3hA+uuvgXB43ABfXGVOJaSIFgKS42E0MkntfhdeRyH/L
Dhn4R35VKHTYG3PA42wsyeSMhZ4pw1BDKya7sDSr54esAiOmZfFrdKJ4nTOSLD0xU295TFElDnlI
4AgV520ARw75FXJ00AIm+9im4+dW0OsiWRHZkt1PSWTcz59/9W7bA6v80OPZO+uT4r/0GI9/IxL/
7j4OvBrikl2dinstuXXs40coEbFoUzYvTPS0IwMVBUX8dO+XktXNfcOfl9PWadrDVfN7xN5Amqd2
9mRVdofHcJO3huXPMGgd5ak/BbNhn0tX5NxLIZ7GFGtVhbAERET+C05MtXtEfVrkQzml6BcwjBLb
3gYOrX4Hyb3FG2iX
`protect end_protected
