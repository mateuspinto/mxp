`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
ZI2rMgHSa4MMkJFWJs2scIWulBvv/PDoEl1Gs6KE9KMBUWzhV2zTRAhvsLwiyzarCFTzDNwIZOKh
DEL/9H4Bk2umeMk0R/DzSJZX22YypWaGu7ca+IrO80N3rTZTd7IRPyBsC/ISiUZMcz61uUey3mlc
DTbUvsh136/WEU1rHn8s75Hp7KPNrKvxQ+2BZBQlG4p/D7E4k7Aibc9STkqQPkGbzQ6MDBKL+Feg
63jK5vEZmBUgSNeyGNkVblSWlEzVMY1TkzedS5ym8gBlokzc1o0O3ldy5XPkWGEXbBu8h9qDqDeF
1wIFmMoX6YwDc/pG23YyrzfJo/0Kk+Ki0k/R6LeyIWPVzySUO/dv5Vo+1ACPCgMH2R3rtDzD0Sj9
4H9GF0WGAbHW0eSILoLWm9t+QnOr8UyFl6MIOhZIF2SILkXpGpV+FD7KA3VcyfrAq4tEcsh4WGG3
4w1cBKO0wWayuXn+RlitaWSzkFW7s43ECr7XUXwKgFPXiiHgF2YwJNGh6iJLirN+vbeNKcWEe9+U
X339QOuQfdCvtH/cpSV7zOg9ezpXAIGlFOe5nrW/pciNisCEX7/C6KoJBGEmZKfbV91snodMheXo
c1TLvN4GTA/wQKTaoMLXklReNywI+CB65jhTZnR43NOc4VQtW1Wyk8Jeuu6/1AfT7WTlxSI4qPBy
E/oNiT3wM+ORJY0/B96RNgViwcorJZ9F1HvaGnIK6PHEi2S7YAkZbFQnNO9xL8E9X3spMPMy2tDc
FFcPZlyD3FlWSrX3YCVuyEghoSZNXejP/AcUQOIrVzfirWLDFugEV6wIiWu4CqE8K3nTz6FJNrnx
j+4l81PJdfey/0Nu1vqiZYbU1pHruJCj0WEX6k2pvjLhGYpUKpbjP9d0vuz4SFQhlxwkoALKmi+M
2kVwmc7C3dn16qyR3VkwTWnRZpG0H7gXutfsTNLFhZY/tsCH4guOTSkxQF/8Q4a5pTSIOguBCn+/
k+Pu85ZE+8NpK4zWC6pU1dJbmZXvQdlcaWIQ7g6rfYj/aLC7r1mTuguWqhcYALmNRWNMibnrGijH
XTEBbPfc9vjqM+U1hfhotOXPxU8SW7TEHfuojM+xjLG03YX80Wvkxq8Y7blJMXvUdCzCrew4dbGV
59W9DilDORu346kgioGZ6C7/42hcpHMmuuMdj2pcnJOqkg+6q50OmhFj3zuxeJLawbOmlUV7VnQy
mXVdpGZaSXFKuZ5CA9b57GsNUJ1+P/UiwoLB0UxnqgbpAnqiQKywYqjn5jMEswbuAa0S8+Cn/LmI
Op++3XfVmy2ZeBZ6hD3VCRbObS3jsYWJ5flTqVnnwCtca1HE2ipavDMQrSGMSRJpkb146dVFnluZ
6rnVbIZX83cikAZHVfd+k6YoVtBtaloePHXniemP0VsWKUrFxbO5893LazJ+iA0BtFMieA48kVP/
ux6AcbpI7YLtXWrDxALaZ+a8bFlIFmNORXKrSHAkTyDKL+ji3LpHPR0+CKawX6iteSNH7IVA/cby
yKU74AK9KIexiWkbfvdOkYVi3mrIEO/PaBrQTzXYz5bOQ62iLuPrKB300LMnSF/Kg4ITt2RUa8mj
WBi5fpWjY55POQed6eGkI2r4XzDYe58TyTBUQT3gB4qmpkL2j7Cc15ADQ5bM52v4eiWJ4yzSZjNE
eXOESNy6WkBZGp1meIW6ljpLqofI0TfKy7DVVdTSzsTfSzv22g5ot9RAo86yhL62KAjESkrbGpPZ
NES13agEBbN9YA78LT6Wb1DSh+q5QKkecQDBe+lpLI6y5PcwLlfQRC81/L5F0CWMdYMgLBo0Extu
U2tWmpXBTwAKUFVE4AYAmDITNEFu8PmEYBqQzPW6Auj6XQ6cN59VyxI5/2Nw9Bd+z8IxSyn7fyPW
pW8aUas70yRTz+TijE8avAlQwvxniKg89AhMEw9PrwEimPSeOhoHLUsbnda04nS4dpSkhv5oLEgq
4ycco7JbHIEwl0NIGeGMYTS+dRWHdMB3yk9R3j3HUl76POZToE9S87v57Dk2KmvbG5B+zusPghZW
HsL6eufWJPCfpAtoJF6K3f/dB3tdHHfPgEH5GJN1CPYdtzB1FVvBjIXSaQlCdt+DeBO9cJU2Y9my
2IBOjKyn+LTd36rJx560SnpDajZhUe1mMpWluoyVyu9/0NcV9n0WNPy+sg1TcP5egNnmJ7+1M6Wp
tiXCWO35TYj9+e2WE662/LzHprXxYjKf36CK89hRyHgf/BWXf2UJQfIx2U86FNm21HUAGNfQx17E
P5MQJ9vtP/vuy13Al+svwJ09w/HjORW6E3/DELIFEhmoA44w1Z/D7+PofgK91+K05ajlQ0E/QrB7
ntsIFardBBa7ckVhTPmJtoZweO8f2UQXKTZ50juakkTFksI2LSfNgqNtS3Bg/ttk5I3kgV4VAbA4
Xepy+ur/i9rXEvfe+8sgNRvswSjrnNNtn/rfrL2knRYdUcUTHx1AxTjfDnp7beS77H8o9OlZ1oaZ
l1ego1fqYiJyZhrN/I687CP3hLyA5KfkJjv6gI+jlnY4wLtjylVKCq4Gzz/+Gik0MAhqlo1Twp32
m6o+y89QkKMr/x6Y1CN0fKf0R1pg7LW7oj/qHv8U3l7TRHhCDR+UL6kjACZl27VZIOnF6ehN5gUT
rQRz3T6rA+A08fq2m5HiuFaqRH1vVF7eJSvSsj/O6I2WHIFqmvcOCQ+XJQDTqOb6KLYabTKAiI6j
oRKzlvHpYQ0cfrHJDMJ9sdnTnwFLOtfpcHOTluHbKx6gAuDsI6G/wcIkW4yEhWyKO1mNABuqpnfn
dKRnxGva3CQnDdOM3NIHS//QnX2RsYGq7P/z4L95NbbnfBqdhmqJwjrNsMnZsX/bLj0Kb7Wg2Lq6
O/t7gE991EhQ0EJyWyjf4gpVqQx4aBOeikOkmegQIjHvWCs9X8s6mqRoTivEMOmEAsgtG+1QApEX
o/irlSkFAHn/ldTntMfhBHRAWLeCa6/IDygPDxS8Jo/F/odip/1Ge8qStny0yApFilc0HuBxIJUa
bk+xS2/tJmpRnxc2EgwLr+myeHmjlC3Xru1NHM9Bbqx5J1Mo6UbGz//O6aNwLORJ7GrKGk1EvkwY
rTjHrM+jZDBME0TgEnk+/0Pjl3GB20fbovrBcUh3MbMbtjKed9mrz0wd9FWQm7yA67HKyABLqp6O
hUrEeGDo6A3+nZt76QzrfiBfNeqhk9+KbyH/8y/SDWIBh8hBH4FiZ6ovFRIXRXlSZVUmbzeYumPV
Krkh298r7pxBK/Se5a+/QRNUrQ0viQUg3BIuWQ1v4rJ7hNVAd5YXTr6STfnalzh4sfIUAZOsDfgH
Fg/tD/ObxKCpyGUJBnDn6vsqcc1/qrj8VnXUFtHItPohXxPmGUBcAXiCjWMueUWIwdZMCXw3AnrL
5aSeWjJca1zmJvDEZtsEhnXNs+aOR4BL5ZGLLZAKbaADA2Pyc+FitNV1hcVZwaWcMPya00ox/mjt
Bl2n81fP46fyDKE8xEFwBVdCcLzmBcFL551dtfRswHijKjypIhOQqYMiVQ28SSJbWxSOI02hqlTx
vCywVNePPEGrgBbIphu6cxCM6kEwg77Sbo7ca8loWfgHgXQZygWCrTl/d0cx3HMO7Q/C8jfd68xO
43ayruhedLCrwaf+aIRMl1XzYXkzM/cKe8rvQMsoTR3otB003bTn+LnHxdqgSdukTjtAXV0HIlIC
cpQf0dvsBVctr08UTQNE3+yKhyqzkkiiWHnA4VFu3DXFJQ1aTOBhLO/sXPo9NPA8X93YbmYFXdA/
kIKRWhSd1jy4iit/bnU5FyUBxxcjuGDs9dE6SBf8ba8xZLVoS0pLbQ9G5lGcFp+V8d+kk2hc40qx
njLt38A3RAjMPzbqXQJRxN2DAxMmNGN4NPqOA0tvxPaxTYHaIRRU6VxowyWun4Em1mNZSawE2H8j
xlvfuKwx9n9fSKSHGLaULt7SYBYMNH8MkwwSog63dKHcSDvrlNXng8yNoexy+7udD+9PWr1H37/5
TYLMCgOQX3HyhcwoxWugTEHNAEhnjjsaO5YF0t26m/pElSMaksB+6SLYlZOkXssWiAxGN1GvTbCt
/CXfpW7SD3fdW6a2d/nlq7Dcp42/ZDApw5jcVEeLcTb/ES98CraYzsfXclnYGg1tw6QyHxWvYK8N
AtVhH3fa5RmYKiNThrmXvQ+CVcl27bE5qN6UQFCjc5dHqm04FlF4fz65LDNfitSG7xtTbw+2C2f7
Qimo53nXXWKUGZWh84qi5DwWTeGyLHdpogy1ZFVFEH+DFAn03TFfqP1mYBJLOLS8nDSZpTAYtbYY
aadJI9aqwWxkwPzNM1gbA/9ZfcSQ2j3vp69O4U1V2rYgMWufuD6gHn0KC2/CD25TPf41qZkcDrwj
4TZkeiV9PSZ3UOWyhWTIpmzhhmMTL37UffKQJnyyFLykV3MrMXLO0A3srJFyEzNIrP0KQ4hSgqd7
EI8dD3gzUkvO7vJ9M6aRRH/NBFAMI35PYBGCWcyc+pU6wBkjFcHsbMus6x3yoGLPT+U1qq/18r0r
GmW22I2RkJdo/+wA2MGIiEhTCLVf317VSEf77N4hyHaRgKIRTWj9VL24l4rgAR6WhLC+70Iye1ZN
FNunOtF7P0wsiTGy2kHrHBldd2Z/cDNuVeHVl5PQA0k7erAYMlntJuRChVHyb2i4ZfUm97BgMLyt
nhhL38z2erUVb82u10GEEsjP2WDlQeZuEIfrS2E+qpQwTcLDMne41Pc/sS8rKwowejDSFqfXBesB
KTFU6xCFlf7CSkxyOQXw2z5X57t7qfpN8bmVpCDmbyNsAgdqRuyFiC9garQp2FeZrqmY10/ch6JM
Y7mCAsaGAkRf/6JYjXIwHwUluEM/OM/3WIKE5AEz9r9ss9hPwKNYwU3FZh3LITgWSmrucaLb/Rd4
je1A3KkQyr89NFGwaJhq6wTYwRf7H+ul0duCt6Ivw/Jh9eCLnJ8yJYnKyr93DIUsEuLR0KEyU8w8
1iL4NPb+Aax2eDh/mr/ROQVLDQTOXCGVZMnNarbFRpdYryBKrsU/x8m96rFttaYZNeU28PilbswT
KsKkeG8aJ5wVtX9RwDV/kzw0yB30WSqZ5nHllwKrG23RKJlOkWnaw79knTH3zniT91uH8Odqf4da
kTqS/7amJ6ESO/bSdZxt2zciHUKAUyoN2qw8W+ii+xQTYiLbkEhGOSkopsa6CFn8YraNn/Xo7l9U
SWQnEbIXb6yCVkgXqnQ1U32gz4Ucukwmg3jJ8sQpjUtneF4hpf0yU4YVK+flerybZQLQ1sQoXH4w
QySgU97NNIog5riRvGJrkpb6Xzwv57a40XIVyeq7bGGiVNkYBK2J1ENkISTvHKEYRfbfD417ZVRG
2oNGKfhCTwHxRRq13OhU4RgrD5Hssl2QaUMhNa0vJFThYI62ApYAwpaNsR2Ait0G7laMxkdnTVVR
dfJ5EtZC8s/Ff3bIt871O5V6sgC+ocj0jOGye7V/I2va9hhhB7ZFRb2Lx89MG0qC7xAipJAmIh6l
Dsu27vZgQ8fdPLys3RKkapV0Zu/KQzEfD9N2XsAxZAWfRBtpUuA9lNDH4UFWm8nljF49aq5Lepka
6yZLWKN0PRi8ppvGujDg7U/128L400aMG899+SfQ7GSfCgTcJPSyVRAWajYw9Gx+TKuT/BHjh3+0
zsrFEuVq6aHPbcyPn1eCunORU7N8UTbOXprrGPPDbVejYoLA8m93+0lghuhsp7ytJVF8FYj9jfQz
w5sDufzek7iYotZS7ULtwVAFoV0L8yrJdI4KQ7jhr4MZiooCluXFEXz6HNGpgzzndXIvQKwKfJkL
8BoSapHTCu2TRwaB6iVS952tjKo6N5SB6PzmP8xftFgD/ljHSsT9DBHeLeGXhxfIcwLaXFTUuYqe
QChc1Wy1bKYqZGl1n5RZhubpRNfSqafjx7XN1iloMt03i7dRKriYjJFgRJ0HgyUG7GTscBSLOEaA
yBzPTPFdam5pOAOOPSsC4DQrJejMGxi33gLUO5ilKxaRzJfm+3OtIdDf8zbk07rTxPL0PjYQ/gca
nSoCry1jB6GIwzDvAlokZN7JGAYb56dcKXV1O7E2e8qvQIPZ/FFPYlvsJHQi4Kh7tZoncXk9t9yp
EGBLalscIAh39thWFcCpNhNMnI1NAcT+Bmh2JrR9OFVKj73vIZhGNeTCEQjDESbcQ7KfCL9tcGus
fd32TP8W68QFTHRc8zo4W+e5Hnyo6JMESPgcfmU+cFRjNZEh6B1WmrclOdmYB075NS809aHzUNn1
7/LayZ1U0IXAxDUIlzxBaxdqedMKrBoSMkr0nTtpM3oP5ZS0J2ggc28bRilLwYiGuMfZ6ZYxOUPC
nJmdRNJtfQujeVRZ2uk7piMpHqzM7kFgh2PudCklTJJioRWJBcXV5RuNN6ZfvpRMxcnlU6WUnThA
8OcXbJ5LCgt4y0BBzEcPWmOXdlGSlyWjB+C/6yxTb+Gt5ty+em45YohcTkR1gkLscNUVLsttic2J
cu/fQcgyQSmI21LpldUWrLMK4y1D2RpDegK9EZLConZnD6ksPL2tlJ/va6qBmdRSUStXbGEEIl/g
qRl8IZLwXlVinLXfnQscv/VwsXlADS9Ra7sN2YpN5aHb0nbq2CvJCPtDQ4nHX4ddbivbvVC8khYq
AyUpZs4zi/mzNxAMDIov6nfpdcLBAgk1eDTRShQhPf4v4rmsxY68hfcG9+OXvGkxZRgoN/WdcmDO
vovodW0/fyT3LOPMMkn6Osjq9nKkjT7rnZwKc0LH+VShS1uOdj8r/1Zdt9UkKjjl/x6Zd19Jb3Xd
KdOwFssD+2luX3GpNi1oPz7BBqYvs7IS680PkNeqdN4+iKlmK+kfSKj5NbdKJKch5mYkL/00C5cY
bnEzsUNi+/kdH9OPxNomHd/eXcxioG8G3VPE5812vny5su5mfS/ktKYGrUpQFO9viw0HKO2Qwreb
CQtz6HFFV5ytURSP2pBjTe4/b79Q36NdKJVyTxRQJjwoy6enY+MaF7ixrPxUBJ6du9LQlqy9cXGU
mzXdth/2C5S1NmN6DfD3fRCBTJw5XEN3b89/gxUl7SWvKOLWPMNkXgQUcx2fNFdvTfIhH7TO2SA0
ixEPGTzZIpiAB4xaOLiSvv5NIv6J8oJhDUADpq8yuLdyMBebgtwkHYOR1BBqyaLeEvV41WFSCEkM
xmMrg5PG36OfX9s+Zl9rUg/r8djU13J6newCtfiOjrPXOvLDqBMZGivk5ppiXaYk44/TsOm0XT4c
YFnXxMstmMugewRwuSDM7OVi6IbVMwS80bHB442WdiyUYt46MdoXgkIvq4LJBsbYJaMghTRPivsR
7sgs0ZiAaLKTtDUYyJH/G6rsBKCNEqd1T5NqMj7EyRi2SLgi7ZR8H3PHt9llXrLvzovtvLgBTmnL
3YHq7G5PYC05tT7+sObtOp+Zio16GfmrEsQarkTyzkP2YeJD9Z5JHTa69PBztFc7ZtqlsbxcbVhI
nRLajQ2oGYIP2KtSJtgqGkK573W0lMfkhvbFIH8ZRFHWYz0KiutM5cyU5lbHLO4FIh4iG2Tgb/fW
fn5ciF3gL8yNbXbz9KJKEn33IVyOLWaZuaK9Qx8l4uKZ8lGBUCx5pjajA0U3kMG+hPXzqsOmHPG/
jXy1QZr2YCQ8jHC4p9bqxWWH1r5snVWzxthjH8xFjX5DrOeGyhO9HYHBgXqqFl82EFQSV1Efxoih
n+93cMzYsb8nw/h00CEWKOLFM8GYQORW+AIZGpfsAEfIJqcFyjRQrmGhdETDxEN2eU+wTpCN4Q75
5MGAQE8FNMMNuGNwFnFmagFhZ7JKBmNgOn1q0K8CPiWGaaFcr4iABVZugwy8DdQ2gSUd3qCk0i5X
wyfReScKNpxYPpZA1Nrv+4ue7MdejN1WwVv//swgfV/eB/Vb1wJPfpz1nt5XLUI9XTBo4wRHO1m7
kdKZn4PEQplJxtQI/ZXoGubP2lxXuLFU08QUO51K6+4F3W6Wo6mo2EAWp5gbCBaB54vj2wbp5bJg
rgAWS0TTM1eMAowuitA+BppkZHm9ZZFacjVEF0/wxQAzNea1k+cFY2FI1m5Npn5rRhYU9G9Tq4Lf
/6ku0mKqnXK6HTdrvDLiE1S2axkdEmCby14A0C6XsK+1VVCIXjgkMniQEelv+YP3z8NKVU47LsTH
1MaAYi/heIH2FZTrvueThFPGnE1HRkyYUq0D8T/eE68tpMqI6NZKeCKyrkFKDQbGsc6R2IQHLlu3
L+OEPzjmPD6kZ6JU1j0Irc5j3Rt3Dxq4lDeV58whO/LGz9ItF/R7iBKB1W1Hi2frKt6G8gIzKjxw
9nwOjQKfZJPT1tFzFv+eGkjC2z3gFxZkjCR5EGTNGqFH4Ou4dhRLUzzcoEITy1o2u2CdpRXLf0fu
LNxxa/dk9eR32rNaE4zyvB/DjfapuBRxbJU4oemHu9jxmUkNHHdMbd+ufyd3iubAXrgVkfsiN/Ds
X0WDydx7p8mogjiFggkMVQ==
`protect end_protected
