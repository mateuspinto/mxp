XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!K�&�(b��c}?�V8��sy�7��';�`�q�B"#�HXP�ӛ����g����3����'����vH�\t�IP����6��)�UW�;8㡏-&�~� ��k������]�FW~�Qkq�<Ƿa��K�:�qp�Qda��v:_�k��Ck�n��?A�X)����W�]��1WRz카��T�~k�5Ə�:CĆ�$K�S���)L�h���%g�sg"�Sr;~E�3d�a��t`tbZ�������ՠѠz�y��o��Y�1	��ŕF��O�L]�ɪ��0�lS����/'4u �-�ɝ��ri���3����l��ؽ��9�Cđ,��ӽi-�	QA��";w��@o\i�z��`�AI	��H��������6�~ ��$#.�ң�]C�Ҿ�.��KS��e�f�A�������o
�򷬲�GSu�)DLy���T[�DV�-}0p?��g�y`Y����s���Q�r'@�]n[�9AKl�{�hwn4�Ɵ�
;<"�%ʕ�S�Ko�a�ۓ�8x7�NA����X���ι��Nު����tW�_��y��;!N��p@��|���y-���+����s@��aɓ_M�*����X��9¬��r�;Q�v�qM���~YW�r�%h� m���9���j�Ө�-���C�W)�מ�y�d�]����&�z��-��������!l�w8A/�a���e�g�^�� �8+�*LQM����[�p�S~�.)�]R�	��XlxVHYEB     400     1a0��p�$A�o?�!(;��8/� =���ypP	��l����R!E�j(ۈ��S�u�+L/��,/��4�OT�����M!4(d��n��Q�g�n?.5����>j��֐<a^Ćf��5ԟ<�G>�k�y���;��L����Վ�Tu�`0ؚ��0���*�[����r	f���>�R!I��9���j���yl[l"9���V��3�����A7l㗅ȶg�َ�^��3���^�5H���!,"k��z��2t6���r�K�{��"g-�gS�1"�zQŠq,�,��fų����Uh��N��Sb�R��`�}� �YhG�5q�G����@.M`>5֣��������W�,�,m��#.��?���v����+�C{�I���@lMh���$`t��^��tߌXlxVHYEB     400     1b0��h��;7������ƚA��B���t�{���Z1��M�(�b�ޒ���*A�3^�ޞ�+�� )�b�VMP��9�W�Y�*���
B�ߴ0�#���~��B�%gmZ�rD *��v蚐�)�p〤�Y)?u��=���R��z�^�s�z����o�O4Lr�%eK��ZW��_���_��v`��� ����7��ʺ_�}��Hbl�Ӳ�`
������qT:Vo\�4B[Yq�?�<�NyD�p�&�c� s���r�ƴ������Dy��E�g�Az^���C`ﵮv��6��{�	�ߌ�d�Awҟ-`t��R �ac�C��*�����no����;�_i���+>N��|���o��t4��d_hA�~�ڌ���MŦ��XRQ��az�m:y�9\V^߷����������8y�T�P��]�XlxVHYEB     3f5     130@0fw�#�,)`��"��~�I?�@<@S�����2fDs�I�t������0�Omi�X���d�=���l�5��H}��m�3̱X>�l�?�����^{�*�.�|��ɵH>�;P����݋DD!�+l�͘�d���rΆ�!�	��%����� �MG��J�E��|��'r��}8�!
v���J�-	GA�^섉�0C]�uB�)���)�!���~��H�1o9xGQ��?�I�i,��캽l�*S�=�aVh^>B�tʥ�_,eI6[�VC�dz�ms�H����D��A