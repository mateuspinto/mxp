`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CMxAniToRZ0xHdRD7W+oyXNWHmWqAAD754NAv3s5bqh+0BbVre346pbV9lOzcFCszi7oLql4Qq7r
ojOMgXUlg73rv3MX1hsFjdWqW2N5pfbtG6OQpHkp67bTTvUxXA1pHXFbZ7/TSFTYzA+R0PApfUmZ
qcsGF5+1ngzngVISkLhiN9xef5SWNK7/rVvT/WAj01mX2taLLGzZBlRN7juzsJoIEMtpq7Q3+3e6
ck5zfa9Z2IOngzJu0SraMudc2PnY38+3OKz7zcsvJhmI7yifqqN+LVRMmQqZt1PsU89m4tobqckt
1VRBeS8PV4CYUNWL+zO8rQmtPGCCj6eT4okG4Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="rbi8ToHIol7FpSUNEcGIFuJewVmqK7QFKU5YnBOXJ2s="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49248)
`protect data_block
CyTw1YZr1zf0vHoFKd3+6aKMS/wtBivz8BCQriqMYfbETfa0tSZSAgRlh/ck9FxWCZN/YDtho2V1
lVNJrvyJrpRDUMGLN+9puQX1A/Njra8Ql2UNqp+cFRuICBIArqFnoLV2xOrKLuOMHEzHNlobFYcj
992MFgCBXLQthHJjvSx7bhXHd5X/gG2a8U8tVkSG+jvcc/EwLoT2r6/Gh1CV3LKQXwAsuJl7SsiY
NYr9LGOzIgodu2CeRcY9hdK2XbOoMtXRM2NHcdit6evtq0NDJCNZjzIj/ALfTS3wkb/5JjliYu/9
G4fEDx/HIHghJtmi/xNASdlm2bjFBoHGRUBf5XB7cgz4lS+77KZxfizWC94f531+TPJaDYIhlIv5
dm+DZSS6lwoC+XENu2jrM2snnB1nZOUSXfJAaUsiLxlNh7PhkxB8JCdJmpwCtd8X5pbKMggKNh5T
JNZOWG/OKS+OjMMGYnTurolTpNKYHkUA7D7xWNpzGyu5Bb1nZM4aJg7j1AiEETRWbdIEhWeyCvYz
RpuipVWXraGbq7lRvPV04jvnrp4kXVLqC0bbR9drshvF2FTeShUFi6ddE82g9rmC7NoEuGCVABe1
byZCacCwvzE/0uXQN7DAnhLseMY1o5VJvZUwhhNTINX0AqRXLWqGyyRHbo/mz2EP7KNREqO5aymz
vbOnbcEEy/3a4sAHwb3iPUqEo5PyOFKYz6faVe3ur+fgG0S9nTLW0ax7LPLZmeZBdm/f8Nj4MKfj
SaCBT78vS/bHDSFxE75x6r1fRtply5r6NZy6atW9JesMFbheZhtrE3pz78yzN4El07dvHTYpd/A7
rIZK/thPrZtfgl3yLSeVl1D/pROCHMSfxTMERJK0mapU3VUBJd8v+ByJyJuMiAOYFjebWzE7cbto
topZCrjZrFylyCLdYipCCnYagfVNvUx4leiW6OnBvo2tMVr1oudvvGXmyNnk0WLT+1W4bG0BZ5WF
aJheiPmhe3Jf8bYJjbK8c/+FlFbJbyiO95E2tQtXpF3HkfZxgsTFXvGlm7s+GDwcBEISY1mwnsft
M5qwN1aJRLi0bTtysn+VJ1GCw7DIBC0jGwHvGHrW3AviEMFLV0hocYVya2C4b5n+kC5QATyb19sM
fBDI6X1MQLDz+h8d2J4dn0iFKQ9QjpfYbROk7jn/jgewZQCRW3XSKPs2gMBqfor6w2Ug37VN8G7H
6JCABiK6bmWPftSjnY8Vlm50vu4J2KMntuSs5qaBa+9lxT1pF0vS4iCJQHVEvM+ERP2i9222zMg/
d3/IOQK2UmmOzEApCd1YVFLsg8gaKGI9jFArXUsR412M7rQhtGPz9uU0E5B/YCCH+B5TZpUQ67RU
oxm34LWZ+XJNMws8P4dh34aOmKVkMTfBMC4m7LfIz6LPjIlL8A3LkaNo/EhtbQBdH0kCswL2OPFC
WMZl3Ax05y9hrz3048xppVTdK0rpMbSNj63Bjznpepsw+GB2nh0XuBobKlDpHp/U/rgcNk66rF+H
ILA/mAVEEjIbBP7Sa3XfHtIGuxayKKVcht+cmmJo8qkNen0FjDl+9iRtR0SQCDO1ae/EmLcjWD0a
Yhh0maIuHjDoY7E6PFX13tHdX/7ThRQ8kt5zt6VSXCd4JHEHEaEOthWfi7xnjbc/fYKSirAFfp7U
2+eTWrndNrrgYQZoWgHmANj6IP4YxnRb9GTRICXHNDXUo6jerunbNlzuu6AKNkixKye372IN4VOP
T7GSik6DJZWB4N4I/X7qGwDrGAbzoa3t9Ta3+W291P5McpFPHvJ+PhBA5G8FF9eX9g1kisyJxgQd
eztnPyqr/Ild01d7ejB0w+zAW7bp1DTlJQ9d1meUBFqCU9r0vdDBVP6j0yzBJm2owOtHm72V2u03
d89nSzU/u+UQng2QhPnfQuMXU+bqOI/5xm9fAN4XDE6N2lGCnM1jdAjpP2IbqNZ/bKtxwpTXCcRS
iWh6nkqhvGfvyunYnh+LEvBaVXenoPJr/Z3dnWjLwuMnCQCaCt27ritjmUdUOTsQ28dkZMrgiHqL
A4+CbZuuD3HFWw9SWB7UKsMoIPJ8jxGWWWO4Zmu81sNTVgGJHDusOWv6ISPm8jA49kMrs3m02sgV
JSpnfmilniQyTtUmQEDWtPa006L7X7JCDFelytk62uTc+0KQFS/RvantID722/KCRbIBqRIRKtvy
c8jl6ciAPwe9OLfPiwhLVQDMdb8ZlJemlwdXTwH8ISSqVmRP6Sb+Jf0Hu5vZ2se2ZCrgntDh1/78
406Zhw58QClRiy0D5slIn0K38KM6LG3EPJxVIAS8hEuO1LgxbOgFfw3tyKksR1MBsHvdpzOYHNra
qiWN+obE6Hr/pe1Z1z+fa48JSuSNqXa5n8IREwYWitew8VjNr0H3FnDMJ1gctOI2ND2bneGTcCqV
h69hbdIc46HWOaYHM7nEzQ+6n9nQ+ISw9Nzw8r5Ks4tk1PUqkehWnfosvg23jGG3vA/77sCiUjrY
AqyCN+2xLu2E1DSxek3dMQoogp3ScI0hiKlT7xnclVbIX7rrZOXAEoedXuJFxkoy/RZx26Q6ZqRu
zqtc9g+La109LpBePhNp6/9tKofEh6ig4nlUj+D4YxYz5OU20fmV6Nr+hi0s8CiwcbFflc9eGylW
PUU9uvJYqWUIQWZLHaruH15o4Q2KJFBIYvSM03GJgjGAAjHlC8gCcj9wOA81XiM7hXV9+lHfez8J
TDBGr5LKOpFbR6UZ6EwswI17Q7NAq+gq/Co0JJWIgVZqwyjxiURrxpmxj5ISOYvOW2mTHvu1RW49
E2N4wRbQdCqVqeJf7z45tJw7JdyURxqlUNwhhNQH1mj4IiLGETmelWVLr0sWLKt2VR3Oo3LnI8ke
DyL5d8RKh7M3+bmR7IhI++noDhSTMmzIj2H01IGlqEI7ImfXNrP6gXTKYWASqN4c/0c6Xp8b+Yev
coejGpMqtnPiTQzMEXW/7eCadKya50MYUechdC2BniUZcxpUDXaRbKJocu/16MtRm98O5GaHau0O
p0uf7WGESAJXrQ1Io4UEt2qw0Yvb8zgRAdqkoqpGXkzhaCuBzbjGJzIhMVvE3IpVXF4TRVaIQzWA
mO/inrp/+oxVBSzijHjTjEVkbBiKc3E+KTj4efjrVsDFeDChncmCcivcmuwT9lVKdPoE/rJkqhm7
YbXpVI/RSxR4OaOex7zHaw6mk6G1HNmz8I9/e6sTEmsDgICoUUpWWbgu2PMUPLmaZ2RL8MgagUTc
2I0WF3/vLBlimOWccP3E/NtURnbw+TtK85ztPgY4YeOj0tjwltvIC9PjOaMYJvTmzFRss3zZIse7
hH/CN+3E3fyWNLg8/EN/MS4Q9/aVxbLSu3M+pSDMU7gCft7ZRo3nodbLL/UNJgH/TCDquW7QwWNb
NAp517JVxUQ1ifea646kUkENkNTjE2Uc/93h2s7CxK8ld3cGH741O3MpUdQqr0pXhIkgqPz0YxVj
ZAp8tcpMF4q1flbZWlXPdloSq3qcQED52MTY8rDkBqvFXk29PW6saKHrFf1PfezRRZarzhk/VMRt
pMK1YmMFGpt/fOd2RsGdfJVYoVgjrXTSvTrqSkvBX/Qy7MuA3Kzl69egXhkOzmM6jR+1jOce79SX
57GGwhvOdg5o4HnBP9CHe/nrcp/jS/td5gXNrw8qN+aE4e+ccsx6qNW1UxsqJa4p0EUZC4TJLI4K
Aca753CWy+kBrqNwfC+vbXsRKXD03hypVX3fe+uF1JeQdvQRIZQ9ckYPV3M+hBQD1QXoCNqvQev+
kBoI5LDnHgZaTMiHq/ts7hNdvG2yLgsO/q8B8/rnGQsQgc4wAw3JABc0DchAAjzIypX+BrTL8XPH
3ogQz6JS7twi9RcTPJjn5YeE2+SwDD+FgzglOrDpMs8j3XnXHaRem1+3/1BW3/MsrEvzjkmBBgSt
8KGOF5Lzv020LS7Z8A/AobalbUsPVAB8RwBh4YsxIRpHgtv2n3K8u6tZKYnBlxJMIDhzmRrImDyR
awHcuTe4Fze65mNklyvK2yj+C2LUpQRxRFK47T9YRDQGg+5agD4yoVxqoUP04TKbPQ/NLDNDpy+7
UretqAGfDgUbCl01i6+ZUA/EdtePxKAzarW46vzHWS8pCC50EK/bujRKdn/xioTnqtoJD99pxyrs
7TgE2Gkb7hCRprxIUtCvzxOYztud61GCUi8uwLOnmSPgey0urPxTnQ8JBmLVtmAjs0s0BXjcVrs/
x1Td5EWajpDRJNyZwN9tVcB8Nh8NBPYrZjdYIfdHWotS+Bko/8qk4aWtJJc8P8zBydE2aNDlNt5U
x3JUR3RE2A/v0iYOBw7Pk12tR/HPH7J3AGr/+GItGYQ8hrzp65fMqjCTlOb7cunw6wTxM0FNcWue
XUUi//jmr7+a77+/P9NihPf2rkjpqcKiqL5HhDaDqRBpJFT3ix04iXHnp6xZMWUtInlNl1AsSBPu
a1oaZ+5Gg/COb9WzxUUMvvody/Dhv5mGANjmW08GjaarvTd0aPXJj9J9o5aZsTDh1cO6+z0w7Php
P5FlomKkcxwd9wjKVvt5DLqkkOPf0uUeU00p5A3blD205rN6b1pG61YGmEPx/vSB3Nav/letbZxR
/8hbuydlo8NV68QE/VS0563R5svQVvYackNn0+0qHFzdB8Gp7QNSRRzqHimH4uJg76et1HFUZLuW
Ks6M2ZTMdZ+pVNrobQJJ+6Q1X1N/YnxFbZIuCDWvgxwkAa9JRTg6Gjtp53zW62KnVGa0So0ltBX4
h/AbyDehe0AaLg/daSkdrk7V0i87epw2tqw4xTAXkmik31XAlEaI6modYfqED/UOlmJc3vxsppYg
nTJqa2Kyx3L/CPjMYWqqZv5cVrwyQOsLSVj1nONJfIqrMfU9Y+ik4mm1lLNv/Mk5Y2ndVMhaUGOy
bEKX8/WtrfJB0UM0fOycKz95nTkVLs1AfLtIldRXbtis+S3hUy7eaboeCG/WMzVaQ68FbKi4c5J/
+MW6mJaPctqoh9ecu7+iX/yysA8QURDstpC407UlUHiGmzLdOPAf1hifD2O0LP02VVIEc1z2w98J
401BDcN6mKB/McALrz/wJ1NPVWF60AB4LnkOclhR+1MAGk78DCXCaGJyanDvAsnufFMl4Gz2AYcG
PQbWcz0lHcncob8vKluIP9RkGtheS1O145Wt/sEccUTm2pSY584+E4wR/QXyhy8jiDfm4QCgIj5G
HHohWvD9aI5qnscBnZw/0tc1fOFliZy0iUa+j0VlLsdQh5UOJthfV4fkWbLLr/HvN0ZiyeA5nGBe
GnldkMoyxLvH94OtbHT5ExElCT5xSeRtjpSOPTbiZ9Te/PNMvJZerGtsEw4TN6TabbupQx1AjdKm
SHHDzDnYEuV5XH2IJsJ+Gq3Qw4vkHo0ZxH7oo9YlioCLFCoKCWbyYtV+YUrAIulVipOUWipvMMgZ
kOQNvy6tzoBqzbDALPIXkaY/CJlyM9AfYqrABgXEdFa3fsI0r/i6s3qDvH/yjIm9d/GavSR3T1NF
708rBykY6gXRsBBKeSiTWCmkmysxOmuZr4FyCpVNAXNSt39ARXS+xAhl6RtRwnKLyUharUi/fOVy
KjJRWlX5mfy77dIH8jpZPAHZHuB9bI2Uqm/EKoF/SYuexfrZWkvvYztONOYyXDX5jgkV1gAXoEiH
hT2JiwiZ/bgSnqN5Xm0SlPSN8e1M0tPFPAGwZcvLYQKgay685cmM0yp/UPcE9cVuxL28ieGfUq8s
WS1CEgfE+m2Na/1UvnkTnOYpaaOsl5Bivv59IZJXim46JgxHfXATHgPUQL4i4ND8GWPsBtL5XyOe
BNWsvC5/V1FI3VUAu/yhxSi649t9RBoeO+slVMohwjnqEZYXUA2c8IFobpKht+mT83mtB5jF6755
n2EREXuJs6uBkUtM27MSZO9c2u4dmQo3sMc76yXEO5EnLcuJLYXBN2hqvP2ZWPTgR+/AII2xNCH+
KFJcbXkolgjsXQx9XHGrBSuaGMGa17djdPAe9LnIqTMkFUc8QxYED0d3U7m90rcep+EwjeDFZYJz
3IuVxtYUth9cos6FECDOg2YmRw2wLWoF0FEoZcNEDelixs2FZKA2TlyLsxw4lFAtKmwXWpJec18f
g1vtr1y8LNpdfI4JBnRgB4Mrfh3ydUlGQJ7rT3SZvbcxFRWuLBISZlXl/lD9r2kf9G4fXDEsTUFA
gw2/MWoDg1QcWliQCHnyMrHPEo+bXbiviuVEjpF75nFMQQ4I9aZ+1L/k/cHI46Lx//xsdmveVaXg
8ANjI12UgVA5q8XcZOAnnd7lb4TdDv2kc7PunfjWV1Gr13ODv9ww8WQ7dA3vF9J87EkYAota7s/z
ZYNeNLc/wGU6+7nLx4dz9hjQC0Oekf4rpcmmzUIUaQWcHtu+DgQP+XDP0jiqbrE1Nl5XMLiaA1NZ
JkS1T/D9SZEerrsh7vnpEeTRc4vkl3s5jTJJWoSAogDJCEJEvMedMyYcXYB9REgX6Rb0thVo955K
0WqcRN3oojntG+NK6gHtqToUk//9JT4ErQsPXh1G0+O9qTmyXKc8bmbFT4adOIpCRIdqwMqRxCNM
+cG2Z/uWHo0NKjC2NFxWCaMCrR2eQinlH7vd7NDsZ67Gb0h2cUoGaelUD6xVPYuiAAhysBbDwdQF
RqLC5j9nnpVsBZREm6bHPguTUUgPc8Ux2gqz9Tu6uNC74bAzmp45XpSrWwCZI0Cvu8CG/lNvwYi8
cHrypOR81Gn1HYIYi9Rup321GtH7w03S2eygRfrL1HKlJpmwULQWf78eu8Ky5oB0Gl5q6ykhWIID
VxKY5rhTi5QmJSI3h5DujFlSbokXELxilH/8A+y29XVpbG7Vgfnt19RNm6tfDKXHK6OtZTuQ8dEk
WXjcBmo2RRjbMibaoXcmLYZIsEKZN6vaTX2ZhKEjXTu3Ns/R1BEYQd8e8M4P8x/oWie+MQFeuR41
hUBedsXSbbu3crV2bwip4EBUbwBqmgM7A4qRumv9LuopOI9gaL5DmAoDa69HYgKcNO+SFHOLNiYK
2BV291aMW8F/xvPd05e8EzgcNuzERCNzxpjD/6dSiE3J567hzVQ5hOC2XY/NpEut7UZsuEeRGWcA
Vv9zT3Oq/wY650QVK0tUT1C0iFQ2if6M/+vqa4OrwX+zap8DNlcrgQE79gK2+dMDDMG9Jlj7VIvk
vydA1K0XXuig5M76SOY9KlAfGUUwbmGBb48H/JFW1HReU0Epr/dKsM4yZamRREYuxIPCPzDEqQ6C
eO/d1gyU2s4JhtNnXnuCBNfA6Y+cpSG2x3EjXXB+yedWaLTnPNxLhC6B3aamm1yWKpy/vZeWUPuB
mvZyEe0xOND4u3ruG+MK+1136/nDrU+ioyrPQ6MjzDmDEhjxbBYO19wkgyFM/BAwtA27rpapaLtS
HmMxIB2OixaAKog8NtM4QmxHFw01DFr1FPRMuSAnTi15XnqsgJ1WT1dgzDfIkmsFw+6XxQPH2XEK
JZZW1VVs1CE93QbEO365Y0WLBhE+cDhdp+2/UboKIZeaQ5cfjughRVFrzk7enjMLZjlsSm4pxldH
PhutPfQ4nxY3E/+Gey7JopBs09qBJueIXKF2okNRDsZIYDSZQ3m9OQcYWwcFurqTmFcQLg8mlQwJ
fJWqwgceMHgPTdLoBm0r/PJydvxEpM+IAPI9U4o3ar3wsiLy0onDn4IaGNQg21yXCNdOBF9c+Tnu
kHDBm4hb61IOOdCCHxUFPQF4UafKwiPah3koAGN6qshGFTkdT70FOfKLW3G8LxwkdqFbZQUZ0Ywv
FRvTipWlnhdfwUnN9PcUExEwAQ3Y88NH0u9g7cDVwmireLSGQ95cfEzIef1DDr+plYd7cYSnAVY1
lCDLToH8ud62dKtjGBjMU6Uce4q1S2dJWhUkOhHsJvh194jUKHcFmffbfCABoHe1hpPAgvE6v9IF
Wwqpid/ZfVVmfqhYyqPPzMIIwkkhqqxXXqtDfYyE31MuNCEfOjIW8CPcFzRco4jOrrbSY7Y1RHih
4hDIkxEu8FkJ25GwF3GMKt6ThBWfV3WVrnjLGvRlp2NGjaFqOuubFBLvi5etZOpddQPSFYX7167z
W3cbgXs+q7YTKzYK9T19pF9DXL/y5CEclivE/l2TqGjNddQcW44LynDx2dprhloSr49r7FXJoeUH
v8tbidV8j8lm070IPO1JG3+J61PzbwjbSxvnbA31BV8i8rvlR4coEl1Eh5zGCiWyJ/Dl1Iyu9K51
qiJxuPe1hwK9Z6i7FBGQgCN/9KiNNJGQ5JWK7WQ7I++BIdcvAecbE2pi9vNtWnQ5aq+n4OFX4slh
6pTvH6C+2nHWghsLHRNh4RDFcrA3/SdCQzrDFVNpn6xX+SMF6n68bXGeB4l5o3XiYD/0lF5TSN7L
E3Lg6dlynv7uGlnclua8lOi0octS9NHS8arUK9wO1FOhQePfLexKZqJ7qPMiRK45jIH7WilxNW1q
VN4iYxodePaZF76Sti0qf8a3gugZYfszdrgpvSyr7s+ZT01J+6VHD9lnjO9mimfhc6u1Lf6ibeTI
MimOqD6FJYJXMsExA/av66ay4M4GWU5nV8TflDjln+EK96zQxGWRHnq8a3fQ1D7u0o9YwkaP7pXm
/pFYO8EDbe3CysJXlNN5eKq/BRgeEBaQ754eiiop3xrp5KDEIRCfwDllZ0BUT/W9cYZyBlPhekg/
uUjdQMoQuO4bnx61QKObvvwIel+D0RlTBZmrqdmKgdcaQNpPwShwggbT5gfZZ1EAqAZqFFNuPmuS
fYpiCErlW0+1wAm/Yy1OGi5R/apkDWXY/FRYOI0BqsUPWv9grnqXWZp3+UtOEhNzvebyQ9bFEmmO
6Lq8imYzT5bwBsDrCTgyi046CuDaDo/YCNabwHVNB18iPbdo98/os4SRNhv0fe87B1hOdqjaRHva
oJGKvGhzhJ+wYEuOnHOEbmwfbOTT/f+Lpwdf/rXfqoySYLy+YCFYVbXT2ZjaWpiRw/UTpPs537Gl
rMO3WcBuooCBLLDbUlh1/tOdZKsEepHwyWSs2A/Pp/zzIy0Ssk6/razseWxorZQJN5CywO68P31d
f5neS7wiHDuYVXQgxf/J1twt5gK0AQGEDPp487/q7tiUT5GJLL6RnpJO4Zlv75Ac5/8oEAloFGEc
zhsWTSpq3UMnLh7v8T1Nicz8uzt4AX9gPmGPL0aKs1PEfCDPVAUKmZ7LAaMEWTeUHxMSrRokW/D0
GEcOXWYhVpTd04g9lGVeCcYzL3oSt4oQEECK/4qOPUAP4LDT/9q7jaW7/tq2Pgd7A9AFs4FQCsX9
wiafZ5boyoaPBZqnLRgmL6dt6ofWwDAsizZhHaAGJ4fVHSGIbMcqLGCJekQG6zUPaaYWAotckHsB
DCSFGSb3xuazbG7N3Mx53I+4HwOfwvBVusLYYOqDr0678gBozUncTsGus2QflzrcwSM6hUjdgvxB
rNNXSjSyyxrxdI3mWT4jle3DKD7GQciKC93yj42yAqAnU0K85M30bpcEIHRJybDcMFp0DOJKXtrJ
mJOPVEdxYsHw8m2OeBQcwDO0A3t+qG/OrU4E9HeRZdjLGzVjoMX3aVlDFFIq4qcIVFd6CXnPy2Oj
VvQQwJICZWKUmnHdQ0AdeXbE9GnkyrxVzmtWUUePzhi2CUiUSczFnOByPZ/RCgr/TXJgxnSSzs1K
PadpXbWdeoyRktqERoFhB6Z1MSTMZGc6iOHBwlQhnqNOskBM2BlEHZf43OWrT6WxXnM1E3gCQaY1
yVpIRJoyU3Vad6SDWKRHKLE4YbFP1tpQekXxGTMoZSgYzijbiaoFXBhtZo+Z3rizjztgy4/kPGl9
UNzwziFYFBDGsVWx9j9xyQujGMCdfTvFGwJE6T44uzY/gSKQ2FH8balTeo5iEku+j4sqF8ExROiO
3jKROku+Z9EArSQ1et1Da3+LsaLp6Uuka/gg6glAEYa0HNjs8Foq8hZOwZexVn47wpoeTJgxCYbn
SnOVoaxDE16r9PAVsiHd+bjeM/PrZTuSudqlekbcgUwvccGQkyBFUaYYomLRuW/k5JfecsYJssmb
0pcmNKndvmOc24BnSvyxPNO1ZPFbFyRbur3zrDKl6FhVq11TuBGNnI6oqfQlBra1M8MDiL/P0zxz
tBDg7nkXcxkAnEOPLedOm5FIKbs7ZjNgWlC0tvIxKSO3r7HEtCOEUoqr+hr8U/hAKKWoEZ08eMQS
rFSgisiQu/tMszSDwcWI1go/dhoDLRoMAQzjyxM4/WgE29OCcUZqw2gZ9tu77ahWr4X6izFluKjs
iexoQjsyK1nJSgqZyPx4Sm7Vt3AX666Juwegk892b5vGj4OJ9l+KGLOaPSdsz+4YVwpPjh60DzeC
9FMbtnwGMx38Iw/+KvSxqjk+TUUOKNWfS85ix0qfxXabFSRop9eGonQAR/3yzZP2/hd/sVFgcoAc
DZvBcwI5AuvkpttRO9znWaEJm2g6vCk2ldoZxTuhY3hgNLqIH4H0KP9rXkyoiT5fC2jUrgobm7fp
lC/J6JXFYMn9qfKvCVtmcXYtxiDgoup0zw94Rmw6T7xPVArL4U9oOUlVCfXJ5lCyHWbEWITMpM4Z
eh6RWY1ajXhIESd9U3kJdwNYHb8bK8rizYlf6QGLKv5oUzV62mFLtad8vd2TYtGrpFJimpzg66y9
JACXRCPXfoxObIHfRdPJYrazhHqTIa/IINHaijohF+O8lr1N623RAAW3HzXP3dCP1Svyo4aaqhri
RSpXNeBk1vM9uJqtp1Ji7DH+Iu4xz/1X/Nw1yY+V0lkyZh06F331vzAiLlkpJ4qB0M/QXb5t0qd9
z4/HU1oweOb42bYnC02PX1xjVzn4wMU51tIHYEf5QgzgLPzjQIzhNNR1hzqRPCnVqyK46yb6opU5
JQHWlvrCnFiace/pNjuqkCeHnRRHGzZCKCSHJWPlFMjEiPy1dIwcpTnAX84CIqvn+wdF3HFSuFTW
uadlx6w1eJn/VLlq38iNqpawpGcFsqDG1ZGYOmVERklAFPmHUHiwIp+xWBFVa+CcAgik+WP7brzD
Nd3cmn1NSKeQNova4f7gMtIVzpjafId33tCIka+tIgSLgcGDFHIbSz6yI6/V63A06RwsuCdseeUB
HHLgZBMnhJ3+v9s8MQjUmVtOU8UYyms8yqpInLniwMY7I5khjuGY42uMBHK+/ByDGYyxslnUTymw
w8xgrq9xXSYOS5SI46OllxYkQHnR4UeL840yQdhtbdMtCeTgPMHHsNbOBppqjTzCRhpmXjNh++hI
a4vT/8WkqGbQWbUY7eZfs5xr6dho3U4gWk2iHWLAS+GQytbSJkXa4hg5oZgix5Ib5QHowcB06DlI
3YXskft0q1Q1pfrJYGzAJjpf8xsNWj0UWlBZFnJCMveQWX0slOJ7/wz12ODWkDBelpRSNH/1tLj3
NguPWFsds+xyzj8i1FrGJ2ET0yXxrssXPpEh3jskydqOnrpjIepE7HSml6Z2Epw0P0YZXbRmzL4z
9IyPbOaJxwCTLbI2vKiO43LC05Re+N8G6exrmsUy0ub292/2v9bsuec0adn9DN+bvBx3LEu9myxc
nOd59ZxPGSCN6fS377ZvQwJtyIfVSYVOIJxGlqN1Ak9tqpOnE0DYYxu+9oIMctIdxCqC1p6/1Rg+
cbLzOwAMows/bIAGQtP2GUrWILyhJre4/VJgIkn1g0fGwyVFZTzc4m9IHre2mo4Zg0GUE0sQceBa
S/6FsuarDW1y7OFFkiTUBQw713+j+pa8d21mO+YccH1wP8fNg6B4AYRSHsDTiekXjpxN37oOFyQY
d3iquk8CXpM/hEjexiq7ANtYSsaNGqvtyLxoy4kQ2VgP9RSot/gslRkosT0/yjiiAmben7uXhMNd
bOFMLrOi+RjrF1yhlzW/ix1LPGwifPjis+P5YB23FpHWkbCkfJ2ySH0lvqr6+6IAO1IIaxc5zbCI
IINqvJArbObdgSDevgbJvkZu9VsdGJdByfRSGUnjxXKhW1xuuYBKiknsZ7PVIj9Gl+mSazIE98fl
yMu5PRUOWQ7Fx01NOeDg7mxeAmdeDrHaTiZy8BRajRceV/bD28w/SG4eOT8I9wKZN7XaEsso8rGW
rmw85FhKuEe/8bYnhNMDOBEIGuDSBUCTWcvUbJHYZqy0oKBtCdWLCfYPSRyGS+00FGrQCTLrPHph
p/UxS5P7bSOSHj56+3ayCdd9g+ubpcfEz3z3gbzohh8KAlpqGbqZ9SPeNdOZSNwGKPeBB2phhe1C
X9oKzTA9knXyBwWO5eu3ybuY0N4ZN9igMCQy0ibaRk7vjGp4Wcz1cbYcuHP9LWggO23w4RFNvhW3
E+fyMjC9iKkzaCvj9aRIGvSROUULCxz/gqngOuphwpXJz1u2Q7ku2ixgszaEgIrLdveqbR+S7DMn
e/wTM/RoXHr2lsEuKmDaYCbhHsk9NSJJJiQ4uLqcPBBT86f0NvWXRuMqirGgz9i/9vsjth8yE2wj
SVtvIVf0Qd0IW+RftUuTRCfA+2tMX+a+/2EOjidk5l4YojCb1RhEgBGrjDPC1IDzJfx2Ug1b4cvY
EjIEiMrkUsrEwxVLjuv5dGObLc6+BCeYJnyoIbuGyjLmoZwKYsrZgqApDpsum/9/dnDFWXh9eCJW
EcasjlwgrXWijYFYgnB6stP71Sw86eiSf0fDaGTODiarkvIT3ijrAO9VquIwTLGm6fNwsanrXe0w
rqizRTZluleA7GCHiaeu8YmzdwKA+Jo+7dF3pXVREtgWCssJe9QZK3HeMF0x7PSxdCDq6x558Vnu
ThKPY9cF2Ag/V9KJjlM43pJ2FXV25VotPpqt0VGYSOGmRXl1l7TR8XiJ7cqedRSrv68rb9DAREXr
XKxkZhHaggTr52ePfGaEw9tzlZiX54sNZ/BQP3Bu6YA1tp96ltoFZCKqCyRYTiHdxgLH/69foYhq
4KjxWEozm0WqnVoRw0P+AvUA8DU22IgIk8lCzUyyh4h86UE4b143RBrVd1MFRHQy997jF6768Dr2
+EOV8dOE6W8cD0ja9vIPZqHYwv9nm7a3Wjv6GloQw4wDMEGt/oP0KEs+yI/3zU71i3dTvrehjmmg
e+DHgRkqGEhe7db7bIqPXoQzhBW2/1y5B8Q++XpJTCPjRmsSUzT0G5u2IAfKIuk0znjauUknT7+J
vze8sgd8pDq8pP7vwPwnZokbJWGHSjaIR//7dlUxL0vUJSIw5d1qrbpaOS2YBZ0Xm1FP52ky3+Fi
IRvMDMe6n/W8Bi+tmhP0ahfmgWSlwcV3RlsBAw6w0MOkSaMP6JmNaEdnmj1u5kZionQ2Lk81kuzh
9i1cz4m4lIeO8nLkLLpmrX/qQPc5zDCfxSnKcoTT+NjxDUbhUOGlZy1nG9yZtrdCC0oaYCYko0Rq
uI1E+/L14JNPS3GdLg2ItFt1sbya6A3VWLku9idMgmTAedHzPxQXj8jSEaYfSMVAg6yjjqYrvq68
2jWe3FFuRCAtzf8tdHeFA6deW9gBNB6UM6q/9a7kXk07hk1yTNoJ7XNzZITeF1zQjJgBvnBeLnli
mZ6D8/WiNeeXToxYZ+hVjSBvthkyvVmh/iU6nil19NYpygYVGCkkxteGF4FA+YoJHDXe7pqoCqQ1
p7poVA0gXOA+vZVDnQhEDjVWpuRV1ALW046sjmbwmNo388f/zw38GtzdGwR4oK9klrR5/tgKzGqH
52YRwmjegvuIR747eozWlFc3iARrsq8WAuD/x6eugpUC/yawlRPbYJU6aVByEKUK9egDi96LGb3l
BfEPFtzafEqnLtWQTrIZx3gjz9pIfJe2eW4zEXo9H6M1QL7kXlJVgQ+rLVXMF7vkqor+pS7YqfFq
Yf5MvvHR3jJLgqEUaKRah6dBwAETLKAunwk/LJeAEq0y3d4SuiecEk0wsp5ac5r4Cpein97GzLRh
tu9FyqfFTeGsQyh1HuJflTi1UKSxrOA/1BgVv/TzoDNfLsZdk5mc3QNZV956TuP3XlwX0pQTXrJX
fFBL75Sr+71dsDTjp4ieifASRD2cI8JbPbibSpyhy5mHaMfDKpd+y4u67DPLRbY04/oMEq623t4N
gzOZniPq7cYXhqRP5fQgdadMEZ1hx1w48ek1Hksva+SjpZ10XyR8RQ8ErDEYbrjoZ1J8e6fF6ipp
OfhJE4g/kGueW9Oh38PAUHXBw3Pdcy6QD5apKfGXLYwuMPYjUsamZryOTH96hoQgJpBkVlVamOn1
gGNXCJECiPT+DuX6173e6hNe5tJLBvkslv7Z8xvVP0h8uQ98mcRXZyYPe2FYKq5tOXvfKIftUar3
fJpvGs6oDIVpLOHYMi7tl/lsjez5D0e1e2EFeUjhX4wuN0eq0Kcgn5NHSDqhPkjkFZoJH1bwr4tt
tEtZN0HC+7nu6dt0d3AZ4rsYrlFXvMZtOlVgM0b1polbujcaobXE77Yc2IyVZ3CWOpw1xk5zo0pZ
5iG0axx1+ytSUEmxUCtQ7rmuiQHO2Rjvx4bbr/Q/X5DMFdPrP/Jkocs6/lw88HIs/G6VMXKa/Bi1
BpU5Fl1IjYSJ83icFclVTmhxjxF3IXqwBnx4rfCLiy8YZZ3hUnzmEM8JNtJLNB464wpOvF+uwH5m
5tPWZteWl6HFNrx/lyfUDPGR1QYiZWSyaYlrWREGD06qo40+eiU4DaolAEZxypRKzKtWuptKwHYz
BVVBE89CckKRRJxslnBseKTO9jxmAiSkrlHWeapdbt0o6BHuRrWTO9X8KWHgpXcbdS6vF0NRP/Ws
5fUJzPyZDImkNbZsVM6o1k1DWOT5H1LMm0KbS3Y6PvVyBsCYT4FO6GQg8riJ8HzDmT1nu7i21O8i
0Fz1U6MYfmF5D72SpiccF1XX6GMkt6wZf2PTgZ6qK1xZBZqQnNEkSgNVY4G9rwzCIbA8vLL7AUUo
VVh2DDGVxqloQnUZG1PkwbXJapgP9RhO2YQBpf3QvJW+HjuhvslM2fnOsQgCOdA2qIezVoRYu9nR
hXY7D0SvViArW1hkEsdsjLupfq2Z+h7g5wxh4QshGz5c4uCHumdNccyjzgN3r9esgQFCUHVeQfr7
qqEMmQOwv+KVWvt3e4Mf6AkzHGzb3aQ4jfp9/lG1MsPo8CN+3/E58yEN70CIYV834WoOZ3wYyh3+
7S8NM2OZtm1QWXBq9f/EWgDeSHDiQwgGWO7ej0Ky01uiFwJO8k6M2n8wyTKVQ3vYQxULdNtaXHAw
Jvm8tHlz/jbh+561AKvKSB0HCXJNR2h29sjGRaohYIxHbIrXGFY4YRaWZ5zBdjjb70e7ZaSvzeIe
XSzzpohE9c6kc3dtR8Lf35UQqO8Ijk2jhGsuOmFvFSax0+QYWMxtNhEqIkMMCRU9ZOxPkGqOV85o
OSKjCmY2UyZ55jzlZ0lseVd+oC7x15c2czNf0e8EnoFVWq25ecPsJBKoZpqxAp7/AxWCMdvmH6TR
WLadxyifJD0+nDXOZe4sy1cRC9l/QU2rgOdX9NzPzgF69XAPGxmX14YSGyjI4nYIpmRJKqiKCQU/
2a7f8E7ta/zFrEjpAsBabvmvW6yE8Y1VEFBH3NMEYVUPTp5ZGCr+fULLoEaMH5rYP235VmU7sTIN
IUgX7zZzB4gi2qOMdJ9UZcDF8ZNTraau1qzFGawDfkrM2QZZcbAo/99A01Q8gWx5TBFKVK9jFl2b
bvKrLtSbCTnkR5RyhaqLGc16YB92b8/LARR0oaNb1fogCQbHdT2SGZAlnzWo2MNTYyZCpGd+yvY6
eoAn9teXIglg4qPHCiod1cL63jh6KryTeRxH7VX673UC2JtIWYdIx7JRDKk6Iw8yhkEAzE0QyUnC
5LtcNYm+bViw8xAbvqUkfJLW3TbJ4PB7wveFBV3og2KStUW4XWZZC1QKdxJfvnnO8iP1ab22W4fY
6AZk/AzVG1Xm6HL3SPFN3AnQ9p7w/5wvVc+/6zKi7v3wW7OXTxNBcEseYEQs465S2bHgimOdF4vI
uPF8ctbCatF51Bl8ROh3xOOlvXDZbTAi0uLdixh0z7k/qNpQMI+dN2Ni+1RGaZpedrLNFwwadv4E
+7ObMNfoyrAmZdvJ1/1ZTOED8kEabyO3d+mDEKvgv4T1htDvkiXA2RQl8E6yNJFPP4WvuKKbyrp+
uKtvJFlDYsJTBI8c/tQ0XpqXbYsvA0kafvM+1GFNOUuY3rlHw3mPQBQxtO3ILgXNVKoupJgWN1xB
Qve1cB/T2G+Ir/O/pa7JHb5ECtVcXhLImhW4oFrOAycqEXdmf9uqjr4lVoFKlz1P+72LUp7Ytm8I
Jc9urfRl6cLhm7hAsRgCjhoOq9NBsIbzb0f6xhy+GQODQt6R3tRXNrbaSIHarpxNoqYuXQH3t+aZ
lYucJHlCR8B/illplpaUxXuTmfdUh8ETr60+nJfM8WGuhhJmY4R4QXe+/Cyss31RkLzgxFYs+iUz
lVEc9HdE6GMdQoJjmNOoCS25B1/cZPD5qi1OGEpcghdR1GnPxJAnQ4G7YAwSlPaLcIwJzamL+aHK
B7VFpLDMJULQqOZNq0o9Bi9B6pMxzaEDICMQk68ewWwynWIMmxEfndpaBfvUMqcf60xQP8UH+Q5S
QEVftcLIg9SkA0l4BQe87FdNbPrsaKGwJnDFB6NxRGHGkMzHIUZ6nizZXVXHqITgcA9Z7YZM92aa
yWOLf56tm5qnEbmOdJevFe+8lOcwcDrSyc9EkkB6mVcdh3phMJ2zvsLKyJnDylmvzKN3hMzkheXu
ZgdPDHkx9p34cSoVjImBBsoJbEXfosLxuxe17UMRZE7OuRCPBjim9xjaXmeAh5y47Qvyi/X5Gsg3
B6KwjiriAARf6nTBAotrA9GbzKzz2pIjJk0vgXIHtpoYq1x/76htXB4FPEO1K5MQvqk4nEjREgxt
/d/as+imkA3/Gk91qHiJ7exo/usLTUvUv60RFKNddYKMJRyU9dO+t4Dg19mmbJb82vbB1bLyD2vp
Ghy2pudDxYNeALQJweTahhzNdylsPWqt0JQgOD9KGKhO0rkeEYE8ic0HZJkyGvbuIRYyiPvsCuoh
M2oq5EyIU59iGDIMJZopFJUy1vxRvY3UOvhqIrzInIQmhzPjdhOq1qGfBfuIuYun0xvjlty0m7T1
AbnDO9mqX1tOUBMXF3g/xx8KDRK6gI6T7BPqH4kbrPqUlSkfEeF9I9+xVuZEEOGEsbx0h3XZb07V
ALcVZZzVnkuPXSn8Vr9CF8f39nT9slv4YTLokIcFgT20+6qDLSqEx0OBnZqOmiUY1WuCUIjWMb8i
oFsjUTuRVZBvEPV1lA4i3w+Sm5m43yVSM+So/1apCuedTQKveoJaPXpx6Kr0TPlkn/aKzCHFYdmb
ZuMuFcFRPG/AjZFkICgmXvnM6vTDW1CdQBsnwI2zjF/faqsTcY3yW2pCHTN0b1D4l72CXyD3v4y/
fJsmtipu77lyxHxis3htGfajxJVsyVuohTFAAE4y1DnO9e2UmXZAcCdpA92tQA7SZbb3Y5Dil2tm
94WA4wVdi+5RNhooPM8d2mHpmVueS07e5pBe7Kx5KdZ91p6ss7g/ubRNP+gGikUmnKSmo4AX9wMT
aH56n4zB+sPR30rFwnPzGAZ//22B1dzDFwyUH+B5MuewS7Almj+VLh14ao28pDS1FwP7I77y+Fd4
MAyzcy0m3AaO4XBn+hSsFV40fJgVqA5aiKRe6en1fsoZCWpxmr/FMsnXFrwGSLTTv1r6SKLbwSsp
YsRqouJnK5ZnVV5otrij4Deto7F+BkzQj2RG7VW0ftc3jGN58gshT2QMXUOo1zZCQ1oW6R6ZcHjd
szkN8Yw2dhv0UxzdIjw8Bu2VTJR6gHyJN3Byvdj1XyfrHL4lLcUD0HSW4NrjcWj/JiB1qal3kcm3
jGVe1u3T6wp+otR9fpEaiPZYUxz7933GvHB10hOZLI1loHnY30oDRPGt+HwD3e+EiMrXEq2i5VB+
7gCNKAnE2qBTyqRhTXDJNu3O/uzLHxix+yx6+LUFLyrH0KjO0tpoODJ+pbk02GwRQCmsQZCrYPbA
6khI2rb5OUIkSR4mNFNGbhSxNmt33FEJ2xXwdb8o2LTwmtf2w1iMRsVXTxU4WZLfLa20gTT0m9Hy
46vs/Kl8FRbAQFeQqTJR1DSsZ96d1JlGnXdCz5FPP3eTckFuMEjDCe8Z3+8y17dsCSIco813cltI
LTajlam0CQUQXoz15LslSLrr3LA7AHatq6KsZuh8zKeDQeuxkuE2Ew7XnCp2e7w2t6HvtuKcT1f5
blmh8g6qC2Dcn7MIh7O1/ggK5PzzWnC+iRNyOfSV3EmDkQ5Z3S5xjVCwXV/CQ3Gd5Or8/diuWWDb
q19hv42mbUOKLz8RlHaveeuCKYvm9PCvXgAmWTLBpftIEz83HteYAgv6ByBsVf9Ef6OiyY6VIDFm
1TyuAzT58NnzYa/kUZJJuiwAYb6gDBPtKaGNtps1olayRO35+M0GajxEDHvrwUyhf4OGtfw4ptqD
0QmkCTJk6eSGepwikANg9yLbwkotKahpl2EQAwzL8TFzywifSa3hRDfFMmiSfUI28KHzms111dFT
tFaZta0hv/9DxG2ZS+v0swlaT/eI/L1kexQyedtLHVxVpqHd4paaaImBSR4GLPkURpjJqYpDoKIV
rt1+6nx900n64ShyHzJjsoK1Gm7ZkXbAo8Fsl13O2ViEKH9RkAvtmPnXfWnG5ySCRWDtwVKPTPi6
Zpkl3eIM/qW7MEjmA1niBwF167aO9w8naAdLCi8qFir54fvc/0P2JzBZ+doEKVMbchE6fAt9ISV+
ShBUkjr4yxA4IuztoBAW0sSZQZbfWt0qRHmY1UHlHYaJUIgm/okyGVlz8ivbsV6fmZmcgZLN7EZL
+NcPVTptYZja6qnl4SK8JX7fZ4PjTRZ1HGzj32VhNwufum+eCHT7DRMXQPA7yWNnYxLaswYsipD7
aBwc1x4/Qvn5LnBXzJnf4XfV/wJcpFAEgTEtoED/hjFsS7/YWxGoyLctqhPmJtM6Y164xnYUDRro
j+HI+r23Z3gK/qn2quU52VCbL4kypG6zGZGKr5F+StYxVAuR/NBz1N3B4TE7xUEaljdq9VdQHp00
u3o875mLRh/YL0UgPqX4QUOM3oVqGjHnIfD+DtRjpczSteh0DlfhnCC/lCwD250+EejvSnJCnL4j
nfWByHNZsKlN5JFJ5fcA8TgjhwLpV3gRIshgSXut1WbspR/Bthwtp4SAMNHk+argYwdi2sxWRvHf
O3N7NMP2ZIq7/nOcX+5a4wHygH05jZFdB8bkqAMx+mBoXDq9OEifeSxGOKJS+rhkH1nzp3TOkwvU
eU1yyRwT77si4n2uduGeDZe86FXK3f7HLON8PpWCsnrMOFZY937QsSaXZKpz4DfIEXyEaZQj8kSR
mbqOZi+uRAExMGokW4gTqccU2cCDje0AqiuSVsEIAW5Xeh6wY6BitfrGd9JcVkWBJPznuXcfL3EG
++8Brb53DJl1WPvj35OHaRRPhDpG8o0WkbAm5yMbhOEO1EQRFD1oFLEk2A/wT5VF8SArzM2p3pbE
HbTCGMaCm/NwTajj1e/2lZDU9h0wtpiQMyFLGTxU9T2H00O0QZL/ehRrCoUpHPF8eIKezeFS0NR3
D/DNOPAEimsQ0JpC869Bj9ud8u+Hmb2Ra6z3hrrINNj7FsbHp1Uux6QheaAIIrmCpUQB74SZS3A/
6E2fxXu3mVA8QDfEZNRfwtMLeX43N0xwI+BEw+7hbZT/gxPagU8aZCb8oeRn/dy1oPFgUZmwdYwX
sx3tJ8FJk5EdT8xF1qRjQz4ISDe/th5YjCEZmTtAIpLHW4Vaoqrgiaokjo50tpaakkgKlQwJ+oNz
dwr4OY0p/YIS/6Fb5yybcOKsW2CEtxYwPXP6ApIXJt5lGjx8Tqaf3h9f0PkP6b3I3n5wezD2mQPP
+suJgUCHcpqoNMsel3Vax31uhsbOFTz5HQ/KKuiFif7GeRAOTyCAzeWYnf/wmZ7nL+0zKNJaKP6Y
Qv0DkRnz9UmXSp9AOhSeuC8st+tFUOJSPSlNG/lfmVRlqKqWtogwOYRQTys06kQ/GAAIvdgXCvOn
eTkRztJMEqlrro+/WyWkHOGKOa2+vhukA/ioXA7NF/+8sZ3AhAPKyGX55qWmv8t53XZGh6ewuGdD
n8UyZNzDSpOt3YkKTqux8eMckXOh3EzDaF8NunNjvRtZuO2nqQnUXHunSvLWGqzqDaDu3kF7UTWv
1iqr/SKQ4R49ao2BORViOgWpULVDajMS3//+cLBJzEkBOGM1/l1XCbcG8YmjwNPgJlZ/YFLz9Hv8
Fj5X3211l0whzNxsfBAYYqFGGK2A0oz43URh+iXeO6QGdhbSPCJFYs603kAzMM/RDeahmPLRBJAj
LvKNWj0R/5q3hEWHcAc9W3GQ1a6Jjg8/r+bkEsR0kCY7rnz0KmZHQMSZxcBDsz+H/0bONN7CXFvy
PBdUdYZPglGWOGbpYj/79PnIw6AtxKADlF/1YRHaTB/6VSNNdxlmT11T3VQfBuuTb/ervixFUOWu
ovKedeHls1SExvYkLJyOE2azJpWNToXNcU1rhO8jM2rhoudAHdng50qyUlhTxLcpUa5QW+k1Y502
qf8Txo42X5+IlSNNbtiAQMOUaSv/J1trkmy0ly7mXCzwXYW5qsac32JjqfRvcOZwWmchNg8cQLed
07NFMHwkbQY9L11i+moydX9RGMzMHnRAK12k0QkRZbzDJwaHi+nb0C0PG5SF0B28KbAfhvx2o98R
kjL5Jh5HUBt+kdgNSw5GxqLfvfgUkuRDGBJKxwe8SqH3v7yf54ubskIpZFSPNvGvw3DiAkiddWys
oIiOFcS2jHBYglQ8iKlef75hLcquBQHC6NuYIhfwUSeU8U1J4xZhMy9fM580rpx5josr+Hop9PNU
CnpQPFzxjruEQk118G3vjAoReAmypQNb9Z4LoHFlk7016sysB2g1qkySbINQduy1QGtcqlPZty4I
7pamqv1LbXYhUbigiqJGlv5kJArgTKuxQYEGjh+xhq2eY4InSBYNrGReUx5MGiuDXYlGcVUdLa6S
cvT7opc2usCtrVNFBaDgosQ0Gux1vAS5UQxTi8YozOlU7Nn/A7d12PfAYuHIG6VqS48Psu6B08HB
KIsGwVwdSy5kNh1/YJsqNQ+djVOM47atkfU8p4MwMHf8EtQT+POjr+tmtaykoNiUKeGGLtZjTXdv
asxgXN9ipqjoGb/KEV07ot/Ppci37i8V9CBvOe/bqv+cEpHTwK2ZdO8ue+hfGj6mjhbBgVeUgac/
I7ensfvupeL0dh+AbDIYzoGeUHN1oLlxCIQu+zWK3cnEpiR1nyWvLZdMCmo6ELhH/kgp+2gOSqbi
P9u7b6KFiyYiolMNU4VtmV9apIg060W++pRNog2JxEIUDQmoyN/o/GCEVxRej3IsrFP/3rrl0DKY
/vSTHyPTSC++4Pj3ZqVJ3xW/L+uJl3T4XWxe3+hr/RtKAbZ3VW1laOnFW81g9lJYDrdNGqBu4UV0
P8EQwrxOn7eWOswV5t5ygQ1TkUdfyxrpqYFfdj/Lhyx7Sdg0kdrZidhM5Ss6+vR61PBuqmZolQcB
GbkdUtDmELef3QXaf01K2h7H+ycmkuLZyOF3FxY/kEy8aYM2pPhznzHSY0aE/JHUT+Al6Fh6Hct/
Arv/9d5aR9/HNMR/A3dnWfkKXGSvC6bHAcis1BmUoHDrtpTHMRJiNVUVzBfBregprq0OEKkiwKrZ
oRq+v+gSO5nWbsYmEcC3/LLRuIcDj5inRaL9zRMqPd8jH06HakR5EVE1cuuneMfNjM5WlijTI+f/
8DfK1zZg/yLFw14F3Hc7FEk+ulOXFzZlB4hx2/r6WnHWYAssk6ay0CqvWmnhsWsy1a7Q5MJNE9yV
I+UKk9occ4HHxh853tt4aB+ZR5zCIwWp9wR4cer6rEctWUDTrWqGc8UKmi4HQl7pVX83qk9jbuAQ
TT6kdpGRa6ezY6C5034GS6xKRsnNDnfMIfXMvy9gWgsgAQveaFX/6veIdcLFMMou1LPBNphjFGnU
4xRYAPl3R/PEUTa3Bkuw/4miIaPXFORhp6PePUNzN2Kb9t/2mihavA7RLDq8//9cYadmA3x2D0vc
2dhK8efuVg/Khu6876nIP8N8j80GEP4+Oknhg/fF3ZEEHcYZVHtzO00WLDBYbLhcT12QLd4XXoQK
t6/M2xkBas52144liT5rVwdgQAofjIrl9f457ERHr4lvl7AgVf2YCO6mHIK2sR6WmGjcDLSxYAjJ
eY7IRJRbtRb+dBVTfu+htJcxLDeX8zyCNis6X6EMAYqAQZrAUNZNPYZ6mCzXWOwaDERW2ZfD3GWM
pyKvEW9AoB453lq9i+u5pV8tT7SJiCNwFlXvwnMWiTfAvBFjUQGsRQYEfZoukgtI3UdWyf9yEzZc
wSB70hmIzCi35+Lmz9cgDLu1jp2HanvhUg45a1W260mdsrWhQFT5tGVLiGpZx8zVN7cT9MFAqk0y
WMeby9MflhDR8ZOgshI23Rr+qkBaMp91RtG0pudA0zLQM1rCuHcUTW2R2XZEcGGQ5uYm+ryptDml
e9GU8qxb2f6ushuyW98nU4jTyl3/snWCqf9OElfs7Xyz2QXGymD4UC0wa7kZDVK21byokZeeX5lQ
z/vrb7deuCWge93ZB1EFH4UwHyH6Pdg6jDg/wH7C53C52mTqDRD89kTM5x05bu4Vfvy5WYJa/3MY
1bDpm7F1AfSE8ZNtdkLHmijvWbcNGjAgNOKLhh6fc/gW0ZZBlHdI1hNKSYMk/EYNZIPOxmwU4i9s
qPLqZ33UlS1YHpZo3lBbS1cogr/WT9umbry5mIQiJ1O/YcTee2DffEcg3f7R3ZZXxIXduPKxaGRY
H4NFQTeQREhFcAyALQMC4Lkk5VkdyPXzu8oVe0W8eiki6O3uwJhRQ9lsK+FTZ0u7NelvHQBYJ5qH
rfJ7YKqW+BO3ypwr/wF8vhnithU/w5bQPASvshdZTQRH/NX452GwxMpnhgmfSknQzjL3q3Ci98U2
prB8Y2Opk+0BASCFe0k3gAcUbqxIG3cNjPFTTm33RRB7hLfzurp88z7mXz1ji7t4I9tlTbMiDdA9
hKxWkJXllprRkDoZ9AUprPLjYkEhiSsDGM447gRNCDxMwLp7p21k59L772ZLw9oD5SENPW3zOFPM
y5BjAtQtEadJTFQQ7PnTf7xTAKQsO0yjkkzpKqYO1rz2LzBu/dT2r6t+OGYxq0rWOMuNv7mAld+5
buQVA81EFnTDbOw3NqlWtPs1gPxqACulW8VZN9laTxafPk25jS3udFmE6Kmfifs6BQw8RqXqlGqY
99/2eiksY/wmamj461lmAWA7thACsI8zenPu3rBifWx/AYjbV9dQZ1Ez4Vfp4z3t446S8CpsCbKk
vLa8CrGUikX7gx6ECdoxj1tgtdj4LM1lwQ/KelGQ4b5G8Xe4h/HWoS5kF1ohCIMqvdNQJAzAvUTm
ykvwbTO7mOsfhB779heGG3Jwvm4oAFBEnPDQUF2fO/Ch+/uBRIiC7UzoshQif6btHhMaMi2wUQdS
DjpQ387hZyvZaLVQ5LA7aXgqfcffEFy67iY+F+EV8Pb1x1Lr6enA+FL3EMhR/3Yfx8rB8TjzVq9E
Ug+ysJV4BlnBA+4win4Rozocp/6tW8rIEc3Dg+Zhq4gglYzr7uNfTwTHnaD3i2vPiv9Fdaynq1OT
Z+5iFXP6HGEihaDuXVnhp2tnz06ibiPXPTT/JmlAWt9CEXTlo7oC9U8I9r2ui6WW20UK/u2GG8LG
BZvDm8KcD7eXmcvuipivDgrmDvlq9qfD3fzKd3lT1KACeXKuz5XvSOhbMqkoZyz4vsIhwGIL7Krb
UhH/2cYlYLS/YrWEW29uK9VpXSuAjhYjq2qYZzI1/3ouBkBzejDxfnBUUVBFW9P6cnuqueYS05Me
x0pcWW0qCmPxXwPEWS5AM4FZS1odB8OddK5edfUdvjyR38MTNqrsYSsVXYw1gLq7mWnl1SALxFbm
iO98MZwCNTFNU8YXMQ+sJ7VPjLPLDc+aJ05i/26k8PpTkvwhBmvzBbGiOSwMjb+pcGyGbLirtX+w
FCzJ1fFw5tt/5VAbpzO6UaPGO/LBoiKaQdiYhoRNJy95FhsbAe083svbJdudX1NyW6vIoB/8MlVu
8R2PTZq4EtpqqJRFaKQWX0WCc8jRE+Vms8O6xombdUwUmRcW2VbmkbFeli6xV488oXsj5CAcKJm3
ogd0qwsI74ztT+S1SJ8cjlGqLYTH0h9Zs607VTmX4EgvzwtxE9OmIAVagdxnPQ/YBT5elpimOgyR
CpYP+lXL+AkC1W/pFC9/yGo2IzH5Qy1k/MODWsbg4XlTWZgdfMi55+silpb3vdOpGiSMxr34yWOo
UZrjrmpEHE7+8DcCFPcQRNXXqhRgdhfWuUE0EDJAFOaVYJZoMbcMvNdr3oZGTwxjaKmG0Q7BBOG9
w8/xzTrtseuJXaSOYNwWyhfbs2iXZqBuSoknN2SHK9OZ/w6ZwNuB8zHCbkrSHSEarQ0w6D2fdSOg
uGxqgg76W/hKqNmTqeGV171qTfMXIIqn053YKVMVJ88H3fI+Jeg35J6kiLtdXYKIbpCVgqcXGiNa
V9wZSNPbDWsm5mhlJOqUf48t0OuBJ/caeXqGucdUkQlQkF4u4tXIUduLaFF60W/352gOxg46E6Od
WG1BZcedOuNw0CMGwRHWyyNTHlGKQ+mCkSBiEiGe8WtKTYvzUNNwA3lg9hiRhQBpriAJLTtgwJEi
9jdBU4RIl6qQQaHOcmUQnOpqr4i1PK0MqEdAXKvz773MQEzXbdw/pGFBv7ReS+k29eD/eKCjnp8k
QPkyepoDLBzH8pFWJllvQ6MzPqdTdtcgn+gv/ZkQzv94SaPNR4XFAR2d6JiWRv+a/A99BvcwsIiH
PAryXslZ8TrJFsZjHeWznUKYA0g6Whx0Ov3sZX0FLFMj4B0EiuIb4fhakWa1CpF3uVjtvl/BId3X
CRBHqMXbSw/Llx6pgwfysRnI/PH57br8mv6zmtjG9hcrUo4a3mr3zdg0iNLAYswtrY2UzK0Agy8/
xsPnJjomA37Pyr1eJC6TAfzg3ER8DldU7JI7ty8dz44Cwiv54o1/OGqYoJ+O/PJ5OklFJskzu4wr
5L0hbV2Wy9XVmgunNREw1+H8dPWpCUrO4N03x7CylEpJg39K/TvUpl2v60pbUF6o7Pc9F40K17Cn
GKP6gxSPxKO/l+PFj9ojbQBc1omYyAbsC83OXO+D5qnxKRE7TAstbqaWZYWeeZSQHq+5pNB9Os9S
h0mSuuM6/BPLC/o52RwPtWO3M0fSbMJQ4dkxzyQzqnRFtQdGi8bYlPhVG2Aj/x964emL42/QXSsB
qajDcQh/FMI8GTlJUUGHYusl2AA8SKZ06CSRMNqK/I0BeIJa5V8JZWh8Es6u/Az+fSYPofnSjNtc
meZUZE051ALsq/hjj/m99A6jrmhMAXegj0x++0ytZINwlbMwqfdB0PmDKAIr+3dwK6lMnVCTHSx7
jX3Wrn1fGDh1/T46J5pJTNYHrqj/n7M9Yoe8EF1i+t+asB6M7q6e0n6XGY7ZAQAVTjPmPD73DzAP
d2M7h9ypgM8lncthTArLhoOArsKPteHQtMumLfkCCt5hZDdM+AKJBIuJmQ9qquVlxMt0rsa9HKxT
3zhppRE2lNRx+Yiqibn+ySCY70zY2w1Jc1EfKddUgVW1Rwk3eFJ8LaWgdg0qAecrhoz2Y05qI0xy
4c8QuoTC444V2+zI/YCPr9zYdgiTbbC9llRiz7RvJbYYYVCKEPDg3OhP0DKDLevBzBpg1sKZmutd
Xo2xtGgeQyoY7B+zgON6i6FLDTj/ZRePn2bbsG49ulUOJ6+shwx62V9gqV/UmtuPK7UFHFS8911m
g4YkHViTpIENJKuL1oXa0fh00yvOr5P9BvuF9LmiR5FHtM/WQ/SVedRq8P4dG9ELnwRN8TAqiXIj
ZgryOwS8k/HXexPBIhebk9IFA+SwvZczLqwcae44mS6aq61n0Tl0ZXHiIkjEa+8j7rtjWyD4yuU8
PfAJ5QrY1JLSppOiFNEqUu2fz8Q1yxT0fUtSL8b+Qo/JoKROA8uMFwxYpxwAOaGZauURXDPyoZi0
yt428NLDsivn6h2VEGprExmiJrozc8XR3c8Hk2ru6cT2HgRJoPGoZmmkeO+8vaNWcblxwa73eUSS
dMtBv5yt2rqKvzAK+eZuW8PvWyz1o8RhrBO9xbOkEEVZitU4/unZbM0U+PiuuqGFUm/9Sp3jrG//
YGcgU2OJhOQMAeE3iCmns8xBgUyke/MgX87PIaN4A4nhWAA9Px2TqBz50EqNpUJIpKXZFcVPIfxR
Hk6eu5yhkCYxS73NSh/CwurNLTAF+kMn0CydCML7rM+KIDeajkrimt4iN53OZgnKucwLzYPfQ7Mq
Mv5k2jDxrROgtUvw8bqr5ysOFKZ5Q/aFXT1I+uQ/YHzzlZ9U1ERR+ZWulqgr/P6oi7gzRH8j8nXO
FBBvB2eMrrZ828BoiQxSkoCJ+C7VXUyIf/SF53VwCmXg0dY3cQNrAUoMByIvgeiOhiYSDuxjFoH7
szz+JGK+SDfOYfcSrr2XzanvwbVOfW9GIjJkMe9yIfKHdyE1GTxkA08/h2XYIErJj2hULw0ERB71
4ICeeTStHxffzY+WLfXjrrXaXXsMlzuty6W5LDRzTxZetnUwAzSMTC3pHsKiifrKtRKRrIkOX7/i
xiRdXM5gR6rFY8SilK5lRewxBRd3JWPWJIDOXIPt4PBQKNtdmHi9FUf+Yeny/OrRY9MQF88Hb4tg
aJ2NGSNQjT8hg+4lgZyIs2snP3z8Yekx7YrtGswt1LsmCtuD5MMtlaqUrUGnikWkUpa20Avyj8ot
MFE1Q6PRi60PXimGbNgqjVzYibUQ1cUggD3h52vFHu44EPQ9Izr+OI+rUt5Oxzuv2e4Dhfz5fKex
16jUqu3iBELJ4IhCNuVKVrJAfAJKD2vkciEBZXKaKn3MYsS1giblrkO5oxhv+WYbEQAMLe6qSK/C
IIrC8L4E8XiB0ADVrIWUPDeL2cbyfwP8Q/Cj9r/e83Xig+tUmuFlXHoX5L5EWvpzith0NpASpLHW
/GJ9WLDYQVgOv2ZK6Af6/B5tx3TDFP0Dmohs0zDkM7tjHQ0ma4VfXvCBUqHu6mFiA5yQSTscZymw
XCPa+GVZ7/KOZGq6xZ07ah6HJ2S8/kXE4iJT+npK3VGvpMBRDfe8mnklO9uOJ+UEojOk4Tb9lYDu
GPsZfkDtWfoRPW6lk3Q/PGnEXmPBXw6RPdOU1ul20P5OToo/1IRo9QkOtnBEjekpmLSqkuxo1VQE
8XVpX4cqI3K19fYc2iKChR+nBOvpg43wxytqd4g1rN2QsC/ZNKAbO9+8+kr/XRfDyh4CUczikIgn
N41BidPvhvf1K/wrGFxfRkN/+Yb9Mwnk6+YXEWHRon/L47MDju9RpdFoYSj/bUCOCPUpDQavZLri
KtmZqy9Y4hk3zpvWOpUQpOxWCMrUxbwk5knRCkvYZFS5x6YbOu+Vgl72L3kk/TKO5f047/7e5gX9
qIeuAyPNxkdfTqSSqDwmR8tq8tOHWevgclajzOkDgSBwXXPh0qZrWX23n6cZg89P+0EM0YuD4XMS
YO5OSQeky3aMt7ysA4rPHweCUZrkL8/RSX7WNnp9qZVhUWK8Y/gwhpnTH7YPeeNVSmtOMHoTMv2Z
GyUTC3Dwg5E8NJb9adrCJLWtRazzHCR/6M7JYfft3rY5fT87rSqq1lWHRodu+ZWsLbSj3tnBFBQH
pJA6rbrhcc9Ug4pBMBBpUucUic/IYJVqUynNWRIMbbaKV02FHIdXPtuu/isq9b4ZgGrtY5xOtY0L
mFM8VT7TpW/Rzjtd8AlfnuHWz45lN3cxWHN1OEQOcVNaV3GIojPCrt33JhqS5qZQYRsLT8ePQTEd
pBbDar9yh7dxK2VeSUADBJ1oaGdZgk7IsfCSZtL/kfb9oq1j6b5J6wGJSFSnlUUC4RNUQWx/T0RK
MkBoN3CVG574k4SozAujSbf7uFLwtRqT3j2EH8VlUMGIC/zgaeqD9yt7VyBA7EN4+ddUY8VVBkv7
QGPc379zr0FiQ061hdwdbz+ylzde8ryX1WkhXHhgyAnByZmK8Hxohlxy825Wyi7N+2Ii6ig/ddc9
b7OzTAqkYzHPBsZ5rUyTdCs0wyzHrJu4m9+SRrZchDhlZW02YWqZLgPylHtnWzmfOPwnBaM2pPDv
rNehaKcA/6aMfkgoBH4UxGQY/MgIb30zJJmFYatXVYlk7SgYB05Y7UGKOfdu6VCiKNb5QoZ40k3r
0yXHyLVMAl0ODzAWbXleR5A6ac75TPYn2m4VOu7jWqK+xS7a0MaFOQJczFJkw4wGUrYroXeq1HRv
a/p4DOLq/+24dC0o1532rqlEAtAXKKSeJq6bDLmjtDVlawhwslE5oexUlvGHt1OoKBGI+yehebs2
mKp+/LNq4HX3vVUgKr6AseKL42ds59zdT6gMwdQMz+yW1EBB3gnzd9cQsb00FaUQsQ6749e/RimW
LzVj8vSeDSpKokTf/9gYLF68XekQNVnmhNZ5tr1hVM3+iE6empMDH2PfAmLTm/GynF5WHWwz6xFH
/7ux6ELmqQjwxFsnCCciXnIjPcNzapGpql+37HWIptUsXYo/JstvzlATgKNEvcyVidxTTeenHFYR
DRc2Ucyc3jEYNeIL6DuBhcPxKmtyTYO5GgCPZqoOTmxR00omMOLuPx8kfLh67WohU0hv8aEoiOT+
iTvjTGgt+MHlCZdcvebtaI+B60CJvPcsbBtGhPljiJLcOSyRv9m2iEb2hS2kiWIwsPFyipXXKksA
SfJjPIuDr/J5Lyd5ygNFSZ38y4zUF4+miNaIdHaVSMDufd4qwv1fcaZYyVulhqidedRQuw/XbABC
0OhpldqGBWq3PGXA012Kab/gifVTYoJSQmmo+rfgay73F8cq28IczN6gXsxWdPwFyRKFslZY1Vhx
BtOjt3S/nRbhN9SFsUWDWWPwZ3Cbc24NqDxpYFQAAk7uv8WGGfmWLUoAbjjI9gjwOz3BQNkJ76x/
puTbmdcP1EUh0pRSxj6LdmnpcKNpB7lbmA5LBqA8pvCC+9wAhL6HGnPn/7e5w19Pt9i30Yo5B4av
DlrgFa0RQzE1gJk22eJq/7HCNVUBpyqldseR4tzLUPSwaQ2+rhwe740yceAewQD532GP6/jCjROm
41wFU8g3TS5qdB10ir+mFXySYiayPegLaKd2XqO6d6pPbUR/0HRmdevEQjShaty6V/gPWkVBlh7C
y4GAbJHAgDUMMGq+nO9G/YCpYBezRKB4YtqTmqoRYZjMpTFWQTss1fyg1stN0eeKyXLKDETzOL91
iAzCBIYDey/mMdWYnrOXwIdtb9q9kwDM5We4j5L7xsUJf5DD0Se4fGZoS33aJEKnfHqPxozFpS8Y
gv22pgGin4sD9yz5ZbG3F7uy36e98NZSBkJRNg6Sgdu1JImNt2y9jVAp07M/7kZcdCpeuIMxM8Hx
hPWtKkpFGEi+ZcI/PoaZcjXZ90AT7FJVLgGzphBVRtpugeJO5VGqsZAbeQY5F4F2VDSiEdOlqn4n
mcMhYPIYOSmLvhVbsnkoGdaw03azQM8emliL/egDeQom6pybx2MPxqJ/3XmGjR6LLZ9XYP3UFOqV
S56jnQnTor9WhraC9EU/P++MCpU6Tyt/FPmTZo3Ipyqt1TUFuZAGL0A2fAF6x59PteLjs4fE4Sap
DMQ5SKRMlIjX9tL9uJqjDvXzqPrYcwWbvev+XQgxv9Awhmi8FXDHgzLtN9fVnpXEJ3P1BIn2vtBC
YKNetHUsz/31nInYVFvExld6gqUKdZaX0F0ZqaduEcviHDslkErTTtpo/XLed4BJXHm9uBdoGd9n
Zqn+gZ5tbB2oAzmKsL87iM+wAG5eNSz7ZqyvdKd7VSKqQaVGFwQ9kT1xKBaF7E2DlXeiHzUrJh2H
OnS4U0FBCaHYJ+N/M8c6Db9CsABq1IBrQdIuE6PKYvxsStsW7fwiIB2Ps0lTg7R7+bNg/8eLRf8a
RAvmPOps6Z3rG4MFpEZR2kuYat8RbzG9GRgSFrDecbJFJExqvBPfPpcT3YfXpUT2vWUXoXE6XqgX
t4TsNKFKVwh8PAEwmJbEJvvbolVfKUV6Xz7ReZQtMS6UwurPEQL7sbS1FCK/35i9QCop/xFZskRE
fKNWjoBBk4LEcq/ngxXM4p7xb6N17KuhR8rKTqtZOLKvXAqDZiOcWVsEyjQI3K1ln8rW7Ib1RrPL
nJXqVMS1DxI+2eCV6eouo7Ldp7kFIWobVyp9+yWW7tl6UX0HrZlKGffQXhm2xbTN6E8WmlnHDTbf
oVwyoIj+jJe1kRxWwAnjo9LTcQaK2czlvibTwlACFWGAaK1ZriQi32Z8mJmkjPIXhDjCqVu3G0Tq
e94Am8MTIIwRgf1J86Y05NIJq9vOB4yn4iKRBqF1DmEc3+JFm1bx/Gq1b6UUjMP5a5HAZGHloQkA
Mvx0KIMCU2hdZftBs4tI3JSjL4SeiH85NNVlnsmiZSmJS1FmEpKRRgPxJbds30xW6exUs3Sz2kIQ
BEUvnFC2WiZEX1W3+BZ1XJNK4c3SF9ZOVr7SecRBAwTcbTQ1543hUAC8nIS7PGT/WLbhuWskNeLi
UvUka3PppZxrK9XH0iA+7T0Z0Op2XDj/3VuSu+4bW3ANviZBCPE6/DWo7KiQNNGvmLwdotwnORL7
mOCgC1HSBs1F/XsW85oRZXO6zMR0Am7YC2DxUxf337hsxwTsOf14eRy9lHZC35b2k9PSS2H5dSYd
ZbE+r5a9eTmlW7518LENEcaimZs+9V863bZA3LG5rRXQWtec4UpioBdlakMZz6ONXME+LPNvwQNR
b/3m1Ah52jjaucnfjXBBzQbYv03DtqDwey35lYsZDQKuo1wEElu3hPIhLaqMtEm7qGbvd47shNAL
GdUVBQkDgkov1Dwk9S014MV3QLQZe4Yyu4/YkUGSbw3u7qFMvXwx03VurxtwJGUFO5NoEJ2S1Efh
b9njzkMs6xwQdIr9ipslc2kN0RmXwkDLyESY0Q5DBGSaSNzhjBSF7EmWj5Zz54Fl+N6I18eLqy1g
2ciNUCSsIkGThE16eZ5bhi0WOjtQbRLXZ/vAAqvl5Nj0KCojf2xUevv8lB2bgQ9fKBHQbs4uXJlk
wAo3UBuvQ4jnmxRDJprDmc17fHwinYtEMGFdU1uYTpPXvo9wgCHABY+zkd9K4tzELm77iyt8t6AE
nFRwUfOYn6Xb6qXbYrGuD/O6XLhOcfR5LwPkAGsYDfxxphJCV69QTHcxrzm8NkMAQkKLac5CDGxY
a+IHR560IVMBSuE/AjD3kClh8w4++lrjqxyvshMLAdEpFPYTyKMTVg+sSaqRMmuqY/+2ff+h41dG
2m0DtzKxNrA7/M5j0E44qZ/9oQUgNdw4k4XxTmBl29m6Lw9VtAF9tV7ZzTk1duc+y/ub+ahJ3fCq
eHTOijM4/onKBrwUvIB5ApsstwvxjRRKblrG26Ky6ot5LbO0T7gpHN2I+/sj6vtd/fY+ittI6nX2
PQ6DPuHkIeWyB+2adK1AwECwE/8kAWrxe7Gyg8c6v6bY78nu1Pr93Z6tSSvD1VL7DrRrfXgcudqA
teenoKkxB+HCTLmCnRT3gxYn7nL15MsTe4xzNx5pBL2Gh++vTT54+ke+cWzAo3xr0WdaL5Mv7Eo0
e3B/cpz5d4om/vyvPn+d5KEm12O5W2d96If8eri2SER4H65GW/D5b4EEsBiGekP8CpAHr7/U5HVc
pEtEoK0W/LNTE3z6V7MR3HVVjdsCEqUixN/dPDh1SeMmQXW8rgH8bPT5L38U9mWsRy6TW4xCgvKb
GDz4cC4VAGQBtts5n3RvlYA8NJalZ7iLjFLv76I/dmQGVIyu9YPiAEwz+NmpQP1IC6UNl9zAu1tA
UOTD0iC4DCedmOvXeorZ6Ml4qyeT10+L+7sULi5wMW6mXSyeRAI2Wblk33n2Zk0yYjCTXyqrzi6C
/7lsNVBohcxei5+17f5ytcikRujgMo0aam9rPzqVN6ZSeqOhdWO18q3od3yKaisSgKRQKjKdNlV7
mUFwc74YY4j3xV65/eDeFw8bj3vbp0ibttzKL0To19yhR7nQek5qmSobCQG+Ee/y3uMamiMwNE0p
AlQYVRSSSqWjsDJvOdpeX3w61XmOGHnxwyfHZ1MX9XP0Vs6zGEPaQw33Y19XjOVFaUmAA7i8J1sN
JXPwiV/FrWrINsLL29scg2aVprHeA7e6my74T3j8Vbz/46hIujTWPcWsKqkkWqMih4U4wFzN9S6n
w+6iPOo9rwG6o7iEFb0z5q+gOKdE1kJijIqXsgpZ+9fkwF4d4Ew6BdpFez4B9cq7x3ImH3I1ZEsR
OIVRtD78lt0B1xuWGIA3fO5t+z4fNRbI6ao/oU8ZqyWqmVevH8lhbvRa+90cXh9ccUuinpcUGsXv
jDT0KjcySJQwHVeVN2oVYqei526QhJqEzQ+0i4Yz7XNJXROtT7bUWI4Yz57EnFXrDJr0EKY5RKOJ
Uk429U/6L04ehlB/Lt3OQzhoZFgCXqaJbW8Pk4BeD6H0OJ03obaNn02bLrCvA4lfob49j5KLaIQU
lHadxiSV3qeeYo+xuMM6Duf52lGOVGAaaBNsNPrDwVtCU9XjHgNSGzKYGErcvFtwajQSvz1VpjxP
xdfpWKvo7Pgmquax2CCwnWP5xYeVu21VXxTHCQpGFKx28ZOFe1xS4zXvcIugiLN631ZiyF2PMWRy
frdOqakuInWLhoxHt0QPuWvbsZ9kyswhr+IWdej80UjZ7TT1By+r4qAHvtrRyUbSSPKKPLMsysgu
3b6xs7mnMnrJysML/6zqRTAZgljPtRHyKSw+AUD5SbXTJzxWSHQaRO55r8/r1/1aFpYZZnlHRwsN
71Ux1JYQm++06CSbYUkYRQMUpntq1PitkprDRk46sFezdrR7Q4/9I+sCwWncw1AcrbGtkuztm0Lc
WhNzSbyJzaaEYdnKCLPpgzc0V40rcZaS9Ymh5bd+Of77Mm87uqbDC0cAWEQG/v9SxvWTgF8eVcpg
CB9mFxHdmh4R8Fe3fVcTjj74eQNsOHRD1Yv/B5h1JwLKcN0aqaAhRwYda73FK6weFtC4C++KqMYQ
vkqVcRV3RCrEoVnUj8bVJflKztLfFImP8D/daiQ09dazrsYt2Rr+YwPIo0+yGGOMplyKyTzF6k+M
OcvTK4SrcMGTmONiCg+/WL3gN9sXJ6lPuPnsA8F/fJimOraxftrY03zKi2CfW2mmZuLr9wHQPysV
rDFxi4juFb5uv1S10Cgnzhn4rA01VW/1vw/RoeOBoK08V7j/niMecS7/SHiu7Cwn8+MxpNLTFgfh
dAEc+MoxJD/TBDDwuEIkfv5MgZaNT9EqT2NSOGXUPZo4dSB/GXWCdjfmDZjJp+V4jmR6Z60Asg9+
x3Qq6UbqPF70hDyQL6yxOaFv8k801PdyEh+IWGxrsPDr7wocAE1tsqLb32h7XhThwPdg3C3yWJM+
T5AflkMMk6tQ9HJb2NNGV1j1CvHzUGMVAOnco3Tc4EG0mLuI92le4+h+cMxJkYM5FH+S33Or0mYc
8itJF3rz8yejzeOWz0ySGOuprFCGHG3dajRWCjmV+m3w9fjshY6MVH1vDwbAN5zH2iCJ2a8PM7xl
sAgSTL/fmg4cy5h5e0fbY9BCT7sdEqK2supn5RKvNIzq/gNj8fbgjW2l8sBpLirBXBSvzVdgm+Kh
iTMBcdeVUTNsF+2cRHlpxH9BD9nXLDJyfsQnO0QhWloyFishyr6CH/ZWjrE8AnvgYWigcZnyHV+h
IMFuGCKnsscaIp6mqwmUY6+dvySyc6ZC+2DqqZEPz/lovRwNiLSSaDpEYxVTAQM58CIDvRVZCjOL
OV7vbZ46o7cW/+lvwrHZG0tdY+ZDwWxNfdlV/dxAEYLPaORI+gIXLqXICHaAixDEHy5Cq3m84gFo
KdzyRjhYCxGfgaoxlCyQMkZxAows3A4XFDi1uxeYT/EEkgyxsctqB2iYzMAM0wPZ5EAkYSy2mXID
PYM4fDS9rKvsG0hC3dYdyUZ2WOCThkheEzknNgKqFrhwV15eTLoU3XCk9ciK1dLv9WsKowd4l84e
3n0fQwidnwNE9/PVShrM+D/ukoHelqgiBYuAcWI3cy6QOx4MKtaxqNQCDQdXjK6z0yLUkRx+3Eej
kFMkRlY0DaXPHclLsNXPZP1K9mGbg9ThrISQbDa/LTeBRujqGtQEVWvUOXC8CBTf6jd5DK/jL/pP
br289K685C//JTajwCNjoJymazGk1AKNk/tV7aAJ90sJbBaRL/bq7vURavlZj84JRRPLm1O1j+QY
c8V4xzUPBiFFaZTxIgqkIzevhTAUHIJDfrVUi004R95Qj53zKWWkpSzKk7QA/zxSi73NLiaGDOEn
jVN/TabKAtBfY6tZ5VaC7UTif/WRNdqaWVH2/WIrswwMJXDEIHLryw4MOPMMY6t07pHFb1o8dw1q
h2A1fePr7ZKNSkZoFFSr1UhNueUn8zFUvTc2La1yRAmv+3xQfmoGav3nUrWwEOJ7APTWlW5KcJcs
ELnfw0xkd0q5ZJ3Z8d6/ZneyCrB2z4RiJm/Ww29ZEIjJGAvlqHrikl0DgA3ib9b4L/yoKrxT6mlj
Q2pYBDtgDT1dDiRjr0TlqR/Xn23hd0otJ/ApxZIfefngB5tX4GCj5AjEp1Zu06NWe9I9tQLBgB77
JHo+P0MkoM9OJdjK50IMlSlrgwIRNSpFkZpmTFDnZuGS77THcyUdvmTNQW827HRPwmcI5RQEGdzy
2rZDy50/x0D92kKbi62eE0oQsuY9+1G8r4W3DMrUHkmfW3kTR3/8BPk4aUZFzBQNZkC2qH57Lw3r
KECXKnQB6XwsQSpC/Vsg43WmvvGnIMQPpWyBsqmD5z/nGxgowdzwtF5Io6BLTkMcwkZoBoRamWP5
Liu6S0wdytrax9yGNkPpir7HA6I7oItvItUD9igqBaV6ozwpvKZBbSb9yGtI1TECaQ+QE7vHFruo
Fu6pEFg1UfSV34E4CFtoUoPpFn8hJeFKR2jvJAU5Y4B78ibS+p0LSUoPLN6bCaAj28tz/NakeYmZ
z5Y2v+Z15AKyTwq9QVWJzVZKSnjMPN2RCId55g8YqR37vklBR+7qhqhATNbh6MfZECCg+NHsjghq
+tCEJkiAdw/C6YDVM0qK8DS9RrL0oejRQUKR12HeAXN8cnSVEPfaAw0I6o1M4WNWGvQoWI3gh4zW
sxZ7ptAkCJRAOn7hl0PLSUFXQy9SvALcDWnpinuEOpVE2PrmkJvWWshqpT77LG0aJSTkUVe0B2ML
YQCuIWfKFGcaP750VjfsOYorMVlSPO5V/1W4y9OJgXJjg7meU3kFlMV/JD05d3Bu8gOy+wNrCzA6
UH4AqJkX6UVbERItB4MSOgeVEvWViLVycrD/I5Zj5OkAv2ZN6Mqs94yJPUG2kyX0C3bUTAoGQkbq
wud10cLNGKOSl05vbHdOJ443lkCoRW+qLQTA9dU0OScqrw5z1btOOf0+2okmfU8Bbk5Ne4zy6Jrg
A1ZPxJVmqRwxnHUa1t2w2R/I8MxtTo2WjHOJQK+xrRhugdzbhhzigZfpkK43mWByz/e1E1rnwfbC
sZxeP6tPwy+xtVSNX2YNqCyeV7GEenLB2fNw/9fek9rAWGujcaIduSRsPpdo9I+GRyDdG5vAULjv
mpeKp0mKnvugSJPtg+PXG+/KShxKhgHnw3S/rwsU6eZE56mraHWZOIDDL3MWqNIUGOTjT/+vqqr1
++l6r6Sfl6yiW0Gm7EUfgwKfqvxyu2YSFeTuWXRXUN4amxTqDdGsGwcB12m+mY/B6cn7jt9JwX9I
ku4JY7edwgAwca8gijJ+d+D70hN6+w/K2iZHCdYN8WGNTBszjkXhGt6q0cKYDyr7z1P5rKyR8ZC8
sa0G9S9tAQlpTY9cs4aPBgaZN45DST0pSQV/t0rEBMxt2W8R+aGs6PZmw8jN7h05vtYDfH2x5V0g
by1whHbm0XRnv+aumMgLh+qe5ZYTxpQ/9oE6hYoqV2hF2fKRBrVU0WeIqHrUafHCFkPmLdTAB4F2
cCsacLvrMHXQW641mIStE6ExOFx0Mkdd4JR26CTtOhyeupzIJJRcOYTqTWh46HSMQ/ycIdU46u7y
FbnPSHM/QxLRkb5tEgUlMASpALHJKP8n0Kf6VbUZPFOuxZHZEbHx1ctI1sJNCQQiquYNtq6BWOKh
3aDDkZ4GAk92CIYWgwc95OMPR2BbCvzjGg1CN16+ZmUiqLIBbVFP1SrFH+iKNW1dw2e9xP+mD111
y+Q55onwsGfLXFBSfhVgMm3Su5jqfbjm2lw+BWABy1Tz8QnBnO/koly32xhEjktnE5TD+rv5BlOJ
5pAi/jjcPtPfJBu9b9btNLSBf7J1PRfUYV3ya5qU7npv52mmHazN2N26Q7B2lyifVPtLL3N1vKYu
fdkUGY0iT8I5ZHDuyCNZsa+ROeQwaDG21M+VFlka2yfCAHUXd9U/GNJUmQyW8m1zvhuIWw2GAN4z
qie7BRnH1TRDiqCKxPubkSoZ7XtSdzpIZPGKxomSL/3LcbjlSwQ0DyI0oEdyoKiY9dRYhasZBaYh
sy3MlgV9tDAlrmWUeiSGP8VyNwDpPobdQkvhuSOmRsIDtGWTTqdr5/C4GelCekcmzBRGf1QuH6zA
31sfZe9Bxm3CNnfYdbDG9LS3CDH8EviLhE3k7Eb6u7mqaeJ/+Pro+1KdsZcOQtXYmeMYiTrCIjI9
uAx7WL1DPHYo4PDXTOmaNSHOgE6Q8nJSG+zyRkLQBT603XolwWNnwtfxHULMEndUA4og4nqM7Qos
Q8uwBgj1Rx2KKJkyrqxUiRQItQ74L6PsyKFKuXIy50LnScOmMcESqp1c8+Iq/ycK7WvhTnNHXAgB
XuH5mLKy+wHChCTuQyu9IkPzEceIE2sQN9ydPFSi2XVE0Zbs+HCaOVEJcSbtdY6YPe8thVxVs2+8
uUCx5m8qVWSPTLng+p7OSEo6eNbxgaOgY9kOEJxv6XDPTymgWTd3p8lHfHYubfwyCOt2S0/1oqWX
mfgMgGheO244k5mor1FsmHtrUJ4bmE3HWyJxCmAl/o2Wn7WFeOVmicD+IjyOpEIKoxG3dwQOOB/W
2BnpuCwxhSwgOMDYOfhQ71NxlnJEEWylZJFDahkGSuvTvRqKX9tqfO3zOiZHT4PReBg5Cqk/nxWE
xyvuTSumB4a5g65LCluHl5d8G2rGmPKL/UlUyp+MDAeBjCAJ+pEcAOXJLA8dA6e127BNC7rMJqDg
sXxj3TOPquMBA1QgcxFQBEeFEiWQRb3juqGw/kSIBEUCHFgPaWOmlLE3alartW6FWTHDP2nbV40d
C7qmq+pGc36YJlZJG25/rpQwK9wYejEK/ePkZ6QQVYVMmThIkNHCHlnBhRODopU8qJDiwrWK54Mv
bsoPJT+VjFZh2lHvdNkn9ZCu8VysXTPCz2oP/9JG0n3K7hJ139/jAGKuXWrGyJARFGev1CWXwMl6
jguGcZnEKJoaMfu5XTXDShFFtzn04bxTNJQ65QN811+FgtAWH6JiH+cDBp2tiSbkS5/bmCdT6hpr
6CqyCBb795O8h0jwQRh3jd6PLtna6NO+cwa6U8uJkLicW8Lm0p3SCLNA2m/NwT6m95hsXDWpLl9c
X9U62BdzResOTxZw1yca/N5Wd1KImppn33fPlosFq+JFIK8beWaIl+ULGiuvMBIWBB2s2XfrFnh4
YXUDE9D9x+AbtrSeLGY2MKoFuGRerGGMiZ0YfPtAkNajaXVu443XqNRy7nzmZQVE8rLnE7Z+3ePg
tTVer+9V73AtfuInBUE+6elgivQv3sUs6SK/vzE34CVs8L46CJhDhv5PYI/Xmi88mBBJlmOcH7Vx
ARAezez5Zkgw2IsBycva0DnbdObXYnMkaV70VMtfxrTZmxutZRNTVMW+ohEZz5R2dg0XWz0ZAx4C
DUk6KyTFk6X4jvJPtgj3xuqWyzuFh4r2nU4E+kjCM14vhVFOJWLp+Cr7qHcJ1JYHdCQrmoCulHW6
GdCfw0zh0pc69fz/tMjaOczde/ld//BBoL5Uf8E5Cc2rlIfeGxuT6seEQbYRl7NBOopFiY+fv1+Z
cptpuusNHI+zxJH5t59iuhunha+hHjJAQAr4ggV+bsCrJ7LJ192QTPisUxzUc1Rtz3lLiPaS5sA3
U2KG9mmjLZxKiyPoMh3QBMiA9j969aIss4aJJtzxyK7jhQ2scGr+3/N/hApT/SoFXEARUavwuLub
bFTDwAduO0grDIJtdujN/X2g6YdLJv44md9axR6n0fflfzvK2HquqfiPQkufmxDhsNJ1jJqDMvOz
iK88Ej+BPcMbG2cMDUvG+frVSsWIYyMaB6dJImVU3nmr0Fwep9oLW0NI+RHdWkv3nc5iYJkftu0Z
bqOIknN4pEo5AqjNJKoxUpWWeC8ka3MqCv9BgbIuUGY6ZZ2GXPguD65Nt5CFAR199zRetrc6HL7y
qLPabEr3PURDZCM3H4jUMOfH7mfoo8gmp3Wni/BrtoNTzLF5bHKHabfc/1LImR2a7aiOw/XghzMO
0SosKiXnQjlsKK7FzKT1IybfAosxpnr3fuhCajhe8pKLg4mjHiVV7Iz9qEWgfao4B7d7AcUmupWF
996Z9jDC1ptvuyd1xyt22KTKtmebGuPO52RBIso7p9fkQdvncVc6mcYtczyMD9Z2UmMxq2MzCHFK
+CTvCh7xyI0WAKavZ77YtazIDB71x31Q8nDvU3JdIeZMqwgL18RCqj+RCDmX1QDI7aGxHRTAOoa6
jnMSdZbfStVUkJe6jG/ytqANm1MN6sO0srr0U2HTK88TSaGEm73O/VbmkqZNimwGX+l9Q2yy2qpJ
+6wFPpfRqlZ8FbeIpV/gJxmzau9F8JDnvR+DE3kxJ7d7mchjvmlqUWEVgnCMYABHtYWDeEn19PNd
ftsvrkbach7CIjXhOwIMiZOV4k/a7lIg+zZMesOWAdOxwzI57sEz+6jSUNveOSntrKUcW/xjwlo1
OTZzUbESV8nnYu0y+baq6rOb8e4VJgSFLBBwbndXrkNVq57u54KsFaxTeuDSObw7JZm9IHHlSN3w
6NRZQoiLAROUCJcnQ+w2Ss5yvTEFa3B+VX9Ylr07gmzkh8geXLgEDpODbwnuHRnUyuFjC1WJS5gl
U8V4SXUjsOihOv5jx8RN7Snt2cgrkvOvJY/If+aBwY/DUoWJzXdJ1Nc7L8VgSbOkn3Z7uDTybKys
J7o+N6g0l4d0m+uhkt9ow7spCx5FfeAwIAZHDCw33VMHw5V2XlFfCzDla8/D9Q2TCQ2Lhc8fKHTV
4f2VEBQaXhMdd00x33V6mZCnHxfEXxOvBueHuPr6gIS8EgSzwPBgDAW7jVW/6iRn19wZr1a4+YNq
v28hS2O0fDnydKnRotVoCrta4GYMPPngnIv8+rjXIxhEaSAwaHfpz9eyoIGddKQQHqZlwf4DLouC
mf+yiUig9Li5aOoH/DwI48Q5ugYTNCNuB3VUetXhM1zgNP5JgxFunErZ5Vobuyku7dotjwK2F42f
Byf47xZNZshUqxtr+nlAveagKKjICX3tTrz8Ayq3FzMbAU2VyLqcDg4cxX6L7u29DevU71R21bxr
9CQ7PpNkew6QnhxMGN+3KDCXNzCipk1oJS9CeKbuCWTTkVCnOhgr4HbH5OMS0hhTwi9OWG35XQ0z
Rp9Vx6dWZpShNx+fsgx9YiWz5sqf8GR2mq4kElmp2t/V8pVDVW0yoeFe8aBHmrPEhJI253ffQQDM
/sM+jcNX+Wl7FdS48AUAasgnKKM6SzmN+F2hJyGU40FppLHIuBy1RjWh7W4V/jkKQKSDL7cQ826k
rMD/+Yc8GKfeL1og/hJ2IpAIL6rh1LTQwcq5v/3Oj133Z6Ag2vlk7+P1+Ac0HXqLMcfaX2bAcIe3
TAg/IemPJTWO+F7nBvy9Vtv9YaX3tbc1aaHfUK77r70I/0fH05bgavrLXHxO+SM0m+gNQkHEWXr0
G7e02N6GkLPK4oeOB+pUsQjusa3RMz7/FUMG2SfLEJEW6nfLRFurUjdoc8XljnXTCXGyJmkYo4su
/5ztGWierL3IUaXzQUBWyWReQYtPWjhcwdfbrYstsylg+a+bscAMmKzfBWHnh/HoI8JtK37XtYXT
tcSJ4cakqfaSfLaDO3Ru4+Y3XHaASMOl1Jm09+HDzd97sCY+qRfy0h71+EH4Wxp78TT+imd719JO
3tD/+NHjCZ48ZzwFusvv3Ee0xGSvTVLDYRw8yNvmdZLJYy/Dv9sfavGoyIBFjK7HAGqGxXkNOs1m
fK7jwNcoxwjuu2/Rc/ALFENIxZSLV+G8FilS3CH3hIahPne8rTdI1YYo4VclaFGgLgyorLl85R7v
93WCo4nX/1T6ea4rJvGLRwdMysUV0/goXTIzrMOqQEJAlZ2c96z4nbVMGUwg9haKySZg7jP3gYY9
lFXoBnIw9TkNDNPe5JyWHh0I6a/nl2S+KeTpvXtWniIzwQr2S/k7194ChUMbSH4gGUYwiT62rJQr
gD7uXOrYAZPo4VSqHWyapHWIvJq96RtiW9AN0DwEwvfy4EeOkx2CFUOPCLCKVesFmnwPbruI5z4K
tMW2CDPNDVpenYZ40E0vCIDWBiAsDR12EuW95nbWKgEAai9skFinBJAzEMsyRbJDKwBrL1KBiew9
8PgIQLSqw7eBuYxOklG4GwLKjThSho9//oi3iQrLghkUQ2m68gS+gmEhseFAA3tzR9tpqmoNOame
hTNdx9JfFjwrUUa5Iu7EI/OyjoW6E/E9tAljkEovbxXUBRIUEiMoelxo+UP2mFvYDtw/rgbhw4Oe
50ZoNjD455ARjrpLcaRpTTnTmnbwUVtt7KpvNz3ZTwc/a0oVyrkMzOgpxGRvbwYK4OO8hmBgmx5O
u/1RCvctcMdjIpmq/NRRCfMTMpDSL9qg5pLfS/KRIqO2YB78c9c9n5I7drgKOcY0A9E0H9mvuv4N
JVjD8/vsl6IuvrNyYKKApXDWF3F3HK+o/yJtCWH5Jtgbw+EfEZgnpgQeGTPuTwTtSb1i7tpQpW4P
ciHb6W1lAdYET11GrY4LEyetraBeqCa/9R15y3Mhx1wUKIvwfl6iRspAm9FmhwHYOlifep3T1rpv
Bi6jTAN6vst6nS8Zx5PWvXtEBaHr/tt6F+AfoKfG5RVXcpdDSejxqkhzoAVVNa33Wvu1G3vMMlQm
AeHLiUno+fUGxqTuucitMZ7NVBJIzYxtXnG6tWSjVInUcJaiqT6xbXeSI4nvgl1E4RgA/QmbsCy/
dXy2Sn6C2CA95827yzrlENAb82pny7U3LtbkAShIBeZrbZlNb8Ib9fk1Eu6CkjUGZ7myJeMZf7NW
NGZh3u3HhRcF7AY8eq9EyjoSn+AkmU7DBgA6DwT+lOTfN7O8cS6444enKp+yxn+9uqaToWRJWT/n
ThztV+JxZEOCWVvlQE8jLdU/RuJOrF6C80LmZa+9QzyxN5keb46fJxhmAiFU9+rWIHhhqckx2J1s
pXTqPtaOsiZW7/kSMCbFZeqFdVtXGIqC0EThc56fsiZ5MijMJwtyWQUo3MwMyVofSEK87T8XiRHJ
o2ejik6H7a2r4ovZ2uAYyLRwI7v8a5zkB9dIrojQTPM0zEiS1F9unkkrM5NMqQ9WNY/155c3OdDS
I7Ya30dn4KfkC0MeAfBOK9nzXRo7dm04ilP5Rdtw9QLqL46nQl2brkoD46lmvI3HqYl6XXkMRxJE
uruBmUrDyQaEvJRM1rkpSUMVhl86WkS3615zKmGFE+buqrLk+bD/CZjJTd8U5NHAbZSCshekgJIZ
s6HRlK7tFNeC/DQ8qcnkTxwf1V+OSpu89xJg1E52hHsoWGU3uNuq3oW3HRBzBGl5VAGSv3ugMs7S
VHLxK+O8QbywcYE0QMDQ4XrmWhTt2omxn7Dx1NYdZgN8gZze+FbSyQBz1gmWn1/uifzZMwW1gR55
bMIDFNXa6JYIja3H5uuTYR3txapdZoF6lY8zQPK/Ijd044L1D2cFruXzgNZjZGEEWdVCJwmyBZM2
8J26glycN9dFoAyugpfcpvs0y03CSGBKyzAPkj/JJf3FRF+mRUvLrNkK4SA+nGzUw/SNxB/OBPbk
6yJm4PNiGjisH9zSqicHQ+bEY+LHswEvBvBsvubvyUi7pPeUSEFS2K7Z9VvkxZ/7XGTcdMXb2PbL
BPn+kUt9jW3yKpzCotvusd17mCP1aQhvzURca3sVKv5eAI9BhAxg7gBI8FTmP5ZSJtc/WW85RROt
iXPmkjcrD7g0/YOx7zzkLeJHjo92iLDw3pHwnluyPgDGJ9VAv7vnwA4vpWW8XMbT1+2YgHmJ+M4Y
DMzkltDqM6EK3LZRSgvgVASCv1yOLjZ9DWoLZOz6tyJbHQDAw1/q+MBdVlKcOHSegNoI8WGqdYDd
jrGeeyVDBjWJ70OSs+Gz3BKlrK/tRVFrklxbHSnBxSQmJBc26/Nw2OA/DUT/b9L04wxDDu/xDIlS
2grNeDJW1OQpe8NvtEbOVJDgRfadag0Js4J/99YAqNK6WtYOGmCOUr/frmvgGiwLu45p2KZ7UgR+
CF4Fk6JapbIA05mB9OqGUPm4evVJ49x63r6zoeWilNq30vI4NHGPL8DesaQxEZ42+lxadiFVO9JP
5I832kM2ecavbwCiozl7I+l51lxbuKsao7nnVkrtdeMbRd12wDfVTJDXGdDFhpbLOqRL153khQq7
ziupfDFDF0BzR2e1DsZCP0gkj0H5u/zvqBkSCJmzeBgztLjkYtFqGpikCYpRJbSZ2k79RwJdo5e6
A9JgfB25MjWRUtBQ1wmcRZIp6XG5Hzm85Lq3lTzCoqWSrcM7H3mGZitEzMWPxdDitp/9yi5ALjp2
eJU1+i8rO2joE6PvddCr0JRtpFsAqKfUyaqaXeFkyObgNYmWl/4T8es0fEFjfh+ffz2MJY1wGG/i
ZrDlrP/6NEvJG2E1lkD4kM/Ryzx0+DZI4QxwC/X7+jraIKIjSVyFMLc/RW2Ws9qT+YiIclcYyE6Q
Rw3GNdoZ6Hcj4jPh0sGHFl64jFtnjh+z5BRu6LImdo1h49+gh69u6MnPEobQDMHE0O9FoA8UvDSe
IHB/YpAdRfCu0itHIF1aPQocp5Fs0lRlfCrcLsSOwaDwBruHtVXELtlhlTtXZ3qwELV5EjmXZ37J
HjWyDIaxGu4YRNwQTJoWLL6J2WOZVtntJDJthDXwg812W4K5yd5Nww8XXr0jCzP19lm4zgTURKQF
GPRYr+kbNX9bOeFTodbHecDVv6qFeZQosyy3orv1mSH41C4ZhKN0gDFP/Jvp49ClP/z5GoA6G/sE
6chVJUyn9PgUdpO2Csrh43innQkqoX0Loj7djiBKXfHhz4WIc0LdVehfzNdsYLgaR4V8vC0M1QFq
142A6G6h9kR+GdDlh1h2TWSfpaIhc5FLBH7j1Y9bRep2S9CZdzVmlZESzKrFQwhvajUHUkOxqf+i
wpjJUAT4PIjTT8w5aMEYjO/TRbVzDaXMWuPKot0Q2z7ENUbgKIdS5pa4iKkiTBE/R9SGU2e6qQwE
dMp3wnYHlL1X5ivjVl5gOAylaovu3cgP1PRpABuC48a591/MOBw9CXFRbrzoPT7vtiyRW9oGzJjD
0exxE0tXK2NVqi3Pix3xSSramERK1jJdsP9MD57nkhPWh4Gkfpeohx+UG+xIB6hisL2WMBzPeMVs
oEmIQIi3WPxa6pEYyAVAtGymXyTIyFCLVDM4w6GHnXoH3q01FTSkhfVHi2/62fa+gbWK9LaDJMsY
tvTn2iHYGUvNhQvza/JTTV4c0LL+2Jq61lNyqsQM6VCmuutR9qS/EQzma15PLM5DX3+SohMZ3y+u
QTDPV9TiZ2cXwDjtWf4IpZouV2fQbibAwWywkuxZW+aPaPV7bwvv8mp/uT7VBLgn2I1YxGUmrDEO
P9dYdwFugAY1flhK168nvQVRnDxSLbSgSvNi7Y0Rb3Au6xJqt7b7PsTe+n7FIzsYIBvJMAvPtjzL
q0KFPDFljvZ1G9NTSX3iPsOtCpBRinYP8g+rUqyTdIN/stmBprY8oU9kZ17z6d3lA3xuxh1fjAbY
mmaAjIFkP60V258medqV7XY8sokDyC+rk8HkYRnzhWyv/7+/ng3tknCrfjs30MA6NYSVVe/+5q7W
Fcd8VJZrSFuZSTWV4Q82tD35vBv3FQFVwr5u8BQ00sGMWP7IHeCVvKqil7WyVtH07rSchxXdwKqC
r8urSS6zfiY9nxWwKfrQsXYX+fMpmruU3J2by2WxXuwsqGvFZmVIR+i8Gl8FUnS+zBe7gVSSQe6F
0YA/kVQEpC29nuoE9/INHBsFxAlXuxNyRjaQIUCXO+erqw+QMxFUtl/HdCiARQzzJpyP/RoE5i9C
+3gvauB+UgdB02BmJz466sjAhtTtyyXSRVYfx+TPxKNPHm4zWk9rwaTIArbKFQniaM8RMXGIeXv2
RQY+T7EkZ+fHoOq94CHJk8QPXyFAkqXUD+2UOeGdJWp4mCB3xb3u7bx7QGQptTPcQriJnORDabuM
iDistKscibJHRtBJbET5k0wkE2/6kfSSE4/CnUr0mvAs5meS0ZniLctKRB83ppF3k/n5qaUCjnLp
8T/bOVRbSvcAglNya09GTDMoUn2ZPzTFr7uv0gdxZkK63oE2sWuEyHAY7C+t4pbxLnQXwQpLfqMh
ZkixwYzXuqK/x1nyH15uaSR2kQj2yHrZ9v/tG7oJUTOTZ11TML4vIZhwQX4DdS+6N31RH8yRKZEW
AbVRoAX4f1U61FDyf6dN8ozEieSdzFZbzAWcnmUkWRxaSIs4L023QkliXNkaeJjKzDu+Ay1R2J6J
l6ASfyFdY93hlT78G7+lYXlV56cQHU3Et+NVgwvLv9aQxTFv5k6MjRKvbotH2oQj2xrVu5zIw2Vz
DvHWgQaK8kUoQQZR5wMimm9KoS8N5e/+zA1iqTxmAKj6FO1R8vdqAU2lFoQOTNOigSNltgYqyZyg
Asn8TwqRWCN5HnwDQ0kdTX/uVTM0YGbfb7nfmQhd9bj99HnHLCLnu/Y7AgHuMqR+gXhmZc0Yd5wp
rv7TtKICDrbP9de+GNEEj/2JOAgiHcBZLE1qWwP283rZjQftlarWNu9ihS0Pa0l3v+r+mbUTPFtP
N5/ANO6prLUyp6jMjFL/SBdWBOgWs+GsbYHUg7yxroyW7JaG90CXWcW59pSuo4UhvrrQVrXea056
YP8fN5TvFeGQJpURFKNktkA4dEzDVJDGa25Fc/D0WZ20DvJnsriT6OAEzKi4R93S5b+4QAywhbQ4
hpX3g7jEnNGmC4yDKeYwWl88DerboUGwt7olex3sps4fs1yXDVQe16DrNTKayNGrPqRZWg5i+bcD
PXQU09rDUp2alQzYVzpRju9SpN80e75oTdOfenZspwv75V3UhLWQnHc/4fAxb2/0y3PaOxyzrWqu
lwCnqqDG1KmNeadaYfgPQgq0cUyQw819iGhsZ6ckVGZ3R86wKiaPfXG8C4Zi8M39v8hQVxAhXjOp
52V5fBDDsR7sCIVbY/71vAdBil+QnxM2Vh0F837t1MRezGdK0wdcUFxSIYudk7r6UCFagLSDM3ke
DKSxJKJP09f93n9n12rn77ohFNnwFOWJ8GLAw6aWnYiJcNg1oei1xW0gG8vRp4TjlwgnLpLCI4BJ
/txJVmjpJraWcXEJWAhrNDFKQxkQvmJvS7K92e4X405LGNp5kWFoNORoxggceeiLFi/gxvgevh2I
5qM5wfUHKT1j4BuNeBpCmOggR/ypV5PBof3wkY+KY7oIwsWUYJzu9RGdIBTXVMo2ajy6a9VSvfdl
iq9q0eTbkq49qoEsT8mS0AHMtBfy/cOcnqQiGQf//I7le2knY4NB4Ba11dJLmRrxTAN99+dh4kOe
/U2/LsfqzzqdanHI6mFbrok0dMIieeWf1sZfAX2rllvDDCXpCcwRgOdNilFFKlv6RDnjPC6o/gYH
q5SMAxB+R0rvAvJZaNVyfOd/s3KYd65AasSJ0Y+tLxdQjK6gVFu0jrq9avW0iCdFWg4joFFFyi/A
3LqHBZHsF59mLd4M4XAh/nUHh0akz1SEiBQuN3Wntbn9Ts3m7AXnM7CCYNppQ+CI1cPnBdA4rWYg
4RN+tlBNjcM2yBJ03k1a2PWTaFruNamYENV1FPPjCbrQpuuGnd1R1Wmcy9/xzJWao6u/RWp032XF
T4x0K4KCkqow74/gMjRJ0qIcKLOAZxW7zRVf1xVDivvXL3ZbBG2qYPhCT00/GDfFq1PSoyrk1oaa
lR4JkNC9Ykp3zoLYvW4ld9Bb7iD6Dzee6sknn1jLXW8tGopgmYolnqYalqZUW+H1dELGPlQwy1VF
LlhjQ7fpH5uqZVTXsMu5zxI+eiLPaf10aa0qygo+/jWFOjw66AY3BbfVZCGdOirRyDI1dbW4NvkC
SB9REPQLeZnyUdkqc1K+onjyS++jOH5dLFnZFzHPF533dgQOhwy3HF33/6qPhX5nf+f9txtzBUEx
PN7m3GtVuDWqa7zmEXC/KkPkzF/YwugzbaRVtKZHu7E4UvTziyrxwf9UxZjgCodrwOkMy8vPyC0u
Hea1WzyW2wdLwGe3aw+DGSy21IR5wOVxcHlrxDtIU7+gP1LuNFVoDQhcw0rw+YVBsq4CpHoVsW7W
hPXTVXzUYu8i5w0y2Z7bZsai86Rs7nvb2CsKQjSZT8tcWyOaT3McuaYd8/lrLHplkZpo26b0U15b
hANEe3mlUbofw8AICdiCiE0vzbbigEjsOH4GtKX9GBXDxdRMbIZbBxD+mzwxktlto9fyZnFkMgWV
GoQzYk/FB/rGdjCRXRZeBSPalGo6c3t3AgkHhwhqBd7vwOckjaErXdeoQhzWbJuZaXR/V/kvPsXI
hcFMWrbeGUW3LFrefAuBXnsmjjQPPLCYxKL55dWI8os3ArCSZr/SLBAjAAcPfFi95/YtMfHG60k3
p6bNXAO7VzpRuvanNIXEqHTxXm+bLboyR9Ggah8DXyuSpEJFlqF6nwxqMxRyHL+gJt3/1xQHf/2e
GVcReyF3SDAoBm1Zx337AuCydiPHoF3+ZeRBs67tSoApWGGzj92ASZTV29fEegsERrFw/kZOdfbf
+KkQprrYTph70MBOrUP/53RF2JSGNUERVGAowsFy9P5xzrRiiFYAPEyfwhckoh6rX5gmUUH5CmUN
GfSHaoH29vSBNlHl+1+gIpT77mB/kS7HzIzzgX5srdC/e+HDoT1HrIyDtwU8qMiXYmUKIo3GlI+M
cC/HG2JMsLJjyZQ4cOjmVUdNuh084KalNISQTawcXGWqXbZHljm1aH97g/UHadzTWAJkbjCThNaX
pmFw3Pg3p73HTT4tBM4AnvHCHd38ZOp3PuFQ0zmkKa0PHdZ4aVDsmW7HFKx4jVRKDcqEdom5NmtZ
2iXY7FA7Z2fFkXyWzhveHWL9RFYcTa96Q7mS7HAo4FetyImGQ92azSMYD3xo2KgqkhxifwCuxhwP
Gw6wHc8TgxD2lXHTMkppndozys6m9YemNk14o/jxdNanWiTDx0wXT/ALSbwQ5gLDsZ7a7L8DFdqd
tBZK+bz8QI4LPIEPBCRa+Uc7+A/MF9v3YXsKHGcIli/Mcd8RTr9mLPKfdXY1gB8E/bGD/MuR369n
/o6RAtb2/OcwyF976cz0+FUb4ztC8ui1l9uLiT+idsuXT52rRf1IhFOW4UNVzNTo34u/36whr1qV
5WfaqQNeSoGNtLn5oWBNuJRDDRjpnFfScXBa8XGyFdQjTjAfrbKKLjLArXFg47474DeUevpLtYlR
0IuZfYxBc4+67aAP8YkpCuvmq3u6QOOvT9z6j401Yb6Jdaoml+hEnVyU6ue2q882OblFop/GAhYJ
vz8dJEpwekNL0g6uog7y8K7TBQwd0Wbw39N3+m9fpfIM4xZCuZ7VBDB0p985GT0SrgU2ZeZ3DybF
dE3CHezXW6AKzKb926JaH3V18WMspk9Jz8A+GEhrumrT98nCErJ3bH1D5VdUXf+hIS6gdYgquEXY
Xf9y6q7dOlJFzKZf8+rJJgEbd7aWsumu0sXnbBQ3Dhvx+BrOhPpeSjka5/fb57aMtN1XUQTlzIXz
yphzEarLbK+4MfsPDueuk61g0bh/i0KNHxd3nlNUZ6sfvxH9+HjMrWpHD+/vkfwj5wSqksdHVc4Y
Pm97Aurld2yGyMNc0oeeGh+Ig1P7QT+OcHDHoDXNLpjBCsFiNyqIjDr6R1aV+2oOy9X5klrlHXsF
qk6XJ+/zED0s5pTv0i2OBJHdRKYf3jpiblGl65Glyk54LfKMduAoWJ+L/NVFRDKoYcA0Obn8zt/s
eBBq4yN95s8cRNnM3fTWj4vn3Xno77fYT8WqFq/SRmQrmZvVXJTdV2pGoVk4gTcfjAvZL04BPB8M
b2RBv6wtbmmunCUlFxqd3vXt6GzhBKPey0fyk4wOKFHQEdaHqhQJNg198A0MkRSR65fzYWLv10vz
j9syBI8CyitONkEXqSZv1YtmtUszui5NQLBVvoFFv+fEg6nBc+CVCEYaHTiF77LdcWu68vMRh3t4
56QikVmE0ivc/dXM/75dSoBR0RTTVcrQhMcAg0/LBct0LUZJaZkpsdfiB4d3595G9+yOi7UMnGm0
ojdlR4PiNtIVOgSqG1Bep7eoGQsRokdyxbj9XYRgZpS9oP9TpyjJmubc5Px6jURbVrHOFjcwjprF
XR7rk1w0QD1ITXXowDUBIYWYngK4xe+LVr27nCslYjQJWhjluOE/HqnOn0+uYs11a3kIL/tMWM8S
DL4mOWGUzCQNWi2BzV7nqdRdhSNtvHVQyffbYcrHA7fZ90QOXH02tclljf0GsPV7+TJBVoI9xR8h
sLxCTU0gyMfx0pzyT51e/b/GqQsr/7pt669CqqMd8+ZVGYxhw5C5YjgDKsqc3WBdW6EhL+mZy4hQ
S+W4RhhejIWgOF4X3nHjiSTBECCjKQuBtL89AWOYScRf1JxI1VG8m8u7IksQXFUNmySRk722Fnfp
RAkuc6+M/IutdxvjiVyQhr7XKhmfz1EHg0eS+uqIeb6JN4cR3AQDdB9U7wq2mg2ztHdC5UtDUYdF
sSyyyB6VL4e0Z7NMwgshJ+K/1w/syFYXN/DcntJcQcAh21DAhJNozzyXbCIfvCGmOCp6O2gri1P+
VjDQDqhRICcsA/BWwioHz6iCMuz3JRq9HLp8ZEcUuWa5p4uWtB/a5CW+ZUF5e+ka89d26aUdPxff
kghHPE0ffe/5f/PzKMCG1U4XONrFlLmLxN5iIXQTF+YIGhWgwbPuJC6EC/pz70dCURqzw2rOKEs2
1WPOo6k7/4mi2dHo4v2UZeHyTLXWcy5DXv7iITEFl/9RnmmoWg/PU9LfOB1uVp7UNQoIv8CJQR+L
bwS3JuYaqSfCyjhVfjHqV9ccD98/UwBq/bKhv5Pa3mqAP+AMqFWrw8JYIreVTHs/rPeqIiQmUEqR
li4ymYplhtuq+kFXeAMo31FrwY0uSRvTZ6uterGAEX206UNYx13x5h+1pcUh3e4tkTt2ss5MgGQA
3Z6NxqA+0jv/RdzA4kcnzcwcGbWozZY3Nv+hqDubmr218x22AiVYyk9ogQlaPGPrrcW3yKR00Wbx
J9Oqw7fHrXuBynaUyDZVwjj0pxOCdr6HPt4AdEzO0k1DMeYZuQTBbT3hz5gYihKaECEt2nHpsoLp
XVeGYufn8wwIKtOJokUtSob+P98LFvHTc37dDAIwkO+yvqP7lk+cj/gBw2SrF8ySBR/orl0ldMyV
YuBYh/qvWFp7QjAUOZ6VFd32C/cy4EN+R1E+9wu/4mkUSg2iLoeVW7YjEGjD6Anpka1oZGvL4eKL
wn1JoU8mtBw+WHMmyia/bfDX4iwzTjCwW06PsuBRixwit3mxuNffgPqCsjG+xHL6/p0zOGYSVBny
muMX0eZh6MT0P65iCdGHsndzfi6Mp0uUzyTmyBdTrY/8CkR9fVt51MIamMsWnlff2f/s/v0CwB+Q
10Gh4Te3pfH+uRTsO8Z13+qWasbIWxUvLMdDEpfVXPMOBrvzAXvV+tcswYZm8Jz/jTlZGM6XS0Bz
7YylMNsgqYxQPq960jPi5PbZ6o/c4n49OyBO4raQmNE0fYpSL6aDn34Cn+2k0uepFVildN3j2ZBS
bt4pScMGYk38GAi0Vj7UeHpr2ujLVYHh7Qm1JVI8NK9D1eupPoIkwIOv6ejPK2d2yHSwWeixV3ci
b/9Jo+LonjbF6xTpMcbfYeJbAq3Q+9FK2RBDoXK5S8sorsDmbKfisbpGi6cc/iy/2SC6sdyty8te
ww94cP/RI5ed61CHrbElFwKj5DshJsjagUTEg5JEzoaVoyDv6CtsNkFZEC47e8R3+A4zkDpyyW+7
U4HBrQ4xTJIPe1seqLMScuJGx7gRO6VYlS4DiMremOX2Hh6jbucGkmN23D9rH40YbPRP0LTKQd+w
TTmnNYRjCo7zkC4niVTsyvGr4uIU/+TorsBm/NOiIqSSrDO+9ZfSFObdlu0rXq9q83UAQs3rVHuY
dPElCeyKVdGQnM6Rl1OthL2qhgv65z/1UVEXQ3GkrJuRhAJiC0k32B3IiPUZVMsxnBEpRNgJfW1s
MXt+8feoue8N7PM9Y3IWdkeSwOBuIbGMEM4xpp5NvW+7O7J8w7ot3zrAWbZibPNtCbiPza5RfCM7
VnXqLH0VQbHvdg5iFHmx2V6gQ8DrwUETnILRHsGgHaE6spTow5GkILIWWTW9TgjxnXk7vLYIBwi3
Bbr4uV1vA7xQrvhjch2Q4fvbwUhDcY0RhZGn2tBXGPvbJ2IprB4GlLTUDppDwKuxQfcpZhF4uohd
Vsyu568nLaCQgs4BcFt0TaeOvy/BHaZOKCm1RkKpjr8onqo/dE8FhQSn+V8yWpzxK38aIPx0CvAq
Oata1eGIAy6Smclnd6IBB4M1JDherSOqw3OSB0SpP/m2PBhq/er/TRHzSSzz0jXz+nNxoUE7CBGZ
IS8jRhTEHES2htMZNu+EcqM1JnQTQA7eBmrW+VrowehAs3ybzX0IrdiOLNiwjrTE8cEUewnH75Q8
iFHxXcsnjh9hGi2v1Rw+j1oXKb7V/axKuRNo6X6jXyxf2HTzLVIP1/j01Am/LK/Nez+lnA1+l8BA
Ln5BTbdSPCHHOz8MVzFzaYmiopBiguEmRioyR4l9F7P7c0mCGqk9+gaetq+PUuauYL3UPCrLA/po
YEtWjun0WgLSjoXN8pxA6AYQ8nkw1/j8v4TMaSELqpmnNB8CaQSBg7X/kJhkfqfeC9rjMwmeZD3G
pTW0ML11/cPakr65z3vqnMprWlk/HBtXbvC1eVbV7Whdr37LKbtqBLo5sVwvy/+ESWd3PndE0u9/
jaXVSfuVJ1Rmz7fPuJnFTgBeM4LxgwX/eTTE5apf3B2gUFePPvppxKyfE3j7YNikY8/vSRbFUNqR
jPC9H/74KtTv9tElk1y2l0380pv2tCPvAWgny4EqQV0XbXt0+Jppb9W5bPEwZD6bZ7xA836SYVW/
1PkoGzniBXd4ObeZuxLn8uCBLz2uqct7ddcGiIFrCBWgdt/bNfDhO7stg/OdbEZW4ws7GrR03QyR
nlcxrRoeF9+zr36wHxfziCg4RAYOiDAXyebXmExggp+Wbt29FDQYcIjb29yjWV8M999hUL6T2/Yv
cpa0Ryu1lA85KjAFbh/mauNpIRbVzaG8JARPeywyZ3sxHtJWGqXSIhMQuHsngzedlJb9R3I/AzvJ
Vp79w/PuUHv/6OrECASSsunzAG4STYS/kSnoqwuOSXgWOqGSG/BEcgZz2f1GyClj47aMN4lpExAH
6Tt3kHMET1HCmmjK2U5yYdvxIIDRS3yQgV0D+tQVOS3G0J2EJQaHI2Dtig1QjiaZvFx+4c7bZ+lx
rs2LRf/iFp7ZYr5eUvVfPkx4sq9Vd/jSm3vidi9q12lKuzb0bUzpCeLwkcL8TDUa94gePFRP3PDI
UvT1UQZDWFGd8slJQ3Ub+O68gmpjDVB6mwKgt4VZfV7ehFC6oEIBPDUctcpD2REWUCwPgHgvhkXI
HRAzgPgotyYrBMdifuZpJodpAL0s2CHxzxeS4xwKT4CG8AMedicN6443uJ57xSpAMDVe879EUfmI
F3B3Bn51169/f19TVYex8FyK/OVA0OyMvOQ13afy8Yo0JfUGCERhmnmvr0FKocqu9B+3ZMoTSz3h
tGha03hNyTeZQW7vG+P39APi2P5fX4NfRxWP003QrZ4VMMuS7GaxPkBIncLQKPdlggrMRFOvgZbw
P3MeuG6/AbJ1bYi7TyG1u3Nr9fN4IPa6fpMWQrswcmXfVzJomOkHrf4FW/ec80yop+IpA1m0yR5M
179ztEb8gBdWtfOzgoT4AY7OUjOjg16FwwWwtDr/fCJI1ouyCi+MyIfF7/LOEJ9xkgmqCUbT2Q4L
E+5qxnKlS5PBX/QofR/VyfficeUvsfcsmjEOO9Aayb6PmtJMKiSbIKahnJocaO0LDdStsHWlSHa9
b5VGNThCbHj2tjGOWd4+SfBdMnbLsqhD4FxbI6R8UwFH63GECDekGl/qqN0QF6TOcZHkQf/28Zxc
w9QTjlm/TUn7xnAKKBMIxskqhLpeef7OJUMLCXKfeyFA6tf0iZcy7k7wT+Xmi+v9iU8EfgjnWjDR
3HTDLyPxe+IMOpjOu3siwu1/h97ZimlfH93zrwk8No5sUFRBiXQgk5cML5skSxxleAolQ3x+YARm
2pXMHIzArJpAVPLMKjXACZVKZrlJuqOqYjzBy18cn8h8vE17fnE0mhBr9ahYBIgIiC69Wv//W3UL
PYrsAR9LqCwKflr9D15WRIvJ46QmWkteMVe9/53o/ssh648pQUXmq2l5AvHUS0gR2W93E0P30mwr
qhhF/dn8fCn0d1a5Rq3+iqehYD7c79XTnx0xazeZYMKmR5SrAxSqwfnha/SyZ1WTf/RS9Ob0LL0h
LKtmQ2RPvfYwzyRns6SBsi8cNOjE4pMniI+jm+C0OUNjBGJIHM7VhF+Yy2cq5Mby6gze4ZFSOfGb
gYtYURn9gTQClsF0mj1Rz+wevSw24f2CE1P2F/5KzZBB4VsKZUmF3Umi9HeufpTJ0mMNhmE6z5ld
b2nPRiRIh25uXEj7EgnkcC7EsWwYTR6D6QzcMm150FZZfKOrqmpPpnjRtE58zVVWkLeaQdDhk9kO
VJPByup6pvZozpgHddrGJm3Fo+19+OG3pOLWBIk6yRnp96m81VnMf1nIxzZMBaN6iFRcXYqvibDd
Q2nkGbm2/rvVTuehhtN71R/yZMwZtA7sjmihNmzk0wHGtqVkz4eSK1Nw337ckzHeXw8bNIXzA/85
O5fYm6r79xJHPM5zJsvCiw26onbC4AXb/e0HmhuVJxKsX+ZsJI9qVZitMpfw6nO4PmdTU8H6t0C8
S5UhUVZL7TGOkb5yxDqlTioWp4gRo/JV7xoLPgnCwcRA8HRdjRoH63SDy21iAcalyk38+STMDqJg
o9/uEIoWPefx/4lB/VzKoduF+DjiLmpv+AId4UIBDiWbMv5Qwz+CXQWEIc10swZNiL1CY1t9YaHp
CSY3k7fEwJpU9x1CkPPeheWw9B+ZYjAEtKQSW7jSs6U5F6EVZBNz0AC0JHlugZrJVxJ6PDN+XMTr
2POqDJ5Q/sYXA7fW0KeqoHVsUkyg142Kk3xhWV2DzmxoRqfLy9NI4ykOnm0NtydkrKdNXL505/a6
MfdLtM79w1p+Ar90h4m7MPmJ//D0PAyhDiOAo0147pMPqT9GVYXyaPL6sXEYwreQnu9gdAgjWCv3
lRZepYkRwiDQox7uwoof0ss6JK1+E3O7CvP2Sr9lgwtYPyxHq7GO/ppmWPZYYyzlNP/v4Szx16NV
D2P04wrFyb/FU+pbkJfjikL9BVoQCTloLFEcRHtEnea1SURIHcIf/fdK+cM3DWTxK+hMsfD2E1zt
Ad7V8xxOCOlgXJ6llfjCMazxk9UIlYtNYj3ZD2eMPcUtfn+b3rVZ+UuGeQ/Q9qNtGlG25aH2QRD4
AwEVgx0WqL9HqtmG1vfwcLCHuKTsixY0aq8dAf6f3oS6XR7LF0Y48ea80UsBI2cLLRgfcXGn3mpP
2kA/SsMq7Nhrfzn+GErM6+99FaAWoK0SbMvwgSd2kLLfb/NdAN/32JGhdp4vpL2LwQ1L3PUfPTQr
kyYwyQy8RH9BlBAAPbpXHirCNOtDX2LbIVYWwaTUVvlXQrncDqFlHgmZItcebd5EPJWaYFeUXb8p
vtPdgnvKRrrcOGwkFTE36ZqYbiEjCGHvI8NAv9iybbtxqRY6rCiS1boUkq3eafmyT3FmzofDSxE4
kHvu4kczdmx+NgFbHNghp47c+U5GP/+/bF0qN3Ip64gevjQJpdOg3Fjx3F+2KP5+HfHE3UPEUL6l
0ZQqBKqAh2aMgrR3yqeE/tRBErNLKlEPL+0VERAUXoD+3tjm7XmgLszDLwrzBOAKU3wKAPmCdgqf
wCCDX3Xi/hZ0EGeJRDiBfl41MzvnRmVJ3tAk3QZ8ZYtAzAmxj1wMSQNzWXMDBadIX+HGa0/2Rfqi
dUbam+G4vBMzk+URYctb0NXC4NIB4bdnULfph2iLuKq810nc1HstlGUfOCK+DR1RfETp2d6eymHp
46ziK9a3BbmujuT7Ut8VlwIoeSKGAddiXWG9MFpBirumpA/W3Q2Cpq9hpCpWH/Boc1gDfD8S16IP
95lI+fq+wBCQMGIMBrfr+6rE5Wr6jLlQNgk6u7XKqPncey3GWBeHigl0MnIPsjTlcVeu794BNEUO
3I0B+aBosNKxTqDky19IcNiwvG4eeo7bY2Hz5amEmi4QUqWsKhffPRq0sDEo0XVNsiUOYoko9n8F
UEsI3va7BHwsDOiiqXm9X90ppgOus7Tab1sYTu1HF66ndJd6sQlS4MlJoRW65HypXNS6aIOr6L+w
kLqD3zPH9rwFCwmzjNUKH2MS/MB66ob4VvMK6Tkwfs3BvAMxh2e0EW/LNlT/xS4fgAQMcBJQsvFk
m6U2Te5ZWzj3fyirFIZV7DPjvp/bM0ddonFDvqH/+6/IhSiZrIlohqEM4ipSjtKYnKp6DgMajNdw
NkLBGPDT3aIYC7ufb07uJ/EOMfyhV/HaoJP95633KuQvUKwdx1KDPqwO7mDdiN/o8Xu4WEjh0H33
BFL1UQzF8+9zK3IKRXAKimhBibBM4BXg1idfs6O0obhVJBKcHZPcmDjb/3hNyP25XJ27fuIiR9gX
1p71LLCOaYVHw2uUvdF89iB0N+OQPgB8JmiEQGKocFkjQsnmQoC+IrBRP50jzn/7mORSz/+AMmNa
aoLNezaeSMPGmU2JqzvpnOqkO3s8MVAlKMepR2q17WDsf2Zrxh6PWpYlLnr+JbmwkXWYIv8eNCAN
vcIrJTGPnhfjoR6MA2B+sU2aFImg/A1qabBfBNBiW1mMJyYu9QLGGpQ0x77H//SQkdaf+xjpWVSi
a1JqLAdlyBXBnk+IQ8SoMn3nhD9Y8e+CMo7jEIkHRC1gIi/25QlRtYQT/soehKHAeADgdhm876se
Ow1TgQ5vq0GS1rsqsIh43h6r2w1MwyRMy33//2T3rBg5Xfabxqc5IQXBRjGGsFSaSMimIa5BdTa4
ukpMUuXoGxUZN+OTSbmBRQr6TpkAhm/4dxXHwZkfc980hGwNUuk8qXKYrsxYN4Tr2YC5oZh6atKz
auJfb7lL8OxxDt9QhucbBDaZl5ZUuXESPaDFI/8F+D/QZ/EORZpor3G8T9EethUwah2XkYwn6GYG
8VXq03P92eqSR/gJ3cYXCtca0PFPckqlqQEyOBCqNgKdDAhTPprunBBx8c6QgoVIpWzBFFsRKWyU
V6VK0Zy3OR5NyjnH0H3zpf8FcdGFC1InglGyNaYYsOxugOnatZKcucsAxZUj9xjV3nI458jvfxwj
xXftC8p9hHoyV3y/MhSbGyAQXiw5Loyo85+zMh3CQNG/n5LDX2U3ghF1WqaMUppXABjPeeZbErK7
aNy13vaq/AQ46pxZPib72ygGfGBc1rrknzJNrC21d553HDRnZz2ffQyDeB7S/nd+0iOLf09/cxmM
MOveE9S8KXTS8toFLS4FHKihHwFvyhqqmRi4PTuJzQb/ZTyezi56BZs2u5BFWGDdOQDz+MD6TNIV
1nQvjwx08mKibuGR7tCDOkq9GPS4Nw8sXHk+kGnN0dHRREvaNhrn0Ni2ZpjUJoV203es1UJvIF3z
3zbdYhjtsIlvIivZ06LsD6ML6TDyM2DRlM8rMIw4sUPHl/eBm/Xa5khAy1mU6jCGgZEJrtTdRdTt
/3MY3KScpaQxSvlQIfn98EFjy8prWMQNj0FIN4VN89ZaDLeH2onThHCycEoMtYwWVWkUlFXmSk/W
UXbf80kAt/1X/9745JVOPJzIKxF8RPEG1xvG0fhT2kFFUlRssm5BZBQ0oIhVubA52dvxczn+pyXL
9U1225meZgBNG8dGbQ4Oe3NCBzEjTOq7eIDeVSxhjbjbrFpQ3Pw9psSMbDBZ/AfeNM5Xq7FHmuH6
C3YiIHkahvztjNe3h91mzqD5bQzt2AMIPBulg8HFkvppgjEgHaM3gJmO3eegpXjsaL4HIvAUFO1V
MZSomHlWOBuOg13Ld3tB6svypizxBWzRuhtAm/MysCXJ+rTs0zliAJ7CwuupzG1ygZVXzQUB2GWJ
LznAEmkPxJoP9tasZkCu5FrHNFujCvkduXJQMWN4hv07mI2EvkLODsDVnP69ClMdYXPaepx9kOdw
NC6ei3jkcA6yoNlLrB4neYeoY40ILSh9m14R0YjHoKQotd4GZoC5zTUTl9n4PLlAtkrKYeZysD8Y
d1we2PC29XgO42dRHPqmVYDv+cIqh8Mc5A4XRUnzwGNnE9kP3jtkNnOMyJrSYEg9DNmmrvd4+bSD
lC1r7Iv+mLVkijV96LxIjlnMFGwzqUMnAU07qKp9/pJpuwx7IKEKbyMfjFHYPv3tLv0PaEBTxljP
wOzk2nk2jWQmJmxLBd9EwpFvM82/XBsQ6oOF0YLJwjT9Ljvy4BSnsYebHm8ByYae792MKAEjUE3w
mEiokAq9ERwTtECTwayfZ+cR33E94zK7OpDA21Jjy0pxyMbyz6jaGlhF7bswjOMXTp6jC2dTjnrY
6m6j6JebeNWmp9p0d1Pp+DRXqMdqkXGLZBLn9oahIQ/gXrNBE+NxTzQX3O63pE1fWqgFoLdWyuWU
zQ8Ts/Y+pBGmn9prM0g7yl1chhIDNlwmPpP02q02mc9DavdJ0ZYfO6ZMfZazk5LgkgrGQGaCxLpp
7MkuSsh4advCbrx1sBhzY18K+v0PjsDakzYbGgBgi6tHA83VHF+gaUHLRbbpvxrhdPuBl06c10o/
TZOAIY+uWO2zxE5vEaa1sTxVkklgVUgs0Wlv6sZrJRvaDCPJtIzh3T3S6hlVknltx8rdyFBJmRdx
FrSPTS9SGTTE/0EZI/UtyHdkXDDgJRKwBzj/uCEP76NeOvdHAjflFuJmyYd3jKvV327Cviaa8vZy
d79/5lGG/a6HjjF1H1kvw2rQYgEx/S2a6UfIOvJw3dOhO+xBKB+q70CZBKmH1z1yLCzUnc6wZ3Oc
MC44u/Lnth2SQpxsZ6P5COyeFwe9fNTMs6F9DVannvjRqDTKtRKq5yTKFnkNwEW5riBg+xXw5NHp
Q4TX1TOtgja5pLiiUhdyzaQgVO7FizcWot+7Ly/m7GwHNB44iEtCX7eQOqzV+7TkjfLff+FvE4JI
OMH4g4J1nut8HDG+E7wHNh24oH6jiYAo//C0HemFh5I2vWIhljlqyon/avud0UwgxEtymIc/UZ24
FqsKegyKprbIh7bu9pHkEqyu82aW439KdvFP1Qug2l1PS4U5GBkCyOy1B/dx+9oGsvl1srq9XTIa
04QsEprqo+qlLkxA8vc86DewffuVul14NQu0wcqIRoD2KZpd0WAtijHx9Uek+uKsnZbdmxBzO7tY
kFtgpJdtfjJYsRSiGny1FX2IUps1VtYFbSk7Mz7WsWxBdbOQDyH4Lfxl6Az2UuFaIIw336PxC5b0
ZHfxqJAEi15xvGYeQUXJGfeA4jFVYwQOJGjzHUkrzTiOmZwQJDR4O8XiuOTfEQj7VsbSmXX2qzki
zvhrhRrPBS1kKLZXNReRA7G6HYYkRiLJoEu23g7WLVwBZLTnTlhArDsV6rH39A/siNiumfmK4RaG
jWL2oFFnpNmCUssy5RJCVOeb/HF3oEZIJYUNaO41qTz7m0bsqvS90QnrTCjJMjAk+ND56pgqsKLc
vwojW6O+mswR/C7SMlGTYxupiKs1YYSKjhvbrcl7Txa3rKKR5/9/TK6UlGyttbuNTiRhkMf/R4ku
9HJOgihBX++tkVyv6mFmznIObuS9whgMzCtbh+WR46rTFAaSymBJDApAmSYyPDTNxZEE6jOoMCOS
yCwse2f9TPHIozq3evdNkXc6UJcIlO2ImKCP/adACDefjwJoHEZyynvSroS53BMqY/ftEXpMBrCL
Ru65EXjQLko7Ryb5hCTT3X8vV/90o2/tpqdlnNGkX+HgUGTZtd4XaL0ifgNHWsh8bPX6S5EWnWX+
9GLo+OGx2xw6HFHRaKtECDUoJLebkvCrVY9a4iXQ4FHrFvWzdpJ8aRdQ7pR1UBnaqCIGzrCweuDs
KWS99jzd4yq8xY3lY+47EXqQQc6zbjhAuIEapu6yok8C28j1KdPT36QLGshmRxYg/4/vx8o+r41q
M1NI4Ix9NDcrhAOtaL2lF0IQp6FS2BjFscczOmhfOTf0r0LE8AcNozauITKc+IU5Bw5cXmT217ld
MlXvCBwAHdqqkfHM8+CnhoAqVdvsvyzMIa5rvmbXioayHOMUFxp/ZoRAMsYC3AzI7So/UMw78Q8x
Z+KyXoCbNPMAoUTlzrkGw1iHWu8P2GQV0TW5yvoO3Rdp/8R5tqgFhTzMAs6VesqCaLpGRgRyXgOu
4GZ0EFPzCPVlIiXakQwJ2q8QNYtrdy31dHBbyYFWSWNIm6rXhNMteGgkc7VMS2TT8AsbAHgASICT
27feKewjQYArgwWGiDBFBWbF0jzW27+NtqFzoFXu53CiSwxwQzT9Xgrlqt02kvwrsOCGD9ENUXcw
FBgVUxo5ObzfpHQdRcyGLX5X1mdvuo/9Ml0Y3vZnI4qLTspAQPzxecNc8nl95F/TqaNa3GP2Rtl2
zWWCaeKCQdVyLaoUGB0kbDAmK6brMXMePuP1FTTgSF5/6Dh9Bc762RwNtE6QhmEGcPHQAxzqWjEi
bIylx0DjO+rA9OaehuZ5rOIxMl18C1KYpwbo2bkouyuOh+q7OR/L0BMgZQJBanrT5UOWBv0NOuvb
I9YB/WkiliLQsm/C0lpIbnLczaa0uw+iSMsdMewXbf4DkbkXI/TlaUbo3k945/OjVdkJjKXUUzK/
lSSqJKk/bejE0ashjRLIzJ4eWqZLkKo7ZYXeMelworyjl0GQDqwZ+kusugVv+tOquFPU2wlWBobG
DHSLE0vniYVoJsZQvUWm6mggYAQ3Jgc5cZUdvuP5HzQZF7DTYwHAXvte9P1FgtCJK6/DVH1SIgrt
TVCpNIoAT4oJpyeEPCD3+WVDZyTZF4vT/K18hElTGiGv/wGCWQU4U4kbk/sfbpeOW9b1Gt15dJm2
5iM6RGiPCCrF7p3kDuw9/M0OjvI+zdBn5BFrqm4ZYlQU9WeBGuXGdX1zU4dX79rSWdA53sNztZSJ
S/ZzmvvRBchfKfAzF/xogym0Tpj2MFNonIBGn5ZXFCmfKpAP+e1NalLBCGJSrArmdmG9PO1qTMoG
T08AIudiW14pp9+F3u1x7//SdSWznfo56nCIEExvggNIoDH4hbZo2nCUWde1I1C3MzCjEM7+NyQd
zZ2X0cndpymrylARyYGcaM7uFX0OvLYJky0PTKttcm0bSC8gKMUZYX9DaAI0AwmTOZaZ/+eSQVZE
06+QKIVdtsPcnCjZSYPO+8OM1QGku7DJ31pe8jzwvshMP9gHVu687Lz8i8tyWK5BGxWhjrqNc1Wa
ZK/DnWZu9m/xzUQwcpWcVp3S+15nqhABl2a4aFlZIqtba7EGE9nBsz3mhgfgQ2DWql4/jgv8zEKs
bKz9szUDO/LhWEI3dtR8sLtqa5244ziIG2b/zzsRH5vKRVZImCo9JEQcRdUErpArekW41hX43LLj
QagoLBxM88ytQxzcd7uIIsIXLVHZdNZ+bhFRaYNxq6iFGY5oKAJlTlsjhPyBQQPYD8tIxs3RW85H
K7FRaqpiMlZ3S/TSqFbiRzRFhoyusOyHfQdXk4qlZXyALoWNurwCUH8UEZsK+/MJhZMwXo44dmV7
8rcmFhsKFNV+/4mVE4JBWLHZsfK1L9f4wkPWUUSoK/OzC64/CQgdHKW4ggEnR2+s5RoF4oWMqAUg
ygrzBzMFVt2m3vEthAdLEiQq5z2EyDgtDFV8SENOSihS5QBUWkZ4DY2jtbJnGglvIhfBo2BaCwwM
Wc/syCnyNPbfrhpyh2chWQZ9P7iaED5cS9XqflOSQaMRNAL04WRJUslAryxMCXpyo6BiO7zIlAbX
9fytHonlB4gKuNt7PyhUee/P1gh6sC7kFaH5nHj3pMSZzwYAJn8rItsukUDgiFzj1rTiFjYhTtSy
Tf+yYPDaAU8zK3f10wgF/nIEeJoVvxrifCQ3uovUo+BJirdSXbEWTBXtIG7FaTLNu+/SoYfcdBFJ
PHTVeduYsc0JZX4RJXXz0H6v+foLrbObotB2zeXWbUrgErY4AHcabiW8OT9ZWtz5b6X2h5+tf5aj
qANZO6mynKRbOM4fh8k7hJJ7UiYNCGPia+tRbp+KiEusbfhRWFo0zG5sDveOCOIXiqeyx7IQeqoP
/KWLdMDg/1Hk+O0AUcI0CtjDeO6eiSjxLEItu0y5tJpS5lbQqab+Nty0BJdT1S0efehvx/eG+/Lz
3C80BknwoeW3BTMeWBMpHi6wVnOYmttYAaTAf7IGjTrcFc5o2+vUOrhdrQ+yRLWcPPlFyeYgYrsv
bWpeE/9WHqgOXoEvtEdq+Kvb6pdcgOjttvMnFDv1Yb+pAfBwzdonCCt+PsLwjGgnQwbQGPLky+QW
G4Ki9ggW9n/YUhhS3H46LXBGgtjWm1Dp/Z4sG8nLTHxVzx0/yc2jM5IPin8deRcWNxSl/JK9aklV
tr4stBeU9vc8TF6QiQmM3io88EExqBekjhMxjAddZ4z2lW6PFBQ742/bqk1ORKAySrNDCu0aKMuf
sAkADoF86iROQ1mNrLcPxsQhfrDW3ph+fbuNq6NDw+jQCUg4xFoUobtdOW498w5imRQsslitvblJ
HR06PFV36npbbl6oMGH3WnXC4nWSprcnGnUJNzh71ALhtZLMi3TGAgyMSQ0QkCIZ3PU061k8vBxc
WlAdmbwUU7yinYzPYjxlIsM7jkuP4Pd8h2+RUuak6pnwaxAhw8J34momv4s7Y0hk1VNJsn8Av5RT
ZDTFdJuIsPPW/HceHoH49MFtL6x/IqIRHXkmRJtFzsiKpeiwo8RAA2+QPNwmyngBP94rYPwxSGt4
0Krw+JJpmJ3Tw5hah9gKP1khp90rT/MOAEpw6Q9ICae02vqTlY+S/iztgjrSva9wRFAAfHK/2Urs
jCms9ADSCFB1DCppkMV7VwdqkhdDbN+mYYhK6v4VW4NsIcRGYWFNE+iP+zdBT5caSk0Kdutb5a+G
CvPb0fxfOEEDy03FgaMydUM0R4DnLpCPNnPwvrtbcE2Gq0rucfeqn97Yv4DYTQuwdrAvwril20KR
7/VfV8WMS1BvokLwbvpqu/lPb929PO4Mu858jVV7s6W8TvOqu4N+9ytV/aMhaGidB3Aw4hJTAAwM
1ppxeHPZYnKGXP431rvuv6OZvrX5kjrCD85pllwtaziK3iGUJ8/V1I05nyOp01Ho4xZ20sPyLH8q
UHfHSa78UmWJ/aADztFsUwQri0WxwL6zbUnK3RwYas+8IiPYwWkSQoZ88mgcruJ+O692xB5PFuHe
OJWNoaBgW5+ANL4xHBMshrcI/LNU+g97C0o0eC4WZTep4gXy2XxoEusWH6qAdrVvdelEbdLVJQ6t
jWZvmqklw7jZqQzm9SJnEbqw7CY+pxLwygtH4xQDzG5OOiEGQhXjLvX2H10Y5n8J+aGCsa48Qe2J
7ty7Be1UlnANhbfWaOV7jXfJ+iuv2Fh9am5VT2e5TquR1bqs7f3EenXtDvMLWu4jILQXGUqEjj25
+d31766keyrug37ryPKZigJn+S6XhIwmlm5YMSZBJRCPKQZtHe3Pyoia9OFU+L5THoA5JG9VTgLd
8b2nixdDnDLcWvzSEmeJ8fg5Vp9QN3FZuzoC/txAwQwDvOgyS+f5o52XOHfipUT8TdsqT1Y/SYYI
k0ku90kGU+Wx002YaEXUlmFRZCtG/dr4/LqCKWTJ0/aW5hloN8N15Ev4QdRW2N04RT17Q9xJWO2M
9CXk3cmNZvN5YIVXbI7Vp7loFW0hsQx0/8BIdHWuFR81ee1hSt4qYhK8aEKPIIHG8rLRDuCCp/P/
TO/WYzqP6nsfZ8w3GKszGOdSOf2surFTmS+wxYjtjSusHabXcXGIUCB5EZ+I1Stka2exQUOWoq3f
iMZ2eL1PdxNiUpeGWFUv8y04cHl+NMJZZIG4Ra2AFxHFPRW/m26Rqi89ZcQT+0VZpOsOYZhjgF29
cKiYBC5NDhDdXB5umAl48Xzr2UXibLopV3Fa1j3gAXPXbo5iJiufItRt9WfD+L4A9IoxbG/hfIMK
6TCB2QRi5DgatvefScf6BK8e2iHOZEaG42IAL/n+tDM4RrtdxqgAxVibBOXZCMHYkuNZeoQ8kYgH
a5gyOXny5wTnH3Y2fiTuLVPgPICpkE2tOlDl3fACh9v0ijGugckgtzgADpTDr1qFo4QV6thZloHZ
TzysIuo/icubHRK2UYUPVvX/wefJByENpv429O4CXL/8aouoUywzrYEWKTrTZma5Elt8xY6aeUuH
zcjiy87Iaix+1D3sgc/V7bw84k0vweXX+Au3K/g1Buawm3kgBXxZMCrCk5dpS2imnDgN4m3b8Nqh
nK2QXE+QvYnbbscHTKRBOhhstOY9ucacDxHURrSBkPvR7GzziHjdKo0KP2ej6by6/ld1x3NXuPTC
HXQm5Ai5zCjKBurpf+MZOIwNHQa6h/9RSz1m+COpNOOckNxvhrfAWXvbQySb5ACZkGFhBeQ7yUjj
QPE6obUz1428NcLqWvooeBfYsCFuhA9O3ajYSfZ2nu76ZDOjJz790tvAIAKDcntDf+563HT2bX+7
65vmkvt2XH/S+i9xL7vZozf+ttjpwFKVV3q3xm9iieZjqTjR4RydoHH9f6y4pol9BrE8N3q009ll
4V7X2cQAblf3WogjbUnNVk5cMPlUWZl2jzCLRVtneyISVV+zSV6AHN0sAGiPjtTJejgtbAPIXnyS
tJAdMhefxTUPZFwh0G6QJ4QjRMUsMVb6mSfw3iyJT4djy5RIPbKuFeN1CrkoxWcLGjj7eRuZ2XCm
DYaMDUx2PYsKwdioznFpuWjAPh5rkCEr5Za1k3QXWiZ+8IPri88lTNqXuqpUvF2zTtWqPp5yYLUs
ZCVyHsg5Za+yWD0CSTTmdO6KEjplRIWTWB5+WbL4ks3BwtoDjCj4OI9+8W84zLUzuLknl6gm0mrz
mbpqt5tNcKQUEvzQ+SOq5eltf7S5fl+asAQac/FBZN+Gb80QCTEMhgR2Y33vYE8FY+KEhmebz2k+
c1Ll969BDeHDKkENnRKMtURxLgcJ+E2eWBxnmJmQev9vXiUwrR435e+boaUFYnhrn+x8NFSLwOnK
f2B0vU9Hzia/qI6yvldpnpJOcjXFrvunLWdOYNLDe9Od5gzB8oI6UxBoQquydbbCyMkMReF+7si+
8F/AH+/nub5nd3BV2j9WjRhAWqHpl8BkFEFX6zDCVMI/fP4ferUt0Z2Req3MbW8EH9GI6zuaLwmM
CmweBlpmDbIlVjvxeq2yMROBjxhc8+Uu2J7OECryJ1CYvioCSZrYBx/FB6Y/9cqRnExSCf7+XuBy
2pL581HrYxi41R58e4JC3tXTroP1ULz16ir08wGt3xnqk5lHXM5TzYzDSpTxYozgGLssihcS4rQp
wZXfY5DIOxixS/YfWzdfgMqK20dV0YZGRLr5llDllungUo0hZOt3LNGd/DT4ARuCeXx+NcbZJHBB
Zkqdj/1tVMfCyXQK9qyn5ztk0eFsDBsFpW+zeQu5mrCAThfMuooufhgva12Q0wYOY/egaJ5zVfDl
bCmLweCfzGRS1nL7XhFN6KsP6F2QOBCaC4vGi/F3SY92URH4bh4vNrkQbj/6DxyYcuqP1pJBYEKo
gtc28mkKuXElgObWH/E7YJ1GybNPDe4c45LRSNO/HBgwLWA5sCyBlgRs84KvJ3Go1s+pXo92UXQq
kr5jHEaK8JJIztCTc+jUm2mkI1H4srAdIoZZhr8GRZYAjqtbVLhS5sWQ197afLC75W9JFVSEH2sK
Fs7i6pnd69uv0856dH5eLSh2ObtVty/TMevDQMpI9RpmqkGBjcq7Eeq0QHXD0VO92Kzs1WdcfTqR
Ic5pSZeKVtzQXXasza8KYAFK1kbR6Rolv3XErmlttqXG8nauKIskyxsuxwH5MMFvEY4rr6C4tt2c
1UivQdu58T4TXZZW8slMkxHcf4vzEOkeR81HhbZhbzdOaUDlOdhsKmfk5PPh5Y2+Z7I2tSeskKwv
pf7oqA/QWUxUyNfwo25/Y4JM+LjuKipqmIW3zBV/Iwk940dG9wKBFEmqTUv6gRQiBL5wZMCYFf8t
Hj+m8khvqm00t/i3FH0qdBNXgzMAuprFJQqlLnTyB19Z/fWCSiyOvTLLeKSJSXz41vJB5sOMLS8a
E2UVlxgnJuWJBkCMTILfPNVN2cHy5wh3dyuVDoAIIpgzPopLgrdByesVsYHSCO1krGG1ADqVjcID
F+262bMwh8HkR3Zh3CQyIvYuPsKJw4T+w07GvNW19SFLfUZ5iOGBYbl4ULvILj6s2kknFa+i8qkU
wEj6VlKj1kjyvccnkf3J53yJRhzd+N01aVEV8RRUj4KROzpeO0JNkckiocgGSJVKSlIV21l0giL6
70bywffQ97aanx5SeZ9Mge2liTDGMqwh+z78WP+cH+IxWnDBLDkqSWD7FPa4NHWc4IvYrZuQNpcI
/JjhWUP48o4RtWzOFW8RV5zupdifA3tie+aHp4ooff7gsB8AyqFRyQe0BhitW47SnOe9a93JmbdT
Uxf8LEyMhuk0mJA+vJMc4YE4K1zDgDE21hTmSpKF3sUcDgWbFGBBL+CGzeQKuo7CwI4Wo66J6UKy
TUN2yNcNjoKs4hCGL8RPGvOp90q9juM4GgbdMROb4yylDUZiTlfkYQ8jEyi8RmdIDndCRfdo+YzJ
`protect end_protected
