`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
ZcNQHZ6hMAkO/tUpTTZ6s6uB//9JdN2vLuU/FctEaEWvdGtA/+SNR+Ta9+vuevsOb53R960vDMhS
5EWzTGUcJZTF/8gV22c9q2v9RwqfthMlQ7g4Pn4fNDkmDZ/ObT946nfdEU+R8O1RUbre6klufVku
sMTfxgDd9k7IXtGyM0WMOzKxkVW/J5xB9fQM07PexLRD9g80g6YfcDkfcdYqggAa27M8HvnXF1cg
KpMFG2UxLeAOE6CZV0iOscNB00FGK6RFk81QfV3srXoYmCPn2f94E21n7EoqI61eBkBsNe7eil/W
SLjZ/ZIClrkOZ/kRRSKkHqF9xj1N7jipqM+3Vl7gFkImVn58jCcuc/itT6FYrkEtVPxnAQI73Ewc
lDOy5/3ys6jpkyqPWR6yDT0FRaYSejaP0IetxrmZkvB7oJLsA/W4MvJ2PMOZgX1aUN2eEgKO5M4I
g2NAlonfwCRywXrAgGd05+JD+O8R50Wj5HNx1t/n1nIBqldIaFmbl4BftfsXFmFkgNKtFJ35tIVU
syFBhqkzt5MshzoWiW56K+N86PFuM4asB/TA1sqU4bp0Xx45U5O5rYwg3UlbJu5EOdgfpDWvSHA4
cW+uDaipbrLzTQab4OVaQFVpTQ5Z7qC7xvoWPpTZNPiu6AMlCLE13ZUyBxxXw9lTnFThKtE0ZrHw
2AXXbaM9OGfQFBZY5it+dQwF/GYwCMOHqFKVjQMMPKuS3S4LMn/goEmy+eulTV9rp4U6k1HnBa8M
KdcRdNMIDcGeIIpIGvwP2CSilfjJHG4W5tfikYNxTtn3sLi1eOdZ/FKjainh0p/U1Ybs0BFEwUlc
No7OTrzkpVhLG03C+ISRRIbGJ1W5XTvilKG+mvAJEFydWt1sCiBDSPtBxUAFPKHzsiCy28NNLP80
T4Tc8gcb67k/Id1LkkI2fh8ASdyttlhC6LCOUhcXXrTET5ia3H3XY8o1fCkon5xLjEPSoy/WVdBZ
MXPF+p/F0W/bDcJnuFUWze7t705MOTow2CorFNSIa2ehqhmKTzy1mTMSpv0Wvm6T7ylN6FyNzXgY
qHEerCxqi/wInlfH/HJOumdsbX1805P42uB4KBKv3vQkpk/zvmIskEPAhT1k4gD6rBoPJqOTYsdJ
kfHvX5dTWQ7PartVCO94LyjrvL+pcUOn2yHSg/GZaHHxYUI2nwg+buXc3Nw+zPwLAE6FN6BnPe0d
5VvWj3ipcehySl4a7NyDOIexyw8Rd8HA0RJTbNOqJLuA3P69QU5bNLIDBEiR+nZpiCyJFiploOqE
NWhNj9A6MIiVvy7SoSUuwQ3KEf6ORRvVxbiPPa4I2WUC2736HXlR1z16AHpeB3ub3tniwl+E/qJA
bUIZXkQcE6PatHJhnX7vA3o+ZAWIDEydiQ3srmP4d9Se0eI/NZtBdFq6MN3AQOkb+MhzL3RlzEbR
dm4OE07aVBA6ZxBa6Qlh+vMcIG/IdIkVTiIVyoAYqkepe3HKltV0paN33EvEIp/McxsxqVP0uOsJ
TVXS+vIyEF0eQ8bYGgF5puYBv5gjq/8ceKoQDUwaMERd1uTIkSIFOO1RIDOgdqo3TwRozB1M4eo0
OYu8guVv3j7LndRswh9ugN7tBf2wrvbUjBFKvOR9nKwFOYLhCtqUdMopQkotjlO69CUvFAwR5SiN
VqzN7j0DVFfVnRZiI/1q+qA7qwsgl9Efjn+K+heCOCPy8jHOalywwix59XvzCcrXiODgBoFqUBng
c86pfpz6FAz6bxm/ypGBS2AmeyGm8ZGX33buC/ytHWSNeAcXcTqDzKaUlDpnARB8OF5Us2TULvsB
wLYx/nqyJjJ+PHrJ+vrdINuNU3eiN4T5npUrDE9Wz2lW9GbLrEsogMHC9i31lXsQfT4UCSvVKZVH
1CtE076MZaJRjO+tEVlmLIuZLwJBKQ8xRJg0fgO3VY3VmdFPxt4Gd8kkL8Lz9nv72S3YSzqTst/7
S/82Y9hqleYkDonDa1h/wIJvyhgEA24LObkcs1/9minE/QhdtK+QEzWOZKEuAlCShWFrDQeULJl0
iYnOgtaCtYdEm3l07duKG5LWCp/Lg3ABWzC2VWNNJ2w6RXm6kuyvrwPgGIiE41jFGdBctjUK0iZu
oJiJOB85yzrqRJStwBYWfQgd7my6GslOCp/LKn/EsTRezO3VIIdKoqRS55sX+sHGJ3b8dgJd0Tjx
91Ker3LCxVCOVwtFKHqlzew2lFEEYuGm4cEKbFA8vLMr7fSpPDb2fqtWT4phZv1ph7XEEdcYoQw1
/uAAMxA7TCaCQg5fXlDjL09q2J9/8oD7/C+9mco4YYZk4GBq7MKUOAzmAqeoyRzmaZDETC1/xa7M
vd+QRpbjkd/MEs5tTAEIvZd0sspi3rOqFaTubq70lOxNsaQYxn+Nqxev+Q4jeFd0iAgP/i0fBajG
M4+hIJ2iTT8KyFMVn0whr4wZWqOdO/lipqrsREX53KNLrOpIvkI4L+C+G5hYhSN6L7WwDSWxCIRN
sTDifGBHouVV5DBh9h9SGjIXc824bcT2com8nCpjxUZmvpdbywU0tWMgr4XIn/Ryq/0mlybKCosN
c9lCU/VfvXct5mQC06on/s+Jwr/PX9RuG0/X9HxXEcT5X8muQvZp4/CSQmFR151OD01Y+Vzh03FR
fxQyJNv7VvaSJpLufFdUFxLEkwWcvzcweYeHQyAgNDZDA25+W45ytfUOiMwnXiwkYc3URgXRxl+5
Oy8fp9iiTOd/vUdDXT+i6OcMfe2L/IAlaqzKJ4rCXDg+EIRQHDcHHq/WmuKY6tY3yVDPrw/1pexX
aVXSrSnK0GYC7jH7/ZS2hxfJ1ohdrv0E+rsciK1fMrQb0O9g7sU6nr3JViEYR02sTAFHiT7e00HY
tYIsevCp7038c59GNLOpTLrtpsS74dg5eLBzFO+DW33elMn67sw8Yh2p4S0bQIgAlL9XP89eocwq
LabXXbwr0QKezVa2lV2HMTI1QW+Q53lQawbK8TePjiE54Q5aJIApqqkVBKG97iWFh82Tz563de0R
AiAUlV0o9ixVT1iuMP+edHIA30MZAwFjiJHADi1zvT9v8ShmXtTy8Usnq53ioeIgqcLorrLWbL4s
rj3W/QT1UQM7aXwbGT0PpE5VoAwWUTMYruG/U/Rhkq392ReaIDhxwNGORcqSHdrrl/J/awLCxUE5
kIjCmuMQxlHv9Twclfj0AnQ+0sTzx3mLMaP7TY2JWA6H8psOr3QjmUGfcPXirMKbCDwJGR9ubYCt
kKuDxLF21X+2HUzANY5/n5gsmqC97jzlfeWMXVbfIJKUuKgyX8zf/dRd5bSLKzoAgAFUNYTBOIb3
YS6Oja/cxAgrjnbpkcVdOLvNDxtI9Jc3/4/vhg2q90UElBCteSBnWh3ZDedPm83lHrYJB6FYnMDy
43+UqgwYbRXRZL288otmWAz5N7qIjZx0mpe4ojQMi4YZcJLNkSxm+pTzzKed7942ZVh1kvUg9BSv
Vzxn/iOw1rFAPbYvZ4CdraQf+3xjVxhRLtLfEIO3DfFdoEbB6kqcv2GiOHvaMGfDDrwtQCkdn2Fg
gaYZMYKtOIdWPjpDsuXtXYluND3uh9AawgkiZnf7ccSY9cvAABhBDW5ck4mf0fP+NdMFnf2T6XN2
U2YalKhiXOQq+PXIGpdG8bB6INiF/5j6GVyovPTqugq2nYmX60e0S3++vyRIi3kCnW1CWlGLKA6k
yqba1cerFSpkVnbs9jEj+1aUWALMLVWdz5a04sILV5DmO2BRrOmtxrx/l1eVDMKkw2g5+9ftKER+
SfvF53bpiYHUBj1Hrs6IPd1vaZX10x3eTrjc3//QVtfHtD63hfIz2W+aphTIOhq4xhGQ+q5HG3aP
MtTlDHX3Xze20lcmqE3OFQi2nGX6F9raBKcQGeqRf6G7me7c4JXpeLFw8L6VY0hRNPhMuuUmnJzL
Lui7qPkMPA+UsoycdM0mbLpnE1G90UILHg4H6iNxHw6jdoj9a0s+LtZzFKek+dQqpxKbHnuqxV1u
dPMdS7cigyH/SUsFM9sj/dr4PmBisl4C5R358BsWWRtqew095maG9pG/n+K1y+Alh6EWOPZ7L0b6
52DedxWDhuRZP72NHHNtrOVsvj0gL6PDBJ91fIiFeb5Y7A7vhS3EfkrVv04JqzCjM9q4tM+5Wgwl
BWNKe+V4VyiaAzRzxU3Btbw9qo1QcfFLiGxf/CDvGoVYDfmiyo0jrb2lvPr8tOzUB2nOeKtnz/0n
DO4Uf2NpPkYjjtHakTDUmdhgje+tEC9lQuMyPHvHjXHtk8eO5Z98tnY2DpzIvlLXd8pJb/KSNCk3
CmQGmorl/8gahJU0liigoeXjUAuXBkzB7u8357+rpnsK9ebIinuxChgGLx7Oa7Fi5+DeBiIvJBO4
FSC3VSsQSa8295Cx4O5Po0QUk2Xgytsc6Tx0IFWQsfFBEweUml2CzTzhk1YfhJNqAx5PbWF21gS3
M/77UM0iqTFO0IP/kpLPFUL5qNPyvsqgMgVBzHZJzB9bO5mzowOxliWoUFo+EcP+mZBm2/KfsPwD
B+jf2vTLC+TymOd2qBieGDD5Hrp4XQDoVVz0KBnYrJZimY7pPcVJ5Y837RZgc8M0T7sDz55kZiCc
oOugPUQHSU1AGsBq9I1uZJmOt8Z5p/VPQ6v9cD76nIHMDP+OFSo2HFcRXzCGdAZ7hx25pGPhO3Ab
hApVL40ND4fqnWuwhqAN4aV9W+MqHBwS1gqTE5Yc5nkNws2/7/LTcXx73cOQp2I6XvL6DlNJyQi/
PByDG6aNaG5PW6T/MA8xHtDBtUzSPCm1zkvXPCEu3QzAiS6jW6PQtlqhjuJOFFhxxg41pwDDs4Wd
zMk5rM42VP5a1z2liH8dMmyyHfxm7PxAPslYgdVcZvdO5ZWbjFto3GczOmfWJn6UpfNRbtpwQADg
iG6cpbQV40IydJ5JUc4sPkNYZio3IZfJEpdgHh39PehRFsJAmXop3ufqZQVKnqnzuqwdXBLlF4Fb
9wx/SX3/SBjma0JpyAxDs5ln685b4NyLjNsPKv+sEylvFnair3WjfoWswWAN9vTGA+OuPfFE8mDQ
lHqmq6IN3/3TC51JTDMqiSw7+YczzhgkvbrsF95AKxD9kXmBaj6GdePQgArLdV/RhLr8/c15ZFcT
2x7kkZ4dlNviJj3j5iyURbfwuxyfzgPC4wsNT+ctiToXtoYMD+rkRueTp+zBAFEymSZi+JOTpJyg
PL9wz4MuSnA3l2ifT4xffMatvQ5t6pUyrjGcCFVBVK7fcteREp93yabnQk5wiEDyk5XABsLLayDi
+O/N2LwCQg+y8MdeF0Si6ZOblRCxCc/0i8ZT1kzVcVkycWXTiaSx4YVQpwUd6aCQGFVK5ozJ9INn
dmneUIWto3IJQIZ1hxhBE/T5RjRCvrPSJ/lPTt8KsGekwE1qkvH/I7VMPOYnE15Zl1QTWKcgoD+A
fn6+u4u1JjemNdWa2lH/+mpiiPX6l1wbUrigUpnaqT3nDrPom1uigRxpGAxmWeRcxR8OpeXj4QAx
55XzoSZAghGnW8DINjR70fMYzaTxbn99lAWsnoo15v/64tn2cIG6bKyOZa8BhkdioAG5OsXoZ88K
W0zS4EC84ipPj3XMeZMZf02Y+FNlDdM43CwvUX9IQkulvfU4bX2lK42LtjYEgxTCSo+km/Kwidiw
MufwRv91vWXxHRnonZMkO3inXv8/ohmmk1nssZk4UAOKVc3nADZkD8Azc/hFsvUjXT14aKOGCFDd
oX/sfv/3TYpIQwQ0eRTAxS/aOtf02zRhwwzdXBGfAklIc8mwnrEWU0/jOdSxkuDcev2sPR6Wqthr
/3pqX5AGPOCUb78/B3IntS99oY1QYi0LyzmixbUja7sz2HPDb5yeaHjVYmo5B96Wy4zFJm1lGwM1
xr16zW9r5w+w3qR6Qbu1t19ZO9bQ8CzT6+529BQL402mGrRz3yNtlY5S7f0qtIfvK33+5RiIVdT9
K0A3Kr2EXwFYpLqHUgVFcrotnNso3N82UIn2DqFK3XBpJMtczHMYqQSJSKUNtPis4QkBb9tQ8Cu5
DWlZQ4KSJok9IZkr5ML/JBQN0BmcegdUH0dBCoQr2R6uX4hCLaHkrzi0AS8lyTl7ruJkeLFTaZ15
1tsZzKwzq7tD8aPjFNIKOIIUd/Y0d2MkhXYSSbG+yw4ttWvH/LlHXaqx3GS9sOqr+X6azUxlwdX7
0G1frtu5B4ASyKSJOuPYSmp4cqNXym2dazeD/LCHiUg9v86iwRxOT1QACdu8lAYFemqraw8PDWrx
SxfQEKRg1lVI5/N+qnSZVsxCtOde4pc7h+p513sICbjSXtAmgU4ySM2yTWOqMn7NITzDA7gOT5DS
K6NtY86c23tI0KmjI/YPW6jXmEB61jswV5/LOxS99R7rqBOqRW+pO55t8zXwB2jRnQr8hQQFr2i+
6U+WLEgb+DqpYP4z/rJMtXjQQUt/JBqlKa33/bUi2/eyobDruhobX3kAZfPOuJ/4n6yx/5FHPCI+
j9KrXtjwMaxuQGJIBVr9tg8l5vk1HNwZmM83SGE6o4jwIOCq1K9dMLasx6GjwK0Hqxl8Yy/hwGJ6
QZnA50seHjIE2k5PnmAN1LBH/qFCFJ4xSU+zTieqAzGk/b1xEYA0HKDqR6CStBNufSVuqMJ++RIr
yDOwlOsjO+4LuPin7Vijt8apMzSq3oR1VakAuEw10bmmwdaBjxbk3K0dDh2e7YeEn9bwXvzxOHM1
iB26/11w3ihtP96GrRVEl+ifiseUiEW0THD7SUikGDhuNw4/RAcagx2r4U5bujqC6i+/xB1OZQfq
tw5E/faNcmxXuwGntTsnweS9hBppy02+/15Adp9hoJvoeAfFBwFvcG2ZXbPauAkoEhIcHN5EQHxJ
pl6gUOxPnuTZ7oPULqP8jImJw5l4KP/3R8FGBzf2OYI//t+uqZzVw1Ls0iu4+Gl+uNEv+T9mTYC5
YYQWVPD2Go2jgf91uNPv9X8bayLMvV2fDkpfzCzkQ6qvK8TDb1n5roOmo8IfgBqRz/ueUqoyxWXi
luH2badTHo8NOCz+ceMZyWcj+erB2YyMgrGtVQZrvZSs1BfLcL3cO9PgVGr76o8rPPaV47pyaSQ5
HdxcizfDuFeAV4zamLUZErrcx287AE4xJJy7Ion2KsfGeRW5CgPL4AW3qylKMemis4TvyIGV4ckM
SoimNMzxaq26wEMIhln2M0xk9ot4AeV4fbRZO8rA2qhhF3PGYM+o/FiCS9Qo20KocMm+kmwa2iyv
VMcIGFfCEAGzyoEqiq8jSAeD3yiI7IN16ylMDbnrue+k7fYi00GrAnxOpnfjD4OlBrHV/87C+s7g
3p5ojohri8H9bDo/6vRupKMI3UOHy8twNg8swnZU9/DrFLMGy8kv81KrjU0aAUZw8W1L0l4IC7s7
1Xy2/HWV+6oa129qzJZbq3MqR0/WunDAb2JOBAXg2OnOoVnxInvwmPT6525t9HR3TYv/2hIfc9OG
ymMPiIgph0bUVznzuurvwChVOL2ZjKp3xcFXYlRsGVc33tDqHKrAZSrwe40FqopbDtfObrZQx3PE
dvRJjSEuB7bFJCmG8OF5wVmNu5prTEBhK9iu/OOFDGjP0fdV+bXplmnVOwh8RDdXjTQ9yZ8YcCLP
yiqrROxi5RymItBF3DRaaMTYyd6J45Sq0me34YDkTXAzIz282e3MXfhqnKgM4Q+BiFbdfbtaWxTs
+V/8vMyL+KWzGl4gjtouV+wTsRfoj1TxsR1zaeBskloewF0ERuYwnjUniHUhtRTkD+ZqyiiGQ/0G
SIzTK4r0JoJ8r5IXQAbXI23C0NRm6FFGnfKDMzAqoh0oN2qjXMzdL/2GDCYkCdviqEcO0LcMMh0U
NonpYP0M7K6Wdm6ywjfNbCn5XCgXfCqvaQVjJSMPi6ZqEPw6Wm8P0bZqxmW7up9f1jZEDdggjkYt
lgQSxrnLEi6aHeq5qx71DSipoRvt7fsVa4aKB9tf8R5fxDSlRcrANHoAfbK/zXgQDVcSXS9XVRlw
UQHrRutzOvEiQF0McabGfe9tRbWR2agN7RZ10VeBFrglJQHnrF7fMD2sNJW/Et31e1dPSg+X39W1
/CaICUUI2yuzYfeup2cW8hl7xIjtjtln/xm8oYOvreqEuIyAdpXIQ6Q9xP3BAu5RyCYGaZQAkuY9
LK3Xe16fPjIh0BmfxIsDYTU9ESOtDWNvpBwCM64gMtYzDs3f0vgxWP4leQe5So1T1ugoSIp2QCCS
aald/O3pGfA5zNwGHuEzD2At/TYndljDaFH1yxakFpcXNdibNjh1JSRxf9HzsN2fRBOk5uxdBdhT
EHH8rC/6PJLtmk/wBZA6oW3eHDnRJhsrHnRQbBneg1r6Ud755WXF3yl/O/0CKR5iBrnHfBVH446S
p11Vt/NupMBYja9idio6dyjYG8ojiFAc+DQ3RX96eaqfep2UChjbScDctBU2ZTcbY0CO/b9+nllc
R5luG1xhIQctgZC2IngRLENLUY9LoZ306cqb7Szd0Cv4jXDjcHmguOxX5zmTRaloleH51YlTnQlp
cVdMaYG9ic4O1/ad7NBDruDc0LL2EGQ3TtRtG0VDyBPfNNHsZex8if+GtA/motcB4enMH7jr1feZ
fNRjl8UzMsnLGu67NQFJ0ZT0/Ua4XlKjH+9XJxJNgDLaY44UwyyWmVEgteXpZdVw42Px6lilYBUD
TbUO96yxAqDdP3GxQYyWrLhxfknOR8K0Ww949WJ9T5HpA0QI4nAEaKW8+0o1Qjtnu4qIP8aR6rM6
2HFrIEu2JdDzNs6ebstDZ7nB/ME6d03eFBV8IWYQLyHclPpI3vWvF2gC8hzz5to1YKv3OLbVOc/j
ByvhM8pOFCqxmKDGYuA4+wsRnzl4sTdXTVoQy9+HuIQDtAdFF5G1ZiTU52GgLIhzLHL+/1rrrx97
QtBtCRgpbVWxyn51L+yiw6Dj+l0/+sZXYr3zfolTsvSMkfXz/b2cRivAVNqaMyXNq1VFkAI7C2en
wfd3f7dMxRGkTQOV4TWTUV44HEy65JwxxmakzKUD8+sBt/p9t+q2CXYM4uuI5Zp52zLqvVx284nM
caVJwoWtn6RhXgzeQf1qJIQIjjSXCHDqCOr+wSLTD4DnYuqdHVHmyGGhwjWUhTU80CBt51E2eWfN
p1Zhg8aEr3rBXBWWOaXdacHBSI17YAXvo+clfFjHHw1gHAxeS27q/rwrzBXRz8Wbrm0gJEHf6ZWK
c0Nca3i1I36Tx1kUPwkWDd15ZfRgZDxZ6MsA5yZmzm6PM+o7Gsmg13SN4gckUWhVNtW08WUVwGzG
NEAcDGT7ZhitqzipIfN72SU0B1Bjnq9D3EEtyouEgpa6kTvH1r/D9jUba4UFVYb7i3tX2ZH2dV+J
tn2bEQG3yOZP3QC7PPB8gmfMad8AsEfSNmNHUbbEgq8FBZApxGPl91J6ctEP34MIaBH/a9Y0T9pG
hD/EMXkNZucDuV65qZQgtNY4bDmY+0H16ChIj1XgcLfarpBVCFURv0V0qOMPCXYDHLSw8SIgyVeI
45mxnrELEwAYwQRetxy3MjDXBKH2LuV1hCw//I68ASUmHza7m2/pvNULR7kuQzRyoxgGuTsM+X7Z
nUAZlyCIh3DAAsHspIaJNd+7Z5T+izayVpfElBSQUOCNyGKhLcMesSlQNTl09jqCNvey+rbXaHb0
jxvaFCOFpA47FObgdaGUrcPMP0jDsmOt4QP393L2g5KNkLhhr2RB7ehmJbIZ5YkjLSnBm66k0Twc
7KL2V2psAsss1EFj3DJM6uhiqgmXUebCGqKddYOJD59ccJD0CLGXujD4cA2o1lEgzqXo/mv1eoSp
kdsKkNV7k0Qu4Lg82NHAnZxxmVZaLR56c9crJF52RUYKRHw3pAsbd1lW8nraHD/XrRaIl5KD5WQ/
t7+nBfEBqfcJq0Ce91Yz9bhca3U5NcEH92kcoqgcR7ItOJ1ThXyIdrziTo+31gRM5ZiNXllfI+QH
BpN0Yu1UKPuw5EnHiceiRsYjC0SBWTyEnkdC9z252LG2Zv1qZsENdbrJB/Sn+OgqPW+qcfAKW8Ka
Lrx9eY+2lExgYJv7GP1rz6und22oQcPr/4I063urQm8mIT98ltJqiSqdFKPIsAGna+VSv35UuyPF
mS9jaShzt0xGrq3Zm6XZEXPklO0iZ1G/MnGHmS/yGV44uek43RFz5PN7gz+gWGQlLwS73Vba0PP3
pmAknSQAsXUie6pK7ENeJQhzRiEGOgJKSrPqKLb3g+6baZo244XvlRcvplaLM1fC5wLkWx+B3neE
sTXhq5iCM7IKdcSHjZLUQRYZz0bm6ey7HylRmARj1ZC4zzntWZ26TXEiYlRbcZEkgVoefMHq5f4H
P7knWCbTxI1WRd2TY7SuHQlqmdS/KlSEWrpkAq9Hti3KNAmxYYXZlymcBD1YzavMiw3jWxZ0bXPQ
iqO5xNBBhE+dUSy+i8T6XFjnsYj/ayg7qUbNae/7e/m2SY8Hq2gqhk8qU8WKVoymykmOfrmlX3S0
ygq9V/v8ekMndhQIJHMMi+1iLA+2DfuliLp23CM3YjIXhgxUmJiiBHAxqz392DquN/C6pxpZGC4N
ng5AIZtsDGC4R4Ybs7jCGdeKiSfjUV8fV5VZVEJmXVk67cuUOPvUQa9hDsps18mZalY3prS24xc+
FWrd1J2m6OlO+GsLemh0UuyNgpIf1pZzxIkS2nlr26ICuXXCCPUJSnMXA+es2bTt/KWGVEEgHHpH
vpPifNOlOWv96rHqmnchVDv7OVEkIWKqo1o1UiCZBnuWZK7NAVNnBZ6KQ9MAwuqxpXSWU/M6VHkw
86d/bo/CeEc2aFvy8bTCwTbfFiVBhzT7uJfqlKLSdg64HdCZRf+2JvsIY8iJ38on82tfAf/mITpn
GD3qkjqNTGl2ixT5wEccJ0pyD2mX3WIoY/CPNTbN9ktXgLU1C/S4xeE2zQxCncy0e9fAdPANyWJ5
fGY2NZ+Q6c690jbZTEHCsCti2wQnQCZUq0h9/1m6ZquPBWu4s2ysovtBPSH3OHT+IWAObWVSbrcw
9djqHGrW3rW6JO5jTRaNHfz/3SAAjoR85vQJMriiuS+7x868bm3HQPQFMHYX6upmp9/ZWxe4MJRh
2ZeWKOZXVVFJ5PaWvZkvbbmSEOJ3HOrbpoyHqnoKvHUH5f0p2QFE8ERO31A+G4wC58Alo8Za0rgv
DSZOy8nP3bxYpZN0xwDfryYvLalAIJM6hRI/sVRb9r+My+2BlqJjyzUcs6ynohB1duW85BsPq5y3
jtVfk76QA3toWbrH81ZAzkCRkWenj62vNxss1DFznodfEUPIScAFpqYdiwuGqHyyGcVLAl6iDx0a
KB96ivFjD/hsdEQvaOYTVfHFFJWXYVU1iXwJC9ItxB9l7DKbDp7LCVs3zF4BPQHQU9YKlCj0SKSm
riTv8tAFKwh3UzWhfgYH7v5Hy/lSej1eF/CiMiGeGW/NNz4EoSweNw77MbhyQXoHoCYuRzRLL3Dy
7l5idvuhpFesZMk1NwjiYUeYL9x48ifHf65V4Km0+jPd/rzouwe3Fm2a0B95Qvg9FfX8rmM9STVh
UfJ4Jm2lB50FKoStsk2lmUasXDiswidzuMhuLetMUgQGdcySJ/YXR3/iRI6ApUOCiXdsoBRPHvwh
3AT/1rgUTH5FbDnMXsd7CI2tM5PSEHfMnyR+8RVjSeYcr4ciS9+7PcRAEBu1LtXzcRNMb3hmY8wo
vi63kLz9UfLJQLeb/dR3+DmghAFHvOIWbl+AIAjbSAZ2RIOzVMYFqu1JzHi5LauRbNUXjmZH5dg1
l8Sl8ARunYfSdsyKUvwOkJotncVDGZu6tyei9maMcO6fz8tL2KRPKX9cCMSJcD6jsSOyhUcB2pN5
ys957lcnPMeAuIII7SipFk8SDp6xtpdij7MhERwfHOhD4+ImzLzrnLYMylJxOhfgKrYEcO4G60oA
lEj5SPRSUWOY9CajmIkvm3kZLQR0ksqihr5qd9Y7en14gTSvF6Zho5/S5dgehWPZBKkJk28uAgqz
eGxiFiMJDxgAX07Nea0HgBqhG3T5Maw7O6VmGo79yO3VzRPSkhARurJEMSOUP3m15ubkZW/CM2JH
d/Li3D6i8e+nscCzOYm4U5VWZZn3DmvO667wgFUhCy2l6UT4PilxmGU6YVHgzEheJ4EFGcq+xsBA
Pr+VEgBAZzliJLC9GY5vRPD9etkpDwroCZi2HNXSn6rEs+WiqXceaXHKDBmgvrzEZlrNhfRlf0G1
FgVTWLGvrEUPPebVeEchNcK0WBMajRTwXvBbD5JmIwU3TEPviO66RZWJnBKlB8iK5IxRNIwJWVre
K5rdq9r4b4BVBlnMprXrrUITyAhg1vfCXwQDs91qSbjP7efOOguN2NgRGbYdFDkT0nEonyxihIA6
C8gJikcBhXDTQ79H0XTVWHwK+Qdi+lK5BTur6I1g8/G9EDhrkTjJkpm3fq+JMFa8nFkiYy+hrPmZ
cVtzUbc08fZnB64NAt8CYv28yDXNT0wxx0P0rSdG5ycKHQEXbMwRXY7nJgoVp5dgD4kpfTWo78fA
Mwb+kJ3PsAKKoNKr1e0hhgk6f/rNa5dr4oG0mwCsVbOt3O9Mk+2dRRgJBnCAaU3lHxnLsLZkA+2E
/mVeBWoxP+QwvkQhszcbSDJVUN2GtNpHQJjo7Ua/U3yiP/weS7lH0NRdwHxvVR8hCz9wtIJUd15g
Vlbibs94Zs7pHpx7smdWVxS5iuiru8iGrHq8Ug8/+aL7bWhxLbpt6dQF4XsNF0Fs3pkrs4OQGJJb
V9/0E7q1PRMaTjBg3p30+9iyuUvaQLJkOEH0283Yzc0HqBy2rXaq8GjSwxn607RW1KD/pkqBclVi
c2iiMojA1P66z5ALQbW6XZtmya17KZNlXSPe0KS4QwkVQMuWAE91ljgZX1w1xxKhOsY/rlvGFrqM
LGMSuIlUmceUxCxN7zTMLW8lYw5xIw97lFMLlRCg+s8CYe7t57yDNNjV8TdHWcH6EzKBd58jyhVu
ZVNdi03govvGzisOAmw3NqiyX+T/z8vVfTuCcpU/MjLDgRG2BBFspNROV0X1W6tcBBc2JWrwqGYD
va221CUtJ2sVQrKKHAs8N5bw1zqLhNTFzLyqZ+NT0wVNROjHr85JgEA5n8MZ1xTySrdkCMps99lW
Z+qeKpdE3TzgwyA19XVhID0oIT5ByK2PXSkmGr9RG3/10xd41TT6a//EJVjE0ouM7JrnTxT4qpU3
ceABQv0NhNhyBaHDDMRtJWw3IjwWlz6fzdILlk7booQaq08KZDo5kap8oD1DEkauOQ+i2OLgfV4Q
Far8/zGudxcdTsXu4IispbmEAO6WsVdIoqXkgpYUDEIYafJ1y1jUdHA3tOUtq0EmzpSWdCPKFF/F
yCqAiU6JyD+Tqg60zVvWHr2mEoN1K7jeub5kTkuqXMMDy6dc0mN/0tPLEPkV4Rwod4bZ6iVx8M6U
cy6Jjo4mE4Rr/jQH//b1mAu7+W1frzi5zDnnRggr4c1jZLwxhbRa1tgTynMuEiTZCW4mAAjUKrG0
0SD5drD/SCDy+LzNtiJsJFIH+Cj1HA9pqZ9m2bZUh0KDCunTsYUog8PysZM4f/bFVYmaR3wIS41k
fx59saFtFeu2r1aaJi66F3fX20M9MeD8xBfHs/FHTaRPAne8hCQsRUnVIkMslLTS/nfl5f/vY5Pw
SDk/F41CWLvN1S+xQeKjFZLpP/weZY0XezA0ZUA5Y4R17GvAKOcy9x1+9P9gt81nrCEy/lamLLtN
K4RryrY7U3+lYOqiF/M8JkIoz2yKFSVSoLlZz/ArJRCZYHFKRnAJs4PHGoOjyFAdFXxSLVMN4mKQ
i+VJHQg3+MVqwfPK5KJ/IYKHA00CXQuwN29ewcleXTpaGsqG3f2RuGharJ7YY1jTB7k1srnf2Dcq
KlYosx9a9msaqnDBDEXIy0PECzpnfad3COnsSDnZECgBI5XylFnVehEVy7B6BQBAvlqF2ElslbeC
JD/09Y2tAwh9ZEBGOkMTQ3i62xiLIhPztz2WclDYv/eJcEvsfPcHzy2RglkOGjJ99DI4qR4/LYXQ
3hMJRwq9ouPOmQmEKbPUaB1qLBhNwmwsteSq70jkYY8iHKU3zzySnJ9SGDEdsJlk4p5mz0902kqx
ftesye/BZc6Rs0bdvbhhQ24KAy0SKHdmlVc7kC/qtAdK0/oO1jMWFQk+/zIdjyPv46gaunxlsSAu
wX0MW/QJx0SghR1zzpL7t5uoecGIHPSnVVW0xhyePwOIIj/Z1zL0iKqMFF5m9UWmoFdaQz6tGGqR
8alR2rCqPy46KjuJGZBeNhOKHX21QQrKdBVQ4iH8oJKSDMOKtfd2j3IN1+zK+lQ5Kr6dKz98QREP
xyou1aAoj0J7JBFtDGWTCZXudlvnfaQRNdmw93qV/dj5WE2Poy2XmV770iRHd4VIjqyF0NU7R+q/
hG0NxnyDeBkVCJCwQ5KUFAFXtauR8sb7VtYx+fUAAkhdi6rZ6bKuhwl2dHFohD0wkZpvIIHhUa81
ze1SMYZGBd+5O1wrm7dtTl+2UfI/BFRo1e5gCygV8CVqqtv0s+WeeIcUJd02AGqwCpRQAjB6lczn
1eBp0On8ISxDaSYovahWStQmSK5eaumw4+zOfvGj05IJxF16NojAd6BDzMn6qOxBzfNo1NMWLxkF
0jPVJqN71rPd1fNQJUZPS93vN+IkuT8J0vRVkpFjJ25rh9K1LPuj8hASgAwbjR7XMb6ksGE9um+P
TGlfWSTt6RCVdzbKy+R2sDDY4p+iPRFQfabr9VxYWxX2stkvrTGWt6o5UasYzjsEZfLEvmSs90Vd
QmHFi/ekv4zuKQ5CZ/lDmSR7D0MVVIDMtj3D4M3XNzilp61QtJsiJgembub7+F4BfbyDNH4YkObK
aTa6DE4osptI0arNeGpRXrGPOtMX94jsSjz6sJ/Uk7vpCFJlJmNV01uEJSoz3zM91f4hunqlzGO+
n4K7/s1njAC1yiDMgDEY0onfouxpjFoLFJL8GPoHO7FJZybOc71s/MZ3gz5PzckaVDCinAlFOD0p
+DzcsN7Z/yZPTUP592FyGZFtELeHHIrvcXabFUjHL7ss1TW5WNf+rUMGYBNxC9fQ/A4tL/DEuhMf
vfrCWNc/9E1O4ZetHoWF8WXlwE0zIzaboIJl3mCbLhDc3qlQXnulC+ArwRFNGnNxdjtVyGWVJxpN
cPQ9I1GHaPG1PMXcMON2WvMRSgLywzWCe6TKqVTCp6Z1VcUwAhnZHw/0eVPlpYtsfLV/wgZ0vy7i
9+ZZmuWx6rqvZtfZvvjAhdORLzgeFQBVi7yeE/M8KroFlAYjjKhMm/f//ru6IDScUQWedZfT02lb
2pGJyQESHTB0nvBUaGcJs7dmgWu5uisCzcLHqsjPmQb/USNDFBAYSMkcPIwdSpHGNvnYLTryvx3N
xdbx66lIIhAW04M4p1XXjsKD8PfmDa56Ma/v7QaHaDI88pUKF671dHJ7W0U1uPFkd4Cm6A57Z8X2
5IUoMy2wWMqK2U0uU+qS4HgOAix26dyZQ4vVPnneYIUMVnJILAeaALHOxGC1rTY35/eioJh8g6sv
vWZn2AC25oHf6f3igiK+aMkK7Sn1Y+s+2HLkAELEbVDbCesKYi99RdBZ0APEC3TbZ97+LHMeLS4v
QJo+ynGLNxNBnrYfGyPLSfIk3MT7c97qWEwJUA5f6+MB9BBCqL9cB4ObsVXiU1ycJt3c/pEPPVgd
pD+p4A7dylX5NznyU8P1EK1zD2Qo3D/yuuyIRpdkwTxpkW91vjcW12QKd8sjbAgZGw4maqh+Fh9/
eN+OFbkDJ3tQ3vVIfovdw8yk+PiW1Eek1dpxi3sOKiA7K/8Mv6U2Hq5rchJXlgL7TUx5B8nOL21h
VAeXmBTX70tbfGRZyJ9+7hqTFn+1jJiLyKKzdRx7kY5BHgxqPNPwSOQjQSz1XZRgw+8+JO9IFI00
XxwFEhwbSQOYkaBmui+wjArQrr+2z+ufFXQuUpOmfgrNJI1mJ7G5r2C1JMGtVOE4dhINopqHzrM5
DwoIQA5aBshpKviykZzbFDjX7YzB+3/WmuLNVtH7sFtM9Py7asL0ayOKjKM69nPFTGUhSEl/43fw
BhiD8kHWGqT5XUCTu0hZ+MIw5+c7zHTxQrutWzfe6uUwH6Cw2S+XBQCMLMo1+qz+YdHW1ngKxoDA
lvM/p55xPdmEM5eEcniLYovyU2xuhhQSLNqM6IggPuZ2524ZwSWoyiB2qDSvI9x4IIa4T9L2mrWp
SkUoVOhF9VYJlkibF49vonxsT8cOT0edjohn8f6XJ/QIhaG8J2EyKIeJmw78hXOwDQMRVsKsCmjs
PcgogUBNMkOg3kg4OvKNEOcLYAzIMlNbNC6lsSfbRO3VSpOYWUimNA4dvjvVEsF4hncmZBWfDB08
EhGCKW96EW2OcVYoPuByZ2t4ou4koSmesuOvhS0vF8HAHtuTEwGamRAxpjUegluoRuP1x6POCmZ1
Kw8WyZZFoO8h8DVqH7PceCmIcYavGjfD579OCgnymS6BDPraL5nmmNn70iTflTj5Gg4m8H/i6QJI
P591QjWZ0xJ19z7OVgGPfoTkgXEicobnKehU2TL/of9hJ9Q1aTPV2E47GTE8ixH3E4wERlbhzBJO
qN9yUzVw5XzyGGBHg/hc7jiTEnp92EwyEdi/vFeh6UJm+CQGYpH7wIGCXCZiw8F8rX4DjBmgURqc
RE03Wz1X7mDsdDzceynzaruSdNhQhez7pZsvzOSF6vr4FKfC8vde1rYH0xcPfQsKbXzwUiF+44lk
6bLKX+eZZqf6MLgG49jV/cHKTrXw3O/FCe2grGj4fP8DZnPqLH8XBx8wVyXpQGpksDBJON212HP5
S3lHuz2megOiRhELsz8lrruhbjs4f4PC8GX4DrepHhW4WI3q0KX9nh8dTmDJTBpXtZErMhAXx1Kk
3lmsf7Iv8oLwr/YLP9t1v3rZetYN65YidJR87d1sb3EOlqfC91R7Erv4RIVY4UYEWvJBP3zFXD6T
PYtkww4iGxXtyYeKcv7AAOlfnvarZULiFSZgltA1IkUI+6yyh85xbtHCe7pnfo5rnsNknrMATtzk
vVFh7u5JKEw1Hf8NsikKUxFIXardMULdqu6W++NzJJYuGtXwOIeO9mhrjhhi3eUGcqN67RTuw0Kt
17yezkWgTgunZyV1sp1d0eQQwsPrGYgMIWo0IL9mAELVCjwKlgFJxVK1gJQsTdmZOpDP/qbMNPvX
PgmQw7Js5prwkQeUKAPzzORk+GpFrtpTj4iP5CHEJxACgFxJOSuMZtmZbF8NDf1sacinc7l6ic+N
1Hr6wGM3aCFLb5v18XcOf6QmoHox8mPSISPNifV9XpbAAzePENmQsGifex5OSxv1r2htJ7+GPa45
S8p9xHK3tKwa8pgbL1XcpesksiEyX27w7ivFEXuSArPwRnw8aJf+FVth1PLmj+uiQd3Eg1etmmem
xrRctRjcrn+zM+6gsGgq5jlDmJ++Lr0Ouq1pILCnDzEnghvozju9+lAInmShQJHRPpyiyTyWoe/h
JbgHCeu0P6ssxkd7S+jLiSpXNx1YqaylM8nFnBiZlVVRD2x6CqqYh1vAoTIHSdZ/Xm2DVJNgxx84
r3lZ3UFi1rKVqQCKw2vNWpglm570+lZfLf+GfgT3vzbpcmMgKBoUTwQIgloQWLk7HNQzI/Hjf926
rHqtEJf5V+MLRA+j2OTEINQ6fEY7QJegUV3OehEjKr2omhjpLPTS2WHOw0s4Awbumv51z+wDrzi8
VAqJ06opVUPdyiOPcwlypqgopyL9TOtAO9vYkF+7bsD9dpmR0qXS8hXZFK4fWTNLJBPZfHK8n28y
MRJun+2nJqqb3gW+shrFgwjNwCkKIPMvlkAH1JZUM5wNI/BhGTLSjcyEwfZi5CWb+/F3CaWF4eMo
is0zFYsiuy1tj2NDjVRzYgU36ehfVkPlH1Ut9HoOVPpdw49BQ48wpjuIa44BF6FwLQrXW1DXd5Wq
v0c/oY7WaL2/+B83QWylVIVThEsVGQafHxlkrkudY6UDSOr5Ytz2b2rPff5dJAT3BTMxetQe1mBm
E3KZlQxXP0CZbH+yZd3y0GXWpTnZB1pIE6pAqj4fXp7AnylihLiCiDq88tOVjM8OZ5qVZHg+eG4B
IU6ZLhDfvDERKwK9LpjaorQ6diggmiJqndYMyGMpVvdYd5GSYlvvjzTviCS+AIUh4QKiyJdKROXA
uEo4hx6Z7tDpnV1CSFjURX39gTL1YHSXmf822kxV/+UctPHRb5f2vkXEm/CfwLiX2vfClh1D1KY8
0X4mjh58YIxYCv9GD2NU9KUMYYCciWMPMzhollQFZa2ku1kr8A5Tf/jH1HgaPF/y64bC0SlxIajw
wzWlKFrPIJQr+7Y+CIUJpgyivbW+LrtgV4+u+6ujvC8fQARe+Q/dCukzsJytHoFAuaGij3OARLIr
8e5I/R9O5HjH5j4QTj4ZnY7mv5lJuQj1RBvg534ryZem89FQwGs60UV3w5/VxEeh3Rwv/8MNvhP/
UZsFt27oEfQ6ISP6eEh8VPTIo8bZvFEEcLJDSHN2hqwg+YWr0rApkrGfuFzjzUfzXd6veEcVEcCE
IyOgu6vhB7E2KEBW620zyZ94ZxRwe24jGTRSfNhb/6rcPdF4/ApVWX0gsAYcAKiLyF0j1tgN/dNj
siNhBFJzkxdpIQnplEFSEJy3ph0NCn4tlw8AXzKkLSszcgqLW8J9gGkyKXephlT0rrhEq9y5lJsm
BsgM/L2CD5TCXFuyRZKqTeP1C4szPAelaeId38J+Z5nFnTIGkWaRx+83q00EDBRBfF8myj3DyAek
OAC5S3g2fkRWXg7UBvVQ8skK5YgiJu2lkJR1gzNj8RSVdNbX644IqTvtt4Y80lUcIk+mXnW8qKYC
D2V1pGuSgjx2IV1REiJvMEeVBPxA5Xssvu/qrR2IH/lkfocWwHIs9fPD+NvF1qTWIHBRbtpOEt2l
MbLISbAoilcaI0VL/hqgE4D1Sg0wtY8IgvUAydJn8ZwS0ZNOLnkc+gKLDKQaKi5P9hoXXCJhouwJ
cQH/DZLoCCjZdrLXamLDQQBEqKTeYwe999Lkt3I6iiy+zSq0p6zizwXXxSzeIz/dnII8GHyKhrFg
h+U5Naqv5eReUrpBFzCyLsCKBfczeIfAxLTk11ixGG4QAkTirGA6eAue0eF1x735HiBZgao/TZq0
0Zjmkt8T7eoHAw4FrhQr0n7GlgzSH8W6FoggjIgMl72VsNVXN6cZWTLrMu60AZJL57jgnDMkdIdN
YGMfMLbjLu1a0dq/YNnuQRQ1ps2XtVBPOQeg9CHgQkCTgcrd7Ul4LwkGAJMaYQk3efjb7rCxCBoQ
FKHs3uaTiJgucL7FXH0exLZRf8jF8vn9n5ziEPDlJnTrVpb1ziWq3Fob/E9HrbzIYEwfu4ptPifD
qxDJyD/UdGpvraRBsWqDf1/Tnqf6etQruGo2lYGcUpwxKQwpw8UZkEf8VJijbartvlb1E0FLXsYX
IDiHuEXaVmpR8xbqGk5fdOFWCzJGHutnoy/EwLZRZDj7UZ83r8tD+/JJNfjN2zo4stcNwtCE/7ou
4fg2zuHQTryZrwQUdvZmYnVIcDdD4sEhV99cnpDvveQnkDUse6/K4X22f2m2TYhWlKqb+xg0QeN8
CMrJVqElbhY55Jn2rxesVLeOJdmctWV/tFa3d2aSH1W0ZMTEZ93iasdeRniNWzlevXm7Cg1ZlwAF
8HQyqhSihjjcphhxJ9QtVTao0NFysoDrCcVkPX7IpcCxkcX4n7JynUHF9m1bhtb7mZGE4bX/K+Fm
XYkqgfbmGcsG6tOymBLMDjvKO35Agjb5hb7ccuQdGeuhuWYm0h+lxv7u9QAJ6m++BpTcBGScJz0P
bkRYJceyPlTsk7cE1MRH6eAzH3NwF385FRZjHBvfhk/c0SsU2G75Vw1sV1r3CaTUYKvKWrsPRrox
UR7KZk/fN8rtijzLHTHiuWZbLi4AQP6y50pnyf166HhJejzSJ0XqEFnKl5o6BNgibqZe6ptg7i6t
gVRMz42YNM3xXPoapXotQLCHqgBcmNkKhZU31AozXZ9OVxhvnPBBN0D170cHrmVVJNFfQb92FWBV
TK7UlUyjMa3oeEpX+00cCuuvhzgHObIpOxZQIDdF5l704aXpI2TwWxMIehpipgMJi0pEigMFHLZL
F+6sTAzsjzpmFewYiIGmGJfTffoPPDjB8FdfKfQkjze2QvKZB5MRtvx77SlL5g9KypeZmigtz6Yz
DAodz0vEf8ZVOlb/zdA+yeJnSV1pOqermL7UZ2caH+iXJWW78wHuEhTHMOlvBiIlna49h4cQ1Jy5
4Dk4RkIUAmlJOmkaZhq3mUpS8g8F78HObTgjn6aujAABtDmEfI0VmxTD3XAS5lO3DG+bK6kzzEiq
gOTvYz9s6sPfEJVA3hLbUQDgDYXpsiP6ugM43VwMiOZk7u6+LjSVUtCUsQgzlkz8ydshry/GzScd
ygEBCCjX5+44guItfg90DMdSJnskDEMnyL4Q4/i8TyrNctUSLPqqYGSSe7VFu77t7/DV1CiWcWog
q/nCHXggV65jTja9n/sJSKLUbiddhy920ax+EEmmlfAgfJMplluNLDa8X7tpSR7UTFjen82+r7xp
MJpyB1WAaLeFW7T9qQBl2g/BfXwhIXPdhxzHE/McErbYgm59nwNuFAkWgc87tnBVUI6X810kKb/7
8Hqx3HlPbFDX4LMOnZyRMQWwOy3MKOurlH83aEpCoCdsqrdO7Y2VzxkTAEtvgKvCods5oKKMIiZZ
FcxV4kTdEc5a5jBVJj/9ZOl4iJ9O5XU9nIBBk5uskr9KIQs3h1NInRZtm0mWlPWpkbHW4dxce1lR
w5i/3Ke+xfwL3mtwE0Ueg/vypVpX+zepys+HTQ86EQ79jmJxZVoM/LktzsKXqY1gpaWUlEAJVEch
n4dEZSkSDNTXS0BD4ICjpIuMGDm5IE6/EVIAII/3UD0bgu2O0Vi5xoleOIQ43yRXR/i84+/V4smM
3VEUo5x9680Ildzb8fJ1NZTuA/OADZRmmjx3OvFfuPdfGNTMoD9cGDEvcW7H69llZ1kr5aCcXBZS
nC9wPQXYHgKhNIRCr6NzLgzGSx5TLXqMFCjeufzlBTotvXHzA8aMHx+itpKQPFk7Jni3RBi6ozfL
pvAVbs5usHVNWcGKXjpfwYk9XHdKgnM+8KY8v0nvrT9NolZECMmDSx5nX3S62ImByvbkNEJ9CjSX
kCdo2mSCDYOcsy9/LW1EdrRuM1yl71N/RkeGDgR/ScIpL3mW2LQy1JtNpffLls9MWPrEGmkHmlrx
w8blrvfrwc0TPN79BgHPGRaPGRyh6baof9JA2KN9UfFBuSL1Y5NXmIufKjqb5qhzKpn4Iwht/l/o
/7+5SGCPocV4qUMnmxUq0MHX/XlAwrMSDBB/z1IiqKE5G8iIRpsQnxetu5HDiODySp8HtqFDxDfl
kN1HuCgttf91VU6uUJ+ohwgQdeDJ1kn8QmKiDDb0kbmVp24Y/WEx4v7CQtEfhgP04VfjCLNOgQd0
wO3XtBTzlUy2ja1ORtRmWcoxPi5zmLXZh1pGATMOO3+9p1uqz+VoEeXLoAupfIt1zCo44OUjO+fj
dZLNg43XvmiUexxZoAF0CFcAWfp8Tlh0CZzYI5AuHHQdOZ9irP4yyaBDbdBu5ERMToyNLKLUoWk+
jqZnO74DEPAMtBLyldcZ0m9a8HQBe6oWFAlZJswXvRcVw7HJKJmWFF3VaRTUMhr/0cu7x/wOsEGl
QeufjcqBuZ+C3VRUKDyuR95NaCntayS3CkGExgp2cj4mwqyf08Xh1Du/iBqj/MSZJwfngb3Xp6zM
TfO2fc0CnBv02NT4n7ciK02IPkvsoSjbvn7f5GsuT+D3BgQ4AbU+1l9IeFUMlDY6UgdcSUwJ8tOK
ajQ6yBIoLvwXW/3f1THyZn8YLiCXScQPTneMvA46pn5QsndBMio44rUD95LbmCulkZ2KZ9ZncV5z
OqnbxUCfBh0k+GyG/g7FCkUIyabLvG1BCmi4xmb4jvHYRm/9rLdLKYXtxLGmJa9EcAP33nJCw2HQ
6ew8YFcy5IL3yNuuvnGk3JwoJnILZa2p4lU/o0d9T7w5DCJzJcUttEPxRoyu5nX91mzjIQ2KT33B
GDgxpq8dxEhjzMC9jfxpmlriGKJAJJETD5cvjxAn5i4l97z4zuNzm+rnXCFgmIdlAimSvBWtmkNi
eVKudE5ST9zYoqSZYCihrWdCvc5G0QBODGt6Geub/c0N9Z8q7eJc4kjV30EQdLMiOCUA3R+nyPN/
z9g4jg4RDyeNMhVsWx0cHnJ77cKe6WkjYnfWWFmj9E0WEm7J3Mz5H3PWIQBGQp/kYTPMPaiL7wTi
lcKrkn2vT+D99lFYn0TqO1lr+FCp8rbBXFFSy4lhWc3bc0p3MWbig5VJue6/Quqf0p9R1q/tcg1x
yslcA4HVson+QiDPBFmk1VkhXuumiCd0J8XI8EXIyndteyXl2YBMNjq8JtOA35HoGZ4dZxzzBPQx
Ig2vNqlgU4uQBb3nEVMNN6in2FopvUrBgAE5mSHBChicXOD3+M66GMUX4SXXeazinNOXQh4yIJJN
MJUK8jEwM7Y3q38rEGf++OThblqafAlqGoMxlCQE8c8g1I/K+5SDZWSf8E30wNwlhUeb3f8i4RTw
D4ol7uAw4Y4OxfSAa5KBFUnVYM2/CJ3Y0eqfBhYGfZ7UPCjz1ZPo9VCjGSgAsNAXXKTAF/Msn1LM
Trss/FRs+unSEz8KvG8ewrOGUnELwEDwULcb0lINtKEokQCTK5E2aWoR1iHcAlvnHfYUlYnSvlfF
92tZMg15aOMIM8qajOGJtQw0ZSZ7BkvB1XhE70+QTcJbIw6eCOFHPw/4tnmJoAfkEBEEGhCS77fK
h9QLFVwhhRHmLgJC5jEQbljOP/X1lsRk6zhv+3lC1aBlv2MFpq7VsDAsX7YzChG+vQsjF+E5UuOJ
jxMfFkDiNdtFuGj9bISwaD7pHeFRNpgYFE7AFSxQt4xznhqNn/+2UXgy9rMiq0S0afqR9qglXFOx
bCDMJtqEX9zZ6vG72o9b2ZrEKoa/QWENiy/NfUfsRoSc6LnXkopUufByh7AyalNY89G6CVAI/NJr
CQVSGPKV6axDToPGAlxLViZmVx0q0zLp6e/8x2ao0+XPga3F4SqgkKy+mCAUaVjC/JqUxKUG+9ia
mQ0ftSGJOeF1+WDY6y0Sw0b3+iBnWxio3nLFhUAu7CDzI/ZApzsab6WMCzFdMiwqEsQHl1QFPOpp
QYGj9rSpSytQVtlGwLwD/BAOlM+k3FtKCg76RYJ1nCXxJ8NmgI7uPmFcktlwq/7b4fxQYqWiGU9h
nWNR4zM2V0EJVS+GuKbFmA2mNYF7+O7dWKTW6CnFR5crXXC6ofDbck0DqZyqKto8hf0inKncUk6m
5LIzM2s9+ymsemv5hs4hWZDR7sK0g+c7T1+gopNT8TwOz512V00icTBhWYaqu/dSURr0uXLpKR8r
HQj28YuhDBIBVPsUcSZC8wuIXAzKUVtvv4ekteLp3tyi2kiOHUX0Ljk6j05kCxAbR2D4GkIa4PyR
io0ADMCRpmS8rEzA7kfaXrvUWP78r2He+fpIVbsi4PYnKLHJE2YMOahCUJZm4F5q9aLtMx0U9w6o
IDVg218wIdjDt5cxHJq7nWuFysSeKNNQTsLENdMzE7Ysnu4edzZ78ZQ7Dpu/xJKep0goWjy6j3+z
ArRj1lyTAbrbVGWT4pUGU/UH/jhFJTDBXIR00XPFnuBz+WTFtiQi5PUXB7T1wrgrDJFQb/Q1aX6f
1MksSneLY4XMoooVhecsIIcMNCqOfn8jtniEmMas3eWJXrG7elAeZSqTDJpifsbJZQ/u6PmObYdT
dmD7iP/G4xcVpA012tEC5f6EX9YkkM1lbn1Xb66TuYsR4ZNId5LiiHTCNSKano7xtAGQ2twrcY8f
neg8VpC3J46VF4+UcYi0NsWVuQB6zHlQpA3crt4dAGMX7J6MjJTo50TtrY48DNhs8ky7Cqcabvx3
deudAIBaGOBa3rOJ0s1w+TVp1gxS6fkWshkq1g/kbZikP+X8ZpLXS48It1+TJoKeAhArAcl16XG3
DbfQOyZVTYW8ygtUxkzHOih6xZCz7VIHHsGo0XMwP9/vVWiywcYWGZJ9MmCfLv8Z62eRRsLiJMRt
xQXVXYLB5yMzKdXxszmXZ1rgtDtiPYAd2jQWZO3JXWfzD4E03c3D8DmcmpfQ+3gkvlo7Q5HzPcYh
KmwXCoWOYwVRF/0/L6cV+W9Q1Hb1EkvjjE0mSXg1izoHsF50AiNSJXGabeTeirMrwGCRctu7RFJq
22Xtld8aXSBYOjaaq/ak3RnFFGUqsO+NCgqBuHf6+gcY/1f7/E5bU2Sn4m+8tsGhpbTy4BtWohIz
FWOR69k1Kx1esI+AMJ5w1hKLCDm3wcE1PyPAhMcVRUXJ91OKHi+N0t5Z0/gWmMlCdq+gRv9AORNO
gtXtMSstxmO1q5c5mpy5Zy5cTV88+IVZcCC6EW6oWmopBAwVFEOV9yZsH2wMpZm5MASot5Fua6kU
yHcl2+/OS9oOpmaMEZiAP1gcRfryjvLq4FndV34ENattu/3z6ZZ6Kk9/curytFFLRefC3ZJ5p9Md
4JBpPMCaywVOn+21iGF+At7/M27o9nILRQL5B6mzJY2QtWxhddPzZXM8kv5c+LDi7mEg9dmeCvey
FgCWOdAbZ1V08PNSJQT8jXCxO4J4idxdOXmeqbgbfJafv2IXZl8fEbrgepr0PjCGRnLf7chaPjhi
4BSkJshu9MoN+/LDl6kM39v/0eGlraHpcPml7cVkfgwQ120E8fujyNAV5GE9TaW6RU4r3fCX3/8W
t0yzK/Up1cfHmfrYsaFgAhMs8Cra3Kry55pkMkrQrseGpLinnRwkwAZd/JRpdKrZ9/1bgVn5+2MD
5+tKYu/kXsb/iygB2SYrqUZBdn0AhwzNwz4TfajBFVcxJdd43d7BXrX9SG1EqxV4tNLQ1OZ5EmOa
Q79CEyw+XZl63RUw5jrSKi8mw7ce476ZErla2UG5TRXBm11DrrxB8QgUz9324VBeyT5np7yWJMqG
QaHdu5lKrsYMAqvZDsilZxirg4zIBhP0582SlAh2F32oqBNhz26l0QlVNAUZjSqHzmOtk3+KIUnJ
+1xEHpHFLkCI1KMEK6xAO0a92rtzmmLzB+uEatIRwk2ZtKLZok9qbnPlmEz73PbRvQ8DaQrKnH3y
lVWQs+MjyCWWY8GLeGYNolmGTwn4BXWe0BabzmVc0U8ngh1gVSYSndBjZXhJCrOwmtMdunNC/sX4
KgXZtvdA4mASj5eCqeMn9yXFoYcpPvM474YF+EejsCC/KTF3IkFIbyxY6m7aQbIWYcD1AaWffGp5
NTlRClduQXISoPnii53tl6B9floUle6tzl5GO33GOCryYHCYKNqjkjdY8f+WaqHOsoIdYVTey6+b
FRoQ4JJ1FJ5cowesqQYIzPra0NDcPBhyWuCgpSZCM66qttPs0ZeX0oIFuXdviqQiTnEMkU0DccWA
V8mPkM8+c9kvzpUTzjx669vIhkQKjd+absGtY4GKPyyyy+gGaoV/YgniT6XPOQd0Kpor8ah/9W/K
M42DM/42wswoGOxe4pMjV2QQhGpiKVadieNmn6rPti11dJrS9za9YYaYZZ01s5lvjpBYMZbp/TaR
z4sldnhpFHWk3lqE6iuZx1/s13lmhPYGfobKZzYcq5mhI6AQB+li8Mj53E7zAwDWLEcaS86kg5G2
VWz0u7ct5mYXuhAghib21fkaswtMiP7ehviKac2xlnrvbO3o4p7okgU6P3h4sbJGvQ0VIo0VYhWs
UDeuTWKexWOS+tPbpNFC1KlnHlDbluVa1X+wxrPSP38tyf4wxaiGd0yJQUk3/t38QybDPUokur8i
uISSEMzzbl3Jk2PE2BmcKQzBXh+BrXlrBRrlJ50Ko4bPXhvDRN7jZKXf8NBAmnTMPQAyMx8YvrQv
Qi9DJmYB8ErpUXjQZs9m2XcQWtk/XkJn0OZCuwBOCkvt+r6Gq1kdLtwi2RyM2ai0NehU3amqmLmF
OKObCdIMXo5r63hdCfWtzQwCeYK+RgrXhRutieDd/wGlZdlUmy1eCvqcCihRoWvNRrLXA+LH7/Ju
IUQhNrSBlI8dBY0rTnyWvxCSoxy+gWBB8UI5gKoLT2zR4+kmqPPsBzeEjbDxRdGhgKAu6IV5YZfp
8vL9PwQ0ZvWYStZl4Fj0Uw7WoBv8cVo81zDJQL7gJQyjhpyk/ZGI5jA3RG+GI0D2DRSRb4y3nHpk
IWDvyLfEmh7+c80RnAsy2Yysmv3MKqi4XADFJ1JPM7I+dH3Nw6UVgQzL1lvSkvCKc7YayPDLfkN1
RqXptr56QLlTUu69GlKN395EAe2gSwxjz37c7yKqhku/SLiV1VyTJmJrOa3dKB51HBHfTFxh9D3P
stv1ss3p9YC6F/ZHy8h50Fl/KAMupx/76RLflE/dDMFE+BNb987VVrRAoeGUrIivg8RSjm2q9fKS
qoaw3GekItezPF53delYxpwyS4CKOXbXoHwMcVPfwK1J3yE+XvwkGyHpzNyqwT+dsZZ8jUBGzquA
O9pmnjH/jJIdssD4HBBrydIYDQaQ4oX4R+OE2zYu1qL6ZU2Nq1kxN5arcgVj1yn9KM8l/JTUKLS7
O+M3aUZz9KokhrSEilr9N5mJaE0fuIhjEkGGe6hsZEOasqs0nQ3rEHcOfeUNL6RV5ir6g+f4wJkg
8qaLVk0TBxrFOisVdIgggPzHaAJrMM21Ni3Sww1z+Ha2lc5uruRcxrcycRDretmk94tWbMALFzV7
5FLUdcYMo7vIWd1LijJja0oXbwRq4M0rOSb3DHpRlCaYaPt3ZLuNMZTvITQ+BieXGA2ZSGSUV7fU
cGHiIWutgb7nQgSdxyYMqSkj5AtcqUoFd7KmSpFiKt91j2CdlBzXk9PM5cC0aQJ46iKYe8WTKz4X
4Ee4zugxUb3HJmG3JKG+X5L/pgA/2ODvm3qp07CJ7655H/TSMMduha9hrvzXtSa5PJxd/axs0rpk
jj5HficE8fk3LimJjU+JBL7CkH0JWZZz5TTP+scb0gWO0hlzk7LEsL/9Zsa68lEOxmpoCyJrOhyF
7Jw1geN8VSxCJS1nQ9r/wVX9kmACF+LTNwk/WBG1cbZEtjaM6galnfkpB9ZL1juHFt6ec36XrR/y
YZiGKp/UoteurJhC053gT1gVcJDNnRtU5HJe5VS5rb0ORDVNoqpfUEioZ8v5AEsGlbYUcyPdsKYu
c4oiRpvC7RFFNieUPC/EZGTrVvRT9YzJ0dzT8cNamrJpIMHXmKwUIxHS0pBeT0UJr1jwZp9KuMHX
Y4CoNrAbtu76RKtMHBBl/+y2gJhHhRMo9hJE/mYI+om1VLK5hd0Uv33C30LUHMrrnavMZh7GKjKg
8Q/0zcLAdr81Wy2iHIwzex0IF8hv6V7OcljBmngS3EhLcOH2DKklryufLYqmUS4xxeddp/WRugha
j2VAYZUAWHrlqRtDha0P1dNs6lkYs8IbwtIdTYkaUovHmx43G335BurhUpJb4w0VnkQqomyLBP+f
lu5t2H1xgB92OBBcCcxOVCayFpqRB5XE1tfoGUgf/Ceh0qvS4WoENivzAHu17sZckoqPbacoYRJK
JDtvG2+/LkYLFnK+/gFqvRq1/6B3pZHUw6HeTRyP7RoAy/BFOmctv3QmsO0Sw6CC/DRxakRlytZ9
bekGMAmSaATZC7JMsZGK55stbwIMcX+XmE4Z6I2blsOZxc2Nwxtx788QyVNYZjfqZ80ouKU6RC/O
WhLNHD4XvkDY2BbmavE7cZjXQ/v1DFCEJrQ7f9IXh4V4iYHmbf7RF0UXU0UZY6Y8z8RUIAwKG58B
08Igmsiag4X+Rd9IGtkTINyKDWQYPQJYYuKPOR0ywVt/AiJ0h2FTPBVcMnhfoug3Rb5X/hk3Eopz
QB6sDnfb/KbFOJPXybZgPbQqdGR48L50peyHuwsK06ACOSEKAT36/hbfFm2hX4XtpdS9VOptinSs
28zNVOQo7Jy3TIuookTrNcXQe/giqDtob+HwqGRiWvp2Z45PMQp0sBrFW2+XKUJZzpV9Xtd9n9hc
Crub1HbcgNalw2TNVAgXaiMUJ8p6LQ5rsePsAbD3hvvYzadRHp1Py/5tMM79NtkL6zcOX6KNLIqs
cveTZyLCZNuFJFdrqHRrMtTkGl9o2pc5T4Tnvg1cFY2AnmXur4BvOErwdOgr/79Kn/lxug3mdpa/
IrI80YinMgCg8zGSXBRd7XqXnFE/6mvlDUj5QG6EIQdjG4gAIfalTkpNnW+JRNPmoU5OeuuFz35o
R/mS7tndlbrg4GWirdLUDXD1XQptrx+TmHOsneJZjstyV626jyAKsU7pGOxPvWbYWuTK6p+wzPX0
9FX37/J9i+XPgcy1WL722uDCsstEqnMgQA2lbY6WdbXN95iV9OjietzOVzLmSrhx2+QAjJxPXErV
759tfFfQKqBpjjB6i+/PNkQe2ZqhNUh+7Ub5V4pjpEj0TkOQDQ2G66J8BGIb+M3zR09jNDhbUA2a
KpxH031cfuGzWK/DSJD1mSK+ZZruxjTZll2GSHiiEgNZbeel30IY47PJR7glEdoYepf9iFfacRur
pE3viYL6PTH/Y2h9nWmH85D897EtSU6JDabdq7CUzoJyFhNtSD5iAHuhGZcvm1neZhYycI7iZot3
pslZ3U52pRUj6pWQRqNH+eBHb82GhonlQlpWvkXWF0xxcnxFXS8MAydtFVxfF8D8vRhX74mOwTPo
jBOZJEO9B3NDQknk/qgX9fGqiDvfbCCHiGdLG4NbbnFLghvmNO1FuqDuVzKEeghowY7837hUhvMX
nJG6r34LJ7ueWM3z5ul169D7ulwqIuVp+BT4CG46MgGfZ6owPrbYSz396G1sJgwgqJU6HG8fsQEe
9QxFpjoPqpMErFIw9D0x9t4be/z1W0EI1RMJe/Q+EoqLxzL+eUvCUlSWUjqn8meDoTs3pGqgm3EX
E1d6rqVcju0UTDDp58cqJTgWKrULkv9XDqwo1RZ2Uod+em+M+XPvboT936/SUo4MToLAP3Bn/AAj
E3Xj3/UY0LzZuPJoHJopq/0Sa7jgsGqZnqbpR1//KteXZxz+NDFMn9dH9d/Xh7uzI3XrJrpCBHGJ
YjglfB0Q2jSGS/eIK0AuGTrP+X5vsW/9k8Q+6Ki/kEog5yYu8gGySjvhtGURLqoLY6ff6jlP51D3
W5O9OxW+hUBxl0v7yDaFdtJhJssZ4v597W7pupV8PnIQ8DY48bo9+13+J/jyKjaFIFckG8Kek94r
0IXZDd+BpzGnCNf7Oq7zGJek5wLl58eQm0h1l4EFz2J1lyOggbIFS1YxtJS8NOfvve4hKI4dpkIg
vMn5DEisDnZD7w7pV2CGA6u1eqKr5lbbgHBeXhZ6Yj3f3g2bOvAZWAUP7WADbrUUE6ulz3UH5Oj6
tkCtSIm6A9h9qUjuNBwJMgl7M4QS88HyCPCu9353vZFrbAlw1Q99PO5rQ+oUIuo3TYBAfzUxhCrA
TsxqO6ht0f6CvnnD0GH0LeC89gUV9hFU6SzrvQOJU+6kzEbens1GFN2bo8O+0XxhHBO21z6jFCU2
zH4PFP0SZzyKxUbhdoq+Ce2KceILjjB8vkZ1fMEwYA0jev9EyfkC64YeRK2IIEte4JCddbBx+36e
bXE7kzIC4gSjz/MQw6X1BqyUyRhXEoVf7kU9YBU4PM4lC0Hd3MOKHz6bkThZjb1DZD6HQAteqox1
l8fvsoxwPTooPbHaaO24UsGyizuGEkk0EzYx9AngCl49zL//t3dlI+aDlUE6vx6wdRZaa+pjhJXc
eoRz1df5pGAxPwme0acbgb2a2JrFR6UR/EypKO+vQyl6Q+xuVG3PmK+i3eBgmwKPOYg/ByZfhaTZ
U9i9hzM5ph3G8Hw+BEcrjuxEb609ppcO44cxz4o7FEFCKZSI8dWpBpxQPRXCsiHty3guudlygjJf
U6WMwIRMu8nGxoPjrKRHy4/1DNxh/HqD1Dc7+v91tnYK5fNlp1kNqp5xy4yANyGncAuf2neyc/1G
dA15MjbiYqXbV9xhfWlDwOscVogffk/7m5ztx6oPx6s3hU+zGhipT1HdsWAk6HvJFvntFDK8agAp
W7h0XoPtEBqjR28JlkwgrqzpdWt2Uf+hX6OEEmRytnbTOH5Jw5oEtmFQ3Om7R5Szq1egmiXnPQoX
UwMN1T+8omlVG+LX9zFLfhGMcXoKuRbRv0cfsHwo1sV5SaIBMeZQwwh42Ke5yDe4Nhte4PMSBpC1
uD48hpYHksPzM+zb8LM1FeQP6hM/+ZRLQyn8DoDuFaZ17np0FgyVowRqIjiFNVcOB+6OESjcBDn+
qQuw+WULqhSm8+slehx1tOxCe3L7SQD2eXjYS3zeoDs4TFDnI9zwEenGmAtJW1L+p1mRlLlqOSNt
T6Ui82ZHS8bRI5W08ajjX8iDtNLFnK8La2hpV7NvpZbygM2dLZ5cf8LfiPS2C+FI4oAXlZkw4QFK
/5lvJSvuyuVxrAdCrWudwTwXtJVmEhxKPNsmhsKrwzibJ4rmAdOZXmA6mdO3yxaJ9c4mb/bt23V8
F7G/piC0pKkovly73brXijWyNCMjq/iDG9Pw2AX1IDdO5gVISu15cp8N4H4rSRrSuN4W4g3YZIT8
lPPfkENzik013raQsOBimYr4rXA9TeMCIqIzknqDc4mvV/FiqpsepizPY01A6Ap2mbSMEqZJMktH
YLr/na2lwHvcq6kXEBshv5wBQ81hzFoHDvhlDMqgU3Q6J4xemeo/N23CUmvcQ4QtZ6g2VIY0gYCW
+tPGdeSpAeiG7oh++4mMZ++ROdt+QDF+Ky7mGeePh5ds+qaj/jG52+74gkitaP52Ez+KRI+DNdYg
muCMxBe3Yx40ol2FcgW/e9RN79rmwsq7jXdrmc1wwhfPFdcjFEicBA+PHnICpSUYSH/rvOWObC9e
gMkqKkWkc1YLb5TSbQ45OBA4lBS/U10xTUm76ooVhrkA0Ypv4vneVqDgGS3j+zPLBCzx+x0Ul8sZ
LR3bOjc/ilAxhROrl07npGhyDVUfZruTS2xc3fS6iuWAO3siC6RaQ/MtL7BWDHR+b3KS4XxT8hhn
7PKuL38gtzwXQGJAcSp6aoVE3DavnQPwzshAoB/0phoZENkQtOJPmOoAjS1MADuC657xXM/9tzOQ
2bpJf6W5NOE4qEUdymwsIhE5D/rkI/4hXzgFF0Gt00PhlDG7WKnQKacqkqbKlH8KMEwVGFaplywl
lGZEAaHASym1M40TwkPWFAjOn8ep0c6dlCXC3FpbUoAH9zdyV+m/DSxCt1AsT9uZKc4QUMhXd43t
TOgqRZGQZsB0Y6JWwckom/nEdwr73q2fhVMq4YZ1LWTyR+yf/f84i5a8VfGgnFH4o+d+D1hyCGdV
ypyFbmigeiHjoEvz6TmkWEZ8bYHCXmbAXfp3pVIJ8ZoQvAFTuAFsP+GiZ3xetqH+ESsDo0u9IgsE
Uz3FO71J6DUOCgznuwBXi1DK5kDbhJbUX6c1H15l9+5qYJuNJ15BoFwLjTEnJ++W3p2hGq+edyGu
zsyoPn/uErBBSDpnPjZ7dOi9zqFFAZNZylwYk0WjHqEo4W/k+wfyRQcv9EZinRPEZXVhv0CSgQ0t
LJpN0PbQDb33Yy0+fhKQuVuSPEDxbd/V/SQFcAvoOnBXn682WL0FeqEQKH2BowuGJyVSVzazyhwG
ukEVYet12uR5iVFCPIIi+KS0xlYlSd3rmzGfGXXyfAEwZapl1A1Rxt4lIGXyQpAO4BCxW/MDqOhA
kO0+Cz2EQqhZu8Ew+vAhcyNy15pGd+waR2Jr2R3mj4xjHwNMBa6gtwTR+VRsBdx0KXXvc0WDyCTt
T6zom/31uXxHEFCV0tcVt5f3mD0YkiNjNwAa4PlNNPxvprQMt+H+4kR9hnqWrI2MLn27HWicDrF0
koenNucJyl5gjIE4LrEqvXw0Eh99RBlEG3nHteTLKNn62/TSc9fHies/hwlVGymZhBpR5Dm0yL5/
kHeYbRjFlPN5kTkU2rShJ5OR/PFIu1yP478VrmI9QbU1rB1wDY7vVnNehArG8l8hDMx626kuw+Rt
BtiNA5qqLKYgZrWvgnX6IpuhgO2moU4NH1U5VqB3RD++BeCz1HK5iMMVs5XIDhllDjqdK+5tQ4hF
Mb3JHU7sACFqIbB2B9kbbc7cjIDmdoZG1Pru4JEDYQWwqJE4ngEp7ZSS0GDBec3xqDOJFEsT9K7W
7u5IuIku3myuDRVEzc2bKa0enut35XMT45nXtdrhZz8y4xtOg2XY+fzx1W4IH0gZ5/c7GvG6B90s
GQi0wj3NQz34yla8oTH2hbwFBnNiiossZD2ANDAUXgNLnOHD5aKKgXajs4kVijq9Fms/AMl4t2Zo
CMZTGgzqqo9aYf8VMrgEipvlcRRaAT42eLpBnxuqtd+DNq8xDPhnWfArD6udLATpRhsjabR/0RJ7
2zb1kvyAIXh7DyAv4X55PXbGACyj+zWuLrDkumHJCNSQH8hz2yHktGSBqXl7B6VVzUagvMuoN46v
YVQf82oyI/f4lrD+evlTIseOLRVWmNa2uF9u2AwbU6Vd/7+MUgtag4RUeRKra2YAEBSdxyhAs5Au
NgDnhaCG1ycD5XsjXCdY/bqrUaLG9eL17kCKgpqNGyrvnDTwXrZo4xbBZ4yfB00DYQ23zBbn+zCT
QoyhF6q5ANsL9Pn56p4v5hzUtJE3QbDXvfJFKvsgsUgZscl1arlaPw/IEQVG00HpTETpDYJXTLkY
PYHTHpatN7pnR0eYEqhBMUZbpKgdrMcGvROMlJe6vqAXUOEc/FeSnKBs6/a2NgaVwd+oSahuWXaU
JV046AzrtEHX3speYIQzC0TRzFfDiAsQXqBLa/VzLCgmM+Z2CCdP4W0hepEVFEXBXpVepgYT6Bef
79KRKsrHe1XWY7dt4fDXYwNuYWwPxfeRGk1MPbr/a93tsQy1Cl4JN+YH8g56QN7asevYtDYyJXfA
2BlaLDxL4C5moYETiFEJUaa/3hTMT0uWCFS8b+64msF+lgrn+PtQ//W9+5F1kLJSCX1FB2r4FH6q
c11fVe+DX3VWJYmFUFm0ySCmFEfT7Y6yW6tWM1FK3auTyqKwf5nqlURnaLrQMYJ84iM9EVcdRYjc
ga0dhF98b0AwHaQLeTuaQl/9JlSE8YbuIhJeTT+YPooeu5K6C6Jbskpr6g7gnydpfnH5rLVSuK4/
eFOu/yP28TMNrbdNwcJFIc6iosX8Je1XI5S1eRUSrCJvWFJVpAL+NGz4hgaKtWLCSqkUAjONFgwV
8sAU6WIXucYh0tWg1OgUm7VbKMgLV+/aS/lVMa5RH6YIrLweZqJWY5i7PqaahQOSAEUlzxdqK7+9
KObmwyqSeC4IaVoYHWxMdhUK+tlhnK0MYm7FTR/rBfQ5zaMFf+Dp4fJ8m6I2gbPnKqnlHZ4GyeI+
qGc9EKza42fU/L0z5w9S3nI9pJOWXJpR9dGWFA0dpOpJau/pVzO984gq1tVqDG4a5cT6rMaBf8Pm
i9mOvEchZiu1aR693EJe4FQB+QYJQwtVMAxQFjhXrW7FpmpFzYkfddd64M9LFodtB8eIlDS0o/hu
Rt0HYMQyduaMLd27pSoiUicmOzfn3+V6FhOTHmP3P6YM7zgd8rMWo5OJTROa7R0lsQa9FD+y6Ni1
SHs4kxq7pITK7dfzWkUaB36wuw7WzHQ5tHCyzIw08RbUES8eyMQIxxmc+RAcqo0x08uQEubTu1lK
qROGeD8RoXB+iC7BihtCKb+viUDWirAKVCBtnuKoJu+I8aPG79hkipNJ94Oiy+qeYBz+LBWM/xS+
V3Z40nQUV3E8Ao02uhUiQP1wguZS0arELwX/3BbDLjNAEqq1/fVF3M3jhePo37RFTKxxKRq88bE2
A33GLOk75ZlEe1Q9qARSzOA/Mf86P1CUVBzTlUPnT4JXKTmL2zP5AP5FUJ3rZm6WoJtLxlhiM03h
x7CiV1EEz2eG61oXyz6gCukJ8HQDI+mVqsjIMFWFBQsI/hsO3EIywfBoCcsUO3rZJKD+kIiHWYhu
2cv+uRaRZdUznpuhvXy3w5cPmpPY7vLTqAJJaA8FP129SVjJpl9GQFfqD48Ft/wRSqhNsqS0dBB4
DlbRstW+pQqwoDhWAOtPIElmvYfY1Ro/vn/owac+UciZeQ6IHVldxAkcNkB9xv/40KnWTq6Gf2Kp
mR0ETcfAcPfEQXCO3F7sfFeLnjPg0Gjm9zP8cM2gRnSlaggyp2cjGl9KcEbd1KSWAr40Iyq4LQNC
Ct9dYTQ/eayBxJjKltCWx8Mxo4lK7TTeijwlIHKCeHQgpTX29W85hVW/VajRhHBmaxcLzOLnNgqd
y2EqhHRGmuIA7b6LRt3XKd46kEaN81aCVbMD0uPTfquOxQhDaUhL5KYjtvPdOixBEhZMOP2Se90F
IQXxcPkeR/Ym3BcTlcoRKVe+OCyx7ZjtrVixwBkIrueXmtMRawjJ8fT6OvqCublmt8Qflh05f6TT
2mNG5M62XrxVD5FRZ0vPa54YiAYNZZcHJzXbKsL9CiGM1qQZ8HGh3gwbbO+Aig+IE4oziHj8R1Yq
F6z6N53l1FAFfDin9PTSk72H7knxNghq038SqrqIDkHDhZLGoJyQS4yJhQd37dDhbgezkY8IeMH8
6clx+yTsU44gy0Sr9h1kZPcfRVOEnBKUMWanXmDHcSLyxT6+DrUx4z8XgyECta/Gxk/8qjJVwtS1
010hAJLwt9PfNudTYB3euotAAzrUpRskbLv0dlSu/UAozHnojkhvjXg83A012T6h32NxJ92I/EHl
bhMeqyMLholjA1UuzlKrx161HETWHHKst88EPevXE3/jCELYvipozUh0ZPdiIBja/oKdjGD9TxGb
qHUWOvvKj/wF2vrLvwAYJgPppe2ssCbdRYCwdF7qsxtxMXjBytsSDDXeCLcVnp2477El5hWh/OW5
ZnpWweh7snYouLNeN0jl1TlfHmoTM7/fqzd+lBF3mZA2lqtsofnm9sDpoFBxPqB/mygSAF+Xr2kw
WSdXf8NVdJd36dOi0hloCpCOMwI9COZ36S1JMwv5AeRsJ7BPNBmryHC0yImtAX9KgdDiFlyPcvS3
OVAB3I30RBeSOlbdJrcWXUi/VBkQWmGAgxHiyQjewIA5Xn6TlDAIFz9GMUBazJrHjXE4Fk3K5rOW
d044a5ZBqIFlX6piWBGLJJ6IH1/5iGhnzNolzvrBdaAjfXx9zOw2cTFg1TE5XyK5+HCMVvg92VxQ
ggKcHaUPpBvtiAg8JvoSqLiGOyey+lN8//3mm76jWFiD32MDxVVmXP/6f2arteHgQ5Ojnmo4rYon
xPKRB02AZhdAiLA1nd/OlDg94iVpdGlag4PCzNFsS1Zkh71tZktU9B517tZCB8r91x7KqmQc5uYF
dAOVKFITqcN5gSE72OR46GjkjTfSq7G1GBGuHTf8nwPVlBdWmciB/n4tQ7InKWV5voeD3xEeOGu0
ckE/c/vYg8pjHrdgy96Dyeiiw8mUAFnRY4JJ7XcZBzFUx2ZAcPTiQdA0ZOmdq7DHE4T1LMAzcPMU
XX0jyMV19/jmKqd236OlnVlTYlG5Nlca35hMEAMss7idwK/qswF/IfMLFJ7vzhAUZ7IPNTIO4vm5
Wd7YgF4ZplvmxKhb7jOtx2RmYRbQUbiZSEWrr0+vOXEIhsqPHS5zzQJbI/XmJRhkT1+mnmKRrVKY
xJzN6H9uAbci7IEYVLrA4p+Nk5YkhFnAr+lHYbrY4WT44cYTw1Cqzi4WbE2bSzLITJ42De7+QnHE
UCFXnTbEv5IOacV3rPngj2v7Bx6ulKaFW058e0ioAN/YyKwDSP8J/VspGrn2eMxtZ8XARpj1n9ml
s8mhwKHA3I/R338KySB8V9Zi7dO7FRKB+gyrhRUoCNYND96JOYTmWpQp6yl1R3AC5tmqJBBGVcG/
TbtfVcebJLJD4HOr4XwTtY1Lw+FK37BDWHHdTEQenp5S5zCRZLscNRxN8AArR4MTEes70bT8/ZfP
4Ox/5vG6tnNPR9XsKg2SYwrbC74r1vrOmkAo47Xl+D8U92t6BjpV7S2j4Y8s8IxvtWQ6m8hfQv9m
pGBuIyXJuZNV5p+CNK/qUbqZZyh35P4dBHs2pEUr0NBtsHuky4d7lv52uZWf/4S/TvOXkHIROWrm
FuA51MqRSYtbH12YiaZCcHuOlE6q3JcVKkFPH3s7RfqOIbk7291KO/pVZR+fPB8nO+Vga4fGIN11
4PHvpZmMfuhczzw+Dw/CjpNSVdV2MV3FIV0+k1bCLVCl5jeg6Qm0BAqfD8Qg2CXhDLr1KmDRijHv
oabht+NTahmghto0M74E7p3h9a1JjHGXqRP29T/RJ+gwijBxakRSiyUuA14dlb3dm6wu65fEZqhT
Yv086QeVaiwRKogUtUC+104WNBV6/Z/MkHdG6vBHoLkEN4ZOhU6QxE+prWyx9zppQxoYVMMMhAai
nA1iBPBtvROrO2u64+i8jcngyBzEywdCzzsP/frahnZme6BSc3qu1qasvF6ghGjqSg6ladFhe0Xn
LsuL5k8yLkjQzgJ831UnYbPLWzm1q5w90xKGT8Nim6MsqJnChOuh2dL5ZSeJvYjkKcV1/AKOYleh
4dFD9KmQw+LLJ04p48uswi+gSwSzImaVbXnILP85UY1iw+cF3rKha3fuCege2e/fRyK2DMW64hIO
05zf8/S+pN37nEx9/1bLp7OfOoMFc/QMGQNrSrvy8WD8HKtopmTs98XCeqDRC87kSPfg/U/5w6zR
2VnuCPh2LDTlnZ6c7xvhv9ZvCab6hzjNbW2XLT+gXKNeufLyKeyGk3a/RFHAUHPdw0eJqKxNJ7PP
RWQ/poMiEdQIWd/64yvk+hl7N7O14Wv+hlGM6Cb/SKpFdEBHR7F7CKQn1mMrF5Hm6dix6MAU6tvt
eMo9+zAMXlzs6NgUfYSqXfeScfWqZNCaFjeTpPpCd0b+fZ8fZU7AHWLlQvKaN5mnlRccrDVKpiMB
h4IXQgqLM5frHIpASO2VU8XH9LgMJJ7ZXEihpTFwK0Amc/R45PtNp1masg5zty4ri9Ohjvxw1/ez
3ul6Z3nTkHRYdOW9y2g/4sUF1GEW6pwuHa83wkE9LlMsNg/SuyHUghKwnnD1711BZ4l3QBJNoq/h
L5FnfOJeaiUZ+tppfCNlvKvmZ9pRdYUhytc26+Ons+hjMDXHPDKFvVlukyBcb3yW5ZvUXqVxPkpO
6DXGJn4aH3JGy6IsimtNE53tkTVDYLpjgwnhsL3pSt3yokBueUe2JE74KxrurpTDQlPoiRiZZqxF
BuQfc/FyVxA/85ru+4eYYp4TNGZQ7o4E9WWsWQWCotcecIwA/3lMuyKMS5Q2u0pOSaYrB3Lqrqmn
OKbu+rU1h7e/wr1hewm7mzA4nxUsMvQeGYyL+7PBSB/Vw4vkPKwZ69rEKnq359P5hH/wqSlzoXih
fFgrVUi/511qqQDXULKoBVF4x4lyFW6uqustyHjd8fojuHEUIloEGmuq6Mu8ezy3Jyfr5LK5KIpT
X/+prqAeJd1puqPaY+SiX1BhyzHFSfPVtTWKIr9tgRZnY0J0ejALdhMsri9M7RJ9EwMFD3lsvBti
7PzlsULQG1KZu9qChf8ynscA7ErvxIO1aeyAMjaBUcUYXvsIxCAlN44RpWZ9Tr6fMamuttGyieiw
Tar8oo3S5yxwmPOjIrtLuvYOIMLgoiGmVRyKVkLwYgkt1z4HsdhQTkS0RSDMlVx9I0uhS9o2aeAa
L5aj3t4GCg0cq871F8oBacttU0KQVCSokIx7qTzYW9jQqWVaSCBwD0s6Mi5w7WYLtAMEvZc1HGra
xONRYDUdusimOj0ywb7nFdAKvGpvc4NqwtqcjFDSXqI1FIq2khcx5HYYKpAI2+GmZ5WuONrUyN5K
g9iQK6uhZtR74Tr0lcuaUc9Jnj5oXI5CW75KrjVjmJEibdqbr+8XXcq5P7yIwTdIeDjw4kQAuye+
amHEd6fqvU9VdJP2TMp73aH3ZgnidP2b0oD0t06gpq5/Lp07DWn85R1725WPhwGvCxHJmV0BC/d9
g7dR7243XgY3opusWaIXw+LrZ4ZlObHzFCsK05m4rv0GGPz8OhzSi8wdTN/oIgDQ1nGrD28ZmP60
uTbTtILJrnLOATACdkSYB5vfaVV7+VV3y5YIgnVSlVSjY597UtK/gZzfiKT5IrMpwTQ2/ooUxRwF
cinEAEiQp2mItMvRGNO6j08o780vfvL9EhMHjHhYYohiziiiYrorJJs9dcW5IV44oppd1joXe1u/
cQqUu/7aPG9B+WDT37fX7J798HH+yujICASI0usoNCbhhjbpQpHzUXfiNEqPCZohgib5HqM42YW+
vwkOLh1miqzJPmgWRVWsnM2PJpvPOzPoB4N5wHzlCETYkeToXtX9ru91B48T7727djGB5ixSJD70
/5PK9E/Xk263yU91pcXHucRhpIPMcBzXlUBnPcg/MHtfm3RolMtcOZrQr9tXO83jzPz7mFuywxPt
cbVYwn4i5CxprcX460j8oMtwReaCnOS8ie47+7/FUJVbcBJ/yxPWMZVnmqtKVI196bRmVQjyMOLl
Iq+dPUe8g5NKSozWQzajii36FeWvUnuc3iEIvvV9EB3ELTr61s2yQJQMMSOwo/Xy7VrCDA/siILG
QegObNYRoLDhtwl98/Sg6rlxVAd4OMT2PcJAKr6PW2PejZlGr70CVMBvROjBJSO6fgOwlgkE/h5f
ZoTEWCsAaB4Bxoa2kG2uZEbSbLXe2h2LWaepc25jU8+ymMJcqlGlStzl7dx/qQEvSreSw0/ii4U5
u5ifxht4eHh8JYyVcu/i0KGcrQSt2v+TSWtCAIieZzyiNY509GViwLUR19Yj9mlZwS2yNnNeNOzd
GMfy15uZ5mmJ9Mn4Olvi7kGYvsKiiRjacIraU03Q/X6IuNByFqiL+4nF7L3v3yFuiN02/nSdZZur
LVo/KCVLugH01zMQvfie3hhRozTivttlc5NE2kr/lkkhEp6LWmVbq8oBxl2ZV0tDQ3tqxW/XjiwN
qiUp/KgmZCqIsbZI4+u1MV0hXBttWP4YHFxmsbRlO3yScBVCigHcpBESEpfOhFHoZdK01z2CGHnd
0mQiYnAEv4bSsMb9dgkMjMlgARinDUK6YHQl3/wOSK7O5f61Q1r20ChjhddqKKxp2Z36JQ/Iqv/s
l9znbJG3SZipw2fbbsusKs9oFZR8pSFyr3jh/yUIavZRuUAuuvs4GFJbSn3GjitqhN6kCThWMz2R
+BXrvEYvpuJZ9Q+Gy8y/8QjzqGX+4YapTWoJLOpnnXV5HrgNQtdn/7fSNL95ATHC+EMsKAo1PtJr
xfDJbp0kbCMOML5Mg3ZLzttIIIG/tUiZ6Ld4bpWPHry3KqZANzW26zL1aq7hYuPfiV8gBnwgE2ql
YCwtUSR+6Fox8dc0Jls8AgGfSMzxkEspilZc6IDCadyl4i5OI2t1eY8l06qOvFaA9+gSWnhcdQ8e
HXGZWgNVolKOfYZHlUL/WjsSZ/Fj1oWNkIQprV36uTxK0cbX/yGrNIeX4mjt1VZQmPYQFI/SjH0g
tUAPQAHnhRfSupKZGaWmoLeN4dLIVAvea/MtaQpPX8KtI1FjIOtDdwvLZcpgzpFJaLpRdsBOQQn1
HTS38etmuKWwyn1hMvIqyG0d2snAudbAw6KyyxaYHujAhDKps/GBBDSbWki56VloV8J4iPtWobyy
g626ax0qGx5OS/FBp5qwE/m7GkEDX2TUuQzUFzxL5o8oAvJm0+x/fRBhnQSoK5Gbd+1ww1PwvAI1
zVm43h/f172IvgwA/+qgh0/EUAf+VVE8lhb7UTPAiZ2GiNW+pvCE8HgeLkbAQuxfr120GOWeO2k8
yP8Qgl4kmVUMOZJEU7Y4RHVWRouflLBdu+FquU+SGOm7aYwoGXSWqYCF3oGoBGIz5CmNEXCr/Mnu
jA43o1TRCT+3aCzebMFYF1QjYZD3I/rnTOVVLUWnwf2vQm3yFsGz+sx/E1tyQ21G1YhJRgK4ZiM1
640T1UPfC44wlH2zpJgKO89HIkM80TbkyAM7/psnOpscTQ5WOVHXzIsGPEUjC7xSHkJqvZW9ZvSw
5SMDh2mscakyIKd/3aepuaCg5qwIFp7kL1ybvW5U3W8r8E9/UDSpgngbWZuwpifE1uaAeHqZmeiG
D0rv2kQ6dU3UfXuqHYJcLrFq5HpdsidMFNJfbQWtM61xvl0r5AxWXft/3s3rjA2c3IDCjcnKTsVQ
rihjGSAweSvysvGkbnqQvRb8rSGwpXhwpAKe09JTj7kmg7+oouuDtMy/qrJLG6sTl4WXljmFRdVC
N19L4ocvmIw5EgExq4gJLQrNR36JTlcznLhKzNrBdjZOXCJ1NMcGOUG0Tyq9XEjshOm6HZgMs6qs
frG8ypaVnIdMnuufeWQgaz4hhYRPMX+pkswtrVS6nzGTCo9YIH/5yaKCmDgzSYjc9iq9u93MryNE
CuO8/cWIDTCkkauX969lur/z7qzRAQ1xBSByJlUjE2/69Ab5Sq+g8MvNnpgKgGj5+Nk6oo+cliq7
bvwtgZLJoPrdpGftXHqsHN3tXuIc4ySj3Cs3ROZv/GYeXENRQQbVxMEE21/CXuGwqpl2/4Sd6i4b
AG3bcouJTK7aKg+oX/gWSiBi9a4gqL03l4l2bNhqs5luNWwYf6OdWJbYyFDQjtRSXDKMcVR+8BH4
kSHenrVTZF5eElYPYwmwsjeBWtVI7QCDGKo0ikDhmuu+ewrTjHutPzsS2wfmPS2PgWXzASIM13Dt
mX3GO2xxc12AWuijlUm+N58uBzflOukt97citqXT24x+3/Ke64aqAzslUw3e1rmH7FQLyzaNTdX9
SSQ5AFoPgG1fi/PVcD05A/YxLyZM9Yzh3s15ohOd8Bsw7Ii2IuGYHgJMX48SYUixTA3Jet2WWLfr
5bXMb8DgzKt2CWLEpSQaZrOKlYJM1ehcw6tCVq7KdH6T3CxkfDR8Hy6w1vvi2HyejybqTj18UGAs
KG2jzksz8pgEGinObYENQMhMXN/FkngOj+yO+kNjjZCkONEFeZ4mmhCVGoK26g0XUD7QiY6qnDjr
0ReCpxUNsp5GevOcv2oZ9E3NHhhl6QXILXZffTZt/aewN6UVNw+5bCTnyKt61grhG/v4j/nC0Nh0
6WMnBJfSXQZgFWcHwa/+vXV0Hd8bYyKhZsZxYOoaOfwKoqm83dbXXT2i1pnfBbpMgqyi0+Rku5Sp
kDhi7PtqaOqM1mxzOD5D1hRfBaAvynyjJvuRKAp/Ae+RXsnbDP7lkXkEMKaYD57OE5WoFfWsbzmt
Mt9odeuXIkNRwj2YZsMa8dbwFMcU9KqA3QM9/zOhgMw9O26OYjBqyiLmw4KmR1pBxWiN+FURvaMN
5GjV5xHo6YvI0LU0b+1LZM8I8l7MQYDWWyYUjMJePkCHyCWmnjGjjxd+Wh29NJXA7n9lsD0OPCjF
/Lx0ERDeEc8tcRsbi2Ehm0AN18ra5CkqWkdklo12V67yhjAADzYQIXFRRt2eCcJL7yWlJHDy5ZNv
Oz5l2PzdwWtJw2fTOD39OqIzXRalTljfq4IcVN0t3JPFPVEnsG/uxaJh0XzLkh1TEmqOuah57U4y
XpbevU5xZ5LzXZPRI36sBSoadmH2qn2yrQfZ5mI0brk6NFlWLWARlgCktp6/kf+vnRLlPWiJpLlR
q4MA7x05sFFhNGB1pYKRdnIroLejxo3GLS1pHdKcb05w6qVNwqn5aC52LTY4YJ7Lp05oJVj+jm1y
pUH/yjhQ5N5lxGiltlYzSPuYBSN0EoqE69tYdi3n6oZEVnCSk8RwOk6qtGVd73nA7AGaAuFWo2ti
XEckfIuB4gVbmOCwLQVOdr+eyJ0+tEep7pIKxQC+iSOcoWDu/+35I3bPfS3BvOlwZpdPhELR2r+W
vLKE0uS0jL7UQrcwKSNB9uVWR1dKjV9/p+IxqXSIfj6yPEmKsLIw190WsikOIw/shrF3L07d9A3j
pU4VSSkyrSBIyLPspx6ymKhqdDMUELqv3rJ/x9ndm8qXlBNYU2Fm1oxmVg7UGjOv8jv1915vIb1x
UOb5MAZLY49VQ/wNzm7FWGDy5oaJQJ1hD0+cPfqXqizgzSt6oVrZhIpj23eL1UBvyo6Hgcm6LV0D
iI2e8xi+Ou0CNna7i2t1Gb5MNIyx6EvailIWh/pOFe2+9i71BVNED/cCP3bsgaQhTABtURt3apTl
/Vt0gHWCJReuAq3jCKM+Nm0lv0roWhob/bpAvMzTNBppc+gdhM1ZE2+Uaj18iBf8/8QOAgK1WJsP
JvXSFBjFP0mL0UQ0v5wUXOc8S4S9ZGQfX5qxa9rCMo+9DX0U2f4hMbaSPxCKQ3M6476lQnLGPeAQ
V8hIqBj9y1Oo+HORsHClpaoRRjd0wblcq/NVTczDrgkEMBisP2hn2KUb9y8ej3dAzlwHLjQmVtsk
FdpvlFDQCF2a1fod4EYP1IIeLIOW6EoerMi56gluJC5RbCXFsHRKzlEpoKgUdj7ZPcXJekX0Twer
k+c5POwmPWum47huP4uSMssysUU2uUqQ2YMnLI5Z5vzU7d9atE6Exu4a+QnGTbw9wLUEXQZkIuQZ
IUE+KvkYH82Mb4BYFlW+I0m9v79x7Fql5OE49bRe+f8wx2nCM9F/isiF/KIrNwbcrqymH6tSjxqv
oIkg6BX03UnoawYK3HYRm+7LSakqc+bbPv8KkmXJueOP+krzKb0jcLjxrbfwM6JCWSlTRbw+sixJ
AzlWiLenFqMFbBlY6YmmGSgBQrF1M7ApIcgNYtqqVtYo6f5rqjyUHMqvoMPYYID/Y7e/qjmNNQzT
3EFgCu7LwXgtDuP0NUG+PC2BD5xBLFv01CG/irJVPIoBrjYNwUBPZw5IEF1WYOusadH4+nA60Y+A
Sfq40KnQii3vGOPbl5E3GGT8obS3ZoVqIrBjllIzAZjL27lzdosVZ+soyMluKBe8WOL7xf5KJeN+
4F0zr883GptRS7l2zMorkyz18731fhZzHIPQEle8ynAkKxjrjJqXBNrpmwcfAnSNdVJF4S41XacX
LRJta5QUtmN3bBjIyRDCRwJPlOmk4dreiqIV3qCZqGHgUW4d2gnRZf8D3OXOYcKuA5lY6dIPJIhF
UatzJmr3nBdKgxexnhjd6HKTdXIL7S84VcBz3eus+khfVb12S72LY8gSXH72BZLqBT41z/CILHJA
eMdmRSnve59GHSF0wguKPK3cInwBeNH2Uu3OWM0INbQWA24VJsLZ4EIMpsAA7U4ijoPOiVoxjYQY
NwBvFSbNnM2S8Z2/9ReIAREN9ln0T1WxDGNeeedSGswqzuOB1+r7JhXQZdeTLkB08XiuJ4Uz8hYD
qCbDxi/KoL2ziUvOrbMbM5/CihFBGorris4U0S8jylQuolfTC3T5ZRuiU+RBEpKUyq35Lfc6pq7j
5JePdZTu7Gg2RoKoBs/RX/pT3tuLiHUQEzyeXAgU9Fkih4p8teMq5hx1m+Q7DcfbsXWb3/w5tFqb
FIT6JWEITnLE9mPWzlmZwtYZv1UbizUIkYzRLrWE+z8FokrHaUABi+6rudxAC+Wuubzq4Zi+8T/h
7ikypcZkIsLPT/lLW+85XTJV1q7fN+yhQsqbcqETmMj+RjbQIyUhFB2JyWEwSO03+vjkEgAT2cg1
FRDUpfP2TxZILndANtpoxatNQEBGZPGwOscUWbzDDrJfi/nQoB5JWkJwZY+Ki6KC7luNPLExNxKX
UsM5/ITs4ZXQRjUPmAxAD4n553GJMFKmvzMj1+FqDhSceEoGAPPKApY/k9I7xqg1dJzbDd28Z+Lg
qcwQbTwQ4IWspJRdwHuES17zWlK9UTSJIRQzuwDLvYxFO+B15f5Xh++Oe8WbDYNJ+Y9pSkGFbp6/
goayKMg4umAtCPGNvn4w3sHnor8WL//w5XGcYz5+InNtUz3kVDQT4OBPfHVfJlA69vLGkGdNZaEJ
JzLqf5bDHFTVgm+aFBi/kKGYTNLFI42UnEuzYQx3baHg7n0bAMMboaa2DP/ec5kIp03VZvhJWWXK
O0cqB2XYJHpGrHA7hehSWjTI2JwmRbm9J95wd+f1yWiS57MwgxOQYDoA3RFL4sXvkm22f0lmLzFi
B/fOpgXCnQlr0He/3AOy7PiydcYPyvjJhn3wCg3OSKKET6vs1x9NwmEcMqU4BXgZwcrTFEuoLnOy
eIgVk1WocEdDlJ0EjIb9JcXKryRxq87gL895hia/0oXrE3BNiA/NoSDfFxT8L4Sl9yJzaD6qyW2Z
GQza8Wmlt0sCA2m+aE8LGnBiVj+RfCT5aH9lH+iQdHr9siObU7i1WT3o+RG2oTGdsNNMvN5M/gyW
DhtX9UFMMB/u/E6eTn0gf8XeAdb6tEacsBlkxD9MflTJ/XHxgIx2YxmmDUBK5qKZwQ99QKewOnTH
5T2prHrKwI3DkDRvD5iNq48Cid9fYODLtgL1K/29J3GL7M9Ebjb/gTV3aCvA5ZRndQLvx0q5YKsh
SQ4eSjs317LVFtwPabj68z3xYJennMESnpHynSjzvU9vvykTpHMFS0t0kp5buc9jYjVWgF4/wzme
WB4R3IPwovbzFZTsFvFxeelIkb58FCfYVw/RfRH+zjLpoqcs8fIWUO1+mFykUhPFx0v2s4463lN5
E8GiGDVoQAzYXVpGB+ND3+EIGYt/S93mSeES+8MRE8kfHnqVn3JECIP8C7gz9oZnAGOu3PT3Eleb
hWSxGrQoLL9J4TUI9uSYJKJ7aK7raFmG55HMjMNRPFa5GPIWWI5vA6dsaAy0qZj1yIDbWtYdPWXK
K2VwpqFTSzR5e/l9JJ6NkPykoLiqZIgQuIe4hobyseWNsUzBVhRiV7xnOZDkODAC2mJeYGBqsKOu
LdNj5mWLK56AOcFXQqBebti6VbEPdiV3k6smY6sJpDeXRYOkYCPBFHkIJ/gxiCDORGn7mWWlTDcQ
UngZ4H3B+TXgB2s1ceE6SozZn1yLkApSGwY/Fb2fCsEE3MIsg6JxbHO75k9ho2EXV3pBKEC+0ulV
zfqN3ysglAB19VllpGdWmKHzFedtmKIq4165ZiYgrREKZxEeFWL30uoEPSSvCeY8HrTjA3liXe9O
jVb4Kic9bf+aNtYrcxzbvmP7PXYN5S7+wmY5LnM+N+aV0xp7p24rlvRwx9F0u6IShehZLQtGOqBC
ipgSISulV8Kj8wqtwlB/KR8nOWDXUe3mJs5X2IHx13PO9xao8s/iaW1NeUlIWiLkd9BtM3q9LupL
SaqhNEmxrNmA/UorX6XZVTEwAtZpuyXZZUzwy+re+iBTxqA7Aqd26oDLAvmMSGCSo+VkatlnthSB
ZRVY1qgsHUNIpLb16CS680BVI+VrlL70MYcespWOu81ywzuZbxkTyzknaCeNYzwutYiKENvB830s
QJYsz2ZDrjCyy5/cyPS2Bf9xdkr8rVXv58E2G9BfZLSoBt9YarxSkabbS8lrUKcqh9C4KXycO5ja
/4gyiI0cRC3tFe3DzKCeAxZP/6ry3emF4r0Pz767Acms32PJiWPifZxCK1gdIM/Itn4QR0JbpI+4
yBtVWx58YKyWFUfAAX1F99401brEPTfGy3gMKopjmlYFVlRsIRXF3vexlbC7ZmeBKJuHZRd/A5Xz
ZJ6mFGF3BUEvetThz9y04+YEPGEI8GovO9oe8SOUkvHb0WY3ttd6NM4vEXyakazpVw/eLZpcVOef
AC5zdHdUREHrj0nS8rdnESg1KQ21CWNBHkuYC2yjv1+ABGLo1JRGcd/lNZvbmThz1fyTGmuqevpG
83REOEfxk3l95nErzKcp+vK9/1IctWu4Pevu3J0IhX/NIXFhMq1RisU4vS7u7ZBM0HOh6bOXl8HK
LkgeifTh1fO24W66fx3D2tuw75P6XG3hHA+rcp5AovNlZNYxAuYsELuJ5n0ABVt4n1k/af+lkTT6
QxmOuLZ9EORAB1EyoWFv6Z6jCqnGph1+gpCJWzX5Kj1TkJU5n72AhXYVbnYbTmO3c6FHB/S2UAEu
n3Wkf12c4bOwsM+wEwDze77KdmLV9vulWA6LNd3FD5wcI94Z8yx9M66YO00ApY1fc1nxDKqe39ig
nzrrcNh81VALiUR+lS1vEW+pUFwtfhjSzOsU0Jqe1Hwxa2/aTqlvf9jGn6rFVR9v/JIl6zyz0wgJ
irctoHksCkH7Z6YDLxIUfpBRT2STn/oAS6/0JmbDd2tiGtsqi+QL4gfngU7BAha0H3CAL6jCb1qL
ptyPdyM5M+f7Y32GIuLKaEvwLvCdEAk/Vxu2NnmvBhTu/plsuVxl2ks4YHSMAqKGW4m+orlqWEu6
Kc+3j/ww5R1FNI5EUV7nRrVCFKROkznJGf8Hvhpg651o9Nj/q1wNTvEmp2OZlYR1VDR2v9ihmo2j
xEDa0kMs6dI0F3ND7Dk8SwQ6ciEvjjLiisaVES0ZC7npkDYEPubtwbbD0SIWBNpq9n4MlZF1zOKV
iCFtA0kd22rl0JhHUPOq6Oz7VoEZBrfGn4aR1GQLdmRXVhHGQ7lewgwfiL3Aq3OCeIyXn/2Gb1Bs
ApY44ZPXXoyFFcEWtjRqN8hkCNAYh0YvfSCsgGBtlLzbaB1LspMc3upT6e7C9J38CdDaMaXOctI4
4PxOUS9MaEDLUzeb4nQ5CsaDWy766QKC5mjAVPdBf/gOoyX0DOuZKzkyZ/0PjgQDqRFhM6KzMLdR
EufcxzyWEbUGSnPuo4DWGHp5UKfzioPj7PoSLdSIFRUdn2X/34X1FNTm1Habnc55IwZZxaPv8bxS
jZmFKTK1995se5gzSW59dqw4WO/D6N+2yHiZjX3dkPRFQqazX2xqNl3EvofaFBh8F3sqKMXooFSU
OTl0qAZu0lOAyqHtjRYbAE5cngjalVdOZOPTExz4TtJqu+9pR913JSjOqjnjTfKRBZklYA5DIEgn
Db+a+OXrkbnJ1o4x/MWgmScL1oobgD9LyIKVHeBmkzlxs6giTnRvkPre/HYxu9v3XrjSGcQdpaP1
VSnRWP2131oOho+RV9KQEe75LHKNc6PXiiMBQBlGQCQfpzHrLF1DZACRw82H9VBMRQO1eSc5xIJN
BO5ufd7a8TXhYomr0KGIVo8zABU8tKfsVMO4lqROlNc+mqcBxwBroKI08iEY2XOl69asq+ujMGlt
v3fhbSbMzTv0u98/GHBYkb1+i0D/Zf/eM14Q6Dz1Lz9DypEGb5uXjtYlE3z4OOZbONzXdWVI+n/H
JSwNxhZjHLAtgd5MYVsJatk8RrtACCs3rqxW98SEjZd3tFgAMdSJUuPS7lVKaDjKYtKlzrpUZn+O
QWa9R4g7eInp6BAiTOxrKmaczIXKChCipZX+aVp04+v6p7rdgFK9ut/KWkgQomAiBXPsrpF/8dkg
+TMTSO8Ntv6Jt2vPMDQfdaW0K5YBNIX/NsKh8mKliqyznsw396RonYtfRkhyLmXb8Tu4/fSPhs+z
LuXloiF9FlY9RPvmLQMKgMV8PybpX+US2XchG33ip4gcklmyqxgYmbnMNhrRGBzjA4pb2T8dbEsh
tRDUAQIzXICQqRoMproh/MIAjQM6afd4aoUqrXk2afuU4yV5oVzuXxi8cuKkW9sfrLauFpzx6ZFe
HmCPXO3+WuLi3NPv3emzr8JquPq9lIDZoDB7H99UT+dVX+p5tLTUqRsTv2/y8x6NPjbSxCn/+P2C
uda0RucoNMrMOi4jMpEBK0JQkpHm/IcS1OBL91KM3OFElWsNQrOcFEndlZgAUlifvcaN1bhSor2z
5Jtzcqudq3/4L6Y02EBsCQeUvBcanvpVSCJo6ZMkS9jB8nj6acbLyoN7gGIpL0mL41YgWGqAHaeM
+hwxUmCXI7MGfFRYhZjB4fBGWmAjgqZ7dFmb1NZCP4Gf5dMChYPEiBENVZDJWXqW+C8nzuqcBUwf
SlkAznn6+PpH3/p04WqBKii58CNQ7Q5FAsFt4yI49vZgjCgj/A8YuCc5eSSlf0sC+D8q2L0+9wak
hyfzFCfmvQ3coDhBEH2Ds/5pHexKAgo+I4ZiCAxKjy946MuJU9PHY5NHw+D+7L4vgYZGutRCWr8d
A3ddBOWCCv3EFgwgrSMh/tcY0qVPWzOT93YTGTiTYSOSy0fOkUtnFofss69+SyZ1lXPIK507XGk5
ymEzEmh7rJMmZFaGo/lAcmo8IdctiTpxl2iblEHjkMupwJ0FH32WBscVdwZUgqlvnImkkAacvAWl
ZQ6hWh3DVow6KjMvQZHmjOjuBAuxqFWwyl/0/S3e9ZZD6qWJqStVhabGEcE1DwjSV9lbI3x1bWQR
xQQXyRf6WAlWJR5tvGTrf2DONaM3uXpNN/UuiHjyZxeQ57Z06h49Ogd/9/Cnotymjufn6+MyIKu/
nZffL2Bx8cgMURAkb/fidi5LnmkQ3LrctND6LYdjpkVitRMsXfdkxCqM0O2U7DaEb+DKu4qWISJr
sG3WEkihZjWB/jLNMxuw9AZ5qsDfd4ROpIiKPhUmR/T2wkxWFqyqufaZYGsgZc1cZG2QTq5Nv8Cl
oPFVTEC6y8cNZ/4OXCKGGVaEeJ0zOTxVO/TbJ3gUS/OuTQyEYbecms0+t/jEPsvXpV2aNjtPnucx
LXvmqyhpIcz8/V3CibSEFTafAdhl8oYp+Mfmx7/1BQAO74jlRsQiOgonztsI+LdgpQPys5C+qCd4
HjaPDpfOyiDKEhaWWvoW/O25BFnoBeurgYiTD6jWk8GZ9lh3H1rSXUCsNr4SQarafDMAh30j3iiN
um0lENHnfPo1LW6egJtjRUohSDrNL1CjzkPfQPoKoQjfzL9lvzIijtVeOMTKZJjqglnPjRnevV3Y
xW6FT/ar0Ic6dFhfT3RQ0UL2Y2un7cDCiZgynJ+DQaNPfLR4JFjfT5lOi5F9wLgDl0SgFMk/XV6Z
VAthKJFmbkXWiIk+g/JznX0WdViYJWx22iQrdCRs2Azjl/dNUsGfAPMGCmzEt6NpV4smeCRXZd5N
+3uV7aIHxnRG96y71q3I7ZZp8hKLi731BUZelC1UtxZ/hQ5f5Yrb9aSrZmpx7AaxO2RJqu42iQpx
aQdHIHb1PxIEJnCQp1yIl1iYowk1GWO+KoNyEnMQXFtAdH9GFnS9t/cuCtunXz/RZm42CKifyZ5L
xhdFfubdhY2KRHSo9csMiM434uBhtV3+2wln1asXKBjcTgx279doBgZYtxQYUoZzoXK1yaL4u5pe
aRJDa9UHdVfoejXaTEckPZpoliLWXHdGA2SpdI6ySbyDzf137UPde1VknfdS6a+lkSHy+cpHTZsS
uPCHnDkeXZ0mxZQZSAC8umFdKvUWOEIyhS/YkvL1oZgaTyT1RMrJ2yHNVvkp4RzM9/98FQI8p71c
ELnjmbh6bASGwn2pYfFmmeoiqTLsTs/COR1PDOmnmSQUzUqpn0j780yRG0skwkq1D5r97GsE75Nt
WM6AvzZ6fd+ZbybL9gHhFXk/+gQ5VaLsQ85tfvw8QM4UN5UHfvPtVBJrnKt0/ZrSnAjdRyWRU4oW
KyvE6Df333EBgocALs0f5572hg1wcECRKETjT0GuRhhe+1vCivBpojd8ww2qwWuNsyhGmnb6P1bv
vNC7vEpMPSiXL7ilr20jcutVxWlhDojGM8++U6sKbuXZE9rAlGtfW3aeMIqtwrOuvooV9JimSTm8
cB78p1Mc76s+12L4JQ5LRcUK9LOHU2LHyD+Uec10+nVg4IrLEtp0RW8wmeDk32pI9Qh9BH0a58hy
IwrkKddzR+WSBbFLOAyjW3nCVYpNOsAFz5jbHjvHvCRPOqo6YZV74Bdup42bpgk5ma/0UdT9mA7S
Oooou6iAFv7+EETToZ1nA+u1ZDwrzX+XuP3aIGnpVDOB1nstHF+B+a0hLaaNpX2ekbMRqwMK+BGI
sZMBeSi9PnsnbH1QmX8X1ECFbBWBQiYc329jozAOBLJ5zWVeLbFkgXf1bQoBaBxg4zM+NCTjgEX0
NWw6gP0IXPLL4QjnRRolC1spG+o2t61a8FnqXo6jYT/2VqkUZq2427mVjx/RFpGbwRXdXN85Iq0i
RmjuH2ibkfI+dkOkalfBAH742SdACQ295CRypOUX1oNjjBWG7WfJTOnNxFRbk22Vtwcn6/I2vHEf
YXxH57yejOq2Ww2uWiUHDcp4uRmJBA/se4FA3uZqC+JvWlgM3375wQmTUCrOvSl9pcOoA4++3NmX
QiZObaDxJcmauxoTJ59ZuZgqVo8fKhlG8u5kTxV8QPvBOZfCjxplpWVfW+3Kj/vWLB2zZPZxtQBY
2jV8rCnmuV3VFVJIc0QNoaAirp6JWInRq0nXoW/o/w242lV111U5PvIFvnHNSVMZoAopfQrpZ2jA
K1AzvUZhb/LgTnbDkxqHrDIZ3jVlA7MKhaACJujLyJ+9SOm0Nn3ZZi/oZdCes609LDjsFN1D2IFf
8mJQEsBg4QlPea+4EIyHf54aAZHKcjz/h/19vvWRY1dLjrM5urfExgBovR58kl8CKtG/lbrARuRv
5i2T7VJ4PPJg+HaZ+20ZnO/XNz5riaFRmTnD2zUBQFkmghXtbyJjylcFqR5Ndhdjibtm9ToNo/+j
wUCE9YpQQ6NKciOc1HjD5UOjhI1MSv++M/RGGxKZB5rAIteyspcMoSjB4S+MdQUp128tSDMW+xsg
ImEZmduu1vDTd/ATmOVpAo3SCELomB2DjCKXN+6kIqV2SMuOQkba/XjAZaId3ePQAzoaO2jnUmqg
nCumFSkeqZ3luZh+gQRhS/yFYQbW3b5oicdwHYG/CnudNeX8n8DjcdnBJ96m1Pn8d+xVhQfXckYX
AbAV0cdGtj+so6O0K0ZNhiSMiowwO0zlA0vHRbC+RPRfd6BUZVcCjLGdGe1N+rXto2a96ziiBGf4
y9FNf8/zYo315Wa/hrktdi8qGeJVFu0ingEfVV3e6qp5w2bEKAHrynqvmH5+fFkgK06cuZjEKazO
Nd/WH5fwADPbM56DZ1OvuUEiBS0yZU99itNxnrniEBZTO/POZXxWegDoYrzvcEazMsf4DD4F6wK3
vvgOOQUehl+oIOqV29Vuhp1Hjk52b6pMVh1W9vOB5xuRRqbPbiOErR2Tyf1+St4oSArpQeTm9trs
QU54xx/R4c/u72P+Zt2MCwSrqO483SlL69wOK/tUEWA2rpxGCxwU21M80tC6F7MghKInHnWpcEzm
JAS7xus0wJ2jGv0dey9nY34pZt+pwqrDHkZVvsKDDaxLBnVR7SX6CTk0o9bvCrnV68zdtky144zL
BhZm6v4EATUjR3gzH4jE1mNku1HfYZqmjSiUTz7woYZ8mhpq1ze7jiAsKQZX24dijvcQ1KFZwnFf
n9brwaSfy/Mf+99KNFM2CqDYoEZJW0mGgY1Mt/3GN91faSH4YD7wkcWcG+aNxtACjb6wefn2FKVv
fVkpW60NXDTQIttjn6vqyc9VEHIqnGaT55OsCNR6Uv8/lfa7PMzla2vjm38h64eMOqoLUFt2EzYm
vA+XQPKIK78XcGKxf8DV2iQ19fkibCNqGdv3jVHQwfcfYjUQKcfQtszXmbDBASdRGmA9LVSjaGIm
6nxbFeKK+1K6zgjO46RzXAcIw6T3yk1jJssZErTGxUz+VJr2C1jZ1n+fqeUgDGbso/yqP77eK+iJ
taRdaiPAjoVer1FrqkxYuw8VDNlEpE0xTBmAzVsGH6vTuTyG5OuuWKgx0mX68iRdkO2dIi00qpXg
9eE3yXEEoCOE7eWOLWojp4/Kz3PkAvrC4o0I1YTkbHziym4GvqCkafOguvZQSVlYXFUOMTsBPYEt
U5zPiihvUwiNLUgEA5v7yKbGZArPK8OApV4hXeIWoc8XmLQaTWFae6SzFGMHQIZrKxs6FY2JdGXA
M09zw6YE99NYToaEYlr9b63n6FwOok6Gup+XwZclfH3gDYwji4JuBDOhi2P3TvOJp5WLvBTcxVGi
J/s38ScZSjq1oRsOnF98wbilqUdO6g6TRmRx0k+WsqrUbiD+tjqKZcapiQRJndYPCRhXIZU/5XMW
r377x91fhd8y48x8K+ynxMtCBPZtFhmWr52wcrpPBDAsbn4Tu23ZQBWoGy7gvFllh5X3GU3MoyND
AxptA7FsBQTEVZI8OKxidWLhaVF/QOycrT9/ThFWacVaeuwqfMS5ALQGvfrBk5/DtJ+jhYyCZDsQ
y3yfR2bcj8Q66nG9AsspAZG2eHeOyNEMZxzULOdnKc5Phb3TW4ozy+ctJqTCaRz2+1y8kVmQpr9V
DeZuHp0DNczu7qdknwOOOM4vRoB+szknTtFAVsGMMF7Zf4Za2mUfR9gHpFIt9LV37x/2Lb0Hck2n
zFo2T3HboV+nwlR7p9QFSSoUxoZtXgSNILhrmFxBaNfJdAkCQCUAXJkND+aJ+V/do44OyWUzBz5r
K7qiSMj7wD5YR+z1ArwEX2XxIACYZBhQ0Idl+Zj1rk5YdhqY9mVs9LlA5cR9utD4qYqiAfnUydF+
lhOhfp+T/07c4zL2E8nPj9gZv/gtmFulIDI8kkAxNQLoJszVrhBx9+UzjAzG7H5HykSl/XfgbSLx
ofl43e5pfBQF4ZkxeFOZsx84YMuLPk1VxZAW6ftRpGi2imfM8VWbm9wUyrCgT7WMTrTfmgoTRLI7
m6VirY+P9QEC0MiKMRlNemSTG7EQBaxONzM8MbXrI9lccOo1WCZuTr3EJ5QZc3uVOdD5AqnZpaib
b6oC7Jy1LIaCa1C1SXUKvBbn/PrWO3+3GbvVpydyDCzsX6xQDDzkqHw2EKNSqqs0/bYaFOrJeXxB
e2561my0OJ7NYkyUvcwcMwYdCir0oQm6ecdr9Gxid1ihNsQTMXawJymXZwiOmWAsOnuaUytBUJtP
5rQ1e+6sAtF10c0zbWo7OlbAzqR5dEvJ+Ug/aKtSusfW4IAB27aI6/RfL2KxFvmOImf1LIxgRLZv
o4TXYLyb0bXuI5ZhD+Hy6RlShOPpAUF2E29ptRrsLmSdKtlvOOTvdmAwgKHFIOKzpCyfH/B4NEkE
8pivpAm10PNMXfdZKyOS2/p7mYmH2nB4PQWrikCX9uFtnFTc5I9L0i1pO/FPAfQt6eP036KgBU22
2TJwWXW6eHg9eICVJYAAW9eV6jYzPS/nJdvDraNjhcjOroe9bAqOtLN/I3CYIvTnNBaOHDyxxIiL
WJH0e9TtK9IkF14e5/lI14gROxMe8AM9dY/IPeu4q+bas6WtUZEqPuFgki2LYuXZ1AR7r/qb6XKo
pn3UJg7Z2zzlZGFYtcJg3xqAJj+t7gc8CMPRfGm6kVg3v8nTTPpLDfyfHIio3ZOJo0Z2GyOwz4+m
keWQgYaPNnOW9Hs5ybwkgFE6M5Do63lgACc604OVZxmvDEYsicxDe6djySdFY243qqruFYyND9m2
kamjd1+MLL3URczfSWOASUoqb7OJpXuWcZt+81Ct1Fgrim8csMtxyIM0RVL5w2FX6bj4OWXblCG0
08HTnF7IKWMAi6qmJonx8EP53ghR1NZBgBlcWaUKs9ZPCIuKwTtOCxYhgOr8FaJ7g+BHYgMYq7XA
jYb1rx7XD8JXGGZl3hciZlj+k+AklCHCstI01WHZTIBIdPCB5x8tXsiFQDiG/2cRXr+Oa+2FGDHv
3zRHL4oOVuD3lzTunJuSxs64fE1qogIImLwECFqXTGeWNQVH1ARS8Aao1DzRVHXgXK7MSeetKA5z
+h8OWhBAneaGt0awyy3jm7pCXV44ZOFxD+5lDwzs8SjFHHVkvN7Ch/4XIp9K4ANqfDgw3M+gKV6P
DW0lng4Tz+1+Q2MUT/y8LdhGKGz3gk1dzcopZlJCXreybYKk1eYs/LLF14hgzFQwJgoAayg/xj8q
RtVWfg+oqyrEew3JySoLcVRx2xNbE6sWg9DHecPVdmlU+SDURgD0QJ2gzN9y9LjZGWHMu+8mtEKX
Dpio857VSukqOklSQh5ArKphhuZYBKAw2vi3EH0VKUHYpy22teD9YUwLGnLTvoXDg2e6j2hYJb/f
AUrIUze8HqdgWUmhe3y7AwUeDmpGYCgRBVcbS2QzUuHT29QiUWP7Nhzdn3hbqZbrGhcg+/l1Jqsn
p3zCCCvr20feGHy2jLivh8uJOYh0mli6yWKJkMS3opqQ2DoHSZe4xH1VRCyiSEKVor2Mz1JoZR10
gJhcmvWBn6Ol42jm8iQqJD34z4icHnWdY9bRLkEYWTNKNR0+PKE4h6izbUu2vIBNeJvexUP+a/rf
p4/9I8Blg7RC+hRoIxAv5H/0S9cAYsTGysPd0fw21uXOBcKRw1tuN1cVHkL6wJFxKXveAQ0ywIfK
CsxES9GGSLAjNhws6+3bNGRxvCc7MK40lzrAYxW47hejsNNgdJvqFwcykKg4Ea56uhxyju6UvKmQ
tbQA6VT7RGOCqG7hB0zRAEUx1T9j7g8zhsfOhzwG+ojnPN8lWDl8+c1dZoUB42EJ36vDfF5sPAR/
4otXCEOJUv+meYuuOjBtZNkuVag9xgOCQXO22wbAi1IdKRFREinYCQz+woTPnJXttEsgu946kiDJ
5V18ZbTSgvzSiHrFdFRd12ZNIDsPiiEP1hkDyjERT/h8xLOpvmBZMM+yjn80Jmy+U8ZhH2ZZLeuR
NHNgS9rLSzL4KTZX7urTtVc/ctkR6jSQqhmtvJzN0bo4IElwBeTBjDDMgDOjQyXsvLeur5oad106
Ae2BaiYzhf2mDmkBcbB/gGFrd3tO9qaxbbEdAeUTy5FivcSriepyz0iLPTusOMQSdNskqAsZBSj/
mrqKu/5MI35pHOrYwKS9owNSYvyT8q2EfxKceTNfNGHuqJTZ4CIerlRUvdu1+85SUdXwVb2FVyYs
I4mpahvJerWv4Aww4p2w5ZSFn1ygBDbEBb0vLPuHRZVnjOgRpZNg6SQP0KkrrUgTRQpPboTLKyK5
pXb3Uya6nkM2KLjCLh4mg9w68ABCzdnmFk6Tp/AqMg+Ev7WSdD1zPxtWzyjs+GPFiQzFrWjj94Ma
At0TBASXw7D9CXhxILvwkUjSiKuinDRwDCs/UO2Nw1lzvMMVTdA1zcAde6R3xur6r8UDPPCWzJaX
RrfhTer1gKWF1kz10FjYNPaGDJhUoO3pDBwPcsouSGlOP5s0B4pxbkiDOfkZO+zlmqxZets94KFe
wZfiJs1FaYn3yYL3sAPusKeCFIc29ey/rBK2p0XWIgVrYtqFZjJX9HeEb1GWHU+7w8oawQ9gLwDX
eBTE4TEnwQCUrHfJs2/wpWLGShDRm1msgm6wTMU8yVLLo9d8E0fsSUIfGxIlQSzbtziOoVnoFgiq
Bi6jkzC8iJtgQXe985IqzcEt/JlAmdHgjlmGuaZ2KY5h/bzsR3K1+u9xLyU+yqmI+tKuChRzI1C9
LQsZBzJPsX0+YRVyGLF4tQAM+p+WHB00sQUbbIvzEkCLCPr4i1exTI4jsfxVm67HVWDyQkVpLzQl
jxiCstNXNx0O/yj17k9X9MeKkt6pD7sKi+70rIDdn+ns2aj8LmdFf6s2LFIiGStBcCV8Muf/5XdL
7O/owl39nsSZ9UgGZlhX1/6U1W+1JHcJcse5O0xTMu9gQiTGyO6mD/33GB6yLidrNtHdvLu3k1Z4
BdpkntJ5P+170P2ubfYNok/H1HXBui2XGvpJmH9g3QKnyHCRyJ52q8waiGSj9+ne3JGHaPSKPvQp
E6kMouUjfoLp45nHonFQyisdLlde2tDY/+3J3Bx0ILjCKnHeg/NxDYUsadKdwMibCR4DeaM16vPz
tuCq29qJLk5QPJRCv1DcidZFpEipeOzCQnzO4n+fk4524mp59IHrf3yQ4CG1AEYatJXkhqwgqHIi
nu9WR/B5+G8kVGoqL3KlGuMpsOt5L8FI5sw+91gwBkHay5qNv33ir9qyj8z0mzLU1UTelj8nId5p
41nLUBGamGJhu/Tn0OkRniTvrvXrkS1148rCPN+Xhp7pF+qa3eYxuYMZddNVryFHot4OmgXstDfK
h6ADq6LaQ93kyvuVemPSIbhFjlKwwgIlmfxJHrP07OC33X/KEv9SjpJP0KGLGouCds2+vVT911rx
2oYapSFXFoaLzbpPO3jCcxiv0SUTLmqBRGpZRNj+diBSnMvpwp8s/+NuYwEklqd9vWi3wfZUAyTw
xa5IULRAn2aj6hF2iGMbjqSnM74491ERhP0EMKJJq30J/jQxgOayFJjcGTZmhXkDQxKXcE3KQ4VC
2jow8nGmzvXnSFK6tPDjRaEv0ZSU2nt8NdZT02DTF/XedVC5oAMRNW7NOHVYG1RYq7KRw8NXsGZs
5wq63k3S6ZeX46GNJ4GGviGfog/9yqXqPaNlMQHuwGPWcUA9vzLc4FPeZZXcJT9RVg0HBX5aEuGs
pkedccYmM7juJhpUECHxMxQmXxWDvrfB0ShNNHNOEBtKBcR4tbSwxInyUCKd7o86fqxgJM5gYrIs
XSGVyqE8ejh20Y9fpULl0RREug6MfrQP39yIf2oAsW1U4ZnTi4ILQ/PwpFjnc2btxUbI6ogrIkJa
c/hugK/7X6qFd6jr3sEHlE35gHV12xwcWnwC23zHyqCz2ZTKUB2KQlQQoop/lJY4GrNlk5QNn0n4
oAj4mxTW2tnISQl25KsUOK7NuGPk20ptx8gbwlllG13CTWUJ5TOIuEYKdvQ7++/5O1cy1jae5q8d
NPiv5udk90snChDZbQh9vT1O4FMIJsrGVn9a4kSRCgGUO36nFvtMwrUUiRVVhREoNbNLp5nPDmSJ
R1KEJwVGARgC827MiF/k3/4q7Arxx98SqVzFm6rHMl1G15KSjaoc4dtFC+GWMAzhkkgJcCGeGIVB
5MOgTTlxt4JZbK5vLKvX7fPOcvdq2b7RNmMirx3Rnx/I+FGTphnCKD1QOHE5XrOFmuAdiolxQhWt
n+veXIG78goUCxZYV2KNk9jNOVOpI/3rt6xFOTNMevT35JQVsbiWh8dvfHXwmBuympVuvvfq2phE
2tVzziOg3ymDIH2Nztu3nOVAozJQiMW43GLK58NV6YgWB/Y5cbGx1rOcfL87ua8PGQZShO+kt9Xb
LX7J2F010/cadQi+4Fgx9xSnOjMfHTbb3Us6JCBsMmpXFwMCVkS0MdFCz594AyTdT+M0p8IfxgCs
NVE9aGBSOSlx+ecbyL6rZ5E+nYJHCtn/4A1ZbyW6oAbdClUmDrGPWC9p2/LP5ivmU1eU1cCrrKGS
LNBSRVj0mslwYhyjdAvYtePSUjn1Ry3LA+YIiU9PYL8J7oZ5NvJK1//a7oWjf3MsGahds+r+zc44
lidFI50Ma2K2ge0Qi+AjxyysqvNZAWJ0NhHPbOblPPbKEohIh+xhQya0JCk1XF6D0QbWZtxBiIsm
t5oXFobAXx2x3miem16p7wj9e18U3DxFt99h1wUP1eaxC0pMNQJXY/vAE+3zwbbsEvE+Nbf8XzS+
Tbg6u+UqGvXp58h7hC+gjXk7xZj+I2FOSN8zpWp4QgRWbLEjbkUnhefLSSGw0UV281c5unxTKvv5
FjkvUX/cQPfPG4pSoG62sp5AtFEBwj4XhPNncA6rR7CqIXQ1tyc5/27Fihu6AKOgsYaRstQe3D+/
W+4VvOxNu49H+wysZgBtbLHn81MNx9A5AiZK0m+Ru7I//naClRON6X+4HO8qzGbtZ+8TYLgDzlWW
b7U9Dze9H/vudFKlFcuxpcko6YAydlxsbdYo3IcmkCY0BtGmiXcp036TvxLmIiJRH37s5kwZoYyS
zpcZ+F1JT+nPY6+9z9qthMJq59bBhf9q0DHg7NaILK15yjBabqV7VIIOh/9J0rRAVD++ExjirP1u
SsDxit4jKaVENbqVeyiB3bWnFmy7RVMLhTh1gB1rxvik71BSHJFAFQsKp5xrJaqWfcVj0V656oYC
/jFLljl/jjV+k4XGMOM+3RUP6ykMrsDBDzxDPNMY8QfbgGunXmxRspdbO1scj4uJZBbSXkGakO+G
oTv2DXeJBZk+rJuPkEiB/a1yFSaMW94oIVRNycSiTiEIpgiBlOiKd2ntKaXm+0rZrQFNga/Kwqai
bl3fXaaaE6xmpyzb1JlavNVbudBxix4HuwrLgeY8TSsHdohfLiPNTZr+b5lUNHndji3oZHEz6mY2
hCpfyymNxDpdu7M6seG25Gcs6brXF3TJ867i4p/klXJrOAxEBCMNnKmy73agNVpjMD48WwWss06k
v5kuCZkkBRxa5QnGl3Zh+tKJT4P2FAEdS/HSoe8FK7yPh1ruseEBQlT6hrDBRXuQi3s5ukzVfPqq
srQgquGFQHTc5MfmCb4/fk6PAN1Mn8vYbn2ZDvO3iFhQ8/3sLWwBenXOiVeRO17t0zkncALQckVe
KUyzKZFTlEThFKRdxYTRN5TCFaWrp16E5Dw76bcHairDCgpR33VKEv6CCc/E0DJXeXkdzMT0Kui9
ef5iVHqq2BzwJwyN1vMly2QRWFHo0BNsjm+wLyh3eIAWvoyr32/zMPEpeAGTbqkH0r6Pk9tAfFe1
uEQRxk008+qmt7XOWKPbkmQU01HwCfamvnE8VlyRuPW3X4fuvAaica96q4KCEkkmiFeqNgBK8eDu
WTcBkWhbhLBlkrf5PVrBUhNDqSmiwGl/EqLId4cGOPKbcWpo6ThzLWKHlr3Pvh6gs3rPV+xPwZnQ
/OtAelbDUnXFKfzdurvffoWvEb7ysAvsAV1medTp7qeAkgEx5Bfq/yyDrpQ9UtclzHzlrV8Zftng
CWoy56p89bqPYiSCJMOqu7asd6JlakSruZx5w+/YCkZBkcfHC+Z0q7nzsVo/QjcZhgN6b4vyeuTs
fNoYYlBTlQvPuuaQiey6EmtfMmR1q+9v4lwrS3TM28NzHMhgqg1RJLqnyluUZNxiphbGCQhb7mCX
a9VKYI6lpAj0Ocpz+niqBVf3mQQidjRudmt4jt9Kqw+Svzs//GYSw4RxK5Kz7kdNBu/9MWKiOAZo
lBN0+FtJf5lQjhWp3imoallZqYGzv5ATSKrNP4IeLC2SScPLqM2uHT3W5TM6jfuGnTq26vPcyvzE
MZf3/IZsRtEJYK7w5nJA8QscSfioNJ2XyhgSRjAntPATr8zufePD5oE1ugy/VXfe3f+Q2/VVEEsu
cUiseVrYBI4Ik6SQKdy96tkeyL4Yzn5V/LvRhH/f+9iaWxuygKK5+RS7TGGxYmLYLVb+fCwFPqD3
BF2yWHco6CHnJUkK+2+BA9CoCQQHpx6w5s9627rXwzC4lUkQBqTPvA1OTifwaXwcFzPSu1MU76ep
ZJyiu8aQ2n4rGcrYGye23kDaBnTIa2/x2+3En31Hw6ZsRyIiaJdrI6SYoKtNLxGUyr8+n8WLsRg8
SmqOqkOMQnf2dUohYzpzyZQXIcqDGyOtPxccFuFSMbYh1XoP1eT+htEsXAKmRfSiKxZKpa3QfWA7
p2/VGk6FM9Vrx1BGTHGMFN6su5h6tKd8CLGvcoeTVoDmtypLnvbaY6l+dTIsOtnDZ8MMGvo53Hvk
zkJJkP5Mp8WNNBVtevxX0qYrfpysnbA2xzfIsgjoCgz8o+YMbhBbmA9ykOf8SprT5j+1xaGGxvcZ
b3gkP3n8E7esl7C3d78aaLN/5uQYAMxP6W66DYXzM5zR2A7WelGn23ZKnbVGBFkOY+6R5DgiWS+7
+3f7RBZOlRwzPjQZ1hK3r+tjN2xZ4Xyo49FseCnIV5e24mWNwd+/Oa3nGLzbHgDjw0ryeaIDUWzC
AMiV0kx1P9LBSPRkjXCM6DyxCEK6jM+YElmlHjOTM91cM9KOPXkNM8fZiF4Hzg4/No0bbayzKMDL
aiC5MEwpDYx1NZqWNc6CuIgrgTfDcezoZ0TiXruHKcdHTYksAV/TSUxID5/ybwMUWz7b4QEwIkR9
LG7AKx7SkAl/6Ccy7uTu8R6uMsskpLrIrvK78fcFjH+pViPtOyhrNBWPK7xqE68ehUgivc163Gtl
vM14y6Y4WOXYpNkgK5brrBD9lzDRSctgDMtpW5j1woGDQxvr9jnSLGFwRenxioRP9AE8DY1fqzpr
jSH/UjYP2CfyEoP5LgRXPrOiTEu/Xlkzam7waJl32hn3P2SWuw3qoUEK6nFu3R4E/uKmWVUVGHpy
SDi+2oA3Ehq8QvRBollk+X6Rh2+0J30jGoRFfZkNxq2gy56IRKA7oKfraFAgBCm5XwAwGtNljFsg
BS9RhN9anFu4vyc2aVHKRYkHqI5p861q3k774Zkj3xRMIedEP1mgbkczZhlAcBJg3bLp06JMuU+8
AoIlQECnOeOfxoyZxzRqscVUM3hcuzp9jkS+NU/quBSMsJaJaPYAZU+pk4olpuNZI8cLfOJXWwDJ
042OlEsmYpl91glIVHQkjCsSl4dWSp50u29cv3dNr68Wuym/MbWLozkis/iydWsgU3IvXK2cowHZ
kHb1BckUyDUf6HwtFq06FDDCf/wh2hfly40hLtfILY+MXwm7QXb06eAwODvtEzHzysK8ClIl1wA3
tH5DongyJMKdI1l04Pov2xZEMSIntW9LUOg5aY/u9qz3Mxje1mZVEsNrA4un/0PDi+bngOQdbOfX
1JfaLui5HqlnWlqe3jvgcY6upT5BdagDYmhyDWbYqy5jrkt55L/9lJEuwvHJ0SW5te7XszqrGpRR
MbFmoU7/0V41+F8cGvTAy50LML32mDpOdJwasLfp+ikIzt5L6ra0yYxlFMESiQJzFeWwN0fRT1Vq
OlzrEZBrlQYNt52Rqe7aLT7leP9WxDR0gpzpTbldqFTT8b/rvL06XBfyryYWgldll3bEf4Jxw9rh
XhvB/k26eaLYqKf5Tie+GDIOsU9yEIIcxhWtAahorhIPvXZt/YHvxKEsxFbf3gZZIhSCVKQdgKz2
jzn3gOwN8YZdQAPDUXRt3T+Ffgq2/rGEuPx2XylmxoYntG1u0WrLG2Q9tr9NtIdfu1P2tB3CsXdl
Eb4ToOMtQ6QdXbL38S85K1rMGdugT/nZXpeHNWfU5rINKiSmldFeRn51IhGBax1qdomdOZ0CJbrU
y4/4pU/Jrn6ZeOazAgmmuzROZz4s6MDuf6WihpExlwD5eQ/cKR2frQnP4MaMtZ5zlvSN0tLCefTZ
7sGECoLm/J6eZI1DbsCQl6IkmFNrHFEX3+eVPElVjra7/jzm3H7TfrKgTwy+tn5w2ylTpI13eWxs
ACo6xSCgIC9LfGLaeQF3NxFF335KQmumpC5cTINEb8OgcIRzsnckRS+Gi4A0AHK5zuzDVw07U8A0
PHmOu6J0aa1FGgK5AcnGIpHpLYpzf6Gf5dtrV+Q85ybdkATR34xP2xMFIN6VnclP7bVIIzDFV8zA
iw5M1o9ruEnI2JyKHmoMH3TmazTG+PyhyhozNdA17iGmJ3cEzix5yWb18tDLqssjWyVTHZ6Ilszx
MqF3GGOg9HnsD3Cq5tW3DTUsoBHBwNjTQ/YWzYws0TdnqNzS+4UTOwJqCApJuj3yKIEsnPft/hmx
qpdckHreNm6yKzYDhTkGICn9oLNfO6NzdxlbV2IiHyAkp4E+NdGnh6ZosxZ3V9CWMlqalBmWJagY
BiDlTsXE/TdtUXQGH/Bs6DgAj/eKfbdASah8YIfXZKtIaxg5gM59Ryl+IAi6CkPVX/ZzkY/Cs7kt
0E1pPVJ5C7jlP202AqRxzwVGjJNUwy/OrkNauwj5x1cIishU7KJjn5K8Ou3e30fcPRexjXdr0UYB
ZZt8hq3ypPFBcsju8I9h882+Hd7BYvnNte5HY5njdiUn19d6MiUGpH3/Go9l/FbP22xCFIcimsBG
uLRJ1ZKZN9DFyRN8z7lJiwmTJfMUyNG4HeILGh/aUcvm0fuubHdnvKSLqDi+L8rUvBZ/rfcX/KtX
ATn7DioxLMbkKpTo5v9uT7v81L5VyxhnrLRELrEpCYbORu6FMUAz232+Tnu2klos3PpdP2uaJpCf
+s/de3jueQPG9LvlApaSgPaCmMLU3RousWIPn4HQb/83A3He+MODQF8YDmKuToJW19EbvHA39uT+
n5ArkDHiRGQIlNS7pikZBLiKLbjOpuMWxDJbd6b2mzNaL3Xrk7oWj/trpB4jLduWYeeWYGgOQ55r
Q+16l8LS9yP5UH0/YKpmS4rloOR6BNlnFJ4bDu1aWC3TXhkkBE1WQPGuS+n+bS0I776eu2nHIkgU
+LpOMjKK0BpKyq4UOM1KHtXG81NwqTxHM3UMEhbp+iAaV13/nOFiEnR8Ba7W8NqwKOH/7ZLt2GpE
B22ewwK4v7TROXhtdcDT3jg06Cp1rAF33Jjgn/7FAycfZT/h4DxxkTudCGo3JdPsuT5OcBVgPLbJ
ZEP5zMbH4JG3TEPsta04m5cvT/SdcnStMMNiv/jBI+/3WKf/p4Fi5i078SpV7Dtv86s5ilJl9VKS
wtuffSeBp/eOPkbinAfIxYAtu3g6JHth6qMMhnO60T54UlW0mjnKHkjrdzWWx37RJkYtglmhwFH9
8HWmPwvUIvL0wASkIKcKOYdkOsWfmIEQhWO3X92lkptkD/OY/Hi7F5YYV3bX+0hdiYxx2QfktVJ6
EY0yMkC1gZU8PiMhGlJT+tokrVSgri9AxnUPrkjifBJAIDsFQKzACukcZIm8ki2zibdn3IkfQPIf
/29Jtkx0yTLcIGoaQglj1pEl9Xz+5RClX8RFT+ZoZYgoG4m2l6LuU+lw1B8FMwLIdvIUUuvszsYz
GjXLO5R3sfJOlZpbmbRfBRZMNn3DBlHA01HEo3j1XmYGBtF2z5TifbI85RNNmAADR+mCezRECiMi
hAHINKnQSM6vbRlqAuUO3otW2NcigaVukDo+J0nVPOo9LQaY57YtpqL0YCvyptrmNjICkJTDuV1K
aqIHF5BnXgZ0AIIpjJ2pfJp1Ok7ntuiFP3SVo02oqWIxVpNLIZKAZurmMlJ6s0EhQtfQ+0AZk2eu
g/Macl6bMtJMI9/n5G2Vg3zpi4QVKJCYFE4SpUjqM/cXPlnziatGeROJ+DlTD0X4KlXlYC8BCX+t
xCUPAQ3IAPGUU7bDR2RtGPb0sHVEOFet8qblO18DL09lNUzlaybGfLCLzSrU5fhkBundA6a+kf98
Cp3M8re/dSg9VvhZzTwPNvFWX4w7LtP0WFfDT2qn/Hi3/58+EJNgNi9/cHjo1V1KfGvZbuFKaOWd
dksle52ldWnRHFVu08fbMVpZOl1FAcrkWStRDDE7Lok1Ss8hQE5d58+xcOF4EPX/ZNcpZF+fW7/h
92S7ccDQoc8+1EsvN9FOHnCFmx4SOrJToVS6PtIb/suTX2i4FTYggeq7GKzFzk0ydd049MzyuM4w
prmZd6fhv83AkggRZKmEcMjRE3p/RwLutt1diqOjnmx02lqJD6w29BohcTkfstl1gFdnS767PBQO
9zjVXX0SYYPQJ9RI8/0iHPAf44E9TRjIFfjqy5WivFfMXBwireGn6noJjBcmPD1Ih5T2eSoVdq/A
WvyjY8LsHuf+uVXS3pKthvZaDzCaQXiLJGA573FyTtwumUXHfE7IwyiQ4Vp1KAyiNF4Rmn7WkQQv
5PEM8R7AW8Uv3seABJuj0AqpMbGrMAdCwnyLeqhlaPbnIShpdmudKmMQZF1nploYmmqJDzifJ2fl
n+8AvYPtxEhw/Sk0VhWUqw0ODjRt3h/BaOijiOTTL0TlTdwIEHPL6lpA1kFxIxU104ksTdJYzeAC
E3V5CQ9H/gFJdbt9BdL2YoR+W0xWVhhEjjNV5inJpM2zgdxT5NKkhUwc8bYfYteSlu6pTUIGYokg
kFv5kwdmK/h/z/EKnevhzaAFTFweV87/ebBwT4w6uBXOnPooL0qZWuWXrtxCDNBBX7DsFky50fXI
2cQK8Ry06iZpi6gARu5WM8hpmmf+vNUQ6t5wU6amiX7zYlR6Z62aPzFmzYvLHA9R3FI3XVG7nmQ+
poVKIz9kVo8tacVphZbL6oEfZZk111OXJLscTIJyxJxthyNHQhDfBta9gwnRgDHDA0mHif8/RcQP
Im/OZ3S/MQ5g1nZd4eswYqYyug1Z/baKdR5/A2oJCGc8uJ/0LsMdyW9wL+Z26zD2nzUJnZwPjryu
HcM+xWrdK3Ah3HrmQ1buaDz67wAHzz3FDJPMYXTJosjJfoe9H3hB2skvWpF3lLtxB4uAjKadEJXq
D3cBmR8yaRYU1jkVSFcQmarlRHM+WpAQU5cOpTodi4lih5laD5iV/HfVMfuDL4cPnHAj5aYYE0tS
y4l/i4ljSx4MoFsnRqlDuk3EukMjL5ihObw3Qktr0R7odw14n4C4dSfxoqi8PpNtPvqubftlPPyz
siA+gX0lJGtBxJsT3E59i7yXJzwf5qFP24WU+57X0iMsKEYeBScLhAg5jMvngViTV9R15QHHmaVS
wjDD/MgOQZ9qwrQpSItbcWvmax1WV47oLG/SIK4uqj8MqjVkKX8a0MRa+2Y9K9O7mVBgutqgZQ2u
vWqjA/eE8kSjpMaPn/QZ4LoIrRWCCOvOWttd0KAPzd+3gFsaDhHNuUfigMTFj/I0DYp+Z0npdVb9
bUSRqwQKtE0Q2Q9ndUqm42iKXfX4ad8Q8xLdWV6rzudY5pa6lmfN+zg9lTzSSadg/1IYUIhAVYIV
7N6ntcAQdS8ZUC9zD5/1n0fSYKyRyywUsaXynpcfPZQXw7dsYNOwKsldIech85CuNTh4QCmD6mS4
Cb5KZSJVeaThM4X/TLAekjgYnlhuIi9D9mlMsAu9LCnUFHgr9otWlP/9+3moXahEuKCbcF3vQynm
VK8TNvQTbPH+v6FFx00UDukjtdnm7b8EUu210e7tDvvK7m54tXhHuTcOl5WfJzG/80YBsFuUM63R
4mfOGS1MLbFvfu+GXxvIkVYddqPint900yRqBnnKhmkIaGlDPKWPKVdZ1Dh2RlCxlJ2pa+qcotSQ
KMlABt1thyhh2+76wZe6egLaMU4cdSwhhEnNM6EQkmZ5FgB9o2akLxhhTXtoUB4LnjxQf3pcNbmd
YIMxarih3w25qZ8gI6LvGCHIVf4hYXDBP8uLmaaKM71qMkXcpc2r+zf6spTHao+7XYJkBLJAlApx
isanI83+uQgAn6NBoQwdkdGP1Efw9zqaydLSBc0Jp3KB9V6R7VlbNj9cZH/8e6HxFgpsPbORxAF1
nhkrVUNIwUF43dakHgpaWDG/UTZ6ATEph/j/Pigwekf8TST6uy9F8Qu+Va/0U5+ON439R7W9m9Se
J3R/DE1Kcuu4mNHN1ryNzwqEnUt3jlEVGkib54Dk8Ect2tOYDrCg+aTAH+3h4RklFrwm/5opn4n0
qeKgxTOB8G5cNttLn4b78JaRd8W06UhmJt5UuVa6Te4jVIFuEl5/ltYp0LLcHoXwajvUhopbx5ko
CmadwDZmELUpTW8G5nGihrUevzggm/XgP6MnnkQbaGlOH3ygQbpA6Ctg1QKdT0kzkyvwNeHy6C0D
ONSkdZMPsXI2rfmdOSmsyJNJZlfekF65AGx7+qhuegYbD48e4SX/XgLwhzFmkn55EKSAGhK9u/UH
s6G7hg8yHDDx3jrxYMSffwkd713cbGcAc6m354QsklV5AA7lu44QMDu1Rl150t3w1kW3XaDav2Fk
3LVO9kmc3xAH40FE4yCCvuW/70S8Nct6slSVMkf0u2t3y2kOpufdwnXWutt1BmT58o0VX9ewKgIC
swEqWIETJXvipiH6g4ZmbepR6XF75Ic10FjwdDmaDHzWE3ZHMxctVroxCXA3jUdLSKCn+IJb+MRN
djfa9UrR44Qf3Fnqgi3RZz+6CnAUvlesh64ziYMNKDLWTWqHmjLVVU7etm2sAdcxOpxKSBKxT3Dx
dsQcb4JjCHv8f59eFgSfVCp/UXs4k9J3yalMASsxDXy0LUpkC90gZJZDgacLgXDv6uDZYMIwYm//
6IwOXqbc0G4aAy0hvGx1c9Z2wEJk8R47kdYfYHZqgzmePCDbLmagAEAIwpcCzJf0Ctmi92/q6e2C
vvhCYb8ZL4vKKHPFvMjPbfoZ8AlVtk21NQrwDlpfoXqS+W7d9k2GQ4h3aSdrkF9QKQSirZ2lJUOX
T6xKMe7SQP3UXNbjjjli0W6YCS8EXA41pxAY/HKbvjTaFEyF8t/MOUcNy0HKMKvXnVuYMHGFs4bt
R+9H76GISGx6m5khaboVJPT9mnr/BK95Z2jsWZEjkJp36v5IlTU5f9tzgQlof9z0ymyjdTEoaz82
UWAou5w2i02QJD9BfevIz56gHTSosKg2vhMbBGcbrWlkRRXjMbe5bbNjvwZtdFSEFPVwb5bUMxdD
/jBD0hTWuRAJ4sXZaW6TwisKuvX+PmUHffbWfPA98RpgT8ONOcTs/qEyKxpKShebnPPAtlm53Etb
r2TH36gEGexC8K2UXANRiL8a0Vv2P8TZ2nJ11Q+E6XUBhQO6gozPt5M/N/FcOaHrB9pI1s2IG7Hk
bAbtROCo5AfbpgObNMKYjq08tzag1sltRXpnpr0JOnM7VAAjzH1Z2BcU1GMqVW2lzpxmRn1Z1k0q
+bTeu/gGJkLnQroPZUDriHaWt+2TyOPklNAZC+UiyBQw/umZV2pB6mwB275zgMHH4M+Sg1ber3Px
wBriyY9ESQg1lV+eNKSXd2oCLdO4yjWIE7o1oTJjLl7Wb1EDD1HQfDA4OSIeWZm8+ZMvOHzn/dd/
txhjCvI3YkDl1Kgf754RO7vfl/dVddy3KvpAqfb1GRD7S0+AaZhYN4poPIQU2Pd/MGKe/0zBfR+M
NUuXYUYSL1yFBq+zF0x7jL/bKVih5zvgFg2CWA2QpbQLXJk2xQrnOHXb/qa8ie2W/fHfLgxMBcal
eQTugiQXIe1MQxbup0AEAKrR64+LfQxan6ORpid6DMfqhd4aj8hvX6vwd5uLAN226auG8Pw7bn1S
/Sm7I/1aOvA+jnN+aDlIoOVi+h+Ih9Lv5obtATKgyTHloGe9sFmWQUoe8qCr4gsc2AK9tZYs28jk
ocM5FY4U9bm/QBDHhcop7vufzDRDPSA6OBGp78MdKWM3ofNPr2fEVd/GPTkCM5mCKzU8nYTL0rCz
Iw2gaGHhMk2LkcHNRqRFeFrdLZ2iPZWwWcPcoRtSLV2hfJDeDB3YWuVQNBYGpOcOp42DEJdnfGeq
Pqj6pOcIfIiK3cTf5wCy4mCGdLbbyv8fFftyJtj/kbcewe+SRW4jP+S7b4RzRdWSXurNFGE3KQ/h
Ft2U1I0VdAw9P/39ssveLftzi5ne4cmszAi8I6DOXjF6LcnwFDRMIJmew8REtzQvk9mSmL5SOWQX
6dcaQVOPFyv4bZDkxnivcVmk4rE0L6cz33aHkplr6dhoKlyBON12AL9EwW40CG423QENAJ7qHDvR
I7YAzE/N+mDKQywYgniwjl3KUuk2OdE+6JmWUV0YCyXCsGQ1SxiGhJ2xUDMHMwU5zwEwux6Qy+Xw
N8fkcqjWoGPL5TecpO5V6+T22azRbQc5wHw+4je0dM+nXqjjwls1WU3kXSBnXRaRyLhrWOiglN5X
Z0HRgM7brpEGnDDrAZt1/Nm3bfwCTfaeoWC3hQsibCHUg5btn+DGRz78D7Q1uEu6UrcL3F3zBqJJ
K+8Bu+mPvqQze6fxnGm0OJtu871g6jk/gO208wfn4pyKK1H0X1IZgqTHOM1KeTz6+wxbadp0xmBB
aP99yARM1WtRSnVCL3PPGg+F9AV90QPKZwqBQMmKBV5WXCcPcDAzqk0OmDz3ruTF1EWcBhYJv7iA
6X/r9utqCQLoy0JC7p9KKa1kG03nGHE7m5Ogy31ilTtxRaYkMnJ1z+qKQWOWdpe9akNQ2SBUxXVv
Sulq3Pm0fVB3oU98N26RDSwgSX+usnaHriY3LvsFNkkG+MKH7x3dkMgyZHzWlpbz6U6Zt4M4zun2
77y3TsYK3qxm05JbeaYxoXQxhrYjUABux+q5gh81kLBH57opBLG50dQuVrpiIMNPIWH3f+eAmwNw
eClKL6EgAbFHfsLQe304B6V9iiGaFBMm7D76P4nWDC3dkXs3mJWmMBOxCy+I1t7Rxh84OdhHJK3J
GlvG56658JLQEPXFSP6ZAapxA+gCr5Z8wK5MY8VDP3lxqo4U75UYH5hH4VTp1cIQ/WDusulHguLE
OucbYMEr9Ov1klxPxe73TvAZd6/wFW1QZlyhsMhMADVakc6E8jPjYRL2f1XMPXuNCuGwyCe77HB/
rSNI1UjTMrP4VwPIIylXZp8eaUwXRkhCseT2padABWAGT9FUORdhaVlkrSH5GVYT0Q//H6ewoH6Z
cNE081KuhoenwvSf3ZvOTevpMAYGohsy6FVbDkbxeJGQnWU9/HO75TKUNJYjD+eRlvKuVRTO5kW+
EJR6eA60a/pSFGfyAhq1SuFfh0nZv+LdM6+kV0n3v8iO192yZHFi6UkdrzcFaNxSeHcCDdpDdVLo
P1SIHdoOXE33yp/09qtMaboFALU/unPFSLeIRQUJM4IkaHsNIkH7Gmm3G+bw5gKu7nKYyn38BWd+
PeMpo/4o4Jc+7UdWLmVe7LAVKWyVY656Y2UlfIy+b3eryUPP3X8r5UuUVHPtQB4ppNAq21kKYU2I
Oe0mnslfzblSefc+g7/wkiX7CqKal7IIJGy78EQOFCPdjxojl3bWPl/jbCwMQml7aCc/1XXEq1Qu
8oovqcfMYl0REoUxrS4Hoajl3W0PAkgb/8scjKNO9odjQ/RaHuMMQRgPN3Emxtz2NfeB6EEvqCai
O9bF8MCbURbTVjmJFtRX5Uj1MStWxuHmhk6kiavhVGyBSCCQtjkaLGy9xwvQDP1ZfWfGCzHhYK3C
/TX5/6T1nPcoCNzkxvr77AefWB5NmL8h3+uNL5+KbSNdo4ba6x6R8qN1kVrwR5ZJN/wWjBtIsX56
WRPCCwG+NyqHTMJPBuhI45dA7NcPmJy2LGq4a8zTzWneXIGFJdnVE+W3aPe4rnDuEkJyKYEkwQ1U
4zswBgAkGtGyNzawLDG7tvTSesJC5sZeFcJphgVyRAtd1Eesgx+mFHVYYUpCdYiJ6HfHRUO4sPJq
pSyF4X5wnqZWwZW66EZQEMqbwkjjIcMREaSqcFqV7eyXi2idjNlSksdnfV8TuZ2ykvjfbku+3euI
PIyYQ1qyAabLM3+MmhjegUsqED+mlMwfBr2N3NvZmpOWuXRgrVp/5R9iegYfD2BL02MKQ4P65mDJ
IsySimbFkTE8zPbvpxBvb6mI4CE8XtbhIPcgQea2FAmFU0C3DXb5lSbix7NERfP4zc+SstaxCEA+
GNou09TnXJald3t6QnpALFyWL/se7uSM5LBtUfAGt1M+SMu16hQFSY6lXuBgknWbWDk0IDMlf8o6
tje3TwRjPr/zuL4k6b8cCE8tZYP954uO0eHYdrj0frGNjV1lLo9RjcAgzUtXhAtBQ94NM0NflRnK
+uhuq5MS1hSsPCfPT7esOnu1C2kbUszHACUPI3dupP8l6zno4S/6jHX+ZSJo5CVqAl94fwmZnFHd
yWRq2SeN0J+GQxzV8cmUg+7pi8Z2GiVcdKkp5XotY2qigZ8TPphIar19L3aw/60HJxKYwPGrbSaA
cjgizl5fP8OEv03cfmJV6W80IHZ5Drb1FR9gbHdnBmrZV9cl2pOb9+rOHnJcw0779ehGdE2IhBg6
mB8vyNQpJzodCB++LlTrJ5kxeRhj1yUkqw3/WsC5SdLEV8I5LWfqFpVzx4KHwsLplmku+iBKuokX
PM/2am52595X+Y764/UfIgIObQJ1RdGbQJ0PAu0k59zIps6xREdqRLqyqLoes+5essNWWEN88nSN
pQnEDSJnNQmksvtZ66Mwn2ZZspi4jn9dAph1eJhm1oRcxEIzt0GBV32L909PoYjvBUxzbLPlOh0h
cvwA4HklnTLQ+01KbPXmhoUKMl2nOZsE6tYUaUutHnhDlRffR45YU0kfQUrcFmTdlOc2BS0kXtmE
ItBSeBxnMfUmd0S1eAX7ltDqxCd/D1a4HlXdTPx5GSnAE+My69HaJbh+KskA6AF/GjxkiKIcbe/g
AkBKv6Mzyr0nJelSWiQbffCngyor/nUHc2cUpD21vfCv/Ms/G1C9ikNf4cl6oQ+AJRI2WItQXfZe
Ro8LV5AFv64BtoZ3+yWm/H/6unp6lTgDBOd7ELw/TAO5bKtWQtY6dkvSi0nGSZLRg29GTzc89TVo
70/ADhIHR4Ft5g7EoYoGESqQbN89DyJVCpW+zsCTD3OpcOMMcyY7NqJm5aFA/pup7RqoKdWXU6MZ
QE35zhUfKAHIWGmuVot9+CR4K97gh+RdleB33vCsReEuniS7E0+CKSgzV7rGzBe7eKIBFEdrt/3N
TholbMNkC718uI+aOGY7qsJEyaxg9DhKV9Ra5i/HEdw3IWVD9LhhL/NAL8JHeKECFJ0zKgLYdHFz
KKayEaWFSAAut4Krru7GFTWriXIYxF9prVRadT1NCc5/lZM+GXhw9YMVBp1Bmc+0KScwNdMrJH1c
lC5ZrYJJekeZAgJGsyotmaE9EMNKIq/R5MCDF++fA3intGYhHzgQUTnu8ka//rEkxtEVBpzTtK8N
YzrhQGASZNwo1Nl19UFd/PVpIEFIXoTlvJJ1hSH+0w4vC/hO0Q==
`protect end_protected
