XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E���9~aڛ�	����־��WK>z���h(�v��!��P?�/:�����������<�u3c��%gڻ�4�:���wc�[jz\�v�¶
�n"�y�L/sc&}����Bfؖƹ��s�	d�%4�Kx�;e�!�Q�'�̓���l�t�x�Oz�=�V��5�p���rN<�Z��=`3	���P�6���Ţ^���3�a��8(��Rl�=9`F�,o�V:��D^Fh* ���V�R�5 �v����+Q����-�ҁ�C������ÆC�I�����R�1lܧ�k?ש�M�LA#�q�}�X���~�֏����&��=�����*����� ��k�*{�s��9&�QfԸ�U����k0IК���	��3'����Is�!#��̖�/��bY��\˦��r!Hs<I�A)���S"*��MU��;x�S9���Q��w��Bt �v^���gv��@��M��9a��?��4+�%{p�ک� ��v��/��u�zx��i���'QPV�����yn�e�2 ��%d�Y����Y(�9���bW!����=5���uK��-�be�L�Le!)��#�B�
¸���2F��Ts�n�j�w����)h�l@���4ǻq̒����g��Kz(P淓��aR΋�6�F�J{�;��a5�Vu8��=��K���1+>Y8�[��"�{+�)��D�]@5�{S;8&�e��w�m4�
�&��s�rH^�kc�S�gXlxVHYEB     389     180+�T�d�z�$A:��ә��yl�9xJ%��{�a�^7��q�u)E�4j��v���E�[ ���j96Y��Ԑ���qw�E�����A� d���q�|�+��3d�K�Y��F7eJ7=lB��(,w$k�{��g�%Xc`q��2�7ʻ#����d@��ӁĢp����|�{쓳������>>����}�vEpQ���Yb3�t�r�r$���Dm�7�mI뢗E��������Y,a��L�7�4��N.j }ڽ�_�_ � '�w#�FC�|�d��&*����뇻�x�O�T���%o�گ�[6�~��c�BR� �Y ���ᾦ��[N(i���Z�Z���>&v���|�_|����o�����Uh���%