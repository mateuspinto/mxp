`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
WA/KvEdbhMDH+jmWvmGtz7aEDLmKsyHu6/O0Vj3BnsQOeMOBICJXkk4XnImYogxeJgfzuoNqD5wr
NMqQT/9KqHG4+45glRz+1LypOdXIzaJ+EvyhDBPD7XIEZBQgwf9y/GnQ5GgrWF9tvb2NSzWISZEH
ghVoCoXo8xgO4aBvojzX3E2+SCWjCKj+2UKZjXaiOtxno8WHjEqHPQs7kP+ScDNLLoPniBgo3d8+
uYuiUoYv0OYGiwmAaNyF4d/lmdTqaTonmSZAlOrCgSCPVskZMUQR5PIVPs27HyVuekkDaKPzYH20
ciEKrxgyMpUxp1Uy9flCh/TwnQljxNJzpSE7sQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="OEJcJ3CHtt1FXQsfmGKcjOjfF5biLmn7sLTGUvs4aFA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26128)
`protect data_block
Eu2bJvshYYGdWxGFMv84EJWXwNwuG5RXxGfyVm2BURu0ggj2DWfU+b9k0mXWG2/nCvkIvLDgMiG2
GgdYk3B8ZpE+tG/hvv0z/bMuoeNNuxXPN6sjz6wrVboxGBEh9RR2yiDhDe74QLWjO+Lpeegj1fmG
xfIRiJeYef4MZLhzIBJLWtaGJQ0IKgq+6L/utfew1/6L6IunZTYrY1de0EUDf8p+OMIU1vk1vkQ3
NMfrz9jcNbfP3QVbAt3ZlXV96iMBuScEXUF9HC2ArhDzYyXZ37s8OgYiGyCY6BwbyzmaiBACQGE2
SZCiIpNP1xanMOkjELHLTcsAEaSrqtmuQQRcJJf41D8FAg2hGgdN3vWKKOTV8MnszTk91U1I5hDu
QTBR7j9/4PvhCY6WrSopHHmc67ip7v2SqB66P1lt+zAxal6k/aOuJSc5d9185DVd3+np5OG2htOp
5xU0MXSpLebi05SQZaNk5zmu/xywSeH/wVk734tFkumPiE4o2+tXp+2WUHmtIC42lqBweuuKsAgf
nYezK4fn/x7OBt5dSUGjwDGyIxpLJR5LBbRKwsVshnXpXV1243HugauucZL9Mg5vEjYVcarYPSX2
Dv+QqbnN9GE9k1E88uPz4aBAGd0FRzS49OTuCv6yb93K3n0+TpyS4xQH0r3KbmtBQT3KeMTaa4rA
56SH2oQ4MP8GqtlfWKrhKwUXqBu4rbwYvQY1F7kKwmnoP9uT7S7iq7lyRGU6v5MpgThjGj+9Jtg2
vR6wHHAGdj/SzS1DusOkhZesCe1RlD06VYC6nsLCLZkM8/ZzPrcLeM1u8TrqDNyv2g/0qugA+Eql
qCnUeOphB3Ijgivi9RInv6QaZul0zJeZnRTWTZDawdCMHxep1Y9HKwmStHUFuK7+tYvDn0Y8ZDH1
9jqWw1MojvKteDW6/qy4o8a+TEf68MYuesP3joSU+bggGGVxrYyw/VLmNVfM9Zc6WgwvNsRyGS83
q7ErnVeR0uUOGyzaz2WfZJ166ishNrv+dkx64pP0SyjVv01gARwyF0HUeSs/JtLwT816sMP4maTw
bN+Onh1iY5Q0v4sB4i+6fedFqmByepQDWTCCscKAxIUx13tRCUDejLVeZ7K5GfbTr81fW2fsHdnG
Lu17M4atGqxI6jJx9zniUAT6IIkUYRh0HZ8cpoF3JAdzKUxmRG+5uQVQOce+ext7DISGmdCont/t
sqEBImiLbw3YkiTwUzwfpgARDGo/rnBYu/WFAdbnVUivk8ZHUXsh10VkgC6zhjWLXRKNqikq/b9z
ed87um083uOOqicjVxsbvGmKtesJlnWbmGlADXNgtzbQrkKUy9MoH2YGSejzSuIkUYsr34ovHQDZ
7T62f3YpTCOCMQqRHmgDyzUqmk2NLap0+e3GvGhEe0oR1QZTAF63VHar3xfhkBUcEr/oF4GeMX8d
9ZZkNrcrc8O6oCBCxDf17hn77IoOZaCUfvRVElK67w8H/RYfo799oFnNls51KfHWA6gcklSl4lB6
Yk2sYBG7zmwuk88iXlOks1/B6+nGs6YAtqlBR7+LaT3AUi0d0DVWouaKBNuw5kaVUQMYCjVtseLp
UaYGFAgMxFDzMCl50cLrsjOPY0yqL2dUWu2pSdqTdDB+alCFlzBWfrWquJwzywqLWyQ0NbwU6+H9
mUnhLex7q8M4kQuHnfSXtxDRr6eSYsbnK42rFP0ARdwXvhAQOTmcU+hOUnFDh4TAJOwutNhjShCc
TPn8Q3hwqjocE5tH8UbKcoZWx09g+aGjVRwffCMztBJoyf5wuyJTtU2VeJFIKLoU8qtlfdkTLm9W
KIdj1G9pFxPf7R3LCeWBHab0aiTegedx7DAdsr3Q3xZUQ38qiQOZhm4OpQqp/2l9aMbm0ZKF+U8Y
SDvgpQHzeO9QVJTHAVWp+7OGe3cnnYKpPdbFZidPp2CBu4EVdNaE1gcLyB/r3yt7FFP5d5/SLua9
QFq7UWNtdsMpNwCenVj6IlV7sAn+KbAyve2nzcmVQNSWkytVzVaYLRQP6CC+rFKthKaCmZ9hvQyd
1UeJG5ILETcUufbJHCPRNCDsyMqON/3aWb2K1yOSBPuM9lLhOdaCcvu8gXwrnMw2PmnyHdvmqU4C
vGipXPgMRYXbRu55FvqqY6TlsWNmNas2QYTZkO+f+05X0bEPP47zER2miTJFKyi5IhQPTbgDtIEM
bczX3dfkQihkOsAjB5V+2iKo79D8pE99gDEMIbDvOn6LwDaBKaTlXS0MUD9Zvh4f0GmcjG0u9817
g+8vlZx6EpROS9vcU9v69fO08b7H8N1KojFomibwqfd/YZGysggQHiOOwBKaDcDIJZZlqb2WnKZU
XUD90nw8vKVybGyw7/P4IfVjh1zSp2ilU5RSy/RU/9FjkwrR7+01hEtJxjWIMlEbOJOpvAHKH8Mh
ZwteVPKaNUjmhboNLPipAX/e3ESj/fHxMOjpceQulN39xKK4y0QD0Zi3QNvCERpKTK1UcaAcY1x3
QqzdEhL1iTNxQGkse3AQwin7YxK41A5SSkPjclpMSJV+dRgN4Y6r38gFvnmZoi/bd6ebAxK+7Bx0
U14Dm3tbM2o+PXRjHyGuTFSke2BIHy1pdftY8h61YiyZCUvVnu0xH7cfz29Nuv8lUVdCQ9ZFThy9
CpL/B43xSrENOqOs2xqapuyPjMz53QkL7E+pvqMYyBMsBr/NJvdMw4y74dqLZG/jokSE3ePYEtWn
MMCaZYSh1oL0sXOmBqZEDPBD3uo6gTlHhANkY/ggyXQiMA8vHLQ9cmo39mcDhsf5dvi5q2zBE1ZB
6Kfz/aGq52fxpSz1ZFYt+GvrO0ZQkIeQtmMJyrK5Hg+KmRyrtasKVP0pXQROHWLnnuHZ+d+kLEQo
CCuRSdK4/xl8PD+C0lLfdCOR2PAOI8CfDVO+OZuPGQe6zmg8DJent175kBjixciI9JWs89Pn5mFQ
WHS/hAugwqXDHlIz65XI6dyjFzjlX5+J2oQopxFdrMtbkrZ+C2svKIgtKu9EN3avbb5JKCsxHRYl
QWlPmhpkC+6YFeRKMGtMs1EDnCFc3KYAKcbLMy4MCayVndzUYuuMwR0EA0vFIfNOdvTQ5fduFoMW
P3HLkym2ctzibmh7PyMn/ykIrxl6M4ZwpP19P9DN19yxNWTtWe/CXijaqT3aEbSyf0R7LSFUWmGP
SE2JrUX+49pXM3MqbotCtfbr8QGkhH+JkL7OXWfgdcPdRkOuv+icPFC+TQ6aKHg9UJtju56MCWyS
2gTH56gBGi05WDtq3KgAfhw8yzq9ATShmQESbekRnavMf4mNulHlNT5edb9AEaxIlZsFZPg6spT+
eU2SAzwUb7bt/UFzJQ4h/zsSDlaSknzTNHJQfwRazPIHSbdWR9zGRfAIGlGd07bIAqdSexZGqCgQ
2sI458aMZvHt6VXRXUFbxEZmSRneZ0AFUa/XkJ6uZqo/2OUAvriwoP9/SoLRMU+P3LBqrcVsIoqN
p3/4Fpl6svScagN1jqBRpchKxnFi58oc7abaWSD1InjxoYySQ2ZDa8oughOm4B/h0EmBrTnMQ9yi
KeBkbuU5+LAOV0eXfuJ4lHP+aDwUDlHZ3hsyQOlh/SI5NmN9OzgIlrtF2R07U3nnHDj7VA0IuD3E
Xjq19BieH3egMQriWnZGTiKDUOOaD5SWbyXGEcc8UiTo7QpaDxbN6yARuUS7SLb7ZAmpxokcOJTB
yCgJQHHwM6cWdCpWw3nZEccv9euV/MIzd/pMx//SXZzsQ5CVl+W5NJHFbckulVhu18syYBAM8ZEr
iH/dkFcw3K/rnt7G9UraIYUdx7JTNP0iZy8B0Usw2uzUyKJJH4d2sOvvFoihmVrOC5gVUl/262R7
ylBZtpPtA3IuTnuhh4vziNpilkuVaTKKZwhcFkL96oHjmHW7MHrMHxJTxoemAG7wpXqRKYNw8WEG
E8nKdJpExf12SfF+CVSp2O3tY6tZMMkDlZASWXaFrsghvuc/rO5pZrENd8NNyBn3mvTclcR51m59
ehAc/HNCVK/b4jBZU3I49KcuOHWTJdtUQIS2c3ZpbuKjN3LIVMvP7H3s8ctv9FLe524TJSD5AdOP
v0mvhIpufrpLNRWtryhKgH3dsKXOTrwSHVFCw0rrulbzUyKi2JfDD9YeropsRLweJUcCpCFq7ymp
Wba3YANfVIk56cd5KiSVzpGlxFyQPXl7W5gTZ1rAVTASIsWVCzv1javw2bbU78W62sMjcb5Yy3oS
pjqsmV65Zrdul4R1DDXb/Fsjk7iKDhBPHBzju5qyCgUYFIVhW3q3Q9uY5mhDGVeXL3qn55l5W+D+
9F9BFdtlXulxMiAVZ4vY06/G4/aeh8WhLxRMOCxaek023ebPzErg4KUqRqm9shfvHj1yx0dOJ0z8
2M1BVtJiDp9I1f/fYvJ2pFsKCvmo1XYv5wfHpUWPoi9r1T7ExgtyH15AdcQaM92uCqCG4P8alJpz
MvtTSsIsTGjLpyFG64hQ3OrLo/22j9FU2kPEHIuWo17EruxeADYeaW1aBjb0Li17lxZOpEUYR4qA
x9JLDnpjFkzHdd5BxPXmGXa8Flo/WVKUdL35IARuTx57D/cyK/86ACqfuYloG3bhvZ/QcIAYeiQs
n5uPa5cSM6et+3lVf8ebWzhj8vKX2Oc/Vzc1TiMTHxfe6EUXbNzPyJaERL/xpWY3pKhwYY6T6KOU
nhNqcPHAQ/BfAgJU3yeeQ6lik6M4pnt2tI6OIHmHjeiz/Txp1hMgb0YJSew+iKNjcn5mJHTWlntU
PGx4lVGHH9JNdV6ikC8eocFxTXxddoBSp6qzqy0ZIgtgytaTvIAG93FKNbQwrSPExGaKedykCvhX
ihP8b2nn14t2WTQ2fFRnpwkaYzRNFEid3AcpWHAsv8zAQulN4Zq3QUOuHNmyI/up1c7/mlCUccgn
InYv9mAAF9Bq6KmbrbsXGqO+edjysU27mpml9na5ACSafQRBtGtnTHJ7AUCn/Y7HVMfJP7MhpRvJ
gAuYm/JqCQVQbBLKPvgMsS6pB84n9DkHa/GN8fUE2l7RleDVQAFCPskazk4I5VhaDqBP3H0R+5bg
xtQLUKgSaiTkZ7KirnJoLTmhln3+BVI/eiQ2QjFA05689RkO4HYvC4X6NtVEhyqdCmDC1RQoz0r6
Z/1YBNWRn6MUe9ZYErJlQoiqrl8buJO2miipU6uIElu7jezpymSwdjL69HneMqCQ0az3nweF192k
qop+oHUST5rpP9zdYJ+BDpLWgAQuNKnmcoEQcCPL5IlpTnU0/Zmua6nI6EOPy6Zy/srZdQfAKF8V
+ZlCvTFgCnOIvLFbcsh6M4TALUFNZFZ6tjQFdhQ1dq3dK4wlyINFxS/UJDt/fLRRmlMGBbiZ7Cfl
Fc/4oek07kj2nZ6wTUR3q0muOBjxDBYMYngO8wc3hMbA/o0lfnhCE7EYXXPIUKK5RIOwr2URrI3W
NCQfyG4U5YkLQP0qee9/GbR9ZHLKf6/+PFFvf/lk38SPyKXKj5vs73PNvTHl3VcmIGfonMj4dABM
cnHD6WS1/PnCGqDaUgL5Zbb2TLd3WzwXZgE4H2nqy1d17XvsD3QDqyILRzS03U9KbjjRxLbrQnnt
Rf/wHMp+1rojYg3SD0sD5Hx6Wzc9KmMe0scMNYzgemng3JVRAGhx5kJNyPRY/UMakXDRSY5vVeYn
euOqRffiUDXQD3Rw2s2OBHLQIBCPBbENzny3ONminUg5snaCzkboshd2gh6S9e0Rn5cEx2FhOT6P
ebJgNBJ3cDummYOEE97ALNMGAOmndRM8t5eI4mn6g8lMFYm26t+92CB1b9FgiLzxqarCnozyQKaz
rrY6i6MD3gHEkLcfKrBZOdoI8IGJLI4KnJzOLYmCB+uy3yX+R44f3d+kuOeOed+SUW3x/PkawDwG
tPQoZFEGat9P9UtWzPYJOWY+UkRVIcYPh68+FGAc0vfkbJBLuqdtUKgDwIbaRLWx+oMF+hw01Ei/
+jhZEqE3zesEoQS6IdjfrSmlhnFO9CNOfc4ho8mIYxt8JpegkWQCUxC+f7YOIfgHZUuOH63SO1PA
C4CugcMGcFCshmX24ZcoaZGf2GhvSN0jGlFg1JYWQewWEvuULBj7BaJLS4TKODVdXq70d6BXzIEp
X2U+LhsX4bsutbCvO6aKA0n+Rknd+I6y01XNQPtrufVORnXiGnBCAHBDTzTcvmVyx3Vlgrb1Fg5Z
drx4vzMW+znvEds+eZiR2oL7i6NoOvH6/KAdqdbspQTAbB370lkUQN8nrkMheHovAuDRR0RmVVGN
L+3hLRk5Hx9z67d0weLub4lgCQ4+tz3FgOMbJlfZOnpl0DU61KaqdE+A9U8WSZCJ5jZO3H31luaZ
YbN5hSsG03Kh86X/KkvX5kC9NarfVm+K29uOYkfvtGmTPrSGY5r6xWVD5RaOjKyNTYktzxZRLzKW
GTGeFr1817SFQhgWqg+TQC3eVLKIIeEj0xawZ6YNV++pgO1CsP9+wNROU7vwAfwiBLl6rIRV49TM
3RmYqXqfvRjUQxwVhrd0skjmm+mAKS/c7IOB78F+Zn02tBafOBb2CjbyB1yauc1i6StKJTMJvyBR
UxG81VPmbqZxl5VrRDlDTMGPrFoXiEd5xaubrMVHe5chNz5g+FYWDEku9xYsdb+tecb/goxmGH7m
F27TU0DUl0vhpjlsdHDb2RAqQyJ0eC3obcW/ri2TCd7xKj5lw1EWlkefSX0BFXyjozVg2zGxvIGv
Cc6b6bndGg7p2lRc5NU0FXkqm/G6HLYvJDBJaOrTPtpYJPa0C11cht0QQaS81daWIf/0MQ5Epj7u
DBOm7TQ3H8KEsVSiqtQJCLs/FE1pSqeNgOA6k9HqNhcoE7dJP+2hUGA+dCXYSDeoi2fCwHfRrZd6
R+cJt3tTGGxsTQhd5vrIs6McqSxckTTjA4Jy2d/QRKsPXPSh8wX4DRF/Tl4KFf4At6LiPDTe7Jy8
6Lb7Nf0xoosmVgoxLmHhyZV3cNw2oy3VwjglCedzz8zxY1YvA1GtxE+YOoLGSjq3BnrBIx7S2OpH
UvnMrkdTRHq0mkyuxj3VmIRvv3MX3cLYktGhKbViONIkAV0Ixgx1N4noIlGBS1X3WXNeCk//1IOC
8MqaTIPBFeJuC18Sklyoia2GyzqqlacGUCU2WCCXfI/AhvHbJZbIzfzz/TXH6gIgPuHkkwvQPfX+
7ciH0YRUQhGW7NpIo5rUygC4OPoPMgKgVmUwvATDVpNGXQHaPuAl31LzaNiS62JDjnDN2sSss06Y
T4IRWlM+Nle+E5IFVOs7aHY1frXfl42hy08qYCKoHPU+wTSzDDQnt8eWm9Vg9xeOvZA76JfJDZ1U
DA2oVaR4D3wYwTlP13NhOuADMD+9YMMe4NSc5cJlHicYgqsoJuppmbnN12Qkh1aBHVItkVis8PLv
Lid4N7TDcyNt9aL3uuzjtXhZHhHMAZJGWgjSFWy6PYcPHYH8y5/dy0Iwlwr/rB+iIGLZMh0SVmji
LYiTpuvIzK66tUjD5NLv6L4cmybv4xjXfOcYkJLIjSaqzJgJXIa95dXZEG9Apgj4WLMGS7L/S1ik
8oSKWkhaVWApdwmL+vmpaqOQ2Y+j5MBVISVUhSU4LVXX0ABGrD2dMU4BV4keyqsHb2NMd94u9dbO
WcPkJUtfjMEOBPXUbCDdqbbAlnC/6Xt688rrUV4gmRq2er1qbTzWtFUf7j12mEgdcnD3tLLOPPXD
PkL1vjc1MtfMHZh0YWLPsGunafLA1+rzdkcl99g4Qpf8edaqxn03xvJePNhtEyLdcGB306PRzwjC
t8eTasythY1rCgCPeMty3+UMiMX11qo4uyeCIQrEf/RP8REcuAeJES6HKVImag5DKFDmQMJUG6hV
nsV5sN5iNxyBdi1DJhWLCt6voWv8SxyvUCgMq1R8/KnEeA0dVXN5MFJRd6rEPZc0Mx3ZRx1nfxRy
IxZyMyg0xGws4WQQ2mHCyIOkQB4YHw8GNaEnTJ+aScHy2QC5jzY1oQgQRpv7p7FRaNJPj4fDpPZK
t/c3dT8Bi4jdO8XEyON+Z29TKOeXI/c8wURj+I3pn6+u97Edc2d+QSi8jQlBuo+UHf/C7JA9bUcm
aDYNTqRdK2a77wip6dk+QQ2KSUJpom1SBVt2J613fQXAZZjy3g2Cz54sUAzGokXyx+rdfhlszzWN
WwhIr+H6gdn9dkIgli1gJV6OjCzTHKJEiIzOc+tAhxO8bY4PuPS2iZnb6TQIiLiwkJ3HtURL4nMZ
uUNTBwJQ7cst1eyQF5ZzNFcdkL9xVqCrojvdnGiBb8fQpuuyOqhk57UsT069e2y/r2FtjpUQUt5C
POduQcmhg4qtY4lLnkkx9dlEcPbEdPV+CgBrf3plJHKOwB+3b5VO40eC7kvnvWB0rT4Hf4zV+vqx
YZ02tvCb9yjIbamELGmNqHtbaS8qmWEhp+tMQ4hiYoTYMZEtZfv7yr5fAFrDu+JQNL7+m2CYCyhf
YAnz5KwmLm0zr+xBJspOZYElzPl3ObMHt2Rng4g9V5Ed+DbcK/D/EJkA1az2At4geWXIc9dGZD4i
3tJW/1tlX8Nx/rh9C4PpoB+F8BtJ4XSkbzjO076Rl3SNYSTrGpIU7amwchOX3Mm4GWe/BDc6zabn
dJthE8XwuGy1QxggfK9BYDpgFLPeM320VcyxaAY1NPXAjqVv3oo444kKsI2Ih0wmy8gaxJEfTLMb
sEPLpZvYDqhOndgrC2M74Db4apPNcFgX/8lObRJ3dhPkXNvkvZqRXlgBdmYe8WEROqlAs727Gt5E
rncKwjbDfziFrLZgUBZWE7IJcwe+H84xq/8nQFpZw8LpMp60rpCCUo6ribfcfqZDUfQ+BWcfWnEe
ov4xk8X0Bp6h9wIAiqVUQ4u3xQbF1dGOtaeB+TTOUC5vCMk6uH3w3iAkdoh2gFgv5IDmO37MrrIm
PZjqjXeQNg+DSSRtH+4phtNrpB8Iwka7PmlLhPlCe2h9HvK76Shn+izs2MAKj3IYrrqkA4FoFF2A
fDekIx/eu0rItyXJkHj0JcSdC2yobTlOXOiA8OMKkSi/mdn+VfGEpHzWcz/IxnF5dZJKrnZFNkd4
dDyc6STRoKHW80WDksyzbeuU2ET2USAsWy0ghi2wBXJvSp15oqz3kdQYSPSXQwQ+lebMZrcmgMOJ
xzdQO153Z53RLBhVPXF9JRXl1eVLumYgnBQ5vgy9gRaUAhELYUE5B2UhsmjDPxN78ldpr/Z/QlfS
h9yZaTh7GLu0T58eqhT0Ay9ND+hSTLRqJ0gK4Owbb6Wr9MXz5lWEo7lUy8Ln8sGmFPhEKX34Q00m
7HjfGGTMiTstY0x0lB15Yf//hkyxst+aFUDyYiDuwf6sjblu8aT7jJgVkwmYXs412r+uTYPEp5Si
EARpbxtOudT5EH0sHH+/YZ4hUr8cOt8XApqQCtC89ecu6ffLzgDFvsKu8zeq/3Q+ueuqDrML+60d
993dC7SwY1sVTjKvrO19dYcW8bK0azFtfJcITwpY0I01i8vC2anBDehP/eIr0gzCFTWzruvp6qvg
/O9EVAX6kOtTBRFoStG6sKfaJ3+JlKSEdL8H+QyQqLEI7OAqAzvejYznf+KaLrI1TGoBzbLU7v21
86Ky84vsUQiOrKF0810xj0OOlEPU9j9LYkz7pudXYyWsa8jyrJigaD9PC1qhLFf1fhvzeF+QpLIy
SIhy6h2jJcV4vh63H0/P4CgNy/pkAej2/36bwrKuoWGleiu3RKxaPEo/SeNELb0SHbg6/FSK5PiW
XgV6CsU9GWK0H93CFpfXxOuiuHtEH9MpVtOHn4vcdr0AL18F0KYmLclbdSBN/tHWN3j2a7k3LtvY
PYx6ARI6Y8HiMB0ntX2Bl/a9eWIJhkKDM/iBuAshhpstqZC5Q3BcMmxVmPBdXHW8o575B7kwy8yC
mAw0LMmqcumlYlO/lwseyimCSkG/j61B+WjekOww0WmuYJT6OPZzpEKh1hHusTv08n21qJuqsxjt
xpopA/ig0qlhaJSIL+wnD9OGRLHertUlf2bNlWV+wf+HKvSDdFM8TH2X+wf77tKwt52Zo1yisHbC
tbiEhCJ+cJreLpqMuJCg9ui7CjP+qc/t24lWfC7nkU5LhN1A/EK38Nu1GSYyf2B/1xfZZVKN/I5P
WheXtfW+RUuPK1E7ICbiX25fJukJqVDhWhGJgpJrlBiEHpAxQgnZf528ZGGUXWAU6LM4DldYL86E
tu7ROl/sxTl30BMPqJ/hjFYsYNZfeKAbzmpzqv5p6zLDWk/DpH2szR1Xst9HX0H8AXmvoiVWX5Eh
yik/tl7lwetl6v8JKSBsrAZTm+P3b57ugFMgcUdltH14gdrSXeUrnDA+6RY16GLaIBkSMQAXKCj6
+CY9HGF3vd0jKsofRMTpkslRzrXMbLZl1pYKKZL9nQyRFlkpRm9q63lOlIW0kMhPjFfBnztg7PHq
RdAhk6Gdgdkxi8RLIBP1MaeJ66zUqNiQzZMo/mNJAJfxKmGfcgc09qVpygEXS9GEPmMYc1AJoCaO
SYKdNLdQLjEvTk4IUG+jvX/kFC5nbPmwBJ6+LbRPxWi5kQ2uMpVKCKyXArG5TAsIRjReMK9vi7YN
whj8T8qACd4Md8DSscivzmQ5ejfutJ3fdFzpPkpCoNt5Iw+bwurvXO+q3673uNVPkNEx0sr9315G
mG09xEnx7ZIilzDm2V89Uh3DQ7BJAgSoT65eagq92CxDXyX4Ir+Zrc6rJJkEaD40upWbXW4yNzrx
+674CPo1p9wLYA3SAukAaSrJ432fmmzF3UtAhQ4/KmVbtO9L6PNnxR/MoaXSbkpNlm2CYreqZt6t
+fNToa2VxnlaVLkenKF2+RlJ7iC5RV8s7DB7kcVFVdU43X3GFXSk4v0I4xu5TdRZYn+zKM8lwKtu
xDVdrs2EIY7c87T0G+f57pztPXLHlWKBfG+2gYYDDb0OjGGz24FD045EDo1xACx/sLUEt1YgJtZo
TGOYr89XFZItwS3/47BmIposxsgt8Q98aSo0vKlsDm2yxtoldgWvvkJmE11lqloF9nuGi/vlt75U
iaSGa5k4DcCt69d5gxUG9buE479IByim97C3UoCYd8a1Uwqi6W6UdwHGNeLIcHhiTno/zMeSPVZq
JXMMnFti0BA7VxnwRUCPhtD1iBtTbxfrT80oVVjzsVag1fqEKIw5XOyJbYrqSrM0HqrQHDBLACYY
nbC87ol5qrEMDSUOPEjUd3oZWZhs1z+/Day3unE18lRCgrb/L+hP2U4sW2TrcHHD6WPKETwW9625
1sXtno+00sVT/gG1+goR3DvEQSKeEgiCla0AIf1c88URFb2aatCXJqpwObWNxHIT7PTIiZqzDefg
XocuAEkFc5C2pyo/qSmvmp0ndFXH2ONH36tK7vIjVm9YL7FWNbqkfNhCrrUhCVSNn4wyRHnypnZu
VnOgrCKZjyTZFt6NpW5+TJFIAfHI5Y4ZNfpUt3GIqM6JtApqFKkUDle8pUUjYHEH3/q3xt+HdAA3
BAi8wJRGIGx9aBeiv6HvOC839Jb3H92BwPuPxUkPzu4E9IoSU+oC6LIIVQabGMsfeo1seQxsaKoq
1muuh6KV7VfYIFV+ZA2sE+N0IeNzOJp7jK326yIN2jUeXMe9jcdkYZ9Zx9TkB7ozKRcyAicVlmTR
MkYUjuMc/oBQcQKidUjRk1ORTb8NIoCgXerlR41P5W5kHRFqWgLz/icr+JKuBPWNmZNuDg4vAl56
v+cLJsNLaQdQ9IYQ4BSg2VxQoxPvo7yXcvEypieHEkrFvSuGVjho3UuNvtMOxtVeQxUN95YksyP7
JXy/fLmvVrgIcBjyAqmr1hRX71ImgsafisvGuYmgpofeP2iMnScNYxrcJUA6ZoqLoW+hnXC3IdhN
LF/wXfuHFSVuE4E+xEieBxrcTI8n/CYUkN9Yh9zUIZf34Op7Es+RnuoN9+e0PCW+mcIlGkXE5eRu
usHEZKoLm1aMW4Bi10V/uLf5hJfUnhNAfxwoRVh9xKCbCEKWgaTlxZ0PwIMGDX9Oq6tMwOz9gwpR
YYpx3lE5apDvsIpe5Qa1hwgJL39XJSzyNfj5KecS94q7M8EZ6R2IPXRzF3nXeto/QNZ7ILY7q68T
tQMFQXCmpejnTT/KvD+BPBQOfz3y/jD5OTURwuHmPuhAIBPRDTt5HxpRZnkAiZVyC0BSStrTX8kw
2Lkjw3H+24Nj2nRzJ/UZRh4OGax6l3ev9pTqCcecYPlucwTQdWM/Gl9FPWhwGwKcc+lvgN4ZGhHB
hYiAf8qjO24Zpu4FhKOezVO81B5QLO7iCtNclLY9q6NzdNfQ9yKNrDhuciKgrOLW9lF0UYMlgOwo
jz4gsW9IiFwTMaJkwI/UgnEae7VQGm8mG2kb7QdfaJwGbzxO/3hJZkbc7D1iE3TbNAneDzx+qhZk
wtSxZAm+ZwIS1odt/6ecpqhodQbBIoXjQFBVx8tPwUogxLvrlM2noHWbq96nR3u8363Z3rSIzmuh
7DEE1zLcI8y84eli43eQlBLotgdsXIuz+KtQj4Huq3fSSxIwRgFjhJvHQ1NmZ8kkgn7oLe2PE67c
hh/W9bl8P+82BKmcJGpm4n3ATuC335n1uZMAOmgQr+lEbWzIc0afNPSmJoUrnEGIVtZmqqOEUzew
Wa8s7VAKDSP/+FYp4bQikS31cgRcBe1vsq/o4lRLvAsc7JiwM/nL6bv4g3X3DIH3CKueVpdFGJ+I
/zdSmCjLKDonUURz29A2k23k8NscH1aY00WLWy1gedDqVbTwlojH080gZXCa7jQX9CIBiIsXIxjM
+9+pnNuA/E8Cl1s5T7S0Ck+fAD5NE4LeNEtGCWaF5ZoyUAvwj0gJnGzZeEC2PieuolMAPgjq5DiF
3onotHBgKRYjY9W8t1R2BBzwWUVl3kTtFZHMKLhgp2Edm+tiUKCO78aAJHnJreC2mF9JQb5WBDli
u5zHGCakxtzDOJlezVhKcb2//pijLLlItiiAzrTj4Ootj2xdRh75h8lshYw2m7M2GiNZvX5kKNQ7
qCG3vFCxNeNKbrmALbe+wF+I/IB5jZa2kWmGxdDyKVt0HsNdPnnVA3y74j5osU+NTuDKzJrtYS03
Q8XPjgcrIxXe0HMpApPXHkKi0OWsyL34XqFn90cGYyDaY7EtITwVwefitvlPFSEd2uFMiKAc0/SM
V6O7iDZyKTb9d7Jdc1gSH0OiV8OA6lK3O5uPrAIQDnMrJmji1cDhtDhcQZISz+QZE1F1okgSKMMH
DKYt2XhOyglcpsLzKr/gZ9b9kKgi/nmq91DgutOKeu9xbec+0ouZwB15ELBu9DVwAaG8LphWWuHQ
lLkiePzp9VI3/Ucky2llDRpJNralXa2DqJGacksVa4Ab0KQ0UDFJKdo2xRUfvRf7CbDI7RFbj1qU
0WyDZ8cfjeqU6YEbDu4EgL+OYAT6qQ4cYwAqtCTqPFBNbHWAwo5cAGTaChERcJYnsQEaDHy3mbuu
p4rVtraoOcM9QVXAi8vYVUb3HUnJ2/RIgX0YC/sfjf8cyy6Q/weXcEkBeFvnZ7Hw6Ud7R4BdMvXV
IKBStoPwplGkIeuo1X2m27OFfzX+GrLVFxAE4Eqedf6oPE8YT8unmoUekXOgxeLnQv19yWicMOEi
z0AUjgn02NiaPXPpTSqItAzX06CAP4ScNnSdhHrJpleQv0ARUWyvqiGUse+Y999/O07o9VB5HMpQ
ecPdpxfVA+wlH+7Nu9GEiVjHXRNUHD3eRf37DVMPFK+8b/9u7bz7vtgWa095lWWNf/rJhMvKd55s
bbzwYbLJGQbuzSajN8OYsifbj7FuSNChtqJQJkseBAxf8lcx6YmoiUabGQKzZ7ayXOIzFMj6HGuF
FmeKCQnZm2Z/KKTowVhJ0uqz67W0Sy1Z2rxAiGt/LekuXDY/ionBFX4L8d1hydXCsIjJuHZwlY6u
C7kAVFT3AqY3OzOYpcLD0Z5UAFQI+Wi81k17uTME4Ufzxjo3QxqpvLQRcw+SjK44Bq71/7794q1y
rshNRXDLvPYYTtoV8eKSM9bRcBVySaeLfSLTOva0igW6Q5tqRj+NBAVt84s2KLFlwZsTKexZ+wE6
7C92+peGNiK7kn64nYh/rFZUUfz1j0MdbO+PyPY2j2gZNtUWdyZbznqV23EP9DuXhA3+HI5iylRk
Cf1a0y1joGmj53sh+gxhjnhA+XELM+GAQxUjkHbBFCafj3lnBmQUFYbWKBM0xWuOlUO0jbRjdzaU
tKGSnJ77RiG3iLDZLJH7h0dCkyo8Rt8+eXy0VXNQ6mFlpNxaM47KjD0UuHbpECOqMRh17ezWWmkF
UzXbywI+L0R0Gz9L8eL7EqtQblkQYc/BJ5vJWje9ScSJg4OM2AmlMb5KStr0SrUc02uaErBZn/JN
T4wsoJRi3OwRi0ur9Ngy393lcpl35tQ3mvRJqJ5Gc6SzCoWkLGvgm5IDp/fNBKjktxtHaKDWr1Ae
xWxoLbXEnCt1vi/GVbNpDWsPj6HLwmPooanza/lpti/cAh6cUjePhDS8UA5H/lufnkYXZIlFleNC
8MW9Lbg/QdDVlpxrE/z6sSSHpTrijbv/Wq0+bGzqdqFbFMudLVpodbQzhKQwOYlaKYCqBAqUnx5E
NFnxDSWnt+26HJr52gxw53bDPuolLhE/hk/qVKI5tlFJdPzmmlKa/GzxXWeSesfbLBQ4djMKigDf
ypT+53c91FjLba0T8z3Utq4DdzuxiCx7dVApF8CdaPscZ/LIQzVdEs3i27fvyHof+yjvH2MQJzzR
ydvdPWdwgn5l9AwVnQ/ANyzigHIFuZXsbQgmbQNWUkx4UhyURpMl8qlJSMLjXnKdV/iEXuUcj4ti
DWmdF+IBZnPvdqDh8c0uP71Q4/Au3iMzLgH5IDqhVjtwMAg2cEmFgAFFHjkokuutrCKIZYISm2PP
flWJ/8znXmceLz90/463EFmIsFuWZeu+lLYiRK2A5cPCwOBN9bjazqd+609HRslHUDWUTEV9Bi0X
hLt0damOAaXmDJau0qhDap1GtBRHxxLvJy7dXKIQa++uwy3YtuaF4vvXjZGKM0EqIHkJeWVVNUrY
yH0zEuJMpVLe1NOIGVVzn2RM4i79/NmdT4oYpQjlCupoOhJWbNKowcoxZbs8XzCeIqgk5jkm1wzG
Fcnwla9UwnxZMKSirGsvJAsoBKGFrwapuKekY3zvwt/5QoGDrrsvahEa8BXErRBG0JT/Jk4NUSQs
IViMGQmgL910IVSwzAbXNYX1D4jM1QVf/LG7/ff/G6VpUDwokmWULzKBxuh1QM6RQVmMRSPFX5Um
I3DZbJNuymlMt0j2OQozWyR+HaYcbWUipfK4I3+mt6kpc9za0pvsBcT7NiDu36lEX+4N1RhEMaAF
YQgQHjO9mpWIJWFLwqV6+CPHbFXXccEF9PL8/1jN7oIjcc6clIhy8reTJ/tYTB39ZqjV7oGjJ3FN
QSNRYvGIkIQzL7sjKiMxYL+ADnv/cuAA/bxCLOOtFSshciCgeX607x5qyY12BxQvHFeFvp4KVNW1
5eoBJSPvHan8mZeGJ/vktMf8IE4WnOF6ciKODtA8KJINJUC6bWj44O63dcHdzeHnYTU2MGNIx/K5
W1pxXOeNHNfnhMg1soNi1WPe9/yYByKsxFwJQNAdUkyxFD2sRgN2Rf8x10rF0ZKKd9CULyK0OgX3
yl8yNLZXtWuy7GguNZ6699Fv+p4IjcLTdx9KJOlB2ON9vnWyM1Yt6e8CpFKd8b8fgvhCVTIexdhu
6q33eN3zl5vcQBw1uWZLZ/q1fGVHQ5oK9l/B5M7301U7/f1YQyeeCV4hTyBuFMGhkDnYMiVeL/9y
oXACuu59DfqsAz5hPbbx5dYEybt1NKOIjbq65Sz6niU0ZUfUxw09w6bf/uLn/cSyTUodu+HcDTAP
o1NQPRf3n4Ate/oBoNo3AmJ/IkpVvgyM4TIHS3ikZwP7ZYPzR06aI+Kuh+RK69YO/yanxTWF2ZJt
t6SQ9CUQjJYjFlGWU3EPcUk3VVFn9al85ETnxLPgmpcDSobolsLnamIRnX+zCjCdyM8edxJThGd9
j2/oWLfXhs2eBzViS8wxlyJ8BsmPlP14BwKaRYemMXnGn4vAW+Mry6QyThRsHZ8JgGlBUuIrTvo5
fF2lOk/xkKBPiStYaLEIv/Gf1gAOH78Y5EVPn30iXHWSx1cWXEbkZVePx5KVyBz0t7InloG4L1Vd
LycegntVsmlVS4SjpcDfwBTEZYJs74/A8ScwjRldiHiSw7qXnQBRDc8HlQGzKpzoaALiI46F1eAf
Cj+yDlQf5dtApEO6OcshM6PGzC2S2wm3GJezr1ha5rMgYMDRZqASEsVA5SvTHRZTeswBf5PaLxbP
1F/+7rHWYAEdmnzrUmWfgNjO4HVnJNjMfw3ZSEypo/ev/IQUQuEmNo+ZgkoeZ7YdS2pOuHKOJ7yx
c9QikdwYW4FPTeO0OYPl1iKeG4v9e93TImr8NaPGGrOdXpsCx7U0qCO1uo6c807xvCniSr5z4qKj
0XSl8nuQSbPVQmRh+gyqe97kXLezRa8mr5NBqxYhJnSgcgP/GimzelqZm/DnKLhLmd6Rjp6DPOaY
NOa20idmybnAAUDS9/Lr5Z9R9hIMimDKFqpbt5hwYUA0bHj9VHg2izdTfZCRu3oK00iFrApEXoSD
38RjMQOoaeCkUNv3vKzSH9zDv2YddwosoYQiilER61+3wbAlVCqF6VsWPblq+I/HHUM+UmdmFa8R
3kv7LypkgnDu6JYRYj4H+0yOkz5houJxSJ1orgesq8y2F7g136YvM6O9Rn1mnAZqIo2a7rSV9eBU
Ycu7hsylFJDDjSFwnE6zyCUD6Y7MM6kUCtbQ1iKMjPDt4EN5ncOZ203d/4RzH0pt/Yg5DZ0rPurq
7ejUq7xAMnpjxkSzGUuo96UZLBXivlEDloZAMOJD3eHOJRIHLasX0+Z+qSpLctRbq81TwXEds4P7
uVSA+ugF6qz+OLEUtbbN8cKqyG57Xa80cWKHSDaYi2sAhU0gE3y6W+oNU9qMJhRSBKvBYxML5VMu
vkMBuv+cjonSLSRSls8tMApg3LTP/M8nqRWREz8dIB3Px8V1RYEdDQZ9YNg1rZD3F8EJz3z1SZZB
kMR+F4faYsXtSINjqRDJJqTWMb7+dsCPJL1wfEadgztxWrHmKZOwtrcfXmSz3kdVxoXRWJbY3maA
TuZG+TS0nDSuqT75yfkZiufd0wN0aFDB1TtMlBJbLD/qNy2rIz7T+gbkqRJB5SlGZh0HmZJe8DGp
ZgIMW0Z9cU041Owms6SUO8YyGKcHsffRtisNvnM1/MigBdaRR6Kk6n6FyaO5lltQoJHm20JLoo0/
kMsAh6VZgSYd3bg1KKk5fvfIBj0jnDjERQxWPQSWt2d9mpRjW3Mo0QMNVK8W2QG709s2RlcHmGG+
KvB92yke2VhiFLXfkWdGhWIsY1I1yaHGkPNIdwexflJl0RBHdv/S5Zw5/REFHuWed/xfLihKuoq0
z/ZNjQZYKrsvBYAzPU4QuUwF/HB34oGt0swo/Z+bTizgxqjz1rp94sOJXB9MaLw7baapwBSS70AV
KA40PTch0/abUpJX31JCgaGjy7fW+R55jVFMaKs4qb0WclsB0wcBCYp7jUPxkxhl6y3a4aZ2UydC
naaDYdv/0lcO5aRQ6vZERNw7D3FbmTjvEZWICtk8SSEdbU625RCaVPJiPpsI8Ddf5ZEN9GfO2eav
ZnLElFS8F3WLdPIyFK1G4MgHj+wiKRmTGO0fBXobnnIKkXZD0V4Y9W5kBsfd6XVSKqt35sYPIPRQ
KuiOASZSMF41bRtSX7hhkwZ+WX/UemSW+z6WVULth462dPlEPlQ9ojLqHyY6KKbyxSZ/OAYV+SGa
rmZfLRV9n3lvTs4S1GRQme5xLeYTg6o+E+tmFE6IlCZPJHHaZped0Q2qIAYC3kMggN/EpvPRDXcE
thySfO2e1nwDax54VFqfd2pPGXfXZsjZ3kFv8z8897eNNfTLSfMtyUs3bNEXP82Eua8UarI6lxW2
ChB+0uSM4RunR1aCROo8BKMxM81uAQ/O0y5vqupzeycK56WOWk9xgT48FvF1DfS+F0rl5vJZJ1Gb
bcz5hcZkNZ9NIw4+1lzhvmlatwbe1e69yq2jcw0qkI0028Hrpy7cOqEJpLLF0TKbf6D9i5JM7Fkq
ixEjK+RvSoVlJVzlTpg0FXk2HMJZzEOpyOmBBqSeGaha8tfXEa4o/SJzzZtgrZ1VIBcrHMY4Jrh6
J979o1o1mIp2H9x4M4GJ0lvgnv4pFG7GSVE5RkZ9D68fzMUoiZy8y5c7WQXqEOMVqTXy/cZO0xXz
d3ThYCB9bjLue0O9Hx+INGZ75Nt1Krh8wewPy3dBVZ8pUiR3GgWz/o6eDxMcuyVhH1UHyPxXFOuo
gOSxMHdvgBTc/esTgOpJz+yHwFTUXeMGd5SgRSRxHnloc4X28NbMl5JIXwwLFh4muvWm6fFeSZ0b
CHDRHcZ140kmury1KjKwHo2ogmBpJD6fTmMR9MEsxdK6wN64FL6YBTljXniEKAafzP+81q9aMgZd
dbmADY46C+wISqD9siJIWtndclMVmIDSK9YCJB2fSxoVCvG/MeBzFH+c68JYnw2KRgOY8mJsh9Zr
X/pyFXRqLinOk4C+XW0wI9G8Pd9UFleKw6JYYvRFivC+cWCWLBHmfaux2WH5PiDSJSVDil7j5iTK
noiuKXdZNlDHFbYJc8jkXEnubIT8wNhh8JTnZO5OxYJw0B1Lh5DP8Q8y/1UpMVpfEACJQK9IOtj1
Iae3blN5WAdh9Dtlubt2HdqDXwK7GoVFlSzwtKuV0721Z7Q4lsp+/8ZkCBw9RUDJMw7DRwE9n+7W
wHFI7oIjnIxGo/0c0pWDEoX2GiQGWmv5akRa/fzPySx5QbzqVqkmE45BxdD835XK0G2lZiuBD6eQ
9o7retTveAJWU10lTUX7+XfpybVXgXjgbu+3rFD9R8Q2X5W0HlSUg1bLe7+y2aQLfQTijZjO/JBR
qrZAZ1h9oFS/2EBPyNrT3V7MwMVD9s8nIFY/F4AjrPBAwaO7q947Erx4Tt1hfPchsMGPvXbl9Ek3
ACaU4So6IWufM6OZp67kRchL5x6ZAZwVjG0NDhkH+riDTic1BLJf+y1Wfsd5c2trAx15aM+vNBBG
KI1jnbyqmsuNvE6rLSoNgNo9iWSTHMzswrYq712e3fWQPdLAzfE5IpPQX8pD7EaM19EYuXYxEU5X
pM0VSAOrnDrxcpHjSgSJAaIlS08Ty8WO63UEmLmjN7iTkoFWHI8E3h07K9q92scpfY3wfd3jzeof
GoDM24BLM4VF5xec9Kj0mp2aBdDT7sa+vdYVj31WmIUZRnJ3z8bmgceK2J0yykXmdTKrU5+lBrP+
NywFXshqtpwzlVxcMtXZMDEcDd1BpRix5ZBi8fLtusHkVee4cSL4m0lx8D7wVlowhz40tfTQHL9t
qAoxhNZZTzQA8MMYradPe+1G+UymtTzKqu+SyIKTgVZhGejsw/BoiK0dXeD8O80+2R9BhQwIAflO
Pu/6lN5lsyeR9HRiA1vng8ahaFT08wWYoiDvFZCgjrQvlQzIL5B1Yb9Lq/TrQz5WVXGS+Wmb7fWb
ny+TRy8fudmcUgCUjfjsivDXEjH99HwnKb3um2u8U/IBNlDJc9KHaGgkC/E+BEpytijeeyziHC97
3FjtRVp2PhEQyh1jVwiiYRZpNdRAYvaUFVw8lYLlvSDy7Wm9AFdgUObte5xONDp2laC2wO/5y0rh
DZKqutjuj7pCkjz+wLUkT4C79v4DhL39QuI/nZV2jJEvBBtZkNkxotUqKj61K+963zoxUBduRMF8
bDIt2zBJdAnjVTvaXf8RfrBhJXDeKFmF97JVLnFwoNH1dpEADeGGlkntyIQvZOsXs8VFBFJCTfnv
bl/6dy835YJDoJyyglQzxjJxPAWX5eVtQYRyY+T6Qu3hV2eFHxeSJyC8urPa3Qz3FVxzv3/qLSc9
SNA4Cm3wWMvq+o+iE8RJv/Yr5AZJ58DcFLS/mpIQXKCrD9Uh+xVYSjgxya4euTQQ8mlNaSC9O8cY
GVNYV829aoRLxEg0SUd64Ed3ZLmqDAebpRVxVMXoyfKpFuLSXB1i9gkde1R9ElaZqmfyrYcuSDBp
rP/WGQVVf88u+eh/EVLpEVpT6vxkju7QtSkn04JqIbo0VBLsYKlW2EREAPP54tL4Mo5odTtbcQBt
Dh7fY7qbrbZgMqnG2Ru/8fVptinCsasR5kdEBQQ1A8C7+uJDPhyIBWwFch8URFmL84g1lrWqO+68
2Y0/W3oHE6meLfdG9Ycnmy6TO8RsZTExbHHn+qd+CeBK2ElOcESftG7ozdnLaom+vRy5XYvuBzY1
rDBgrhHcjYYETD68rnpT630xAv5UBSEcRhU6QAiVIBV/jdevret4uACJ5NnYqDLZI+peFIetC3dA
AY1pNp+SSvDnHam9xfDfYuXxGoYyacxuqSuvkIFUBqCLeUoCDp9XU9mFttdV0UYEO6+N8RmFhaY5
8CW6VmL74QmO5HqBwkyhYFHmvfqC1BLvs3/HqEr9CcB/SG5aX4V8SthL+dpMRGSgyZed6+RONv3T
/EmUA5Q0BERTG4AUCTJ3CR7nuv8BQGmLgSyBPERks88qm+YH9vFO51BNvisd7OashCaPJRJ9EMf+
Y6hJo1bth61xopp728uAKwZGVMRLPZq2Ir10AwuWNOMaOYaCD15ppCz3gNLfNkJY8lP0r//Zc6qy
v0XNfEW+07GY9pDNnd9i21F1lbpisJhqiK4zAnOztfwBROuPT643+b1n67QDTAZng4uLxBLM7TF8
eG5Wk2Ahmds7TqME4//1weEUHliAL6kthDFX2rRpZcdtIFr3bIFBW/7FGZ7hLJUnlru4tvMK2uZZ
qADzHWOiokQca8RkHrywKx+7NxlgYMNJq8qg3SdrL4WnAJ/w+UHBuHQgdnxWkDKQsM9U8Qc29/vg
vW3yvj7R3fVJfCil2giB55TRDI1YA9MKKr1KBDLYLnZ3vMJ3RbaUlVYxU+snRIX8WeZFP73Aubau
yJs9bpufMzx3DfSlCIbUzwYQv+U1IR43Ns1SMrobQUBueJgYJx32yp4/ynvba0vkBVdNFRX1Jhyb
OefFTtsMv3kT4HPO0hk3Q9asQMRSDtWi22+ZOPIOmppxBIHiHoIzRhI5juUixvToMZ6l/CLtqIdC
Wnq87wl8E3am9cbboWLbAcL0c8ZBYLdeT9qEVH0NGjTZDvJBiXeiFCAWuXebp3fXGlZXTbO7rszQ
56VTHSz06zomeC3tIGkbwO+j0si03smRuif8rVlL4Pxk0Jz2U+6I+ZuTyHKZZrUaPuvRNdMMJ5fN
Xgowm7EElPgW4sGhzntfEDAvg/VaQlMtdZ4fkTsB3VPD9d/8u2g3hICqbLVwsInhZZqFdiLA5Mxg
eVZ10bYEv/pg8GTP91LiFHOiM2FuGfcNAO0+AsvYmkpEAYcbjl87B075OtgH8tjEHF++ReXzKVDE
raX6bFmeCOYdm8SY03Rnh2zAwxKlAH4V3YHUcN+4FzRw3IRXTuhy4yh8raQkZSgMbWdlYd7zuOyf
mDdMRB67YAYpnjUqHu3zc0MdzQuww3zT2JuzalafEhA+qOKaA7Loq8soW4HOlIb3QiOW+UHFADij
wZKB7GK6jqOc2qIjH/MDVwUoeQxCv1ulpzW9gJsskzdi+0Mo9PiYp7qfCJ7vf18+9lwf7ZhxZGyf
+Gq7xbv7zQc9Ez8vZhBB/okAb+3FUWpY3DbxMeit6O7uEvpHzn7XGsLAf+SMzaJyPhISR5Webb7x
QEy4D38d7xpFptrvq3SkuV365zjkGh0VRd5ZJ56zm3jCC37QHa8GLz4+ZEzWAvfuCD7Giso3a7jU
s/uCVQwGDbEegsBn992MqWKwp3FMPl7JB3V2TFaQt3LeHjGQPS1mg0UE97cXhP/vJPmV+hhb0nyw
qkzlfZ2e2+6ghvxFOIJd4XELSKawYemqsA555Ze8mxCJndmieCwrVyhhJh/qkZMLoWaRQMxGbNkF
/De+jDCmWCZAwPVmnABQd9R4t81I8Jj4T2bSEijbJakL/2fryQyU8WJsYpQVef2eTHhEiTMawMkw
dSrXW6N/cA/Vf+XQE9LU+yA0zvSX+5wydg8IAm2ReUbFmkmGEo+FuQSx2iRmOv0TRBlpZyeXXPIK
E70V+P0F4oYZ9uozrX3jvGVT9C5lTmQtigrdXuxYsEx2xsyEm6kzGVsAonosn3yfvu65pVI5Oov5
FQPx7gdNwlYr8uZXUY4sSH3uFqdK+O1UBgqc/SMcmpD7QI9x54a2/+5+j2J56CsxmdqUvk8ioTyV
ISYH+1EA6ZIQmUxhAE1a+dvpj7OTlOKwPjOm37W2yIijfUnDHzmq3KXjxoG/nGizB10JpKHpRNyG
JgRW5KbuiHTcke8F7HA9MXXKBeUf/+S73ArpS0+Lvc0PDKgwitrHkmKTgeacQ+eNcZlxcPyn/dom
t2MYGDfqYeqHs/QhzARzhli3BQIPlcOv93zuy18Rlb0G3+YKHjz+1HTZUrCcUQpIh/7aXgb7NI4h
9Z8bNevHK3S7h4o5mu7nKoug4vHgBkauZG9I+Zs2ZAwHv17Nxlf47LKjPmK2NF/YYwf+BSHevwpx
K282vFxNYeqlRKzR5Sb7fQnNiP5r+NVddryPWU5g5uM8tNspHZl+2CONmUX0yo6bhpAAAYPKSBHW
topxnnB1tz20d/tYAR3lmKWHiIEXyQbf+K3kpLDRzgQ9pfW7mrzeAncMZMHXPnH0rq69OKzl7Tly
MQS8Ug0+IWx49e9WTybbcBE2oFLPZKWErkk8Mp0iN/9DyG/Sf9s8s8f1gOxH3MYGxxXnVcHVG8Ed
wuv1ZH6LV85IzoZjA1GYbVY6hF+SalPkbCQrD4UGgnUeQ8smNYgKf5gUm67+Y/y9wzO7El0SAZKZ
77j5KP8LwAwqJvuxezCq/bzIdJPWUkN8nX3gZHwk8kZAqYTOQ4YtTUC3m5ETB+rpoAoa0CLj1smY
BKA9YzbFlNklsTaHqgbKFaqreIp5pkDU+vPUfwIaYn/a6VS+uTdzgOVDTynMKAbtHV0ulc3L1GWZ
GwyxX8soHBWgDOqcl9vlALqott7Ep5/m87lHZHgEER0UL0hRZhA3JsDudB/WxH22xV3Zhi/xNFAi
l5eBaKxRwgM6q7NWzcOheE0qqCr+ugcu8MkD/DEcnqldJib4H+OLn6mOxYJupp5q+ZCpizA0pXl4
RoPY6jvaiZ1/V8q7A46+yBGvf1gz4gv4wJ+323wKtj/17JOTxWy0yRPVuRlk/x3k4P6jFbCgq7Ia
pgxYy8fTI3TS9ZLr9SvWUAlnrZykM0x3Eqc6xVy5WZl0EsiyOCuhMvKqzEeCLQZDZdwlrBJ1pFe+
K+CBAkVrdqkgfCq4t05Zhgs1Ep75/I43JSE+ofBOQKlQEGTq0cio2N2l7PvHIqYFbPZWIZGgpDE7
mpa0/tBB/2lqYykRZv3G/E20I3OiOBMsyY4lq1ZrYSG+B6XaI6HNiFp8GSHTGUMnOuwPFteVfslk
k0vaGLNTAP2KqhczMdj5oxu6mN1DrR8pjBV545mcTN3biwBshiHaAzlcqJwxSl1m7iStTzMwz3OQ
ChLZeRtmwi/p4SuuyZBYlZE/AkY86sh/jOhsxvPQHh3aUZnz5UUx1D9LyAYzQnDBImhjNvAmyM4X
H0mT50QTxG9MAzTZXO5Dd/AB5gnzzepMympOXJJ2M6he3pPQ+6doviuWL81ldF1f6ueVJO/oUJrQ
zO2chjlVuKNEihz4A8cV8N2UANN4TiCIS5+HmDZEmfhvUUzuhLomRswiDPHt5+hSKPZMKoQ570Km
tDh7cyjC3hmgeWLFW8TmvpWAw5wtbWkRyrZzETjsohWCiUWjqUJ8nFhOx4kvXL7qunRv0WkRWdwA
RXcTb1F7ZF6GjTtAt6frQhLSPUrhT6koBoVyHLCbB/YnsPccGUcQ1ziOlxBD/RDk6THBDCNY9L9o
epTKqJ8kp3q0b7kKjAWt2FAvqY3Uc4idr7wZlMMeZNwXC3sVUrMTnlzFJ5JsoHO7zX86P9FrXUap
1PTFGLRLlINFha0RPW2UW+oIZWDcN88IPVmBeooinXYZMoFfD8J9fRxzLpIAlOKPiJyZ9OEoZDAq
JJT5kT+JNuUOimfaIGjCOq/GgyU22vijKmj3AN4wQavrMiEKAo0mg8/DyCmsyWJAEmNWNSfS9r/7
IXQDVsy7/WnwOWfhP8X/TTQ5UxaoZk+WpqcIrFCfCBOpVJmTLrQa9dVrPANKTrmvoCfaPE3w20ox
8ENTkkDNl6DH0JDmZYWc0ON6hhTinoX8pQay7nuQrAZztT/YbbmQr7Lj5M2kuey4KR/ZlwUszILS
mO13UZEHJjtXsOVp0lsRpuca5eaE3bYHJAhg8ckljMGc/835b7pMQhKeXLNxOhg0AeJAp0HQ5USj
XRgAfpzfWua53Dlud+KZr7mtA6PdK8v9GZdky6VMiV+4BnVuh44FNSBxUtM3k2aRL82ulzMmTAOe
k1sq0ylSiEAgwQrB/6gAoRadPqAdbGR6Y7QomPkBGuQpyYgEEBEe0x7eBQJzZz+/MtQyICuGry2i
Fe63F4RfFuXdqvP0GQMQ6GyCwQc6Gz1i4TS5n+C9BmugFJapRqwih2Y3BmFpFXe9PgNcHY8QmecU
VFbdAYnyIh2xqSSUOwqvZVbBCXCETSyRTl7eZa/QR6fBfFGVvKQRFFkZfR64MnVdp+kgIs5wDju/
rfIHlUN2KgdwXVWtHi5FHahz/lT/gxfYUpFVcdHTgJvaZ1vDYG1jNsZZptSzoXo92m8zg/2cpEWR
+CTVMON4niaHYg5XdSX/Bi4KujElyXPmQPcsANoeuzAdLoeBPK1UHz4Eg+RL/9mEJJGos1JoNjtY
QhBev9Cwax1E5BjdN86/+AErrNHj8dW8AAEvVEj/QZgwnRzd1/rHr8kpzCMu3DKTUqJ7+vAt9EaQ
/j7ktP9GjaLy1pihZgLzCyVURMxUdSJdMU3Amls9LOjaWQYWtcQjXqTXZGDEbFx/eCo6o0U/ULrE
qFydTa6cYvzh7vABoy+J3exsju39n3i+ipwfzFLl4jYF4bWGUqxq/ue1N4VF5VW01CYGoy+ion3H
nA4xg+YnZ6nUVGF4u4pkELCaCz82gQaxoZM0Tnfowq2aBqhR56471yrs1kY/7bI8RsoPQsE1r/MJ
ADTL/QwUgDihLIhglfLlLkSu6g8MlYCzmKYwmRyK7SmcX9MOXs13ktV+Rx0bpz9mR0AWhAC8YmDS
2xhRTCuETGo8EuopNSG9ePYtH8DhzKahEdS1LolGPFw6yI4O17+6PBgsnl//W3DSvic2isfmX7rL
WFa37ifXTOViAdnseN2UveUrdn6Le6OaVW9MVJx7JKKGvxu0T32V4gLGRDVEuXqpRLOZabsKEEKv
V5jRepWPPIV1zYfhbX0HTW8KExn0IJLKCgTPa3eMNJ+kZ+3GG+H4RNzq1IY35djPClK7MCdaoya8
LtHlh03MI2E9JMlpOHN4lmTy++zEox0Acj/leq2KdZ41Y2Op96/Rsak8Trbdw4ubsqxHlNpNIAcG
swJLZ75XQxVEKuLSLkNOrqFpO2WrqkkPSZcRimqNFioyt5nkl6hs+O5Od11gRLThbVJXaZx0wsdz
tOIYAAvJxNAGs0y4fYjlPdYmf1FA7r/RgxbkbbLOfM8ucjvZiXjBJumiUE3+VD8+NU+y6wtd0gpr
OxnKFkGTDKt/eMxxDhjH2wnmzplD5kNAKcvWWsdnBu3Fu2GP14aPLma/nOs4LBpzYz32Ykyx7x//
NzyNds3Jcv5e6wjsRW9ISP7CGsI7xXnyKNYbSMgPZLMVA4AwI5W99ZLtnURWDtc479lr+ACdEauz
crexJZ/O2CsJM9rU8FQ90Ht1mptfy+MJYIAMRyzSwJW0QY3EzBR1jjn+Avp9N6P76bGhvJDb+aJu
OD7GId5WyYfqb8UDsYph2KsNYtsBEOYxmkaRN3EehshabrOeXr8DE0fcApAntDYUpMbNpfDa6dgX
bxMxbPX1fBNHcPrpgp8d5RplEK4qwYXh38jB7Y/C6eswa1yYVCJSbSuTGfc82At8TQr2+iYynBFe
PXbGQYX3h+5zOr6QMkzRoHkagfRAI3JMO/UCFyfo4XNbmMYYB8M/l813t+hXU7lVpjHtGPd1ewsH
1ohdrwYxB7gtK4aScuDy3CiJ8b3zq/v82i/ZM+HwtLtnJguAPIfGzpJ/Zd1Nw/0g8XEfUyWWFXyd
heoce87KZRRDQTKSDuj8//TQyClILXpc/w8SvAdMhYLADhGs0kuxi28vLaOSySeXSxu6N2RdRAdj
NdzlhfLpavmaEsdSU/u3YNraF50x4B8bA3eLozzJwQ0Z+ZpEb7XGJy2eFXxLIvAf23fSSiu1yMcv
SE4nV+qPPqbvY+GLGRSZRAxRysoR3z6gkL3IYMpZQID4T+pWiEZmbAD6bDODxJ8x+Y05cii/YMKZ
E5yWHIe1Whk94zkHnBqShPlVBE/bzau1QRYOQZAyKDu1CfhZW/MQdwXqK0YRysJ20XsasrNPQ7pW
ilok0Px0PK5zKuGkZZccKBy1O3BVGqZRbHIV0MGobsVvec1j7A5HBJsJXVQ6HwYQf+R4jsO/K2Qo
uDc5Rq6QOyRi+bE5KyuGCUr6qmx966morDxlPgUtxXRJ9WWSjGc3xv12CR3McByXfk3L2FZSuapE
QJrCP5OoMe4wobbsPWleLmV1PU5WokscWXOIIBGTkt2d6fNiCQim48wv+UHacsn3/Hy5yE2fCKqn
y32X/6StD9sDyJXtyPjb6x0EmScnsgB8aUNHH0imniBQrE8E6VVVckR5HPbF8AZxP7sZWuL+P338
gKv9E7zJW8CM26ryygAhkrSAc6KuIiFT4rNDv6SJT9Z+ohdcXBgfGDdcRQVY+UKsljtOFrL2/KJi
JZmtbOVySMxMQKcfXZbOHobWM5ZbgaUqm0BfK2SrQfZgkCssEmaGbvihVJsHGD2i9tGVBA1NBT22
ieJFZyh7d7ME6SgyPs5oeTBZCcYzMQ4910CyKo5b9DfY+FtuYfMUxXkxzgua0HExFGwFqfuffmM3
ILI10PSZtc4AebhTf2pweiuK65zkXfgYmN/T2lQ6zqslbf+egG7WslcleSfecpuIgEzZXjZ5xNrW
pKOjikA6tzQNnL+Ar9ssQVvP4ziWwrcoyAVxUgN9zadC/LFOmRDvtSmISB0aSDwNewVKMUT6X+rE
I4y6QteFYflBVx4sNTIC4ji5Mg6aD4dwbUZbpUHz5Ad16B9a2kpIpSjobHElCPIWzGcuJVtDbDOG
6ldPRPRmiHjyktjvGDV/jD86ZJHzX9PgaRhIva+amUqNHuLPb6JTOWPZNht3r8EttOgTAFSqpJae
BKD5JRGrB8f1T2qA3a0G9R0hUvIWaylEPcsGmY64ZCj6dHX2Vx3FUUyvWhIaz15zyFhk4UAr8zSv
o8qh3Szw7zMEnuMWKP+26iK0EeGM0+FU0xb79r4fVwRIsJM97Pqf5xiysrMrli6Bj7ZJGcmWisFQ
d65Nzvv3bQGXs77Z3fxodUr63/iMX42BSlztv8aW+t69F0qTgvps/kurSFSeHYUnB1DkvcEF+SNw
dXIAu32gKOfxjyzfxfnFvdcXx8pWU2YxI7Bd7gBvWol0vhZOwtQLMoG57MRT0PJCMYXT3eaONQDP
hxU0/gxaMgyD+TqfxNB6YfwyA04PzGbFxs+DZBzl7oqSm2Hgc9x7Wz14FM8NyvBFuluvMPESXXd/
rYR++mfr8oCGZw2VhqiW7GQF0wDcmx3Wj44Ox5Bh8+Fo5ud2SivooHGuRBImw7+HKTS4Iiw+jCqi
kVyiJRoH/a87Q8/Un42pP2lyiFbla0s1j6wYzPCZDj7yJhC8zaqD/ym0sd8hbKWXNtk1dqSbt4ms
7YLr7QIjo+JFCqP6Xosx857doSFDSdMtqLiAQLmjDOB1ymuspNwLN+S3Amf/7QA7PQ0UzoFtf2L9
lCEl9fnRxHkgyZ7AuyerOqcs6qzbIz6tNbl/I8BBr3uAeqieNVLIT/8TxqRpcSdMYhh3ZKPH7DEJ
asfMbJVPhv1qeHg6Wf0OiUv+ae7udLyRNtNMXge87aGEWkIXpI9dL3cOF9tf8zwTPKM7Pze7Jawt
elhZ7cLSULKg63/2QvOtZydQGdHM8LPsipbC3nbhCSAFFv11W7DrpbN+kEX0QBLv0T4XSdcAAQ5f
748Py4VYxP4SDuyni3iNDnKScFPyJyxUZh7Kd5cZQgepLVWo36itn3fIGIpf0mkxCvlK2vEezzng
V+5Kae3kiRV6//8S6JcZUQ78hSzzqmz4BZg1aalasDM4tVlI5k9W91c67dHBZiacCR41NPafSioH
2PPD1PN6Mp2DwXqFIEfBo9GkIcuLHP7jjWEJEnslo3AVar+U3vnkXwp/B8bQgeLqP3R4WPBXQKtq
uDNlpi9guNluKWiBxhHS620ZpH3u7DhS9F5xQkKWxuU2Zn/yGRg+1yrYSlmIh+kgVbjHdn/WzESQ
u6LAVcwxXUBaEObFajW4mhW/xqLiB+bE1jrzFb+kITXu/ESTw3mYNI+jShsx6wI7c+6/WtX3kz4D
jocZEA7zR33R73Z2E4b63TqveLQm3uBkpgDEoM/IK9cW+xvsKplNeOvcQTeFKtdOyiSCOdalii1h
/R+FeAVYK1C0jBelrjsmfacfihwjjdkyNmEJYAzJfze25Egcf2mDiZJya5BC3wPj/q+cVPw+6oT7
ImUeOONqHgDW8rtMP0Zy/QTRCOa/RA+y/jr61ff2u45B7JhZkaEYrY4z3cLNATjpqLzNLLQLkVzg
eU1XfQJL9KXr1aRF+pP0cO4B11O0D7+3UvH6DDWYKscy9A3Z9RJNSQwxANjWD4QneZDzEwRa8UKY
2N4N3WqJODE31UuyWTfOpx9JGMUkiGfbRGuFd4fun6BHrv25Mh0seU7xP9XaGQa0it/tmzwcsgR2
USJd7Yju0ScBxT2YDPZEbPOq6u7LoLGjDCS90F9kTYgkwwNgRZylBYj8a6ey/w1xN0bnNIDFt6Z6
XWnYs8MGWPiUqB6qsylKEjnOBc5U9Gm3TtlftR/9CSoRzSAMwhwLbK4/FX1vogHgc0EGEEw6jILe
faMaeTU7JNtN5WzgoM0OVZEEidL9li4IhkmqyDNFXCqdV+ULck+4vgWuyqRP8oVG8id86uNwi8GV
moL1lV1nqkocTSkR7EyU2CTaUgxednZQM0RiDapyOchATFcSCNb45NDyY/Hz5Fy9h5piZFnVssh0
vDoBXjF3o/M4xLk79agUf7KGN8abffRYri1wrSDLVB3ZklnStq3I/xhmMMpEueIBhCoJYKY//hh6
O6RH8Hi5QjZINUHyUOwOs8v3X92knOPWoLkgTQ+rnGo83kHyhlpxY9e9xH7GFx65dRyXAjYiy3U3
5VtAi3Q7XXTqiSpEb6EKOvHIIwjNcj6SnrR0Qbyzx7V7lbGDeGnMPcs2WOVDnGsH3fJ1CoIZDPTJ
9wNXWQasAm3UsTHXrmlT/RDU1UIxyMTcwLIefB83sHpvTFq/BRF4kL5SCmzsx9gBFwc0+kfLlgjZ
+1F8Ml07agOd+HSYuY5r4fT0TEmXcq2LRBq2E54GWLvgnnVP4z0x7qOTcu6hH5vEAgaporyrlce8
RWUwMoV2mlTp3zgdQeCcvgjjsyU71UFdM38Pn1ZaBfmOQcL//LdJpGXZ9H2ns/4KZM6J8SlPKq9h
xd2dQsmlYt7pNfotVJZiH/GmPdZTk4UAQTxqE/at8JuBlCBoolfY4roGkcFTcP8uKxSsArcx3AnV
Clf4lMFJbK1op1HvJXoMgRbHyhiqrfA91GxFHKUkwwp4q40h+p4c3A7Yz0BekOdUYlXA7m0u5rI1
Znx3jL8PTRT7eeGXbHZ7CTbSR6Lcp80GW/80b0dFKqzBQiseKxNZ/lsPBVa2j/LU11wHf7IXfacQ
P71OPvhw5s9hwvgdn3RJ3LbtSkh4Vp/dT5a9zYJTmGPULoai1/r0utnTgqELmukqjENmAke+KEKH
v8UOJ9bGIVZ+7Ait/+ECqTjXozRSHcdSb1+0b4H3Zm4baBmH08cEbZd27Iu9p75uTSDrRunPSUBw
tGvAJA9nXotuorp1x+1sXrwSi1ku4JpegiP5rvg7JxmHVAPzs+zkRu8kNxziwFG0IS/K+zVYDYU8
Pos76ilnvk2dRrq9iwFppHGiZdBs5N1omM1MGEHVzmrKkBAjsWvHwoo9ZPkqTHq3TAOa5S39jexm
dTRbXNzJpKviqFr93WvnDT424RfL4vpKYxfQkkqDxAarbF6cBzXRBYcMKOHh5z5ejDxv7te2i4yZ
fWuDFFh3ZxSyKLVza2J22sjWYBAGiwUWnqN8aBdXoolk8R95cNB3I56lfBQhN3O0eHTu6098SSml
wRJ/DZC6xnvN0JpkTnAyMUbT3IVVs1FqQDPOaQArvzs4Mw3bJqsImSncShpnSCZ1tARmaLu4DYlX
nmOJ16ORYVxelv4YrI+QsKCQsRUvjIhxbmKuTt6hRUA2RefiJbzaWTBctpUP9tu1xOzUBsnjYkYo
wksxXaL9bpmghqeU49s8SO/i4nx1e9mmVEznA4AU49ojzrPlGaAw0tvBNB6jnnslVyg5Zq+TrNLd
+wgd2Lh4fMdFbvS8+bBXcJ1ZOJt5FC4hbqvHl4bYVrp4PoT/oQelPqromKBzk51E+QXhkQ9wl274
xMjkj7WgQ21L81W9VEjCqpYmV+MouYdzn775Y9KQJoma+Gcl56DhaRkpNAJRlX5bIQ+wORvenNjl
teog2j0GNYc0KXku3CsJt1C1k/tLsh8sgfsToHbNYy3slUme9NnTHoH7LP11HzRh2fH6SlrloI8S
Uc8iiTl2XzrWHLK9LdBJu2ah8FFatld+/+ttRbTHb8QW0lOVpY7Q+I3ccN5B5DR83bHYtRAYW2Mp
x4aedw/58YCPbhhtO1Lil3JWBm8sg4j1maZ849od9ocy2TuHKpHiu1fk0fORS4KQUf/vOykaP13c
X5Y68zt4wzKtwgtiXosBqhs3KFFw43cfnbdZOcHl2iQFsetg9+i5M0Y4wzor+nqivVGsnMI36f01
+s3JVGdtJZKWlci/476xt0+uic+z5Bhw9RHXydzHqABleS7CYR0n5yov5NcSJoZM6zlfgiK+3WNA
YLD8HdtXOa+FB5E8QPIr3erFtZ+tWDhuS4x0j6Y4C2Bduu8nd0vxvq5LpSUMDiaqpKnmpbsd+qFe
9Ah3wzY3mY1PLpCl007jWKJ+p9D/sSAjsDQVPSNQG+a0gTSqLcjiYWtno+PJgGYUNaC+ivLCkuyo
DUGdJLf+GaFF81qE6dNfsk7kbYTiQWkq4Iey1+YdvM+Ne+rNFyR24tx9KEpS0ZM6W2a0OMNsFuNU
GANyg2zoC0WQh9isUOy0ZC0k3/MkUSxnfTHXh0hlbPdyt4+gE157FjsB9wYJFEesf93kwI/6ZxIz
CGbOkD10+9Sv3lOrxbZ36ss67WKo0rVie1DN00Jai7bDjHrFIDKL4x7zdJiGPB411B6VhsNyIppi
OiZbE5vJxzFtrBkH9fVmbfLMvp2lPIMpWH0+BuqHfROI5g6YMQ5wju3nPtYfcxtEOdFvB486h/fx
W00xpklTIe6Rkv8qgcElCjIbPKJAasdv6+gWX0somQbXfWS8aFoKt7sKkFSVH++PedBVtTMlOFW2
phghjxV7Z8m4v6KggNfVjHZ5jX/Jzf5eX+wlE/BOfU19pwdcphXItRKCi557xyg2VTHpSBCiecCN
O0E+Mesu84H1wKNM85QwK2N+u+CBw3xwFh9wPgMUOGdEj6DxRsP77+6YoUZtrCGnk9ypsbKgc0ri
TtJ4EKmtur1NtE1hdPJj5AsVjvP9epuxSIFIbYtprrHY7+NXyj1tk0y8JqXmBPUSkIee2C7rQLNp
LCjaw7XuEZ5Hcpj7cPeAXTxB7oPacKBmMbbQQUMV54gfNKFSNBpgMFvgP5cVpbWpXZJQA0OQa99n
CE6pG8BWZ6XSUCx1axyzTWIKpB9NO0NP64iz4W1rlp+/YhVg3hJpahilfO1cCu0gNZuUsC03bkYT
yhjNv2b2idHX414V9iUr/lbqO/szRXW083kTstk5KW0Ba9FOG0vXUoclFN59UBlwz9mmpaH0+h7l
LWpjJFmAt6B5An1I8q2uBnA6CeCmDdEgY6rh69eHmDNxTQQYFAzpsfbmdJnNO9tnAdBY3f9anlR6
llvWwunHiMwgR1QbHrdXi1rlGdwvmqnOXjoczsPFANRFVyCHAyd+mBD27s5b1awhobI28ZH82oqv
V1x/NNoKNTJmEuP7kzCH9SH3gtrWbKf8QbCXX7IImS8FnpDRLjwqevsZey62I5rNN6aVVHhI3jiw
vvmSyH5oE0J6YElajMjS12p6gPXGzzTtmsRgxpZOC2SbMsnq99LGsXM/e3QyDpH0W2qJtuicHq2k
hizUMa7Ukl0HUOwgd1d13tl2KaIx+EnJ1RhwPWIQNBc0KQikSiflIvrL1egodceAViS8eXo91vlw
1e8cBM7bjGnVyGVu0TfTx5mjPUpbcabSGZJdS5JjhXqLyKp5D7gT4DTwrW1F9KR1LW/cUh305Ux9
RJLMDZHP1P/8y71aT7llYAZbqR/I1dbaHOvE6SY1+DrM6rUZxQci+oPCgulcvzb9XVihXnJHrZw5
dw+OxyjtdoFunohTxFuh3l8RiA72jwHcZFNf8FoxN5Yu4HhBJ2HgkYkzbZosaBfu32MHRICE4B9X
dnyYTWZckh8t73gRVjZtSFz3ARMfu4Fnongg6JcLe9sKxbDUoSgEaaAa0qRIgJ61g+rO78xdSjqZ
K9b+tAKKGidtFekfgpo9d4UW5Xu50MBFbp7FCyDrHJPEvhWPi931RnNnHE7C5BPexbJ5jiCMh82t
jIAUaHEkuPNj7SWORq0NvGoFqUWiYtDCTShXltw3XJKAso3n8uMxff5Pnvp5iei/SHdbeifZnQqy
Lezxi/NhmwlOxfjGm5BVcpqvlgAExOY7VLb5NEMFOAPBerK0MX37BdGorYed7BeHzhrXFeZ1Gmn6
w2ORAjrlUdgUHxp1/qGxblP8Tk1vVARUt0n8KQMCh9tew/uOt6KHsBW5cGMPVdx9iVIVOnWav2Kn
9Ek9SPw4EHlYuu0xR/KO3dKf/TFmei0kHdZ5dlpCcd4qac48oTSEC8q8rboJyo96JaWHi10IMp8E
UFJrznMWosjmtsRnBcMrLlEk7leRCRXm+gZlqQH2DZbWakhIyNGk889eoSYbTW3D7zdDlX8Jx8nY
MglW7MQ4fbEyF2QNlg3vBVnprcNM4yUJG6OhBjGjJnW7bDjJoWlQOMl3PhHxs5nLUXU4Uvz7MNYe
zKq+g0i/tuXuBqWA1wPXIwHWGSAlutm9cFdTUswutLjb6HRBpaNdAn8Qp+RffnLiPsoO8v2DLCIB
JWZYSbXU4xsiTZFQtcr6vGoBDM5H1waDURj+HOsqTK58R6V7qi7vctZnbT1nz+SarDvs0BZnsb6I
Wtmz5xHLKh/FceN4/i3bk+3mGHT+d0n5oeJaOrHFOJXGGOhPgGgWEZ+ZFDae8ug+2Ylg4WCnm2+a
34CDYT3tTJU6E9mFpjROadEqIdEQ0TUHG2HCXj//p0xH0rds8kfvMphBB/dun9q/lzh6/2196yNu
NYlJ2ixip5kPAyqIsK61cpbXuNRkTD/Rs93iMrarFwmwUM0Sfj9Hp8UWr5MHp4geBybH7DXCQFfl
IeuZQxX387L523GLKJnfiHMoDGR2Zbe4Bb7b24xDFoYsqwENruFXJTiy7BZ4Y2nELWZc6sT0mXPY
z8Bygm7C2R+14qWtFJNEO/72T7Ltk4IFrbmZ7iu5WcvvcBkdlwSMPZRfqRV/Fa7wV2ZB78OpDpz/
7zFGTYJi1fzFaTtwHU5lJs0z4Sa7aDDpUftYjTDh8zc4fRNsRPkZ2l//2Eet+syYhoitLQNfcurn
mg+LUDbbIrekFVBWvPGritlaLhbT6L2F5rymwlvPawR0CW7PhmYiw45u5RKhJNmfREwjN3WVLnqL
6vMWIoEmcquz54s6ZEP9Cb/WmAGvjOJJKlCazutOIzP6RK4sK9lag7mWAQH/CpsybF7eeIlZE7G7
G6BFanHo579TwzrWGkS0uNYkaU7LGItHkfRw3Yyum7z091LQuaURrHRqWG5kEHBo5OdRgf5w/beV
2wnoA//FaDqwG0QHc6/g4EeAHGP/bY8Pg497V3UzGqkUKnPNGNs1y3AOJFCsJQdcpRMIJ9QaXZns
oWkDg3uuf/d+nT0F5m59Z0fPoqlgV8+jnC9/j4B+yResmyv/0DCZdNmKry2TaxBRdJpvkb3ReEGa
8YR58aEcaWZtEYeYQ+N64u8Kk1gtltN5/L57SyW9LzSRJQOAiyMvDUQYBViFywsYpMslJz14qwC3
D9KLfl71hqFINTpecr+nGZCxvJHn8ydv00RQ2qaD5G+E9GLmkXuX2z24eLarSBGUiula+3T4unSd
5rERMhivVho6he6mqyDTFBKxJctrIiH+eU50JAea7bsJ9zlKOW0wMzw0aDX/Alhc1bHIZbVOEqDa
3COMX6OF/8KH+6BhJP3NBcl15dmEw3sXeeBBn9+xrWvK2ERHnkx+WgCrnmHIQ7xIZdUpSN1gtrSl
KyAwft0Fmr3wxN6rVIo0pYKbEOoJ0g==
`protect end_protected
