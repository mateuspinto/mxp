`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
gsYMO2efp1RTjjP32ZzFokZ8S+sSTAvN6xb7lRAZXvK2QMUPE5tkiKg0deERPrD4BD1p6s1/jN2p
Ca/AwUU36nunoECPl2QNn9eG/6fB6ECvbFC44LEfeqdQDHE6lGmacvxzizZQtvrbR8xsqNgQzaet
KOpdTuW3xs35/eFO4UlzWiQlh9kbZwSASHXUq9J4GsUhHyzJTYftGGdqtKIg2c0v1KH1LiRcUOPw
yvMpkAkqbBpNFDTmfM0Cwz00P5aE9gAph9uEqiJFIH8tlro0jVHZ5Cs/0w5zMgxowvboSHv2fiD5
7tJ5sgYQ2oNyDz6KjxJitTpp/FD/ZuO1HVgBiA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="UJGb8TyZxkl+D/4S2djd079GN7r0bEbxkUMu4YI6RDw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26128)
`protect data_block
GbRitbPvTH8I1bn0AOsfHphkTQBVAFHQc0s6OwD1EsXcH/O2qwdsVlXQs2z2leVYuyaGGXlzL8lj
kaLhqE9PLjvxmhrFzRkSDAvHN0b+MHU6YsHby2++VIX3F++1uVdlQYeMZzA9XK6bZlI5oAX/hUKZ
izx0LAr/7P315e0xLDqziu6NdNiISUQ70RmX4CW2kwU7S73d+fmw0kHBzFot6vVI1Zw1PI+o4K/p
W/vkip/C8imTpPsxw56/ztWRZRwHEJo4HWJu+HNvkWHAbCyU9d5LGFLfm92SlBsCqgOoWUMHYAIt
fR9pG7oPazdS30NW8g7nZCi7RIimepK0YIX+a8KzBaUJreuAZgFrbZu/UP57dmpvwaBN9n2VTpi7
Knn29t13coilGTEBuRqN0jxReMmI1X06EopvqR8qfEDe/vemBI7crJYyR3PYi6KyIRVsGhaT7TpD
vj82iQd2/lu1TlZfw5Ra64h67qvvThq+iSdkKYfC/59FrOTeDlpoNaboSzFzLarrlBDxzCYfQkUu
7W5ExDcVy+MsIWGL81mReOgVOsJVA9yI84Z/WuudjjqueZKXvDOxl9Cmow6/+wrNvO1MeHBvBwqY
oat8lL5kFunNTUQFl5gCsHf0DeX3RWjegwsXY7y18g9xscWN7BzTarprdvwphQlu94V+SAnOcV+/
iXDqy6RY7SYRXaEnanC/Qs6s/IMh4qDyMs5vhnS8+1JmCa1Sx/1UKiQ7LMhRE24qSqpYFb5RgHIk
BcbfLiE/k9loVesWhWVi4X6QIJgG9EOBn9R8dcaiHpbWO5QJvDrNZOiklzLtUT+BKfRkwQtfXi9n
CVizGIM3mRpjnmwJSmu5B5nI0criSx2qhwBVKtqzJOI38swtxGX7BhMLhTzfsRMapvbJ1BRKJEEQ
/d+jEZh99MVj/VfIoqi6LnKD43YP8gjKuoZV64RvS//ORBIIghuC8902pBNFoe5REXH9oAJ4pP4z
y+H6brCc8uElwbL4icIQGoVgtP872gLeHK313jxZXvm10YHdWxNM0lPxbFqWK8MCxpfFOi+kXLKy
echEZnl95mXmcFqNp5jPedDTcw0k2/hEH3BzzVf+Mo9KcCDgV41lnCt6NRDwsuc+7mU6I6naQrmP
NB7Z0EXIoswfECxvleVl2Wcgee7VpoKuVJlRroKkDAlgvYQ4MwE778SkoNXAJM9jaM/QXYrUk66U
oF78NhfSb/dJbQ0rb+BZ9sVddlhgXZDjIPA4cRm2PFQUAaUm4uAiwCTqpOC7fQ9rp5h4jaIKc3wc
TotoqA4aoFbq6trkMXSlKMeUrvqjOYUoLx8y6Hotluz3IsyFUtq92FwAQntEMXiXvctdWR5XLVlf
KLcpvmM66FN0LgKXvi7n/Xg0J4EVFlow1SgW2L4Bh/obvbVXphD/LqiUqxmh4IlN15Idbw9UIcMb
Z8RZW8WmseWuhZ6Adlx6LmbFsEdQFVFHOmcuXoNbmC2+7zZOTz3pW5Rc4JFR9xV0VynwoUqH1mKA
VixXTG2i5mMlW18QsJ4de9xmDnuQQ/fVaVPIcyFLCxRSeAvACE6YkWe0hbqTlpkBshwf/HgAGxXZ
Fa4hCF/mlPqcAQCyBKxMPT/GyXDCBYdqpdTFI8j7JdPmwuyT+XeJ76Ak4VVkitFFpRB5nInvQ9cX
EQZu+ufwNivKzpfRZyZi3hJkWunsonqhD/pMWNX7XKEV5ekVSVo4mxKPBk5xqC6kgyfbDbce93mj
I0zOghGe8XXX2P/+yxvnN3ZuoaqzhnHMqkex2r6G3xKg/vaeinu83apEVokX9zdeiTlE8dMRaUoU
Pho1KxOdfK6KOWPgnbC92Wyee7GaCSr1iWeUFjyrl5ywqJJCTcUBWyXDEVSDFMLqlyapXWqoRMxK
cG9LdiuXzMnAxsLuIhUVk9vt9UYwva/kAWvqkf/e5XcCBAzhKz0x0nCflbizypD5pzi0E7B4Wsnl
AU333M6P2K6AoSLeDVdmAcqY9mSiWeR5R/zbhk+wC3DA3YJfKq1rMB4G6dZ2OyidsJxtgz2Y6KED
ip3e9+u3/HUxLjtmbXLId6ALowMzFYYx63wzOxQXsRuhTrL07NzAFKECOQd8R8B6tnhX1USAkyaE
bW60dFLDDUWYSQo+QzeFlSzqA8eNascZgQ9h5Fd8fFR7TBM4sMQyRQWms3pM9H1ima5ftI1XVQmn
0AIyyKZ93Tnm1u+tebcDTs8SxwiupNffyNk3JxuOKYf91+6O5qphf2miMcDcfRtsVgYbieZkBwjX
Cda0USjHtBiaaBridjJBsb2ekbEjYW07o79Q4EsyaMD5AEbDYgPB1ia8ADnTm5+c6ai9Tn3CS8If
6ltaHsV/TOz7vygyqsMy6H/TXfa4mPeOExOmN30/UfE6Khnu2EsoKX/RqNxRzMljfiyAzTeI8X9C
MAiIRpf5IDpza8YAl5fRCA7L0a8zOGTszUAHO4GLt7zofgVyxxVNKEa3lzozgvasY72igvYElCli
hjPuxc3f4vzz3lhdYKNwp0sLSILayiwQElSlFNVChWS+uO83Ffz5bUwNkFu3bSaJoidAST3d1DoE
OoGUxvQPuu3zx62cjgmB2y1RhYLq2Jw21fxG99QmJUdPv8mB2Ptm4XWRJLRFS9Ho7WJ5eNAP4VRQ
nheWBhT2zpii9/V5xuqFJZudsnRFm09VI2Ha8itJBQUqb4cr9XGvsFe+PF+312J7/IfGg6FWNzkf
Cp+Ie3n6t6vONjj5Qcnfd4TmrFvGOK+/n7ypvEq310M4/0m146ANMJzGtp3uIB/qtMR1aaTE6XSE
8b3OhUNhu2nVHFA3KWPWwmI9GsiYpdfrE/PTyaGkaN0qdRhY8k+cKLpptYPGNvUsbxaTAU251SrH
daJE1HY345W47rU1aip3lerqUmKm6P2o0AglH5aEajlSEcJmqEkTi1KZqTgULwWBzKB5ylXvn6Bh
diUGG4UXVcmtDDGyNsKbMyGr3PrTh7H91soPd+fNZkoc4S9VLUYhEcLNSRCemVrYi4aXCOJVWrji
ugKU56nIEykW8PB63ym0h4R+XuFWTl5bLVgIUFgjFYfxwyOStFhxhfstRyI4Jtf5PoNqcAbugoVL
GZiNSzaOuiZLgOnfT92aRFGUVdLik3J8p/sXnd7qT+pBcnR3nQgNstYs4YkXNMkYG+mriNwHWtoL
OTub4obPKW/EikodXVIK2eYjiEY03J0j+AxKJB6dLmrVrWLmoqnegAX7n6ZBRjQDH/Pk0ekIE2VR
2fHt3DnEdNgbm84upLnbuX1/CuLFwNfRNM9554CysGwO5wUK3LIf6tNZWP268k03nWYXIBLzt2nm
zHZSQrZnCl8ZDwxGw88n3ADkb8yn12oWAS33aLms2tjsCptT4fqWMrKYojN0Z90mjXEKQogJgw79
xoPco1AXHcDIbVws1UPzmP0kRHInfd9SmNhXc40ckGVhLFmJg8VMd8M/kRS59vdPNAsLV8SHRNer
qmXIzSL5RTr1KV6bzQtJFlFZ7ZMfA383tNikeFhIlSLY3FxDHvd5Qluuf5FKUvoRgphAYCQ9EuhT
E0N0vwwc5ZeHWZ/79loGSlMq2Y3xUoSazyw9VLfGOLytP4Y4ptsxCjX70lpn7Dd97hhXAlurZC+U
13urZKEAMI6B5USv1uS+5ZWQqsrvYD8PV3dnb6TA3FBSCNJsJZtFyH1vdw8clKa2awNv2V9jLB5C
K8TAh4m+PcIaTY9qv+NLqA+PoTFvkdcoDFAbbwURSOeIxDawQdGpZpeN53ly6UyAyXp0JS4tXG8D
J5KQrY1hlMbJytjWPogCnUWXDlAFxf1phA+RCKyvNARI1r5K7uOwO3EWpdNONx2duVtQ4hZO3cxb
IE6PM5A2K6PWjOEU9XF7tGho2mPq0eetwjraHsos3VXkltotDzz774wowQeOU5z0e7yXX3VkAk68
LQVFV8rr5fie9MvYy9/MBxGQ6gbki32aeTOUJU8DSLDsT+xmtqjRfHMvQda+ewQuVq85ZWQTlvRZ
iHu/7pAYjWY9Cfy2LR/ecv6Zx3q8MYXJbIt4x7DcCe3MvVBKYF7RNmF9pJXvWUapLBaQKPCaKsg9
4JfbZ7rFSAh8Pk+UyLnz4XoOFCv7/2TYWssgLrGMFSTh4KQOVg/iIAHcYEqf6qs4JJSEGWWyMJKk
MfNXTK9sK1doP2Sih+XeC10QSAwqDc722kIfLGqlt0Wsy24SrjcK5alJJFhXvLt8OYv4ek0UEOky
b6x7iLX9riS26Tz86NPZ3NB4pz7Kwn0+xymDDh5QuF+idFagCfN7uMLW96Aeiv7d5RTj1VfC4ZUL
7/bInTw3NDFkvJp23zETQmatp6RBfsm4awQbqMPVIfaHxOt37J+46V3Efq6iiMbCoeqzE3vaLG6f
qd7xTTs0elpzo8VZGLcD3IoF2A+013ngstnzq3SHDSCSfeoc4En9HWZmsgeSzt1mV0wXCrdDGbYO
IiAYYNtae88a/0Lbds632fTBRXgLqXFvtaogZuIOXkq7P/B8L87FLgotJ3j1LW/Gb7b9HLLqYsV4
zQCvFtKkkL4dNDVF8OZIcv0Ajqg4ITysfyqo2ziU/vgFbDXM9w2+ABQJnDTs3IDW9gyKSSOXOHyO
tDr09ST04LU+PLuAOCl9Sca3fyov80Qq3VOo7Q9VSEIQSF+cQj2sd5LSb9zf8N43d486ha/i5etI
Yh/NUvx9fy86w5zE7Ra3qPIbGMD/3+zMYXv5RqkJ8VBKrPvE1dx5IIjqVLG4yuh7CpScrpFc1Dgr
RSiDQntxJLCVQbyntpTQmgaEwq7Kc0jeIJP7vqMWqOtfpeLwInXPOlHthDbWwhtzUB/EjD59YJ19
wtQzdZX8iM1RczEufx0uo1zAteqFXzAgu3rKxt+/FG5CRH6m2UhK/JRz5s5R4kucXxEmt1wedmuk
mbhmT+c1GbrR+HqQr7wCt+ENYRopferoSfgclPmEOcPDU2MSYxsBo7eTTrK/foLngy29Ww8dJoov
GRrbTheGaWur0KkyzcZeLMLV460ne0y4VKMLZPKQjP7rEUk69OlT0yHAmiLukofpRZGRfNuVA73Y
QRCv7eduDoKomLOvrHMsXcCLlUsKDoIN2SqP1pFR/jFLBEQsSpZQq03/ffIE3Xi73ySSiGZvpHgX
XJdSji346iyTmKEh/MlsqGvufVv/LPtQkanaJNzoTQUAy3LEZ+Vt0n2F4rg06PgFJmwu1wiBa2Hw
8PQozw/tX/lrqENPkOjSysOhdyKkWPGw7hhiBgJ9QGMwfWahYVqpCWJokkkHZHAe+CoyaqzzVLB9
3l94YhB9AlRu9LnFn6m+Kdf+3RNPbeqXQFCQvR0+EXw/cW7vSb1OUYUPU/RB386igL3p1QvTbs2B
gyGrXa/ziKaO8h7+A71egnrx+scj+6VJKFu0HIfEtGNuxX6dYwKfTFzNIrS7rA5zvvPMyldFz9fH
41JQz4qJhfvnBZhoS2g2MIjLwbBWRYQiIvk6lBvxBmcL+PJJe576DoLgtsjg75a3obs/fs2+1gJI
Dxy9xmJI5qCKw7tSvVH+oFBiCc5qoOWLgodwI1SmMY7SjUFmYtu96Ee33qhFtXVlpatxsfXyqsk+
Xlu6na3etHn6dvckMClxJIpxWVRDHzGUNePdYCGUUxoSltlYAh3G31qYqLX0LRB7PKzq9KBlz0aB
lDcGo2ZHztlMCOvnhIMrD4pI0cm42Cmjgr0vC8OmWkb4aQEmcc//4bAuTRFcUK8NWBb3vNpDOUJW
FaiHLMwbYwkfzTz+eumKMHD6dLiBCYG39O2Hai2TvsUKBFFMssGDGfv4OrP5bmAhsFfa/a3eT8jt
Jw+hOfcNcepaijHtgHIE0L9pfrFHOWGdbqmET8V/XQmwKFbVPSPkCp17TghiH0cZPYPXpnH5hsXR
sNcGKP7ob0X0BaQf+ev/f0JzzudmEqT5mVjfWMhh6alvXVc2Fd0WXUd/hKId7ZCpix/oTctHOUZy
+/QT6haHorqn4lOuStX2pwNxbdkurY/GjAsx/5u3tTDdKVOSDbtY0N2ppdTmAuoAmtYxYnBVfvjD
wOwhWLSCASxd/LuwyHiuJtxxH1zjago6I2LoNzNogGR7GCMbY+sP9dcCuMiqxLX2VCpmDhg6T0Rs
8j7CUO112L6AKdSJoI/xQ8/ujQveSD/7rASmGCTAruVQfZ8QX+eGzptH0Ksysuaz0GsQWGx7dudp
xdBDVHGja692dHH0VeYb+bNWcdHG+RiVbOOhPRG++r7IUr3jZN6Fj0JD1xKR0NnZ0IMGnUmGDM2F
Lcfg0PmdRkUkc9V6N/pVVWRvhp93o9yKiSlt+fyLkIf+lUDWWsEveTTjTDcCah8NJe0bmk3modjl
swpRq/cfhWFEsTbCuno+ftYLH7AaryQCV4Y/vLUyFKrRZpvqXedLiKYxXhxIoW9OQk1Wj/yzbDiw
lxlYLyJ1Bzhet7CRJjCkdxM4wQ+x9oclD26d2qRa5gBfg+xQ/IUupvGOUvZibAyRK//LO+B2SePY
cTnRP65uQWBoMr6R3lmmgF24ZICHJGgO/2gMg2YL2ZSpwvl87a28UF34PHWQ0X2g6K2Kjh9GdXl7
XIPu1IpLNNcd38q/VMecBlnB9NSwloFkrKlM3Wk+ehc3vT6xee/mgZEU35AbxORP7pAi9oK8O66S
YXbCpjEzPcaCZy/dUKXtJM1o8C52rnETZ6WSDzGyu/+wdo+7Zrn/VnzVidEj9mMqEjCMRoAA/OTC
f3QaEO17ZCOjeWDe0k+OZ/zD8k2cB30lQ63DfE7lDBC1RjN91FVMPuqdc6X8vZDkj1IOlfMvJztl
K23oi7GMzT/V6xMQDds/wfQv2stnf5OspsO7opZszcoxMoou8yepCQbkX/PddGZ/LyIIyalw8fuy
jQgEdibDERi0F5J0hE1Kw+u8l+TF7BC5m/7ofcgJFTKPEqvSR2qKvQARujuA9mte4akcdhVDAaFH
wkZ2Z3U2nyoEN+I+qEhmg2mRbId76NRy5mlLNTPwLzXH3WjGDAQb4eClCq9AlxIF0Y7e36d4Q1dj
22ghyHBHirA1yLG+d04yJpcWPXGOIxXj5CUIjZAKI9lLSHEq7RHqmWEDO2/bugw0spIkF0zo3lSm
74/o/keI8PJBOHuNdAxYzom0LYJ2EvO8zFJM6h2pWvjzTNGd1X5bsRjpitSaaGhdpicExMwvfd0K
hmAutYPMJ1e/UaBKKgPIr6wLDGGk+nHFRdDs1ev+Y6xLfYUHpXKCsmD4n8Izb7zoGpR+5GGDxkVm
OSe/xzGpkFx0ZeW0MtQQxFxoAsf0+ty2qnRRQliuUUWPnp4UQA4vCiEz15te3xjJaD2resdz7Fom
gB++boq4KFTrmO/v6bIzpkNSQgMQvckkvn9J5ayzuIqlbO98B5Yi5PwfWkTRAXintumJkTD+BTcO
KpjUmwO1Yy49GOC7jQrxRHODyrV5KtgY02FyguQRcETpeJhSpyUOeNXWqR6BGag/sU3tQQsZ3yuU
0lDWM0wTKnf945fdr9r5mfSxzUpjWASVk5VJ0u+wnZ438+R+jfHcWFoGOM2sW12IXXHQUG2WVhi+
lX25bLF/2tqanGvn4yZU3dbY4zZ529wM3WEiOyAouB9ewgSjEmPtVgEfCT/lhoSK3xwRrWe1UVcB
rALc0UFUpuuftFzK+80TE8JrqTwQfNNWyWrew/8VPBlOGjcWVmSkUsf62cSvsd4EuWj/Q18hp+jX
PdHxG9w62LFGfYCtMTgabwbGdSMdr0HMUlZKrERiYsJLelp3Bu3k4HBvVW+B+2GGixFElDKWwv6O
wpHlfpxBYWpOASkxYcD5DFFF6NeIZzZPZweQTOk3DwLLomJZGZdKJ05hs1yhs2XSNpy8j6zHXXHE
mEWcwY2QmTnE3qiJD2/YnpN8W/7KZl39gn8a2pEfrWRrF+2GDc2dxD2e0J9uFCCeCorwOhLvBlUK
TDremJOy/ciskaRFqFvYu+euMr9SzAz1BHcKNbs+Vl6LVPmCnUsR4jvmhWi+nVQ1JUeaXXIHcIw/
joY/p4AItbRvFKWLE3x7RwdlOiuNj26+AxNsHI11h0bz8brmRx8XcKWJFQawJS9h6YlnisMFo+ht
AsIdH+qcsfEs9QGNnPFzx9JI1EPjW1LcOl5c6y7GPs5Z7huEb5440YL+OVwSJINKwNjNJEc7xsn/
PX8bmtJEPx+uuSeq07CG0iwd8dyge2Om2BQ5B4jURXPNsrG0NtYrlFO+7cB792n3tASw7XvQB9z/
sRWKdkVAEbH9qk20AIopePcMXH4N1rlqE4gbnQqd0rhabFJCA7IExkmf5CYszFTQCWTJtWvYDaHK
VSOTVD51AU0E1SuH7lGWcTSgGmxkJQ64uP6vzQK5LAA/pfRHB/CnCnjhqPBjR4oF7KV99dkW0rM4
CMy/Lm8zn0BX0KTcrRmNsVH0LpfKTVXGNntcRUmG3Fp+1FBTfB5X1VGhYFJgVURY0ZsI1odPzZMm
K1LLf3cdWzKqC5FYqygxeUNBIbQrK6Q73aQORBV/rw2ipYt1kcSCjzVFF4anCcmC/iN+k1hkFdQ5
lPXwdj+6n53BW0zaLnyLNZMYZj6R97JRY6Ip277+thbUBj3R8kFlYmPCrL8Fm/I1XNquDnoM1J3P
lpOgSGYr5iNKhhk4J3Uq83floWLshf4dUL05rpLuk/3RwoQ83RvbkwR34w/GnE7xKnWiyd5ocVfT
+aElhl+FmlImPMdnJjUcUR64LVhg0LOgDCcRyTGLGqFF1sTEbpmx8PmkqYfAbPWWppfTOoXaIeGz
ahPIAmm+mlAJ53dmIQDL6Y3QKbS8JsTOrG7pfKzWKmdwFtLjoaiqN8nv8N53uf+MGf55xw7FYYAy
AG9asmKZ6DtCU7OoaJhp3T8alsVYGqAif5BUQAdC/6XrXbLsoANNMfNeu/AOy6X1hLC+y4vaYgI/
3jHg0QR8XyGLH0GLjQxkp8y7iF0f45dmZc4ujh3uFhkpPj6TQuAqJV8wgr2REljaeTytrc2HoUlc
213RKkTFtVgS2dtBs2hrGGQ1y7UYon2yQHpsGK2qHVguZ3Y68/KbG8KgOCXObvtsOCvmy41Jqzpi
dnAiZ1P1ILq2rWtg9YXFe2QslbxVe7oBWqqaO3ifS3hWVi/QlEBtrZY7JzHW6HMSMdtkCwW41dpG
K5beuVrieeVI+tJSyjUzje5ofeEwkehVutO8afWfBdCGeFUbbsD0vCMO5GjydSm6UsnlA+CgvwL0
0CuayM5znZoVDmR54LFNVDKTBn48/lo63CqXzNbnF6rZu0VdbZToW7JLWqjg7igrrtbnf8Br3O4m
hTfiXvqdIInaRIhpT1AgpmHUMJm9ug+cF1xEIGPaW8lSu0bqAnEZkWah+LJARrT+KFMcul3q61TV
Sk3TLQliqMWrCx3MLHLNu5dPaKI8nosTWjbvbu5vab3T+0AjZKTKMnHVOsmwLXjm6J5BNoip2fTd
S1zJs9MPDUafU/M5EeHQNmNsrWEvfCTR/d+LEd9m2UZ/w+9GKVvX33wIglEm+pYrveA4MTBitiDm
HZxpV2gzvvJddvptortnqK3HfeezWk6durqkuM9tv8mCSwHkCCsVPY1HK+OWyQNuovFc+Zc6+YN7
3u3e+qj1JkkiV+teMTPl0uY189Jq+YhTsI3vVl0vDwlNATukMNyI9tPM/ke4oCQ9lX/3x1XdfGXu
yB4H96ux9cFwHvYzs7hQ2nzn4zyjYJD2WSM3tqMnybYsmnuAUIPO6gcfGmH43KcnUa23SpIKQ4u9
OfdoFFyncowp0ZhdnGQrEJ3YwvFW34kC/BCnB86PgzaXVxJfvrXpYzbTIkDf5/PV1r3EPfXAp03g
QWZ4e3EEZWjejVDvfnSeD3eGSvc0gPlyCGfdMIkyKB3xeIP9qMeMdy0uSMCGF9qoaRzA9kmcHO1p
AEHSofLX3G/7laOUt6z+iDAD5KdXAdyKFEQ3Pj6X0SkUbx/8Q/gSwi5tbh1BTilfs2Us3M/SdbrC
yRWhhNQMzJBjlEOQ2SKFHs+sCn8iEn2xq9OwMjJmLMayZ2O3hyw68YKEdTqAySkmTmbNcf8+9x1R
4uZOnlCD/WA9GL0GYEs8f1Fx7ZdSQ47WeL4ASbJbqufhxxbp+ZkjjnvZAcHjj7PfgyOF8K5TwBfc
OLGIHaDbVNZBezvkmAlt2Qe8vnsLAqiPiuWj2ndUHd/D3VlhN01tOri9Ip8EC7c5frJYG8zhe8OR
rF+U4R2Z/Lw28imiEO5xMbJD+dNsHmhKaUfXS1EZTFWLwYjVicHBTQY3W31nA5zRWih2aUBXav0V
HTXsUVJey8edx2uXV29zrV1vaCNT5hRgBwOr+6StgnYzpUQEUsyCWCU1Z6TTQAOS3kfgKMWhyEEX
K44bDxslrl46O4rhDpu8dUzy8KSiErHgiStf4Oetgm/QNe84YWMIygZHWSlMTm3e5zjWeCVvCUg4
pZ8WrT7woeDaDks2Ef121qSzgnEfBUc/F8o6sphATQV9w4rmy38t4fIuLGXtVie/qsVtbvX7+sIB
RVHwsHmg3esXkzAJ+SkEkadez8svVa/JUKUy7rckl7rr9aDMp7N4hg6XJg5nD/7jPbzdCfDRifDQ
njhF7RqnnOcKX3zErxYQePLQk/8QNNmNl1lUMNoPnbHS1ILyvIFvNOIY+TBFjsa3VGM7FebNYPca
VmuSCapjUoqBUUlFx2a8grkY8IcysVB00ZFTzWUITNSxlAbnoeAymFW3JWMdEykkLfm2TiXDHlEx
W567ogaxGaPXmbgRO+K/fa7sYvT+p3yEGY0GX6D4kvJNcBR22Z14WC7mZwBZ7Ww5B4ztDmOMxTbT
zosAqCM9Qh8KPPfEBK88LufPWYqyxEKE0+/Af2liIr3zFgboBHV77gA2SSJQ2dquZ4JJLOiU+0Lv
etNLh/ihAepfqK+JIkNnp0t2cG4WUrVBm+JAcaMScxTFECfc0HcNY4bMO0tBLCNR47QZYvRpr1Ud
A4VDugdOMtq46oKlmlu+gxpnViW+EziJXNzk9o0ZNkMgaugLC4D8EWkUPzRSfHfyWBnmBGzWqGZv
0XbYOU/Ay7VFDtgW3XzRCJpd3Di6Tfash2MKrkHEdfRpBmWAxM0qvAjKT4kA9vxEJwpua3DnY7p5
/cWBt+fwJcEToUSlvt1ls914dLlRZXnES22jJhd8dKf8P3IsFDSF4UqjoAQP2ka67iHiq9zOtsag
6ALX/PFYG7YEvvORLWr4m9xJd0pxTN87F6zeXB1tbUz2QfiVAwTxHZqcctSpDl7phbzTQojhmXBu
FCg80qS7HKCC5RIIh3Ouh2WZOA3urrth2lC+fiWG8X2pG1rjOSntvlbnbLvEsVzqmfjtSt1dCFMt
b96FmgxMqXTfD1zTQ7t3yhxRkGUoOJCWNYe6BHV93oegNItZp/Daz1VjV0uys2MhCPZCeSnDNxLR
oVxpz2tTmw8+GRqNnQ72KvEcG5Joo9CvkzAIi96QhNK4/WHptIbuIpCapxs2qB2LMQhXehjbMS3N
7cg/R7jz5MB42ws79yCl+DQ2CBZlQ+usxHZrU9iW6udbBP7gDc85cdLBwGDZ9ecMGfujZUhadXSA
PcOfZ7RIychGN95xgHHIUGqs8t9abiRqLnJquEb9VZE1ftlNirCL1n8w1XZ0NvGOUVUmuUnCYC5r
ZCd4MU/UZOasFZcbGhw/S4WqZ0zu7uhmZ/Vpa7juNas7fvnhYJn1ODGTt6oPZfyg7f0nxcYuaqB2
MXZ7je5PgC6gDpHJ1uxNI5T2a5E0Q2RNxF08Lq01cMLrZcGp9p3PWj9unc5+5iPUUfSnpGINOmR1
F9BZuEyDRyzsxhune7QOo1ZMxMGghV/fIIv2APFdJskko2FzxmQ09A6lqEEmoS9TkEsCSNrewF4u
oOtCEoG6CReWHoSLg06bLWjjJxICX39alqGaWxAtpT4P8kamL+wbG3DQCnYcTk9C+inOlv7da4aZ
B4dRCBC1o5MrzipEZN9KAeyVkA173Dv0Hauy2+devvcc9hR7+rFtY5LqUzZk4l9KPv2rg+0OpXH1
L1hDHhVQzRjAq8ZUy2f7Hy9L9pU6xhElOIpW3hgYj2E6UPLVSE0vCldI+C8rH8+otl8gFds5WJh2
IalrbO/BAAVn8Sbnek2lWyY+Kc8UPH8RAEsWIw/QcLZe1Pb08H/nGPqAikLDvFj3zWp4GqRoJxqy
1OtqobOKZzUjiJqKot0ll2GZ0ZIsx0WtGxb8uORZ78N6tj68iVMHmxv1OB6RSpbflGLsTfeNSg9N
NuxeqLY14WQaqtrRLYgh9UdQiVlSm8tJCjsudk1WQTcVgBOqxrBoOd0j7aPdPNHa1fIjBwXRfTlO
VWyqLVyz69Zdo1mBYNfpILxrytd+Acyl3bTMlvpw6ie2vRPuk82apjkgbnLzxJtG4ILevFDbd3MJ
7VchTvcOVJu/I7hyOiRyvqdgerwQZRlhcvOqEtmBoFXJFPP53lzkUnKKDsEQ75hbjSomAMEAKzKi
KcCWF2aScE7dHEbCbdLpzFc7IFTKwgFJuyXKWTj10IHG2iznQsGHt6YWH2S4Bywi5fESkRKYZeDQ
fDX4ugkfzgeChMNSQnDMOE7f8RDSOSiJ0+7fW9fjOg1zYU4j92vkXkhOlfgPoeIP99BEXv5KRnH1
wtbU0peXE/P02FaKEZm46/O33teBA9pOY4s3HC8TxvlxrzlIkL3A5XtW+ZmYinYQkd/u+Da8CFOM
q5rALTDHxqTJFhEEP3VzjrOgyH5kooKEh1X13Gcfzvqogw11MWg0i1KYi/K/i11sg0tfS24S/mmC
ICvTPtO2GDqqlXdpuNE+ajuDa8xLUT+tug9oR0VVRTm4dcKquCdYk0t1YLqC1IoqiZcA74k/Yqe3
DcVHC/K5LOqkZOcTxqQIDuGb01nArCWylofsr98V6QirDLdBbCxv0+Aapafd7ckzNJTaQv+NNXIE
8e97ERYomX0dF8r+oDs7z5JsN5BzRppJRilIPt6257qfdGDIZUBuDK94LUFDRdQeiG2Lhx95bsn7
vn3pEFJKGbQNwEdLHx92dUprAOO8hv0+x8p0UWLxMNJ8NCB5ohnC6yIZcoAB2jton68FA9975Lzy
pq/C70EY0a2jY9VvWm0J+93EI3cpii2xSzBwJVQoxT18ASp3cMVPd7DXRNJ4No9vbktX84Uzk3JJ
d+yp9CoMrrJTfXIDKSSW2JQI63CQu5zcrf09qsQB05t6W5lDpKfuWgnrMkIs7ZfCAxBXBhCpK5xn
BeNgxTDj/GHScfqg7yFK3hP+HfSAu6+cd+A/eW/qwJEh9K4L/HtP3RTJoDCyMWj/0l1onO8+cap5
AEM1coOwBHncqAy567ESY1zcVgJ7Ut79avwH/ya84QDpnc/F89UNtySSGDviffG8l2tRbeVBISHd
dleNYL2ThwMIvt9G0AgpAatKfkM3iSKhnPhCMsVRhK8GtwWoTRcSeg0MD5vz6gKW+AEbv5JrdsWn
ZzbLK8OE0vs9EYV6sBxNHbyj3Vjccb00W/9BWlK440hhs77PexMWaCtVaJdKsutycrb47NEDrFry
hm0tIkMNiXYQ93hfEqyaHbuP7INNyUomapLxjbZ1AGcML1dZtRaYNph0EqZifcb1ojwmab54ld2z
3yBzw5f0Ww75Lsz32oxFcok0lXY1I6rhPwDjnGw2RFZqaPfqZlb02oy+Qi2YSwGVOXI8MvIjeC2F
/W77S345leq3zTIs/E21ErvOj7rYP+asfJVVC/4BQJWeznTQxd2bQcytyJ5aa6JLHJBRo3oXUh6q
bz2Zp+pEy2dGOkGpOAdmgkjpU8UIqm2Cv3YUEPLso8kicm1/OMwRmOcm45ncTM13QUtxEmF8Jjvi
8q6gyn+c7ec6GGdYp9PUIFKA+f93VMzcUyXCkzn7J7QYGIKYE0EDqoEyohX1+C7VO4CZTCX9MbA+
Me7IB3ulkAtPqW2NEzFa2rk+Voz0lyER+esSh47B4KrnxRUPkaSA+Gh7ZOjeo5YsH+hBLadi8gvU
6FssQM+ZSSk3f9KcmR7vuNOQJbeazpPFdf83neidwmBSltZHMrN/+I4WGiT83momuChw85aQD5ve
xLBFvwt7tAG46zKauGkv1a0qLS/MoE13qSDDPCisApr5rnORXGjcV9aELBIwea83dzdNR+ZwnW3w
kxzE3/W0QoUIT+UM9D8tyQGfzVCkn9PTcjvvgIQys3henS3FhkvhO9HLMXcWhUvzS4yqCe4xojFf
BAIIPBWnkQQJyTnhBXYH/hxqOGUNqqU0xQ2ZeK4cPGLDfZRWZTRZbVEWAEc8LL8RottHvtLirfXY
fTgXOxqSoi1oPdoj36Ziq3TBddPu8zltdS+ts3Ip7BcYO0cj7Vu7jDrQxcpObUS3Udc8zf5jNaWw
PFXW3nD+aqPiKYOm6KBapPbkCoCfZzTEa1RACxtiaxi7cYatMEq9BK5uQ0MhnHTnK2FvPcu7NNn7
i/nP4QYWfaGg2uKw8KSZe66HrVywpz/c5vX9cxfxfzZXbOt5WJBi/Ph9SahyY45QJizDVp/tp9Aq
0PMXCrkZH4qi0lSEk5ujmZm03rpEWU6cyQKd2bs1jMWOB+eFC8TUhGvcLsdfa7+roBQiGF7ACVVs
JtW/Bvn8q7EOBjTNjQPlX5iKZvv74GxTSI154SlAuozT4+pUXmm0jJa1MZhExLuE9IIen3pVeq/u
6EOaaVh/nK5zzEbUPKtTAe+AmtnMbthLNGRmrNpohqKQlS3LaHHdJues+wrXXhFeK1o0rTK9cOED
4/7ePSfMhr+GWJSjwTbmveOXKoveclJBUcS1NwEZhGrVgMDt7UpjRuFeBgPoWJQttPfNDM0FxmwG
w8JrgbOHYEzPmcvh2+/mhb6mV367Adjz5Be6VhG75BA5HhI0w5cotWhE/YYBDL2NUpPgJ8D/qspH
zbrmohc3p6Co6d+B0uwcegGt1twYgxGvlYbzYexxN32w8WwmGWHSRI5FeDDb4CREtKKw0RbPHmYw
I1OftVpdAv7El2DsgLLegpWLgDw3ybmwOxuP/rDB12V5snkMFuNPkukkjiTExFeRV3ERjrmPp3y8
bZf8X5rIfiFM539YBP9eT2cMxjrmXEY5N/k8PLC0UGcxWKNP8eecxogH6o0uKwxHvfXWlWCTorMC
jgRKxCwt51qid0WrPdUMPP3l9qYkB0prnxRqSeNOeQf3inLjqMzemzm1v2WhNURLK5PsXPk5Y7J4
HBha6RxXN0vpUrBi6s5UWBZkv8TxdaIpoFm6fViTlkJ5cwVUTcgq1ykLdXmc8Uhd3K5/Ewo1ChDn
niCSg9UkcCYzNl//RoDWY1TcVFOZZgfpJ+PgjHoFRW9QPkq2CCDiTlM5mkOLvrJb3TD8seKIJbZb
sPFT5vZfsso8kcS4hbMOfNKDUX/DClDL0cGTG1by8LNzsKptE5fANWR6ZWHVkYPjV8K4ZGJH8wOk
Ca7nypef62DvusZpYvFqqqiLZpsJ5XkIuiBYw5oClr4FFjJpnb0E6QHp6FFeNoCCNJXfalT5sdFw
j/mIzVQoStGEB0rTjytHKzOOQa7d+Nayd94je+IbUelWa9xyWtKnbohg6fWlZ6x2mIezZgAaUSbq
qkwQQxMJTnUyMK25/lLhY36GkJ1H0eowdXC/Rt7i43YjupNDehCJeWVRZXQGG0Wh2ZPb5L9/+vau
jvx0MVSc1JbJQK6W6mXFsMMXXTktqfOuwDWzw2b6lsKWGuEB2bijeNNCjwujL4t7hLXymWYE7LnU
6M5GtYM4OncKSrzPw+ADAyHW+TJyH8jO6vNmFryicMIQ00NL120Ui+7QkS/G96jVxB0fmR+jqHlI
49iOLebKcCqCh4jN3K0loF/OVR/dS1aUYecSI1PhC0SKM27tgsTNPe4OEcO63XGoCIacBfxe7sHi
FRtIC5aHBtrQOc5yVCNSn4VHBwtbxWofT4zbsfkRaseTAMRjnenu3jOmw2Z+lYqdgAYcVJfFJfnP
PaqFL32gSHD6drp+nXW6oRmMgZuEa67Wb9kocThwK/LDaWumj0glLjq72M3+6h4E2uwekhbYdJ7n
3W0rpx2q+JFg4ejbtbvVC8rVteainXATHZC7XNvFzoKKortOhmXtcGjPwwr0ojUcqIh/8h6WHd3r
lShi6X+NuiNVFYTvnmBg3Lze4Ec89yeoMjn45ttAdBNjwYPpsjrL2acnHjhwGPy/ySpHtVHibsgg
w0Ve31u9tkWK4N8lIJKiSHsbjfM8RcMUdfcgFqXn+FQwAqtz7uPe4lgHpuckTyLIZ4a0/6d+QgPL
Vvykw+OERD7E1EYgRQ5W/ymzch2nOdmmiBE0OiYU5zsq+kTfn+7dpfByPJnv5q2ELo/J5ova6jFa
V//vXtRmRCKmVXYkK0gZYdATEe2YAoePwxfBYkEM2F5h61mXLW4CER8y0YBnFOFa2B5HGy9MHQ78
2IMBjp47jDigcbG9KaQxSxr5aC0jbRq6FNlrnqsegkYTRgdLD7QRJPQJxgR/xYKVOGeXoXJcy7xO
odc2rhlotp6EP3vV/zKtZEZ5X7wHnK6bJyuH4qmcjpvEUVW1hwIE1WUkK+4HHWHMFv1465bouyej
Jd9FpubJEXVBGpLK7iloq+eVJlHwEBijrfetE53FWLNEVIE/fbZ2r2iy4VdknkhjD5yUT5UUoxB6
+JdglRhV3IBxs3KEGGHTgAegZS5qiZKVUBSIx9M1xFmTfjUPedEF4hDVxkxZ7Gwp/j8YgoRUEW+u
7Areva58kljktkBbYIrT1EFcDXPPbrLyDi5sGBpYasnVM7a0z/nTpa2PMU/74hiwx4JlqsRLFK66
2twf/cu5J59DWlfYzgcRRnbwgCvpNpuzF3OQuXAfMnJuFlh7iRTPGV+gz9uq2UIaBNlvveYcr/YB
nUcZN7Ov7VM5u26TnSl9aNmAzAfpQEyLklNmwboBNz0yASsJ1W7L7ahaMtYaZtlnGODglrfJCl7j
pQWVCLLJT2rawr8yzHBpU+e07ZKKsuHxFqw2rn4v1047UkJ3AXwRjEU3Zo8mLXRXoHtnZKoF4x+f
sxHgjTf0DAYMbFXZlphD8q9X/zpq+bLZI7k2Nfuvc6xP3L4w8Mxxio4qORIgh/btcWJhUVFq40VK
LyPwBbhhtGoshSiri8AGx7klBk4cDNN6Q2X202TkMcVfxPWM2YsTNaayjuERSdDaXhLSu6z+ofKl
k8fWVaP6hbDtiE08nAyvIQJBkuKh5KOc8m4dagGOzlyISeKHB//0qIdH75ha7QMO++NPzY7fPSu5
PFyOlEwyl5ako2aItWupe7t5SVIcfYhjPUArVWldZRbTwtJ/W0BKLitdjDRyRI77TmGTC58ZqTKa
VcJof04uFlmi4Wb7aO+NKL+qAZCyBsz5ikpku3G2HQ6qs5BwdniIPMewTfHeSR681Phau1buKo8p
ZLJvUd2PR/o6hRopRDcqwGrsH47YOxvbkL1TjTnaC6F+MGc6M7ly0jCLqN/im0h7z4xePXje92ir
A2OLzYaaZslw1dnq7xaqWFZ1zPuVX9reAGTdh9LNhrOMO7giX/uPvS/bupImP7dnETUvDmskn1Ru
rmjA+fKi7doYnU0JOEPkQRF927HYi1TCPrK9kyqRqqFyjhNXLyQ4FuyLBuNqDj0fseGG89K/QsPN
4EfeBQcXvxeT7RfKAkXrezHH++OBhGGBuKC3dr4JxH0Ga91b2oMm0MuNzHjDJIoAY6/EA0QyvlIV
oQTV1A2qL6ZCmq8CEeGyO0bMxr0n8SSSyyj0z6WQq5QVsyA4C0QVX/YQpQgrtQH0x9LN2hphnNEL
LVz+ymwVd6DAn1ZAioMEz4uMrIG1F2N/Ubrjww7FeBf+dryC4ABFFS+gcfXDja0g0JigfStODbFN
191A+roJagt3b1kF/BNim+wZovtfmvnAO2dwo89QXnckCbJL+w0qis32fU0qvznZWjjmtYWNfXVs
3PgAGCLSrNizqcVnqFpYob1kLcLNHkLqUmGFdBLOglRC6rr9LFlPEfW8N6wvvm0SdFB4b2WqgMLA
DrhkgGDifWAb40sNH9VO1+HezVG1Itp7/n0TwoWKXX34pkLAAZejCWpZUZ0EgQ1F94DLRXGXFPUE
ayxzmjuO0gG/yjMcJC8MXZI57vTYPJDWkayO10EUPwxy4bvhunQ+CVUi/wsbNuIhqPoLCMhJyFD3
ABptlUiMFGOANVI+imEiuF/lRzDDIv4gU7IVZT4loGpP0H5Ym9wjX+6SXMjuV2VX6giZEJVKu7Gg
KCfpehBU9Wrjrv3UxdoKURh3jXtoFj2Nb6W1LnNR2UITzvlm/05lJeHxV1eTn2NjY0cmilkOKffB
I/sf0dTQzuyx00XOV/SDkFF/FRnhkTZsA3ltZYmsMVxYUuoLYurZkmfU4/gafh4LJFImfU2PX0CR
DT5ElaSQc21RGsnFbg8kxnTWXyABF+SvGQh1fIsZ3MrbxFhm06Q20LfMvKhN6jp1cAYQPERCdbKa
Az6wyr6IgAAzPz8GL8qH9Ooxa7y6wJ/lBMFCE7IV2sLyAhnvuushm6CVJeaCeIeWw4QIcg2wahd2
Pqq+OjyLcJbLA8vbiRAJhzWJiCALUpEKGYZaCHKxYgPN5deYnQAinVCJAnbWpDx5DiaaqvkZZR4j
n22wFPz18jb3qV6lRxPSnLCm1elYHtONNtEVAqXsmOr5eHOq5jxVQ9qUXmAA462dvwob/1LcEPdy
pcpYvNf6Dplw1pQ7MhIbV4BBV+DMq3VrweDancFMXuOIre2BlMrK91cHnsm7w461fOL+AD67wOBs
M1ShXEUTBR9jCdb/eMEill5bICGM90zZJmygdPs0/YaKmriApQlWDUWWvd3EWKHebNShIUv2xfiy
mrMoDbHJkWcgP+UI6VTtCJd8/n1FRbIUQqxM42uR2PDP5m6T2DYLM7GYmTr6uD7WDlmZrvY4rxl7
vimq818iyqvT/GQ57HdHLg8v0LGopoZWY58kM2da2yjYxDxA+8CkBpieSzyZTz7gjirz855+FTki
ynQ62EladYCAClFthVEKKmRI3JZG3wWT9eiptLX0YFGPLccgD3WLhbCllGjhF+BUHbJNd7oMaAWi
9bcz7txwPx41wQJf9IgILmjoFhMl4StQ8h8xCZxyCSENrV+buQW9T6JViyw76B9JZJ3NY4pvdnZ7
c6F1tLZ7hhQrTHgF0DoFAkToXactpFqimRwL2mhcqfCMhxvlTadnuN6rUC5N48jJ2H1G6GRilULq
l5M3H5q71jw122+16/fnxsRiDcoUbR2yR57+DJnLUgn4FD/Dd24oCZsQ4rx7kRGji1w6fFPEEVlC
DIFT2h+BszPkIR4SQlZUhi3bTpBUG3UPiSDFMl8IUjcflMKm/RfjoM6EcFX7xnB8Ka6odIs1vxj2
njqt79E8uiRq6UaSCX31uLBIZisx+vftwsv/exnunoEZOYrqw6QK3tkUaVsU7T/SzKA33tR9Y5De
1TmniZ2z0yDSVON1OV6OE4Y0BOYWsP3yOZp5akqqUIQoxiKgD3D23JesP/fB8hCO1FstvRZU8tCa
UmncO/G4ytCoWGqgJAgtAtcWbXj4xXUFnS5KYKXpPqqfXHceA4BxYOLcxUc5TAYnrHd1KL7f1Auj
M8tmEtgpmgZUJHdgQIKSIZA9gjep57Ex6RmW8/18f8Jf/5qE8rOy5iMkSJ1RTSZMNCFbyPcKe25a
loFdMsecFGm++J7AViMJjkj/C3AMNLCNxZ0P8BKe4/h8Z6mfyMFGyJT4Viz6Sin0FUHAzMOF5yJB
t4FZiG7pQh/gRA4Pqa1eywsAj3N42YKSGkfWAMeWaH9aSNiIulKHN+t/ERTdIcqnR/lASU6dD39R
13bnn/n629OSLaohdYdgys6URHAoZ391UORnpJmV3+a4aWbF5GD69wzjYRxlHZL+7Eu5cqNQHeeg
OLL5FMBBeh6AzlOeVvTFQ9L0BsQ3lKuHMDHU8VDMFJFCMS3xJTVL0tEV2Xjw0gpMx0pKAr1ZqyT4
P+8XQDlYDv6T1BguGXwdFdxYhrr1axUf0b2fI5YaCDGGt8d9ynkPHhd3Idaga+6AyF7mk9rXLSEQ
myMB2mBsZOdjTeCrSJlFZF5z6fARJYYShK1UMM47tibBF4lhlnlw/anLsyJ0vnwp25hH9eRsKr+h
JUHrvVb9vx4TF1MvZBWQrbGTgsD4fufCkSvtnwZSHPByltbP1Owqiko+sLdMvjgF+j2DFhbba5+R
abGy6QNKBIvcMM4m58IcY5xvy8VPGSpDDY7a4DXxUJmiDgZh5B0MDgS8ezoXtDdwQ2BkDoSfTOD7
PfTn0nB9kiZTmpibRFpoo8huQvvhQluZA+V81IHzIhoI9YBCqPBH6uPXjUAj9Xc+14pRrqtCYuv0
7iSUzu/HSaEq4pEJLd6yezahQ2kD3em5GK6Eq0et+sIecwwujH56nCd6wEGwk/xnjXxlM8LZ2ZGK
00iMvzSqWCqvbNcdHITDTldKDf4vyzTl2YfRGuxNLEPqtENQ1mqUIS99FPclEd+rsnF43CdEI18t
LkKEokdJM3LmU2c+NTctIXPUAoHCsiGFQtw/HZd2CDBrDVMtUrqZ/5/3rSHPU5BHpJ1bYkHfJnfa
kjB6sJEFV7OvzTpqgRj+TBiawgmdUw1gbK6kMkgGCURB2xhnhiSS/Xb7hS5sO27d1ttuuVyD9Nhf
07FZPTpLwxRwbIFt41njEg46WrlZxkLu+H0WfVzBknbT+RZLyGBQenRTHnLXrLFIoENvIzw9tgj1
c9Zmx+69fDDUjpLC2defzS0XZg9GI4XllpdXLKI/kRWUS4bDNrmidmbZ4UCln4qQe02WrzkVShZ1
gJXVPbd797mH3lW/+eGb5LJjU3M5v1aIWk/DFCWfRHbMV+5g3QUqm12UqQgB9h0Nwho48+MFJQRN
yczrjqQ+UBj+Y2zmwD2/JO6J/lsPkPumdaFJ2N8mSvkVCRqWq6JxMD0d/mqTg5M3LEXCcfSt0LB2
ONldmIm4oEbBJS2YtTLF0EEcRdGWdg0jTeQ0GxeMIxkBKJ2lhwkasE2jg7xDMQZpKlYFLkA0IPkt
wp17ul+0QD4NTYfmp9CWFtZCHopBW+FamgosU+GMm4beJ0iO6j/wRxlHvZO742ngzSuPiSDJq6Dx
bbrb9ATfu97mmruc8fTxaKznK8j4Gm7+JM9XOxK9iYqnwF/q48lNxXnwoJrhnOSdbTsiJDvuaVnr
NrQ04WwC3IT6FjQ5EcNcCMi2cmmQjSBTg7qeH67qthsY14Om9N+/P+LF+o2oVRcKB8jnrJ8ginSv
kJKBKwZPphHOtr7ZEx62EGoUYSuenJLDC8YjY0+hN/W+l3msNYy2K8fbFytYeaNlvF36WvC/Ryn0
vmS2mgN3nOfna5EnQrjacx0hkdxIUnw/gagk2Rsu8hI0aY7vL7f1qqL06XgTYOO837yI4UjKjAK7
e/tZVE2nygAukK31I08s3iG3kcBDzlB7eQOP4oyC3Mrl2IcfZDbM6UCZHRk4xU7tPAfRMKGaBtJj
97GhrKO9XvIUG7V82+TaP4c+/s/sRPJahJMYBL29rF13bnuCzVRSbqLzlXNlBErZhjC7vJtTd+cW
a0YaqQA/hrP9pljO1q7SXBLmWEcxn0hzLV+EzJEcJuyv7AmlL5xB8FunF7fVPWu6e1YZGvoeYLCL
n+wtfMjqAsQpEdJzFlhF7iNrq+wkZpQ60VQd/RpF5/xfNoQDiGjvR02+72ILYSFYS7USh5whCALc
Aqu3kQwYfR0T6RunmI/Deesg2BZgbHjzGfZxmZE7Tkeq1BHrYay27Mrp74k9jQ7bOfDoLep8HW30
U+Iv+PsxXDMeT7Cj4zW8jx2qFrHVtwx6CjShF1SZ+OaN3gqaXJWLhDvTn97nUkRlezAxtUQ/vNJA
GDhF+SoopIt3KXqn7yYcjeWOkQGNP/BHGIKKRw0CRxK36QP7qenFLXYW9QplmD5Ez4Rt8+7dq/wg
VTh1zDNhT+vWvxmgmQqIHzzAGWCWhXrO2HV0EqGVVyh3ipNSZ+aU/1CXHLx9AIbfvKHFxU0kRXTK
MgLQB4xdwOpN8+MY9iL0NBxMkyNHE6xw+ynSE8+5LeLA0kter8kKn5nAvvcpb+aBX3jYOpIpAd2p
C4TKp2r65kIYgOK8dbWzpsesfGU9xU6ZpatjFOziRzLHXPPr8gWC6QSnQtgxoSHmjbnDtu78FBsl
k+gNCc1eDhsEzMY6gr5NQjSDTHiYgKfNb8/m7foaDELmz7yGUt0htI//n/NkUzS20uQTgroFANcX
h0+TdnnaCIw8OQUd2JboGZOG7IH6zjaVM152GlB4hRng+IGm0lF6wgk+19QaXRnUeKoJXU1/JjFS
5pBeGOKxG9wCR763w2+2q8nwi1mmmxNsAGuqz4IsYMxHfpWDgindVQyiLu/j7ihprwSzhNFkPdKt
PfCE9toRZoLlOgxWCyYdPcL3r2D8z7usR5j8zJvhAg9ljEOGLbQA7ApdOzGvna8Zlk7tcjOTSKB0
6JNibRYCl4JTiWhPv0t5r00Jh5zymdRzfDL1OdhEG5XBIEcfcHBZgb6zSvd4ZyEcII5R5fxKdlMH
vmcmdv0o56031lJ0bwWIqbqNpgypBDzG2VwrDkluMc+lbzJ4ju4CLWFMbhHzG4BBWrnpXdXsOCUD
sX1LGfGVfypKPWCJGvHdXx4GUU/HlNxyckkoZHZJJ2rvclujgqhZ9/r/E+j4EfgcBsMxjF4lZ9jf
P6tUkf4KP2sUhbgYQP7Q0YXJAa38266+G0wjkdxpdFAN/bOEXfXunYXephauT+9ChwrJQMU/ZIjJ
++M/l5mcwvsWKxpSBf71+5OYu9vEAwZKUIDmYxEEwamW5AA5rnCfcRqADabvkQg8je9yAMwpZ1xl
VrG7kW/8AxNnFXtb5dN936zwu8FJH2BT0lXUjLooDz/9LhhZ+QFLZ5cCfu8VmSyLxT2h0aU96G8D
1W6/9MvBV9HAsikSeLPNLP1/y2bMp0mr05QtavNqiazAYv3WT8FCaAlQQHDalBlRz9ohXsvX2xYz
ANFgBlqa2lRURlF7knrbxLB3Ou32ymqtomdW2pnKRQD0mQi2BD5Lv9P2fQsAcqgejYNDRe0VASmh
6ITpOZiQzY9z0ruGY3JWyoQzsgn7S+UMSqh4j/VdWcw8lsz9z/w8+mqIxStXtP/O05BGbPjZEtRQ
E95tAf9Tf6blK71IoRJhmGGEkJFBOOdHq6SXlj7BZ1s0xJrvPVLTprqcGRLr72RAMoktsFIKXUlb
UkFljjEDMne7i5UorIsdMDFX2AuTWedrExT8G0QTDl/9+U15742ekU+Vkzjdl3j5e/QF+ho6dYux
tt+T2qS5im9LmnKlnhVgQTvnLq5voPpz2z6M28Z7bHhAlr5bLicUJev5qk0WJ6gLRAB8kUa4ajGP
wP0T/PypqudhnK2lwSaj5buZHuwMVHFpwn22aB8jaqsB4j0YSaEmmRI/ZjEdFA2sLxvWOmFnD0s9
qZzJrfnYKBQytHJyNzkItHmiCNs7UpvfF4Bobs1xvZ4j6N27wWcUm6aczvv40K/CvPfnMThjS/9V
vQlN8N9BvTNzbn0PXwFjY6ybbqpYLEQ7/HTnFj6UvJ0ClTWw764YxGTkBzhRATKJfCdX7aAHYhPm
8vE4aU1/Z8DuN8LbXAYfafgFbl7h5+2Fv+H5LKP4qah/gvYdr3VqF7Xn9o/UNCKH6UAlZaLyiOAn
9YY6PH8AGhwduH82nGjBesE8qCOuwORAk8anwqGvl9Hh4+NYB2HEsIDcunhL9+aWoGRBO8fW8caW
rVwQWbBdosKx4Ud4gapp1um/UnLot3vKkUut35vNvHl+g3AI+EGbr4jENuzFOKEw42/KKIsG6uA7
301hL6jurPhagzuLYmHeA4TLUw09qtr/IXe2I/ay7ZCl1fBbrIpajGFriIkPt5yf0ZRqApFqGPYy
9Upt0tfBTaSJcUwk6nfdwDn/RrBLEPqWwVKthIwt6fv7aAQq1hRMy6Y0OwFXJICE5foCxHeWRgxq
XIPkXZORWsx0+Tsa/QuMbI5VA7ziQ0oben9RZN/Wut79hVzS/jTRtIaoJVx/ANKIo8v2ybpDhxa2
QhkGaPh8gfWnyFHCgFMFj35uTFRzgWdKtkO4gE3LdcfYlWQS2qNzg0ATX2gTSyzf80P38hCkmfQV
jtW2Tgop4p9AwXL1jFhKt/qgTIsRt0D2cHVmk3fXpWWPhVma2GAO2aplBYNUDIs6ZD/SqNr2Ua42
rFdXERQGhfhEi1lOcWXgXImMO3/kU7c9F9+MeMlvMRgNkWDAZiQ9V/tnx5oXDYZlo1AXqGZyNjbh
P5QaOefdkZ08FZTVDHhMD6D2GyjpA1BMFuP3arztXw6aE+nihZKxuJuniKaxu2n7plo42XscnSa7
fM4H6GDOrQWihR99jj1P4bwAFcSwJu0YWMh/JyPadaUk57KazADySWHmKjl/B8CjjGjcx1ar2kDp
OGaanhnOua/tpCCRSgLIHC/cbEu/1XDKEs/TCmpVRbPq3gnt5dOuE3W4//bpMApG/HguYDMABK1k
i0cgIQWpLrVmVHXohl4GLYpsfaS9zgHUAcU0lg8tC7+AgB1k5eBfPV+qfw7excpwfoLWPimFTen6
dm1iIB6XbhKn5Ujo4K1BVH+Gwo80zAPA3JuQ5hpkYY4TQF4xKh7JTQcKrVI7ruPzSJeGcpY5p+Pg
Pv6DS74cUzXzf6nJ+IYjFiVzb54ZysR1S+sJr8dzw9ol4JIr/6lgEdSYOqJgSQ20J2ukIDVw35oF
RYl82ahO+9VmG2rhYr2SO/thsRTgmGkeSgxIVjX+9i4Y26emtDP9L7FKIL8k+GfQbvQ9KKoBPTzK
hIqM/FDDqBDcb2XiCD+aI8WV/WI4gA0diHtADmEwN6f5b3Bqmzot3PrfEsMUsaM7Hb61kNuM/Kax
tp49E+pTGcjAAqmLJy5k81LD2bMihwi9xVH42iBh1Bz1etkgLhVtJJumF+HJSmE4gPrWNxLym0O3
Q1LMPhCPJrektxj5Q5EtoNINeHwuJNWEJa1iVhg2ereWn+oCrkprA3NiPpPMZ8u44/HejwVHaF2v
Wl8RpM24udLgUmLSuVBbJrrmuFyKytmqiThyNJzXP1csEOroRHLtgLo77xj5akq3G9qALzzMyWDs
QQ0TM2Vb68vcaqM5QYfF4/ZRA8ajzSRrcDlNXk3gtw5vUlgXaS8d4BTr+oAUU/siJDbPt0ceqQbn
Y+rEHC9wKF1+cDKxWA9pfgGURlNWYQlEhHqTj8Fb9t2UEjGahq+OrO+5zbEpXKArBeCEJdLzWN5K
c/V4Be1j9RIBHeAooGH4dy/4yVzHZ1fyTd/G0zgL8suzedfIZDUgDTBOdtudO1B0+bKyjTIN/YCP
BAF7lzG+XwY2A4nEuwbjkTPif+oZGjV/FvUdNynEp9/WEMR86LeAZrNt/coig1LdTkBEPTuzoeGk
syjjKAXVLzW522k7DRP5HD9MRIQi9V2GR1GRy8uqIePfFuKEiLcpidcCFfMpVxB/Tcfx2ukuUxk9
jmxRxleHGE+ljRyJgk9fJlSahUm+TmPNWyS8cNDF/aDpReXWgWYK3PdlRJOqed3BLJ2tqNsgOK2D
uXmnrgZqBajbNGwV/vi76qU8uYc19JWvQmiUtMSCUS5Pvc45521SdRci/PZYF6at/k3snU2LD7P+
2FxUnUuol3K7V5ZDs0F8wsMzCuP1rULX1vPafDPdYYxGHiyaWPSK9BOnSLzHXMBVM6qI/x3f5cUf
l6AVjHzEetlOfFPbejD0JpV/8myx7XfmrTPLQH0Pdk8QG9JCatjrPs9Q1Dc1KuOEOaiCZYsi/wiR
ptcq165ktm77/ePkMHeQpWtTrWjcmIMT+nDSO+dX5LXfA+eFaFY+gPLBvKSoOn2LY1FxHhBc/pFe
8ZILPjc74x3fUj+DB4Mshx8wBRCihT41tw8vQ6OGyAbRU4ZH6FBs3/e3INVHsPVEm6r+vpY4L/1+
ZjXraNG7jJyTc4IGDMNoMty0xd1lTSKBc7wLEzP+k8ccF7GIab1JTy0riUclWJkORrzkYWBYVC2/
9P/3yVh0uyDgTAF6RIiqSkMciW1HdgtMzpD23p57KgDK3UwjrydHOFdtCvhCSPEBTsy6iKdLxdOb
zR4qAhjgZ2ba2krfQwtJX2NX6WgX7IwJs4+CLKPlauWcyoN9i1EBigCNWZm4vbKITd/w1E6kM+MS
bG5XLlPSqzaCrF/HPHFDrSWHA1jAMqVAeti6gi7mpg+Daf5eSAWMhxlpInX/NwuWeXZfR89cJuDk
pSpZkL+hTv3v5lXkuxhYlCfOf4NuC8V+xp37fFCK4XJyqczgr8OdFNCNnEMd0OGY8nhc+p/j69tZ
t8C9xGqeIg7t698GJ8sm5cqBYARH84TYIW7SqvUCsB5pKgLw8BvHeGHfv/TLuJ/kd1dF59kPb3N+
jnzhlaRgFHmkdqzTeGyR4XVaHCgR2W4jSL1metznOv9eZ01KWpgkcl4o9Q0cDDjD5Q2pwWYRq0wT
Bv2Abc5W6E2951k7gHnoUZ8uAsJdFmUxiZ022rnnvzlL+4IcTn3QmQD7vwiGCh6HTLCL7FXLqQpk
imBeum71yjEd24obPDDxyHNjbW04BGHZfToKP//tG4EnC5HXn9k/C1h9NPXh5SknPPoFrarKyLaV
Z+CTr2OeG7ZL14GBat4ScXvwyAzW6a8BdB/uGTRE/bk8U7ctPBZFvFpbPmBlrVtqNXVFVJdViyyv
VddgyBAwRkecO3/enFcO9KKFuzNUWbZox84EB3vKPR8Vr98YYQu0Y8Mohaln58cO21Df00bRb6mu
XFXaOyTSFqHxYNhqOSc7LCA8pjGC9t5qk42xPZCO6hV2eKpZcBDTcvScKjqwfnXvxibgsbXPsqZ+
gKUk6razMAxANZjsfsbgd7IaE2H2jigrHyeeup3wSykb9COKkXaRa2dyi0vtRaIMmV1QzJA7haoD
LCk3e85ceeakDyPDNrW4rLtQSaXX+mSJ9+woxH+TmHekJadCEWOxsMWbky6NeTdfIOfyHIoPetK6
FdflcVSHeYndD9up1FQCYOVi+ks4R97WWk7gbTB5Tg2Vh3d/TkPRXmmpmHMQI+VrW8/egqLESKzr
nnki3wCXtxLjVU/7srT5Q2efupCp396YoKnX3APwa5f8fqZKK3rHtnJVAg4i98UL/8K7M/0thZOr
7fdAWTFxViHLP4km0ll/IUM2s1AEdWt7bvLNyUdPzNBRlxmrLBAQk63nqOIkG9qDhJopB5iJpm8j
u2RHAurJWNTF+M8DdsOIrufKKQ1XJZWQTXsBGiduDw7yn3su6Vaoh0/QulK1vh8nPo6Xj8ttiltr
ESn6mOV0FhYUoUZun5iaWBx3X+P1+0tllPjcqZyo/Psh4KLEQN/6+0dONJeklbsDt9egWAzi3FDS
NQPEUq96pATNYUIMQZ23BtSS6WASR6FTuRc+bErVWr9DtQEYal3fOetHDj4WePmyz/5d18/JmsJ0
MTViMIuAyY/7cGE3XcpJX76Nx1ZxuFopwh7ODtKj9EYgXsrgp8AqHGRwHdpFAEaFDU9MXa4sDm1x
mPtQhFOngu6yriFjCMUjSFzO4UgwVEWsLWDDkBrf39nBsbaJiUG8azfsWeIRhSbroMPADr55q69E
toRHzjDstGvXKZ1n4MXt2ifewNP8F7XTJmFWccF4VYInww/3gJRun8sWms26p8mLRrlosSy1/Oww
5suIoXATVMU0trMzHPPPGpXEwsvXYqBsc68zRgICQxd8p6yIKzGgLBQk+qPVAro2hR49iRRLrgrm
DeE0DRiUn2QbYFqOlmDkP0S6+eCgJfk31tvE2QKCeWDJTdTo2rTQqslNJeIM6GvlBHK2vWmWNypl
dZtrU20RR3nLA0AXp/kqxbNX15X59f2DEBPpQb0ADGk0bYym0Gio4YlSWKw78plETAxO72B1ROMy
AHw/FCwhCjdy0j6f09li04rHGr3WUIQZN2A9ERn2KAvSgr9Pi935cAuQVRhdFc3Uky5XN0vGUKc5
yFX6cGYPwYAJd87NtoLaVcYqlLSiXvoRW9mTl1N6EUJScbX1i9Hmzut1+wSD1BwBRYJyr9wAcsRS
5lKrfyhM0+/mjevHc1DfJv2Md/20TukZpJIFgNJCH5pmUVyjMxukQdjemoikaEx9BKNvpAOv1bEJ
/SX+c+24dSHLeYU/at4Bi+zPL56QIsDxOV+F5etY995vGaopPvatfznk6C3YiWUBk2cMfiLgSxfp
O4WP6YR/mFphOGSo2qmJZnSXHRc0OEL/KuWXSKfrXS7tdjulX/T52eklS9cA6z9Jno2xE+8X7pM2
MSFrJ7xedXnQzoCpTcN4WK4btJw5RDOEwyCWBmZ6GdKN4ngnymiQWT4UlLJwh/bZCAVZxBBGIdG6
d5vDWkUo8i2wGHa3J5eDYi7RwXdu/u9fUquYPSdKkj+J2czPhcfSECmKrD9ga7KnB2bABveeogke
0/lRtWe+Cflq6zo0TJlGAURQeA+0dfWVCBri1v7CiAEtZQTE/aq1IuToGh7iFtT7d4p5bPvxqYW1
zvU0Rt2KImY4scRyNK/W4s9yRj5BFEp7iYRh5TWouEp10em9nCBOaO1KTpU2wbqEDUZ6yFJvEpQV
BLolnWXYV7iWovxPJnPMWgq2PfzMJOIVc5R4E8DTs7Zz7K+MS/REPvdS43mhXOkuJ2ePoxqUQj6f
rqhmEVFvzlP+9bVdpu9syE9Qt/a0PG4j6YSGHLHHbvwwn6ZUhIZ5v3ZegB6shK4eL/GgrQjikwRZ
XCWW2cFElxZAN/janmv9cpLmBjlPqsXf/1MZx2ODnplHLpiPu4eNjAcxRAykSHFzEraA7fLvbPdG
Ui+pVUy5LdbN7D0dmaWeM84Ly08EmaXwppEZYFWvI4dJjQCkRu93mx1UQW3wivIPdbZjqrAHqzik
8fZd4oomYlRquMcnVX9SztrxD1d7TBd6bgBvPoohlFovZcQ0pFO7LtMDr6VoXfV9AW2IBqvXBLqa
c6dX3zjPuFbIlo6Hh6PA6IUFwtCmA4W1P9jLX+RaOstHEIXEia7yxiZAJooSITDDXGe3vutF/Qdf
UWFNRMPatKFdihARfga9dvOoLzM65zYI4iJSh4+fnTN3+qXNVEVsj6o9q+8XxeI9pEJlx0cOvxmQ
YoneodUraqYAqUmBlGVVWdhrwQBM4MHNtCe4Y7F5PlqInGaqXLrBxPuTQrRwz/2J+z/AS7Xt2OUO
cFbnj5tSu/aL6Wt/oG3YPiK2OjZqDHutA6QweOt1X1cw1L69vLvbR8vbktEZmvZuGxUZqK2TrOIk
T4dg+IN2ywmDKurK/CmLpwg3yp4k9plRyGYBLv42vRyrzfspEoJm1+3hcJ0xyf8nIjjrzcsc2u2S
7ySbFg8CXnrKsBqP8cy9jpC5Evxij13CifI6pK3aNrxw9zFMKnm4xE8G/fyMz6YFk2lt0w7l/qAI
4bT0zwr3Wkgpcc4gJpFg/seUiFlSUFMhMIoZXdIyD2+NsPLNXNWetQNRLVyxEllE+2g7/Ff7BmWy
lc4Dku73sx502Pw/vh0SJVgfc3TQjmmW7mrRU5r3iMhN09jHeVgh+BXmBgdbHnazGm0yyK7toiRw
YXRw5SbYsQfFan7dHsxhUPD9MtoY53FXqpjggioV8u7mDehJX7uyzsZMXSMdd1JPx0RInw6cFbhY
HPpgOiCQy8LKc116KCcHGVLAR05cAxy7aOqO9r4mHwn7U50fLAtZBW2m9UEJbKuuf4EIwtvmHSGI
/5Qgol3WDbEDnSGRwU8L7NGAi6PGYBg8FepnKHBZpsDVuUeLc8/2GtaXdPFE4Ks8MZsP8qrx5cnU
QRKxKNF154n2F+7AoRvRY6WdEHemU0WxITaaE0WOOP+IsjQWkWXJNGEN3MNweAe18yv7/sjtq87O
SJDF90kLmwDF0hrHX0lwUh434LS8b83+IwYJabWuSaKBuTp9pjVbWEnnCHumgThKZYTx0oscxdjf
WjNFmwl48TvRTVsQ2AU4YtltY1oBwr/Zx1tzXMRHyldKpGzGPN0x6pAwi1+qh/4VEnRX8rCVqLnS
kDUy5YUjLAcY4uswnruAgJ2ltlHIJSyBJzuTX/TfyuCgcGi8mEAPNt3in5IgQ6CpUseeJtPM4btI
jlqGfJiltD2G/ifQ+yBKTz3tlsrRSfx1RhXTls9atNlBIgM87eZPhbvtcgq5zhZdoNiBhCuoNccG
tZ4x8wCdChTpV2gRxufaGbH8MSnlcOif3IFSzER4wWw/g0rsU8H62Zje35ktExJfUGfxjC4AjBix
b+Ew2RnAL+Iy7F51tX6gkHkJxW+5z8+TbIAp1o9rScBmzAC7lEN6dco/f3C6Q17DvSkpjPLXFFSC
dt5UrTIyZI02rMKPG4zYKSTPPKMcKnMIE8Ewr7Tzbv6WLiqiEkheUszpbH7gIYjr6Am4fQlMxHLI
TIM1Og6BDnPjw8m4DisgiPFCoJemqYpMDZNwjPb3Q0wv3acf7M6SWFqLkVRXbOSCrduQgfJclf58
6c1RLFciofj9+n+OrkrBwNJnCEETusf5pJYt0JPqkmSgNKq/hqV8b6f7vytfqgmlWD4o/ksS0MeF
WwJJc7hPH6RlfyRIZWh8MWL+rXyLTA6quyGVlCHW1z284H4zcaTijdcDe7Q1Xeg3To+KQKxFXObs
ExVoVgDgaCNEMDyhleWUlxvij6thMZvU8JzTyqTzw/N3vk6ryzWusgMw31xwEm1Pp+LTDY4JM69f
Sm0WsMAqHMGfnDTL40XNbUw5rKNAqTpZYAYzPNyNtGCA6rH4gc87iE0NcZ4OTcYUo9uWNjJDsz08
aBLRCdxDibRbsnGl8eqCs7ZQlX94G5bAMSIqFriX9WJOzHCG2jgMqJ5g8H8UwiaDmA+0kH0qZuhp
tI8canwQ3QneEZqJnFSE9QQ/ahCaq/a4aZ+x1LRsHpQIeZFDPkp2c8ljVPc82VfZcW0XzQwnsZIQ
ZFK+OgdvW52ZqV2cUanqzeZksJicz347wDJP8unsQqzBdzaDWvD1D0LdGM9oLGTds16OqNyI77z5
AnbG9jJ+6Mj5btsUb7eEokzow2DDH1Az0TMldc9LflI+A2JfayQbTrE8Xt0IQjNwCFkwsCvamQe5
meReR0X2ZQXwlTKcgwMijNBSh/61DyeGxnaMJTnnkQuwZ9n9iPgbRawAs56lSRNxPTSQzLIidJJA
k3Xc0ZsVtN7ngMPpM+/6ao7UAQqF0dab33gzfvIHvDa6adfQYmf+90dkGqdZ6c+S/u1Cl2jTAwmg
h+gIB3pUhfvy874Ilf9FbXVdHUgCepVqOYLvw3MGqkBKE20gCpZ4NEzayvlRDfLYs4d+Jlbme93f
m5Yelz1G+9n4SgsEl7izOohh2sQlEtWpYXZ0s2L3Knsg2Nk/H47ow2Z+V2DMV+QwMK7p/+zfoqei
hU30odetMMThzZ02Q3hv5JPa2eQO6wwuEkOJHK9ai+nB5U8P+JECHmRFyF6ukqRAk6n8OY56a54p
G/I3V/+XMVugNbSAeoK9pWBbL9CkThShGdLo/s+3IbZp1JurByOWtQ+ZQORYq+tPh4xdBZoRS8WR
Fti+vKtv6UJ5+a+hurlVNU8r8bJUUBjquUGSsbfQ0wsmfvak/WWuByN1guJGLpEih8MXBPUfXrbO
uGPgoTVRquxDws5rJZ6PqE7DITXHcl/Lez791aqV+7UTwe04UE4FeEeg72pXKnrDF47aYhYmIlUD
LKszXQKmz/jmmpHGsaY1z0n5onZsM7XKveQ1/ekSMmecviWtOUS2cwIx/FWhTagsJipyEC0DLNUu
7NTB2zAnT9k9t/wVl/V+vCmjIa0QQail34hJ3se+eZL70pK4svuMoFGjmXJA/jYUsZYziL9l2wBC
DF0vp/38uST/dXRaQSamm3k581uaoys9w0kvgKGOWjF5PNnVONGq6wLx4XP9gmwnpcoM/Ig8XoAp
wML1u809cAonMhOCTJZs/vQN4MFw/+O67bO3c0tcrH3bQBGA7Y9wEaWzlflv4QyuZnt/sS67sN42
zDqfEUG9myRmkm47BPkutTVsppzPoyJp7GtSujC5lMieWdIy3ohsgjlUOSVqHoL8NUg07sxSO2B4
Psj+NXzaC/O8n06RR0AHHKT5DO3mnWaHZIDBixQfFJ+AK2A7PtQ2vPqmZyzkNgA+ZljAQB/MSV2O
dnDKop/Nr5I1PXDWNc//Mtma6WH9SquhwOk77ZItCZ3XRc6CwpcpXJ3K+Ko7a2Spz/1ruTE4WYrh
unMF31N22F9p3ttToWX1/J099v8HIrRQJpotX4Dk/brzaGk4N23LrzAk4pgXO1mReDD0sx1na2Wy
9vG7Y5/w4tzXZPv37e4H9tc1jUICX4IjilYl+GmzSW2N0pAfWtodp+uYFFaF5GjlZXyOCR40Jw7C
zEpAss5vx0NekGtAL0WGvzOozk8AZx+pFyANoWIX4hzWWIpVFLZf1RigStitU2nCfStjoFVPj/lm
1AEr5U4QeuKtak5LL9ttjr/ok6YpO/aKD4ulvrDQ1tE9wvkDUdfFnUkyfSqvRY0Gxo78CMUNbHrG
5JqOTuWMrjX1CSdcGe+6n4zbAhCZfSfBhkxluNiCUvLvXSvd/OG6N3uyGcBEv+3TKcx9ko8jvq9C
9s3f4EKhEvjns7l3W2j4YEoht5o1pPOv1dRghAKhss/x8zrg9GciShVp/vlWVKuyR7IVimYoSoGN
BKKJfkeV47CO6kykuePFbTs1/7uRWeWeaqI8kEJ+ECoi2i2GGqeQWxA94kaCHjVbNzXgWq6UTMvC
+DzlwOYFWN4LBRvFSe263f7aLMPpOOdGVzfZcaRXhZAqcSGDj118LfXLUiPhdESh3rafT8CBzyh7
EfmXIdpOjNqjY0y3Rv5KeZ/fIiRYZavgiP0ilZGqIiMphrcsA77NaaWC9lbpIc/1B3iovrAttb1M
K5F2yNpbc4pgHIvOc7nMNv9Al15yXS4DQOl+454dJRjCX9853+vvFqpkTAYF/2mHFlkKU0mADFvg
Y1PngTtwarfMTKo+LXsRwG708NQ374aOubatxeBGlQyuSW3Hw4oUtuizBXXQEdwvhAEf2zdTVS56
7CzelE+6ksds6nsDtvlLzeFnXXRZO1QnJ85kKx7fRGkdhy857LCYhN0rDpEK3dUL1BndfkRYFp3H
WnBv/IY+ocB4tGuwpcmCFnjRmnQStP9jYYA+8VgFtzl+XMGfeItz12GjbyoCEJJ28Q78adxmveOJ
kCQUlt/hsDOIUQHVQxzU9DX//lRLH4LMjQc4FUwAkcXvatO8VrX4iYdUSaEW0tDMUSgRWqwGAmx1
hdEjg4gOUbiyTH8PmjDVy/KnvcksyKRo7Jf0VxZs8AN5cZFLNgAYuQBo9Mb0ZUL528DJNvi4peI2
o1y1WlG3qjmiGsCZfO93ziijOUGoMbZjKzIpL3O2h7F3PdnT24Ap9ZeHcUoIMMbDlAQI2UMT9Wdh
eMdi7kSVcRsRDBprhjCqQSDHPSxjnKk0XQ/cjc1MEpMfbPNU0y76tw6FYfOsLx/VLn3IthKMLoVP
aU6hQw3v+x+i+qtqTJ0TEdSMfi87jNx0RBGgo6v78VZ7F63aJQD0ZWTAiBd6RagKviRA69Bt3o6g
GQMuyvlwqdJCyhQbzg9/Fde6OVs+rAFE84xBMQ/sj92SojfJbA6O6F4sD+zZS8Qm+aYNVKiG8c6i
GslxC3IBH8uX+ACbY1vYFgoySMCR8ZXm0d4jzC/NJWydKagrzZsPUBKOfsynUPQ24DECp1xKoj2h
mCOvjdOn2BG7QzvZTkVqTkRFJS16UqUW0s0NMowAV31mlIbGf1m0TePIL/JmNcq6j1JYz7beP6Zs
4hwaqXJHNxYi8AXiO8CNVK+K4A6/TVKY7MgdOqq9JQhvr4Aip9EOm4mcvPIeGGT9CTKkQWKZyjVo
lu86xA0hpE1ZMHIsXnJ/8Jj8moECncN1322acWaBayqICTWAD6EAW+YBsa/RIecsaMDcBb+EfXzk
8r/nmXtfUoB0aUqSrqfPG+PApGPyMJP6gc9wWa2odfdUFzFVBPVeyGIbra+nXE0IzKwaLfg+BQiC
i7rB6UVoQ5yompeLD6QeCTQMWiUeck63O11TFqPzkR4frrO+52Rg199pjQG7aXf0f/PP6ZiglS8+
a4TX6h2m31cUfsELHTYMYiPdWQwUIH5AoXeNZbzyQ9s1yfh+2sI0bIqvzhXusH04V1GX0qsaqV/+
GzDR0Rz2uFzTEISgYBdN5y38fgyYUgyuJRGbBIFl93R/X5DWWPauMgsQXUKqAPdYGnSmLdsq+mtb
U5EthgM42aDTZsAIDTqppLBqj8teUOyDeOSyn8QplFDw9E6M5lHSgrivDgAgAop59sLxPjLEtWdm
3Vaw+HXaxOUwNr5Ra8BHa6+lS/07/b9iPveQtzaBHUwfCoiLEv0aB1Qt7NVHe7Ke0kXAojO7gCJx
wZjVQQ1I9PeNciZac4P0kOjl40A+8/X2z72tgLJt4Y2Ilvb9zX2L09NuknalPS2S98JXbRGMDbZ2
kZadU8jOau38Dq0Xx2aqSLzc9ZmaP485lJ1Ktxic8u0NrY7LizSpHB6zpHZcmrAeReXkeU1csWSo
RBOGZADd6Pd5tN1b5NL71Fo9yFe9YRFptMrsfSoPC197dCQKIVDqaCYI0ASS2G4/3jCF0ST9cnRH
/vmdaBSMOrj8xGr8cOASBVw030f59w==
`protect end_protected
