`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
HHXt3hRxl09lVdg1T7gySnfuKR9LXVJERwsMgHyfYd09G5KVIx3zFKvVfw2G9iY24SzuyalDpJUS
hG71KZgdc5Fa3lzqsmxTw8I+ebjKVNotySJe6sjeqUvYldaMAwIHbrEGtdYjAedVVfA0Eucs6Bmd
eibAM+XrKV7+scDi70lKH2MuXxFTkWF8EaKxPir3f2dbZ8GUBNKNI/xaBhf2zJtqCxc5PLYnLaX8
f6wnqb3c+88hvDNClXCCwX4hMP92cNATkGHAbue8EuI/i9Qy+I0T5F14vUF0kobYey8rtoUmIgSq
XI879wShlG84/b+sUPk3+RxbOCqSjDKJJHpRFeyn9VxZmnFjmDQJflKAxGmTTFUwzRNmVhzWg0TL
MLbaEBP6cbycfRGROdyov/18PO5ZlcEw0ghY+KxLa1f/eocvowkcS+nunDNTKSqCvEz80zUkDY8G
OPvGaj6nB8XowJfzwSLZd9P70iNjS+k64Vwq5KxqMSZn3ESThpHIisFxLfvdJAT59ydCTHUIo+If
wFws8dGY0nBtbmSRemeEpm2cKu1WU5eiV65CvcPLI0HBoSi/FYFu0aPJX2SvBsW8Lw+cdC11rg4R
cyL+dY4GNDaKHYhdJEKEjoD6CKjqi5cuABeGyULTS6bMPlapXumwuBBy6CxI46pDOoKub2cjUden
QftLAPuyUBFWtA8b5Bd+q9hyJQzK5MZLtBYFqg1a1i/FlmZBvtT811G4WyJv6uRYLGPXWKWyfZTi
Nx4uK5tH8yQROvUky6WUA2PfqHogwNqnq5ak0A60Etk34ezpyhBw2pDhXYR+XvrBHAEmv815+ofy
6z2auzpebgZrLeGAu2w+E7mUt+Vwcijc/CbVcrIzxWJYRz5zyeVcXGG3ns8LxRi8Rfl+B5iYlOMR
JBfV8+zMACL8M4KzBlALw2PTw8SpMry+fA4ppXDnAA99UN2ydimdqWcyAD147ycHpeluJSqpee+s
qv/9iCRFAVm/47lUXyjAArv8s+bLbToM1k59Mn3xwDKQ6hiC1E99zVg9nZy5iYZ4yhJ9SzJt79fP
+3EzANbdvdcJEFnMLiHjhSCtu9pTadX0VomKaQIkPozCF2TZ0gTSTAticKrYwY+yHuGNGwpb54bu
n+EdRIipP0PwAv4f5dSq+LlMCZG1K7xYdbjqeCQbjC6MEMD18jdcAfvl/kHPafTMhqEhpJOYhrxF
ScqLgqEmk0FwNf8o9B2WT+zIWzXNY/y806jmQQxQy8QnopLnwWtXMGc6vjVvJxesxZJJxaCB1pPu
a/wo4OeI70IMWwj5CnZHu05MVgkDbilcyBom/Dc3PXnWlvXEmR1PK9lzP/tw1akMmlv488dNPQgs
CZSRskmVdZsqHY4BZRz2M536+TWQ4StVU65X69GEL4y/4hTfi+1l3l83jKIcaxaVkZdZxlIZrL8b
wOqFlopQ956stxsua7aeZBbw348FKblzZnxJIsE5UI8m4EVEGKb16geM6tSsZhnoqa2DyG+iXu6J
nDo0ciEAYAa/qfQkiz938FMdKIyDrQUK7EGD5m4x0D6b9m8ARU0w9OgjSNgjkMalUyoFgav7Nwz5
xifyXwemWvIdWFW5a6+MEwkQ7x2YJ11d6gB/vEDgy7dsiPb4gpPfZ3MeLhLCRf5UN+j+Jf0YntQE
zjzSypdvmvZZX2tThr30fi6ObOc6CtK+CNCNE5eHy5uaeNq44ekgRCNx7d6ekfWG7T6Wrg85P/Ow
aWKdKQlPGALOBfAqaSFq4fz6hAcDMsupG2AZylx+FbgCaIpHoR9JBjRKr529FrN4Fm/zhogo/Tai
mut5WUypfPHbwrkMk33/Z/84CzgAi/wvja42kIVN7vH3I2NBxvXi1WGbNEP0nRsT89u76bs63ys3
j2/Lr9QHHxYbMMsiI8BiwMecJHeqigS8qtaaE3rF1u6whvLoPXWN59VUSY5dhVtwTWmYOisooLDe
hJln6po6aPdOPZefuKz9XrH9noc44z9MUeLxBx/v+WY21EnKvyCc04wH1a12QnuikLf5maXdOg7d
Zg/OPtsykspLTpqWGRcX5jCkFRNZ+tuMGF3VpPYFLWsAHFcFjHRA7sb6i2BpUtrnK4HSkNcM+acq
JLzX1HIgh3X+SU/GB2GRoqZcEstXC6E80jz2VnKtd7SG0IAtILZsZ1EraI+X0f0+ZCHPBLPOTq7l
AJXxNs14jXOStgRHqgiod5AfLwe5jmKWokEL/3jBV0t8b2csplJvtu89mOYeexhwjl2XBaXU87s3
kH8nCNwSzZgINY6+atDNy+ZM1BJt3egG6/dt2HLg/C2pNczxrJeV3/IEkk1oIyeNYPAldFxayM5k
01+vV7X2j4pWhkZmoQvh3JuUzeQKhgA986/xiaxLsJF0VeSdkTfiIp6iIto76cmfoFBzR7ZUgbIZ
8x3wANREZC37s4bXExLP3Bhj3gMEn/fIBoYW0MOxSGlbz5W/liAZfPhRBQehZBYLubRXdkQ/qLVv
BseiW7zyjTPigCgiT+T0gUlPQXA6YmQFJblj3ElvaGJL3nb+EW9gau3/cTw7fkH21a6p5USQHemt
n1nLpouKJNiArjldZGskDRQ+euc6SVOCnaaMVMqFCNGYNRvZKjhqrlDFoZ3018XtlOGSEdXhwBEh
AdgWeo7nWY9crgKtWrF13oj9/xgPSjMyZZ1yplFcsDfpyiF8s9SIKlig8LvmwiBIpOSux68PBer8
CCl2ocwmT5xzTbwBzfpegF6XVMM/l2bbAeYCykzacn0Xdp7IyzJNZ6bTVl2XQuTKZ6McOX6Do/rY
yeDdyrg+gxObE+B+xGfH9t8YrNw2O53ecbpZxP26GMHiOAErfsNERzbw0jLCUzi9r+odoM8zFRmy
F8x2FOCaV7vLJ8n2vBZTdWM/qwumqxhvGskJA+cthI88gTMub3s7jz5jAjgaUpQvNXKEz5/cxBzT
Gp2TFcf2IjhTmbjnbIJUZZ7GSxaH9jgKnnwG2nu/5VTd2JrEKWjxot8+VLS8pIuWaPfmRUqWGQBe
sO816OmaEuS5aCiFzewMSl53zOrNKG0DeVZKMa1nTC/8GJAICoOdve7Y+LOU000AzJOtEeFW+TY7
JGWeedx+v/0fbVENH5KIzeuYbFUxbnwy2MKEd9P2TlmdtA2RVrf8zmLjJ4xXw/SJw2U/dELLvUFR
IiTPhMyvSSJ9dwjjLxQBXAJDbAxMoUgwHGgsyjmHNiy4oKOTZOeWGEHD5ahVafcLK8L9YcrXoddb
Tlf2YkvtJj9rsWRsEnni25gv98PTAxcFPKzEMAJKtmqVqcIVbQpr8YCUieybc5Svn3GJGwEtMNrB
8itY3UReTR2UvKGcHtevq8707VPfXSasCTQWg3GEOX2ruApFCiQVgN227vlCU+QojBmG5sUxJyj3
LtStLiKYy3PMJ7Z5+/Yk2GFeX3xO2hDrn+NAeteJuelggAFaJoeECuptjkhZxJsuhQRixrpp7PCO
3JZIxF/FS1KWxNwF524sEFHCNmdAtnUvHXH8jGCX0g75geNU/XYnA1u0tn4bhsralZ5fafv8RXla
6W+ovLww2qw4VoJucc+VWrAtgoV4cgfe8bbreK5hXE6QdzzFCml5kkNZSLr8T1gEd2FVquxwWLS3
i5QZ6Bz1b/UAlnw7UmvEZIbBWUlsiu5cCnbzA4waRVUVFBWN1LQHMPTJXeYQdW9wlIPcaEsl8I1/
vh313/ZrSDgT6R3Lvb8z7ANMmgg6uadm5CtRFRpbpa91VqCgRmf6n9Jpl3WdHpmbC00xTrxpGBIU
MViuf/Ia9BY1P+SlKskUI4hyXAMCHkZspk9zjCRZPyUctJORK5+1GcK48VdGUovAdmKDz9dTUyxl
e19qg8qklelpyxVO0GFbUMYpTyASBdxNHxU7BoPcqtxqQrQn7AKZ3ZvD0TtbeWnTSgVt9gy+pjJz
iBJmmCsAhpSh2E79nsBXl5Qh1R21POZWEwfOLC3fUqRwlEsam+qROA8779//ucgS7zvqNBcL8fdw
IkdhNfZuREjmMWbEzbST4tPI8+hOC9g+3M9kxA04QwhlWMiMsff+ZPXW9MNTBmlAh1Z0CV/eHLDS
lNcuGZrMWg+XtYdZ7gdRerlx3g1M3LAyf222njMOxn5JUGyEfFHOCZicR4/CKRiRrSw7x/2VcbYe
Fg46joJq+LFJ4z8h8++C8QWsZCDi2i4RydTgfeWhJpVh7jAL0RdiqsZ7wQyrK4D1gpbsDFUwI2l2
/+igglS4rqRpvFhSfvHOM4l5ea2Kdk9DmUjUg90FZJ52RavJYFeS17e3XTWFwBJ6ixQvQX6NZpoL
zUpaEG79ASVUl9l/ifdKn3nTOrE2qsfmItI4JfnTKs+rnsXly9lX2aWCR9mGEzoEdgKKobOrCJKz
8qD0ja7Br81ZmvxjOnI84TH18FQxhPDo7feKyN8ATeK9I0e5Q8FEZCPzMobivI5eQAJ4CligXExW
9HN+HzRHJZUpeD0izXSKyxGCG2YUTr89MDYJ3ntZICC94E+B8hS8ubeVHreAjIAx+1xe8uRYQCeU
L1HoGNz+iOgzBXrRfReuJJW6K08S12KHuydEJirgD0uj37lqi/nr7biedt6ukns35LomzMEAPJAq
LB51D2g/RWqcajRgbStGh4S4rYAS5ef+lf/rSaOmyeTC0naeNNVA2BzwFO9tQRSmWBpxtzAKATkc
ncXQ1os27vLqriwzWcXcIe5sFnjHjciGjELnZAE4yEv/O/kTzXSN3GO0DSM1kGDyAJfYD7/U6C/Q
fhjI84B2AOMTrHx4SPboLLljlx/DOXlJfW05nuy8G4ZexdEQPWEqQUDOykWpl4M9Xg+N5cXzjVhx
hqEM6VSRj4LLeEu8OTElpKbErxLWkltB0PJDI44R+aI6ecQrDgz1Aqjc4XG0uDTs4LhCS9pkRPEk
Y+djfQJBBwUnUwBrs/iWxvvlclN19qgF4ozfYXAf73EzudpzD7LvqBKrSPEaQx22P+VOT5d2DySu
S2cQ2QvoV3z1/25ydkBpUq8Q4RNeoyb65lnEnfW65YtCFScCcJSrAmEavwHyOU8MHrz7PQSBFNWV
7iZZxBE3Ej/Q1v66KNysKWKVS+FwyUFCEmmsgPX0uxXQl8E3i+Y8rIg/a6IZ6HILD20Hy6pbo0mB
MoUmNXsDg//leMjNvLu7psl79j8/pHb/GolhHk3+CE3ckQ069/jxdRqJ62aKNg3/cfg6xolxqSKQ
Y/bPDCLjxPssl7uwEbMTMEkVm7s9GRjOYOQ1IAwK2eBweI3hZW1aU3gylEh1d1rDZR1HXI5A++CJ
Av131uipfUI0ARIPCe0nzjn7jQm3+/elDrWxPFvV7bZIJltuXT02FdODz6HzVcfSKjdZilUU/KQr
edx2lhfmdIkseGVXIcB/pCoKtLtkKHtvy1oZ41BlipNKd2PQ130Ez0NmFwD8qrZX5iNa7KUOD2iR
ProLk4l85DL8gpq9O7LCRZKKckAsAjiLsjw0ZNcdELsMfmX/7u/Ap3j+Wsfgp7OZxBceuEvAG/5E
p6yF4iWa3LQLKpfgr8gzPnfd8glpeijQcwmPSW+oeUFzCq4OhUzeDvTvN2nDkysZy1FOjagvG/1o
3Dr+mEJcwo5VX5qT+56r4vt6RsJEt56pSPrenVWNtUaa9tbky7R7sCFzxKGFIRGtcR5JNhecj5gP
WATpeX5U2eW7cKS5c5DShCbG5AhDJnJq2ZBufJP++iY7Jm7DMD+MEIuXfJOf2TeauyHCRPDMx4k5
zEarWRJEHmihANdMZXW+lSxPYfJaXK+2BNe1GkhKDOxAblX6AeqmekTKBk+bthl9sqIHex7xkPgq
hP0uHSWPHb487yktSchl5oyWIif+EBHrGR/QmzndbsoSsfU7UJZcHaYQQgeej0oQzj7D6uHyRuWZ
eqEJeNQkW8C9reVZynGjhwtnEHrtxOImp+8te+32zWEa4VPlCLxxav+VjBPJ1fNyv3KV+La1xw32
IdO8GRc7SWDDV/EwDyk9gdki06dVAmo2Oqx5yfPpkmfKzctTOdt0nhdnjHz6IXJYtyICQXPUwhnL
Pi7R1jD/4pMZ+Bq1pxAzYZa7myobRGrpW2/rVQ45GLugKnFUzl4qnRmpxy1KxBsHnHtnev3VyPAa
tF8Si9HNjHp07doFA9suKZx4XmaJSzhjfFi2C7qSmCWoQBfuvwxgeRChFhrKLzwD/RR0zmTy/k15
pvbBQpnD/GTOsLr3BNK4zUe2ihwvqmTgL2lBWNwzMPmK92ltqMCr3QaJmpI36Y6SyKj9iVyx49Ux
M6tMYapIPCHLUi+AGcF6cRhwGYzGmXe0GflfLrXOHOiwRaNZtapjR4lzT5AYeNNX2wI/FzsVJYC9
+kJxrQebWt/rRPDjH3lTGjUs0kKm5GzdDpovHXrp0SQ4Q3zwXfUlZsEzfxWWDgN4ESI3s0IF5anv
DbVhuwGOhN954w9vas7EyCNDrWtZwQy7InQxIINs8ixMnRi7V9NivMqQoJR6kBKCJlSX+5LBlRpz
8Y5FQyFVL6iyQUZF9Oy4By2axhh1M+IjXDhmk/P15EWvBaR4+ykoyXbZ8vu8Qd83c5ktKktb5gt5
qzhrCuqc2Qlqm28DE4dFfwm8M5XDKnXf88Hnv/tzGQixUzW/iJLSj1ZSX6kmxNHDxNpyhJQCQAPA
Foy0YHwB3kdXKcmmAcxjwyeistcm0XUWbBw5rs0s0BEMWauEu2aIqlwzvL/6D7yxJmW35MUCcnXN
LwbSex6ASgPYfXOYKHT70RUdOQT9Omp3Bf3RwXo6JFg7C/WNCaIDb+rBBCUW5a70VpErKQanIzaf
0Znnx133Qwt+Pgi7tA8Lzq0Tlf1rOJV2vGf9GfumN91/A9oTwWUL89JoEz9Lm8KesOkhvSp03WQ0
AorMDQPVxVytJwMwk9IWCNzRWdLBwfc6t6mQcSABdSDSkl3ay5NsbUAbhwNEz91f9UCn9R1zF9u+
gr8qE+nIZe0jt1PFfCWcjcTxsM0O3kdy80oeoMmV5alaIfY0hYsUuNSGwiswQj7dLT0ucI1u+JJL
xIlFIvQZwnJzCsQBAekbriBrbIxkli5qBA7bCB8l/4p2ZhwkjJY7G58JW5tTSSrhrV1W5Bv5B144
Ujs24VspWq1QRvrY6n9BpK8ZURsjqrREQqduWLDOffU1KDZgwy+zbP9XhO5s84Uosem9Q0hpOre/
S4R+dnbzjV6sPRhp8BTeE6614nCmk/Fyirj1XM1bVBShG6/ry8p9b8l9FnJYV/5Wh+cGsj78RVQe
bs3NFXmwHmFZeag4V0XHw3YWabU9UZdT08UzM5jCQ45tLgb2EKjVRcWuGZ+0LA0okX/8N9szhtiL
qzePFank1OGNyHSOGUoJ5qW2caRn3BR68xOrXIEane+gafTMJcMzlA/aX/6XGq2sA93HeIWMURSR
VXuU3g+j+z0u0TRCLBs0rAel17UMZGqZHTrb1bZ33gu8BhZ+DANl8GiRpFgOgnLtOuhQpQKOlWeO
2ePON3Bq+AH9N/DcZBiFbhc2ksgdV6BWiT9DrtQcTutkl8SJ8/MPRS3/B+BrSFFYoSNheHtcRcJQ
fMeNLWbQxDndQvAZU8+c/mRn/e9iODbupTGGEueS/K1jBPUTKwqDeSk9Yobd2gI6k2/3Y7CGqQ8c
+9SzHcqBm5/fzRdylo+4qivFIwiiZxS903TJL8lns5dx1gGxTSYAdAF61wFFFxIMXeCTMGIZZCKb
D4OYUeRFg38iTUyAN1ijjvid2uBncJ2y3fts/cGNU5yUjZpVMbYo69dYMcDodf4Lh0/q7KdetOJc
It10/uGIkTsf7blRsZQX6JdyNaPs2S1LCRlptJv4rD3mj+kD/2wWPsPUs2Az854uOUZCP94PlUR/
fbqDcQlBe6t0Wc2ISb7TWJQ/+8OUxww4ZL11OoKsThHkSKI1mgLygHWnQOCI/gQyotsSmz9j99/7
309VaQOQigX5kr7jjDzuK23lL9+7CAdhADPjgVBtEJO1RtgHzt0qgDQKxE79nAej30SvMpqw+Yuh
baIvQc5A+cC+kNyxpq8GzPAHa4Jbwn0yviIVaCuN19g5SL4c6vwwbMioms1fxzEDk0gl4qRKqsSc
W771rwyw+HbaZsyjtUVKdAG4A9dUuyM0O7a8NZBKKN0VTC7lw/125Xm6aOTwL4nNJOHPE9Bxs5//
ouyo+aWDFyK3ENZ5s5eLCeQxLw66sYpTw60tWUg3cmLhmg1Y+W4FwHJ5gtPnPp4AjKvAiPOmxajf
ffy8fxrD+OJF5W+ZCciQN970uj/NrnsQkVABagNF3zBXgLMOMsjC+94xz35SBeB5IlKpSF+dNd81
zAhWAasqBHkVFCJ1tlB6yJ4hYfLXMzUKJvK/L9F3m6GU3d5gwYHNAB++2YBSpI/uDIbBSkIDocRx
f2cmA/dAPnWms1Rb7UGEVRMmVVspOzZHTzjuXCbYacxAK9UCrY/CBj0blhMvgGRYw9pD0UbnXaFy
8QzcuLPPI5iMJI6zh8uY1p4RXxnwjPHiyIBJ+AoD52XPDYGCDD1mz5t6vYmz19cENF9aLAxjGNuU
gEQ5gL4+OioBYRhbhx2uR+4WWScC8UJaKDQlzXRm4yOtlm47aj3gjEyZv2uwWsH+C5ir2WqEhUZV
otU8c3AKBCyu00QItSQYe+x0fIqNQoDtHP4HeqgSoWzo7ilOUDioFX0qrv16gpgSXp0VXg+6mqyh
tyq8GpqYIF5IgYzicUYWqVnJXgqBdOPeIZZGwnJgeRixMoY3YMXRVUqcoOFuzTkhEKjaUgtiytHX
LhXt+qA29fBKboTxEiD4FT/wtR5Uz7WI2pabzHS3ZYAmwYnI0EzjGrjyNQxpfthbiSv6y9PWw+66
cAj66A3slgs4b7Xb5hhJEhvVdmJzWz8QzYOhfSB416vshn1adWS3f3qH8SiXiFLHn+su0C3jX7Sw
QGNBVosKV88UJZZx/dZnwRPMrsjfQtUhVOGGQCvPEJKwLRRJ/uUfqHxuo4zNkX+oGzBn/rwFVvZp
qvTNPFug6twuysQzu1lLRHktlFcOs1+WuwbhBV7BU4kkyslQhfXHVTbYTWNTLq/be4OnFplfburN
N+IRr71mtCXLGuHRqjc3wcyiqJ8pB45G/X7J1uSr/1WAZmyVBzOyJvp/FrOJPRPKdKln5wBaPB5G
fxGq35D0N6XpyUye+DeZu/o4IYZN+Q9YWK0inE9Mx5eNBawTFYMQUie3VE3uogRSBs+9vssKCqgh
bRFORA2VI7r9PuD8O7EjpCStiBNVMsbTVxyrBfoL+qA89tGcioQBE7INNu8i7MkB51stBzcS4yO3
HakeqyzV+VOdism5UOtK3l4abAdxDXYNzuqg9bcysslOI91eXBUPCuiPi2oXFooGcYrHOInfm+nw
xvAFz3DunEShOoHqpA2uLshlXNziQSl0SOSBezgFF248SYcDZgLuoVVs4WatK3oQj3sa72tDNMMn
cjFq8JYo4qFbBuf8gEJGwJFOJSch8xrE8xpYFGir7StavJUhaQbjNZhmKB9qqQvgFoKDzTGXq1/x
kQbMfDfeR6hEE3J0wqnTgIfFg1Jw1C7jJrDMChZAxVv5X31+l/b3w4hN54yfvt7FzJ/90rlvv1np
FKsQIfgFYmvY3YUrzUQRLsFu4Sdv8fputN+mdIAb7Q2cD6hv2J/gzMthgdMNzO/dcPOa45XndT0B
G4EXeO2fh3B5/QYYdnHbczHwVj4tnKhJwEnsJH3OvkPWWprY8t7RHjffyhH7629LGbGzDRNWlz1V
kccU4K2cYdUJqrS0NFa9pLuWJ5GaxK/QFopS4TP2W7e/LTijLHJmA1fz7hB+HhV0/VF6/GZYoy1/
lT+WvZyT47OZ+4p+8/sL7MvdtdOT/4qiSAool1fTD4Zdb1dQQb2bFNEtRTGWnBBXZf9m5+dL2gKJ
8l4hK4psbtkuFLxDv7KHTzonkYRXroUlYD+b3gGFv16wLJY7y6m2vQNQZPn0LfwCfj4hqndHSwD4
cKAaRYbotHtQU7ga2GYPHtXmnjnpZ6K5rnElC/wp1WIdneq438gvxuHa2LO859mPAZH6bCUKpcJs
Kk7WoSBxoe/NLU+UR4R5COlCHzY1ejZNwiMUrCzS9tp2ypE0T1xvJcDno/S6j+6aIu01twPacAJ7
TiUn2yifHzh1829riHphj4T1sQJwZq9qFc7axAMso5ONfI3CPLbdROkm9NxDlp47jAqqLTdXrH3I
MnY5QOO57nL/M/YxKQ7MOvOzEScgEb3Tufv4J6VkY1PvaRVg6V/lO5MwCbRxr1JNe5nANtjPE3bf
MKQc0rrWVgeLsjqc9lMEN0PkEbbvF11pkFnHuC0iz+83ORyeOXEi8g/TesTMCW/laS54OuKTATMF
OeSPZ9kVEdIBrvnoyD3Cim9TM4P8E/85V6ZuJeGQJtM6SC9oC3BTLIlFTsjP6DvWpruhYNEZwqEU
jwivNJaExY7/lL2TbhN3iJkjygpme+J5nBNCYC8ihjBNWd/LlFjQKRrWVWIkJ34/nvG5HpggQggd
tDO78Yqd4BieygzeNnBq92TIbzlQUYlLu+zK4hhFgAWf87jvH9beyi+i+8dIyPDE25me+xAGIp3a
9nOhXl12y8RCYUWmA8XmEe3AeAHtXqZXxtN4vTgFJIfavI8yCM1qre13TWWOqRWKc+2Gq5BJrc3M
Do1HPlMu1obgiHpuf3A4EppfYe8ZundcLAPDBBgWZiso/YC8aYPRAEWq3+AWgR0cqZoJozYlEugo
brgY9z9Rh2LJ1Y5SpiGLAYOfoOOg/ugfxhOVdKJ/eLrTH+b8R3QKz1TVYoMKNhR8FWrbhES5sXxT
8jIcbUdh1I2QZYudNziWvA1pUnoyZs2NJXcDW+7SYc+A5/PYf9NL1HW/Nqx+l++qEidYtmkb9wWt
+bbVwGISc5/g41gfSdP1ha1vGpYnrZjVq3/NaWJmON8+piS2wrzuUUMe6M0/hCpkihNJvrYcU+md
bELHfhOXNU5WejX5jv0eIij2vnjzfmkwxxlyQQMw3hqqGcj90luY+q3umF2R6hAZhNUSsNBwLN3B
IsBQyFTIOgJzu2BaLrEwhCNB2BbpzmNlPS+umk9nZqW+XTKYnbxOf2AMh/eLZOdctItMbAnmsgVT
D9mgdNOYbS153339p1ZPtHmXnXD5wKxt7lJbm5RYmpg4QJL3RHd86yAdIm0JMFrgHp4fXAGSqNhh
wq3CEfqBtWhg6a1pUtwNMkLaZAX0crpc14LlwIKbytfaB7fbDrK3pteNAsdl1Hti9voSIZ9vp+HC
3bMVOcki8vnStdCzotXnP0wedWDDms12DbOb2yQlJN/HI9xjd260unH+vJigDzLHB3zxeZ+qW6qB
vKcxxxVBBX2VmUGpoZO+KE3lVgGKYTDzxvnJ59AlG+PeVRDhxi851ycBTLvW0Q8slqXgZWPWRraq
X6WTSSmzCAQy2WTaF5MZ+5y8EdqFO3UNA+NF0WRzTMK/FUGCgPUGxJem9oXKmdXz7Bo+Id6R4xaU
TQkizX/qH7axpHPL0diE/HERWo9BlHFms9Qc9IiEvKZhHc1/socOcTiHj/o4Kp1f45lGsJUS1oFG
KSubaxXQhAP6oKaibudXHvjXbykE9a7xAxuqCvnqUILQkYxWGzErmGlt9M5Ct64X+6f4XXd+eRdD
a/fcSrxwzpfmb76ZaKhX+QGRXBOAnI5ISxkbPxkjtl6T0OhAa16KdfUV7ztIhW3bnKqehqgMUztE
I+2iV502I6uAlFB1qBC4CbzXu31rmYvtbiezhXMxMauoyjsmOx/kpExr4jD9aT51Md+e412nrDuZ
7FcR1hoQaL5vmJgwkr+rt5yoK0pbpTHuIQNJIET/cGdzGeFcjeQMX8Hybhao0PcGTrD5YHwKRZtq
GoVsTLQSVPtBVDZh/IV8cD/nDm7zc+T5fUNT+jc3nU3flkwdriTYGrfJIWKdZcGpR0jU77R59hBN
BGJv9b7gmwrv5g80SyFbDjwV7yz7rEsXJ0/EkioEd9oLKt6KvnV4SiegtlYUBqPo2KJTM/PTp1PA
nJe1kFTrYyb1ZYM3Z3Dm5fAWVpVoFxnVH39dMnC7cp66dSfVufeCfo4amsL0t0A8huc3O8ETynLl
U5dcVvuwtUzKnXiudhKhAGoNqxZzoBKGF7gcEt+jJi07QFE4PgcDxAKPZY0tWSc6evThqKOd4OIb
+yMtS1nhkseHHkVtLr8/TNxajWBGKKngQkYhK4jzXZv0+5v4joqfSu4SrKPjseKTufPTRh1mROQr
CKJa5nD2dDwr9tGKm6zx+fauXOvu46sZwSO4nExZjnOq9nsGQHDHKgoT9LZFMpwhwWjY+rslCFda
NIej7NCQnUaroBpXMUbNMrKsLPgn6OYz1e646rB3DbE8X9+z+IM6vywt9npvKNi5UUVCfK3WCdGi
Tulu61r+2JliX6ZTNTr+Ufhenn8x09UgST6w7MDSsQcYl/kbRgHFTmDApVtcJg9rrPRVZkvKKR5y
27r1UsxiuxhKOiPnCdRbNR7mH1zhRyfNj0lyJYKg0IZqq58NuUM50QqyWXWflt+AWqXdXN6mc97V
hxdNFzw2xcMvyJiAQY1BcIKYpkECITv7M0tEgOMrZxrZTv9TrgPuUbydmCZMHviLEkCDWBEPPNG/
84ZeKQLnsuN9fdIw/5ALw6Zo3Pw/Lpm8CQIXE2srn0Udk4KEChn9b4amIqNZt6sRt9enS1fO5R1b
ba1xmkHo6aGxtej557SiGvfNUbgahhN6nzBICGniOAnpgOJMWZ0qC7yKon7QYRSpEBHCCI0TOlac
ICixAbRdMkkSlRoa07GtiwJ8rrVB1QHLV0un1znFk/845FvRRfSI2b0jcK2me9XMPWgBkwOZSUlO
YkS9DY8RKKxE6fsNq0T1BBXoS2Ff3UhGjP3lrIqy2LY0r2bHsoBupc+ZYU3C6xICaKjIu1K75e8d
PBqiqEDw2TuLl7nUZvZqcPaA06DYh/jkUCAJ4CDt1CWiKq48avOGOfqDVrL209y8iFgw5PbbFtFB
gonHSDMMqnMXOsW2FAew185YPFYTL/pO6Sw7op5YCrQMGSD8TrEYDOTYn6H5AAiKW9vROY4oR0DC
4YukwHHUrmr1dKj8kXnKJapmDGUN2bKCOGj/6OnFUVhvbDR03xddPHKnFPBVaLuYjV84iFwYn1Wj
k77QoFPPm5jQMsPnwdXANapS93hAbpsXC6J+bbFaWJ5VYO74gnP+p70Kof6T5duBQHcnqjZhzJwz
YRF0+fYCbt5EhJ4yqg91fgRyWpmg6sk4+bAuTUbuNGL6wjn9NECpzISQu8+W3qxuotRVXsXt9OJj
ojU3EINu137IOXb57sLefCRtKsuub0QoflOevnOeC/bbWWzZAdv2iMTnssZL26ITVtpZVKPNqLHB
JE8emyiPIIzmFwi0b9HYvBkh9i9TZ2kGMNIsqL9zH8WGX5EKEM8LgrJAJDuNVGc+nDDD1nNooRTn
rFhIhG/LfvQcQpJda8oR7AfutgUZZ2el3PXX1tPvs09QAwt0anRCOkKsQaaOGnoVYna/Wla4KyEK
6e1TAPTrSJrnSaDDW2dVoZiw74ZWge1u3giBfMmBLjC3V/a1IKiC1wntDqKIdC4Tf2GSIQ+7/mvJ
esEKFdoPhJb6f51JplChle2OXBJiFR0lw4Dj10W2KS15jnfuO47pubOVBhO6A3WAJG3Zdy8EVWNo
KQ6b893ogtf1RgJ5BNrIJH9DLcfm8JrgfQAD1niphTjHEWgQa/TRm++Xa+7UHUM/kfDVnqYHpa0u
UVhN4K9l9nTf+lUjHRAE6O0VHMjaVWpIkuf9Fv66vHWSDUPNI3XpJWG0ftzt9nnz7RP+w7+yP76F
y8220G1TWaXKTe4jQFnxBUse0gmSIxSLocMYPjuMNd5CnZZZbbqf0XBjjiVzaCGqiHHdpC26yQRw
ww88ceMINvjRZa/QU8U8bhOJRu5WsSd0RS+qOauhJik76p5CLmh/gFWXNzsQf0Ye7IdcM9NcjHW7
aWWhnalv1BA3VitIHsFEqfkSEjsNN9QtWL043HdFmeViCVRBehh3XJ6JFf0kPJuJa++u72XAbpMA
h6b5NLL0UJ6XE9dwQ/rdCuY96ATd9tO1CnLlN1J6CxZMt43zEMHyBD2Zwx8Z8b/omR66BPwZruPD
i5p6qCxO6V5cTq02mdcwFpeWZneY2c+jHXwRzqSktgEOmyKnmEmnrdQGrptpShlUvIFMfpG3wP6h
XUOIj30aKig4HM+depCIpJqouYW9dQZH9vqY/x1sSWrLmw9mr52lQ/BqshUtv5J8qIF3fnuhBGwU
y9HFvJ+51uNNOs2sp4V2HnKjdrAu/8QHlf4gnlTAegsEOtra3YRJ15v29O+Fn4uUEU6fKkY95h2M
xQEeLb6KWFLPwZu7b+GA8cEmJcAL9ikQ398pFgWUZI0QXwq0DOQrnSdm12A9bNuv+udqymbJL0Vr
Nba0V1uXjhZP3GBCvtHyWH5ewlxMT2x/LMU3cgx2uMGvQTxCClFHJLAL/z+2Yd2dHqysGDa8+d5C
9Km6ZiGxw0MmvfavyNbupkTIW1TiGupsYI6+Zj4aTJ1jb18lP1rcsH3ZkXowDJBEy4U2St82huoF
Y5obMbr3lO3AMjA4K2mO/BCJMReaKss6pibXtM9XJUfluGjUqDS5x9OpozzArbWQlfyyp9S1rA70
RkLPELz03+q/Ui4elPHtTFjd1LtqvsYqNiz4jotwykfaFF0489b9gnAuGP41bW4UVGdcTtWmNGzW
el4hADKHB6/GyuBvAfrZhkzpNQGOfgZV86MTUERNMdOfklGyFs23eXn/H1h78T9JLzM0IS46GbAZ
4hpzPkI2dxvPDa0fiZlB3ofuXdFaJ2xbMXZVnB3gXsH0nq95eTQ4s8mfD0H+0jlcMaOgjlx9wh9/
v2mX/F79smO8xO9O7UwfukTmgsh3btRaPYr3bnz7vxw1Akv9AMPlBN3VmtLO8nDmAan1dIpM0qFL
o+pyA/X0DtPwCqjsHMUSFjQsJs13+t4McFgDfl/VCQhSRMNzc7mksYJCGfncnF79QHf7kKGecZbx
JQB+yxO3XoCa3xPNEXKs9sJ5HjmSudgstJFEVel5jpdG0uZRiS0RH+0TKUjbXJM2XS2rSa/7badr
f82R8aVw/nd4aqInRu2LHD9kP0zzd9jKFH5JswDj7uz1FEimORGRwGz+1DkATxlPJLMsoasHOaaI
UGL5X6o3v8JvbYSNm1+gEASB7/0cMNDwK0xvB+4cmL/emmemd/djl5rMG91FB7P9MeG4crI1vb87
r1lrp3XmUd31cw6NwvAQ7s/XUL0peNnD/pei5/Of8b+/RHs5lDZ5xbaDb01ggS9oxBSVs4iicJgp
Xv1dXvS83GyolNWTGecgtxMrvAdZhWu2N2lK6fJPCVt40+yjGGa1uKtBYjI+rZ6Cp6KNSLt8lgo6
oyMJtAIsvuPT/Uy1bInXCb33RRFPY5QTr/IkHNiqmYEH3cO517j9GoFh0GlaepAYXjgaH0dSryX9
ZIA8w9+sLJwEq/KKToWhxoo2+3phEedydvzPUioX2a1oqui3KcROVBI0MUOIxMdihXgRFaJH7IXV
EONHhY4wXtv0n+3v7Z7lfGYOSeRI64Ba3lQtwmCb4kbr4+LnFhk+FWH4GMxJMSX6nQFz1fly0SVT
ptiRItJjs7481TT0pK6jeosB6/5olxVB/Bmm8i9YS7uYbRz+qi6v0zVj78d4/QeQKBr5krpG7yyD
HYt1n+wjItsV4hR2NUk1241Z90atfYUKfYIuI2AvfuzTWF9H7vjUDagzJRVGV2VeGTC0V3SinMvE
3tH5NKkSFS+Y5Ui7jZdxUszeeLthZwcLA9iWXgXK9kfKZ1SOI3fqbW2q2JG1JqaR2drBvJ9ZI+Ra
5GLo97djkm7hjnQ3kJnzk5vV+F8VNb+JtssDQRHZ4PmEl1//5gk7jQml9SVtgSAQo3NModQCdEjO
3GNlNIuGtFFDPrRyjtDt8I2UGhYjjSpk71517n5W7rF/ylrGdzxtaWhTL8ZBFoT3/BFrRS9mbypE
CVsqbNCQtKs1bqOUxho1rea/z4rtSAwcxNwkHmGz/S9PHax8tAW4pdrn8CA5RLSTwd7DuRdMwhQM
RlKFHTM5VPCj6It4eG4KkHynFzkZOOiRR7CTiVmlYelNBTkdfAxbLeVDy7pG+UFUlykS4ChlGnNl
9bYyEw7Ws3XDrxQU6mG+dy1vtYiC5/Dcd2bQR0cPDydf+427deWTOsElJOnoVQP0nysAGB7MOprM
F/q05an4cVB5CdhZsaCSE22qDvpJiHXlfLlVz7jq+iK9DtQkOaFIFwPBQNZNqFv85P2FWt7PukAq
BcDliFtWkXqgKjNqPfB9IDqr6oPu5xpoO1ptHqnnMICLpQrPeMhNmNgA241NDHl8kLX5hFDbZjrg
IP++oTGdY1Gzu9/zxWYb8YPf7uM/YgdT7gU2EojIIpiQeQOfR4UPflXCjQluhti9mMTNwVYaDhjv
RUY4xqr/w9EXpTD9gFzmBM8eG6Gk31MxBDu/E+FJ0aou37ZZ937wvjd8Mjs+qGZvjumMCYpX6E4m
9m76Yba+maHyQ7T8W7UHdkc7tW+A0whPXIlpQS5tQh4l7w7hUWxLRr3Wen2t1iY7bn0yRzAa5W+h
dOtZt3r4B2+qHvwfZcyQFrV78Vc00KwTNWuK937csQaWqn97n5s+nJ9BLAFApftkukKR5KIfIsC3
smwuT34rA3wFptorSx8PIHBeRM6AjcDFKVVpcFy7R5mDaVNXDYgbyhV5PYrV274Png/ONs6eosGS
Zd/YbwkugTLCnfR9BXCmQOLqXg10oW7SM8jcA6Gij7eAOa4V00GUg+rkHhihYdZ0w8c0nY/R7UMF
3Sj7GcBxqZbkxgfbhstYUAdY/M/RbPI7Ds05X4SdtBnYgXEalwypye+HZAQW4bU5P7Tm7r7tIqGX
pVjo4tSIl88s6vGFeUyOkwZpW8RyNJC8UnajGph4m/Nh34/FMDoXnc4a/bw74/MHPkrclyngAVi8
++6S5RQk3WfCzqkc8Bo1dWCJPebDK5V6QerH5bF/ydEhrZv/l8Py0cINbYrf4KojyL4Bj9dGhOqJ
57k5EgV8e0cxXwrXNXE3DUwFVEVJKAgA9+r+IW/PEENJ6mpMLbefWWiqixMO9dkbnHal7NW8JZNO
Y0nccGRMSftZbnvoh1N4NpBrd88Rw1HN+abq4PTUJr0Tk12+BzKWxd9sVIg9Z7onriqTGIdRSAX5
XKF61N2M2i4uS6a58PENvjDf7sTq0OfUtoMeSBK00FEUXUqsPulZzRWFVZuVrvQYm+b9RJ3C1QWv
aGnlmrGa7znA5NfboyVXDZzx8Na6+1C+1uZGhlMP4qqbPydGFoTv7X+ISzIJ/hdyttZQdG8LPUs5
HnKB2R4X16K2Jvd3WsC+YIb+jkkboM2+pXb8otDwe8rZ/bpeOjT5CDL/p3N5rPOqMxWjZiBxHKk9
M10lwwMOMN0XQtIpm+RTYepQkSZoy4tKC8I/RFrbJSK/y7YpH3R6+RqMmcylNh6BJWxQaNIG+lCe
N0cuBGal9DOgpsi+vIPylMJaskmOsEs9SihEZnVhm2xJmJ3YO5lyhf/g1SudtDlgq/liqOCLaEQv
nej4OGvO81k0VNoBk+NgwJ8zeBpUUhgFeivuz659a8XHVysSsRMhZZq/YdP3OEipp0jbeBmXbKhN
BDCoQEmnAOFTqk0P3eIJQC3eT3U5TTv9zzWHpuZ3jwDt5MltbUNhu5oUtJmVqxOVbavDWXYpjaas
wcbMNAJwYzzHePXh1qhRSgC1wCGcyqdHvlD8zhM3RiZV2tSJVUnI0qs1RRxrKxMxbTcPIzvgLGd6
7PKt3LRXBMMaLr43DdtkAGzSHelvKrdmfqvVBRcFFFAleh7xsUDbR4rsU6jCQXh45jH3maXViDdh
ahFRQw92FO5zxunv/2Az3F0RcN/7pHO6ZMSAr3VJWkIHRzKWaGd/wYyVdO0B7ITdmoDEMTD/998x
pvXr9pc2hnDErgjuXAb46x08BxmSxJczIRI4mzScN5S5mJijjkQtCnBy8omOFR9G/IuUczvyBhiS
JzAGbCkeUzRcX7pWPMmbdU1KDKCnp2DvpZw20vtVqJhTtgjkHLIInGs9StE1W6qObx1VmQkjVmMz
TaqoCbsmtqqevI5J7ud3/jbIXhtbvyAJoxYbHmpa0ztu1m7wSOUxvyWwdIhE7TY7P2QCn3y3bHdy
Qu+NLHzVNHH2QHe4fYQWdUOhrr2H/u/amsdr06m7IqgbC4iif62tiKEvtethj2IZmLQw55yY9wzi
tzwQJq+pbsgrgAQlOzpQqR70h2i2WnmBTTq1/ViwhHtNlEMYUSaZqBEpdUInxaq18T8fqg6ajEbg
Qgz0zr9NnKhHIkQp4YGv2QsGVSoZ0zu6q5qhZTCXjT/z+pD3AscNMHwjnkDxMXopiP5mytaGlEwR
G91MN2rX8M9/vMc7oue74DdhYfMTm+LRyk1bkl37DV1U/NVVx2jXFYFXd6yW3HwSlgZkJGyoO5sX
FTkuHpk/1YNbtfOYtluAf7RisP9SfRG1SXIpA6w1ll6BLTI8YGUQSKj1bylytW+zjGeKgQzXdIi7
T8nlF9nVzuHLpx40H3xhSpVhIpdRg6NXPJISaRy8IzPN9COd5HyCOIxR6dKcKNwDgwbzNkhlT6Xk
RQXuVty62lPkQ4xiQ3uGkLoW5CqljOCaUkOzqa7PAXF8fCzUnzhO/lgWp55UXl+JDnnznLjM5ykz
lWbjKVlDHtUPn7LZWrq68zisckuvb9N25j/DAz2THy6O/QjKwEthcubLQMAXU3i4RvvrJ4l+Cr5G
+Vv4YjenODHkBbpcEujBXNpzQWHWArMybAfST0TXTIGgfR5PYssIiG/H2FlNl0ZQPTthkhuk7zfE
/m3iY5iohUD3DQXBx4P1fynPp0sB8Do4cKWMxmyhBSE3Wwb4X4zvhgNbwl8hrt1VPzqp05U+7J2A
5vyjEv6qd+x1u/Ccvhrrwxz+oHg49mKZk1Kcj/2+xGmA2J6luVoQEzfXbHCplSNNU7Y+4W48JTaT
Yu325Nn6CBaVlpdV1/ctfO8jcLery6rnXxSt88wfRIFbSw2N1/FXbxvVRcV0u4AW4zVTeNj0HrYa
Xk2WCIllcbuGn1spITXfV/WbzAatczLYPNKnWvZ3ftZ5FGW2izWjcTPNEHLl2pdhnF/m0LHGdPGw
z02TUcV4Zb/MO/Tu7w/Gf7lwYvhi007cdkWxgyAD0MLlTYq8LCuqbFogDfksnEHdk0R96rw5eQWm
UsWf7+XoRJf/h/xgLnhlokQI++3TynEZt42xKk6WIOqZz6ssFdzmXxtjoPZ0lcHsa/u+9y4sljJP
Fvi+8mXGYlWTezAE2nqrkEOhIvq62mKWZVf98/7ITs0vhuQtP9mdeQzzKxxKp5foV1Rbs/azzTwL
P5SoQgpk5iltHsDzk6Kpn0NTDaDuMqAKUpKr+/TRGUPGDF52VxoHGMtQj64E32+AP13b4FTOGwwm
xgKu4dzphw6qwyc/fjMqu/IO6cSrAz7T0bV6gX+FX+7RfwV7Re+77lcykbz8u/IPHg8cbrizQmeR
11hreIAQq+QhaSxlyImSDE8WNTLBaxjL/Hyyq/+GyZpJYQnFCQMJJYLntAAG5bhZjfOjPbFyEtdZ
Ft2B+/SgrGbD5/ghu8fS2rCwY2YSvxu3p44MR0dq/UW0IfMr4N857WGrnlya+HyWln6gLGdgiBQT
Sw7Gbe6GEynTQSdEANas6Kji3HBcWnaQWoOdmOIcESWkAfdnlqKpVQqLEdiPE52lOpjP5VaQFmtE
zbDx2OzFubbzuvy0kHkGdi9nbk88oFJ0EQFSFx/Sba+6OPvNlejayOFiivqF+HbTcKt6TVhGhspl
lQKmRaOWbfrrHDhZGzD6cNhEKRL3nt4u2LLfgKWRnHm6D1RXekJFkzlnPqepIg7rqEWgRGwq1KHs
tqrecBTeiTRXvrU6dBmNKTs9XY+LrjrHB8p3G0n533piC/5qA63v3zBdRP2OxVfelDuYMycQ9a5G
HEbZdHFrYWSfEX1U3kWOl90g1FuAIIq+2zQ4QWr0xlZKAC34XHIE49hsTa1/hWedcE4xZDlkHV8a
jFfhi1S0uOG40uvERyotf+yJ7QKPrVXbx7nE6gSBymeTvao9Qwq242GUU2PIhf3zMWL6wIN8NS4v
2USTDL14CaQXfq8gvjvs+tNRoSctySLksRUYCTU3+hzO6Gvl6dhcUJ8VeXmu2zUdzybaovxWkmbA
QJix5t0tofJP58q+lazWDU0l9FNUozGsOqxB9px1+LVfddMhdKpS+xoNll9rnA2FpzyKpdmVWOU9
mEyTNYfyA/83awtM+VaeO/TyXuAyNcOM+INNrNCR5KSBbUMJQj44iZ0YQUugV5RZhu4L/pYefOS/
uAxyKY+dLDHYCy0W70L9fSrbb4IaWvveLhSOitqK8GyO9UTXbfGlFeU9d4aIROVvYukWPdptCm2e
Ybz1vCljNm73JdksHyN7ShqyV+KKSs/h4ErRSYf7rz+YEa3+onmn3DobsWkciHZ3zLKo/IwTdg6g
nMLn84NaEKo2qGXQruDHF6Kh/lqhwI0Ko0BrLVQUY8+j13kZF/TRN2Ihko2iry91FM8jibvjh021
vHYSIQSMoHQ3lPyHcBtCqiCQBc5wYdo24BZoRmEwOpft82K6SLv4cafLVAw5SiJERpZzaH6yLroi
RPVO6e0zegsYUPwMSPQbm1u4l74naITM6jIqZU0wvNBAtalBxuFi3g4LAQxDC/OKHkOZj4vojTxz
CD9RtFtM8pIdEWUcvb5aeAwqNyg2/XpV0MpXWhMuZMCZEcCOK0+CvBHOterO8eGjtiZ/Nj+SRtVZ
UvVCCbiqNeOJHrFyKl3olWinvkkl6y107ih1xO+TPdsvqAMs98W+h1Dx7F2CkGgymPkUtrn2J7oQ
/e2z69V7DTWjQOtxDL7LFLYTPCp9pSMqyTULlmEj1oMMVQGHit6b/eL8cBgAezuD9MRizgX67EuW
2nB+NGVQsZMprusSO5hKY7d4jsuUp8IgJCvpAYoJD0WjZhGljJkxIlCIDAplH67tj1Ij4wFUuKeW
9LIaJZIehzfdalNsn7FjhZb2RD8Ds7h9UNAPwy8zuvJomK1EPQTi2vWbP31PnWq6epfmCrSdA/8E
RhuydMFUR/MFS5vzy6cO0vNBClhx+CRvq13j3+0hXIbkACSX0reBt6c5h4xDIhZUhhkuLAmegHRq
cWXmBlo0XReWJuwPpVNhWjUdYlEMlYbSZIhMSp1cbEvTwCzY61OmU/CvWHGNUcRe0oM3sfS1H4rE
w0awj1aKcpJpS90szmi+kZ0EgkYWLK+qZCFMG8FatI36PC57lOtwL09dGyQmALok1F4k/QTB/EGl
MeLUx2wFiJkA9dUY3ozHeXke030A8QbVINi4ozjRuz/3R6KMezWbnVeECHDeCH7d+Rt6bpnobEYy
nBS8fgmkmYioj5bXeIK9FioduKqQMyHA8ygFaDx79DcMuTrMZOZ1NNN6/vWysL8Ed0K2thwq1nGk
3hcVsN5oENMNBEKwr2xdHtkx3vuddF1BQNMJE901LVxgishZoMVfYG0LpJUUfUm8g582EPL1maMk
QXwQp8rkKcGugmne8cZBzvTS2YEhhR+HEhzp4pbiu5RNIuyWCyx0KuIfcw0BYGD8OaH4ihq1a5XC
grsAbhnR21HJz/DT3svaPjvJ7nGnm3bmHr+/aiTljw8Ld5RPeoGKn6OaYQjWqIay1/vRHSSdu04F
MsNr2H0CetLpeQimzldLSGnJAJ9PofMwYnsJ6d1qSQA9VP/6NKhnuBtJA07Tl0sOAzQjvhBUlVvE
FZ7TBRsVPBFazgivXwl+qATWytsvoqcOmrudOWF7G2MWOrPtRDTt5+jaHrO4ZWRgfEXAXPUfPn7Q
o7dZOcQGOkRmqcpLiAw1YQpjE12Ghn1uZNL3LY4prCESGQK6XOwCvCu2QNULCQkRdvZ9HQwVnYbr
ZLe4hHSsfgCzUHveZCNQ1AD0FLMhJCCxwkNlEB6m1g+ibOu2TOA5Qj1t5lyuMT/IThQwkJZhtj+m
ZWC10JqmmWDx5RCDB+XkiSf5uokBJYqvabix8J/8PgvhGR2XuiqC62ovguBQewBsTwcuHfbaXl7V
rJWk2yOG97E4RLfHzy0FaJZIA8GBQ+zzqJjecyF/L+AE4OQmjJOodaqTCQcHdoUCfTMhjT7a0U3O
NTUNd7qVZXlbF6oO8TapCp0Gz/su+3oG420rkNCMJSMvBEYrFipUkK5ZfdesM7dt13IuPCY12qFO
mUerujE5LOOWtX32T2ONBtAj9BLD8M7jyxtFLluAKIv7Yhn5dssxzLThEkhP55OexQylZKSHRt1T
O8P5cM04JltFAsiRsBAi3X1P7VkKHBC4aPcEcPvkeUXz9E+Z1SJU+drWNrQIpucTouln2+hxqWRG
tnfUz2QTpm6PujIluh+yuqukdsMFG903zb7Ox/F/qrTO6pRApKyp17DAiL3pDXPlDKoJuRbB13kt
v7IExqoVVDdp226vvVL3fdtMesWt5kZHdjBHG6Mvvs56HwFDAzS/obUCJEAp6hNKDEHezwd46IB2
GXcNqqo/CfMLBGQW/0N2/FCWvhK2rVDC0SRrdq933jllVYZ8/lmryF1fKs7P+1SVN6gDRBvIKwOX
xK5cz0gpJ6Bl6c2+zFhU3znoeMIGuBaTAL7gG2GcSy6O+V5F6Ituwez0FwWQbv3ZOGeqw0kBnm6h
FD/v3tU+eoKOfhazubbrSOox1rZ4v0wAa9pBFIizBZY4g+SPkSpAANz3063KEZuL6UpoEUw4t5kF
hveTLYQnXsv+e7dp2pUpnyAJyvqnygeahqx2eKB5cPB2sa58F0Vz0fm4uE/TnmuEBKbKz2WN5nZv
A1tn7cPAqnOplEmM5UNbehrnEu3fz6O6xZb1JLHpgDNNF9xmCTaqFaKiy4+56JNRyjfO4m4WhXVE
tQUXmsomUf3XeiOsYzPt9bB9S3v/EGfthETen/0lc4IWKPzhdKxgMJsam78nE0dRbNzzPNucCqgZ
H0xy0l7rxDw3hlXN39BaBtKBVh19Z+zqQlg3x3PEWKeHPsUbg8kxQsBpuBREtMt9AOKpdMcLuClZ
HiWC+jH2gCKrNbSXKx282thmd2Uux/iyPcwU498EeojRuRAPFmVe7wucHJV7MzDDLaKYCpyfRN1o
82O881LbJ9wRyi126Qw02qoYSNdb8jR0u4WmptHDFaosf+LKxIpGTX0hkwDPszfsmutW6ypyztv6
6wwNu+869Z+mHcMyp68ADkCPC4/wKEc9R+X4NCA7xhjtFtUvQQ5QzxfBOEOPAj7hsx0LrFNRB8Dv
jfEfn36M1XLDLs+0BYP0gatZEuUdSaOGhWFbo0EUbWyTuTT8/+5yZNylfrfka9zxwI523DgB8nxX
0EwUsDiud31TevID74O3ocLs0jewjtR6zC3vpd8Azpyc7szUFpSLzvjbC9pY4pSA0/42icK9QiUO
nHMNNprINlOO++QVdlDlhtxq0fnixWgjeBmozOMNqCCjR/kLGIgph99v1K+GRij2sOZ3INMxpPUr
RDhcbpRARYRRI41v9+52puoNRZWu4khvg+CJ3daNIlfR2cs2vZBjPr4NifR9NwhqfrQZRsexAhll
TO/qD8fJKLmIzHu4ZC85k4tYCFB/xG332FrUwMg2xAH0+zF1UrZjUwgkmcFp2ESNIeBrF5hB/cJ6
KIXXwh80krzfE1G98gW5EuBPK+2CtgAP6Io9wfVzo9m5GCMHawtYZvRFMXkfHF24JKLCpZJjtDml
UYeD2vKNourkmkqL+gvtgXeZMcBAaWH435qc/Bzy/R32oVfSyYKafmLDHsqYidtkeeklDvib730N
WToV2QQSn/Hbya0SjdZRJpp/fzDFF9kLlZzjiZbyTRQc47RMUK4cbjVjYjvP78oWVvn3MkYeLdOS
2fQzxMggcROT3Y+yxTfyrlPD/oH5DxhxY47Prax4hxCvAIQuT4ozWqZbLILS4xsVo4fBMwfSgXhi
puTq1g14ByHD5tSGp1cWW2DkztCvF3kQAcR30nmC0sJih+HtU/MeyIWhMIJCxsXKyqNexK4xi5LO
4Zp5mxCzR8msNgLsHOuyOoX5vk2vXWq+9zxTWWlkF35uHmxRkS4lcoatGEDVcXuof1+ruk+EVRcc
BjV5FjxAWvcKnEPFhvrIKcaNXGwdRdDlr266HARPgmHhfNjivVaOtwqcPreEpy9SJsUDbdf419oD
GTbBxJQPeFbVaciK1VVxk9IIr+zRspcssOiKhJDapPUQIW+z0N2Lm9ht7NTCjFUD7MoCJQE5BQBj
x3BsPoGpwW4OaU/yb8mPTjhCVc28gCYzq9kT2Swwwnc0ekNXCe5Wpr9eUHh52IyrpKdc/iljaJtW
JjGhxFEvN/xd0yVMGRDRmNnf0MP+OK7sOIj1wcF+S4nMevrQuRe825aLl0o6Gr+TwCTjuYhfigP0
yFY+PbqHEiW36aQtkQZPjsYXbPZqpx4l/w0kks9JLxvI82yIlmHZPvnhgN39UbALL69oyz87bhp/
oeV5Ra3Sw+j8FKRMa0d83pdmHmmkQuoNDJkspAHtxWGORUwB/Wrkq3pBbbjvej49ikV2pWZ36f2S
u9vUAocQhSQoiRTcmK+Yklp3+KECjdh/NzfYIiCiPEe1IDfQhmDET3NceSpWPKTFi12emRV0D/l7
ui3xkp7XG61yZW9DDR/BPCw6fGNu06SaB7xNrWh4HH/mz5q/DKM3Fv5AvMTBP1n2IJc0HE/1ferJ
r7juCTWg8qdW55Yqz2SDXk149gyExnvNIZhkUwbjTBPs2G5GF51Bz0XfQzqxSAN0PtyHlFY7rIEz
aJgxMMFPmdIK7R6hL2fJTbsIHv/eAANm3RyRvSNsYPqwP6CnsnX8lrKwFEgp+ks9URsqvcAfEvnM
6Myh8nzmm5fcDvKbx87SyjDg3YHx+VyiYgEdSD2MslZ4geX5lnNo3wKOIr6t0FcNh5kNMIP57tcf
znhgWuy5Odh8LvQd1QbUwk+hsjRErretlcyhjMzV8t2gDq/FwN9vkj7+HtA364uaFb0fQgUBOZlG
ZrakoUCwe6YDstcXYHt77A0Vzso0HcQUXn/nlvUpb4IILoMpgQSv9MDp+bEA4RtzGDnUs0ngXG83
ASCcL+OsDC0Tont2rYn4X1oHSRkNzBQcN7ETNMkO1lO2qOlPNiOw9tDdQkW1WlFJhRK7GStVkZQm
2N6ryXLaAwMIRrkEXUH54wQbzJlSJpqJXxtgjH2IhrxPvAKhSHMulVbcYP2DQ2GUSKtoNH1yOHye
aubWID8AeTHWgfUuTzhMlToDNcsDoGvgKOGFpzgxlND7sSCxYdi++dX35Kdwe0AJFB7bnpUiymv4
nCTmSoG2COOzPFLylYELh0qhRfHV3HrKvOQbHSDOtIV2KMM13DN3WasFKTVsW8Gqj6uwR3lGTbZO
TUhuKFedm4Rknl5IEtnBZKHEnphjnYPvjtr2K7s/J0eomEqkBJrkINpbi+OHmkH3A0woekARXzUN
dFWl9ij+cwPAyCTHzJtnwFIQ4fxirhqgzfWm+LtnnmfyACQCsPHS3dkR9r555TmNIRNkCe+QteeP
Gvzih+HodvMd/bXD+ahvCK1d9uxPkv/7vhiy+oEsJCBTI88FGGYskAGb75HuDHh561itvdbxk73V
obP1d3j1RIWK5rU3DYGmG62/cW12Cxy732HBNMODVzz/1/JzLwXZ4+coc7Bduf2RaEi2dE7tdW9O
Tllw042cA6tq3l+0ZPCiYl+DX4a1Tk+gy2dLwR97gdlzyhI4ExxJDb/J1hw3lPAx09yFLgHCDWNk
todOEdBl44iE94l98yNxKsHagqJEU/N38TOTfLKUawbje5xHovs1YOKEPktmSHrWli6jcvKx9+3P
6Uylov7HTo2/sZNkTYv0X38NGBYtSSacoKDyOM9BWqoRQA9ZiLf5evvl/AoB/XtWW/qrlVJGmy0A
bCvaoHN/Qfj0kda5kazvebsQWgrRQrPf/V1euvv/10oyD8IauNPh1ws/B6Tb9guuvKO+i1wZxaUl
6MGjo+IsBad0S9ZsyXVoN9iO15ws7yuu5Fz48OKe9b45YUpSkx+MluSbUB0FOVpcSuCdStKz6VZw
JvR7R5hJqwq26whRUCAxY+5ZrF3K9XU+2/4NxWd4QXxHEehIO2lIp+mx+NMyG7gxLRF+H1bMNASl
tvTSygeICEYlrLuVe78n9GJlbZl41Dnv/MMzohmA2nveYCBi7coMKdcBilE6+pzfI/Xcy0qVK2US
yhXDdE5bf8vhiG0Q3nSCV03k3KhGwI7+5Q9wYKIi80N5YrA4uX0PxJHl/7WWeLo7xLuiDJG0MFT/
NS3fGHRV3StPIbDeuqWA5wDOHoIfnuSvUGONYuxskJLbdn6BzhVFEJ3MxRDDNxgq4Jvr1/JX6Raq
jgSIHqlgydA7m/8QhzKyCzy9X7tfnD7gjA0qb9dw1FQnK+tbJSg50EGd8DtwJsw3fn4YwNF2Y6jj
puDUDvxtMHg1ji4K4BQnCvcXxkziJd+t+4szSv1Jk7e4cDWtpdkSua/I+7s1Ul/Mnj1Nb7MgD5fk
jENDADgC5aNzCcrrpqILHABOqGLbaUoK3pW6FxYtV7e375LxyA2TvkamyagXBKxxSKiHRKjqZqfP
gD69GccnIOF/rxfVRexVRxYxKqkYTgdjgFEYtGvmtF78PIZpklv50Y8t0TZEapuLHFP7reO/98ui
jObh0KwPhbFhKUOiuWMCP8FJ/5k2O6AQL1cFTzaJWk24u/AaJBrHoW8Edg/OGXCNQDrnJcIJyrGm
KL0kDkFEBfuhcNclas4KPlao/uUpiRTx4SGKFMlkkd+utCKJ8QZdxtYSCN9CunpGCNrsB/uNQII8
viZeR0egAEJXtLS/APMVx9RVD+Nrnqi5okus6DCGwrQsg3c2ZCLyHs0bIaR1s3vmXknPmEAG+nzv
ouwxWBgimbTzqy1boeIYf1Z+eGCDnlBoE5WX5vT5urgjcfaLSQws5lWKq+rYqeop/0x99G5Nv6EH
eu+GPe6Q8SDvcS1rcfHp+fTFDboqp5Oaz3Mpi1H59yK8qy1JgoOiqwW+0M9Xdyk0eV7Ac9n3SFuv
TAAYPLD10mgR6E+dyvCqq4Jr9vGF93qnsPAsthNqvXPgej947GYcuHKgDFnlRrp68pxQF4aSdnEq
mwDs1wjhidC6uiq9dt1lgLYkRjvVslGcEaqiqqEgqvGVVueiI4BBRhD3hwwk5DfvnCQcRjztTsA2
8Y+IFkFHS0NV+7sNhHhpdSGD7CTRP2YEizf4igCB/zxCz79fXCyH1MC8we8Nydza8+sS3fWOs1oD
IQXHARz6LcSScy38E8HWC2dswApr9NAlCj41Sdoa2cQzO6eT22k+6BHitKnUiwXUQFh7ItnhOCtp
nDsUAsH46IBuGFw5aov9Ix95+eGY2tAMv2VH4k1mV3jxaewtmwvAU9aw1m7iEp8slYj8GVzz1pv6
nTJKojskwnebQXsPd83ioJocNVXfeoPO6THZ2a0HN1lOgCip9G7X1/kxwpK3BfkCHlmK2//MwqfS
uZr6ER7NFSBRfftS09uzA0T+QkCUQsZ4krzcn0hyyOnmX9RBsdEb8KryCZPxlwNq0MBs6naJQDOV
jROL06oGGLL0KyY8uZ+s23OtOzn8PKDH7BQ3uS+SUaHgdIdLDe/Xu2GSyeW56t5gurAc8RjTQFA5
NmJxiqnJd2qASUWj3R28FJ5D4BlH0uQ3wWsGyKBs7oXm5F72P1vGZL2Fi9ps0RBZ3JrNHEuJkMwh
wUS18wm6+7B33Aulg7r909LcuFc2ftzZUhXRnLjDTTbqQAQ5cEKC41b0CWkGC4Q3Ipwzv7PmwOEl
WrwXzqOMccukgptbQN04G6Eu9hC8t4VivyKBz8lSmEJ6YzHFDSfmB2JfzlnU4gUCMnOpNPNIf0u4
8455uRd5Ff65ElRlq1uIpaiOI1J+KlFJ0b2MifLdBbFptEjt5Q3ss0gFeUjdjrLpVqqzBfnKWkkQ
ZfxCIsMH9LbZ31Ozp72t+S58T+AKT/I6b31Ns3cFRhHTvLOwBU32O2StFARLLG/tonsWDlQRfq1t
SkxhWIjLb4745hFLLUKUjm/IkM2Yu0KbBu4zCz7IHFAoktNDk5dm2s3aPATiaTvRCwORBU74Z7h4
YImpIIsrrvmf92g7ePvyjezVw49psJ6KEBB4qDilgY48dePHaJnBSmsdkTUclFF0j+gY2itsUroJ
6Kudzmqq45VfiazZUpJkSDYs88DPwEEdJCQPDSvpnYxSiMiAOZqFbt5vIuY+6MqsQ6Di/AWrG9ZR
1tYjM2Su2xREi79wIMC212AOTo6B5h2xu7x43Y46pyq6RYY7SPA0D4lkJFYF8ZTMtg25O6ANnGtF
2yzAP8gkIL07Q3cUou8lO/E97c0GmifLKC74iTgLK6tp7u62F0uPYL2bGTUJCxDqT67lpqUBDTuV
NDjHon/qGdDUyAF5O3jEObK7HseTvZ7j4jlaIusvmsBEpqeerhUe2Es6ZWWYSNI/y3isNCPzNrxZ
B0H+5dEri2An0qWGv+KRYfxoChyL+1xN5ALtxbX5uLsn9YYw2Gutchb2Wxp5PX3+o/rCtDbdrF2y
d+W9fOVIj4CA7ST2AegH8S1tYWO09ASvRWMRWOYitLmk/faQcnsOFKbf4toMwJom323GmdY3k5HM
wVL9FxToBhyf3Rjg4c0ozOE//aLXp7Y0Dmv8iwxtA2uY/tY715FtxpbUHCruvphUE8fvYPvfibFV
QRIGhc/+0ta4VWCVUa8Bgl+EDPP6gYpaGyR/ZnUzrYVv/U8o5ou8Y47mPZswG9BECTwiN83QwvAg
FzTvJc1kiADjXl+MA9ckCIUZqw4s6IizIF6kH4ti9skDmwsPpvp8wMElReYSO1FklU7Frwp4aPzt
0PTeH3DVfpP+MOb3WneSbez8EWJBHTDU7qo5zmjGy+tFLfzNaXG+6AtQWNoaIjp7C338skrp176G
hWtiMyrAD8uXPtWsBmfC+uJt3YEbYGHWGWoEl0gYxApFBvVXL8nN1HtSjCPP+z2tgxjpAcFMXuUI
cy+kJtLAYyIODbBWLX7YbAiSnO1ZVxhS/0cMt1odyRVJ/Wfd88cKFpBg4epItR5AE3TXwskc8Q7v
oBJ/ykYULhJvFqPR05bLgzRJVJy93rpy3NzMOxlnjg+P5mcrJbHi0t4G15gCeW84S886sAIaMwbd
d60ANZdZ5S2CYz3DHA655kv14WOVTPDXvhABaQ73pNhN5rjSUXiCBwW4iQyL8NBN+I0ieJNXNw1X
XQG3oUAFTqtZ88e6Ib/qu8hz8U2IEt2/+b2fxUNfzM5FBvvfj5XEm1YhsAr0KT/ReA6hn4YQzYa8
Dp7/XWIUsueGZ3jFwHXmH61UcW/Qxps1JLIuKC6P9m9f311VA0EFGmwLOWvMGkSQVgQfWzIyCsHl
VUmSppyo9xujlIjIUxPhomrvi+bClDyiZuyaPSW2ZsSxgM/lFmD9agPm56BqcFdviPng9hfeqCbM
V8kJ49BOy4hRPH0qaDys0gvNUc3WMG7HY1pCotuv1KtX6PtKTdWtBsd8KLiC08T+7p1ZofAuXs7t
FVgrjnAmS8wp4/gUvAKvRfuUBxxA9EYjq7JwzJJCHDOVz+qL6jUXglHVH7YOajsO/yIpkFM2PRUi
mID9uOCl46vRLqBsC4VAbjjAyE2XAFKJPtSHbP7ebZoO+pno9ZPNLVVEbs7VvanMjcRv8GUbAiYZ
CNbqAdUfpaFQxiPosXqm6i2aR0Zsi66asYhkwsYhNdOaRkMcxYdDuy8PgCGJzngynfp5NeouammI
TS2ssVfmAJNwxCyWQWtg4lIKT8FrV8vu+1eF4+4+7c4Uc8COymUFk+PEUFCvFYjcYUJtu/LiCdHo
8lCNAiuuExutinUclfW0Q9Yh7aaMIYkPK+m15F5Vu2GbBzXT486Nob5Km5Pk7u3okX/49IHKlAoC
WRljaTINm/0l8MDQKKJ0uWqgzNDnUztdIx/ac4NmTD8VN7rpT1qTk5rJ9twJivuIVwWCxFh4on/w
W+JaHyBIPJ+TewpM2Tt9mZGt+viCYJ+bd7fPnFiTs6LohsLcbKbC3rzHGZAdZxkwoGUuqvAVlKIX
enlzXw6xrxPNzrco6Vr5YnEwSiiQ5LZ23+Ajt+AjXYvfi7mDkxg54/EtJFiq5ZmincVyh2lzg2E6
HDSO5Mu73L7KTJ/P7KR2bmgUg6jjHrsjyvvJRsFnEaAYP3mTAZqG+l53ghLGrkWaV2HHBTdjSZ4i
/Kb6oga9zE9tjX1GGz11tuB0YP7FZP4X7uOIovLcX5/sPzJrqRJxqbDrjUkFcx7Jngr3KBb4kS4e
Azs6Jtrf2/9Pb/jrOPeYpx38nOa0xUHPLU9NEe2z7Oy8ypBMyGofMqhEGNHVlNuJ9zcV3q/ZPHAc
8xaJpIGiH8mQ76ldoq5RYaio6kBYywyE766A1TzGIs/VVYNns33tZCESbZQfiNL3ueFzjVVQMC9/
aUjva9dP8oRFstMkZVNzU1rlBPLPxwqCAGsSmkrTu+2aECBkW21+D2AdAVJCw5VJyRFxM7foCem1
fE9OOgqaxp3aPENYNPcWHIH3SMTfGih8VcQuyAoR2TIbL6iwY4aQeZrOfr9yp+2sKojDypJMCSTM
0hP02rFCsFZ2TM44MNhVMetj2SdaUfr2PEz3nD0ah096K4SAwaZmzU4WQlhE996UgcsFXuYxyA3s
Cq9x81E9Du4J8WTsA+jRQcoGTQUU/BtgSzKVHRx3mpOvJhzUJ4H4naKIgPCW9vtSinMB98iZGbzr
j1LUp+azp5yhhhgbd6OnSGeKbe8w6TWwUoTNQNHp8cIb8rXGL3De9QecBJT3pyByIBe+EkxY1Omo
effsIfB+aaGoCyO+CJXcBktcECECTb8ErddtnLHtui+T7q5soksunW0tX/0md7Tu8PTb5MlinFzZ
m/8qik+UcbWgxDwbMupm+GgjYG4b7f0EJkP3E/YuIWCL3bYw0LmiweSgrRu5iNz+c4UGImKMuev/
4VTIc2EwDZaLOLhXzoxG1vR+7R56PpCtdBBWmrtJhpk/Ef3LN9X4NSuiTmI+SK4298w4CJMaMGcA
eTIl1RbwevhieVnF8JU26ceJfGOvuyPom69vJuN87SnozHYsNHwFJAeki2hKWAbeqnKy9zWNGAjs
CIXcTZotrmSFLMFDwuCMDZs5In4YOR+phIFy3X31krGos29u78/8Kt+UkAQkGVN8XrRVEuULzYxg
LbuZrsY1+DxJQMdRn+RlHRfY3tYut7Vew9aJFDsGCnw/HJdeQ7TQhN5MJhafcHmTkFlFWGgfZeEU
05WCHI/ZvU9jv1XfLQSYKe6aCTNGKtVJh9ihlC2NpZZhZ+YIEYsCYD3gOARHCeRcL2h5i9eBMXKP
sevz+fSHNypVlUdIssBrRcDcsHSf8xEDedfpF2obWxgyhGrYvJn74AmzsjsxPCu0RxTsBKvXbMSl
AaILuVOEm1WmHoshdz2hsirfIinyvvvmvHpf7TbWW0rIvdqw2L2jD6sCOYiawlwj/W/O5lfUZU9D
g3iSwg17P8JLCJbQxF0l1cYAUoS1R/tSY5kKySreD8xlVrPoKUecv9mTmsteA1LZAhuV0eWlu5Ja
GnSTKVt5mLohns3lrUDCUPgteQrMtzWNP7aqyoQ/q0av4brW9PgW0pWIXvZfvJ9isHhgrRJxJtcY
zqqt3maRxSutzpdYsI/8xR0k3TgjgEekw4gCJPWOtUx6+nTsW/oeKZ3wZhuUx9/auA4+pkj0If0I
mjvjYEnPCw5VzHz3nDkWuR9T7znDoaF4oeMIkFhFAnbojElpFuyx2ZQgPvEMQ5X/mym59MFzh0th
eiBxI+q8hDaJUYBge1lESmyzMXCZNsTCNYlrtfQ13eZx9irV0U+m3Zb1Sh7mQK0zygcDQLCmA4MN
eSzGc+LNYUj1Djm1av5Js1z/6txQAgHeAIGeJraB4ZHQnu6F+3XjuwAPG3rvKcLFyPfjwgxIlWWx
uHCUatLRbIWJJMtvCmCY0wmUY0ZA0GUxX+FrZHp6TERiep2LD/s8R9/GO+Z0GeGaTuAzx4EeuhJc
/v8lqu+Ut3A0abLSN6MfVq+qTlib1z0thPZZLzJ1he2DlrBpmM0V4XOoFG2cNpZ/BqlooPc322Ic
FygGptEBqyjH56+XX4EArJryfsNvXu410GlB2rM5KZguaWJw2IrqtTGq3HRVnMZJJOIwINtS66x3
wvhwGARfcSVHPpH+GuQMH9nSTVpCBzi1mCGZ0OP6gvvSZZB6T8F0TTXhlYhGkshmRECw5yMgZamZ
Lqri2R+m6sRadh9E1gcr4Q/vGhd5squBSvfCZr9/2MetYIoRnxEc14NJuJnY+AJCtzNedupSsks7
748Uj3r2D7WX8s6uP9vvPd3NaWEgznF2kDGLWpvQriK0kmFqfRnc73d9ftww6mCNWoosD98KVUcB
DB0u5xxCzfOBPZyxJ5no8Wv0A9Y4CzqGqrqWt9VmUzP1kcNLiCawLHF0B9oN+q2wAHgtMO3+dmoJ
CcZfUUwn4V+FjBpVBdrbo83npXkKXtKQRf7CrkXBgYe19y9Nc3gFO4JWiLpa78bIBFvoT5lPjncj
giXh57IGih9MfwxXB6f9tBb3z8LcJVNpX4DHOTc+HsWInIFElA6D6KZfsluhsT/94cik2d27J/kT
AZySP2Csf5ilqqipqGQmsEbVWcTuZtkmnd+1zCHzQUUvYcX+kfrT+nnAbZZ6Nnh0EDq8i1vtZiAT
9l5JE0lIl3yPgZBldEMvhqg3VbnebmkUh7sbdbIhKqW7DB24CAh1Ga2FYTIPBMUWOZxiDZm9rwC3
00PxO+smlmMGis2FrccAMmbgbvcdDHaUv82LLw1wq8GxDtYH92Ea2R1BEAYDiuOnfGS89QAEqr3W
xnu7WaaoF7bvd0id+qZEYqo1CPebrRENMD/C9keI5ZXdzHKqBOt9q6C3g8uGHCN5sjiFWoNtYKbE
GTFqDUKu315h5OCPFrlKVaqDI8u76TxHglqpgoc9qW++x/pt0nMd4NAoFW3hQWhE+DAVo1Vpcl4z
ttnOCGHbgTdztjTA7/ikxTwUERkGaOU/LjAcnWBDfMZuNTY3upvAehSm8gole5G8vOBwR5OPTOLa
Sly9mmwG2LHy0IVeRfoCnUva72odsscerZg8oE7GZzR7nQMZyKIJUHGnMF92pKUIP/8lHcJd/lro
Kq/9/8RihuzWT9pIlR8Y6wWMfORQWuwDg7a1hoo8A8BXb7snqYttF/k6bzFEf1arJrVAaK9aVxH5
chgrhZ4AMbqUpVlSdrjJg0GBeQpw6FshaP1BOULDdw9/x4x8kGaAeYfUIxis6mFJH2atOdPUUxSu
i/hHyTDriTXzZDpKEa3Lc1KYb2YV/ZvNRegQ78LYh52WgFc9gw4P19eGK85Nkb+kclYsxAE92k/I
u+8SyibXlfdxY+uyT2VHhIEQhnmj/OfUSl1B/1zkEJhI2RIiHKoroNTLrqANZgWchhYtO2l6XDE0
1p8OqU47fS9llFooMaWIl0GEFdNhE05Kqpng1QJhe2k5PbdKc0K0Vj2jctB+VsqF5iBW8b57VV/3
qs2k0dMp7MTegZy0To+z8Qf6oJqFDnW4Kj/KdvG3r9BBjgVOowezXJLMNYlY7akDPXjxGtnCDggn
DU7iMGULGdvd6ZCswTcEmmWZxwMNKNfTPGMRj35i8lfHUySrKOYAZbPkiDykMEFW+i6ABNSvndC/
cHQPS9I8Q/tzed48bFxN+afNjO5MbsM1l2L+nOB/H3AsrrbRJsh5no/Wl4sEaHxwHM8+gw5oNO7p
8eI0BWnxVAJzMzs491gL8E6v44z4jUlSd4pv7Jp5IYMUivcP7WnRJBpeFTH2Fj2+FfLSvrDSDRgB
V+sBqQu+UBLjk1SGfPa+PkK63XjTG3/vga3LG3wLcVunag+GAHCBtiiMFGZqWzP5lBhATGgDRCqz
I2GMMGnURDr/1ufCmH0zfD5smYBFnvEu0CKrzm2A0LmGZTyOwo1vyib/9X5YXiQMKgnqG4snmvYR
wJbNlVRTCD5rDe92IpGuot3IrfPKWVwgw2KoTgvcrZAMxpAl0d1i9oriOyvG77nSR1RH83sEuTBF
50TVF8UG1YOkYlNWjdhX7w6s7y4HZn1h8ASnS91oqupIp96THGwB/gmb7KEQOzECC4Wz34k/mqJP
kUW3NRD+Rpaa12USp+lPBnryHBR9r33TayJvU/jw1jTfqbRKi4s+YzZmYbUxuiKxnjDexY30QKz6
ZOaNUgwKFDwWVH1tIfU0q3RaeUpgMwiX9Pbf4i3Yg9ph4NQkHOjV7JCF9l0W4kv8KXGhXxbCww4I
uA+d6WYw0YcCHIbiQ/yj+1WHjo/9XhGJIx9FFdZ8FkHgqhCwvOePbZsAXdRhEs4vD00lis9avHe4
BDa9DDLzNyS8ORjFsAgEWRrawm3VWRDC2sZqKyKLHHqC7w58bJmOACyfu4ZRogb2Myvntn3URsU4
kXPM7WSU1RQqOV/Cf6Jl9fkZrlpC/ipVU29LZoYUPrDbajwqJ4oUjMW2mMuGL1+VcfRjHP6i98yc
ptJGsB6EHjRE5N+h+WW5EHfJE0f2Jgb8ONzEUtL3PsvA0Rgxxt+gJiG/NIYHRORd6Q02Qo+94n8T
stI29b7twIOdlW8pGVjpBiXGylTWMFioekfZD9Oz2rA8s+Xwp5o6UhEMTFE5WlVze/o033V8P8ee
87kYPHB9BcE6nCPvqzKl/zvqcSWEMo0d8SI5skrofLvKacWsyQG/t2htXmxiGDwhq1irGfjt1B3/
ZUK2XSmEkadjHFHPk7DY+oGZocAkIYh7sAV8WUhh5/sX8PcMJbaHHJXqx+G9VxpaFyAlvvT9wC5I
TsozyGg0wRTLRkHUZDBEsMCaSZL7K1CocR0tzfzTVRFGxTSNWSzpNeEjrl7kRrOLLlU15ly2HNOW
EX/6MyC0UC4GeaF7Iiy23gjk/MZF+wX153q5F8OihtZNzErFtRdtYWF5stT2gQ+rFoVcBDTriHke
On3yoK9xiT36G65Id144rg204wRoJZ6pDsshtY7T93s2c0NWGo542dTeGqtActKXwOFqdTquCEtJ
Gluqwugjkt12lNZYNqXugPtgK8h4O6ccMEdH1YHv9fpEoI1W3myeYwK2pWiCxAZ4zKPxLFnLYjRR
MDdwKT/dCzk/1TuyWsw23/7f0pJ7+6LJtiILe5JVp5I3YOhiZEBXb1vDOKNsG5LB/+m05ojRqlAO
YlxSvoWBoFmM84BfZPDHR1YNM89OFp6ER1GlfYo310TDbWPJpy7RFL0q26ukZFQ0lrBrxzKvWug4
t6qR6FguSHin2VkQ2X3BBf7cANzi54muuyJLmAy2ZTHGTHNarRfOoSCXevq1Ey7vCAQYda/p7Hu+
7/xxhUnT/7S1f6utfPgb/dFwjpHT5WZ1KtXMvdzvXPGjukW0IoaIVUfNeAl5DEe9g7jk9YrpG5aE
YErFLNU4EUsOceuVgeNGBb5nojOw6sktMP6iGah7tpfUEaSVe97AtKWYSXB5f1kRRCyD9Mm7wt8j
Cq1/d2zi+/joazmGv9ODHooJCGBzD084CvpjKay9P9ffjlX9RcoiG58nsZDzFnNnMy3G3G8qsYn6
ricsZzA4jB3s9iMWLCRELoDSzYCeIVSgGQ6PPzMlPh+IB7SWPoF5NwVtxvwKyv3g1eCIr/r2J5Dy
Cja5UM0iLipBNTbSzERXOJwWig6V0U7GoCfLYtTRPnAeW4J+qU/h2pv4fpiioGpGSCCeMsxy/JHf
OWNlpFbe3PRtsyZrzuZpnE15G+SA89Krj8tcfRhXED/LK2muj9I+i9svsYlu86dAGaV/TEdwbZoN
RNVXMi1ssFeOW/6nk5otbB64tqTC04RMFEcQNOMO341LpkVyXuA4rF0rU81kxdjcwRIPgci30tsh
Ufn0F6a9u0VbuqclzgdIfVdW0GLeKpYFFZep3G3OoRWl6yB8diasSdWl32BXh0/6EYA0mS5lf5Bu
BtH9sCWVOEo+ALGqwULOZj362p+6gGz+WOzHwQAmLYQ8EcWzPkQ2VZXMG5LSzQ8sdex8vKmB6E2x
VbdFnU4AoAT6KJhiS3p+VVSFr01ra+BGLZzTbYKmTDkGirF1DZCZ7MxAiH72oBNscnDpoHA9Z0+q
HKv1QRbiEajddB4Qp1gm5BaxkVlRvWRemHVrwFHNWD9/YGuJD/xN5BUWVLq63nFrzzD9r5V/tMk7
Q60oUOnpI5WjbkfI011fpAtWdfilccai/ok2j4cuUclC+/2+bTHu2+1yQ1zSA4oPQEhh+e18ASA6
ZiEAR6P/gcf4nwv3M9oYOrMeNEPrtwQtdDa0Z77X0/azkCxPvi+pX45xXi7FWTKWmkkCGXL62pU1
FAY6JAoSfFxGHzfna0A1JWyaDKKG2gZAcWbPmfST2/phb0tUQsvwiqOeJEsIL59wjtZy3+OXCGQA
5Ck/kBX69sl0hVPV3h2uBFXc2STaaKLmTgzDT5ZzI1SKwYIi0DU6NgRH2D6ZOysZn/2rjgKMCqVT
xlcFsgaDttM9ikINAVS3r0b8lL+JBtI9BhpKVPA7JyPCMLRU0NG6NQa/VC5X8JTtpm6b7Apymkg1
tlg/la5OZiTficXtgMaZ6j7gvJWpqRj8+KpxJJz2s/Vyb7HALYoAlD5g2i8EH/wVyq2KgFukrBPZ
baiTN8TkHspP5+YXd/npfXO+2gMrIvPBTGfIJBqpyTdNWM32QVDkrBdJsPti03HLqqQSfcOWyYuh
kgXF4Y2HqW0LWfNeI99tSr58UeH1n5dNTe5TqFzq2tjtFa6QwRmN6AGoyoSEwHeWl/KLF1qJF+dq
16nK8cl8JTC0tiJDmblFXtegeXW64l7FpKOgdU5ECi7rBopB7xfe/AISDkNOwPWVs6ScOFLsKVxB
HwSvttcW5mGKREUCk6haoGf+6kbykkXTF7oanhLNE9bOQj+LxH+b7yiS/3ts+rIYRF0prQHXNP/K
AH97bUgbmIAcZqLcVuGezGZgLtDeJMkIeX7RIEsCG5uu3piNJqzH86MYR0IV10Bq4EfgtHLoo7If
9fdbpt4t/ZIF3TeFYiMMbIw9Y81Us4E/Un4jPx1a9vnLRrL1E5BbNIWkDh1RjTLBYTVfUk48NEOf
ahGwn/zYHQ0fLCak0khCahSH1TAb/ijMHo13C7Sx2to4zjR+UobaPPrh8/eXVU+be+An8xgEpv+a
3lB8tjbtnmQW0iVZiahUH8Te+4jZY9+P3yIAlQSOKsgOdr6fCTCUHDpBhLo7Yp1G7eche9ALMjT3
kHRMPymVPe7KIFd7b3bPAW/OamtRJpKlUBX+QWGa5eera+pej1ZMhEPgSs5dPRIK6MbVg1BzRrk8
6YMe8Yx9srQcYoxE1VZTBsuM/b0IRpg/IOsawQ/luOiLsOC7eWENtJ7zL7h1NoyxyMYrrkMn12C/
EdRjqwPClhaWPuJhVqFd+riyC4J35qLnrnvWgTGPJaMM0RtIRF+KVkbziJ7gq2FeEsjSPgFEos3h
uoIneBkVNuaGCa1oDZw+hDCub3s1IdGewBOtIpAH9cW+mIeGaq0XpyfwtapltBuGq+do5RPtAWV+
p1v+phlIxDfAE432CKDKJ5h0ljIziqzza70BmXSiCj9l3Nrbjgc9Bit/0dBQpqGcF00bBX0C0FWv
3rH0euheO0Vw3LsFLzyk9vZgdKUiDa63bacgUmBOannuAaGXX2+0PkbiAvkC0IXbelA9/i90pn2g
Ke2B0RRQxSUtEi+WqML3Cwag+o+Vtd+ehFd/2xMApPBvvqyRMhm3wGoQ0T7SWWd4lIEyUmX1ltVR
NkcG3QT+TTLzVhARB+3DYQP9OZ4N9eJiv4oUJ4/DYCP79p2VJLxsxo2Ocmn4YMIgBHB4szbk9oPt
mzKDEWN0e/AB4Rmo9Al52mxnpmTFc/7tFxf3arciUqSJPBaQDapDYsPsXNngyxGOy1dMkUaRVZmU
LZR0arR7IHPvKkGAc3m0FvyhdRhyPnPOJk0PZbxYegY1fu7bWt3tU7aPAa4S6u5ypKv6AewDBMmd
fsvJ2IT0z3zBsAcIgfTf1/WQgJr4BecYjLNXJQzB+Ic6pR4HJ5zGpqvvWjO0AxLhEUvwpcSNA76i
0MEtOXTeltac3Ild2uZrpcm9ubMQLy1a3Wg38ldbtfgCFPg/Mt5gDz1rnxWqgmS0p0uDgyJU3xRQ
iryuGDbZ6aDrjodWeRUR8x0cS3kcotzPSQ6NEZ8R/bhcEnghK20wAFUCQ/UkusY0fmRHdR3EvluC
dhueI+oue5Y945u3hlc5gzOu0HankVQbR6m6Bty+ER9UkW9AWdfJ6jHvFM01BLIcIU+/9vJmH2iD
jL3BoZGS1Z5nglwNKaTuGaCZodHMULu2GUy6iDHW8vGWdh6QFR/qQEWX347/DEJV2gm4EG2SZH28
Ns1pJPe9xJPFWPDSnLrpYJHVli9PiRRnyVFDz8ajir0UsxMm/KaDX9Rj9tNfoYI2KEVekBeXi3T9
dr9xUyHbjkEjqhvV0sDvzdsQJPjXzSZPYHR2R7pZIf9/HF2GF56DCMdZXeHrMkyLtejsyPJ5kipy
SCUQEInN3yuob2wOGndUO9z2xCPD/r4axvtV/xIek3TUcJUdFXrDsdF0wgiCCNDlGMhM03W9EFtV
VNbJ49bWpYcImaSDl7pnJQGN6HccZxmziE+dGyU7LBlmKjjPEbAlbYHpaxXi9GhdPFnNumb+cdmD
HTCuMcKj4ACSoaZx394zeTfn0tN5bWfCFSgAkA795q4noP7neSLJenwe6NgST6dDPMsiHIACC52b
4H7BEgf3v51I/Kn7WZTwarOsGnRU2KckBXyJgXz5SOG/FKNa74CDGMOGv+jny0t9pvsBzk5ydZql
Q2UUmny7sXLcMDW4+rTPNcCzPDpnqZWEAmiTvcd6WMCIBQE+UiCWAFWdVXXdqjHdUpmNZGW/CpPf
IgLwlveR1vQhbjw15HispzxE+UBFPmAoHYOlchjcp9uJFzpD3aLIYVz1fBqAQds/1rCNt++iJe/X
XCio1tYkk9g9ezmhx1186yUugCiqYbMFsdiacycUNRUeRXwGJ85ILr9+wDH2DNwRanezqWkHKOU8
xRGTYZr6wZoCeb3ZmC89jjEDIXGTkCbWOWb0PVwPwl+44g0W1epLkdH3/vWX27PcygUrM5ayj8dr
wogMmuTQfJvQ9QzOFoB1Zd0YAEkRtdGVxyRm+bchPoVsgbr7LGdRZtNIHAWADRqKat4YJNYOEqxM
kj8Ne4cxNUqCB5qI9WK1nhGGESRimV7eRQJjIH+uPZaZVTH+QxWVKNP69CC374DSMzLL9YYeRjrd
+EHrpFZ3OM7lFUB7yxsxvke8Uo+g8WQl6CmONr4dUyKQyO+CLKn89xpUdyIHVTxsHxxiuzIyn1qd
sxZFPv3Ybr8ioi0HJLFPPwWrRzOJ9upRMJ2V89M6Q7RHxoDVfGC82flOlJl6qyHagA5N2WKBfFc8
KcV5yS4i1VvENqiQ976n0RPrwVhdGqXGVRZuD3ND+EVD+VZcSQddiD3zT8bGpFPPzkkLCokkJK7G
Av8qQHrFfG6f2pRlFUjUJ2MwSLnrSrmAEuCZMMih1m9Ve+AuVAzRb3roMGIXzrc+Iw6P5B6KICHr
7cjAlsXkt6GaXwPMaGHFTI5BOYAQNpbYPi9GeyoC3dD3JvTJnJHUh9f/s08/f1/xrZKmMBR0VGtx
VUe6VMcHkmX5NEHwmnAI9hM9E0gEHYrKBzlVCdUSCvil5IxxD16/9VPhU1fsErtyt/dgE5qTq4hw
lRodDCjcXRpFNd9FvgD7syD5E7vZzrdWlGloDlF98Cd9l6axH62oGyJQJ9HFQ+up6qJlc/2EVoh/
0OWWkl287oS68jBVYQq/fGAHZpv6051x11UPuFbBVDJgl2+oGBJ2znVD/ffx7vgwyI6xHKxf9gth
WwPKZTcRT2ClknNzij/PacR3gzp4ym9/poCoddQCfpaa76C4ghqZXPb/dSOGXhdy/0QtsvDpW7yK
/s6Hytq/xQNcf5DUN7DweFWRQjKEOkcYxIA47CdyOqG4N4s7aFjviSY9Ubj3wEgOUbfKfer3KMvT
931gi5+y6jeJqilRkIRkTX5Yf0QTw9CAqyrlQKods8QX8rQHqeGU3s47ZDbSUIYQmYKL3AtvGP86
J+ATNMLBeKgH2gU4jHP9poX83847vmjs+MNMV/dX0ZAy5b5oHwJE9Oe0VmNSAqYLpdShxGN6XCJp
mT4e31jOGvW2SuREAM98KQ0iQ8xzeiIdG61ql3rz019Zz7emI1IyJFOIrL7fxvwIG1y3BWqpOFKi
/wHpQLqAwNyys4IdoKEXInaL5dJ7gIGJGFoomqG6nzOQWMbWxmTMrosineujplVSsPNBD7RW2UD0
wd2vRkeAkzeIF5pAEVSDLpCzFdpjVssnDj9t1j1Qp+nALXcIgAUuQ1C/1OSsn527TcZVoYXOVJsO
/VjIvhZ3wZXX7Hz1n8gkcrg9bqKDAz22pdz6dZVaZUrQw3Oefjz7nq0huV+IjfmJ4eCbLwcGiHFU
8QJP3Jx43XDnRWZqfYkaI09roStCk3e9dS1/2rqsEFa1sUaa6sVE4Acoc6nV/YwKpMm5Tzjsgi6N
jFpPFVLHMvb/LnJkdmebuRO2xEyEwPnBzXQqu3cyl7MiQxlLA4ouY4jgaVVIlNf3mIaM5M8V+sbj
APjwAr93oqSexYpan5wLAxvczlXqRvErYJ/uhEYd6OLDPvw1baOJdyRr44eTNmXJ8BHzEHtU1aEP
CXyOz0yjmKgwiuuvc5XLI0d3z4bjU1rgDr3ehGOvh4MzwWlJfjT4mg6yfbzsmdpouK29A9ibdnXa
6XQaJirKwmWP1v0DIlZx2JTs4ov2Q6QDP+us+1KCOEuiYBIBAt91+arJ6MlzAXCH9iJ0W+QpZLts
3dXA5u8hnliuC4i8B4+A52AH4iSZaanqJd+fZ/pIzCbWsBlXGyH6nw2RE5Ho0/cgJKm/mAwpseG7
lQYAiUOlXmVlXMcZO2Gt2iCr807T7HjLni7kcNUqVZZs986gK+Q1oBA89sMJ/V4bEJf9hPzcpicF
5XIKbEglIV1h/2ryJvZiDERJdZt3VBah9b+GTDkOJ9CJ9MIFUvM6pA6wrF7PHX9w8ZYyAPDZwiE2
8rMJyKjLGX7lMPsNsg6m7G0k696GFrKiX3lpFsiWn8QZkcBhswJjN1rob8rNvaSZ30U6sDzGJMIw
egeB57RIe4KrqsC6/A1j3ZThToaXjzpEmnBTj1hc+X4ngYPd8biqiI31UMqz825+ipDz1i1GkDhv
8SKzL/PwDEQuXsVZ4J1CKKZys/wIAwwTWlUXY6Y3uRLVDZvnuo/pNFSx4npSg41SNXuUlIL5aSRP
lOoDFc0Dw30AfFfngf/DmfgqXCaVZXzVlm5/Uy8R00TfMmuVx3rfP1jFQbgYETZ8V6xyjWo0FSa1
hd1aSGvXSQjbF75qZXoiJVeaxSppwncvKVTLQD6Cxr8ljKtutlV0hIoUIXpwtG4jiHbzoZjdxO2Y
P9nJAntA83k9GPyafATiRGaavhqn/aaWOFN5m99COnAZxGRZJf8jXF0a6QYPpN+QFwLHN2Ac+VKr
xVpPqOzbt4VHOKVb6LJ1SVmf5z7ouHQsHIDxjObe/r6/jylS2P7sNSFchhh2azkWohMn/x+iKnOh
J0zxOKQRVQFRe/t32t2S7RcqeDsovp28El6bXFnChroXxzdCFHMTtKir8Whh2GtWcQw9hu/5i+iA
q/NQTllGxs37PmB7yBrO238RRMw2MENhdFBbucyKbLOkSMM34EugxfkCrL5RFYh2FflmkTpIzTW3
I1rl/wkLW57PyHWb/EU7XctJj9ka47R/lXFnPqidTkFM532T5jQsvQd/5X9pl3yIVnzE0q0ZgqOW
SONawYxnk+DohSUUGc3LvvjqXxOMc7LDQrajKSgY7cI23wmz2/oHKdaapQeCMYBvsp2MjiT0Fh+0
GhgCWnsBCPx3BTEX2fQfdrOXpux5byxmZIWpRJ8EtlMwCsijkGXD+tlQcA0icN88BsIN+6BSKF9z
E4y4JM1cIAfZt+OwEQx80l5JZN8/w3tBInPLYmqnT/Kp9z09jnumn9npv/oYs4CDAovpKgSTPT2d
eN93HDOaOVaS9F8OZukxYg+EPTmWWQbRJ92fz7NAGmri2uz569q5pcOJ/IZasdWqbg6al6vX3rYd
fR0zFsfpvRmtNK7q9EvhjmEW5zO/ZCd7RFCAC2wBT8OpyzLLvWnN0zEr4832WDvbG0KxvrAy9hjp
/aU69+M2Hq0ebFNRQOwmisrjQrpA89FqWpmc2XTzqipgWZbGGRF0ep0jS8+du14BhawIKtiydDJ1
Xc+cP7AG+2sexKKnpSMCrZk8s4ZoS3J2OcO/d0EvF7tofB2Vg3nR3uQAIhJh4LGQoqurl27Z/znf
QyA0XqSSc6q3ZjSELiOqz7O7c0iYN8Vch2fHJScYVyi5UEN55d2e8KCnVecJ2lq4LAi8KfMTVXb+
QwP0/JXcSbuNdlrjiKWyB/I6W1NXHBtrXxt1yMYAuqNzaF4f62W6LjwcPtav/LS74Rbea4e5GuGL
pOaSulkug26DKxBZwiAhzhwxUf4RAC2DhxkNmV+pK6DvH9Q+wDBYFD9Bf3AX54Vcb9JZYJMbKsPy
PHg2VLck/O5On31gEGCY0Ku5R2tXrOXi1dbwsB96RegNVa28jIDDzjeJdGMJ6ECp4pLd66BY+EKz
eMIOb1sEsZQ3PE4TWKcZhOZYuIHPsHNkw5j6wjHKQW87+9RN1fuKK22fQWOdD9jqF6sNNE97zQZQ
IgvQm3Cyr3i0xOjsOiGVA6JxTxd1712EM5wBGW18Yh+CezsmVqkpHfO+ySv4UpNwmxWk0/iNthHv
2oaN9KedcVObkRTX2EYLatJ7ZoxZd+aSg85A2AIuyqr4OG++jYQrjCLHMZDGtFF3CoNeWw118Ck6
TIQA4Tf+FMh4xCSBoVDUTnvfNx9VvHxeN9y9Iri+1q2ba9/wxMv34QsSzWKYHR0Eofwza2Obx76C
GRiQ+mdKLLYQMj4TVttc9s5Ddgo8RonvW5G9dSc7HD9do267HR3o7+f4krvtZ8j2O6uF/rfW7n7J
/W0nHMTvdJ/BEZ74Tc44vDLjJudV8QNsyLbu8YNOCRrLV5imm7PKiwvVgroMZ0q2NU514T7mcNOn
spx3xGgwfXkQVhUyxw6gAsCqXNLgpZ9S2grftlsj+olFt33eSRKMEQKG2Y5MePoTbabDtip4H9Ix
jGwrYe3JC5SpSSn2XfQ2z/FLVAmTFTGYBw1c4fhYdaTq9jPaaV9HXxvtuy1sTtBpbsUN3UeIc/4Q
4vgYyjI/f81ayoBOoUNJtYHmCcvQDNc5L3zB6v2ThtF9LqOPf6YpfisJWR3XjHpo+1CWXYtQiLY9
qbtfG5cbCziimsTtxwj2Tefec05mApicUIJ0QVBXKHZvBN7AP9cOSEkIZ4hnb06V4G7aeaBeA/d7
3bD2hJD96gc3Nb0e6H1XjbilIFnPdFe+8p/g92i6FKAyaXLRb9V153E6hzxu9PGz6ZsXER9Ib2wU
maUXsYwQGeyt5DTkKj+L30Lsupl8m5Emz6MBvFfwhakb66YgSTVFoURYA4X5J/U+YJqX60HTYgDw
dgdLqY/bs+kez0+UphLRrrsULcSqAnQRg/i6EgBY5SYORWaVa5reDye7t3a2TEbI9lH08Jk8FBGR
hfNNansdpN926BhuTxLWt4DAlDS2saP6EqwDsCr6xa4AHduj7AN2K6FcDPQoWTXIjIQ/gDx7Y5j6
Vtl5zvFbbplWt2Su+/NgQBjYemVfKywBv5DWnaNymN40sfs6Nprb3WMpme5znjzMZKdUgL+fOLNd
e0mz2XVMksKmwQr/hsr20xNF2+/Wfre+7k4wEjv9WkezfiniPUWhZh+WY8Yw/c/y6PDUenDlvJpo
7NU4rVSF1BA9eVRtOA+M5SwOlNAqY9Qp8O2esAwX0/hOJGKYz8ndFoW5yG4SqB3kK/7/jRnva7DN
vVcFea/l+UabT3MBuRqBHiSOAtrj5cAZ1mUJA5MbHZLUR0fX5QE8r2IXD6Dk0xdUQwZa5sKp2uGl
bSjA7bLGLrhUOGypezkkTuxpZYb1IUeI5ZHnM6gq4GVxZvQSDetyfljvOVK5bHCCmP7nxpI60JvX
RyPZJgTXEk+8afSN4yGI7Uwx59LlGnPbOAxoNb8mSPR4Zy250wFGgUV7qi7fhUkU7mLCWD3BTuO8
fQbyrgEVQQuwU9cdYlSE8CQNkmo+cCrgA1+JzyiSFTPurXamIrm+EWe9Yok32hKqi6wG9ts9dvkV
jKCvEb8LfhCWb1uKUUOtn83RFdT8cc/p7nIOvLcAMZ3HR6RHM6c0/q7rFnJfkVErXBtOFvAI/NyO
CGLiyIiTRW+UfMAWOp84lOxF7fNl1AISNzC4eUf/4uFOnd8j/jubjv+aoaVuDRRi0RkwbVnrE/y8
ik5rM5LzylyPpPtodrt0owM13C2Y85X9ch53mluo/hySx9abdCtQqTSOjXKy+I+xg7uUXnlMma3I
dLXQJguNkMlPAz0G2zF+GGkZpIHjyVGQy0XVvm7dnTSoP+PnqAlv8UWD6BVsQu9TE6aJawQXlRDD
MgWAIZXmcYYKrt7oZXesiFLjUyNzely71vQvTdphNokfTZ7A8i01HSAaxyTOJZ2ONnYx0ex0xaT5
GYKBOiddbM88OTe4OG+hidzLsFzTeoJUiyYWztwm1BmQSIPdLZU+ch4FWS7dQ7ZtL8rIhi7N9NcN
PhwX76eIwJauOlkrFm13Typnnr9au1UJ3utDY71x/t8OTu8h2yykgL9WuVwKzR415Xph76nx9paw
bzHdeba/cCUtmk5eCqppmi80tSzdP0BwXMsW9INIfPqXa/Bq4Mqxf3siJ19qvt+rb9Cb4QSLt39d
DGOqAiwYx76oI8gV2wtF2Mm9R2s6VQLGfotxG4Z/HXQzad5qFhcv2sWH3GDKq7EtFo1kH/5GXJPu
SpvpJLDeNkeSZjuIpYFdX9InVYIjHRZJ95KKErAdHb1UyckUUbJvGPmy9U7ikYdiq/OGsTNPv4Gg
hIM38O8HPyzOKTvKMJcJ2L78P3+4UYsbzUg9KRW5pxkIhQp0Wm7tsVzTptfnEObRBDtzsxmHIXqF
nrRG6OvfZ6RQqn36cvuoTi7M4EZWoLhkcDYQmkbjI6FmeYqDsbBr1DN/bEdgpwioWHKZru+bIKX7
uGmcIWP+OMTx2O0/CJS0+tpSAikV/CFe2yDyV0FzasaGzwaODynoA8ZR1giotgeODVAT/ukkvbig
GmrQsrQUvrpNjCM28rrPBnUrZtYYE+thvY1ehKzdN3w1Yo0gD3F7LOgEHjCpOLt+Y+68KTtY3obj
Cu6YH8mwOA+KXiLcIvQUD/Uu2lZKBzGL+EU3BEuGOA8jZmaLRdAKOjuuiFIxrenExXUjArlNPWYr
YRdEzyAT3wNtki6R82fROYDc7Me1MU+Qu/bExJmLiMuesZEgbqK2IS8vD2qaLvkUYZrWj25Ndifu
akKBu2t7A4w3syiuj1o2OSmcaWJbe2bR5PR137UwMzNR5ikS0zGBG/zC8GVdYw/ieX6eux/ld7+x
uN8zjYohsBnKBoaljoHFruvePiFT4tAVwda+ixRTOS2LK3I1y8RJryWtiWDh05mIUKA92eqku9Vk
wheuuhKvyss1HDlLe68/RxQn4zLW290dXJ1IX2bNvJg5QryUlRD7i5Te8/pC1yrFHnabdDH838p+
eAGGHvlIC7L7maKXdQeXAWj+Pj/AYEJzuWpOlvLhYunE4AwQ6SRmHHGkRGkvYGL4bni3RckkFBu9
D/ipWjd+uhoiQeLi1Qyi3+//f2/nHm904Y078M49ofnMXpAWOgP50XDJEmt25AIiboesCxywEqAm
vZw8eC0QYznGu3q8YJK8S5YLdkeahOPyCy4Uy490s2saGtI9HWx0ggSzT7i/OKaW5WpNpoNDpVdi
sI4nYYdByazqW4RUUDEA4udIZ+oYwOjsJRsGoCqSRdeqoYwnMlS1ECagY5XARfPCAE5X5AxWcf85
yBgNWmVLQ47pZh6j0upVpAjIVcouwdk8H17oQnIGDbEtrqk0LXODQ3BAMQZpx92VR8j99Rv7wE16
q7HD/AOvn4y+9D6LD/4VdLzIoQuppc+mspWWMvXt0RVollGw1Kw3Lw/hPlD1MeunN5KB8dK7c6fv
Z5XhuqFLlBlT8WBbW2RaR/vCdEHND9A/mee8LvF5nJ/UCDtWhJqB33usQiHVKnN9GqeAb3wKLWWr
tp4/kSGLVNrsW2TwjiDaR2r4UUrEQnwDCtRFIEyNr16Ol1gN10EDCKWbuV66CPm39cLQHGrR2JW9
i+urvZJivuGNAvFmy821HMdGXIjp/vaYKGv93aA94VdNwSRJ3tzRi66BfbOa099cqIYg5K0YE48o
wE6Ed/GemBg91De4Rsg0j/eXv54pDUgcGI/FZVciIKqrLgpQuCe7P8YWAjX1AP9ny9LiQGux3TCz
+iKuXQVXNYG4pYH8p8SuGw+Nqpv6IjPIiH7HzDu+mOb9vn3Fq5T0Zc3L2HPDnGv4RAkfV6B3DRes
G/axuCU/5XD8e6te64nUu0EUTOM+HAMWLt3BSTHWuWrbijHby2AANHRzgfATVlnUe91qHCkDwzbP
VG+R5BknnlPmHA3jXqzoQQraQQHR/3wRL6DUXvT85YNX72CEmuJloPAyGRXjKRb3S7xL0ILPiNvh
nOR6NO8jAF1AFyn5lrVxn2Pwvu65pX4P8jBbs/qU39XKphpZcCBslk3BwR7MFygFWVkeMpysRlNt
0BhGXOtKEtcNA4cf6Cj4MmaM3vh81dK5s+Ko52w6uGjtUHPxMsZHzcq3IvbY+pbJAq2ZeLtGlUf4
/mDiHl46ll6eGEbyOG/qK2zOo+4GfjGMGFsWA5af3d8CpVbvpB3rw4hg+Twh4VsiQUGLG4LRejTK
QwCrJDoRA7u+OXkHE4Qh0vWOM9wtYfoMV3ae/MkUQxmQ599iNFRZBUTq3XgrDZ9IGfT/x9IhUZbI
OpPqTECjGBtB3jR5QGcAcAZTtmzGHQ/X0WmT4GOKO6ZbY2BPskA+X/MfoPlhF1ChEI+gBoz6IZQQ
dMTroyFybpWBe5pSiepwxq3LSNxqA+AcZKKO/OGSc5889xHlCfRh+d9q38ZTyhCK3LQSwYR9dATB
rPVmTvT6RMShlJ5W83vWGgSqFN0Xg8O2W/1YuPUxxfG0DiCMzACC1HKIlR/xRr/HJl5xZmkFwJdt
CQ34NQa3P0T/yIZB2wQ+FrdVIqUiARt8SQ5L0iSMDLAHgQRSkV/Dco4rqgmBrDIsAsZmqCsDzLxH
fl6rumeDIgUJyJRtjswrhXWooxnPHkrw3YL4ZeO354kSA3UMsqra68U6kYW0AToSGEEhL3OLqpnw
bnNTRMbEwIeP1A0npzSa8/AxDqNvz8y4OMYqYgJPvVoUc/UC4GJAT8ZGdbcf4K2UCQ1y86mZmtTZ
0RSrLwVUCZLv65DFZiC3917uTGyNd2rCvRZamjge14bmUhfeb7uMwnd8d2fejbXJL85BHSkGsjrn
60VQZDjEa9BE3RPkmMLOzpgLE9dHI0yxzUN7UjF4Q2LwPwVQpYjaWccd3+2obS3ETsxCL0xYdO8u
R1ISAzdl476mnPss4tvlKEI5W4WH1xWkClFUrGKljQZZ4J4XKHm4MHBnNIAiQguQmOz719x1Jmw1
jQkilyeWTpE7/+e6l8Db4smIfKp428vap0tCkOPj4o6aZK/cZ1hga5STvZR5xizVBpTLcxaEKDq2
4B/mVm3L/XJ0Pq/xGw0DnkXgr6n5/CJj849wEL838q8z5LbyCkDb3Q+UFwjVqSaGuKx8QIO152FY
4Ol3iFyyyEklYPGvBlrJJWrL4GtoHqMyOzBFLmoo7MysqmQqxBG3v3eQ672JFKqr+8wGNIuzBR2o
feEhCrVZxZnJ7ifJi1sCyoDon30AMBMNpt6o10NC3/lqgFi4ZofJelkr5JopcoS9CQcHZ2Va6zsF
LFGNtN3XvqPDp+dtbE+rdMgPygTSIadY/r8sO/CD/+pZ/jk25/AU4cKbBjlj3ZCVh3KUZHc093aJ
2b7fdsaviCDEOIpptEKLLamkfc/IRRKg9Bz/4sCuZoN+PY9uKZkFBu3AaY01RQHc1lpIRg4Ap/no
i2f6XmPxZ/ojiGNEbSx2+P+m3NjMe++h0MTuChkfwd2OT5o5QISW2ALiCkapdsaGB7TlN6bXCEmB
jOz35E1QktokJAr7zZrOyECoQ8bKAMe5aab1Dm2qGfFjIW0SGKt1qTtzTtiFR4k9jNGIrETI82bu
YiukXfz5mKQdt03Ni9tNKvGSAtYjF2yqMndGl/8SMsCQ8XxjwdXKcRuGdR1/U9ww1Su455YXVkYO
XpDTsSSN/DiBp8YszQqa+kTINofYnCANfDNRH0y0Jl2m3rQapBJGFNXFcZYRgoYkSxwAQGACtwZa
aA4+VA1MUpWJIQLLIK2upNWqM94k5+CMSSCiev1xAdoLVb7xLi60y9hzSWuyE9ylTThpnTJiKiw1
GWlMN+T8aWWqbjNgvSjCWCDUG8knlcWODk8vljVPjLvmzbM1ijDpPv2RJ8jTiIwZ3kJnL8Y1kL61
zLqNMmnT+Lbj44Gv5P2KYXDt23mV2eYqcWjEjS35YSH4d2GE940QCEppYlDTXOb0Z7cZJhhGgiJz
VOEJI6gDUZKf1A49BsQpLJoTwXb64O+jol2klvplffLB0XG4jcO6OwVaANHiWKnz8boASN8BrQ1m
zxYO36VVEVH7ywnmxaAMQvdIMTxuRG/+YIOsqZeX5tqIL6oNB6i76I+iuZIgzvG1VOeSlktzt07p
rFyvOdjkdQ1kVHHoVfxZxTWr9sgolp/UHisT/dpO5md5eqjag2hnUsZJVp1ntN75gwBdfQr/d2R9
MSpvFn7brTYjbLU73pIsIAGAXTf95VUayotZO6HtT3mQYtZQ85lX4noezXBmUhDwcuZW2a/RTdAe
NJNHsRGtbfQPFnKr8BggWCs2CKeAIk0qZkwEA2OaSOMb6NPjI43TVx9Ij2cFweIKerie8jHP2zgd
LAkEpLs1IvS3Z35si6ICRhzLl8IIj5mSJuefLgNR0kxHlnPBoUNBn2d5Ja9ng5bqbo5B/98NIXs0
5+eTiz/pV66Ju6txhx/2vmL1RwaP8oWDAZWMlHAS+x2wk6WPexOUj6dPYb42d5dz2pnIB51RBT5c
NptB4n0FxcYubPsHp/sb7Av22OvLBj9fRt4eI4jQZnUwjg3Dt8Hp59K1wKO8K5M6MdTlRjRfKyuh
NWEwqZhokAcj6SiiY9oZJXuOWLcVn2B3aVzYD7lsXt/CtI6gbeokiFPD8nKhALlMvhQuRFMWFkaJ
jVjyzLgn6oIId/PN7CHRtaFwPklAiIrz8qM6dCdcwhahlIhY0kYq6LNCyuhX8ejAD1Dg2wArzsU9
jXqx3pyF3pBVADaVlzCdZwvuoJnmABxq2Cgx/bozKSOhhieZVEh/r9ALMPqoQrzIbatMzCbPoz2i
NJ0gkuPuhjqmDdVHHnKRI2iQACv4DVmjaUecM9/mLOvVVXzaNg2O7EOrBJ7Np01cQ6ShmAuoN3pq
9xhu3/1JlVeuaViVw1aq++jftym5IqsOyK41al2wxgXZF8ngjbcdk57+4G9M2it8JZysJ/M4EiS1
T+DaUzIDEoX5yZKbPl9zP46b/wLr42jAFPAMbADNrWljrQ0XbpYO4zVUoJL3mIfvaaePzSF7Ffba
KyHvsEnH/LP5sbOXKsKJ3V9SkAuHgqN9Vc3yKqiC0NZb75dSmAh6W3H74aQtOIuUFjlHQBhHTKWb
C6CavQwO3R1lYrpFF80sEeO4AcyV0ul3DWuTshgMPnuekHOJmVUOXvxfi+r3fNXbZWRGHN7x0OP8
tXwxw0WuN3S1+UvZkucTWrBdB97Aa80ObENF8JfkIe+Yc8WqKiMuHO7H8kZXTkG4NRV46M4wtpeP
x+YxJqC93ZMvVTbXnVGgUV7dFDvqLdgwPRYBVpENF6AYBl6JmzyBM/oW/phYZum7lPS8v3FwTZEp
A8JC1mosu4FuM4xjbrobwxKp8ceYGzHwYcPUkGKrF3iCmpR4L/x47H5KAWFazOMmbDBkDQk9wRUr
LPcMiUIzzTdlG/6bWux/wgM9S9GubAGALrkl1g9RFgFYfg0QD4mmc/LK0F9Ty1DpUCb0baeinUBn
5Z4N9aqu72hl3XlMSWM0utyVYGcKbbUxHLmGTpaeDhqdnuff9ZduYTkriaREkpEiq97GmAlJQJwJ
Ag6EZ1utrScvg61ZZApo+tTKsP9ErXQpiNe5ISWhKHDfgEGAF5h5YPxACHjxi5tw+f6vsw8cgtnm
iYJIiDFSzu/INzQ1zJXF07sm89sm7Qg6CrZli/Nql4d7Gn25iMdzwOF1RW7QvStq5b1JqxRDPYVm
qEO9pTlUdFgnT1gbe+YUAH46iwYyx0zPcE5aQ5e/1RVDlkkFLl272VpFlx4LIkzhyuBnWUukH/Jm
GRpWZ91YV/YJmg/2z5387XRTHTcFiylgwbsle5oNSKaV2p5MqJePeTh97sLfDwszonAqKxX8Q7hw
WV+biH3ri/ZhXTu1AvY/29YyQfjgnj2L0Qie8BEoGUfll3PRZRiF5qcQeyqpeTVb9prAm+sqLmWu
FybMSvp4YTJTWv31cfzLnv5nb53Lwk23x/9IZv54gncVREUDLBBaE8VjEu1MJcEBpfw8PuVEehgO
K7Phz9AjLsPvqVkegnberEolEbUbLyyjVU+VYGyv87eEfV4RpTGI9m2R+8LQJ5pRcKAqoCM25cpd
ifVGoGbNJwC+BgkF20J0zg3Izy6YuvdXk0YNQ7J7DoEk1GFhfLAcczd0V8njA8VQlSX6Zrk4AOWc
BFSr9iioK4UjH3ewu7UQQPo+NLN14JaNMYdqECXAQ59bhmSW0+GId+fHowFdHDsu4FDtDtZSkJ3l
KTjlrsqCfULX0R6Nx0Tf3voa35LFvoPH7NOpfdKRnbQZ9GCpJw04ObpeVPBL6VRwbllKLRtlxD07
Zd6wuhLMrlUNSX8ZtN/q5KwvvQLH37sSd5I+u7+OzEnoSUCi9Hkr0Yjc4917jYbVbNlljKUwIwiF
KCK+CUvw5ULrwHndgClLhSYRDYASfeVPpS9Q6Z02URAUB3r4di+GeBO/6zdxAYwa/66a2PMjCtOt
JscK4FLvzjlxWlCWDwoQ4flxx8ogXmoEva3dbcPkg4A4EXjwrme9vjZr9IGVaYPcsVvcE0sz09SB
YTF9XSFsC4RgrUx4xDlHqBYroNXe9JtI5Ure/xqua0kNclgnFdQeaJS1UjbOh7wnlNbPeei/g8ah
WE6iok+M3GxNMOQGaS55l7UptIZTlHcBqDQxIZdNOJVeVwRjcB/fZxxWM8cRcWT3rYHdU+ZUyH3K
KpG/9+9SmcXEtDl7scBgCuCxLOp9NKoWiwC3JCDmSadCv+8Pda0aZvCGDYpTp4Crsfd/ZEKU2ksq
wyUXGvbOEP1FYDXq/mueX/rewubySWwLOvN68yelKR6obb99z7YcNBoTQWbDfXVv40ETIjX7hHt6
SDjN6741jomtXsKrUaEQOJGepBv/Zbw1l38f8S4VVfhEk89LvGfy5PBtTbh14Fq520/GbRPMRReB
uEXp+zbj7hKXnNScI17Js344kBEbtymmAiJq2U3zNlZMQQjsryf8S7tgngaBkeEdJpLnWvJsf+2b
wb1XWSKW3iY0+hdkAllF+au1gUsQF5loIZZqfTUKUSEn0L9GOl9IwK3LQmuDfQeCuAOHtW7mYiqu
XNq5n1aPR2xM0CMV+Z1BbVHETT19hLCHMmh5HPW71rZNZeDfPGK8DzKX5O6cKCRgCemI6mNAiVkk
/nPPft+THBR5JmqUKpNvlCbQfnf/sTdUqt5T64F6rFtwWDoG5ejQjmYbsHT6/7Nqb+SCgZG1/BnW
U0mMb4Yj5cEfjwiQBXTYF1R+NBqFg9bfvmmrdZ5/QlC9PmIwDskCOXubI4UtQIPypcVPEgJ/Qqho
A37+RiMcyKmojr2csW8XPvwsPNjOCzmYQQ0aelLeb0pyCZ5eJhesfm3nJZMyxq0y566vCgLqWBMU
YshxtVg87ZqZBUtNIuT/kGt5EGk9bmoeeJxzojXTul+1ZytLq4j43AC2+UnR0wyus/rqQAFLv2e1
L+OYOk2lZ7kEH/morYNwd1pw62GLQY5DFeg2SIlCQt9NXhE2XBWnG8TtyOHfzAYmu5SWO6m4ncmM
boU7KECtwRv+NiU4GqedQTkDUzZecmqlazZdl6a+BW/a3IH2c5cn5wm6OXF6gwpt0xAXRauI5MrB
uhxCnvKJUoKuMpT7+sw5nAV3jWeu9w3OCmVuSZ7C5JmuHHLxdlOYkoNHF9orVcofxDtKUlGf81Mu
lOdYq5zr0sywg6F+tz4lgp8JPK2uz6OS9xoX3bMNVkeaLqMGRlGiu6oz1i5kFRY/55Ka6zNAVApI
weJk379ovlIgnDMhD4+zK+lLZGVTbXdLowsaIzdxVal+tD18PFwPXz0SF+n5xnZ4SER5iHG2mVKj
Cska0VHGVm1ObPfAqw/ZTp5ny5fz8M3vvD8lqK+5WoTli8EEC51WfcPjAmFlvWKfH7ldoVVEp9vN
bs9ykCWzSi1TiRKaeQfhR1vMYyvYhbTWleR5Q4t39YX8Yn1DWbZAM7bgkVhg6zc0flT7A+jkyyJN
cfIFLx+2Yo3wU51AEqfuwlhVoiKx2k0L2PZFp3TyFsaWUNwRhCYOWQKgMHo2a1WJh3C2v3NpPnp2
FsjdyDOjRDyIe0uQgTmGmMtZDs3hiGm0ygnvb8RV38BYIqjnUdBmxm3Wqvcy/t6Lm6ClotXg2l+F
MewXBhmGLpOIHz3pjzenrXB9OlGsqZHc1m1A0Vos+7OEVbCgb13nBCr6ob1K7kshkah1VNMOSyGO
I5DkJOwe5RR6A0TPbupLlUydjdpA9rgeL+1fctakPVowc1IOQLKK9BSy12KkYBNKbu/Q2LUJUmaK
k150G99m+U2nHD/kr95HubNppPQ2ezG5KHi/hCpGZDvW0rlipS2bospfDdAPE/PNMzq8tX8eaMa0
128ugDuBoLmFIIZoY9X73eFIW53O+Dgj36aObOznUGjQ4M579LicXauTIAowy+ePVFbYHGAMl3m+
LxBuJ6uKs+BOezB4cTKV3STyEJ6GKPNoH041jyMSsljgPLyk+CKXA198tW4NB4pJxfj3jKV7irSn
RWMXGPDZ5KCu87RXVdIlmRHFCR/AbaVixCam/djS/Do0wzzjvZi9iSE6TI/J90mFEfoTmW6ZQipa
1V8GWDmn/sO5yNCJAOQ3ZP8DmSVpchQBjsYDtB+sdC6JKRQlj/vcuvc7ac1LZLSKDUdxn9lraLom
CNRmN8NB53LrGS3oyuPNDS06/3MQ6Btg8d12gqNs06TUrvLy9TNsbSUK7aZ3RvnfsM2RoytM8U9d
a78dfovXrnPubiHOEPZyIMRtlk2Ugi2bIxhIXyzVMsBQTWLMAO9Iyk0/y+Nafju1WjyaYg3/J8ZB
0IzfxD6lWQKvqqyjocKJ46oBV23JA6d3n1sbrMvFNBzukdiD4FI1SPYd+/infRzB/VSlGsEH5wG0
tkKVcOro0UixBrMep3BspWB7z7yy4f64CFJvO5ZkeGz8CoFS/bt8sH86jh70vhTGPaRC3t9LGyZV
Vh8v1s8EayWBkFk12ZiVqdTfB6DAy1gEDFaXuKs36+NRdXZUZvX2ffggOD8Qm00RvF0xMMaA43rX
aq174CqCc6u9JzbBVQwwxU1bBaf7iKflCFsTdWBSlNQdFpv7tur+MLWtDW902fRaCMB7pg3qjAMd
aY/5S8oQGPZqR6xAxSTd3yZOdE2jibJtjdf21ldQIsWoJAAQs+wrDSE993jnWZAmdJf+AJLNx1Da
R74kgnbN5YGv/9pw9pjUX9Zw94GyvnZ3g0iFmt3zaSyg3z9qEplV3MxdXdEZ49v/eiyeivgGGhA+
ELp81PTn14tfq454nw2KrO4I9TR5mWua2ufU1YHrwVdxlPG4KN1EUDS6/FEVCUvDs+5nuOzFr3mY
bq+DYEXcnY4bTYTga3uc8Q2V2DdlDQubOa2YU3UudP4tJR0vRfEbgiZbhJMuOC27USf0OkM1Bwbs
kkMoUYzDa+hzLB5sJoJpK2ev1RmHDpR9OuVvEYH8LB+4bZDiO632SFkJN+ilCnAAeV0WlPBu0Dfy
AD/Mqy8hGICbaU7x/lzEyh+IC6usBkP4BxWVazUfrLnhUX8pJ0JcxRXhDEApOhAcIGU3cRqc9Ssu
OyboX7t6pVJ+wwhR4BAET8p69oOuDm/bHMCZidmQb1UrP7lMtu+ZXWBtXQXTYScYnF5PP/fwOo6u
FgSBRO7GnSOdB/6eOrHD7jLAE3Q6fmzOMWQxGzXPBuXN4RLCdi9qeJO2L34YeVnvHZ8RQ8G3c/AC
FyBwhS9dxM/l4cx2T/1mnHXwXDogZ9JrLYAZFHooHHebBBuPy2jwjLJbYrEAMnSHRubMome0BmBX
jbvfpf9/7bEaHjWWcbDu1tJLJZcGu2wsPp29hbvW/GPkTn8YI8vBfBvH0k8TLLbD68IqSIYhLPBO
r2cEqafBLdT7BbV8dqbTPklJ9oRaGjS+t0gbmM2++ErrN8eQ5Rs7JDH2+rIEJdGVvup+t6iXRPE4
Z8GdtD8SqvKqbJ02NdCo/m6BNlD5NM1khwbEqr+twPCdhn0hu9t7EUQtyvcYkuEJPZ7TDYXRTgad
596GxEA2WQOf9R/lDlUwM5khE4ihsTMREoyzAp1yELU85Kh4PZ5QWrdHZiMG7bRIcWAnc4PLICAh
ZuUQnHK8spoJV5puI4cVeToNA9ZQbf36oisom7Cpj0hNC9hsjnhDvJ4MZQs2J4iJQ/glfqCnqd1l
la6k+tPYblSo0OS3cbQEHXOAMVHG2b/d9ggcNkXIagXWaby6CRsvs2Y2UYDuraMSqI9MLfVLLGYr
pu9XubwcBO+t7v97FFlv3I63Wew+tmgCEccq0HuveAZJvkg/pPSEGOlpNc+smf4m65/T7Bqra2DA
VMFWcejgkqLxVm7nzuWNZnbdO8vXEMnfXGqeSJt6cKYyrhw6P4XmAgij3znhDTrMhEInQnogQpPf
vVIIwBKWNgaxBcixUrgoZdkE7we+ucAXbubCyR4JoiqXJFPM+QoH1zxHJqckvd+VzC7JEnavWDey
TXe6edJcE/qQHvsHl0PIxZkaweS5eP3cHsNlkgoPUx4HMXhzKXQq/qkHpQcEX28oQkXieYwBOvYq
PqORCeLBz383bknoD5filgohlbYJkB0OhQZAb1lioikxehO5sNDarGCPANW9fhqAbmJdaWNstIDe
67kPWbp3adVoEmeDhnJNFL5edOcICEAZ+7V4dECQchaKzoWErleHQ7PkJmbSuFtQrgaD0Uswsl7Z
qTz5fugzz4Yt7nuWHYRPoCGW4b8QDLepuu795wcY2JeTSq3g9mT/LSNYARye54Tq9u40G5lnbUwT
yJDMc6sVQs3RZrQZX6DaP2SYEPEuH5VWSxVNc8rXymX3I9LhXQn3N9SBi7nrGXW7tO7Ad1340+z/
9m/3Og7L7PeS4FsWYaPTk5o6ermAfZgfVSwf63JlPo5n8SB6yXu/IVq0Io6jfKXP7Mm+p0VmMlvk
cW+wMc9+nwJ4GFaNHWvYnpGTxMoDlHsHXWH1JkJWhkEba7FAXgLs2FDdOtj3im2Q+2cFqjT/zPGa
aT0pVce9PTM0V94Cqqgm/b4WPtV8Ox3U4NfgmEGhoKhESxqgoyReUtnP+0SveNDOGE6Th6S/OxJz
T6afHnnwKQ2CcWYFROLbO7gat5X0SUiBJDm6SDjUZ3OAcQ64x7K8XewvBXRpO6fHbNeFYmOJJaMw
0SYuqi+Nf5g6IPErXAPJurAUNBO5qxhV8M1b9orqoC5PC+4PnTf5DMS06glEEn4b8QVlbKYma3Ob
Az1LHzKsjCQ7oIEe9AkzQNseIuhsmU1w+dGps5JIhPs4tNLiqdOi7AckBSA6SpGhXYTqdmOU5+Cl
ZXp+Zd3wh7LnYHWcf4uXN0wzV/BfuM2IAZUS0oyTBfYNcZhJNE9LFXcEDnGcJ9XXArnWnl7Rs+zl
ucrStMzBJeQsL9MjAyR7oK71YZYDJ2cXvg32mRdr3GB/wcb5fjN3wgnFTLh5tNbGLnlIOfEAmjYc
kc2NGTqZ6DfVNAldXKAFvttKcUkUpGPjXZOtzr/o4nP9mDgvWUwyszjpkdHocberLsbLqHjWUUN/
zEjQILtmPR//tOme8T6979DansL8kNw+VQ/G6kbm9GgUHVA64fOoJ78b1ypmWWf45kO5LnJ6P7C1
Ps5PU46HN/Wo2zlpFaKdUrhSVVOOGWAo9BYcWNHzM924IgmLlfBCDhb+jcqIihAUfBF8NKafhIuw
9Ged5K8ItBl9Wxukf3G4i5TNbDVJoY7SbsLS7IDztpGc4e5uq7F/youvghl6tE7lPiEX5WktQCav
NpXRSXJjvVoTDhrmigHh0DEKbP1r9aWUzqRW9lz0ydnadSejbWT62hSh2Q3jvu5sh7B4GqdeTVav
FmsvIz+3rdF2UjFXuy0ptuCsLvDlg+XOJcEnC7niAItZx88LSCo2Cu9Nps0sP1Zl46garSU2c3FJ
0+LRXXUqs0VcU1wmjX5m5AvpErHo0SnZMLiJAWMoAGNylGq/ein8SVRrgD+nCJlKSudg6736C8bI
kngiJDKPtAgYAZu6spoTnjZHHcGpzsq9ltKmnvw0cx7f5odmdatMxiO72ZbaqSox+YyI1NBSMTQ3
91n4UIU+7eSwT/tOI5nzPcFRYnrzSouTQh7kLDLuAkeQI4zY/f5Iwwys/0SAVELSLKLPPRLCafG5
pPRwDdgjiSA5Pcz/AKaiVC9I5nC/OPZcayBbvhkdV7R1VkSXhjcx8/JGktdB7yfxm4RGaT7FqHxA
+P74yD7ur5R/Ge5s+VyCmbFwdbSZS+W3VBrjPlgCKPK/WKREhKununVmszl05mx9JG+iuxu475z0
TRnnIvLY1kE272yhXM+pgmw0sPw9GoPiYhfS/a97gOjEEwMyxXeZh4a5joHB70meKECSdHyFDXHX
/jgjGEuSdzY7ZZPpSvPgx/tHU6L9amv+SDXz+kiKJSzUEb1Xcu3qno4Z6dhiHc81p4rpw+/ni9im
3CDzNGapfDilALdQzoIm/0OvmyWpwO4fcMTUj50ONdqmjX0oL4ZhYNeDs7fqZfnWCA9ATaNn7eeW
ACSUbyCeSbT0QNLrAjs1W63GIGBfXyp+u3HDMvAXjYI2Dsw4S78MrUX1FHlC06CWvEgCHFtBvamY
B0BZfIOpsyzq9lCuB5NXkXMyz4yhFtjj1oIgFttKk4E5N3snMxOw60VIdv/RNJJk2FHGDWsfOBcB
XRVOwHKt79u0FnfA5aJQJc2LJlJCS4Cyh62rDoqvgxRYXZZ0+oHrfE9KafLs5mY2+EjboEXDIaNx
WySrAp2RvRXOkDHTG6AmmMsP3pEP6vhZyLCz1zhxvGgZRN7MEtLJRFKj7IJYorR/GHgBzPXwnG+T
YctsdONKNw+kN4m/xYhTbVA8X0djZCQNmvWbZaQwyoTjXil6uGrUxZ1Dozwe1uWNnTUFXcj/0BNV
7LY7Ec3ksGcbswZ467oKg1YkH2VeALtVOgaVa6DS0d+LL19bRy1UW+HAQmQseR2IXWbAIWUO2cIL
ygvpoSKPHWbejRO366RTN0VDbH32oPCnY2VRjDPjXVgP4jBTA27CbP/0UgxB9jXZR4ps60Uxr5ji
yfzOBSOhZWG6Ukf+JVi1LjJezfI1hC5nVLZusrUrpWA99nmyv2yHHMPs+hEwU+swS1bEL3SqH+Vl
KKnM7C5BOhIsZx9UTs3UjbjdtMkf2+9iELj9Vnj97u8Z0KDOXGdry1s62e6QX0mfGRQVx65fTAvQ
ez700Wp+SSAuCu0eep/LC3W4DxgHIFwtlCA2PVUx25GprqI/PjCRXcdDN2evH6qFoMHEtHt7Rpjs
0V/ptF8vwXpZKFWMJvg60Tb3PPD5UoQfUhducWJERj53BqC7yfq+KQGrfe/RZPU3IDj+KQ1sn5TZ
SI6owLsm/fW+kPQvtuOUzREfH8vjw/t8priknnQGHq8wwfPon2zr07fvXZ7G2cLCiHDhneAtf03g
eADay4b91HKY44R3t88YSc4krcHqhhkwntOj9kskUJE8wEjTuVe49+X26Yym9TZBZvB4lR7yjbHw
ofy2l0xrC0Gc14bQoIhd5NqmvtSDpKM9hIf7FLMcIW5CleTr/SHlv0YgpUm/6j3eUglYOENUAN/5
IeEt3DiRu9V1mMGMWjk53rwuRVgqhvzd4jUv+dOb1gFSqaWfzi/f04e573cExFRELYZ9ePW0x6kZ
gY+HaRqlNY+ION2NIALAvddLMm250xYZ4xcwWCMF8WB9fBpBdX7dwH+qvb5xPrvzcLp9SUB2UtpW
Vlqc+zdlBvMTUgDFlbYtyuIFgDWDZK/S3BqrKu55IQ9bUA5cCcJZZcykWIuCWn7WgMeHhh2YLX5Y
7Gp9afbJDPjix3P7YzpmsqIP4lGEUDWPCB3CWvrifTcop7CgprPxCYbFQAwQfwGEI64PPrOP64Av
Bb00QWNQ03o5G6O6qMS6CJjQHnbPZGid6kNjnorb7R3w3K4QcLxTmekv4d682K+TAep6tCXJLW3U
fdJzx10KXzQCtmaAFoXwiE4W9GCFBWobrGD45wn+Mem/kh1IlrTfEA6LzT/amNgauYO4WTcwvURO
DjUw/6RYLScW/Z9NEmvymp0qBWyfOGznS3LUAbrhA5fAq6H86aI+5X5mD+moepaCTjnIswfVobwQ
+KraNRK5Q/pO80FJJzR/uSzdtGS7c1vaZ+AJj7E+eoDg2OmX39+8ttiIRlH1yIZtX6NE1i4CU1RT
QV21CydJ1d1V7Fy4SjmPmY4kjF8PMPcAecAWPWQyt3CiTO2pTL8tEa/6qnedMayAYwo6NbWcQHAd
HJVWYJXv7LKsp64s+rJP/UGDqMhpsgQcsVefFz1SVKCiK4hA6NnGg77ZI93GrZ+gWj8K1aAJ48xA
MnXKU/i2c3w2K4LLhqLYWLmS2CHsI1HYEv9KFH4DiFIrhEuEc7iAJdE8GT2d/sK1/ZpafrO6SPYP
p0vLNHDj6TzMGoF8uhjZF38suZCh9QifF0TWESYphbU7aKtHVCyUSnR4yk6Oao2sXR0VG4WLJUj/
Bn/whc8k+CKaTFN7bCXrSVmlfcGov4QrsWYleDqv/Yp8l7MrDyxk4JbiqIz1ndGFM5bGILXIsA/8
9QlqFDDQXJHuzoZGJPVIylr4AueqU1oDQhEJn1vOOXnEoAwhAjp4bMWDK5tyAFWVwjDiF/frY5eu
iRa1B8ssQY6+yl55fTg2cGIGx91ZFnYi+B+QJDDSiBGWcuFIvOOp1vk0bsCU3hFoFFv4suDdE1ts
p8XyocGEd0RPkmZ2yvHdunB4fxeV18hRTf92Ca0/Z+2rKuqC1h5sV2cqlGTxBc0j0xRBtbyNF1Ro
hZsAqBNnMhE7qcdClDDzdbIM01UiRD7ayYYkiRay7cqY+2qeamPykaDrHWbVFS7ECdgZhuWBMDZT
8ZNBAe9eRlKvH0ZoXgyxMDnEsWRuQcYOX3Oh2N4WqrUCyGGACgt9DRfqKFe+2ZeOlQE3/5LMyx8l
Ocaf+q2i534l6oGqRR6RCLTpKCwhMfI2OnmTfxmDr3NlW+J3NeSjf+g/z4K+XOFBPGAzGekByx60
X19OLoucGdkIaoujHZLDl3o43EaSyUPFDLaZbaXTAkc6NYw4k2ZUMQH2s02IoUXYTTOMTBdkb4ts
lKxvieGR/BgCzsMS/4zIF/6Wr5vm5zSRFOwcMLQ4OCeFEnG8pbVqHFFKb699VhoutKJNOC/aFB97
7fr5+0NArsCM1C/uF2cgiHqQQkUObFmwi5V+NZv6ZOLfFdJ4mNhbBpRNBT+sLn+Me33zP2yH9Hrm
vVC3RF6tOp7FV8v11Sda16zWH3Zsp5N27OuPrlSNwbQ0bBVvD2oLtHjen2L51KrIzy+M+XX6QzTC
jJygorcFIAuzwLFDVtGbZV9RwBK98dXkgnQ/xdE1C9Ie6FqxNDDJzfneqhn1kINvks+LvfHKWOm+
Pu3ClznXID/hDsXJUaYWPfsSmJJE0QoYkmUgZXzX07k5aq3bU5roWu/xu5s21kM7PwlPWxKo26i1
8N9PyU8dsjeTVBy2fWYJo+CwK1gNhBnqEtCEzC9HxRL44i9jTLj2Ds08pxkfZ78TpDe0dW5SUEZp
CYttKz+A1ArpvXlDPpaErNmQ9zdy9i0M06JCroc8+OcrXP+vM2RRBYDJVoZ87MnH148eEdT39C0o
1O5hXB87iRwNRvyD+TqZB4rfCWUrQnIezeiWexC20xSW172YF4Lg6AUciC4NqoqI4FFqhrnBvBH0
o8uDxvKBr7VeFIL0A/IPd4KtU4tmHhjXQ26XhVHIx8IeYMff0xav3s8NWccDqZ4htcrVQtl8o0X9
uTSC7TU1Fi96mutvuN9RLQBoKXtm3tS5dWNw/8w8kozAAJ8Cu75kgLF6qU0HDEdApy3hMyMdroQn
x7045459hUW/kzNgfj0JSWX6tURh1e+lxCjZ42EKioT1gNEjjGaHAapkcTKVEvSpmKOKLSKD6CMp
PqOAkBqk374v/cGp8qtVkqdvkRHR5sPCudRCSlMUj/xXQvIw4r/7jXdaOv6cFY+WC2F2PWe/A8Ui
ZvFEtqn6oW/j/cahwAjimg6wdeLBlL62Gfejr2c830lDw0pTSzXlIuwrAMrTIbdJiixmSXcJ7pNo
lxqABrNa8l4A5sUeQ2p4nhioAFxYWmkulyl5JaMjqif/m4YDgSq6ryigJvF54WOmOhAvGzNBazzN
PHG8tyWkL+QmPfSLIH8ZcE5aeH2Vj81E0lxVPU6g9g3lr4nTBBplpb0hpXLAq1Kfk7g1FzziBFP9
OFBHDBKYFGGf70QR3cTK5MtegHB4rB78gqcJZEzWtBNaDi8s7cvlWwGstF1QD3+Aisr1HF+qm8Hw
/mM/6f3/dpPSUz8BVlIxGYJtm9uc7L/r6EuKqv5RRDbSIawzLhVtQuUQuIRhyhujlD2S8cNTwXtQ
Iknfe22BFeJsUShgTA7DGkYHSRM+AZ7HQDbkk2cipeRp9qu/zmIrJA6DB1LakDRybFtyESypQQ3K
+3u44+ITMdL2uT4LQ+iJANk8PVF8bADu2bYppJe+Z/lEGMFuLjIJWczfbjbpXqVmnT/1Sv+Y2Y/O
f+aEQqVPK3VLaNlef2vMYxOo+uZXVld90NhK7XueP4Xca08+gNcsbiWgvIIir1IXfJezRB/eP1Z0
OSypkoE0m8/TfgEjOitysF9GTgYCF+s5dehlwU6189uSMatogCkgEwYUMZuiySfobdnpKgcFH9ys
IKkxWwFW/OLpM7SPlYmxXFp9sz2MwuYMBZqxbGAek9t1HoLrxbcBz+I4BRtbF8NCi4zOHXu59kyY
dlcTkEp41aDT9FOcgE5HOdyOVb6hl9/tC1/UEcT0gDaN2s0WMmp8T4FnwYbpw3Wd5DZd0VGFeu3y
7SObD9bhs6iMNX9DG/TI9kmdb+ArJgjU4XtQrnNjcglNXIwT9DeaPBb7umx95Mb2+eeBu+m80pLk
Ukp59cncQp+gGKKxpaEaBCx+bxDvaSMMNuzTaqqqFkSg5wNkRuv+bbXYQ8IpgkIQG7bnj2QIFCg6
VkojjaprFWR4aZQgrLvu3dT3lBe+6dfPZ5IvfO1VXRi1emS7uoucjV6MzZz2cmrqIrJwoCRl3Xis
3nkc53A9eXppyqupvrts5RqPNDW1RETg2/FwDjqSjvLI+Nw7YYJ2FcvN0anaDPDJjd6R3KGa1jXY
kRLcRv1KAITRFX3A4cE7tdJmDXQHhSdfweu8aEWQeoyBOnO5OtMB2hHuWcu4v7WA27RJ1OYOyNbn
17PW8dCJyeJYafoesXPAeVkPUhepuN+slEwYmmARcsk76lodlEHMmn6GL4c/bCD0CboWx/bm30cj
tljUdtW3AGuUDc/GQyi9ZjzPq+VF3ucKUY4VXdV0M30Z7VSRBLP3MQphFGHOEnfnYqwD59KTS0Po
RCOPWb765NKkKUqQXVZcGc2+u50wL3L2VV5+ICqEQvYZcP0VNS6CgZBQPb5bS3qURSY1K3v40zRS
65m2fp3dkGKSQwRPzHsDM9fDMLEhN1fbp0biJTb7B3wwNqn2rPhjOsxirFNOGG5grc0GJbIUHX51
YcJKR6GIpAWoH0W4StrTbxUwMzu5Tc1iOENe6N/jNEtnY2HgGTrFrDvc3s2ZXztH4X+0p7O2p6lv
9d/iAA/N247RWX2rKXJQ5yyR7kt2uUUKUK4SPUeRLLyo95lV156EdrjpKJyWnkpKJLV6Ur7O1ish
2rE2+oo+ZaOIrw/k7NEQR4k/vXI5oiMWD7dgoOsXQtSoKU3u3eM1Q6PcWR8NARNYyYoaMG1txyTy
I5iYgItyZaUcb1HsaTzw8TlfKSuHTSQ3wNHYn3fwE8ebK/j5DqY6ndXWhZ0djc9BCGc/UI3iKSI1
e25Ow/pKQIQP7fJGhKJn0O/LP1O0q2UO/bJ7sIwir5z0ivETh9wbIz3o4HRqU2MUhhb+hJWn5n4z
C0iwYobaEOFN9wdKBYfaOLwxquAETOFFygG28ofdul1U0YZpECQfPZm6+4j93rXFc/1UmtdFjqVT
zPmUzsaRK79j6E3bttvEvoHRTTJVIuoDzmkRw6Z1b/QgPIw3h34Niq2zDFgJm0O/S65lsY2U3Uia
AkjzoTTMzkuBW0YI1x0PPHR7qVMDCSvrQGNFpIWwZf2Fpyug7rKPxSJBEblRERkRqFVgvGoZrTbP
K/pYi+bLe7ixWRrXvdFNACcMlRFxvKFpZbaN74amFbNyGKEaHsMDl0uu5C8MZAt8XqEbRbJLl/pU
UWkhGobY6U7WcrfvqbUMGLzC/DtU0U5GdDJpVYyZRKkl0otmdoAUu0O6g02CWyaNiU1xgP8Yssos
J/2qtzpaOp4tXvULcMWdT56Ef40FJBUqaAH9P6fwwxybqG1PTyn4VXCap50/OwfAuiNA0rFQRoNF
0XZlfKhBx1UGyYnDEd3YdGwYwNV50CAMj5niKWb1kFKk2+dB7JfGjEIFT2kRvKnFieRSRpZhYn7+
IUxqQY0AviAp3RUV4Y/qaHkDejYS4Ec/NsnfQxCJxfy634GyYkBxFNdtVGqnXPjljNRcB7xbBEiG
n6wCR9zTIfb6URYbccApk5qJlxfc7z/bc3f2GI8p3POtXHLcKSfQMS6A6ufwBp4HQ5I65CVeyhoQ
vBDvCiZADMCnzepI2AEOLNsxziT1fjYUzl8tVGc1Kw+tNw92mn4IFVM2v4tLPMobJZza9tVKnvuX
YMVpafllxL8AaXheu+Gnr/9N3ZujUwbHwZIZMnWiaDqUU2FeX2xXxzYDqhOSlwk6LLuei6kUqlYz
Gjl71BHtybSgZfEkf6+nehlUTFCKz/JeKuOsZH8NDX87WOx5sKSM6F4xtJ61GONfkGFCjicp4A1i
+G/2V96tHLTvbWMsditxoy4ocWI85wIaqrz+ZsRp3t2i1NVgxi962YR1Fg35feCyyuRHhNXtV+OO
vTz/kkpB9DwRxY6BLNRd0ctoZX26tsBRqCkDwq0lo3/nRaPpG3po4QKH4Per4mnsRU7lbCzwnvP1
3DCcBc9Z89KB0D+LBPzrTLaOmqZRhodtYF5UCe16d9ENe7RU91+wxuNfspN8iE/UC0kp3t4Das/J
m6UIENLJMFBtBeAnw77GsDsfJlb4ljPzg8JU1HIyurvJWB31tXcVi12MA7xM01nEYXA0fhcpInuJ
YhNTzLExWXS8JGawNlvEisoTRuTi1jM99UwLbWKUOtNFlhA0+kPsuJw7KidduoYp4yXBoijJLEmk
0zS/SAEHRamp9xMhTmAMYV6eM1PQvDzQGGZzY/2vV+4lhn/uiy9UPGaCP9Vlje0GKWafhUb0YpeM
eNsT8cHnle4gpgCLBkttyk8rKDGt8cS7fgIo3X0lLPVVdEDuHyah2uc+IvemQ3eiHqQWLQfYn4hw
j8qa+kHkH0FjsPYt2RWOwEQ3+dJxNn85AyOTyVlw3AB52dDveGUMMxdYkpGH9VJgHJeDlr7JxVSb
c4YQcdjDlygaJ9ZW6WvJxzsgm0xiQepc6IcV205IHbC3V4edMr1TxaUG4bCi3iSJHdqaZqy+faa/
xxlNpfzICAcflKYnOqzxb7h6gqFV2raVWmL3cpnyhepZB71Wuzv8gQhCoXNiRoclxAPKLnfKVRCV
1MRqpTONiK7thIo/84LhF8y2QdwheGdlekORSdvvdcDa2zKeHzJmkZLLXMKvg1FXvsoI4nIMgoxX
QO59Bzdbi2BeSlC8v4chxMcjTaC24dXKDlwlXO51f3LuCOG/AkKMWuDnMCS/ZnCk50ZvE1TFMezS
VXLgsGz35pIldg4d2mvppXEc0xInQiwRb6FvB6G5MWJJOBZctOV8ZwLtGhCVjOaqbjfPYhSczqHN
iyMWgvZ4KfvEbPabWsqehoruQyVgWcYYTi4NSZunQbG7/Mu5UhU0Zic5y7rXCw9I1GF7WWU1SWDj
Zyh6kaDIgwYA8txIFBXc6BEeDyH336SZN1tBX5kBZVXEhEfec82Ik7+jLndTumpQSOTLoFwG7sZP
ojz4dYENXB5yY5dCuUI3jPkp+YiHHQgdwbnLn8WIGmHG7SwOMJgnwNnQ/+tEqEoUkYshK6piUSGd
EqvBW+SNJrAlWvYU+Kje7ElJKOM7d46x05RK7O3+fbnZ3BLETmAoRuXZ4JtT11dyirbR0OIFGQTE
ciC/0w6GnCnz6v5NYTk0So6u1IXPqHGTKR1//inJwnMX2+C19TsmSUYZJQJdxMRP6TBZXiEW9824
qpR0iiv9IyDBDlX5KMjedjj1lp9i0PcEgAO4rmqbn6pB+UBLQlkVZwPfqs8mb/ItKr3fec5qc7LY
rUreoYZwJwaCOmBVZb7XGBlQocamwDx0lcRRmFkFs4fcsdBxNNSPVZyfdtz4F44R4sqmQ3MkNMAQ
f/DjKtma67afMiApMlKDnPiySpblUGMRhZE9MEs8kTvnELXPXSRkcgLbqzFuqjfEqNlJsgcsX0Xq
qRR+Bi33pAAwIhveh89uaDMrRjYY3Rjn3zzoG3Jyy+LhpPcHqeQ38JGX5xBxlYCOcqEvM455/400
yCsrVWE0oXhQUmUaNqlDVMD96z4xtX97PU0Cl0KE1KHMpJZl/TA3gQVIJJ8aAjxYFUAd90o9Ao3+
74FA08LlOGx2Yu85JDUQwYgo5hfP2OFFCUg0rj9XKgcARP6akdjNVIQb+144Ei56KtTEoOANDSUa
UK5IrmDsYPKjeq0xEhjZk9XfEOILr9QhOjBLi9Q8j03OLHBUXQsOYgHql/nmaBQiECHzX7perWJI
xHbNEfqN6+cLtyu+P//vZRTJwbHcHcLIGwXm6GHERffyhD6fi3+Gz8iULEenrl4z4Uxn+Yj3p7bc
R1SxGzT7pMMOPIeZ6Wu7rQ5ZBXXkQVbtdqASlLk+0K5iUSnpi/eXS1jA22f7//CWMgaSYeu/HWb1
6wFw08AxxPolz599PR23hFoLfhH5Ki7e+yvj7GKyBqcD6iQ89U061w0jq/SQTK0AwlrxepLHhbqy
OXguV5h0VoSPdK3YBBZeAPUgoBaB1Wa154Uhbw9Nyztq+Ld0wcRZ7nQgufmptiSVnFu1q5tuJBkZ
xKau17SNjLRb4eu9jEuh+LgHmD//l1kKXoLQy2AI9WdywKLJ2A8K6cZO4Q4zozhwIWI4/9oJE/Gf
42RUp2nVnsitTiDHt4x0VSQYJTYZtXEmuVxtnPCT3pNezgnE8DycBvkddITP4OmP5ZMbAqhh8gAb
wAnOloZXxJ38dCLuYe1ICA464yAYoxAFTdTUKfG40BDK71i+lxFY3i0En4x6UDl55m+e+PHEU+ho
kb7skiwV2CxdRmJ8GRnUQIQYPimAIZdGcjt61gR6plLH+xO80yL3RJjlgpWW6ziQzTCZ2LPwW0Ch
TXms5En9lcz3ntgZPrUVV1luoBhgeckX582gPiJoBK+83XEkQpichXe53XpQN7Kt1uEIlNWLBSLH
55qaXa8p796/vKuh4nZL6+swx4BfMrkHI6/XjO6zbmgZrmnES/ZJ3QHEm5S45IGexBi0039w/BaG
s7zZFSHfFUgbB8G4QTJF1zNj56zeHPUiHQ3v5tZxAt+Lqk+wwIfyMGfRs0LUSWjnOLpF5fy5hY+I
RfA+KE4FrXs/ezPPgE6fIAetNzZ4lQjVcX2tVfZsWxgQieHWB0zoy0HycyvJsogNoDZE4XNrxJ8L
dOJP1C3kwIPlYbUk/UsTZtinwGDArs3srmKQrcFRsa43hBZhpN2gnuoQXo8o2wzxv8Hu319M7qoU
in9Raq17dIrWjxznZU1wPMo/EyZFUMGfsPGOgxw9aBFUTnogPGebG7fHInAthgHPP/cRCnn+9F6w
k1xdMzbDIV/nMf8p9XQx6utlEZUPaw7Y4ey08B2hfRQ230oATyLQT9tNsPc3YRv+PxBvFbBOgQe/
N2PCXVVNcvb2iWVxvFL14iP62DSxwIOkQjnPODdqamFrooaIV6nmOdcHCIyCGy12BHBNd6ldvDQQ
LIWNsnJce2EDy9a+WgJTw36K8n+mmAg0M+zEtHZqdbaZfs1kELNOom4oAhey2SUfVP1GduS5HzYc
psSbu04SNLk3RwrLMeSbwmGJCLlGIsScwM8PwXDNIiTiAx+46UdMFstjOURboo/2PxwR5Tg76pi9
RU7iqxMfnnunlAfNzkRPdOrA7aLAXgLV9tjVM7M1gzlqo6yYEaINPCtb0WRyPAN6mMVBDhTQ/Nq6
yB1XTgs6tiUKmjXd+oWDSz7yJwe2rinP2P7Uq+KIRfFWYKIBYf2UO8Ny2o3elAjgrgUSmNCNHT2S
dNTWYAGjzm0PhdDVFdCoK53ciSTHeCp/YLl6rzP99FlS3Rw8kUvXonmRc3hlKcTtEZyg6/F622er
x+gd4dHlKEytuBiXoV/DmkGkPorlnPwA/7HiTbPz6sJDu05ShSIlvdSjBJGvrW25cFohjQz8lNB8
vp3o9UMNowb6WxLLfXQAwIs3K/a2+8MAAv+MkqCDAtjyhgLYrClydBrrE9TUry4ad3Ce5LJ8Q+xz
HemfP8ijjZmTkvu08lY+D6qj3zTcMu1SAO4u0U1UU4Ml3c8ytiGzT2XlhyO/lnyFMSKJDR3Vn64S
a62QH/++fC3jP52iDIz370cBepCcfbmApz380wssjf8ZyM4p8qV6IGlMPmTWjXqYRuTAfNo8FZ5d
GkxdwJLMzdZULtgmk3KEF5ZH8DrKUPQF9/2D2aI5cJp5a9h16XgCn8zIR9gtHlVmyGMNeYBsBJyg
zDtINTZOhOG1bfL8NL/oAEKC69VBpFHgI20Tt8rYs/OWs5cHUFFpZuzyDUbbzx96bFAvQOPUq+nQ
BBPInQo5KHFDPzoKvLHa71IFQB6uAIkqXumqq/Wpa6Ma1wHeBq9shPgNvoqqJQPzpN9gdyjMhiQl
wwpA/WO8IJaqkPPDRmjvs+Cpq4IeakSDuBD/AsvXjpqwHDbkcC2V5g1QL7MBHUCqTkvusqXaElLL
Pzx4TXJBjeHw49UCosOsAlMttzjb0pfHet8cDRbeAxaltGntQ/kSDa4oHITlyfGhu5sm66Vd4RDj
SGPKWX5oL9c7eGDhSrF2vrs1TWQcs6kKWpJa6RcuzYNJ44Zk6OpzfQzfSfz4aAlvQCMwmZVlUYUy
5Fu5hWwzraLB1hwQQDeNxBRvFqQUoOjdGK2/3ccmwON8igby85cGyCow8Ojfe4mJVSvBbGhlxLE5
wlgQ3BhYL21+EHkX2eSPCvIvc10HqIyIJdvghT2GTOqA0pST+yrk6Lnt6W46PY1YZjr+8ORppFtJ
P2tDEHmz0zqIrDggelwmH/k3vqsVktVPS6iOY0/4rXfwwFVZ2kvmGB8KW6hXoc6KWS16r5jfUrGN
It323i7Uhl2iN1m1zGO4LR0gWa+dplgBo2Dk1NDO/hhfKqHRHazU4aJjC5m9Im8jbXC3LPVE8IwW
zrTaaBZ+8Meu56TOcNDnpurKnh9ySsjtR8V7rBkEmARszTxCg5p4PtPYSGqVWgCSr0/ROmVp4Bez
XZYkUfVjF1cXBJBExOsazbNybrZP0o6AaT4UY78WwxyruCaXZ1gUNsU4tumUXvOa913usQY4064v
6e4R6jnLHLFb7lX+kbHL3gq7pOSDEJeSGj5GVPfCiUuZLGe2ESCJO7tLhifaaNGyjI4O2AIakJ6Z
tuXS3Qbdcxj2f2fdFGRflGb0ypGtimUsnAqOdfJg9jdeMbhVWHuiL86b57/xYQtXBv7Z1XN7j6CL
RrrudGcMPsOBtH9R7H/kC0obLK7MRaebuxb6iG2XO0zDNpsX4IY3BWYoFG62g1Fj71QWamMJUunp
7HFXiXfMlDIHUyxNyhlonbgQa6igXtk306ElwDo5DkBWPMDJAgkjThNSabooFjw68yRgF+k96jsW
Y0v0lUCoZeLhWNUBAq3eFMpJU7XWxw9E82WqCxwCgzJ0qziejmjwW4IE/zkxnq2fuZzKGLU2KuAE
dmLLCBdYYoezw5bPGK+i8pAExIU1qVgDlvfAB2E3DNb1VBH7Jb10tq6grcTyOG1eq+0yEfHNmnjI
EQtbvmVP8TMpRXTHotxe1+Qh8dlDaAEgA1cG5SpYO5ORhlM3WzgIfIdTv5wgLQa+mkqDCU/xqNK6
0n88b5BkYKEp7bCqyU034F88q8dux5rCBsUsLMOij6alLOm8ugg+t0Rnyp5K813+2gOf1ZOR8SiS
jByvPivPc1d71z8o5vqp0Pydt4qpXi7BRdbTcYuK/LyLbLYJmbBd8Nfs528JOqh5RJ5G/pg6zD8U
/FofEPHhS2X5XcuTVdRj3+/gCBTPANL8d77hWfbqeIvi9wWGeZ6VLUVf2TcetXrGce4chOi+7ck2
1C/MrdbHjohXRchMpzs1DYMeGFe1/wlIyDxNUycoNgiDOKQqAuIB8XxgksbVKfYFr/lX2Vab0BEY
WWRrVFJNLjXXER0WbE0MDOjQdhBg6v8dYWEWEhpgcZ4X6vsYhpyoNsYYLIIf5GdIi0ax0UHElPf7
EPTtJ1J4mHeZWJbz/cHyRZKPSL00wSygThJExpgkA3tcjPJnXKbwqPkMf9Xlm+vxdkkSpMhhuhzq
086JYXnV1gdUmYVtioKQpXzP0YFb7W3zjz8qafGq1ZD/KA5KSkvoFwHJLSw9FJ0pl76K5DVn3avk
2LThf8x9FceZNJksPBtcvHmIY9NrOvjiOovv+bYve1NU+ipNOmAFa+d4+pJwXwzKcyWGnO3nQDsi
ihW94F2WF1GvzX2FCoIKvCX9E+KV/eTkWlIqoTUOT6leY9WtK+AiOQUPp742y35Uf1oR47crQbUT
3iu00jW1/3acCwyl15cCyWy9r9sLPdTVk/AvLu71/GBdS++8IpEwp8sP6DwKnAYR1jxPSLvCAy4t
HOuAx51HJ4BYbCQIEH9cRblbdfsNwkS0v0xxg3DvYJCjbp9CH0SLniw2NJd1Sv9vT5fJzNjFkLRq
6b1av+H+IRywiN9XyWDouPzRbSSCtWJV65pNOv0hCpyeL3JfBdX3LNTGepj08JjM/h12x5XqARc8
On1D60WGC/catHEsw88ctjH//bH7BPHm3v4z0+uEKnPqR+D45lM8dVdi4cV0J/YzA+Mc485yfd3P
+OOhsyRcnj2BpM8AMJq3GUfKiovitDXwUQqd8Dnlsj7UVoYxiYmPb3L6BYjjSQmGfh4pa1qNcigk
dHMGVgbLOlI1rmph1SCjiArQVcLLAtb/urGPT4Vj/kGQQcQALHfBHELnUDTCtCkb2/g+JqmDeBqr
D3jM+tr1ODJqbCZuNQbmKeps4xVqsuGqtUjJR/6YSTvIy9TXhKEonGcNA0UZh7DwA6hGpKbnqApy
DZF4l+SvhVimv7ESC8jmDBOH7Yu3dk7ibadqZhRVXJtxtY1OMsvZck5o1QUpFdShNULiBJ/3o+vh
+iDUmCJcYBj0CsngKtJPoKoMXsz8Wpq2r8T1n/43oD4MBAK64DubEpuPXv/PPJ6hbmXarx+ZT55d
8s6fALEJwr+DvbBvx4uz8YL+PmHOaV0Z6BGkbXnok0twzfKWa8FjN2LItY3bb7HLKW8+lilDru1m
VjNqlQ3oGL2xWIMZz14qV8bJQmCRnnOPedkGxySdHxCL+xNx5Hb0vL6K0QgSHnkEKeSk2sOBZVR1
QEM1Oz7JbNY2ckUJ7PRUfOwbVni9PS3lVciC8SQ0HySfCzAx8gp2efm4D9ZgEVERUJkM+HOmNSI/
NeYcJ8tl+hTdF+jUXxr9LL4U/AlrsoGO62Fhjzwk65GmuSN0DX6/ib0wzOkqlUBUK7mP3uoLvKBV
6SLOVDCE7GieDZCtkkpQEb3unGuPgp+PlFX8vepl8mkKDbSUyq97uXSbXHbaUzTUBWAwO7VJLnuU
NDicWjWmTgnCAAUo0GxpfRFVhSf1B6UOILNeHYh34kRa6NIF8abSLDbgFHJNWtB6nDTg0LqDQJi3
1thOd1xxj7r406AebbjfixVv2hgYUfzSX6QQ2Y6as8owvWbusynTc8PVI1mH8L/YYaeENk3Uw96+
0aMlySA0Zy7QWq6ZDMpnhZtWmkdlAJuSDf1Eb+sRXER+QighfWXfZ7pl4aLhe++2jG6jHcYwD4OJ
68aqnuzgOT77rPddI6ulRWan0hoDsF95fyptmALwGPOxjqMI2MjAJ+fWUUhaoBwkGpKg0jrPMgkV
ExHCh/w5UAJV3IZXGyPIWS5qSzQ/wGkkkLMuigLj38leN+xY+hVbEtffpMfZhyHNYn9ZWsyeGfOd
+AZxSt/DowC4l8s9IDczZ9u2sz9WMBYEvYmIoLqyvfIGvv2h8+AFLERHK3At/sxu8esSTuAHtvE8
EqGKLm69OOBQc5xiecSnDf9TO87CUCNJUCzWZlL+/jNy9p7LN/1wB20NA1eWuxaa+KNu5zWisJl5
XZVEVkwaW3ojdOGwN8ycduGKOxBSa1svoONjhlCZxLM6eay47Gw0lTUzfKKxRg/31Pz9pD6DveyT
28cIgn9HMxCZ7toWTQZMTTHtlWag3sQqJkdDdZvFVRtBDb35dzQI8haGRfBQ6crgWeiOBRuNuSAt
RO/+WO2gl3miy8gooQRTBV0/js8wMPGr2z8nnPH/jIUgZc5Dz9FOsu+1ujL1jdbWLtlewEWNBFyZ
MFl+kMhs9fGHYNdtzKLAiOfb/V/s2Gh5SDdpx7cyc1bHPYw8CtX2a1JfXmzYrpsx/Uggkd/7ZKei
ie1fk88dvWxZlFn3IoZwraGW9PbGMhxMiAj+YuII/VGSgIsyix/PAJxLHm5R6mpjT8UwHItd6t+S
cuP9nF1Nb0xTYnR0ZdYFWHNbz5ZpkCLMNwVNj0yJDcfqdbJeasdz47lcl1bJ5CUxVrCsynh8C3gu
4Zk42hBQypy7TIoB1anv/V1S9gwZWIRFdB9eceU4HGTpurxwQwTU8NmrV9chfszf6M9JoJHIS/59
0mTH0G3/60TzGP13qRZcvR53nuzu80qfsX4HI1mFkdrrMfvufchqbgrTXnBVGL8ejd4IITrtjVK3
9nbhRfzpmMyncr2AU1g0zN/KULAypCeFIsz2g3xRFk5UWhisAVbzAr2kQrF76jZalYL4H43j7DXM
cqxWu6o1abwghQ4JcD2kaLi1S0I42/4ZRXCtc9wAoCQ/n6LweOOonboAs58WF0bkWrm9crAj5M/j
gLce9pVCAlNyJ3GlzcH7eS62qakmErzq9OA0pKfRxxsl5qESZJiYJjOsxkHC+rB9el7yuNsvqc00
aTCEgZC5OnCXpXntLlYM5w983wvjpyOjxU5fpGGrhbQrHZRQMoXSXTFh/qDcCXMeuMoCyjkE51QI
L2VRVNYmjsnF3zEKuNQl58S3UfstGgIDya+BWXxMcr8xE7g3Da150FwFIOZ7CfdWz83Cf0dZjJy7
rCQNQ3BIoRPUoVy2s0aqtxqJXAKXKhIbsGSNr2ZPi6kvIVe0ueWFWjLdThe4h2Q0001QG52+5U+3
dqvgD0mxJBcZHwbVH0mOYFFDMn6WYLJ0WWrqiIsHKq5u6eQNZSNO/t9UwJz2yTq0OBocHbTxxPoU
Zx5GpHY7lm8AkzxvXVC4Pc12TO7CwXrKABJz15KS7FPDTZ8LYJFb/phuHJmA6VDMOfGsYDj/5N6B
Bh9Nb+HgQHzlSAov/Iy5F5tDx7bus/hiBfIKM4x7IOwh9DIhoktgSKpsc6jYOIfgPPzcDEaWsYIB
3NsGUuGcvcxIzaRHO2BunFXOye400xVhegzHvvxpsvnQVlR9pm+0amqF0Jg1BV7U7xhDLY9x6QvG
SYdH4Qpt/d8c+qHGJvf5ccDqqzDD0Dn+6djE+Xoioz0YYm6TfoNaey3BodNty2cdSa7nDVx5oSds
jcieXGrp9s5IRM78bjZcgQN1SYvmvFiU7M0u6ktYxIuJrdrIACKqF17PVFHzed3HtU3ckxqLmw6Z
8tnjh4OcxkkLWZX7rC/aPoDfULqdBPdXmvEFmD0fzbCn+N4JKkKhbh5D6wZep71LgtPJHuf022/A
WHRnRfbS+lZabEJ3fvVmNSmHAaSZRYqxBE5wPTPkZ3rRJDGLWW1GrCAAH8r07TDHgg27k4AosDDj
3LKSNis51YtG7J8IRB/ICyfUuogfvkLGdG2uFG9S+co/ZBErBssTQGwL4sbHrZvj0yoPqplOy/4X
eTU8pI2FcfLnj/rruVgoIPFNNRdJtzPRKIQYBdhwBSC4W3iIK36zngIN2ieCvbOBqkfqaes+o7XL
hKuAm18jxxrSliCpf78pA7MicXIvRV9xT7mIMioxapAAm+430eZ9bk0oQHvKGJvaN/tHk02NlfHY
niotXt3wp9w1y52fI8CNLIZlkNMzDptejFW1hMLtD7hZ4RdlLWUtUfTicZ/ZRsfHz/n+qG8n+Ehw
0PCRS2EVi9CKezk9qZ+EBwbbTksX7bVU7/TRigckseHqhxU0CIEuZS6RytHhKnQc5lv1SzHDAH0z
l4wZVOkWUWnwPUp+3ltcQdrv52xQvrJO/s5kd6z8Ap4DzAi7W9XySI71W/E8+2DAZcqUL1Xg4el5
OvxWtOEnvdJCY7Q8EdrBQfX0IaxO+ghD1ob+hivgk5wTL7oJP7bYFT8E439agBRI2sMA42pwkT84
JE32A+ibcoiGFJku2VVbpoPQMAFlLu4CkUmlz0xb96R/A+q9kvW9krB7/eCJoUXGKvGNKBncmYpi
UNw60z1G63KpYyF5lViIni5AKY9JffvtGyrt6u2EtyGcM54RSrKN9YOjPaKXF2yLYWNfXulZGZZx
sfRNMX5kt1uplPUOqKGwES07/ocLa5YSasdBK4M+LU02dBlqGO13NMjJ+wqo+SL5xou4gpotJLmt
DjehKJJ8Ons/WcbIok+mZhdJ3FRFrqbjTzj90yN+rFuvyV0Va4EVD725tRSDt2ohP7MH/y1Vz51j
7W5begcUqPrxDixVOYDW9yn3bDU0A/xgaSrgAsfslS4lBEFVeTEyLUzpo5WqE+UPlT8Xc6wAGAr5
u2982om8l9rdZK/G21kgMXGBv2F+Hn/+HZeWpDpySgPdDfI4Y2Hm0upNEUKN//hQydudDZPK8sIR
lI8bNSjeFuDRQPx5iMgZ3bmLhw2Mn2DKQX86bcY7H+SSOXPUQP7xkTwtHgtsYzQVjmuusrWnu2hX
7Zl7mHv6Ksygut3zMUiJy/9XMRGfiybrg7zryBvTioW5s7mtsSPxyQwb05oASa0CtOqp6sCoSg2w
pFTWnguTDKO8NJE6Iw/uecw84eYKAZiIDT1CWLFv47hGJbfM7/a8yJBUceB6xhYYlYc9hlNSqQDO
gpernrZLc/Y686xJMR0rT9HY8JxpQSUxVNqNe93Ac7yKqcUGMXiZDiAHxTWyTyWATT5uje7myeWR
ealgFAVafh4kar47FJbH2FbABRKkESGRyJo2DAHOP42/Yy5G+VLetzNCAYoTHEiqrlOSNVdJB7L5
XXWqER4K6/LVmbPljocYBNdA5oFdc3xQjzkI4V93lkQcE+o/pbVEvEIqm4s+1jmttKriB3JJcSqg
e1IdfMlmjSIkeUu1cSFvEHUuL6HgYqXzuSevBxgW1COd3jyhLpXgXvmHzBi72x497w69xXBrOw0L
UowneVGft+mBh0aWdGNm1toik2ObjOmQjQLZYgcf4JsnLlzkkFiHI3biCSxE6Mqcqx7+KgGvUN0B
/bX1mf8hm8rS3RMOe4qoc3dHj4Jk0PKi+0DzHluK/lIjhpcGmSePgKDEIRZ+ijSq8BJTo1LHI8Oh
vE4ai7Lgo3HWn5VB4XRrcuR9zHFf14BLZy+DgViubIXnkQZT2chJL9PtaUN3om9pNgZOx3CX5FqL
l5YHD0lsxFe4ID8fpH/dqhCxr8LmNypk03xfnTdt+J87oVGvEytWp4JVwzVxyaf/sh/0rsF3MMaa
7VG6H5IFNHdF9q8T4YEpy2qGYvhEloWmjKsgam10Bzx+R8t1A7BDzh04zLI3TR1fHC21FgxW5nbn
UnqzjQK5q4SFQh028E8c5Cn5VlMmy1tUxakCxw8liaDiJ/yyRPCjG1hlGLADk/MPq/xpQqcV+Q54
3cb8nww2nt+WnFGI69NosaEipJ2MdBQr3tXy8+zyZiqDIvIHA9xPFw9yw/d9b549BnKK5rSKJGuc
7ZVy8qlKAZI2u3f51aH2Ve8vSX8uVf/Ip9Mhn65Y2oDQZdlRLE4IAvK/zDRy7JoDfOD15IjxYB1F
qFuugHZu1gC3uPHecEUvAQEn9nFt0hWd0wQvH5QeMd47yh/xT1o6p0LRHtue8pFfipcVBlR1AWlm
dazo1rdy5rwNBK4XM6LtN3B7xEVbbAngUIG9dyC/GqhP1E82Gt0diMk9zd3r8VsATC7HIIzmJUdn
sJvmLyU7nAdk0jXSjgkowFAcXlsDv+9h/yZ5kKRPYnTbg8YhU+S9dNZEL2DC/QPmAwsTUzhsLJui
VSWvxn8vBtcWQ2K2+n92UOhqNHCVVqHskwoOWLixGXWP8WBI0lWeLQbwaSyKmTQoKZY/D8vGjVox
ykVW9QlK2QLEkUEI/gAwcLmeOeZWFC9fiev9MFZdQa4CVfZUzQj87JtH6x5+v596pZIy6ZCR6aOY
wINh9E2yyCxiKqoAp3bwB58SlxKp5h+DKfayJd6uUU8PCvuGMyT7uIZqRz/Ga3H0GbsH8+PCpVYP
NDsJplhYChbSORH3BtuD6kdqCBqk66LIJ8e23DB+LFcJ3BweJUdlHWa5hP4rE/ZnQHmchji7hv3x
FtT7oXTLlq9F5OCeXsLUsZxETZrymvnrlKDypGXE1eb+n3ociZQp8D9cKmDff562Lhoqx2uuEJVA
cJiCUYNvksNJIfa/+9sw01vdA1OmW8qVv74DB60gXOZWMvN1kyUN9ykEClzm67bOgFu9pN214CMy
Vm0agNTdKUYYqF1kPptmxGfPZ9LOkM+WhR8h23MIEmcg9YFMP+RsYfYzoSV7FoHT+GDzW8LYZR3R
vDZgPWhyB7pYeGnnBxG3BOUzrEaGKgD8RMFieHPUT3836ux/QVTAwJnGojtkUl03wA/k5hgmWuuJ
kKSERzh4zQcZoIpKHQrQQVBaBBXDTR9Sbjjpjuvby39b5Bkpi+Cw/ZJIGxk6cluld56GbeyMGT6T
E9hnqA6hCG4EP/b5UIrUsBX5t+T0V19JMI1FEnVjqJQgB9AMl5uywJj5WaMDc196ZvOA3hwCKgh5
ahlE4+pdO/vA3BVhFDWwYM7hqxQ7F1LoKBIGd1qpbOqJrFXN1OaBMM5XnOg83iADOoawd4dayVGw
YFy3+JWby23oXaGWaCMI0S/ak1p+T1qdw/pJouoh+hTn2dA3EbnUbXjSozA+BpO92qiS2dahPUWR
ZMd0cHZUcHjiImAQjXuHCgMk5ZutF1iBD82FD0yxkx7/0AP0ZsxKb4AQddryQmV7jBXY37Rrnb6M
62dbIiKw4v1HKGUNp3kdMN9bC2I9qIiC5ToS90wt4Rsqc0S0Oq8PH6/nTgXkez2oTwNCzcQSzEP6
W/FeQie00jGIM7jniNtjliQnWZUYI0gBvBCzJNhmKQCyUrHicvVuvuevWThVw8VvX2TKGiMD/P+H
wJRGt3gH7bKQxj6nE5wIxV5szYem2W42K4QKGxMNI1tnFbvuNIUx+eLMQXqLKtvj9Za/qfXw9Zds
8Q+y2jSTSEMPCisEC/241fnr4f9jN7EuEi0GPYokI4HlFqwbYHPt6+2O/O2QjzlDaAyvIlDtyuYJ
8CV9R3y5I5lAOrHJkQjgV7QruOotykJaJynj3W84ksydazwB/KRYsvgiQiGqEgnj8BTsgXPIHSd3
b98xEl1QPsdD2cigZhaZfww9LnGhdw3JzOmemzH8IBdR7JGNZ+t2xUp0KnrAZz2eoeZyLHClbPag
K2Xswl0wAyFvpifmtcZWdEkLbn/w7PO5veR3YxGB8RhpcbJ0LAlEUfNxsPZ5+KjtWGcOLEuUlxyA
2KcqRwJMsw0zoruCL10+vTfwaqV4U51nQy6PeDimFKkm4k2k4LHy/tDcV8fpu9IGOYiU3PJyRCVD
VxtJoWHggXJLhgx62J2JzJNCAhS7nk9Ax0oEwcjwLtVT4Zm0F+a8os0jfNiYp6Z/un1gdr0+XViX
STokG/ZFNwa+xfyZuXmVQEMYT47P8/J4BXPYuzOMYgMxbsxrx/8Al1Ix3tiRgJ2OgcHtg8rAh5VB
4A8v85+PVSH6DhTIs6oo1I8y4ne7peZLuSR2kGcqinkt0okDy+z41AiC5REW/AqUsDCddH/7ShPv
eoherDGwdRVPOJ0O4PeTvO+wZ/5xixnshofLV7GufGv5nKJvSlbPL/8aordawOroAnnCCsseOO6d
p/ql3+BKCLR1T7760XKhzrTMe2ROzhAlS8Gbc8sRvgMKErHAciKS/Osjt5JMeX+WIgbWOUXfzrie
C9ZIV7V3zIgd8Chz6O+RhNCLHwV17lqHC5rDCb7G9Z26iZL93/I2x6XrL8/lLCNU/SHJO7JmGjeD
VDKpw5j1z+CpSL7WtTD9/NqhA+8Oju/0msSMzTf4a0MDIpd9z+PQQ2i+xfKIDVA7StONVuV9iPyX
6vK+r5jKeYlk3JR/h0/k6M9x45qusm5gzZ1spgzaXAzuzhPVcYfjIFpUBLhvY63BScNEr8WrP9kQ
OujlmJ4qm0a/p3wNlZcNDx4oeEgIxyYKNl6uj9x5ij0PjjWTBJNes0W+dn9xdLid3K15y0u5dmAA
DlUD/85OGckZx9ZMHFgZ5WRjtzwaG2LBpG/EmtIxng9o3eNuXXAJpnd7cg38DoKoxkciIreBNalq
5zmwWhYDq0GaVbRaKlukV+lk9QlXGvd6Gs00rxkYQFWVknLtzfRTc6v5kjbKJPGFCIAJCV6xI3X0
KrTSmPk5/vHOY17uIYdz+lF/+f2xswkWtmTpNRMF5eAiP5mZ1JnHXZsP1oIW84Z44lEoG6L/fPHd
QxuxgQYmffNrEdtlwYWIqOuz82fGDht+PvnWPri4PIDb5SluLhq0vpukgPUfzdL3ebzNOMlgrnFO
ba4wdtuiPB3RHt34+VszY0D2rZ71fzONitx4W8HREDwMSJk+G1y70WnfmzF+00h610LkL+dMYGYc
7sQ4QEy7Sm0LWc82hLRXiLPfucSEJSI590xCipKCqjnQIDq6/usNOxv7YKMuLDW2/AP91ys9Iy2O
RTRgwG9tPTpgeJHpuVm7BtEaCRzwzFNl2Hj149TaJD8T26I2Eo4CVNc8O4FNo1iI1kwijnYOLYy4
d1dj/F8UUIGheTp2pu5wmSyWPt1TrygDe0EoiLe/bSlkDmu6woM5GSPQ3lZg55HkRhMJfjHcB9ZC
uE+VGjzU3NtR++hKHGOtwGB9DH+Y9gfLUUiWXYHjyLoFdPlVInslmmabIyu4HJdvfvRxDA4zaEt+
KwHy/WzwzSYltjL6AsWicYga3LUp2qDtXRFig13ajZeXQ/sUaRbzD0qVUbScRT+MLgDFgKGzkANU
tGRJhPVJGQOWXD8+JOAlXexBubksFG1R3Xud58zjPx6JAfWUkExu98hVkqyVhRitGBQz7+tnZYN7
evmf+TIt0RSsH9oLG0x5a31q2oKQEqBMWhJrYMfzAHNipToKEOB6PruM2DS8WnwgG0apx19b5G6M
IJgDcWmxwzCT1xdAxdFZbX3k+4Wr+UhMtUaFj3bhYxLu1yZ7F/oJ+g8CTPK1As03TcI5BI3XfDYF
7Rw1ajUXQcxqA4HclGe79bYuzPCSBkjBF2MJRhuUtLC+DXnhfvwZGd5xABwIzkjSj+Sez+sa2ldX
eaLLiwGqOdU+6rwmatM3ts4Hyz7Qe2mfKyVZv/kCrXVUccAoQ5Pnx2om5vBX2DNYMVUCrrBHhzjB
rhThXynDXv6ZKD4KKMiIrcuRewjRZ+3rCVEKp9OuHhgJeOsfwE2vdNqn4g4S0xZQ2y7WKk+lOsQQ
XGsqd7OEL8zSB+r3sFrMFWZ5GVXTSnJk0U5AedJ2TBnBsrkb/2Vp2IlmhLzEwMrMZYBGNTM4gORW
dskpLCQ/d6g8q9EzgSweMwNj1GveE+0/haDIMHJb2aIZY+r2S77WH5Oxssye1zmdh0GkyB0bVJaT
m4ixrB7VfmjTDxHIdYyytsrkeS6fo5vrKp4scfyFjOq+qxAqClFeu+ox3yJne5YaD1HD3GY6ZBV3
FpMiwQkrah0flZyMKMmslRMuPdVJkIBQW2uXY0rVowmJpNwehi9699Fq2/jWpw2AJMcAVLKRvsl9
HzjCkgLFv1VVJQm9jt4jrIF/qIY7s5l0EAHEqUt5953L9pc4n+rbAgqAR1vIMIMjuOVFhujtCJ5o
7PV0nOtzbapE6f7pxnqyIiH2PAESafQxwrhQrEFf587ew3Q6LYGFB8gGnCTYndPNtQHBRvUnCBNv
YI2FHdyxhpOYXDUD5BWueClFQE2YkguDyv4pMhCdf4KLfz2fLjdajnMjyzX/lGBms43Kndn+5oTZ
w5MG9fF11jNoUP+I6zAH0AIBZtpb/RRwsw+uF+aNylE6DrG79GSIsJpM4tB/gbq4FfwdwpTY26Kc
6BCJTkDzV02WZmA2jjFVjK3OY7lcY6x2JxFYk53t2iA2EXrUSP+N9wjooTBbaupVgUUINh1Xe3ig
HdvwrDV/Tf0s4q4dbxhMixfpR3LTECeuub7/xo4+549xDpbteRR/Q97yjmrFDu4+OjrfSyiR2gVq
XBn9uO5g1X1hIOmIl+ozc8YoeeWA/L1uqDW6orLmZDPP79q3/ZYYy8opljt1tRZ7jcvmPe6eBYU7
hB7PzRMGYVWDfsv8TtobyOfwbP1ilBpwoEdkgYQLdlqz2AXPLoqY3iE2o+veznl7HJ0bhCh1txif
4t71+8M3AMi2omxnCvPHG2UT5BQ5qe2MLbZ7ukrFDE8tfA9sOMCIdZIUnBbbKU3en6ZBCAnmvh7d
V/++NiPfjZuRzpJmctJ1237/Y+K5PUkiW4oBArwiKLpZugSPnA59SuR4QCY47q788alDNM2SGThV
Suwa8IcpAVbsuUK7UwWJ4T/+hZx2Jf0WjKYaEElBT7WEfW0hA+uWxZ6RWnzcup5Do0N5eDOi54qX
L6Yq/z+FmUOjaIZvSoAewFerKKDVYHaD7besDH+ku+HelTI9wfCHbS+TNgsn0XbH/XGRyJpj596k
E6FkkJvV1kX9LpdX9Qy1+YRkNHBL6mRkB5OAAJAAB18gvngsrn7hwqWiLvycCGEvskhHt1ICBXmh
oHfI/1x/Dboy2bDhsoyWUQ03sH2m9vmh1YhSy2vLP/Tk4u7B21EkEB64u1q4NNLUO81tugLOa8sS
84cgVdhgN7Xj4HMnZqE6OnLEXVfOBI1H7FQi+YzvBzoOIKruoqjWZTxJ4hmlSsvBOE4UgnUju9A6
u/quRgUejAdQzuT38LurUFzOVMPAXwTbvQz5ZOc/tDcGImMSGE21hUHA3N/Rv/DwLtTERSNXmd23
AAl+aiOH38FbfcX/oUrjzCQYWkfNBufB5ChSzAxskc2l1L3rIH3nh/vdzo+lF+lBYBIKJTp5iY7c
HCDDKfLjWTKv9nT6OOWP5fhsxBRX3NGPuDyLnCB4vp/qvk5Z4RcjorirAygnLczj0++nZ1HsSzGJ
mA8jADDvYqTaLq3/ROCs8EygeE27lLWztOrKA6WWh8Fmb7BJ2Yy2gwEU55Tjm2iqAmiUZI5KVHTg
ou4tFj8fWozlyOK1R6YEvbLdYsdlzsZoAoN86zhvdZ2GjRQYpxDIlBRNF3wJuChsTzu13z/E4+VT
WBcu2298KUpwxcCSyve2K4JjKgyV4bFZNeSP5NL4lKYkkM38NWodmGwNLZ9oo5Tet9j3nvfJGn30
ggjjEailubO3SlFcYoUvz4IttqUALASSLlewpAi+59LGPucYskn/FUCNOLMtToZfsyNYMtIDxnCY
aPZwzWQgRxXXSV2jh67e/f2s3btcu83dpKPhbD+1yN75Q838agzwlZRN9Iyv8qeVL4hNaJBCiQqy
jOxVOd1hz+E9MpcyqWyHgwRnXgJOL4uhKWv8qo02k0Xf0rQYz0pCgmfwjmpF5+J0E6QJ40npUjbr
V6R1LVeVlp8LoWQ2f0y93Vsh5/mRpVSkomfl7hBkihrh8LbHV3mMrsvhpF6YUGzKVuWVZ8vX1tVe
2S3n22kB1IprHMUpy8FsfuHHf3JrX52mb+LsXi5jQWqWCbUp3JYRC2r8DddMgghkaE4ZxVnJlnSf
HZFruybuVbMEaTzM5m8WKSTxTEwOrxsPkAPU0eEsMv/XmFu/lKxgCrSJV7PJvIgi4yPR8z5M8y2m
tsZc7p7viqIvFwi3BDFnc+NnsPjgTfugJDPjYbyMQGW+sGAo76I+nSSKqvaQU/xXLG+qBf64xDl1
MKKR/pJaavGxWJCC5gbDl2YJuUk0cTizwvR+H/N1gyFJoiAwBrETvKIo8ywCbgNh8Q6tV18bmgJh
bZ0XGq8Z2D3SgRn9se0SJA7ShQQvChPfvfma/ivmBmUKh0Cr5oyDNyVslZXIqV8hrTCQaTHr1VRZ
vvLCnHNxFcwPQepYaWX97eXUDBwzWWul76sPZz3Gi1GaxsfcsCWRQ7VqDHeE2RCbnZHLx62xZOxT
kFiL4dtvt5MOMc5TJ+CmR2YTSgeaKwZ18irCFiYJkPi5c/6KrNdWy3YXGBs2Z5VQMJ/GEQfwd3bC
mE6BR/Zc4m/4vRPd5MEABOJT/aEXCBAe9SEVfpgRBuVyf2t9qZJ2tG5aXLVxN2GIspSh/s853d0G
UdHNF0YjSQiD3s2kWyTNa+sKppyHaZBpYbpvcM3PdnirvuI2B+QH9Z7k8OimlDU5ADTqEZtkVXlF
1VM6h86tIP9/8D2fugQzNekKoAIs3eqR6dmgptm3Jeq+t9tbGPRerS/MIQyPlCgpc5Svlqeu04Sy
WSkVQj2D6Y8z+SyhLqytTLr5Dm1nGfLz82bhnroppp+gnSI0LfuU07qkpcKfdL5JDmp8GUP05CkR
1uH4uzE/dIXpmuclxK60uTVbCrKQoEZFFg750SBKM4XUG61vUFispItKOO2kkCDmuldGkKcxg6f/
+Eo0wC4GCewDEOttc4PR3LvyTezEPrJo8p/rEytlTCPAwgGL7WC6KfHbWEVSFOkxvvw+2BFEGfU/
zrWon8oGv68lhcM+iJbBFtAvbeTt4z3+CFJm5F3OhZooD+sQpCMbj5cBQZqolPQpRAnRLcyeESVm
DjXo5VYeTMViyohOJiXkI8R3PQzke6TiuL6k3gbmuRT2Ez7/iL9/YpHB89UywiMA0Qp0FRraGl2T
Q3yI2YP3IBVdednTqjeC8w71evOJBLJxepcVD4x+l8Qgt59dolC9Hz9dkh9STBXB8Cd7bSMHyzJE
TQjsv+2cYvUE3C+qZ6D/bQLrwy9BjJ/tsX0jPlYe2TFGZqbj7JHyWU51rVZ9mVQWe8/i2d8mbkD/
DKemgb09l1mriuxNzEOcqpSJ8Qq01ixYdQAUEXswyO3CHMGF4da0hV68DL47CZDqtdIjPG3EJpQj
vtVSjbtt8jbClxlkWmE58NGIjgE48DLQmMe4mVM1oyHWKFPxw9V+H/8q8h1F7j/CY+b7g4aFlgrb
9JdUu1vqBdW9WiGkeVTvl7pWYBITzAneeM1AQypepF/uDEMERR3wx735T6aeEAi33IUQdJkh/Q3N
B0IgjNfIHu78ahmR+4r2Iap06obYsDg8Fhy7ATJav4FI3ic9gbxONH7YhpE8t38v1f5ljJ4ydI2m
1Qc1zHtArjfStoIsiXVg98A44FAS05+JvZz5xt1FtiTh4BBElJa5/RF6uJlrc09A7h/uVsEmedN5
1LwjgGbsrJYTzn+peVzTLy3aZG3Lew4MK/Wp5GYAvGrutCTyo7ptPela8Jkf09PEDza2cbWgAPZ8
KZ2Zhsz7iGL7/sq7tNHhvX/nb3K0Ql4AdHU63eH9ECmorsiDhG0wn3Zw4lO1Gi/rf9im1zgivhD+
0BrZPYm//AY1vaaLlegUIs62ii4LNMc7S+eO0vwmwauspb1aqkedmrSYEqDGi7d84V4ZQSmNlycG
1xY9Gl3RynY7AwE8MorAuUPNpqO7m/Cd6w8qIhJjdpvBwXeA4ztm6ITxvVQlwrSae869ttTToTI+
kI4BKjD/Xbr52NczcO4YIWAurZDHUt1xPxVz26Cs6bXTd086r2v1mr+RT9OqydxuDw8tenXPB9W2
UC6ZKzGZQOtarOqQonMfhKaBa1+1FFDadWuVD6tXFEFXa0cKSSU0w7Ui5Cq6cVmmDrEOobNg6ZRl
b/FA2qjHTXKYoI8Aaf77UCdGuv6Cn40rbfVdvOjjOOjSk2ntNeEu3tQcK/w6ROo82JlgrS54oanv
e8IypSgFPUkezaXBRp22qI/i/Bd9ha7UdL1Nzwc1INllkvdPPzMK1LaGcwbSRymV4LEW2fl/BOl8
Jhia/BZcByu4l34fxgpZoRdHI++uGjYIM/tiJSgn7lmdjMyZnxSt7zMpbvGx7yL3qBn3gRv/IqVY
N6Gb5CbN/MaRIMVbHvxR5m1gzHKicNH+D9WwNVeHm7eSU3TzEcKZOD64vh/IMQFBy9/1gq9vDN+Y
1N45gh+pHC0P2dFSJZG9imAk7Z8MX+oZf1NqV5/So4+FMJw+eQb+wVDhB4QKDkrnnJ34qX5lFi5m
Qi2TK76R0HoYBoAab+WW5725259iNnpVkgAekPXFQF7T1bI1B/eP2R3D5PazBFpX7l1in2gUUc8n
edXn9q9qZP6uxX8khRzm5EIkTqHizRwxbVlMG9MI2Qa8a3YYH4jZhbs3NFpv0qTx8Sikm05/B6gO
Hkf2k2hkL8/KAUDBGTphBnukQBXxKv6jDtKuT+4z1JrgpULMEPbeTgEvr/ep5CMuRR+FtFQzdpxb
JubZF4C2qBMxHRjf6IS8LfdWgVYQSO6cOw6QAx5VQR9QS1QOxSb4JlTSAgcRq+XkY9aaRVtqFWRJ
fbhPhc4UzimjMWAAvpGjwerVRuvEOCZ2XPJ9oD62q7ZpYIP4kv/IR3pbCPkplhwn6b8RerieiZYK
Dal81ziduZd+GScn3fmdxASul5xSGZfP7t5uz4atbjpAo1me71R6X6xvx9AL6T/uZNKzDax5s0JL
eTcDZhoULemLwAZFPRrpO8v7VFYj/43qw7W9Rxl8TYRcUk2ka79GDl1eRSYLMT9tvpzPd3Q7/0Rd
7lCQz0d9TaP1LqY5jUJm5gkSZet6+MyS72DxE8R5l6V7+FuXuJ4qa/clg3EyjYcSrAaEutpfAxP3
0bu8YOOVOlOv96LSaOEPf77EEMl3clUsh5Pb90w8Ipkiv2ex2TwKAlsm0uXChIZvLe2rtGXj3o4U
V+qtnWyKT4J5PVF0Cvh3T5iU4/aGPsBbNHiWL/dgwRccWLxpdtdXQzotVjXEn0cP/YWgO22RrEkr
lITclY3lEs4aMTWNx1kwUBUPwY8/vVMQwBVFaGqL3lhw1q1+Z7Gh9zQjDnNLZwLAyMzvUZrv/D+h
7XgxYoVI/s0TjqHxsn+F4r7JClILR3n6cGniDRt1i5ElyuKS/K3+z6cQNSJ7N5R/UB/dZVinh+E+
+JguOOFWI7vLzzVdj3MspwSdTuSw7DzJqCFtkmNhCGXFj9uQnDgBmULmqSpUQgkS1PAPSGbky92j
pjLlJkvbMsYzM4/1/fGBMA0e7Nn9bzX04euoyg7OEm99cHKAT0GBoq7nQ+TzXgmTIm4f6i8zQDj/
CcuxavS9pUDF7rCH1qrs5tYk+1PwUXfxr4omNHvYI/O4Na3P9o1RK22OCjdrELoXfFvpfMjhvRI5
eQPOOfG5/75IbhY5LAhvihuU73DXWvqKDC22aHQtUSShKl+hShn0ENJnsPigGSoyZ9G6B0QOGnCJ
DoNelfJ+S13oFV0w0+h48UrcwTHSV+7b/IxTWRX570M8RJCXc/Q6IZ8+apGG1I4z0shFZvdOS1H+
ElJg0eEdce0lkTv+e6Vmg5gxGMlCyJ9hTyK563TL9X0STrAmcAMmKxr8v6ahcNXyFLtWv8S6HC+7
17+YjbR8yIl0lhl1jeVhtvwNqQ8jWIMMSk+8pVVD09hTgCk2jsgAb+cuHVnRjeRq12w+r8UIMlqJ
Xq5ToTojpIN39xaOCJwAyV3XeQW/zIUw/SgrCABljmkvCwb3+sC/DjQd0f9kp6qiUfVqJEMTPdOL
HH4w0jrzBaawNJq5ER+Gk8yMTjLyqha7zvmBUvhi2QIU2qHNE4zPOLLtIcvjy/9fZMQ7tRqyRep8
I+/Xl7JKlaVf1hm25seqM3Afts/u1cjKG8qwPvnaEXERqr8P5nSv+MclXZKVE5DXMgFrRGgC/GPb
gfQ6krgnrVKb1dOyEGNJdVlgB6lp4cMvS18fOCAyrJOvlHw+lqXP3vwS3pdSZEsSariamSapnUNi
WRJfEn+asnzabZ2c0to190XgcaIFl/n0v0tYfYQwbnfOT4uDsLjn4nf17usFqOqsR/crJF7Ey9Mf
fh4uD+8MQF/D0CC+Oe58rAYLI8VsiNA8Mk/V6O/CGOt31bkVuAGbGHwE/JffRf4Xqh4OghqDAk9h
ITP7dm+KD3Y0FZQCh5G+VsR2rlp9DTNq1549aXqKrvqkjPPLwbSeBBktrRkKy9YN7De5XAMidvZ6
NLQWwvJoXgRqSceSkCKW6nmNezrN36KgQfjNve+ZgM/XUiXmfGm13Z3Xw+gXIhb8uzMynq5FVDVf
z7pr82wwzyLeadPxe5d87bb4VUCBZrV2zGHa3BKtxQb9wt71Ey+G+DuXsHPGFS37Pidspvjoqaeb
guaNTS8quTJtcN6YCfAXiFwC5TVjhZtB+th2d5vhhSElK7iRsvMyMaqDyyoOfoKsrEJWz6L3bhUW
5BhQtj91lJprfuxa3GW7SbWAwl4duMhqE+mf4zZFVFuqwBu9sRou6kfi4mF6jICrw4S2MTX1cf+M
7LQRb4NKPoDLgH2B1UV0pzcg5WIavO7Oyrf9ABV+dJ4aBDPDGSgrSrqUJOjNeoZQ2GOfz7QxPtyy
e6g+A9Uj91pJ63TxXd5VGHUK1zmCtNerkgsNCY1Q+nfNELqnpmMJHgMCARs6kElgkwbwOo5+drjG
0g2pC7SHw6IaSvkIZGyUyEcHAIX+sMdYNpSawjQUZCME+xLxAr7JbzQ9FePvNcRIWxxyLnSK3G1j
cUaMsgl8YKkAnwi0CLMYMQ4YUK0B32cCKrTypGiwOiCEpphp08sYbFeWN12+484jdgKTNBLT3J4n
en30V1QjS5HZM+443h6tkwiUpWr7mzzcA9FHMRgYoNPtZvo2jAhF8teqfZj6pkYJFO7GcNyQ/mSm
/eqxx/6udxBhFhoZA2dTycNrwFlq6QnLU7q8veoxtH9tufK+byKHMcatT9VchdUdThiRm6IsvCnS
WEElHV2flrKC9fpRlqwq/FgrH65wc9tR8HnVF49ADitN22uoSo30BbcalQ+ImeVQouhWDE31m9aT
dIS21RUGjIfdLQ4fwCEASjPRMuAY0JQKHgMzubuPYZN2U9CjSTvoBfUR6R3NZaQDokjSDlZxObmQ
i6iv4RiwemiH3VsJCvcEk5iczWF/DtLRb4aoSubzmv0ydzgkFmqgTf+A445OQjAzK7lo8JFgYcGN
5A0QykVuWnWVHDhzhZnxY0ew4k/VyjWfAvGTm3FTPkt9zySgHyagl0k9s/r6DclZmooKQ34KkDyv
4SU0+Rnqv/WbKT40a7X0sKsxxak3duturrVCyhfGFBFVZtrdsdlX7HSsGQ4dg9jLiQJMJrXe1xdR
35KF034foqrq/hdIpNL6zP6n6FX9sVSKpenSnl26EgfsBokh1uWU+uaLreZv1dXdapvOgmOdFEJz
EwKS8ZNJBA9oTZI7jFVcsrsij/xMEHTfrUaaWCrMjR58k6mvKkqHI5/qF4r8TVZjzD4wgXNBLG3h
FI90APZ7FhMnR+jmGI0QmQabWf6rKaa5JnmLx7bIaCpMfGi/BDroLNBAYAm9ZlcUtH7tLpD7i2u/
pLR/fnIdRfi2lhUpY4laOM5MUvw9q1qFhc2v9ioXiNdnspdf586aBH+uhgGt6IDepty82ylpJIxS
pYagnZW2ogExQdv8scqTjXEIenCoKtpmirDqg3ugx7ztAvCpH8PbE3ZtoUmJGAdD8kU1N2t9hlpX
hg+zGEhh9C5n1Y1ioaFbCFjeP6p/G6zP9qmjp+3CojrL/dzV2zeibMJ4SqD2YNy5p7a7SQkKf4Zi
vqLkWpw6OSJd4A9yVVkKviMK56nDALcWd2D49OGVoGWvk214z5axc8xbdVV2spQ2T2qxgVgBv4on
SwAOtovoKy9SHl+BgR07qYLIv6K25vwNeQ0dnq4JYQlDsA6I9OJo5rhqO3diZwd2jlh34IymqfS8
qZF5Awu/zd+fEL1jOg8J8JUPqzpBBeco5DG7X/SdKyfBWBKXdBdwekYKqflh0uhfr4z5W1I845KW
DzGExUR0zzw22BrK1szyYhCjEyiaUw+2I7tCJrigfu8wh39pt95PWHjoHcdyhUFqOiuzRMUNa2RP
J18h0UFm+7EU2W21oi9d/ayjsqwAvUu4nEt+GmIWUbMIsgxKFAfGo+tfSd2upZN8lf6RQokqb69p
XCmL346sKZyZo5kTe3VzYhOmS2b/vst3RoknDfBy95OribD2HoQghRa6GenMe5j3VJ1yMCOj2JWh
k+cgY2W0nJqwi4lhvvClvnXrFkd4iPtwAO+QTPo4IRs3veEa522HbTlo89jxUlV3JOnfN8W5lYXW
sDtioiQXU4q4V0XM4xnGZi5u6eRqfXYybHt/meGB4+AUcEpl1n/LwPFSzM7vNrEBgEU73cegO76G
oODyAsxcUscrnTgt+DXFl1zQsfxatpfX8c/syuENkENfFFJGrBQosyv5oENiykecdxq7sPs8zXXf
/mTK9e3DRRxtCUmZETBq1MT19p2F55EZC/8NH5t1WOsmHx86scXlrfRXinyLNWm+uE50caqh31wK
ICvgOzRRMVuy8q3CLFPeLstHM4aNERL2LwVulIzhvlHag4jYHE2Ts3Zk1IdBOQdAiZdyuR34Jcbb
xEUrk7ilne0B57CcBF2cqG66uBN5nVO4QVRTrn4zhI+rT0asPEoiWZiawzQ3cTkRgIxp9SEEhnEC
TYSWefq8sVQ/33bopf980tpCMOKUkC2of5dmsSX6UbFw/YFo2bLuCYBrD47RL1BxLoLASE2BtWq2
BJ+7T2GEqBIdomwr9kx+JgfxIbGykrRDqJXz7oloQgQ5N/QhK7yfzM443Of+abpZVbOgA9X56dgl
OMg7caIUG3bY0WntQIuDJRzkHGHl1bzXGbXFNOky/loGfLZ7hliGVK2RHYsFXSKE8NrIKKMYGkM5
WtPC1HbmwrPtmdYrSycU4eepTb0ZkbIUHKMTHWMYWv5T6jHySgevEsrl9STQC3kHti+LlIRaL97N
fwpKUKD/ka54XDe6R0WEQ4KPLqf/sT9k9l9yWizodA+YWoqSLkiTZKF8HSv8HWevFQxwjLg5NNx9
N8hFUl6LYGVXjqxQK1ceBZFqNZV4LayNDZx4ejsarjiN1NuYS5XrdiTRQSn5NrpKO05E1UWBD4wk
JnkPdDCOOaVyLMGp9wavg1b6TzP5D9psUdLxMJXlWzE6ItA2dqF4EY+MeKcQNWr8WWUdQip4k73h
Z7PBHgUT2RXkH311DTU5EorDa9Htzq7C/VoDKU0mNr6Tqz1v06QMvUOASABpc3MM2Ix3r+9myP3X
Pe8/52dgjRNJgpkTKrSWOaamE2bKOLYAuvOQCmpidDK2PlJmDy1uLvuRVflndELqyY8PfFU4lGPB
K7X3hURmPAM94rbxEx0ORh8asrMfEseuFoYDWWFuexYMynVURh9TQiVn8nQOzyl+dFE3wn6KSky3
Ia69acz1nm5/1W8K5nStyFGFE7kl43YqlkryV4z83t/lsIlo7SbvzvFJSh1V74yJarwR/zOZjTp0
3WdsW96zjqtuOVmzIJRzbQbWtU5UdVRZDWNyLkgZGS1d66gP/EKik6ujEo/CqEtQpmei6tsauR1v
W7YWo2Wlzwv0J4N5qNuKSsYDY4WoECLF0XxrehRRwAbYJBtLNkft8Hk8OdlMIjU8kyS627Bmyc06
9TKVOswUuA5b2IraXNgWc+T/Q5g0LzW3c7tdwpp5Zm7bHajaqoEJIZg8gAIs1qWGmJwQyfonnL7y
4vAyfLj7aoeULA5vzaX/l4gKpGTQRrQuKybm6C4eYlcN3K+pCBoNxk/d4NekW5LUGYpC0BE1jI89
6GSe+nEeZ5RTgyHHfu0TycysV7aoiiJG/iMwZXZaBPsUknu9LsXECGFoR5olR9TogC6JqkyuH82t
1P6SI7pj2DdUaJ7Nhkhp7fCRsyQL40cJOx3y1H9/CiVfAFQwY6gSSCjnSC7sMU9d0ILhsW68OHb9
BQM9YPhNLLlxcoZrFBu8tRTWOgxqYUf6aElc5gAZ/Y9Yf+M1P09dUVlmrfpilXVg7+E16MkpYoib
y/kpAjTBrXek8zdwWgg1V2NHmm3cYHWYjVycmMnhsA7GEFlyge1Mxzp7DMhiE2mRI/czEtCucsjb
6fKVwpJ1PKm+3TUSmOY/SSuq3RMn4+bLmsU2bGGQ7Dqk92HmQFNEyoC6FeK+BoSHxtqa9kYXo3Ld
w51Qh8OkaKKZulOwBYF36B0fkf+kPG+tQCUs4t4ozphusoOWMZD3EoiDotojSvt5IkJL9bhC97wi
/lFXBHr5kRyJiBZBVFgprHEdkHJ3YZXhqczRItoREG7PtZXJX8kaZ6AGWhyqxYs59QUdeM8N8RJc
+CXOtrJRHCh1S8XwFyR/tAgdLzTvPTHE0Qe9PRD0hYV/MGP45OxATcylrwMcn5sQ44c81R/Cbfgm
HmoZEWvwAh+ppuc32HPEnpTX83d1bmbtr93eu5ca1v6OWf7BPZ5Iv0qKt/ZvKtwjxXVU32QqwdnN
4HfP85PtJaCRG6tcWxWl9JFukLTUYqcmBJ1FgZMwQ33y5Ns5fbDLeERBvs43iINi4KfaYbe78I8H
8F/d0VkKJ5wpNhx6gcmQ1RzvvoUh1YOlj+aEV389FYPBf1AkaSLKmHGaPuMlLmMRIc+ts4o/DUU1
9CkZ/itXCYXrMmqp5XYeDfZft4IDcOJ97XRDRisL6RGDmiHZEJAp11E1+omFMk2MOFbMcmLmPTUT
7KdIc+JINZ9N297mMTs6fyh3XRTVDqhnJhTg1CcdkZ2Vl24+hiuEJf7tQc2FdbBpn688SZos5wL2
nzVFUDLLCq4nUlAYOKXp8SukWtnI6sysmwA25CmmZP9wEHB/BpMUhVhkGp9oH13CaiIK0G5EAZl5
hLDOWrSL6NSiuheVIxSIGGqGwmpUqfrVUezhC+N8gOc3fdHIqmH/xFUmOyPP2E0jVq6e4cwNygMw
Mp9HyB3W3RZJsV9MrKxSLIz7Mrbe3NrTtXjWiv97XIIF18gCINOnA7Y42JjiQKtryVcSwJ+UmuRB
Ef/f3CLrCL5ydOs/yXUfdpBLPcQiMN9r7dmmQN+vQM2tjPDGm8mXLdRKlqqWQz+wv0O16+coC3IR
8gXPLQTPCkYsgtU5A5K52Ewx/Jx3dmanGhzm34NXAUFzclcpYqWQR8ZHBCzJfqogBYq7ouf9jSFY
ZRT5r/I8ECx7S5FqoUBNCArdU+UOBM+7ZqHjGwZcY9hWjJtxtGLFKGztyPu/ldCTop5R4bOI6xvj
fQIdJaooR6sHzEewynf0goTF33gmjOy4wKx/VVdhnh+QDSbihgXvLdp/D6UlSLFq0NE5Uzz7fp9T
/youoMX16HOUrH7hZ50ceh7mILzpaKhtHoAigVIZ4B+fYd8E+AfQcOqDqyk6Vx3zzY9Zl8bDT/ul
UwN+v2tR1kpyh8UttWYwFb9b1A/GYtBCt6Knc1N22JeooWchaOiIR93J/9plVNVk3hn1Gm+sF4mH
J6bJJI1+yde5dVru24JSA8EUThc4GUOznCiex8097b8nS2E+c4+hP/5yQlk1PWlNU8kDAtuHj9vx
Tc0vAOoeXWv0Vf6VQG3Lr3kby9nxq8PFMOWISSLHjhSSmlOhK38y3+tYrAOigPTDh6U0yAfFingN
qqhANRA1/NIbumQob0ipl50dAvXDjtBLgE6PRtBLm6fBGztzXoKfjh1J+gfABz20GEyXnagiA8b3
jfGHT1huRn9mTsgZdrIOlI2qFCN/e3XmjKhx6pTqF3nDK4WEMxr9AHMXxD84V75EFUNgXSnmPrjI
xUQglD5Bxn1NddzI8OG3cKREUD+afbvrxAY0tQqi7RC3o7sk8ncy5Y9G2nY/E4aop0g6YInZHJwg
7+Dkkz72fVK1ONHB/bq/q3oOiM96CKi99is7Szsqhgvb3oyxzA0MZgdcR/tlJ3P/Rahfk/y/XZ2P
QD25jkJx5E/ugfAlTQ6erYyrZDTW7HDY6kjLFDZvqal3sDiyss2O6dIPDLz8mcviRBAqmgjAzbwv
6sZjkwH47PMoy/RJOLmHZB0C6JXpzTxnOvfzWkPy0+9dcnnkwk/eG/UQQih0MGpJatiUdiuZHXYi
yA9YeHCQ9/wzTWusy7zMSnEK30BkE1t8sjirP3NZvX4yxWFFR3nYPVEn3CX+NT50mueLO8ojdrcL
kSQAgOshI1YnSJoNGPBQ8B2di9KXGyfwuJSNxIvf2M6NDkNXQQfpVlHz1bY/YIN5XChutzgqFJgz
erhFw3pSs0X/Y8SpK7RxDqsVT5byqthqTVZSikOt8rD4hVvD8Rrr8uxtfq+1UAAOkf0QSAvJwqpS
Nl4hwXtaDAPlWwYg6axoHIdHlbcSvtTJn4xycWF6biSowoIwxrkXY/qwf8rIsww7TS6Is6NTwdTv
SLZ3LTmLJoAmcENY8gEshu/GMvpUh7T1ffEhzLJctvFQ6wmBQ1clAc76HKU4U7gSo1zvxSSlm8ra
HBNR/tFJDctQQXJAe2V6LnZvtlupXzUQajok6OOmnbT5m5B415Meq9wX5aRf/5SbRaODDUj/CF92
uZ4i6mHOGxEybFIHp849jOhP2ZAAMkyS0TCff8SFuia5viIWYRMbichidMEID/BT5rzpyH/0KeZf
sD8lRPEESszm0/uMG6/sYtCnAekS2fqkBfFuvIxGJlAmq0Q9AV59EmLhgDTKudrEp5H4n5fXfB5x
uO2cqegsfsf+s1d30GLZ+uNP1U/NDCWOGRG7/jp9e34QMAmMAj2yGYX3lYqBU5H0ypy2cTRSAYBQ
q9MR7x4XC2LmYwob8I0k6K3coIAIzO4P5s2PyJn2DnnHc7vpQK7o/x38T6NOpbWFfrP+M4IViKnJ
OccMDM3sqDrArWyel/bmYOcLHDW21s/H5Jpd/ldU0pwz7E286ak4xXIF8+GricqFwvjWWJkXKhTx
378bJxWLITVe+oXjtu+9rD4X2Yy61m4cI6YbpB5s7gFDW3yB0S78dkJNr4svMqpZUlW7wJN/HWy+
fY+UBttQ+wnlJW/5sxM4gTQ03kBM4QZ1eyV9W+AYXm+9CmoJ/tUQILdVXa0W9g/qHTjTaCi7L46e
1x45nkjxWag8IKEKK9JmbrzF4B5rA/o8F7/abVDM/3412tRC/nDhmKQdOe6uSVrAUBIGm5fi8rv8
/ZU9KKJKZCpiYUa/zvFCyfQJUZRiqm3qXHaeruElTnjz+Qdr8SqgptePv9dkeSLFdcFbvTuUDD+8
PoTby81tTKLKeLoFuta1mFbDkxYej9iq7mIdJjUtmmH6cuCpTUSZky481Ayrcb/i3k7JyQKGN23I
P0wnM/QjyElhpBxhoT7oaqPBBQWDGPO2ZSCW7Ya1wzK6aT4PkT/TIkItyhjymth9uArXpdT/M6wy
862wcGa7edmES8iIohFK6S6PiVNs+829AziGOtAgW8TOAVsdrvlEEUouFVwtLwUsVE5iu3tDTtQm
yb9nwwdKGrUKRpqsMi7nR/VR5UQpH/FcvyWoJ/Slj8dkPA5f/x93gnDSAg9h1uV8GgcHx6HVfNpm
jl8IKyq7Faye7IPmTPvh3D0EzOXJon2WY2dDRW45pG7/bJxkZFTGCi0u+FEoe1rQdx3MzWMhzKAo
Y9kbzz2sVtAHLMMJJR7KRLwJz3dJf3+zflAj8+Flqd/r5xk6gPcW6XEm9QueEsGjRmMhRB2dwD0X
Zy9xntNEK5ch1j6qbQRe3YPI4O7IXp11/HDgI0T0N2CflxfAKCL69/xdPmzPMkYle1V6rolWjDoz
2vBGyZlw87rnrQpy3R1oqfbni/gz0KzNTlpf5UAiU2MBqd6kdu0V7AjwuiwJ/oAEvnQEFvKXlKjq
vHsYyN96K9kYyYMRruOPQF+PfaZE8PjLo3nRDM13x6sJ/4DQmFSEPh2kDEWzaTbYA9b3uJEmkKqk
eELwiVXkFzx3TIWuy7uSWAR2NEshM1b+hORdn3aCO0tVB5k15sF71Y2LIhhWQvfpvmYnZv2UxN5B
O08m7h9H8mNKbHn84mPuN2rn0kdaPHtr27Jm/FeOzm/6ZxpKnXoP/xN1KYE6Ui/69jVD0wOlYQjn
xKV2fB3qO8/1G5hUUseshcgHmXNAe1riZEKNTFwwgZv2xIhavbdem1N3pB8qQnJktsJDr1ilAH38
upR202rjlL9zvI3YC/wgC3Ef6Vm+Qxcg2hSNHMCodS17oIGxAgFy9fsRcH96LbDlbDF1asniMcoR
mrI1ukhaXmzGjVeyP7ioepWqar770U+F3eDc/MamMQYXTZyXHpArzKEkPyGL9E0zmcjB0qxlLyZQ
PLg77ESeBGD1sr7rCQ4yC9Ac5RupoAIcy/+toOODCSK6v110VEqETr6CiewXCRmimPJfYYfyCJlR
XFRLTPf2ryOLYhDu2ozaVSA4pwD/eEi7K7Nc0HZOsyigxh/Sgh0ylCRnYqNwX/vUoQLkc4NTlYaK
hs7D90w31w5Omqb81LsN01u9IdJvusADm+z1HY2AaZa310IdDPg1yebGb3JVM5z/jbMqmuX+lFYq
oGTlQofHjNa7JEC3kxdY6zl82omyPDjrwtDYBQ6X68IwJ8wAUGsiNAz30+xjRBCa8UXyB/X2Ld/P
+tR1P7xiOENpzfLcB7UHwBwPhIuMQtdFluv9VziwUy9JDya2vdVhanU3wi5FCkVas0OUjt7BTIrL
wifdn29D+3qNlQ5VNhJDDthaiEE9kE4euNZECw0trWI+cNLywklhzG0Pm4o3ljZg0BSvTAzoEct1
II4fToHrsJdKRKW/2rQZjphqdNUaBU3JkwTWcFugB7mnV+omie+w9+JIMxfRY15yvO7eCgDoc+y9
eb2wTmVjc2uST4H9irs3rhOe455Vcd6Who2kEj9jG6afCvKJIOztnaie86JJlEtmBIf+WNn4zWDc
GPD6kNnjXgklJIPC+KXjWSnSCU2n660+5Exszzn1WLEz0iA9xaFK14iHa/GX1Wyf5K8ZWKlcKDoT
H8U0nGezb6AnuVZTgceyMmNOVQkQHBSq/yV66nfomDAcYu8V3Umj2uxP+em03A0mW9eCE3lMElpy
9ElvvOKWQWyHY68xlnfNCUS3z5afJsOvmWEu5tuFO/a8lDOWKBd5DMvWAbFiI7xr8vDGvzDn/Mxz
LRfTm7Nz2Gj2kI+gp7iwb3OBbnGV26+G1XYLxZvwateagKSiKEqep1lCW7rzPTDKszNjwWUZgAlg
rV++Wdm+tYsgHh0eATn1UmAo0S8qPqg3VBldUHLMnSQQ/aDyirFLP1LJQ8f5wjuUqwF9x5D6rdmW
3vXjx9smkozhxvH+oA4IWDBbNvo6CxjN+74QTU2eRHuLK4/AmXqSOYVV3LM7Al4YKySlm8nSoKcm
b7bCrARb+/zI6M5ZfI3KTbCIBT6vQ4cfkS09ayG6U2BzEiK3G4FXzj0TzekQzFZHgUkybXvWjj/f
UDRtRJGjt1fO7058YI7fskKmSbWTMnvtAvEKRKO26fvDMYpRjwb/dddqmXwCQxQBOd0shQbIQ/7U
RV1r/6ZFR0SqGAuhtBgTTn1phOSZL3dp1iskeNmlJCfZDs/abgbl6/OidLHly0GEfgbwQh57ZbIf
tX/OymQhric8Hco9EQYynyhC/1PUAWeCsaNLO/KPGzDGB0z1g+tDMhAb0WxyZWWO7vgsJdgwbHl4
nRRKmaXWXbj7v1rklLgHAxuDSZOMBGlDQsaIu7OlDDuiI5q+NCjCXUcIgNcVagHP8RLdZi7YSXh7
PwulMVFaw3/ELW3I3DDrTZWjj/oSBnpj8ioPeLiI8qYUezv22JrmuRJ0SD6SmbjW2fpSyr/XKRgX
dvb7Xu7t1gDuJK4ZNmjD7vENNELC+8Gc3ZjAXrjUGkaJiTlRy8SHLAQT0ASBmlqZ8Ot/O3O882lN
Wv+as5BR/QCNyOOCfBNIS+kJTvtaz3YpdF/IDO0tA9Tiu6N9pAKd0TmmLBAc2ArD17UaKmonEddN
4gAFbS7fNIC44+J1qOAYYXXkjxq5hUQDIdQAddNH6LtjxKsQl3DShqYQf1xP4fBT+89HLHvCrsNQ
N10A06oFZ6u1LPd8gCAGY7enDhpDZE8KjzMxwEdKFTu3Mj+t1TrdXVmkFw1aOGpP4xpB2H7YcFuI
5s2u0dLWZTA9Zt8RxRFcTOOWAOql3yCiqcDeNZ653zfFReTlTyy9EI3UZUNfipBzbunWF7geBXCK
NOFel8YG0LbnnAFyCR9oS2BMY+QyOGfDxf+VJ8mWVavmuNsuv7VH+/+krYRCKqEC7nm5eUQQbZdw
6AwwGVYc+LTkTUehhnu++KUIwIDUAeOHDoQfVnxysMLLYOlEDCnVnBE1N1Enh+PwXIgfa+wsbC/l
sGT94u8AtVgAuMzidB3bffJmy8NTim/i5uS0Iw8u1hIXL7H89S29H5cAgn2Hp7xqJcnrMQEZo/Sb
374BkYwS+wOLycwkMZbB6n1u36SZRZAmSFT6l4PG9aUDxZt6/q9rJZza5eJMmDqxWNzmC6qg2LXE
SmKB8W1ZvsAObBxdoFvkGMJNg8wPDNK/RjCFiUabDq+M63MPkHTD9k2KTVexJ1fs34Og1iIapWY+
AhjthGW6CsZ+FKWfy8isrIP9Nau+IbF0tYPbpPhpAK6FJm7ovulpFZGx5VeXl2kXrDUFCuNIKnHt
G+E165B2xowTE93snRc1p4g2NuVcJ04AxCI7Gq3xjOwZvHGQgNo5p9HvPNiboJgFdRIHimFZoJAc
f28xIE8m4TeJG6GVtqi18CjvbOmf4fX5NGOJnMi9pLc/h1S6PJurzYgNmVRPBZq6UqCjL6ntSwBo
+F/sgK85uCwyPu3jBk0UhOGoMljHDqA9zAoDhJoxT4D4I61lagevOel8E0kovCsCY3pU7LkTu6FD
YCnO4Omgz0MJx3xKUJUTbAYNQG3W3M6cBD4AJLoCs71BVarJp4BlBx2o4YlAlx+KozyaJdt651cG
LVxaVcjoKOlVtqtd8Gbl16+EWbhljy9+hd0nQ0ZpYutSSqMkXR3XihhHgEnt+IfGvpxU3rfK2oAA
q3Pb8P7XGFH3UtsFPo0LLcZ4IOG7k5SaeICcSjxfnlm8E9mMJQMI2XzP/XZZn7eCt0dV1DjBIXpF
t/Op5nZOX0qwkkWp9NfLqBkkWY2yILL8fNwyPTlqv8+7NCW6nY7+g1GV1WWYmS6qm2sQ8IYPCHzs
U7SMpcRHvSRnrDmBpdp5Tr4AUBHdIKyVC7CIq6QR1EMIlWtDO7w0MTrF0YxaQryVaj0dxf8BGpx3
6U8fDToqtEepD8t/9u1Lsf6u6GISuC7SIoDFENUVAAD4F/pMH+x5/4ejA99ZL0HOIAZNrjomPKjG
R/HGqllZ6ablFUJZlLH/IBlte/jeFHEkxlZIyq34tsbL2+ODrP3aVf14s46XT45bY29EP+b/hgcV
TJTIuTVC5NjJbxZcteFZqgqcFt8+2yuPcFx7nujQdRUtQOafjGbW9xFLLlWZL0OoqfBIs3mdiyMd
tQ9fTxBtTXvBLEiKMohmmd7RYBcxy00hw+A0y6L/zGUPltIHqbo4bBpAfjvKMD6AuPMaTCLG5xMZ
dp3uEzUEtNuCoaaOW8Od+ymSDmW9paoJLIsdtIPK0jx4goQiGdWxb/KWARAHD3ZWAR8hNvfHuhDy
FDeJwO8t8D/riv83ksa5vyuJi2zlOr1ikJ1MgSR8d4a1AQQ9yPxJuLO6soVM0H1fznKdGyAM+67L
Hw1HiL0357cJgLgpu9ysrudjW3UFBqAmCyLKv1oKotFiv8eblK8tJrA5GZVCrsr7v8nO5ZLJS1g3
FaWJoqyp/S2ufKTgv0sZcHkM82tRu2FpyMmPjabcPr1Wo2iatOALICR8gRQVFpvv9LsZzqMsLZIC
7pwXW57zvJTNukggSEx6suTR+TlEvVxVaUHGLsXImwHu7OJ47NfDtigndKi8w1S8fvNKkKfBKiFh
jKKa6hPLlDvu+kQL7VPM9Cw/Scy0cTqU5bi8TIWhM3zxE0R0U7lroVqbR9brs8hvJrRNkKGxoZRp
sUNodnznG+CwmYf4rLgcEBF81Rmnra79qUsrkhq/x7DzIYrDXBJhmKE5gWifSvDxT9mBw8gWRVgi
Ibricq48NNPfXLuGZzcKhS+YCbY6LAAaENyvW3AP7JWNOfHlRIqKyZYWt0sYI4t7+9nDOxqboiuy
G9kBGhCd0bJIw48+/OuKak1Gr5XngTZUBkUPcD4ozFfXCSsxawuA2SpylA6TW9B34tdJgv0rpxSV
TPFLzEpQ0xAH9RWJdNlIaybyQ+7zqTi+1dM/jVKZbsbe5Ae54dx5YAPy3IG3b4KuW4HgIOTqefOP
3aAeD6yz+Gfzq27RjlwKQqYP/qYpY1ronB6a99tQ8xrESviiXprgegHGBCdmawgdwGO6+OsowFPI
r1nwIjXt17yUyx20vxQmmFmZYNqCwI5gdpPgRtNcJL3vPkz2LjRADjZrBAUrIkP7QneVXd5fXaNH
4+fUCzQeQIfzKp0FaUfKJeGeWJZ7vMBiH4wdnmK+ELWYurHFZ5lkDKcuQl0cm+I9Nm3UoPCVTgXL
xRy6xGVYKIpD8Nlde8t9dXjn+NVKs0/9WJEK0P+OJjraCGDGqDRFj5Ezs/i2sG66ZBQLIZYTYqeE
vJ/EDJ6ekAPpQiLXGMKgHUaP934dT1rGF2TU5ldPDALjnd2xXPKZBF8+W8U+phgAskcHl6sW2taW
G9yZMDZVKNMNBoUF9dFTazFMeGBtLmjah3a2zQkSQ/Wh/qJgTOwuMZnU62VTCH9qujJdJKYOjKdn
L6GxqyBDBBMyLdpw4o+kFn3w0PpNiiFSmKHL8KjBwiyZ0ZLu97DgQX5TT0kQH0baOZw8JnEXYzuX
2/tYf70eoBG9hEwfk/O6tMGV4UR7ZiJIHVX1SZnRXOm5pOb5d+ePZmuxsTXIWeaN2F4BwYPBpLkT
n4C84qHPgHUdftDv1uAF9VtwXTBsSsnW21imqDggvy9WWt+PfRH25JFJM0XDA3pyPAUAJpFPpYXf
C30gmxVP8UMZ9TTMnCVwoQTePB9RaV2A4vFS0YdidvayKiwd+BgE9xY76AMGSBS9XXlYPOgjo+/5
t+RerzcJyBkL14eu0EVBm2qeD1Z0t9eR6plan8zjFiUe+gGLDSW667nUP/jwM+sWVYY6mscmOBqJ
vlq5LeobTqX23t87Z8FyPxYelWwo7+ZFuAyJRfzp6b3HfwDCkTzL1szXgdFZ8WwXyuZFi0FibVao
YaPFugBy0cChxV6+ZG4MN5gOFLYCpQADd9s9bxroPIelfsG/diZFj/9HiNSGm7kgB7QP6uK1DO28
z2/U3KHzAXbFLU/MG/tAfKJuLIh1DURD//42uSfMbghX23LLfQODRQOpzqGmIjoB6jtLhLYafmPD
NDrBqkkk+ph11OR8IldgH15FPnWRPAOCKbhweGKSEc0aQwQf4bbbMXqApDq6TKcyQv7k3TaQPZYk
vEWZguE1/AWOTq16yXYWeUsJIfe1ODjSQhX89rHx+ggX6GoQuWzJftvVp8efuQP7dXFmali2/QLy
eo06K62VC65EcFS8YgPRBnJ9VKOfRQxpf518yvQRSFPOgi56Rb6xicfcANTgLz8et2cnO7ywlbJ/
CA7cnnvM5wSJ71rK2Tlwl+qsmpBxERZyGpDufxv/UuLE2XRK3R+aJhoWFnJLyS1rMHTictGp3Q4q
wFR3TlNDpDbc6a3L56JY8mkBt5qyvNSTpBac6ZNCHi+HADuySn+KsUVaqyfX+749hY6eDQTUOY0z
75LFWwkC6HBcvBj3frOEhnqgEt7R4Q+qGxGxJdgp3Oz5X+qfxOUwEaLEtRE2JfkIbFVsKDFPfoIL
6y5b9Ci2bgzjFwdeZlFBjNe+l7ptdLogCGsw0eSz+uMSSvXZ7DQ6m1gR9uUHdOhjKZdqXCdGJA/6
21Wpr98Nd0lOXUuZiSj4t7Iege89HB5V8NNeVmZH60qZcbI/dLgAi278uflmdMBGiTtxt1zQN4YI
Wz1H5K6dnhpS+NAU93lfuVoTZjZuyZOWezzzXH9c4kK+yCYKR6e353B5+CbKez41lxpI4vfW5Juh
qxA9TRDQeqLWbieKGXLuxPpvOh31uMVj323zJRAZufEiar9r2XGN/DXpfSfM8W3y2Kt4UBVCWstf
FrJ7RpZDW6H6jomSkhEWxGYousTM4zUS+YuK/kzXrK27KAh4lp25cpllefeixB93qKrRKtcQzmuK
NahS6uhU8/RMjbvcPgj42WRoNDynSyrgvmihJXIOMBbXoKXmkNyfYmHaZarRatHjvanWBMKv+gml
T7dD8fTj4nWmedFQKLbkzD6n1Vcv7NXCcc9HI5jKU2mppJVjHvy0oFYmwdPr4Bun4M1B9XfCtzWq
kEDucZ9nVjM9Mh+CLgCXCuiLFpkyoIH7Dm2YtyzoYBVa3ldUAoljPcxqLe6q1UnIGTT9Xsowp/fs
pm2pkuiInkyDaEqXsj+XK2VrYiEuZcXOmE1Lx3rXdhzvqRdBDk1HWkFtPtxFuxp+J0BVurYYUjX4
AUP8U5B/uZyJcNNbY7FLAolsd8WDdROgz+32V2XdZb1AJwmc201sjc3P9gNYpjn41WDNOgCQuQzu
sPtAuWhCl00Extw35jDcnKQQpMj+WQqbZledikAjmSvwKzoegEeXQ9T8HrIh7qLGEeRzQp6CD+ST
EGKtIBHZbD2jip24yUZG7ICJSCRw/bHxOG19GUXTDkftCpvKpGV39bBmX12d2EV550N5MP17Soma
OGx93cttoCRP2GX7OAMOmxQl3+z9Z8JefeNnioo2v8rg37NDC6yXyRR4H59qp+kAFiSSg/+s0K3m
UtarWAM9xpJ3grqaSIOCcw9hADgdSYQvG3usdljW8CpK+iu6CJShD2HJ9XAXkFBqwhUIbpWR5gN/
tlr/TGSsKemFSdz1JkyDqmL/9InhUPine50Fcwsn2mQgpXPfzeK5Q/NHJeDPZkhvrMmSQOyIB9UL
wgnWwEUFGPgcpp2UOV1SV/GYRivcGdhrfRyDhORyaKzT+uukOvcFq7n0uW83gX0Pqy0Ib8CouhCB
sWZJm3YpQgyGqPdiP0PDGMc5KOqed8X44e1Eph4Fp3BjbHocfZPZ2M9JiiEDQTh3Ij6pVz/5foDf
H93bDSnRbuEBbsfXYnmQup/9p6KebFY4+VvcQS2zdqPMFT/+1qHMuVG3coyaZHxJkDA3K34VqgVr
mqAAIIOcOyPabRcqYpH01XW4x/IdpvEpRU2eUDenojCSduu7N0Dw2/TRjAaOeGc5+kZ9RjxAdC4K
MXm5kE/nk6iuPi/dG3lB8S/HxKHyuTrORjX0wOtE/OylRAY2CYriFSRO1JM8eyVftyoQ+Dof58kN
V7edltO6XbD+ewNUe28yU4TYMKB7VmEq+xCTRzPFe8EOmKENPEL/R3YEgGW1T2UaYdZCobxA7eQl
HAo4vnLdZTPm9rLIH4C0b/aenKvhWM4c+9TrRFFBXNOaU+/44RmWrq606hWcUP4dX9y4ERXioyGr
Qj8VExTI3KcsJf7ZZFoe4BIb4gI4mX5vkczGicgsmF5abOhr0G5MLP9V1utrvrjmYZRgtZPczYHE
WHVIhluWPpSJb4wRnzS1b9GcTsbcD3TX6+mMCB0VRw2E54aQ2GZKEw39cVTD5FHWWZ66GPvfjrhW
6msSxS4pWZA0N3vUuNw9TLWokzcUkXZ26rFx/3Yk23Ip46cKTwHgpivhgKa1VmocnpRy3NvnjPiP
ygtKgy08GlYo5rSvAhP3FxaUzGq2fAemCWMiFo2gcnzvpJT3ag1xP+G3+0jlpvXnNOfVgcRJx2OL
nNvOXYrv4GrzlrX07nKDuz4U9aE4wQI3J5FN674LtLMvGWgagvCoKkAN6wlX89MU66mZOFJYpzo1
k0NmaeNRN32coMWamlpXRsbS6Q9+8AHwiduv39oaBrgKBsK1CtfNZ9fznQhruVtyGQumdTn2Ya6p
2JkuyY+QQqctf+EIV1NiRJXcnsuqCZq5GIiaGC97wDJyH9EmRQM0PTgipPv7zCrNXTZVXnHv/VJu
pV/ke3bE+WUT8W0sip3n6Nm+hYzmGtF/cZJ05YYTWWf8t2qRyDV8WZa2wF877T10z4nNBL5l/9UQ
vm6XEFxqN/WOnG7ZQD86vSn2EfzHoV8sQVcQ5T860TbPp+FcU1jenPugpAW/MysfM90ZT3Sqt1ne
YUeSVnUhXb7xIbJ0B75YU1s4Ze/o5mTJhQSkmj36GcxasLZEghxgpbLbltbCOEn89Pgfu9czvlft
iMDMDWmt0714kO1aqDPsOEJiDLAEtb7YiT1k7/cfHcoZANjtyYA/+XK4WRYSkIG6hQ0vjisayBnX
E6gWQwc/QFjgDAtJkjeNriBp0pJCaq+tHalXwoXMRYX7mdkis3X6FlMcL4C5i4xHS578L/CGMU3q
6+fDNuwWq5D7o54V6yTF89vOdysh5x+w1CbRlspGqATp6JYxz3VMTH1PMlsugx5KnM6ixDPqV36j
tnhmfGVwwfprINQAaqjPqY6B++1Fwym0Q44pE56eaY3XHAY5QimDD171A0ziryqoVWd7PdQARikS
b+P0qLsEKPSZ1n14u8OSk4DLm4ojKtaNgtHMPfv02fZ/hbaSMn4k8fhrn3BxSeQZo9V435WMr2Yq
q2bwr88AaiI38V2PIkTQ1SMRSQn6VyB3tDqFEfKklGRj0bS9K/dtquMplqWYO7RqzpEBzo6Ls3Ea
6AiVPOZdlsyPE3NLShE7HOj/8US/6mRRQzbfP2C1h9kNfOIGCohTHjFPaIMMZOF7txVc8zvWhAz6
En94LQ9SaOwU++Ixx4QnZ18/v5dl49bPHRLW1kRyAR05SaiT+AEpGZcmiKlzw7VWoB4icWlbvSyM
Y8Pj4fv+vj1Q8z4+gaTwT7YUTDrNlO/WV7jyyE1X06RV2lU0xrJP0P2TtLrLp0SvH8hY9kVU94ju
Gc200Jefva9xfLjJXOb61/IBM6l2N6OWctyb7BooxcYk3EUoLBjjohmtoYcqnMkTk7bXTeBjJl/e
18WDjYqisQRfOiQkljEmVAB/r84pimqvilwGOhj5nNp0Xh7h36pEPns0vDgRxcC1MR59fBJRZO5C
5UG2qzMLfEYtK2f1YDGcU4B13jbVLKqF0yteVK/vlINwHLUXuO7Bj0IGEhxGS3ibFnK274JythQ+
C0glrV4+Qf7NvpnzEZMfayCh4qLCKpHl3yw2V7SOKoOQtbxvB2Nr0r4GfcV6215Q/HLJJR+Z5c0m
Ub4EgurEqP49pHVDlYMjo2JvfWHcdFBCrFnFivQMCTGyNi2bW7/nP9Hh80/v4AMoZ3gC44xCNN+H
SwqFiQWGrKq26JocA3axwKRUieFyg3BMIBBry7gRqUfyz/Pd936bgVmnufmsrfm6Bw0IGh0J5N0s
aFvxm4t+8/5Hexgt+2R221gGhGaiuLlE0yX7zUMrQ74BBMU+Lqpyc/Z0nMeJojaJZh4JNuENU9FU
flGp8QKlWIrs7GvyFpm5bcR9b/aR+BmnEs8aIWABetwIDOuH8hnkMZJJTWgchyxmR9KhNhIthWE/
aM7BiH6KISRDohqXJ6Nk3ueQsCgaErp8hbbBPSA09bfWqXV7I1jxw+0b97eOhMoLEzSF/kCfO4k/
dkevpqKUTjCtytjPJhK32REkxy3tKJHZh9c2ObZeJXMQeJlKcr32qm/bVBDs7I+fIl4PBnGT5G3g
DW2mTj8KWQLFF0Z1Pzucupnw0P+vSi72MyHnTljq1I9K6gOStbjU4hbPRVBEbtwFbC2+kpAvJchV
geQo0mqUKHdGjB82jKLOjbW2sx7B+TO3Po5EsBam93E3929yWqcwizlA98eAu472mPWWJulkZLi6
MiMWaky3oFtXgF7C6tC2rHOWGrWQlUDkM33/Jzdhzw1zM/slrFKxr4usbYYcQU5SD68r1mtHMFfZ
HSr+u+hhQLGflX1rPmKwW5yWAJTZ+z+UWMwRg9DWyGtHhHq0Jw7bhnVQ98WQNAedfPQM3nkk7Xw/
kLFP/trBj8uxLCJPJcXCg5kuK8vwqRoV03UKHF7e1GLFCtuOLqyQ7KJWRpbspbiVQtLNkZfwDNmL
Xfg9IyrzPFoGH0fniwsSR5b+OrRSHbDMYbXgcAtbsXWBmq1tlqpUJ4Xj1WSBKvLCIWR9PTsHz0VV
90TMK73yCfjyOB2zxLaxkFxX+ScK7YfXaaK8Xm64zVm7xW2vnyqUJiDTqX8Czz8eLDdoELzQt4rl
xAIKUKRv0R76YNJJHfussGQ181ChtZRPanIIBmv/rozqunmaAmiSobCz3D6q2erGhoYHp/uB8d3b
SkwgyRpdcsXVM2GnC5DZQj2UJft+9ql1suY7edpwXRnytDP5apyUEN9ElLPJ3o8Vn+PgH1LDwDxy
nIwU7ZXi0pOXBYbUWy24PXaVXFSuxMvAmp8fZj9MlL28nNnNGbRhGokdbhfEAQE52Mc1ycZ98f7Q
CY1z6V7AWGBNHGaXngpqWYXOeboGy0fVEHVjyS2zSBASA9LFP/RSnB1ARrk1TC8+4BncMj8mDGoB
RaPV0jbV9bccrT9rkeUKtqr93yE/piQV88Gd1uInW6o3uhz7ZY9JsGmwCTg3kjZ9hEKHnmppoWs7
flKo9qcHIP14ssxjxDSbITlYZql5Ir/TPxc12CJus2D4s9yQKfhSmGWLs7stLZJksbQdaerNv8nQ
fcXoJ/Bxr4pJbk0hOGGsA1h+8AIvOb+orvANfWF2aSWLWiNUtaxhgL2mb/dgzB6VOvfKx55gbJlk
u3iUN0SI6xG69SOVGyAyi00366cCyGWcGi0WBQD20LmV8euRbN9NjQa6JI0dj/rzKhgfhZJE/6kc
rrfUI4H+suiNlvqK3mLgPOKPYBg0psA7N+qCmgSmf4zbUib9tu9NeOYCwMYBArnC3Htkghflxd8x
dmhDMjwV/cLlG8Pj9hINBrDtx7t8S0H14HDNxxu/Btp3flqh/enr04GkXFXM4YS3B/by6E7mVW+C
y38c8F6UlDNlBW6fz71SzESp35Ttuy5slluConq4zpJVw3aZoEIEBGYZXyaumVunWXh9AZ+wnR+j
gVdJSBIzk6KoODNZhZT5w+CK/jFqjaeuPo/IEOj+o0vAbB+NwUDrf44V4RjcA0A7BFh28CEB9QkF
rLfBsJrL5JLqXaXTnANZzPxJCvQhFjqCqcMuMmAkWYbgeLmvihiK6OXnNXepMcoG0PUFkjPJ7b+T
CQ9WMjMow0SVf3atezrx6GXCL38ytxeGb3v+JUkyGcRlIh7YAjgu4vt2qXdekUs2FjyohP3WJYTq
TrV4+gcgculwBI2LqAhbx5g0VlB7okyqf3XwFW/g1G3+dbnBvVNOpTusbb1YU0+1T4aUfuhIB2vE
wmq2I3rFp159BFhYkvCdyycumuE+d42ypxfgdw9JQ5Z0np1hMukB7nxPUBzMWezY5D19c1cF/fzO
2SSh2NTNo1TdEcvcpUAj0cc04HeXnJF25eUqt482ANI9TLY5aiFrJbziE4LWv43iQiyTxkX9KkWf
qYLbEfrXgZwOr3/Pa7xKgt0eV1BRuPhWDCyiUJSmXoZq65hXkO5weqgmLNmUAPWLCUNFdSlxtLhP
5WTXPuf5/RQM/KO5PlpAUPGN2/AOsOX+YTBYTUSnQ5p70rzU9LnLHUzo+ualRcg8FEB1GCOcqx17
QtjAoVw8XcuJmHmAOdzxEJXGs5gG9/o3l7eSq5uDQ0MnwLL4rhAVHz4y3ebXps9aeGtaMwxO/O5C
+WK8rygtavIA3pe08wcwlVtH/4TgBph/a1HqaVAicMcTkg7YZkLR+ZVnsnslpK+yZxpHSx02WMTj
0z8BXWF1MRboas1wS9IabgZgvNOPwV/AeZUqLkcv9LbEBW1Nb75f4U+vj0WGpLIe/2ES52JM5C29
9cLorD66Cl2IWx47YYG0FZpat483QnOwbRDB4TEpB0j4fk1xSpawKhQM+oC2fH4/GRxmGKFcPfZL
NbhzHGEh8Vax2D985+gsVFqzlvR4O3RiBfGY0+YR05N9pBjkgOGHAed7JU3RMjf790SRrgZM03y2
IOVPX0Oruo2kIJvpbnwZbowGey9mJPuGFnP0YCWma7/2WnlZ7QK3wWLZnruoEOLAhJccbcdVoKTo
dIMXA6RgonT1a6ln8PdouMqJkkBCRqX9d9EsCpd4zZP9mUcOat5Vke4UmiFuePutZ0Xv1DSMtrzT
cU4IFYn1FmtfxbNzh0UrEWEH0NLiUVHwZerBVMptUVWljKuekvwGaxpRSeJ8Yo31oSyE8CcGeGR7
x62Jd/fFxlqUBF4H6SUO7OvVuswwoEKZTx9kkAv4BjW33zYACeYbax+EfywybCBHH+1I3olYQScf
VLJBAK7dZs8soS/HSmkRtIXN5ERnqtJpnpumOlRiZm5KqrcwFe94YkWgUY0tRSRPEQ0aq0n5AwK8
iMEDmysMrp/Y3TbMKLYGRvco/zRQrp6AWjksOtzjE8d93agReTG8NJlzkoihz/DUIUfi9bSsb0km
qhlmwcMe8mTda8ti2isxEvXnF5iejbnkcT59fnN0PKjiD9atDCALkoeGb7OY+O74zENmwm1sPffP
jsqX30FH6d5y0IN1fd3A1exaKTrfzL6Jroby6nTNdAuP3P6uMwkyqEP5LFmr5XXfUbfZ/lxxodiF
MMXII7K9lY1wB9rCV94x5FqHwUc+CJ9+PQ4lLLzTBUeloAbHiEeatI6FEwMLn0uZnhIX2YcjL/ue
nhvZ87Z8XuTsetQ3HWaSxczihfa5oI4M/bTlNV33IGUGAZdb/3yjs0SgcDb6bsNO0tANfLDiDZUh
mUXMML0gtoxTiyYMum3JrOdNBqhhd/FrnogZJxiXyKY09Ia7V+4PfDpflDbm9Y7aGp1qTZXBeRyM
pRnxEcozUl6XwucPOdSUEUIrP0lUscSePKhxHiyXaJNSzC3KECqhz98Pf5KFojcXjBQCM0P2Oa2l
kt4kelesPgXRaQEos1gecT9ZZ0mTezerXU2kDk3kSS9ZLYUK4fKVuScECE9HTkb1YE9FRAS7Vu3V
VKz7FYBwkG+WEfcrBQoXv0phW04N0eixCVJClnCt9aEaAV9puBDNEs9yKWZg6aQk3Lh1dgVJHoVi
ndLGMszrOGksi00hZlalPH63MskcCqplyB6cfXQgU3LqMZxAXzzUvzw6ZAqGstVvMhywVsL44KpB
VJ7STRr6vLM3Az2T1tWTsGVZUPfX1QNq/C0eia8fJLE9Ptwpba8JIYd+J4hpNu7yK8vmaUFz3Fpp
B5P/ARZ0+MFG7ybfv2UHjBvqKLkDeCx/HLKcW61QO2nzvIsD7vEO+ro4dWmOd+rTIEFu85ulmfBG
pVdAas6MxWoQM0c4//h7s9Q2e27+RGNEdvaPtMffmmNyJ4XqqSYSmGJei75vo9cxZ8TSYy9woN82
rPgXuTIWbiBW8slL1oeaMgd71cYLw5PFOtbnkj4v4yEC6bd+15qEDonmJVMBteYahprZjeINsVab
7T7KBflKE9jGQOyne8xhW51GHfWImU3ohwsbuNDbeQn3eX2HJoU3XrsmQBYAkWizpd2NIWTPwjJj
DThwtPdo6RUDygAJmk0AswVdbvJA51UW9YPQdGY4vRM9mViWYOhTx9c0brF2F2mKk6pXG1ohJXN+
gVu6kZORI79DEwGTzHagIqdt84JC6NRAfGbHJhen3nyRPcaL/pH7ISzacBhr81jHpo2QswBvE73s
/JHHlYuaRdnnh5FPyXgt4LcOCOFUhW17VW/gVaX8ZpXjQkhe6jMzd4AgD92nT+aVNkFR/Hqef0DM
2qQT9Vb95Gcktk6hFOAa8wyAt7RAH53BA5ThrI7kl4itlX5EkphAY6+gVZxMie7GfDDV3PIVJdow
m85MRQ8bcnTMBwHmyacERtvvwL/QX2vRiXRyqJ/kSZXgyJp4zE+/fkh6OHaqmVc2qeUG1MIuJOE0
M+xMT7v94pJsHihzk6h0SNk1sGbyoIcBZl6FCngBIiM4PB/meHwZXvAVYSYSXRlaExYDkyIdFhdl
l2YXcfs0vGOOBS4+4aW8+sKVIGrEPoKs893c51EYpLzcCJM++rQmdNarPGr5xbpvz1o1S0MzgpCf
WywIo+/OPq3p4o9DIa38Nj7ObZU2JupJQ6l4VHw+z9AfMjKdpwZcbRJ6XTQhv3WoQXQl+XGZdNm+
WX2YQdshQNJUdBQtgwoyE/1A5r/uDQdxeiXkCzbttEA7YGy9CgHPhyJDYIWxPpM5Pefnl3A5pZz5
5gCkUrGfODA+wlNO2U1mHtW0FDqWCmU8WYpg/EZEn8/MD+/IsU7/ww9b1jl5AZPbJdHenoTCIfKv
FcGB15fKn2kvNANck4JYZiK8jvAToT/bD7iSSZfS2WnE/KIzD9XqmMfXgCfZOT8ZlGcY1o+a0Hpx
fo4gI1fuVo1Bo6UqeUbj3F62mgdBh3jQcPIGZDbeguyMUkwf3kv5uJxF7TIwFNYjGTbqBfjgj5DO
Cs79yciA3X9DXIuAANTQBC8pPZVkXSV4VdQ8zMtj3GbIMvM/yi9XMu/bIQHtSy2OjkHmVreuqtNO
tbCrCiRJU/bEQYh7VMICV4ie/jv6nv8jBWrJN/BHaS8JAW+6GDvf1SIfKpKECcXNHoikkvbQOUOf
+Da8LHww2mf1LFu1QtmctvI/0IisrRNICjNSVdHdQ61hLdhL01GLUiFrLUtyevtOWCtyHxZFyNUi
Ykxivq2Lq/WjxDG2LzFCn1LZASCi8dCAxiBkpTXFLgdkeFcSdYECvCJ28bXx/wQvC5IZp1ixHg4W
iVSftqHTe8ORvOD7GkA9gIrlpKjaVBZsNBfo5n5kIIrNKw89emw3mhaH/v3EpjRzb2phGpcLdovr
sUJjiIWZKUE58FJ7qzVfhRT5/riO9g03Z6NuQyYod7Uz1Tnp6IK9t9BZStKZz0OSU8YM2kddfqM4
NUvhLj9MkTIqS2pla0oZyxS3JC5RfOZhhxrpsAxP8XHMxQsfSra12fwGZ6x4wUhxo3qxTYwFgvf8
51JjDwrfxlzcSUc4vfY0/Fz/9vnXLiHlKRj5TgZ1JQGphO9/O9Om9njjv/kxuzEgTChDsTgbW3RR
pyrU2bLqwfKKcc6RbkKgUCJLbzgI7BEx8F8qqE4PhkT8BnGnY9U7SwmS+hRX5T1za75e3ic0KuYJ
+VBHG9OeiZA+AlRqduzAJjtELyKIC2qMJtvnVm6HGdzxZrmCTO6c7BL9dDc9+b1SJ63ncgCszuTd
A7FVqwOmZhTMxkqO2JH0tUSWV3O4p8uZlxIHTo+WkYYPGzsf4m1MqdZZUD8q0UZUXwJXI5QDr1ad
QC5dfHq+oglu/wN6euQu9exnlKNGQ3D0M6hOHGfE4bE+NmqQF/0pqBczWkta/QVF3XYtW5IsRxPH
DaKzOdBlFBLpxs0Wfp6EMlWrQKICNiCbD4BFRf9y89H6gWoydXvqcQVCN8sex9FwvS8fGvWS8UeM
/pJ1GUAO0tP63qfsWViOs4H64m9BbojNclR5i1HtqgeL/ZHjMa6zfOmBEN+Fpl6tQ9fks1i6hxNO
l+jq6+zRBvc2PQ44pHybMCe4WYaP495MgCTsh1BYat7bk8bNLtsaKKHz2e1D2YdZU0UXh4Uew9F/
WUtg8si1reMx05rVyecxQkn9NBgkq2yuWNiRIU8Ft4SC0wxDCs5khTQ7DoVHc0U9PgGuolC3yDvW
V4nja2ryHwPgqbAAd6JXfgRLa3RJ4DzieZpTrZxbqwElBBdX/HvUtKgngwX+y0ecJ0BB+FCcjwb2
9lLNpLp3NJVZMCeOjGMP3ETR5ynfWILILlf8WaMnlfBJ8PXiHttQ+jv1dcUze9ZyAZVuOhB1dzk7
EF0Tw1wZRnuv6IcbUC7hEnUBGihYHxtZUiFj5oToIbQQjbkytM8NyPKo4YPOxSJG/zJvlw4L7siE
Bc8CnXnq+RlTh46bqOwbks6qw4zMZKm7E5wQ5PCA156ErQxCTtHCf3Lj6M4j1bt48SfGwfbc8KJc
hV/07STcNlDXmDf7h1k7scmLpC7yfJ32sjjS58Zh+PfdZ3/vtWiyoxD5gjiQ2Ba/jGmHfB9NecO7
IYxgdVPstCSn2NPhuS0dIFlEoTFBJyPIEdwsiv2zEiMGuoRorSS05xcMyzEQ5yKfbzMtoD3UTVlW
yB84SGgDnbX6+9GYHSUjW1BMK5YEUnsdpWi1PIiA4cr1qENmgifeyleCQcwk17Ryk/ADnIHVWzob
jgN4bUGupdszkae17VSyT2Kn0bUv5nYXQgtogmInPl3Ya0O/AsgVQw+fFy8QWkhq96or/aKgjSh0
//iiqPP89Z6mMtHReoslTMbUe0LwB9YndWIF7mB88eFAD4mpaQNMP6uhINTNR+RT2zn5LBQi31L/
mmT2cqlB78uL7xw3xWRia/aPgq71jcn+vSq1BZ3Lj2QBjlc+y65WYTue+vwu2lgo2FRnuodfEkkS
MVlveGG76VkKPDR+M4I3rMlk5n/HvUZWYIpzOdHq++KElsEnNzuNu5Anzb7Dj7R9nzNNM8QfwsRI
ApyaoiiCu3nxFHBO6p0oqmu4NZaJfYIcCZjrqPLFzzGOOicCOYPMKNHjvFdkq7GSj8PD90W3yEXB
D8nrXx6SevTnFFl056jnqm/tFauZcMwjCV4YrSBcIb6KmcWsRAPH53QplHH1pRUtEhHlZHdXWuXV
ClDN9u4EKUFc81PDaDbYY7XLeAkT8VHQ83s+Wjvtge0jB62CUs/Cl/kxdE+0rvwpflhZLEG2CsX2
d89tsZNdibNYtFC5kxUlcVirGoXCnov8hz4//H0CxZtLobe2riY2DrZbbd1vWtQJVnvfJiEcO8C9
HJt5kkG37DI2gtr/ZQACqL5J+D2RsrT/7otxPtPws1cBKwfoF6f+pdqNsMea96QX++bwQvo2KPH6
sdBxOKQvr9TFmcYzidguVjK3IfV+IL75A+LTK00CuN6WRXvmBpqzei/HrZ02iqHG7NYwP8pDwh9i
TJfMJgiUI6gf/AXCZoDu5krNL6pOgME08e2rNl+yTjeye43r4AjBMKThwsV2LfCLy3ltpH7SR4IX
d+EDkadwE30AynOqstrbed82VeW4SREc8sg5ujoYe8exXYxa05kjX9G8g7WgZqJEdmMPWLkVGWmk
VuMMkRf5jdPRAm1s2V/k3BAdog+HiAPVEb7TV/JOwj+fBx3nNSsd8Wq86QrUGZuySegy4ELYT9nB
rql1ATjol6FV+MccoTHUhW2TTolIVIQ1G7qtLyKEJAj6xsSjddJFMVfawjyjnJ5I8CbgyHQG3QW3
l7tcdipDBStMyMvuvh2xGQAfFHjbSAfCo9cCucoY1ogANNVdckiajJwZdx2Ijy6tZRd4evsL3D1v
8yYWPzGVkPiFE0QHLSvK0M5vABtxhIb86GgbyDHwTrar4D/I8X2Rjjks2MNnEr6YGwDkdCs4NbSL
2fGi3uIoxTBdV1su4bJJue0AUf2g0xdPVuUxMMcz6oe6usHAsThVpIAdaSFUHkB2pjd6if4MFAQ2
R3FPBROka/hMB2UeCmO/ThTFBOClKtfdzgfQivP1RpnwU/H1fkuJfn3B3KdE86b5kplNPASwMwuj
VKn3E+g4nPc+biSUugAEmrd9RsKghh2jvQ/bmNDqdsk1hzh8a2xIc3Rnh1XwjEDwp13fIFiXl62T
KkNzJ7iCIGLvgW8q2iNDgaBjUMmfviUc0InBFzIyFO3Z9BL0PYBm6j2HENOjgTuDDvwB3UWF5ekX
fzIqJuAPiTAsqstYq6xsh5HlBGlxVduRj6OuMx7OnaxJSMq8HU3JW6tRK926ezr5E8jsCuU0z16+
2r/9f/DU+HWPiYKTrRVLPRvvyhT9aE0AkO8VOnEecwduAnWnLD4ztVWBSeZGK7nXS0Nvdw/Iv9fY
7SLG69OC++XO1RUhibwVcFezlyfVitIiGba8wfRk1UHI7hAXSNEQs4wIsHaqp1i9sKOsNp/igjho
JhtNW4dOjNLRWcYMBpwZ81oLQquhCr5n0N7iYPcPZjxs0tnJAaCxlHG6z7YJJQyLRknaBl6Yp0z7
pwhbfXjnu/vdG/iaiK2/b9AM6Xjw1viIp7IW1l0QiC4mPId0RLUjpGYkNMpTGf2IMtiRbyITYNW9
V1HDuINy8ZFveFMLw6k98AK8jmH7xBkOUyuYY/uz780iDKN5tvs3muul5vMom9bgPRW9fphP07jF
eVf28CzqoKcXlMofh1D2Pl414lxOLpxDr2HqKq3d6qbmzk8QtsisUvY8dzw1qnMn5IhjW/ExPui4
4HUoSdJa8cH2TorhV8zHsx65eCbb9+y4e/YgsjxhLGy58xZSdvlhAK8y64oEx08ozHGPRJ16jCZC
q23b3Ois783JfssZxyaOC4e/iZ0A/2V4RXTKegOHC9ETgOflMTAz2h5G5S/qo2/04nl/8sZU33G2
HYanfG7AV3VOcAgkD3hhWuFwwW+I1Hzj8LHod7SGVRE/rdGw3A93EbMIy8B2ZRIppZ0Su1wL7lws
iMq9xCcb2R/PmlBWGWNh8TX2K2aBPgmKfcYaUL540h/HGxeEoei5fQJ1jjY/f3+Ha74wSOvAKN8z
fiUgmsomgc/ZtV29Q1mKHFxHfKfvUTB3CINMCGg+I+Av+XsNWHqE13gW7QiikiOZ0WcoERjwyZzc
C75w9R3HZgnN3ud62SMVDy0/jDNRNu2kNTD2cN92U6fcGZ8Y8OHYVtbH6QbyVcy58AAchKonkHKu
vBLvDSsO0z/zAIr5UIB0qOLMt0zr6ocYDCy5poyYrlSEeQYe0EQBrlUnvsms6djVdZr25jkoOd8b
SMjR10DY+F46mxdfWzyvC8IqX9QoCRdL1XpZuBLXzn+cYbOQZYYQ+A8O5qTqD/4e6T5JbIn67ft2
3kv4rdSWQyl+w0n2VK/kv7U/gpaTCdCo57SM2aeguvNUrkM708iNVpLUWqvB54GiufzVypd7sFEV
1bdnuQOllfSA4w7Qiq3CwD8vrLfqvT15byRI6mJqajixPV829+hbiMYDvrxfzq2RisZ0LEd5BET3
nuKsqepNP4E6sHLvbMyZ+VkTQFhg2WjfI+gsWwwtxQnOO3zPInqHkAmr5gHnjCLUGsnc5jZHvLn3
FWuZkEaAc7vLovlvdgiXtLaCq0dikWWkXRfThZOKlJ9ZJUdgUOXMTePz4KCXfGtsR4gK3DKBxtzF
GCyKVN2neKq9c3TFt9LzM2U9TkUJp7phPPZ2vsiHThoe7pn1JhMsbXRC9g9mIiqAJPj6nX2ULU9W
IjdngvJ13hh3VRP8emSsroMugYKtgvItaoCGDPPLdsKRNj1nuipWqxCa7FKcsvTJzv3b2Wq/AoTw
Je0kSGIXURaHhzS7bd7vFPEKRbb87Ajqoa/GGuzmZ02ThbY0kdVSxBhqGie5BJYtji9FD174/0qP
DvsjCPmsm9ji13w7CtSvAmpXPIr6IGVtEnwDMjHJdsukD8JLossCky7eVp0PYDUW8nIKRcRls+fT
MW3Q6d7tofezxibQYoKR+Q1eiF4gtABSeusk6xfq2oblvvVZtp+yItmunllKsS/Bk++I6ViQcK4H
PWUglJtX983YzB57C536YV6qOzqxkSkutth3PZCYwoCMIH5h3BSJsGWTwRYcuLNS5ExQP30sJcz3
KhBdPXcLxM19kLJPEus8284oOq+X6Vuvn3DkzzthWPmp7kU5ysmKtzHYD2/g5umEs77p2XoBmWtj
iNeSljE+G//k+Q+c8nH/2sevjtxsKB8Un6GHYqKdwgLsWR5FrAsb7ep99hKa8YZGsj16Dn8XZbWq
jgrNYtfwfVsrIOispl0VDNhI57yYugIzrx8IbTQKPqsEbuzbbZV6yrsSf4k9dvecT0Qq9irWsdlH
I7EljN04y27A+z46bFyuulF4N/jJPX9G7koZAgym8JQJe28eJ7qAJAJRvf6NIR2IYRNVx14Jt9yq
DPVxT+87r7er3RWG1SS9//zBwV+Zlp5fjsrtZl87I4czwJisLaTyK32JQkJYBoVXcV4Of/Sm08gF
1uaQlcub/8JK81fZtj/KOWiUDKG+cURRFhv7L2GDUlALf5iKWTCSBMEjuF4LSR2Ohs3LDJ9YCNrm
ZT4DQJzeVzFdU3dYiIQf7CsIqvpWaQkuGtgPU0+vJkxINpr+1mEM+RZU7EUkguE3wajIQemlOYJH
bs615CNmSj8r4cbbNffaBUKH/pHx+V7toEmrinUXG7qI9VVuC6Cpam2rq7dqG2JsArMOTPHidUXK
WMS8LY7yIVRFs6TTm9YuGcNsjnHXfYKaMufdt2ZhHuSO8d4z99zc6MOx9NEG14CUfwNsEmeLCcF+
eGwpkYuPeqCBSltSHr8p7be1G1eoLFyfSzgfiB78HJxfwz0UfHTGh2n4zHE8rl52cBn30S00es9z
eQ4pyEWc6jZHSMPdKSUGfnDfLCaiPt7Dqclk1IPXCYVUp9/N5sdDa6y3OvuppQwAH8Gk1WQnbbC2
B4suymUsTCmPJEfNQ3nrVnWG1YbZO3yCZUrzxFIYzw3kK/MXyY1OCOlwF9q4bEycKfLaCMMZBFjO
xBGjaHgcjheTpPK3X3x6zeHYm6RB2rfm5Md85OvBxjFy7jxrnGvPbXBBQMAaUQuWvoyLLl5Nh6mx
hDOuiYQ6dZlEVE0H91UR677gwHSiE7TT7qvEGuirDZ0rRN/r7WYMXJz0hfCDlyW8H+dZPt1i+ME/
OqWjwQQLchLEsOCd7wy85TzStxmR19EDgktAi4fcHUUrnLvh2SpkwdaEIozpicfa1LzMN6V35tuS
okWwbQ6lWHBBvZbsFVzjdcL+ebSPhNTCvzPiVsHXRpz2n6hNFznZfJBfZEzi90rAAaoPiMRriakc
xfactZWmaSTgd9C6GXy0nZpjvSack2aqe8iCwx0BZJYdHNRiIE4c0O7CEgFg4jiGS56gx3d1RWk+
G+mN5dj/iUrVn/+kRRO23U0wsc+Ib9vn6BboYmtGqMQwoo23aPyoJuBy0EsKMak6FAe6QrwHDgr9
UVOFq5nDk4rvaDhaBmhgpWWLqWro3sG4vfP90gQQV+otf9EV66u4wtRmQxTKWu/60V6HZ0w++KNY
lyta916jZnMHJK22+zuY27F/w9hk0F8pdm6vj+GxzQqyRxu4FA5W86mXaZaBu/nzEfikV8Rj6HiI
hWTRG1yPlEhjK790lN7gCsPZwnowjwaQ0exIeBGQcyXDnfnPclO3ilBAXD+rbMwvwJhkQUBj7PK0
cxbEGXFLkqMBMnTGHQ3QG7OMnsD+wv2vzqFpXILj8ViJkw9pyRFNzp0B8aBhwUaNOmS81nzA4mDK
8JpTEJLM/JAgJ8TLgnCtx44a8344VsMQY3PKxwo+Dp3XTflZ7DnlwNOZWi0Xh0lGfCJrdXHFwkdy
Grmam6FPp0J30yfOpR3Qf3L+n7t2WE885S1m0mG/F/0H+VwkM02Q2Ix5jVQA/eGX7c47I21MwbeU
6R3z6KvxGtNLoolJzsdHvB2GskmrmHTyk38OT4ue+8Y7zKd8OWOqmYMr2qNx2GodY4PBpIs4ZVe4
7mYblfO00lZxripmruUo/adaMcLTUmw1ZCiUbgwQYI70/mkLZhs+3fojHN+q4T5PJ3YT4N5R690M
kiKRsvwT86KiQz6kun19HT6bNIqZqEfjXXaWIjmr6hheXaL1DFP2gXzfC+Ua06ytEbOLRx2C8qZ4
+a/lnC79mKC4NIRA3JvAQqZviHDLNmGJIeiwQmtGz89zAjuqfcAqpBTNFUVm0yDt4svTgOXHCxs/
gvOJYttoFrr64vSFaGAEccoeW6rEc8GLBGf6Kj7Lh3GN8g7bbAkjA6+/3LOFkyOCF9M6UuuMVB+b
eKf19AkGyxfo4VAacdJ3yuV8cKMwFeYtLmpgdul6C6TjwyxhDIzbtESFr6T0GrHFJoim89UUEf2k
HE8yEvxSVMF6bgG5CZWkY4D0JO5L+DdpmyHcgy6+XEqpHGdasoMsZzDtArrDyjJjjPyuZyJsR+1S
HgB3bJ0dDh8ssQxClwjyECdLIcZ8oLC9DYB2oJOjh/MKKxuXq4N5vFj4nqavd2GKmraJ2aKm5/GO
ol1h6660wBz0t26vE/pXRp+bHtIOUR8g7O0hmGqRXVwoXSvj+jGFRCmELT9IAlXtBBS7/iaevlZb
v/KHPsi2EpjYJgP/DQShAuzf+Blrdf/cYQCoVKeo3NRSbD7PRb7wY8YdzEtR91o3zNL8m4SQiKNg
iZCkZ0IPK6pWC2P8D/JEtpq9nbkldQTDDjMTPQyVtogp17XxIo726AhG7htozozY5ES1cVNH1Nb1
yn6fkZfl+3W3rGr2EVPjjbb7BxpDfKQIoBAWON2pZFx3wj0B4q7ZBpXeQrqfoYG5SZTYSvifg8Vv
TthOpsmm19Q+l4tHraa6WsSlFuDuTSLvSnYt4Ace1+e5BbQvs+DKe/3ziabePeggHOTBjUd+kGuF
NpzKF4KYoNDW/a3Bw0kGEhFAdpgjgI6RvdswtBOVP7ugONBSVh0jCi8d6+c9rbTWsToIf1LifSfD
aVsncNflvmfUeSb0r+el8pxQXZ14cBx1dfZCJ08UDkO4sk5vhXF58DE1bczSNrkFJvzF3fPhcaV+
AstYtTxa7qW/r+DdfOkAa9STzZtQ0Kuk1nn6slc8UpvbQVAFfY5CWPopoRHrtsQXyK7aa/CExHmS
C3JScALinNrnp3jRAFk51HzDBD6xWiF29NN0/MUmY1TcAJ9ty3herfwnY4KTpYA2NFs/bdHA8YBL
5HhHh4X9bSCxnv1ujto0M0ORIZ6sZZ5kkG3b10exGpKSXdBzj6Rwt2yfJ16VNFn/VdGVMI5jdA2E
d9OE2SSoOIxMhppi7hK3why0ioE7Roq79PuMTDolrbhJiWPNfDUN536FXQFA2SV7pIzaScezyNSt
k0eNHfY2O72PdEbi5kUHrU+uvz4SufCjdqG874tFdnaURDMkvtSjfMP+9O1S00iVo8PdeQmw9JN1
24oxrOCQ4u6IoKSiG3YOvPHaq9B5+fzNeC760j9lZpk/zGj3d/nUVnSx6Qh6TaNGA/qyRdDPazQD
NNqFn4TZZVI8H0wdlDmKomUwIvckiPk9FcLQsidH7xtS96ml82QdeHd4sTpCJSN8ew0xroxNzE5A
0+La/4HdFDxIP5T92AptNhnZLunhcc1VmsMsgZh+Nt/RLY1nRm1hecBFbfuc5qDczn27mfYUMYxD
K4HpzDZqzQwDOjiVEhpEiBCCL7YWXnJABLUcleo2r+QPukmIfnlMiHYa8wHyZrblU+seU8g1duKr
OnOJMeEdrN5ZNC1dWLU3x6fwcnCPBB7hO6omougZhobU1/VfRhDgoSsbLvg9yc2V2pnO4F1FYC63
vlYo1KSrCXntNHS6kevjMIq6MPXvGQrxS0gmqyUKZHYe4ky1l3uf2Jo3qZLqjiFCAQT2/tRkPvD9
ezELWbIVteeHAb5c5O09+KvScjaIWaJALGVBp7z3ceAuigpCNvRXHcaPN+N9mSIJsRA69BiIs9+Y
HYDW3EnRy8mSCN+0qBG0JAaCf5/GdWSMYyf0bfqb819SmmbP99G36VvatBeIGXY1yDtFUIxVc3nY
N+DDZz8C3rRN48LLWPx6/vVa34qbT1AuhR1nUFC7M+t6MgYTMUqlyCvWSJGG8PL1A8qnNNiS5hRO
Sjm0rhH/pTMGJBpN1mPFhXtAfar3NGmhvN/rQg7X4St3bQWD8AwXcGVz4Tho7zQtJOhqJ29iMuTt
LaqXXvVEpzIPnORtSr8l9U35Gyiz+21wI8kdQUD5YGfo2zysZvoRqynPwL/bxxTXFI92ZC+Ho/8b
KnYcUVBs+JX/xAnw8YkubByjSeRlaDOB+Hqy3fhTxV3tyRgRAmiXpbvEzOl4pvV2fIgn4OTDzM42
lUPu8zz3ElXL+OWVjlqoNGbhkJS66kxoqeT/gIQXY6oYKWn/gLcS8/VLgwAGC2fujDMqogTOOI8p
0YiyJmAxuwlO/Etb00r35cGgb/JqjqfOAKdgJF0ilvZU5o6+oBig7+AjiY6qEsSAwO9Viv+W1MO5
rRh1oEXGFQhJe8T8gVW+3xaQNAfXE8PVxnt9VAcoFkhE/Qi/cCvQ6Kq8XWFqeXs+CWwkfzvZ47ne
PvwlwGjrvVEsvab6RTJ4AjqILQ7nphRsm8dyxu1tbTX2r0L9E88//bMeVBawUfisDDGqs660iOJV
viaecHEo7o0xfhAqiI5y1QcA5Ro+OKOIp6Yx5WPUSjRfYuKiWkwKxmJij3VknRWuhTb/rMJZ/wuP
OpWZxDCnJ1x8rstrCFgOLYSvfAwSIYw0tcp1wsB96+AXQUHtAJRWOwzXvCWTVkhzTjvtORnuYMRc
ylQWpY7ocghYy/IbYves4O2EFgcUOghOGSNd/sgI+GSORDMMrk1jDXJbE+6qNGkJyCUMxuCswryj
FCdjJOiIvLJwKMvundk6l8GoLVNfE1vJ+zVx3qdPySKytTgCebtF4z0kg4nGD1IerWHhQR4BKOer
fATOXy2v8xsaLQo0V+LI+sef6Q+Xx+FJPvuaZJmTOLjT44+HsWMIxRXq70p49AOiJFjfTSl4W9gT
nvNA+TGgyOJYY462KIU/jJDKDfL+KbpS352kjLkMWbyFB5eKjiDYE85p9ZYjOJsaaCk/LE0zAEoA
08/sG2wr2w7bW9tUwUh+WTt419zot0klQR1oWTkybIfiN4Mix5VDAwPAaCHRiAp2CExwWZowMYbG
bVRUswzLMYhAJppuU/xTwayAVRRa8eXwYCefM+hv0jjQ0gQ6WCMoEHvuDodiWND+Pcg4XkwJy47o
0GKWd0jMhV93PwzEgkw55kNmiMWkgxWHmQrq384UdC9qelUDYlmL86tu4sTprwGPYMRKv8b815sI
tt/CFfFiMKqz+q8EBgAJL81Q0LsQwhJeS9z4pEUIZ3Ghzwt1ngdNkh2BefNOLGTFVcS9+0Gm2QOE
9W2yAjM04pdAf6YHPSD7CA4AhcQNgybm30FJZxI5mefIUyItvyRfyqDkNSikgH92MsImv/bOMVjC
wEcSO6f58jexpXC/sAXszllwhPsqE8jIdcdx6A80HrntqIFq2FE6/KwLp0AX45UC7OKRI42YXLqM
IoCPJosWED+U7xaCmNgvL0Fm25NcxLSlqVzXVMBnaOYtNtGK4j4/iTliS0mpWyLNXLtXpjfOejs/
e15AA4iZtkGH7+oZTzZgJ0wI7GnISRUynjmi8VOb/b9ACiV2GYHjlw32WEmT7uXblU3Upm+pBaFV
MUuqziQkm1rtGaCv8PW9J8Uqh32ynLoboW4Fcg8y+87Y11o+aKWhTMVf0eFW/gKuuC2uHXlT8z6a
kvuMc9zJ+6C/pOaY7dtqMtomMJFiLTQ6jtzZPQXWPDn7X1dO8bZqUaBaZkyYbO9+EUYVV/fVBX3A
IWaOqGt/LfcAHp/K07dvP/p4X2y+0+vxpihqYMrgfRNAk2O8SygGRlYlbd5INBr0Hp319MSZcaW6
83KStCGY04cL0l9zNN+YysaKc7obNVyDu06EuYPIXuIlkL4gI17p6oeU/kP/GarH7i79mqnlvlug
XwqFhc8nx8hhVwVZFPZOtceBJZDuUcm52So2+KAN7WAxrpO5lmO70mqfVdWPvo2xru8wKIF3D36E
LfYUV7izN/4kjVJHopgiJqqldv+0HoX8JFjVtLkyC0xXt7t1i++KFc8v2kHrjOqkb+Ud5OCz5l7a
zQbc885tAJiLq+oEhy0kY0YEy6Mxoq3IWF65ei5LwOMESRnRmvCNQKkY+PLJU2Zvbn2Cl9wOQWEu
YekncK3f6zSbqFJhw2d6MGVY6obRgacsSSc/c4edCWAm+p1l8tVEsEehU3sEMJdZg7MYVKI9np1Q
MiMHQSSAyMmCvWDluj6bcXolcIgJs30MJEU7Tv+Pen8nnVshXORMQ7mC8DDj8jQ/G/ODoneWpxfk
Kivfxs9p5JxTGWN/yJ+aIRWG4K34EYAvCNhsiYJzZtL8g8NEEw2AdDHybvT/kzyARcoiWF7GHkLM
8e8G5/RxhJuWE8gWETJxRDZaR1/RVlA3Pc6xQe8yUnMtDZOuhZFxFJqvHc9OlAToGHtLSZraooq0
h0jWtWSmfcC54rSJO0RVM2rqci+xZV5qNmUzZXxgOO3+dbqnXF+x8l1gtCgFyWYCPP8jBbM2jNuJ
e9bvbHjHRCE8/VJlv3SmvJKvksxKp+pjV/v6gKIC0Ly6pTIsumS08cwx10QILeMw+83a+HqP2ke/
LrZ3HfMqK3VNr+IVnGiMqPTt1yYQ8j2pNdCww1LNGodEa/d2ghu0E5BAZ2nCP60NwkC/8inF39ee
VZabuX3AV+6WKBdPSP1FcafnjuTutppmXekMgIRXys7W+JhGsimEZWfOmfILNR/VDZvBKwuFA5Cq
zQxC2w8c2mrQcfe9PCHcjCur3ong1eZ/NHlU9Hl5LZfdMjvKwCMtu5YBKX7hYdaBs9s+RU3vDijF
E57FIoms7Pe1b67zHrt6VJLqkV4cTXQx2NCkVttaetfNKT+1RR7yHJex+jie5n065jARNxMV+cC+
qN5iv+5Y1AWk2tAPPmbobKXT1JA0adOY4o2EV1R9yxPC67B1gWlqSkfqKIYlktLoxY8FOtG90Qfc
ti15UonnGR+W2LSQBfAN3QeZBtZOOcAX0I/YkIIj+mm5LW6tgNRG2Sdbj+zDYhFmMlamRAI5M3wZ
/sKb5W7rusSNgJMrJPNy1uRSav1GYsMwpnYMFB7OQddhHqR99H6EiUFmniAPT05MEgDgAtaGW8Qa
0kB50jbkisVcg0UHIfFHOq07djQQsCN5ghX55MxNewWEYYJoE0keReX0Z5jnSXNhrnvjDUKSfW3X
VDYdEVbD0y4Ckmv0QtuRk3yoYjFSB6hQaHBaTSaBmVQUXVcsxOV4N8CWK9hPxK9f6ieCPv4fyvng
VZSO+1HBKLmYmGVDfYbvTXfpL01UVk77kQMAYdO+BsN6PT7spTK6Q9jg58mrnyNPU/CtE605viWJ
IrbnRfYwXeGMrqj+8YyA5V6rt+gUzvziwaOdn5nM9GUxLUq1cQRFdirzAMdHKDI8pngzT3BthLgb
IcXChbxeXqsLFwbj0kSb3uIuwxmMRFnj0Mrtve1CFaNkbY6TopxEn/qd0AT930B1iopD9BV9ARhv
9i3873g7vk0l3E3ZJXsNkt/3mvQzKf49hBlEFANCzOwNWVNlgmDYgazuJacLziiF7scDM+v94z3t
u5h5Tf4yv1Df99BcYY47R7RSq5CfZgsFR1Ps4kFwOwYrA9ObITrTv7EC3HtPt7qOMlmirGZ/XnLZ
6FByx24fMjC9ZnKj/fM9EvMzYZvS6QDe8CGFiODE9mktsJc1KExkQAizezVMrsSlRZLXNUwom5WW
E6vnlsrcRCy8brE2zawMt7eYH7Z6aMzVHrNJ3fQ5nbFzASEgk4juXgNJx/SS/h/oOFTlkpRqskTK
6nAc7oaiPerO6J+iD/iiOQhSfmkrmnKuQ7a/ApAHIgh7hzVHdp101fyFIN/tNzSoujT0nC31gGkU
XUWrWpd/cBDZn6ylRyZJNL7QCYC8fxjqjluKLja+z7LrPGodB33jdFfEq61ZMNpyD5IsrEQpbVUm
w5f/kcRmHfzhi6ucKv7JVDClMS0r23OkR6s9AgzbxKjgq5ZkT1e/w1qhfSEO7dZ1cXrwDpQnIngB
NeakQO9zC6TKHEXLi0pDOAE6mH49fGISEBnWDcgGGKyyGG3L+sFaU3Fp1fSziw+wTmRQglt9WOAR
8t8HbyK5FN2RbMTryLDGMQ+CABKmzSRRX2Hls+QegV1ujdRDQQWz5dg8TmxfoEWCHSJutShtNZej
BNTQ01hmnsmeGsimhP0WLxJdITzCEWvacfUezUU/a+W8pHTmPvP8Fmo5yuYn4+9AblhwKr4lZZZ+
x+KyjyUib8GrV641Gr0IeHgM+/6TB7rp2fS3Oi0777EVP39VJtflBnNLQKDlXkU5ze9KOeNcx/LF
1ndfE17cppSPn+uLB9Po8Gu66hL5eag57+ebGe59Ph0tedCQa9fxhq82I07uXi8NOpfHOCZFxmyw
3LHJcdjw61sHJCyZ9jZQ4O9VAxahl7E+8o7ItCLj6xy7tPv1jEUZz5c6pmW5FWVMZNRP3Nx0Xitm
MsG7Zk2dv0o4fH/wuIWXKHK0LR7jb/NhMdp2Y8+QZ84yiC7sPU5qzi1wvgGcC7Pu6XCn9+JlGulG
zuGZIpwUbBvK6vUvSbMvPi4I+nsYPfNBft7sw5BhWHUOnM5wzW1j0s4j3Yry92HSTb9Fj46NnZ1A
EGXxF8EHGD5tsXRKpS5eet4eoJnXTy/2n+RyAaP96fyWS3w3+JYKJ2Toy0YnplIkqLbHePDUsDtP
DNVh/i3nfwveM6dD6KoTCfTHNlIW5960pCDtGNs3+pRNTOizeW0ajz+6i88oL1HZqUaWJudzl+sP
kzyDbDmJPULHOn8DKwDpZdReaOHtl5eI9ix9CvS1WsfhrYbWLeI10JGw+0h9v8pMjsK92MCiyMuq
gclx4FophCBlhg1bfwr8qfWueFYsOXDH5MVCNg4PL4B0Ede8up53AsuNDS3+Q9s259leT1frXF+6
WPzYEpvoS5ZyukOcx14FfXZluAjIp3lgaJMOlcK85H/V39oMbkgWx/rO78mMi4YnoBUCqjvwSCw7
GUaFyOQYzl6VblGOYnuixf3RxD/oprPcT680V6eg26/KrwIAt8rdyOQO3yg8JuCIMn1YaCz3KTKa
QineWjvGA2TNVxETvaPX44mBe4mLiILUjflCiIj7xhL8+hYgRNysp07UYZwiqyv8R5QOnCtSKGXf
p9nPFimuNErlhsGme8QRmVhPYNdHUdPHRplQ7rPOOTzhZ8wvlOPkjreFGzl00Muzivj28QnWYiDg
59c9bjAsLvs9sdEWN+E+3yjOHkTDvao+zQY0fAy68zgp56T0HL4BxaZaYmUdKVbulWecxniS2g48
MQ2wrPrkvsGJX2kvAcSdPHL4PiaFiIVflFN/7eR05fdtFBWXEQNENq3wEvyxLLEZMS6ckcJgUjVo
dYyqwsyjG6ls4JfQA6tJ3B1uIG2skgvqb2vjNNGR/GK+5VOdX/aRPhKLafuiRoGXq//QEKnlrilh
MHvZRSwjJ0JAMZyVlfhZbxrJya6K0YOqp3hBgl+A4Sy1x/IqnGyb5wveYTKYqjLrMdQbr5lnZdMB
dM5HwGfUBbKMpaDWhhx3gdzN5etQ5rAMDTnWz1OH8blaLFLVwp9a4wu1ZUktlnraGZCtDjF7RBOT
I//VrWxB3GJW9p9kFB8ugg0INFadyEKNq3PK3iKtOua978XHeR888kbShv+4bENWBq6Wlx4DtNSC
wT6bqs53MR6ItkOpcOGIsynVyHSwoCI0mZWvxCPqV/gbqmVTYoZDm6p4mUai/meNspHFQmwNYmv6
YBXXtB9Akw1HnuKBVeWq3r02qpMX+lQ2o+BdWoeeJK396jGD/ESMPA250RYjHd3lsqrJonaer5cG
HTEqh1d95o2nwb4XZzsMApYqUbt6xFogZpiVusCWgyanogIn31RqTSy/pDJSc1KpLA2qNz2wKOen
H/iJlV7Lvm/gY7c7tJ9zKPmuNe1n5aIn5alp4oqngogwgWmjirck6LrTBs8p3ijMOIp1/0nr70py
c/+sQuhflE6SlJIFMiybo562ZIEOhtDTXP76OlV0uQ+k02QMZjUCIia98EfiarXhtF0HQaZIgcv9
CAgk1re6Xx+kPAiyRiKbxhke71E4LE6csaMxrgRNh/CY7bRuD709Tqdxtf53J253XE3X6AfNxnpg
WronsxZE//CRLTeRmbDIZEx2stAupXG5bcoJ22CevfxpaBrvCYrbZd85d26b2iwkFnuHKbi+rjg8
YA8/kfqwemLe+NHjbuWBSi7BGLo655217MqlE/YdCQT8bx0Hr9U3/ah1j7NfILN/kYlLlJKd85yo
Hpk+bBI8BE+cFTbrsk+JLsEFkSGEF3QpqnnPf1Q7eEbK0CUwg1ehZ93NTRQCgtx3AlVU3lIshC2Z
MRF69/YYpU0b42dE79nG9EFRdJh5BmGdiqaggWan4jTa+rnRUvoxYnin3eQ0VvrAczZhyr9FPBnU
MqWArNoVdNTkmCejMO78xDjBtrPjBu2Q+qXNPLbelhlsE/r/NQUs5n+Hs3glokLlcBEFLZ1yqspc
rghoCiY1xRkQOai1iy+PM0NxKW8D/69ZZLlHOcr+Ojw6lpYJkAQxYEQp9dyTW9MDEdDxW/pwP5m5
ZTUHdfkQ6a9rVwrkmUVVsWoeNhOUsk3WDHwo5pAOAPyy8g1nej4MSkd2izCWIv32WeqpeauERYXa
Mj/oJTYLF7IYjdT++1CwUljLdaq7Rpf6YhBfrn6lCXUNojnoXPCZE8nxta627YvZ8n3IanFmTyfS
g7+6PsSygmvdO/jYDwDhOGVTTHyEmG6RQanoTNt8PxnBhxpBJ+9mC7HVjvwwAHVeKR10Z6Qfyby3
IwKyMRh9fpjNzxmiXW4AiN5hsS1PoP/jaDZO7ut+Ge9mS/439AmyrIWzTLKJ1TXfQ88z5frQoYbN
EIxjs08gIdbleWCrWpDMzxKOjjZjp8ty7JSsu5fXRU43k4q7Nn68NKtdivvIek9F0J1ya4kek89x
2Q5ga4VbvYVWk3W2ee6dlSBOhWtgTGXyWj1oQpAFGzixrOEUCZ0GZ1dMJuNb8XeBmFyITAE+I5Yk
tugJMeBs+95qU8LrKMnR8z2UW2dcw0bBR3/e/njBql+IkPlv5LpezvrCtqvzFxl65HZYTlOo/F3N
3d4Cb8aIOn/mRCMdhN3u1EQWgRTOAsTb32tBqM6ami18gDV8IQjw3Xx3S5Uo3SUdq99FG5JAUEV4
Pch7n6nQp7xUSmO2+iRaCAF0jV3oM4jQKtO8xcaIZvWuYAKwlLuHWtvrbRWXg5D6XnFSfHsjCr12
8lSueh/cKMDyvR8xUFH/j6SKbwAgGIwufrfRVYkuI/sTzzn4TkTsVL0uFPZXiDXvi8ljKK1W5Pw0
ZhjWW0yIiZFk6opBA86vaRjeV9N7INDszLSphr8QIMYRvNbndoJZ/SPWAv/OHu/1gcywS6PYdK3w
JkUCBvICPwCcCNpmeda/UKPMSQI31iSMr/46tHJLtaukbZpVQF7vRQNBslzyCbXKwXAU8aVQU1tX
5Bedt1BhyfGqzrQd1S+I08/0A1gUJp/Enm8t+k+6MUey3FSsywfnQ+NvQ2qgzRE1FL1Tg/PRp78r
dvmmIcbZpnXEXKgw/2W8wxt9fagtQmA2IYlHxPcoPCPAfqB4940zjI1tFuQqpYVMyC5KMYPW4aHk
5bKh0ma9zkUOUd3kAQRIy+LjtzVRcjd/RLxRpTxzejt6iuwtQ4xD2yTN2cBcFjrWRStkGQ/CWvgs
aBBs8fohCXPzRbjsLBxyRWswre/FEaFRVzHUW++/p8RsuK6/JFwdjGQBWjNCd2tH3I7jKYsb70S5
UhsvIFc6xP7CYVcGT4PoO3HBNjwY23i68LQXRgatH7Q3tXbQ4A+CQFBpAOpvoqjeR0KwIkN6GcG7
JkkLzUTNRPXJEg3TFhx9Eb/CxnhIAAGm1RVgXdzHFWWSTzrZSeHY2JWxJtc+JUA16GEV9wrqhLY4
HAyMqzo4SGspZGObJbK/a/e29CdkxoCneFbzgunFsBjv/2/7vgeX0KKPBe+FeeX1sKaXtUPJwJkf
eRvZprHIgpl10UzZ4szLSwpOP9fmaSb4Gq5qDjg9KYswzWAAR4lRRtDqxuoDAhpltjIWyo2Tf88L
bTF4tPFQUDl1t/hYKsGvqtLGpvLJwBx1OIdEM8sI4iMGAZTflAGQQCWORmZhJRMxgdmhq290osju
V6o47tLb07vp+QTD9Tr26oB8kY+Y7di5hG2qi+AI/sBaDk6Um2HP081EcXLL6qZNgpmvZV2EJjRG
5F5JczmrBg58HMX0BIcXogLXI0SfYVCyr8/kB4UtzXRtl0kfJMnLptDddnBMBXiGxiQQozjOh9YD
7utgViD0yrJdR68s4V8KceWtxKiL9VOCyRKieGdFQSrDKKYBzXhFtY8YjChmXZZjzif33cY++hrF
flhqyZ0GnEXH0W3cVkqfGjMy8Q5qNRwrJDqLTgL0+KvQNHQ69SLNIt2toQufEYhel0jEY3yibXGm
JO+x1Hq9szNm3osQNwYGH6mCAlc1gBDJLwbBTOyGsON0/YbpnPe878WJClJ34iFnsozRMFcyB784
iHmqZfvi5X8bnNVdTo/EG8RGBT2y1GNNLd8fYCMfwvD5ot+6DiXIxi/1Vrs2ZVRA8NDLNmKJTn1J
jIkG6BScnPW2hGiFWyxTHiQIScrvcI1Bn92AbzeB6cmEqaU+M8dBbAX40Wj3jZ0D+c5/5ILE6I20
2z6wmYVjYaISGJo2u8/iPq8ieaIx9qDsOM8q5vDfbsFzJFEWu8bjuzR2EnLZvGN8ojlmqAa6F3ZF
hW0A8/ioaHOFra/u4N/S/20BpNfE18gwxSZKGguXgL85aGyUrSmI5V2EhsPLkZ+qzIPeJK8rN1Rt
RZ68v8omcdEyF3FvTaq5gfGCeCgykaouvm1+KpXee+MT90Y+HPq4R1JHybM92XbpdAwh0hDt4pSl
dej/hWJmPkDtjl+Hqq4NKlGy18SvHCRhx9dP8pUeSZQXRuy72n/vL4W9CA9wAWED1sX4S/6pOaZw
z2KyrsLOVOvPXHrkV9SUlid78Zt1247UTY7b0OhBvxOx7r08WJqedV3App+mH3UX+xGo5B5JvUO6
wW/5ZbSIpeb5JQoxdS88bYKYwC0EVkJGWs790JyrrI2Ttnxe8yOsx3NkwEFbuLaHX2D+Uw+YTfoE
6j0tIqvVz6cpRqNJ9NQHmleEGQt/oOqKIoiLJvFyFQC7dn6+IH4GbYY9uNkqAdhHBijfKg3U8yc6
6IqjXqbbS3MpE4ToaRfBcUYmJpmxUNRKpKK2dDgknU2AuAFZr1gkjX9lYQTCZARM873wh5NZtHzS
MYj+5IqFV6+sPJlfMEnfabmhacF3wS/PETnEShanov5PpU1GMOGOrSLJtnJlZd43x2lD36mptYtI
heSNdeOZG9NQeI2q+apqFRJpTsiU39zGDt/tSdNnWZ7cnYgxloY2TUNLS9kO8HR5ldlxw9f9Qaf7
8Vee485hyj9dbeQLc1+qKRB1+ttUQg8P7tMuYrTmWoYTnqy/CTNxwCw7zPYIRet0ryVULaZhs1XA
z5htmxpro+cGwd011rKdtVnSQVd9wDuo3bUEw+s1spHo8pRJgEvdXb8ok+Sy8v3Tv2dgYUUSK3rd
sXJrt3CWvLyMqjuQXA+UCmg4jr6xDwAfyoTsS/oBVoUVRm4on2INDkP+VD82wkg681KwTV0+uNB6
+/1oPm1Jlb4rjVPieng4AqmtrOIf9wWPSTVUivE2q/+BYzy7BxTL3iXaMOV4q5T4BWtyjLCR3+uE
/aEQdosfpjKbRTrzNCzjz3KDajV5iNGtuHx+ag8dMJ1qvG2ClfqUoaUBl1hLX4M29H6vL/QJG/+Q
E51qrkb0uUlgGEqqBqedH1AV6ybd1fQgh/xZu5q9Ox4MvqodIh5JDQBQNaUmy7o3+ByfkPEdqeW/
+Yqew8XEuenuWED6JLKMTAYOwRoa1uy3O847HeGyUPVvlqpzeuxFUbzAo5rQpvTn/xQEdq2VfpbW
VguA8A3kKPdqqDxVaVopFcN9YC/cCWh/d8VG/s1E4uZfYpAU+2B01UvMaAArfj3ycKxi3Q6vicTD
AGIGY+LsERV/1Cf4OAH/yGJJXAyNZAcXuC/f3rdju0Qxskg25Uojl8IEtt0JzDuDZPd+FDXbhhwa
tgQKQQXgMtn231dMVOzAumA2SYjp6Lr/jw8zRwg3kSeNcTZZlONgvj3Xw79UAWlh5lzLxgIOTlDG
FnQsBTdKGqwSl3TFPtB8A3CVNHOl6HPAaMe7uiwN2f0M/fyJKOGf0tfJ2awGmT3FxnEVx1kwIW8X
G8zAZkumjYJCs6f5SuLdfZaaICekbMV2g8EKeOD+/UFKhQnnn2/xRLCgMrt1uE7f7Ubfdy3hrzeF
SioybAxf9ReL39B7HoO5wZZJnV5hzP6jUxyTcCNz/5s5XnYyk8EG5PVvYLC7L5oMOOshsayVviGI
uiPZTIU3TlbMpBIk1UjbJapn7kZ18ad9J2VhhBvVCDN+Kp+cE1nKBmkxbQZXxshA2B+S9yznayUq
5SojTBqbdKaoAoWpPo2BVTkkiMUvB8zGOoijZS2/OKkezkjpR636ozMCGb0y8o/vrjgmrqG4apJp
B6vfwu3/MpbSyLLIKa3j+uJD8ldvG01JhA9SpNUr4E0eMZwI3Z5h815YkP53mvmW2WQxenO7DD9w
jQi5re4Zaamvr/bn5WsTTe1ofHZoFBNJZ5vL8c6AJK0X+sCHjY3KOP/uNtJS69+b4huBCgyzIxe2
iP1MXbKNez8FdZPsnKi9mSOA47HluuRojShQwn2h5mrmm/uevDkyDlPZGGL2CUy/DxWVShRl9+Mj
GmuQUwfH7dXjTH6IyqNJNOG4ahjPWBinE0lLovqtHJAskaYN510tBAWoL6pkxghpQfdvxXWUp3sp
BCmivE5zEqHivICr64DUisUanbVBqqVF8GTBu4ssNS8KIjOPz5da24+9RMueJPU/edhIyFu2hk37
3jcgAF5j1nBoj1fu5DC624VB9T7DEjlG3fJnpVrUFr7SvQrAkwEwwO5LiE8PutjKrSQNciy51elN
Bo4h0vTZF6Qve6xV5Xlnl7yWlomPSQzUPWpIwor1kgPesrsJ5+vioVVg4q7yoqZ2K7Qg3RSOPFQ4
Zc2vUzBVzXzlclNmbnzgqnzY9XhTz+gSNlWA/FCm+atQ2xNgdw7SEw7fzyNmBbpWLFG+AYtY9KOU
Uyoi4iN5T7AtJp/Nt7OvPoOPouiQsvNI6ExGXoBe2NMSuaGuulV2b2p9bB/pg70peOqy9qGMNcgn
/rhB7baBdtJX6wHl0GLnczumIrtR6tuAFBdNu38p7lsCAZRMTwt9dClWsrid1CYdm2l0jas2TuZ1
ZIT2JibWaUtTljnxMnIIcitvPX5mZEJRDcQ2EOqXQXCJHiTMS6PXo+/0+3FwkCvnJYuPczYgPlU3
ZYAuH6yx+ke6oGaS8Z2pthis0ov0ACYtVaHEpJZ8hZUfI8PMfVBrhAmoF+Wi1b38UuKRwqBJHg14
hPj1GQnbnmZ2ijpRBIowdE/FfzgvoniwGIeeKTmfLl8GSWlolPODlrlquwaM5dL/RxT0VyAiL07c
OCElcFaTYoBnOYFaZMv+AqWnCCk+HYi2u4ijRsBTkdI22JTF4UsNElcYXmi5NJme+Esm44QGCr4I
/gsmzY1w2fPzKrTdzmFkqMtzDhJN6HC04Osz1YCDLONIQupSnfDu/wVbxZRleFMlELITMOkY4XeE
YZuf39m9TtfW8dmPmDrw/G8iH/FueAw+9BbopbY1bp8vv+NH5OHyarB/V3Loh+L662jQw6SkOtbg
rPS3i2Vk8STc2QMavI3FNU3ltr8oDGUxYrMD1QTeUIN+xm1Typ/Z5CKfRvJLfIJLXWU71PM6lUk1
dNISyTQDgWIswie8FCbQ/HDWUHahpMrhZogEDEyuCtsHXzdQy/l1sYghUhf0Rqf/3tWYX+v8RCZJ
KwecPZA3VBH9smRaRsezgGIlRQHn3PtyAai4TTjLKQz29F4ebFkJJtHJpiuVIPX3p+MnLl6GiaLL
WViCrTfjyWt1dE6jyJf1HPKZyG0Tm5dLiFN9ddsdbZ9/0Rczmm8f9+QGpkVbPFbq3L88zwDLIuyM
erMWKp5J5OefVT1eMPq+wCUgNiYmSFQDOq9HpGB9bEJVN6Am9hzr7HB6MnPcYwwuKPTjQA6LnK5w
w9mNVx0f7kVE5crm3wofuzetEwnKxzlYwvzJpcRglID2Af4kmf76EEZAIOGs2ChAbBlk18m6EUQO
fAqQAP6tUMaONoxjuz0zIiY0yc6uH7Ps1hXEDDH+poQQ54tMVtnzPd6qv7d6+MREkx81sbetKsJT
nC4hIGS91uVwx3izj3iq25Op2QrebEnQU359EK4z8r2gB58S6gDRZ0DR29CoMe5OyjdjcHRdAZXm
MBnGr5MoM0Sn+98s/jedJSFnyqyShFYJtXwXCRGOVz0EUEfY986AjlciDiHU4Uro6hUXz+Fsl7JF
FrphNTx6jPLFwlB8Rz7C2Iez9YD6NaLLhA130iYyVnqMGC05EEHQrgwW2cMtrWOoTd5W1avmlZoH
iJQAUU2WpFAWb/p8z0uO1gmdVFCX6R1B3Y2vJKY+dMHHiUpwMlMu5bC60GU+SSTW/zwK+SJ7Jrv1
9E6mmvaLWs3ALO1pNxgCx6Ery9cqgygHRlviIIKdfOKjqfr6uPZAjeetUGjbrbtjVG3GMRxtaqz0
j8nxxsFVr+cRqdr6enB7Y67KcuoA6oDQgrOM1npFZiV1fTL2vmuzWmP1UqiBCWtgtUXysQGgNwqL
/OJeikeCgMbylDOb8ru1AdXFbb0MMuH+tepaYV/oGJCguY35XKuiuj9UvMVRsy4rfApwjg2NuFxT
n8zN5dbQ01v4VnXNKyqo5lzDO6fefvlVoHuwL0fhjAoGcVMXSPfTV854KewawwJ8AIN3SrSLIfWQ
zJIDNnSQ0Ufa+TsL008ZN4xwW/pMH+gWY8tn7ZkxUDfM5mTR0fV83vQg8uTILygSsfq6lo/Jzb4t
KmiqDSUqoaXBvT5kIW3R/7HuutqTMAPQKA198VCDq7t3k1Z0xQRGKUFrpZFSzpQdw4v/fylNCFoO
VwPSthoUxIyIAeDJnF90g1j78azrm1jdCTqqiuJTFktJYghAgf5ovTEhXHnUXLcDcTugvCfBUTPy
upVP0tkrTby05Z+9gNpXDmP0sOZkL9rB+r37w1jLmz3k6N5rQWHQ300YiWK09bBz9froMo9JJA1/
TUaNUd0zShRXyACAHga4lhQxZWz3SrTTF4ccmXrZmpigelGizY2jxPoWd9fNnT12kxaat1QGjVSl
8pe/YoXJ+Uh8pL30QA5iBqTKmg0RTIUEQw0yftbX+8yXlB0RGqU/ABZ411P17cdrMsexkYAn1e0A
D0oeP9HkrfnIaISWMatP3aqksp6QP48bxqj2x6BJQfh97wsPBRN4YA32FbUcKTrJl/nxRd402U+M
P1UDgI+jGLc7dE6FdMM24V1fmrG8bpw2CirzUvEVSP3P/0jT8JTFGpoI3ViY6lEi9txQ/p/PZqy4
81hWFBGlaKrfRXcZO5Uq5IvOEMfvffOpMGX8z4wngdGPviXZhv+aNNgiO1GbawRhH0rpSTu7g5wx
xad23vxZj9o7gSSjaCCtyvJj3Hia9wXo2xHJH7mW123XUrW9/s2z+dDFfeBiVYDs8ppNGwoJVHLe
IuPb0zj7oXCji+EGOTNfR38fGH6IBvJfIGoeqBfICY/9Hn0IY/XgeTnnZTztOaWyB2Yk/W5DnRwK
pUs3YHfx2obyAhYHrweVnFmdQUGlT5uteIVhVQo2bp0E+4SaFAPmtwF2E92N67sts4ijRCbHHsv1
Hl3VVfIeBZTeajfVQ70ioIB5jm1cOuSE9Y2f6e1vlBRxbd0HAyTki6VjR6HHN9ehZ7PrtMonEgKR
RefQQKLm9iJhcBRW5DFg7rchWjPqLBYQYn3DiFyWGFfM/PX3LHfJv4T9vWsz1b1ATKbDs3qDYDr3
5veR9v6ezaBQ9Rv7wu+HMLYnyWdkJd8Rujr6lEiZwLgss5yFKrwLXankmMRbGVvIzBteaqR/GVzw
TQlmc/o58g4BRS0NmjcW4QK1zXU48GRMUzpFHMM9DSfeXmNT6wWLNj5hun6Bzkug0HDKuSkp3lwB
aQP49rPnqO5V5vs+kb8D6pi+f/U9b2iP1FzkosA21fdl1v5ZeRRowGHIQ7AGfEvSYBr2GG6/yt/X
FbtYpXGZ5MSyf+7Z3RIndlPRgWKWC4LwHjLtcYHDSjhmS1QKKk/e0s8G9HdOhk/Zob7cpnckSB1y
UC/WZzeZKfO7Fuee/aWD1gMEabWRPAnBG4d8RpH8kZDq1WLy0hHuZ5SRe+ti7Wdeiso5yql+v7Wc
4QvLjstXDCMXOVIvs3wu/SQvTEH4qUu37bKbgPLm/LdxliVn4HJ2ORX0VhMz1gEQ0pwiWrTWonPQ
5w0hxC9usbAH+kXR62X+WL0ZKUdY6nPWTMafnCfYBZ65ZPwqZkPW+gzdVpN9ymVIHg7DKdU5xDyl
9+Cj/46KyPQtfz6QDtzV/yp3GsEqSaamd0mRXGyyqEt4dQMH/RzBA2Wj35dGWg4j+GcDnWmsryzl
btBXi42QdUT7vpZfpgI2jPIv1a+LwGD6mL+r76gCwXyJzeHgihtUJHkuwSGxCQbH8BRQKydPFjXU
eyvZef1a2IlnTVXz3yyv8iZlTV/EuzP8MqWP4x7O8v2txbvRCrAgenTL0/BOQIBa5kVhdMd/nrHp
W1HTxaDOy+NSks9fe0MXY8SvdiXDSjPqabqx87JgKHhFqRFyLOyr4VhlZwu7MFxkn8go3Y/1cb17
51uzGpsJePLEB3L/rve2yyfJy4P++vFh73PS35S2mdY1uFYgmkscjP9EGRKKaY562jQE2p9wQYKM
CryqvioVePw314F48cjVpeqoW8It8o3329Fxmy4iNyJ6Um+fArh6p41Vh3aSsUnBhsR22yR6NFqp
4Iz10VttbVbgOfZTZcWiSmATdeGD/fvFE15OsnRtjn/uVkd68IDcKBxhfUFnLv933U0pqUx0MK7p
hX2C6cWnk2hgws33eT7f51urZ8C9wOeNRSaPk07c1qixHYBCDwgsuwTzK4X3wmK1obf+3tcroEKA
1Xi3IQGqoubZ/h6Xe2ni7McFVTNpXV2dJT2NPcYCvNHLfD2ScNsBmYaNoOM+WXLxtWbV9QO/OZYh
q8A2ZJn+5UJkGXfkFdybvl4kz3VOdU/Zz/1KS4XfK0XDspKcXddPwjPysU1n5ewQZEnBBCfz7eO2
Yin4jcdJx4P3pI/oXbxG/ycGABKezVenDKN1u7LNJ4qJMxh6EBncQ6w7/vDTvuOTUQ/kkJPdH59c
jXF6caGpcXBheesCj4yyUFdsN5UxhZrrtM6fcRZ1S9cCAMwLh4pnZpo2eLZblymSjfdV6IIBc/KS
ymLAsR0ImaZttWUGv+EOO7AXkMvC6lLRydSXlaggirJltcpc83kCfICmgxmfHzd9+rEm73ApOLVL
Epp3jd8DIKGOC5nlgDLsJzWM4EtZ754DQ+S2L13M9/KQQkp+ia8/nsGecIwYacP3A8Gl+7FGEHv4
IAAY0yPIFodupjFksPjWFqYMcDBGHeHJyIbrkpFt1ZlJZdbQsNyEpd74i4L2XklrV2N+1TsBxyK5
Dwiyk7zio3tFweTk2N2sonk10ACFOCQ8/jbYokr1WZaPf9yBEqUX82s7wAJscZB2CW+24vEEH+HJ
ufTuSh8sZpRh7/LZPvS/RCvSE7lM7zx4Og1FcZNxCTzEzaXF89B73rmP7bW1R5q4m4CL/EzsKYh3
rwUlmFtvoJZhQG75co66FG3Q03V1ChYnqsy51SL5LneGfNZYjqO3ni6Y2ZbSPEQ/RP4T4zg0qOS+
fVI5i7L+Uh3EqplWmc8mzTcxQnFJT8JGaLoohpvohpgkZwC6CUTtagwto+QU9vtpzp3j42zxLSIR
aS7ZBxo6PvN1uJPGyX7py5yWDTgbyuRbnd5jXQjxupsqcIZJvVBsOpNEUtwk4ONEj2USgV6WG1IZ
mEl/XI/dj0n1AnfX4Iag6ql5WtkcVyeCtPkUPUANCK6U1Ku1+d1rVTwjZFqur8Cdhainy18X6GQT
Vo3IXfGPeBWRFrJEz4HXSZNcArOGNTwH6GU3l9eDE0bs+Sn/Aohx3wAmsbHGbnPTX72O1RowwvRe
ZByetK+vcP/JFtqMu4Mb/xt5Rl59moGvFzRIBzPAJlPvWiJF0E/1MJf36CnCo+qSpBp0O83YMb3t
E3NV303rUAkUmxCVkgsCQLPHRIItk/rfATRD
`protect end_protected
