`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
0USWSUGxovGsyBJteYpEoQMYe57U7EVv4KgCh0gNmqL7ISdEU5vCT1g2t69dXIELm9FPt2ujZh5y
sShmvCVBNBbTOA0b+ysoGqSZz5dJp6l47JuilVNYKG6UTE3/dlU/d9L4bsUQJL8uD1xhUgWNc7W6
rbmnpQGvUdWMj+k0FeC+Dwlz98mDXJn6i5SUp4WQegOGPpB9vIpWXSk0jbpM+7LVmmmgDzmaAKNM
2NMyCHHAt/2ZahaXwMkf9YNCHBq2tzknceKKL3SLJ63+D48dr4ZdT9pPZPhsqDm/DqzEpKM5WxGE
bcIvVXyvqGBVMM4qwEOkGPlZ1rOeGSmOqQDtHxoOpQDr2aJEYuVrNFOmxE+/J7AWaSy0q3Z/Vmty
wdrdSTs6hcyGwMPuhp+SahUf/tasyt1LozCSYHJ9geMt9gG0uDiY86dQ1nNVihdCimIjO3MudffK
Rfq1jx3ovndkbNxIquDTX2kCTFKsP+nb9jPjjLr9sxS3WcsojRbnHnTaIk8vcq4qvIuzl8rAq2nQ
AkOlX5ifZji717B3ujHyCGtqnGrgULf6FmWH0zG1VXGMfq4XcR1DH3+ARdKLiwRuWJT92DTtyBkW
yJ7tIseMnepP2vVmbr7v8b6thwPeEM5MjcGiEv3rkJqhrJoDUFZxVWwczGCtPhMSABZpaZeiSLPu
rXrxwsaxNMLcN16AUbkpIvxp0Xf325Zy2mdnEFfNLT92n1Pt5XNdkvBFmcKI0fpWpz956nom5Jw7
EndoDZK6pLXr8bvvZ1urjRQfXuUI3kklU/kb5dNoA+8LBOCBaXvNoY+I9gxTvRnymuXp12yHZqcR
Y8xXcs0YwsQ8LQpxMfn38pK915FFLiKm/T+z8hvyY0Bjy/SJpEbOrl5Dd1U6bbhZyrysDzj93Bl2
f1rfjG16HmXblCx6kN+ihGXNaDZKBWvvGl8231MmqiIzSKRwlUaAzqQNI7GkTCI2gQhB9mlNM3pF
CWw166jir/q7wnsZhTG6vjAKaexDFXJnDV2KblVHfMsLTWcRUM8x9vWDFoYlvkT7JqvvbqsarcW0
i2BfkgXIFFGJddmsKX0h/mMgVtlWUSqAFNNApWNpA5H2q8dFT68DaAiHBNaiUwii0iL9E3693q6w
tSuBahrrb332Ky/sRSQ8lbiyyBhJIHAmNjxJcsxbRMFC7QigTFlL1hH/SU3B9M/1yc+MksqJiX3C
pZ6MrGn8VZTKtIQGaqd8eEK4LopbOQ2vGuUKFyr9Zc7Iax13cIO/55XHg+uGk+XPl1zcaxvBQiPX
uzwz52V95luWXGJhBqkQmtQy7G7CNWJHaRSbo9d5STQwzu6/DP3DgNQn1/k9mFQPDCYT7L3B+fTl
9Cm77kkjl7sgGXkAHkvN8tZNy5FYgoqRR8j+p1RgXTKNrC7azs94I6GZuQo6tdKZ5in629AKfsfN
ltbzMilqFat1PVuXRJOOupwHPcCb2XzR+HV6b5TSOXwAPmcSmzu93D7koYbmsGa8+Erw76opXwik
YrcXlXqcXa9stLbVxyRm+BknGKPdXJo9akg9udTtxn1qD/jnP6nvMOcG8t0gCn0xVSbPCnY2bjgs
OyScMMLFWuBPmj8GDAFTjeLnFN+Cj/9wvKYyZeBkA839idtmMeW4ULaA2ojpR+o6EveKp58pbRVo
DappdWsR0yrobimUjb0kQ009IStzB8C9iFPZbvlnlJ/zrzMEfm3QiFhSrZQdC3fwQONechFd8DAT
/gr75MzvqrmuR6iY/PK2wA45+cW6AXpyeTwsN+0anKDvReobt2tds1BvEXZOpwXH+K5Cj4eUsObX
pURhx0GEo3XDZw5Q9zQWl2i6cRJfpqTRRGv3eFTQMpRo9ZO1vPxyyyjbPuURJGWocqVrS75Bw5EJ
DLlHUZrtE7Jl47cj5uGi2kfEl+IkB1P+S/LnMKA+wbUfOimTb6qWAiQTC3spz1gSh0MWV615xEX+
1sXdmO63UNt3yIxpaHg9Z1BWt8Ga8pahbQ9Hu8FUavari8L7K7T0uU7JlhCR90LIa27C0r7hQXYC
VNPSqnW5SY6yUVjD6kd2c9kxdvnLQSk2qt1mOpSvMF6cfMAQ0GcsXyXlpK7RTVPc6Z6yvcAbs2jT
q0m4BJV7X8SSU6clugJfqzYbUIyrU8SEsk4JRpyaWxJb+r+lyYLQoh3xzgd6m44CRSyYiHK5qehn
Kiu2oPcCblNlzZrdgPYv/djACYhXQ67iyT2wi+wUzy30OococuSvlqr/HwD/RUBAIDkx/VZC8W5r
63Vzw34iPotMG3I0bPDTH/knNDKUslUa6FqYVx9R03rzw8NzFef2ka3UgiYGoRNc+9Dog52TiwTt
TxqNHFROBTQQ+ptRnffy6JnVW3oOD5G8wNfdT6G4/xZ8S1bDjMJ+z1ujPEwzfzvvhtnSHAAwMHjx
CXnqxjp4RxFI0S7z6sz8hHsUNy/IXyYyT0dgFHRS3OD7bsVa8e7yMQ/icOXiZLCDVkGG3XvVyEtq
88D+VqFQ3ukqF3AwRgAuHkYf3yDmOkCqCG5c54YlQ0JV9rivRXm5Rn61H8UcuXazSlzd1lMFvmKY
Ed0PCgub7cx1o8WBY5ImgWu1CAMbMck97QDbq4TMBHcYKxOXbj7hQzZlm8NsgIcppl0WCdBYeUrL
GAh8f+0ZMzUzaK0utjCJJmW8BkDwM42WjjkulmVASPwgPFfCsyPHxHPGGvasAum6QTfk3y41oX5E
WWFySjqtMG+PtEiNcp5Bw9y3bBXrLpBDinbUqxALcwA4A//KFms81MlZx1ZamnQK5985DDmXU17P
Y4g8/4reT4983osG9BsZRYvOdy2wzT2dR+xHPpLFqlsssLSMurE6ZeJkoGxVEpCuRKwxL7qelUqb
aB9nZvaxg+cZdiPyjW6O+k8L2J7NQOTnWFTRYTTYdSwwLazQwtw77wIg7NUaxCitiGjxKOfv5/iE
WzzmdZkvm3I3GihaNoR70cXwMHyKc729XHNHPnZ+ZROcCuh8NZkXRlIqXhyWOMnBzlevGuf75tc9
/RBYSprpq03ZauRFKAjNVTxoz7hOO97TN6I0RYp+0BNG+KExtulsSllc7UHac6SwJovsgctp0k0Q
y7guZa+OtJBtJFBWrVdJ6s/z42OSZE/USCwbZa+/xzVXQZPydW4G5LkqvavA1L/l0dHFJ/UXsgiL
cm9GKWJjndKsiCs7uuHW/9J80m3c+QvAx8HgWSxp7KQ8ycWmR7sCRe4YzgTbwKUwRyVNh1luM2cm
+nLnB0Az8nuZNPJe/PUEZmUs9b6EsO3X0/r/+Hbsas3IDqntrsvl77kBHxXBcu5TC4YVXeuQ6UVH
Yn/pGmhOAHsUYE55E6Uxy7CX2ksb7jziQ/PdxNNJpLWichfec/W+0bU48f9jSJXbtKWTw7olTNnI
KTjhRgqOLuhSnPnF3BhaG9nlSzEfFBBBgLMf+DujXYDKyAaqjg4H+M4o0eQ5MGfhrDmfT3ut3uHJ
jzis01ObioUk2ZSTbTn1lMEAi5XHg08BZ2O72xem86n7yn+ON4oi17smovdLY9bXYzGfAx3NRg7a
Kg4tMnVrI1FaA4DlnNjSdc8ITMEodWe9A2jlGai/YOuB7ZmpqhN0iN+nL7Qvf398WnSx7lWlQ6zz
5rI5jExFhZSqtzssflaD0DO91MMm6y19mfS4yzgwpos7BZssTVy+lMLJ6JpqDl7AQGYilosnQ/Y4
EjXOlRRQyc662DQicGmwidwGmq5D5stDnE7/Xh5l52H8aYNC61gxW1s6JlYoU2yFBV7366Sk6ffD
x1EUsXrD7ufzHCepS/w6HxxwUaMp7ww8gwOa3YOzw2zk7168FuuovX4mid8npzBDpVxYCHJhyz0c
MXbWKpNJwaOouksC7NIDQX4HgH0u75q3bqGIrMyQ3xaW7mrJhd9MfANbrUKE7gEjbGNgBQSpoeuZ
J4KLjA3RamR2XY5ao9Ggt55WHfZ1KKdFQTQ5ivq+kPFJuQA/VBtNq3ZyF4RUcARZApV30F4M2jxJ
lcGYHxsNSW06pp9BvYz3JZD5XB1xPX97C/vFxEGZvO2C+LXMDFv7BjG1cmbD6Si9klaezonmPGYW
QGAKG3NwqsQbdaxIMq+IqNuKcEFKGu5ArXTqZTiBONbIeUMH60zwmrd8sL5OIaWoXJjwAc+00Z4d
tEZZWY4ohpI7lEIJzoiEpK5mFJuopaNEt+7D59CBe/JpkA+owAi7jVIdXkcqc3fm3WOyEtvS3Vqq
AHeLIID8QPY00pC+249fMvd6qIp4kMNYpBcSKlkhft+tu4URgXbor/KLnMROafynJup7jCFmdjjh
KXOR4lB05v4/BoJGU5d/w5AeuImd7DhHK3cP/JPPJc2XABjjq0HA/ahve2t5iMLkXHww1IDti6wS
OsRgFJ3Yz+LEg6kSeSZBquCX9MlXAM/A6gzbYIRSfP/Fj9fdWSO1cbzPs3IhHjzTD7Blpr2N/80Z
VAFPJ522kh53MX2xrSoev15OXmBQexBupow0zo60rYunaD0wJMMTpqxcOm5Z9jsGJNgugeMk5UyC
s9u5DPiiq3jsgLNMPYMKO4Bu8MtixeSEZay24kKv5A7l5cr/VmgyrTcxH4Uiv5udn1S5LR8tI86X
nmOApaofVcPIFc85KbCEBk1lSk8oL4/c3jJwU+v1VHqK3Kjn+MTOL/eiNAyY+kjY5u5KQh7fytv8
dq5MgsVwe2B3U7KqLLd/0sX3K4Oc5Lqpu1brQnTYUVRFW/jvtnk3HaEHdBmZ1AhjqoX6h36/9Tub
zXktwS7/pDvAHWsKZSXjRRj8JFiDoquk/0PXXUMSacivsJyp/CEAahs4ITPrkXMf2dyGfopTqUKc
a84+lOa0gU2wclCCnof8LqlmtLXqO3wCKOXKQpkKF808TExrsCT9tQIaM/7Pgyz8p07SsPqF8H9w
SOKtYW9ErTZVNMOg2L8VfYVHjCzMS6jEefLDSgl1TLQTdvwyaXfCL/GyidIZq7JsPC+p+T67ZQl/
2AI4ZeEKrvozFZ1RRrXRKNVqVCEx75Sok/fcXd8IudvejtOJQhnGBJMZ2Ucq+RobPVTsR9yljI6C
Ek8I0jhrPiHKr5KOFFKSfV+mqVNC
`protect end_protected
