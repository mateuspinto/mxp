`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CXFLE4opZDij3FJ4kD10g0Dz4fpNcwp++DGK7mEwDLZ2JnpvEDzhflgZ4UxUJGDQny6o2b0Gz6zw
BEuRD4EAaWi0P4BO5Yt9n3RUHx/BU8A6oAs0l5is0YkSbR9wDZDPdW626kF9x6a5eWU4mo9LbqgY
VE3zD45Vd3qO7Ed5LhSiFvRqZ2rOTKQJUam8SlM7NP8JKG4PB3Z+tbT1+7mZPoXBWsiEPmjGfyiK
no5qHLs4L24MeIPDd+pUAu/kcWnQBOJ1hEGWFS3xJrbyjDrWTSZsaUeK+2rNxdjEIW0xYwu6/tJ7
r3U5QfgeNT9fGK/WxW+uoy22dxZIGQ+L43+AIw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="5/Zb+64d1C/PtM/0CNW5UFwDqbHUiZQiLB1IDUu6opo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
x8QKkxg9QNxPBw6kYirur9OcglazrqCc4r4db0IYrizy6OlSKLTKnKPRjFrqoOyVNlD0P6ltWAiH
mLzM8Gc0AnNK1/PhTFoukq+6UxtFxhyAlUMmDI1RzMDqXmmsZX0821UFE/3m/BAQU3TK0rXHPcCS
qGoX7rFX3IQ91j+wGT+nA7NfH9xJd3HOaCGVojRbn4/vyH4NWfs8BnbI7nnimWtSkb0OZ94zSGtY
k15XHfVikleoeivwXKj0zfYpNkNXDOnfoa/lSJBl+7K8/fzwZhlanqrR7UAx0qm7tolxpRawMgSW
XhjsnwJHubJCPJBxBbzDDmUdNUVwe44cyUDpHcbq7n3skVnDBsmQI/CFYGbQneRM2N4AA1UVgrD0
ntjWTBYAmE9otWleWYAUmjXLsQVSsvsNwIfIBEUfGVg8pKyviz3EKyh+Dyf4YbwO7wSmqJQbH0Kc
MOEyElkdAUWx23Xmh9NeTg7pZgh8CT8W3RPXIJpzePEn1qkJbndqrjCWXW2pGIyYKIki+yMxm7cL
VUR7tGOAj/tL96JyMr+Uoan58LgCRAIXt4AP5TbXSbie7XoFy0+KCuikAN+C/0pW8aCUUb7+s7j8
nYlb6jUdGyBMdj/GOpkgjsWwM19eCy6TaqpRmapFfvxSiAXMEhnUIHx939ivfi29dfy8XLkOZ6iO
4kk0ae+VQjoOL6U9J1EbQYbb54mjmKej2lIoW+Zt6Lo69+d44m1sAyJeLnAUpItBNINpMXzAOQ1/
dRtmEyJ7si3U9GtPdaALpKQhHmT8ovrOTnSzkUpavAMkMukqPTY5fe7YyOy4dv4ycWXZt3E5Whhr
s3rqr5OryEGsz7PEBX/UnmaPgHW/AUOfCFH2cuEj0+DIXll3o2Gm8M5ltzRCQwaqhH7GIS4AR0Fm
uHyVG9tD74vcSPuOOANbIzv/rcu/VdyUPlQycYPVu63ecQGCey4eSgM/McqLsxe97QxSQ2pGzMVB
do+LvCSPuFoK0dyz0FKwdcl0KSXWcq5bAscXQsmRDHUCI9Cg65rv0s2w214WPJ50jJOXmtFlOq+p
0eQyTgAav6jUBHyx4+GrGTU4BnXqyZRAGlbO+8GZu5vzvDj+Wn8mYEuCTbkmqg3yWKk8XIL0yobo
nIhWxpG/ARCCku/QiK4CFj/2+tklMaUKSxHmosFbw6K4pY4EsrzUBVnT7bb8ql/ij0rKdovcpFif
0orVezvJPjsPgGcRSbRNsNq6MOg0CMVwmqVCzuhE1EmmFhtJy/6AuMBVjjjyehNgqFu72BznysGS
BgCmp1m8/EmAT+dumuzfT5DKSuMV+CF9KtMjtlOJm+fO0tJJGzOwdCAozfRYGYXzPPosYS5JfCea
6tMbdEoEO2WonljHJMmNEso+nkjaDamc0t9X5E6cFQ8/xk4s0//fBFHH6X1WcoKLMV9MvdehEqru
AJ9Cqhq1jV+BUFCDzFPUGxzY8pDe4kn8O1E0/JTYtw7NwvClaTK/yM/7i/FA8GxoaacV2GlO+3x3
k9pkcQ6m9K3QnDHc2oBZx1YS9p+ATyWM8xXoKA65aXYFI03SXioZ5gU5K3+zrLp5xiECU0LrZrOy
+uBdcnng11tIhUNFqrptWgVphxogyraJNAmRpvMkLaedsl3vVEyaESpRQl4DS6fdiG7uhfneSRKs
As7Nsv4W/Yl9/FLWUSAEvDPNe83et3PYfroBLeNMaVC/SU6Wuh+hf2Vlh7N3gNG3ACpsqwxQDiqE
ntpzHkMqc4paqdOzlCrYO64Rg6IfLWjT0u1Ba2xRhHWe5DvlbiCPxSq2Fwkj5kf2XX4kXPeNgP6l
/a1PdB9rKLUdTXB+qcR5pzT2EKLOw2/NRjV/eFh+4N+pebnEnxxey8clToFVYQ+YDNNdTe7u3mf4
tAJIT7GkctDwLf6vES/WZ0x72CkjRkh2SaEzpcub6RSmjBMnMSL2WWS86JHiDe8ojCCismQfWQ58
qWJlq0RE3zBcmXOV08u0U2TtiI204iRMR9+v0e9BZpbYG9pTuWLWG4lH/4yu8vYWbclUAHBYtT9F
ZxHKkENo2VdMhHhydtnRCQXw8yetivBKK/HYDPMt/t1fGp1Mfd9WsFm0zSjaacEYdJIu/xL3zTtt
twDE6TOH31jYfWAL/fRs50/9w3YHPOk5znF42vxFce3jvRoNxmdDBC4YI6oPHrofOBBBGd4VyLRN
t9L8TT5/dEYnmIXI7AKOVrwQx3zqdUPWbfbQEP+elZQ5RmGVwKgGuJtBc/SQV/aSOZizkgS1S0bl
j51+tv3WENkWtiGVJcwJPi1dep/iCQz+SSZ72iG7dNoFF8jwRytiA3/QNmPDuyi1rtw3fMJOmXDA
YFvBy92MdPYgNLaKoI9tgZB8PNAsr5e6r71A1mIcTIc6KTYkKd+hsjQn9bBZtdBGZ1lmN7MujiaH
vrY8VsBEIq+Dyfx33yBgEpOQ5RHCuRpwERWQWAFGvkMaW42aHvL7jeMQ0Q1+xOUXN/cJ5he6a7uk
gGtIItfathKpYs5PRYGsfdgoNKVOozVWZEqddvk1nSDkGs2Fxi7mbQ93CHrywHorW5ggaJdXzTpQ
kAU9UbbJIeFr6dyNz0K29z6TvpILMWIdC7GFQ+MtfxLkA/Bsi3GpP79QzeQoJA48CGl74IxzbEC4
3P4q4yLXx6tdXZ1N1nqhb1E/MJRZkLlOYCwJ30FJH2KTvaQRGXn/YfgsL3RHti8DVzcjAlJUg9ad
Qps0SX6cmE/dRSXjahcsLhrkqqa4GcARswpzaPGLhUzrxREL76pRQiiDs6PnuDUj9D03WxK/+N5t
52M1uOjO9aY2AoWNLVd2B/tvruCX5hu2j8YInnogkCGs9JqQaeuuUz0oDu+6e64m2nc65gEvN+DG
YhSavSLs6Qp0knsIw6HtGAon2mwfAlhKqQl7fLn7O3G8txZI8+rbbj+UfA7TiHlekJiH6Is3yvxx
48QvUkhsD958U5j6mDMV3tBzkU/bevi0d+CjvNaqh339i5Cv1WQdk75Ym2ThrcJnnclmxTimPz2e
xnlYOxeeZGDEF8GEe30gzKGOu3edE0DoLJLy1GxG7NtCU3MS5eBj1LX5/1o4uZQGnuMiOf8wQgHa
9W6697oR57YqobiG/tkuuNhwzAQXdIJPU2UsDzLEvsnaTxJOiUiSpmpeSk5YXnL3NXDMV9j/gew/
InC97GFZ+rMDBPYnOLngq2IVOQ17fW/8i7fSI3hyQ+tORRKCZTMUi0mMSO6txOmbeUXHGlnwRNdh
DKNuqvoi2nF//9afDc9wvOBFb57FRfehKHtHsUZebtp9kk4M0R2Qx5ViJ9YE9P5gnmsTEzT0b+nL
HJpm9J08MznptKQ9jCxEe+KtFp1uZEIqkDykiYX8uCGSPTi9icbHEcslgc9Lmt4MZy4BwPMaE0ht
qm0bkyLjoqS8mxH7EHKRt9/YwVxEfMjguxpPLA2ZsrJ04hvuMMrJQL5tvYOcXgBj7dn2LhUjAqEq
hXtfDmAYD15YH1wy5JfE35LTjn/ucFx25qXS1uRf+WeXVv975kGxxvZu1tNrTSjxuY3bvZkZICXu
/wcpuYY4H2iYVhnYRPw6ujCgKyKDi/PEcom17uX8lXLNtjI0ZFzi01PCfeR2+woVvoGN00rfXJSn
saH3jihZbP9WW6VDTIif/PY1WmMItbN0bWooW87xPZHh01kri4RlLSFtULJk86ZTkFf4IvMEwmbJ
GaFCSWjqTCzAvgrkTcZQvIAKxgyoC6qcIBEa68Qo5DhLEB/sGO3hSrv8jTJD4tVCCPG7XcIZzW5u
1yjF6AQmhJvWMrYj7EmRhDF2xlAiS4imW3pQ2wyCtmWIdLBqZsXDyWi0cOuanJhAMhlVh5e20m9M
Y+aBQcENf4GRP7ymStNAnzeYtaHwOPGXsv3hrPHkjBmmCFqD65G6faZ/v4uYYUDGcZZq9+jPXdGI
GX+i1DYgfQqdthiXRlxUlwOAt/znLHY7i9KA5dzZjH0fZG8lioEscxiamjTNZDcQgoXGIAYI0sb+
hxmV6497dKgZ+NH7RDmq3aw4Yb/FBCm0mIqbA2NvQi8rNz4wJv+qJU3rUF4g33/E5b3ExpACRchq
sD8MUHtFCN8LF1mqG+Yc+l69LNerL9wVzsbIfZ9dglmll0rKmLYCHkwCS9LugzaRVFYKtiwe2LFr
wWapAVpUYiK8owhlxuELjdryacpIDAz8j7w6gFGXrQClCoaBWgg8fADLdNJrTTesAesUC/r54YnN
cGwoIjJyjQUrolWATP5n7x5sAOs5+vn9eFY+mihQsXrIasCC89AkSYR2NlYEnEpFNJOVYh1UiOt1
DcYh6D5ZJkzA689fwA4Q4JTUZ1HcMRJTyKRQ/waxkhWhwySBJh8vonIRJ86dXfBEC9FMbfU8SwAd
01m2hfrBcUFCJJNCY6J0ka49e7aO1NAe24N73SaFJEHNMOLsfokP7oe2aTK3ArLOT1N5Qd7fI/01
ucoOY8KnlGCgts0/nI9YMDP5586LHlWLj5hvPLY5k/5lgIg74Til2cdSri/dAGbqj8dGvStJ56BU
Yt02BHSmglN95HmH/Fe1jgLCyLRDAMyK05PvLtSA8YunBEw1RYHcNFt3QQyJ9ye3s8Mfs47Xx7co
IQkjoUJFHk0yyKVSXvmh8imswcpLPMxU7lYdXMqcDAV5IfbtssJs5zSUe/j7hQsjRnETT5G2bi/3
6LKilVxzKqxjheCdsTboQOt5naubbiC+fe1Dp/77Ylo9DE07MtMAi3JM4EvH4p6A7+C2SmzjgNvJ
mDqLEwMq1naHk9QIF6t2+62ENA1Cr1PaRfx04nnWp5O3zkaPT7wCTTERouUyVyeBJsx7nKdpbyVU
WtWKW8s39l8uIVV3vCghrjJ2UG4y/wtR6HBgttjtuUC9Ysulf+kmd3mvmaDGQzwc4ynyGbr5Q5jG
AvBzKrtlmXV79DPkqXletJQcYuBDhGIx9ubYhs9c3JEA5It8Y7SC8B6diAbbn6FiBv0hG8g8R13e
FNKv5aCjhaxlFQs+HoGci4H3u+/h7Luc/Qe3oSEcTSb9u5tpD+5s4+SYQvdpdBgpVRc34XqXJMwy
41vAYq97/TUhcFX9P09/TuN1xTzg
`protect end_protected
