`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Yt4PqtdF5ThBw6efxyNy4r9UlpPx/sTkYh0LlMlawPfYP1BE7zE9YYBvm1VknNrxfGKgLJqs8rZl
g8b6WS5reOxxTgDfoGEIudnJbLyCDX8LzoUxp4/XFNxAsWt9fQFAU+q/SuwWKzEcC85Jwdd01QVv
00oRS+LBjhJaxgm4HAoKJ05xRk/ZQckZQ5dHNm8MAgUHhyxBj0YcrvsrsAkKPOfcHUOf4mRD7oPu
mM0RJ+gU3tVdmtnMoZ6de2ZBWau/tIMsTlwguocKjIAFQaHfIA3wez0PzjAxbqA7GGOML7IDAO0L
R3lGh5DY9cWyc2Dx0FppGLMPIDmQyxm60WdUtQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="9drkZT+kpxTCB5L4YDFO9yMOsmpE7ZNcLhr135e8/ME="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13808)
`protect data_block
yCldZuUsHqwzF+ZDwjcu4po5HdV+TFh0O67yGxRvGLn/QUYIpNwuAq1UZfYA2KLcBrulim2jFJKS
wZfVD4ITLG0D9+VYO5WDXdLf/aZGcQkXNMCeDRN2PfHsk6pT2BBH3uBbfBlmDVhKbe5/bmUmwczZ
V18BNuRELdcy87oZ4i111bLzGx7troSNUo7lNi4BocBlNJAmXtqCQ+0XqvLi4RAsBwcrZBSqadU2
ZQhlWORQAw2Gu6IDBZCYff+W65H9vIv/NxU3q60qkeVtfJAXnsAron/ktZXOXgW1yMOCsVx45D0W
oi3pkSP3f6aMLTXXsH0X3OlFqkFoGz+sqR1StDQUJt3LvT0wVdYJNGLHVe7ZZtpW2sEvAh/6HNIX
sXZvDzSfWPy0bFYy+IW0S6qpCRhJO6TFBeDK5NJYTQTNQD9NHBw6WBP3ALdS9Lh5Au+Trnqnh49w
3AZYdzjZ2PiH0MOhakO+8aHgHWMWrVOOsdvw1/A+LqxbDxqjfi8+u9nEmRV+ecVqANAmm34eViT+
TKZ7sNDfwm5lBmB4abkqwD6/Mlvbavty2UTkcJs5ksYrVevsGwn3myIRMH/l26h6irWkO1fWCFWj
kdaH46WGiLA9O/T/NWR/TWMVwjtpdFPYMESECWPmSOsodnik/HnJPWNUalXxU8PegdwTM2WxQiJJ
2GX2pfK51XxQFpOv5sMCoYIM2Uft6trK9kdhNRrVGQa3BgN3sHa+fchH35VarA0JzQroFBVKpegI
Mc299ByX+5P+d273yS0tewk0vI0KI9dq4IrPzqIh6i7NYrSjS9TdErA/blV9MiKQO0yOmdijTPOG
ZW8zDCZ4cjygRie1RpXiBtOZmGmeH5S3BPOO32IC6wLBOYQzYjRrCD68j2dzyD+mOLqsHGTiLWOY
Ei0KnW2hPE/VZQR4YLfNBfwinlz166AwCq2TAWi+fIpQaAsmk9Q8Cy8BZdcgqLv+qCtLDAbKTDY8
IG0yYPyg86kIkA3nUJ7iDfTuk7FEUbdRGYoaUwmrBb/AkRM8A6wYDNWQ6cVWoQaM/3taq/yx/lNQ
kPx9J4oqgjDDzymrO6cwMAGfNVkihvODxv86Nh5VOEQgHWphmQRAMoX2vyq+NsDDUSlMSE9PqDo5
uhRV5JcoIs4CbQD+hBohfaIr/j+CWPefdMpXTEET47Wey64oLyYpPk06sdhGSiRSQR5OkapHOs4W
aEMaJ7HMUjmTth4c6qJ7egcPlf65rFg7cO4NXXBg/+DubY6M1M5egGz0BCZlycEMHuTJsXJZjVId
z+Xbwl0VSee1mAYKgjFF3Dbl8K7VTVmAwGOcq2NEBFZYlM21DQJ54q5FmNFhbjDeyPxUW0Cf6SQK
hcxINF3igeyLBK2VOyBTS3eetd76wfkKreb+P9cfVmnGQbzp+lU8AwKpB8oEzA9qi/j3hIqATd08
ALK7hrv27z8DGTEsXfRjOGh640ILur/01Z+IHCmKi51q0VkrOMJFd3LfThRRcfIODDD7MYgroWP/
5Hxv2yUkAMbs/3hdc/YY+zO47mL6jBPSyCTDxwe3K2ewPnuo0RBecuJ6UHoBhM/Z0VpIXt38Hifu
R+LSrQyiOaBvnELyI+sRWBShAlqWTY1s7Cpabd7ghsbdq85z2Ls+cmpu8GEFDqW+vle4c0UTJqAX
YQ1G4as48xuKk97C8n8dVUGm0ScscMRaqHZbiaqEfSjPSqNV47fSUbPBvzAYBT2Zx/ofDEsmejkN
wLq/4AKEYwy2T3YEBZC+aG+TsqnNBEJfEOYjC8YH028zT/+3tFoxh1k4xWYiObKNIWOr8lohmA5R
mGSrSOmyIy9WhKJPyR2npHGdjPKITlEoyL/luVrvwdmOSAOqW+Rjc5Zfo8MUSoe3otbefBE1NF7Y
Q8K1SvPldYhr/7OSRv1j/cneB7eGALISB4i5DQgKgc/Zvc4h4jqfHwjCo5lZUpHm1LQK4otkS0sn
2dVSa6pPTkucLkrOMMxvWQC9Fu65rQzt07o2tctBEszRkRsaRR1eFl+oW36JZiCQyh97FypYJNFa
kMq1zCOxLXNp2bdqc5aOa1DekmJmGemWfVZFQaeaAyMvPnAB6/pvNCr5xD/clnJ7/ooWjMpRsYu+
wI2fONm/Dz+G6V1YyB8HC5Mqc5TgQ9Xch+wwnq6AIxADlRaV6ad5jdw/oIUzK9DlvdiwavZrzQ5V
az+QhiC0QS0u5mcuHB/RL6tFxnNSo6njstbdfHqTrrf38XUUZ1P5MMK+bl4jKz5apkTr9Xn1dzCS
yEsUueCE6fX8X3cFOAjw5QJkJB+jwf9+XRYbA9hF4z/syVDRM2DjliVPp7yaiYoxsxTWJ8dmDPeI
9Rvn5TtI9qf7zSpk4Ki0m5ZLi/lnJnPMkbr8TNNqVzkKf5LrfCuQeW3tPA/sGbMlgv5W/lClA29i
I/td5vdeoc8P9GCmFFxVY3O6ZGCDdvBEcwY6+w8VPAHsRqtTS46yfyk7HAN2/3HMk/f1cqc4+PXQ
+ZLcHvoLZFxuy59wd6m8ZinOEQ0BKc1VV9GEYLiDcTlRKaX+nSkv2xHMVTLs7eQoDYKtXabfolq5
AaqwjHFxf2qFtGfMwo+aorgm8rPyTz1F43RNFtEm9QPHGbGyDdMgqMTvuJKcXUxlxrZFKZy7kxOy
Yf68cqRvywuF45YFNAegTTPvEKaW0xRncjfUAzDUC0xd+s/bJEiruQzXQ2RJChkxsuIIyq8CWvbn
9Xp3jeXHZ6a9rxi+dNuOiwglyaxVIx0S98yem+R6Rh8CGuJCYRZA+1GWenUw4h6Juf293BBJg2aW
6WgGSuGI4z2doF0jfFACWzHoPJzyNVuKilxpfuW3ScX4o5BOEglF9JW0qYNm/vmW2h9OfZXW5yL3
p4Tof0QOqr3EmaKOX1zvBW9xsMfWWLqkMOPiz67vrvvk2agNZYuOZx3UNsafDySLHzapp/sAWGdt
8m6Us0egcjxqDU1NC4CVmpSCUPJhnsPwnACzOxun1OyIp172qmv/CuikSQjhcp8oFjSBpxCI01hI
R9APpU0HwhqS20zHVkMdrzjdk7MR1mb7bUGmwmxB+jx/i7cQQY7CF0RFQXGEOFEd6jn/MOgde79J
MyZbxPSOmGwcTDTUJ82QhDw9rBmQPk9Z9WwtlCpWerSLDt7hYYHWvcSCKYt3Q+4LsW+tLBTixm2+
t0wHShar/Zbpax4YXvjlJVPN8cW6hXTvwiYiaiHOknjoe+gwotuglC5Oo7KtPa13V03QGr7gr+ks
CDLMYH2c7nByU5k0ftNfGkpzm8lh+UrKJftJtQL7AASgi91i/xitmg1qroNteOKPWiJ10+fSVqMY
FpbEbhSCh6UPdqHNyqc/ChlrmFSFsPJN0cjXQUV80//FV4jarG0dr71S3b82zByRaie6tJyBDHqq
0ExSLehTwc1Fn1LZMe5+2zVUnKZy+cG5TpLuUN2kRy/nzy5IDCgi27Dvzf97zWfui8H/F1oUC2pF
fUXVyBDCqStkU5AYJQZOgd9pGyqbaUK6cUW77Sx6Rr713pZ7Pl31RitfOrzn2qO+xvb+L6uq7njL
EAZteb6vTCXe/xmyw5MG1caHblteFeolGLYYzzpr5vTsz8zkWerzVL7VtIJZ8A33nw066MlCcRiW
OPwjjw/tanlGfmaZvTiM8pyRtKqpEqaFIzZXODnJo83mS4XhKQLE5tPzY8btkP/AZ4pwjvuZ7Htt
CidDQmfydy91hqVkS+Ok5d8aBbw55lkgr30NPafkTGuDJEuPH4ECgCqD/qQFKEBdOzIRFjG3pKjF
tfnWUyvEMPBv8/ET+WDxIiuZ+aNkKgZAJ9RPNjrTyPNKYs6Rb0LPmzHPKnLQ8BlAkb+VP9iZU3+A
sMxED61cy4z70imvl+W27jIYsUF//a63SpdGes7WfjCXZIEmmssuHwdpJq603vvMC9WsL52I8BjP
figOdikLnOmFvuOuUDJk+7hqyWj/mX8sNAKmnbB5NUaod+4Bry+iGMaNSbEUMtx+zMmO5smFlfVu
L3I50J9AjFg+6k5YhgkRGENmAeRnk6e3lP0sNWox03Cnyc6PrP57ES8geoAClgc9hIj6SaZlsb+I
HMUcL7tLfk7Z/fcxImok8sYlaj56/GEZsl3iRUR1YEHWO3tz4ZZ5SMH7Uo6BrY07TwyuBgS6yr8a
UUYjCEZsK8xOuF0FklAocgDIUKR6hei96AK/rbrO7W6slfNrJyGSsE7x+xMkUUfiwHgnZN+gvT/F
yIm+HgvneEVq+9kjNZ+xH6Y5rCzfyTSnXbh8Cf6V48k+0sxvQwBY/hWfVRXjF9ctYGRkJyxe1p0d
qshEtdjIcNTxn/GznfdwwmjDdaq9Kkvk1F4fzVcYY+L1zxmY7byXleukzMzXYOGhlul0WM6q6hYq
FQr3W8uJW87dllCl0rDXmbEHlLRCS6ZjwzQvJz+IHJ0qEvvsVYXdZiWwP6nY4+WFh3tpSt0+Sa4H
D0JnVoGyn6dpn77qYmzoNEa8KgCrAJBj8gMD/RNjuTI3DpaHKY2RIZZxexhTPxsBccBWQG1XsE0N
1H9gOTCF3lhOPSajhCmBiBy//h9kNZTx9C5ikbZXZuUFRB1MVReDhQzETh7KylUVtxs8gvlZ7bcX
mA/Fvzyi9hwJ/Mg8fAFvjsqY6FdKQahXlooYGigK6UTrAGm0wFcfejTfB8b4X8TLy/GGySjam5RX
5xLJKelk03poPltoeNVrUE1ZriF/p2eDEpnqklvkfn6kntskB4xHDFDKoWVeZPXLVYhiVw8hqJjI
bWbsxdEr92/iwCIpz2PpUmzj+S7N3YMpOCp8kIMHgrowLHWE1m/pczgpeqUMmynP8yhTqvY/gg5R
uDp9kdb70q4Aw9uHumE0hriS427olHqKtEpkaGTpv++Tx7gSgvoq/WPM6X95qpm3Mt2Yu5Mov7VS
PN/qFS8NzNWDe7O1b3ReWvZ7xkihXkWx3oEaW2zKci7mYR8x4Jhjy5/4/GOTtLJ/khfU6s+3cqy+
Pbi8p7DxCqlBhIAClpIHIl8Fd8Z0NXrFgG7+9XrmZiIy7I24ZX6N10iqxVAZrUI2bXPhow4ZX8Pp
R3t6IlAES0nDYyvY8iqYRa2H99rMv0IM1Ed4jaYIHrnMkfEKLSM87vtcpSFY2fY3/tGgO9TAebZL
L+VxT0BB7Z+kno2xB394OFpfe7ZAagvk27wGw+dY+mKG7iO+ImAOO+bvaKML7twcbPv/4GqNJQeR
jN3jprypEvaT0DgzjW30rTa0KuxGycnKEvZuAhPGQwy9UWmH4lOSQT3FR3kIGDEfcxF3fKZxC/lJ
v3Y7D8oxkR18WR91B98sBh/xDhq6F3oZ95A+zQAOcYR/wv9rwTYmSaoheWyxyVIP+ImVK0r3ycZ+
C/xOqO2yHLWXtaqG2Jhatx+81lYR8Vp8eDLDNrDyi7jxH9obHnzfn1TGQL8WnWKhIr5P98rSCnyk
OPTyKXWtuDgzQd8vinIIybKkQIMA0dmRBoLqvf7ot8DFhL0K+SIjDfmUOemX9KEgwcQ+PYcvy9Ue
jeBeiHp31zlbHtO+eJfEyiGz9U5lZhHXn4lt6MniiiZK8GK71HvQDaroLH8wd+YPalzRNCPTsZ43
ihbsguwQvxFV7VbrCExcCVBizluTfNd4gDaWNi0tZQryGGIajjGiCJrUHu3WbSZIhegpHXddnqJN
KC3W9ZozWUSrA/2avCbmdSO6awWSNPRKUMbYhRvbdiU/m9HBxm3phDMt6nhL0cTti+txPcjOQtp0
I3SZX+CqGDFF8CvRlG3MPhLg+ZUFckFfgzvX9Vb0nW/r/TpsbqOBZlEurid9QeHSUelKSoUe3JhE
oXBR+JRmFpreTcW5ONgTXUqanHP8P8AwFGpt86wGJnb+fA2ZNmshnv3HyExZAJTn5FW6yTDhi8hc
x7g+vcwtx369TUc0F3q+CcSq4p0EhSyF0aTLH0CQMbwGD6zWB2A9QAQjeaPhVhkupC6cAvS3LLC9
0hAMlbCiOIrB3r6icNK3wjU5tBR6hWnZmkv1IMJl3QjSo1zGwas2idXgKFdzfeEsJf8rUSCqEqIT
pxvpH+JTL1kXJXhMVVPNbYJEdCO76T/Yf8EP8qHn0NoBMpQ1aEdFplyfjbV8XXjNgMOawcpBF+64
0BsOQtUfE69cTS9S7SLV+fT92Ecc10qlLCsFtxzg/0kCn3cqeFJICeioq6t1ErwgLKvonsNR/KWD
iO7y6GNL7+SlDsKEHeaCEeQ0H+2MziRoREO9U+55nD/vbG33RnSN6crWJHytUOORfcKAdRTGyRc8
14aHdNAjaIuyKKCGBDpRMx1wP0C3FP1haWGtzacvF83k/0kBOE0uearMMPaQ0AI//KeOmf5LeEtD
OV0uVaOaAETIaPWzCKXES+hhgTE5pceYc2GrnkncvhLxWISVPuvuF6YxpRjPMZ1xMjK4a35grfM2
a+B87hvLbjj1ait+kIuT+li1BdAlVPvlJHJWpA/zQUsgWjFYBcHHaquUH0NWKB6fDGOz/eQfdAS5
SpQEuAy6279jR/x3r2zQ0OGNgL5Uwa2YYNHByFNVXHhD1WuFRWOyi/JldV3MDiEbwph8Q7WzPcf1
rFsxrZQHeS2P5gH2T9rmxtZptMIv3rrNN/ut+nOjR1/0bO96zf8SJYVyCMa+uD5Mff+C6JiY4K9O
H7fPKgxIvljBkTHxaUf6l84QFwxRl6i89Bo7iEF4dFznoEZcF/IKyNvUXHHHx+fsfZRkHHja1ebJ
gqtQGseixSNuBgkJemytDua95Zdv4BWyODTCMR1U4cHFfMJmAptnYnnEKfXDzX5wIOT59ST33VW2
A3D/g2WxnP66gOCYVCIKHLJVUjTdlJoCSMwQ5i5SYQmHI4pxYJxJ/ig8a2UGlT8UsYGTqYYB9zAR
zAKuDjqLPNJaQkSguJE+QB/0syFTg9+LSKKCq+RZ10sPFRHTpAaSGkViftm42DmRuD14Y/XbNJ01
YpYrP/FUg35HvrY69fURBvTToWnRKA++8yDf5O1zrF+jqu2LEpp4XYWlGvfENeQQz1WNjPJrZJcV
m49lSyI8/vPkyVjCc0/s7eGFEeTCW4Xno9091L6cFIqluJ/h/LJhQJBIkrTb3ucrw7fHddJragD9
1oi5kHGZZNb+xRZQHdwJkL2JfLbRNKRXMCSze1mgv7un8YDN03OYuMceAVBJ9nWMgeuNjri2i9oa
Ze/YgxQRgvr582H0Xj26z2dSs5HosShVA0RmqfhFxNd7pPNn1tlwTYDJUa1HEhBBeN9Dt0KnyvFw
AHbYcL3DFu+hBwO9ad5dIr2iBuAt8vpkClv92cM6Cw+/iMCMk/Q4cBP2ESVoKI/4j6Xrg/pzfccq
ltuEXUMDNrh/AXigrCoS/yFvOfHGAxGZNv76+jj5GQY7sdEIjfwOyiWUAJ5OP9vmqQihgYpTdI7n
xKR5aodtYQh458W6h8othSiXR+0IheC4DtEWvi6OhUV66YfbYmHLSGP5ViuhzwJffrMZXTkrcLrE
VJfqlc2qeoCnTddOFblwCWbfLQ5/SydCA7enBME5hWuPE8fnnTTsF4NAAFr5lkJT2JgyJHSUngkI
lymm9mTI47UJSSbBjxPzzPgpAmmwpoduXMOjWuCVjFNT2ePyWpU/ehOlbTTnls+1fUPosdYsuikJ
wDqvb2uCtQhkQC8LCfttJeYZbMkOIc9cAV4OCjMVIdJUWDlaXg/67FLhv1u+9wNlJvqjVVtjpkwW
PFKyhELJPqti+kiE2NGIWQE8CrK3qxFKm2BEtpieyArDd8aZzBn4ZSRBY9SOFaR1IkyxtswmPee9
m7Kfn/brfnlTr34KC7CkXgEDhdmiHiof0AGsc8VAT54slEUt+oSvzWXxVGxDO5PXXP6FFm0T8mMY
oiXHZqfa3dXlyHIDCNH2FDr5oO4V1ZQKOdIK89lzNzTVU4+Yb5Y0h84xLg146Qx4zzYFBbZ19Far
VeWNy3k52yY0aZEIkSaM5yDkYZi+7AM64mNGUHKZjWmRO3W8afMpvb5BKbOkbnBe9ATVZPo6lYtY
6MCWvJQGlrAIqLTNAuIcrEJhd0cMlpeE4PX/cVWGXwR/xuoT0G3INT7q2AEJWquntNOnFGdcsVEM
gn9r/Idz3QZ6MVwnv90lYiNOr53cMBDcnisZNg5u8v93bYOgMVzk4PBan0pQUS2sEkj496iByGqk
hq24arZj/OdDEAdsBp7AkFEo6opTTLjt0fCGqBHF1gpOhObj0CVqVzBGigX0a2b4SxlPJEtomljt
7EjnJ5vrTiNQYYWRsYzkwQlSgp82lVTQcuePMmRyv+5E+mQEd+QLRQR3ECWTBpew7F+0aXwXB8zr
vFGJZDIqeltXpkibmKC5/H6R86eJU7FKVcpjPrMuK9p5IsS3dNjKFJqNmgoXcx9aY1q37n08p7bf
InGaqkS/LPez9nODUitsuZHr5D56ROxGu0swz3Mf868i89ABvsAgyUNB+LrmZsH6mYrIKjFjFQq6
FhDA8b1CUnXCpA/UvizrtQjA1CN6Djyvlw1s2KWoo5ze3mArAIef+3s6YwHhKHtuAFLe+YP86pCS
DbdzSDFUqhb3rZ0QFsde07r9OWwef+u4b7J3bcpDyMy9wslm8yMVrjE1rIPuP60waaBNfppHLOPD
03kqtAfgoYtS4J8ar/0F17aRNPqH3zP0BniBy53aHNnVJsgOOuyvdIkScLXQpNtu/9U4HM1g3t2A
boDJkgGjLyoYNVXKK/Qz1zDEZF7ufTIxL9uqBXiuFhBx7PB3yIzoTzvdCYpXD9hp324bS2I/e7st
cHeIWRIO/+luRqhcNqTnbuCGeGNqDWAk0/tPhH/Rvk/Wdhxr9sZ6Th8EDFsYGKOxFvUZYcbOzPyL
BCkBfcLfwvYnelCNTF6gfWk6vAy1/6GaRZBLgIZqk+DEosq5mHevi9+ArlLRe9rZvdQupQRcLw0+
CxIDc1mlkrZEurMbLL4IaadvECv9mDYFofH20uFyZedhT14/vHUIFNOJFaaxcJuATdXIRjI1gb/Z
kwUEG5iQhwhdnveJi6Vqqy64nHG2yQuin14zyzYHphGfmF5Zq0e0Z/NKZvI0hkIYMmxqF40IGMa6
uL9uYReyxRRZ5TI1LdMDvj0Yb3WcHKkdZnEfh/PvVGMn/LEVNbLN1iEuiO/65uJPIiZn2O4Y+9pV
g+Ni0xAoXDf90BR7OxmHpN1AUhBp3l00qSLiN2i+lH5xhUjjAOwr1cbsCAn3nmdeiH5aTCqYCrwC
OT4U7zzSCWqHyxXuYnQEV9yx9Fplu52E/tWsv0VSr7YZR7T1fI91yYCk2rwjKGquNCS6s3srvOdG
iCbmWPfEhMBGJF4QKWWyUtKOlFkVYFQFSic8ZjEvKULJP854Ofhjycvr9jRFkX7ct+RSog/fDQTL
C25T9a0cvX8Pxh9KfTxnsk6oZYJibaLEyP3sEJ0cb9JSgE+Fys5XVdA4Oa6sFYer2Jvzc/fc9iV5
WR8c2BvK80GTVS/13s9kQDoY/KcE8HUsfjx9YQSwHpP1RFRDxCpVM/YfSDqJUaL+lFNOoMsNnXvw
86kpV6tHLjAqf162dCTVLOtZHMIOfLsAWg9f6Tr1ahIxB9W8qy09AlJHx0UjMO1+oHd3mmu1/NvZ
jBW82QfdhAGQsH4ZMyeOjJ+Q/0r5yEtl1CebxOCuU+w8ioP8rRnXypd6osOextzAjUQFNbNi2IeU
UtdkLMLgUFYK3L9hV20EAxaAADzGDhsa/BKZMCHo+j3jZBdH0uCTjmQGE/UsRZinrz9LH04emdCV
9JhBupcgR+9Lq20irANiFclXjZYhP/V+aNVJ2l3sblGLt9E45JyQxTaEj+Uy4dEy6QcpLK/IF9QP
19LyUOekfFlgn00Yo+IMlQ1iRcvW2euUWVAED8x75+X9LSzxsEC46nJbN32Z+EQuNeaZQi0XG8NS
ZFVK0KScm2ekU7hv53C0vScCaUdt4QNvZwVTPpEG3Zo2hGRkfv/KCOYpbYZuAXTf41uzxmYl9m2B
bkDzpLbQkxRUJ52R6yPxxTcgOdxt5qHBsTi/b8PldZ1IRydfly1VSkFlvEha38nOt4PdmHHlqKQT
b4BZ53r+f5tq9XRnOIY8uHVeGC/iK3J2XEowVi7C9jSe+rCqRJRw9cU3SpCem02p/khkZUvIm4fX
wuSa/PSpKOzolpzXMPCm/4qIw62grRybIfivSc7qOgnm/YcjmdWqgS1a8EndiaSfEz0wWQLktE7X
RlLkPIaX33tJcWWIl+bih4pAH4JqZjgD++6acUzwD8FAXhL9GG6bQOEyx7hZ92qHBA0hXmwmQXoy
MZXI12/DLyY4j0ShsGKHxahjCgc5MFIV+yamiG0F/mran68FG+XRwGdDJUACrUBq78VJ2KKburiR
S8t1i9QPTKKynfvVcs0HgHEFoRvi1/fpRTBa390cmy6KetKR7HivxqEr12PrwP0MIQ3Pp/KdW/i3
4DnMm4xaAqbCjIe+Y7ZG6V5r/hazZ5vBVMnmKKslPzjJ6wMB7V/mXRc2fk4pgYuP0Yh87bHTM8e3
AtzpkoVxDbN1PEc8V0TupUrOpOB0sEUu/9CGCHRaKPf4uFaNF2/su1bQ02Exsu3/z1fvmJWI0Vix
hS1oajIL19pJmQI7SwkmSfnqGIfYlDWa7kP8cwfiZ/KmvKcCASlT6b9JyMufLPyFuA8qvLS8dCAu
nKspM/G+yx7s/6kHddTEM+njeRZlEKnd26/A/pmzSIL/glDB+2Ubpr11Q2pY3ytW2GNRpMH8mYop
U4ev+sR0c5PZ/08CC507xj7dDbiMMzxcNXAakBF7nkaOocudfsWutFSIEzCcQaj1EWa4MYWet0p1
gNtkoNOZne5NQTLfnPeaubBpj3mQiCqGZqLQadgyrpC/8QRTxgb02TKGlkfkBCO970mViD5G8nC4
tCLWXoc4TpN2P8eGETRslsUaX2olNPaeGdwuj6kSQbem1KgxjNSDOztkTA8K6Sh0SXkDJPd2qkXy
gUzEr1WYDqplJaECXCUwocAPbEFxlUTl79Hl/E2fSneCuGKrqiP2Z4NZm/2aICfItvIOdkbCg4s0
fGng9Nlo42/x3sc4h8A2+tqYm182wTnQgdNF3x/15rbwXhhS7DwGz2l2+jAP0EpDiwzTQ1tQa2Mx
rpMv0avMkI5Qhv9qeaPxGLdByxW80da9MejDX7K31XO3W5RZ1y+wZAWfyBVSBwCiHDRpaemacmeI
NvJmFgsHHZmq6CcHvXsbdU7zwNi6JknvkG+HUQNjTfxke7jTtPjgR5wcUN3cZlwfbCePGZQgN+8N
V+Ltb50VinRWHth+07rdOaRGo4sPCScBjR4eI91hdwERo2mMIy4DHK7l8PEbGibdXGoFYgCgvhbV
3OLYQ2WD2TmABIV76YaCmwbEaV0SGfrT6okTeX9Ryys1eTaE8GOvPvtys9EgHVZ1IZ3UfE4LFjl9
2hzc+b/DfzvXrEItnqatCpFberK3yKYp+IB+br6Wuf2mi4j7sNIvcBbZy4rm5bempsIrJbHWuUIN
xQUY6ZrBxgKtTt01xR2O0wZoF6hFnP1QsTquWxBFMWp5MGF66+qUWCd/IPF7bdnumL2Xo1+IDNKB
ZLGpxHucUWCtlLZaNA6MZJ7MJy8lwvmP6N2QekzBwW1yELdpxRMPQFvvyUTKMAhy71rHBCnC0TG9
a2B30RIYi/lv323sk+RG8D9L3s8CtG6SudduiHPJjm33QJwZBUCLNqmsjVDropNueh9vVnYi6O6D
OoTL6OhBZDw13KhSf7/nshLxd2mgiYx1OZ8f0m2jfIiabHKqnYZngRShURU8c0qR7c/zRakIn5Nt
Q2CGyRvCimwSfVPgFzvunpScnUkLReZLgqGD9eCJWDk6UB7Lle2rkZ/N+xVny3DvMWNuKZ3YmrGR
wpJFrnsyjRVYY9VcrUX2v3rZ0wi6gk+ASxa9M3bID9oWKVkoGVTE0jW4marJ4dogerHdQrtaVGaQ
CMEoAJXFIvsZ8vXOIxeej1lm58DITTmO7Gamu0CAtlp3KJ7PDzvPdIfBK7ufGEd+213eEI37ueEl
4hWNASSBfTAL9e39ZEfjd2PLyA39KQXtVsMs8Bv3lNJL+AU1Di5qbegCUpfCsmsVsvAp06r3cu37
LNzUXAGOL9v2cskYpKsOXVdxYYXgRJZ41UxNToGVJyJC/7OIWWc8Fps5v+0J75ZguU/m9kI3bUJo
SY/lmEoblKq57zFFQAc+O3IYKwTHffaDpHTmfoNZTJbAXCCgtMfyL0ggcCxnrFLObiM2f86OU8FU
hIj15BuBGKfGQdIoaaXBO1aCllcHVd2sOXa42zo+WUDpvGNwfqR7l3+7/lNqSJnvS167xwq/Apru
w4HaPYaTqRAXfWGMA3iwsnprvrMU1YLNE1xwxO7ksOJOpPE/BG3Lkzq2ksfTH329FSUoPqY7fZlD
lvwI6cS/3y9y8MkpE8+kCxhleTnKIO87qeVXdU8XickLQmK+B7oHpq1PsKbCM4zBWMMKD3gxaENi
b0UZPai0DsixIpkYH5MN5czsJlYn47kaY/e1l3uPImF4yVw+urRgtkwNPWcMhqi+PBBv5JdrdEhM
SunOtCIAC5ftm34/AS6maeDLHlK07icupEvNChFMAgLuADKkJ2Vepn146QsU4epI2hvmMYTD7pa7
2a81raX4S/gP+q0OwlgPSvF6VMc5iqbOIccl+OZyTwIYuPCnlgIv8KsQAnGMp99oVR9y5UzBFhay
lz5UcCtmVEhLJ1l9mDMyrJwioFrOGcTxYEIPjxWdW/a5aIJ3JNqEGe51iKPlkhQj0ejIJ5pYstEY
0TMSUahITiFJ267+NgyvEj/S/c7ITAjThlTGi9F+YFh/shdWDPwG2isaRAYg6OHGa0l8Ydq/QYqP
ROb9HRsz5TF/BJfC13U6gE+/9s8yyIfo1skYV2Fc2vYXS1q8T4F8iD8+Gr+bxDmSHgTGoMHVIHTB
li6Ji1fAkL9GDd8/rf6IG4CWeHZ24A6WF03bobL01GUGrpB3RuL6clmB1/OByNINJq0MkyvF75gO
A6WsEDNrMWtaXD678puH3LWlyTuZeM3Z2K9nheLkbK/mC0Sxg+qXtYu9tc0lRYqSDXtXn+hmW5as
UakPUpOibCRNXrDtMbw7CPBrZiv1DY5tSrkpBBwaE0PIFAG6Tv0vqRWTe04BL1E8pTirw+HxJEq4
K4kbU5MFDPj7As5VsYj+5Pa99IIIE9vWetay04F/uHrUoaw4ISZPqWQETdWvw1L1jNqT8wnIBcrY
JhqALRGVfSlu6uo7Fo7RDtiTsP36RYmI8CgnirXX2v4JTdBhaksFQ70Huqh6ivx+MO8xb7QIY5Yi
uj6PUqPQKBZi2ujaH1AvWRT7XKFYgLWRyvVTxzuq3dBK2zR39G5KRbp3oQVvmN4U1BIr3Ha3LFRI
vD62rQhkJcvvqFEkeBiPmIGOdbBl04kuXUzSI5QIuUzJF+s1JpUWRBTY2zEklwp7V9FWseNummVz
R6bAGnJa6LMThOtyJ9t5yr78LR6CHUXkNB9FXnxjftNcE5QTgUDjkvrBevjMRLWdL0oDesX76FsT
pa5DOCwddhNlta0PINhFZOHUB46rV+Ro7g4mzvnFjTDZDGn5XlN7BD23WFbolYWCtV0KWUwCTaBY
SmOapgQtrF/LTv5Xjwtwun9yW38R4g/RUmp6bTrINqmks5aG7jf2uPCN7NsdRKRa/AAs0vGzkpVD
o5vh80e31Ppyl9EOA133/ozR5mupkrKMxGW31odUK6S/9zy5aSGQqds0dyG8nfpNiWaGmCniOk+N
nK65/gUdr880pUxdx4Pk8lPvz57xLQdWf82wWvahiiuPAPjR8Vrs4BP+yBWnMr3mrEY4doRj46GB
7JLMDhX6HQqf1Ifb3BTOncs65UfoSWDhEGAQctSMR2s4casevWQuyztWzGZyasok6eaA+hr5YiSc
M4ZPLZRb5khl7ox+EmJjp239O99Wmgyo5QMzSzReaoHXxfa4P7DbZ16Sgg0iCRaDrKBusV9MOoHR
pxxyrDpRVlHffUb+DTkiDPRemMCJOAwKctPfuqQMorFZ8Ejgw5wafZGmb83ogaZoC2kTb/XdEJSi
3zmqQ+dLSrlHpJ8EGPvFSWais9yasOmoQW7cppxwHwA0UNic2d1/Xi7vXk9TzEu7YaUgP6A9e0u6
NtoiIB8lBCufiQJuJ53jLtaHtjQJB0kDbuTTHjT1mvmHkbn7oeuMT3Ge5nLyCroaFMtroHNBOJ2d
VqYcm9N44HVsD2hwpXsjtDTDM4dJU3ZYj4bw0JReCyLwa3du3297To4xkwP10uSfuJDdPrsZVsHp
1AM3IaWnKkcbXEzhZnhb82lIjvlCpcozXT6nBSkrJslWdgU/TKb/lNpYhw6us/daIDWJqmQJUoKj
vElmEh/E+Gu6hB41nh82tDICoSpe0hCeXR4A9cVRI9PLDofXE7iZRscWlh0wGrFHQubHBb0akLgx
evZgllXwy3eQiSdC599L6Z8dBgfkDSO7Tx0NyNy60SfxNU/QIcyS2Sh6wVsrQzNDpvDyRDxxo0OZ
oNtJGHZpKa+uXTTlDqKiMqBx8YJ3XgsSAoW+Q3n9CoQyc5ifnZ5Z1bm3dql91Szd0AUlywaJH6UR
Vm5c5mWjpZ06TycOV2P5P+nBie+lP6NZAC3xt9CL8on257UgvSyo5lUs+oH63xqoZ/ygSpiEMu1f
hqc3jdth2ro7JZOLsW/KxVCs3IGxNDw0TujL8GbgQxXyo2m/Kb50hN9PUakCaPhglzXTUNuNG/0A
3DjzDZmIq2yErSOxRHbSed4NAUr5oJIzSOhNktSL0DpF8YaGrPnQHULpfsUBS7v7nlqYA4Mv6n4V
hwPPj0nYPYN2KXg7xxN+ijFHiB8zgYrIMQT3fmphzyw76arDHXAbP/EwJe0PzGTaJlSYW2nohSIy
4xSl2Ovg+mog+u8xc53s1MW5qTwOicNzr9U0gxO37VzpbgL1+VA4gjL54DT+26Gu8u33IrpuPHVr
6ULyFOhQskaMsf7gFiSzPcXb/aZwjCLrRVxM6kjYQrr1a8Vepv0onTWavekAlxznjXtp6FUrC28w
qNS687gEIU/5ccKDvKWdg8vpo1agwtPIL/FT45wMtt7mWUKZK/Bt5SOVMDEgu8jzTLlRd9z/jAYV
foDW0j5IGp6IKp5PFLGYB1ObtrsdIZP3gh/jKDySLiq8Ln2JicwUxQqDX6Imaf5lHlVILES5Rq+P
W7E4Tok1l8L5kcCWgnylYD675oJOeuxo6EX4Nz7qC6MpGU0SQj2bSzgjFTB9+kSvaElX+7QO4Oc0
0KOJtgwH2xLpI5lQjxy20Hzkol/BA6xU1HLdFTSUJBQfbVhO8nwQLPahwUUb1N0CH319lg/y7Q4k
EnM66sFkXJxu+rcs6d21eTFC3+8GNuqNUsBfCsKKiE7j7Uu2v1ayJh7usvLx1Ll79KRsjtJoAOoU
vZGE0SiWSrRMUsFet3YVhntyKriOaR9jPa1pcErOTUKUlQa3gUImOOo0RnBoVvsJu3DOnb0YSN0d
QwkBDMbiD2FbN8hyUc6Ku/y1IvAZbWyC6ZeNchw1IFW60iZtLFRMDwFA2ikR8QWIDBpCd/w0Mf3o
vVhfrErfCXS5hwUV+LG29hJeusAniGNBkvyWu9m7x2u8j5SlkajEtG8Gn3phRFp2cN+GSZe+CVFS
NSORwQw6Qf4iACj22dXtEpG/UyZnt7U/7gDYEjLUB6Gbpt5WWQ17Ar4qOFcoc+XE8maPiWkqlWPK
4cDKR8fU7TCUHQN4zVKMpxYn9bVoHV9fQ0lAOFCIRcMJ2n53G4Mq5rgx16b/8EzN63aA83RHT5kC
ydI6P950Rze+kwZz+sbGtx+wqbDuqU5hGaviktNnz3UqH893dQ2+fJDbDuWSsSMOS5G6Pg+kPBU4
kx+uHAO9MPPkIPPfFv2CY+WqwCOQEFBdvzSNG1/ziitdsOgc8HmMGa4a1OACUy8WAHLDzCmRONG5
pg7pWZj3e13LgH8V2Mi54rLYKHXUvG+/vrJTYzpITYLh4YmFg5IathYLnNgrUZpvEoswsoow9Kor
jFEE0eKma4ARdweCUqP5dRdgdI+52GFF1Gzo/3Mlt2VyPxvtJ6t8wJX1UMnLy+k8fM7ag5eAwz+6
OfVWhxKAN6aOHZy/Rez/ZBtKZbfGaoiF02mtMRMl240g+Ywq3OH603VJbyhf+xYK5gM47C1859WM
MDb6w8lcbk0FkmTB5+K+vZFjdeMrE2EMoroRSveieUWAPFBidALrHsACxJquNDwIaAs8wYl+DcDe
2BdxNmRJOc2sFrZZLLD1jEUdY/4dZAxLr/Ukg6vYFSNyymT8tJdbLbp/m4RQGPnowZuSgLzz26Lo
oxg6EW/Tj1YJL5VNXUkXr5eJofbOkns6OhmheI0VENe8TOVHWiOzWhPg8/a3as24oGWCzI0MD4zF
YCc5ljrR3MLy6dEut/k51CGWUqNxzHM34KMyHUf4dLSmm2SmekVJJYGkXUluwxCwffqXZnaZeQxq
dAbr3etIExNSp7nKWTABRoorsfAyQXytYel9hj+xxsRd3CdS/RGAC/2QiTA0DOnzRwi0t5ofcMTe
2CG6jyRAT6Y5HqUo8JU4Qiwc988RJmqeC5l5j+vSF/1OFMsxAS+OQ2TIhk25nzaRML408IZ9wC5f
x0tA8dFtKw7EO/r4dIDDbs2bti3BWo6RPqDIwV2uKs446q6RfRHwitqEOcKkF/Vqhlqs1gq/4eZt
tFjJuxzscgn72deSDR7qujmKsb/oJiVbjNXg9QPEvsiCM0UMoWQV48ODpUJQoRWANduxVwQ3/99Q
A5K7+EceHUEssnmKLGn/38iMYsN92GvXO9EW5MW8BaqT8QUrdbdLDN9GgqlNlaFRkPSkDSlsM1VO
i6ze7/KH03kuplu6XzGywC3ANTjFu7Eaq2jL0wzpcxda0OaMwcI0kcpKtA4zKoCEHtKw80Frr9Gw
lrbIh1PrPXn1mbsNACL9ZQg/97kZizlSVLQibRfdfcSc8rHryHFepzNi/z2exVhm/onjMBFno8RZ
m1SnC4VRFPxsbUMzOEzAFd/Dkmg19y9D2M9lqZ1P6yTVWnHaarIQjMsneOBeqr4/lOSpIhZQS2O5
MfqK0wZCrHf7wBlzb3bDZEWXwM1yS+pHg7wYdKdRi2FpVZLb1RWx401hpqKhzhX9nqMA6w04iPJS
P7E+gtwyca/nCKhDXATU1ph+MWQnSqj8ZRu+UmnS25gu1VPzvUGkGS0KeHwsVwHoR4ttRgIG9b1h
EVonJkA2MVMKSMgWN2Gx79A2PHG5yeI0CnUvEWH5zYZw+3Z+SLfJDOvHxya19hlxZ/SOBVdOKl+Q
Sk103ErpzMj20LhlJ1G8PskvZnGcu96/8Hv+UxYvb+8yFey288cuI8/20pTP7fDHvvPHaFCtOShv
m59MsiN3bqXOVnJSM2hB7kyuiR/CMT54oFSe5Vs6x5bQUwJ3LVemwQ1ulJtIvZC2zZ8erhT2FCZr
wtp3wFu4JFCQ/y7ogrJ+uB1sfpMjcxIrVmkVsFSXORZ2aiDGMJoe/EVHUT0iU3o9hGAxLsidKxBq
0LKMlOweBu2pj6ujMJJS+PTbaa4Zp6Hiu7gAMQFvd9l0RTJaI0HaJ6ici1TTtA8ZMXAtMyc9Kl6P
qn4N+iwhUJNVUPveTYuSKXIyZ+PB6E6XLy0Tzu2I8HrvglkapIhjAwOR84+O7rqNqp7B+5s9atLJ
fTXrtOf4VsRc0FUS9eVlfjz1nRdQbe6T3vK+XHz0KgrFNGyBmGrwkkTn6ZFCZAGdmUzZgV5DPZgB
1uvBcT7YDrl9Y5r2b85AT12FjpwTkUvJD8ybNjHxc5GBVmwLy1O8a/JAhNAfFhj05bXGxDaZcq2Z
CNXSyiPRuFhhnkLDSridyLCzi8/EhXdnmaZ+7YWBx9OXNAOHnUmh/oduCJUJV2pul3OE2PQCe6rY
vrXswTiEeohMXYbvppEnD6iLiaMvRxUmQghuuwNg+EDNia5x/pkTnkccUVMSvzbEahhF5gHcueqU
BBDnVtQSO2Oy8emxh8bFuwRRo7mhs697e+HI6ThSq8+HLsXZ0yQ5eoLawmVV55axN3QuCyDRLYiW
RcWu9dn8cps+URzR06M/63VAw8/TaeyjcQpEcP+DuVZbi3tVDFFutyyE/XXYR+gEfsj7FGio3An6
49wiJ7ByO3wBgc7xetIyiqTuUSHZ+vs4My8nNzC9KAW1cp8VezTrD2LmF7DiaQy59zyt38/+QPtS
GWT3kmnTcPiz6BCKbD/cxudgwW885N8OfUWyIlZGGTistyl5wG4LL8Qmy+9qOyHo1ihi/DmU7yYg
N2bb+Ek542nmCEkTsCk=
`protect end_protected
