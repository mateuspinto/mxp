��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����&C�o����@X�;��}�)Vųp�mb]4�3�^f�LXAJ@�!�Xh�����\���	HVVE�9�XָP��`��`����{]�3-]R�K�����7-�vI��b|�l�mm#ۘ��
���y�}[Z��G@��XxxŒT)G�B���3Ͽ�=��;���f�e�̬���3�i'y>	0�!2��@p�BN���Um���<;is�X����R(���K�;2�.�����jx����
��nOPhX�����a��Gv��T�<z'����Vk�p}_�������yR��ZkP)������o���x�CD��%<��8n �u[K�?4���%��!�9B����2`(���|{��qs���	�-�P�����t��v]�4Lmҧ-��.�֤������0�"t�9"+�>�V�n{���̝�����tV���E�I�AчN�VQ���d�xo��Ȉh~n�`?��M;3?���[E�)��}2��fjMW�ɩ�������j�_��p>�ӊ�N�yMu���w��b}�$'��pW��|�.��i$�ZC4E�-o�������y"���{~�q��%t��K�"� �o�	��h���E���o"���ث�d!�0��%��<�qs��W/R�+Q���me;v�6U��og������K�(�o��,$�����[���0���A&��Wl�9d-���ϐ�WU�c�Ժ��8SQX��D���$
���94���.���K �	��N݃��gP��ô���X�y�	/�!���M�l�x�vL�Y#֪8���&`^`
�E�Ue��>�����E��&����<��aދ�>7�zk�n��������c��n��u�r$6�s�D�[h�P� �UX�(��v�Pm��}�]C8T[a
Q,a��|�h$�	>�s�s��KSZS4$����Ih﷯�������V�ʴ� �`%Ll~�7j����7(�B��?�)���@B��c��t�'x����m��=_9B��gTn1P��:'u>���n�A�MLr^*�o��l�أ6+tH606L���Y�]؀��S�5c2�&�Z��Vi̳�K�h;�>�������F�d�AS��y���&�P+Y�U*��9���GG_�0�P����6z~�#���z��НZ���*
���7����A�?g�V*�����%�Y�ݣ�H-v�c������2;?c���`�!a|�O��6�Q���e� !X��<2���增ɖ�Q�ٌ8�C6�)��"�_Es�s��DT� �J$*t��l��(��T���l�%IF;���5<l赝���|Up�4�-$����#�G�x���Ǚ�^��@�I�^=����i�? �)fޘ�͏V�y���EG��/�g�/��c���'C����h����IgܳZ[>��������X�u����3������P���f��fR�H�\0��"��9e(�j���R���a8�`����0���L�`�'���������J؂R(%c�_���zDͬ;V�f�`