XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R��Ip�����/P�q�C? ���3�+�cN��u�HV�O��u���s?�{vڬ1�Uۥ
乣/����"��� 4qF݆c#ն*\�QVw]�Yk��������t�!g	��OZ�Ԍe1�6v�=��f[�������y.�G̷+Z�����	��cĹ�̦F����Tޮ�1���"����;mN�,���׽Ζ��ץn{;Qf�J�0��� #T������JK�d�*N���p����>�^�*��?���t��Pd�a�xI��,c�T��<I��k��)����n!|�o�끼A�|A�;��yl��0�?;Ṍ�կ|���+���ݱ�+���b7�{R��r�Xq�%��"�����30�"�y���g,�j ��_p�ئ4�gpZ��_��<.?�4��y=fK���/��'�v!��
JY�U͇7|5�l��"qůCC��������z�7��s��-H
��Y�\�V�J"-[�N�\Rp�7��λE��
���$��XTY.TM �WƊj�P6���xi�н��<~��y�\�MS}aJ��_��A���Fw[^.����$Q�:a)�F�����]rS�.����F6�'1���Ǟu����&!LE�M
'qڼ�~̔3
?`^�I!y,!~!+��J��]^V��L��o�6
2Ay)��9���x�) �ru�^��Sqb�L1 C��B�V���>�aJ���HL�eV�NUZ�k �,��������&)�A��6�
``F[�TXlxVHYEB     400     1b0�J(�����%�G#%�8U�n�����I�H���)x���N���C[����t��og�U���m:�o��ȳ���� �`Z�1����n
YW����4\A2��׵��Mt�s���S�C�1Q��|Þ
P�<W��u���-P[0_��A�[1�G��
B�������L�Sr�v����om�<f5��_����F�w�#��Ü�qOWDЇ�$A�l� P%���~ �����!���S�fq`e�q�_t<���?���������Zx*�_"���9�,�m���e����,{���ˊh�d���6���?� .s/�}�ӵ<�X`�/��5�90��P�*m�W�oQQ;��7�Ct���M�+TᲷ�^D7&�}
�j�p�S}��-�.r���L�Lz�����K�5�ߘ����Pf@XlxVHYEB     400     160�2����	��mH(w�Å	��V!��a�݅E��X�5`<���+'֭�D�
sC�*p�	��g���[Ux��]Ŕ>�����M�,�#�@�~&�K�;�:�Ϻ�2\�%�2>���Gh�c�9x��*I��մ���ngT�N]s���Zbw~�@A0�|����6S����Șǎ�-�O�bO��3̯��w8��8t#�>��qz��J7�a�(��)�#Ji|��^�;n�ʡ�fI��,�m�JuBn4���{:0���ybC��t
n��.�K��m�9��pp�n��
�Io�b��;��^�BHK��� ����,H��\4�Wb�!��Z�V`��&�\��S��dujsf%1XlxVHYEB     400     110��d1��ϔ��a�ڒG���� �}���Ik<d�X���<$
�|�ߗ ���
c������U� )�;ȇ�� L�J�sǘ��E#<T7S#i�w[%܊��[��	���j���ػ	5]�xɩI{�ً�KIc7+��hG��T}�I�zA|n�mad�e�ܒ"芑U���3f[q$�����"��l� }�z��N$(��_�#��a7��A���E_\��n�r@��'y~pu׃����7�׃�-���5��?XlxVHYEB      42      50ې�}$fr����;��B��� ��4�ыH�!i�Vg�-8";�*#x���L�� ��[C>{���,���s w�O�p�%�5��