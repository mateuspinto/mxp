XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����sG�t;M�2g��N���K��\�t��g�?=@�؋Ոʛ�A��Ҕ���!d�i/C^�1S���Ki	G��OR�"02�{��j�H�l��@,?��Y8 È���&��7�̌K�.A����'9����ۧh�<k���Tc<������lU� #��}	Zg��B����(X��`'������F� +^� ��s��W�2m[1��?r\�����������2�������(����Z�-ի+E[��5��J�֠�K��4`v�I�Cm:hk*㯏W�����J����:ZL�Eᬖ����s�� ��D��µ|�-0��~:�XC �f�JjǏ52�9��ޡ,;��F��z�h�j���(LF����8v�H��J��u9Zl��-�ޮ�޳�������ך�&��B?IY2�9z���1�!�6��b�]g,ҼSQ���]=Jef�z?n�\z�EUtW�tn���h};�,8�t�L^R���GBP�Q?��*-e�8#)�7�!���ǶO���z��7�z���#���H��b�_�J�J��a�E9;'�� �1�lO��9�I�cɖZ�=1�
`ѳ�M��)b #�Q�}jz�귽΂��1G�	��<�\S�C��(�=6K�z�7u��`O}�n`�s�1܀)���-&��-� G=v����u�FVю�\𽉼��N�x��!2 i���q�k5#@	��&k�A�S�`O�Q���J�^vU�XlxVHYEB     400     190C��A�_���+}+D��dD��X$���6,N��kZ%�y.cd޷���ϜJ�A�}��g8.�w�FNI�����cb�I��`�n86z[nCn%{X �[���O��N!@�P��+P�I�:�.K�JûdE�`��C��]C��h"�M��������|X|,}��Q�xq'Xy��b@%Ŧ!��B�F&��#s������F��G�Ð���X*`��R�:�A�;�ұ���"J�a9��v��[��C�����9��E�X�g�<q��`�af���*(m�a<�dI��&g'n��xS� �c3��Vl��*A��O�lЙ�y�p�2����E�W.ɘt*�1���K)� ٨)na��h+ʐ�?��l8Q��<���>~�F�J����s^����[B�F=�XlxVHYEB     400     170fRg]H�
��wҿ�6%2Zӕ���9w�>B���z<�_������J/��3@K���9��D���G�a�����gc�ƕ���(05m@����`�J�>w�F�����8���E�JΣ���{�` �X5�^-�/�~�nX��K4\�4D�9x+��bs{�[]_4b��b��`'��x��g8��D��$�J���)cr���fP�>%^��0��&�U0�C�v����Grg���hKi�e0�C85!���n-���!�]����Xq�>���!��TCŜ��)����/�5L���a�ߒ���F���w2}6�,��WPL��n��u��L����"N_�]�$4;�K���V��������4XlxVHYEB     400     180d�h����R#S�9�؂�G�(�\�"j��Ykh��1_��ky~�lbl�.p�A���r|R�i�6p��7��,�Bq!z��߆cJ0݄4�`�u���g�p�"b8����
{foC���(�B{�l��Yr��@�OZ���!�Q�{�;�����5ؿdK�b�Y��C��,�<��?����\�Q�ү&��s��
����O��o���&ѕ�o�H�!�J�°�"�����Arf�ػ�|�Aď=�z���y@3��_���w�ǂ<�Hh@���lu����̵{p�>|VZ2�%�%�s(ʿp�atTYӜ��qX`�0��t�|XBg&l���t[٢L�'��U��Y����9#w�YG�phy�L��sWXlxVHYEB     400     150�!�?����~�0<��`E���E�wiƵ����߫pvPz���Ec7	��#��=��KA�(����1�A������M����Xҕ|���ʕ�O��1���譁~��-�ӗx�/�|��B�dE�����*A���x�,�b	xh!� ��(�w6������y2�Aw.Ú;sd�����<���6�-,@ć�m��T5'٭1x|<�`*S�y*��s�s��W ��7i�G+�Z$��0@b�Pʣ�* "',b���:�$.�F\��@��N���}���߃�ۤ�r]�
��ȷ�A��|7���h7�����9�i舛�P�.�k��XlxVHYEB     400     170�ɧvZ���Z��p�PHJtvL�,�g��Z"����4�9D%�?��Y���Ӕ�E�㥺�\�I#���7,:xW��;�� ����?~� +0���i�Ӡ&����h�
&85����� �ę��وj��6�*`��ha�>7s"Mh��'�j�ـNv�2�*�Y�`'�|�_j�H��I�si��Tm�l?E���W@�ĥ�T�5_�ꥤ0���}]���A[�����\˽�w6��`u0�@�F!�eLCMfl�N���Yk�� ���Wo9���f�rYK��9i	.�G_����ɯ|q���t;6<x�d�m)� �	<Huh6���r=r�yH��gc�|�K�SBU��`XlxVHYEB     400     1b0��kq�b
�?�`D謀��}� �({\u�q��iC���s�~t�{ۉ޽[��N���
d�;�rH�/�"h�g�,��0I�~���ة�6u�K����/�es!*���K�4�@�S(���OV�>�� ���PӤyh?�l�)	b�K_�&��K�B�S8�T����T�4V���4��S�����Jޝ��'@������](��>$5��yEJ�/L:@��Z�ʃ���L�].�� !5h�W��q�`�K��� 8����,����6�� }��K�{*/��2c���8|q���M�9��iH�L�􇝑7{��+��t���{�#�!' hs\��(Q:_E��l�]��r����;�Cٔ�����[�{m�'n��%���a	 �K��^Y��0/	=���ȝy?�SQ�&idcXlxVHYEB      e0      a0xk%�9vx֖qf���c�L�"I+f������Ңu�J�i��?����UoE���k������D3�Q.�n���6TTPʛT `OuH�^N����!��({?JJW�"g.�`�l��� ��C�J�V4-ƒbr�a��=I@���Xa�I�y�?  BQ�