XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��֌����<{��Z���|v-��'z�r���N�Z~iX2�__�ײ�Kv�KG�1T
��c��Z�hg.Å��]��XU"�R�l�)&[�^R����]�CuJeSdၫ=�%-��p �y�A��*Ure�'_�O�I9ؐ��1���0aG�P}�,�	��җ��jG�����^���*Iå��\�h�T������b�H��v� �4����\?�����@�������ӭ���m2d�1�ۮ^	�8mǑ$��-���}�;iv���y.�;= 8��8M@:��q�����3U�U#6�Ԍ)�˫���!��wA��Nh�T�o���t$[��vNo�{�r׼��;�s��H�x�{=Z͟]�8��0îH�S�4�Yqm!1���H��i���v�5�v��l���;avd+�즷p���(l*�N$��������u%���J��d�d������NV@��d)�ܫw�_��Za�W3(Ep�`��嚕Ɂ�3���BD��n�{��o��@6��9x��N�Y.�L9\#w��!!*�0�u�.��zFad�q�97iTC�f���� < ���]6^)l(�f�*w�-ͅ�4��N�Iw|����z`����s \� ��\T�%�-)H�%3��o��M���+���D�ҫ�B�㾑���
2,	oX�|&ܶ�����P�7"B#���aS�O���?�.�>{��o�Q�^s�օ�Gb��cO��O0 �Ѻ��9�ǹޛ6����V����wpE�~�\>XlxVHYEB     400     190y�5z��j��[|'������ۧ����ִP�	膉E��`��C�3�K�����+�h��,c'0T~�qV�Z���O�Ç��-.����8������gC�F��ß��P��i�����y7(�W��G%�]a�X�p��7�����A�6�\?�@7��,T�tC�\}b�����%��բ�(g��ű�Xӣ~��qe��Q|Ɍ��e�p����Ϡ1�5�_��~�d�O�܊'x��i��ͨѭ�;8�U�=��6�*�Fۻ��g�� ���D)��=�v����O:�+tj#��{��5�*�y?�j-ގ���5Z�!�?�`�I�%�{��pcH8�ʦ@)E�ᴚȮ(6�M��%O�K��m���2ڈ!��m�U���ˉ��\aXlxVHYEB     400     1f0��m}U�>ȶ!q	a�O�Z ������bX������hW��VS���������uy�N�3p�-�=�����#����;�e{>`�>�O�]A����0�RQ���s���:�4�un�[XrΑu���D�OY�I���p�������b�K���Kƥ1F�k�, ���ʌp�����N�]�#���)���~1D��Qx8�B��f/�������o�KKo*�΁�i�J�v����!y�ƈ8��I��&b�F���TN ]�L�L�12�&���%})_:�  Y����M~	ǚ����.Iߜ+�W��L]T���8k���scj��MZ*�.��I�A�C-�PM� S|�LjI�g������%j���Qa�םE��1:p�9��ay*(��� ���q�!n�T����������/M�2ݤ*へ�>nL._B����
Os�3�B���Z#(pMc�5~�߫�rɧt�x5XlxVHYEB     400     200�fZ`ꗉ�pu7�4&�¶��L�T���iǳ$���4	,b�~��c�XSw�l��I��X�D���'V���l��f��/���VT*�q>6�i��q(dհ�p���>�=1������]���t֭A���oРS����#�S�
�r{b���^y���w�ŝ�+Cb�v/aݲ���XK>K:���,.��KR\_w��Z?�iū��2y�R�qE�N?��z��k Y��U�]��?&F����}�������ѧ�]��Zab�!��ւkѩ:�,�����KCN�ޛ�I�QZۯ&c�;�ܦo&&+�و�D &��>�B�,8(�J%Ѐ�������umt#��v��e�ut8�g���2��s�0��tW*���n�B�K��ή4]��w8������83�m�3�j$��/���u�-I�e�����7�8fG^�w%'�(�?��m,jgn�׀�΄�F��\$�����@�>�1���%�G�^"�XlxVHYEB     197      f0�׼'�7�*�u�B�;����X��Y��5����1�jXɺc`���*�����i���4U����/C7�=��Ya{����v@y�YRJ;�q\�`�D^�vUC�>d�V� i�MO?�S�s:R�~�R���1$�c��.����<��#��:��p��ޫ0ը��F�R>:qx��jv����n��˹��Z�G�j�ͺ<-�#m�,�=�+ik1��3~~�W���ח*�F5�?d=��=}��