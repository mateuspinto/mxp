`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
QF6KfCYYsZxu3OHlcYiFtLkbArIGhdH1c3Y1nnu1/sRu98Y/+JhSK6X0Sp4VwzSHpn94CiFse3pH
LZvf7jnNLYaqf6aELrSQOl8RHaddqAreky3IWouqDSvIIXnFKHRj+1aXnXGFKFCYMSkk7ZPzcY5x
hETcV9cWzaLCtr4dtaCbiMNRFFx8w7g1st7npxfciKZnhCG07D3E7/LAsR7ThKOpl9iyADd7GNPP
Tp/DlTIuaxQ1HlZPAeLYElK4qm9aY7Yv8fqqdB9PM+3Ks3NinfMj36h4nhBjhhFJ8HxLHLVJmPcv
VRw6oXI0TQK8NhzK8PrjOmdMk5WKDvWzQWjUT21Oqk3FuMGUakqPQePT66yvrchFuA1U3RXLO44c
XutflxhV5BzhGlFxrH1U7qJe4aMhawdGMLxBNBxxME5nOLPlFyARtrjQRjGHXzvoVjzff2kj2NJL
UTRevkYQe5rlApDK9nTtv4i14kNsClH23zjTTx2XaJ36S5PAvSlPlOnHMSHkjugatq935vaE85aG
KBbw1B1M0hHBnClCKpnu0x+qQLe17ABTTadKRMM6ATKngd7Cy5EzX5iAAquPLL0/ANykUSgpKqie
P4qxEaAuLgWJvAGH5rDDii89wTsk8eMIz5WzjtH7WTlVZWREjwawrMeXdsHKqWTqUk5HvnWcFxEA
P6aFHcvxoh+8wAR0AHPrD5aO24ggwqvjAdfZ0gBDPKPmcsL3nuHleAQ+hAFqrJoLx3EaFwiFvZBc
0DzqB00kiayRatBwegUbi8bptgiDcsSA1rTq5qpN0ob0atXkipuvWaME0Qhv9KbhpCwTSpfOiw9t
kk8ix1DIUzA3KGQbHlfSWJtuegtTsE8t8zvbttOs9WWtx9g1UjeVK9wOe84F4YZDe71BGEjGF5Qn
ci7vT9Yko3IfgYf4gzIQp1DWKNlq3TOEfz2ZKZfIm16YYQXSzWijCqLMOb/Yr/TbyV7FnPhAvR+s
pgKWCLyg/AeKCEH5AXA+IlFk7unOFOOjWHt3QKo27ZL7OAQtcHHXI87AF0Cq02A1ozsy3b65EIP6
mb3u7rxVP/LgfrgmCr07vI8HyKeWgIDKfiRlbu6Y0m/cXKZ2PYCpfapPwFcX2xRQ+oXJgldd8qNp
wXhXhBbNloIksp05ba2V6FmyaeIDSsZh0PcjFnQ4FHegM2aOKdi84cwSUOd2mnrr71VvJiBVBK25
86JquXkBYOiyP5xA0FuEfagMEMQYt8dduz8vJhy2Hcjn1Qzc61AQYjxCyEJncHRJfnKKaYlHkciH
PHCQVNHaET9HpVzZybVKgXtYYtEXNY+oxZcTJct89AF2VNExHL2bZfOUXdNaHvrTm2agIrjuY2qz
OI4y5FJGXeKvxlaMGBv9+gMLjUQ5XV5io3X19hNxrpZFTfU30ByQEO/U718pTwvYD+GmOHon1h8t
Fm2ZIWCDlffI3GjV+KFs/atZk+ZyhTfAPBXN7MKxBT96dG0G6okWT0+/z9uzQaBklSBcwsJGnYPb
n4mk9OlDQQerC6UeXCvWMPKB7blL0+X++W+8Vvp9/O3nKfd5gLHCSu6xd4eFQsh+brzHtPeNUKW5
JlEOULAr090eX962QNdU9Bfn5PZ51r7zkdng+9Ho7GIJYngu1BONLZYZpv65IsxNiODyyV927Kob
AxLbnSIFSk7jewvRC2Funrbm030d2zH6b3iCXCGeK6L368ViGstm9l3vwMGpzpyaUE9JCvgMui4F
qTnNH+XO7uo55NryAohGOXethKHgzJ5pcACTQp1TGlP+mau+WB91Zq1Jg/borkPrcYLLtpstMOXF
srhW8vbnWwvvKHPpQvmmvzdNOtIouo1KE0ud9yYY1A70mR9gurowNzC/6/RpHEhEi2LE83PilRxp
QZ3XmxdU6FVnrs743SfqDvJZrBLbLvJjSWUppxU8on3d+i+ky4X/O5SfKS7bown1+DsQ6BBieF1b
k6i1YdHEK5hDDJ7I5C8ENH9hgPeSFzVQLn9NwOACWPP2XbTO3HC0za4c3gsFGfZTZOi0dQHXbnWN
jYn1xNXaU498Avq9Kgm6tODSQMBe/1pA+FgSwiJ+NR24BVNjMkMJKL7Ml20V2BFfNSdIgnY376E5
vwiD/h6O88edMKf9sT6U+gZzRTsKHfmcC3HXgZs9uqTdSw/fORHdw5Pg/blZqPi+A/g2ojXy1LR0
tNM/a2qg+MgXrtmU+wuHHWHt0hyppIjbzbZC3dG4Q7iuBL1ZgZ+jZav7VkgHagzLUC0Aew+6ajpz
ZtYIPG2qJ7hsQO/76M2K48xYnfxmYvKa06+Y18wQ8c0iiJZB3C/jee1U1s5dgtXuqQ85mnSTB3Sb
3CbO/jZ9wO/FcGEUCcr11JDiSV0ylQgJxfMO3BikU2gm10r3Vd3GpASszJVCIJoIgst8PPhOaNU2
xymsfEj6svfEiAIQga0zD4b1uGEmVw7gHw3BZJL4phjOA/Dy8OMrDX9t/TtKAYE7lJg1rf+YXdXi
r/3atY3rzawljSe81miebDk2oPkkKW05QpYJbB0P+U0qqHVigBy+vAhBQoiBba8wA+eTWVHfqbUL
EVu6uA/cAzVkNttsYKs1pg/h9IgDlfQ9qFrTvQZX4qogAPnw15YcktLaF2v/siO6zVJdoY/hPQVg
lSM/gS29sum1DE26OJli+mlwJB4ufo8JpkYF8rKj4Z2sA9erosk0PkDC2tw2bjhKMCWLL71gdnXJ
ZvHHNddFr5TXoK/BVistSkoxge3Z5xHN9x1tlioj8uQ/p4F1wrb8ysYFSyAMxay+ciytIAS2dPjH
0CjxKt4lSdC6U/6gZifGYyTen6X4bbErzIhaAGcHOemzlgCkp8/JlOnHkQju2MwM1taIx21GVWYC
CQFzhPsqLoK27I8WpU3ijIhG7XmU40Q6cqFaTtxu3qYFOaqVOFQ7lVAXepc57IuQm5AudfF0Fp5Z
CNgAxkiovDd04lLtDeGEAbz/PAAo723BLoFzMoZLdC4jzK4+EdaVv40CpL+xqxomPJPUe/Du+Pc7
IygulYtCqm+u4rfRmNAKZXU6bNwnBN5r+EZq7y4nGr9krlVrU4MVUYuLPzCMurHj4LDFYII1vS3C
Z8VMIQ/+QjgF8XQKA32LMAaA5ZL3DGkNJ85yl1ibPY9VGWwXSgNAWo5fLwPNk5xb1gcy9JxSjXm2
6yML/3LWdwh/YfuxzjIkyAlLb0QffC4tqOuYYQToTMPVkv8qVb46KmWW/RJ51E9X6OXf10A1wGSl
BBrjnf+L4v9NqSRXCIG7CaUm247FjPvORJYuquZsb/ApdZfn6GB8qNZRikuFSHxZKSLWwxkQp3xI
V9VKCNF1BLKCcz452iimcK+RWkX7OzP0m+1GdS1NDWmsQ8m8KMkEG0WY4rG8uY/THcZ5+B9jtH9/
4IDNo0nnvZC4cnhMP6Q5wLx2ZpnpFQ0kRcACihRA5TYkR7MreqfwM46yKCXnEUPidJR9isFdW4EY
VlLSDE1ADAUj3W/fvv+Ha7afk93R8f68jE3q6WA6y+l4V9arRpdn7+uMEf/Q62HfdqXEEOdJnaHY
fYZDpsMv2cpZfOg45TebbQUeejm6k68ppe7lY+ow6T3UU4tpRH7NCQU13Y51SEalVs9qZBGN/7ew
5XM9rdkrSinGExWcygU4bsarCZEWz3d5mc8eWPtqBgiJuVTif/oSHFEZbJhEX/4yDqy3TzkDxJuW
mgiet0oWO2X7fmffYwVM13mioO8tNmza+3H4M0M5SkiF9gyRusjRULb5D6fvdvobk5R2bLRmJg8A
TcmN2t9xV/3E4mhd1RbLXkjs9HL1DfkuFpubQr4q+xJgclr9fxOfrJIwJGArzGbj/SflG8yeXAbp
GzAuYrzgZp7k26l6JciOXxDrNXYIHzrMbwAQNVyc196tia8ry766yHIvv18dl0jKZSb1mSmb6Mny
KCfUPZdpfuX/CPK0BZZXJU/F0l4a5NQuiFwu9z3HWLY/TLqzfZE3QjBVe3ia95t48tfABO0+v21q
VaYv1CIDn7LAJ9nHQUnqveUJly+nCIe9k03oNo5JjaVwfP3dDhDeQMTtMAvf+30NHnUg+3pqWbvt
dBcha/Sx1I3wFmIBKVu1YQ9ZcPP2yVQz/IFZL9uDphR0sfzD/doC00l5ZM2XOEWMd1AvHy5iZhKU
DxkBLL6t0teYD/U8LgghYQDM33wgISVb6c8133umVKOnPBADfOVtJua4JNI7hAr6DK7px6aI6lXn
garDiPVPS+xQpPurbkpIEnyXEEgIa4HeRwvJRlaqcWmZ3sfGqTHkmWx51dxnWnn70vVZqpkJeZ6p
D3lFlfb+pAxn0XcNbXTq5t+RSXb6aJyeiYL+HVLZoC01NXmwd9/wBusIOd+PMceGz5bvffdvkC2I
6+3ope00b3vWZYXv8vwTJ3NWELX+57JptfO/IAGy7Kii9+P46l0HJipImZXVBIlut4EjbevYvo2g
MKujDWwCYc+QGH93vvBUrSybtcWnp7hfuN95qT5HowvuT7hhD9Q7ASQ4qsDmxMfQVU0VrN04URX3
I0RO2E3i3U6Bv53e5FkMaUIZgKy+9muWedDWDA2xMLAnRkPvKBLb3BNDzdmj7zWPhpRNvrVgzpqk
MJ3wPl7AlEKgoTIqKwjJc5ypjIx7kMoOM/xKqWS9CyLQR1/O7uwTnLW/vYR42IL5qQqgPhxSqoyC
CRD6eyLy8xm4FdARIW70o2QfiWjxWDjgwCZnNY9dqljk2XOtFprfNnytMu62Yv2xHqSNS+VRRlQ9
hRNtdNycJqFG5NjvV9B4zfICVhK0a/PmOsBlSmS6SikMGY2IOFSMYn8EUB+uyr/Bx1LMinFCVFkp
mwzAPG31DWWKR2ZkJARKpIMaP9ZB5xHGBg6XJMVHPbo1KFGpMlTDIOaUEuWhBQ7z+u3/nQd0ak3r
lon+O5prPxes+Nnwk6YF9f57xobciE6UZg2/8H/Q2xcvv1T0DQjJgTX1YHxT8olKOp1kvutIG/SW
8ErP8Vn52YMTx7ytJg4rIPvRdlaeFW6Lpfns7exppB3Y0dpFm8lt81eD9zu5Pz6WBH71nZ8hEUT5
Ex0zsLDevwu1nw4BGrFyc4J1p0ar
`protect end_protected
