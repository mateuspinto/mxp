`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
q8dZNEUC9SouomKLwjOqJcqDGudkV5e2ehbLi94eVgsRarMHwGq13H6AyJnZWs9pjl7Dg+2Iahy2
o0rWegYAZYKz7Qs2IjrolmvNwfwlZcvNwo636+SdgIEM+pr8ytzLeZIGprk+VFbPFakEYCZlxcUE
ioDVIWoyu8GSDr9HbOsXCtXLkPwD+46F9xw0lX1WsfK4y3rSXw7bn1EHFzshTFr6dwQqyxDyJgsN
qyWHet4O9LVY6z6t+0HktMdEhAwNiJRCF7txJP0HGgdHrXR8KfLkxLvgOQW49C37pjLIYu5YWIrM
LTVxIZzXc4yCHfEG+4vHNqvxzphnjqsoGCSZs9gepwo2btfZzid0OJ14l6nXd2aZl9StsOWXAt+/
S60yihP3sY9nWk8cYUN7aTi6N2PAUWTjNYv41+G4W9spARl/kw6KxKeuwUvFHj7jByw6AY8no91k
fBk7DBAYZ6yqV882jw1QQA5nZmOUGEb3edzyrI7GlIZDPIBYz19hlB8Huvn3eAXvfDGiEMfm+xZo
tP4t7AaZHEDeKU6ayh0AOBWDm+MTXk4Gp3PJ5nTOGMX5bLCX2tNxZFeF710I3fQOstmnrl93TSMC
jkEk7gi6p5hR+Tq3ruFm7dPaJbxK2Ckl6OGQOftWQ9BhNH1n6qIrqCj/RqHMUsQlkVDg9gIY6PYD
KBmAdx3A2uffkU8VZlfH3miYKxyfFH5J/Qdkzwv7jZ/aC2BVrjv4ACVHfzTEBpculj1mmKtqPoeI
dDHNF3W/uDNl5+MhyYRFsqLm2cMBL2FnDDxp8EY1/VQBDFkqlrUZ88sbIGrSdjAW6ymSI5ydQsXO
VsnCSXwzpinqD9iVwoads3WtV+UEpL82yRR7g9PdwTbidkHgaZEWq6hDClvURz6lRLnxgsEfxTxL
QqMS03Zoxyo8/Rsjiq6sy484dYLEP2u7tfdxnWVVhtu2v1fY1BtVkmvD8FLx5HSdANTY+rOPPRek
oB0jwZpSpqaEty4A8F1JgCryEcwGazStSLSwJ1yckLhD7Wk6YdwGRh95AYOsniTjPmhVQ0X60d/W
mPWskVRfvCHMkXFhm3B+arTCEiiLru5QyoNvCQgZ4RBy6XVL4Tswd4Y9O+q/qcspCAOCLNoIrR+F
ji/WrOPXTEcJc0y3CSR1g41+NMBUb6ZmvvVXs3/D6y3VIcyBmN3Gt2mOtSvd/u9XLp7f0HmJgR0E
wxptDmdPMGi5tBFaXAMduCsIFDjkXltkJMgg20hyYGtCAM31u8pg70OSe18XkZ55ixHyzKIYEv9L
UWDR40jQirYTf+5tTgWFgOy0g/YvNT+WNrjWvl0L6crcr3y7doW3YEUYyignfLXEAyGzZwpih4tj
u0V+vPrxAycQtiECGl8tccKj1hnIQmi9ZRc3iOsdHK4f3hZKbB36kBH/e0vl+2iB4caf6ZH1bzaY
vGruDvzms+0lvEFUaGPTIukzcMwey7LlpCQnuy3qN+BP6UalcXD6zcQyBhyZnI8lyTxAM4Bkb5xa
zGT9OhSh77f9o11FYJQU6DW4vAwBOwDts10gw1i8RbRwZYMYQAgWNgvrWes1+A4FKmWQSB7zskK9
BWliSGIgycmRcqcLID/tfyECDFVo3kGWweCC8A95Ndxavakseu6xIzZ9c+YBDjYORhEyZD07CQz7
axv3LfHNHPcFRVO0GWEJ7jon2BtsWJDqi4sAq8HmDSVbB7PzIkx892t6gsWr4QhBMQ6nwYPkG2ge
14pgOZsuJme5dfDsGUXBZkeeCf0UQ02VZflwVy2eX/LrhLbKTv7BCRG9DuowcM7YiNbs5vl+Kdqz
AiBqUPSg+Els7qytYlFGTXD0Y+4jv0mdXJQ00EdRq4YvKAQR+hW4k3qHti7eg70OVlGtkiD+fSBg
C/q7l6BQnmxsbR63LDNO46Xd9J0MOAgeyP0MirIuaqAUAfsavgRdocY/sVVd5B1S+VMlQg7E3pUN
tiWRNsQP16Qj+B0mg74KNcNVgDZDFkOYos5knsHUIr4c0Yi5T6PEETqt2bN4tLhdnjQzCqDsQNcF
z+ruZOm2tRxSR3DWm5aM7pi0a2+RpqdmkmEiRdqyiDB3I3f/I7k+o1PpmC1NnZRdIhNvdkl5rZZ3
pywlt9hyIx78c7R9ONKYHcaqu4jWSLcrcsIABtk26xWeAhtZqI98vSNm6X963ny0mze9X9vkZMSJ
EjdBZbPS41ZTMfdN59BZ5AURidZwMsN7SEKTLWdgXJU7SNO30PJBpkv3szph+KUV7xDeztxuMGvS
/8SIg6OXAJ5i5NEOMDxzj7VRPjr6m4jcJynvtwQvqgMUz3eO+HJFpKHNbdrciz9p33NJpOl44T2O
g0NgE1HL2XLoonj1yCg4NQJnUm77Qim9wdfJU6st3VHcVqHxKhUMNbstCe1oI3ATTajF6fCVRZw/
oUKSgNefQ5ozuv507U/oTQ8GchpEuB1+q8tejoNUTZunuDgBHcqennHlyTSxs9ARukaBxCNflnHN
Rk/irXhdXifGjVyZmwj4tSns14oRwlS80Cse91381LTdaKJ98ah7ZDfFfV7McIj+BhEGes4kz8rU
SOtGkOXYfiAQ3Y4lbbxgXMyc8bx7FlQo2rOoJ5/ynR45/9lQiSpUO2dFoPwe15tmAWL74VHODegy
Uzeh0g4aZjyukQiOmbQPILHjm6wxN7mL1wvuZfopvk4kKFJIjzxumDdXB0vnMc3RYbnQMTvBLhCF
haS9ijfBHImhvqqxJi7X+sTy9WOi6mcY8HGkYR61jChR9Rk0mCodMpR1HPNOsKhodMV1wqPOqnrj
TWhrZeHnHwwhArDjERXuasa1ibmNK9J5lqiEnsIc8UWTMbMH8/O/lviHAzUTDCx+TzlRqWSVrWD5
D9W52PRyNCxdkclxLd9/9Y5MlmEkP2fALi+7t4mOP3fxZHf9We31f+q/CcXJdzLeTnRVLUUe+lmU
jct/ycna1N7BPErnJRM9xdMLkvVrR5MSMCFKUyB8EV0YALfOdTssoE0HkcUPnF4caoC6Kj/082JF
DfNQv1cMh2QirprXpAemU4+ln2iqcAvKu6MXn5L3e9p7g5Vn8lDtEDneJRWInQ1ATzOXxd80+XRd
X/w961AZb1TAoVI0Tnu1nfKlrLS+5l2cfXcE1a1WbPs8dNowYxo324a+lFQyS9jGTFC8iq9tYefz
+3K6JmrxXGjPkMqdJQRQS9jzkXUijTPVniSD2RqSacavneAalZFo8v8hvnjPARWv7JbI0cKgWBAL
Z1WtAV+ycmZ7x3PKCDZq6OF+cnKcDdjeA3nGXQi3ykQAg6iv7z7xq1uVg8Rs8XOKjZiCD9qf56C8
/eTxfhzZN8ls0UDDxHfMjaMs5nAHYE+38n5ht11LeWNL9eLtlmpTRwIwr7CH0dM7DzcZD38lnMjZ
U8TIJXHQod4y2HtW+wmwIGPMTkSNk99ZOsO1tTDGqB8KGQkp+EeRFO7xgFSWunmo/1iXwwcGYEqm
sLaADY3D7W0RJTiRIr90z5CHMZQ0ionHvlbF/N3JdIU4CZdJNcVPsIQiRBAO36OydsEWERTc9jwb
LRIwc1cwFW1ZzDr43o1YfYD1yVP9epPDibM7c1vTsZpmgE411OOffYyk6Q8UNCJSoacsmNHjqlWN
+foxgN/RfrxrYmpAMZlxBtzQji86tXi0QrPz072kYDnN+2tXBuw75fh7Vj+/64srE+syjlOZevqU
qnHJUbXm3g+s8DxYaMsKAj5GdeZLEU1G0oTt1pDjpX7coLeoMnnRPnR9vrHXwGp9J5ozvXwO3Fyn
JxDfG0zVA/bmjrNh1yXR+ENTQSNeelMCbou9ffBhiB/kARptoEYkdNuzbkMRXAiAFxzDFBxiF8C+
PHk5K9ySqBPMPO+htEh7/o1MGEVOjqVxYHIHWVxa0+OubiwfqJfOq0cypW18UjxvICaSJOJC5Jmc
388ktHjyLerSEXxeFMxhNbtf7ARFI+apCUYDmcQ9UaaywGahJvIoonUJfNqaDM3Ry55nARBfxGjB
ISRSvnbO6gUaYNReZG/UMcLUneN0KlauS418I34GK6Ff+AwVR4H3aLJ1/kcoksaZLky7ZX0zb3SU
9zZBqzNZ+K+3G5LGjCzF9d1656i4/Hl2S+AHwWqKI2KKIxY2mfmuY52fXlcYQ1jSKAqdfhZDziTM
DU3WAsklIc/qo0brxcgc9p2vQevrAWHnqtzOKKPk3xdPqVBBla6cKTaICHaEetntZnSqrGP/Q4Xk
iPRfkXGRdyExtESiWuOdO60t0I1QMpD7A/KyhXgny2rBX7wJl51vzNovsQFZfio8FaU4NndpmaE2
rgWdsbgqjwmZUhtAoaEs2AKDyctpdTTH4MFfpnGjE6yXYajWWT0zrY0W/nk71UBvZvei71+lVX1z
IBkFq8EgdUozAIV2NFSstUNG4Ly8pMQEgDZJHjqSBuFnT+aC+FPo/N0whOMzhk62xeH0QVQaTGVt
1VD8PgpuxvIVxxPMbsrCmG/GCKO08JU1kyaIkbMGI/33CsmhNPi25l4+ytdDhbFCfCAgX/wnD5fz
7rzg/EVQFjZ30IzuxlMlsTfYwSqIMALZEjSEswVTGH687GmhnpxnCXppbmyTCDrH3fn+W0qOdAP1
uPvjRHMuiBJLSO+67YrbPrtw3DJ9ny3Sq7uri32J6YAc2TP28yQ34NkeiYQ5HKwFyqYS79X7nGCS
LVLfMvxZHpsC6HYAK+wGW4hLjvz/zJVO9BxE/5GYrxZoXr6Sy77GcYmo5D68qA7apfoY3V2RaPSX
ESmxx7E9CwDNmVYmwYopvAio3g8RPfq+xkS5/f97B2wXxO1nILNMhSs/CdxzkE9cNiIruCFk1+i0
snJhCUMfwl84ToQhaLNjcE3zRJ3gzeDa5na+JlYWuhy8ms/SOX6nBOeSydS6QwTVl4ZXXZp8ycHd
ucyEhOsLKSCRPEFSDpOj+iY0+YcnR4lEKcjxtUxlNcAJxtsnvByT4dNNABULmjINIXmgVuCALCIM
SF7KifDZMqnybxgrBlzsiPFp3CoBwwT/1gmqFHUqYi9bUMYdmik8rvBZF7jbvvALZsi4bw9oS03N
HywQ8YZeAV8sFuQVJWkyWMGqjAGyIfQGRc6JddH9tYN6FDsQeUcpT/mBAog3Kkiv84kHpUkXrzBE
fgBwcpOWYCKRz66IoFdc8y2UDRhIY8QxptQZyh5vlpBFgACesTfG7uv6QJpsGEIuVSnDtKgzv2AA
JZYqLa9wUVzscW9ou+mWYiMQI6qyTon/hdjwtcMH3aVhvvzIIAdyYm73+fHe64u+knSd7Af/X1yA
bboPSwHYRZ69GnchNt6yUM9B5fAOuDvhODafhBSAa1m8xBqgkrdEsKN1DiAA+LJLiIYMn7/HcY2J
IdEoHG0tLARBorlhdfCe/2T+kcgKyWx/rNWLiS5yIWbc9n9g+SRG9Xgnq+2MR02EsULMlnPFivh1
wP9TLBe7toH1pZ+wFCykNLkjfR0/qAJ1HcRUd+SyRBxwwebyfV9QpCrTmwWBnVIE/15j4Ei1UiMM
2PMaQX3zhzDH+m+vNsq4TfzIUr3MZTTfQ7Y5P/QPrBx8SuvxEBn6gf23dDVCihgXuCE0DpilsIJt
MF02DVZ2xG3elSdv3LlXFKK1l9CcCtxGikNqNGdbFz7gVmg7t1AePxmZH2HG/Vooydwb3nMzHl1s
UHUzTq0q6QxWuZtJFsl8ycN5VioE1BxLkdnozMKtOqLO/HyV5do2v9WIl7G9AQLttgXMCfVlOym2
kvOevMO6j8zGH9ZJX4zYSYIhJchfOOH4oNC8DmKjV4oYwadGg/zAb7BIa+KwkWeygPjli3hLp5Dr
ZxVvcSuo4eEIcKjEFAq3s09xK9PXoF1D8Kk9kWjM8ViX/5fpAoTDoLnjBPeYmicWhNX6xqepuk54
tzvceZVboH++LGQ+yB5mQnqQY10yllzkZcjK4KwWScGS/zeN24/vVG9i+AM8psIhYrWn9TmcxLne
ofWb28HPYbMm5QpsrAEq4s3C3CBO2gnH8c4X1iU2iQFpYZTg6AUU5u/sDDHHEGqcwQ2YpJCKoWPA
MCVjEJqoVujRyPC1g0knU6rbWYpry5XL4g490DJpVavYGRIx0wwUiYat+K4GyshM6v8yxtBtV45Z
ruNf5YKNJj6M3larJ+rTltRwxFlAG13grtV52dfhb3u7o1s66sckFqVMXBIP3keqqNFevl4oxNFs
PvttQ+2z3SgHxvEacY3tt7s9dmFx2b/QStXhJ19uALIxHwbU8cmGkPLg2FTzF0jqM5XaOdXynplk
TdEAhHasBumnfo0hHcD+DKN3yjmY2Dkvm96NFFoVZfySyK6em1Axx/invbYa2BFMOI9peV77JpKg
QcDFCTqzSFEHk8ip4nDA6vuywrgW/UATQlwu4IAy6WUz5e/LLIPXZuJObZQL7KiizSPfK32yxeHL
nIFfWNXNTKjA6z5MNA/Hx8P9+J5N3tkNQ3Hn9ylHVpRsRIHLsW5U4qFnxK939t6sHRDqCE5Iw71J
FXC79XSlPjsgkhN5TUejR207KjbnVbGbL7iHGB9uIpAxCMus/tMPveAWg+KlqkkT9hESnBahAPcI
A2BMJs0/IbwFi4oSeR2m4CFilhArHtsMq7QqRBTkPtlDeR6qCXIBiT23Do+qylhHdmhMyD4Rvp3b
AiDIfItqaVfqajW4+Vybi+aTjgoH3lxMoG8LHwAYfw5rVbGtYeDw6qDw+k0fsVxutbda0o46Gd+p
aSiiW9sJHfTw/nWpj1pupRJtABvoaajwANrLeYavOixXpl3eAvmfWjozg/d6IhHBOOgff5ocCheX
ZG6V/iPABZwtiiUZuP3HzsdKWSXyH2uHqk71DM08ylgnLo71LgXwcuHT6GTBTadtdiVTdOFGLssB
sWozCjCUqulEMDNk0VWDO7YBzNGgcJY0QHlbBB9hiiEvXTdgf53uJwAK6TPhbR3MEKhjQARAXMPP
7ibC2z6d4Y8CEyxFWyM8zoMkHXxRkUehUNNqjGwIGFXwJ3Jo0SOCuCmp8ws7zYX1v35LW3+VbXXk
BLxsEglAZxBJxvJduk8GN0ITEQcXbWpM20bPGISsTz+sJJMehvpcRbt0BvjfHV09SQiLnL197mBX
5+r+OQO9thOjGGZNLR4hKYN5QZhdB82R3R2Ya4PZ+oqfgTAYOC4Sr0yL4Sd1MYagq1/GHjPJqTMJ
d/1K02fqrX+Yy/aqOh/hbT3kcOq63c8T3IzHkEAEW0l6LviqiW5UIdVze3qB+g+ArixzXuFgww2A
jPduRODwcfLk3wbVLk4fqM/iumqxP5eeGOZvDveceyd85wvTF/cRj69ODifMgiKQvz5D0WRvMNY9
bh3NTVLzuC+AgqYoHIBkmPrt0H61b+/CWBPzUb0K+7k30detlpk9mfLrY2Xf0Ez+zkcr4HzuzfXR
bXexgSNc4bA57JIRx2GJ8R5M1q82USFePg50qPIf0vvBO/UHSsp0go1KD2g88mt7XzeOWrnJ7Pk+
Sg2IMaDBm4FiowiZ94nsrEPIk8QYIUNkbemlWLfBZL010sjd9eFY1vv1KhD+H5GJgvS0UOhT/9jj
p/xs7QFjx9tPc6J3atwMMmFwAdtLefRLA1hzUtshbZ+BeSKHCuoM+Sgzcrm67TUr7zRT8V8sgRv2
e5+B4GQsmXV2r2ItsJPkkGIET7wWYar+NhdwzOkPXfky+ujNg5+7+Q6o8zIj2jzJxZ7wy+BgivoA
ZAxjPpGJ1lZOg80xOSKXB8p/BfuaJf/rpyQnQcY1zyq1C/MhdfNr/LEEeN6DuVJBCTjwddqaxnKK
bKwBG2tQ5gThx0dfqfKGlx94HIpwwSnjpqX/SCrvQlLV6tDl+ItuLuujy0aSyadLAWkghdOXSNsx
GNz3St7vEeWcfqYwGDI/jTJVoERsffc5iPu0dXrz9ZnZC+2XJCmSLtHyCKVY6/i8WxdocXhf8uaR
8iTpFwckVK4dgP+1zbhciEd9kMdv9Y4rXAXRsu4eWrGhf1SOMSIFKUFigp3PKaOPst5SI2utI+xe
lcomWaa2vUdUFxhbtTBmzH+uAY75+/ycQqqP6dUGzoCOh8GO36GCii22CuOmeQOe5MA09bdm8kA4
9n+hzfGt7UhWx2QKAjRkmpmY8wgAaL9HVOebjhxy02dj6scBvfcX99vj24GH1t6CZnAXAn+Dfsxc
p9U0ysqW/1HSG95vXXwfz0ZfcqAAPt8fgzGEB0MJvFkYwXJziXkrSM04NM+54n8dOpk40YANSqCF
DyAupyup8swzCeC9FIrdOh5rBgMDDaDM3UcthKszgzn3ojxXJzVFwQD3N7I5fstdUKTSBnXH1YT0
bwr/RHMl0GQjsKMw3bEe+ba4ywkVbJ2UrvpGN6Mq1P3Dh8oT91W1uXSc4Mw8QNaFNJY5UHL6vUR/
/BsQgpa0BqqWQ6V/nIhxkCVddPYrs3pEizhEyAGSIfH3jm/o2TNqoh/twxLfXq7vA87v3Z4nqiRo
GfHmN/mfZRo2Y4SgMGCE1wm4c1RV0oekEefkGnc+EClJwM47aF7Lb4VuvSynX+n+VNkSuh2oY84+
RSVUPd4fIJ0ERkzo69fVMn3am9IH62sylC3297TRecHsyMbynLqpw9DT8A37hBmv+jpxbIbfbqHz
QN77D71x9ll7E1UFpHqfhNtBduWf+yQPpHE2rivwW84OHfkjEEGw5OWo2b87JlbMSlrkYK3cO/NB
cHdOGHLxXyu0yVOnvsMZ764iw4jmkZycDH7MtRPFwb5iJSf0wHp+0WqMlnwR4a4Fs+9t9E7b7fw1
76yqq2QKBjSS0eR+h1rWgTrMS4adeNlPOXyOkNieIOVqS3XSdJRw/cVzLg4agL9Rvg68/1aq/j0Q
eZ9BmfVXciTTcdDH9prdeTirV9RcuHwLrBLqNuRa5M4Sf8sHuRrz/iBP6EQY9S3YxZjR8d8Yx3w8
X6xVp646c53uG8jdkv/eXDQ2ME/2e7Pq/T/dZNsvhcMdgfZ/DFxlMxR1Gv0I9W5R9r4+3fXN9UWk
PWXMjfts6fCgGLOi928qZfYgWhTcA0OUZKHZsKAHix2UPEM1ksiexxbKoBSJuLRecJA8C4N4GJE6
8XV2I0rbQsVTU1jRXJl3m2cq9WtppZ+9BDl5gC4f3eFZNH48fF0B6aqDCEZiSBvkOiioWDbqDu4a
e1vWVg4rhK+kQUf+oaJI0GxiZ4Ts4YFLEUDDzRVpj7DsnrBd49pK6TuVOoJGRkUHAdzHFTVocAsi
9kMd4XB+dzxmP0KTjEniMCThtwLsgidK3HmNEBNDmpeAop1w+fPYbXIlY7qLRcDD0DOEfepSizsp
AJTWcmSfHFevATS9yaCEqmLHFsyiwy6A4EwMr3mr5cmDCsF+8U35SMuQqqVVqbphwWBqQkGSQ5Kp
UQjclHKAee8Xd/6mw4vRPqbsj1weOAfDPX+TV+urJYq4WIw44VETXOVDMZQCR0zTWvJws3Y2qfOT
be5SaK8g4wMcm7XnqwudAUQG1w0CybVKjTAlRL7kYhg7AIN+Rudi6IBQgv1vsbODaMTYjiHdNdnm
DKXhznyOvXrTdFCx5ek+0EgrKffLTRXNOj6AYjhczbQAXkDrxlpjpJCNfokPPGZs+YOpZJzw1zfL
98aT6s1QK7dKBVX4GCEfgmMrnuRGOJfXJF7H2dcbJPwl3o5OhaVW4vpCm9nodrGbXH13AC5hB7iA
EuyUIbmoVJ/xaUA+dF+ZlsXc+RKiW0w8oW0Kf6SGCXfI9XPNKrAnYIcwb5aTBfEEcp9QIK5sIVOV
qRpufRYOC8zdmUkHfJ6MYG2WSMeeQmWg4lBe3Pz2ZtDUIqAqIp8YzFHfPsvw5s3ravldCIUlR02e
mMhJVFHbGh+xgbu96bBG/wt0EpkZSdyP+eF9LHd6pXBWLYrnLLYfI78ErESC51Z//bOS2oqUu1LD
OyC+5/ocLmPc94Kjgzq4UBLEwx7DctL4yjgMaJbU2gTH6zNAgaBPCxqMta72Cx3jS8FW4Zt5covU
jFAlmhl8oWJ+F6Y5MXxSje2pZ4cr0fpjCiVCV3CR9tuD6HttuYqxeeSbG0LwtxRf+VGSsXy8u3Z5
nI9G2Q67nP6PBhlKXSKdzd8/nKS7Svul9Z1K+deUQbinKj+lHWxjvddhrxL6UzQ8BcqmL2GA36+I
bkcHCrgAcM5Sc7FwZuhBHi8FTtDpTA80fjhwQ26x1SrFo3hnptyW4QRVwtCA4il8Wo7JsmhbukjX
zmzocA25qA+CDZk/1ba8412YKPNTgTblI1gmdsi04BOBuB5WvO25ZSyOsX5iCnjmL2q2LHz2vUML
IiJenSYb6BAjGt9WW6PEujPdDC9yMfZYwTFLIOvXZbtu3pP7xvTtCBvUrI/PeFpinbwI61ykHgX8
eHN2/DR1pAStDC3WGO4EBY7hH3KOjnd7y7TG5SSP50/f5AWPkJo3F4Lzi69aElo61lwKkTpzcJi1
/3j8sCIkURutUgKwfY6i739Lo5AmCcYBXgVcgZ8PoW9FlrLCausmPx31xChtic7Gk2//37zDtHBa
BEUdTMShHjHDb44CmCA+oYeWfRBk32EDkGH26LzZyyCgpw8meW6Dt9NXG1Ccf4XM02FeyEpgBUMA
CPXsamiQvhFMv/Bozqinc8YKoN01UPMfTI+baxJv5pCg0y0TJf0o2LI2aZ2Q+TAz1DZSR5gap6Ll
szUEFiUXH5PJnrEhJT3t7MCyPIsMbotYyAzLWoBCt7xJ7+yl0F4x3ECSMmFqgnJdFN2W8kJRoO7q
0K6CMISm5XlCatLEna9G3C73xRgLxlulr/Eb/6LjaEFCpfcWZUuV9xDKeIH8B+/kFua4/0xVM3xQ
E9CMj8ZB5U1vNJLS4WUKIUcqTu0c11ADI6CN7Z5JSjpAWh6tCzWfG8sSkJIUyiXhUWl7mwMAKzTA
ii7h5jSQ0w6kCZPeB/RoEUxZWAZmnlewM0tMXqUXzIGBnisXSxxMi7zhKe77nxEj02QMjQAxYWTk
7elST/Bc0ja1cb819BjUPul0pSzEdBWMcw+CEEF4jypOQwep2UAZcYi8lL39azEgdKeMsudNfjMF
SvkO65hU9b6DFnMAmg/RpGtiAZ7hbwt+jaBcQFK0N2ZslsvKbBoQk3rSaQRjedzqz4y4UBHRNwg7
H7rHy/dKIdoOnwUY1S7gRgBqTDCEc9Jus+M2BRvn/i6FKF4/KABH+3AApYKs5tDxkZK3BOHcUrsH
xMASanHFyS/uK2KkhyHQmkrlc10ebqtpTP/1BYBEs34LMilYP/bX8yJkT5Jt0AxpqaByTXjTTNC+
3/9S7KATXt0cboJ44mGqgB1fnnoU5MySeQ02idvE/YR2Oqb9f/DxZWxPZXsg2R6y+lQuU/HKQnYl
znXcbKniEUQpcSsEpU1h2AsAdZbzatDO/TYsvPHSb/D3i90uyRnnw6jewDfoJoUxfJUzRwZdzCPJ
Oa8pjtmEf1oAOgHvFeaxHUFBnkUiB7DyZLM4RpzcDwBUf3PQmrWmvKgSbtkX+TMlAfyLFu/QyEo4
lwu3Nf3uBmgNg5NsV/ZhqP4+jIU/I3vrKbVCoT8DirG4PitxGYtu7bxTnqZrgRpo0ucVKnVRALna
2rqJkrN9DZ2qk1rN00cq/kQTNerFCfA2ZruHC/E51MC32p8hSqO2YJPcqrPJ/POI2tgyPrcQY46L
uxq+9oiMdWevdrpeTetPrVCQzfIKbqqwf5+MD6odEEblTPwpmAfo9XH1BDim5LNgiSmcEEvLmAIg
UUZmlo/nMDDNFWSHqRoy2R6pdkFatmwtMMIpcQuxZyMDmnEQnZYFUyGu0gZmTrwxNUBr+yR8yKse
xaB58S5ljIlCDk9+lWUVHRveSBp72sb/sZRzNXo7HL/m9IXpvXxm5NnSvxHUBJg8Y2Ugd7DIN6PH
qGRii+qEBbSm30XGMyNWQwAgQZomAe+rPxyHptmPFtmgcqSmyuniL5SSS6MgFW6Bxudpl5um7FnA
gP1n3rCuzL7G5LavSk4BfIxwllAKrNpRhH87PSccoIIWkPafg2vtHT0s3e5IictZdeFgGIPIyLBS
TQvGJpaPZ0wiCXUruOu52+x1++er0d+We+2i3bQHWZ15phpHFtJm4k0026EBREQT+QqyS8bz6hKm
fAqzwKeN47YKxe1D/TXXUeQyb9cjtlZPnDmRZY9TuIQ7iIHuZnHBoP1mZG8vWQpjyOExDS6IoUeq
PIpzuzMlmRTxfyrEdPgs/ty9UWx7KiA01Cgj+cKGFiS/uWCvKTiZ6L0zBt/6XQ22yDNTK4PIYdNJ
sS7RSf4DuawwuCa2qv5bEudv0RW5wamvXG0h2Nceu2LlCUvfYB6nJO25RI64EqW7CgcjaY2MT1q/
fByb7B1yysi0sZNkY1qIYxYTbufWlBU1OMg/rIypP81U+rWvpH26oI9VodO6733R2HSu5uwOhqmI
FFrq7VRPwtIk9qoM1yPMMNt9wIT3KDnQ7xGaDLOu35WxmDPEkr27WTDfdj5fWVKk0LWakwCEbjfY
CmJ2is+QQQiQBM+xy3g2/U7yf1TfWdVkXo+SZdBPzr0Z7lxEVNt3zOu1ASskdhDVQoZSvFDPtt0z
udgo+OT6czjXbEGgBra4OBy0gIsRqNZNa5QRaux8ZYER52FWm2sQfWnOT+zFxfSX1SbvPLlCaAgL
u1xWLCwcjxYcdFoDhkP5cW+sr0OLGO3K80vVDuh/a3+Aj2FsczY9HFCt94VJl79Cg90IIZnh3YyM
ghxiJemEsDirNfB3vRKA15K8wUMVYQzq2AMzskhfJEkKtYZAfK20Uk8Tn5KGZPiO2QWzM23s1Uhv
mlDtmSj27vL8404uF4tjbkLwMdNE0qlS24lVU0EcHz8ChQmQF/UIrMOzgu0qFtrsme1YCD6nztbF
m65TfqENdRlGObY9ry5dKiGpfrxGaIQQ2DFApuJfvomg/3x3DsGOM/sQ4zfqYfHIgRhySzPTMcke
Did8Vip5oro6z3kBf6dfcIlCZfcx0C+Yyw4GLVmJ85FWYeyS9BbbldjqFjJrJvGecLCXALQEK6/5
VI5wmTzz35MVzy2AsSrsy79k3yH1MJN04OsSbd9TAPjSlVgYUHz+53SzvhlYhBUbieCzwUEbUVuI
CsHqmfGUJotmhTI0JgEcRJl3vydSI2Zs2fBViMq1NTGx3JkMa4G+DsCMQC70xH/dDz2qGskg53Wr
QOCJoC7Yypq8U0Agq/03FIR+31jTiF6dR48tmZetAsSy+grZLwFcXoljurWm+mW6iDYzaQyJtuSr
rWklrQBGFVhY6epIP+1R4Xaa+n8ZwuEjFx+m9nHpPSDnL3t8cq3KcLKZj6RZ7w3reIMFgRRb44WL
T9tosmX+/dgaAnbB2diK//3qsgmbNEkij4QUDvmWAHR0BlC6XPZkPpeGlLNswEs3ylNGLyKCGWKk
aYboO6DGcJGjrFX2ybCrwBotfH+JeKtIqHoY2ZGNI8thAkN90HuAeZKiwoIVnBekV9XiirZRskRi
g2oUroicfSfGx1a2qaafr2oKo3Hf+5pQ2M3I81Eyr/ooJfS9syL3RfvwjhiQ5CNh9/nqJ/jRFYvb
wqbRwhujhgwYGEDQKHtvJFiljSaBbRsKjpW4YmOLvqgKBEDhzfC8gj2b0oIB+MeGtNFyYERvALYx
J7XvCj6miRtqX/IaKVPyR1DHpj3gSZBp/TybDRes3ntfBICwljrSYmnZSVqT4l4j8zrhHhG9fCsf
nYkKPJX+IKXYpxGL5sRYb+qezLn6Qa9AfffkNTPvLqeEQ3eXszFuhqueIcxtXVUj5yb+FmY6uPZb
AVsFwk9MJDRnA3SR40bRe3mEZ8MfWnLqoexxIqbv7SLFMvIcaRLVa6YIbBzaPGszGxb7OtyHQHDD
fwzZDuhSQm5kLsJhlYLXe+YdthNbYTlUMzX+5lDC4QXTmZhRvEk5hSGn9/K07P/61jvTvKbmX5wr
scdn5NDc8oWicHL6IXfoWVhq3EKHvJQsT43+c/1pcRUfztt6XkxNPnfvtNBGj7KusY+nDXkKndVU
MjbpTnVxLGsyH3Pyjl9xDuiFx8iTtLL5k5R+2s4Ba0Irb9uJbkFADIDk0vf+aP2EUBQQStDe0VHT
bt6ERv54R6WJoHYWOlKMHZ/cRqXjWaSdCq7NWGi0WlNQI4ebMhX+IDXugvqsHemxHQLuCtlCAsQU
GUhahYqA1LFBzDUhDwaXWUo9EqG5TAzosBCQRw6kOHAuSsb7zaOY1Qnqzx/G3hEq4Dy9vjpjozyD
neF9X34YSEKxxu7hJCWSG/vgSFw+YzFdQ5EEwwixeRhwpHiIdvKbIaY3lVHEMJjst8VS6v5n1lrl
3MnkRpqKuWvCyGzRGBjdaOJO/Zx+h0M52DceQe3VO8RSBkHpZqTeshsuHxtcA/QV5o/71c/BD0Sg
p9XwL/jf/SkBvuRPvA1gzzpOCYNN8HFIR0Dj5DhxDExiMQPGgFTzgDGw/oui5aS+mpR2qswo2xlb
01ieoWD/Z3GgusBll0oS7/sea3q0R2WE8mb2bAmaiy39tr51sDubJC4apkNBfEq2VN1HpT0vCVf2
+mQRNIsDJXgjmqmESHAmJXPd3/O1N8W4J0sNyQhuci09dOcK+PTbPrr6snQhDkP9SaQ0Oqj23Q+3
gVWiwXsEYx+stOmqV6g8Y9oCyuz2zB/9s4qBiGAccJLMEKc8PZ0r3/DHCazMIMwuF4g0My2TcG2w
U9Sg7wuj1IqsOf935DZETKpyvSK3PVcV2yEgbvZbRl1sub/A31lKR5YHX3EMhfb00W+CBAM0nJgH
uWAWAyvWCxTEyW/OfQqRrZM6ca/MRXceSNUve07nmdawbVFygqpHmaWT8cKM4DI1lJlCVIDaBz8L
UdoO6RzwZUL0e08H17IGFJWl7smS7dpY/b6MWo0BzmkVDCTQjc2GSCnqtCfEPg+uUqTl0faGQv8t
NqqCNkG4Kp+HJEbbaws4Go/x2F0WQ+l+Nwn9kO6mx3RSIJLAG8USUa1MEa+oN8B/51msHtbE+HUh
pilv5UsLSLIkoh24XnpLIfjQi6k4Gsn5kzKURLhMHHzrOxUECXjHl6vKG/pcv+HyeQgoBuLa/tg5
FSfEqi+GxpqXCN3ABefDuUvWYM9nqLvbboDhyqRokySYJm4+ntdKASEwg+Oab8ZoStRguVli+55c
XeI+sWjXGch3JrG4A1g/OLBjOheiNHYdp31SR9a6DZPjoqt0hb5UEnKN4DGlPHmqaoW83pYJ4gWz
obqWFKitiH2nKbyxabTRX+m8EDkWM/JTDr/zZHaTqG8Y3FsSfxGz1bXcv1XD/AXnySAMeYxzL7oV
QDUFZsZjHM0/xeMagGuAoF7HO8jbmkbqnO9l26UVJYaZBfmhQ2sARx2J03zApTM8BlEcYFiqA1H5
2C4wU86enztymPkeewSmEp5gvwAG0DQ2PBql6eDNk3tKMm+O+8viX+2f8+uWFUwvJQUe3qZfdFxC
U8byfz9Jjx0M6PIYMdAGJEz3+5Nlu8Eslt2rR49oo7kpgyG4u9OULdnaWRAhVhaHK0InkhK7x9Rc
xSrLlSiFAG3dp22mTJHE6iPFcpUmYJVYE0mEtY5N9LI4lUfZSbVzGRB+jFFiI78Ob9q1JCL2Rkut
lPbqbMBnWP/jB6dNfMPedRSEAurN7gogAzbLnlbpG+K3jWeTniE+/G4IQIx54gqPoj4kP2+iMy9M
2Hp4NifxpYUkCxgG6Lbf/+4c8zlEsuAF7pQKQMONqzPh2YeOPinCxjYwJxuKE3d6a22S5ccANZeZ
xVJLxG+RyG7iJtNjYezvWqmRpUrlhyeaU88SQ81J0p7z9IHWGGO8FQAuCsdrCW0k2E8V0A49q5S9
Z/pI1BDz9o2FF8J7x8u9ty4mHMSHgLL07iS0TAvnKMBV/wbf01aZzs4WHraFbD2pHPmvGZBdJmT+
5n2EECTvNGMchyYSUb0+spBBgPdNTsS+4pdOYNgDL7pUm47FzOOFenP4JcMxeCmbS/WVL8s/DQp4
GL3ngC3iTCc7GkriGqSDeUSY7V++mOV1Y4hrZoYPmYQZl0GE3Y1TDh3mNDjv+NFOdnL+xnGMCRpT
abcc9vYC3XginDawkKZ69z8qgS76D6YC9+rhQaC99o+cCO6olxg/e1yFNHD2mP99aWu7GDNxOpEY
5YY3xlmqK/Z5nTz1w9mKi/uZlZW7oqnmKUCMKV+q3EGnOCjIuyk5t+7G4f/a+kU6etrPK4WnhpYO
b9hldE7or8i8p3VVBBF5KDrkB4/dtqIemKx0FrHH3sEXLOLGGiLZ4Qy8lL6SbxDtnnbaAcEs57JN
USwCSRIjPpy1ZkgXta6TdSD1bblHvlEBEqDheSnyCncVjuRSmgSC+5U9Uiq81vo0FFIPen1ewDX4
KhKbwHNSwJft53qf51Y/A0OEOJPJ4+RBzkUZNo3xxubavFb3GM81xBavZgTyDJMI9qkIPv4RSAAM
lwlv0l83ggE5hP8v9GPTu1kzwNHDK7W6bF8edEQh/cKPYWeqN2UnIhtdRrPMkUFzpFSAgClib6yF
UmczndACp7BFEgC89B15Zc0KrDP+k1C5VG/PL8ePR5VRgEmL9e01I9aw5c9XFf7SqWsBIchxd/i5
4Vay7vTIc+a1pHaDqPCvFPQM+XKv0fHwXa00+TH3G4JyQjLGPUkGAFhceliN1RQD3FLTCs4ffZzx
Trr9l8ioH7jy7vHCKXNHiRrVAtQE1sxnnfxqLxuH0K1JaXB2IwGMPourUekhw0+AdT+hpQ7RogSE
D3ZIjKKIt6rH+rLKi32ucQeb641pgnxgEGNlpdXorjeCrdgRFBPLH95/GKd+45S10z6cYw8yVmQm
MktFG1dGvFcMwdJv4Hj6J21zHBpsBsxCMQZYE9/nGmaCX3SGMRlJIYqtLuM45oEYqsTR2TFVGrDR
ZmqM10gwMXPzhGQHQCrsfcRYM6fOP1y3ZaTbwTAs9UrnJsRxT020mU76N99gC8n+Vw4/qhZ3hUMr
ShW+mp24KHJqv/Kb214gWKc9TxbLlfwF2dGlxi3If76ADhraQzuNUNLVyzSn1URYQYVnnkJF/Fri
zwcjAHWppZxLHSvTuQk9HH5Sjllu+ynhv8aNN2PjcSwP/nvBOs/NfYQCvN71PuPTdxu59QIxHr3J
Nfttt3qZLJZ4BSAZpFltyjR2120DrzHmIHBpqjFKETRYUwAI3ucJs8GOKAiX5gyNF/MXbqd+9aws
2cA6M3M370IDyFeS3M72e4X4HRTXPY/JvRHS92c6eQKjdSFGv5NqGl/Ewg9+HSxEnmOoRTIoDxYt
o2L1B7IPxaisM8BOGcdoEAP07lSIlNq0MxsCflH2UWqtoEb4Tu0YcT6kH7dKBGs/3KWbsM525D0H
LjaIRL6uPyxfFNPBw8mE4ljevzRixSQVd9uNIJqo3a4URxpVZX7uhyO1V0dgfQb7CcAKkQdfwIom
QmxB4Fzl3j99ZrPoa967MqR6fYmf5pMLWjRi7ZgA/rJZxvyvgobR3F+PN3RfVm/x82eJTPc2QQSH
5e+WS9aa6KUy7+3dO4vCY2ZbHLMoPRyweGzgGzA7js2yxK1k4N6dHe6jraQjZY+9xjzNlvnBHn64
njnVHaEUUVbhfuMp+LmhrpZxKkz314BfHKFdLBx63N1dc8c0R1ve1ZLwquXQqZl4WIJbCqFKrAKH
k6OLlJYtZWkfgTyjW14ouu9W7QmVzSppKTObK/Vof+UVbAoux3v1NSib/FaVGIN7nAyKVJ++aEQM
DGqbll0k80cReu1y3LbozIMkZgXTGuwyhLa7rqdRFU/SNdCM2+JncGsxzLK3ctYfGAPfOqxT/pZA
w8GF5onvEzq2exChuN56pULFQqhbmgKSuZKgUfHlffvXhoNk3RHqlXytqJu0tpt9DmkswGqqZKtV
C1KFnHsn1KyIv3IfiVIfuh0YCgkQ/QWgN+7FZftkbKXOLi7rxTm0dll1JOGlsTbgwSVSHyOQqKam
PQwr39u1OAfl7ia+fESjbo+S+huRgQHx/LhpGp2kBpoa8+F9PPBUeQNI8I5EmfqjnejOQeU0TGA/
VUUo2dmZY0B2lgLjf/f46Bcx+Q96o6U3NH0VYzKO8bpU+XVPvOFUilSmDQJ7Ud58zWdumM1APA9F
H2qmHvAEqLrGwDmgLDOEeF0wibRkwhjm+uH3ToKx/Uuc7ojjSM9My/8+7cxbA6BDUgrx8ND6Tw8Z
5WZ197oUDhUxqrq0UtSfscQTHbmn5ipgUXuXQGwAGsQF0SFG9Crw2KsStbGXSgh/pQqpCWvfieDQ
NVtztFKcB73N1muOmKEH1V5ryUsmTU9uV7Cfn7PqmwFIum9V+1x+Vj4yjsrTVkiZDgGHISNeM0v0
Vr1i5dYsRieO10xeebCttgRy8ish0Gc6SJ7FMBzSRu9pS4CSOgoUI3jPKlB4lEFugRyUiDyNbe+i
1v8t7XJjOEEVz62JmxmuS+7KpSt4kjGjuwsYetJpdcfMpj7lc6jq541dF0/XNtwkryLFr5+2gaVw
UeFtQfR6bqfqdfE/Vynpl0W4J8HClNtnYQNks+99bgcqd6XfGzwINSF1hLlSnl4HzgSf/p6+Fi8U
dzCj52qYjyLZPfYNFRHR9PrycziIYQPphzvo5OuuBgS3/daTqWJwNfjeeDRtjcpTZ8G1LrNLQHQO
yYJjHc3qIJmwSSFnZ6jYpvE0ytjS4v1v5m+vFltgkdqvK/2lCnZ7XM/kIu8AThVUGwBMPc2xM47t
svZbPH+OzzEb4VTdG0ylJJ3vMBileWs6/YFHJdR/LeXYn0+yoGzQZTF9qPb1bq85fWHUeC7gjXN+
alp4lcZ88ii82eB7HlJ22AncvAwT7fa1h90kwetAfgjy/Q+0OHE2rwIjaLmmuvxVMAWxq7XhdM8U
HqXhWrSKoFOTBYxaqjnCrkdzKZs6CocBBLDouIxapG+6t+A/L6FNUn1ThitDOXJ8PlkhJyZyuuVc
Q1YfuBZgGBzkVI/K8t/g5eno2b/v952JutktbHvf+l7/agf80/BC9T6XBOXvmf64lmpZcI3fzy9Z
JuetnY9C8jBY7SK0cg8VX356uPGxrwyXM/HbnfZptXHCpdnarD7giXQoAYl3UMXPIvsKvJcgPbGS
j1GZ3PorkEhI/39owXq6S+KMriOOxiHwseSHehnW5lO51wpu8zYf6784Z1AozOa9LS5KJ5u/dyDV
xq+w64kjYMIyho+tra5lF4CVWfG63GBhw7NBYnD3HSlqDKUbJc2LR08aItlWTdVY6wwL68nliDfS
vyBQyUgfb9Dg6lfdG6q7mpYN1vL8KQAhRBmY1U/9xXwhUCq80EZBKyKph0Kiy2VoKDdTI97nMdej
nsND68Y5oQH8bMQ2NjgSbQGts9EtXMWImgidb6vpy+AqCaNXRSMxUwI+njZa3xLm2C/YNhezfz+5
qFeoSOhjz3JE3lNNL7nk6oiYgn1nGG2ZUqXsbPhLKAw1ViON76ZAOGGxhIG8jdIpim7T2spMHxxY
A+9MLNojjbHE5/0WrLphL8p9uKQ8nnHDBq9HUY1GjBA6C6yhAUdaG+Tsv9FuZ5CEmNXfzmHS2tYB
9Npjuz9M4zr9HiJWwyiq0o/CwoUT+ya4Jl2ljdzBYPMjXFQqv6g/bw2lglpeUm7DXR77EUb2ajg5
ZvcZHFr4RkmHuaLT5AIMTsIXDoJP1U14pKIy6/Ozzvc82OU8EjyOXsQxrcVJjc5n4hJ/PzSzFWK+
f2s915OGn3PrHb3qIao+kcScX5Uu18L5ALBzmlL/t1qX4DqAYg8ZwfVKpAH9hO+aDrmO8da9c5WA
56jlCJPwEJqq5baim+nNChE8QaFZhma+0/CZwgaVt4U/y4g=
`protect end_protected
