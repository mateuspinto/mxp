XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��tT^%��\wdX	�P�a��<[�,�2�ށ݂S��ך�Io�S)�S��nZ���2����(��J=��|w<
UsO�f�'�fjK��a�F
�Yl$�i��D�E7�H�{��P��*ܑ�I�f�{>�@�c �K䕖�O�`�/�m N��9����s�F�b��)x��nbr�k�MXva,2N2������;�X����!�&��P�s�����?���vUfp>����]��	�,f/�T%kѮR�,��h�E���4Eduzo����$�6�CPz�	�j�l�<~<�)�����R����j̹馧��}�sm6G�%���ӫf?�K�C�ӑ�2�AX�2K�H>����+���k�5>n�Y.��Y�	I	�""��uC>���γ78��\y� �SS���D���d�ߙ��٦/JR�}
�C=d7��I�p�ţ����^x���\�\���a�T�-s�\���E��7<~��?�\ԭ�L�L��o�^����hzT�-�6����;�S�B���\M����B�	�i����,�c)k���"�xTs���[7f�&�z�H��ї�^B��1-������7���(.[h�X��c�zw�v �K�2q�e�[9>y=�;p�$�g�b�j��{���
LK1��C2��kLsDq�ս�U=�	�vM�π��$6W:T��⢦��W�}-��I��4( ��~�'���C��̿�e���§�V��Z�/��G,�=�E�mK�.<3TT!XlxVHYEB     400     190t��J*v�4~���K��l
m5GCn)8p�Mַ��<��<s�vu�����>�M�_�87��V��ĥ�}f�j�J����ُ.	я��M���d �В"�VŇ?b��A�I%$��3)8s�o,���c���T]J?��?�la`v�<,;2?.3�J��:�).��F�X�_�^ZB�����v���i���� f��.�$��2��F�-R�T����2�Y����AP�eHK��$�5sB� Z�� ���3���{���}F4���T��������w_;����V���;|SWBw�&�~�x��Έ��]��9T�Z}Ϧ�I�d�&_�����y Sv�:or�k��9��x��gt,�����>�`�1n�;&2�>-�����P�pj���XlxVHYEB     400      b0��Қ�ٞ,fl�n��
L�.܂�K�q�r���64��kk�˜�Qs@��qr�:��|2�Ԗ~�m�u}b�r{rӉ?:1��T��T�T�����]���(���0��~�B6�P!����`�X�W'�w�L�{���ִ�Aַ/=�}��F�O�Ϛ��.os�����ȒrXlxVHYEB     400      f0��|�.�R�Ė ��KX�͵ؔ_���;F0�Px�/|�?��'�9*�CD����
I	����_�X�Sw	< gI��-�ݝ���z��oܢ�G�EA�4~���6iՆ�W~�`�s�Wx%q���A� �©�|�8\�bG��V�MR��T<�X�
bV*�9���T7�4$:�_��xM�W���5��Rm@4�MR2 5�.�h�M��.��k>���4�]>��+Q���@z�]LL]zXlxVHYEB     400     150����h>��)�0\jcR���͎�6��4��i�����9�wǒ��A���
�^�{�D�|Rc��m*�h�kc���|��ء[���Ox��,lb��Ҟ�{�8��l�^��=�@�Qh�_|�9g�t���b�Ys���A$�Ѹmⶨ*b�g�~�kÂ8���eynS�9=4^��Ҟi�X�F�۹�0���n���<�� �r2HL�/�Ъy,��(���%e:��M��[,�4�tW[q�P�$w�0��뇊mͥ5��\Z��X|]����k��[��=2|��\+n���yy��ɨWU�FEi|H3��S��5(f�XlxVHYEB     400     160�p�}�yi#�z�ո��b�u*��1�@���I}�x數��j&	;��ݏRJv?�c�EVj+$D~�%���fp.?'�g�u�kkm��J�B�q �o�qa��3u��N�_j槬N$��o�D�w5�Q9�j}�M9�'�G ��tW��L ��e�L�ˎ �i��7�x���k-H|�� ���S-s�aj�y^~ߔ]�І�&(O�s����S*h�X�~Y�Q(f>��g���ۍ0���Z���FG5?R�#��ƫ�����Q.�]�A�R(g9�EM1�]0�H!����ہa�l~"j�	٪Y��:羯7����]��/�̅�{�yI~�XlxVHYEB     400     120Z�H	����8��[�L���iK�v��02��0�Y��l��T5sd�ԛu��Z\b��.����tb
>t�;��+�d�;�hr41kkU/�{�����Z%b'��r���.@G_0��4u'�����\�sGLl阹筱�~���Ę��tdA�r8���h/�B	�CK��l��P��ϘR&�bʕG��f5jE!ݧ��թ����!���}،`��ƽ�<@�Z��F?(�-��"O6AP��t��c/ᥗ�X�c���]��l�:�ן+,al2�;�n��HbXlxVHYEB     400     110�t�����|���G��-!����Fi��?4[��$��Iֲ̻�D�=����z���j�V���1���d�I!����U����+N�ma�ml[��"� #� �5��q�˕2�����CG%3��P?�Sچ��/hֲ�>=� ycxD�w����v�w����n�l��g�#���b^u<	���rC��ѬšF嘥0eqQ!T>���� ��q'�V��>;\�\RlP"�WZ��0H���n��܅��JGff+&��H�s��;��h�z��XlxVHYEB     400     110P6�������wZK�͚�'z��$'�	���h��z@���T�������L]W��k 0T�T5X�5��x�a����ȡ�{n:��SSj����.��\tpЁ{�BeA����� S�9]v��$��`� sJN���3o-�!����wA��B n!�����|�{��o���y8f���I�EaLX	h<��$]�m
��Y���[�3����]�����$O�Q�,{W�#���v1}]���]�>����L���y�i�mH�
XlxVHYEB     400     130�E��*��}Hf*�^����{�fR0QМ�WTn�AB*-�{r�{/���ߐ��4$����`Bc��:�)\����6��@Ix�"�MӲ��l�dΆ�C�YB��ݯ�NL���VTkkh�/B�c;���s��C�ߑ,N�����G�x�ofvG0-��D_N�&!�A�b�0�w�J!*:P��/0�"3��EZ7� ���s���~���'����^Qm��x�?0p��yF���PuC����
=O�K8���X5h%�oH!A�m}7��j�mHjgm��F�����ꒆL��~ɛXlxVHYEB     400     140ދaD��RQ=Y;a�%q�,��%y��

K��s��}:���)"����6��&SS]:�Y��jxL��~��T����w]�^�8�4_�Y�A25t*�
dH����'b��J/�E��^�s���e�f�w�7�$�Z:֐�hc�L�#N+l���$Pͧ��{�jL�&+-��P�k��������*Q0���'��O�/,���ԇ1#�J�L�_���p�[&;�ʛ������O�Ƴ���N!�A��ŕ���T]�`(/N �4�����h�q9�>;CMoJ/��8Ag�9T�$귅MQ�N�8y� FXlxVHYEB     400     100wEa�.�Yy��9���3#)�Xgb9�}��k�1�D�\P	^a�y_��y���3�7��>�ճm�ŏD��j<[�p���̲��r,Tۋ����6T�������k�|p<��e-��q�1���Ķ�3���'?�e���2}���7�-��tӃZ 3I�GJ��]�N��R����g�=�{��������rj��p�(d$}ͮ|+��&���Z�%��%A��u�r�9�� C���c"C�z:ϢK������<�#0�XlxVHYEB     37b     140/�iXi���E�Ͼ�o1N��sy�;���7B+�W�]-&m�A��G2|�Z[z*�9��T��1nO��t>�{�,����hZ̯'�p��.z:G�a�`*��J����F����vs�����E�ǳ>��T���ʐE0+y\��0[M4@lMNW�m.�b�h��U`f6��Ԯck7
H��oFS(1�De5���i�j�t�P��.M��$�w�U@I}��9�ä��oq��R��rI[��	з����5�ok��L�x�j����I��\�Arנl�6���-w�/r���0_�����b��ʽR4��P���$���