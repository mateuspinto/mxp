XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&~�oQ-H�N��x~X{��όī��T�1�L�2���j=�y�w�x�M��	5���/�h7S�%�x���x�U�!�ǳ�!7���N��VS��R�p����z~}�rW��9��dzl�8/<����n³t�x����&G6��3NHBi��36�kz-> `LPt�SAW���o*(`�]��0���}����>O�=��{댉��H>t����t���Hq�ZڟuSk�ZϬ�|.�'Rrt�S�����*6��L��T��a�
l����������\bsn߱X�v��	5�ғ�}�G��]#�zWBq�E>R�w�L	
s]~IGǡQM��� $-�7���/���d_�،��L�_V�~Q�E�:8�T��k] U6A_ƙ�vM	G�i�y!�8W�-zx��
��_��N�!=r�d	��\����g���c'���e Uy�>i���,hk5����Vj�w{�u��3b�u�9����4,���ҁ�C�:�D+��g�PYMkQ�B
4�p�*������P�,7�ه$��g�q,T�.5�m��x�"��qZ9�!�Q%��o��P�q���N����P�[e�\L�1���u'�p0Zw�Ā	�� 0����߲Vٻ�b�Z0�4�Ө�d�A�,�%`�olfx
�y��L{=��`�*3��} ��c��׻���B1o�/�|p���ˣ���q3��ߴ/���ohQ���/χ��9s6��:������#.���*���H������V�>XlxVHYEB     400     210&n&��,@�U��j�@�g�� ���_�|O�:W�ݓUs~�?j�ڋb�؎_l�V	���X�&�䒾-�ר�v�&�������=�,Q`�cs2t��{;��������H.+��+����=�����&��/�]�ߠ�D���κ���hz3�֋��S��4@Y��\ZQS)�)^�d0�!��Ƭ�Q���8�Րm˷2�/C�ؙ��<ʀ�=��K������62hJ��o���z2$�U���8=���_+�-_�E4M����8
5��۴$&v�~� ��s	�0ݩ��߸JQ3=�ts���7n���MF��U�+���$]���ߞy�A�9ux�8�����Zd=Z��ӷ	aˠy��XI��yW)��Ս���_�L��6�k_�{+,Z�B1iNK's|hHC{�M�����֔�G��~�|r�1��y]�;u/z���1���\�-��޴��#��1�Wl��Ǿ�@�<�M0*qm޴�S��7�Vdw-^k֓��\Da'�ʁ�XlxVHYEB     400     100�kc��F�؎��]�-��Ii�1��{�����Zv��Z2z�?N��O/9ema3�	#�l��
��q�8���aJ���fd�R���K�_(5WH�lN��4��������� ��E�w��犄��)����'F������j��N���NTT
�0��8@V���:٫�_�ed��� G<c����� �z�_
�˳9�VMu��E�S��A}�<��(���̗q��<츕��f�AnG\�&��(�XlxVHYEB     400     1f0=���0T�cE�6�Y��%����kC����d�ϛ��9L���d�{�VERS&�����$� ��@k�q�z���pX�^C闱�J��0��:ҩ�e��-[�����ht��Nб�ms����o�_�I����1I^��ڦ����|u�xJ}2�N���сCd#�5ۂ7�L���kB��y�*Zq����?���@��~��Dq#8n��LX.%:'E!g$��ص�b)���U-9�8+��-˼%�J����b�*��sN�"+��'�[xfp�i�����aS"j ޸-���w�	۸*�k�d���Q0Q-{��|�6�+;_P��U�n�.���;�K��]���3d�������/l��w�s�F��x#{�������=�ž�iϻ� ����L�GƮ
Kp�LW#ʿ�y}��Iϒa@�kHj"B�a�E��IЋ�L]D����"���c=�A\Q;���(9�������>N��WyXlxVHYEB     400     230K�+�t���;`q5w�7S�Sz�-�_y'�'�
_�B�q�{ѐmI�>�$>�&Q��/^;�Lu�9��<�nwĊ����Ԧ-G#\rf_�(�\��y9ʷ��+�z�r��Wh� �sdOR�,O�y0�^G������t�Ga�_D�i�4ǐ���g~�"�/�vm���?�}�V���X����P�N	z324:�<�d`��ţ7�x� ����� u�xv\U���!au�3�������T��?�a=��P����WRM��5�p��?�NUն���j��5���{x��r���g�3;�����������(O��Y�p�:��`����u�
rG�Bն�>Vυ�%�����݊5BwO�x��z�DË�}���B4��x��Z�?` �����F�'+Q�{��}VʧD�2E^>��}9M�u�ީ�<�[k;^+���өj���(�a®|
eRW (��)?.�,C����,#��{����$O�}�-ؓ��}�W ���0A�1lr���:��s�⤏\]2��� �{F�f��r�XlxVHYEB     400     1a0�^��cy�w�Cu��I��Eg�Ͼa��y�����'��=�,�&��j}s`D	/�p_�����F�=?K��>/��l�Q�K��<��^!����M%X�CN���.��H.�>*��d������� �&Y�q@ٍ�B5A#a$��rb5h<%V����/�'�܋ v����u/-�a��û,���`J�L
���M��BuƨU�	;AnK��C4'��:��|�?�ࣁ$����	�hqf(Y�~��p!@?���Ѳ����y��g�$3�5�6
�k�M�HJ=K��A@@�(�ُ[t`��6]����~w+S�tN&Y�wʆW������'��jN<��+!*S�N���J�{���"O{��@ϊ���Ph.�����JY�F���@c"^�XlxVHYEB     400     1a0f��9vV������d A���UI����x#�m�% A����UNe���)�E�4)�3��aS��"�Q���ƪ;�]I}�f:���s�����}E���P-�I��D�+?=_t�&�\�^jF��w��j�S-��{�7`@Z-#�T�1՗lQ7�Eߔ�JA��L�����<%��-�>�b!+�mk7��,9�x�+G��;N���(O�����	ϱ1��ج����se�-��^���!E�o�[��<{��_�7��n}�J��*��HKh�p>��{A1�vS�HW��Ʒr�x�&
W�g�w���Y@�nCk�~��-ϙ-;ݐ�;��=&��+��~��$'�+�T��(=0X����{WQ/�\�!�؅�][�z�^�#)т۷it��4D�ď���L�pl�XlxVHYEB     400     1d0�m��嗃�;�#3��KFo�$�I�ȫ��/H-�`�Jm)��"��܆�������!�T��Q�I��k݃�ZWU�Su�H:wQ?��[�	0_쬊�}o����qS��ʼh���z���|�Z���w�MU�I��P�uH7G&u G�E.�?��iUc[ԇ�bc��E�KM#�����狨���Z�BW�fK��'�$�u!P��y��h8tQyVnLsM�1a5O���w������w5Z���f�FO��E�D���P(o	`���HZ5��X�����Rk��G� ������ltLe?d�ƶ���֪8 qؓ0G���r7�h+�Lv-��ZL�2�*���N�5��Y����(s\7r�!+�\:ҏI�s��tB�Ċ�mR#$<���_�{x�7T�%�1�}f~ц&��Hډ�=�HU&'�y�E���P����1�Qc�4�����tXlxVHYEB     400     170eg�@��	�G���f
�%��{�W��ľގ�(*O�{
���w��QٗM�>�1lv���A�.xzߏwP��:J�);��K�>mB��l��%���bU69�1�l���eJ�'��c&[=v�0=쥺(���s��[93f���O��)V��O[J�b*m����0;���ٽ�0u
�e�͹�eG'rj��y���;n��F�P��X���R9�96��(tX8q4D}0���6_I����y� {EY6�ȟ�B���Y/ʪ	�Z��8&�5ru3����1{�!6�����H��]Fcw�,QB��USe���Z���o�]6��4W|��M���?&+u������ob�bH�=�����$XlxVHYEB     400     1c0��<��dD��H�a�7B7:����
x���| >����N�(���N�4&���(J��3[I�M�2��eq
���}g�C�?	3������X�@��1$4��:K�S	�y�����q�"����t!eM��%K|�b��Fr!�6�� ߈���� �K&z�"�:wG�n�d�jCQ��N	
�����xx�b1�.@ĆiP"3�O*ƣ��te\.B���U#oZ��`�PF�@��vJu9��f�hE�W��Xt'������U���2���?�Bט��_(5���R�E/�?�!w�� �~[|����y�-���n���#����
�C��F�'�ĕ�mYץ�<���f����}���he��9���߶�8	�)��%7A���"�����z*Zʍ֟N�����!탥�^���fאu8l~8�p��]׾.C����XlxVHYEB     400     1a0�h�J)�^�?g�638X��z%q�s���#��p��i��w\v�_���0��/��E���e=p%�78�ٲa�zç��8�*+��= ����mt�B�L�.On����"�@s ���Z�]����.T�u�&��yHl�((��{���&9ѝ7�3Bh+f��[E �;CR&�Eu�W����=ߝ�Ht����"�
0�N������U-�+�����C\��cth8�oGY�=�B�$�s�q*�t��"!O�?��kЩ�`8�K��w媔����_$a>~�=pB*ī�`(�-Ƹ�B2s?rF(9J/X�ʠ9*���b�NZ�.l�4�)����wf �>����m�X.�
�>�%��V��4^~y��^�?u�zt��HU�_G��U��Gy^<�;:=�3	G7�B��tӨ�=�Jl�I]XlxVHYEB     400     140PM�_�un��� �����ɀ���q��	�n��F�5a���])�h)(8�O)��SWy�[���	�aZA�9ECo����G������7rIK�]�6�O��}�Fh�7J�~nR��KP����Oe$`�]#J��Y��uC5C�y$��R������Z�����,|���+���y��
��GM&:��$���k��l/p�,r��Q��/FG�{&�;kSF=VT[` j,��ʌZ�u>�q���n=�:bQn��l \E���B�-�F��]��ѵd(L��Y��:�z�v���b2����g��lu�gJζ������XlxVHYEB     38a     1805jW�w>*	}c>\>�N��$������Z��c��8���������'Ù.��X)����}NJ�?��VY��|a+`]Hca�q��T@O3�[�?���h3����o=TĞ�b�9V�2!�J|�r��W�/���I��Z981��Q�$��j�t��l�PO�]�.J�߭�DV̊ɪ��撽�����]N�%F��%�V��?�Eh���R}Wo7�T���f��������ʒ!t�G�������ޓ3@X8T��r;:�ow �,�����C��E �[3[��	�W�L���~��RlK��7cۭQ�}�Lq�_�ə~d�m3��v}��Lݗ�	%%S��O��LO���mr^��Ѐ'D���Uc���J!��