`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
FJ+MfRF/7LmZLhsrL+VRv3msCr3BlLCzTk+idxKs5HscZSlENsPaLdSA2GAxeO2y/UxMlSjt9wfq
X9tJWVplaRkzJ5WdT332IS96Ap4EJH54RBXPY/ddPPyBNsvQsZ8fHcS+9XdNEyXA+zQBKVWNDo34
YF5cJwtkrYrDz0IJmTyUkuYctgd1B9MTGnwA0DVJb479HYE2kPhP0rlofnviN03d/6drMQGhkcHK
iuaAaD2vRB9n4y+dahdUztwP48ULB2KalLoNDS3mg4hUBcAK/oShNGSEjY6qT6j0Oqwg7iKtNMJb
Z431x4Kjnf56925Z4g8P0K8uK+vTp7QZVJPdjQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="EqwN7j5lZoGWxUK+PqOMH/m4Wz6mHEppElRWSlFYV0E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 76976)
`protect data_block
abPUJ+zohSGIcOqZYzMvK584xxcQGE//INNZGIU5sFMYJclyMtlxau4wWJOCThOHJ4PSCtssWokY
KYVVqaQt2ijbyWeaplhN+Ku7I2pwu4yCQxy1VXDxpHdLv+b6LvZcJ9ICzWd0HsuTZRke5x9SNLgi
Fwm2hgYkytsb8zaZoaIB/dSPOSz8g8oTDR+t8cWZyp0zpndmH+mYmH7rl+AaXZKy+jet/B+MBXi3
rZjiGMBbyj+LY0BW1YZAqABnvhkoXRsM7rKvqs3L2Y0rK5ROz5QCR5jsWYjcWjJMT/AV0g++uSSa
WlcxJ5GO7g2DgXmiCbbvRRuxgr/AdMAm2taxwDwj9Fty6hwco7C+7LO39fugedGXEjoSXEldu0xq
J2hhEp8UILeHYLceSJQGgYwoB1V/wWVaeTTznKypFn05XrGlTGr7212MaNQwKCb3KX5ZCObUarDe
Dnk1Bz3Dgndb+yPLHFeAVeHvz5B/B6Mr/9gSQA4UyzoVXBLELyvaQaL5o4V0RZRk4ytBkbxgByq0
9IPqaxVUPrR52tatigVRNP+Zh+VeAqX4bygzOij5PjozqBOMV/oMfnxpQyF+/Q8fLsNItEjCABBw
2Npicb0EZD42n7OgFOmKFCKj+tZZR1ic8peaqV7Mr/8F8kOvZ7EOcyPMkQUuie4pQWzEzNVNevyC
AUcd49n/xQTzQEfF8LXcy0gZibFbwN+BU6Nuu1nLx17vDLplLn4jR4k34t+8RxRCgkSYno8BXNdH
2SgGFHqoTbwmoauwvTkx6XPdWBXR5hbI69HGQtNiFMY/I0ikfz9OwLwdyoW4RLY4vmDKKyBQONS9
7Qh4NBH+EgJ/dtS/mA+TTw2w8DJOIu3Y0KXhHVT+S0feco2uGCUciRpQ6zzG/f/aikP4L0e7j+eh
IesHwkZRQtyF71ddQJeYc3hHYnNXSf/UCXMw7AoTb9h79JzqyxeLVEG6sJUiUpKyyhc5/kPRLxFK
XNryEBZ1vZ0KuwnXAR0lddBiVM/3Y6UiZ+z8U5/BpOiS2qtMJpbU/83wW3f1eTF5FM8zPJ0ptiEF
dQrW1qfKVhNx4o5eeAV99WAj/bjys5sJHt/cZqhhMuD20WlFNJ9Xl+VjuydvSWon2++HLqxlkhIE
TQ7at/yMWZA5K3TSdZy4pU5KZVQeXPiXj5cIGI6N70CBKsE0PlrFEsIjzO+rItVbTkShDHT1vBY6
SRpFnlsZbchciQUnZhFl3iHh+WN3ZjWjVXWbc0VHfDkOPgHgtU2tsrxulWy0WK0LZJiYU8hlWvqU
lLXEYYHfFE6ytPKIrJWeDakyGNQ2A9KLlioB0NMuEwQ3/aRrZH4wTynfPga2n9suCdfzQqydeCjn
6uZkVhSbg0BiUIW0IOF8suXxvCN1ZlKEdR/o6SYDNMfrE1sOXP8doZxg3DJKEZmYqNEW2IWojCrR
R3O+LiRfqzRCbKTF+yM9K0wVZCA/VaHdaDoK6/Q2/7+qjyKKf5eyuo4Zti1FWM+HjCU8iKzRBn+J
6NFbVVU/boy8cUvB8JJkgSBMW8UTiDw+4qWLh63aD+ehl+7CtR6CoWtLlrcBv2nVD3WdcyFfNhln
+rC83JDDwwlSIHA5Lec5oh8TDysaIFZ6xEKmbkIIweKz8VOGH7wWNdHPnlJ0aZxj3ptpjod1rI85
CaedmOOcMZN7fvMLmVU3EdzrX+I5E6H5850zKyZ6gEdMCU5+AE4HGIIfuZW49zSi+KxBWH0tMUX+
3Vq2PgvGRExeNEpURpj47Oiu6sXJ2rxIhJPxdfiDPc0bycDBvnde8p9zZovtBhstt6anzR0dI6EG
K/vIDtsobBvcF4BlKEdm5A4Aj0fhLKDBjvtxWuB/knYD6VN5t/SqjtgvLLecOUpuTONyk9mtqh94
MCEMNaMgGMsRTzeTs9nq8gpw3euHPRmnszgaOi9cfq5UhwH5IQFqzOk49KQdJnbSB8vdoEZ2DgvF
ITkro1kPA3H7g1wyQoAZKAGnbWqjF4SL4Xb8J+RICtjD26oimlxLmrwU3Ws3UBhcDO8A4ADMzheZ
NvTgC7pr3MPRXlEY22PhKis3DXOUXBbGkN+B6RGnDHX7ikK5IfjmCI0+zH0PwH5G44iRhzBfCGOz
+kjH1xDbLCt1a15osnuGvGH07ZDjlwE3Xkiecddl+HeFbaQCSObJkSdrjnZAWwRuP83M8AVjVFhw
ibXAbj31MhGZ+4g65r96Ois4rPn5OCLCh/9L4p3U1usr11XbpJafcRlYbb6JtboGqDianK3pinyb
9tHALvt0a3Y3mCBPbnugcxtTJO4IL1yGU8HYMvcYNmrnc/zEgdnY8luDNHeKD7o7Hz2OvNlKkZUP
we/B0cIAX6butGTU32qy7zcfIKAy7KJ6j/OxOpAy+DaUkmlItsLSfeOWJgdWYu6zqpxMjLNsI1WP
tGAesEpTAZrtsUmWVFFjOAG8yVCpz1oR1NWM3NMYXC95GHi5LPZHg4F5sExtq5k0QeR472CwWbUz
Zq/2w1ffoAGq13GOEwMUp9oV9mDxpe/u6Zj55gggGFlP5b/PKQQb45VmqLZyxo5/DKWndHJk1+aZ
t0mf84bO8N/1KiZE1I6sOWYxc4gN3iCnuGFrcvzRNBiH0HB/GPkh6EjVLpY5P4pRDQnqKp4kIYnX
8eAiDucf/Di4yMVRShf5WrvJcErECmtRWiwfE9rfaxKJ9IwMIJVhLHsnuafy0l9sFsGnB7cjY70x
tf0CUa6kmMVdWqFGMc6eVObNoqAlsJfohj8wELILz3uPtELyY14CuxH4RxC1tMAsjkmF3hkd7+dp
cMrdMo4wZzBuY+970MNslTMl7hGmRs+YcqBEqq1f22z9iCxijOwihxZUaCpXxpQ/k12MceP7frHA
oBb/zG64HeVBEGx3C/3zprxK/LVbPaAvpSna9hwFYg3ArxLDfGSQB+MXslQky40Hqc9V0ZI860Tr
tzpI15M0gtyUinpYzQszTquOuoIz9nyPJ2shlOTbs+enfRwixpqoUtsbYrrHzuDYL6iSrUbkv4fV
f0DMTCNV+829m81vPrO/OviYfiIJS+Wd5vej7lcrSPyazysPCcbqy2ZB20cOFJvkKKHRdEk3K3Le
0cavgEqb4YiLuk8VB2HO0pmINwG9rFUlMiTlEXmhcTpO8O9pvOMrPJX67kkqP7rfaOpxY5thkTEj
IfEq/ySIy0hGniCqpIkQDY3fZKyzYOCrq8h5rJIjhHkPgjNueK/9jpi6i0ryT7so4qNs5nzC3+FO
38238fVC05NgoICmy2U8CWxE06u1hYoNVr0/7KscEra4YVP6xcfUmKNXl3dRB9j3jJRee6T0IR0d
2r5JOWzPhJL6EsClLNUB5sOIC+eegWfv1cIgAtQySi58x0O7FSjDnRAFXVATseTCpm4uPnSiMwxK
nd6j4xBMMFQuI/gjS+2pwj7JWOSznOAABVsdzpKapgWJcSKdpvNV9/3f3AnvZQQRSKIm9oe2D+w5
moKnq++FKmQ2I5wO/Gkv3Y8O6a/luygrEmBMApj3UuQ4dgrZzzNEiWb3rHRSPE2cNsXn44oPl8bl
ciBkA3crsMTwRIDEvZKOXYNa+yGVPG6CV+xY12UdzHEJBPqx+46hy0SaaP8atXqq2r2pNqxBSJ4h
Rg63rc/mueEI8nkZ7PJQDtK2aCJ6DGXYwD8pgMUM56V2krt9c4CZ3Ia+tg+25+qQ5kOtpNndUCh3
Iv4Doe+S8JHjrLlMMfS//50AY6/wQLS0fJPMXD3bHYWL6FYe5ZRdbmCmKxJ0Mh4jRpnnz/UWAzJr
zzmqG/2r/xrrsRgNBOHNadVCy1uRbj4jGEtxhicIdtHSI7/yFaCLMfwOACB3VdtaBWw3iR50/bQx
TCEgVFYIGYtoYtDw8iMfUGqt5nOBVNcM/EjtoGCKHfIkRYC6qK3Sjc1jl13h7J94e/yXWujlmAe5
02GHcnrhU7l5iahhBTdKUb+Wo4czkniXpoZrK+CsFWZBxK38qv5jFSsqNKTyzvVqBUTrBR1xpoS4
xGEp0rGQKOk9Ku8kQaD/U+Mywo23fGd1FQ2fOC+2S4AsI1UiV30byi744dNFcyVrn/YBAvyMeg1l
jZV5TDaRE9L70vf42M1+Aha2NhCunEx2KAEMypRq0Nbt0isVaQQWCt4Wiv1ivHT7d4H/kT0ojsBl
azNsK4XQKa8S2TyWFnLpsbOhNlXbZBi7TyXB6ZpE0D0WJ5jiM+HblP4FxPo5QYaje+xwLcsHfcnl
kt7EYJJPq7SuggZD1hZMUQR6vG0vz3PE9JDYxGtJm+XwxmSbJltoIGmf7F0pWsud9NBT60DhUmO7
yLYqthEaHhDBT+tuqiucK2lKERgo9Z5Qc+FNXi/CkSUuXAzozYWZwmD5Z52F4VPLRgNR4RwDhiou
4ZyBA//LJmxprnTHTlS35U0ky1nKEF91Pp/rtlfIlo3zBsctuImxdwGipBrjMGZc06QS7LXRkL2H
lJ6vCc0UcUObOYze4s3W4cdIyFbaS1BIy+/1Zc5JbHrVsc3P88DmOKFSdnKQCfHyvPd1CFHkrCWZ
QTauyVioVIQCvJ9GcgayHr1OzQqgp8A2DGUQE4VHeNJnNigDChov/KhZA5BEOvs4URAMZeZvslYT
r2ilV9TQmsztAK6j9O+z1t138sQvQdtrPSiDhDDYJxKWgU7v84j5PzUKwXA4lhhOUIwxhTkhPcwa
94ou4boOISHovRqB/Ycz64bCK5NOJuhNCyTd5mzN4GCDy6TgULugvWT7qireGhpSRpzTAabECqs8
tt+d1EUrF1OHcNGoD2cptftpJqEGF6Uuo68Xl2jPU+5vBYg3Bcr72jrZkXaU2yn4IlG3X0wvrzlJ
dTgIcAve+vHaTeTzqoiDo8+wGTixf8SwyIoAfU4ccgVT70U5BJPfPABZXff9sKk8FqjBbT7Agaet
brt2O6HzPqKQrEYZzQxhkk4ncffdGqcrJnQ7WruMXbvmt+NZiM836z97NVdeXrAR6AaJyxdMzb6S
DcfdNABOIgcH9cCQZgESfFq54s1Hl+D2XFO02I+m/nU3obBhJCNFuTR0qwHQltGyUDQffnCAKPWa
xbtM6Hju86E7ZQplJsNnDmsZCIxcUYfvjP1rGOOKMZJiHJw0iYyI+AmRDFCvwe0+4Uv/uzyy/ZPO
c+1zzfiE0R2U2L7y5ND43qCykCbUEE/3DJSVt8gNNtjYs6Uk0BQDIYHLce0Mm41dFOd8ukCt33H6
s3fuQ71hn5F0hQP/823GQshFtuxhoTqzwkFKFg8K8S06ONiB9j4g37txCHeBfv29GsrrZMRJtrT1
646IRlWKaPU5oePRJ9g2f9bRU2pL1MULmDb6yezQDfPpUTw4+7YME37nX8FjTUKDUxdUE1O/LQeU
4lKRB8M+ZFICdzfrpyaxPmocC16so4a3P74MuUNdc47jz3kgfCby8yUV41y3S3pvw0+J2KePMD3t
6fx/6YpoyhulZYQshPEitwqm07M+Ln5jpYRUQNEXsZI6/vaXvSMyLtYQLUOnBxDQdNqFQY8A5EEp
OtaDEbTRbaHemEArvhM2+xlCtgYUuDNR+wjjpZpyTcguEOq1nz0F0FO5vJiGSBAkrlxNU5+RXXtG
vxjfADFSJ2QAU+ptsxNZEzuvPk4RzbVgjXyC8vNaIoSUJeLM/Lm9Mne0MYBnEr/jbb7nPbgVhm6E
2oorfrNbX5FC7FVchYFf2X+65xbf5JeQOb6CglKDj+S4HKEfBRqwN4IjwiOCGk6vmfO7sJtOqq0w
zh9d5jX1OYUed5xizgw/KKbwHzHYtzp3pujorCsnQS4MSSa21nK7SgulDp4V3swKDNCGbRmM8Hq+
u+B9OiFFAfQIrcGS1nz5zPdrN7C86Ej7SBi4WAtdSWteUFjxxdKr6QYHfVIPsK1is+ofpKNu3SSP
A73mbyUJwxLZooHk0LrPzJdabD5Fjegu7JkYPYU67ngSEFFH3m8BY8F4Bi3AzahLzWG5QQUARCk0
RjxYgSdoGPWLOCP3BMTFHQ9tSjZ/8d62KSRIvyl2EXZ2phHU0V+8MDSnTPZU14C0GJlpB4GuEuUz
zJ4ocDw1D5toLzT9PzQeJcjK0HZnw6l3Un9178jmCCaoEWQRIaqdb/W9z3RKS9CucPNbK9uyfH1j
ER2p41PWBtlXI4Ox92QvHK3oeTLBTsrX/MbdEuxHWB4SbEtVw4sWfZnIvUxgMFM7NHYwUikrx+Bu
RplIEqixCZHGWDEPFnokay/AxViD+uc5leXtnu3BE41gnYd4YF9YGmnR+hA8LVThoKvqCj4pfkoj
5HfP1wd4sfmSa/ZmXfNwMOCgdYeTEYhT83jDJ5EYht8Ihm9IW3YOijxP7bFfO9h5X0S3MIMGO7xe
ZNdySf98R0T3Z3OMAN0F6E7oEqqI5uua7hcTQWsfJVNhnTmBaW7clRlyX3Y55Pz9CP8a+tNQ+0Cv
qjTm8CXlKGcCZBs5GgjdScYWnKjPjdDw2v4YGN0xlXJCTo7fGkveeDmuD1bgIizuib55UlHux1LA
daVmywkECK++Wj2onKByBGHjcpqb0YAuqhOuUvPou6e0kBSdE6CwPh8DBSRNPrAKMFL5PXWJQaQu
mVQDz76x5k+96dJHOFjEAS0eGAumq31Jy1/QjJRqm/K2HN8LSt/uwpK2RT2pB+qUPr1x65gVM0U1
wCI5KEYDC2SmNbjuG5WayW9OCcSGimz9nGhfdvyhCRpL5Djyh9JV6STVyMNTkLcQDcwYdaKfoalT
6DFckc6pmId1a0WwIv6wizTh7qzyZiES1DrYLOtS6zf+LeYYS9X5z7Q89EO6mSJKwOgNmov7DaX9
PLXQG0rOSKvPmKLCb8La43pRZl0I7adA/THKRra8l3doLIFvXGE7hJrxxGvsiaOyLfF7anlo9qxQ
DCQp9cm98ScDkXYcO1MebO7DhNWSmMbTKs0IISWwxB2MPj1xLUdNr4mU4YUvKVDvOw5oLMWPO7LZ
jopZeN8frKZKsODfKQTQ1x6+8kgNdr3x6oxoCtU0EYIVfsA7UyKGZ0Owo8XZYyFuBb9dIMoJH4Qn
w9RoWZhQNWxqSS/OAFBZBsmJESJ9ah/uZRNs60VwjNUzV+Mwikr4TWtkcJue6HCKFp7C5++QYKUr
J9zb8/d44DM1tNQF2gW2EfA28WzhL+5J8NPu5vKDEGp/fecWxBx7OzOo0Rz1Fg35LJZumsvPZ4v3
ruMf8ljelPAedcXa20caRRDoHcHlsyaimqkd3m+UBgCHqDRyqXEjfUjuVV+NSAcXuUZVX8rcq4Ky
4Bx6xmAyLWxXfuMSQQ1rzuT5ya6kxGlHodM7xQ4rmY2wFYCgwT955T/URwGsu+xK9KeNgBimqQRQ
PneK49f6pB22hi055gjibnrB0wO80soGUwfdT5WvFSjCrdaiMZxSy947TbruPbH+KqglDjt2Ps5a
rx6V8IpqOxF0rORWxzD00z8O6RD+4EQ7ykukZB4GiR5SUFlDcLjxgHx3ypuI7bU1o4jTazruz7eq
jve0z8CVp1nqVDpTd7RlI7rXhc/AhB12z5iN3v1BvDBJaKfqH694WcvORvHXDTTIRZpNF9kr+DBm
C62ecnRAO2E21q1bwEFnwj/thy+ylAPFOOYgMXwv1OAaFVsPN+Ubg2rZaZqqqsVlQTSWNtoFH/ri
Zv48wU2XU86rWEAeaoF4HWpRGb+XVgFKrch9G/ISkji70iqDAffNvPFZsRtOjuhq47w/P4XHu37e
UiQtFe8HJOJnEDePev+HT8FxGv9+mo52HrlJuATIUb2cPMmLibWaNGAYOoxqNVF0ohc/eLTkacoU
Vxl1UIV2E0cMk5I5aHgbjORY+Tzmj08F51GBJ8cKPvtRWVv5U5x83PRZ2iaPlrbYqYWLPYwMB3Dw
6Pcza4FyWbFcar7weIZ+MtZO/kh4Y120rTCYpojzth826ci6Jh1c0TrExRncRSmcwkWQ31lDXy+b
M4rTFRdl5bLy6UW+iFCwii7c8JHlgD6i7pgpPgTgj9LdO+lh3eqEe7gUo1xOPPfw8FNqWMYmps22
q0QymSxY1l4CiJZBpyWaRvbqqqNWQJZwUY8pVhlKS8o0qzDT/0JXr9bP2wLr9YKV5ryz/DrSNUlV
a8oWZUUdn1VuHH60wKwMA7gJlMhv7Y0y4eMXfL4bFFJvma5uvr2HwmbGUuCYBLQOmoVydKdG+oST
GhJ0eaSqrYTD+EfjQQMAWJVOnVl9kI7ys/ucPnKNkPRjnet3igjgBk535lsaz1KRjRA9aSwb2LBD
K1NCFizk5AubfxuXn3LI7eNpCjveVPBo5Y/v2gGE40RQ0qilUBlusf2Q0Ci3BnoQ7+SuKMymKLOW
gyhe57d58xe9IsDy7JV3e0kAwNDd3Tusyy1nuQgqMxuzHCt/IaSCHacVL5AtpXvM6IrMG0FMIVl7
anEqR60lfbOsqwLSOzseOQKGuSQhamzJAk/aknxNmTAI8RrsoG66j40qpg74oVy4XU3EH/17MAMv
dYIMNiun+jA2Yz59GTmC8fbVVpwTJnzTvBPGxYed3wSkSQPtDYcFzMngFIqdfFrUgxD2V13Myd/2
NXzdDsMzaHlImAcZvC49Pemv77dxUx4op51/o71TsHLv++G5acQVPUa3G3llAWY12jGwtBXtyqP6
erR2K+6gh4aH8HOL+AHOBF6lyAM3s2LtpwzqC04QUu2Q7ohFSst+gnScHrT+PoXeiWFt4QsyAyUM
XyM4JzUKRfTJwQ1EOyBIXssgE7a6W/90FBh0wYggQe9cydKigQyvz9s1VgSPYxRqZvdIK07EkCpf
LPh8BXjnjOV88TQkbBZCg0R6NY+CwKGySrxSV6sZ4dU7F/8JRhK5mf+V2uIODZE4uW4Ij9JGS7Ed
qFNYU6WSgD+y031hBW987L2Sr0EubpOpTL3UP+gJuTikynr9ZyyZpNraKgI523lp1Bv9zVF5acWA
cTZzXmXXxHzGLTsOhUBhqzUAk9w02x6ynNqFi4I6bQiakIWkbuH5/xTduP7/g1QL8FWgsrVZwiVd
qHLqF/5MJ8+/18Y06EuxUt7eNO/rR2ia2Zcy8s/IanHbh10bDFwHhisA3TkABjS1r3JbUvp9f7kJ
sv3HGArsfRnUkUU/vUI9HTinQ7e25C3dxoti8oW+0rbXpgJa0dDBG8eg+yKjQGTGpGMQJQK1hrSx
eHmICUOaIkHpisEA+JRzh4V7YXR36v7eDeAZrcM81st+ZhZ399Py/te6Ir6KW46YWexW3kpDuhKd
314QhyyqF/pD4+R3w93/BJDES/EBFb9xbLe54BRBj/0zK8wkDMze5izppKTxDWzOxPmFNsMZ3zE9
5rUBfsNspEwZtSiyRRFkeqjZKvEJldNyrsuEXCA6dK2Bt4K/gKKum2X9hQbW1sTJk059i97bov1S
YjzXqkj8aZ8gaa1Q7Wy0jmGpu9KSimbWD3snnwQaE1KSVb/5IwHAjN6muwQ7pwtlgAt+wiY7BCOK
SrU0ngL+6YbmvhEmtF1FCx8blNQFiChdg75MoBO67VSax0pHhXd4WF8sF03NxiU1DW/nLMkgVpfy
eO12ppWSltFP//5jR3Jcb1I9kUynGDjyY6s5mjefb2SJ8TF7fvR8y5Nb77M86gvHod3Gi+z9o2l9
s8A5/U6FKrNZx/P1YO/Q6Jp22Zogq7DYGNm9b1oG7h0NflD/AORMrAkGZS61ZHqKBuYqV9Vdxld9
loROW0q6UYQPRCdrzTwlS6kSnTcEdz9KB1nUzKRLIB+zNLghaWkfzqZLZz3tHB6Lc/Fm8NJHs+2k
WRdTrLShyQb/8LL+/1h6NVU35yZrR0FD53end2R86QjWFJpL/JmCGozWLp2u/A5a6q8u0Pc45PZw
zvOj/vkCdgL6A8xCJnODt5lzbVAU5lAsaDuyL1YXT+6v15X5WYVRsKHS54zCO+INNcXMWvcmmJ0z
C80O39wqs4EPEVz8gJcXg9CA957IQuwUlHfkbZeGzgBYF0ugj5+hxUNljMDn+IF+ghgku/235r/q
2cz4++phc+c9vVg8s4yrpVSS5jBK+1cZHdJ4bPxSeaysD7Eg37CpsEMluLKFDtljQL2WB0cBatK8
yjg0BbCTDR492z6czcKG3E5hnVFxPRs+6xOo2L613tDBwgY3skNEmCRWBLvHArDyiPAJj/eD5YVF
5HKZVEtUkOp7xl4ISJwXQJp4BHx9YSgN8Mfw22D8KsDt2s7c6GBSWCUDlNfWvqV/ObOmO2XFb6DI
1IIqYC1MzKPWi2zuZBKXNJ17LskjPd4kB5CDc5mcyY9DEpC+kvZwdQWsHx7CKVWqbdLbHiBa6Ozu
w4xQ2g+ssLEv/NSIOBM+SmAwYjfP9yowxz7FQQ40wKoNhDpgVtEGamOK7VYnxvR5ool1ODyrsosN
5TU/88JckeS/X5NXdQr2FWhe6PAkvi3/9LGTzb/OJonjsoIQc7I0LlayChiyAFA9rDpd3SfQ1pYv
Wo/gd8YW/dGr0tOmO7r4WKnoz8po0Z87/qPLxuEuKl4jcA6MLyQntaFDGUbvFqlHXYltguAMjo1b
1IqvsCJ89pfQd4spuLc6XUCsRkWIcnq0A5g9laIX8B5dwMNq4yD/dqCW+wqM0e4ZBs8BV9c9n7+z
of8103usUQWYmNppHVK1pD2W8CdbvdHDDfHm+TvvzpWYXBIzryTEGTcJaBBS80XghWw/G5MUkajt
PFl88IeAZvv/BDuozPFAVmkPHaoafVmv3SWKHApVGMbkTpALCDoK8i3LKy2/B1SOkH0chTWO5ZL2
4A2twdSZpEV+r5EjWIIIR/aamD7vw7irnUAWGCvcNzAisxEvTGXaoD763SgNEnkbSeoafFoFqJK+
EouHped86PX83kzsFnHYHOXGODo+59sr27xgmGgcT1fq09jElykboWqg1u1deB1l0LXNTR8eZ8QJ
0aRLs/MIC5JVyd0JSj2v8RpNvUcui+vJtYa2qJ6C4PwVJ4itKfRabSteiBAMCT/89WoVlouhZ4Xv
aZWZsCDtau/e5GzlkMmI+xMAp9/LnRiTZ3MbOTlTfwA2OIF2nsi5bS9MkWXeWUsxk54mq0ACDRc2
2V9hZXWH4GRBAsyv5J4j/3v+cuzUoF7xV5AKcTbqtk5L1Ejck8gk2g45a/8F74BKOfwkQl3r26d4
cEiMFabz4SC5qlxTCUZ/JDzV3tfWZLnHc2IrxoIe5+EvQ7JFMcZvCUskglKgzWL2MoRlCD5nndGs
yZu5IPq+7QU7sDe8vvciAd3MCz0FlpmuLLanOY46NFDpAyxlpAdVh3ox42oWn8pZRGaFzqoy0qxX
xlxtCb7S36IXRk9jp/WzJ+8rpgFY5UZPgXcCKBgOyi5V844Lz28C9Lp5g3aFXdWV1NYb2odByHJi
cnTmZyTaQU6lQ/FyqhMIyblOQyF+76Gvi8gUN6qq8ziBXX+AIt7aY/0fjRLLTBIiQqbOJGibcxD8
WISoUfMbdXeO0BgVOf/t4qb8iy8J/SIgHbEQzbnnGbUxgmA8dvMU7TJLS9w5A/eaIo2XdyXKBk27
gv5F9wneUpyUqa+RMVVg5EFwRNL5MVQqwSXBYP+AGF9R+rp6kjGmK0f5k8YC84aDn68TO/zwopFf
3AH6AvP7kK9Lx5r+v2pieuhXIB+VS+buhnHHIa7I6Da5Fl4IoXgq5vbex20b7YcDsms6Ba6pdW1P
Xlp6/grMZs0+aPdRT458hl9TR2UQa/O2raeKU5rJD/s+pBPphYZru+XWClMxCez+FlldPi1Eu6LN
cVKZWTOSGoZGbgjOqjSpQr7U2EFWAywvrVqM6tT+Oy7hEG7FSlsgOxCwuef77TgrlwY4ua4MolE3
8CFwZBFzxZAktnEsM1uQDJLmaaCDp4Z0ddJD9W8byctOh4W1mhc6AyPdtwwp1CLS9YOzd3Z4p8nJ
Z4vAWVbQWsComJOWJgLlFJhkHhBVSMB+cs7FOx2xlj+2FALO5+s5DhLNx7rqV8XEelKAtuTxbeVM
C+7MS+WrBV8WRloOgH9KdDBcQmT40WodAtu+JlDKm/BpKqbOaYnsKNalWHaCov3JUw3bict1F/kP
UvGRQNRmRWP1OdDLKijIzahh6YKnsNpB1gnPMXwDru8AWnNLPtUIb9noZXrHJeZSgRQ6euanpBFI
ks8dhahinlKfyBO82aixjAIP5HFIa+9ZtbBsp3L9RmYrkTnhqfwQJwQGkRxUpmwHgF8oTy6m55mX
Q4yXiMcda127a3l/XDoFMtMEZ1rQ/HbhA9Z8RDdvug9wZ/RAH0pFB+Ba4dznFjza5MIitsNn00pc
gBHwcHE7aKMQ89pAkZtdymdZmRPNwi8u4VuOeo8DNmBBPeAHT1D5llN++yPdGVI1wXHT1Ed1TBMw
M8rHSlRwH0zeQfFOGKoCxmGV+Vh3YPP0D23EwEck22R6/mf0wts2fpK0z1jETqtApUhfPpP5aFn0
0iet3Y295WWaHpBwHtUfPnPDTbvz2AJbH+38ASQf9ii5VXUo+5w8dN586g5Zu6NWaZA1Mmf38I9c
VURF6lWdsDJhKQb3j/ARha8L/3vX+3S3QShx1PJBV/4ww7elSJG32WTZBnE0M/tWjIrXfGti8MtJ
5VMkYqYWvLm4/vlddGj6YtioyNa6Dx4Ye6KDl6m66hHyyhsAbjnidwHd0ME/hZOKRSWTfOUspJkj
C2ZruSlYMKVhtKUUIICgT2WifiTPAS/yCv6Ve6ubDMMfYKsjaQlWLHNGjY6Ahp5OhJKdwgHvbsJB
+h4b78vW6+KZuyBzU16Af1hsDFWZN8CYiiark7eej++uTQ4aAk8lj5i6YFpo3U9/hv6bP8aRPclq
XkxUySPEDynYXUVWggKpV/biSiLBYdW6ptJqgDUKWeFHKL33iuAfL05wss6VvfSxUEf1vzSdOIq0
TCLWJJBoa5sWEi0bgHRLRPFxDnkOYb7NeSit7czxLnm26eX85+y7zZy0wUkrmlz8StKWv8eSjysS
69YT6UBnhaQOhUfW6hnWTPFyg1SCq2+89ZHxuqLia1n9f2+MLMwsPjxzYiuxXubLpXS/yP3FDW4p
3Gn/aQjyzb5X+wgsmMR2wiH97BDE5ahJNZtXqjii78vgql96ut4Ew4Hvrav8q5wXRzqoB6tldZzs
67K2UrSdg2OZn0MblbXdGAh7ALN1dQlzb57EPEka7txP1Eh2yS63OgA56SfSt6SwVJtpl1SRAxWj
vRWcEOnMuhNI4MOfOuvCyXw6AtdVMYz5+R31hFERIIv0vjLIt26cqP5NLoZes6Se/0z0opR0O58R
4XuHl/5khy1jWzTU2jcW8xVOlbw6LKnUx4lTMflzFoAK2c6fwbjG1gC56ZUbQ65PLBm+DrgtmKft
xXnxWceKJ1/qgf24VHZHtoEh12Emufm2fhrLN+vm0i5yHwZUpv4/x3BEKt1slxZ5u4JiEQS2ouwV
AHgqOva+p8DhZ2b4ZzKlSn9rQvrEaKEgy11Tc3GviEkDcAFB9nxJMKSnQVe7iVQ8+4J+9Pg7/WGK
If0qta8zJV0AKmGzZROGmNv7tl8WoEyFUW2xPCfeIJ11xFzmGOXnClta+FGL22/hxigvr0MRUYtM
sC3Anh42z3SHXEtFjJQj5apKMNGTzRxdrbSzgsow4jPF5mHJQpH5BwYyS3g+U3YlsBDGjcmFiAnM
QhH8ldpdbX7FheN2Ejt/huh98nTn+ql+vNcuBPAJSaOIfPPpdYmmdkiLLgX1RjkleHlsvFS7pB10
7k3qn4Wu1qVQ80Oo15+Iv5CTHfQFeZL1ORh8HDF/B1XXf4PxYqkJGTsIUTdnbpGDgYVfQzCeDpoE
44ANvlUwEKgWtdRrXXm7wpUWFjFr10lTqEGp2F+FeXNB5F7KhvOTXB5a6KYHqYsQuLu3783KU6Ey
8Ct2cXUrJ82KEw/5NukbYMiriooZcW8+bNAQv3trhqLFskJOUSdbL39dl+aBa/mODdfubRD26IPi
fZLl2iQdgFPd2R+KUoTvc9qihywx9TwPneSyFi8O5APuymoeCu9RgYTNwRnMwRv9VjG1OZSlA/XG
dKgj6OAEE3X8b59E0Kjtd5qadDaGKwaRwlBqO4yPFFWkHyBpaYMHOcu38iwXHnMM286k8jEW0rpu
3n921lOxxEWwv/y3E+x+oxXJz+NnxPB1ytM7CCt9NGYiMmmSoWcg1rVsWpoZHt6UxDpjqXxqClaO
yhB+c5TbXgWR1GnGIS21hL/j9BsgAIFiHz8aDBeM8SnWg+4iTTyyQBPCTJXT3pOV4i5Zx9JM418E
P2Yd4yyfAuCYJEnKpDl4lrvTosCrm/EJHE33rEff6zXLmftQxlt5w0ww9SOPP/Ciw5w67Hd6EfVx
RoSE/c5hYZuQLWqlF6HDsYsNGj5/kMm2TY+EjESGhrol6Uk2zK8CYT6CLoj9cS8YhfArQOpeBNsS
BxqaIj47RUl5vnVUWy7cDosfFBhs9/MsiRBvCtIhJMMIQvF3S12s7Ng9IJLWmAk64wYkqirEXRAk
2l80o8NGcmro+4c2ozYfBzmh0RCx7p6AeH17UcoSAZf9uHoHJ3Q/+Ys/HSN0e6GOJ6Bi8cGqMIqd
m8/pNxTcergLzZfigcZqDFzPU//KJcEjEzkp7jCUMlXYZFJhWHdQHRPcRcWdz7nhXO//tpQsukOJ
R7BmsPDXJFAFxNjqfwRxvPoZkx7HUaEYN9x0H24QiW5LiEU3Eyr0utUt+W74TP2DjAlfMtgzrIQ5
6QuxyFlLNVpMLeZBn7n8dWEk6ePED4UZKEmj7BXcH24ceAC7pZuWAirznSmuk16AiA4vztwl3UdN
VWzJuw8VchEjHz+R7URXeHFGa1Ms2teB6Molwuknn+VnkaQVf29oR+mrsZ5WdHmmIoHIXK92E3Xz
RGgDZZX4veUDs0tjB9jv4NFc64lb1SJB1cKptcfDXO47Dr0StPqeVQHvPTE/YiG+iauYxqfwEr+C
Tz7A0/qmpwGR/O1eFmT/U2hW1KRjJa3HWKpDR6eFhkuFjtQod9Epp7Ra7ezAtKONrkVlmqvIpEaw
EX93xIePkdUEDdbdFxw4/p6KOq/W9VZ8tcKpSqWlDyTtysiAaq0J9oPF4NF2owwOtTtIIDZOC0iT
2TO+NWiI9q0Vbp6LcCTpccfPny5R+WcFhUajjpdHs2BL4crffBZtlIEYnLxLzTU6xDjt8oTrWOPM
UQ0h8oxVfHIH56u1m/gRrxf0FrSPlTfZg8KzA4Ux63De7v2Jk0HkG30UODYOjAJFgLMM9JovJyFP
HEaSvPxFi61ULEojkI9ZvdHLCEw5jWm17S2m6IaTTI7sdJ5GCpYfOSXG85YP6Y02RrMNbJu/zNeZ
kSEUzNOIvy63qJs1bfwVF3yck/9tlR6L9pYJlTyLuJeyaJYq7Iv/2O6SqVweLwyaOHkTWbkKOpow
bgEyO1WizzmtJSSBifAVAH9PDsV8XXNMmuKSAB8JLyu0k1wXnCuYN8Z2yj/1uy/s2kHZEoLU2EPE
dvbHJ0e6rQvQ3fUAUrSd6DTASBV0zX7Z0jC+6EDFG0eWLk7GsMtNO6gphF+JrBYAtaWOI8ELaEdj
dq7stlrubdLl/rBuV1yIdGoPuC/Bux3ZXciPRlKNVPReKPMBS9t0B9cfL2Xmwk1Ncpjiu6fYRbQc
wE13jJkBhumqccYbNI4Y0+HZ0CjJSlCrnTW9eQiIIdWd0kFdq+BvM1pIaROo1HtBtvSSte2l0ism
7pqsC95oNlxckUEX5RFXP1xa63Ec6mFnHRIpqPUfAd0KPxSNtynBDzk5a9aBZ/S4Qy+chHRc7mR2
DDc2T6qxKPh0PnkRPjbAx3P7OTPy4Hfz8izop+zGADx7joJ2xhds6ezaOrQ9IAZZWPoKWFGNbxfa
e/rag5llYQSxzKh+rCfo1jOpmngvbmYFHqkKOlrgyb1I6UBAhlk7kWzINJzGJZIQqqZm9M+3x0Dq
XC3cL3tSYbfa8zrXFTkGB127E2+gzRukgvwtVV0Z4pWXSbD8gc6iSuhr9tstyt6vox3lK1BbarEZ
cgNL2FyV6pkkmOHhyL1qpoDMAG9D0nGlpbItk1cI5/KK8YcP9jdxyC2cD7T9LmToE6/gBGRPWaRK
rxrhAWHu2Rh5nEw737yAfgWJ2sFAUootqk4osNmfyFkseloI0eH82EqcPE+wG/HD98buINXZfZ8N
7rfR1KUiaTIb5c0u/3cT5cErO7ulZcS31W5xbcOP0Q19muq5FdOTIt+0GrSqo8jVjLzpcFz7i0ng
j+bLJvecm1pT0rogzDjLSYE3QYhvdEhIkZMeMRLc3+XVi2yi7m0lTaVOKMuuR3/9wk8j3ch+Bgdv
waM1Bwqyj8GqqeQJSKD9jg6qdTv0xngduEkLHdE5zSDsruT9g8QO14RGoYsS8O7n1v+WkYgXiuCX
LFdjVbdUMDUCHRmtV7LoacgrbX3SfQhMXwFeKZi//fj/qHFeKZ0dpVxae1+2FtmzP0MsCeNdS4w2
IVlR6NXxgCD2kW7ZzCvylofjTuKN4MwtZUhqBgILB8LDRntb1DC2wDw3/Vc7/i5Yn093zQ60cWxL
SYoL+T+2+X7X7KfFSJODXsRAruXrEDgFEfvJLie12ClzF2De+jc9mEddkUIsy48Bg3Os9FKiGT88
65hSMJt48PUuf3uqRILK5adAkanh20DbWeaFTH+LzOu4CaKzZ3n3AF3vG6nhPORB4UdlkFNV9inY
RTp7xtzwWESemJ1fslCQBm6VmJIL/7bF+rSwNW1FcigQlfeeiviccwTTZD9rRFZX5OY4vSP/0Ev6
9yjVEzu6CYtc7SRA9tDPF0busAahOnUXDZ86rVJ1Pdc+JjGm51gWe9CV0JmBq6qqHOnlOLk6uAdw
yqOBHs/Ta+pNiiOH6+j3CVdxzI9ISwug/kQaPsKHfOQHIjqBBcA2nJsmhYeQ7K/sGIXjZpiGpFjT
hl4tjkz5mWO6XbnwYEcz6VT7gycMr4/vUujDg18ZHw5SMrCWK5QIDQ98LoqWx/eFsxVcxdSWG0aq
JCnPSZX+hwBSEHTWli0w0TtUF9VtGkEVgCsxshIBcQjNxJoUAoW5mHWh7/29b3d+6CJ3A8oaNLbZ
O78EtemAVYY/yQlofHybKM8jydb3j+aYmfwR/L7xHukBdHwFeGto/5DoffWmpU3uy+9E10pV+H3f
pgJdsv77vQlLuiZtTuXrMWo70E+645Cy8qdlVxze2xKk/oQhAidqKmbzxva71iENpz1Vsw0uPJ8j
b5X5u4q7jnoAz5TBchmKasD4RgedVg1YMcVuqxwe6tCn3me5PWAji/RBqAGVRy/q/mwWOeHjcj9O
JovWxp/nR8iqqUwPTbsFBDVkD50DIUQ0/LKPJT+PI3DT5fYcuLNLJDd61f4YuiJ6Rlra8iI7eWBe
HMYbVeX+sDLhKX0TdVnN+DDC/SzmWIOXiNtPIkZKEQEZUbK/pieuZOcOKwezkz98xxre3tB4rQqw
ZDE7dF9khvEKkqZg2YYPlsS+A+FQ4DyQDJ33orhfA5K5AGeiHfp+bvBCCfWrfzfYtxrq9WKyAV9o
ezlytXBP38b+us6j97nNNr2liTHGTQRA0FegCKBU+desjJ7vbVwb4qjmmHeiXlkFz/xeDwIpx+ac
Pk61+EJkcaegx92YqiG91CZK4SF9bGiN7ndyHJwVhTdxp8zJmziIxjyWGRyE9Q693fjwGm7ETBvh
+LJaBDls0PLKVVunc2wjw4Q2O6JGGsTpt4gycWfeEMoiveJW6DaAWbkb2BwzhXATCYYs7UjZVM0Q
qPIM+8e2Seoux9Y6IiqOpzVu3+vLLI9dEdME9OykV+kVyNh+GdAoIRqQioUP0ef4QstHd0RixlPp
vzbVidvthuo+Yj5vtHzgEemimjiBBDqoVhw85c5vkOM7GBnMS8T+swBV5usgheIa8qixWlNKVz6q
r/GY4fYJNj/4sNhwgpDa7L5Bd4A6AgpjtVY7POYumaP/Iyw//9nVIpYK3KxqrUV41d95FW5NIrT8
iQ+eDVsVPJuDQgvpZ7O7OxZGJLWYQWpBzJIOsLKi5mO2faMInGuO5sLdq6h7FL7Xl74Xg7baMIwp
0ZjxZJlj9PFnmU/nOd9PqBjlkQdhobIXV8I4Q/gCxZtCdDPoDEXDGaWJIw8qyCji2R65hO2ewG3x
1nEh5hdQbXNc8Qv4bv4vMm80lX6EWNvHYdLv026mYUXZyWdPzellMSgzlAa/v+A1bSa6XNO/BaTb
6Z/4Ytsnkh6BpbpEVuM3EOA2F9kvF0YSeaAlUhER2S5UwFcxqwkShOW1NyMxLd+5aGc3dTtiIdY/
CQdbaY3K0lqg0p/4+TbJCL2E+NpAiaf55SYN8tS9l+4CnwhMrjEHu4W5m53oUbJvMX2V/Ch8krz+
BtgVQrewH6cYNyjDivvSBnIgurz6FU6N9u2geo+55smbO2zuz9G/lU5rzBdCfOio7AHyBqCcdcd5
Hy6pAL0uoYwxV9k0FI9XqDenp887QMxu1qG90rdwvrrBFKtt2cs+Jak68neklBM8zBFRwxSQskmm
gXyamu7MMivAyLbvbqiXne/6qs6Xju9Jjl+JMtnWApo8XF/XzHhRAVzOPWF/9sH8m1Y+VgLcVjQo
k3Ac6LS13ME6LlCbLWQX3RfZXhuiIfE0MPJdHiti23qNkp+qBDblRt+QYzZYWHiz4LCaVdDT9Occ
6Var7wRn+9nYiGfoun35lJcnf0RqGoo8wvG8v9Hc+Dqpe59/UcmZnowH1+UtM5yvy5hnHQs3wKwf
lppB5f0WNIezYHXg8sXPi3AB72N2QAyjFU8OL+PelOnE+QED9bPerNH4ldooQO/ctuQRJVscm/1C
+6m3W5ukkH9j2M/XodHUUSHmjXav9qh5biPS3telq0OWXLahQ2duiWlLaX55nd7x3DltoFJm3TOO
qj2Ue17MqygLs7Lg+Q0tt6htMv+AuCYJg2MK3Jt34jAger2W4Aa8btf6mpaRWZR/b1OovmrNgeOA
NTvVwkMMbPjs90sMtiZmRDAA6QbE20IlisKT8g87Wab/gYeW5ozT4BhRCKHgE6e7mqpPYnQRM+9r
JIkLGnYH+mwWQ+ys1xud1pPBLAnO0uQ/16Vd0lToEXoIzRLg3FqAFRe7ZrYgsJmMimuSxaB1+qCK
Xnp+qTRHVx5J3YfgFpxZA73pSw2STfc0fgJZ5x/qeDo5aSXuHXcJ45JkH+D6hANRW0CIsFoqadg/
0hOop857pGtSVhpTUAaaimX/4l95iikxQ4rpLh3hqp3XsSf19vEEuVdFXkq14g5DS4z8lwEeBZIV
8mMVPBIcQaiDpgoOwwYKZt6cDgSB6RMS03hL7dd5Mo487kN2elBhFqOFJ22L0t8S8wK3ys4NjLsG
Tf3vVvqOV2OmJgEg+5bCeZFr0U4/atB0ECNhqDOWcWPFftXOoNt1+voy6cEAiQ3M7hZMweCdXH4a
k1C0NN0nGpfrJlN1oh7UuS3KOkGz2gfPEx1PrifYRMqqCNSByCdME8+GNi4mFLxw38+sfkcAU6kQ
B4uaa8qSR6HVs95VxJVt+U8KY3svA2WApgbxGeyob9UevBHkDIcyEmVcbPUYpnfzVM15/O5EJYW7
OLXrkeh9DlncleYJ4MwNQZY1kbhNYW2a4L5fmKSJhs4rAIbFCPuftYW84P7h8LH401UHwJ3TH8Yq
DchC7c+niTeDbXxtGo3jRAQ4A97Lm7Z2gu3VQuh74bBRnPdOtGQaOntU9dJ/fXjTtewtqEG6LQTK
c2rKr+eSf2Fua+DIPgBBKVCiTCoCDuGHWylZ6pH4Lvt7mCSGlQ0RL6kf2u2xOvkvkEozqs6nVRLg
HCHnlG1j2sj1XenocdRIBClP6aolCAHZKPcu/fY4VLjTbSW0bD3HI6+MhOg35oMdq/3N+30egsYR
XifdHc3f9g6fBpvv3wPfNKN1ad/F7lrFN3721gcK0es0tmq6H26JPTTqo04zo8MZ8O3VSheBlpfY
pv4e2S9AiQKBRQ6U4nGS2SkD8NT0R+q3Hq1doTG/JrR0VJa1QLm4qx8WbM6EN1kwqkepAkrEDT5X
J9aULZKhKm6F4v5Wdz4Mj0TAaMIsIblnvcRn0y250xRuOvQ3Ap/e4yNpwMWU3KlLX5A48VizEmsL
IUVeN0lB66mokgGFc7cLVlMHOUcZCQTxlT5AS7LOQpz0yt3xPwlDIRtlFcjyZzKHYQvhsvzdPxln
uEMtVSaMnin6OTm5kiM1XxyAGIqNmC6D15Q5mQ0IAmb+VTimpwqKSRgCZro3zOwrYdRZ75nW4Cb1
XxPKusf+CBD+SNjl8EFnGh6kMfmEChWN//qGy10VtAzi7Txm815A+EE4W64iivv9IBvmiPCq3Fg+
SlPw/dtPE2i9iJlmbERyLQRz/vv53MNHJFiphZOd8hHqRd5iQf47UG57l96EFIPvpNgsi3dqxc09
BA7OtGmiq9ENVteY74KQrUIMKkCAIV+a3nbLWu4TdyWlPqmyeRWNfRLXFIoSImpww1w0Ro61UM1z
tmJy2XdKw9XtRSuUsOv7QwhAZtLjJCWR+hKMXJxnOw9+OSHabNT94xkR+lyPzNjCnRECThVZ/BuI
mULxm/SapiKFtFSf0KQKREVWz+LnTKLPzz7YX0oFrLHgA8b5mz25FPWo2uQ9rdGtYO/1UwN+9Hja
4BdVyzVIUvYPH4IJI2EJyE63FoXOETzZRvJ2Lm3M1+9kZ9X8918le2OfnrgzD4palEjjgLCbaAcn
L6ztFQIDowp6230ONQLN3voS7jWTZe8H4xQ8u9aZFDq+juOJz5pHgpenTgtSwwtKZ2tJB9QpMDyU
HB7dc+AMWPS1xc/0b1vS34BXlYOXegvf8nfBlXQF/iMC982KvkuCFKpmqjMb34JVMjY2V8fvnXW/
1tfGJp+z6o3ME/I+hApsMQ/2KYJqBeWDOCkjUrglujxvM/JBvrzm6GF1UyD18CeMvhkfmbrviKNQ
V+vqBugr6ll/G54BqGsehOrI74CxCAS+darltCvItWWXct3gpPj6uvAm/UUfkZhUMUtDmVzvbNP+
sRhGUnfqhZPI8yXdunn+9ZQnrKN5+JnovhELyh78TB2gqSB3qcfTWH2ok21WulWj7XzC7hgS7xm1
tCUcwHTbrMD9ZQvfhSSKyY4kcvfYNbkGdBtmP3I41vOCzgnCaWCAF2aeAdtLWUKs2GHkUewBGplz
ffi04EUZZtDIlQBTvV342vVPOpO3KIEFSIAnGL4LXPERUiuw2KbhaS2SQX78iOokhv+FWslotg/V
8zIyDlb8QDWLYCMrNickHKm+LuSZODBnzclGj6RFocqGSg/V+BLkOGVCVWulrJhzsSgIMvuM3w2K
ya03XXoQVKpSfSllumI92lhGG7lY/SgQHpNM+Vt09G+zcABhWscjjJYjeiscW4vot3a+BSYB2Yih
kd0OL7G8eq5ajvDi0XCho0fLGeJNzR4RxoiiScFotLVNg5HXAvQ2EJkqu3qsrrTXdvI5azw1ZTm/
vM9p0KQIqdpZWV/WKi2p2vZSmkwQDImsasNi6WSU+BpzozQicz8sly5ikVd6JVIwjBBktQ6fNkTC
EpYjPQtuC6p5N3cmtVz/mQgOKGMSVg9jLdKI8JoXbCvdDi2YL6ivNEFo6aNAZoKv1LkAgwlE+vdc
4zu0Zipt98PeiqGFVPI3GMkSOCmKLcRNEeSUiPagz9rX9FXVpKoWqX7nz2DghvOkDlnZU5jhkB7u
Gx4pho+RdknTKpo/ZKetxjPVMo8doQ41ojt3r378DpxIAKB6TdNbLmMLto5315fjveFoTpgsDBu8
G9PGhK5VBAcQm6r2m7UjvEw152mKRvcz+yrkpwtrpV6wd7o92e9xGzZ+ybGOcaLkJ4iTSDVP6sTy
T+F4z1RQVJjloNTRluARDiePC29oD+qQ3XDTO9AgWHbboRNlMb17FRtAO6k/+aF/CeMU89R1smlu
Qd6i9rgReXSr8w3QtrH1wWRZcI6Ppe5alv4LD2mOk8V4Q5llMaL0mYjEVzFiBVf422kPkFpUM1JF
3+D/tcSZY10bQKzrWP8qjJf2jUlUJmoCSrotD9fn2lNDXWcVA5zxLpTojQSutxe10ivuzYQR8jnq
IvqbHjBNC7phvUi8jpM3STaJGonkvn1jssb4ARPQA55zOmQ+3fgNez2k/c4YuWDASd3MkFE0ttDX
JkcucstgwjqLWscduHldcJnnrZDGP5kia+8KuHZAI1Fjre2BwdY66Hp+OKrxm1r4TAYWuTlMnGjw
1uvktyR4SY5vPL6IktiYzcK7yJDpU1nLO8w/esTSXPko3RNRp4lIE24BjkY1TicTmnpv3cRxEM5O
gfhKxGXxU2YhjUp+yvJS5Pp79unL4jaxeHBfXA0g6rsVyDrZlaZCFjJW7SrtRGi8bmoP3mJXB81r
jicUVQYLcNR//VbIPMzay7dOhTYgIfmRCa66iYA2ooL1Q3hZlapCmivDdEL/g6QJwAKXW4wUN3lE
u5wCuqollY+STWGG9VyY2wXOJbVSboyc/4E9FIs0XJG9uI1h2KsTLQoH8xIc8YQPp4sle7ssmYD0
ZyLJHNtlKtnS9BkKB24lHtF8oBhnhlAxIz9+ubujFhJEz7HEwc5/kygHBjB0VgVNYfq1oMoud162
EYXNqp14ZYFlNK/pxISwy9m8KgH9WX3pKMjo8XdFADFPElqsorQSMYEjKDJ2tImTMtdpeeoVXGOV
vTSo1BvwxHDl/ycypVcme3a2gDFhPadZKYcxL/St9HKDPjdNsQ31yw74xcCYod5VKXBc50aE5zgO
MhMIXNczFQMN6HvOy8EDs2YpineVvdn3DRZkQw+wExDZ3kgen7hDW2G1UXbtnzWWfuhz1nPtva2Q
2v8N8Jj0XnfrinGMP4eSYi0QJbc5rGOrhWlO4LjqD6CCxXo8WN5ZdMI6adMh60WLLooOrhrqD+QG
FtIt5kl0W+8oglFrs5u9l7g76sSS7rm2U1nuM90yYQVBq/8SzIIjuMpDZw58dvjp6BG8dQYl+mY1
20QGGslpP4vT3X/hHJK9FRASXYxgIjL7QU2IQmVicfYjT7Ea//D0akqNnm8wSXlZhNddqb/CHiz+
lGX7gE20VohpJFssTdNAjCD8YKK9FLYm6eOCwyixj0fVyFeBFV3LjZmjogzFaMyC+/cxtmWSdy5J
BPAnJwn4/nvOWYoSrvo+r9Ws9oOTd5zeS9XYGiLU1qKCgM19RqRg2MPvU1VeGCZId1XEztDN7Ity
U+Le1j4Vc2OHN598qp/UHxOTpkhHYCvtBmfK1//BFC8REsHZww33c/GeDTnvblKHRh/4CQ0PumMb
CpFtfKL+YCFnETpMm1A+4j50K2FvkqK3fw6PQ1Lcp89uZ7sqQiwIDKg7RPV95fh7kuS2ow75E0Rj
EqQsJNvA7u/sCdz7mh41b+pxXVZWV3kwIrSxcHcBkWoTGpzh7HwX3MCFYJktrnoFMkKLNB36PPna
5aFWig8mkHUrc6RKKPw49Yckw/hG8u33ntJpHLrhT6zJocnwLVyrHJjHUsp2qNGAsDxRdnJmw/JT
scat3fXegPS/iu6eI5cy2lEOplzEk70YTvFmVyIgLfKuOQsBizIPOwxUPTTN5T5LXI3c9vJe31Mh
+bSk6OSJgQKFc7LWXvYuMQzeJ/2usEcgWhWLkrs+xu2ZvG7Kuuy+62DE8dAjTNwrbheegghjKBHA
nt2svucB9HVKpdXB3O6eMzDuUdhj2umhy3qiNY/yKdAdVEp1trmqK964IubN34m5/EusEzvxqF92
FAzQ5kYEr06SjVXh8DjTMjfA6ANGnditsvEtZgAL5HCjMGzHB6fjTKyQz8StENm/HZiK6guojRci
KT6uZ7m5g+mGjZ5hMSP8+6Le5zKtBH+IpyXj1DlyI+2mCBZcZk0dYQENsyv8q0t/gZBB3brqdsCq
YMsStBQLjKZj9JGhvIVaWNcm5mWe7MdNQ8oNkjWhpD7V2wgfdodpR/lUfuot0UiPVHBDqTOckt8u
rByg5xacA4LT2G7D1EC38fCoUGVd3P8eNLnBwus0r8dnntdM9msXMhT24lqkTeW6eA42mDSXovDm
aw/WlrLgBXDCYYPHsfVZv4pB1Q/ZjhENqobI+xz5FPJ4C09B1RKaEjbSRgr52jGylBKa9umqbkjG
HJ/4cizJqYYeD3O4RMveBVbRkUHH30SO9rIKBZ++DnbgocbE4ZrvCFWm0CS23GKU3dfOkvG0jr/y
/OABHZ1ZOf6FIpIIHBHJEncjQfiD1OtxUYQ1lpKKq1e8GMDEwwH6nv3HVfHhTX7MRlrBHuLDfhJG
P/PVyqDhYYMEKSZMEWVMagK1NvGsbuRAgEWapJMvfUVtBhCh3rnzzc3mLjQ9G6em8os141GQalAS
p3lvKZ55of/zryYRXk4Mi9jjnRTDWJI8EcctCmt6J/UbOEmwV/2xP1FFdCBBXilZK1SS/ZaQJf26
X6w+AlrcpJBPiX4+3MRYI6/+t40XAzezQIFKbD1iAMNdHxZ3t+E676cdMuYdjyVKxnFy5WaKM2KH
VpQ/fFoFhlgqxvHewbccVvOKP68LDGzXcxGUdcbyPXQS8kOFPqxZln6altTVUA4hVb/1W42lqG7f
77vboBhf1iF3Yf18+VALWF0vPQy6kfgvTxOoVvvdQQAxxgwGAsSSgR+bi8s8OATIOWy+zNMV1xfr
Iznpz2H8QEKOroN+nbYR7Ky0YJtJrD9s0ajKQAzYp6rB3XtrZ6jBp417rXZCkNL6bM5L9ca1cf6X
445ZOdjLnzRGBtiVCu4oAeVlZHSQashghDN7DvWP6zeyyh1MvDogisVIcZ9HrhuuiJ3g5XtG21sU
bXgC3XkRGolKqnfnkKyaPgCq7uiKajtHf7INCzmTZj+G90/1bSWzSvSsLvL1nZSxULhBvcljOVSG
pZacZNGuF9ibYPiZJKnUOIq6BsmKEgn1evC5op/oiPErwHM+mRps+bHb6Q579J7aV1Ux0Zm4UzGq
+oWw/DI6gfM9xVSMr8wIx21xfs+wBvw8oMrNvGSSaiG1IqIM9y40TgpY/xjAuUM7ThGWhWW/eC1p
Wap3W68DjQ7M5yHnok5o7a4zgWCIHr0UkH/UwO8LVVrXDtKAUZS/D7xpEE7wY59kY1vU4CtQT1MM
U2HpyKyfHlSzJDDVTYzUtxDYq/7FtKp007GnUe3vDzRTkX1sw3ZS6QwdL4DvPHVIeufAnC0+Q7sy
+h9ANCGlxSMeT5RhkMBTE+rdiljN0PbBxsEMGrxQYzyNjr7vM/+EmRAtYHZ2Zqg4XEa8SyR8ZTIt
tLgvCci73GDfvTvfz0WSDSO187JaezPiEhed/C7kfsq4K5a3I8zuf51ZBpv4+oJbH1ws8m2D9oiv
YIhUlQLUuvsXSTzKrxvtX0SGoelGwCzVtoQQkvOuGHzxws7NSr0Dqxlk5WZd5FsriBD3hBTyaxI6
FC5W+areVw+1rOOzh2esDZfg3w9etwrI/BTRCRRjCrdXtk85ag3rFuV0/HtNvKxaoAhktLNxnDmY
NQTdcd2mQHfjngSqqqg9ZwLovXwWF3L2jd0ruWRc1DiINOcD79+PwVONCd5F2imsy2dSklrhGt4R
jH1sdPSuldwk3qTxy9mIEGfxQvkhTfRdECizCGPXdGb+ZrUhMrh6Y4FLyvi1praME3Uztd94yZUx
DsG7zJ5n2J1PgCbKbTPHy/AW4JZaC+fnSeVaW28M0DNGjsKy0O5YNWkaKS4bJMyUcO/pjHoAqoLq
1jxbAydawIjaz56sMzq0M1wNdhpvm2P9tuVkNr0unQTU+iU75xkh8lZAcSe3TmORTmsWdaUkohB7
9gL7gg2tmT9DdSwjcXoeTGYSoWIqCZ/SCXVedyz9hzhJVnLLKLR2dw39zpJDWA60ZrvyXRpqkyVz
17hRkr8YxJUsP1+RC6v6877XYAWmAXdL9SINkbyjdVPUvaDBdKiHNYZPGPd721Tagwo57PRYDtt6
na8PyRin3zsl3lGSi5JHtEvIly5kRYLArQlzFxeNsAFEdAhdvi5KMydIjj9bXhPvTYR2ZVrJ1SdG
sYFsEy6cNoTZaz00ajnHg0kIHAsrwJ4hrvE1lWCYK2WPjp7MWLV/ikzvXayCaRrEg2PNtYQZULtP
SwTTocd0ET+lj3LruvBVfhQhit3+uYjG3CEr0lCGzAu2u4ZGGgZUa4/PrjmY83divivJr5Zb03bV
Y3FXxqIjgFf/SJuZ+Pc0BpwAMpz8cQ/MWsomWm06cQrc1L3Ji8Ic8Akznar3YC+BqrJHfukO/iFY
wJiktdyzXQZNrJUEA1fbP8mlv9fln16l73pnRP3WRGP5WN+7c6D3qzbSmOYWfxcbOfU1+X7qbGY3
V37S61UfOO1UUv4jx7Ae9zIPZi/HeqcUenlneBOHBvNi9bxSpaZeYOpJMPclMiq+ySs8AtVd/pW8
P4OUk2a1ilWpn5BtTbrogf/0VQ5I8xhsHq3njxn9aBS4udyk+fXad0/Kdz2S6eZP9Qgqg1IzMDDl
ZPWrNv7maddx6pE7vS7wQVODPv0Z46jjJ1puVkLViLvmcmBCIaCxeRW6NCib1OVEtG/VqGlCu5m2
/tYOk2xJKgl5j7+YqyTHtR40laxM0iMiB0ovRa/NwyFTjVAF5SA+dP92gRx8VPXYiMMJ9BnjW6q9
cYQwGG/UIOOTzDWMLEf8fWtJoNvxC2UqxTQdGoLO3ityyEJuBVlE641MVzSk9ZSY+lK9febcS7rT
z6svA+2FR6bcnFd2AuUWic2IiEn9sCXhoTR0nzH+TkjCdWwTxlrP5zsNqUcwo66hDH6FHybZcBap
8Xkxy1KFaz5nkEH1KyK/rFYPoAEcr9YyNo9dbUhLdwqvZI2M9RDuS3Gksuf7GHGsYaO3IP/7jW8t
DylEVHYp6NfEJzUwstGXwS6vQbc/rFgx9ShCypRB5zZm0/yrqOQjfBkv2BiC2NprNznnWteVi44e
kGIVs18uEkfHUD0MKTrWrRhEp19hyu8L7Tfif0xCUB2BIM1gUZCdLpIlPmwxQY5S93w6espayF4o
DEEafHb/S+xdFqdGtWNZJusx8QtZmI4XkwbLR+SX5S4HCQ0Tui06YRPHWu9xb5/edz9Xe5HFxn82
0RVEzvlDFJ3kYJ04UZ9cyL8ZPF7JLwoia2KOK/f2TD11+0LTjypz2knj+eJAx96w+htCzTPjC0rf
pNWLH/+zyjWErwNrllICChvxkzJpIt+YNK3LusSOYuW7VRcNJ4zL51EkpaD0vTG2qQxhqoRS2oJx
+kcCe+f4SqPvgb0i8zd8BzVfGwwB0cOdkuE00WkofJDLo8Y06zudUtgCk+wMZEHNpnu/rCJY6V4Z
igSRby6YurcDnDoyFVhTU+DBrh9DNlBag+K6Yz0n1gMSYkGSybHYvmnSQbYcKTib2uuSaIkYhXWM
1giiV47P81Bf21xLMfOgKznunvblFLWExjHCfYhgzDRgMzkpbdd+kwyujodAH8/YsfgFmjteXf4g
M6tUulfGSitpVpjTz1mSNRU0BawyaAoo+QH6gK1LJmwkomWIzwQUxJbKTCOtpoY7CAXmw+MCYglh
RhZY12iLTGREOL6ma1McRbdwEBKLeZpSCYXM7yy5U6bSpRRRsm4LtZMdQiCA2ivYvgY6rvigGOpZ
PxmQswsn4U2y2UFZAOpzdpsPol4O8K3bvL4x21sU1lGTUJPtXCRVVUJmcD0c957Dei+qn1HEnZUh
vHwmz2pDJZt+wMM9tfCKj+6PyRkRhmXzWXDhatzw70WV6wJEAE43ozZ0WD4rln2UR+k1K4q7b5Ah
whw/qm9Q/8xH0ilAL9x+AfrKmQT37JIscgLByVmHTR2NJfYW0syDyfv9advf/f67FdIFdukvj5ZA
0WUCFWZx7U0dv7Xdt6SB9YT5GZtygUTjyt5zhDq3cm0OWF3etxfDJa9O5pvD/ZwH266JwaZjoz+l
HPwl336dBAiLBAVeqMkI7iDf3k6Gi4rpHk4KcZC3/zhwjRMyQb/RwTIXj3lfe3Ey0g41sIRdsh+v
yGErMYweApr8lMmjSeqfRc6E00Rvea5gHblFwTeS3sSqZcRFcWW7Phtpjj7Q30o8yuQruFuJjNZ+
4XoS1JzE0nIrJULoZkOuDNK+GLAUz8J+bpyhtD1Jf6xkBl+xH0VOvpkthwS0jri1zix9PDA8dCcm
Jq8jxgyUzfskgkoTTKpVP+dTnCWvw3kkBvA9b+1HlbWMQ1mRLcEuDw91wuis417WdeINm2zva7tF
WQQU8+9+zorN20aMGruUNkPBSS+wOjMbHeY4rrsb2iiH8eofkiV9E1z0AcfyZkW/xTk2/jR+DY5K
EkO/+zVOsIx068ZgEKhkcTaqDUyZkUEv6T2M33nSNz/0IaZBaCVMHAPJYeIVoA2DH2BU96+usabK
PmRcmLYAYfjX9nyHpbpLiLtfuWM7+DSIdwuo3/XWhZyEFLKKh4vNMGzLP1vDJ/sSlWI4aBYlJfM5
mbvdwx48XEbndFO7V5vxclw6kWHDB9r7FR4kxv1QoGPyREiQuL64VQAE2Q2NwWF5DOm7Vsl0lX+o
6KxwWqFudew26SoR4aY25GPIEgRcbiqLSYvjeI8cTiTVxUM9rF3+u0/WNZVOuFWFvvLB5ccUirXI
uBmTA8wGr1+TEmTEM4iwPvNBsfGOaHnLeATrNVqctJtC2A3UYq0nVXtcDoysxuFdszBfdoootZyV
2C7gkeCeRJGKAvINDDtJlgleJKa9FwGWd3ynP1FOChSSaONQ1WLcf74QsPIj9Q8qBLJPpYMUaVf0
kjeODTwb1BQ6Xdh4YGsggiBOBhL/nzeu3N3QJvtTFmytzOoUUBqFTEzju+YdaOCjbND5jDjc6l+V
TMXfCKPfIlN9O1iYJjQlAe/jeQH2cqoqXboaEF/79Tl7rrvrhGwXUy26cSw5VuR+Cb/SlxK7Rkde
9oiioiLrauV1FblGOgCRTbwVW3IADa20+z4Jm05I5/nqxQ1omnS3wg9hp2UCK6CEFSNi3iBxLEof
MZGkcsxR1Om7Nx3mOHEjZ9v1OJoHMCxUV/KePI5MPgUKL7Ux7E4vrhQvUuPiCku/xjXLaeRfZgLn
I3nROkrutd8WQ7+S/PuqP81vb5DZm5fok2OtIpYVnEWeNqav77EWjJa0dbaCpeNjQXpbxNEGZJB6
aLKWvged58tSTyeaF8iF2yWya80ZJJ6Fa/KZh4zZC4ax+VzoS0Vyd+0Npa+mCCknVEJXdWb9kzsC
P8NfuWTvYz/PQpu3c/Sc9QBpV3E+2O+TmPJSpyomU4ANcHqMj1zAWdVSfub3dCwrcmHIinul3TWZ
13hBvx7S/1dAVXVjaoJP5pp+8NaWYC1Xs2o2TzYsNuy1Ug7QKoNIXpOHu/aHiAlBLs4Kaz7w47Bh
0Hp55Fn/OX40HHw5JHCtbGV9Tr1Mw0qI3hjIKpGZzVx974gXxLhakAPWMAOUubRj6Fz7FZg4XrWG
ixWr9FYe2TfaQDCOkCUTZVSCj/0++mMvPuAQPwfUGpvRNEto6n2+q+zmk3idNoO1hWFG8Sdm8zDs
7iNbWoobzHoXuoAfalEZlNWFaJuaB4pIOZyq0vWKpChptVlVmsHDnPScLdvZaOH/PF64UrXoImnt
yxypiBOfUZpS3eM9DF53GXcGmqvbPl2CfvL1yKncRtiij5iYHxemxXpymZ8DLLhSuh/F3qv0pR/1
0gj3CZEeUv/idAXTxhBveBLXobwYQCbEYKfpc3sk5M0jzKu63B/H5HLHgAE26psQrPDbyuTtqHGy
n4ze34oqqNSOpLys9BcN1hLTlP9citubt71Ue+nXH0oA6O1lbmGZo30ZwiEyoonJU2MRuksDuIpG
YNXSeJfJr5Ua47qX7hRXpc0/sp+P5qIK3buoEVaxzmvsMOo/L1eV0mEB9GpIF3WO3DOoxJX1hBTw
yFfuSK84wwNZwO/eXaTuGy2zKekLvGATFSRuv4/nm2zZUt3xBIKxloTaRiLHnp8foSqz54ddFBYB
/1pGHJYKkyBF8tBzumye+AWwrAnD2jiv1rjOZMBJowqgUeZo9ZUPZFBnZ9S5+7HBxe4DjbmX8EYd
gzWal++EAimFj40an5B0yKQMwRFM1ux5oDNfOaYdK2FwCJ9736UpyQ/2J5Tvc1Tjc8yoJUuYORXQ
KMbdSjT1NplrUWHY5Ptat4S4PVeGSUTsLNs8XRCUW7B6ttcr+8fgo7ExUnbNoghHz8g1PDX2LZVD
fqqrOS7tVyLi/xRDFJwl/OYluPIcQ524sKrpUWh/ZRvxLzuA8ATzpR5pYq8U0SHL4HTiFFiZDLFZ
mw0CvECrOxLl81Khq9rFj+p1hbaC2yIt+FC/KnlGI1iIHFTmxlP18s8+N6u2JlhSoddxsdknJ5dT
kXGrvFv0BsCxjxa7f3xRUoTIf0dD7s1WtR4zfMo+8E6VulioC7D0wb7Dxp6c/++wxJOD9Ga2kclY
yIgwEVWTQHaBs7Q8UBT0D6bK24sYSc3wJ/YlQ9uUXz/M0k67zosjBfJN25XnMbkrs+GLP5JnFStt
ktB3b4ZLWyhNRaMBZcxA8+KpQXsfm2d4NVvAsa2wwmIg/AZMoGG7BitTwa7bURLWoGaai5EVxQ3j
uWFKZeC3cTW8XavXe3LD8Bye1u4+eKG3iNYBj/aCF5pcWu505tVahDnEKozBR5W8nyznzSvTsTpo
vWL+9wrTwSPV3M4uRvD3kK9x5kbDZR/BeSPI/XKzzy4eQNRz8HoCn+Ir7c0nxbMHzqFwbZ3JQtvS
K3EYbkMoPGm1uhUn6Gw6da1BwBKSxYvfV0luPSlVqP2JFr+DLW+iXSxfmehsAbZ/J2oUtxGb1sO2
ffc8pM9m4px9tVi9zgINza6ndM7dHubfEkzNxw7cHhNcyePTi4qaJ6q3XRwhImv2qkiW8dT9nzqM
SvYHz1pJpbM6NAWvzRWrcb7yI3JGMot4C9t7XrgWXcxsoKjLeBtN16bh2Mm4gE92Ru/irdVBQKaL
MpG8RK5E28hb6l7UXbeDg+1lqFAo1qsQGBdLofiFuMpxxgtQOCZHDduE7TQGEDdUAOp8ebwf5B3U
MpOw+UX05Bi6ssbTK8Ir8/JvuyhL8r56ZI32niJfa8NBJ/QdrbAOC1X6cFC0vvhDtNLgIBBM2MCE
avBk+3MVpwz0JcAY1WRrBLJY+RNlDPug4Jy/02Em1Qb+xohhCc3us5VE4SnUEL5hc2UmQoEB7ske
Xt+iELyWdul6OgWMAlol1X/ohu4hce8tjnFGM9xNgn6BpfoqYyMRpgtoDc0o4QXHcBd7A12FfnS8
wtxxZZSya55Z4O4zMFnu7TaEB/ytjp7xvinsezDKo7N+HvOu/LFMsQIZbL3PA/iDMJtU7BKnATXn
WW/rpVuBJzEjsmCAFdDAMSQaolFtTYBusVC6499pm74OTGj7/MAm3nCGP7IH1cSzeeF4SKRI0CtE
Mq2NvFaiztAWErMi0iMn8rd0CMRklWTwGrWUbo2cW3vih4lFhJiE5XZ/X2eB4EkAFH9Q9dATaYrm
UXbPeGvb7QVamJXEQpJC21cizgX16kiusPQuln+MTZUiu0aOEehb5DZnhf9GBJrmZRA78Wa6k98B
RME/Fhfp9ELg+nrOK0xDO6ClJHazNRhZtyNUrFrpXQgRy8cEENBlVOL3kr1kSlVyzCrPmONOBgWK
y/R5TubFxsHm5gTu1LOpL5kHUagMuWcANGyiX4bdO1HW4Aww3TLZ9ZxTFFnEU/9WbSH1YKV7bjae
5xdOF5gamF8MtCviCmScIGXg3fFORMt7RLKSYCzk8DQmXBc460sR4/V/yHt8PJPhy/EzLUi0ZV/K
+LAw6Wvhu2xrwJyykZb2hgtMC9hxxm1uhxJKJ4GR/rhRPZZliW/eQwC8UGEPiA9EE9yZInndbJWs
k1fQK43QYqSgxLIjSvco7I/bxZOu0aJWGGgz6pXsuc1uNhdTDLpdj0sxbRPsX1ev8jhtO0xGuQIS
iyV1oOqiU+d4qjbBf8d81UYKBR02XtRQctJsKVBSmWf6kIi23RjoqLrTRc/zbT+VFrUExfgaGUGP
1dy/Z0WsoYwW6NRk/WbmZsgJXlum/CCZYiSaNwGG2XAeTY9fc18QnO5a92aKKRU2P54WHD+qpMIA
qhpMMos2sBB29RffmI6ClXJ7XBNIDAw6xWoUhs225u2m5hbD4Aisws+Dv2PHjqQzRwhh023DBTAJ
l2pnlFJz7wYxy8ym2gd84TLqBGoIgPMv69+w4Sx6Z9HQk9gB/7ELVTZVDHO8chwFNWj8wyJPni81
y7uL6Oo4+PK/R9HDaiwTxbmhuxqlky1bqae1Xu09p96L4biKncplZTJJucdLNpbeH1dZ/c/F/yXp
ddms+/WNgYtsWbAS2wYjoUr+kFZqQw82rpTmXei3wKBiDtkE4FO1bRd6sTEgNJ4CE7rz6zDc+Kid
BZzgJj/Z+ASKAYOKlpUTevQaIquv52uAbITx+3Xl+nll0ddAmQWpicW+Fiww8FpQdcicA7IBAvXd
16f6mrRMFzyihstBfiguZW7nvnmW7/julmafKZTXNxh5MauSP+mGU8xhbAzQ654hDzPCS7m6rmOW
6awkjJC6QM81UGZh9Rr46HD10tDMf7s17AZlqZiGbwqhmK1AmOYDPjd6za2EPK0cu77QBp7GkkA7
9INNQFOvuj5FcpFaB67GHb4Fv7q5WVidy99o4FQb1Of72GNpZ6q7ZyTswrSyTVKXIyrpqNyGKubC
Scj5NEKT9BOrJ3eYCgrnshxuknGcx5B8gWM/L3x5QDWKJiEXNElNIcHcldRjGBrRo31tqR3sLWp4
B20KDvMF4Z1FOhbdQJMcz04+cXtfvefucAHi3MrFXlx8xyEGnhyCBlKpfCYlSMWDoAIWX6o655qA
OT1k77pHxZqiFkLZ3TAwQ/cxkIxPsKYPq5GJ1IX2n2H2fCLLCP4do663Kr8A4+ngHFZzVtXvCP//
6VgeS1zCMnyb3gDN1BVvN7ixUxLbxxJJL9mGNcWhkgJwQ9D/tQLOPUEVqnmKrMpuQY7JwJJdmqu+
DOwGOBbTzywAX2YPVpsyNfdJoPNHM4KkYneNvNQMPJVv+dDpVVgypEftjXqnkyLyZa7d04yRtXiV
lBXThbjNdQHGqX0Ik3w9Eh3OTDBGJyRSc6I9vD1m6x6o7kEE5nMZpZXwcWYfGLlliY/69N3FyS62
Askt6b1cXyhKcLRFyV4RZlkLz9GY8KkdWs+H0Z9DoWkDUDadt7TacP3kkJLx9lklA86aFuamqg+A
zdMCo1gLjd1qmtiktcA0O5iYje1b13iBXwQDZWDRle+Q9w1yPhRun8o0OLo0L05eF0LlMAepwc+e
D+QLebd0HhYHyJ3UeZUnbge1wr45+IOjjIBRE0x1k3oQ6wBMBlGa0E44Tu+okK4WEdA7Bdt6lx2w
EdNyg528Np3pFBZ0v/ASscGAtIGWxJ0UIA0IEL4nGH4cR+Q8h1Wta7F4Tqnsl+NgHc4RMXIeKvvY
UqGcopzMjj6fLBuJNkgyM+vJTJQC3DC+IP5PSPL8580mGrNAb/CMgl40CcTstG6izzY2yrOPAVzh
9l36P3mw4Ix4pHOBh2kRFTcakYIbdn/JKFsg/FBBo5QOijXXtCq2DDihZEew1RxbJqTqvc7RcCUj
gyzR66oi+1XA1LjD7LYNLDsGiaO/31WMgHEKEyKkNfJOwXfp14vkpONCEl1sOtM58f/fe5h74x1w
XNS3LwaX+Jr77r2CJCcNXhubNUiaBwtYKIF1MPfy4X6iVJtWSXKh+jdDGGBrNajREar3b/J2JZ6E
WqxXYHKdCmm426mU3SNQ+I1DfVREpjT9sMpfoy+XS+/NQca0IKLFlUboac49zoOmDyzn4xIIh6G0
c5PqJiKXO2iB6nAlwRg3yszgX6Q5BlnaarMu1rS499vUvblJMleAWaUOueaMndxfsZp898/EIbVC
2o+5CLEGZce0+vvUo5R9ZCUVlJTM45RtCP3ECoG+OcYk4UsUMUpXAlPTUnu2RcUlhyqWv5Fk7ETf
LqfJQWAxR5pnH+y1QxA1EC6Ak0/Ous12wUZRfafqCIsnxqb1A31CDUJrya4hUSY78tSeLmgkJENe
4gNm5OyHDP56pJbl4WzdqzHzsu8v4kMX2REu1Ho8gw0dSDjzrKLrZL5k3w1ybCcEiwaVBlYoZqnW
CYiddFBa2pDgqHiMYarOtrg0cQ2XZPC0MZcWX08IvD7xQ0yDMPHwcV8WhQtJB+Ekrx3b/Lh0sB+U
1ANVHX8MSxjAN+ZcMcd3kVyN2Mbf9i3+6b+uxpCiUDdP6+DpmDDaVzZ7HF2JLBTMpJ6oVnmv2TvB
KEMNhr7C5U3RXmYj50bhiwueHIu3GbUQpFych8CPaLBKGiBGVPHE5Hn6kaofj5pe93sfSh/mG21Y
10ncHVm+xo/fIoXYpdJcRoE2Fmit/ohRMtY8EzFU0ER0THt786FsAfBAw9weLpQUgt0b5XTVa3DU
0YoXLooA59rMuquBK9gu2e79LvQuI5TPvkONfcMNYjhR1a4Ylq0d9oUKIHJSTYcDGJFUO4QeeXhP
DC+2spXTYLfzdVnPBkLCL55bctHRcaXHWggXOwNIyaYFNFz5xwhDEP4j6IkUVNTgjbzRhBkrPZgr
BZT2+Xws1TQtqZnpPCeYw7fXVHFHxABcNgucVdBITjq7qsncCnk1yHGCxm9w9OruK/+6OZSlZnZG
0EwW6VB11qlmESp3m2USf+PCgl0lFUD7KDvqa8HeDYSwnYyNczozT4bha1o/yB3fqwyf+Pds4bnC
x4JqNJCfxwoOD4J13WOcX5BMIsB8bqbGyEmPTCHg+VVWAu/d+SpGO2xPORwKSOFrHKb98RJkW1ZV
hJfOZj/JPuVBiq/CSOsqfmHX4BMsJIWOIMgTTX8rXy3rB1KbaokbHo599G7iz/x0FyH/yr8oYA9j
W8TuLsVOLG47cE/b/IstBiV9J3XM08XGBikOiTKyIAbj38gKwCNM5mGWmx/zQ9UhvV03hXi3OGYX
PbElU7g80no16tqKf/2xIfIInoyQvWj+RWAsrR9kBqpiQ/hvrdk/nWdh19lo1KuUhJV0D39oA2yk
ZJai+rD0MgN8gJPb/NKktgVuQrpqUP+O3f11ZXsOZdWUVHADOVbD7GeFhyJ+ya/IIiCDw7jkWBWq
kb/3Wl2XaaF8kNxHVCtQiH9TFJjsPipSSofDqJtJTwC1siqyqzWECj1x5L9Wuy25qfjA8f9bybES
7rcorAxkheCGWdtiyLo1EcQVv63Gqx3xJK/hyl92uDj2Wg10nIbBAQvNL3o5qwnPzGfZLbeodQbj
9gjiq+7GIfGfsZBcmsdEKh0BrUUd4cJgsNXX7b5Dn6mava+dcvmDHp1z9Gz6ke8tE9qAp3V8aLdk
JEIAXXzKjsnTIMIWdDmWxi+K7qwjymltBN7zGOdMBFweni9cUDIdjNm+vPNhf6rlM9rVVM0q6a/q
5C1JCaM/Szkq2PiQJvqETBu4rT0mPiZKDOMAHTRI2dc/9lKdagm08hRi2KQvTIns24wIX+LAfASd
Z4TY+vINaB+tnPSS2V2Tp1+Wqld5uDEaHz9wtQAEoQjtjN4T81Pmj59YZbxTaEA2nXC7//GbBH3y
DvrhK4bGJGChzXUKNO1tfJDVpNYKg55Y2G3TCGdySz+bNOTcFtJrTqRIFfwW/vbXCOnbAPd/O9i2
+8WctDRLuX+DOjv7RWLQaEvferAGUEes0TBzcGwfV6md8Kyh5xNlSroaiFl1Ue0p5LtqsjuW/8XY
ten7q9HtwEh/vxsCtdpS0Sa3D9/ZkbQXJt9ilBvUJWwmdqSyxEmMXFXeO8m+m5BsXdX7ajbxDmcW
nvuQmc2jxxrxvUZc9CNNSZD5qWJtNKrpAYBHjnjqID4LPodyyp/OIZ8XGxNL3nfFnav9kew04dPG
DJWkg7ltz7QhLPVKAEB3ateJWGwqptvL6cGnr3LU3kR18wWBzOUzHj6d/SgH0tSQtPX8lsI6fUAC
Fi3cebn4ddUwlAzUmXr+u/csUC6Rzv1wlO3OWcXTJ91iqcBh+S+RZfmqYh9RZI4qBTsk6UhJu7OD
jRshIA6izgdruh5bsZjb2q8yG+5hWmCcYGVxJxqZZ55blaSuAJimstVE6d06cas4UAo+7sDm98MV
B6qY8fcgf4O015RRN84M1HzkAoH+jOisTj/Ll0vajpJYCXyJqjdbGNz2L1OcnSANzgn8STbIVMYH
l6JAeEctaDWwfWlwtYwvz3I5ibiiSJj60mb8f0EwY9+aB50cjeoN2VeGFTPELAW3IIL0O21/aISD
Wt+ajXBcCbZmmoCvM6oTdcaUaiLQkrGuuUMuTIoJsAOltgrCTAtNs86w6h7DoBV97ZGS7fQU3XnW
0XcvNs9QHtR/v+sQ7Vg42/jz2277sw5pxLzcretF0sVwohnJ/yJeAsyLKbtKgKIeE1/LLNodS6l9
wgYTUpWdsze2JIstfXFMluSG+PO94wFp1eXhDJqzvoaLT42+JouiJZmYAn2ZUcMyEbocNtoOWatO
+/66vpOIuLNNJnN07PhFXiohaS7TNf8ckCnGtudmK1HbBAaoExLwNsaKW0/9WtHEv6Hlll5YIFv3
tqW2Zdb6NnapOh+HFwDGzs6tc/mnGx3wruhH4T2WwximLCzPYqbJErMDlareyI8f9sL/zFRaQP3Y
ntMd7ex+RVOife+TCZ2E65Tlwz0hqK0VBPRjsAM5TpRziXtVNN47u8WRJe2jZmpCitTrQGw/S7Ah
sYP6f6ipYF4BylQC17lDm9n5BrE3K0ECV7UKHDQkV6Vf1iJo8mT7hQlmQPbxHaDR1aGOAHR/3Cz6
TjjzEGK27Cl4yH1l+9WLYK1bTcTEk/nNN3Y19qaFSYAQ1j+3GWrjyDngde8FlFOifySkZ6sLMFRx
bzqlEzGj9rMx0Yc6hF/tQ+qSizh6PtvMKmvH933B6dSdghfHiy/OJnYyORXXSCs4EcwFauCBABAu
ignplxjcIWSDxYVpZ4drgW2SaqDcol4dEPoEPwKfee4DaRHV9Rj6S5rBc/+/I/QHLPMKj9vR9Tzc
N8Q4zSgfng1Ja7MPXhd6nSaFwSORHD5V+KeVbk49TJYbDJVzY+o3yKDOHB09PeTXX37LN9yPbCjP
q7byoIfUXQ9NAmzjf1TIqPxqkDrqucgljEUyEN3+E8+S3DacGRkDqIekE9dx52jCg5ogi4FBJscH
G+kVDHqjDo63CdkTlddyuzItjhLxprKZ0SBbD1/W2R7wCAJnuYhZqMxx28EtDd6LTqDqmXtR2Pwd
r5GKLyOdLKJl+xnm8McquyLInlxjbP3Jkkdgf5VEN8IMyzGe8dpkO+z1/fpdxP0NQH2bklIAHwx3
v+ZmnMncCul0ANKrvmFWPPOKC3RP3VqCL1VqP2G6YobsbCmfnGcy6g2kle8gJ/JjAyT4q/IN4Jjh
C0O+wMR724YykeWK5Jz/oa6HAvqo1HKOdpx3B4K9uqrCHc8Uw3hq2d1fJrIkRmXAaIh6rcK6qIJ1
q+MX/Ws5GS/3eP8/qSDp7AGEjKz5YKE7NrPQ8a+gK5HumKYWPNHSvFrhX7IYuzo5o37PZHjt0zrD
Ga23QB9llM7jrNg8iXyeVJnSqUX5yVZnc5kXyj9egN+BxW8yvxruc1NoqQiIQK7WFyOoHUwFpXlx
wSaAESDqp9DLZ3Dpa7rWimchLStEwMtw4GKee/KRbVrzVWQC8rDqmqOrAgaEuR8Esc8lIPabQxV6
QxUQfNoCvkGJbPtqWs+V6ulTjjn6Pc3EUXI0Q7V49mW1BI7fX727MNgX2AyNd6BK9qs6ZbjjIZ/+
O9W8gaIRRBoQUr6i3oGf607URuaUQID8/ceDUsg3AaF8Ht+qh1/kXSnEuaYeaC61sSo6jWigJ4w/
u4xFwE4IU8q3hOsDJzFs1tCcvkgeIWiQ9HmfIKWdzZVcU2+Fusv9+QP4QtNwcp907sYvldO/N9iV
PWW+kns6npOP4dHl95rW00AxjyRIUDHx81H5ZM/S+SFjOOEsLgQapxnrK1MaGvJ8M0A/FXosZjmA
nrIPqv0Zz3uD+lCkYZeTPQS83J0LSecA3ds9DZeopZJ5ovbBKnZq0u87YwpD7JUGKFb8W2aOYNlY
5qLRo3+tdXzRsZBg0DifIQY17l9Kyn3PjkJL1bEBTulTFM3JQCPGKB7BlZwdZGAt2s+UwRhYSVUM
5bjO4+fNR/aEkSH51MdaoxgRrciZhqSmBG7AFgezOHqutmsk/sYl/nYluJAF5i3ycJUoi4eKhman
2iVMQgX5MkjsHoxWRyx1Q2LT9xs52VGqhXO1UxjZZ2k0qcEHkY3dvIA5FKhIobpWhtjuwRMKTZx8
h6Ovj32VYR/zqI6+3MomxX1nXHXD9jviLunDm9cXaUObaRKgZSvltGhTrxE8UrKTeqnzMojuYCBe
sTAHcuSbUu2of7a7YIwCDdyOkpEtfL0TdLb9wIyqNjbqUGDvs3rDHRvOX6S567LIBUgevpLtnBl6
NZpVskcDqDeN2ednAW/c6VPQzRmtUydonNIPNgwC2y9ZEncah+WLFuL0/Zi6WKbfZBaYF2mfv2kI
w/QsUglpzKrKxHRjAmts9y3Nbm040J3blhY+p9V/UGLFUmGI8PB3qf5vlJmvwVnWMIMlke8GA3jr
19lk9qvEUPP3MndaYY6mey+naRJPjKXBoFHdr5OYfPxaFbcewGQSNx/cAKosNXkouKqJOSGaGJMe
GQ+Eg576L+xEAqKgEasCJ3WIPBSrM5AmFBVvDsrOmzVVESPbKkhv4VQdyZWy9762SP6axXvkzaTK
9f11Ql7fBkfOscpdAePtZh/RudDt2QUW30awejHSOEVAuqHKh03MuCUd1/kOLffRHjc6J5+S8mwv
NQYV0i7/ioPrI5Bq7HGlu95Ah3dHKyHkkWxv4uaiHmB0aO3e8Gh6BLajQLmbp7l+HQXxVRI+Yx3+
R3l+bfKIx5/IJWTC/fVaot4+rvwHXpWp6MDZLbGpxDOMRErovYJyiLmhdkHVLYLmDDPeOg45fQeC
NtAbou2nBqbMePLeYKb7nU5qpx74JMbsCsJ96SLmLm6dPdK8qSiBgkJDr6VxmLhRKPAdLJk0bfw/
0piRWVpr23YegYvY3HFYESAHk9l8ELvOGy5kriUZelSUQL3Do+R9Fy30KR2qoztnPOqUfk2ZTzas
PDjiNYxOGbji31Wyebx20unhOJH6d3kVdfJGdoH39esORiayFMiYZtFaOhqcs2f265SFTGcRT4mm
eg+Kt0gJrGhT25tO5dPwnl60YRMXO8PxkMjA66r+D751Aody+NZBBrpA/Pirg+8vWIse0oQ2HEdr
DC9Cr5025jbH7TiWcSCx+MdiL+XqkdvkJFUEOuHT+8AEui9oLqH+9st7E9iW86YV5OBAwdQuSR/y
GlFWFQKrUg3rcllmWzxu9PtuEjjkqVWt7kdLWkGhIKYSdgzPP6Zqb+cWOi1C/zpVv9qXHdszuchg
JJhXGbZFZsQFpwSzTkKqEGhlkq1fUxfuog6N7PsAk9OAZ51wfKDJ8nZzwYAP2Cf6LqXsFtQytSB2
cJ8X/64GvNEbOGERzYYZvm49ObRxKNR7S4OW/Irp2OXZCzuSV22KXAoPBCNlGfqxWJe48zG38+Bk
I4Jek9BdqWWRfDl9eERkm1VkoPX7uerph4q/iNpM1LWFqkTbWM1lezU/L3FH7FJHCutV3xWAls96
J/BnO5xllJ9lEhUikCMC6rC8jhaJLPaBNSpzHsJB1qNIOaFRwnkKVDZw4DBBi1Zf/Ty3Fx9S8w2e
Jgm9S5+hh3wlTRAsCqB45FssPVLhEhb/EeNB3N15waWMrQDGvGlwvThV8m8CHg/UaZzJiRRmxkli
xH/xfKq74RBV5WibMPL3Oy+0H6cDnLot4dy6+bm6I2TmPTDyGX7Z1LoHb+86cCHRxHPTJtifkaP2
MkMrH2/DjNAN7UG4vkAb4tTbCgEOQUxMALZGKfz+EIry8Cwsn3mKkEGTcqP2HnC+oN7vMgKkZGkc
//TkhhoX1qgdp8rg1331Uf69mA35YKecH4eIbGD99zeHWV9J1b4l5k5rtJ3jv2OoYw1ufwy3mlYL
oDHlwlTYRbgGc90Mbfz2iVErNFTSEAUOGPMPe3bqAey8J0ganK10mFOGT0UPuRCwh74TOyBw3dNa
sqcG+QSv3oD0RhKsMi3oh5BKT94VpiaIJklz9SzyGSwEzuVgVzJL7/n5aYNytwePUAmeAKI2TvUL
93W9J1LN2HCrazfv/WJ6Nx9nF8JpuHsk3F1tBwG8N21d8fGT70/sVRtZIUBxy94318UgWSratdV+
/jy85qZ4JzpzsKHb/t8FqhtQJ1gT6RWQiQs3xm8g2BdqTmOMlLtuTRPqNWf38H/ySiH45qIfsTXE
+vRC5R1tQBxerpJQcgxDJ/uARJQQPVE/wQBUT1c32Unt5hq+0z+ODqpv5bDj/8VQD8y65cgzAXO7
v+woO4BgwaxYgoXN1JlIwM6f3ajk3JPdnBf8hTo3h+QYzl0sQW6wfXnl7csa02qqv2bivvVAs5VB
zX123P9yYn24oT+M4xHTSe+QRkMwaDv5xi/zWzDWiPP6cYu7a75qqGaSyTUAdHiX81UpAvYiuYVv
JT/JmTvhwYy+9ed2EagIspaVGQ+DMg/YEdCyxSpz2EYr+1oc3Sm/BiCRKngy2bP0u3pEB+aDfIlw
x4K1QGdPzYzMaXE6lCZ8amcNISJ1Rz70nPHAePteF0x6gH6z/CGuaT1Gtf2h3LVDsnaru8VUYWMH
BSk029AnnLRgdI6pM5L3ekPnDSK+26ffU0DgsAdUjqGaI8rt0fJk9fgt/qE4WngSUPyvM7cwvnY7
jy8ATgKbI8YRAeYsUArXGEdlyceayoN35sU7/jlweCzK8OC/0eWx36HB7pF4rwFyLT+e8yswfcyy
/PxP4G1pGWd5+vrWWSLMcD7glGjeSzcucGzi9z7VKbQ1r3v0W86nq9GuBKtTZWn3/InNhc1XA26n
ujGJU1CsHt9rnnZykwdJE+nQ4tbjSz2DrujMQZ/PqGyKAaoi5nMjEVKpLHcI406GunkD+qBJt1bD
kXnbEjLKNaTprpXu3Fr8jJTeDbJpkg9ox8wHzZy6Hy4kkZlNikb0pDiJukWtI1akvVFcxdDlG5Dn
23hF5eXUIC2z246ddZIYJjFVRBsaCbBO4IwNdIALT9p38g/YlcSoe4PZ6yaeEerZxeBnTM25SJHv
BXH0NHVJ/RI7b5gHYNOjhTcQ2/29QoWGSN11Ao9tjaHXk8lO0FWYUg5iPQFR1jJen0w1YS4ijbpd
ADAfD9q59iFKjd1fScwM4TxgbmfFwWkGi6qcZE4RjSo8eFaJQcJETAqUEUM8P0o4kxX67c5Z0UsV
RTCvP0OnTeZ5a6dFEEDb9rVyCeacQJsVzZFuNPIchbVoiRkMp+Ah1IKUtmpbXpJAgh6W0xBHKbSl
JMqAwFMi8KwYZI18T3NM5FSmAGN5+waCFRN5IkM8uzB8Tt8xet0+/Xh6j7jHNDKq1A1P5LJx32YV
1VXuHEzTRWuRnVz6zRCRMTUFh/DNBA84EWtCNkoDdocGVVV3gbgHwlTrO8YiWu7FzV9LfY71tCTa
axgvrrCcKwWp1SeaDb+JPdamZm2PtM5fG2e0/VuY0Nf41o0FEDq5rqoAG10rFc5CRKwZqHvBtGtw
LFm0O+ctC+A+lyRqH+aJX2FZgHsEXpMZ32sFjMhsDTMyfG0LOp55u/5/JjFZBRXlv5LMy1Ag5gRw
qS/4D6rWs8rq0bxv7p9ZzKWrs3RE/diOe2V+dPRpbDJ6NvTwBCH6USon+DCKHqOrz6oH7xo4Wur/
AeNoit+rTfWy8+LWpEg2ElIhXf532vC8lPIug4xkwt2ojVA/KLZEDZomEMVFA2YvYnvBcwzexCZg
XEssAhrY2W8JN5WOMWdN/jf1p4FvTQD8dUan+t1GY2UGnSelMuoGW5CpVzDZrwANeeTk21IqC5Zj
5WZCn834nqwVh9JAgc4wU7tDL3iv4k2pcs3XJgbGUtzjN06uwvqoOxhznp+3cQI+ZQTy93I67Vro
Y330aJWz67ZBPPY/45VqNbLv2RzQEX7ShsGR/s9Mywe2W0vjgoxIpKnKGdNoeU2e0vnuZF64g1aY
XP78KULD/3k9kMwcBTublHppmXFlNoNx+3+M8dgyt9715aqKHuGvGlVI1wj/4GEyL0oY2Z3o/Ip7
AZem8Fbl85ZkeiUt5eiRqOKo6z96Lfpd53wh9z1CwJX2w3wBnSTgHQR4XXjJB6xxDIKdwnglj+Yr
Q7qnjhObURrNfwQ+J+EyE2eA4F0NSdFyUpyx6NTD90TFgemq2YPZ0hOqu6yfAumibZSlGZbr9Sya
YCAE1rfXsm1pb9DA/J3TxfinRY2FPwmiFaGgw68Co2XWvsxnJQHfefvGBh3qP47oUe6MK1ZrvSus
sn3nHcLTeUGKGOtZ0yWEQPW6T33QdZF55DEr9XlfAE2y+EqFVdt/4W5mK4W4WF2xWKGBmPb/WUsG
7haY+OH0kK248cmPOZ7i7e0YikWGBFonlPHoP04mCidrVVeQNRgOpXZer6HsD3vnMB36zzPohwt7
+Mwz/Iu8GRMHtfAbgRw5+w2t1fNH8WCwz+mN6lNus5GNhE64QeBty2ySF/dVDS0pSWElTowPwXXg
i7Ff1Il1r9+jwLAo8hWNf2Bji/OnJz0lKFMtIQ9Wl+iZDMsV+U8Ph1qKGKBJUZ/scIAIOCMHAVO1
KdouxmrFZo8sSH4BDIvqwrCRpMuNADPznO9zLS73o6av5NgrN4ahc3L3RNVYAfvFs1d9871derc+
i9WE56govGTCcdPZlpL8awQYm8dezuWV9k235sYfxY/cHDeKgsqRPyv7LaELChJ4Szm4jaZEUY2U
5ejsghLOWiYgKraJHrWIb4xncAIz2OlVBjitn/sT8EfnBAWl7NKEAyerei1E5XCjklsdGgfUDh0F
fpxqLeVoeh9hzDgud0kzUNakQ699TTXSBUaZnYK/y0aDTh7/7od9Ig6cwt01bLGbUj1UbFAS8zem
eqpu1o9HJj94AvgzFMdndNsxC8YQIEHghVks5dq0r5xJzvG+f5gufiTf+C9/tRvZsemhchDBgQ2Q
AoDxhPDxNcEQTibhKVYEN6VPC/EvaKm8xmCq6VcLk7bgWSskTLT2QFTo7L+vRgPh/p1WSBg2izD3
y86mSIYHqyHhfYsU6ttb23xT5dZOG24AUht4VerdJt3417vCNnl3deObKgb9B8++TBM3wuO915cB
ViQ6hdydPmfZsOBqK2TGKyZfcEUVANCF9ec5XoQLxYmMrcfPYRG8ORAEwiVe0foRQRyLWkTC+V+Z
9JBf3+hM7shfVRoK8QOYxYHCXtl3KLgnAksqGiGrkoBhg7QyCPPxbvg2GvZ+kmVg1oOuhf1QCUDt
yRncKGJqZzYi1xL9+v9+P7BdjZEvWIj9bS+BGfsU46q9DURSqecS0x4YaAnkBVtGGEpoP+m4q4hB
t0pvCUPs2ZQqnb/P7TWHS+U4jK8cHhpJd9190wTMU9D5lG5+3H4kcQfK19FFnm07+ofAl5l/4Mx4
Kn2+p2aosWXuTr6BkKfwcZ/cv5hA68Lu6mPwOXriVo8U74RUTt9PlpwTwI9y2r6OEG+zEYqf9wUq
CUrSYB1I5LWGS1U4HaJ+Ugw4iRuRgbPQFRngw3NIRBIivgblt5UWT/MJiym6EKUXB0kRHuBm1dVQ
16x2uia5O1oS2whCwhuLXHdtl2r6Pkha0ZSL6T2A2/YRzZtjIuImFVvPZFKS1jHUWjaSztolcRgi
d1XPiTyiBQKT6h5bbDI/3ID3u9yS8ZXncIPJN4ks8qFFIFZjf9jb2QQuh3/WllOza1kkdFVKHy7/
FVcHAm3mEF75srHFWCgCeYfwyyCbAcXv8X/kIi/Hqkvmx/ManKzUCa7bA7pG/pi16pZPEdq+GZyH
2QR54p/bh4xpWFSNO/h1wqDxw4k4JZHfzIfZKI5UMepaGxfJ9wmhkHqfByS+LVNZQkSMvxc2X8L6
wioegvaeL3e897vO0NYlNUAbHDwm5olcyLSm0ndT73HIo5pmu6xeHlrHvtNMGJoAfhXxT3g3fC+m
KDxyO/DWhMdcMSqHWezEORHY7K3PsT+sIDJ24nBt1LrePvJ6Vbs2crV65otj1FusMpC8rY6iReDd
pAAMPDsj3l7FVW50i+Yje+uzDIv3Nz/lxjFoV58b8q9dhfaI7DKxzUteyBxHkTUO8Qq3zYjLPw4T
xgngeFvGe4L+EV8vtn1gZ+R+mB0dsNzooD4TzgJPnwJWKGyyBa+/t9FOOVFZQXe9885p4rBKuIi2
jd1jIG56BgAvManQ+/4jsk/dvPQt11sHmgCP8vY41ZZDRPVN7TF7trqlfG+jwjd8zytDbfc0pqzu
5f4TChe6lxFoZmfGZ5qOuJ2/42JFlQ8b99RCDphzcwkxtG7gSCI8jXsvdcb+Gs8U71GIhK0bgPbA
/PAN03akFokpai/wZSxiEO/m6ihXNgEN9ErsaZ/NA+8Fn4Lawoj5naaZLFUJ9EuBZwfwxebyNWxl
465YyC9tRgkv/DCYbEhFilvlFch5wTdpR0UYjEBRSF0vsliZJW2oA2H39hB0ZAtx4lZjVlx76Fhw
XqeicqeAxnQYJxGkIO0DUJElxOz0zzd/3XTqwPdyxuUJmNo7+g2xkgnh+qJvUHC6snygGRkWuAhW
khc7Wo3LBQjvSlTsrtawJVUob+HR7+as99KgOKHsACqwludFXIXscLfnkl+glwKWUWE0mvrlUzO4
svREi8ECe6+UIyTaqhQYKFqhdDi7pzHO6PuUK4RK9jjqRDrJk+/xtUCg1d9V6qMtV++ga7dP8eZV
AOBjiSkAorTf1U/vel9MUifavzbCEx6nRqxSH8CIXUYsm0wtLaJsmyoVxCNH4lrkRBfSKfmhwx/Y
HLZ7A4URC30sslQi9OoGJJlqpD9sRYgDidcuiG6Dn3AirA6PMv1N0iSkCayp4qUXsXSxkTP3kdVP
WaOgaR1EiA8PeXuMH0fTkZjG6AcwqayCq82X6zrzSQ379RL2e7bpu9NONc7J4H3T/R49P/ogWNg5
xXh34e5NwSabBeNGJUPHzyNBYBHD0i10bAkRYD10GjfmY9TY2dA5ib4Zpv2WS2i4BIDI0Z79s/2z
tRDyK8Hrq1QdLCxQtekoSYTpxsjpgreMhp0YTBoASFENn8mV/1QlY97pl4kR7OMSVAgFjjFpDuix
sZk7MRJK1UA6lOFqlHYBs3rsqFpzTSBpD1b82Qnzhz0Hmspx2NwqlTAaUdMX2egPNZAZcsHuZc2Y
pLCaBxJaU8ujHSTlrBguEvqPuNXXzPR99KTMyJBcL7Zp/PjnbnIqwr+7T3IHtrsLLAM4S9DMP5HR
Q4b/X7GN82usWHVsFfWnImmafWPNQ5a1Vx+I43+2uzPZfC7mes1OPssW6uGYZI92iLosoaZj9g8u
C6mjHbrepex67n6grwFyCos2RrZRXRbFShhmjhJ9pjm0Q8tspYUx7AcZeK68LsPHZeaMXbqu+ai4
/HdP9SmEiGuVWHTeUBkDYWyiuXPciLti9n6/OOMCSNwOXVR6cofmQz3qszfRHt4FgHtgVgOjHwdM
axxaZJUGGbHt8QSzR+vI1/z5RXu8wMkpYjgwBqVckAvKt8jtVTGb+e3415tKckCkuEG4nvJy0ed5
E8wzHYpDMKFO5bPZyjn402eUdq2uaGAfF+f5/24D2iadeHQC2PWl+2WoPeR7j6t49Vl20CifbuHF
ApkldoJ6VHjIOhZS3bo25+gim4kCWwE6RxDwNWTBiSrA4GfnSVAlArbT20ColmxyGxiSAElw7lZB
IgNn/IvCtme4y4kQX6enMwa0Mux+8rDlNT8LniB243KVQ2paP63p+Ddp8gAghiKYDya+nZaLGtFg
aJhDsVgY+OHFsIftjfZstqtZtfsnlofAnC00UO99w1PB3hDq+WbINy+Kbh2wXqxKBfvc5MXXYUOj
pHKU5zDqyaYm7eAvDggnJmunMCE9W5KGbwSdUvXjgp8pEUe7xhwCwXCFUad61LIjzXaM0Y7XkkBZ
IKHVnjYfw4RYve3kUxKUHHK3i+m1j21BmvGM8DZ9syVbGFsdk0y/7oKW6Cx4Gc/WD7nDVMyOJc8N
LM5Le+OrybUjJdiAdovBRqFXphOKEbTgsf91RKx1zI3YGFxFAltKBMvVfeAvNT8mQPhXBR4IBFQa
y4HlsaJoq3omYpjH+DwdNER77IlVJRCZGBgmuKGM3Tjy/ni3tSbT7n0+I/U3i/zF2YzsYTz99EO7
PYMt1kgLRNMghhtLVks6ldK7LX7Vf0CKsVjgRn/HROYt79BZbEpRJNQRQip3LeKgHAl9C0kEmUxr
tBDKHWLn2K9hTx34T0Is9T0yDMbGCq0VIAJZMbO/fWAaBx83Qr4q7mb5iRUPvANzRnyW+SJqG5VO
xwk2msgK7ANQoNz+dGaomNB7RPol0zt4UqADZ7cXWRalUtojigzR1vsbYlv4IWMjAt2drS1qdpL7
eP76Bo0pTDWdwFLg7s2lIq7/DhjKcXAaAYibJFuQ7bS/yBjhCxmMghTNAXWNYkW+E2XogLV8wcC9
0nvb+6O6HpTf0KRzKsNlciRWKtWhYY1z9YaO4keUBi42aAiqmqFLqwmdi+3jUbMEVO0eDxJx9qV/
U9Xt2IbIr7x0SwoPY3OED4sMPR3/R0Wv+RyDfneF6T5wWC1eqrN5/zaxMMuAy/7Jwl4nGF/g0mPS
EVLzgAUVFTdO0UfF/f9EfRRJbJieNUTla0TPTj10gR6EQ4I2kSy4QaAoA7T/GA4uT0/Z/g4qoS7F
KqHu8CcUhgKcRqKK/wORy8TTb7DtJpXD6Xre2x/qJ5isNW+4Go6tp3E6KJv++fN3DOTPebufwNiH
XqKd5J0CTNcIJyMqxVxiF2A9jwgKZEarz+1jBxvFfLIMbQpgSzvBPSCCWl0vPhpbT9abyJFjB21J
IYSez3sOU/Cr1E97mu6WWhP0LzZoPbGHfufWF0mYhOuEMEl3Mwi+7tCTmA1+U4J+2d8xcAeTWrJZ
OzFues9uubUsd+vyokpYPUQQaTI4O4oOrCTceyuatQvdWMwnQkaZnMcylrL+PxfyDt7h2U2x+U2p
kz1gKrWGylWJkoRC8eKJjNE97wctUF01UM+cOfU3KC3J2g17iRxG+3T8ZARcctrKp5D3CdG6Img9
eUu56+/pD0dKBhLm6tKfzg+nzFBcZJlpTPCNnY1GJlErJYP8/nfIkh6CHfZQe/wjIxI/flbrTguO
95PakkMYB7/xsw31HtxOB8eRfXAkZ3/Ir6yLf/v9+sNLPA+uyHGsGBRnmoOPuV5DMYYL1DCGUOge
e69R8h6ZwRSAsnrP8U3gFrYt2qsWoPNlssOxf88oYugsHvNeIcWSCg20fsbOFc321p0Byrpm7fTd
Ln1jWwZBgXy+KQVhGKE37p2HRGmY+TaH/UlnfF+2ItufvsXr6zJtFoyf6mgRiYMH3bYeR8GCI3bx
O7ogQ/FdfulfizgltrkVJM6+VL2b4yuowojDZV5rY2Nlpk3jrgWjNXO2B7iWzgZXkRJ6z2pL1o2z
cSZlzSXCzALKT8e4GF+PF1a5U9Kaogm6dIAz3eMzAJvWZv/5WDbOQ0UZH08vKrkzeutwZn8kDXDd
H38CUo3WIW5E/YfoYuhNbCxSJXX9bFNZBGkSkH5s1qBVzPolxYIOueQreKMUdYN+ev8UBGohGF8G
k6ztZn0yg0EOCQto159hBR84iTX/gMnZChTuHfYzgiNPf04VbknIIqjvuEsSy952HdqP91g+MCDy
8W2fgh4aSKNkulfI81Xl8VWJf0pOpRuUX8d7vYWf5VQXQvdaaNfDhaCU2lNcNNdg4aY59NVVMMi5
8yiNifX4YZuggm5kknHBBeJ+LalsxRkkq2yBywjUOnNsGGdDAIeLhTIlMngdQdWe59/Py8co7e7A
8122vviea2ZTZNQRbDUJMmyW7kyVsb8qVm6Y1gALa97sQgTeCTEE6qa21QyaDhChR+CytvL+qn2g
jZV9zoKgGcPtqtiJv8qYgZ/iP1muezWXZLLU+HHXk7dP0dprRlg/2wuxhe67XdGBAAJTwJVoL2Cz
+ZvQLII1f0kmxWmFM4ueGLRzfdIK1Ppdbw745McGPy9uJUIwEPN6y2d0Y20TVF7C0dCmj7hanAHE
E7++JA/ouWajIyJLOPiEEy3h+FbGeREHjFpW8U/YdIbzfbE8pKHih/TbqNkYxbV5ELPpElvxqQxy
PAd1LPx95ExfkHcYxU7FBZs/OdnKCstUqMY70NoFQwW3xTz9sVJm29OiFX1MJ4SkCSDF74AstCq/
rbuf9xVyE+djwIjnRdJMcZk/drlqYg1MA7MkyE1fhyQpnntypvL+QeMo8P/Ric5SW5HDDueH3X8M
QkG3l7gFSpwdbdIERC8QpvYsJIRnFJ0QiK8tnGf9/La4IwtcDiGr8px42hscxRCAkTQPOA/U2q0y
Gcts+pnkNmhMyBd63Qn1UNhlhVo+VES/cPDoaEuOnaQq/eOGQsDqHFJ8xiki9MocUUAJZxk+3v36
CCfWo9CuJb4qfaTj2cbvhN26P05D7jseR3My3+bVNxXJhAXIGL+sGX794eDj2EPiW7lk5JJm59R7
YC0CCgAMJ96584JFZesTebux+wVcOP/pGf4yJ1RjUjCSz/4w8s21Q+pxtQmsaHQ1aSb13VFUOeiH
Tu5y2o4Ze4xndtXYMR41hJYr8o7S7UxmwkDXa5USskfKEFrMOQfJ8QxAcu2nJAoCvbEDTQ/u6AED
zA58dil9eyCVbUsYKZT6SeTs761VTmjFAqGPVNvTCnLi/hq/7f6tpdILpxcoQlQNHeSXZ4u/NnS9
AhhqQj4tX8hnGlqeJdlfu2GQh/roumzR/cggmctNjdou2xW0duuVdIXNhBxWKP/7FaRwQLAatEJE
mKWl5n24yszlKKOFifwlXX21zDb9ym2SjwjX8CP6B6zZa4/ITfO9YLUIpu64wr5RssSVVQql18d6
YmhgGygwUaJ8fdDDCGyfiocY8t+hNyLx1/AUDuWHUkCfSrzSs38Z0kvXom8N2SUPv/Jc4hyuiE6J
eA1G4iNH2G+lGVQfCkHsKCzAWBj1IIakQMU/I6lVa0zPftfkB6Ed1KSmOSELvNKmRtkbRypFaftv
ICtTfMUq00HTCcIIYDCc0H+J6V8yIH52tPc/448E9SL84M9AR1DaqhWmbLhiNnWHKrPvhcnCEd+H
ZHXzV3kR8GjdCAcVn0+qkW3bni7o9NISdxH6gz5NZtPofWeOkHIM2uIdkDFxH36Qq0AXjgXihbax
2OYSse+l1cvdlY0Q9ipWQhktr/uUyvpRZmZog5DQqxH/y8NQXDazcz2krH9/OHgiQuCY2S1B++VC
WpAkNQ3l4bdUXzqrE0c9dRqg37/hN5bpi/xXiX/9akK86B+p3ohbXb15BUqxmZhPfD000iy+bKzL
kyyFhwEszs+GqKQAxrZeY7LU0pRIiDU8mtMEM/nxyrki+hZe4YIrLxae8IXw+qfeRiZbn/diJoVv
WaReKCrtwpZtSCZJqnMl3RFUMXrySsqMb0jlOonfu6KmnJvVcT3Ms+NWD8MH7k1bxOQQR+pRtgl7
8BTcaSzxKh7BZaz3GE2os7PXE8BiPmgkcHn8aggubb/0CVTRuB9z0VcqUZU8LIlcAvzvtJ3diHHX
AkO0MvwggaDJ5IzlNSTIGL+bqbBfhiZqs8KNwXgGxZKuDXA6cBfZb0/OpUjwOs1NVfpSpjI8id0O
XVfT3+9qBm8r3kAMl8duS6FDCUXjygoxUPh8DSicvbklAE6OB1o7cSw1VQ5zz4W2dMoUIq5B2Q9f
qrsFVsyz2RL8CKnan42Ra0wCfjZRh3rMxu+bKMRp579oZtjLlB5Jy2HO3/9fuBMjwDmSz97LKZ/m
4/s7g/79reFf3j9vjx5hi6Yq4QWZI0aujnnGBx7La1uN2YDBtTiA1hcp0M2w5XweknSDQpLv6Iyr
dBcMARab66yvDl/0QsQ4ycMBAkVyK20rSkrueux04RTPf2JufUs/TPnwUHsT3G7J+dl1uwczFlWp
8oWCDDFryDUrQDSwRqOer94M8Qsef2nOC/TlDht30PJzyrX3vcEgn8tPWsPR7bvnhQp6bTrMobyp
q8/Ozowpy4PoLHt9bc9dnVpxnkI9E+TZ9I0MIR5LgpSMuFOyLePi4vCS7zTUAcw1+PqSSbmsZma2
CE4JHx78Ps56nP/xuvAu/4F8TX2N1ofV5iFnfLlZ6Q1Ru6cms/eK+TW8G6Znm6za8a04wkmPTQBb
m13XUkzNVsDt947CZvQVDEDhx0mH8Y7WAQmy9uNnd5JSM6CAjcseXYWqZYJNxyprwUB+wxDsWemK
MXZHdG0wZAXCTaffbchulwkGoA9S0VU+ssa/57y6FdAP1Nyr1ulAhOWzIPvGktGKf+Xo0HeBG/ki
2MHYKCqRWL+6PkvC6rUMHomfZZuwsVD++cmRjkjeKNjWbN5FmCZKczcW43nRiKnqSCM8YYiRo2eC
OvRM1NxIRov5myqiike0QeU0Rsmxz6xq0oSm68+pTQF3QZpUYQutvJjPwZR7CBntBOrbS/Xl9hnY
/aEHpcB+8KzbCKItAWNt+37P5pklE6ED5JFKlPjSdbpcNclONYnvSLKnmy8KlnVZESekIJ/ddfHf
8c5Ai8BHPVhTODn6VNpHmW1w5di+B2S5A/fdf9pR/SaQAmmQ+5p3QHCa8+/8qbCawJ+yfGLUSAAZ
pNBpuHoe7HfgbUKZ2RyekNpMo+w0F6klv8rofka9EbuOQ7mN6Uj3PJnGtbON+EiA+djuxpMVv90g
hqFFLBo4VRik30cH2O8whGJllPRmctfoOT1kheN3ESU6+sIxf3SUjg7arE+x2XMlVXsBkJ6IhYRP
NwGzF0Tt9al653hguBlu8eKIQ6HxDLDcS/7p20gcc/VsAUojqhiVpfeDllcsnwKaFu7evgVbzKAk
iFn6y2kHZKGso9Y3FfgZb/Q61SA1ftNLQ9N1cE41I5vGhjB6xff7xImoq/My39IMzZ8qwO4QThNh
uoEb6uLVBWq3AUjhlLUKrTUrM//W7M0lwaq5dblRbQSf2SWVj/9/vkmViOuK05ldoj4+tsG8EnoN
ugtlpl0asPXV+y3DXjPC3jfiLvXGqGhNF9qx6iaTay8XguhYo+LCY3MDzxp9do+CYu36kdoHB7wG
vVKM4UkpmUzxrr3aOFagEXA8PTdKHX2OLxb6qgEBbelzN1KnqNGzYw2U4aYMwSDL2gFteECrlpV3
OeNjk7V2wu0tlMlhD9s5Np8ucwmM7GBGJySvtEsBxSQQLiITCTNlk5D8pws73aS9aRy9RCngKU4+
jvnvKf/DiCtm9P6Mtbzu1vhtEg1fSxb3HLoliAmyyF2LjogLGBfj4tXNq1BHfpgiWCPNYEs1/eqG
rVl0C1YHUJiGRpL/Q3sIO3gFRDIlswa19y6Cr6iBxyaAQMvar+F0mXbl1JUWEv7CiD2TRJd9Zjs1
BrnY1AENAap2zZ/BPG659ppf8ertfrnCzOP7MXjMrZban7cQ7cNEYCEdjk8PQhDuSknYgALhFqsD
wjprUrTiXsqnmbUUg4sSvVmJTzwPQATh5SJIwNIomAjIc0D1aBHJWLRZ7s8cHw+HwPcggvSAUYT7
EM/XXct3Va+FWBiKp/t4xpgTOS8nVt2gOunbkhB5PiKW+p4C/Z/tzkjlvhz9FHQzMQc13N2t/l+f
V6BxFr3Typ5I84ha/Qhbe2yr+YGGz5YmIiq9fdWCJY8lKXEr6F/DwCnminvNftxVuKJOBBA1RYmR
llFPfvHdUzW5PrOdx4bwMszlSBKpn2oRqJs0fNVauluf6Qi/j/kO/Gz/EuYhTD8WHvV0iF00jq8T
T99v7jN9zqVnUVu4Am8mx3PDFsoJex3vwxkNg4rav8cSgThzNIpzeKE9TL6f9wHLpiYvC4KRTK1e
nCL8JbPEXN1ZT30fV+8ViNyGyUFqe6ZGvvQ6+9bSnAj6ok/UY05lIu3BmsZfDEH8rT601EF6Ya+r
c1wubEJQDKG8agd+UbINdeV+Yu9Q4YdUap4XTlDjT0741K5d0AxJlo3H6eljqfj6c4tXcmGhZkKU
sgEd5pJtK9C2RsthiHqjW1uQDeqQmi81OtWaSgkur96r+z+jwsigfibacjowi4HA4CqTqNfcIyyP
cMSIHovFJGaxsxHyTOrWjSxHcRRSJbY5JMGGMdWC0zH995rmCg3gyOQw0rEUNg5zKk/n5PEeWLGf
ozmFbr9S3DJWYRfFfIjghoEfDRavMh7YzeOPlxntCaD31QADkiPZuXg2MEh/c+P7g2faMsWa+cL+
JYc5fCipXwXtxtAdm5yY9a4IXErcml3uitsFkgnIWiR91ocQZ6sHeIsyh2IRLEb2cEBLMUXqhG1g
Nz5vnHEIk8VOQ9Or20eMVECdvEQJFL3I81FsGR1UwqKMRILJ3+RCU/OJTLruWqe+sICWRAl15/jE
S3enY4SddHMp6dwYIPAjlCHY4J+dI1WTIGxWBY72/w8u3umVn5Kv9N5D6HlixcyGaXSlzesH2EGp
hd6d+o4B3ew+hdKcj9XwTKs+MCyYdcKyg0Cp1dTZvoJEBdV38N40NQnOak4pFNyY30t0lLTaLlSs
3GhNe1whoij+pWa+xAMzjzMMjM4FutOzHU9sc7O+1w8Y6yLxWOzithxonU7fiYpYvbU5YfjECYUx
9mOm3EFX4bt5uXX2EwunjTEKTJ0wrbohIC06eIdrfo0SUgaseFJgUsfRRnGpOCucROnU2Zfhbb7o
WD7LK9lI/G56jYPGZ7kbpN+1sTC0GXfJfgwAukiV0oDTKLWgY2D6JCh5mE26h+vM8dZ7YkiOQxv8
kxNmwzxUNJyvWLkqBTFn0E9V+zqWUqkDz4CQu0/HMeEgW8RkNdCcGj1rGw1caIEUK1uItuXi+Hhz
o3FVV2BFSsfvj8HL56/VH7QaW7g36s56H7ktrQiRxaUGIq1f8igbxvuG1kbo0v/6474sTeQe1Oox
3B8sWJ0rRSytEZK0JhQ76o8GDuU9M2gPUIPi9H+nNZyc3iU+sM1WiugrYTJXbIkqWec6ko69PAbk
MJi9upTOzhMh5afCaYFQufCtE3AhchzA7g9Du6jgL5HqohOTUdi18xYVLLVJxqlaD3n+QqR3q18Z
RaWLg3IN5jh7a78lZtzBKucHuLIt4usF6RuVMtvB1yRrmGAKbr26Ggc5obnMYmopYgPeoeczTEVp
eCo9G+jD/zX0PthGRf+HEzK6R+FJtWxVMRECNzgXaFonzUlCpXWZy41kRVNwMp4KmSO9YzB33iMj
sVxl9WJCBVNeCrxABCp+Pp9wDkYIt9doJ8bmQwIyrFKWSlMc4vEjgyXT3q1lKjVXxeAS3gy/fhMd
5s637LQN6Sp5jjGSCIveTw7AytyRMURBaeZWRlvpfpnbR/1SpzaGCQ93e2sYLXblyCc5bl306+/m
91rJouGSExIOyI52q0ZeHaf5W5QLDe1G0VeHnMF6X1BaJY2QrN37PvwqoSI6PBVuIDA06GSWNQfV
HViGGBpl4krHC2ILKnT+MxVEzBqTumVca6TmFN2cFuDOzUSNYaQNOe83p/DDjVKCXuS9gmkEH1zv
jaKDiBpRScqWfr0moMo1nFr4XZxuohKPvgyrFacM4SFGqsrg0XJqz2oWiX4r1c3HuiYzBN8ds9sJ
5TgarCDJFbpNR+iO7pgaF2lew3l8xSGadIDiHWLOuh6qkf4G+PL7zYdsDOY4dUZsEohIpjeX/nbC
pxRnmFsH/hDqZZyKk819aoG1lIO+O/BiSC8eImySchRH6Q4/nsuCFlfY9TysUPs29gdqeZioqZPy
HFIOFsXY3QKB1wFTm9F1jYnthgTljLbL8ybsv2QQjFe7zMAE/e29H2S7f+yapvvVzjN+QaUgIFht
Idp8VFbbbGQRtna1TGDY5bRB2Rv4PFusOkstOKt1fB6k9O+NEmo+HU9p8KZj3dZqRGDV7PRddsJ/
KfY34lMWeShAkgpSEgS/+joai2pEZCHexPq8YfDn/9gCXxyepfft24SiF75sQUmuiuP2O5Al4qsz
Jyjvvg+jsojJ2/5IB4Tu0jSVUm4x98u0UeOP1e3N1bjy0o7RuvStmB6EORc4TlI6zTi0IuDzaVLQ
qHwIJAsd99WXILex5QqXIU8NQMAdahcF4MJYy19GCWZASqzr8GUblXlhWeoKZkw9sI2le4CR7ZeJ
jouWrNAX/sp2m55bk6v/eb2pcl5+SmxCebgGO1kgxBtaLmNq8RMkJvcUShCN5IKOQFr9ycBbsHnb
ejF7Hj5FuZeAScmIBlAY2LNPSSQKyrIG0sCZNTiZ6AMDWKtmBfCF2GjOfNdXt054wGzHCysrs7Vn
LC2fo7FaOYdYISZUnOy6BOwCZYW01TQRcjNXQDOmaGFmAUpY0EuPxEJZOUiIr9j6BesQU8hwDO/K
3JnRMcDw9ZbEnlZakwTwYl3oVM6CMc4NAV8moHxPXqQyUfF94BACS7Bi1CKjqkyNJP9PAStJn9R/
pF+1uSBmmYeZmj/aCLCNu1t9GTiDVGs62jKseDQleXzfR6H2Cb/zkcYmnU40gDY6xXn8WYdpqDxA
Xueqg69GHs/i/Y2WXylDceFXM+rC4PHgaTkbE/cix89awKJzAEWs4xaSn0dtfjpdANDK2WkILO4X
lVvkgT1EcsKydIYlcrLHAiwj3+1QOXPDxfbcjHtUZyWKsWP2AhJS7pUwuvGT+LogdWubELTShNaX
Dtmk8jNlvLRhzc9bNp3JOFMcaMMJ/GMFl20yEtEhMjLSFFbk9hGoXnpxk2Aqyyp1PGSqY3bzXbWQ
7EWDBdjr3Uy8QppsRxj4LE/MXcSgo/XBNUR1QP5RfZ4kGYew40nTSQjas5AmEfelhMH4WhdcwfU7
3NLS24sRR8t9upuvs943EksSdYJaa/sBeY/Sv+6iEpRt3uwhoXzfQzCi6koMpUOMcuqJiX6NBIYm
e0FFeauyE/cDdbB97SCGafEwlNII0sxrrC25hTmXLu2rPoQuWCni4X8rS4Xq9x2E/HXsvyInA89o
3QA/mYiUVZV+Tq0EQCSZ5Qm/C1anyaCTeAUsEbKw8CixNDl2rRriNgvZztJakPwQekueZdV+ZRNS
tWgsgQFRJCjZKOKjSyq1sh4bjHduOK+/8cjP0vaDzYU88Cu+bo/ZYxNi48sdf3SlncH5RxEEbvzX
6KXZ+fksKIzP9kN8kjc2vh9te9TWgSV4Zn0XL1sVgPNCOwOr3Z4ZEBDzn0CCOWZOeLMOvSb24jFK
aWMLN7kn+8qHKQUa3wCnA5rYkmo1uMMI85YjQ2z164fDURm3QQUIcr8jo3LsFD/F9kOrBq0Twlzy
QgQuw+NuhjA53dy1+DhTBYu4whGCOKO0KDkW992V/eGsiKqJPyGryAco++NwBDWx53CRmed7WJZt
rw1FJli6kM0HrjepCBxezVAXzy+tGl3R5CtOOYZCZlOqo5tGN4PEtZFV5AN0BM6jWuopk9i5TlN+
fbmSCxvMvuVWQQcQw9iL/g2bzwfPlmFnUCsYz92kRbTjzQId9XQi8m60voBTN1ymLlwi8SXejKpq
9ycZIrOrJ+kLXW2NyowGIyw0bvvi1FqQtKlkYbQe1W8zTbhyij+t37qkim7WwBRdTqFdgtYnc3Gd
N2h5V+HTXv1GuOhkCNLCehhO860nfAmOO5LgIue3vTV02SUxq47UvifdkSCZKLjNQB5OnVdxKkVD
HpYhqjA53L322ozbX6BQc76SsPK0oiwzWGBF1khynE+WHHgslA5bGHn9zP+Hmx/xTpiuXAK0pQeB
PKAD43fp3w1VTK4kXPcpNIBr62H0/NjAkkuOKfgmteiJnIiK8ydmHsh8EXyS0YcHcSOqYfhoTRg5
OXuTd0FHQrKYPIv511fDGA7+41q9itH1W+2Gl3kwMQ+qn1IUeizeAFRkpCJMZKXAyqPJcwfZjcDO
EfAaeJUITYiQ/PL+7GGBJprFxkAk/nP5Vjy14ikh0dWrf/ALXsX3/s0WdpxNbIoivtOZf6BjvDxw
98DDq3lr55ftc35H+DreeqlRkTqbaXdQaZgXcvq8dhn3NyPFi3RhgmBhtrC8YiBhSSDE37HvSzOG
JUtF0BA0WI01vwnFgx85MXuU+y+ZyexMPb9q5UM+OVehyA/Rlj+v4hI/dPOiW0PTeF7AoRSmp4LJ
XVRpWwsAkFCBrDsZrk61iMaijKXxxHxC7qfIpYdHNIGXaVNEuiyizPclXauSe9cdu8Jta3/dV0JV
f8ojjPrVCMEIDzcf1kMVyddqjmnC5nX1eLzvJEeglCmuFUc+VZnBtBx/80QwDm3Yu1du3AzZ+Ix1
elt0Xj8MZ9CTmEd/jN/w5Be8ZWW2W5jfidPzTVBKYjohuBtL4iyT8QUD5Hqwmpmsl8kgkY5nIxg9
NBNdFMuVjKpRvfDnKCY0lmgqNHJ/pYKl+4zhEtfg4IrDToklgfpvN19BaY2QWcU187GfYa3mROqY
8+QUs5nnrial4l4zJH78w/n5ZeXQ8zBp42Fo9WeuqxGANa2MpGTbx8gwEs7yfXJOjHy4KSJrCAeM
vmfgSUMCfygkiluvRR5mTN16OclpaypkuuzVOG3S4DU5ynvmKZWrGdHzVNWrUH865B+8i4mw9J5z
LZ0ui0ppOK+XzZ2TJzSANbKJQ5vobzlRloN9do7Ys+WCaDRlC8kpwyWni8JNa0dI1eLZU88oLwdp
amhvhPTxzHGj2QsRilb/+rVsNC6jfYwYES0rUd8hYUjiVlnsoOOoGb9mjuv31G5ospznBpSMkGeP
C0oeG4iwfI1zMT0DCo96Bbqb3eFm7/lZAoHWbfYa0HRdC1Q7nJ/aleyqSCw3XlD4zt03FiYmXWnL
D6EuSVxwDJLAkwkULF1YQ2tQT2ChXvtxzG82yX7o03kYj+v9FHGVt9L9ce/jRe7mRGXQH8VgZTQF
Fqpn41Fx1mEIhV3kAb4HNSOxOGqGWXbqXTPls04EWe9T0lUDQ3/iP3I9CMvTCYEg//UUtVVT9QJ9
v9OTo2gab0eEh8F1XrwfuSNTbV9A05aMTQV58ADSYG6fZbkM36Pd/YEi58A/Nvc0ELwTEVM5f1b9
Co3PpxrCR8t1xsCwaJSSjpTpNkOOGhQR0eLTnn5GKrNdPPNWoRIyPLA7EBt6H7wS1MSvfZivppzr
SXzEE17epdIq/NGvjsfyecKdbJie1kKeRAOqVwCpvSujXUoHhgsBabqlR3j7kkm0scdh6f6rZ5KC
q0DxlYHa8OD4nBRQF/0oXBShqAWiWucd8XhMF/JkXvON3xz2cgtjmlRFtLmm0ojn91DuHjQf7aQW
rEV3/hJXLwtiI0jUAz+iYy86OOCXoNM/Gg/PURyw89y50lH4Cjp4hR8oD5NQd2kCGZKujaw2N6PB
ztg/RyMiTvRTL3L8Os/LslNp122PNLj/eqWMEktbA6LmAy+0svxg/Ufu64OUDIy5VeQ7pxh5ZL8n
MDnjhDFpJIoN67J0yxzgon0wdP6wOpcfV4NpZT1O0LzKkwcXEEpDgTeVqrfcQXRIHy1iu+1ov8l/
YqUQJ6s7cdvBdBGR4cLF8m7zB2Ib3GxP3II2mru5eOYYLJ6KDIIarOxpJV0BPU1arcFtFJrlOWer
2pX81jePhGeMik5MPZHuFd4wyN8kLj9aK/6174peF+L3X0/NdzX9DGN/IiDxcQf4ttUl/Fk+g5OM
utJov+1pQaAEghukYEksXp3dp8UOjMKMy/iqoll/oud0eY76YJoYN+qP46wFny8bQsc9dWu6FD5C
5kL+mHo1LzS+N6ov/MwXWfj5KMnLZ/jYxpposJHoO2AZWDexOAIZ8gBYsmIsL4Pd+xpln5EPJqRT
alriGeaU3LGYrpeNMtoIBShSGJcfaVSzI1sFvoUR6J88fh9ziGKDMbSDBPJ6V9ESuqHO4qUsTWY5
yPyWLMARvDhVVSxhNXEJaN4ydhBc7buIS9baL2TwJ8FZQuTm4Zd7CQRvTYJhO3uysmMwWIVobLA6
Barvpx9MNw1p8kdBZwf9H61GIj3yZ6D1VHHPGmDdfksWg+vHrgmtb/+7noB4Wg07WE7rhP7w3u4z
zhs4fCsjmd3cAf+u023rgTRvoPua3OzSZX/D43yLkEg1APvjjwSMO2lIT3vgfB2c9TeIDou7HeHw
WYs2lEfvq2OAlwc/XBdtElFhd9AuQYcYpGPV2G1FgB2aNaQnYdXRfrCsH22QuUoPbjs9vK7BR6yc
nRLqLM7bj2yoTF4/wIFc0B2feZilYBVOU9FlEQ3Tc3MDmdMGwA41HUweuXAPLL8JfgabZhrRau+H
YXA6DtV1dhcFIdO6tbz0kqUywhYwnKRxmr9m8zzANQrpwo0A6JK+Ni+hA4ylpLkkEMTYyYuyxn5p
6K8Au+1NwedizthweVAII+SCBRAjAgHY/kT2CF1o8YfSz7sThiVXjS1uL2UacVFwON7OgxkRfP0Y
snZoEfTnroGnUb8LYEV6hB3crCtpfro30TwX+oP8p3r6TC5Vr+yBWltbGUqmQIQ+5f4WwYn72sl/
eWmdD8TFbsjvzDozYTm7uu/LlUHNVj/M3N8y1DQTvKrPzOoctnudBnY8+r1+/DK0tSTd24how9Sg
QMafdGMAhncUJattzBNL7q5OO5PPeg1/aFrwF+MQO+lLXeG0imRmvYuh0oCWcNT4py6KNauodqOs
SR9cNTjqzFKmCkEZ6eEEPwi6yxyeDm+0a+S5w52HXeBDFcdkBbGAQkic44McO3F3eMqQ9UNRHrbP
jJcEkD0YciH9NSRYX0efVYOJbzVyYLXoW/vJ7evvSjERkHXSsgKDE8A04aC4bcoQlVaywTh2AIde
c2KY5kWcrv3r7JpIW9FG13Rd+oW1GbCm5Sy0+DEE9ZcqforcBipI+lGKnybVN3UCwy2R12F2fPlW
lO30U/EWQAVesBOtScmmL50Z9UkYgIXbpA78sIopIHVtrBf7CBmyaggDcvepx/T99oNcMlE9JEL3
HR6mD0loJtBfFA7jUK0Jia5ZkpWMv1iycPJQoMapbWvGs5g3n7xckPgTCw+G8p4sQ7gwf4DMhagW
B7kUq8hzmm+9SVw9HttHWXdwMnqicVCgJOMvUIdaYVuMSEaGT0mvlkRo4GILj1Weh9ba/faFqFq7
ygMT65DzdkVRTQ9nmi0/1VJ6DxQfNu82bV8qoMO1dLWPJtx/5boDreF27WDvNI3qy721Zb4vOH/b
UsMh+kcUrZUXlVUunDLkXTln+CjC4mQrbu0zmQo847DRvaAUDfgXvXGvNeDh90tTKg4ZPtoeO5+P
JPEodBQL37/oBqSvDzad9GGFsnzr4RCJnjtB9xyKoRkOLPBeDmQ3IsdzWk3wDIEk61Yy/ZJ5Rqp2
gsCgJTIYMCX/2jzTbpIeaYc+FPRvqRYrnbCMAIZ14Wb7oTKzDPKC1VY23J02YBGV/BbAi1+dTGss
GVi4Q36rNoQjGHcVCyADf8/FJqWVp2+gu24MyLpRCnkvzQVJEpu5mzyAjzzBv7VPgUGjbcoeQV3O
qW1FhVGQxFxX/+5Z2omugrnaqtp6Ba1e1luYo5sr5e+RGnX65+eXGIxUNiSfT4IF3uB0qi9lNwt6
R3/M8RqSKhl9dNMP6nSKuD5HqIY36DZ9q82dTNu3ZNEujmRh8u/g6pKo8WC4QRueV/BFzD+zJlOu
qNPKgZ6BXBhyIMcBqaxqdtqGrs5rmyoYYw1FoeI69cbA1nyao0Oc4ptBCpuOuWtDvFN7AQ/XXoyv
ClyVdbv8kkeQWE2xbtPuxQ3lw3huopTb+ohvPkg87M1pGSc8fHqV3TyxEwEnPktb6oLL+D2TENBO
fHACQxzxxXijllUldGYicJSzfmV1rldSx4D5lh1YvXzRoNBPT0oLiNGIITc/gqov1c9DaLwGyGhL
Vpc0IekYYw9Oun7xzI4f8Ia7VgFrUsiP9/EwBvfhfBt8ZN42HTW8jqnsSuBIxPHtYW8nMXqhyUzY
dQXvHB/NrAF3vtLino0LQ1xc57gQXh5GQGvJNAS3DFI+mOPEN72eAVUBN02D7yaq9BWhYABleQz1
N6MQAm46wh+T+OUHHQbNEkF0GV49poANBsHG/VWWD294Ek1FdvugHRXwoV1+gr0kJPsS6nzQWN1l
PnedxECklAMEWYzb9jkcnKa1eXfw2mIK2+L7E9c9UTy5kIQgySXmSaAS7NI8FBjiGxgA2bn98/Qj
IwAcYBVVb/q1GZaoePUv97S3Sl6d2cKbMXA+FSf3r512if4RYzE4ABfamj+T68iuzBqR6uECSfYg
Dap5RxsIzObEZr45yzcM0xziGc3GYLUktpbhuQQBcE3nFNqH/sVWEVZLug4dH6C79qnySzXzcQUn
U+wDL5QDkWOkis2KSOO/T/CQjzrq8f4BnNw0qeCaJ7177e+paA+fQSOQHQFdjNm9muZPIC06sREx
heAB31DxT7hIRf053XFn+7Dmpo2n8nZ0WiTmrg0cjtqeoEYdOFIuk+oaBWsr5iSs8VsQm9+U1Apk
oob+HJAHTmF8OpkLbgeUnGYR8xogZ24nyy0N3psEUykYQqOPjRw726hyshFNLAtwJ7MMuXgDeOZG
hCtlqsd3R/szxbKFwjKW6KiIWrZFuz1SWrAj4oMWIeLlvezRuT+0ouGavADHv7ux0/fHqY7HqvtE
l9AZJl0UJcx3kDPSocvI7SRe407+S/WtQgTgwgrIshTt+mwo4bmJBx0Hr8zV4YHMQs1Kux4rlatJ
GPft93iX/N8txmoK8HutzpEoLXCN4NOPMQTZBYbrS0p4gw4uLEU1Z93nZrBHCHM1s+dQpjO0V13G
s1HY3PG5oFvJxsLJDn3FZl5rqaxmqpsUCBqbnq+z6QVfqXSXUGa39qbnQlmieLAHdaR0DeusIJLG
jccqlfWGHmKCxViypkB7oBGFee3WkVWH/6I9+lgSfI4dShCItYtM3R8zSiilqqLk1WUot4h97Mvs
qcwxMex119onAI8emTN/1TtDSEmvAo9iPiv9oNCBATM5mwjJIHj7VmaJiSENImTOseGbizNYytB+
aHHBz9cP3U5vVc5HhRbHDfyueAz1uDyW8s+Hd5SgZhSVfemymuCZ5EOFT1ZsYM+g/12osURNzI2C
bvqdIvBjmE/f+pSYI3II8cdlzLNvrq/W7WOaOQoJeHix1LLj7MWdPCfYWDSlGpxq9NBPWR4zb7Ik
A62MdhlVVWg4KPuUtUzZwfyk+0J/C8Y0+0T4DEdkt4o2arcDeYh6xpMxIlhHLp4yDm8a4MjmIKgU
KLZC2CGLuZxPbRbcNxkGIm/QAwofpBIiHZxCARKbvO+nzE/AT52yI0W3EZvHzWqyEaBxDtK+jFKT
v15FaqGIQRCte12Smi5aKc7rp+BqLRdqsMyOW5Krn9x6JX9bQq72paEzeg5g0D2mcON3nJtAw722
IlpcG3mfojIwVbwXM7fh8boczwn/u4QD4iXGltm75DnTSdvJDKPZEq4ZhsLLbuiNq/vWR2x+UVO1
F0jYitdd0uc82hXgwQSMK0Dr4OCr17KsmTXy4bUaKfoontYnSvwaDLiWunJPCdvZkdxNMi/M0RZz
PDBAJQwV+V9zAtFUvRjUhlKtwbhEy7iUb510oGOP2AxuOXfnjsC+6G34iP4MN5NZEAl/KhBYt+WT
NOWq7NjJdYXzLwqkiOfYbyy7uUa+B67AutLZ4Xct2Q+vSQeG+td1fLpat15fuROn5SbQFlqd5v4B
osNEglJkRe+qMg/ndTlIor6o4jTirYkfumrkckRRL1wctzjg7ZX+gRqHLoUUltgzvHhECRwbVy/u
Dm7f7ulOitevovdEnNO2jJbv83//LiRmXOkn0qNFbn8aAH6l4FTMQ+V8L1gyg7xXUDZgmo+g9dC8
uKmm/C53llF6HI1Ai/VX3jxW5Lh62bAQczPhxwaf48eIRc3fiIROfwWMk/+xLLW9c52Qz6Ya4YnB
VgEGzRrjeis5WL2ZF0tNt2M6WyMk0VG10epWg6vMR6BvHiqK/WDmhy5ben419Fh3uj+hHdaVisoj
qzOhIaNogFmHvuqmjnmnQ70JCx82j75CJFA7hjDEJ84gFXjfMkdm262mzjrA+BEEl32Kxu2y1zcz
gF3OxHOKIowg53AB1mEm5QgMpSsPKQOceZX2qB9czL1r9xRvPBD79lQm+hoq8fHMk3LVWfCXWkjL
2mLfLSz3/8Le18lBuVR1c67x/nnv2S/H4ByU1WpZMhwEMNY1U/Yn3dDX1AsRM6a4Tly4BOQvdErF
4vfnjLFCmNyQfUGSAtWoF3IG5puCtIFFYICpPIzA1jokFpeEZ80nsL7p31nFV7/PitwyPTdS39PH
LnQkl42k+CMmr0Ib7On4RdY//2EO9fh28WxIQvqHaNpolOvLQ6uwBBo9wntEq+1yccercuUOuL9H
BLJI7X5kVE+YV1NF2jh3J8EPRguNFBRbnrvOM8pekI0enOqRA2FLlXdRkRsk5hGrpmsge5VFTbR/
NsTrxoouPv9jdahmiQmdiUY/cw3l/7FmqmbS0x5bNezGhgxtAbWoYGIg1EP10ORmAB7cp2lyhqYf
hGgN+IPaly61ko7KthQv+CYXzN3RSjxZvMWAf7Vn/2Md6v7nCBBFdtoB5lld8CjoQvCWVjcPfriM
nwectnai+3Buq2sj2ACAEmHi9/sWOL8z3nJnwOe2e8X7ye7nz8KWMyGGAUlI4s9rupFQKT+kLUGL
oI5b1jrtF5un9xVOCkfY1qjhBWpqTEccswTKVoePAnjNvAnDDjjRhX7C/ySt3nVfWHA1Bd+0Wbtq
EmOvHCtP50nv31G06KIuN8m+wuPzng9At95Ay0zniUmir/uRT4uoiTAV8keiSA1tOAOCkCPsShNJ
DdM+2OIGOjfbW+ehO2oJrAzEM9sAaBL9RSlrnAm1vCycOyTtshHwfwozvJL5z1m/kBXfQsB8CEAu
kfWIZ9BIQiIe1hL5g+N+JwQ20uT5/mId3oS9lHBOw/O1HhqiV1dmtNQeKCDjMpxmJoTakS/92T/i
IUMg3hOY8DtKnVl6YqyNKWpUbfqumb1nLQ8qtrSstQgYUCyC/YpvTpc/aK0a5xpkGjXcKCUGT98x
hcxG58JOJdfIlL1EkYJKzrjFDxYxKQRbC/mePc0pWejrObdm8nl43Dy1zpMdO0zIlD7oDww2luIE
rAo6vBsPNngLqlY+gvOkg1iF4pkeiQUIGVU2q4LGtLm5+eauCd2BTL07grkaVWFzS73SSSImWgyc
K8s0vP6kY8IyTSVw+MgSmO/mr+virRbXmF0B/58oFNV5pIjF0dOkH0iYAy3zPMjaDJB83f95N5gN
qbBhSq8uJ9kHDl1ydw81RNsl4eliRDvkPq2IVrEy3idHWY+GockZJSng4zOcXY2uGdNnSR6tzxqZ
iJxeZF8rR1BbjbLb8rT0b/eNTk5AChXNkpiXcuguKEiz5hs5B3NToR6BbuebMHiabd2UHU296wEz
VV/uP0Ec7BuGybrau9mNQ2y0+cl/RQjlglglCfgqlEx4KjrZOLDi7hjP7cKsO1urYEgdSw186U05
RONVrxvqQY3fUHZIOJjhIkul+mgyFg2GBZGDT33d4JR7xa2HReIbiGo2wNtSFQEDdOGGfmO5F+nE
cyuVxgww39ch9uptAf8S0zktuOKqo6nPnAMmv+8p3U1weVoGlBm1uqqpLAWtyycKwXIke9zIlFkJ
9Kz1g1KsV0MG4hUnZ5LgMsEkFY941r48Je/dZNRaxk61IFRrp6AZAcRTHS5qiWZerz4Ugytd21LJ
ytaYt21GIhRL9aKTJmUm9+tFThLjimS3OhyucdJKJzPpjkWZjY+tYG2OEsHUMspuhl1GweIS9/nC
jLsZ5dIzAyQhIvxE79DWyi8kLeNoMHcINZB9J+H7vwMXkWW4p/lZZ0GkcRsxyW9+ei3k2PJbF8CZ
tEa1jz2q304Xe+yOU3L2K7s66tL6ab4g00mm9+5FMmGvbxUvWDif0P0TBz7pdwD2ZoC134Cg+d5M
D0BUbbZZowW+r7xQWI1fhluSU5IlDIVpYHM5rX/s0A8QjZxXCH/1l6usjsyeq4hPF6TahdeDzOxU
Igx2GSFOAs9iA9UwkO2i+d5YivHHWFz5bKAUGZESUBjdZPFL2UvvBZ2hG5s/86ooS3+NFUefFfzN
dY1LU/gKuJptVecxmzPE3EN23QdaQPo37JkKxwd0fl3Kk8rwlogCS5QsE+HZVli22oSbIFzMG1k7
yAs4gF8YX5p1cl3ApzB7jyLBTYsY/Z7sNQgtEKl86mzA8Mu2cLsnJXy4b/Qwmi0kQmNzRsg3nMxg
KKov4y2yCaAE8U2d9+gzgfsovGN1SglJLNr996jjy7p6Xz7N6XfCuuoIhsA2ENlR5y/Gpsku4oz1
uysGjSnppFrfHAOJklPFP4KvS6vuFeN8o0FgVEzOJ/n8isNkmGBIF6uvdbrTUE8Fcx9XFgan9PMV
vo0fo/BBaTJX3OKWCJX70UDbval+cA+s5NCZVWpJrgK95/sU47N/0vULfFKctp9lX+5pUv0keYZ4
8Fn37JA7y0ynG7qb5qeLrMz/kF9mdmqhHP/1dsh5TRwuyjV1lRwg0GdPUvdYPxsSpqedEtOM1rUu
8+kNDj/L6W8KOqwrojJoMgn3bV0zAZqGqat3c1BjmSGO/FAtAZebkW7udMOiRCjbfrd9oA+CyKfQ
fZVVgYbW6T2/EaxWZVenridxlQcg9UVVDJRkhoM+DjZLOnNRiv+P+PyXQzcFvaH0lSv31sdyFBgf
8GizJUPN0WNM3pc5/e+rKXiqgQXEaDXOooOTLCXgSCo+WVeqZgSBzOSrYk5aRaVB+HzX0iQztwOd
fp2F3QAkYs4mc7BgyTDca/8XPRWHsPR4oHUOsx0g1G2Pe+zx/ZrXHJLU/OHaTW3d6UrI+0i6P74/
VUQa6Lz8YBtU0/Z2MUV0Z/x7CkT0FkDp6aEPVnsK6auLFBgrH/UQHi2B4fDb8WcA39gUFikAy01T
6H8BCBKLnJtIl1dshXM3wJh/zdGrGXeUV5E044zE17diO/VrH80kMefPMC7fh8dNfT0USwwucMsz
95XsOVU3naeS1Cqq2NNQia4IpKzzRK55m2bNA/ePsqpURqQ+tSlXVb0VIRIcJBw/WPHzyLHfrnO5
IRrN5hUvj4N+ECquWDp282G8xTyTE2bjoXOOWjAzhizlhGs5+Vjao1zs6oP0e/8bCRquNHQo7lI9
VSFD3xZnqVDkYAeUXMDB/LMrUsAiZ+K7U7hoWsu2v/Pbv07dySBK/d7o/7aG//gMdlJy93uRGx22
/ljXBdT9CrLY9Lu96WkkA3KNoX13IodstZLUDmIG7ZOaYfertyHd+1QjUHgNw1/y+H0C2VaKCx7f
c8yMDUfXkWTF3A/77DCfFdeI+TgNV2rNNER+bCJ8v0IfEokSmCNrCUuRBvB+gNXTVN7aSB+wwwJJ
z2JK3VFfWyPVX6sJWppBEVN0OQ9AGk9+Y4/7NlIBjfe2KSr6Lhh0K/Q0zLfJQEmrdq7GDOACvbKU
nVpxwItDfDmk63GLH8Xg3AffXDeT6MHNI8yFnf5GOqQFXHXAJuvZnI6J/bl1TfZhDC5N/Q9N2REJ
blXyTYR4Kwm/DK1kBvsCw8bRLZUW6+rCfAqi5gFOdV5HPrhFm2lmRb8X4hajn+1JsESpevpBm/lG
3qH3khQ4xlELZuOQM8QHTdcA50O0MVoIXLOf2jvw/4S5IRkYtZytdxrnL/X9zziFumnjQxtsF3j7
j6umVkK+RFBMGunkw931xqHeQMC7mylSqVxtOPHXSqsFRssNUdZ45CzWk+q+KIh0C6YAtLpf2sym
3giPtDalXdlwAmssi2VCCX+d5be+qSVyoSTpu8XtJgFWx/KLHpQ861tMCjBrmZgC7pGbKu8uA1SI
dWcaapuK9kKQNlAQ+MxQRngnJkJ78Fkcx3UoV0oOaERIkKOkUmUUDcKtJpV1CFUdGL6CgrhAxpQa
BmnL9e4bjyWp3lOaV5cxXMBvpljZFjZMMj6nRn2NUXINkit9BrXeeEg/PrEp3svWz+/HrPhQdFu8
L4TfI92c+afntQnD/NH8G4HRy1ay9QlnAN2THilC4Z/MZT6izk0CjmE4zjWSXegxcBoPOoU9/Iv+
Uh45QhYrMM8VmUB45tVeXlqRyzZP+RSCofU61uJ0C6ZxfMk1Y75K/BnrIqGbGjTMfdKVGQNBdgYP
d9byT3N14UgPY+V3vRCrB2Rvbg2TYit3Qr0AfH8zl+BOM36gWKEu5O23TxCN6yF18TUe8rUCKBcm
HJugQejnkzSo5svQ7wS/0UVhaeXvPY8mLqq6AnvB+Nz6u8UI+x36PnrtWdiA8NSezvt8Io42biyH
RuVxBH5FITDaBVtrG1/r/O7CfXZXVssVJC019d959emGxOZIyHfbLzHxIFpdCoO/2CR2GWSPjGyC
bu35oWXR8nr4gtTQ/Ol72CjvoGy1byqTO6ALgcK6Dlj4DE/f5VfT8Y3+PFuDqvSI/qMTjSuMjxt0
pZ1etPCmlpP2qTyXCQJzM4JM6oUDZYC1LIE4Sx66E2pEwLk4FHJvRAY76Bs7Bcya5B9FU2I838k4
uXJPRKj2spP4FU5iASqiRbANcRHrbg+3wYMF5ptOKD9aDuApBLajIWTBpzvGi6SbsigKMvFT9xmP
1ItK6HDJdu2ovQpHmvkLPlYOd/MNoyadpF69eSis6kq1nUKibPG5CzYBNBTTbMQPcwGHOwXxdLpS
v6Dfamvifk4v9NhtS//Bx9/EJdp3+9BuMfDIX7h0/sOtDPN+mKIQPQgHo0bwNaBG5y/xHLmqqobY
Il6+qeSVQGLWh8IZqpKXhudB++4tVFMaB17DF5qphBy6PlZUGfgq7wsUx9p11SBc3mY7Muq16yXn
XbxvJRUOEqFgKslrFdJVQ5w7HIfcxM7yP+ScILitkvX5HA5UH7YocTf4wO9zyfGGaXpcUie0tAGF
96ze80w+tfEIci6gQdMRhMmxxgRc8trydZN6oXICdKa6y2iqvbwg9nRMg6XqlWV+jTgJ22cSYRCV
orfiNgv8PU6/eaLauYp/tkTsHysJad5uwv4caETzYfy0HEyHKfqquG9Zd+ZGWBpxuJahtTnewjC6
q434twfeg5a0uPzUCs7UzZMQ+A4VNtjZ4GK3ImzsojgAYX1S/IzVeVwzTOh/r7eGa1qF8RAWaTs6
7XmoYmNtwyREEs0nUTPqHV4+77r/45lV7aMi8x/5C1KW6D6TZNjjpslrjSEODhNXEsj24cQsnIS0
Df7z4y1b9cCWhMgZRYrEY80Qf/KThzafizViYfpZNHyPK4M9DpogppmWe+rUj1CTAxLhay6tbpX9
d7D1U0Cp25GzCzLZ4My6pXnGOXLA+85eqrXVCJ2JHbV4Cp3skdnGNBfoC2KsbktdVq5J9xCR8nHA
XPVCWiRR1L1GlEROILBvoOSTJosb5Z88QfTltN3ZTMEiuYGG+kq50mq9slBZx55eHJtlL7/MN6rg
LS1KAzn3hXS3IBLOQ6Vm2QaTqE8LZOc8pM6T+zYiIid1N29QVngrbny8EEbVgakHiBBnjLaCJXFt
4oxIs/gQDYmjcbuFaCtEttqduJ6yYoEJKfpmEzA9g+F7/hqy94n98keDlGMn+Khclwfvp0MZG/Tq
B7sND6v/8M1Mp955KfK14kuVN2VlFyPYkAFe+jqrWjduvdmrx4eDdzbLt40VMD8fNxJm8thUBEy5
bqMcn14R7QrIGyubiSOQoSWa9RfzoRkqG2EwmzYEp+o0FJsSJvXYSKEwWsOCRma/kxuapC8WclyP
tVEPAlEO5LYE6rJ3guC3Zcplov+gZu607l+ejB9CzjGfL1XYxrXpzL8udN2uFzUecAaKbq9ceqKm
3O2uELHICeEr2WVF0adp6hUMFA1gtL7SzbIae8rRfgwShyU1+oXVON3jLuiYCSZ+pEC613ACGAWK
I20GQaW/qaUl8lc/WdhCpmyLpmeAMceMHaPtBCLmBnPXEuSnukCF6hFyrkunpZA4YuF3HWQ+pXNf
p6lbbebuQwvVUhszeTiaRx8ABV21W89b+8tW3Avx1mpx4OiyGxf1BdGZUVHu21keUtiMIYZOsG5q
+sBZRaAG4NRyY7JXTrxqypFsUAwtSgvzdN8g9igKP5VUvWO3EucQ+Zxh0zER3j/UVIbp9xTU4cop
70Xg/NwP/0O15QlHtKEL+IQj21FCbQoJepoJB0gCKifd0JI/gIR87J1DIGdgjkqoS3XQ9wxbDGVx
OB0tCOeRGP/OsA9W6XhJ6N+vUJ6nNbMshlNvFR2b1IrTMVZLa7IjB44gLoVt96tmi52E2bIBy7To
EstGvo4nMRwdaqFLMBSZymWsutoorMaJbchJQHH6HLDWzPiBSx1UsHG4C8ePmQ7BgTj+EUYyPmKt
QkV0L+Squ0vuGH+cahk1Tqp2eHq21YUYbbSPe7uH7Wc9wUTF/Zg7Re5VEgluBWyjEAdNTtjtVwiD
9Wh0cD4Lg/Oh+I8hnYPzFnsXuzMiRpJmkO6ypb/cbXLZ9AFcoLpRwtkvlXo1u9EP8jEG9VIhk4El
whYYCcl/qSFrXcn7FDDb/XqQszr/aTR4/vYEXgVXFu+QpiSiZTc9K2DLM1f35StWWU9fFykBNEJJ
/SyWJsEnv4y0BC4WsbrPyrOs1sgXLSFZTH3xSFwHukxTSkw+J+Un7Zb8yI4alVpwWIRyrPqCO0eN
t4OqDaionw8YJtBHB2ezh4MLsQPLihuD6mzTD5C5UrL9XyUZtt9CtqtwlyrY60rO+jGAmHCfGIf6
ZlgyCSOS962BG+UgAWcN1uyNV1GKDg410rnXWE4CD87sfhm+rrDx3hAWnWUiAAW0mafcCV5Vsuuq
UATOIuVkfcVrGRM8BF1jtGEHDKLuJA35d5Cji9OyKbpC8+DspLwyA3C14ZmT8G5/xNTSmWjPDUmG
6ee9H0vTo/RvOc7RVuGUFtBkipjzAzUiYw+B8V5WDszZVp9cVcAFvAp40wRNw6WDLxlEDMRN8woB
WTqQ2tEN3+sQzOM0IqJbbMyJV66VZFwQWBkxz70tTzRfvNqOxJkXpByT0DSy56RBOLpZebNOdqk1
QrNtSfrdIJIfRNKO/FR5SA23ttjGNs378gq9r5N5bexseQM306C6dPxroOULC2+dcxG9VTL0XrGI
7VigpxElnt6KMHgWzTTat8CmT+WUMgVv/BLtNHgbg4Fk/pbBvvaIEeK+aAi/LM6WiY/oL1yC8K6y
25UpaCHNKggpzcOrciLl+EUvIbVAznO0kVMfVw6UqvI98yBIhUI203RZYGQIkFhV7tqMpHBD3obE
MOtoT5CE+96Fhyu8PGXHo1ypYrme0yo21vLSFh1BslI4ENdlPWvVqzWKDsDB09O+9n16JlPz3NKB
vveoMcFA2AbSD4xm1PDy8PYWrB1GevrsiWRJUJ2gatAlfoI2HKvGZOPtouM+qGzu6pPzaU0tnB4x
w/sdpzqjEaKDmOBgxI9epWtm7eu9V2/VgAAVbBqDfPvqIk7Vu9bDfW4xhRS9NoH+xjBGTNZDBJYN
Pc19x9VNr+9LwChHpjH51anJvgVYT4VZ25ogxyj904s/Rw+LKXf84bLFyTXS/OBWPhnQf8wOw+FT
AjGEId4J0/D+WklHBK4OuJyBGA6EEfd/gbeOn3ERjE2YbxD/cq8RvsoBx8fqItZBnXfimTe6335p
Ge/C9eKABwb3lFT4X5NQ6QPl1UQDmfGh6jZi8oIUjiAern4RrVlRSgZw9lbwEPmFwwgm4Q5VZ42s
qUfcfWajyeG4mXEoJi8acrj37U3qvmPZ0t3xcM120aGhAUGB1RvtptoeR2k4qVW7gtvA0VLMctrl
FfzuTt9LJmVJ/gl3nxTRqkwM+kkm0MHXrGPO5OEt3CEVHZOVDnCmohpjYgSuvORzr91MxmxvtoDb
XwS4LzOxLkch9UBTUcIkQGiYqYdjsjIA/DGWgZhQXz9+aDd6fINJBf5VxXjbW5agkM5oEvj1EwSA
20nT3OXUkj7AYN98V1cSwwuvilRymn+8nF8ZJ7uUGRAJFUbFK9/7cx0Op/N1q0dGPyuCkEaBI5Oj
X8PrxB1jeN0Ixwws5PHOt3vwDguM9H78sl8MHkdcJb1OQ4NUh7VO/d35PWaBsSiFar9PdsW6pfTB
jmJLXSBbaszKykdZxJvz6sgFLQ0AZCIohhfjRDsaXn9ylWFIev3tYTmk+JpMp0IoEfNkJGon2TKF
1t/vz7/SX3n4UtvpRTGFas84B/ndAdW5XpV/5HRHZ7Zw5aKFBKtAteIUqAbOmUxIYi8f9epudGf1
COlCJv4yPPg689jRmpuyxPUqhIr++7lc+10r95/SjOQ5cxye/XRzMOCat9XyPcz2oMT5ZKwQAGgj
jCBfvtXK14Gm2kdGeQJ/haiuepxcysAg0m4jDZXzaS53jqoFserStdWwsdALq1E6XZYK6Q3U0zxX
9Gvrs+p2YmDlED3KGM26yI0rF4Rps6L2YrClpO0UOaRSbHA411Ok82piW5mfBEl97OJKwgZlekMj
1khoyIMu9DmCuZn1pRZrVf2EKJHjs9hrH1TdkFESOsz3sgmDV+U5gMbXyHIOsORftwjbKijsf+w4
MsmJe6OaI16OVUniv8f28Z9gIGRqtUB6Ksdn1WMWlRHD7Au8e9FV/4bUEVtC7gaM5KcWqOBUW/ia
2tg+YlR7IHCGkeswP6WyGUD7qGw6pha55rzIecIT7Wx0E1DRqZR5TYTSkImQ0rzohw0dzdtFGWYP
8sX/Ri8KvSHDdDgjv5xBD60TUdryRMePlbxnbBNR7p/jCjQD5cNF136hf6nUpQPmerxthq4Zjtch
s6P5nGsIEgXu5kvZ2fsZFcHKtUfHH4SjZhYP+/qBCWizJZcZIg0YifZ0P6eH/SFwuM9YfH4SYzEp
X3xPyuoH2arcV/9som9SqUU0eN2HMCKhRLs6d0LCFRn0NDeQPtkhBUQ0yu559uiTwmk+bx4o1Fg/
OC0TbasyIGeyEri5kuKkWetzlBFaZCrbR6IDUMYyzRvXE5wZLVgoj6YQ4BlHkE93ZsY3ZIF2z7ke
4Zy+JtMCFmNv57YaiYAz6gSVT229KB1waHIm8IfL8enVmXMlmmKcQMOMOP8bpBOOtd/JIfmewK+3
UaoC371UWA0NSE/KJLf3haUFpdGONsYzP/HWtsrgDlLOMgO5sOjnmyid2VopaCK4NJON7atAeKfE
vShKdizBBCluajHfYf4mfRltm+/tiSmUkaqEVpxAeJIKjWMLCDe2aeIETAK2AXKikPq8224iFU0w
sXUXN2o6XoqEArBaUIVCfSjtUrrXiN/w7lwqX2iuamHtbgWGOjNqVdvg7Y7FArV2UEiwxMRjOUQy
uu5YCURzhmXIdXCXxR5YWtLSqfMT1dIHN6DgGucynNujHUF9FhoWtQQYDiFwQZ3tRsa9uyKlerHf
kpM8xZCU7s414bpK4Y5ry6Oc5ZyQwTmwVt9F5rXdD3f/LbpSmoC3lsd/cjvxueGdeV3ZAS/8UmzA
MIXKMYC3Chb7FLmoocmLrEWg5seGgP56dZ/+pLLocl8WLJswoCQc1iSnxdS+twVBWuyqxYb9tgHM
LuPL4EjbLlp/AilpaXtNscOoYUTmm49Ol4cBgIs2v0oq+P+qLB8pB5AoIviIUbphOQXrP4mBxsqX
bhVAPITb8kyT5DjOSV7OrmaAn0+2Nnlni+Y+wPj0Lri70RBFaESrVtQhnODYnAWQ/cg+O5RI+qTr
s3J06l+34Z9LeBhzzs48C+4jD+xOChp1oLvyGht16KHTIf1BkHs2K6XKBrNG+rXQU1O+vWriTLAW
U3VYtfho0PVL6ykC9R8T2858pwRjOHTMZBMxKIpZq8mFFGJ8umoXqWLHmCHi8YPzFhJRGo2I1vz9
I7a6IiRtlBOl+TtYcG8AQXyXCetAtsbyF3+d5ihrsfPy4cazjOMwFF4UvvAZLFl4dE50J81DH0zQ
/bmYMR+nr0n8RtELjovGxrxsboqJIiL5tnxgFLOuNleno8CuUjSUKFJiMqxMdGtCAaErHAdW9yCA
GPTapRG/AuZa22Q19nToHMZNTkjBYfiwHH0KTEiYeQ1HGD3PbFiOyDRoeu0IF1KGV17AAPmYqsVI
G2Aw7kpkexsQrFOMZmO2GzYycElDrWesU42CBUZWJ//b5LbAUuk23yjBCrGh80Z6DlcTrrEyKX9E
WwaCmyCzfQwyna8aL0oo4x0n+s5t5TYo0JiL2ECh7YccGtWQjW+qbqZjX1non2wBJp+fKEiVysZv
RX9FO5GX7A/Jw+7o+gqmIT5H5ZULUszdf9kSGJPQMHyW8o4VHpjTOXtVcn8piFRvyzHvNN4DIp9K
exSIHdb1jeTgXWPHq1oSdpp1kP4FFOYRysVew2JQd2hi8jmd2LSMt8MkgpTE5OElkBNeLR+DzKti
/RxEiok67JiLQwG9EelF/vT6UUzVct+JO8hZMgpyeP/laK/aL7soL7Ax7qLSfVEfVGsZBoAxJAI/
bz25BurwqNzIwcnxuvzLa4jWAPeG+ovvZBVZeoMUT7sPkvy6DKDNxHlyQdlgUP0WDJrvKST0w5oD
nRti8KqrgkFIslz5RmLBOJ+7vjTklKgFh6sPg1sDd/gBEhyLG/vdWNE9mb+RHoCYzUMohV02Zip8
6lZEsVOFCIqsRni4ociS7qODJPRA+6TrPxf21zWBN8Xc3QTz8hAPBp4XTRsSpUqvOjVh+stPM4dM
Wm71w0940n5ggY3n+vPrPnrQexpkPWWZ8/NMgKQbSPCX8pmXsfA5GhP9ZPPRnaH2pg7raiso8sPD
7rTRov1jv7+WRTgmFP6pMOyeMlyay/G7r0/iYsPy3TTl8F2PacorG7sT9rHDyPGkWNFlUW93gJF0
yZTdWBOx+WaXt/X+lVMMM6NAqLRd9LMGcuKLohD9B6DXl1CZo8KqnPEKx8nnx5YUUKDmOR7dyo7n
Ic6wrQFxqovv+G3Z8hCed+TmITmjJPNVhTdIqXqUOjpuKFLBmiwbwHYxhHStMb5OjFebmsLbcQQW
CFpk8dtE7SflpDnWUHzGHtnV6rqcc4KGFs7M3aJgQ7k6Wf7YHrV6A/EzA16mpAAW7/vUhXhmiEsk
DXQQB4jwtsGx2hlpVI+TVBTyqESqsqnNQajPUOlIPZ7iGRSKk+8OWzf6vb0iT1cyT3j3lnD5+hyT
SKv/IV+Kfxk11ZeXGATMGC6X2gBHOB7c+kEBe7dTsHi0xXyZec6NcUU2rjXZEaM+Gjv7HWg1+i6G
Wmf28+DXVTZmePXRYY6lHKb2lLsCEIEJnM0dQg0mb1K+Uo1Be1ChCVLylMolXBVUBZOrmhpJE23U
oKdhsXw93l8EQ6cIhtKANF7kG335B6VOzRffslviF7BMp66dhxTdFvtLc/VKqG/HZ1mfHRgkgndL
Fu28pkETAlRIrfWjPPVHSXp7CBY2Ge8nNmbPx2ky9Cm+ZP49h4trvwOqUVtM0jHMj8hddOe6SsrT
mc8tYcKJIGqgLoqsNB7cz9NDeMW+1iewiwLwWtvaK6cAR5WXJ3yOnlFmVxiNqHQ6M1/XIDpoukkR
R62c6GukrI2zAhkuaaGRtyP4hwpm/Qj6z15rYYJoI1NDKUKbFeiA7YrqPrqSlziQ5WhOORBpcPtx
cJL5+gjxJFHZ6LZl681HR1YKvN5YE33CwwUvFMOFH+7NUzoNkbEA9sTHnUoOGEteXS/C3F2U7+5o
1uibS1BpJLlKR9tRKGMSCKRwshwRo3j+k8oq8o6UDNPPj1jiHbd7VnJ9Epij4bwD0V6tHa0LANml
tFHjrVCQtxDQ2w3qsCDPKpm4VDU8oqeEfIWUCVvcqK46JJDFMtKb7hsD7LUUBzGQVZ9f1kXB2/nK
rvtR47iI/mcAbNORu/KNFLEeDdkbFtDdUHtE+muFEvTovajR2pNKu2llepdWGureThYDDj6YGWtu
CXsljD5k4zNJangMNc1U9YI3zIjXpbLE8MSjp6f/lmX0vSy2QL5DaJ5t5aeScmOXLJtZRwZJrGr8
yJo414OUFB3XzU6VvMLcTkrefxUo6KwXd3pSYkTAsGRnCIA+CylW8qqwavw6vX+ZbhDErjKD8Iv8
CaTthWbnh+ElVq+uCxu0Ao/7EqUjFjZibiWrt2m8XuPVD7+fwqjYEM7EqkAsqWXXBOuO/zruy4Od
54nZvU+92BCzNBDlTohav1wauPvAlWO4wDbAzAoY0+wiwzxMfEHzwewnL/46tR5QkTXNtnV29WKm
osqjc5jVFBvpyyaRL3nTygS0WnkIkxBGCzBy0Ez7wQuomB4FXsNYmuYA/nbDN5Ampy+PBNKCxmE9
d3QvLz1lkSEG3wkgMxyibG0j8J6+svfRI499GHjAdrk/OkEEddzYqy7gVccHb1wcktCcQI3IYfqs
e6oMb/bx1vcM00YH20hWZL476+7+uzpTPB/NK8i6n58ee6MNpUn5cwbOsgbGtjpO5MvXyOImRsC4
aea1jd70ah+26N405s6gt3mEuEDP2rpJiHDwv/8fsAWoajhnlMSE9sawYNqiObyjKqGLAGeKvUuR
N3oFcD9kKgcwgNC5colv/f45c//OI8U3wcNJYNWIN8/KXo+RPE+3fOhXtOCcQftwh9eBTH1N33ik
wA3zbJqo8kT5Ls3hRV4wb+4n2a+NAoBQoJq3Mpy5Ac7CTvXjUuAPBOSMK41THdbVYQBXJ0jiYDW9
Rit/O/0ksEfkVCfpEMCAZTcY8i/wee6K3N1Vzd+7v+VWGIf/mlAlOz8lHJik+paaI7cqrt7cnYDa
QxfXyBqPBx0aUMZerAxZzOIlaLFyGG55TAKFT7mxl7Lc9NQQDMu8f62/ANU1xgbWliLIU33cW5JD
u0OIxnPBQQ7OBh01CsO2Uosf36hVlAJvrP8tk7kDpU5Kbn5MKkRy9NriJvqny7QFeweZDKFrejhW
FrfBi0VSg19a7y1+MCkQNJuRffInFTdkYpvVnBjDfcFXn4qgUratyajCrSugZn960BoaF/Yxb1uo
AkiGcm6QehdtINzVp+8RMT+qONX5iBV+6JBmbMvO9PfvtDwHZB2nUa8//NhlRLRo5wn+VYSvbk0y
95ApUJHIRvRr1O3oae5bxRLu1zqAKC0tsUL/B2yBgqVsHBMlW4Z5/BiIh4CfV+jeToK/MnxRwROm
tqa08A4ozv+w3G1S3cnFZ0bxp89ymSKzErz+XQ5i2V2fb0SIoFSRDSU1gS9zJmlEwUMiSBAEvwpi
WYeACiGsxnWEdeDM9Hd9sZKX2vjx2HYwDpt6B+JWsGk4+UvZvYVsGhvsuZuZ3CwxkfUn6f/o+mDN
+g5vw4bEDwglnGn32/hxfZ3KubnpCNSrbXCf6kPlVwQnTXwxkaHFLpCjDiNffdISiXEzXpgkH6DW
IWmfUBhTuBLZgXc8eRSLe6twx+4EULj7JeQd/1lQ4afhv7FYx3tYePs/v3UVhR+3Hvc1sj1u4tgZ
lLTmmb0Jtk/4SreUTLAEG+9GVnGVmvwEUq7bohr+f963VD3aZDy0PDvRWSLDAFGshtl2LDBgEzU4
MxdsZHZ4zm/KROVcZAsF1EJg1GMxdtfO7j4BXGdUck66GZweoZe/S7ep8K7CtJmesmKZu9N667ga
HT5hNZ7Yd4quF13NzTsAiUjQbCPFwdP23mo+Dgy4dJ6RC7EwqMQVA6WYrSfS49BzNpBUml2ExZQB
LeSs07pJFfqEOnEAR4OOZ/dtwFX7y412NXnVJyosFExIOzKaCzHiS/7R5lzapeu+ofob95u+1XG4
2569Sz6YhD3hmgUNqOIl5jlc6zD857EeWxP6TC+NR2jeYIqUahuUlH7B0t6G2pH9uGc597Fpw6kS
1skBZaJWogIhREiXKcBBkVrq+FC6ydF9GG+Qw4B7F2q7EKfVcSBCFX0MhUsQcSf2pJW5CSxY9OG3
elpPmRWF8YdTAK0nQ2gZCqrFlUBhqtjxvz3Xv1kHRyblHtpAZYBJrS/cL4zfYqraF4KDYEyD2H62
RN2cIXtPyramebwIJmdO2RQ9w5jtWURRXYu/7TYW/SNqLq2g62e3CGJj8cX9rfBBzOCpuHerl001
LgeRdvXPJPEfzvrPgE822wg4hw0UzpBAvBh97siOoc12v9GPyeHKqlil/IR8COK+I3YLeW2sqJFy
a45ZZfY38Qt7sIA0/j8qxVgmxdDvYsMVTTJChfZj3hGdsq5AXlH4ur3WGvAVEjcpGr4iBtBGb5k5
NYWLEmr7JqaczerAPjpPNpmQLzQ8wYJ4fL8LoBzDqOsy1VD9tTh+wJX/+Vmry9C7wP4DL8deClVy
xx8LaxiyRwckC1FE+RafZLHpZb3RXI4PEXZ2XimGBGLFwQhYXDFe08onWxx0TZ7vC5SyKXs4cWA5
72Pii41AHGq5MZhocnXHV51/Kxx56UnpVeP/DQ06OZ02HZKJz11BQpr8MCIOwbhw0vX6UbQQW5tP
877WmMptxgYwBAmCCEcewb5uUPCg5CPyy59hG+JG2Ywi8JGQWtU9FVAI9g2/c8dFH1pfmduCUtDr
P8LaXMH0+7UYhORqxktX4RdtJ1unjHOUtoOsTqRaPGzxlfV953YrHsFsWZpHPLU8p9Yud2mj33hF
0Snm1Za3mqC30iSG19yJv5x3MZh7wUNh/G5qp3laDGLUZFiDBO+cwsTb3ATIiSkRRJBjrtY8e5SS
8F1+8F0EinrCubYvSWpkqgVQ4AeE9SkarIGjSAA+Ioxv0AHdiQAJeUYj6WitXHlgxiVPIjCnGzds
L0ruMnBFP71x02XcYnbru7bdDqS7ZhFH/ZPRpx3uqD21ZUkWuReXzQD+BfdtbBM/Fel5lwFYGUYa
C6GbW0k+xYyz/ysfKV98hHYTgpYlkWlb/fdeXAFBO4LhL+4TTp02806WnRxp6vHw4TxTclz47diO
h5Pkd2eIdbUKvIAFBCNUT5GktXV53ccRcGLmiPBe6K6X+7YkcbKZhcEIh+RvoLmBv+EktRevXIy1
iANo0HYG+lV1zM3MCVmXu9S/RJ0zImopMNnBDAyH3AKNu5WPygYSseStw7mCLX2xNCzKNS2SXPEr
mL3xPcFX8qhj8BAxmEhVy3TlNchbfsRVgqVj7O2R1UUePKoxlPRWnn59A4OsYxzgwOAnm0JKDOaW
GtrQZz1MnJAuDIUe84d0gW2Ycj/dM2Fd992gq4GPHIZrTErrpNC12f7dNmzeCnmfG3eN7Szw2LRu
rh2h+fcmquGj48y5B+mIODgxoagjDECqMUoEGY6XlzhCJWEd66yaD8SwGF5Fr60r3Z/DwyrIQRW/
Q2folXiMo9WvKZzGmh+m9tRvsXbLI2ajfdBhnEARzrU5jAESq7uFsMwASJCZBM4m21LZfc7bgP8/
d9ug+mDjkIafPE1JaPVnFA+7huzDjjEJguLFlbYZvPvMIaNTjSIZ9WJbQIq6O4uMA5IjKCS4vePk
LzOF0SfLvS1SA7BY05Dfgm/tDTgJkh2DP3liQp9W1GAq8vFPE/4/98A0XW80BWlzTEb2KI+nghHH
YX8fdOMFnSZuhdWUugNexnIQ75u+QSnypg3uAjaln2QtfieraI1Z4qq/F/t/YuwFY9oGX3MPY6s/
XMthw8Om4vtqt0VrryIfwqhYsbhHmutxkSfIp/GgNUSokmqhkbaa+J3Q2ENtmuUGnjLr2gK201jZ
jE9VGRB2HcXHeyXK92XyizNVIIYeTLnK0nklT9K610B2qdh8e1RdYCH+B2yHVcmwEjo5DUIDTKEI
7yQIy2nloCfG7vMdxVNL92ZaLOvgjd3oEdpKFNz6ttRQVqqoN9gk10s6Z0eJ21AlQGTVeP3YyCTX
cdYJ5e3ejDYsDJfxecWEqE9DBtH6lfcQUvctjv1+IwRrUOdT/M38Xv6FzBLUH7j542Ss3Je8KwWm
K6kKenEqhJ7xQ48FKPBTuWRXPkfHh7Gz/oSGZSz6uIkXmRglTaIhHfr5IHUwfNEjuHM73yknvOJd
KRDx0b8KlWkjaDmD+XIlmVLkly3BOv/RxoUVlwiN5ecsWMA0TUpnrNsS8xF3ImXA8dwKiUOPJuL6
DmO7lLWnTEFbi7BpRqjKiBq/wZsuvSK5bKEoucSSzo5qkMFNAAF/axrH17M0oY60avyzSb+LLI9v
Ofmkptd5d0Qa3Ln5UvfK486chV7wbMIrW57U+5YQp2kgpZgtDRwzZZU1igYkbwSk8wW9I/UysJgp
U1+QeHMIbCyTvwX6SRvkp33e1E51T7/vzNs6ZSBn1JxiAok6K33I1l5bbAsOyO67OWt3Tzs9NGr9
OIyCB1VP9OxA/gZwooohka7BWIEtQcx/I4Xo+3vLtJdMdFKhTcCaU3HvYAyqukPighd4SspUpVDu
1NxqBKJo17Kh9fXya+WXuJh/rlhJ2RomMpoVGO9byKYe+ZCpMrPUboP5o9oIZbI0TZiRa/f1Qp1S
gnpiCGkMxXJMb9QY4F4JoDXF7CXw8EUCIPhQyUMcg/kz7ICENr0dsC2ykJtvMnm3TLc1i8Jtw2J+
IaihjWmODAjh2bHpi4OpKTGtmOnQhhaB5jjMsfcveWlkl8pZxuvUa7uZWZ44CLexiMtrTMrFQ9qq
xmbW8KMugebIMpOeMtVGFqTP86PnYo5r98hyRI9TCuaF8I7WLiZ/I7GSdhpziZa6D/GziXu9AK+X
Kfce3GL3dtxsemYa2GYkgVA33YWoAtcFjryCW+CFoJoxb4koTq8yyCJcpTGVmWosIdGZLXey1Jnt
VsyTGlznU56WUYnueftWBw7UyEjQnadEOiTlFk+qpzyfhAABmaIJ7WHB0rKKrSXT8ADkD8ymFVsk
RFMtig/+N6nshrFav0Np1DBr8kPDunyj7ahQuP/xymLEycxMu/bB90CqrjvhIasUgnb7qqEg3m7u
lw0XDFErfDbCiGkQPEuoKnNe3l+vnj59lZ1YlUSVfD9cc4Z5NnjAol08IWvCRf0Kdlqdle1kSbaQ
x11aDV4XEL9bjEAFCZYaQJq2FoExRw/+LVAogQeS80Fp6yn60Gfq+oyV8bW33ciusNKqr2iY3nLM
afUhg+t+Sq5K2L7zdPECe9HsvBTahrbuUbmoGW6oO9WoK3bUiaRl/w3PsKJ9CHvyAKZcHEvEhW3o
QQfe7YSwzFNFLXDrukCacM8aF0N2fAW4ILM8re+GcHwzcxTsYOwc7PYG4DkaUxEOUYuvlydQWGrT
dzmnWqYqkkcY1fTSYZGQgcMEqW47SjF3weH4lMYFYSGFrEtsRupfmuYDczB9oc6Wfu6QoZtMdfwo
rHv/g6RfLbV3IWHarsXu3z2RR1N70kRNMHj30kH/2hp/ocQOHaVZpjlBHpK2Q/Qsb6VC7y4pEhyQ
pA0PGHISJEneNAJEexa0OI7GDnFumS3vxA3MGxRer35AIOGt/d6SuWeFSiLJ08BplmuUl1BbMH8U
8AIfduHjw2O/2gtJWJqp1x8Pk9rdFhT0EGpkA754b4nKdkeNq2PKF0iDQ/vebZpl/Fq1YLVXd5lD
RukyYJxXC4cUffyMGaRFKScAhZ/byaRlujygwUVWcBZ1Lb2qnPljCD9kXb+zWLs2aOroVpz1iWl8
A9osSP568qffmpmA5mDELOXK9opp59JyBlNXYUDuWwwB5Xj96luS4o9dr7J9fM+0m/WMw85WnjJh
T2LpBDvnMjhU4nvf7yGountW9aXItK5r0ymWhEBKEXkqaJ7K1PnMRs9tJWsFDdr2e7XvfYFbXOXg
HbDmUTFctqxPHmfjeQk8Yt8/Gtqzh8GWHhtyb7XgHx+TWH6UUI8kC7ofUFDt/AIEnR6wp11N6Mzl
5rVspcDgAZPA2pVd5sBvYF7RMGcISeI3Xik5juy28Dgv0CnwTWodglWSY3rmjA2tuvHw2nTGh1vN
ZDeMfL4cuekZ2jaMXXee2efB2nVXQseNM0CuIUtRFvwLJt3cmX1xKZSXf4rDbTLuj83+Zzx4gD99
3v0dGmwJjUe5m1Pv4oG05n+Iy+MeoJJ1ztHbkJRccU9YWoifhEnK7GhiTTUi+IC+Crrw4QQiW0WW
OlGV+jh9Pq2DQZHorePMSFxD+2yk9cvWrlmEHAaYKGk34TfCeMj7k4aD/Vc0EcGCK0GMYxyHkEGc
yVxCe7q0MEJeRv8rg3DT9KIANtr2YaQoEqlSaNUWkmx9UMoHS3fvwHS0+KvjabARKfSRXKvggY8i
f3NxmYkEWNVxoQ6+zSd0xDkeRD0gU2c8wx8VR19cIBu+N99g/gzaiNAbMxVz+LzKxp+LCYgnunyM
7Zd/Ttt80hoB7uxPIwDj+Jq23bszh0HVqvAbGYLawNaxTv6233/eqiobjE3yX5D8h5IbjjueGjYi
VpZHdxRb+MXluYuZaOlV5lOBF4qiYv25NK1hI5U5/EnVbKIVS9L05YmzddMF2uKgK0484qvte90Z
hxUvy+8IWeWS6wA2VprzJmINMoSB0XOz3alshoZ/I1O4RvcE6uoRfKwpzEjNvhLIfZ55SOJkR2u9
9djH2HiOv6IqYxmti4VxW/hcv9tnJbH0UuvXoZs0Cb+zYEhWb/ooY1rbyuY3YwoqTTP/uivMoRDn
9+kci1cWNe25HRB8S8rmOT3Qqs6SN0+zQ/D0R3GLKv/xkllV9KvbwmzgYab78W0tzW4J09gipmk7
5XevrlxpPQSvIrp+Kpk5L2FO/q7p3+QjNlT8f4PycZo5AEZlOt5zD3Qs7AIJ4ggmV2thk5I5Vy39
HJMDpPDIZv8MYRWyhDe8/IzoURLm7v3bNW3vNs1LBkUWm7HtauLQyEuDdpGp/pbEsZwXWu1RDZ/i
zE4zOTNAxEUeqtbocyruFOJdAG5TZFCC9RMBk56mUNy5/d/1NUZZyl7HU3ZAt69f6Pufn/Go61/Q
ZQOm6gMXyuFDu/ZaDcaxNBzJ6jDkPOEFiyCpBNnCuW+vGLwlyPOdwN3aPKqyH5S8tB03XKEvcmeN
9BELHwv9CqBbAcCBrvTouEzm/wp0wQRviR5XoTcztmVYXE5/5uHiL1DJA7S2Vb68TsLAZ962Mxla
la0km54S7bsiWu6uGgI8ifP/NdHQ0YvNPQY/H1oxKTxEwK6bnPg/nuNmFvv4z/8XYqjaqPhI1wFS
aMfDuYoOMRCFZ8YKAiMN63bavY+yCPrJ+kQAQpGWZyYL352uwnRtFHlRZv3QFOkja4EtaPxZUxGS
y1OEKtiT/eLPXwIHllSoFwYIg0ZJ6Sd6mlUhq5aHfPGG2oitqw0xt0zxk4yvQGTlKoeLMxXjJrBr
LUFUObG02n3frGl72IVDWOUO3PXBHQGIKJY4wpNkivUovUu6MYoxn2a0E2Z3IuqKAEPH9G+GTmPh
hLOEFYg1dhHBgBcrMGixLWAU2+O2zOBXAGfIgV4PHDxbPRD3lf/AMuBlHIgQUX4mbV6GvUHWKQY2
QIZRbl8xuFy/tgMRT2inOJIFQuKPYJNYvIjoI/Y0OZgrDM91xuxHQRTWqshq6Pd/OUST6Km+N7CO
BvyVV+Pa5Zimk+EFEI7nv8yMeCh4EJcZUoNbnsdY4XRipG1ExNTxXecksNqT9300jvBxfqASB3Ab
PC99wBA5LcVHXh/vXzP6IiJBvOCy7ll0wq207kNQeCO5wEwyEeKRqXUFITmRk1MO8NvS6jUbH5bo
V5WlOe/H2E3K2iB4hfXuuBWmhpQdd59LI/7fFceg0gsVnGNM/GxLooEDQXSdVqOwKdYQnzUGQkuX
BbWI7INk504Rv70y2x95TxUEznhPWNz1WsPSj4cN+u9/xm0DqeDLbWOSyeRmmqT7mdNwaKtV84Fc
gjLMF14cpYbsIN7YRCSElu89QIT3OW9uXJylajK+g4Sjqzf0hjAOM/46Upa9M6OiLVgpPBhS5+GL
T+1IBfeCfYOuGoNh1y259r7mkO001CpJ+LXdi0O+dqK6E/afg4qkItdZ6ZbyagdpbXxrtPhAkniE
acVvl4fa7NtQQnvEzxma/73pAcNvonI2zK/AfuJphhfVtLz2MBl1r3/VyH9vh+zdZ9t1Xgkk2R9W
gojlrNtUZ0lR8Yp+VxM5lAxEVhQNRP7GjrnFDXNK5DDXRqdZ4t8InAJiQ8GLh+ASM0eJsQeSrtFR
mJSCIdQbyq07uYe8eXE083Ha33K3OPU2Re4k5rb/lrO9kIDjRdHM3BSlxm1dDoFbPICQbGRQMkGC
8Fr0ygYhS1wWjB180uF5yvIjcBb9i800YT8JconJRqcC26oK10+blESV617E5dUEne54k+5WnALl
f6/OXohF8VdF0EUAM1/H+QxU4dBaaA2xSI//ZwcoNaB5Y4kull7Vn+Ndg184QqqvqmW6gd8QdAhv
5SrZM73Pxdj0VodV1DORmRLLDQvNHYAhkJj+U+ZDZrnnicIyrSsX+IooRM4bWDDRnJnJkL//ZmAA
fIJuj2wdPrkiNnl3zhdNl8mKHsReQjyArw9X3BlKjwadTlbmNro7xWbLrvCOeDD661PF4MC2lQY4
QN/gmUs6iRz/1eiPs/yl41iPLjPixjxAEMxO/vNPIScv0+MuEa0lBW6SHI9/9ZcQ07bQ53wgYJkX
2cJCkYKdRyn59II1hglkTEaa1mGI5ojZYTXGfFGaaoJo9AkJa2MlnyspGWRRZKUdgYAvCb5HcnQ0
j8dV8w6EVtu/RJddkFRX9EIwlNKky3nnTAiX0DkUKyc2rBEMZ17BZ8cHKVdWEE2k2RwKusgGKDN9
DEFd9gP9zKtzpuaT0QDMPBpsAEi8Xc+hEmUhLOKSo+oe0n47j+pZaHe2yq8uildVRsFQ9IWZXz2r
+gVsM2Bol4LU/sXzhiEKqBCDLieQEkcMAuQthGrSQaONI6VwKwMwtoCxRJObbIQozYTjmd9Q/bOs
Og76DashpwSsqec2T0yE0Og5+avbZk5HYItd3N6E1Bz9RETRjQvsNFuW3bRoIgCFf1oyOUSqxilP
rjUszoryNoLXmjYrmTgdr3rKDpa+N5msUg5GhOwmIkbUySS+7bfgZ6QuXo56vRYGwuK8ecKJckE0
21yH1f315uvF37pbi+Fy4Brfxc3LKge+WYKL7PbWfn4GE7/QxqqnJs1ZMVXdRfrAdRVZ/8rdrbuS
WtuM6RUqhAH7lL36aYxSDz9uBMtyRalUP36uVTfIWJQJcTtlIYGsoU06dIkkrsSeyntrkfAqoLu3
LLW/yj8PDeUHfu6PmRr2elXLp/ThMr8jIvLkIG2P5Jd1ecMIq6ZpUVSS1I9EHzrhEmWDiVbItBeb
SZGMRdTJsul3qpuvTUY0pDmg2cTck4JKQT7Mo2bA+NWW6VckGczBf/9reCkSJ6o4aNcjlRhImOjk
2EoDPGXChlcoa98LJBVyy2keCRMLl3Z9VtB1BFD4B2at1UudJaNWyvRLwKnUS1X4gcGxnRz6MSPQ
HUzsKFg/W/oGuA83jJttcG6PfptsjkkDnQqN02pznMBN+latsN8jZMdcXY87JQtPz0QunhRZShXb
7d76oL2+azULQtIjazJynxwYziWlWKiphjZJWKRE99IhFqTrTwv0lU5DR8NHDh2GkdNmdfx7WgZ1
VuC22F51K+0aR5e4cpSJfdOeiXHlg06BBMpftUx4kHYWEWE42y6EKtDNiC01fehr4Ds3UVuQ21tb
3s4cF7Y1GSUDsysRvTG7KkRGZ+0N+W7BSHBkhBHK7TgA1+GAsYkhrZxn8UuGbgBrKjBjMTzWaqX1
6wtHc4065jq3ipzktIoCr71lgx7k2MJ9W2fEcflkWDW5sHxgc0QXIWubLkEpvcSPohK1/XTD5/Yi
gkAufRvw3ST/op8fqO1GAqvRZAOkFPbFcAZxM9zO307XRVWVOJmx88fXixTBvsu3gGdDaSgSY5t2
yLGzMFzY22I9JgwcgwlyfSviJl9QxBqPURhxLOQDB/f6NWDEdxYUDlqn+vJM8dBdwhuEHlhdugtP
Q0osbRHksTlkgUOaPpbW+T4gxr+zm15oGgma3CngUq1/w1PgxZC1fuWt3NIeZHASVZ7PWKmOfLSF
EG6+wUXdVknINZFFAt5fexg2rQvFHfRfxaC5VUfy4pUyyRtaoquOewduawO5pgXcOcFNkadQXWHw
4S5ytAZJ2Rb00pNVXqccINHgfj1cTTx7885KSuURsJR2DKMtAdJjx53sCKdllH5xymNsB+BzHX7s
lHutbSZNMbv+bcztetWWzYLy9gLXMhu7l6Zan/j2LfKRUZKcsbghfECfqYWf8StttBJb4IQvs0K4
+5SZW7FlL1aHLxtXaDn8vKh4E9UWKJBe2byYiotqTGi46H8EWtkybZIERaVuxdRoWH5hMqaU68jX
ayWudZ4Dh7s9VbDHezMJpsXs8ysKXU72Uu1GwFvjYLhIDyrFfNdFERMviOK6uz2h5gJplpXgakE7
nS9Cn5H5t/AgNW0oghQbv34rJ6XTqgPq6W6N/SEP4sCgZnyiANObHzIh3ViS1sZzAqI+HiqV+4wa
Vkb1UJjOiRaUZ0iv5aUDNCaPWAAg2fXDQ5ZJTF9asQA69Pt9BZr0gLJdQGPsSDsW4gHi/9GXiilx
lR3okpL8peJGUDJkNeNpjl6Bgp97fJ9Ksf4AeNm5fqK3CzUYsKc30ASmtFXCYLBH6BWnKXLYGWaK
+bBKHC6vSRPqbI6cnar/BKbxb4yoWZ3/jPhdv35V/fJ2ifa49ZDZybByl8eblU1lkE/RUCSL5LT8
9IDH333EUnOE41YvC8qPQycuVa/HhKyN282k7y9py8DQhhayCJAKCZABZIerjJG9wZwWKoiC0Jzb
IgfBR9l5VyasOH3kwd9h+4nsbGjLkQ13LWrmZXu2BgUS7rbaHjHwrvaf7wvhL3XViLuVGucQmQc/
/RaSI7OF9tRn0lsFoOJRIMz3eHM55/JVOp7ViJE5NWx6yO4w5cOU0VQBM0LtS7ViBkHHZYOXK3xP
KZKJ7BH9ScIhQCp4bsHjzVQ1Ja2aJScSXxqXSBKblbWm/Ac0OvzmBc1HoEp7jnUQrrcHRr98dSvD
Sdwa/a/z12j1NFKNfqYlxVce62Mxa7v4GkdvuqhihI4wjO7x+6Fme1jFIBxlbsKLcluZRp/KHcYX
IfNTDl0gCc5+HpguRgRUy7aSv30gmUcjAaH1NqkAKRDCViJRwhhGWnkMig3wZ3GRKYnV0v62bj3l
W2mWuE9F10HyaUfOMqa3essTgKkgqafdYB8S3HY2vDGhd3x05FcUSkOhNX7zw8eiJ+Z+2lQhC9ee
Gykn4h0q/VUd6zMIRHxSWQUi9q8CgCiDF1J/DLHF75dUZ4/dRSTqkcL3fEHYW3/5RbW/RwI1g0U+
uNwVz7k2KqwqZKQ1ffl+5gu6pgshZz86vB1BBwziOnm33mSuskM5a3XR8zYInYVGftxp20Oq5N/2
ZhN3wzenwHbhbZDGb4ilyrmWAjmGCRtMByNC/GndXwp3/+f5JFIzRnuIs3z3ypKygCrTw8POSbGk
Sl08RJt7fkkloX3noQ6axmbwJvDKXZCyJonEJFywBXM+Wa7YDQInNiK+QYUlU065uxZtAv0eGe0K
AvkgJrAP+pTBI9MPdbWAxOM+TYUkYQRFl8fZgnK0xjiC0MNqk9YevkK6ygJAaltzjgqH4UNDUpMv
7YSB+7Zg2eCsvi2QraydqZEye97ePzPjzij4WqAyRIqYdLLsF3Hd3cbPDsK3RCPi1vPqlQyRf+qQ
yGFFozauDlqDTJBEc+N/P1zz0ryBgPBNeFXnHdkpcjpJoksgY7vlFeaWGa4dhEUyVf8hP2y0sj9S
Ek+XeCKk1tirBaLJQqvTAO5FWr6LUZ6F/N9UZel2x1ff1MdadEqynPe/Ibpbx5ZefN2Tnx7lnhd4
S6bOREB0smPaT7AbtZVk3Hton4esi2eQOXuejEDdr8U9qACe1zX2TOOM2NSdXV/i9U2sPvrVonz+
lK+wHq3KsbgmJrRP9njA1vKj1cv/ITSrgRwWaSN/TyStFJs+MzWehmweQ0sg4FPDw4EJdgLK/rRl
3JTEWAcp1fY+SgufvjYgGVBCfhTXRAMlSYKvhFdHU/j1DC6NGN7d4btPyUzIQWwqKXOsSqtqMMO9
HhNouoiwdcxjenLY7XqGswuACGzTQoqkUVl8ku5QgLgjzKRBajGARLgqkPuxJDZqZBoqdw1ZIjeg
PetmSTQZMHNiTrdmVx95wmeAcetS6cP1sOxCzQAg6NhLw0iS8tVMG2UQ7Yh3GcrEzZB2KISEEdZa
/mhiF7UbGjs2W/86vH+kwI0FBuJyILBvWuGpVZbjzDOeLBaaaBXzMHEz89iB+o9hwDdGjiboTTv1
OqASS80V6DJlZIdAoCydS4dNHvhpE+wUHu9VZ0AzgZJjIEH3hb1CZ4sJxUiaJP071Y6s82jJ+CjY
Z79UjrzBZE6lsde2PdCHkEdsd+1Y/vLKUxsJZ6+9lyDJpv6w65ZYEOZisDsueJb+acR+ivv2NZYQ
aT10GW7i5tG+lRVGod8SGYW5X/cgIsnbLtLTAgI+NLsY4HuiZubTOyK6vbCNhtGQ3gsERABv5SAm
P1Te/UAl94FM0VtNK0G9Ey1CiHlD25oy1nsZoJ9ju5+vaXRreapoVFvYAZQRQAVuNFIZEpDB93t7
HFK8rz6NNlbNQve6JHwOGRq0YKoP2acgT9UAGBFOpF9jJal1l3JjMWK0wOo91Lkafy0DuAhnnaQX
d8Xipa0EsyP3ZgIUlc7ib1Ww8gebC07dqWEae4CSLORApHd42T15uGQSjsETyVyaB8P5Fa3BGzwZ
mj3vKDnIXMApdlrwfk2NFMmGzLTbBZBLTUAaWe8xQAuiZmgnU8TqmfONnHwbD8eyxF8WjWLf9pcI
2RUWMA9OCawWKwg1FLhfAnzGRMWxOFe+I8WMr/NsxGZ5uOsl767BYEjvalN7NIlVVoPXfO8dNjR9
gCvICoOYCk0cnc+KbCme5BO8ECTf/NdY2MYKW+jib3XmIKw1oIUz0TdU7luFJCeRZq8A7Jol1GTi
G2s76Ujo58OMDLGhVmGcqbXXgOU6ppB/uUfLg3ebL+L2TZchOwckCtj2HMvly6jkM5bDtQS3U1X7
M32jGCpFksy4b9hiWNB+xudl7IpGwZ7/gupbfFckvVq1GHuG5fOUj9Z3ZaABqSk3i5KRfuq514Qv
H/cLQAC5wUQzQds4IuREnkYz89rEV7JEAE6rLoAwQoLzEY57QtuELRFCvbVsw2MFzHeK4wW8XxmK
390h3W02xX+wTWNe9nKgag0rO518QgaA4IgQUYoJuTEN2XzNHbtCV7nCUCUqVohhaiv0yxaDGFyb
ZA40wfDXRvyTNiDMgcgkGlk6srExBvfeIu5FFqwYmx2Qbu2ow+nPbl9l3ZHHi+NpgIeRU4pUKC/Q
VjsMaY9I2lmVU+q0mpwlpD/gwBHRJuFLLwptlereB6ky1bgyS7tSVTa7PY3lpuEek3sbpQwqm13p
XWXXsMysx9niihpBLS7XcLCgzU2nV7udfZchamqjghpiTKvNgyx/d9EOCkoJbGPR0shGymvvYzxd
a+/PIviQTKwz5atOVFnOdt6hBqzl9jVuUFL3GqYgApQHvYy9/56AmfDe4z8fqmH+mzWNaC7hZEg7
VOPDmFzuYBxK7bSZc++P3KafjOH85EmU0bH/I0Lkj4YNHpWww6j8vQNJyoRUVlwQxTGQHq18wqx+
48L/uMAzwAWRLO5Hh+XWuHGeIOnDuRE00+94gAraF4PxeeAF3NfKHtav+hJstOuaOdy41A99mxSR
oTkRHX+ObMDnyZNCNKIr9CD7453rR641wowOmd+xjQnQkFBjy9TD8i1tfny2Hxi8KZonxLWDPiWl
Levy6y0bq+WF++MXJ0M4W6xLAi/0FU0TXiH/qxA3sMC2cRHmzkn12Xow8QI1F3I5nWPayFSAgHu7
cp+jofgGbJLmBDhe3WCVBlIofdvt/FIFHK4SoRXsKdx80sgM1RfihXtyYUxg0dUFsIgdv+Qqgvdo
HKsSXg/wTyw1H7PD3ZroAONIE8J6XRinjTXsKae/oxCFk4CIHjw/WIkj1Ade+pn/+/yffwu0Zsr3
eHyvP3OfMbiEOh5OCXWtqLKL26VzsgBEUQEAfRgH9XdJUbSIWhZQpSx0mSmhLUWlsX8T16qlVJKG
nEUik1oru6CNMofU3dJvnuDvgDCasRKaiwIserqdDgQdu9tegklD77+Y7+WSvfC7VTgVM26bd4n8
1y8rIwHcJSbRAPnAGtEbtlq8WqgShfIVsGkDPKPeyAedqMmKdw3RS13Qh8FWXdNPYe/6S2TeHLC4
kBuAK1YQztIrEGf6LZNPWO3V2horYlPNWAnamMzOmPhOD7TquxXaCdBJig54l9wt3rYkHSq0sU0c
4gCKM74ebI41AeOvL95R1rUmHDbtTAns3hUYIn6IGyeXHbUFJGRHFTGbTfyZLtAjQxXlXe0x7iB3
Mgvj6PYfj2OkcXOID9rZt2ovD225vdU4EIby2KzwkxO1WbEweFkHdmcgA3uJWmsl2uuwVt0D3rgP
4e74P0MgzV3tWMivDjL8gDetP48+AlpmQAK5EbUnms2FXCw13YhBbHvTKRArf6LsceixyR0q9Gwa
k5WUISCqqxermdQvezkWFysucudtWBPMSdHWB4WUpE+zL9KSXll/+wn8sbSNVt7y5W/WbHZAK6S1
H345sAKzM3Ao+5JIfBS+pDAuAgBwYJl9ce4UaIhuSFdAX4wev8WD8i7DWpiw96rwU9Jy573M+IfR
x17TJNOrYa4NiaFi3lI1teLy2ItfUM1AvblTCRO1WF3lMuplf0inUQAXqTpY2PMZ6HJs+RCPCjIE
Vo1juT54kqdETuyg1YOERrwpXWX6/890FI/LJ8CifuO7Hm6iLFOJwyXnikGrA+N5/fVKD0VrU9eb
TIRMr5l8OVe0RmGDKFW+Nm6wA5lhrTddhvPvRlxF61qr6favxjikUoiyGGfPywNWjHxFzTejj/Ba
FDl1eC7VBhgESEfFx0WFTEc9HwbCOyVA7EQZMXn7ML/fM3xLCdfcyF7k4mmb4u3ZcGp5DMIIWsQA
cU9dH4HYAx0EAp0UvQHdCqQlEogaY3TC17/x5ggVe6LBy6LT93dAReLAyh3p1ZIBCtlLpByZYoaw
CUPTabz2TRH+GGSJjFJul6NRyn9/6EoLrV3JBmiGJdLwRDz1BLalHLHK1m/Nu9mtX710G4lXnqhW
ejH2YyWJKR+nH5rL/S0JOHPI5e5pC0tK5CogCy2UXqlnPem23CqiHztQb670y+vwbO59KKXLhj+U
jmwW/elk4VAV1bw0VpO9svMczAXqzlowuM4bMLzPARlMGYHews/GKttuB9x+ZQ/HtcSY6V13ckO0
oKkZNdE5+Ij8ltVaci00g0WQkdttFdSxzVk+GSnKDQV9qKEXp1I1Di89yFwd7WYFAVWr1rEFXM4a
bU6MIl11JOAEJW/MJp2rMgSzfV3bhtL3YLgVlQiwKDihsaw+i1DRO1RA2sP83NLBk/fDnfNkppzs
c71T1cuTe+ydaadYJ+E8bD6BIEfFQasgvna6LgW9+lFLjcVh24xf0bF7VZRlOT/pR74QSgrXV46C
liAeOEV6oRqhVVVhvJCCEXSmfKY4vkdM8csWI1Jj6R10oT281Iw/ztO97XbZlxAmUb8GYbzmXmmV
7W07TKc94clygIHURGtTmd3Y1/Vgt+FiuFdgIcjGLeKyyBFNllyifgWZQ6XNgqiNxN7i9chxNVRg
N/8mSlhViynHUph5UV2TGIEptvdL4AdJgjD2fpqy0rJ7HxbUq7naWxfZ4PgB8pAriX3nNhZ4CWSM
GwTWbN5idxDCnKXlXG2KTXH/IxR9tpuxwKLw1akIztcjQJL2eLTd/mmhn8gT4jaz6BPQRCgcw3dC
+UXJ09BNen5XusGdF8f6ACGR4DrTPtzc0wJciIUy+TcnLSooWzyxWGbti3rVdjtNoWX/XUl4nsCC
DpisX1KOQo9yq5J919fYorqJgjqjO8REcy2eVPG6GXRsoVfrXT03kiQdA2O30Wv24WhaUAxJh4P6
C4yBQUrJC5AlS8DwI9mDnC+lEqDnvSbQbhr3wmZ5GqSsu2PHCgyB/ZVH2gS1Plo3A+qYh9h96d5Q
xpwjz2Ze0Vwg2goTCiSsuV3bcG9D1SJLknrtvzQLs87Fyo34S47CI1CWlKSvaeYwwvkYm44KFncL
NkWizeWGC4yDc57EDYxOxc1WXOpDM9++wFoUAWUZ4UM5AQR7P6lj4C43feGJ2m8hT5OF9g3E+Snt
GgbEMT/W5K5OgWBNUwkeyzhRG7qNdXVofJqoe2Eku0sW48YFnarIjlXUgbtBvlHEJLriwp9yviGu
KLfOOGOifpSRnpHM49N9YbmXyT837iJyuVGFCwGGz8l3ZSNh6bnWdmchpKnmlNo74TQlxVHdanz2
Kn1qjoFhJ0X36jm2q+bQ9ldGQM8r29LvUMekjVl8sc5ONdIAf2fwbsi52Y6oHisBSCLp55r12Fo0
WULjKWV9rdjzywcoX3jtLrCSP2DAxHkuqnT3+mmPTEXxGzCko8aUPGM9q7pX8kW0CG+O1JNAI3SV
dMX184IgxEWRN14mtz+cN5VzNvfWfe8J0W3aOK9r1gBp5A+9BX2Me28p2H8zmpbm+rBcbsWTQhUG
D7EdoHlwsuH5/M1iVpKDvWgcToygcA+tUFQWN1WbysHNPvXq8FGC35arztKaHeq83b+sQs5DHsPp
aryDd6wanYXE/v+vF3EWSB6d/lph8A6axQsrR4YotGp14pQF1h5KdjYmN4sjH71fZB/pFmD4rIkC
16tDcn5ZCPRv7Fv+Ou1oe084RsA1rdf8PkRLtNL26nZM/3IMqOlm1WX52uUBC7e/Yc7h4vFb91jy
iN7o2hvVxjUqMwX3NXTMAvbhMQcPute2vMBQo7p2AscOoKs89IXc2wMC4ex0KeIBVwJI3cwDBVlu
GfgvGSCNaH/8NFhqcBRSiwwBkxRtHHumi8wk146BGEdE0I/XNKDTz4hqTVo3n31rxsFyWQ9K7FzU
KNUSV1xW7RLRKkxS8WAhUYKw8AbLh196n5C2lHEnX9j2YUuQCxHO0o1ygew8b+b9yz4LxhkIN3FN
r8rfc+D1JngKDHQIO41SQ+W1wHHB0VUWmcS+qmbM3Lm++PMeK581Ur/RIC4eF9YakuCWG6T6NcFy
ZhX4QTH1Dwuv+gX5TeEod4v+y1AwoH7+bGIuUAntE3zThH0XvCXVCPfqP/PEF0aUxjbzz4ex7CUL
YlL9qN55yxCICo8Y/JVJuDiAfTh+6iDlbeSku4TqNTudM1ZakkJKHekej3wb76v9w5UaQZ5QolVT
iWsD1BaB7B1teKa0nw6UI2eWqKJhau0yuAS7nWruhY8Ozddp5QSUFQLP7g5vZJfwgnq7VR5q6MKY
ZWo6l3HyUNXVWCmMZ+6bauUvCEZ1ZYXccJ/6cKJ8RY4qsA9Z3sP5aoXpYWdscaCFsytlss2TVCu/
uv9KnrgjEAkDRvO1c2+leLIcQA5UM06Wau6YzpA61joBkMHXOFUhIO485SLl76SvOn+u5A32WW4K
Pnw6ijHVKHvzfdvXkGX/lyfiDFQdB/LA3rENHnlSDjT0KsGLx8G1KnL6u3PQBqrqTYu1ac0Z07uq
XERAfm9xyITTJo7NqgoIcAWeHl2EDoK4360Q8jNG23Hj5u+I65XDc/IYzNADoLNPgTkoV490A5Vf
j7HAHV5NOqmG7aP+Yy40ExkPoweYJho47TPaRyXDoaQBXLFDR7fTTJsjt99P+uyDKx9OwQDQwzni
QXyus7uYRN7Rx/SmmkzDT3pP+uSSyVSxtrHE64jIyZUX/R6aajHzPwuljrqqyQpjL3XpAPxedN1A
lz6fJEkkFxShTu7Il3xCPbMsGKh2DFP+1mzolWesV6bVyfgxV7+2XuX3PpOBO9we1g2zhaft0Za7
YKbcWOIOqpBL52nPFMSDzM5aLwhpq4YPvp3ROmkECXMTO9/LXA/salbJ63Q+863fK+sH765qwhL0
0K5ue6P7MBL5aVsNxl4f4zrx1nthostkmh+SIp1ZxLF/pW8/qntwR49iMBi3nXByPPO9lrHdysi2
kGTzZ34j1PSvOS6Frd0HE/pX0HNCLxif4VVYCklJy443NjY/sPm9ymXJMTts+g4udu80AWiTpX4s
TGvCDVEXUDdwo5+5tdO0ldxL5a7pwKRMTgF8ryZk4oMTJqsUgAmGqU+Z/JdbYg0L1AP9WO5ufzyB
2sNHVGTx+0Ijkulg05u8qZ64DEzZ58OWySexf2nsH/LZuNOzu89NuFQzwjdR0uFKQiKGqXdb23XG
eokTjsIuM5jvAA6SwG0/8vcXJc8YKCLGrBE2A//9uwaAN0Zx5qZ+0TYXydVKuVJo+U/j2nZw37CA
bB9+Mpz9zf82fcNMaGbuFL74k6l18tCMON060Ch6+Ykfn2zl74otrkFOcGH2lN9EWJ8d9E73yfHF
Ot7vroClmCMGl+T8wH9KKc51GO5gP2iiUYYBDjmscMQMgcxiNI4v0EvOMbnGt0M5iwKgU7RnBSfG
K7XQOpWt+HuPuekMKXtf3AQS2Nr8LhCsSw5z5fgnioKEZJ+3MBZFCx2iQdS7gTkIIN1OgvjM/lT0
34JHUxr5ZlGehT6Y3VQOHfIIA+zID4VDERmFkNOTynnn6XQOsoyJqItpcG//CvLgsWBZIRsP+7N/
aWXz6Q9d1jEZrUIrK6UmRdYJEp/6BxXxn7TO+qhiw/dyQ2HGcTiURsSYn4AjaGuxXwoFE5aQ75Pl
EIs9QdcCKmQHgWzH5VZXVPT+/wQAFdyBGKWfXMM/ypns9X0B9kHdKR9KQBFg78Hx3lV/DGTR66ad
FevtfT3/4R1gdtHEXQUp2VYwxCMYEfLgCDubslwj/7/dVaxV2P43lCQFqEQTALjCXvVFomiB6bW1
ECj6Z42om6AgE/bJcNhFXhTJAD2e3eArxP+Y79vcspApLuuM7q2y4aPOlmNWYnATFAcaGgdyEvES
kA+qBMoKuHwMiZzyVsjbGxyAPvtOGBRiwLlgznJ/GjFf08vZjPvZDrPy/IiRU/Q9XreIkgcZ9Y6u
LlDUKyEPWX22O35rLKmPczxhz+7IPk73DwrAf/m3NG5pt4rpamtx7Jm7BeygCs41ehuKoym3FGO8
XPTylLofNjjds4sGtLraBH9cR0pcC4BKJfotUqbeywoKNb3skTANlFqtN0nlKbe44DBCw/ONXBqy
gK641T4oLqLFLWUo+eZpF6lu1yVSr5mXthsRI2E6bpvl9S/yPSSjGOf+eDbcVPCw6fi7/SLEpxdM
/5b5nDGuv/YmuM5sJwqJ6jNX6L0jgMS1U6gCq7FNzwpJTMwaVgepcQMXJcSSIZ5FQVaMk1CTk5in
g7IosAyEYzcIp5g4jFN+OydaRNpVZR1HRt9nFgj65wv9g19fZ0x3CEXhmxIH8NMgjZc6VxQlABT1
EedlF9JdIcyLQk9NSnHJu3V0CFGaKf7yTEsJ4MEU+vZcZhaplHI7+6NrKNyFJADkdWbVKf3ar6jB
imOuXlLLTnydanctgfvkJpzOXqymq8zBbXBXZ958LUrYLBizyO//V/oembaUiM3Rqgd54kISv7xc
+Qu/nqrWqy1oVORrLaRUWDMHmK1ZrO7qHDYz1CJkp83QO3POMDa3dL7GQFoFb30kQRdpgCq95Rsn
+YEkqeiAvTV8OoN+yn0cO7RK6hOYlubhlW1l01Gp4aVxG7GgciNBStSqS3lTpnCWiMWj0jPBoAE7
ZlOgm4Bjve21zYN30ZF4raLGaB/GRWDCZQ60rUJZ3Cawp7oR5FXeXBOY35rRVSc9NeH7jJMXZ2OD
5xtC1iiZ2haxWGAoUgX9RVLWpSQCnMNxEW/oBRHQ0rHbgb+vVcCPfWILdWVkhhq+faWBrhOP0JNp
w9ZHewOzy2qZBYUhQ29mT6HtSQ4gaqiQeDpi1o+XW6rITXrAI0kM0ihcPpJf6nHjWNuWkPOJ/Pf3
CK6zNLmH4k3cEPDnB3PrS7Yd3HchhlNs9p7M0N0bqa6CGTqDBI5VstMLhGF+KSe5q6121lDHVXk9
69fwmSxS7Ng+mkCAFLKdNKZuKZAECCZktarjrU9Dwg4YvjOLgI6GxlTB/ALmQwVfNkDXP51uKOyF
zH8vxVdYeVRW5cYMMc3+0z90Wh9uiXK+7mhkmjvqyF7saYac+zE+gsGLY8oUWexohj6KZW+qLPaI
79SmNjN9wfQDOdmEUVnFCYzZEr9vM7IQ5BsUu7GT/APoCJQRcN0iVWjnrkxDMM6iTLUDXqooAYYb
MMhgPjQsR2/6c6szaH+v1BovfSJoiiiLqOIQB0MaQfE+AhF+yoTy34NDRU/fh0qsfzFMVFD+ZMjs
GYI+U2FN6dJuxY+l8W8TDbCgBpEK2iPeEC+icpNVX3CHfKOMfL/0sb7ZtbsTy2nyN6L3Usbnk/K/
L3XLM4dszYonsPJWtxpn/L39yazy5WumUZYAi5ub54WIbq0is0yVI7fsNqzV5cXCdD6WuJq4yAbJ
OcvEEB2qjEuRRbPyQp4pyfgMVEHPySSZ+y1k2b1QyaM1G7epVuHbl0gcqlNpYajOBMCE5tfUTb7g
CYLpS0E82PkG4siKEdcBkhVG1w211q6/nqhn9YleJGNn4RdetJu+Kd+E0PQaUT430IICgyFp47bo
hiy3qnBSACTGpenejfCLYIeObQHrc9lJnT5AQqCB1S1qeQE/ArAYy+98Xjp3WZQSh+sKNJrPK4+A
kqgtvFhy5aBlHw4ejL/+wYMu+8WwU1KrQGE7xKWhlTMFIuqL5DbdRaQLPxMSneh0a33L8dfwK+1q
RdrxxHLT8RH5NzBmCCBth1+hmH2qY6LWxwaiINeyHLN7+N6A4rJ97SYZTwoHiMLeAh24qJ0DbGHY
HE+43InTAf8ZwOGQBbblGOCg4rvFlNesd/1SBKQVf6BAcvcfCtmBGx0qiPp+NeoojItYqY1fl5IH
W4+k2AlNX5a86W8yZko6qkbZ9ntBEgoOC+enqXnPaiflMSZavBkEsh7Lu0HccNaSYo5Ri21Nd4rM
Tjf+Oy9Ksb+IwZJjMhnEWGL+d/bnq+ELdfIAbqt23wF+tUZy9BsPh3992vNg1h06e/PKbDa+X/qR
CNC0qzMjQ/Xi96BU+JhZ7BZz24JnA1GHzSya8flSTAp80Pbc/L8ppgckMQIIMN3werx0ou/d2XZ8
RKbEG0jAPbGb5Jd2z13mF3S53WSsUAxC4IV/ARzd+ozHqaJhA8Rm4NV2xJ1P891foV9SkdoIqs1a
kFcSUIG17fimMpa5QYx0FtyFdcPI7KCqY056K47AfINj/1RJvKXWXqyzo3OTW9XdQa4wgp3ytara
dPEfz2yV7p1IiN0XkRSquv1TbpimmY/qk4y7e85pfHbExGTlt6VOpTT75AqZrr3hl5xbI8qLfAlw
K4NqQkxNqUmqkq5ytW5sw0MA08EY4+CbCivcG8UKTRqZSLsT4yrP9Li0s+CaK3Ku1sudxByL51C0
f5dbceiuOCQjAkXyWzvh266Ns5hHNMlmwvomfmPwf+wQBJtUlgOqL9UU06jG44/bGAdoR3tr4/Kl
ohPfNLWoMIbGI/kDUDuJNx7pBbrSLl+tiQcHVrFR7hONDXmOcJ5EB+A7Bu5S7uuHdaJPfpFWQKMF
SHtBxoJ22+HMKdMdH0PPVYZR9IZenEoJ0wwUgZh8K1JLZc2g7NXdBThHesVZU1wdBZqHoh4TB6iv
As0sVq709KsBaoGe7PCL/MH+i00Ije00qIau3uLRjOnBKjgfFGgOr+/1DLfFmhb7U5/ue7By8Aks
6ts3ykwXMblPlOWzwOSBAny3huzlre7YnexcmC+I4RQ99Abkvf62Zjl1GfzGyU5bsdgIIAm2HAfD
/VO1rjn3b0hei5CMI8oGNdFhNWly2z4ePomkmg8c9mfHTjeQxwjl+9k7VsFsgv8V0si2HWM2xWHc
3b4DszKQ1rJkX/VhKOlJRCZrB1XCN9vRhfuNrBQTxdxo4RS2o4K/7SZS0mA3QdIEEDWEOuObBbtJ
kFIPQn86q7cinhFXXZGJ5Evc6yNJTDYOf8pS+NJjS2SsHqfuluJRMWn8o7Ai8ZWxYBN4EIbpz1IV
GzIkEDW/10qPT9eBwnW+YU+nltcov/LLuwelKsog1J5wElqrf1C2qJAkvntk9LjsfsU4956wHI2C
TGNGYYG0GCUUhJE6WQUVxCR8XNhen5OxzVNc49cqWSOlmahf0uhtFXKjDYTrI8++5e/zGVAVW7jE
nQ2a+rw6xuT58+Tu4neSBKTFVQqNvmAtaZthklpYwYEoFDfXeGkYj8azIxQt906N4R4pbT7/rC8r
5MBgyQSRaQ7OIhnW1ygJa1ZYjZAPCe3qX7/wx+ZU9IueejvO8NQI1Z83jl+0p7TwRaHWWCK1WW5A
sZrMEdJOGmu7KxI7Yy26u0H3F4U/S3cnsuQLH3/paX4yD5Bu219JCLoB7Nu11K5RYiqTsAfiAmPm
SU8WoN9k+lIW861WOJOh0CJa/nVqKOpZe63iL3YNLct+ucjw5s1Jpr2asH5A6nucLLYEEkj7UzjJ
RJNk9Jp6MWLoOH0jSMZFUAn0v1HOsolt5PQJOq8v/tno0jjlqs39bdYyPgRbNtnED2k152Ji1hPi
60woTns3WunTPVGw3T1u3b0oDmRHBmFFkbZ7BGAijCSbKC6eGHx95mKdmeoXKQZNpwfclhd43L6r
0AI4jgbjK5om2x0sUL+gLxOoKYriEF2mBgpI3qHnsWHljR5Sv6ul/NoHugKQONmA6tCltQv3HG1M
l7X9uB2V0r/4TBVJ/FcnplAOiBIeRhgtuUQ7xffvk2HgCp9uV1OZVi99bFC3PuRM6mzMoPkCNmuR
Lb6G07zK03UP50szt1oYcc4ag6L/bZeT8RpvT6L43GnPqMzQjYGOrjVgM/CU4fhw8p0id6FDordv
vUd5jARzscvbT7EC5UnJzkKTqXXFEjnwJIBKIHSXPg3IRPS8yXGbieX9N80NlQzPrp19Ycd5Eg2C
wmkphfBdVUYl/2TwX2xWZ81JYb5IT0bab665m/bceGyRRfGIZ8U3QK+aZ3Sa5ansOwKlePnOCZEZ
+ZiOJlPgxU9rt1FywxEYo+QYPjMygcwIOLfkte6h0e0mT/CD9U8o9O6gxIWFioh0tQdJI6Wr6VYw
88VTbfTHVaa0eIkf4qcy8jfCF6d2ApdFhhjkAl8iWwJuxDPcWFR3usWww8wpTlliEdeK2liEkGZv
x7j5+YDwbDujZW37HzfFzbiPmZq2e59vNUDjvdDZbqvf5ecjhlbv6kGF0are8pm9Hwhdna+sZgFT
0xvRNwUFh6xRArb1AC89pN6kxyEJ8mi2Pky3/JNj00tmiCAlXf0rs62o0uIH3TaogzzxKSUU4JZS
aIDrP2X1EUHqXfidv5m0n5CdZ8mmyXzTO95A0t2HjF9zvNlz5uQIperI084TS6XJnTCiEKV5Mt2K
IfahNsNxLQw1JH5Kko3RU+JVoFldqgmkg0LpnaWPfR6ZO044UYHljylMQeg0WaRKCM7s4SuqH91e
GPmN1JeydI7M07KLa3kjxUsRZ1yok9TiRw3bvF/ddlHhvF5v9L8qc01e+VkmRvCWfiRMav+j12Ou
Jqr+qMyp8FaJlSFvYN2/s3MknCUjvbqOgKRvw0hvRJ5IRm0I2CZ04d1gZIpp063r5Wfl1YDk/kmZ
sgHXGZpWUjkt7ITDczBpwCI0gUgHRZGTZecyx5U4QVULyj+tetNDjc+7uqzocYxCM6YqY50o7jJJ
otFLC0uvJU515O4n68T/HGr+dnVW7DvWcB7v8fyfV22c/QTnCx/ioLd3bDyRvbsgXX9gt3Cb3AFj
s2fHN3036U8Z+ABCguFwyOXhEJpFYsKcAWvungqyJxlNMtRx2O784UQ7GCgFbJV1TmJwnueKMoOK
OVSCgX04Aj75fDjnYUtk2Gf81DIgX9kKZAN2fUm2lOfPtj/SycN6kbbHKhwFYkqeL9q6w0gw4hTr
4nk1gX3Hq8nXeZrazuVPpX4JRWG/6NB/BWwsZ34J4FkRo6q062Hejcz/z/mXCPRCaFDF61qBXAWf
FJgF/azsB1hU7ioWudjwX0Vg9ksYGzFn+FIAzb+iijcJj6FYMDr7UAJXrxaWv/YmUezLj6PZpZwz
fZII0RLaGVPHeqvHdaBZv6Mcru9Ft2MAO64yf2eFTucOVN7zpsQtMQWzky05Kkzvu8zPrrP6p4Fw
vHTafIrEnBtF8Q+cY3G73RmnXSc1Utinz5cJmttBRTyRwXFuSgXvJ5g8SQNQ44JnuKAt2LWNeaKg
1MRbfIO+BpEvWQIbc013mP8fGL9wr2H3U7SCwCBJKwNq0lpq0xeop+1k1dx3ns1M0X2enV/77iR0
br+ii/2XC3cvnKaQaVU4kSam/2VxCwWv1qCGyZvo2w6SXWPtmZTQULmLeqXpA1VT5y+cs0QWiOzA
M2boCqKFy3YxezZtNOIJYWeG1rs0oecdDXN5LdR0BL1FpJWQQnF7Xlnwpx2FJLEloznAaXMezrN/
kxQWOHjFnBMUvODj9x9tsfrPKc5hKcCOv2tK7Qe4uphJ1zpKRRpOhSv67hpLSsAfy/EIUrdsNC+8
GS+0U+5m+j7MqQze9YUT5LjMKY2tEC47tI7QAfYCK6AylCmyCdq9cFFiFICdCBe7Zc0MMbnRxOEu
aL8HFMKzqHucuiNbIuqTHzIXR560AE69HLdasbkdtm+9iDMo9/QRR5o0F0G2dX5zviLoKhBO28ou
xZz3+xrZXVEx5cizWz7p5RuYqkKp1mkxe84HnqjwRdOSqwaaFBrd3xFIft2fgbjdOWLW6elKJGBC
hLHU3QebliK7bhfizzZTIkmUj9essjlGabTzEXBRdfK7xAF2WrZMgDE8888ctEF5ZI0P/+C6knoE
ruPMhH5+ELKNqFyVLy9/R+xbpnXuhGx0U9wLjdFIYXI1Sa5vdqQ8qknLzLxt5P527N5YWjqYzAQd
rNJ5XlcnqteqqkNk1rNrlcfT27c4RBm3XwzWqffj0PyJX37pR8OGVPB6geeo+D7mBEqSdl/C61SH
U6UvVxnR5bFA5FaiiAy46bHJg68Y8A3m4MzQcbNOA/YqJHrbu9TbWFKgPrnOSQfGJwnAbfEzIEpc
zT7oymlRNmLveb0o6EUAtihvWrffVG8bbEVQ+gtS0wwCshXTWFN1pfic3hQQ8W+1q2WFPbieAAYn
Upc0XZNgyC17Azybg+Dr58f/dsbfGoH3ER3FDgGa/bci+fahd3iLNVm6kwg6kx8wYXS1Q1hLTTsF
J8T7zJO13YaG3jhp8WAwsWUfw+PmiKCb9QfmasyWFI8ghZiBCXCkvPcGAbCWxRZRRFYvhzzLpoOD
VflJ+fctDkE9ffwKhL3yLoA4oybJSrXnbtGspKuhw49nyepEQNDnuNxlMEzrPY6XQDkAfBXIs8KJ
Wu1/Ph9cX+VsWE6uCx5ScLuOnm3fzsn452cq5tXxABrZBezQr7tIWKFfgH8v3P6pKGOtyVlOfDOj
3jFocjnv52sprWPGvz1zTsLrZxAR4eQlopBTVO9IIV0G2Kp9R7Xh4VzDn0/0A+woHaMFY8S6+FAl
BSoDpgIOfLxtP8+59mvvISG5LXHv8xqkplDK7PMXPSSFeIHOVBVvRZtIYxDkuR0R59ZInVKveQCp
tJd549mHS2PovQOuSouKXFBzmv7WEMVPt6AFbzc4UDOFeOcWLm5TjfrjouNQRYnNrQPvzYcHmGXQ
eo2/FXN14Cxiujhlx6FEArK6ANmNP845DkZy8P1L0xyUDwn33gj4z5m8AXRKT0d4dvtspxnstnlr
kiUE+BJFPQiL3quI0yZ+l4rlXWXHKsmTbi+Bi6V8tlLVMBCydKjyyuRvF8U13AVpN+CcjLviemk9
mKTcL4w2L0CF9IRhPCI+w6gcNmaO7bSKlU/5TsH/LcUfDmJfBTzMzaUIhqUhI4k+0bmxwRFuiKDL
6oM4Hg8b3UxC/LV32n2f/TRrP6mHWerEyL2YwXLWAIuhRvZ3fGNi/XNnxUpQA3dCLu0cUD2/qSkX
hASbetqXi+rgShGtqQYKDE2SVse4fVhxnqrOnCmAZhZFc7SiF3c5s0sCu6hQrBQlZ8XZle0phT6X
QrPl5tzRWdkcFAdDP00kpRQleJqO0puGqcXYA7EaELT0dHl60OBpDsDvr/OXKiOW+5BiVZwG/WkJ
bjxw+D0Sfihie+tp7WKUfYFWEtjGEp2+4TFw034KIb8BWqKhD6Yjj1T0gy4+OZlZy0vg5i4Yswji
hEWbC5FxH3I1r3xNFa3M40pxtOvDnA9iC0ip5R3Vcc36um6c5x/Zn3BC+0hTgX81wiYty0jhkC0p
mQwLjSmYvb21E1zrLvUK3bwxZNZFb1bTJb0KXiNVNTyMQpQP4aLF9ct9BZfSRv0dKiK8em+VJ73m
WjR7uF+h7Vtv9NQ6slk/RU/mmGmaYOG6140g73UdHfLIGKRGdVYfzVMv7P9VuE2Z+wD3+7ELBEXB
5oLnwRWhxh26kobyQ77JvAN9HBQGkIzkB61ujT4560VU5tGI3u28LeqyBNO3Lyfsnu2ClwCQb66a
6G/BPOKVOYab9sOVNU5fK1EY65mK1xftoCZYs0UC9+h02sLpvUg7qSzrNR/46HGxsV9sePTRK/J7
k96syiOPIR96k5sI0yZ4/381G2QzvgAQ97OFJmb4yhdBhIr3OXltqY9/eX8Ci3iPYRX/hNhBMRGp
yVuiEL3Dj2n/4fnL3vQ+FJS7psZFxJw5C6Yqj4HkS3GdAMM8P9JAYu1asalxKx7HzgDm0Hhzt2ve
KEE6c+VXSMqSrPr6afKeRBH1XUVdo9Byh+28poY3MWorScpxRCzLwlV7K6AfA+xu8auyGP0RNgO3
EcFaE/YlU6VVcOvYN3XGYKknMTacP1LXAmVyHDN/tQ9ebzAbYU5qkUQ9OmI15ykbZvvTYdYIfaT7
0ViNl1yxLmjtioPPUSnUxo8vGnzkvSCevRfwFztTAZ1QXA2s2HxtT1GJ7Zss54D7H2mxNqfihanK
6Wq6kOtA4kvoaZRjEaJM7+c4nbHyiqZ1weOX2ljFVO5LdoA0yXb+qUlxRhbxFd02Z26gX0LASQOK
qv81v1MG1SlCaCtropNJ2SZluVM/REH6+5HEqRuF7QqtYmysQYqmOE198qyjofje2ZKFYgLy/RYp
hoA0lwq6556yFhYuVuqRYH/DbTK45h2MqD7hseanfNduetSrmZNCifSTpSC/g8k6nj5oGNGau1Z9
E5Th3PYdSoGC2sceYW/yFCcEB/ABIkBWarqbC1BQ8pYwqAAI9Zmc8ry8O4IoWios45AN7TWyQUiM
SdGMdOggupygAgZdrYnEftTxMHjlvT2+FxZ3SVixztaKVqiCOa/IhpnbQYrVMEVKN4FDfZTQMvpp
IyYd46tGUp/Jjq8UEi5TiO3nRDbSQjrcyp99GFOxfM//wIiTmvimaJ+vwdjZF3QCy9uvIF2lwjKi
V4/GOcASkK/WLNPYs49BdEdydwIZuciQuQVm+ljEZ0PsWwDbvmmzcShgITj1nYBrFzUm2EhTrMOW
xbpofABIFKuvAgAHO7o0T9WIfitAfkb3fnLQyk+/17zOk6uN748MYEHT3/j+cLzGNr/0plip3vSM
gUmUfAA2eg44q3cBt8PHmuHbi5wDMue2Eo7FpJVvNbOfjJXvQJWm6aKjWxBsL/9xpUNP1eN28CuJ
/UBVtUVpGTBXDflIm0aQ9O3e8+/r9gNFehV09Hk5cKl0JoUselsFNy+heSdUVcGt40UtaB1ShOHF
6P29v5Cr6xe6aTGMwGGWJdLmSJbm/DSHybST7M3IFZ1jc5cLH5e/AldEB+gQ82hBMtgqf+Q0eMri
tPtA7U836PaqGi7evxzKMmvqlG1M/kzrI09KVICkS42nQXxEEH1pndrAh5RpMuQ0ob8EgLl5CUq8
DieVvI0CBvQUzgXIHhKDbUCLC4oYTT4YsU59Z6YkiPltLKPu+GNI3/6hxF5HxCPLEg9Wwkzve9EJ
UVB8ysl076zsI3+pHIUaFVvC9eTs2XZbcn9DaxSzNKNeIbsoDGqTetIuMtZIVv8+QrA2OLvMzowH
RqKvNZLB2oqbXRaoVD40MkH1VHjJ4trNsXqp85WP7VRF0W3BkqoPzBEAZeLlRWeK2NQgkXvb/mfd
q70rbrU1/Hy+3oIjJcAjcoaCy9kO7cbLihYJY9825gb6eDU6CR1CW55wLwqMkTKFjJ81aA1NPtEJ
/ShusdpDf+5lu++OysByOZVaehdN/h8hshNq6OoIPbRkiwonDFFF1kY7/9Gr9W1bLdCeaJxLvzk4
Zi0eF3DHxQgORCo2xtLzpcCWUKL7lBwT+RyBCieogaoVgg7VsRijyFbvNjUW5cNFdQXysN3zNCOo
cobSxYuM68K2t/d2DJ0QvzRga1I1SUxmwI+FkQlervkXh4LHXmdIbcChi8vRAZNIYFBtJXJc+K2A
Q+ljdSh88kGQOVInnrkYpmBGGIgukdqEWn0=
`protect end_protected
