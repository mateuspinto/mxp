��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����l/I�b &+,��r�"1B�̻�SP5��ƗH_��7k��D�/e�3��C�Eڢ��`C�Z���>�渳��_N�@O��EXu��ٱx�7��k�S���Ude�V(}�d��@����9��&��ʷ<����'b߅s�!P��v����`V�5�8��N(�[���tɞ�-I��X��NO� ��c��%,��<=^zR0h�N�����L���h�:q�Rڈ�I!��B{1J\�~��1Ɔ��A� �:W�qI��<2�栕�m]u��?���݃X������+�<9}Y�oI���"p���n��ft��_�?S�����&��lD�M�4/c%�@��%��A6�іR�s�<��E}�}�A�@m��*d	FMI�A�1��7�k�v5gHQ|��,v�O�.C������c�hN�����cϑ�R�)93��h�g���Mz�o��v�X��S6� �h�Px����=�9���&��K?^���F"f-�T��N�B�H�N7y�8\��_�ʤ��Rt_b��^44w9����ܤU�.�f=y�E����M�s���:g�b���`����H:��jBU�v�5p���>�k_�O��f�H�y�'�בh�߬�� ���d�I�ɱ�쥷�b�[��<%�W���/f��^(66�٬ȅ:oAt^<C߻���%�EoF�ȇzv&�
�uP��;Ӗ��T���T�Y���P��"�;%���ifi��>�PR�4��u�&��<��� |j��v��%�V(V��j�/c�S3� ��C���{{����_� W����k���?AW��^��n:W�
��] _�I7���~-��1�3�?��&�{���'�	�]��v~H�*Pp����(k��h� ��лE66�%���5Qx�-]�/%
--d03��ek��?2�}�ŋ)���eIH;�R�l�fJ4I;����ENJ� Z@'�]Y���pϜ��P��>���{�՞x>�y���_�-pi�z���7\VWyA�����o���iN�����"�3���͕ړ��2�;��%Ƴ�P�>�<9�t��U� �J����ROͯ��-�Ȱ���ZsZ|%T-�q1���EF�� VX��%�s�x+,E���:q�a���qS�i�(Vߤ�bi��LP+>���S��C�Eqo��e�v��>K���vC*�K�|'��'}�nU��=��S�*=��mطn>vן�f��sj��G��R�85P��B�"p��b]�ߵ3�:�*s��}�|��o~�
(CڨS�k� {�gN1�[�xx���{�J��#�&q%�)��6ryO�J��P�G�vs�x��Q��Z#�0n�9�G�F��akZeD���ʐ|萷��(x�-�!NO���O�s\L�M�]�Q;�ԂP�G(���|1�ǉt���A�Pw���������k�:��2ڜZHh4���^^.���� �K��ƚb����>�� g_��\X��blZE��o��'�[�7�҈	B�%6R%:Vs�^^f�xέ�Aը@�Ȥ�t�o� k�H���|*�ρn1)�ZO-��bؒ}9����.P��k(�'�M�:��ls1���+ W����}s��*�L�~ם�\P3�r���`�o��XJ�JO���ƬF�3��T��7�˶W����p�u��,,��j���f=d��C�x8���C�3��q��+ˑ��]�X���E[y�m���J�|������D�
���?���"
��:��Ƕ6�\�p��/����|]�m��8�oO� 7��g����R�)��u� ��la\rv�MGiNF�⌣��sSlW54\ːt��yld�� ���BeȨw<!��9��;돿���	�l'A�z�R�j�#����Gh#��8M���G&E��l\{� �!~�K�ir���/
�zO"�m�}4Ja'g�[�]l_�3���I����v-�� �)���y?#�k{N�'`hQq��۵�kQx�;D#k�ŗ��Z;ɠ�N�ß[�~�'�V�����	@�9(���Хl����g+3�)��Y���T������9�靄z$�N^';�A��������B����O7��/r@�YX2�;���
��`@�ٗ'���+8���P���Id_���Oѫ(�U�2�0e���	�@���|*����o�^�jvQS�#�$cZx/���ə>_�i�����#w�;��%=ī���i�:
��OWX�	�T���^��5IjZ���'��&���g8vsCh��ǝ�1��s�I��Ge�`��R�[ɯ5��TO�?3w���9��ꨶD�/������[3�"���쫥����z~\�SIo}�Yf��e��v4p�l���d[��z`?��u��bM����=c`pz3���W�ڧM�O8�z��"�%��>9�"�JTLk�fq��6�5JH����x���-� ��x&/C���k�)�~LH�ﯗb�0��ƣ�G\b|��0賔��?��������,}�>���T�G�$O�q�g��tw��@�օ�X��w���μ��!�Ĉ�Tٰ�!�a�t����&l@J�ӯ㤂T��[�A.ڛ?�t�k��^����?���V^��~���(q�] ٥�Ev� $}5+�∃&����5
���5�f�_q9�(�h��[�pҿ	YBG�idZ��)y�ם���u)�]V,�fۉY���m��Q3�ϲ�ީ�V9`�i��qg��!�Aݙ2#�@y�s�J�@I%�;qc�L�%k�!�`э<.zsɜ�.u}q��	Vj�f��:���D̩>�ێ�;" 2Y��~��/�ǡH��Xy+�q�	:���8^��t��:��&��C-@C	:#B[X�u�4rV�ו�m��9���q^��Bb�� ���q�� �M�h?kF�{�����#=	�j�	tH��í�([��QVcؓ�$^b=��si���Yy�q�P����o�{;��G�x�w��z���&w:U�
��ɍ]H���üQ؏.NkB�<�"�`�Y��H�&�.��D�:��<]N�`fJ4R�>�v��1V��4���$�Y1Ph���h�������݄�+��PUc��
��@*k2]�=��{�c���'O �:�m
3�s.���j�^�h9�S�M�,F�7CI��*�+�%�W����0������<qc��9S��8�-���]�4�u]*2;�l�7X���gԄ�Si�����Tx��κ�D��-ǅ@������:�9��Ґ�-&��r�`<�#Gл�B-O��ћo+�N����w�vp�O|��S��פ7/C�3�8|�I���J����螐~�R&�乣*�Q���_����pX�%W�/m�\�l�Z�S�>�]ȥ�$��O?�
�.2���V]g{���yR/�)(w���@�hUs,���z�w�b�Aqq��f��y�\!�V�J��m.fn�C؉e�1��I�t$$�D� ������>_	��y���ZJ\�*�q��
7MXFG�ě�%=ͧ%�7D�X�&�H�>�iw�P�r�B́ڱef �>���
S3�oM`�o޴F`ؗ@����<���ރ8�����.~4��8P~����+cpG��$�;�qaE�͖�_���k\��!n���$�!||U$O�BO�ȥ78�Ժʡ��∐"a�+��))j>_=r��u>BB>�|=V
��2犇�(�G+{u>Z��#�G^%���������}�,H���GE��h�HK�"4K�aS��/�(��������Nܙ2�@��'�wo��{�ٽud���?@��,&�{���{`Q�l1\�y�"��R����m�2ݡ 0��Y����?s|U�-aΪW9����7��a�@a?�4��Ip�m����ȱ���fkS�Id�ʮs�/�y�
�]�a(�� ��p#b��\���Dz:�t��6�H�����\��3��n"��qpd��&���hc��Պ��غ
�(��&Cp��GH��5|5^���]��fй�vyC#��\�k��05.�A�˜����LU�]aB=ե��4��׏jOe��ǂ�²M�sx�u������PyyA5��Do�&�-)k�=�����|�|o&ˋ���2��d%�Ps��	H�\�.�F,���@P��g����$q��3_�*��2]a�w��0/OU�KоW�v>Z)�����V1Ɉ��f�f�~��P'K�5��rfC�U�@tsM���&C�Z�)jߕ�@��qTT����M�{�����Nܔ��Q_<��J	����y��+�Ā8���J��r�����FP^3����m�� 6 S��jM�g������ɔ:6�.,�����2�5�6�B̐_�(@FB5�B�Jqů����U/�i�a|�F�Cگ<��o꠽f��e����@�7��L�H��2��C�N涂��p9ԇ�B�"���Lc'1R��O�>6����}�3e]�_c��a�������-Vb��E�7�CA̿�}1�\���������75�/��%�U���@Z4�~k=YJ��Us������̀���+F]�W�*̤p��όZ��t�TDF�ie͎7�a��&$Ԇi���\�Hp��<�=	Qk�}�NG&M��So���$۱*wg���8�R~�������3��SY!O�!#�3́�4���|����͌�;���������F����\&	^w��r)*�?���u:�:�Aݟ�'�
�QX����N������U[�Y\��q��{�q�j�Ms���"eǝ�_�I�ǧi�^�(�%DƠo�1C��W��U/�P��r��j��8����` B�>n'ʺS�.�~18 i�<�$~�x��)I��.�_ ��sI̡~emK+29$	v}kip��J�m�K�`��`Ͽ��v����L���g�G�.#�ﯝ�F���A!)��5��w��<b/����Qﰾ�y{�k�SJ��/��ɮz��[ZU�"�����i�S����ݗW�pt��$h����]���`}z��i�����V�]?��5y�'g��j�a�*9�P)���Fx����
�:��+�'H��N!��48�3@��I&��d��ڭ;ª�{�����ވ�Z��X��_�O��C/�Ʉl9��~��xC|��dҞ�L�����ܒ��1T�d3l&OZ��>��^$#)�m:�\@�������	t\����73�L��v�+NP�j�MD  �
��a�#"~��=4\ա��jP���\X�E=�ڄ�;;j�D�D���[K8^kd�Ty���n����9����7b�{�ݾ)��UVO��kF)<�-�{����2]�_	�n�
k�z�A�/Ys�9��q q�Ɉ���srW�ԍ@�|%�ߕ_��(�Xr�<rYǔu�"wX�S�Z�:��-��K��S�hhZ��4��Ac���e�j���P�F�����:Xy��q[����]�W�NxP��A�b�VαB6�!�O����(�e��r��9AM>�3jy�[��y�%JU�P6��6e�#3����z�2�"b(j��Y|��7܁�T�hD��غP��� �'tm^PMW�:ô���Q��0քХiV��h�f��J���O��x���*�<'.������ހ�u��&��5W���$�D��8�9m:�D�u�%����bz��_�G?��u�L���y�Bz������:J�%�sǞ�e�;�&��;-�V	��E�	��� QbuY���)8w�g*��E��`���0 �64�.��z~�s`]M��W�  !��U^�j�\|����x�閲�Օ����	��v��ҳ�A� X�3-�yMwip����!�#�?�fs'd���5U�D+9��U7WW�W���Q�T#O��@wg&���>�N=��.�2��r�*��&R���E!�*-���[�5�/R((|�E��~����-�p�����ԴB�C=z Yt��Cou�ם���.P���PC�`ێ<^UUI�y�WWHA>p���U�\�D«d�H�0ӌ��b�����TH#�pHj��klS.8�e����twv}��ҏY���V�fOT�Te�]��_d�=~�����V�aL��{�n�k���X�=� XDs�:�Nu���i #g���_�c��r�>CֶCW�6a��}�d0Ɖ�~A�������4�mλހ��eH�Ar��Aݴs�����J�e���$�����6Ϧ����a���ьcH����W�?�#4%��MdVxBC�#ZT�K�쪫���P�f��ۓtL�G\55��q��2�kA�:4>-����=^%X�� �4��f�5�^"�3��Z��B0�%dZ*��(7YաD`���1@r��2��5у�b��|F���Ђ�X���'
���J�U�!�w���@�ߐ�ڃ;3����s��O	��q�����\�1NS���H�Ǭ���By�lzkTx��1&ڑ \�͋�'�����)�>�Y�|U�u�����QT���*����;�W�Կ�2��0���n��	���9CҎ�ʷ��$�v�r���q�xխ�Ʃ��Z`Id<�RQ�W^lQt$�=H��۪�_�G�_|BCӰ(�)oMQ�H1��L�}�X:�F�����^r���S���˂d��	Dqa�����IdZkx��j���|�VNn������ �j�ja$����T�ބP���D�V*շ;R�ј�+�>�O�Pf���� ��]Tr�5�G 3Q��
Zg
����$��r��L���I<#ŗ{k�V�&����>l���X���<�,�F�9�bL������<9�N�98z�3�"e��,