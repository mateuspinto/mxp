��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���f��|�DL}6.� �~��پ�S����䖙!Tf����z��ݎ�����:������_�-�1� ���<,��N�-?V���20����P�-	ɓcY���Q0��u���G!�5�ڦ/� ]+|��R`=���j�i幝曡q�F􆬒�*=*�l��DK!m1�N��j�#��E������]���<ch���l�B�j�9�4&�b��]e�|�-K{�rhm���"���*a,I�3�+!0���=��G|��gѩ�nm�����@(�11ST���ƃ�3����V��\#nl)��z4��+�6�k֋EoF�Gæi��xG��P�����l>P����]������T"���1emjy,�o�ԒQvk	r��i�N��l0o���A���F�j1i�S�ul���>�A���0��LE���8�ȞG�h������pشS��<BJ|�������.iR�|a�#��!>�u���\XV�U/y~N#���N��݃�6�����|2.���+)G�ս��!kRc"�
��̇��p_u��P���G���@��Vj6�w�Uw\VÝ@e`�Hyk�n�./��<jNZ���w~��Z�|��~�Pv���T���}�!��(��O�D�Gc�2��7�~�	Y;!g��;��-��Uqb[<A=�!�|�ht�U��`)�v�c��bE��-��&8�	��TQ�_���h�ut��]��c�!�)���ׅ��cHm��e-iΒ�Ę�ė�x�*����H�VD�X�dt���lBi��%AN��B�v��M��Q�������/����uC\�C���K�M8���p�Q�k!`$��<���C�Ԙ*Uy8�ڮ��Y��(L�j����qKb�zd��c�$hDrR>mY�7�c��;Y�%p���"�.�|"MͶ�(N��k�]ɱ�&�)�3?-oiOW[����M��~5���pN�VRt ���1tGF;�i)��d��y4A�{�U�ꍛ�!Ҳxn����!w���!�J1�?㫻W�[d�U��w���"�>�x�p�*�G�CE{����E�cBٍ6?:�}$>��8&��\�Nx�Z�G�SjKsfT�6|5���;�s��㈊*h�r�����2a��B�R��ZR�=
d�ؽ���t����(�������fN�+i'6t1ˣ]hF�x�Q�\Ƌ��m�Ht��ZC`�{�5�O~��05��X#���4{���j���}F4���L�h��Q����
LO�g���1%�$�M����V�$�R=	}�}*40Z
Z� ����d�wS2�&iu[A���o1;�n&�Ģ�oCT�A.U�4`���Qײ���
9���9"���y�L�T�ޣ؈ߓN����\�I&v�4�G�p-@zz-��n]�D�G��z��Q��h��'�ѩ%�jO��CX�E�
���4����O#��Ր!�+>&��s��T�5�<7^٣���
CI������vf�R�j��{dg\Ȯ�NZ0��q��po�9������[%�gQa�(�2q�ԑD�Q"����&�֌���.Ce8d��r���龔
��q��4kzp��Y�X��q��7>�hzU��KL�M�I��W?	�Ur`�&��k�%q�7(/�g�� ,��ʿ��� L�r'G�.�k�Qq��Uux��;,v ���D
N�2|?��+� ��D�"�.��8{�.�jr�E��L/�֎]3.��\������/��y�|��:��U���W���7}�4p�j��7� �o�����~y��RQ�V��~�[ds���'Y7�Bp(��i��11f���^��J��7��8�Dy���7S,��2��:E�I'�L�i@� �[�vz�b/���B�A� ��)e��#;a��iM:��6+�����x�?l��@#�� r\�/�\�wGp_���><c��{�D��x�0c^�j �eO�Ľ�4K2f�?2XO���F��+�2�ݲ�C��z�=f�t�\|E�N5��%=*=:���V�2xX�rF�sL���	�D8�~|H���BY 2��QÅӐ�}�7lo:L�$FvSj�2��'��˨  o�[��<r�����o�;��g>v�4��U�:0���)���^�dU'鼈�jY�	�q����^O�}�m~a�=~wjfk�$@��̽XmҏIv��ZC�p K6�?�$�JQ�y�<�~I��ơʐ��/Y��a-�u��ڋ��f���O�~B~�-;/�'�-V]�?����pы�����U��@l��46������q�ׄ��	P��^6�����.�>15*룺�å:B+p�˅(�ɽ�ȒR��`�C�>�Ǎ��E���襉p~L��0�k��B��:��Y:��"�f��@�h	Q���8�C@��@�L��֊��m:;!=�W}8�y�m�A 8h�>L��%�������.�VTM�|�^�)���Y����z��Y��'�8b�orI���2v���y����S��$��a�wӱE�AU�*�y�B6�Y�Sz]��#R:6�+�u�6I�muj�����#�_���ʨ\��-�l�V�c�����5Ww~�����t�s��W.�&moh�7�/g���\,̑�CW�$���?�ـ���zO���.�J�_�;�������k;Y9<��]6X=Ҵ��T9�j�\W���Ud:�Ì[��K�u��y�Nv z+�6]�9�J���1�0��٤�ٲ�����?��;[$�}AF�с���_����L[������[� ��;a��<�����5X�PMs4w����jZ��� �.��'z��p b�2��8����I�r[r%*�)v 7p��qHʭ����:�	W�3m9&7(������H��Y?��;R&]����^��9�=U���x
c)�I�冔^Ą%��^�@8���Ocb����]��ә(-S�t� ����b/��N��S4?��H�H�E�QQz�dU�D|O�dK3L��$��W��n��z�@s^��C�E�95�	��$�l	7}���S�2ɩءh�4zDE����F�;�^�nvE���E-��'���ѲP���n ��s bը=�G�?�.�����c�:@f��@[��rO&�N�-���@�����#���S�)ץo��T�(��WM���L̟�k����[��fH7�فD]>��"`�����SvChN�I��⮀� �o����䠪��nOM��7��,���%�j�3ч���ϓW�!c��R.�z��+�ߥ��Co�v�R���!��+�v<6cF������[[
֤$�������&�P�
���ZX���Hц�K+�1��Z~4a����Ң�	f����h�U|�젤X[$���m@�hy��ќw|*�eJa1(�3B_���5+#�V[���&���7�<�㫜d~���}b��	�ܳN���|ӯ2+��SLR*(���y����
�pNԒ6P��M��`�T�e]qU���.v��'򳍂�eF2�"�F#M4�קU�il���7#Dd�	�`��ye]vI�5Qx��x�ڝ��U�S�a0o.��'u�X�@��E\�C�u@O�g�+ۖ �p%\ߖ�&�:*��[_f�"�E,�>J:^:&�Z�|�/^�3�Ame���&��'ɍ��$4�(ţP��p�M��V�ͱ�ƙ�Q�����$t��W[��Y_oiA�͂��M�YZrp-�(:��ݸ����_��D��<��y��tᡳPpv�����<w'zd}�mGX����Q�0ޣ7o�݋>�m�ɨ�ːvX��汧�_սcr����s^V}o��A��j���lYEl!���%��Pe�_!`'o���M��Ɍ-ˈ�
��+/��a,�0M��Cf�B�ջQ�j	�����tȦ-$�H����� qDv�3ߕpd�x��4�^U,|���
;�xj�>�iw��;,��L�QW��9���zu�t2�t#���RwĮ5�Z�v���Vg$��(�Sa�>����� D�e���}�Bñn�����ty�2t��)��]ql�=|�n�@ڙ�KP�,@�ɪ�b�<[��s������U`���QL���u%0
�������eܝ?9O������N���b�<0��#��M���&��uj�q��ߖ|i,�'�Gu�c�'�6νeŭ��a�Q��H,Vy�����J��������T���v*2��M�ypO; �l�[l,/.�R�D�����:���Xs(LYF��v�OiS�"�<$�?��"���}\���;{�>�v-�%��Z�
�Nݫ��$�JO{�L���G>ZacS�Z��:1�9�lb@���5�'.��4�t�J�����Y��ԫq
k��_��z�w#>�����K�,k��xgv���&Oow��spf�yJ�-3�]���/�q�����6�����U��ŕ�)k�Z���.���7d����Iw���(�7{S��:qP[�kB��e��կ�˼�,�]!.y�Q�c�۵T���)���22ihz�ZZ;�%d�q�[��=��o��v� c�e���4��������o�Aj�������=tI���[��Z����
��n�"�B��N���K��� qV�R��S1�B���->z��M֐@�`8������וh'`S����F��?�f��B>� �����|\���}ĐEІ�aݯ�B�h�]`n�f�9�]�!���n�A�=k.�)�������.�K�T�wL�lM���SB~�P��I�G�*.�U��FB�',�	���P��V�r���/��|��-�7jh��U��n��l���KD��Qz��ʲ���(�e�P�`�J����m���K��
�s�$�'������HTU�����:)�A(r�� ���%��)�O��c��t0_E���B��;`b���@�b����m^<�*d~S��y/�AŖ�L��8dD�`��?e�CD�Kyb��Eg#���Ub>Su?�q�\�Rqț��{�(H�Y^��V��
����TH�Ӳ����zB�mh��i.��֩R@��8�E&DU�G����r�q�t
+=�P�C��-YSW��Z�X�Yyn��0��+]���\O��5��=q������؟�����bǺ�Q=�=#]c��ڊ�H�V3�gJ:U�f*�ijߵ�}:���r�6K��'�-G�)�+��s��q������&�"G�IV�)d(��L��{a�>4�BP�[)� 8�Xp*i�Ћ�hrh>5�E�T��] *�hש�68��>d���b������X:�q���S�"�LI��=����4&$��>��\ْ���u"6K�Ƒ��{�A�Qz�׌��Sg����&4���'C�n�wc�����3n�׋�J;�S\���ʘ��3��4�z�d���R���t̚�צ�	�ŏ��@���)�w�����W ���@����n*���n'Gm�&/*g��Э��NA�F�U�nD�Y����8��dѳa���[:�0�@vF��N��h��r��5]jj���'圃�T��5ĵA{�0���.o�T���E AC5���_,��U��N�D��	�Ks+�^w���*��q�Ee���Ҭ��g�XhH���c��(,RI���/
]����&KZa(��p���d�CD�0�&�;ǚ\a���e&���a��Gi{b��������bX�G�H��(rt�
8:�W�I��]Qc��W�tx �,wT�QKI)+��G����x��NZ�q�=R��j��j�]�C����1 ��ȸ�:$�� ��p��+�m�_��h`T."0iHy���A%65iI������ 7�=�,��� �+*r6�k����Ǩ���-=��_�G��`�H |k���5�PɪU��؃���4#��>?f^�^��޼�c��^�� ��[��v���b\vu��k�ԩL��G"���٣9�u��=EN�'cխ����۩��(�ȭ����i^�"$�����)�v�b߁}uii3Fǐ�k�N�dS^�|b�mG&%2x/��d0y��`ˋ�i{.������:�������!�xm�>��
��F�"�z�><	 �����Rءt���Z���.�nq�"�ȨL��Zً݊ի_���;拭&�5b��_Ŝ41[�+�+D<պ��s�e�3Þ���h'pg�wWH#)��
�����P�D]�񜬔i��7��Ӵ�d�#�gH��\
%S�M�(ߺE�Rƴ�pS���ؘǳ/�%��}�A�@{t�1~���Q)�'N�X[�*ЬX��u�ZX=�����A���"���u���>�^B����j/W��'6��qFF;�+x"��|-���qO��t�M��@� 
��#>�h�F�8��C��+��)�K��V�u-�D��sOȹ~�U5Ëى����C��*�
��C	i)�ٵ��F�^�1]�_�+�!?r�,�j�e$��>���V_%4fk����4�T��e��2�N��w~	L<[r �-QQ��T=O�;�����E�tm�f>�E0�p.��*ğ���|����!U���ASK�A>��)���%�GD�&,��G�������S~����b�\.beeRP�AM2�b���,��>�wa,f�C��}� %=��4�4�U|3�D.(*7�_K�PȱI���=���WHCP%�X	�*��8���,�:eۂJ8��J��CG��5&h\.̢�:$�4���f���?�\������q~�E�8Nxσ�
�I�W�F�/Mw��?>��b�ǃ#�絅��d�$���wb�e�,z;%��:V�[��ߜ�}}��{�.��R,{�Ƈm�L(	��nXe�+- ���9�S������	��6�����O���֑��������� �QW}��p��W���H|<R��g���V��P��`\�(�E \�������o�T8�K��}+۾��x���zP����a!)v��#L�n~��@Ƿ����y>�>o�m�����#we[�G)��E)ކ��~W�nw��h����$�}��/;��������/���(���X��{�/�*D��ܨu��&��5�Q�ʴ�����0��A���N�Wk�P��k�PO���X}|�%e16RB7:y�H��"��
����E.[��`tꈘU<��/7u`2��C���x����A���W�b6�,�О�ݰ��p��};N�Qj]�G���h�l^�k��"�a� �>�D�R7Mȉ�=�5=��h��y�&%�z��)���y�T+�f6Y�_��L�?��^RH�1"�g��b���rΔ�4n����Ou5!����yƭ�A��O|�߹f�E�S�N�]�춉�G �d��`]DL�o�~�?}&�|��9��4�8��=Ob��<�g�rk|�0�� l,���Cϐ��Z��0y����}���#�}����w[�/<6�,0��	b�[��ƣ�Y��
Q~ۘ�k*�Z�}�n�<}Ϥ�7 5��׊�v�pǤa�_-�.�V�y5rv-��U����y��]��ԯ�9��	`-⣗�E!�ЦMa�.M�#�SGT92GT���Q�t��*E�P)��h`��{[����^ �^�6[�qP3c��s���^��ڔ�='����9�X��f)p���oG�O����1G���W�0�z��_m��}�����g��#/�-�ǿո�
�"Sǘ��O}� �F�7���(�d4}���!�Tq.���!o_� ���y�JӲu0�bw�ւ|P�l߾���e���n~LԨPܥ�毡:�>�5��ʖ���b<[���ߑ!��hK��%w�=.~��
�+X'y@�<�0��XVaB�A��t�y��׵��&��.�#<'t}@.�Du)cX�1�4��^ӷ�jQ3-�)J�X"��5%��i^�2�s�=����]��B4̾�����ڞ�{�Yy/�ǘ�>®�o0$�L���h�4S�����xaD�/����D�%�Lta�2��<���B�C����ieޯZ�`���I�/�[;�����L��i����ts�����> �L~�w���<5<*��"|�/~=گn�+)�n��S:��Җ*b�"�x!�����h$�)5o*$�L�	�X��ӏ*Ӓ)�\Z��%+f>i�\hO�B��AuqRź�_��8_ʍ��)!��x��Y�4��ݙ�`i����a��girSD���y}z�!��F�Cht��� :?��{p#A8&�m �~ i8�?�/��n��h:/��q[}��r�q�����2Lh���LTh�nՋ��Y�o�U�	~3	�q�Pi�Ϙ�~�</��f-ss	�a�oתF�BMq7@�h���8]��V�A{�pE�dU(���
�ȧPJ�c�bޜ��x'G�vF�ٿNp��_�M�t]�ϻ�)���so����#�_��@���T#cM�Sz��W�pN��^u���x2�\>�6��ށ�s�&3(<|�5�|�mD:�s�A�l��}�p=��~�tk���>�D�%�R�� �Z��%�Tį\����b��r+�����a����<�����WG�n���K��k��n(I\�q`l\'L%kGH�C,���y=WA�Ci_�kR�7bN+
B��,lGEp0(|�뛭�����m�zF�#���jRK�cش���\���񂦽����y�V���t}�+/���s¤	���q��/%z���t@����2q�3}�]'�"C��'�$(S�8�Pc�a���G�Fk!�]îSLi� ���v>֎N��:Vr�$��r�ŻS������_�������
�$h_�s�5�"���0(����[���w�Z��C�h���W �[�0�I�2Iv�OOh�Eb� s�H���`J��K0)�IwȒA2w�2�K)��d}�]8�,��+�G�f��A!n�]S��]�#|�~��˞$���r�h7�IE�
�jQ;r���*�ip��1.��-��V&�h���=C�!�>����Z���S���fB?�;̅D��Da=����|���x�M�"��>o�c*3����;�p{�T
�����+��T�X����2 �'jc8��o���k[�R��Z���A �O��W�x�U��ms?�̆�3�8�un���h;�Jb�_�)X=/w!�L�ACf*��b)���A�Xn�X��L�^������yY����"���yώă�� H{��~�qat����9�V�P��e�mzA�
��)����u?A�R�������2�