`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
YZ1XI4y55CZgce6GUrUYE0dIPB3fuLTV2Sg0DdGscBL58wDDnGArk3VbDJql9CkRR0gPKaE7U0Cc
bvyiFhAY8LHojHQgGgUu1JdZVQdmLgHJ2GEm0doTbI6n9dnGAM0VBaQ1dlIdPZ/hZ03Q+faiCU0l
6xzrCiI15dUY4eEXOdZn9xexgPyS0p3a3sy1NdIWOcP0qaGq3fVOrxGRB4D1CUCPVxedC3qf7JtA
unpybSefNhnIJ2jPnBB8lcL/52XEV83Jg9wyyEFGzQ4nE9pj5xvQhJLwid7zaRGK3hmTH9lsvwK7
4jfoONlZxi5zVVtWwdP91wdHNuhWFBL6/D7DZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="Ki9ftUD4T16DqC8L+7tg0ls4I8DBxRXoPeLpd3nilHY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6528)
`protect data_block
SUd9j6RQktjWsLMhzsdWhSaVFCbTeczkJxIBIPNvT2VJU4+ZKgLQ0f2Pzt2DvHa9qWVx1SK/16jX
qzK1cBEz0RxeViUI35Hq+FsdHFu6k6d+PABdSmYOfEFu6qT1U7Bxx6UeyX6D4nS7bN/nzKSh1xqc
dNFicV/ogmznxq8C+GQCX9pfvw4q5qbisQDpMHfbqRubUlCTSecDJEGjrmRaYJiaZLXK61PNJliO
jN8DSp9EPbQMD/BDIyI77FUnjL0mtTx838ly0MXYG/rLeLAIdKEUSR0vxpsZHb08Za0UnLrqdroV
NU9/+deu3RmBPWo3zSzeqBM25+29k7XPlEyreAlAt4ZyvNum4zrZY5fx6zdxj67is8k7VmX7y/3+
oKj7ilX7IW7R9CZP80sBNTwKKUycvh0IUA2YF6D63cISYhRSfazznrXCwwnFWpvLqZH9FqnFcfv/
qTiiGfVkGFv6fe8HgdtzaO/w+ePx+/9jS2/gj6L5zEnP5qdhOYUROlZ87XKZVSPdusXgJgfP+Hnd
IkeBTha0WCyxgKDMU12m2DMdnHFVCA7k+kxss0xKxkhtD+RIsDzL9SY9ldLtsUvy2cCyneoCQstN
IAa6ZgxvxP1Qd2SPBFKQcbA2FV46rGd5HCvaq3afwcuAmkMZpU0LGkv3eHKDJuzAnoIA/lwySNud
OlyQK7tGyXNtkdTx7X8NJYfqVE+rbhL7I1+csH4leV5/saCwqEF938xLxYnFoGDcTIgk4RtGqj3o
QgzXtAqgEGq8pqyuQeJUNXwl8NapwOGMJVLpGDpyw1iUHoOKWH1k5U4lENb38nP6883mzgFBNci+
A01CX78SIDwB9E9W38dU51QX8ZFW32ErxDaM9Yw/Dt9BKvwZaCD1e04JWyopJIvwagvABH3+IJfw
SAPDomcTOOaAQWL3q1/IavawCxCfsQj8P0K6Iq+rzK4+AODsItWVUzS3u5seSbzbSzRC/WJMQF6Y
za4ko55j8MfME1CfLWCmtLTi+mAxX+L0XntMz7tpkv9Hw6k4NQTsNnDjeUpfwPQXfAby1qKGGuwL
Ky997gyIfRcXD6zSFIln8UVVOFczyaiwrGfFpm/OfixjMZdIqWJgjTyhmkaauOt8IrhGVbRmtnR+
wvUbbr81ivp+id9Fgku5zrVt2BXS+/7ea+nNUfglwRPnEl6YTf2NKHH5tqxDVWQjR8Oq/qByjg4G
2DBqJ3hQOh6GyQ2H5+JoPTvSJEPRuFG77h+qJLJGvVYkpO97PGGkEuCvSqBZ68PMWwtepvjJbjVZ
ei+sjskanA7/PExfogEVx9Vn5kdidRPJNIoiru9Yzz1DarkTDqEzOpOM50Cfahkn/6OuV/aLZRcm
gpSCBGx8WOs0qyLMFpdtDVGuj5jP0N74t3OisClHdw0MYDE8067FkFO+tUf7GDZ0XZsfHmGO5zUA
+wPuaNI+4zNX+hGgdH34paTd/2WAwsdF6Qqq/uC2MUDRc9ud/YOcKdz3ckPRHjVeI8WHLHNNUDVH
pIvZ8ovGykDgXIRKesR0RslGd2+DdHqke9B12d9QLO0iJzecuGyGrdhkvMtH7o33LRlnd8eIzo57
DgaA3Wa2DEzVqyNJJlusu73Ptkkq1i297gGsuALfppDrF9u4SPJ5YT3mX4ou4Pe0MCGty7zgbWZN
BYpoKGi2ZMC873/wRYTKkNWGo2AnSky/k1YO4KO2Pl8syemCv+msQQqNnIMwrek1F0iPfjxUAy/S
dDcDS/3YNdQiLAgDhHd0pUsj1qBZsIY5URYPLGO3bSs9U8KSIsPCGWOSikGqflXbYUVvjfXpnehF
CggMU8upy161pWNXFbQij5yDmE82AyLR7CN/NLlDbv/KTP2nXPNvqXWmv0SQRLrE5ntf0XBuD/u3
izhQG9w1NVHYmMHnsL5pc1o4gHHVXJ3HBjlTgGrkltaGabtcrHik3fBVlH6Fm8bwEiCL0vRd3PJ0
BUN8A9Pc5Lzzq8e7kEo0Ia5m6FzqotI0nKPIykHq3gu1Fj2zV8eCrCNmO7HlyOS0RuRPCW0qOaM3
qnG7mQimgwt4G9DV4YnHuzc8U0oSeEtl+lR4sDKk/za1v5UuFjMEwZqP9bbpKSXyXfKA9Mt6K4FZ
maVUwxIGQ9ffgKX/lxuenyCE8Wodzp+uYX8/uyfoY/RU4lJ29lFtI1APtxLuEzGMk8/s4fIxpwHz
Nu1X2JTG3lRFy48ZM1OyIgQ2ckU4TX06qrEej9NecwhcY27fKKz0cdargLIfTxGVDTsSIMckl9e3
EoCmYLlIMu1dc2yL2Fd/MzSu4/vcaNd2LJx826TIsnerilh71zngvVdnFVxDML4t4xUeqfr0aCxi
5czUByFCSe69YaRCt3vwr1wSs/oM3UTk+8m/WAh52Z9IlkP7Ozy9LyWyFwxhHapwwaxMN56VGy3B
M+rnJ/N+i82PdAl3TeFc7xJ6TuUHhPmGg6SrsEO4Mcaoda2rYyc9fcVphKXxvLJ4GV6mitlQp/5+
BD2IiOtFTNrGp2Sy51yShjiB7HXt9lXYQe6KjNzdGjPRkMmkjAIhN1H+wbxCr2rwphJp4b+v2qzD
uMj2Ys3QMSX1WeTa9ivpadZ5e6+kEMUJXrIqWtK0+fPhobtP01oGHGwxs5BX0YM3zf3NG/5oA8BW
dKPYu0mYytOFkyo2Oy000AuU0W6a9bDXwUuWAF7lYbJ9C+1XL6P5Hzx01JalwvrF7OSBEM+E7roi
AGkAvfhkeAhQ0rjwZm0X5KUC9VvhJWqw4wqguSlmYQeDTHDwwSYeOdZTSN3P6iH48lzqlG/Vi/1Z
VYq00bjaedTctaNrsU1uZvaMjg4R4ucbsZeEtygb8GnEVPP+t42DDd9LfptshrNzXS5sdJHwyXUT
XwOUpXkN6yIKEhMgVBOnPTcW1lL2ox4ubK5riSnTdrdrFKTTGIxwmS+qNPXVm2/r9oTQS6ecKhn+
w88RksGAjakGtz9xO8V0mY+VqalfsAJSMgVQ2WNmvp69Onn2chzVVhKSSKZ35Hox/3AQBYE9mMmt
NPbfi+RRWLab/TjgrAeXAxE3tjZVwLg3aWaExMMp/t0zrN5njetorUg0itNdw6/bzCp8pyQPRZQf
YMfIx3gprQj0AkcAsJgft6PJJ5lAha6SG0MtpFv2wrqGWuiRjdKZxpjrnXHkWaBbF8C0uCADHgMD
qnNyBuhvgiTW5IeWCZ4irxCO2L+qGywPirD1YJWYXVvS29X/F7Q+PJzgIUImOBRMpeuoFFLeyB6I
pUnGE1xoxDQ6x0tMJ0SPemhClPSPqobviQ6NNonkuLEicLXV/Yc6dvMBywlaKFI028PFmNJ0yZ37
d4w63lekcGPxpofZAydLvHdamEQEa9o2h68Mz/R2OnNHDzsboGGGKb92CZR9BGbfws3GzK2t/PPp
NyMn+kobLqgo5nXZsT/E8FoTS7d8zJQCU7HVgYTJk84oelN9X1qZ76azunz/PA5U3BNQzxboJYKA
2GI0Tf20Z+PAPrOo0p+xx71tSpfYKF938HB+q9OaP3lTY1iqgRSCwteVzdyFeJY7Oabs1QkhahLt
Wn78lSC6g1tdLehLVp+blRUsRClyx+rW7zEGb6RaxqkmpmRKi9bw2mJVO0i4AyIag8qIHCIeFVyu
jCBxfgCBkb9jAj/WALSSQHbuVgiVorbk/ZBtCOtgN8XJpK+QOhiNaDwLBGYjPSEmei61wE8RfcVb
GQH/l8VrcZa4Wy3x5Uxmuo45d7FaULDcmOeHlePPbbue94pI0uwDazxbinEh81lAnKfwh6+uoNZ1
xmGfOy+PNesHDXE7L1xQ/aBUfZnJvP2nu2MNkjaxsVL/yvPjp6bnLOKxRgEQFsbFuV4+vaVIzQTh
Dw5RAj83E+CkO8U/vPCdB+gJDm2STXJFvJriCeTZLSS5YC9URmVnyFv0bo5pc+q9gBpiKN6q1keH
hfzM60ro78HdJ3FTs9jlQ+beIoPe7VxLZIfusQBu8zxAkquKbyWSTckJtGR35WuBk0MQiRipk3F6
WdneTN7ksmVxp9JrCBXtWxCW+5Pc+9iwzX7aSX/wrxUgSPMIYLB/OKWQBpTGIW5LmhLT4GM4cCJD
YIXyNSEal/BRouo6QRMs86Nh65Nmq/NA/F+anwIusoTYwLCb6jBh7aDEOjoBycLcA1N0JwhAdOvK
ul1Arj82qeO7TmDTRyNCInpnuOK178Y4W3lqkbO/EUVwzivPrjXi0EByj7L5Si1QRytwYVAW42qX
7IUOB2TDGRYLqm3AJW455+D5j8tnUNWATvpnh4Zl6J7EItwYt5uzcmXt7S8X1/5DJwAWfJjAW1tT
c2oo9CbW5YdId1Y5nsxZQBCBlEJ1guCL9UtIhBvA4eLeNDaH6qLhvqR9DBYxEoBJonouSo1SmSvV
uKVah0tpOrMuN1FVNhu+EcxoReao8gZoPfG6QW8rx6nIFbW+2ONGwLEd0QxnItvPVKF7e67/Beow
sTWztyJxzA2hSiIPilVMe1Y0g9Z1cfb94X6sm9iO+JTFba8LpCUW7Q94rh/dqaOhEbh5T3+hlF9h
iNjKfzGREQGX6o9oav/FCjIsFv9/CM0BrjkNPFwFFQiiH2XBjsNAE9kEHsUHr+kC8Pi01ig7Bx3u
hpzz7nMjlon8yygQTpev69QB07mc6W+rd3ZBf80p3fxX35M/Zdc2blfi9UadQSDWlUMR/k/7uI59
hfHzpHU+rkqPDOyOZn3BVPCUZYX3+IB5uqX4p/wiXj35OCXatbwW13fi8KxVs9PV7gYK1jb93Ibm
IABnYfpbjFOPsFnzfhzPLthtNi9nbh9/rOPn13wFYlozDjx5G/kn9by8ozl+Rqt0k06pBP3YqFhl
rrhq11CGUkcOsOb/qs39jwkTHEfYWUKpFQ4qijb99/0OToo1fOmMW0ZhYUIfazzh1FP6+WKBmZzB
EgMQG6zNccTyCCA3XVxUU8LFp0+Wz/e5/ntKIRWWJPj2W6esyIrLfEHY86Ytoc3+HfOaiJflamlO
wENYYrbCV++KxTrEV7XVMW7Yqr5x3gPfLMFKZRjkzEjQf5fRYNeuTEsqdoNsh+5+JrztUEQ9dYVV
9icPG9109gjPwTuxv9pxgngP+cgdg5BIPOGKmV/kE464fXNB56qxokeYildGT7DQysnCPpsYiLln
an8pKnU2Py4QgPKD3gjQVwVMFqetKKTf2X0admzTI3nX7qPnzaJU9a+iRZ5CLnrR83Fyy4bq5WKj
xWtt+rS8fkvB8jMNmoOPihcBteI+xxq2GcJJYIVKeX8M0I4fasSrXLsBh8KVQAOveX+iFibLcrbG
9JdV7iSEJs2tGeYm911HvtcvggDEI2eg3a1F3wN9dunhOHXh+e+FrOJq5KEhIMNnZnRWlbg12pwT
8F1xJJkoNRBFb/3f9h/5HUcREG85Yj5SdhQxMd8FkuZUrwZc9Z2c2YVzuKpLHLrh9yDd69U/uWfp
zOLYyCoLa5aK0aUp+FGgMNDTTBRV9iou8FJlZhFv5j9XqtbjT41sKxDHdUvVskWG7EltmGvOvCX9
Nid3Dl8VSwMgbzeMYdmA17sXhjgNQCqV5tch+QojppbpVtnpXxv8axJp67SPEC+gNlTX5ZDgjayK
s3UhDrF3HpAT2h1nQm+TiUHxIT1SaXSa5JQvn5e7zynpsVC9cCMwzM27GKNe7tF2XnJIO5ZyYWGI
VUEBENErGcS++MhtJii4aDYtJVU8QBEhZ5xSHBFMyh6fwCv3sq0KjHv49ajPuxbp79u/GmKQJlTs
5D0P3KH41WatKT1CBm7ftn44UJyym43ej5upAeP3xxhNmgt/clZExP9T9qfMeGp2lUvIvcVgjX4a
bgeWYLbj8uoX4wRw/og6ob79N7Eh7ighXc+WwnoydU8hRKZhL7IxLXHSxi27/B3PyZPf01vk111R
tajASDA6LeBY7uEPp/OBRqNfMvUoAB6JZHR2JiPPWHylBYBeQ27buxs6puwIL4tfIruktRsq6pZX
wwobmOgJ5/uhEci56LIkJQOuMpk8YGnW0dG7wdYhqpTNDv+g0u+CxhY4NdqZ5L+kSrLeiC3zgIjC
4poHuCoQRZr60cKr+tLaXCaz8z4RZQ2cOdrawAgTuhnem7bIG6V0bed4ZKxnYmPDLL+EKRN+jkme
E0sMUfdjr2LPXikZ8K3sUM/1Yd8EsqY31GLm/ECIuwZXIXpIFOxUy1C293YX5/dUl6MAQ60oFq/5
2ccIRt30qSPpU7X/Zfbq4gn9DZtqKhiU7XsVH1hfLvOwNTK4Qp1/11fI/HyM5JQ1ZEJvZfc/QOl3
hFCqgiLzE4Val8kAp32X41FdW/DFNOoV2zMEvAsHVXNTMPUiyGPrnyaol8x1UKcbmXUQRTnS7i41
GnYyf+HeYVO/TRgzlSWfsNyuxuqmTivKQGDh3QKuz6TipBO9Dy/9LpI30DhDRBtBsohUd913rAmr
ccwGPTfb4GkrfIPUuBwaT6YJzbFOko8ijF1NSr0diUe3ixSLyO+pSQXcJyGlnBVesdLOu/XhJ+Kg
YLlTB9jyDaMfAz6tyamz+za0IONswiOPp/OecWFCSnzN76sPTUyskBdpB2f5A05z39oM011zr+pS
GSCcIT70W77hABvSKX+Zifi30uSKBjgU1p10oOzMPD+5e7WWcExok/HuOxl5GXh5aKzItOKrREuF
CJx4xogYS/LiAnJ/ZmmzwL9i01YDuVykrGOP9669aogKw83PTWjV8VkEbpEgMvKSwLvuvZp+FPuF
XHvDpyIMnobbjogd+DCmnnn4INOKQgf16Ctukj4oWXuYDpNPb7sLsDsZd9SCexYQkRZTWZ7FiTc3
eD9IUYTqxQ24u9v3zSt+CHfZ7unPYnESb6IEAXe6WmK2yrhACJHNYHRjb/QPf+9XgWlfJ3VPP1CF
i71dCBzbFDZ4iTf2zw+GK+t+WoK2MLHBxWeFbpOjcSCKEZxvUwpoNIguK02Y2yvdHWDvo90VF2to
iLGnyPfn65uSdBKtmw9TffSUa/yz/HZQEtiMREwpO57FsXffFtzyHMRgvR1pQQathNwb+VVUzOIZ
8Wvk5n6aXLUD7NQA59affo23L50Hfy6laOn4MXv81jUuq8N2PYCepDT1briCmbOSzAXmPMadwTTT
w/KdxWgcgffWRggqTsxecjgk8Mb4cFfN0CFLGjQmAzcjrVp+kmQ1+LaOvmIaY1xvM7CaBFj1xg/4
KFUdXz1eL1hc9tmRjxOx/eTbaLRH89OQYCzsKLFm3v6+/dKoMx4C/7lZZqz2zHmBuYYI+eHuR74K
L1o8NZgqJaMw9wxx38I9212TE9oK9NpKaP/cOwk50Q+mayZ3v9jgyGJ8kPg1j1xX25wWZfgRe39n
dZhK6/CjyNxOcLDS6Tl2Hl1OwahaL09VoeM9w5iS2EjPxDhy38UdOEk9MBBqa7oxhj5F+fOOnm/c
9O8KT7zJCplDe0hJ8y0/VR5NZlDApdZ1BryW5qR4BQglHFkqoVQg8xxSBAcez6OluVgPUGdgMCzA
l1qeQ+bnIOr/eqKII/q19GGYfuRdSCzGnvc7B6UqOivaKiTWtkdQWPELYPfFVKhvz+X1bRihI1CO
mHlNo+DDteIUKWIjtNyTyY9zlWWO/lNjKFUvPYqrIeDqpBsBgXshKZT619QuHJv+EbbdvUUejfEZ
AV2eDCmMSmX26QqsEqZV3UtsEwM4LXEOSG1db1blzijfjKe/4ZsE0D6hry/C8BHhIbwCXPmr2MQ1
yU3LaREX4AdEh7qjAqilEzw26pdI52Lunb8j4+k35jUzKlb6qc3H8gSXAPWdCkqCQnuLhXrPb4Yf
x7DURYYyxx/CXBQjfIybDWd4Rre3Yi+FLLwNJeYeR4l+KDzFgrKimT2NFwUn33FtDBLSzaXs/Q6Z
MyyzDId70ZBQbcC2yK6gTZTVaK1f2e7CLHVJQr3sXMwGZIOLhwivy5p75iA4Iu/cp8EmNx2hxKTs
KhGW7Pcoi6oD7X7ah4zDWwprpv1568floo6v8ozaUeetaSro4ut6rGwd6MLlJvdr9ZOKjct33jyg
ztmY1lFapbW6J1SXne7gjNxg/6FbHM4goLl5vy+c+AXKI0Ic35BQ1HnPBIkSqDCk6Z55iiiuXNHJ
Di2Ot77PO5oGMgBb+g4csncmr8eSlieJOQ72c+SdxxFBIJAZaEYK+TgxEfk2C9J7ZMP4jtxSDB/P
QWrKMWeJbIYNhf4kavLIW1VIKTcZ/+TsUnUGVVbg4ibDgNcRDXa8y+AaZCowkVuuAXpkZrSy0DrN
Chztz4c0TalMuaMOXt9f1Z5+rODMeuXL7RIbn+Ro+WyFZ3lg9rLj3ofl0H8yRxODxhKM0jLYw9ej
0eefJ0SWkHaI0TwzQc0mw230NP4TOkJY6v7+4auNYesC9T6fqS6eQ1TI7PD80gAnkqLTDVTtQP3M
XW/EQRvvYqrujMZRtcDmdQl3ecuVlfTWgU22MaP9vEq7g1Ow3PdQ07uOxKjzQf3HC81oBxCP+Ojf
mSZIqNLMy5uD4D7izUzunGt2GfYI4EzA6LB/btI6WJRRIbISYavBqShqd3L04zfasQQ+zg5qdDW1
zRbb0OURYNIaDROZUUOHukAT4JXQv3vKNT2zYtAsqwTEsz1pQjfEbNKB6oaoJMKc/YnrzILKKFOa
vBRhsxVUAy3qT7g1oauHnQwUL/g7ezyyXbxe55EX
`protect end_protected
