XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�q����FVp�}s�#���ֿ�_�E'��!.�����l�K��κ{2���z�*9}�w����r���P��G?�K������}X�v��o�I$�p�=D������l]�����--��%�2۰�y{$W䩘��,I\� ;���ҁ�%?"���h�u��ߐ�������"�7{Cm�	�P��^As ��}�g�R�/�6ف��a�Xv���D����L��6��}�F��&�u��d�#Q*�C��.�K�p!�|�I��O�bx$���5�%�RP��n�m�X(M���g��Р#V�f��Q��s�0��4�+TM|������;���^l����E>ٌ%[����)�� �BF\�T9%_Qx�QK���� w��N����cB���\�G��q��S�٩#�K�x ������g�2��Q"dz�\�e+X̝�cJ~\#��p���$H�D㫩�����~��ejw}x7&m|����C�{(�`�(���ݥi�H��W:RN��ⷚ��%6�B���J4�v;��u9��{_��3J��dH�p�]P'��*a�G\� zFJ��{]m~��4�.N�:�� � �e�c5H�M36A�P�k$s�{^1G-��d�6p�U�@�w�2�����P:��#����B
�O��0?9�X�-����c����9%�.F��d���~ �dQ��;
�-Dd��1�q<��*(D��B���v]-���)Ќ.k��<~=b6���ٳ!0��R|�_e3�d�XlxVHYEB     400     1b0Xݵe	H����~q����[�ͧ�Ro��D��N�Ƙ��L=!&��<�kՆ�
�<�e�fX���=�=�Pu�]Gu�&�+�M��������~0�\�:��?�f��w��`��γ�z57����S�tb�0I�cp����ϫ7�4S(����4���6�_<�����K��I=O�<�0��E5Ƈ��i���{_�f�������C���j���y�Kvm�09�|��_N�w9s��l��0�7�~1���xV�|�����PlTA� ��^�,U�l��NE��nȝ�5�0@h�&7K� ��|'�¯�����+�#2�+ش|�,���Mٌ_A�ŋI,B�Zr���1�nOx���J�ZG��I誼 �4TD.��V��@�qU^�m�rӢ1�
���!hTT�4�7B�\�㞏�%c�?�A��&��ZvXlxVHYEB     400     170��l�j�2�3�.,Pq�!�2+7*��c�$�_��ñ��6��%�/��0X����)��Z3'�Z��`_7�g�>e$��k��a⟚������8D�jK^�=���"N��w��)�떫��r��O�������n%i&<��@�����VD��<;�		a�����qO��4����� L�3u$����/�ߑ	;��H��0�NkY�T�I��qV84���s��V$_�$���W-�ћ+I�v��={��l�-2�9�oY�J�)��h꒲������i�B��=��y�ЧI��Iyj�Bi7	^l�(�d���4p(MzRL�s��qL���p��p����'�`^�������|��L�L�eXlxVHYEB     17b      f03��~C<�D��p�	~U!�����9��C�pd2=�*8hTd��y$�˹jqX�
�`����v��Z<@��.ˉH��	�t�+>p����X����53��r�*��P
�?�E�,�=��VU�ϔ]�wp>�C�ʟꦔ(��^ 5�e뺂�.�!4G酡���q+�nL��39n�RU��G1�J�wv��F�~<�z�,�A��)y����f�\
���xJ���"�"E