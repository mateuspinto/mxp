XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Wr}'�i��eVQڵ��!�Y��@�������}���qDD�����Á�[P B�7���F�F�L�rI�'u�+�RM�����	V1AG/]6`���zZl#>��*���["`?��M_���"�_�t8��@������Z�q�4T�tE����g#k]��>�@�j��c��"�I����p����\O��U�f���`
i�;�uv�F�T�^�!�{��Y/x�L��ږ�:?��<g�����`�W�k|��ZH���i2ߚ.����-��F'` O�,���*� -��>/@M]h�B��K(�?��ԗea!���>�S1ť�
 ���h�W�Y�K�J	�(}3iYO���ʕT�k�FL�<�MI�v ��oo�>��ۢѱ�]*�� �t��q^�R���_e�,g�43s��D����&w&����_�``����0.��H�hr���j����â�%eNY?aO���$ӝ��ꖰ�{�W";&0R=x��bGt� �↔����T��4��P����S�6-�矮�K\\���"��7�A��Àq!^�&,�+���7��zs�`����)��>R�FX���|��CY�h�!S�>��_{ڢ�W����/�_�>�9�ŏ�퍦 �(vZ�(�&�G�����5A�8INi��0X�x��r���D�0��� ��V�j�"{�4��_.�7�u�y
ìͿ�4aR2?�>h�)�e���?���[�p��W�J\�2�IK����XlxVHYEB     400     1e0�G�r�/-��(�vQb0m⋸<��֪GP�)���.�9���|�ʈ#�:���v�?v�`B�Q:뤠�̉6�B�2�{Z�.yx£R�vY���D`SP�J#4�3�v�u�*9�Sݯc�
���h^�-�������M�{���:�Rq@�զ�7C���9��L]%C�4H�G��w����ȵ ԍV��_�9�����.}�`@�t8�p�\[��?%b|BL��m6Ac�f�� ɌK�t?���Q���a�m�;[�O�����Z�T�;���M,e�ʝl�XŘ���34�����Yq4��?@�g�`W�`	2��bC�X�Wb1~�%�H��U��&��,�����Ȅ}d8T��Т]J&C(�����¸����/��5�6���If��$i�O�|U�@,�mK����)��㟓�BN{�MLA��2�rA���r�'dw�3�lI��2�x�}�XlxVHYEB     400     140�8� l�z2�[��u(Q|'Y�-��]Z5X��4P�� �!��U�Y�S���3s5�6A@F�49��j�U��6�-��H�B�u�d�x�z��c �$=.��rnȄ���?ps؅�3�0f�wB���v���m�#�`s��Zh�H���A�Dg*N)0�4���G�$.��3�Z�!#�=lf�r&���".H�f J���O�Q����"V�1��k4���לi²̐@}���X3�`R��Z�!Ɋ�9L�Or�G�¦Rli�-�f�m/�Yԯ�>Q:��a1*�m�JR�q$bgAYl��E����{+F�Z�65�nnXlxVHYEB     400     1402�Y�w�?��hbr����qI������G�m+AE�:�����J��o,�C����� Ƅ)�n�ʖ���(�8���"��f���c@J=}58f^{�e�K�Qw��P����8����h&p�����ي_��İ�ǅ@n�٢67~�&���5�K����')�k8��Y���%l��O{�o]�u�����9[������꠻���j�6bg2��yk%��lQ)�*�P����~w�6};���/��FvyrW����G����
�2/��hA��KF����b�Y.A�EfJ��{Ь���yg�@ ���5�e��XlxVHYEB     400     1a0�7�QY��6��C���^Ȑj���#���=����>Շ?z8��n�ay[�R��<���A(C������{b l���6*�.~4((�&���L*<��|jL����F�����)��l��w#��QbvT�)�֔{;����M�	�gf���	�ӽ)��*# ����$/���	U.�A{�V��a}W�e�dH2���|��S���L�R�m�]��ʮ��S���zW�W����;#v<�FH���?��n}2J�L`��ʌܐwb��@�j4���;�q���<���V>�D`+�{4��ε���)x@n���Q#]��;��c���В�;�>"�*�ݮ)� ��v��W��I��C�t�u} &����Dǫ������Ы�}�*�b.mt�K�Yl	C����Z�XlxVHYEB     400     130KNu���� G6���E? ������������O��X��D��˴d�r�� h��*iM�e����@8�[�Cn���\�^yΈ��de�P�|��U��1gU׺Z����}�ҩ횋,]��E���Ǉl�ҿ��� f�EnQd3�*�aB�(@t�&�e�r0���a�HGۈ�0t��<�m�n��@�ׂLOz�M;��V����2f.�'K��AU�&�t�>��pbMϔ�ȣ��[�*�wPL���O�G�Lh��k\ ��g����jt$ٛO%g�"e b0(<(�% �-Z�6
�ބXlxVHYEB     400     190'O�w�ί~��<����
HJ���fk���.s��[�Ҫ��3�b�x>�hй��YHa5ƪ
=��D��(�������6�|戂�N���<��I�4�X	:I�aS�c���.:�5ц���}�bB�E������}_�D���	R����f~�G��|(���YvL�R���\��veܴ��:T��S�|���Wp8�vigoT?=�n�L���+0'q2(���Î_�!m_�O�F��2�ɶi__��og
X�nl��N���-S|cX�"���%$�a��X�������GM�w�;����
�^҇P�2�0�:~|������C迁�H���V�E������i�"��OΓ.t E�/�� �~MS85��j�R�&�:_n�E�kXlxVHYEB     400     160e\��6Q�=ct���*T��S�>���,٥���@8�";r�Jm)�\2q3TM�E��8��5yV�F,�C_x�)��"E�蟗Ǫ��}˧P���Fϟ����7���{͞�ST!�[zoXn�kM+U�sLyMh��V7�� �>���u*�|p�E9[��$	����!��L�l���J�K?~z���j����@�BU�:`ֈW�g~��dOGw�VDr�PvZ�c��\@`G����q��7տ�%�N��9����v�HP���`0��j@�[��l�~B���l��6 �<g嗴�Qe2%���B��J8y�%�{��Z�]�M.7C���Nfx�}jw�W��˟���W
<XlxVHYEB     400     150Y/�N�X���W�2 b�NP�Y'`��n�RJ����0�cN�o�fߤ!�J���4z��]��.���?;�""%v� �d�>�mn)���R��L#}�"3��]k���b���_�7�!�{�p�0=����:�;Ik�TJhb5)oP
ۀ��������J���_s����R��9�q���2cќ#����A��(�%��9�Q�g�&n���|\s"�����.�/d�yG�_���� [��;��D�˯��~r���nmĝ��|Ok s-��K�����Uj\���6�0�����'t��Y�T�a&&�R郇�$�Ꭸ����ӯ~���XlxVHYEB     400     1b0���G�'T��6O�B�%�ɮ ɨ���2R�P�h�tɿ�V�Tv�:N�K~�����|;~���JBʖ2��w'I��$@޾��)�u��W����R9���y���?�����S�D��=�S�Ö�A1�Oۉ���s2<����	���2��,�0e~�{�!i��Hs}�Y)�Jo��>��^�j�Ό��gI(QfK�rh��Β��� �N����֔Z�t8��{�g�CU�y�
��Kl��c<8k�s}����Ҁ"o �~���Tl�����n��'����_ݢ>P�ڍ���qO�;�����A�+�\*��3g�f�/�,���[[�o'M�mQȽnnUf(d�r�p��ب��RL�D�zuE�rA�c�\�&f�/?�2�ec�6��ޯ�4�O����o��V������+�5C��h�N	�)o�XlxVHYEB     400     1d0S���7%}�tC����?�b��B�sR0���P�������p��I��&����ASro��H�d���e��$�� ����fۏ]�����[j�l��躞���{?E��?G��TsO�4 ��2�����a��W5u@��P��=��0(Q���T8�)�z�;y����z��E�}�f��R��Q��.���Z���o�t)a¢��%���Q�W�dWK����\����,#m�)~2��҂UI�&l�W}�~-�mi�`���^������J�F�ቧó�[ ��24���ę��y��V#~���4���
�KJ�\UpKRl5E�IDiimI�J��CG�w�_�̌�0_CvƻG�UVM�5��!p:N���?������0���1m}X��F�<UP}X�h�C��I�#/�K�q�8�oz�W���㓨kа��FuN��o�`�XlxVHYEB     400     160=��8q~9Lk��W<��\�5n�cKNO��� ���B��dN�3U���
���]���3��T���Ɯ�����A
S�>�F�HߩĮ��� TK�3�K���^#!�+ݔSƢ�t�F\'V��y\�߼�V&˫��=~x�v�ϝ�5�Gˊ��hc���$|�M�"����,��O?�Д+yQ����E��Ѥ7ͧ𲋮�_��ZB�!^Օ�� &�sv�[}5�߁Q��¸��5�d��̠��sY@	}_'��[V\T����Po2nd�m,���n��H	a�^t*���v��t�V�! ��}�@���_)Lȉq`�E�����V�M~�KXlxVHYEB     400     130Ʀ���2��������#�Z����X7�x��N���m,T�2�A��ř�^%r��z�����yX~t|��M���C�owv�o�s�����b�,�%u|�|��t���^�6���2R8`�Y�Ul�>����$!�A��܇�4q[-�c(��樑>=���ҳޣ���n��Q�(�r��}�L�\��2�軙�������-|���Q�D�ϼ�Y���-qS�t�T�C'6xߑ�[�c��6���q�r�WG�%|KS76�UR�{�4ާ��CN��[.���V[� ���������zXlxVHYEB     400     180�1f�E9:-�iB��m#9o�~����Žt0��8�N�8�ކkqnXF�UJ���[q��d��AFO1���}ظ4�3�G�A���HJm/0sS�88��
Iˎ��4P��I�Y��u���YVǸ�҂�i��b�M��.�\�� }�tO�	h�����(���s%���H�&�e`ΗŴ�*O�-�Ni����¯�`P�No�f.* ���n/k| ������E�~��ʌQnl���QsH~��6�/R"�ޘ?�N4�l�/�jW ���v���o�) ��|5^��r��)�À遑�O���_��@'���#J����U �\���j��%�u	|���;�v�EeP��N=72E������<70��l-}SvXlxVHYEB     400     150h �0��S`��/�������n?9���<
�@�c��OҒ�Yĭ���cxvw��I6�<Ј#�U.OH��`�t_��K�Hh¢��H�
�|�34�1$<��#��<>R�q���q��GNj(�I�M��dTl$��uX��[t�7K3�l�A����G-@�J�2�"��/�H�I�0�v�q#�ظE�% ú�et���ج��~�w���0�+�Ѐ"�M5�b��+�u8�)<�y�����y6X�#�s���8!&sZ���J�]�ܼ��X�(��+�=�����z?�e0&%��X�;	b��;n7�5�����x�XlxVHYEB     400     120!-��xKWp&��7���>�6�	WK�ͩu��c[��&�Q5�8�b̹dqjQ��?��M��"P?�|8S���
�`	$A���s�i<͝���в�`�v���& 2�.&w�T��I�
0�-+>mW:)�p}�����
�}���5��D��ź�GPF��LZ�Q�s��3ۮ�v�:b��bP�QmSMd�`�	�cZ9�p�?���RG���|{xR�!.��e�q?�K=��EG$��Hԍ�(�����P-���aӟ�Z��d��Uv�E���~>��'XlxVHYEB     400     1005�8G�T�Z�����0��V]��K�v�CY|tAW�Sz����z%�]��d�h�`_��Yr0�� I��8��� |r2|�<�!)�M�����y�I��v����#�JY �ѯ+GҼj�%���5�B 2���8�`Ϧ`��2��/4��E��0F��`
�(n5B��tG�8d�	���g$Ԙ��qJ�5���]�C~��]���!~U�_�x�]�*��Fc\�`a�(��/~P��>�XÁL�a���b5-yI��XlxVHYEB     400     1a0�}�T�kJ*�.�Q��y�{$�����y�+h�;�-� Zn*O�{���<�7h$.��W� N%\��^z�S�Bu�N۝N;s��%��ގ�[A�F�>��Ʈq@�����3"�iE�n�@g��ν%f���Ä�\w����C�mE@m�N�C|,{DYr,
��k��w���Ϧ$���E�%K���`1����t}J�B���e��-�K�Ip��}�s�&b�G?d�RC�9�kFؤ��#��p�0�bλ�Af���0ģ2?ϰk`l�̚����+}��{�k.����)���b�$
��@�����)�%½��.�E�ΰ��,5�9��08~;꼵�'�n�V9��m�\�������Q�I$*<�~�������d�4���(��&��5	"K?PQQy���FFYh^$��XlxVHYEB      27      30��x7���.jϏ|�������#2>�y}F3!�{��Bl�q���^�c