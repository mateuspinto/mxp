��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��в�{�����2��͏	�o(>���A��R!���qH+��8�Z$5x��(�;���n�!p�]����e��:�ׄ��Yb��a�gdM�:�Ƚ����)�M<i��vY����fJ~��Z����Ѝ\��1Qr��U?E�r��gA��S>�lY�e�ʳ��P:�gP,!���W?9��KAe#�7�|M�������\/�W���=
%�v��ɿj��0��Wp�d��wbu,S7�nQ]�P��F�
țvՈ�g�*>����X$sP{_����mY�B����}��m�?�'[>%xNwk���ޖeM)���b�R�f>ԓ[��
�Z�\g�p�k���,ˬ��2ӻ;w�92~N�pte�8Kg�N������?Da(&k���<�y�)=�<��>��zE��
;�pa~��o@WKJu}�ds)�_��0-�P*E��j�ݨБ�y��Ȇ����Xr�v��wx�Y��S#�=�c��V.j�4}�^��z�!�c%p_�G���D��<�9�wE�����߰��N��۩�Z�yKϋM�3~g��ݍP�Ԁ�=��Z�����O��#�m&_�r�8v0(<pE=�PV�-(2��u��29�������j#�`y�ߪS�%�b�'<>9����d��	LW��6�&�����Ls�xG=��W�
�@LE�B���~cgӇ�Un۶s&y& �n�8�fR�@8e:t���,@�Y�쵡"S�t. @c�֝~/��@�b�]��<�Y���\g�/Ё�������K�:�5��"7�J!u8�PM�� z)�����^�`��6#ON���Q�O!�M��4�Ju�LaXjs&r��4R�0��	P��ɓ�_�;�|XբM�
s�~�j�	��~	��(�����a�d�6�B����#ҋC'�M<�@0u뤾`�SH�Й8[��t��J\�1Of�~�5� V!����@�>�;6����������_3r���e��Fl&ܴ ���WJ��Bq�eX�l�R�=
Ԁo�O���:)T!(���8.��).<�
��gNA�����PYA��3LY��#��M'��!C@���x��S��I�	�A�Z��sN�:�Y^M˄�8�̦S���4��v��9�~:ج���%Vこ([/ڞ�+\k!�8����R��~��@-ѧ�dO�f[	����t2I����a/�e�I�!�W��Te�5��t�+��ּ�b�g�ky�{��1WH�f��@�����#�cM9�i
�^F)��$N�{��c�K8��Bj����$�@V�ቂN�!�lSE�|�}�)8�T��p�t�K�����*�
�o3����+#��t�[O�Wt(f^W�U��Je���WA���Y�yg2����`�� ��6�S ˔��L��5I#�,i�[KR԰�v���e�P{ɧ��j�if��':4J^�3:`���y�V_KP]��Г��3^�����V�l���1v,�A#��$k�Z2u�O&�)���V��n��p�'e��f3Ps?�4Qi�y{��O�I+@����>��s�i ��qh��_j�7�D�<2=&�)E>б�M�wUĳDFb��0��(�Y�3�)ؕ��s�nV8P��GY�yIx�˖�;��#U�0]*�\����,�T�`��|�^ŗ�����V��-ew�+_S��jF�\�s��D��������8�������B���;*��c.����DZhN����TW;(7ŷf� ��p�MI�������g9�`{�nbd� ��fЉ?�e�G�:��%w<��$1"
�3�`*�e�z;z���Ń����C�^� �h�E�}Om�}��%i�^&��ֺkn�^qſ\[��AXrÐ+���,�*��:|JB���n����e ֽ��kQa�j�-Ƽ����dw1���`+2W����i���(��������uH��Z�b_L4C�B5��()�}9R�Ec��,��N={�ϴ�)����	���\���;u�vjc�[�ފ�����?}[��T+�2ln_�͓�=�KO�c~��)*N�/�����w��ߡ>���G˭A���٨kl�-�8T;�`5SBt4�4;8���[��A�b<�q���P��z�� ��xx�p�iѶ�H ڮ0�o�w�Oe]�y�S��%�ʀ�N�OP�a}'*>�#�S��=����������'XN�iby�4*����w�Z?mju�p4m�),�栢�Ѱɨz.�������a`��wNib䈙q��F� �fRϴ���#��?r�e6�4���N5�!&$^���y�3��yU|��k�k�_���l��;)��2xMڅ�Ց{�($��Z�C��E&�_��{�E\����/ێy�[�b��{v��} Uy8�W1�`u��C%���<��M�'�)�dK�2���={qA����/���9m�H���܃��N�vn��
frVs�;j�J�8��R� ���v�������P�5�)u��6�������d%��\��L�X�f��܆��/A�D�P[�CC	Z�ǀk�g�nn4� l,s��!T:^��ʨ�a�=��#����r�l����?�[!��a0������{�q��r�O��f���{J�����x�� )]�mL�z�j&����ҢS����Q�����2���;]e�m0ꜟ5��9��y��%�@c�q;*)BLâaN���IܘxG���w�W��A`�6����SS0^��y�tu<E�|�T�)Q���?`����(]2�֡�O<Y0�<]:,�s#^�C�@�,4Ж Ll1����ir��L�
B�^AX��VS>E�%�T1�Q���p����l4�_%q0��۔gt �U���o�dM�q��������7 Vҧ��PQ������|�ܿ�-��>@�7_�U�L�X�9TJr9�X�ŏ#4��ץRoc��>�D���.��I��U��6��P���=�¶�n����EK��̋�*p�����_*4�g�0kW %���+��Ĥ��=�A?U?�ž,!������v�6̴)��z!]>	ڎg��� ��x��9w���W��
d�Q��.�8z�D�j�X6�}S���lIJۈi+�LJ� �g\b�>��Oy��i��M���7�<^�OD��b` �Κ��j4����>�i�@��3䯮]o����	.j1IDs��X����W/�4�(�k��o3[7�8ǅ�I4�!��v͸��y�O��k���j񩶵߀�Т ��k]d���e��v�费�2x91�0	͇�����Vm����gIP�h�G?ۘz����~]r���3H��o���]{�hW=��N�<��9�^PH�S�\��z�t*[��'�.���J�k���m<�C���U^7B���4�X �6V��qBB�6q�ARo��PǸ�8�E���r��l]!���A�:8:�1Y:���]D���Sq-'tC��8d��9*2�ޙ���p.z���UT��.�	��+g���h&��zY��`��p5���w���h��]�kO��燆;���j�����m� װR���<
��d����6� 5�BR���=�ϲ�ss���Qm���Wd�Ҳ�w��s�`�?�B��nzq]e}76	6�2�CX���8N%j���U_?���l���,�K���q̑�>2}��s���/UN1���rI�F�x*��r��'��+�����y���
��I[#Ō�"훠��'��gA��I������Q��K�a�dF��zEl��h���,σ��C=}�:\E厵����/�k���N��I���S9w�T�3QT��.�)��e
��l_�}� �+XC׹���L�NX;
�d�e�<�W�\�Ax�����L[5ܧѵ*�����ΒB���$/D���sB�@(&`�!�(m���+I��RK��s��WN�t���Ox��BK�G����S�p�y�����Ġ��Ѿ\Z��,��q�U����I�	Qc����Q�O��uN:F�k��JFiϢ�b�_��O�����5Ib��g>]:�~F�YĶI�`b�'a<�������}P���5/*���  ��ʊK?+���n����� �j���F=4����z�7����:�YY58��l�S����4"�q4�U}�a�נ7���T��E����۰�M�7�^�I����+��s����!:˭�Q�W�T�-�6�E,J�uƙzs4P��W�d���쪞�� �68!�[��J���<��H^�5�<��3��EQy�Z�$�w�ф��#Ů7T��m���ݏ�Ҝ
bK�X�6f�b�uj\7��xY���@��N�w�g�s9��X��gݾ��7��JR����#�Q���vB���Si),X
'���-�5bbH5���<�uu(Ө �^�=$�k���TQ$��p��]���DBQ�DX�#&��h�4��Cr���ea�AH>]ׇ�ȥ��b�f�ɠ�qab�Xq�����m�TU!c�i%��
��g��Z�Ux%+]�QO_� �cc�i�̼q^��"���*��zV�w�Ǜ�
�U�ڲ���q+�К� �c�Ke�b ߉^���>����=�EH��L�B�
�6��J�����3n�!A垡[A9���	���*`��{$K�T���̬�貚bc���b�n�)8���j:�6��1kR$�1�ma�0y�R����P1렭:;�q��/�(0|=|�XD�q$H��"?�ǒ����"�?�^�1k�fr��D���,>
J~#fo�\+�Z�zU��`- �� a��\���5�v�P��x�K���cǜ��4�`�w�-=:�O�8V�p�8��!��� @�m	g��&6ܒh�C��cq��x��PK&@�q�E�K���p�w�.];>���ژ���gm``�Q���\%��T�r��n4�����w���C(���h<ā �$����E�Q��.�\v��������6�r+6<�K�z�q�4 6���bs�����
��rx`y<J���#�d\��LR�#]� n��\���2�^���݃��u� ����wbk$$���>�{ƔV��TXg�:��x�jy�ď-5�:��n��(.��Z��j���jF_�[0�(1����-Ũ��}r<:eC����2������2��'��T�Q��.J��=�ZY�`���X���"?ϝ!��@���V8��XL���0ɣj���P@k�Y�C�YH�^��%V)���&Ǣp��J�����+�4�]�G��zK��=���ݢ�Q�Z�`�p��MЉ��;���5��`/��fD��+T�q�cr|2�EO*Qf��/'�o6�^j*�.f���+<H���n����ӹⶌ!�����j��Zq��5��j��6�!]��0َ��e�q4i�-����_���ih�,���R%�~rCë'*Nr(瀫���0gp����Z!>�D-pr�"��D���b����I��Ѿ  e	M�.��pE��la0CM6Fĩ����DO�a� �`������%�!��A���/j0�<Ț'b5�Į�8����G�C��Io=mg�:����e��Q{��è��PS�F[.ɥ�9�*����4t�nT�lel�q-/������ `h1Rg%o���p���D���m���CU��>g<�bƿ�)V�i��D����UV���l< svyӍ�П�?������*T��]�>���?�`���{����m�nK�췘9e�a{���O!�J��×;k�C��9A�&|3vefH��ݐ]�wv���������5�VK��o�Dމx_4c�1��n\�
Vs���5 vl���?n��s�΀*����O��[	�s��J.�D2p�1���PR֏����~%�e�x��
� ��F�̝SB���W�_v�J��J�t8<�L�9&����k��Y��}ɽ��"Ч�������0C�S�tמ���������#�[�� �%�k��ʯ�N�ڻ��;��HU��6�,�(��6��[~�S��Δ��w2Y͉?�2�&���x;��c�֜��/��tG�
�ż)[0{ ݳ3�s��a͸�T���}�!�Gz���u���I�E��tQ����/�JuЩb�z��4H%篦�RI_u��6���U�H��ׅ�P�в�Q�0f�M�qáF�N���1r��*Vf"1�\.�6ѓa��b}�ƽ�SR�6�[�QH[G5"�zi(e+��,��Ye���?���ܭuنÎm2j�z���ӸM�e(�2x�<ձ�[�ٞ�e��o2���X�<�� �;[���Ӻm^B���L6�a���1-���Z��#�"�}�B=	@���~ȪE�v�A^f\3��4Vb�V,��g:���[��*�L�4d�	:���IQCr\!0���K@3��Z@>���ƴ�K�ݫ���
�d�'�r���uf�5�iQa�LbtUj? N܀�ܕ�x�=�!+� t���Mw.[��Z�X]v���&�(� _�����k�$�l��e�����ƞg�u(+9n���]fOT�Bj>=�%y�{����v����k�r߉NKH�^�t�\���������������K=�+I8Ή������g�����'����xGW'Ч�����>��`�E���5� ����ҴPq����1q�uT�|rqƇ۴���4�	C�+���F����;P�+��gRX�4��-B��.�.ڱ5���^rй�e�Kb����e��ƭDԏ��Nm-x�Q^� KVnh3�� ��cdzT^�%e�b��E,jU���MB)����� l���Χb��O�w�]5�E��_�����)��=,����Cy�S�L�=��]�������l�ɇ�T.�+�כ��NG�Ǯ�/F�1����[������i�ɀ��o�;+���G��I�l���  ��ɒ�~��=��L	H'ZPcaP+�=D�OĊ����'s/L-(U*QI�}==�H)�ZHҗ���,�I�1�����A��R���|���������LAW@9&�r���ǧre��J���c��_��k��?2FDbK�O�.qn�0��H,���^K.\2����:�� ʗ���l�k4��q㲈�I�

o�E��r}�X:Z�[���ai[+/���y�Ӗ��-������� ^t�9@iSrll���Q�c�Ɲ�א��͹@�+����g�ڢH*ed���dLM��bbh�5���-GX�.�sʇ�<��9�~�8�YLr3>1q��a2�ܨ��Y0֏����<�ky]q�1R}��3�@wD��^ֆ�0��{����O	11ƪCH��J��8��-H�����b�����T��_�@q��y;8Wκ��٣b��*����4	'��o8⅚�!�޵���ܓ2a$����ɳ�y�����4�9ڝ�gYI�A��4�����Y���1�ÊnViM���7��J�gn�w��W��}�LxK�I�+�҄;᝱{Y��2@��'M��h5���2�@�y��>֨"�(��G:����Q, �
�εoo*/��<� ��6RcŒ�z���i��c��9�#�1���IGg��6Y�\B���4*V�p)�
ޔz�I6����.���ͮ3�%B�I'S�"�G����#w��e/�U���:���c| �	��y.��[�o�N���Gw�\'2n�Rq����i�K����3�0J�[���)֭��^��2�|ex������.ں ��pԖ׈�N~���)|�f�P�r?�ƿUW �k]e�� v�Š���@������z�9����̎�=��O�[�� F��Z+LK24�� �ce?i�6�	��2�����&�}!��bu�?+�7�ű�Dv��7�߁��`����h�}G�Tj�Nһ��3�<�'�*��f�G$���^]��J2�^����d��XU���Z���6�s��j�BW�A52���)�	�w-zɰ�̚�&Z���(>�� �a���DN��=N��W'��6p0_�?מ_��q^&�%�E@����Ӎbicx�PM�d�,�Z6���6�mY�q�}��zVf����	&Pg������'��3q���1z{���M�S 0��<�5�%C�-�nN�+`�@���M��>F����TMGH@��9��;���J��u�]qΚWZ�Ӥ͞������X�"b;����2g�%G�UA��l~] �$�ܴ�u�D���1ye��!�6߂���=!����d]<�h�Ҡ����Mj�m#�!C��	>����P�UWbeA�7��n�?@% 91r��U(3g�̞Ď��x��W���5�_�u1*nA �6R֒;}��:�-�j<on�
�
uB�H�`�6�o��>T��p���-�K�E���F����H�iY��� �6���]����+�V�aT��l�n����[#2,�y���Uw���N����5�ϯ���Ζ$	Ր��?�9��p���;;u�33�Y3I�:gζiP�X���� W�@���u�o��09�{a���11����p
�`�8&.����3�����ӝ�2w*�G�r8]�q��zXw�.���$>2���h�]I����d�����y���x�+�d���zD��w�^���fz'�	�o�PGR���[%@^w�
�x�B%x��rӰ�
{X�z���u������������X��v8����!�ԍkC�߬r�zs�]����t���od;��+x��;��8�I��
\əHc�;�xL]}��ű~�

����|_ѓ�����ii&韃��mԞ��
H�'dZ�_,�e��:"D��L7!��4/r��ĭ��"�gd5~֗d
�o��2�؟#���u�e��z��_0���Le�qt��b��i��D@Xi���_��]y�VN0�Î�k��=(���[�N�+���=�26B�\����s�X]���#�����q	{��g�H���J����Ų l�0}�����3��J�'����_P=6`H��(�17,��\g|�i���;):���Y�]U▙E���?pXjʰ���|�820Njg��sfP�ye~YU.vu�eGy�0�*����<�*b'C��U:?h��y��n[��;�#�v*=G�����ߤ
25�'I��-i�RN)�?ƶ�/z#���;�k�թ�HzOC�簡s��pΏ�j�<3"1�xo3�@�����	;7KY^`�ISD���V��u/��r�IT��Bʧo����
��6��@Tzw�K`/�֏�##��^6�5����n)�z��k�?�O=�O��m����T|����AB)�i�&�.�BG�݃B��,�\�72�	�����+EA{B?��	�|��(�: �'�=����Q֑t74A(Ow��=:	5Ԋ�z��&�r:ӟ3�Ka�lT�̯M��GO{~>�F��Y�P��\"���ǆt�� U��[m�v� ��V��u��f���XC�ߨ��!���)Q��_W�MR��d?He���(U�:&;��I�R<<�ĐC_���?�C[��� �5̊��;���q�d-A8�ؽ���k���HD���ɴ��*����
 �K��Z��a-�Z� �`�^<W1��jl�KnF8����#��%�v&�ʁ����V�&��u-0B�}Z�WiDg�V��2Z`c���T��JXq։�:��q�x���V�*K�C�����l�-#c��i2,�^:^8���9��)�:�,j����4�lq�UV�����/ꒈ�í�g-i�c/ixGڃ�6�E�L�S��L��p�)�:�H=n�gf���N) �����r���k�f���H�qɛ���s{ i7���3<&<����+�/���ԅ��0�bzMc�����M�e�p-�3d��w�Q�Bp9VW��.���X�0}g�r��j���(�Un�:�x�Cg�m�K!�
�G^l}%�i�M���gi��t��F����x��-� O�w��m�����h��dqz����·��c~<��]�>
�2fN�%'0�c%
�k ��yk�%��S�,C31͒��N�{!�/\����{�7��F۟j_�e*���dW�N���3��:A��W�I�bak�z��zB�&���TAZb�*��4<)��s:w2��(�kV&�r���O��*�M��RúF�*Nt�ǖ��$��Ԧ�b&眏�w�AL�ύ��8��[���i2�����H��$��9�w��D���V?	��o��*��tP�I�IR��/�>�(��K�OR�`C��3y�“�_���R��"���Sm>��L����������]D�H�?����B�*~+�oWl�U%u{��\F���(�&7!��g9}��%��4Wg���i}󞆨����	D?y�I"8��!��E����V�wj͢v]ҷ�gn��2�U���mi=Sq��X�UL!]~��H	t)��3Q�s>!�[�2ߺ�`쏄� #V%��r���"z�Lx��ױo�OI�A�#�s|l�A+��UGkB�c4�~iܥۧ���4�4��\��0�Ģ�R"���/�q9�R/K(�f��S"	�]ӣ>�k|�6&<*�~P�^c-<}��n�䮊�^�|hҞ���; �`���h~O��"� �tY?Kɠ�����"�9�hT�{�j��C�`	_4�CN�K��yہ���C<���Z�OT9�M�K��١���B� ��rY-#��'�~\��n��ƬQ�3��M_RINi6��'��	�:��e<ua��q�c'n2�?T��!I�|b�>��iJ��&� �u"n"i�r���S������)�m�BZpю�FqL�Z���Ý]�����5f��	v5��{c�+	;��-f��'��5ͦ>s�Q%.�R`h���x���jV�5���`1���{p�Y!�Gb��C��.=���Y��PhY_;���#���Rxudf��C���Y���#FO/t���C`��<�(�׈��1Z
�Sr' �w���*3iA:��71�C|2-_�;	)^-'j+��!�$�v�2�,���#x��<uF�8��,���"@�9��t�EO;�4��r�e����Ł7I·�L�X@�F`k$r� ����X�Z&{�&RxEyF�b*^�����1k����t��9�)t��A����ހ硙ф%���V�.9p_w�'Jc�l����M	�v��xےl�9q՗�QR��[�n�e"v���{Ec�#!���+���A�J��r˚��w$w�4�s�z2t�~����6s�%]��N�鱑
4Qg���[���d
�Yq0|��4^8�va��V9b��k[��	��� gh����#�֚����q�;? �&��ޞ<���Hۤ�y=���#3�V��n7�3�T�1�q��۞���VA�ȝ���VmԹ+���t�P�?���n3+�\LGɏW�+#�И����Q�'J_D8Gc�i���H36�G޽{fn�c��G:Q�H� 6����Q���?8�3�֚	�!\��B������:���7c�&�҃���L��&N)����_%��#^���z�k�YC�p�PZ�����	_MPic������5��9�Ex�z�1J<F#�*]y���_���{�໏�vk�p�=��iAt���aO�l㯵|��%�y1�9�`���h�v�3ߡU����}�c�v �J�q�e�/@t!RJ�_�>�鸮X�am�ƴ����L�������p��W$&Ae�/�^������h�K��6��&��q;�ݘ-J&W���M'���B������A���cAR����ͧ?����0���<t�6�D-G����l�`\�� ��	>*��0���gQ8toq�����h�-|�4��P8��#�9�8������Kv�4s�`�,]6�Ru7���=��2��Z�t��d������9��-�t�֍��hʝ1�ؠ�y���[��=Qýa���b�1�kE]U�1qhW�`�QB�ߘ��fT/7��y�#*�\�r�`}!�ʎ���͇aZV�Vlf��5"��3,Z�ٶ�=)��Ֆ�)#��3��Y�:wg�7�b��÷eq2��5�i��O	j���6*R(en���VG��(1q�N�:�Io�����n
��P
,��"�V>�x�.{���W��'4�jױm��G��դ9T!�4�7�mU�<:��z6P�Q���Ҫ��_.w�p7��f��̝=ָc�H_���mvQ�HP����t�����C��Is�)�tN���&O����ӕ�����˥Ql��
�t�nX	��s��T��Ť״K���1�P	��MY��*Ve��kW�@�Y�ǗQ�b
pt�$}�ۀO��JH���T���f��r���@�"\����SJ�L�O0�������(p+-�ư���$��2�n���xh_�ӣ(�'I(YC3P��<�e�Q+V�2��H�޻S"�ܺ�i�5�.�����{.{��u妲�`y����(�zIQ[�L�j��%�[BN��HܽCj<4�x�0&���f����AG�ki� N�~'�!�<�$���0�&���`�Ipן��7���D/�jef@�^�峘��9��٦��^�y�i�� ��n����c;�3��f�r��瘺9�<V� ��h)�k��A܊���i��5��慐=wcGJS.o�q��ΐ�L�Lb�F9m�Ǣf@v���e��骊`ɂ��R|��K�#�#)������)M���9^]�]�1��(Lƺ��$eoũn���p�����o��h���틭6��]��۹���G�u7�5�u�������Y8��9%�]���Q�v�\���7PJ �Q9+��Ň�$ ����rOK�b���'�Y�ʆz���;�j�a��P��7�/#I}l��ǐt�JU/��+�����'1���Y�V�T���؉�9o%1����Ct/�x��)��CUۨ��vO`���
&r5�F�z8~�м��'�͙�iɊ�Y�M~�/k��T���T/�#��|n� E�0�3[�Μq���A_���}������ё�y��A��8�Q`�+9ּ�l�5�M(��PP���uh���� �N��y�@�R�
B�
�vY�>O�gy��Hx�)�cڒ��C����E��2qAtc=b��bb�=���||� �<_Y����1��}��[q�+��N����Yr'��J�A�"���z�[��;�:��t]��>[�����(Sz��e�)_�B,eҖw����nlOp�`���Y k�ϑ���U��V��~�4P�ŀP���W%�w(E�t{�y�!@�س�F������K<�Q^m�����+�!3�bZ"DL_a6�Wߕ�l���E���EN	���D��Loc�����g����	�gUu���=[�!��j�A�ċ��cKe�mG��1�{�"��L���~��E�����c���'8Ӱ Çn���y�����F���ֵfU�ܨ�n�Tm���tA��I��bq�r=b�À�1�skdZc`����-��_�kIy1=XG�Bh�"��}Ћ�,���ã���~vԯ�wݙ^�㷟ҟ��+-4�1�0ت�M�e��I�Nd�>c-�XHh�������%N�&�؀�����,a�d�&����+�"�
�F[
hz��e���l�;�y�L�Δ�I΁%v�J00��
������vyS�%S�ߋW��H�� �ѡ�i0�PNe�-�~-տ*Jڙ̢W�;��
���bLv/��;z*趩a[�d�8-���1�q���Ha[��-&$�C�$Q�L�;��7���	�	lqO)0�䤻!��<��x� �����thّ�~V���q�V��^=�|}sV�2y�H�ǜ��j��Ѕ`��4�[j�����P��7=R�h!.��<�IP��V.sI� �� ~ߠy���+�#|5&=kn��$�2���8��@?a�J� �ڬp�S�PE?=�cAc��0gЯ;�'�hu*��M�-bu4Fk`����GE�`��H��i�
m�I��O�Eܻ�UY��e��+���I���ܸ�*��S�J�*�W'o��ޠ��5�{�* ؕk. �Y~�d+\NfYvj$���fD�p�,^e�O��u]��Y��_�~��K�74��y
�-c��	��"�|^"!ïo��=u�,'=��X�VѪ�7K�����iC��l﮿��1� 0஥��ҋ⃭�)��.A���B�h̴���t�8k�Gj���J�Z�8$،����&p�.�*!	`-���]�ԯq�DL���20�-��<5�c������2�$�TU��܅]�?Y��o޾��r���<v��b��=S�	���gns�z���%�QI2�yt]��6��Iɏ�
F�>����l���A�L̕���+��@�P�r9[_E�C�uY�9��$YV%tB]�7�5#�Ə����Eq���70rN>�'d�����w�f���J�N��Ԋ0�ցK��D���;�26�Q�!�8�4�IX�j1�q�`���,)ހ����d��䄶��w����Sqw�z�eHL$/@�g@㮈G��⻉���m���$�_*�"0Y��V���;9غ��_�tl��sT���A|�_�J�W���v�v
g�;B�[��ﺦ�hNW�j+�I*BDh/��-$���ig-�m��u�$�7�
ǐG�k�����G���Z���r�p��j7l��v%��^��q��}��LR�鉾�5��o��\-���PL��i+���t�� EPИ.1�sI){�B��e"[b�P@6�Ǡ�d��Fμ���!����z3��|V�X�f�o��)���R�4�[ǝ�&)��mx-V�o�`{�ﮧ���!��5H�腭/�V�D��-�.^<SY����Βt��k�翱dt#��活�{f����fwh��UD�אt��W�.�re�����E�
���$�m�[u�
Ɂ�X`t<f��3fo�H�heX��|婫�9ܽ�xBG y%[8a����_\m��;�b�S�:#yN�@�g�d��_����5�z{Y��92=8ƭ���+�6���R	M���%�f��^_�V��}dtYr��o��y�F�K��-Z$� ���!��Cа�G����/j�5?�<���N��B=�y�+B��}�TČ���'��i�b�-�ЮE߻�.�=X�i�����;����T�X۝o��pr���{��a�Q�~�AA�O� �"��[s���x�X��%R˱�t�N��U=�t�`�~7��e�������9��W^��W���D�h��󵼓ㄞ�n�#S9Ǹ��j�\[m�`2UO�R�Ɯ;��;���������w2�r��g��Z���/PkM�L��!H�r~3ZM5���Ur�1�f	%��_�����;�~v9�T33�V��Yu���ƫU��AC��+�Le���.��M�E��E$	L?�s�s\��T�*3���'�%S�I:�f�x����<[ݓ?�d�K끪�u&�A;9:�g<����ek�Gx�5�]�#:]|73�jy��@=�֒����=>O�1��5��=���S�{�'�t�|,:��n���p���L���d	Σ���M8� ��fA���k��W�����k����9�_�]�U�)�D�0��+}A���%"~cJۊRl��~�14���i��@�d#ϕ&�{��聴2��-�J_I8.�le��e��׃�,I�zK�;@H6+��K8Vr��UZ�Ǒq1��'�:"h��`GG\D*r	L0D��
)�!FR�c� �>�+Ɓ���M�C�+Ʒ�s~�%�o���9���N�\t��x����r�p�[d���aJ�� �Io�)���r}-�ӽ�b.$��9�����n/�p?�B�N�,�M��PxAeg��H�Ae��_�ʡ�kB���'h��ܺ�ХZx�`�g,o�	�s}4���u3��B��'�+�o�J�yqA�-�e��A /Ll���X�d�ť�w��W(�+�N�<��%��D�̢:��n��֨$��}i
	���?�b-�gh�'����aZ���｝=��R�E�26�G���P�m�k���{�*
�k5-c�~02�>��������V���o����:�}�ã:���<��҄�4&��h����Ƶ��뇨�to	��B����r�q���p��[<G����g�X���