`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
7zAJYTED5rby88cHdYxwHX/GKPLlsMO1XKnm5mQR1X6El2zEKIWMguwzYYVoT9JzZDpTPUVIlN0h
80bRSzMDJ/cj7vU5Dh/RY70X9b40dxBg8C6V08L6ddUFKOYaWoM+iR4brstH7v5aBZDHa75YcoEf
2pfBFUVR1QU7Z4d+HbSO7cD3IA+PrZiynGvo1C8na4VeylU8roaXLpyxuP0TnOoox1fY3ONyLusI
jtpJWb1r/3XqnzHB6YgWJm4xVGSu1/Blih2nRw+DnbDfkXkEGkfAAYtVLqnL7SumBk8U/hnC7aVx
hJblelWbmOEg1GSVq3WvwlATo/5IFfsDIZodP6FNjy/QGZvHDtGcbIcb8FB8dJrtioJwGp0x32pl
xsyOL2zLWqPmTJNWGn5MNO1qZa40Z3nDLTWVVSNohddnif/6qYl4KoxUCeqepzapx4L2MnoylsSO
i/x2xaznlI6TTJCFWAUMtHxNo2xEMMsHQKfOy5Ua+1qIlXaej39dRdnivNVQQs3rcJ6bj9Gr7epL
FWjHGJ3uf2faCeZQeeHeVnfui/QlJpLGcj3ZdyLLqE/i5pEEuQSFu240HsumvjJ+hiDVLGw1OoUz
yhBDJznzPUXhWuraj8y50YBkg5b7qdsTKpfEGp9EbFWKIv8k4N2i7O6JNmCYoUXiFSggF7C2wB6V
fFjqDydAxw6+5s9ol+W29Am7e0w9r1zud4WUWKIBjWb8RUTYL5MD7lrVbZTj9y7bPChYaXc7h5Ch
OyD6OblJHnWOnZZpgljcHS/RI/X4BG7SGhz1QMQ2/sghIzgxPKJqCjlBALTDIsqrxtOTpPUHQ9v+
CuCQT/+Y8ZK8ew4HttlK7V9VVgfBR0hJvKd2J5wrXozT4abIlhT3fKJ1oInHeD4Hj3LyM+U/lLTN
1yqZS/hmR67PHf8q2e8Ss7lt00H9hHKWkM4iQg/LIGmUfHj2+LqQF7VMaimG6tkDB7PajcRZqnIm
dS2G270ALUQbX+w4u1oX9Lz4VBc7KS6CLC8u9uL7bc28wIrQzZoIN8UUFcQ3P2o6lruAVIlxCovb
V+tQjbOD9IXAvkO9BYFT8Ex7eQerr73vWgN6fx5WSUYxm6NHBQwEIONRgaZ6LD+UhQlY+WVocASz
XdsgPG76MjFnWEgwlyLJHrKEyh/Aql3oV+VuXAhwRnids6Nmid6fr5Jvvcm2+em6LhWHpfE7gDAZ
gmNZnmZTZX/HijUk8n/dk6EMCDwCMqdLzfq9M1bDQjruBkyOl+GnXmT6z7a9kX7yOLSycs0C6/1L
VnKiSHDTT59bd3PtNuLJU4HZq8o9J7vYctO/dSt3ezT5Nv67R8cLDZNNN3wKSeZ7oDgAbmu6gCB7
rJxLRdYhlmKRrud9H+/NktYe/0W9SoVvoLgbPUs9tbIVBHxJvySoHZKZR6o0SBJELG7XdM7XSMGG
S3CWe5HyeJ4QNEVBcvZW7rYOJPSymtOQ+u2jSERO1iJO5LhdBj9W/AUsy7Q1IlLCTQqM9uEGDnvB
OovgarcFGLn2htxScyslHCGiFRBCmadZU6M6UefcpK1FxuVdZswrlRNR+b0ka2bVUxfnGM+Md0rN
b3Y94ON7hgMIY5k4MIn/w6A1+VQKDRK8fjCutdA0Mc0qQdkU60IpkIpSg8BQW1IBlvASxLzMErfL
jkYbWxcPQFHeaFJTpPWwZFdczAIO4Vd6/vagZpnKyeP+F46hVbZOLd+w0qlfcBIb1DSuVG+TA1X9
3f/Rsred7OCCRPhBoeWfWkYIQNMtsLyqRYpdvDTxlTBWONRkyR/Yy0cEZxoz+4n7tReQiEXM1tUO
greaGz919BHLmfWylcNcygtEWw1jochSpWd2guMLThmQw8jFHHbPryFKPqhw/WS7NbahJuwMOeZN
pqnuHvRARyRaMzQdCeOUdo5a/OOHOsZ7bLUewemphFU7My/VpSTKnb6JBJnvDPRKblUPPMXQ6v9L
K1ktVrlVvPxa6L0C7xm6rH4c7FrGUhBqylO2iRDk4yDaLADPLe6fiYkwj5Nnb/dRrae80iyPnNHd
RuByUuTSOtQGFsh8pZzCV4wuRnV1c/uJOdtqLHPg8qoSUR0FR55myzZcQeQ5en35C5yx8qQkPqCp
m7oM2YWsUbMnI7hGfcruu6wSTOqBuZjzTF0i/ZKxA/5bmIuoeZQy5GakNnmYgLwZsWwdS1oEC91t
zmgoNIJRakGblgYPM6tHEHReuxbIxePQ5gnJozeR0Tg4tuSMs4Kv2COZSCoOLeWTsJ0ntqiBCeEt
H50ZJKYp9EYcM6c1ChMMSFs/vKk+HWy4dAOzqeHEtlO2o17gz9wW7EiSeco7ZmeqXoIEMcmr2heP
E/Ri+Jm7PPMs6+sjVhZ23UErDiIIHPBTPK86nFwiI3cfN7olDUYXhJ/dBsIZpMAjSot2pT4UYeA4
LSFIxrcBUffteLT4Qa6Z0AYXa2Nv1IAcf408xDZAN3I+VoH+A33u0qhIe2FE++1pgDBgnmk+fjGP
PCc1C5DHbAvWqUw2BY+v77E68ezR7M2N/g0FU8LPUfGR3olYDCoJiYazNtcXw/0xbXvJgVKaAYKS
eZsb+N+DwnHnuTBmrgtmIvUH89Wxy6r5QKvFyhGtHJb66xWytBLG/kdc1EZedncu2DYpUFddEbQ1
ngUzFuVq7ajFLxcv9qlCDmiHlLn9mqDzR+7CWg4gZwJK3ity3WgNbcvjK76+ccb6wZRZOLs1kmjd
bN7MsR/rFJgNBC+SOSdByFUJ1hRbROXOZwOlDzJrlsWWZmYujvDKWgSAJlU6A9RbEBoUfQYQ3xfc
tAeamkx+Gq6nc9NiPE1aq2jytg/kevXEdHgQmwJ1al1wxqx5Fm8hd6Ocr9lQGSFWxpad8xAiwxo/
8J69eE6ytBXaH363ood1pdmyXiFLtpC0gz5u4DixOCFYTEydlZhAOFtCGbVJd7j9XRJpy89ndGXt
FTV5agn15fZK/IOezkaNmfmfUN77E3qtv/qs0HWbUyb0H2BMNDFo56eSi0n87gU/MFlb6MGZrsaX
rJhikKXCbHg77d8sUnV0To6xQKim1oh/laZ/fUQHFUbcRGsEQ4biLhgJ6duRoSXyFocWqR2PWmOu
/CfC3VSgMeFOBmf+DCMEwBO9GLfQWZjCDC3JrG9h3LCcxVi4ivkuEkton5TfUsT82Dlyc/XwIHqs
NuxcDv/PBz0lN4qBnDkiykiG9PEOq3Pz1TfNwnxiqhy81Kov5UsvdGdUifGYMY3IwMvJivhzziNl
is/DPTeiHqJWaixeg2+oNR0j34ABQtTdOsGOCz4p+WxBiyilz32aTSwp2gnqF3SbL7ycyUxnbHkz
Pg1SpkupOFhoM11sqjosuadtEVcCLGCUpu9kzdgRH7gkfD2cJNCH7rDa7zfCX1rYTV3FVfTT2l1S
0uBWZe5LrDfR8uRhyU00wzDrmGldaHXw0S8uVpKwtk4HAjFQgmm3NBss/spxySJ0ukPPgUQI27W5
bqTC+BzQ5+Bxeh50WB5OaX2UMHB0f+QjHKO1lBSlApUTQtbjQ2/B0fPp/1XwqkqnJDnAgOrwhNkv
G55p+k2Zc+ISTgMef2koCjOlvN62GaRglmTp4I/7qMgNLGAol2irgw2/ebPiWZMFkqUREQcvPgPp
RUl3g72kkq5blmclxK+xW/8ruPNIfgRaxDpovAEhs9+EqcyPl494zNw7T4f9H7yfV1TWoDLjZ5L0
xegkcKhKOwZue9+Ptv2ra43luFrnx23CWmlmplhRZwWzwNZDiq6C26WvKNe3ReMtCOaC+rDCrXJN
j4MguLnBqukdV4yMJ7uxoe/Ah9wW5LZl+rt0yFvJ8yWMcYDZOior4mfYHw+v5u4BGIVBlxBqPqF3
5djfy14NWVvsuxpoPKfTIuhbEKVTtf7g15+7oTEVmcRBtbM2Hiy/lX/hsxzLQqmm7jefHTINYHoR
vBIZoqJSUw71LH5TT8m3CvcHsq4nW2KXXciru93L7Dtk1UnqXXB6pTIA2Tk1Nh/HCaO1wAAG1vs4
p+NPJeCIWtywhBnruvXS6G8kefTl6MbTAuPEx9/k96VjI9ts7c47rgLAGJISfMgmERC5xavaDeEt
pqY9DA203qkwSJgFiKbq6GDUk5aXoKxr6YSSBh3T/S99m7TIwo4+qI3wT6a5Z6gxtReHbKTzcaSD
4Q4IIwhiGlxMdu2N81SvyITmmB3uYgWSAMVgVCF9WjUQT3dAE6txx+tFBSEm7+T5Hj1QsNFT6ZmW
JQ1WDIgZrl83xtyz965vLK+HZTor2ULxH34IZBgjTF0NAarueRuJru7EvDa7OjTyOy3qzSBNLxAW
FcmTWPnG1dRU6vVtwFK6EkaquIqQcRQW4dkyUTKUyuIXoGJPux1oG2RcH5Vj5Os9MZXE3/9iWTFO
5su7UqK4+8fewta4i3YhJFZswI/c3c+MwYxhVmeI3UMb7aATRweJeXki7YJV5NAPbGG6chLS3whK
2/qP6qLI2mVXNjpt0eu8F4LM/4L6lg1QjLAkXp1oBqPv6FKnuZryok780jWLvTNx+X00zHcIx0kQ
8vdsGM2A9YijBbcfUuRnEa8fEAx062XpzDwUYJenxCEDVoszsSQ94aNnRy4z5ObMn8vkmXjnn3mD
mtR3tVsXhkX/FFndxBemZ6JYH50R1hFzEcVW4uRPA9hrBu0VW7JJt++ynm/M1hH0llTU0+JcZxx9
U41jjQT/dzy1Rcuxt7GH8RABTsBU9INmOSxkYlcCfynvcQRXTJrDwz13BPE3v6kwHpDwykRymrOj
UGRCVvYTFAzoR/1n1mxjVJTYgf9UPE+Dftu1nXcidNhTGSMg25pwjERJ0lu3QzK6jWFykEThia0C
OEPKXHY+0yl1qQPFh3WfCWCgZpZYUU6cusk3Ly+5ToOTLwKx8Q2yQsQiXoZdNuzhli70GXlfp/O2
GdrBG6Wd5OtTrsX/qlM4J1aIA+O7FuR2cMSVs/xkzxZaf/3sFvplv4+B86U/5yWuGec/p2psv13h
tH3PjBM9zORoD372al04JRK0cgKAWnS4igDASeXLQjkcg6kgone/v0oSiT4cCjAIyUyNKjmihodI
EEtNMMRC3sxI7f7psDyDkN69+P8+j/V39GhejIiXLE5VC0CEfchdirE4CftKKctGBd9TP8HU83wA
PWBEFqs4Fqcbe7If4ty7J7cASconYPuRV4bUaJBrsiqv5SK+RZ2SZQe1Gi7E6/Pz5myu4ezd438y
ij8+mgJfdSy+FPhKoki6PJswzCMBFTwOj1JcrEUj4aQP705pjGW6OAsznSrnOc6FYgIi8QTb4Oef
UHMn0lebUSkoZbRZhUzyuXzon3xFNA0U12c3URyfOhq4VkGV3gcOF6aU0NLjOm/DZ0asfvh6CWOX
AX9GfXBCMs00izkFZnveW5ZopY9I0rsfBeGaNacMILgi/nhRo/noRxSK6SjgFjk37Ke1T1meoijB
hnRWrcpoZGM2yFk9MQEtykSklcmWOCaPsyhAdxTfZCcfPe7ZFvCLW2nODYwZtju+kNaqCAJGv/EN
9nINO8Hr5NtnMCr0ONOYE8CJr6Q7rS2MG7kVyx5Js2nuY1FNExDRxSKDG48jToFPtM/A0gKVEz3W
vjMUbLOnU9iNa3Gi87+qql8yVK1+myyX+xSg0zJLdN4uhPg8AzS6O+huNIWXg0Ps5DW3b6DC54Ri
lKEMKSORYuB/pPrAlA0VcxXXA7mBPBjUGcy0YExp3JJlvqzwpaUX9nIhxot82EnIj2ouR5mHPjiS
S59xLSVZgteRssRo1d5Z9WYjSJI1+Lm0TuqFnyN/5Iy42AHYl1vICFqTfqPk0Xgqj5C0zWjz0BDY
JI5ibNfJbBL64CLBhtAQYTUtkdv/lDN95lHZD8kgj84CSuerpYiRhnu2J4/FFvkHNj1wh8PTGjMr
3IcOZZ4XuV09ijm5x4Zhbw8EzNM6DRsaonllXICwDzWhjqv2LsH5QCRk9/apM5wu8DSCID/b8s9Z
P1AHdGeN18LCloRV/7vwh/oaj1P/piXyyvSC2LbiOA+szHKp4xdtuZaTXi3HPKG0ny2juTI6UEX5
PsXCgIu1DpbuS11My9kaoi6ktYBYbHAlM00SFmo3T+u9WDBEIyrwrdAp7sSyLopqzAiEwT1aZ3YI
eLCtmZt0Ccw4Qqe5KdEDnu7nYObkipQdEc/Q1lODbknI1KQaVVHoEcufdQDfQc2X/oXme2jCF3dL
Cqv24kJv7i4o3WnymEQppNxxV6oPCtrEOAtYzjwwPyxhHGpojItAiLqJ+LnHttpTzTz3SdyrL1t9
BcdSkc5cWVwHFdVTxyzcMtNfQXbaMs/IZFfhPZwRiFfeLIrBBUff5oN9kjaLcIBhswYheyAvfULS
hrnK97BnrxLuT+CoLNU9itaMfgpNE0ng0STpNh8I/YiduZ3W8Q5bTnjgfiR8CwuAQYUkWfBOZ5g9
5FCNakInWBQ9b4sI7RNwp9+pQQdX5vJRdWXADTJpTXwKSB/wHe9Q5YJcgp5vfDMPdEo7YyfbfltO
6uZuosBoLhqXs1yQxM+KMXLaISPqFTN0qlFCJdRGglJkEaGVf5ya0HITzOiYtH+SIZjlq4m4D4Ft
hsGPSMY4b7FX8FJZHxfSa6H8O0ASb/+5QYLgzf28oOkblBMKV9Be9db/K8oA9fWLzeUo/SaLSU/G
j0vXCftYV1hR1RcvjoT/Gxc6Y8RW3r6oaE2mKMfXetKPjznLW3heAL7fguNCcKn0JwBiWIoiLO9v
5lHxVY+25zkDqob2irWY6J5EMqXuFUW5LIwJiA7v5BvDZpzu04LimfFRBsXy/Qiy6GWus93DZwHo
33E2tKQiuJ4nIiU88gmHtenU6yrGGaoBPCWmCeIFANwOeMrBfOyHfPcu/xKgWwFNonWuKaAINqV2
kXfg1Ilq8/G7IL0WebF/KoPgGT5EsUBvGZxzLFS64K7hFAI5uv0TIonz6HBjsc5L6Aw010vnCPcL
zmBs/x8A5/pOyvJqbmD+bYLcLeQgUAbVNP9jCVgPLolk0+d8hY5Un1kbo/X+xIKGenG/pvnuMDC2
TIeuNVMBwVHpIOt/aStTecWEUAQPiuoKUlUOarzgJuYs3qOTipNAd+2L5ou07rRtHvbHhMzNeGlR
cU+BU+An1PlhIBH0vB9Bted+ex4vV74yKkyrJFx3afzPN5Y+QnX4jlolUEHcnvNHOyZrdWXmOOZ5
yvsNoZL7GclNs9yw0WgYWOGfA1gUOdD5aQ8NhtBuYDQUaWaJo9JxUohwSrvcidL6aC/tyJpRxdrt
ySRyRQbuKAEwBg1trPXifi/eApaNqcWeKWV/u00soIZAzpn16b2+i+aTlbvHzue9y8J1fW2bT97j
LDGtGx+gkYOgGN5qgnhgtznMp4+eN8njbWFFvuiQ7Vj7kZiV9gz9ze0J2uoPcU8vN6jxSfI/eauQ
KJDgzAYylLQtF9Va2aeFmKtwAEJ1tELYqfExri7kPwUuVdhtFItCiDV9TM/3GBqLlMTQDsZeG/To
D1dqBj7j6IHVaQIGcv14wtYmTyRvF4GMZzwQwUy8wN2hyNfpbJb/NPwZ9A1saaIrs5XEEi5+Dt2L
NuJ+d0wqwS0qFQf9otvtvYxpt7z/n1D8nWBreWuJcrkik6JpwFz8EwvszVLygGjk0XPt2LqXvCFx
36Wy+gldMDQxg3RrAnfQ5XbBznSblWq4ipqjoIVCngNcBFhi0D6ePro/fXunx0KSH7djvHuisEWl
TV4CbSgXhIEaBjGqESPpH/eHD+8V2IMvBjprrR2Mhkd3SJIiUUCCs0nqr98CqfkrOaBxr9ihiG6b
Cp2LP4sb+dUN2f739s3195CcQOAOqW86Ha/+QS7xbNGOGLgOX9HmmjnXLfIX0bawlhcAUf0sBiEt
scXfr4+303+vGHuaPkhxNqrQjhJvDIm1c71/0XnDlZbpJijZa7Q/zIAUjiYUc44l5vrNRpAHYB3s
jmJEqwKnTX8jve88B8uix4njHEovGmiQEELQEGx5fMZlSL0h0R1dYGSSjuKZeIB0vVHq+MnYeNeZ
QQ4FXpW9HVLOV+jiBjGiwnmIeJVrBnDXbHm4FfA9Zl3nITKirTStviyI1z6t12HU9jk6u1DwEGxA
qClHJpfLe05/oSU7hwB6NkmnIl5NDzH7vRL7myP3WSjI/mpXX7pZe0BOx1gWnLvnK7QTRbV9R5/r
BD6zrXLwI9nvgpIBnK1/kFyx6ILmQr7rvv6aMwDrVFXX24k5LFHFijkDteffRBTvkoaWmEz5W2bP
t35YSKUVOqiil7u/A7gswcctTHH/5EmNKQaIf3Kt5uEav0IP/jgLAwo/Ytacny2/a3nMLGXFiuFu
t/Jr3TP5tXCpJMDZXBvhLgDC1LNhzwL7OG/v4HdFG9ELU6Fwl23WkbtgCts7cDoYhqBWwdKd1uA0
OIz3Eo+QkEzP4jPU7OTdhyzQ0vnu/wH1W6UA2y3jGgutRUGWdipMA24/9ZFoErvNIs1qdszQ3IrR
cAVCPyuWApoq7k/P9LttEKuYcEF59DR8M5xhCIA/niWjmXYOmOUNlKTzsYyGShI7sm0VVLTo5ubQ
bnUHrTSG15nbNDF1CVF6YCCZnf3ZOBzwFicaiq163n8QiKvlYNcP9Ccf2X2q1pFvZyQai0vp3ce+
h4V4+zB4a8BGpCz4SCR9h+qfPruMcKNY2LPU2KTBLcF5L26FhcI1oOguZN7cMK3vbFGZUUfP1nxj
/sCy2+ZEW++wJ84zEv44I/ItieJ2VYkzvmQ7fLwPI8FXsbv95IV7x8z8tajdcADQqIqKdRiC+yCU
v6lSsFLLnW16agQkREAkbXY0pK0u7zqSF1hb27GZdMqHnLjPrboh8W6y/ijLCCpd1IvOtVq10cVY
mx+MZ3Wd2iBQQrphMKUo/Ez43zQmqBpnVLgupSgPqXIgsIhqgIGxxtZINs72ESxYXhUCgXhnZOe0
mddvB4pArvfIUxzwqZ+8+9LkIWvnhVoV4+Pp4l1Jg+58Ssp6eNhSxYF3i6aISXd2qXYranmY+Gff
4uJ2ow1UXnkmGexmAMx25iB6wEcw6O6M4d9AhTtYJUESGPte+C4dOGytkPxuWjRbi+Jt6q+XpXPf
i9Uqivqpwg4RwbKLgJr7fTgzbcrekoYCnP/rn5z2YmCP93lGH8zwjyopRLLiuH7J0MMQt4slqswW
UPWohJ7do9LZ/Q+8sxs6cTfdDTVEZHDhvfMymvqh9x69VmCFBmmMSNBT76FJTrJSAMUs4OSom2iQ
Lvx4R987i0abYbikwglCNYDW8+0zW51xeL392V9RkaV9vEGckA4wbPji7yrrC8ttZS5KobL+v0do
E1ziotB49gRygak6auZv0VKte6bagcKJxPgwGUC0hweXsFSKKnCJmlV8MkMpmIu6nfWjSDuBBf2T
Xu9AdtB7hmbH9gVM/0J0BEDM6HJiWL+OTePrJEkQm5KkmhQcwuCussT/0mlj1kIZpMn420wj6M+v
ejrt90FiI8qcQBQYW32NIG0+HrJt6NHLJIJqzE3TiFk+8SgIKKknmpW1pisqyOWlpKoAOrLXOAcH
a/BkOj7kfEfJk4BrzhzdUZ34g33+60Q/k5kqjOxTCs9q3g23nWLN3oQn/2vsLUc1VqeejQOuNOdr
9mQadigseXE3W7iQGT7WN5Fk8gMk3972UW4AViMgKdpKBpr/Ky+r1IXjvxhxG+fVfvshQ4o9f0tA
7+AytDUqseRdsNUWsPmia1Y8GQZpykD9j6p+rPJ03oKQW8CgJImvegzjhy1MWtFaOEKc+bLDAZZu
kqIeUlPrIDZsnupZJto7+s8R8TCoq8UDmc49jwLKYEVSHYU4leTyyosdxkVwlC2DrED02TuBnXg6
aUkiVXtjMGjJSm/HZ00gxvNQJQR0jqXF2O9s5ekm394xzg58srOv+yOw7/bAq7BqZXG7vL8MW18A
InjonqVylrjjz5J8+vQHnWL8B8hfUdOMJAMbpVEly3ds6jM0mor6gVr7FtN4wpXOsWCVv3zrqxIT
gSkrgY0TgVYLuj4e/h1HqysQkqIvhEO1GhHOUUVoA0xSb/1sJFAqpO9hLF+jbw93GZSuJra1lO+i
1q2WtJnJ70QaiZvsKZra8R7bWmDx7GfTj07hpjw0n/cuw2g170oIC81XQD5jpJ4IVdxG39c13YhO
t/B28FAPcqiOEW6h9xkQWkeHrH3eSnlr4Qi2y3VLsh2xNJSc7VQAEwlwDo+hq7hC46x6yPbmmkVc
qLMg4Sgbmtg+p5r/XjYYslivj/K60p743Dh/zF9Je+Z/WWwUOBASPnNAcDscBCDgbV1AlJKOAl9c
YIVwP+6VnjdAlaBG4zBSKmrl9yBQkQqoxvtyLMQ9ajz3PcgNHXm/f4Rk8ouEpbXtJcfrNObRKvS8
ClDmlhq7Mv5K71WKO4oRxbrmEQzT3azxSCzIL8lS4igECWqmdco+1LOP2bTC/l+pf1pWgZK3Ysqz
LEl8DwY2szATN6XiTkrnd/G/rOAoLEP6IrAPq+nqLoXHLmsDwW/avhVGvNpNt+ZppMSZ6oTHlMqi
ditGHrePY1jqlCFzuWZPcxIQ/RrJOv2CX2t9+zr/k5vdczz419+vwnayCpbrQBeTnlyuOJmjjbBU
sWR04Nmv83ibas4zmxEnrwlCHHtrK2uafDfzE1AWK3WxDBwct+5OSIfSOTurxsApZfbhA1B/zJOo
eTlfYd6BH7Ccjlv4j3ziK5zu+1OraaIcfKs8571YE2oNF0howzeJSGvuXLMxfRJdQ/CMD0PR5r17
RNjSKmeB4fS1QZIUebAqfa+lpcHliFEW7/Zw9g3ztywzP4VOd7qL9S0V/FAKYhgZJH/bP9Dnw3VW
OA335bB0HSBBA9PUpsMV50vHHLni8oZu2oJjLV9LiVNwYeancgzgW5exuS+ggykHoKK7OtL0kuFb
ncjYO2ak025k6r6+gr/cWoj9jG7TwCyC50+Sr9U61OFXCneQAAaCkwuRpgaSUpyx+hVYxnmmEy7+
Y4/FXA9YC6C8zMSaoQpXi626n08etNS7hFC3uCjSYhheI+li2kP5RaAvt/SMAQAvjBfJoWK6Bdd6
u1kV66ELNzSx12mxhz00IPwhb9DeB95jCOSBMDgpD+UgHAT45vlze+Y5qVronC9TExiqbzn+h7gY
ik276CCJkUik4Dv5YSBvJEJnA/pYfIdPtgv3EUSPkdmrH8L71I+Ec1kDZfonwgSdxjg6D4GYvm8o
nv38vHqJLPsnRfImH2MHS1wAyoRycQj3xTnwXRHX/mDrOt2TLUgKEi1C4ghGZrumCn9779FixJvu
qRFv6XT5yGoqn1shu/9r9raMT7rKjmjQnCRux9CWFyGolv5IWwRSG1C96NtKtapIaCWE6vkhgOC5
ftxJnvd8QwB6Um0RzMe+GVY8kvUGSm2Xamgn8zA9OK7u91WPEq4iOW7HUaAmwllXH+jz95hlbTm+
kzzf9yPIXOAaU+UPndiTyr+1z7oAExcHD09uRZA7ZZ0Dju3cOGKG0CEbf2lMBUCzDn5xTz982lo8
uG3kQC5JWHrHaM3mrxc/yUeWtDCOqDOnhkHwhs4YbgZUNWnLnobRYvrw1sOBQT955okJCosXsdwo
dNku6qprugBhEUZUjP+5QDBQSK2RTgxlpi2kZKXLLgO+EetY94HgCGy3bgfCf636mNYY3wUJamxx
CHv99JIgOC24b25yJ5lW+f6MDdyUFppPDz+cXlGKHWHMFEdYk1ubbXiD7R3cvN/kxzdjYiAp+0H+
aslI3/P5yGMLvv2QMDD+h6oSqhtRKc1wOvb+PUaD8tlruZTXx6P0LT39CYOvqwVwgUiP4oRmVt4p
Apm+nxmnCL1+HxAqHIvI2L8/wXGxKDCYQHBocadi3T0LNe455SLjLFK5Jt7hPq01uEtr8BuGMXm7
sgrrPdFOI5eNzz37TMsLItQpKHDeKrl8mazzgbopAW1cRsTJdDfC/+uiEnw0ttsDXwPvI7kvhVmk
OzOGUjLmpKuMF/svYIn3sTuDJwfV6tYXu1w2Z+egbrpK5+maPvsOK5op9fBd/oWb/xNSI79rtTI/
uK0It0oiUOKH5K5nCdH384vWBGHIDbeHyI9aN0ZxY0X9UqYpHG78VyA4sDJOGOpSzFcbFlkpszbs
9JOJwLwI9TF4Xw/u6eXG9/PDC/pBU4snO82S62VZLsCxfACoNOds7VEMRDOr47d+M5Hu2g0AERnN
5FXHEmHJLWv4C92VoWt/uyWXuWfqRCMaMtUM4iv7aA6/c2jE+meKLahHUbXCsaboUJMQvCSWLRZf
ZVVExof6zzmF5NDgKZXmlNGZfxVniPxjwA+pXWsd19upr0D90uWm/cxpE2fx4bSDp3Zpk9IdMrxT
XrxeuZcBKUBrEIdPWMHx0o0dWgFU37FEiJKY11NyqfOGf6rH9g73Gpe3nuR89l8rOVjLgRBGMajA
H0TA0pkitjy6MNM5RIZEVy7d9zsfMlKjZowMswk1YsCzS4P28WsMmLBY7V3t9nS+gNw+pIkknu5u
hdGRR7CnjhhMB+SM6Gll6zVHmkz6AAn+8bAzOHvGpAstiIw6QEx9OQK0WCsa+jo+5kxCvDsifTM3
9d0a1Fpzpbp9/Yk9/3HUFwmiodXxO5ye3hQkAzfYWoBG42eVr/rVSlY5ZBqzZYpVikQFDLulSrgh
ZimmMdj7hsJx7hUNPk8PrHClGjCvbXtKbLH80ba+mGpRWVXdVjLeJyIfR5eWKJVPhUEOlaVKosJv
5NHP7Fk/X6gpSbpznO1t5vouizhxg5Bh3PmTwc7vZIQP19hQzflRvLMt2Q3Su8G/wmpdUCC1WiiG
pogw6aGmHKlQCihjQYricka4CwK2XfrJPnJ8khJ6W3Yeg60pAEcRhQ8GpeqFgotlJ2+3lvcQRBoO
nMjgLlcPnvgGrcFB6vt3/izhVBdgdoyvT3n3MCjI5Nk/fRJU4o/Nq0zTZbjaDT8aEGLSxKEdDMy/
RLnfPadfGCSQZjov/g511+m2VXzvAWz3UvcLkpzTkxU6uLhUkf+ilRTFN4ufqTdQpUr7v5dLAJEs
MocwdybuR6rOa0Si8CwINXajcbldLw5Zt/DnLBRO4UpZF8F/tT7B2ECvKd+jS+mEHJW/ES1iUiFK
pIqMdb8W3I347atPidTK69TpEXCy8Od2DUUk3KCI4SPmUcj7py+KLT/Uyz1kM64Bzxrnuvun7dNG
JsH82t3f4SH3g0EuOWNyLfSj6Cnc2CK8RGWpWJRPVEKgRJxIawMa6FNv1xZVz+XRzFQyC55OCWEr
81Z13YjuQzP8/5QIybiYTtThYFE+0+LCH0GBYCA+AEOP30D97uOMDDtcwRwaHRcrJZuEGspBxzJ0
W7ndTzyWPKwZt7JjqZJkTE3ga9RtMrl8h7MblW4k/3him18ytdNB97V7xrqOdYgsnxUk72WLQPmA
AaRwdv/eleWkYoe7vfjhFQDGZ0iA3wQEuVA95a0TfNEQJU5ho1w9oB/+yht0IuIn8Ltz2aNIeEZV
9aBkFtSYtBNxysBhfiKWO7yGdrYovm4dRIX1CH47/zo7gQ5RuuMTwmBj2nBjd6lwZKZVXYLhyt6R
KdIPAa24BSgXk4H9Da2W2mYR49utahOErP4+gGrYN6UcpQVqkrfDiFSJR0LhkeCXBXgMx9NSlx3z
DhTy5iVUO+QQLq4/Bk8Y70YCq/FxdJYU91f29QurAIF/agnialCZ7r5W06U34xCeY8RczOdzOzBx
kqzbxOSBQE9ZNmxChN+qrAcpbNILlZgzwSYWmEtt+HW5XoYi/vTq4fMY8977tHgjScTly1Z0NRvR
jxVGiFB7N4Y37DcYeyHCS5geTxGtnKrd+gZLX12IdWjAzUFO8XZMSvXWRurG47PEb/uYhQiYWQqk
CvDmf8rmIOGSRgsOMYpZUdq9PvyTvvsQi13ZdbQl2V2gnbOMk5u96WjGJxLOGmjTMkmzSCXbnWUa
+75Q1QTn+dSVnw/M2bW08dz9DQ7sb0bHYROQRfKdO2HYiFDmfk2Lx9CtdAJfQJgGJlCHn3yNCVCi
FRMmdPhi/LEUD9OxJE07U4oNWhgrk9Jaqj6Q7T7PUXLJtZstk2oeNmeQr0tTg/FaP2Xezh0TKD3L
mh0VGfqMMfm+vQsj3MPKFSi74ggOuu1Bb42d298fS//RDUI+SkMgiV63BScHkKYBfd2bPWtMP9/y
tLvxZ2HPeaBDzYu5ttd92PhGVrLSZylzkApQ/fFICxev2xtvie62ABCXzPriLPwH89/VaSqSjLUE
/13lVf4LHAr3KZI5F7NnxYKQZGAlpJoeBP66N4wVO2Algbd6WY6Fkneb+YAHH29zg7LaQATeeKPC
m7Fo8+Y6Q7zXNK7QS4JPYTTVbsmTbRyoT6Sz4rrsnh3WIc1tqRWwytJepAyZI7faA2EyT2EN4/qa
FN8W8lSZm1rWky2TQmdmRPRUQkLjFiVrVCssS1fN6l33trDMc/L1vaKAZhBoz4G1iqij4YfPW5YO
t7IyjM28YV1W1NSu421h6pSAO4yoYSaVjXAtugGy8z9MqQLSfcHuM5w2mYk+sUcmVi9+tjfNS3J8
L0b8bb9TC3Ea8t6QxfX1kiHFAGXwCOR0J2dfdA9Fokksh0bgVfTn/brPdSlxYqC1nBf71zItzU/1
YbROh122dfgdPHlffvwEkBFGGZtV1Lcnaed7f1viac7+5oBgPXlF/kB3NbWk1hbZDNeqF4B3rqL6
z44lsBer9ABG/Ccp1Idk6dD7GuFFlvLxjzrg1buVpCdotmSoB2p9O9+KqE7gYJ5rUu5hPbznUrpW
EopVplkmSic+ii2U+IPtT1GZEV4UKhXhNBQh8DnoaxkFos4Ly7NVyRQmbQqoXN3y2palmltvdKq0
uYN5714mjfOz363GYWQ3bjoF8nKTdVJqxguw/c1s+fFh/SQOLKhV0xZx1I+9OUM0MnoP19Qc21m2
MAuSRKyLj6NqPrxN9p5vJFZQh4m1nvlW/IJafLzM+AvFBhAb4LI7QfzlKsT5m9KCpEsr1SqteBfC
hdBCr0rZXHwtNW3JeVV0CqkMUHTG4/wfWNuv7SQ0jfSTm0/Leuwo3JWb7MKwcfoF+v56OnS8fbTV
YmqJroobal6VGwwg1bKnagrn79lXCMGbtHUu/f2mQTpvwYR0ujqDU+35XJ2jbkPJTGKcH7FVb0W8
CHSaJ7zSnvV4nF5v0Dma7qHNvSAMwh8qf6qfWZ+DnbjRvN4fZzk2fw+KQVThT2wSlTRQQUv0UCU3
xPS89RpILgJCLqntd9DYJmA+35ZRfgkL3RdOqu36jyHaCioxsDqO1vlKQYBTl4w41waznGmKe2tm
o2cRDes+ie4zOYDHu1LkMRpKggJLU/01/xw6kXZGf5nlaWMyWu17zSUEFSSdMDFT9CUNtMhstla7
Lkbe1Ym8czDdX4q9lf4pgek7cUrY9P9Bw0AnCnknAUFI3hgQQjAQTKy/fP3YDNJkM1wPz7wFEWBw
pkvpoUwB2uM2qHLYhTLgX5dPP5Wdwfopz22NHuegbjiGNb9BOSTF9MPhWDmmp3NuzBWlauOQL1iS
CswEzua0AhOYarXK18XaHvzbUcCPiYIiXQziLT7FtUxOAz5rF31a22y40FhaSoA+lZxlwtz4QNuV
lXlZpi+/V1+BY4M4/5g10nAAdFbn6b8tP6J/pwQXpbLf1oB/ujXPyfaeqi2jOYRNElnxZ2EUZNj0
Ez8cl/q1RsTrfoO8VV/4N4W/osRwJF1QsVHIcdBAuluPLHBOaDvuqDMbIk20+EjRV2FXVUEjekGi
M27SvFTBFtHypoVR7+593mxf6KpJKnMNt+rXI280mG7Dh9n2h3SvuQROX9bM5LS9g+4SVq9EUXvQ
G+OZPYhYkv7qVCkTjPpBtcA0LcptEtwsyUgK+RuQu6+fpILSwX/hWI3yLTR4CNE/fGP4Hr2570YD
Aa0pKrBf3ECu6F9LB0MRXJFLljsVOi2UvtYCpqQMwuwG52IW6DWz4LQNTYZA11jGF4mYjKnGY6cQ
wQOdNyFBBt7CGhzWgo7JyS+KGnu50T1uc128r/buVEaVm+gZ/Uhj2AWfuiesVNT1pfgrLpss4kUV
Yvz1L7g+h6VgYXSZC4Q4EWDfKTM677lT5pxdKgecWaooh7dFNWqdApXbanalHOsuzs5Jm6S3lcXg
eY8z5dDVnDvy9HCb9vcwCtNRibxICgEUpXuNcPGAqR0LVcmB2IlQUahJCpVRQh9X8RT7kM8Pk292
8a/GptRz7YyojV3+4d3ZCS2mDNZEOy/yEJs02bzJt0d4KnGm1p78pQ9JxidwczShLUNOE6UW0NZl
zqL2SAmwwcPRJgQdVvHuaLx/mEFB4+xFLPF1NP5TScgfGW0a3Wsic4FwceZSb4cmskInnjOGyERw
FlH75OIO7K/Vrr/SFoArdXnr52e3LaSf3YKuL3n6/PHauuunKJhPAzULDXEtQYtQrPjLsQK87Twa
bnUba31DfotSJSbAdzpOm9myNN2xAdETSIA+7JU0HyoBjbDeMq3ZBDen0DcIdjKVRkPKsepPpn+K
Ghyiv67y7TLeawXjW5eJLTqEtHW2/RrVYv7NaTq+fpf18yF3ZPzUz3jNlhiL/dC7A7i/JHMMcXXl
Qfu54qMNdotGSH+Ejh3mJUaFhmHnq7uaegg7c4Ol65aVIasm6pwAs1O/r/Mp0Y38/Iv8U40/PWsa
aKCgTv6dt7MzQ8KCpIzwbrUEL1cPcq4iPFkBpTBASfeqQCfZb6QdmbvVLi+OJmWYFGjnKegK9+1r
xe2eYiqKj2MxEsg6sfoqbKDEhwoe67Bp+59NVfvey7OCAXmiYyXwILlcCTCHB+tAXGrmw+U75zkQ
zKpcEohsUlEEcna13HsbqwtZQbYsDZ3QnGCymoeyWSVYfIjHIsrusgcM+DWpz84KAg5qhMNGDMQ8
tZozC6bo+vT9Fe7K2kmHs2Q20BmFg579MctzWr6qV7vHuM8JE+SG6ObdNgi4OhrfP3gpyflP2Unl
hkjKe7R/O1yvngo4nKfStNoaiCtNx2zAS+08pd9KzQZgFkAwfU7L9RFG+gI/bml9TLRsfxev7XAG
3qYqU0U9ORvrknsp7SDHseMdZORTa8OCnmAaGU9i/8CUbg1bZCfnPstVCINiTaz1/zF52KUeWcrC
K3Bc3+LEQg49lh3in3m0Nfd5GJvomzVrBm8ekB2pbZuIfGtkCktRQI9d2/se8O6DpFjCf1bpJR7t
ztdQEhrKXpCgBC3Mju9HHPNLHB/HTMgTsKzvl1ALmZBym7m2kzHsPPS6EyL+c1xM+Jo7959Rfl2N
+7iVB8je/JubZJvfgvNxiJfevfGmr8hEZhR4Fa2HnJaYiAwYOVsMQxRm4GoCCKPBK7bZFzc3vc0w
/3djDQUCwyfq0KN4C5YOq6sKBb/y5d7+6VkjWgtYzkp6WJ1iBQ/xsIdyZ53vfU/KKqzal9HIJ8Au
lFRSkevfZtiY+SJnCS/zntkg82iuyID8CrIxIcCiWxvpVn2Ab1zb6cRgZ+EddcI0GP7XT422a4wi
DNdKpDI2GERg1ZiWuE+P/Oo4S91wcw9kGgtpXhnybTJXPmFj/mQw25YUKv2V7a96AS2oQgOElpPX
P2n1oJxJ7LrBpDxgoOLC0SR0Je7Xog6N21WjxmwSyXMCemU4ucTAuy/0IKETWLMpyDLKjJ9buY+v
l+yhu5iWTXxk8mDWBzO8njse5wuPPj4J0cFutpaPyuueuKZ7MENdWZtIe8DXVcC5o+YRa4b2lq21
FI/i1OdX9se31fCgyes0XDHI/fhPD7CkB8C1N0dT87ZTd/w+R9mbpOiIXOqhu88twqhbH3fk6mV2
8SMwcpqNl63fTxjYG1xNtrd59VZNrUZN0M6LTV0edSBBDeEWDjWo/ipT0NZrsRDIltnrgHdpLwqF
VH1zRW+RItFa8qJic9KD1rl099Kjioak2bqPPQd02m1zdUJGAhncXUhbe+sXDKtdbmzZP9EF7Z4T
jtsiJeZmj9VIbnOoSwfU47IPW7IdwasF5ELyaRkmNljXPrJTiouZ+nEOlVKw6EhxgxBcdS3bCG2f
ymLON6Ep66/tkLyLqpXrQoHp3txxuFs9S7LkBJDn7BnEI17xBAlnJyX/5veMGMDtQHfDQHZIfWrr
EDG9R1JhOJD8S1s735U2boIjL4oFy32Wv9rk9aEenknlS21XwwFFNjxMjLJhaAEbCo024BgDjwRu
ibVmR6fryar4Ii17pAIxUOEihMbnvnuw2a/q8uwBevnDWIIyVNO0rjVtyaQ7Aww6hovZPiDDatIl
g3VUXFHzo7b46WRJLO1UOP4CWDNi2yju18AuvFRs+RLa6VZcpIn63ikB6ha8gt6OZXs/yex02bk3
toZWO3IZFUBuXK67+W9VxFtHpf0ribIIZitJqXxMSUFHNi50CKE73oPEbLxCji1DcTcuuiRaP3de
TWCr6qFvs9yQfX0zLinzrcXs5jOU/aZCBg8qkeSqbUmVbZ9n95GWizBiKEFFu/yd0w4R0XWQfo2r
z8oU7GnkvO0uTPphiXCwgIsYdLr94p4QqD39sX0C08W4+MCNE4XmzFolgY5+ckCN2F3YOFtT/8kB
tZNTFAfiJjIo3l5fYA2QA2iCvDghL+q9/UiDre7sOfCgdamGZ2oKdc7inIaOhK2MMJOGhliP4GO0
d5LG8zdvX8Ik30v7EwTrH1JP0J73j8TUKV73gHLIDbxrwSM/bCr/1ZCUejFpuJpB1wEQK1JxiWPZ
Xs6c1Xrlurm+Veom/fNgxdwJvJEImyPvSVszDgpDyoXn3j7tbOpNgjr8Vt52HCEs6V1fBschRJtD
ACtAji1/+sWsMIZmjiR9Obz1+v3VEvT4AJ8P9EMd8s3m+4c6mngJC1wSf13AhS1IN0Lk4Dil1C/T
aNLPeMFwqzbBSBTFJvWrRNzUrFB3XkpOejoqR4rlOTPuV9iCIHczgTG+qsgcq7xrOjefSEVcmHgI
uSopM/g0Hu8Jw1HsX/4q6hLIiIWyAq8b/GEJvXRZjwouKsURhf4TCM2gJh81cAqLD4XAbZoqgEvk
fgl7+y9BfA2iaOenFKkkC1ie1VOQlrGiRmbXaL7TCmeHNOJhM/qLl+MChXwbdwaGNahvxUrJ9h4y
vv/TEaxEPhUa8NzoJjl1oqPJU8pf+aT68XbqxSFdzIuczOFq8f/mV/5s4q1+LRPaCOW2ONhl4U38
6/9DdFAsGtbcWyovbT9XlUdhwav9Igzdi82W4uaBRhf5s19ZEyvaY+3+0Uh/1xj8dxMfDhxDL4A+
UJg36rFoAH/2/duQ99Eychq4QZ5TFQ8lF/fb7ul3iEDPsASV0Np31v+rNLr2bOMfHhXfcKpT6bw+
dc4dn4uP2/MWUvPRgt4tOMQCICuUbQSjrywKfyfKX68AO6DuWERrsC4Eg03Aj0Z18Y48h4UrVvqR
65K2P6Hri4jqyPiqF/tfAh1n2prhnqZ3h1Jp5lVM5ugOsHTGmF/J2gMQ3EHgxtKRFPa0m2GQecPj
l5pB/6CoQqGPTGo3MLhr5j2vxhwmuikX6FmbgAqw5XSOAGBfUgVdu+kNcLOABJSPsgL8k/UrKcpp
VMaJxKzJmbyXM8RJ6UXD5oNuMZXObE5uKaLlfu5cUx5c+UwyHChD1/MIOpo//BDTSJHpyrh3xwhp
rdI3e/1lmBEGLsIDL3J3YDuparctvSEVh7ClB/eONbdxpv9HIJJakpW8WjjC+WMj+8ztXepe4yZp
bFir0rlxZFniloLcHBWHlpVxKDNtTk7EduJYX4ZAvR0zfU2zXst5a/OSlkSvgjla2tXYBbBAY2vw
yZuHxC3i4DsWUeKMgAf05pWvBinLWGsskCXhNFMRmEmf17dp0OGbsCAZfXruw+x+Gh7iEUiVOC2g
Ekld7CgF23lmnoD05V+WLrwQx+19Df1qAspqHrvCW/JwytAhoz1xDWEVshlb01CTgevqGpb9xSK0
h3vo79slXxCAkomLXC8hiw8iO3VDwRAEBW0PIRCeBcwLcmiqZtxOgIWN+6tNI9wAzhsIEttJVizx
5JBfrl6u3vG2l/WzL5EnhGxI/Ey5vDfn48Z410b39dyjsWm6vvqwVR0C7TS87aWM8de5sGNA2MZF
3Tcn5viFpG8+N6EeqlVD4mNbbYF8Z50rnWkI79r5c6EET2seed7YDpLAe/BDA2xxmi6aVQ9XIeiP
+5g9KQjhSucpPf76LTByNVNvw1+XbLq/Tu619qawWzSPxuz0kr8B0YVBG8/7i1KLn+VAhu+5kCBl
czdmAm605L4oJVIOz9JwLdjnMIunWTloXZTdXwo8YkRICb7S6I++IfstOW9i5tiTTDXT/7CLE7+v
5qP3fwQ5MRRGdNj0vXFUUrYXkZvJDxNP2+ci5jhzfRF6jFGqn8bhxB0fcKMC/UFfnalFozZiUx5d
ULtZyaYF2vb8DzU5F5Bk/EkQCvpAsfVWGI4pw5ZXhg2VjI+/tHGZL1qh/tu0kYbA4Fq+14vHJ7sG
Ai7ngR8A5Mq4xp3fGFZJUGtUy3kFBO65gwgb5OObVonX6fTZWCPc5j0fW8xqsrrtK6zQ4AnISD7C
UPWBJLavDaZbqToN3SAwmcGVKak8Y2tABRILbClQy5lKqmjWrjkNaoYMpJF8tnfSVMGONgv2N23K
SfHvH52nHkTjNwBjTtU4J6BHpPQQt9aW1euzBYXxy3wXInzPqrzMJONPggT7C37kPCI807+jdpxm
VvpVOiFAUaeBHl6UEELsQMGkxmOEN65aXFw6QN/4J5vSA18wddpSKadEzxwR8nVG86qdPUR1yaDi
prGuP5MsekxBBz5pHlH9Zj1dAozaaZ6qw9S1mkSK2B3XJF4NAWbju+r7qet0X7L2mjc8yhR1aXlj
m7a1ugORaW0XUuoComq4jMeiGPFO+G3xmF5Sc/ySzpTKXdePS+1rKpdQt987IH7K/rwwnw66Vy2t
hanQRfvZlEecLMxxySjgwgNBwpcHxWI/VkuggdX+9q8D6WQaHxEouJcWZw/Ay4UtThGL8AvUH6SD
sgFWgLYNlzDGZdS9WiXTJupFCsAXppZKCfxZjcepxohrP1ZTJKs/CR1fjdKXdnAjoAI3UuiZjxOS
qJRhxcw0NEnuBWfi4BcDExo03qnq1b6al3xoZqxQfAL3K2NY+r1MY38oIKnLvyTNmuzV01sd3LQJ
uwLmojSPzLf4yBWQVGi9Hpl1MhDyoahaZcfig/R8C3CWcAUCQIwhgHwjNtQNgqVdlUOud4p9EoyC
0UnR5r8KG1FB/uJblld9AZtICLCe3ymTO3QdJLoLegTyruSSZ8f+h+dO+vwILMy+R/Fvo+E+ekJx
99lNJQ6BciveamCzeW79PGK98KIjYYFNLuHowVxVKTlKolzcUN6b5/FgGyVxSqbJLh3RZv+7uXA0
TgZSvPjumyXBWstS98iQOWx6WdRftiUblyNJKib9SgwQybH741gbfVWOtNt/+KJ281hcQa/Bkm0n
fhBLb18ranF3eriv6a5OhD4jCZxLz+vbZpUjJgYvmeNDzy3akn8W8DOkPIMWgCX9BBy9vKuzseng
cG/cKTRPM3lxDMRo5Gl4VZ0b9kX6pSHUshCnhVGQaAUBCMdy3wBVAx2+9HRYVvtQZG21qCMnvbY8
h1G9eJe1Inm/ImkwwG1qFKt1zbA9nvMgha8L4/EOtn9it/VAOxZOpjV9XkvdPfN6ualOeYNkA/kZ
X+gwidFb9k+RrsDuyotTL1EWr8f8IJARvAhOp3hbQh8qGkE9556k0ZNUYG2qslcH4/vsD/3jmBiY
+TEphc45QfVQpEVejlUymOb92C3McxZ3Rj4fzYl2jvoic0FRwILNr13jHw0UvNWsPDnVnWoPjm7o
S8FAq1cRG3ucxMB2a97miyblbWbIdcsddoJbB7his80nWvP1BvnSk+PltBjtIcb1YnbDWuzMaPIk
wBNPr/HfUpEabuGRkKq++Gx9UEka2bpfy0NL02ZMSpDmJLuvvSW3V7nXyUAn+E5jwR2hs26mx4FZ
D00Ih2m/ZJDLkyoQgeshemiygIUCA2xduoHqE24lRUqBL/tAgClxU9YGksarn4aLEn/ZIQEk1390
QFSjSQ3avKCqjMu4qpNHgAp/KoHtNwNcnnyixZM/6jnIxJUbmBRBTBUjuV5FtWbCw4nY3w4ccgGD
VW9FiiOWIezYMyYVnTUCRCJnT1glrq469sFHkpBqMMZgcO0knOY3BCnbnDfKnbKbcTfFulX64HDx
4hPlzTvHXrRoYruH3Bl3imZvEu/CJ6h4IsOGHeODZqYRDJtWxvyDsUrr0K5mTgtmUpiimP6hN4vF
dsEY0Ak/Sj4AsQZ8omogpR3a520rD7BlgnzKjJH+9dbIgwA4btDMgerjUNsyRo+nzV02SayVABFW
v9PEJq3L96OwfIz+x47hZBjwGhnbdjV/6YRr0QytMe+VuCx8hTfqbezXgNEPsNWQnsfdSQZrrJg9
KzEDfYszISqypaVz+Z1eNNP87UdjjOHn+OaKtygkQlSpSGuTXa7ZcIvVfi8c6D8BouLNfviDmO4A
fpvmLSbd7fiiRZRbOhiY+AL/wnAxu7Gu3Tr93tUmZ+OVz5W5zfBhA9UtkjhP6bD4uyDhpDPe/VvF
wPveZD2isxlJZZA0YjOV+n4PoBHIZTLn2eO/1sd+CRFLQchEyEiRi3RL+6G/23JTtst34htC4fME
4kFyAxmvojUJ9cqeVSfQEzwnEibnsrA8IWnsP9/1QR6uX3+fUdC9pCQpetMbLmfg5/754Je/13Ws
SU3JePEpxwWIH6c5uuGisHJsBSr3DQAfhL8Yguy4IVHZm7NU9DDswCnC2gFix5NlpsyhmlO4ez4X
AqrKrLT1DAb3EpAKfHok+BEXiea8B+yJ8n87j/TWNmEfZ8Nx57hC/nmDxkgVeJ3PzX/xr9/4KMFm
u2e4WoNw1zeqaMclTv5sYIh/2ZUnKrV7raoBDJw55n+p3UxKR2Xq/btN2MYkbxMj02pmyG+1AmGb
NKgDSZpar/hQmVO6jI9NdmD0zS8aXA6BWxaB+Xefl3uZu4I+DQlOrpHYqjsy5+I7JGNRHdwb2lDg
mXLY347hPShQ6DmtSYKlj0ZiGHBky8MFJqSFqzb2/K9YeX4Np3nmZIzy7cPU8FLiLB+Xd5Ey+CTN
AA16zOAuT/kXD91a69jT076+x2hQ++Km3sNbDPJjsoWI7tnDUVEa45Lrm2RZDdGvhZ8F7izKdKLq
/UhN5OqMRZmylTBzkgl8QFwVAsSnc3y9nomdoza4eEncdVzhEqLjrYT+QAGjNfgJXIplXWTFoVGO
n6eVmdb2Htzz4iz70wgOhU0KfggPTzWpDHN148AJm3RVpNuoeBvxa5BxLG0fqfrmqhx4y4rYR6D0
iM2Q3nm6/6QLHczHTsY3TtsPidXxM2gip9uVKXJFKf+Mr4n/HpHTwOxzFlYfglQBY446vvbjSh+W
pF7Ik9ESH7LstVOEcl3HAslV9idyB5Wz6bkuHRnjN1s6mue/du4QHbW7ThaGH6M9b4kGUpgwsIr5
QOymDwUGXMCro/vyPQpe3QvsXUXoBpGcymJYRjazPv9lek76itZ3AIGhkR9wv3T40ohWNkQAiJcy
frdqRsgBdoR/WpWECEv31Ij99QxuTcBvnhP/4U8+M6HpcDDSaNdVuKWlU4tL8+KhJ2RF5Bx8P1Jl
Cu7+8WreeB+9RDvZhTZgD3petg3iAjHn8gVMw7Gub5Gqz0Q3mjUNKDpU2yJ6uXkOp1XLHY/dhhjv
Sw2iPHCsleqT52QTtbufA+sOloJZzWW0e3ffAG4APrV+yFcdIWuPTHZpSxT6+41Z+JzKobXAjtGP
mK2KstSIFmOLUScbXSq0bH25Un3zit9Mg4HSwC8QfwJezekPr3E2AQ0qfOkZwhzBAC3NdpqlIhVf
2FioWLobcquneSVpDgeY/o6mUNYXWmv4BhxGv9rGkLdOsSonBjBdcP88PMWFcKN7T5gwIr/FFWla
NztQhbtXf0/sH2H0G1w/zB9Ne6PemM8Th6ez6X0gk4XvZ1/3U/QnMNEHy7TtBb/oCwipURtHL/kW
F9PfdFIhc7VM6AVRO8rg+3CABrCJYjdQa+M2K6EV2sb6BboWL4zGlWbRxk5txhtMCZuz4U0898h/
DZjH5WfWV+qohQImuPwtEI1fn8azq0VjinpTZZMR8SAmA1TSZnWZhoS+VkFnJ4VHa4nZPwslDhVE
FU9RjKZKAZpV6H9RRpIEQJlBtizVJL7YA0srfipJpBNPtiDgTnLkO5GpHc8gnGqpEJDw64Cwuda8
RWPbdKZ/u3ZssQvt77lAIHkyiM4mQeKwdluvo/D/JR9OXhZkNh6euH0BBxUz5JMvaTA17XnVjQ5d
QrP/bGa6pFCXbZuBKwpOqPWKsXzrNYNQA3TSOzg4ST6ykLmTFONUzqe+Ncf0mYeDke1mplUrWA3u
RTf/Bnz3bdVE85UTpBGRTxyz/G1VQdPc704jG5MY+ygbK4ueJFDImQGQ6/JYfF49A5SpvCXaDRU/
Zy9VkYE3u8xepedNxeHmvUX+AndWXNhJIge2v84rX0VnSBttCZzpQOhHlWKLEDv8pPoENBkBGDUm
0TpLwF/UUG/S1uUOblJcj8TbJP4dBWgxOCRAtNyLJtjLQVgh++NYcuSeA4ePrHke505BP0iv4Cyx
oYiWc0+79z7qk7zFDTrppd1zO8UqLlg1GV1qda2c/GSkLKqedpiIL+fFOidogLRHsVZDv7e0Qs4j
n2wLCghAjhi2nm7fHvgsA5Kl4mhyNi4f1dYG56vxJDc3krmy/tm/Ph/6den0w8CDW4x3NivMqxwP
0AtNYA80z78gdPwEv3QSGFi4sh47lHmTyhVh/bpgNHolCuO6RHOTGb/PWWbnWWpX0IcYbaNwNVFE
iQ8UrDmQK2U38iWaSG1lHAdTTZXdhcN5eDIPpnUp7NzcRgX1MAWV98IhgEn50AY1kpsyE036BJ1q
r+rhpnkTioHtUydmSLThAZFcelC+SLinmgbCdMt584ha3gaT4DI1y9r6ehKNWAscEX4gzQwgWfyy
0eybMPusM1oKlkY+Du6U5qbye/KHmd6uvfdB+85mtBGb5CHYZImjoQ7BeHetfbCCR1U5IKksDCJj
tKOe70mQF4El9ameZ1bL5LcDwiTVyvCM4aucNKfGm+nABakLILxG8GPVX/mZ3HYN4qtLu6GA9XpJ
gfXPZ7qC4QqC3ohIV2ByfRkoEpmoERvRA6havM6UV4RCCIkf5lKQymTgCSFLBm3hArwBq/Wng6fn
TrTkiqVz7xNNTErwESQxolPKvDtx5rIDqIdn0uB8TaZ59kVkvu2MvlKZF26m71717jd7oR/muewN
r3B5A1WQpFFK4gXgU3oZpaqvCzO7TE26c/fHQb0KLAKyi7Ofm2E4I3mVZuiCFesDsu3ZqhaZ768V
fm0ntimrv3+Pao1pF1GEhYO64f3qEv3HCcGRRcWxCqezTGgKTH8Q1/C4a4kwINR/4Ny+2f6nFoPW
98M/l0CEl8liNcrzbFgmgiK7KFXCzBMkheTxSzU0AQp4esU3Q9TvNIu9UCop02vTL1sV7Zo8/dKL
PhUAVgNkTRUEHDOGTpm0KnP+CGGmXV9SLqCGW0TV8l6DnvedqEzdbtDBOtwFtNhbmNtNVb1ybksl
G3V5IlKcPxfensRorPMm1YIKCb77/OpJQCM670zCKHUs4//u6FAtaaPK8oquv3qu+bIYUPCxjI/J
UOkpBgqbsKF24BFPZYwbgL4MKw+CNnNL26tk7ppzNTw7uQv7h8A6V4RFY9Iximo5vB9vBPtSOtfN
0q3w9VzSq0Hx+5Hc3hrHjKXqIq1JOCOo/+ynlVOdEc3rHpIFVC1hB87x0MAHEDLJ4Z+BaKOyNfws
a+xw/IlJKglhLbJPKV0Ynun71Wu/bARaM1YJ9bUHdgLV8UJjztKl9mZBqToyQNSogOYIOCICkBHz
jAkoMlOTt+JaStjkDgUUoe3bLTc4y5fQzmQigjzxM3dmwhluOdxUWLGKv0GU6iaSbEo+AHcECwjX
JoazmuhrFiZr8+afmc+FMlr6Ah6GRDPVj+7DPnXRq700omPAsRgd1r6THzVFhJgXuSG0OEnCTYzb
O8toMUAXx0/TqrK7UTqFvTCs/MkGwO2xtwOgeYdK7hPZRP/wWqrF8PKzE3Ivo/PPIiHrCzCf3qWA
8t2y+iGnW6vOg7oN6+9R6eEgSeifO+xzsj9iV5sHaQ6Ij5zK/Qcf6AMqdVJUVayDjBeYd2dXULSb
VurSaPmkNMlgdf65nAHwFREbeJ1Bx+nbK+5O302drrQaBU4wPIVGJem+1XId/dZZWD/LaIU5hlmY
DVmiKMpZhhdfHeS/DL7iqBTuRBF6BARot19jlb85/BrZQTvhGW7D8MmphLc/g+DCOOFkdXbA/lDz
QHckHrKtbysasRkwagqX0hJWjF1bSzJWmTQsSSdjkohW0AyP+eNCqMfzV4yVkeLKbyyGdVYYUKaa
xiWxUuhZSSsV83b2dXSwPtfaZDom2nIQ4GTeCJi2y79FAx1TnyqAAhN16N3WAXq5wC2dnNrIEUGe
xOU5dwBsdINtxKbjTtRpcW3Zf6DHp/j2Ynqo2pJ0FdA1kW/rPnIcv9YvLcDOcDoo/FrMid2ZSSIC
7VZ0X1sVnEyK5WtNvIyefIuW+5V9KidtQ6tS+L19yiL/w3NttH70AtSXH9/EAhv2/hFAHzl/zljf
OZkzURegtSDAxrnRz/S2KpEfKvoO4bnvQ1eJQx2dLWbojgv+v6I/7LGvYaDFLA9BZP1BnfyYmeXb
IkwOyo6dAraN3n7/yWorgQ4sQ/uT5LcICJbvKJCfljX+Wqwx49qp2JtfwDgyjxNR41gTTTTQMkso
7FsQuNxtQhTbZ+QmE5CzYxlcv3fkCYO/uKD+p/MVs7K+C9Hh72PmKmrpKqV9+RTxlzlqSXDzB84D
PXvcMMmuQK/TVVn9vJrv+awPrHJ+EzFGFLDngNdxDvLXDCahwaWAwT2J1uwC+zsIW5HoomStLXBO
2yDKGfBzDbnyd9UVFinvSCO/l5RwIgN5mLnNLSgEXa7KuI+oPQBZLMRGaOMk1Xd5EiIUY8lVyxoB
/EIqP0Xqof6biWpDnGQhquYb5Sux+1rt2/MPasEolb/OSnYNLJ9G4lywivXR5GgcbbP5WQJK7cRK
LlLbUXK5Ao4b56hnUWDaD6/S4cvSEXU8WTNnCOiIcdmMoOM/MHVC0rYOeVnq7RN0YVopTpfGadkR
GIRhgROW0TlvQPhXt9VwMLSdEiCRJSKXJjHXpw4Egz4sTYlctiTOc/Uj6at6grqUtHYj/VygEAIs
Du2MjzXDgKVr8EeIghnLuy74Cog7V7w+rWEjF3JzvkOv8ZifoJSuo+TzGy/kEKSF0dLq5k90DeJ8
ssOr0nlD0kOplhAPD0ZWJyCZB0OLjcHu+Xv+w/27lYt+JCajOkxAo8lDGPbCDXsoFujWa4zop9Dw
e2PnxIqVMhuHrdTyOf5XuJ+LoOTy24oDcpl+vjMal1QzjaAxljJd6/bvW31a05otGyPwv6MLl72i
p5R61Ab0jKpPFO+WnJ43LxDgvMtBE/9rSrL49YW+QpfeHtUdVmX5MzFyUr+OrMPOhfjwpVKHxKZw
rS7yjVxCNn2o/HIUisO9z0hczhXWc2GbcPDIkv8dOjIcsEjHuRrnq05GeANL2b40pU09nsEKPWyk
BCzts6YJTIs1ZWHq4T9gRwbs+ygtu/V5/dLwhZ74Mj/7f01pdNGZSPb2ImK3ume87JVpr8SXdb6Y
Jddr0i58v2M+u1oCCFJ1UIi4VWWMlJt+LQGAQ1YjYfgtwaOvYPE/sHmFG6f2hzMIJMJOByQxGbZH
e0ea4yHAwMR0omZVp93l0Dlz+OyOl5tjrQlh3UfCj17QR6Fj61FPitGm4yp0uVW+x24LWWFk20Kz
ahPHV7T4W9Okhulc30A8kYf3d6NaMttZIZAT/bRZAxEjVyVZDZT4EVgBIyEx+1Vpq54OUFSe7cYF
eJVtKbqdG26xMnfg6ImsJCTcWOfiSH5s2N9WSbYET6RtLOc7zZ5Q1/Me2ZZzMcIEHzXKerJA3DvX
ItRiZSogJ8R2Td+2oLy7EIwCx+NFrJ3T8Z3Rs+Q1dV0E+Yt0ltVgkFxZ+me6F+LlUCRsq8L9rE9U
Pw0pzA6xN+SVaaDa088TrnYbi4jd7CC7/eQUiI4X4qluuy3QWpNTwfu/C3BM06tNdGS0tDYnqprb
O2ZWvJmjA6YeU7fLA+cEGOrFDHViblnnUePlj+PUGN7xxPaveIcmmWEdOlTNXqgKupCOTBJRTBXw
IAG5mtRvuQi3K7Z75a6n+x/BwJCkNW4Nregc15VF2mB06uICrvNzNx7g8uNghijK9XkiXVx8++uz
omhB2qi6h+kW2yxVP7o0y8Md+sRqZOIsWMSVlFubdeh5WwKDn+uDtvz/R6TY07EtiSRMvzYul4In
vco+cwhkRJVGVVg+3tQ15VPPu2k+GWTiqyyvk67ebqOendS1ZjFaG68ZvdYeHWxR9PNQHkGE7Ufz
HnLVHOLkK8w7MX/NqPDtfwkkHDKojIngfcK9qo/TIWBi7Ynx9LF8PuTh7j0oF5xcLUkCfDI/Ipsy
uW+S/kmmLCMWxYEdKZJQ0MDT8M2eeeblWC1nl/KEtakoRUJWepxWi5m3LKL5XPATJBs4l30A5VuZ
pwSwxFbzfemTHZyK0dsdZLZd+iJ+MU2qnNJG0oABCJiHDrypeK7970mVhfwq42djkWy9cumlMuSj
pIfXVJfjl7CbPgCKaxLr7TURhi7AVauQi3wQwmjEyz+PoacMFxUCSx5hCCxJpEFpwVVLhHf7b7iF
CJxpgtgRWyO/SgNou/WXdALl5H7+WY7zj5A8GQCJf17Iq5Q4oNPIkY6YbQFUD8P3LSOanHBt2sjC
ceV9R7uZFeEyis8g/MyC+D5yIsHJucyuzy747fBgeH6LQ486gL9xvUxkV3YGc2invqiC5WWIn5da
TaSzzKmL7EHF5YDTIM9eaTKnnSLlYu6811tGSnV3gttaTNM5qzqo1gbWAhmdJnckd3FDVZESVxmP
XEvlsYqu8w5/UIgoh5bxFrYJk+rRLMdUuGphcUBfVNXFb7cy4I+tv33idIWtSuLBM3JzX2uyK6/z
MauKKxndp7d7s9sAXBY1OOip+u6u5mjXEFVbbqKuRSsNoG0LxO9IbOQ4uGqpZONqz06MDFjWO0yU
6AaCYN3gSNCmjVB3aUFlhwhDlzxtHTVtJ1glWjHu01u45FEKFx6rASVEFNSKXaZ1XlZn98DGj0wj
qg6N6OCFL/rY7756rO33AONsy4+MQJKEj7JpryjHlnXdw3z7GrhJXNw6CpVIFQOPiQ/5RhRuKzOH
dn7v9IrDONtI+/lNLmJY5BM9MqwHm5+0oYnSP1qkqA8OnUvrzqZI9PXPCezLiAzpGfhaKSOEokH1
+SyHHV7ndFh6JduLCNMfQT2re9VnaYwbvy9+lXjlbInYZcTjNQHt35EvTPncAURCMPsfAMOOuEjT
EjUmr8D4rpSz6wIldV0bhlLw9dwbMIWM7KRcPl/2OITUBKb2VwQAeEQ2ES41vlNEqLsRqeP+k7Xs
emgKaEHB28eF1neA48laJXdCbdeHP8MrhY5V8ssxd9Xu27Ku2ZCFldCBllrcnZuAL5625S5jfMd+
1lIbdt0GGjohmPCf1BxxYUCJGJ/vw/f7BYxgJ95g9XhYGQsDQNp4f3JuszDmzYENgSf/6A1N7cOj
B+o9wDfOhf/mK9SMBKS/TZFfcayUcIOZzJ/0VWoiP1p2R9T/SSd7vp8Qo+THNmr4ZAv0YumDQquY
WWrPSq2nN/ZOyBGb3q1CJtOjs9kqfhykOhAiwZmhlKJxKDc4JYAMvb0pigyx8ba0Mlts7K9DM151
vIQ0nBE9c85wQkqSXI3shVvRKAziUQ1rDZUzX+S/fVgb4SNE9TPOtScgNvTU3uFUqPWrYErcr2XX
Mj6fcGhgXAf/nZxAp+ea6INufvG5MYvpbG3BWnoDuVbKLqg4e6B8lro7/4BvuKMhEfVtL9SgbfgH
un8BWJt1rW+1cHtJhDmImDz7f0UMH8QmNI/FCkrwPBnUgkNIVnyBsKe1Mpttvy3d4dn2fmxjvAuU
+z4gqH5zwlt9M5N0g1yfVNwoVYAPVz6SPVQz5CLsjCZpxo+cWXAiVFd1ic9rggLynsHJ4bdCHqfh
mteRY5XhcCIOF6U0Ct5SvvmNQ2B7QYGLARsmHmAV8NFm1PxJo2o/n7RXsoivgFrjEd6HNnbHJyru
XlFL7QIe3w9dtZKBrfMlIT3CUdkdkpJYFNIOEALt6fFfqvS+Bms7m3APypoPUKlavFAvCgLkEH8r
0CQjNYIa4qUXQLf/TQ8Pg5XwOPLFU+7t/3u5tdkM89m60hz+AyRlYcqz2V/MAxEa8Ng3f3YSN6OW
FDzwkhwFaRr3ZzWw7+4HRbrq5JE9KyDNdtMCmCwEh46q4CoQBcItkXfwU5tKljU0SZ6YsCnqo+BU
lMnULwqTN7/bKHGCIMIz5qTk5IkzD2xXYg9cCgVzr4qb/sGGFjEcDoC0GRbgT8cJpVnWf9mytNMf
eAVs2KLMT3srKhdWk6ohqUbrKsGtuQ3otO7WA20IIi4nDuPY/YwjK9tFHHwjzH/kG9kcKkXljPgM
KcSGkksloUew8WO1oQz+jYZolt2d852G0oZGrppm0Qv1tRNZdNmiitAoRf7K23hpUXjQh7+MA0M4
UvhCbTsIA6sRXyF/VXC69p3lz9BcXX9+xlql0snanTwrLPUOKp55yUdiBlLeYFBxjy0EE4ifwjUx
wzIodr01YbfMWRD1A1/jhPsuBwp+eXpkebs8JXeJ2kxmWHswWMLMVdzX1L2GxJlfIWn9fouKlF3a
AmlFWhnTrSJ//vWRyhsMNU6fQw66vcRgWMaWsMrkTqoFO768RElpXZcvrysxRfYLJeKRotlZie5J
QhGMIpME7uSOX5P1Uaae4F31BVrvzgJsNcKpR70CL3fDx11KvNBKvAdVB7ZgtUucBIND8zpXKHsY
zw1W9c8tdL+sfrqx6pIA4dEDbYlj/0+4UgE9yPW3inAOBbHm0jDfleL+J3MVcWYh8HUhGQ+Y0zgd
uGM20XpY3b0mpvaLoAIbwRTYACsAklMz0O4HLPQzCAH29e/jwgJedGNkfXUmV9nNXEdSFtB9fxqE
sE3RKe49UTBauXm0S3bTUJMurF8j6Ru4s5dwasEVnMJcGTOJv208Tp5j0SxwA/cwG2dLXkHPoNR3
Hm1iSaEo2KUu3sOONmm6t2wjyEHMqceaVUv7+AUu7TZXxWuHEdIzMA/s68FbylUDdKcnfNUBXU3h
SwIHiHy5yJzGF10IKI4hNlPlulI76y2stzvjQxDBbLnCQwqG5IO6SycUcey8mzvmKIcBva8h2Ajj
Q3Lggu/LZgsCp8Kx47riw+lp2pMKmp2fBtbtE0izntC/lmsdJy7uQc/RXqTziWtyA0vmaAZwsdYQ
zL2iuFHnVm1UHUwtJ9TCB5ELxbCOtClrR2iTSwYGqQFEQodj37mioC1ekEPOTpVyr6fn+a9OVrWD
eYEMT1XRn47UJRkw2oUPH9b1hBLqbJ4nPCs1TqME9FS3mXeLiAmYSNqTK0qerSR8si81h1+gcObW
Ytc9DS0SNkbn74Ul1ESOxJ7VytfpO0jyVZ7uKRifT9rN4xIlnZ6L/i2UDoCfez1YklUKvBRR6njy
cXKvSmhNMtczzRUV0eHvfqAEJ8fkzIbsWeaHsOVHl1AaLH27gFjDOoeTJuPCV/EwXG8lRRoX8Ql2
WT/VXMkV26C+nSi8OAPWfyYnd5A3HOojYKhKimFmk+SrYl8sXotxBNRyeeksvgFO4o0P+uqqDjYM
HQ0wc+LTZgVZVqsWR1LAhk7oqI7obvALmT4R47XdV3e9Xnpt1FGqJvobhoAwd8X6w/eHjjHbUXXe
tIANCRmTPMoj9eiKXhtsDiPPz9T8xCKV1lpi/80lM5SfLW1jkwrjbOoCRrSc1E/xIRoUsduWbAfc
w3JNxq86Ppkkr0OYBiJ9Yb+QzlWPLzq3vyv5DzSu1ScxDtkUN1fH79Z8V0ilZ+lehW9MWY9qtdMA
D7VYWhKDr8oao/Ytk17OFG7qSs58vMacGR8aKxXOx2k8C3bRw/Ztrg5l22RAHhf5Xnphp8Pn0m5b
rZ0fYrINJ+qp46E1E8btGoGq0Pj5N9rIIHaRuAGf+9pVFQ9/O9FYzB9EiVrNDfSoyQZoU4sbP3Di
sSStqDXvpAsr6ebMCtPEDTyi49ZjLGABkTdvR0v6GDNX8A+WKCFKhloBBDzwodnSR3MHKxJxMGr9
ZQb98JUjcvCfKQ8GprVBNpLyMVBbaR0iohxWkbhPfMAKZabrteL3nFK7Y7Qhh5+NAZT4DIg6NOBB
MTA/lgwfoNSkwWhzN0fzNo3c7aVED5ulVOiCbk2Nw43D6DDUlVqxBHec0O8dmWd0Dp5Z56v20djR
kDf1rfl4VjKvkxtM8wE0hEt38JQ+CI8OKImbzfVaDgRAQDTYRNuMLee+9hA2g9CKduv6YhjxGGJ2
mviuksuZ+0ruQZc8pYv+DFJXkDfAfrRPsn2p3LaxLrcyVtdFbIMtJf3650rMb/yiKHUlDkjDGL2D
mMcmTyeB+lx3KafEdCCbG3nCYbgLJ8TeS1/AQekVCDG/ME1Cs52XBtajjoYvn1ESQUTjvm5i6rkO
cFUioqxco8ENJZYTtXxzaRGeo/5rGEK9wYZgrBsFHubHI+6F1+KWCr5YaL40/LRhe87gjbZL1Lha
iQ0uBsuSmg/GkKc5y4Xn69bTla357WBKLfWPLA4m4m+nMKe0aSvheNwFbIR3TpzqNIcoMLdEnrmd
tzEYZjCrT458E2R8rN9twA5GyzVUo8mJYxfX+zXYKCkz72Vo4VfpBGeo5BypT16Bbr65uCSvEtHn
SShbrAn3C3aCYhjeC2swnU9CObbFeJFxQJU9IXNjmhJeppB9vKyXdn4Q4K0AGJzS4qsRlM3DOH89
x7RKSAytNimEPSUtTeNQ5qAeteE6rUnBqflXcvloUoC+g1X30LCUP3/Lb2F0H3zBEYzSmq8sDtxy
N5/8Xn6iKfrPA2omtAYjdoKhrVuNInIla5Fbr0FBBTIkji+opHbGPfTDtwj7qEDFhADyVndjVmBk
nPabK3SbB9HLmoHmzqvb3KsGHHnsueOsRNIl5NBZ+xhN94kybDibmwWnPklrbWgKDmNwCgFDo9jj
qSlztMXaEbMt1tHE9AjFhgQW7mMyOvkK77ynLCiX6/WKKwWtP9mU763kexfL6GH4i1psmItItcJG
EusDt0FvsBqwRkDQGvFmE4tyvUmMUCbt6ZMzTHw/vydWSsF7Mq9y26PqwzS5aETXxyb7S9fYyLIp
8SNi+zlYKr5Z7VCre41EHQxY01lq4H9eQkNNxWfeHE79JRwbuyJM0BMZ759v6j4HyBI5htQnXowN
rSpRhaP8/AkNzaF+XKyarlT1tBfaDGXOv4i1DURqVNlG/4Zy+ejx0zY+0NEjtBbe0BoalRutjIGL
TzWWc/soVaC5Dl/Ophp/G8GT86WQKAhmoQWHDb/zBDqELBZso4p41dgz2YesQpZOq0YryAAZMbFv
9PVKDJUaGrlIj8x4beCEpHOK75mUQN8pLTGygVbMer3BU92Z8FQbhIz5K0qKV84P+R5D1eqRAPOO
lQLpHJmO7bLWQRaLWwOGhgnodws53Mf3Ha4SbCELNn5/IjT+cpqqk7OleBMs3FUOh7SpAwzpFra2
Htka91lW8BaDiLBuW/xlbARSA+7UPDmhu/GEQ6IInqtHDDqhUr/xUif25CsItu6wCxz2mb+boWvQ
DT+K7sERVnLxHb73PQ8ro++38eukMtpN0oGzmRB31UcWtvlrHqHAmc/HDHVCsFavP7kawFFl5+iv
uF5+IFQbKpzpp6YTrC4yZTNQiJY7NB6LqGTHZCsgf3b5qXLZcBm4M4n+Y7nLBUCEcnrV4T6Q5DW3
t80ZqUBHgiNQDzCD93TqSxzD5UYRDrbc0zXRhXaallMqHTS2DPvk1xjr+goIpnpYiHYg1Llr97OH
AGyw1VZigJjc6QMcN0iPgFi0ZXH0T92tgyURZ5XPV5IGDLJFZDMAirkYdIOYpnxM/JfFrE3C/KdQ
kgPhG2gjVJa6M4755pIqf56KNCRIukoLN8bcB5xaML9YSMjyk6SexUg4pG+ARDsYpgfWbVkjKFcz
9sfWbmI+95sbq9wmzABAy8CRQvOnau1DxiINPCjDBQUOL8q1f1HN6uzZUlKGAeVUU7gtVpPI+yK8
VqzR2pXnC5LDCLBtqTHChM2AVvbwZro9desQqlnlcmLwbwm7Rc0a+GOsABneXg9gD8HknMqivIJL
nS4DP1mKbcSm9cqweNN492PUGcJVY7GdBXTGmyeJqMncgWBUlSTDM8+YtT1XvxKgCfQxXIjXZgTB
sSH6RGTAElK7dMwPig/9odzBkB3RThesizBegGhSVFVi4FKZd5z5ZPhMtSKILvSY75HGwvMRMTa0
8qdfMC192KAr6Dh5giCDdt7QYsZCqOk/PaV7+rhJGsTxkqPoXt7PpI1CAkstUEtfSgmVgiv4SJ84
0gm+6eRXTYUrVDSFPevIBSLD95g0P0K61g0cQahDGRhqEhewAaRdhaqDggYWWNWqbiwPuJBmzFtc
rWJrmCKE5nn+eKdPVmBVKWAFiY61z+zwvaoD1lO8gwvz71Yh/FRx+0rDc38iHnZKyeNrdXA7WjU9
lfjgUr6X62qFd2LQhUJUc+lLdy3d4Swl3ZRZQE1lGmLwkvjPEbECingDQJIq81J0xylqCwfl/caC
5KcWjFXr1ToLscHKvIXSZQ5va+qk2B1KV0l1uHgy6Ugdn/CTH/SvGjHMhqm4FFGM8rC3+jWpBJwQ
EJFllN/CBDsa0d6xVgkWJep7rV3VpBLTOgbjai5xoVf1OFA8pA/XhdLyL/NHca5/AiQ+Tm4ThvFY
oeEmGJBue4Rh+23SShMqZwV1YIJS7eXfhGkEeglcRtO0s+ddEPBAW25xtjvJdKrkR/Nmu3uf9XZE
x5c/9qlpvL4pJ0luEfkkDuhIWZSPmVw0U+YqjwVjvzRvPgxEccQuDQNoe89XKbqfyMtxwsBr6qKS
jQ4/dJpKc/zKoOhYGOLuqidA8NCyQlJqrrkU8NGPLj5A0jiVU2Oo3RvyVjAIMY/Es0c+8DxZkK9B
wKgh1RoPZWvkTZ1zEBYGuNV2GTzOyO25sv8LxN0yGeHAiBqO7DKvq4VS2P5WE6HNxlKv4abOt0sa
zADoVb/Iec7gjT3KCIBolC27FIVQwvsgD7A6W8XhXX32x2gUOPdEeGt6Vypc1vrThtiUE1kez41b
RYcM1TM+22YC/sZAI76AfaWGMMlCJuwu4ztLa7/imEb9pBDZZqcphQ/Sc/A7L+NhnuFaU3LqgsMM
AIURTkRBYgROM6PFF6b5QgmqGtUxVJkStOiVsGSkHQRTHpaWsoCyxKQJtmJkRxVS4YKZ7PO4Nlle
gsdyC8DTFFqVJUd1dIJanzft9DebuCpPJSryc86ZzVjtmGa22QUN5V6Ihwcnm/InTLwDxoeJ+8Sz
rI3miNmDjbpTLj2Mz6derMZ6K8FeYiuf1i87LX5UvkTJlBv+JBXC4DL4xiEEKVemI/1pCG88L4TQ
etJ5JdE/6Q1xVmWd0JpbQ0CbIWTCbteFhTyBlaIxt7Ac0sGrdx3vfgCtzFk0dYarQtCqOcVfUuc8
idGBmCV3Rit6TTVuTbb1jlaW2z3Qlx6YAZO+kxCb6hSMLp/t37o/NuxOYNAJsVi88eY5CO2DlyWr
V7FeNu96xdr66hNIr1r6v9zwCuotw81Pg/uNeI2qPoO4BrQ7t5RAxfD+CE+foXtWy9HQahLAtUAP
e/yvOyXUVFtP9bwV8Y43l3xxucgkenVtht6cvMpb/QjCAu9E0oQvC/IPCivhyl3e82mt3DGC/LUa
+I0TJsGDxdqGKBLbh7W61kpbQcDxR9n0eoJefAoImBlNZ6/tYwFxnWcqybd5ZIy3SklFKuvglV/H
lt0R0gaj2UrJDpUhRWpx+C1FpSV3DD11r9nEhNNQkLAaKXYQenM3pdToT4P8+2OQIW9Bx4U1aU5Z
tQcZLFPsE1ICLrn9MQlDo9qMuVzzi7fNHHBWkMp7ywOQWjct48U6XrQNt5SzxY0ixW0i7nYPtG5s
OvnsVN/6YNR/lt1ugvbBg4Mo39rI89cT+mn7qQGgTRE3o38kA7mk+/mQvpdvP0PExslaO0nLJ0xn
G6t926rHA34DGKsYZ1LS5Bap1mT0Cc1wReX5v2UQ+4fbuv1KSmhO/q2+IyHbYRwKUDz7dgN6WnZy
a3ASb+Ba7dbDSq/QeXNOkJfmJgKULWpzQGfbpZrXbtxMebvedGxPZxzM2fGb66guLrhQj3aPzOcT
kQc7RgwKtMPUlxA5fZSvudhoOg1WwX2rSM1gGXSN51Q0nP04UZVUeXD+KlHtTkmRqKKrQbG159eT
CuoUbNnROXJjt/H//6I/kbM6phnsv8KOeMEzPjxA1pieiQRt+zjqRR5wB9+TI/IJUixTA0jdDAAZ
2MTUYVdn6DEbxlKMbZQigkdGiANMOOlyZNzJVwZCAZusdt4qCZ8kRxzDwkwdnqPhrjW8TVNwesPS
nnJRo9XESolbrZPTMY5LjUH3O/rAvn6K54AmT4HVXDOU3ubX0HVGVfPBugMCw3yFWxWXrScIuwN1
S8zTcThqkkGSnvqxezxZW5VZH8vum8USTdof9BALic11VqJTl+shUCspdlYrX2lp1IsXsiqrUELA
Nl+whm5IsbP8OhXhZ2nvfthm1SqE2GY1Fn9zwW2mUx2TcHQDhNLa+MNAAfXA7RPgkmdoSUBszZHE
IGsEC0eV4k4GoO/p0Ef+N5ywb5zEIBJ5C6tDn4anUE3UhsaMMI8VKS9n4xrrbcZcV5Acd11yCzdy
pjwdlHG4W2j3xalHUIyTiUmUQzTUmFTNUK9vcUzQBiS7dR3rY2SXxAOvwWbGU5P9zG+Wnj238vw6
lMZhfnr5PMVXkk6R6VhdPG+2OvmUjVc/dKHCvb2qIrsh9wwzT5cUiqpnAeb+9VycZOB7y4nsgjzR
a8bc5eLw7rfVkku8pKn3EEzTRmXZBbvpDyxmEJxu/mIMoabTaRdQbI0GQOfqIoi3FhWn/KlQEaUm
L2qVdO0Y26iCnEU7zX31aBV7so2vqxdpbkcE7XtTB6GkgKu21pDhttIK2rgdg+drxMs6YXCPNJ/Z
dSpYGIyxhAnSkTIs5XZmT02te6t/j+II+hKfE931VZIm6+NGuGjr14CfX+3VnrnGGJ7NzTPU3iR7
6vHOzm0PNNP3w2a5HO3KEwRMAzaSKCkRmFeLpyuW2Wqn9MLnp8uZRWWJiUfT974x2eJH3rs5QJRw
ZOGP5SClaouPjfO5sT+a8Bq9UBBchko8USRonq+/O4nhRIOyvDrpU/2Vqt1tw5TfaIFYT/Nsd2PB
iOAr9fSfeckAIqCa9B6PP1cWMEuMfLahxfTpMZbHCXVhj0fy2q1EVeTt42TptdkJlATjXqGy353k
+t3GpUOu5qr6rBjFVLKepR65QbkE7xJPdZwtJ/v+NWCQFQfFSpqNekipuVDkf4Zmi+8VQ9dqDKoF
3hS37hAzRTrD1ujHog8nu2AK1RnJ/Q40rzNucw+WsUYOiEBex8TpsFHQqEjZ1vHlvMcxGIUfwYqg
I8PZTeW8exBAkKbrkGahUakApyiueX3O7orLbZhcjZF/Hu2OlPXBBL8zq0s7ML0VH6ZRsgvAH5dd
o509/rE39/mzDkGZkSy/fe/TEbXo05Dcyn4XrIBXq2XzObhKJmIBW4X+MF7Irk51CpfQ4NKPAcZa
Cb24OhL2bEgOMAeAhyeCd7TR7hFjIkfmENXc/7GfPRBZKZrpk0SCqDFh+fbxLJCS4Es87UjtUVj6
tLWnSf+NBiEcEANEH6sD1+10b4Y9sgPqaaaP5sKqy5+DQWKngEilc9/255xoI4vw+TnP8fcfQE9t
rwIhxkrt0CugAwY3esEFAelMHW/gbLSuU5yjk8KKueqbPmpQbJg9QyJczN3nmtpYlXCEfgC5dPU8
yXJRAVp7zkw5GcHZbL6Ecmd5DcJh2+E4sgb/dhblLVTENuG2gu4BdMEq/6iL0/+DvJzRNjn7MC+K
k7/qwsRO0UCufw10EGTHo8mxc/enYAmClcbo90NJBVd6+nLjRGEe7XGWuuxUhUqurNyPAD909c0J
aj05KyM0JuOGGW6x2tjlG5pN+vx9NZFv5Zu+BuH8u5kq01UFg9ZTM5VMQv7du+UcwUtU9X6qgmSi
jP8q4qFNGfjm5Z7F+Xu5bGAdFT63sFTI082N3jTNHfRZC407wMlK84QIr/VGoTPBqXxy161VxAIr
pwbgUG7Ohbs6/vcfFeYRVzF+8jvkWGvA0Hj0gr0on7K0hzexgzFyzo4qLJAkQirTPaleoJgBMjpx
5UigzajSuctBm1thz880RqY6X8zYKPWqjoapIoewJRBdpE2s3Kz3bmBpfMYZ7lZXuhpt7vFKRnWW
vaVE1L5VA5VxLAjPzVUj+CG9AMhoM39+h01z8KYysiBZMP7j8yxXUVvm6bEJLoHqGqptBSM8HDBs
gRLqR561blAiEXyEMCReQtHiOMagFtWEKkIVLXV6k7WXklpBP2zjUUHzVAnFVvUFp82bgfPOBhAW
/nNTUL/PGJ1o+ohUSLIFFHTwW4IhsNHXhaB2JM/W1WHF6DptdIVt/WPXJOsziskXt+xO9k6D7ho2
DkTX0m4F+zwGYsuQbSO+Gh2Q1PDEVHyQcuLTpzULeJo+NxouPaWaUFWl0sWduZTCxuNOrQ+7b7H+
ye9Zp8XQaSitYVADolA0FgR/IJXAyiB0vNUa0FK9b1aJgIY5sW9O0RjaFkBD/OvFGZxqSUl3Xao3
ocIDAH3E4Nc9dsqGTHdY86Zu6XJYwB7EKZJ/5b14jzlSrJh/Kjq+Q3W/OeUYKainB+zsqNQv+Fy3
vFf+pD92J+SpklfTMpufx+oXOeFdNUrgCl1ys4KV2zPPQIQ8kctpsv4QOZzLhTco+TTZI4g7lQ+8
eDYD7fbibpbWVLxLPgos6/w5+D32CgFjMXK9t3bM+Zb8+REM+w/hFGg6v0Fanzl76/nmy6UA8eO2
MfddnVCCsz0VKOqsBp1T7H6Qo0RN3YBcVtrSpEs1ou06CBpqPJENSqoNNp+v6u8VoXBzMZRGoAFV
eLV+s9Rze1PnR/s0ihsplK/JqKKQJExylAfyzpSdttV1v9BiKsQc/IIq3VaElEdoVpAc60KlpM/5
WjikUM9tDI5kbTQ2kWX4HY2LCSzyCVRq+kBbcSMZXz2QcsUcAsQ/Ew4zKnXB/GKEcN8R11XKaOSW
ep8DEc5GWnmV4giwDyX7j3D0LN/pY8wWyXKSi6c2cgYccPcbK2CEpBVujuKNyYEPAz9t7WyOoIUp
bL2vksP4Is7lG5VEUj1DC1GK4g7sY1JJRr/j0SQisfaPUkpPc5lw3qE1iseZCz7yw3XourclKGwF
lvWDYkvqW/gHZlUNn8Ec9klIazt4E9+jmsiiszJ4R78OOQV/nibzYIODUOJByAfdC/tAgXNZJwNo
J1BA8Fm0eiLjXrPzPdynu19ruipjrsRt6mfbR1H02L0Bil6dKAEaZwnPsgPvDEpK43hK+FjoeAov
ae19o5ylSkVftQ6iabTSXtfl9m+zfvSerwxxat5dIwqUHwF0gQQMaZOSwg5QGFIoEONwrmHWoINJ
yv+xWhSA+imJTkSgF7B5yTFkjtW5qcACbsl79abCBA1WC4uPmEFxjI8ilfovNGu25x+5R52zWPqB
GZYUyBWKayGMJM14B3+RVZrQKcK3L8KSEBX59DLsqKGzb2TFZn12TjtNFacFt89gjOgoZee+2P2i
osQFH60WSmGZE1vkDLkA1f1tT6ef3ZRjlzGYSYux3m8oV9ylb/Lu6IN/1+LT1vcb4czU1OYgzPoV
KHjb6NiJndV7NB4VKxZFeyM02fVL5QsZ3a7cJZ5bj0fkpk/B1vxIHWvkqrpH4SYYiFdmEDtRmzMY
E4bITrtgdMUFrEEWeyW6Vn90ix9f0fqzueSPaVibPnp+I9Z5QDPSwriaSBmqlE76iKxNs62z0Wp9
gJ+6DwWOZssKj6R1bzoI1YAKTjvmjsXIrwi+Wk3raTSdJWbEl2mXDUoS99oJir7fds22+lQ1+hMQ
8w5/zoCOuwCl2rx8ppDUaLNrc85RMp4KFdFRlPl0y2nWfrQHsqp+Z8ZmFHoRpxgmMP6HYyzFQNsT
uEn/aOQi8r2qTGNTSXA2v2JPlot+yqLRKjuxFzDN4DZJkEiLNm32+8R6RcOoVcEs9pLmpEGqmNJM
1kdvjV2xa+kx4ats4Qa17vz4UUjoKdw5+3/fbOW79Lk4WYUg6rjLQENreuL917mmSIe5Auyzw4n7
oJlRmZGbPlwvNBFoikho/f2yb8Gip+WwiWoQK4orjv0ivJ92o0jTehZlNmzX4mDI78CsswLgRKMD
nme9ThkcG5Kmzz0vHxbbWiWlk5KEsVq1YPH+SZZN8BNpVzTjA86fcZ8h0svvy3dYlINABHyOXcJS
4U4MYwl86SFfSFe62lRQsj8Y33WIk87MD3G1hHtDnBqg+g6+X9p0uF6JNWaZrx77CyYEJsqEIf+B
O+cw8U233Sm1LKULbpTLHO5t01IW7MwkUPLxL584JY7vubxRBulrCNrLGHidnb4gWmQVVLm9tN+H
2PFniQkeTsF1FbTmnMxU6y14n2UC9nT8yYHynbcfk0UezYfdKrXzkgqv68ie0ldzYICw/6RhsBvm
k5PO2IfpODakugTWRhpdNOj8KiW1mywCuQXuSSjFaQgfYWzOqM7my1adCEhLTdWa7KQv4c4RTU86
MFQ5W7HVLugYREDeqRIbYJZW9ytmSgj2eulN9cviHTnCq0Nb/bik/hRg+FnpEqViXjtkD1cIkEIM
I0H6VMAIIVF8FvTZghIHce6L/+Xj53SAg2ypiB+vaxh8Yd07kQx6/YIIatT5GwHlCvHQeAb9NnLK
+/FIi30xjL+l5R5eoxZhcWCZBa3AjtZBe3yhjk0b9XRLQZPoUDhC1qR9J+zaJx29wD6qkDLOCsQV
OlWdfTMRRWKH6h3621/KNP8PMMKG1JW/n/175kjiZxkZPP+VcyqAwJO/fwu/W0O0AmkLirfRSo9s
2p9JCWDCsSpG3Klkds2+cH9znTVezXwedO7AmJ2fdsluAg3Xu9szSN7FxYs7hwcVxD6BezXMHB6o
EdJTFeV9IZK7SEBRadNaFy5iylRNfQNe8xMKjtjATQN6Gj8UzGFVqiXzkvJMHWuqhNEw53QGPBuv
7nT53lVXc0//IscJ+k0JbuOAxNrAH7yCpTFoXhEJtXL0RmVEb1/vxmIIBz9C/x22Vdci+hxOVZY7
bF4k9myTC7QbPTvAZ7z0ZHmSlRjZekw6mS0TF/S71cvIC6xnV3h9lXXQcAsoNr+0sXDkHp1ki+2r
hhnI5lMGrJ4hYkpoyngG6PJLN9tCG5US37UH7mqFKblpPT/PDKLx545ycpxInow75mg/53s1Cwbo
7v/6CjcYBIZmlbFSQKtYc3tiABlD3I9sjoTB54Vd3L3/GRvTyNAlRsU/9bGQ5RTnthmYZZbB8IUw
zx4uGjfo6/bmXl5n47ASAQxjA37YjfSI6ogfFsD4Uj2hNiaL6RqwjReZPDtMV4KopkAym2ErPxqH
jY7tuBNLANi49axh4bjZ2kGR8pa3EMMTwYll8K7faWlAUGvNs/uTNd9kvxSYKa5XI98F9fHybCgt
xpIxJR5z1ygUoqKDpGf2wGOWI8VrvvGlskrkaFjKUzHQyZCW/iVDaIQmSi8mnm8ivU6c2qpSmBm0
eLC4YrnvUW+9QMNkTWBEAmYACYRs5zKLZFhHVnyfrJpX6/7cZ/p5LnEN5It4HGQW1j+JNrcDMyHf
PVi5QGdk/4jHQ7ltYq1pD+KhI1XiTu+qCHbaOSM6Kq2m/zBLfBhfIS0KQTsW3tD+VmPIHpFKIX+H
HjCrkzh7UzhGytczIzjmCob60tPESqRZdpii8QvrBeeevqBKoU8RqYsPSfvQGjSfz1NSfbMN0LBH
dJ8l74lJ3Z/fpoX6V2UdgBknsWt/Y0r0PcKaN15kcWbp35ASHf21poPnl5wfaK4JY3b968uyqnAo
i8NpaakNz2fzeMzntyJv8lOr3NTJzBJuJMctorQE2cokO8uCbduhGPTCp1Fygovs5ZGZxJmWPr0n
H3B+wDXp1fhGfVD6ZKZMqMVPskhiVawUoHJl0853eMEkKJcGPYAokh28U6PNITgBCcgFXE1edFbk
hM34dHGcbokaOrSVSv7R+q1Jg6fUbwyWu0a7V8U84eTyCBZg8JoxiEuhRpWrP05VE9qjE+Jb95UC
ij4YT5AqLF4XRAowDBqmXyx5Rigt+rWxtFrn6/1zvalO/EIh6ZMlVe3k+mF6egWyaYpb97cOtHvI
tuK5QovjW/6b6Fbuddfl2BjohRim5Zz02xrMs6VfkaPtDI1unnJeu21hoYz80ke0oG+7K/h838VX
V8o7B+Ni8o63xSygR+t/dKyx2zF8qtjuYEdbJy3bNVAcp9DbxfAOhd2wpj73OgXQe/RhySAaeKk1
FNAiXhblc94QzV+P2cLoxausro8Own79SSC80Wdno9U2JTWKcMiqaseB+DUrMwW2WGVE9c/jTtsR
lb+YsJG9wM4u/h2xNf5pRwd17jUf04K7TRp0nBlIhjpalnCwNrVKb8fWhQz7VU38+/VWB7V6ogf+
KP5aUz0qdxC++BSo9eoQMzBdLzbjJJtCb96mmk4/b6N+3sKBmQ2ykgG17QKHs0CB/wjn1gXFrlKb
zwsUbSzsrwcAuOTKFMrlHmwJo3YOK6WdMO892+BMazsSwb19vixHQa/TN7jDGPGUVkvreVI4ynsg
Y2mPpVwtQyuBwiK2Vd89dxndm3laiCni51B4T1WYA0+r6m+UOLij2IO973gPV0zKaCnOmqAdiTRg
/z78lT++dsu3+opRrTKKoDQbG279aa2VSzkVBAFoOODR2r9GT32MWfGWAqwlcBwgBuVBqC69D09M
VrHG4cVKWJBmFhNy3hsxdftTJgJg3Ujlp7Xjxr0Fakz38EGbN0J1SCFAlti233vgOZjXnlTlOURL
14/zb3Lc+Dq8W9LAGPGuy0bp/jksw5yizmVXxsdx2gY14MgpOaXrPbkJGPRKUTbTel0I7UacsP+W
c2ZCdyxu9v/NyAlBtD3fRvUTUKpZaWJsMH4iNnR2v1b1Mw0dz+Y2BvxLedMF0313tbiibfNtTR3B
FiiECj3KWLdWy6uJVGzI+PI9wmu2X1YOVzTSG9OK9IPTxP1j+5QXSrAVWS6jkATWkGT6Ha1hlVMG
V96spbAibTPVLyHvxTK8Msyz6u0AYi8na05K1H2AQr1+jUzl/qR64T9LN/u5p3f33ACOs6j1566U
yt23c19/3Zh5gPX1WFcc3zgh7tGHfR2OwRHdKRURfKWBf+Aznu5p/fy38F0LwlfNUW0px7n3nOkD
gxO9KPLZZdNXoGg1p78Ulm9u42+Axi5kTYczooI5elowR8/Y+ZKv57P499QJJe8k2uWGAFuWuAIX
+z+UgbZto57qr1f5PUkKrJgUhKpEjmVa43jLkDgt8FwWbtc3yEM9mFTRunnafTxw/LYm0k/5YhLG
EnEkXddm0c2tOvFqu5/P4U9LDLSwE1FfqESqSMHXNkfWbjtALhD7IOYGV6kY39fe3M3Z1GzUZIBD
o5ivemEqNwzE/xDq7MIg3b8vnY25muUrySqEF0VHeWtcHZGuHp402MK0uFvuEcfebBQkQ1cbJEPm
csO1PBMFM8Y+GD9+M9laI3sOmRzsMrYsNHHy1kqoh2Imn7fmfhxfV2ARlBLzt/wMEmS5P36XnrO2
xhAa/kaW1hrW99q16WZ3eyh3g7nUtBAdd3pzZ3t9HlQWbFcKQ102qa4JePaav01yDI0+ndzACMyD
v54HEEFGInlSzfuZtOrOOxnlFoWc1vR+T+6PFRqMPfjJi4+46m8rcpo6IBLM5bdiPdx8aL+ZIyEu
A51Qs2FtOl5xANIdvupL9RxanYdPO7VKSnpeaA3oU/jEzzvmMnXD6RB9A3AtJEQ8TkTuVs5vqKgc
V0VtNqFUwXef3UqAL3EAAJAlCpvD2myxoV38AskwUdGoIhQmWboQXKEf2PMrJR8M7X8b1pUCz+oY
2dw/6UB0bnlFdWBpHQe4va/s7aKMPIUvbDgYO8GVjP7EXYMTIxDhsdL0whqcVhhFe6UtlNNbtI+f
522c/uILoiElzd66e0OlCop03BOIQukd6EnSRJGznfm/dgatJRU7SV30tY0vT0YZqrflgEEwiEKI
vCbNWz4Nx8S02UGam12djWw6eNRq1lnbhShXeXjwe3zrsqnglqRLC9bjF1YRbYZZgayWoRupNGb3
qat2xoT1hism/2IZnbdDAt6UAbrrU3Rmdf1oGHVJaI9p9+3mfoXXtgVCod+K5tFEXEyXdLApQDaI
kp7G7SeD0hoL0g5e6ywuv/NC2pxWCXX2GWD6dERJ6mEDRzff0r1/BvMs4C/YKjBzUGnjJvUxgkbe
HvHyaEaIafgdJqn2sOJdbxj4HfamW+FqZCxmhyYdj2sIU0NDKNQaqOI3uoNHPt/mm1/VZNJEvdnv
NZbBWUfTRjcFr4BER0xwcQ03jQgpynQ3cp+kRF7ihOZz/UNi9GOtrUvs26BJdCJ62yW9dKHpp8xY
KieDS/uysXlhii+n+uec8eGJndTyL8mea7Z2SHV8YNpjQAzVhawRWknm2Awa4zXfQk9jCWzN+J1l
lRl6RF5U22CnLaFSoHfGrnBAr5fDrN91uqSfv2KU0483bytV0unYrRxv/sjcnPDM5pfh5Im3UZ2X
3fesGN5aAduTD4iV6PWbNtPWXQKt5AgtDq984S56aQ6quH6LDxDpjgILBc/haheO5ObqfDOXAfIO
f/U7Tt/z2uD5r3viy7wI/r/hnU+h4n1iFcOl5jhcTl691SDuQclCWVrIJAaWiKROGcPMVPhTN/7i
l6aOt6QqCFFld9YKKf5KoSgLprB3pRf2KT1yCRfGtRtMo7fpVuBGRLxNdAMrEZM24tyV3dgIqvon
sWEkYS6LwcB3/ViyD/aW9A0mvnqVapHlTNGwe1KvcpSLCY1lWs+8tAoXKoLXWMk3xwT4s/llcAcR
GhT85ADyyfixPe7e5vpm02iQ68u1anjpOHpdp10vsEsw6w9HpHwGGFp7HPIsHlbsKDvAL2Jf5ERf
Xxlrh+jdVpg7nXT0MfsIH4yj/2D34Z/vKm1yx4RF+0rFcq3i0STrntCqKFbbUB3cWUMiHL8+pZB2
oM87yzF/CnAEHIuFpITQ8JJKu3/IQdZkg32qIrn0huY0Rg7Ut0xFWxhTLs5JCZ2mg9jp6tHfGu38
PGpwwYRHw8TbWSFhVwfUeVUrjRXztoTdGlQF3B5kPgdcVfuNSo6BL26DYXo0MtA/g2O2xFeQFrsG
ZQcRNJQhB6Xo25K2Y76bApAxLzpXcuVXpXDb0GwrxJT5tPKDk5iA44cKETK3zZR0pIaLAZX2o3xE
a4kdgKNwBWGYimuYLGN8YbCvgE7dPoiR6jx9E7mY07iqOrBZmE2lVpjHWgmYVlxTzeJO+13l8yua
z163djRxt7FS3aNV2Da0CTxuu1uDS83DDx9rSMUaj9/M0Xh8hkivzoyGJydi9koHe4xUXrU94/uQ
aDl6VeYO8M4w9OOvgojyBHVj0DFB7LNranMGq12pUGjpDVo00fzCqRIlvrlrSbT6aWdgShWy8gcH
moK9rbJ7lUgE1Toi2bMw80n7LY4Qh6j54finhZxP78OMQfFTYVjHoxLHkZZTPW9LQJu1OSIpaBcx
9MfjyHC75XkZh2e1Sw8Pg5EosboKjboZTY9iZMn5JM1FVAAhGJqJEA+/RfAG2iQFEE0YITTbTJIQ
VBYP+oyvnxU6SAUXVd5a2m73/4nwGbwBfMJyp/7z4CcyD+7uYvEaGNRjCEWdvOcRC2IPVAWFKIXc
ZL4g89BVrZ2AouSmdr25yDUX9uTUXybuAuGz2fI1zoQd5hgGme5bouTh0XNiC4p2D0DQR1QvXnLE
wO4ZOsXQxyBSHh4hgMxk+QTeP7CI0Ut1AOji6jk/4Lbj2bVllyrupiHXAyLqncev8V+FqCM3EOb1
eSZsA+rb+QwifJxk7eP/kx5BlnC7XGU9mkDwJ1tbzanuTVo+opog8ljWebyPeptarL9eR1oJ0cqB
UeQ/NI2IZvragstkrggGfBdU6ByL0yghBQR3iVnCvnbj40BsSQrQ8lP5ihmEtFRjQF1+Sj9idhME
9St6a/QyjQ2cQbvXG9fGmATqXYP+7bQl0HrMOCYP8jj2O5gMpY7OUvOnrGSyMANoKcrfU2V90pR0
dWP7wU1jXkVbdLpZLwckvU+b0SQW72OLupmII9qZ6i4DgW9nD3BfUse80pWZ4LeyXlKMl/WU+d9U
MQf5bvABnFVe6rRLX5bo8NU7MNoOgNi7nNVetC+1cd3Mb9wQXNbB2X52xa7oBtS1b52W5+iQXVN6
yvnzyam1RHCGxgzfjUxuk+TUu0JlCgvE8MqoAN03oVoV3GwCXaQkp98FBMpkNOr2svEZhbqiG4w+
xfm6IHPyoWUKXeXrThqpwlh1M+Zz2aptwkgydfajikewoCRY2gwM7GXyqhkupAlXXqHc+gPWN3q4
mXf6lQwLzNfiYqaAitQZEL+41l4BpClbfmn59s30xV1k/4IZTUcCbf+gK7H/gdJvG8mhGEvckx2C
fm8ARdqCVS/8sqqzHIfKOuVQFh03s4hdLz145APYGJKxypNEu8+D8kRcCcMYILFoXRWOKORE1tBu
a3mct1gUVp4zemwqMiFypZdUFdzpB6TO6YILBHlm6+UJj2PrTB32HbBET+3diw6xXY1xhJHP/x56
3FidxzyQgCMx4owfgb5gEn7IwArHiQLydPYVpB9Y3q28PyHuw8vULGJZdvP5Z0uWY/rzMSqlMjFu
SFiQTRcmYhF4umgtRD2wuMxPFXT1OyIQ8uzbkyscRn0JJmyqVa5KRDQNy77ZNHwggNFRLZySM7Pj
DjnWpVLH8vQacKQYR9mUweg9RbhnM9/JI7AZ0b3XV4zy2UyECUW7kP5FRbWbFv0tbaz+7cwut365
44wDQWd/wVdz1oe4wT2JWyZqbKaTsw3tyRFzwe8gJxSgX7QeELHeiHkPWBfbJpdeqCWDIch6DBZt
CGUP6SphXemb1fKyyUDzbeOwEvZaWXkBadazm3cy5zjo7mSSlWtL6MfGnsNXdJIyXSm6CYgswPWw
V6yeE09DEUl4BLL4WB2tcfiSdiOMcHqH6dyLr0pfkWw0DBs5uKjxrLPbsS2N3Co48kPaQ1lRGVkR
M4kl6WqGqluyGMgcE8F02wJM+Y/a3hKk8/oLaur0jgX8IzLJCcRkQB/fvR7RM72sWJJoMXkn64BW
TS+mcF/FT9nu1GaPzqCQZnxXqKFGDtTcRaSwR8sEZHkLcf8BtSAXQGEhPMj9YKXwL94tq5AXl6nU
d4naO0D6elZr2qygsL+7ZlYe0fdfIgNI61a0RgEYcWSr3sgf1S1Lm0oK6C1EDuEU/3a1haONdLVU
e/pXwXH89/vDBlLzMV4/TfHGgkOkh55oDe5aNnTKbroLgyW6U9tTjYxfUUCZsJ9SnBaCLZENzLcP
LTtha3ZcbombvBacSCYGBdHqHEDR237Y5g/qUmn0LnT64LS3lDyxrvb1c7sZQkJK4HXThp+PIKqh
+DdAhzqG2G5p835c/8U6/y41g5z2Gdn7AIFx9408RdPFF6gEqu4sdtiL0cakLFfRUnuBcVc1/D1f
NbfRnHSr4HCZgYDf9Z6ui3vX6s7mfahP/DIriqumcbuUnEnDiV71j41+0WgpGwURBHr6as0d0DHJ
1fLa88TwoBu4GmrSaqBTFSXQtfKjhCvdRXtOyNhIyx4YbpPsQGwOePuX2eKlUPSUNDzl75ZCOqRc
y0uwOZ8LlpsD+gf3wCvmFdnZDPLQt7tnNoGQRbL/WDGRZYQaNGz6A/23cMhqKKO9v3cXUiUvUaNS
SVUcJhQHdL+flYS7zaXyNyyrG0oLTS+Df1P6HW/NlO9ac09X8qKQCIWGu86qZt82HJferIbgziv9
FS5seT+dqbas9GR5MdIIlTMSOtLYsb/kdSEwv0VQnaZ3mfFf/B6J5vpP7AJ+mDmd/7CmKXYiJdd1
1WxO1asfwFwgDevWMwPlGOhvzVfD1EBsmJgUs2JyiIljB++n2UHXHG5GI35xXJtvv9lLuztqxiDU
xf5xbhh0O36yNgJCm9Vw8FJUoRMimkmbRqdS/o8of1mTSJgHe//+kb84dt7ndzEMQKFy52pAqNMH
zFYaKDahgpwKVwR57IJdf36DmOekbj5vcZqcokx5WFyM1/mCYOmOeW4sWRUyx6ekXJiNBCqJFS5w
s5vn2eTVh0jnv/DWUUo1ilhMHEy803bi5kK2dj3CJQc69uCOBdPl7Ojyu8r1cNUkJarjYDJKuUjI
IobLXvH1I8ar5xrKOgy/wP11GkVUi1syVEmParNnoLp01M/LTMwKlqWihB7chdaW9hYUGSxBdpvI
zSPu5DctXl468UFGbg/SqyFHycib56QgDx4ZEGtAaXarVnNvSUddUGl0byW6TkV9igd/Kbo6a2h6
/KELaOfWUWqzqh+1v8kZMyUWoAU6KLRydcPkns3/wJMnSMHs5NT/n/Eg+jmQwg10UBnEpZJPsuUE
LbeA4IKgOpdRi4nUEY5q9C1bpS3SrB3pmV3PIyE6bNgZGBt4AhzHFaVV87x3mV3tLKLThJZMt9iA
FXPwFKo4kirEvW82zgC5l37POySGw/clP7UDUaXYN7UBQXCxlpApxn9wAwDU3wieM1Gb1lHCt/ix
qxFIsmchspVMz+/pNGH3pF7OpD3kB5KdixBls40YZz+byOyTb+Bkx7xMtdZmv1Wc2MUnKJMW33Cb
dia5CVPRT5qh1OCBbFNuULeFuOCBBkvgLIC9H43UArZKLPluJGgX3B7vXzBwsMaPppr68R8LE/uZ
x7Pw7XX7ZPq4og6PKNyJngXRC2WqcQA1dl0nzx/gqFhPkhcqvoYM55unmSNCp4eIKX5pNf7oqEMc
PGoTjhD9ztVsQmbheqH3AQCzO/ooJ5JeNkm0MEj5glczSamuJcWhKToK0CNT8HnKI6h86XqmgDPD
BEasqusNF5LHmdRGWJuRFw554JWcs+tbMZZ+IxXj+Ju9Xolo4a9dnyFHmksno8MdbNQSnSzNwxIM
sTjbQc80FB8VOZ5TEu4gsd5e4hJmb14RFE/yBVHwyD91YmoHUkwGb7LR+dv0F1pQjlaYTBQGKxw0
qGsQBkxSLzo3czQpDkq1KzIAKsmcF0reNfg8oFO64tlFigePXAcJTuJRwQ8552K/WMZFkIx4315W
qGeB/XmIlQK8QOvqCT+FUHkHvCU5BJg7HRsSotkUql2F264h3r3EopbX8MhGLQdBnOFkOGU9Cxpc
AiIz1buNzvdSts/XOF/VB6224dEbIuqCx+ROoFpsA3Kkf0uOP2gHBcYdcoxXsVU5g4BK2svqAzq1
BIsn4xM0oQHuEwd02FeVZIedb6bYgYHBAWNl1eBPjYwma4F7wsFcy4Wtt8vPs77bjO8ZEG0Xn9q4
5Sc5dhWHVHc15fw54mgBwlzO68QacqdmAfkRn5S/ZZOl3BSyI4p23MxYfIuRTmEi8bJ4RIESKZC9
LCvq86iA2MRVhMsMeePiVKM8m+8fjZO8v21fr4zbI3s+TveDo878iOInhXDifi3gMjtyYL7ijS68
s2iUSoC/r9G0ahs2Zm5XVM/mykzAPBvOueD1KpBezf2s8TeDjHU+S2zQOhVTb4D/36vxdaC4ZGA8
iTl99TQ6egpX5RFMUoZAY9gs+wVA+J+5bioBsdhhKdd7bLA16LccMOtl/1esWlt9AX7xwrfcRoHi
7PXONIUusOyA6FdcQefkjyoMyCKGQvI6uZsSCja1+rC3kbWp8ggnXdQR/GUlWW4b4+vJE1rKWFkd
jUXNDFBJ2DjnrCnwMsw96SClZ6Sagj808DmsFnpE2eT1fcQPcZEUVFckFVsYOZGt09d21tE+31mZ
e/3fzJ/jlpQSfHPU6gq0pFx6gPHUzgswBMQlyGiYSi6PozZw3N/8CE8oHOTdFEnOYki5ObFQ1Fam
bgpiQFFDVA4GdpzusJO+PNRSxW5zxQb10WcZOKYSF4Rjb8x/ymKHuGK6Fdoh0jqbSYAwzHTrKTIe
Wtu5hIHzvZ7PCWFX01XDEPWbYM4xxbj4v9GnNSijAqp9IjVxPStfLLoz/l0eSNwxEW4+7TraLzPa
SAr9lsM8pSfKwNr1gLaKXrT/S2BaRlL2wbDN0JZFSE48vgnbephPX0rv8mPDx7JeWY/WC0jwOHoo
o562ara59NkkeKIlD74tHbSL7ipWuod5OGsQkglbFZigE4+/hZru59J2sVoxHenjAp6/S0EibW5c
tQJcxiAx8+JyKy0NFGyuGNLXV5bQKd26Rc5aQ2+j74cSkCkjAjCttCwnYa779Jz4DjoPakc/q2Vf
F7yRAXmDZGTx+9zSCNXn6BFBPi1JLRlTyr0WD9lpk2Shd3IFCn1gnKHWJvlRemeSCeBXQscGKkgq
F3xYryX3L/zQyZf1PPngzWVRbA24tN7RCpJ0sb4ERlllSgBUHseOMulHZCOlCxjOq6o3I7yLJR09
DApA8qpOwHuNHq15lUgACz4ZPuMwvyy4A4FP6/EHM8liCGyJZTI9OIlmnPE/iw+M1YhrX8zbHwZV
T/mXFeaJV6J1P3d9lfYa+d7F9ZEy9dFoskB1+QILPY1KGekuo3xd6QlNyS629DvB7ey/21pULH8t
53xl544+9kwNBiaVS75GzAptLlnveud1mH8c8K124HH3CljlZQXJQePSPRZMen4PJrJHMeWk7xRy
M4JHxK4IH4c3Mi1i2EtkJT5tIC0NHi+XitJFuKeze/pMjfBCSPSgVCFncr/SHMuxq/MAlW/OUqdV
NzxWg29VHZsuSXtA+z1i0fnznx6DshsClgIMilswsXQPQigjn1KscwNndGqOAr7GLlOSu7q1JeQs
pf09njOdtbYp7amK5sYylSYs6O9ZoGVcFDQtLzRtO/26aGfOEvB+m2IfF8O12QpcXdU8CtVgFiZh
Fqz23M0N+uxXW5cQB3pDlGEHJsKcKf9zzbNnnChFO5IdgbvVYkjpQESL2d1USv9J1k4pHfoCWqt/
yrLiggU0+Gn76j3nk8d6xvem1SQ1zcoSjpD+ZRCSQDMziFJ41EgOMTntUXDLtNAhXeOJtZn0z8DY
SAH9alg3TZ0ZsG4ptCOI8qCthN1AJNTx7x4cQEuB3tceY+P95iTlEtQjIE5Ltj/jARg4UoLEQZKG
6U0Z0dI4eRn4mbVMt3yfXmSD7KKp3TxI+MddAtZFEOJgYkFKzpaN3xqKp03fS3JwXdcYiYVPSkFq
Lkj3vd7kf8zdsgzDaslSiOD84m7Vv0/FwMbBZDC1ALzvI8V+/7t+mNfvxdXHL8ExlFJPwOYLorG3
PPyEy2YTgpsIKnn52BOxT1ZJpeQnNHL7SQinecYw2FLL1aavVwfOg2uIEI7AlH/LcLIYl0clGIWn
Bokwe5Yxu8TpERZsfeDpKbpS+3CSVhfq6Chc4vqTpqv4eRe5th91nLwS2xbFTNBUbbRq73ORx1Xb
b8BOYn+yUqK35wspeE0NPGWZ2SRA9ljZsW5ggf+Ao14Rjokf1TY8uhO2ftkMoOByQURWJd2odWQB
LW92hMBOc6zMiKX6rePm7nih2T1msKz8SMQlRRRhTmkp5dFx/lwJzeln3NG2cnkds3nvcdKJ9izi
VOkPGrgfDyjEKmCtSo24/lxxxPzzyNnjQeoSIb0RcMTbZ4ncSvBOhDRDAyhHvW/TJQS2ybnm9jzN
IM2nT9jXuAafMCTV+8kOzqXwoIqFtanNKmTe+Mh0w+AdFa0STNCMKBCnpLNqzIc4vTP46GSStwdm
YUHcrAA73EVZDQLQPaPo04RDqPhIX8MietKfDny02jsOjUFYp1LkUQIt43Kg4s1RV6QBqO6Lfu5q
AN0vh1Tn1vdFQ1U25qRxzeKqT4JFG/B1ueK4Li1/XjPE1GWE5cGGJebEj/7p0gjic9g+oRIpwzcM
ocoBh+qIDFiJuVSh6mfvNH+p/snQwGootEQdIPf1d2LrHML/j9NvvcearAwUcD3ksneO9819SeLD
L+oSPXmi2Cy0o1wk7qf+puEsnbb4fL1soTQ9yzCpQPVeKn2WKW9ZKw/1h26Tp7jPo+Sy2NPKGztm
+qnnvqIwlJ02/FUCCRjZHH0AS/QsooGvNYPrBBf6ROvg2N86jF7GKMtocRYzc76kvEHIYhBnPFwz
GKIhR3c9ArhcH6LoJbNt8tOxzIafgfRy6BOtjqKHgwb7QjQ0hKiPsRw0ppskffftPPpIVjqG0k2u
PL1R2FaiL9gtx2miAZZdjdW1/Bed/ieQdzXHBRwGaHSoPnVQzBjWcAsTEwdOIqHtE5WNvd6ILZHb
p5b+v1yNeaXJKVjEJzT7dE24eOwN8kqyUDae6F539Sn9NTkfNnGs59VQJAN6ZoKvVeyhXqwBi68D
ZYBu3QVCeuSkmSPnQob3DvS9VvQCoGj2TYqysavYxzAEvRewXx16KqRZfwjFj51iNoJt5SZo43NF
9G8u803vsVsvBkrBqH/BY92d7wItlf6XY07u4RldLET/yeht9cbAusNqkziFlMNsvUOg87W0sQ+o
dUcNW0bnoFJHNEby7EQYqKypF7E1TophstaddxE3yJQPbtCis9DeuEZYCQ+7QUlfjD8v7L3ltnLF
drt0GKlocBF+b3HlzfNyk5cZJZcydkLlK2fw7ZTAE7sOib9rcfrsB/WBoxc+yvN9Ks9YZetws1p3
WeQwUOFFgMC5ufoJs7xQf1rIUKSoX1CC6qaNIb5wrwX9PVVnjdZsYAfeSeKFK/I8ZOqy7goDdXnb
FuTJBBlAb3SRt3XdbL/D1W1zhFBSpiNyAs+lDWKosgdCwr+ZXK1NT+98yU0m3+LXemTJP/4rvepZ
CXMIF1QTWx60GnQMWp04WJAw9yYWpOU4ZwisZhygqzl1m+yOgis7qTBvizcrzFBZkuhIsg2maezz
SzEttZq6pbFE32V2msWNJfiuVo7gr744U94ZkYESl3kkSY9X7MBCUBEYTLsc4NyDZqhEWvpugCXh
/m6D6U7hrde+0gIqmbRs7byl5EXel98Q8RppCTn6sgDgJI2itt4lJyg4eEqtxRUW0q6ouLIIdExo
YzWz39Nwv5IJE4CHFheqhHEG9izAvHqnAa+NyoKZmNwBnsOMKQwefFBVP+X7GTjZJcBSpH7zJcfU
8/eF3dOBgtr6e9+5QZted8hb93fOBCnFt6yAkfu1pOuur0A+dfOKfyZRMdKIVdq6PQrPbnHPGOkJ
Lypfh3VUs6G5sSXhgAIN0AOv+vsmw064Zd5Eet84ruBl/aKbMFo01WS+Y+bFZ1Z4Y5nCPz/1LC18
JovKROK+3F/wlMsSiIGM8cxJfnOuelMehFKP1dpf234uKNZgbXQ9660+rzBbV3C+uwTu36pkuE/D
sQ9L3AButeHjnX4gGqRb8IS3uXb7M5e5xWy+9Ae3RSLj5SkdoV3u/digdYdcmwsAPCMUmP0s0l6F
fy6mFGTPHqQpL6jTCAnjN4TUYiSVPUpCQkkLbH/mlY/NjqufAkDcIHsTkT80APJ66zVEiTafwmP0
KZJtz506IK5Gu/+ab9FsxQCXRk3QYOu2MzgOcluSBuQ4Wek7/0WtoYAmEjB0badDXdUK8RN31jbX
LDNPK8PQuNwhajAHdQSG9t0NYWJ0xiSqy2jhJd42y2TCloyQYsmD9OjQz6EuUfyFfaNniP2ZHgeF
IzixdUI39G6pU18Tg5iluqZMDIGpombzCPdXw6BXJhSGyEOWc3ypA2A80EBpSQjYGffLJzpMMejQ
WHrEIVeAUPWMS4cUiw8TSWJcFDx+qE6EHnOnVGUB7x+03Q0fhJT0AHTbqWGEmkFL9irepBKHS/Gr
fgM7RiFM6mBgTdpsRtrhR6fO9GA2icbFMjjHald+wxn93JdkSgeJJ/Mx/C70YZd2C5Aq/0P/LS52
FOPvtbbywjBYmtL0adgNXwk+rTYhkegGMs2FwI648H1QLrqqTbM1V7l+FJCZCARbqxrYdx2YiAg7
IwWNQFRLrEy9duN54YI9hrrk4lqmqfob/2ndCaPT2TGbpEL/7uUsObXS9+x3dF562844miiE31NA
k2YG+p9BF5r0K0TCl4DPeex429ovK48QeQpFX0bqK/JLxnM0NK+T3/88JC18OTd8/o2eTdhI72uk
/ZfWRFu6MYz+6OsJXW5uNxFjppkjckqzu28wigDsXVb0Srz1pC+82dCNJu3TK+kcANfZi8IFwNVw
Ss+hvkOfy48giSJEGBs9943zpBPg6DgPcWotRyKVV8EbR+cg8rn7KtrjvsIfMgQOzr53NKKu79OJ
+LBgpqYkq2+Bt7tc1WvIwY4U8CBAX9n1r9nuCqHX+c4zTLR5zv9F/lTvJMJ6jOKl6mU8JNL234v0
gYaKy0kLPqpiVkTCaMr9/S6EJF9iiNkq+Rj6Tft1criUYlktaE1UvXfHwd+Abc8Yww4NDkan73vA
uKq3axtQiqC+ZpNSdhdrL8bwmvf4r5Rc23PoXby9OhK0Se3fCJHaMDja/myiYplsq1oUyQ9HsXw/
4BDAS5v0KFZs0gnqpUxtD9RDXm1uecpJE9btOd5wIpN2hAMc8gc6GVVsFrWF8zjfQ7mgPlnt5Rjr
+xZjPCxdlrttJomTm4lCH131bOHrMKR6ORmmlj49ESU5O45tjt3bhbdRWwDuF+Zn1fIyvLyi6wLR
5KkY22QwpQSbA5/kqBURifN4eHcoHCtR/C1JtO0BB1u335/JQIlNvIhhwZrBgM5SAPzqJrdLBtSP
SSH2wxAVqyjTC1flq+1GPJt84yq1E3BIsBTmT4YoqsXPEpQhkIH+qylyDQLUbNhT3TBXSw4q5AhT
4CYpU770TAW24wlWaIcpW2FR2YQsgpWjVBiDBgazwKzKWGPDx8zZRBmbUa/1aC8ar+EJY9PPVMzE
mRGlty331uMXXdmL1SjRwTJCZa+uxQtg07YFEmILkzFZNdCqYkq48kOZ17iV2r7iCJUfHCPLoik9
T1GVSlRH79jQ0tuK2FPI+fwf7LLyXtQR5E2uL9U/4NyTERARYCSGDHZVaZMjd72ugIhtPDiTC6Kj
jzBep6jwYxK1qjZi6ngDKPQd88iDAznNvabYSFz7DKKJoZSh2RqnFogoHP/9yn67m9KanqidJv5s
4xrxrQazznED9hYcj3DQ2HK6x5Gx69HJNcZpj4cxvChEXHDrbqgcCNB1MA7iD5epawf3HOYQbxGx
lKACgTO/P8bDFwglOMAiTEz1h0VpCjzeioCFWMm4v+aNrzFQcWyn5DNa+sBBGbxeWTsOViNVRkkY
DeOKC4kWQuAK+PiAMbpVaeTjInYmiOop1fRYrktgWUCOfueMqpWCEJvLcMiEZfwX+JeuJ6v9aQ8v
I+CS1LAzqsGu6eKO3KuRaai2hEze3BjG7ue9Z5M20EplTolvRRV+TGKLIhbflcLn4sD0RLB0TnTi
j//u8oJSHIdCa+fgR+jIy6w4fhnxebaQXqaBrG4+EYiR4aLllfEDxcsjGFlwfdWIVRTfWkkwrgyr
aFvk2NMQTZ/T+pA26fQL7ypwi0T9SMSWjXeoP4D48UhKZCsSOavrls6GEBV1N0NdwCSWmjEXU9CE
vhyKG01tg0ADuH9HrIdu7YCYG6ltVYc0MIvlErs6yCbpRyOO7Qdvs7Tf8iOlbW5Fe/5Wvmo6H9uU
/CdiriBWxZNlICXuq8b6dWFn2D+SnmTQyxCwEGOVYoCZRt5al9RDrLhmT/SJ0cBnVQAoaYHwlQIS
ZajHLkcbOThcoZAnVKSJ5BHwjVANMc4R5C0x9EkerHvI/afLgQVrbEg3H2fdJsRKeqBFKmySRbQN
pd/SX0R66CGSKhwum5rtdeO5dIE8vzVYijjKT5hNfmFTHUAHdzupKL64/Z9Y2WdC0TsJUbLW7lxi
xjBXGT4hM836r36M8m3diXdWKKGktS7WXhsDomEdbAoYwWyBriWaxPIvmTLcAkZ14i08vrplJe+k
v9+vxPbBZ8MkHf83JptkydqMjsl7n+m9ISZOWRyVTdCwlYf9PIv9nQTs50NTkDZwPgNAUlh+oAmW
XDCucNylag9R35XCPER/H89aOX/xtA+GZJ0irg0CBbtUs7c95GowWPq4kZvxqOnPsxHuiJpoYAvS
WXpSkiJEDd/RsCLvdOkocEPb4ydRx3Sre+6ZNuCMwmNQemhCjZjSELY5NSX2GKwElyAbhMo3XOZa
7dPq1BW9ZBLO2e8BEkVKtk8BN+jonJXxfoTXeTiRrixFNyPhb7lmZrSH/zdyWEk/00UCoCeMKdld
i9LdFp8hpEJLJy/rJOsUAfepPKNNzRKMb6/qOq4QdAx7TD0fQfhshg42mfHtD9xGSaBMksS3W58w
jerl9rHNjqn42uW4QmQGhpQ5obmHR8baY+mWojja7xmxDfprDfM0/lLW/u/2+gbT+iKpde98grU0
sz5GTlm7fQoxlZ4WER3KhpBspTUk8/3oHiCIio3ESXcbvixrNUA22V2KzW2IZ1EK/x6m1NCJOZKa
XMde5TJTAUPy4HlMrYqpPhixfVgC3nu/sJPO7qokiaOixINMIgma96Il9PlQvxAVCbMXJYEePsok
UXDD1C8aEaoxJROuSqrwZrsosvgRzWDzxo83t1+1lVnNu7+H7yTVV5WCUkuAxPr90WaTrdlgwTwp
NS9s2wFA9O5tcDeicKX5wvR4u99OnGI1RJdtpCs4hPdhSXhsckjfGar7sWafsMH6BvfcgG0JvwRj
N+aiDMH0YGjCV3qiCJ2gWKSBgWLJosxz1YwKvavXnqHyHkGLTZZHN5aw/5c2A3xx+fFNQ7Kuvpna
go+nriNq2emfHNlJQJ2d8/WgvRfcHvFfQaH9+zenDtRU+5Z3r2ISW0g8Ff9YKXtCwESEMBgtH9L5
+nfl5b8NkornsuofGfrd3xfRbZODzxNnAJrVW9KRxBVmAL9FTNmvdIywb/0CIsyOboml9zZGugX+
bIMa6aqrOmM8Wh1YvN6G9a/rMP1ir8pOQ98SxLsEVKt5upfLMpyBPjPC6GVqLV4gx5SzMN4B94h7
eDwLtTvNCWyPZ+9OquFlWvFDPXBjwFoa6qFAbxuzM+C81puzIG9yoS2WbRXgS+F2oxM4iILiotFT
LL+8aKnpBpYweR6cvmz/95jAEF/mWwQlz3z931hairmVwZ7wYgSTwzryLV5GHKdI1ZmHA8/i4elU
+n65ojDl+B/TkhL2gERhcxqIUuKRdnYwewMygNnEW44+H2TU/4p6Y8sMKrHvc2vJ9wMeEZQDx7PJ
KqORWNlAFi0Aa85BIsqfXnWOiVkBdUWRj+wOjLLkC/+XT61muRuw3aUD8FUrpfimMaZKXwZY+y/1
w2nkDIPsa4Iv/XPU8kXFDQN5rzJdHtmk/N8guC6lLOorRJLs6ovFjgXAcyq3mTBuxXG9vExytaZH
Ba8y2VJ5Uu3wzmz0fuZPhm9RfmhVePsOZivU/bKn3wJRJeDMnX/YhM1FbyHUbdxU3nm3dLUjkwsD
x4XguO1mb+up2w8erZ00KIb2MtZF3OJitsFYEK/JDPiWs+oolf8Nglf1ahlGvewE/4nXGbgIWac1
11F3GAyj739CbqGAlIb19aP8qGJxyAsy4wrNefxJOwfEipUy2lkrfOYYTEutnaudItTwhS2RSE47
curmOS9IO//KqBDCA34O5Oq2klrMb3kl2FwhU4rJKSt8/0kZB683EAimLHxtSOxKqJgSupyPPxMI
Jr78wQWx51zM7scZPZVSgvAgFO2MaLbxuUdxs1CTRVd8G4Ky0xRhGx9t7HekRLq1qfRwlol9dPwE
C59MT9cR30H3NYtmyb6Ujgj9Lrmq1rRQy3SKQ7JZlUzQhvxhy5bqGwcFQUPQwyfD3sRtlzKe3FgO
jmcD31sTJafb1GBMye45uEfO0RUzVMb5lUrDI9Y8LAWG726mhqjb7Z3Pj3HunzWdX/rlTi6hcy+y
F4TRorI1Wg/bApevEiQPdBHgDh7vHeLXyknKJnu3XFmznxpkUzKPystquYpYFV0ycG6JBNA3vHoT
rqIA2P3+cToPomM1PGFH1CXLQOqeKoaOfi3OrqnqbcasPA9LJYsHydy+T8s7JmcnNg2DRRK6Iw+p
hXg4KGfiMxK8Y6lEpBcRY6HPEVcqN/HqYgnPMEcgdIkDKBsq63hBzoYrz7EmncyNbm19SqJoSIgK
ucpsTjKtXTQ2AiIbwjO3SzKk36eE6f5uqGhdM5YG81Ib0zWmWYg70nFcy48FlnUv2SamBgJYIVaS
jIM+Qs/jDCcXJHfBVbEugzRb5S0sJFYlHsDTWnVg8MwyafFG4xqkDy3NRSEkMAZa6wGVGtJfmW1+
zrBh/8j1YLfN8TPfLtuEL1Z4+NY4Ef+sNkBJsvu3udTHY1GSfCB/yL3Lj3IWKu4V3ADaSfVTV07x
zCp1pLxnfagBPjyEGAF0gooIsuga2WGZnM53PAZ0rFy5NfEQnKwFLcLjcfVMXVer7cJ8UDtWl7Bt
fEk4m3VpyPH1P9IVVBTOOXYgKXbu9czdbkvbpuv299Pv7SJcfW+6OkiyePXEtUsWnwaon44zHtcn
4ARgwp0O7YVQPNenDmHNzKiMS9QqJad+es+vIh5RR2S/WLqEnA4jlNZRlR0IuCf3XEcyM+NF8tXx
9OJrarJGN1rNrU2mU8ptGzJlMiUCy7MjPiyB2htgLYSkc7a0UtUq4s0qKT81PGrdu6yP79epri29
Hw5i4YJxFw3vQksDD1W992ezlHYftR0DtX6LwM72ev3eX6OP/EWl1eJYCnDP9lzM6x3VXpU57l9d
st/87Uy6/jTY4EmrV4cDJx90Gd5nkedL1pD7POne/NjWRqoZXQ7Eug2aAZQnCIJrvHZrz//EWaTC
eT53fpsmp4PCO5X1YUmwxCL+FT5nobx4N1vU7/qvMZV37LcaMrU1VjMXQnnK7a55yRoJ+MBH5GIV
z2NK8bcEcsERyw7YbeLPKqLwsk9NQqoMMFHlH6QN7vCgHLGt6Q4Vuun9HK/gKc+x0l0QljmpKG7Q
i/bO2+QqZ6h+MW/ffKksNoEOG5/dNfkHf0IDq60B40ctPo01mav/kg+kMtwvSQ2L9+VbJESHo0tw
9nlv8bQn+0E7eSyU9HVUqQfZT1w4REHcZAQhbg84+iXjihw5v+8L5TdC62rpdkXfnJGiDI7ysAF+
p/vnRF+LA30JWptI95VXDZEFYOERPcfOj/sdTECuz0/InFkmyjqtBC0AAXLZrV6zKhcjYPl4j2xD
J9XDF9r0CQG1mOkIfLjABvkpvGVP8iBK6fE17no3ihcUlVJ9fvs+7gK90vRgLAgCBk+vGrlEoMaN
hnF+4xRCa+uNd9Ah9iHUkI8mIwYCGEbkJWaSDIPvPysoJHmMATQUCJr31UhBZkXo1ptmBnfhhzGw
jtS69FcwjAkH10csFa4K0LWj3og+MXJp4GojyJGowb7431ePaLOEBlwGS4tYr83H6WEb3dAXQqaE
XQhbiVqXG4P9Fcm+gp8VSFihqTx3KK2htiCuKxHpsianxqR0ykVWuAq+S84dseMc4VJaYDmMcNiH
NdbGn1Kcghzv+yWj+lefBw8pLscDKaxr1jMEWsiYpAUSr+SPbiLl7VrG4Escc2WWYc6484BnAReH
eSPk6k4vPJKux6mN0JWLCc/TjjGByJo+OlQMtIKKfPUt9CUOTRnFe/exY6x0cMmnqQbsmtK9YpTL
OT/3ffeeMACpqKP956k9Cu9aVM4jrjmwMwJ0mm3Jn+RsZbt+oJr04sL7CJ4QdTqd1UFMohMDGZbe
I/wtDAi74uzrwS8fPqLKr3H+F9jnlUD0hHa8dRZOpX4UcMmEj5ZEYlVYHqDLYF1ddiR2jKFpa9d6
AKCw+uJ+k3Tt0l0ff4LB6jDm59jhdD0LlD6grpHjfmc0+a/+LhfYc6Fygbu7n9bEq8zCwKevu+ye
Na73+aJY+A7Z1N8YHQ/lve1f9skqWWK6vA33k5hYx/eU7zEUHE5jF9BYXr9zdqQUAUchsm4kkjU1
x9K4+zZETROAXiofKCFHw/xQ9vrGSG0bFQgMeD23QLmyEXkCFdq9MikGXA1ZG+SzokTfEvKBqLrY
1MkFakxt8Q2sKRdlhSZFsu2jxitlOak88DYAzCMlKsYfkvIGzMbQSz2SCgMe8Kj/V4/WQV/kn3mb
B3cBJCTPNHUqtsubN2fdF3ugDlazq5fV0b19kbchoXt+cSC3xJiZ/3IGATjfLpIS4JSSF57TFvZi
b4MIShhLUf6AB+vPFznW4bZakcDWs9MlO2OdhwHClbuQZAUdpVJ4o9c37J6JR4sabpaKASVXMj4M
LXit0JRIpEXKiM7npdDN5HPB6P3IfYjShFavQ88jxJUI/Uz8rmPqd2Fci4lwxwDVLqF6j85XFrfX
/rJxC0PiCN7UYXJxPCaddD+1nKVyJYZc8zcJtBNDPcbEbmuLfIPhc1MCUF9+0D7l2Wiq8vQGM408
GzA3zkhzODwgWHxNtSbqFOUfcBgXbU/k6qX+yj9vIURiuJm+pxxirDHaPaOXLXKus6DssurExY31
fc6Oks6ti/egXzp2NNJmNbsX+l7XGfi5+63BRNU3IRcPT9+T/FTxwQBKwqUp8E4uuqYbX9RgPmuL
Z0KpiRMjvj/n2HeFnJXkN8UrBDjUMJyuoWWFz0T2GNsK7s/cygM3oYEGvk/efLLZSlhZJNpiigdw
AlW/3Xs8xvp+mehq/7YbGPU3TE52bZo/eDwmlcthnXrSdfUMWFxTGVQbcxfEW4ffIlfAVno=
`protect end_protected
