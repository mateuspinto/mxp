`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dBUXbtdJX0p3z0UrEnuTZ+kRaRHbmSDsFJvi1sQAFhfq9jxfxGedb7dXDnG+khoEIUOb3LowtlXD
HDE7q2k7crDVgmoD7zvbVuVq54WT9VOZyKxz1sKY0MlFC3zlJ3f7iNGJbcgzFf9Dk+4gm1HJzZng
GPOrcdVgZyrzvzqAaW11CCBVKG1YTWCHg2o4LopAQpAAu0DQRGR2cbqV97SQSYIRTD7l3s+UIp/k
6OR0mpgjS9CzD0ll+cFLZlcjgR/wKttGi28zPawdGtdFiMyurY5WSGsoGnZhZ3ndWrMLYyuPJfzJ
942VDyitaWPbs+zg6h2kue6Wl3J/7+BDn8F/vw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="B9Ei6vBQJHYpIz86MlXNqloh0NB2lM4J2CBwApzS8vM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8992)
`protect data_block
us9fgN9xFLYFficxbNb9DGgbm28g1qJh/eumx5gmxwFMp30GZrECWg/DJR9dZ8sNFz0mWR+zozih
4IcPW9OCpfaMbUeu778I+0oPn9a/yZpN21WIaUpqlKbbNo56Yn0a8e0r600Mi6bn85WbbSr4uJWI
mbI8gSpJ+CXZLN29rwwgOaAT/7elTm04FsGdRZV4tCHsbszOfUAlpEvAFHAssPMU/m6hpk4Zv0rB
He8LSRaiYoHK/jPeRXlbWxDpKyo6jVJZcIN/suruQJRD2WEhuXWt4n8KmEjhcvSxXfNT5yNBRAgH
UFhbwjaLk16Bw9yWbFGkPMan2e7ZYPejHmcZJzDiCVFl68PblWFHwOB+I152oDzWYTPfOj3Ju/Rk
JGUfgWl5FMmhs4JUiWmVGJ2uePHgKJNijSJLe6YzPpgFU7jSnMkGrFZYWAugm3yRZ3yKD03KtNJf
ISmXPW1iLR+e1a1p+7gHw12teDnv0XhXKtTPheB5w3ykR65MtU2RaAXunK24cd5WPxiaVxRv6Tvk
D3kMNgQVMGYrO7i1Qz3DgJl1ZPy1ngXdSI+yGaz4gshZucWNTPrpqz8ZkOffuxYRKMl91NmRoqCA
YWVgikeFJ3v5N1xMdsbZVzkaS7+vv/A9hlZGrG/B9o+350CQ0Z3jUpw/6dB8wMNZztDcr/D25jEL
XIxzPHIQA/zcXqoPUkDV5Rw2GcNEtE/6cW+yAWveM+OsYrZqmNvkDTCikb/aaLtFhOCMPpD8e3hN
d9C2W4w/Izb3LE3JzRvPetkd7Poq3Z4tb5+ucdGHpWtmOM/WsmYx+is9r6vg0ELJzh08jf70LQux
kaqnw0eaihJFouaBJdRMKJinm9FIB2jV/4B1uUuA/UHERw/66yiuUdVIwj1OvMY62mt5m4GD5EPE
+X15yuPNmLIe1ffUr3mlmPbPYnB55g792VgqRSGle7deA/I83VOjpIFp4vT6OY8leppd92Lj/x6d
xM4ZQW0Zlm1/hkNoUmYgFJLoRvokIUFsUWz45p/vj/9nmn7oC+YBz3gAzxHU8fr6Zn9odwqqxEBr
u6yqfQW1pwy2PAY+49u3id2fQ3AI0+l9V3IGiq6F2EQ2Z8D/qkwvNsBn3NzoeuMe5rWjDOWqzJbH
nfe+H+gJ4yEwbTZETscGr8mR4Va0DPimvGnOW/1WRqRHnu+PYxQo6/VqMyXJDOJpUZwelHp49zRB
TQ1yEbZr9GhbzHanO3n1RU8MVlh418UGth/8r3lw0hzP+3DcBxE7OLA1TVRJL2fZfADVhEwEY7fQ
t3atSEEOG3KU+5lD6Yn+ioGDCoCLjDH36uGJCUWn+qHg7x8M4UGTL8+3gHdmDfIYKhXIuBYLznPG
UXV70GDpgsKY73WajOia1sE6PXjpbOV7rZDTLZpip7TseOPoSSE4ChsYfS25fgB5BUGJl480DV2r
CHZ4T9l386m4WBysA29YhCriRvDn+j6PoZszZItMvbyf1K5dynpATInsLEKxvTcXLu7NKmn0kUnQ
mLvhFGR1C82ZG9bWLHebGmWQDhScOuD9Q+ou2kntErAbxWC/4xPxTBJ8lY9NR+NsNTgHW8lsumN0
EklF6IFZCcSeXzqnasQPKBsyv/40dyaA5PvyApVyxT9AvIwCvUHMXsme6eXzX2R6LeBnB6Pk5mqK
uZVcNN1DMrwE9NGNYHpKBGirIYziJzGDr2yCIH7jX1F9Dxy5FCmDqbyLzkqXcqyiZbe/JgXsHZ+n
z7kG9ee5CSKLKyROx4LkPTep7gQsPO6Ob5n/MXYd7kSjWZlMwafeW8d5jej5JhT6zN1ynDzjHvJX
1WdmjGVrSeoAcnCS1X1FohnB2kTfTHWEVTKvVzKPLV0KpU5ogSbqfuVGUIwMeG//yrZdGznWSPnM
090BQlLrnbh+wf3eTshS/OvJWUJTQDFQm/Yi+867E+x5jZ51XZh5Tc3lqa56ItF0g3mnYcrfQnNZ
5FP0vf9mxUsHsDbWB9gZP57GewLSdNMAwojC8dGCxzKAB4iz9UzU8lf2GU1Eb/oJWZ0/pwVQq4zQ
W6wXj8w6No03dS1/0vFQpbNuBARVsH/94xFXsMGgStgExj5Yys1XZq45EwUvZ2T85R7c3fROm4du
UO+92kMSryiQ0NWw3sJrwjyxHNipFcTohqWNPDFwrkNWt7yOJ3yIxowcnWUp5zD3GKWMPsX085AH
gRjmDPYiwOx1/LBfKayGSJJdshUSA6mMLHsIxGcZ08Tpgkp+6PllVwyenbsXNOM6aLaU4/OVSdHi
47Z+kle3Yt+33SSXE0kb3Z4du8rEKQlyVZCrJWTDzNcltqDQ3TuCS2/sbAJ6Hyrn1pb/AVqEVHiK
I7f6GjBjEqxOdd+PARkRiAJnNCRiFofwNBBL+kATAYyyCzQoFLC1weBSLpipRx0prFUSfVBr3iqX
FZadBBXX91Xe6zfud2MvM2EZGN0mGjrLtOz5X7QSubP3bKzija15ni1nrNRxL04Blo8cQGFNw3Pg
2b/ZSqcqJbc4JqyirXyZl4xy3A6eUwl/92VJD7oWuX43Ke19mx+eZ6VV4KBT+bXpgxJviCWmFW2j
1gf63m72uqJDxzyTsPcMl96hhPHutfjFtOJrC0An8GAeScKIG7z8Mo6IN5BdYG3j+sxH7Fqadd/5
ykWNPfrxsKcqckx70xaLsGzBrcQEgL5vuP30TAdNPfXTa/oTZ3Qc3upJ9CZojf4IiHxUZIUEm67P
dW4tDqAaVYUz/XOxq9kZW+vwQd12s/gyDODTP6wHWVIPdhDURMF5e2ra5Nvazf0gU3RsjPWZcOfO
SDeYmYLC97JFkhvPQ5Zs4mx5v0BlrzMZsCA0blU16wgi1lLv4ga+gEd90ysCEWN38l1ON9Vm0iez
X56X3uVGpOHCbUv/TkgyKKQSKz8qV5afKHsIoFrn/yhnNBRmTd9yWXhjzSycHUH0YCfKwnebUy0t
7cFyz1MP8gF/YBIvZKTHBiyRJGPQTNDMvRpAeIm348T8FNbqGPRObcnw+eLF90QWkXYlXLm0P8CB
LyUDjbtFiWkKL6tAnYST6lx1eF+jQwSyC9D5VD3GlEWIDMjm7SShsK1CsHK8EicT2khArQOPCapu
m1a4l2grNoZs7N3FnVoTulcsy7+ix4nZTfsq4RtyEPNxuYrubKtx0VWdO8M3rbUdb3DZIx7aPM4/
EmQ73K1yA5MLtXh90Xx62t8RJhevV8/LC6pLRcgqGOOhd0n2XAuysMU+vsZzaGogsGdMY6OWhhkt
7FQq0jX254+2SrVyjjAa5eAg7A0lYpq6/MUQZn4D3qS7Wb7r2B0vGfCxRij/lW0D0jQv62+opZw1
raLyDQvycrV5Pual8MM9HE53hgHny9wER1SAGW4pAIYUW2ntumUvMeeDyoBb28y/rnYmwliFONEa
o012hHZigz1L0LDik08Z5oJfMSRl5J59r3Rdz+04lTvzOsfGChIaRhFc21SZpw+ma6lUZVinOLrz
GPYTJSnNWkF5NgEhQh6iFMx0enhLB3L93kDDmvrZCTqnmNWAYZpM80FXtHkvAX/Ct/8LftTbwcQs
x1P9sweQtYpb44UdLSxF3Oo+1KTbVry0nvHwA+KwbtqpsfzUP8UtkIG8IQqAUm7eSTJIY3TEvlL1
HeJG4VGWiSkOc+n3la2a9rNT260Hgz9Cz/yNbGBKDxzae+AJpxIKawRD2k8G3+69yVTj1FKT4SpG
mzSZjI8W3kYbccEHNjTWRURlAYpH2dvB6QT9+m6y08Xq2XpQ7H+6GYCYyBMLkZvoQ+lrqbxYmWgb
tI6sFqZif96ASy1efPu/+9DC7VJ0ZEPs3AAKrEFXPp+YN2vj5Hy0p37TW7PI9d4JN9rKrbKQQ0qK
Xd+DV4yQjBDITQhnSbfrdyvAB0/x7JXXWAtKQS727FHKw9hWW8GPmFsew987naFcQ6zchTIFl2AS
ccv4glqXXD5Vni66+xeQ2ngEsW1JBfJdunjIgKMMHu4FWvsKt50X7jJBAtRiu74AuYWc2vHrqHAt
zXxcqrUq2lJQj8gusHThK/XoNrrUh3MSIb6+OgmNClkLy926LmmBf1WO9BJJcEHTv2jBbq/zDgoR
OYaRUIre/RgCnXeT1pV4826O12qet7wiMFn4Jx95LodwoXEe1XIyuN8xCizhAzbewAhdNi9QYnlG
NyuI+YCtJw9sz9V6ITSUatUrxiLPJ2lIRjwMPMzyWg0YlH9JazDFb6FSwB2QXKe5oUE8eZFRr0IS
OGssxlhGt1A3euikJF0KF6oracfGUGeT0hQ8Mat0gdWGJhikwZiRhSIT00I+pT6NXGUzUiN1eSuR
rW8yRtoN+thpexvnpbryYD/AcapSWeBr+CQckLBPDaE9YtK259fwNtpr4TWbIMJUL+A7M1gw+qRg
WXQIvXAHFulpt2IuCjPMtsv9QvBtJi/uLI1Sku9cOfg5DesSLl26bxgdtURwjQHsCZOiCWa7mPjz
sfWjy6pS7cO2/ZzPoqT/dOJeb3ShociJYOJ/WB9DKSZx8awJQBea8g+GS1dWFvJM/uVSb4pUVRWH
7+DKeXUU2blhyGpYPhMFbgOHS4oO2swz8YclNdqO0idPHMK9CnqPjCM/qSQUdMATZoeurrBy4+nP
iBIPexZQlM7yLLaU57aTLzAQGv2mQFBPamy9VL3U5OdsMnv+YvlseHRe8ukW+XMYWO4JzGNH45Go
GXHLLdRFFycC8tzMpZSTKeLRc1OYYpMjB/n7S5xWxyQgCqRDQka1SWvgmOyFuOnyZq8B3UBn0RnO
7IxmBpF4fSlQpe8Y5JllMTEjtoc18gKtNNW02478tnQqjUx+49yoD6MfDHkIoStit1tCVFL0JR4d
68tdmyQcB5q05190+/r+BcJDFdi3dGcO5vrU6bVT4V0G8NiLE3qZNI6r2yi7FMAqTYP1bRd9et4k
O630hK+hmeNHiAMw2jFnFXqHH/r9n38nPwjevSuDycbIbqCSJzNSuNN5da199kLBVplPqOuHAlP6
L20hSr9Y19ziGBaxPcvmrcANqxa4q+hdaKypPCjOlVRCid/5Fk1RQkDn5gK3HAYMqYlsPuJ4hkeW
ykSZtPiiVsGc97RgBcIcBP9Y58A2WuGkoFKSqSRHa49mxYcCmObcDszuYJZlvqA9o5g/XNGaS5d3
pxq/mJ8BrFmvZYApGv5V37jE4X2op+Cb8qSMLzq+52q9t4Whu1ZKmjpECrZMLu+W1eMqTLeoCbAP
3hceyrvNzxstCsNTHJzU9TVJowyi2lqKAoUs/JIW/2/wdsv1IYhivr6lZrtEjYhIa8sKsK1+R4Cr
1kMCKvRZSeVjoYnRqM3smvOm8bC6o9g7c9lRYlZK3bI6TR0GwCHTtzGb+5dHprwzphZt6o5zUW+s
2ykxgrhYB7CU6H58xQP71AeEi3KntEgrz4jkK2KSw3sq53R1he9FFbLQYOeIZ8vK3efnl7WB6XQG
YWTMjzRDVLaZb7qWg5VZoq1wJSPs+/meW6K/1UK+FAsvgbH6ZC1J2APqvnFPVOiqNRJe1w9KUHsV
MFziyccP9/9bu4Acuen8UEG9uwKyap+b5H3dpfJYw5+ns+cALQDyl+XvrcCQbBrEf2VRg54FkjDk
rn+Ci3Zk9oMaHBmoQMiB8auMwQXBx/HaC1jqE6amcxYB7onWFquaMMt5t4ZohB3ZpI+BQibJ3W2d
8poNpiAXJ3y1eljzBh2F0pKCUzj4aXbltQv0/6A4XR5yZAx4wE4ZvzAQLTvXU+tb3x8lT1x0lQX9
1E5Go5A/dY6FWBpUZugmg2lZhaglUx2LFHnVqjjG7X0ltdeSJPnxcY3oP8lZHmBB+nxahCzIZ7xD
SjOQ7Isx5K1fTyVNkKD/CutEVIZDW1EofAXWvVsjX98ZaWtBOY6mE4SrOuIVluRo0/L0hId59x9k
3e0/L5WQj4VF0uIMhKLtaBWpQJJq4qtnSdz1785Lc/JGBg0gFwyaP/yurJCHFo9acFOJu/LLlR4f
tsWEQHvNOXUlmudlXHkJ/dT77GlNKL9HDbyeLB0D7BB5p/2By39SCE5atHigkciwD3fwxFlDLFId
3a3Yfyys5QWlX8Kqx+gdUzmQy48PLRUJXjMNV0waZnBGcNe078Czi+sy6se3/p1XBHNFf8ZrxTQ3
22qx2jhvlPEhOGERbiIQrNZMSv1cIli0O5HYoN0+ousrF4wLSbhccma91sb1zFgPgcqTsEcoRVvp
uDQjeDiKGlmlRzDUILLbZ4cPYUckwnEn7IV7T6Oh9sRnWhYU3fAMizdYZd7lXfhoceuQEhTR75Ds
93qTkJyGTr5LQSUn234b5qzaPthaV0Q9kmWLEV/MduRRMkMJ+EQvk0Oi8SYqsfMMYTMhPWfijxvF
Puc5czbW8gJF065zX6lL+wrQ4CvRrQRawgFtN6hIpiZDg134Q9iVXf4cIZtKHxd5WWBAUAwdr0wt
B8EEI2NFg3SK/Dnhfqg7IV2nPgXH+xJhl1GFn82MvFT3gC3doWsu+pfeGxnS8XQMMD4yCazwokkj
lUNtn5G3yXz8p0jZYzI6BzQ1rKAQ4LsinykO9zqZe6JsWSw0+c1WPQbsZGMcvowhb9/ME3ePJpRL
zcs/OyoEHF2kd9DUCAeNnr/McsffL3MY02kY2FeuwP2WW5V4BToinp0/mvsnPXy0SrpvwwUAnCJK
BQFyHOzXx7A7C8VbhooRW98RMRoUuIDAgj16iXaWNSnjjIaL0l5qKMYCndWWSKP2fxuCXaW6oZ8c
2bWr+Ga6JsQg1ix+LjV1l6FvoKvCtQAlPg0uVxxhLYWhZz+Qgf0PjZLOsLdI7oleqrzWhfQmyG1l
zEtEAqq7PC3bR+Rtrfi5Yk1qfb1vkNLDK1GDgmU86K+vivHS2IxR5bOS6WdohI2LcShzWX4WCbyk
86582LK8T3LVopND1pTIr8O+vwpVuu1upZw82lclmBbI70A22R2dQVODtI9j08rkIQGNRL/Ya70F
09+M3aSruaE/MBAejCDuQYxwNavkFnhkHC/LvY2PZ2J2lM0Hkrvfbx4d0cE1xjpBaeRw3xUe0ga2
xVTD5w5d7uvFMrj1mYGoJkJJrxPpKojnKpPzU5jBt8LHCXD95lxHEVHAYeR4KfMUZ/fQaWpDWf6D
F3zAP1RhSluxASVnemSJRshW4vMWqZyT8gpeBAP89IUTJUb24zSDf3kqzleHF24UyPqnWCHnuUv2
aeD0/rznqd4IYbSWXGgxSsGqesgtD5r18O2R0+fKSl396eFciyFEfDVQnBWKJ3v+GmgGBelnSuNY
koYzYhKn+EDundp09AMLThNkzRiIU/u5arX3JsjwkgHvCoasHkJb2KLKHlpVZeIPO0NnUDfUxRfg
ml9V2AHx/ILNlSQNOaAfVu68V/N/u2NfJj0fmW2q0HztlVlBuBD2ok6362540TSN8PAV77zGgXEa
Sbo3oF0ZsphHEPoyw+rrwzhdCj47U9Qb6SEedLAtm1IXWaEeX3/oEzFKa6E9Znk1klxsnkG6MIbi
sGt4qQd/B5wpimC8BGKqFGJhZBbdkZYQbA6smYRmKlO5OmnBMm+V7B2X9zrf+Ca/eo+KtF3aG3Z2
Hf6/MWBev59QzNrWfOeJx55v6zRQuyJ/BFn+nDsfINT8ZHDRNYYNdCqFla281CeVYTxrrRFObn9h
s4vXoExHMo14/nVSgbUNoIOoPn5XEbSQ1xXLkBz47BCvRwFr1h5vAJiXwFnMQBUVAHjDaZAvknBI
gERecZwVCDkmQCKVHnNoAlGb54BbzpmGsCfqOdC7x5Rt3zQr4eaD34THMapfjuBlqG59NX89kdbX
sdcNQqgB+YDHOn15LTLbfxXxPti++Caklhy7iMQjxGUVgEY6n4d4eWwoRDs+L1WJRkl1KIvk5fkK
q8MXn3vtkYaPSN2io/xOk4Z7mwiKgu6LEp6nPWjvOBfhOKFLEszuovKDQUpRR3D8vVv2LRfMHWJM
MsUOaEEiV7i06SyUA+XgW9R+eGwcO4in9GvwoKuT8BV3DzZ0yNWbMjerjUg++BQwEtNkm+wtkLKL
RCN3hMp+HhvtTwIIycGcSZlkIGgHMjMgwFz1EGW8m6umN2jKqVNVOqJ4KU9yOqErlTQxjDl59/xb
syv/eNBUjZRBiPIoQ6iPozgbqRjEUw3DUDtgB+yrcejYgr8v43GPxLL5gZcmNPQj0npQwAjte7pk
DYZh+teFI6+cOpdSzF0+VfxgYVo0QI9mZi46lDs0fKdxKX0Wmbv39tMZuMAxAp6D9mTM9DsZVgk8
rsjvUi0VWLAvuqYYzVAk7EMJT5attq69nwq1UEFGLZlcdy/GfqAKxK0nk4SK8PDjc3yx2ufOaRhQ
Ft08iMvI/QLzIqBFW/Uy51rxz2GwgIqgZuvIv3Sn9v3yon6fdkVbckP6VGesofbjQP21hbm5aZnj
aS9yIYPBMSokA0QfMR9nqWirZXJB99K+5nAbhhWdE/O2xrsZg4Lq2XvyXGl/EsIa2J8yN05tbP5n
xhLwgKtcbzz6S1t9UiDYFcjX2U1AtuGSxDyYyGUCUv7rugqLu1ZiRlUAYK9zdTbtT4iRw9nqOEVm
AzgIJL21Q942dn1mbr0jEaLGYMM++m6o8L18oWEGHT/coKJw1bBum2lzOkksp5nZjKvG9rX3qsZz
W0r9einNgULnRzrBUSUaVS3Ie2kJf0oeSUruSjIlzh8CMdteEWzCfPhsjlptM6WE2gU44P1jbq0e
AQagtqclF6DdexyoOdSAwTVo3bS3BQJAYyT1EClBVSMklbdMVrNXskOF3dMbWG45QOYTdN0cSN8U
UfbBK2QcCbzrcT/Ud3KRE5K9kXXCs0gJ9+Wn9oCc8plNxGxVfaU+foFYMsusSab45KggRj5etm1J
2DVi+z3rAmwh+4rfCSFCq53YgL0A69Nt+eUPJHbdJygtUQ6Xez3rE9/DSALNXoQZiwDx38oaOXMl
3fSCYAlgWdvDgOkiC1p5hvDMII9eoqLqsq39+WFu8EZ50cPo4Cw9DzBPnNFeMiJPjpJIiDltKton
lnCNLl2r7xKvZFZQ8ng6q+DN6oJAb9GWqAwgH0Hzo0eZ3sXLXQmpBDeUIR8O3dUqQGfATRJMZouq
vax2CmCJgx53UbZXsTlBiPfQYPCds6OyK3+s5md9ABXTV2dOVsSm60NchuF/4df9c95+DsBsmQFo
qTaVfejd/GT9qm8QC9dhyJXmVw/Yn1ZA6kdzqo4EuiUF5SxU7UwI1TprrA/GurGi1zMT8WcnF1RZ
pZAkWxlFRRMwH+UgxbUmAeNerTjPQg5XgC1NH848Py/TlQZQFaD98EMKxm+9Ggi75CcpOpoCJ6u/
tLxeAHGL2MWp4YPLVlt608M5+ICdmZB5Y+eGSJYIfAf5OYxNxvRhNsYWk9r+ayHF3+Ncu113tG8x
bUf53BY86dNzyMXmi1C16cPZ851I0LjzwanwnrjMRc2FjWiPJrHq/O8Hm18aVZw77VlEarIEQMvF
E53ybZWCYAqtf1mLDd1BxUZmO9DThPtPdbhKzsJrukEyReCOes8xt9rkAIBn9sQi8lHxjZpqWQI1
XNADFZJYCuMNZfPnhHUxDdjY4XqbLZTdlrBV/mDLsSjHOgOLwxv55qiVeOUML+yxND50CMF9ra0Q
GVNsdlslIGU1zPbInTMf7VzJbqpg1Huw9XEegMKHPXxcG5PAvWH5Rbcw2AxV7B4B5leGnwyN6TnI
PATBkitfY2RtsOaCkkV85rzJ/LsU/WSfOhslg3eW+JvDxe/IdZXIRTCG+EGhmTcjKGgjvX7pLrRr
afLKpJjU1h45wf8jLCoYgl6V66zXphzmZQON+5rvGfyciVIhXW0wNvSJUQA+wMCB0cWdpUZWuvsU
R3VZDh0USt3iVkuOSHRnOA4UQDtXUwBNlAUwWZtrxTYDqDBPFTbYlgcCkvrQ5TIOFG/1wOwv0RXs
vgeE3RGZmDvCU7cjeNNtYWdbRiZ+khoH/bajkQ/iqLDHHuvi+QhADe3rHMEkFPkeZY5O9MENSaj/
A+IkcPO79HG83Nzibd/4Mke3rip+DjIw5tEOz3P8humNDTPvIe5Gcla5MzakmKdVJ5sYzWF/pzNU
CvEJaIQamFxkjKlcOEiQME0/CY8ES8I7QymT7JOQGWjqNIBB5jKrvmL+a90NtkrQUemDjElIH7Ht
jGC2GkjTaR1TQ1FqYwmi6wSSVQL4obh2nPcitZyEj9abglOUodqhUw43/UeYR6owwQza8Hmlf2Pv
RNO1/69T0CNctF+79qEhcCJh/g9iwF850z7E3sHlilAcb1BAkpcYJPE1jksUnSEJ5wC6Dcb+TorR
o+GlFwnl0WrLhCKYSJ0Sfq6piRqCfm7UtrrdkRX1sNd/HoDrBDXr86I4WJjvyMiz2J+6jcN71Kkx
BXfj0GMHoi2NfLb62StdevkVLAulnXbY4Hozjz0egdBml9qt8qP/vmE92LG3IeHEsG6Xqh2eT0Vf
I79Ml/8KLEss2MHx9kB7cxWGX13vbd7r2MpCE+DUmNA9bk+Wr9OFO/E2PmP/HJh5eSrcz16Z8ZNW
fXM2FloeMoFCngdmr9gLt1R1O1HAf6JT0woWXaCS/yvWoJJbd8FZrkkAbHKAHP7YZgt1p2uc2fcT
8Jjl17eqEw6l90ViZOHmH34uaJVoTjmLcYmtmJVmAw0ftsSR7M++R03w2wGA0GfMX9bwCqtVOe/T
ob9t2zzkBpGM6rvQSf/3a/bsI4nHl1eIvjFlnlCs8RhC8AU68ThJHAm++G1AcHBaWsDzYUNLiMaf
aKcmUsPw0Ma+k/Gkh9e2JF1H+L6HNG6bwGddZcaH+K5CmcLmECasA4p6vpbCtE9iFp/DWWRrFjvs
oCXzShGOBm+5l92hGUp3ghyYWw5uMApCDbxnTo+nIZTpe+Yd8E22LhTFTMvqc+zb2S+AW8X3deWt
fyoBRMGgQe4B0dZAEyRNxXtELNRMobxIO5Uz2LMPrQK7zZSkZyP+WQMtpInFnIz6APeaL+pqKY2J
oZxSbIVHhH+1Ae4HNdUHS5s5GT5q9p9uZyIgk0BnVjDbWzzU73mh7DdpjWQEZQPEMNHH94PneSKs
Ap0YrW4KHJ6EDMd/+8p2qLOJEMOEIDdC+MoSsyjSgc3LMcbcr6Y3+gapPLYYVC63ZUAGckS4ONAG
U0wlOHT6SqwC6zo9wNmzpLUxKRAGDa/Lp17nt9Z3FxQCtbckXSxzMgVKTNadObFbiueu/DTjyBU4
hiS7wnmlWh3MokPPPaerUviUSdaJ+ULMoUIF5UlasdQmJP3bPch2RUfhLYf/H3oWrj9yWROqe1sF
npPT7m/DPm2OzSLmaGZCwTMLZUwFqXRfiIdIQldIid26Avvh96qzq/v2PFPUCOAdfSTRKmswjt51
Esvp977d79S/aOIj6dwTFiFaU8TVT4LRn00mon00rKE7leDcyPuxvccIQQM9f2gVTUVpA8NH5FLj
GY1Z9QqAG8quvtxG3vrDIUL6wxYCbRlrZMCjkM89O6YxmXrPaZPcaTjjs+fOhk94pI8RiAiH86E4
Snq0JS+szNjH8Sd9n5r5YYjbFXPCxuMvFexD/o03Ad2ZEPOQ/NygFwcRJnKCgod5PBWiAofs0G7M
4j2g0xoUwNFyk0o1CBej4K7k/Ff5sUZmFpASdhcW7nS56tNoL1U4Hj3yTjBALATE2JlAZyoIiBY2
iQazYFyw8bLce+z/r3Dg6Rjxy7aK4ttkFB3fvur5K0cX+W6a9iGLtepOUWHlOMKzfHIz7smQ7CsZ
sU1oTj29ZzzZIvTZYhXmSdIBOESY/Y1CowMS3jdafkjGaCIMHMCVBiDxpPY255ZhnD1FKvy8qoMW
WR0P/oqr90ioEDlAGxeCfL0djzoB4HGEyv8kksTdFmoRHfGcImbzFKsxIEgKfYPv2JX5Gt4/Fgrl
HUWSbphmizn5oKSfxN43vyuLi5uMNglAdTMcaMwU8DJM8IFSVc+68YsWYg==
`protect end_protected
