XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)�������3��TE�y�GtbSc����Z����֏��\B]O����m1_`N<kt�۸\��`c�J=��$��d�f|<u�gI����;g����i28�˻�աb��� U�����Q���~(�(Hf8��7��9�z����ױ�j\�.�DQ.*��9�"�E�4g<9����ՃΠ��~���ۜ�*��-��㤰���0L�݃�J�@Z�j�i�����
Jg��Uu�.w�GΑ�`�.v��% q�Y�!Bk2��i��5�+�?�.��uܸ���B¤>�
�:%D*��T?@Xר���z��nB/�՞�X�u-��;�p㛟�_���n�c�Ў�$��(�)���]��!�oTX �lǝ�d�����7�?��K�o���}�[��3��������v��e����@V�6�<��Ԁ�I>g]!iX|n�jR�}+��$[@����G��������Q��8J��G���&y��!�ۙ�K��LpAtv!���䴕�1̤��9�u���Ŝ��/��!��S�^KC�-��\R��v�v�v�qk������.#;ծ�Ӌ��S��&�Wj���聫�Tg�2}�-���&�J�n��˸��`_uf����公��Nrt�^�7�KD���p��Ų�z��a��y�5�XMeg�)M�m4�����N��i�ҵ2{h%����w����̛�i��|(ǀs�Tx_�J��L���º�*��Z#jD0�l-ܠ��&�|����@�Ll*�7��_JXlxVHYEB     400     1a0L��Et�Y}g�B�_RVY WglދoQ�_8�ZYD�X��8&�/�:%�gx�[����w��)j�VT:�-�b���Z�s��F�4�u�J��S[*�7ͦ����i,V�J�%�ړ&ؐ��O�I�i�Sϖ�I��X�L�,o�A7y'-���.��yrm:���Y�]�(� "��L��"Ȯ�GGQ���jDmdӁ�![=�8�u��;�]�����8҂��k�#��B�_��}� �c��#�	xxMϡA�jSVď@���������W��ݨ�5z��g�����1�{�k=���1o�H��I��5Yd����w.#`L6B%��!�����>ҦwWc�
yWu �Ea3G.�,/���+�z ��p�{pjx�̏89&�i��-�d��F��P�{Q��'�AjM�C�XlxVHYEB     400     1b0�Bɋ�Bh]�ɠdT����"?��1��}]�g	*�}�E$"$�s��4��y`m���}K�8�jU�]���)G���1���Bb������]'F����a?�Ù��L�0���������i:��jm��uj�I���o�5�c绑�ΐ���f� ��(�C��u�G�{ڲ'��_��A=�x�c_˺�Ad�����߭5w1���VL}�:�L�D?mz�Nȿ��mt�=�{탕"z�^��&����p��~��GE�Ϸ�u���~�/�U�u�z!��n�*�Ngv
^�����l�R��GC�Aad#�p"���Č�Nu���dvG��7`�`�}�yUCS���n�M�ϭ�ϱ��q����£���n�v���%�5����|��/��T�ʺ��Z�a
���ՆªF�ήiϬ�B�u�!򏰇>�XlxVHYEB     3f5     130yiEۚ����I��2.�Zo�|� h?�e��c����  c�>��]�)��c/F���X�O�:vj{�`e*{��0��C{�`�5�y�1|v5T�<�׳�Yx���e��|O���K鼛�&3+�����_�u��u�{O�,}�7�uU��z�_��@q�˱����Pa�%lܮ:����H y���WQǯӻ	2�$$GF��lW���{��9�(��{�0�y=�B�q7�^ˣ�<$+��l��,�8�_���:�I���1�#�~?��&������[2Lr�0��Z��wX�שq