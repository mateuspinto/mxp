`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
2nV0vAA1G/ekmidFYzmVA8E0S4HI4FlLt1RP1mfhxH+3J/XfQGiP9jZ8gQJSWAGGsE4heFKMM357
o7I+mPVVYajn7Fys5mK3BZ4wO6WvuDJ8zf2wytipHtV5fAiF0PkPLbJ3qfmJg+iit4ZvbxT7oKfM
+1MhbgNmU7TvauDTPc5PBCCJNOVBF4j07wwwZy7w2NsFnxYX5lEuTLxb4UHaQrnXKhzS2DYeiVwD
TSb09GJoYOSlM9chzQrPKOp9F/u62rEVyHpIAim7rCdcHKiNqPG1yTq7bn5Y3xDLMFM33tEulN+X
hlh/z8mX/gpTCRYSV1a9fPAHMCADsuG9rPB43BmGJswl0eCR79yniAjyOiRBAMcn/XGziHvptKi3
GjNy+jsh5LAqxoAiVB+MUKy6a/UgXakKtFO/QSJBEY/reb9h0m2ub22oQ/haFAyepdHwwKb7oUTr
0fBafVQj1i8FUHOid+0gNDA5TZSbNK+GknyEZFjpzoInTwkD/z34F7cofq8nkT4qRKKLX6fJF4fj
xQCUrshU98Zfns9cURcvdI52geD3tD1786Fr04kEUhNUTFgel5YyLZB349olvdTkinWVeHTpWUk3
uiVZ6jLFEAstF2CKrcNjPBXRVT8qbQAAgblBCnVbuqtf5ViRVyHItNbtkkyIqQbbeJ8pTXVIOXdK
556KefVrrpUEpKm1DsyBAu6WJ5/W4eG9IJfpIr6LOdvXh1zKxoELLpBcG4e556j5anasEu+ghXkd
sr/iK9zEC/LNALyhOgRbcadP2hqfbihlJWQVrDKVswBeKpp1/n8L4OqK9oHIP09v54X/xMY6n0gN
Hsjt3iuXOHQPSz6/3L5MrcbDr5FywkKaCzpfeSZMZR3bVIMnwjJUv5u5okHEFMTBiuQtBIhPo6iX
Xotr+AOfW+7dux6ommP2zlCPiYE6LYDNVZLSfqUpR5t/QF8qYLmZOwYiA+GOVE84tG1hEPC47z9I
TEbx7R3pmvx8zYsBMP4SPtZCrhKslkuMR2xqbS+v5JaWzYjdYTreY98NZB4aWlS9hg96M+uAxACA
rKxR5t/Jz4Wi80+OHfYMx4+rg3y5JylCSKSiqpsxgbVG9te3u09NdltEQb4qGcfnng0bn+VB23DC
e+L1ys+Dnw9mYaw52adRAB2tCbUxOeFctJug5dUJZ8jC6WxMzL3acxdgXvi/P2oBm2OZP+OQxFI6
MtNGWDOEL/FtOLv+8qZ7qQUoKwwoDeLehRNSYLkkTpid0TAuD+o8rbyYhbV9Et7O9HGw2GJossba
q7CCHXBRIKbkhXDPF85d3yHMnCPJQp0Nu5GDy1QAV2xOLRj04xJYlQr9YDlSOY6unushEV/xzJzM
a/xebfPe5CPuwLrwuq6f+XzzZZ+ur96Pi8mo/NdD8A2/OdNtukngxHRXomCwfWhmN2fP+2jGX0oY
bArqht+6/8yepbpxFlsYgcnMwpFKjVEpW9FHFzEgBmOFRYtINbQ7nyM7o+Wi6EMVV3c+kNFifAF6
P3zz8aFDCsWgPxMYVJ/QCdtRYY5Is2VbXelcvMwG6nVNgs1Vqovg9pdyH6nTuV7L4C6JM07AIEFH
xdo4N4nwsgAQy6NeBNLEJpEg+Fk+tuX4kWHD/cc+Nrajl385zx9Rk0E2oczi8xrkbwUxCg09vo8N
TkC7K1oanYjML8h+Qn6qwQ3VCRXaZmCq+O8yWagNV0wixiqH0StsTgTpudEgU/n+eZSo5wuE9uAD
RnyNypB14lZwNSJKs3ld+BHIHw2pWbgrjgZ1G4Gh6Wlf6aPwdXhnnKnmFq4PpxURrFPNZHmwEb/r
K9JsIjSbPWas5KYbHscAzDFT95UwxngGi2TFCfTR22oT8La7QwhsRSoWeyOjtCTe0MUiFAizLKx3
aOtCs5wJ3N4fGpvq1+2CabQfPSgmVqnIbGvvtaP/cqZ7Sbkl7s/hMVM+/1Jkxfur7u+tVBEcFHSh
Vcb9RbZlARMkhoI283UDp66o+4A5zT2toj9WtiRtFiI3v1dGf5riIlkVR69xBtNr7DdIFSjQccc0
FBUTW8sdOFglWtW8JgXXK8plVjStTIPWagOyYwIvhmjkgRzo/Vk7xZzGLtubkz1hPG6ZV+MK+owD
HFO2tm6TlP3KdI/cz6bdqqeRmeYFr+2tGZ6fii89VEBWgHvw0/W94Nmvp+uLj6tpOufwO9x78Ckl
PWBFnjDs00AszLpOZyYUNKcYn7of5k45lfJ60/6X8U/0OJR7v8oQIYIa445wBjFbl5ph4DUw3HI7
zKdhcI5gZzX/d0OAVav6Be1D/wp/3RrRtjqDIVKdMeRGHytAxhqW7Rn3lLbiCMvq6fAHrd27X7L1
TS6uQHZIgaGvyEagdqeOLoAipzWQFH05GjkfcfbBlJD7tfbuKNUABeqY/WEid+aDYRNsdr8nj1QC
phTNWoncneQQn1cL+OvPiNkAh7wGLZDZSu4NFSGjnHDEYZHM8r2y4tFY4PvnUw/5siITQ8gcBPCx
6io2PaGfk9EhulMubIW7jocI9/EbngocDGuiBWAgLImREC7jouzogZmea5RwsiUMP/PaRlBN30nm
NlCXhBq0/MasSMjcJfZZoV+A9uCZrnfoB0NRnQ3MYdiAunay6i53Yrzs2QouspDWUEFtWPGDRdYK
SETpyS3ZpvJjt1O8jBzGJI8PIDS4zr0s+1XCDFUV3SFpJvFVYbgphZwIY2FDzZhF48tiXxfg2mOV
EeXzjrJ3TmUaKRjiBpWWrYVM7it1VNHcHccPmGnRv9JF964sDCQdwvq6tHbUfJKhv7uEdXK0WcQV
x5aroXvZklhwCdYYUw3NvaMGW57tmeyre1q8LWSgxDFVZgbQdW1Y94MyNIj8RxZlG7E5TQESyFAs
sN/zHo/AcaiK8XLacT0sa6u72Ml6mOsWECF9bkvEbtk9n2WZsSKyyB8FIOvIkdySmCFoetSi1cSA
BpAOHV3XdSCInKg35yTN7gEN2FS+KhAX9m0h6CcemqfGnjembWbZpGRnmMYqB04JZQ3kquKCYsg+
5M8HF02YAlsBSqyyEV7KSHNqvoPR/EwyU9cmhHr5OJ+9Piza0+PJfpDY9TR+cV7f+lhmUu5eKGFw
TOQIAwpAngWeOV+yuW3AOU5F1snQgsn1qX0CBkVG9tAvdHxTVL3BGZLFRsP22WIsAnoHOK4EUr4A
/0Q+qAtsK/W7ZubzQGLKCFwzSVJhaxFPHY7UWctFWXv+Pq9opjSbD0niOLLXQ4YGSeG9tomamcLj
P0aIVPN2FqoYLbQvh2qXrbq0EGSRPXhRuUltvGC+StLxlUob48XTFokENNX2Q2DQ0IDWdbr/Qf8s
62bU8mN8UJESYh0gxPcMiEDHCD4U6Q4h1mgvT2KjoEa5Bi/FJB/RLJbon403M3aqXs9jW+/AXUp5
l+1oW3DifLTqW4/+f61VYjMnq/hsxLDD4tdAoVgLF2BiazRNE5AubaUGCBwkWTLZ80gOUevQ8ku1
ZyfE12kioJNf791364wJiNjCc5u0RZeHPYIQuViOcqaKrcmc4J1DxzPiqXu5pbS1hAPxC11ElR4s
qEdd0XPP9OrE9OCICW76xuw8YxoOQzbwQ9XRF2qsBjw24k39s7CBlE4EEGCRh6wZZHQb8M7L2ZKM
3g/anqRVJEA/j+iZNmI3Xgf5Tq7ZeFFxBOWNtzDfy1Ml54OlsoqxqYsVs+aOBFPJcccUvGhwQDUh
1sGzg9IKrXWYN3sqLkNFqooNYbWpnNJFM/rGLavAKOY7lyvUa1LFimWv8WqTN2A1NeHlpDZbQVIo
MqonBeukENH9O6g3GB+PPcO92NWrN62F6V3S+EREyirJuxHxkJwuiAxQ3g7wEi7u6F4c0se5Tt7D
VYGL4Uy++9gb6zs8/45kulAMoa2AQUAwy87q/AWAL7eZfRp3IDBZ7052bpvm4h/2EMFuUamlezKm
2Tbt4oTEGKyRJyNcpo5x+Y3nYciENZjjTFHQPPGwKehJ35ra23ltNaYnFsYxEsb5pIUEtVdfBq77
5iXY64LgnHAtGBhX1jeKLXlk/AFbd8vBCegkOOnnx5+D5wEf+yeCYJ9YOJOGEKRZtRfjdK9LyYZ2
VCa6obRob3sLQkOUJGMLMadkpMCQ8UM3zODKeCSahsYREIYke15zWYPTMj3bUpJGEMaSLG4aGhBC
wDYooTmMvQoPtyI6VHM6Rlb7xVtNGtRxTaVUhEBe8jV6trj11RWZ7mjun77R0AnUwGvdY6S6Tvty
pl6BhTuMqFSCiL8EE365Yx4V4lLOi3+yjxdsKEJ1Z9P859UdqZK4x2faD1NcH9BaJ/+u8ogHrjxg
aaLH/abtfYxAM+/vPoFdIu10Gy89vUIbEiwM8JiSlDDJvBwHRmMbElijKSxn8wR3MlF8PH+6rHkP
z4NuykR8ARFhTUiP3mt6VA1Aie2bTBjsrwedoq2ZTME23ZM7qQJ7SA6MvTz8B6Nowod7vd9FY+fl
4B39HUb/wCc2Y2uWVW++4sCE5ySxLaiejh68CBJlRR9a27eBIfIDnEzWcv/KResn6+XcwpjS2UCm
vrQs7U5t27ZqBgVWDvdQAsSFXQXKNTbc5NAU25SiFnC/QVm5VWc0p0DTV0rkL4VNrbhwJjijZVBB
/2W0KWHjZBny5SUce8uQXEETP9aXXBqi3JnWMnXn/xhyo37mpohVLGTTHL30FKwPPDdoWyVhnD68
/Wqq1JMyHfIKRqKTxl1EEouQtXQ6+DS1cWhVIAg3HrhQGsazsdiZKM7Nry2WZW9kUeJzsA1XhqU7
a118pd3acUiXVrYq6Iwyi49YD6XFVjt12rks3mJ9XaoF/RRzF/VJe9/VMi6DcmU6LoDHtrGn4429
KrBY8zZaz2zYES8YCyAWPY+r4KfR7Qa8Qy6+tWn7MSTGFK+b9BXSncWGKqDFgTS8cQMKVUKfExOo
vim2mO0NuGqj/INz83PV3TNvonBmy2mxacnmy2HEChNmmm/ENBmwQ4v2PRGaKhWkqwQUNgwoxcWJ
QYNuU3CZEvto5HHAnjQZX1MNHA5LK1FWOKP4G2jJZqalFcmPK+uW8hoJacth2XR/UneE8iPYm0DD
7T/7EGUKK98strLNneFmzCVlCPMgWDSGOWoPGNDctaECy+SRT1lJD8gM7+P1o6Bfj5TmdaFW0YPZ
Oq+JiGrGQgHjVoa7iBF4PdGkT2ppXcTV3x7WLMPtZZwDrCQ5mzjwCl1BKLEO4BbNCtVa9m+MDku0
GTx9II1wnPS7uUxL7IRCtG+AxvUqJcVaYGR/vFDgMNQ6OB8ia8HgapWrpbClJ3uQ3q/s7WtyMm5u
HbEV7FPcyOXqQpvf+vRWqrynXn337+nJ/A67CfAkamCEcZgxD/a0uEW4lHMHugLa91ivrbdbroKf
kmKrm6CTcwBlYl8gtIHQvQ+pvrenr9b9ky5IYV2OOD3U7YZQddPEP6JeFHMjsFS8ImtvCoIj9Pfj
VRfIyGXT2hJsNzqTip9DVJ005uxrl4FXvEZLgKsJwFANjl3r1KfkFLENBf9LnXK2heo8PoLW2L4I
jqM11dAyXXAMlAxa+iJ5XzS+9PVMB0Lq2laMPXdqKruwwfdWjrTu6xKEyCORPPLP3os/CowCXrTL
QQ6sJ8iejWHIaSOVNZp6DWG45iKS8HGtSw45tUfDZqTx3EWF0WKc1pSIm9yq/su0nAyPp56/YPK+
vqy4YwE70JbZkj7bZ/Z9UNimwBkHNi3hH3It+TWboHVwXPgu4w8da+a7UjSzpWwWmx6KqtaSdOqm
yQjfHD6CGzWiaGiz7ZJvNwHu+qzs1Tzy79D6R7tQ8Shn16NjfYLFcdIu9D33Sis8jgTY8icepEsB
wZdzz6XXEoXMMnuReIGmRkFng81NGwI+80ib9Utjd9rBcSH35ZiccUKhbgRs56MRUabFsLYrSEeX
UTwD/SkacClzqu/GtPdIZ+UpZq72b2KWcZMk2oob6BYdy4GiTTeeZ5rKHR4q1wOWLMxcb0c30vqT
NnOIZhWTe+YmsfPTgGR0oXYiETX3ntZ+6l/68YrmCN0j6NG1fdsLl+ZhDwKgGdvG6nEjiwANxEQA
kwtFXGfnVYNCG5NcodPkYAH7/neaImBIIUOfy29yiVSg75ZpoDZlrcml2aoPOcRrcNztsUX2IAyn
tMXF37ZnwigWd6pxjoXP7wKf8MKauNUW2VODH9ECkhTzPNj/kP4oIrZv3MfiuWBzTJQPvKT/bbDG
DXx7oUs2o4j6TCMTuaEDNN8RUYQ2UCBt481nYVdMukMw0CKVvDqvCj3vdU9vpk5Lfu1KpnKSLnpi
C2ZQfOjULbtLm8K9qvDsUG7JZ1d/LCikI4l/XHJ8ZKbSfAzabZWKvS7ZAxMYBcSmTscvNYsoCfsg
1LZqgZgj06WAAYeTF3idL1AS3sHWQO2F0ztXEfwEBEnyaNtK7thJ8DdFUno37WKkCIo/4JjcW7/Q
+VHauE0y4ESorD7oMjcuMnwZ3o5spz/NKVlKOtWMWAnL3G3fghvRR9I2oeQaNyriAMJI+3bcnsJ6
XvNJ2utzgwFZ0xdXq1p0cDGdnssEW1I3jJ0CfdwxB6jZ1EcLZoKDtHTnWmcjKrOsIW+gWeKYU6Is
NEQFNWebp5BD1fOfKH9FO7AWdPMwXmcw7a6AlExYcVnVOEKbEm5WN4yCnfWeUke76C30PweCipQF
R/dwnTM37RsVfqHjDw8MQ3taQ6gjyxg2em5XPCUi4EG2oqBRnauSrJkZx9M5ACWjTKzKvzunFmF3
/o4SQwRWN0s8SSUM9W7UXpRHq5HSohwmMDWjTnNkGZAebFZ+g+fFBPyEruq+jQ5TspIF3TPCstyb
uIcNG49hSDJkmuD4mD3vUn3kcw7v1FqXn7bVu1MrA7+e35Yf5EKdz3UppjjwYes8EbYCjmi4zQpi
sq3NJcGy0e8I5DWhnbiF0Wt0YILIYzYFkTOGsZjrzMc+L+bJMyOZ1Rh6HWos5ZTxeA70yN22rWRf
hFVOnvuOC16bhy+50oCbLoMk0IAne/VM7LnQ5Rooe1M9/1zTUy3AmSJIQDbxrcxxQGpGgDFtL2up
miVH7/FNNTF+FLsLW2JZUN2pXZEB9pgdX5qaziGtYG0NE30oi38A/87izAfkDs+CIUOvJw7iHZAr
qXFa2YQ7ijwf7TeKXHS+eFwOK6hc0qoGdJta6FjsV5r4HKYO9ROE3rLSQz0nq9FZaQNrrxo0VCtT
N5+00wLEHJcnkPxHZs8r7XsON59Bq5kC7vNaiemkG14TAeTsxvzEz4wUrJ8uQdEACb1iD9x6ctiT
8tG++uAgNga9kR8ntMsGXdn13t2KFgIRgV6qSEDpbOk/ofok0/3czjyPOl5KKJSTTQ2/uktowwVX
HXIUtyARMQZi9Qk1tGinW2U8i/U8Xj9BTFbQqV9d6Rb0FMWKAHcTBKrYKi0ndwJAkyZvUTQmjwqo
rCMiJVaD4scLQuqz9+smx9rD1U6fFEO5ZyVKVBsck6Ge1fNube1SvXE4dudp2L6oppicMZZemmk7
W4loOsiozb5YoVe8jHPkLbImgvWpo1UpF/fXkwCYVWYSuzZh2JjrLON9vBl5vbydWVaK+4+hpUk+
6PjOtEgkh6opWpzZ4ApO4IlbNfsS5Q19IbETgXhh+/6TLbZf8sW0LFmAW9ipVSjYzBovQoSffTxy
IWeLP/cnwImPnRJfjEu1TYEATjGXxsPzofDRgSWaVZ2JaYSHbr9iZarLuC+C82BdWUJjUb9Lz7PJ
M0h8DzW89qgVw4+KIHXiEF+Fy/2HAhFAknNX3hnqZ7OLvICHlTExVwY4VC8HPMHw+1NR6ZueEEOv
hOnwwnMetTWoB3ou3i8mbdf2r22Hz4jKMLPPmwiYctCJyMDU794xQGVNeYmCf3Hkt6GlTG/UeHMS
0qUHNTTTJNDujMv2zl21izJbfrtkvwaBI7ZGnRQUgR5DztB9CHsBQfvOkAr7uiL+4msvRljZBAdE
kuqztWoK1WMITOsj2xBjIk03zH4f4mssW7fSOoEWv2FChkoxmA9GKHWg07BBlETZXylyMnXsT6X8
CPXqyGoVBeHRVS5u7Ij5Vou8T/zzyq6l2Q/cUb+Nw/d6j7+w4PZvbFlyhTOI3nNfNhcTBLSYv8SE
2EwGgJGlvFscypsEmTAsGEg0e22JwjszqG1gLh4LmsBxBY/r/PzhXuLVbvoalDxS0Vkbpi/d2xqc
NjvwFB4IHED19i7JKKv3vsp+9JBI1Zr4nX+UyRsRN17OYeRECKYyf+5dsr3XtmzxZ0Ryzjrqjp3u
DFcuuJdbajBvcFkZ+jlZH0GVyegMMNrRib++IbGaHb1SxUljTEne5i9hythaE1ylqoOz7LgSEWYW
Op/dd/Wg0WoqXULIA/DVd5L5Na+vOp7wvFkMBobRi4MX7uOcqAi0Irlkq75l1UjVJ8wdoZor2zKH
uZUorg8kBIiQz9IqgpbkrwX9mr2gr0s5/yZnuderabr0okNxBJm1rmcVIiW9/AC47ZcDhvNXQjiw
iNBTHG1ZsbXBDj5vq0maFXH7aDzYtSK733cVMEv6OGLgWuXOVlh4qNEpjNPj1ytTpo9rRNH3QyGn
chF2fl4JeIDBzKARBQ268khRO5TPfKcr7OczeeqnFg8mkBbLQYLY1YWkrLALgdEhQ7zP2KrLMIYR
usGAQujzzH4ivqCnvLYf59ndB5seZ67hfvpLN1P8fs1gL4JVWJsIr58hHg3LQqTurH3fFMfgyf3q
aA4uxInq3ewx3fWvjjpWlZ0GWGh5P7uOLciASGH5CyR4/aJ/6rflVipJPTRJ+BjolWVcBk6gVVku
QfhvqPazv5VTRuvD7ZpLgzefLlAiY5gd15v9Q/3a0wOPj55kA6H23ecGFu4FHHp6vviRlh4H481t
T7OmTuTnYNOYF75/ofPHtyKcjaHAxZ+T4DKfTa3vLnfxif17Un+rjc99c+rNueFv2xDBoI6jv+Bm
mCHrxHw2b+Zf0zmWE7zFgTpj05A9WKCak4QrhCuzb1eWAV9rD10D7AZSVTrFKhtbJXFcyrc8Obco
t7WQ8QzDbd+qhFDXSnXsRq5pYarUlvOvXJEFzp47CCmsOQPfh+lceSsuK45Xrq0ITG8uU63g4P0E
2mSi2BP8Y+/PTG9I99gEKhESx92ES8R5NSntq8fUGI0K8bDhKrEx45pZhJ2Cty/BiCo6cvkkBiDH
AeQMyNr8sRHiolQu9sNJ+Wkw+Xj5qYYpo7Y5o8YG3VZQNdPqzfZpilU8XUdirxlUvhQ6yoDJOnuv
jsUf5EqHHnrvfjBgjkUWNrJVFlYcmMhNB5X37Mh+AUz5ykKS8sH69/R4HKg8fPyEyQoxRUp9PPb7
LSxFH6jL3c77OU71XfCvfKrU9VUP+Xccbe+prjFcxQ7m0mqW7JNJmULyi6RMsNP7z84J/qd1h7BX
tgiqq8y8b5OLhsSTGXQ3oTzLsckiLsFXFe9N0bxILvQYnn4YHb90Uo+SrqZ+3oEIjC1LiE8+BfTY
q5a9LGDGkxfldzcCb4ZOkll5AQi4+j9QTWqTS4yhNkS+nDjHeKVhQYR9ndIRjC/giNPUTRAj5dfp
dAk/9W9c9XmXtRW3I5vLFQN50QjBy1CG7SPhKsIX6X5BYaC56V/YcxB8ZL03kr2aJLBqxEqzDjoe
WwAI024NoimwRxZ3b2IhPfxnlkcJVujvbN6obSplMh7CSTx6HYJLVhEjhcptiPn1COnynKbOt7dx
76M+aCXcys9V9tD2SMY3DFmLldc7p6SEyCpz9HHRQjpN9U3aQ8HiV1N4+elGRbn8uikVPCRc1Hfq
P7HopYbB3hPhO4l45+drKXiACjABzkJkCTMXTe8FUUNvZeopc1AD/STTiPCzzF66FDAu02HtKhC4
3FHKp0utKknkNpp3H9WnHS3U45Eu9j5lRpXUvTQKtRl5SyGWck34nJgaUEFQdkpOw8Lt8gTyCDNG
YwDZQ7JTAyJ3SEVhB+JUUEar5VJuhwk0JlaCsVaxoXuEFyaM1VnQ/6UJGqN5+xgzoK9Re2RlLnJY
Vzjb8zLfQYP9d/R/jSr7IfNQKKHuGabRBOdAdrTtnb5Q5pQfhGR/ZwlSV6DmKjvj9IhrDhLExQoO
OyHpx5F+1Rczq5RZsJxIsWHmD85g28MhQwW1eSk5ZyRxoCobIzdnhz0eB+8DTt0LkO4TesbtnjuW
NTLBPsw3Fu62x+LLG024UXKlX7wzEBxDzabtv5lyS9NkCny7FzuY1PWo5QLAOdmAdLmuQJH01dqX
HV+YTsYConQzRrKRjFT4jte21p254nLqMF/INgxuesAKeUB414t1zdgYYB5K/lMtK8FPW8glpX1c
oCEt4fyKmM3Va+8VgxSqYIdyg0U/4I9UI9o6qFk9mnAg+shaQyDKePSCudRLvbBPHfLiXvYclVOI
IyX6GU/VX24yvgLGa3CtOUGEaqN1P7aM1ZNHQyKFcOejSMVRV3UMasquCankFPXBpa3p5xZUeuCB
LRK/2Psthm97/Ju6gXd60I/q8F64nJ6jeYC1X8CnC2aNsEID7d2WCoEM3ci/hs2FSyZq1OEgBIyb
7D4oJFNXjISkOEMuo8lyTxvlTjGN/KfpSYdy2jopb/bHP0KqpcUHE6UxLphznOGItSXfH6TWSyw0
7yokwAj95KQDeCUxTaxzUgh2T9ro5QwunXeu+JD5IWdRUgUBTKKI8VJBe991U9A8E+vlNS3j7mRh
Kk97mtQK4e2D1GuZxS+1QjjqZEe9yYa/G90yrhzPyW3WX3mT+e04qp/yhsqqjdEj6iypWP7555wK
Cwwc7CcmLfdErj0Rp4QrT9jQImnHqt4REdaEdyOATwkOuHuXYQ6VLd/T/MrumSdJaIdn3qATN63e
XA9MhTE/EnG3+i807iebwg0htiDu9q6dJhrVy8LTBBv1IA+H/d0yjZn2tGMSGfn3a2cwVJ3/a3/n
P9/9suZKtqScn0C1WN1JbHC5CwF4R1BL03aipvKYhrMZBSSKDQojGSTGeYr2LHoNZHPmGxkHvluG
Mfk5un7L6KMwbv/leAC4rCgxYZjf2T4n8yd0UdP0N3yoES/eMppgLEJC6L6Fz+qkDrx5SOtexf+m
YDupqDPKKPc8ULuUfMHBd5ZME9UeZbDd0RuHZVK6disl0Vfpg3rLoqcyycb1fUP9QnUWubYh/BLE
hfEOVjIlqn4GMmNIqVy+F8+7tBB8ruAl41J1cUUIw9+UiXXIA08hX7iVR/nC2cW+ygZy9sdBN9pS
9bGUA4tc2ZIB6hPyRYQ7Xo1J/ulaseI1DS6kCjLXCAhvZmuV8seht3Y8Dr9eGAp2X6Eo+sZnWwPi
aCpsDt5HoDi8JT6uCUJx1+gavawZDY3PnQJvzZrSOw1L/2pi1yP0ve/1PK1M875XgGcE7UIGHkmL
IdnH50yKIbQ43HIURPXmrfpFSymuc6IVjOwfAb4/Zla7KzlD/wJ3QavZTO5tgqcWRhYMwoudXNlo
4i2rxPEncrfcLzxbJZwGB/Hug0q7Z6Or5xT+VlO9hQq7nG0aAhUDe8Q9AS+4UgCT1Aoyri+B5q1o
XRcwvQMQEIa0GLOUPJlnswzHOVe4iM6f9Y6yVYnVVZGeJbe/G2L9M/AkUDVJCJHE7Iw40LPyB4is
EXy8ZdJa4RZgOwmGOwAF/8ZriFOKpzwgZxpKxBt7Q6QlwN3jPLTOt6Qxb72TBQqVACSZxtPWnMN+
nZ01mt6itde0JtdOLJ+kELQwouaf10pr4aN37cIlaB4itGJQ4qXj1m3AQqXGYvhqU50EJO0T0zFX
2bi4r/yMbOgsF/kYKskXc0am4x7J0koSklDoZRuZttq07IEaI7FIJDm8izgyjDCWN/Mp9rzUhvVq
ZY5O62iWmQXNuIU4S+t0+HRAcYilEgJ7IlfjXTkEGPAbyxM0N71H7LVa+qu6neywdjKBy7To5WtB
8eIq8KCdrU7sx5tlWA5ZfIdfmbMpH0hfV5h4s9npbQWvdsPqgb5eKJqwlPDc1hmnr13GERbrUPP4
Vv8PnLJ+bwIl6RPrUp5zuiAhD/HYDWsckZqhuD+UDr1TQdYbFKciX2l9HqZ+4EsnoNhLQ6GBN9QG
ptMZvPto7BSF13ipeokbb1wAylhqshYYY1VPYUTJGGZA2KnYgMyP+NghO4Ww7Muy7oqjkhUjm9jU
U2v380iBZcRsJN4zqnqRp8w9PoYg1ql+Or9uLe0GFuM0pFg4oQguBvHh0Ql1dIxbnqs5321DhAv7
iQ6OcgL1I4CYMgyWs25/tKcKOXZ3oPZwB3G/s7PRODf2PS5jm3HilM3ZLJqW/NGCHIi084Wwr+lZ
dGZXA49KR3WtU7CaRsAB9A6zCivWEuRffvX/lFXmr/tUJdpMTC1jugj54a9U3MPpe2UwR4hiNHcU
HQw4i99Wv81BOqH4BozI7Oos1gTNVdnlvGsz9cihpVDzzkJko3PIL7sNAmJnk81mXTXqlwut2oZ3
UoglQlA9HN+ctiiehCxCySk2scnH484QxeB2QI/8hacmNT6QiBaWBaIkwoENkzZlBQWgxuyDnHvg
qrXbgpF7yLQWnjLAGUgiOKwsYfExqS77kJVLug83FKmOdfRSd2nXa0BdN6Hnt4BBuza9LnlCAdA0
G4H7VwS8dF7As6Qc00sqGkFsHf7Xfu64gGZzEEidTqMfQzxCZNHv9wJkFEU83ckSjUpKsqW20+L7
hXYmApBDCgkl9jVqruR9TLd9jGCxi3Nmvbbx3C9NgvhGtg8pSkkSjDLEEF4KMA+YUM7jYCs+Z67d
EIX0DdF57KMrJXxSlWLkzeSTdDdo4WTzlo0Gh2DR1CrRcwfJpPW7WmpuPJR+aBipgcBfsvoRlj1Z
5Cq0zEb/BqY/2ADmdMgQ1zwgYTSSHnkzLq0NxF7jJqB1uZKn9FMplAqmJakn56NT3gVjz+Tjd5rL
1pBOl8SUonPQMetr4jQC1OihWdcfjFD0fCJWhWO2MPY32AtUP6xNwqpO9GKEBRssMzpxmYK3bPF2
eS2j82vl5EFskFXEOBxlZ8cw/uD2449x+r0ZQ6HjQOcmcnx//uwM7M/XoHKeWNPFztDKDG8kC3cH
6rHSaj1IO0v1Yp+2KfbX+He1lVfe89BcZro5wKgEYGGqubwoPn8zH4sWSTIOA/z6dVDyp3enuurO
ET6wwq2P6lToJcSU5mQ1qPIFW9jHZn8rG8DHXVLvb5NDSyLsvVFusASR7IaIkE09n8xseU3MDLIA
2yH03S3GZyPVU0WQeCLwCC/PxH7hSo6Ma3wRdRclucgnsDJ3hIeC/q6YciJpGVGqHYtn3NQI3oFU
rK/5gDb6rJcHkiM523h1/t9gcQ3HpGM0kRiJzVgwWdcposOezUmS/dyW9ENQOZzqM+C9sC3zk5uV
kTxArjx5aYJubISErOz7+tRtMZgDjR+Ee/mP9x8fJ5FEDEpqhTmJToo7KynQrzhPnco7wygImFw0
Vn9Vr7z9XbfedIIilEDoUvRYPCHjFeBofAgFjw9gjGwCD9hpDOeBTtFztFzr6HUzRJvqVx18TNHE
gBuj1t3TWPsSNEfgcFKqXKUKlFxG0FfSU59mSwmN8j2bqmBpsU8eCrvON6zxhFj26ooq+lzLZd7H
v3bwIZ0bm3sf/ooPfNdcJntIG8DN9kwKoCyLkjTt2b/n1qDCE3x8RDnecN/KbhZcL9I+us6a+Ei+
tzmOwWr0GgKZx3B1RY4iPkYyIis/fHOWOJBNqw6UtFPDADpLEbwY/w252ZW6n+f9qLvzFOjMS//l
6ZLl6RaLAP799nlxR0HjHddcXDQPAC0kyL3ZHE5HjxI83vazEm7nShXSmowzsCFp2nVANbTCDTJN
i1No8xaj6KhoRhxQeUctVFFYOcu8emvWlDSVM6BYhcTiQNV3bi78zNrCgxQQfzSWYjHH1CKivSz+
B0MXA6nbV9vc0ymHdPcHpdqLhzqT8K1rSc1MM3bjKdVL6Ff7Q8ulrir7UXEWR7gbPeZ1WLrSCp/A
Bh//fyYF1jK6izo/5eNnwtrWAFAPzplHc0BwaJhDhBvQuMmJwOFyh4AQhcKC7Vt/uuwQNl8iqFpb
iDKszRJqlGZumsZLqC3nD2tbbArdvF3oZCfl9HHmEYzYuusZU+VKIuv3hdOhRNlI3YAQ+IJfPy3m
9t5h72XIFC7x7qgeioHJIWwwhmLQdU1fzsYvHJhU/38KsJe+7fWo++tBUARqG8+wow25uh7KRSnk
iHbzCIrL/EnHdIEAeezajZEqdX7ymSL8VAep+rSL+V3BePmaCVsKSnrQWyDgLxCe1ZTJc8bcHSzv
n14I37yinqsTs8S2Ah665rJNRm32R4le9Uygbs9TXPkAmkXJAnwaH31Ax2/MSt3B2emIf+Ogqoci
hLF2Z0kodyWiwfLxPAPQRxnXajcWP8qn28x4UN4oUZhr/ybM2g0Cu2h8IbQ5xucX46bBsunP1z7n
w04rlX7kzrKn5/Mp7B9HTLoGWhhxP/7cCvicOoZFVYDRfp1sLK1WsEaclendXn6n2SHV60KCbe4Z
Aa7wKph8ZxMJoBqsSMUhStRJ5dBYZ+d+d0N3tHdGf0OcHxGUnqlpgdBEWMhBd7DLxNEX3leJJRrR
G3pGKVUerw3MXVH5nfYEIxsG5ChQP9Mama1tON/3epf5YmczTWmb8kXxMxlvWpbWUwq30adtL/p3
pBHqUvQb9CpTbzB+Us3ysIDOcGkIWmmDFq/BBU19zliChB0cwVtOQFMpe9zTNMgVAHoM7VkDI+hH
OUwJNEsdQ5sNE/lAU7lpfv9wUIXySFOl2kT72ZzHv980VahQki6oEH5vhYBCYPTgDYHlKmO3/hXo
v8rpw11y8goW1NrzCxdpei+pqyw0vPWukjQbtIMOetoBYAFEaCs7Kjjjgbmn9LYYMalPZlTwDwHg
+7u97df3zFdDiPtA9WyQlRxF3dGkkxdUuIkelRLBUMEFVfnrH81z2dJGLOLpk7R/b6+abXSVm+wz
wq9cTXSIdbyT7UNpsyR6iAPqcY2WFDx4cV9oZUcex4hhW4sw4KD61xxJ0kqxeBaXK1NbEoi0dz9o
XlIqKuSOJngGd+lS4yFcsJcIMkUfrlIBiO5XnDiyZjKFludxJc2Xs/cqltmJ/+6FnEtsBNaeyvqs
bHJkYeF4r6sMCElbrlYZZAN2xsNJ9oa4C0jFdCmzqBnQ8K57s0Ipod+AkYOzzqgmDPXimfey/TzM
5wu3g1pq78ddgE2VjXjK+zYgaOvzIA3a9QXOJZnnDxJTmSADwNgsyRrcIfWrQer9wRLCHBjS67Zf
8t5yCNoxeI/t2qozEjVMJfdjykBI4wEZ7WBbwnC8sMXWpKnEILe6VUrdYZq1/J7VP4PDrMoUK16f
ARQqRdAzfbmOcQFCjZhIN8qvt07qia0y7zY7NgnWRyv273EOzqlcvtUJbbdg9njq3JB64JS3B0Dq
bhkC0dNeTBlLaQHrIzNehhN2BdnSXDxGJAQLjC71rva0L3p0nSFqS0AahrEN5M5h4fqLEaTC5AvB
0QpADCYS1OY1wADgVuLVKgKEpJmCcu2PUjqGDrziDoaLFeZD5nsbdYKAd6DypKZCLXH9jFYkm9M1
7GElNwFlHHO9GSHgJE3hmybyoVofdx48FnAxtL+ZY5t0v/cMgHyR5m0bhj6MNgmwyqNugVZ93hFB
AkTXbPoo8175M2GRY1Et0KC7KmIStjKeZ0fmk93wtdZswu5ZEo95xoPAcsmSjxO1O/yqBFeyqPBI
jZWqz188/aBl3YH3ofBjmkCgHeurJ3Pl3lbj2BGcPpCK8lKBxFGoLT22zOoNMeDCxyqvTI9HARFb
LX/1Ef6srsOHtAIjlFjHuhrsfiYiPoCcMgrAVNZRqONcRp7j62ZNJSkWQOhoVcXBxxMUO5P6FkLf
wkBhRxRCJgTzoPeeZPzN1nOefQeZcwWouAqQQkDTNc0tboWn1xF4Z2BAXBWQcyzN9binbHwK3Xno
OkCzEUVNG68t0OchisaTVS3nBErUWgXVcHNa9YY24IDjDu0ssLGF4RbZ801oPA0U8zJsBjd13b7j
LlTEJQx04iBM/+lM3DpRDPmXBwIJKuFNyKd8HA7LbZzDLDWZ07RyLBF5tv/k/qT/rGyMh7g+1x4O
fivMPeIWaeyhFD/nziSFLluqF5cNEbNT/nOy8e70G/rHe32y47j9c5lI1AFnaHE6WEF6f0KRihXh
eF+5+B4D5W4oqCSKiNX8wOsslundHqKpsvRW5PeDBHo9zcKa6nlFj8LSjWEeRrVBoH9JOiyn2aLy
e3Tp3A4Vlqb87Rk+zOWPJvH5nesSqW9j5gnzX0qUuH9+MVrtAjnCYoKT1n5I/C7Cq+m79ibUvP9b
PSbNBIEJZXmchOtiUtWXwR61FRQhiHHdY99PKEm896nJ95me5m/hkOmw+9qMoF7xknbn29sogwZp
J57/AV0jeikEj7xRlo6Sj6idRoTkBb3MHR1aKyeUowjegb4jOQlReP+VlEbm+l8o/0wLTRBzwk7A
lxlxE5xoqvyHsvArqHszwoO7k+f4DaDTnKsVJkBZ2MDsVp8zbgLcFTidT8eei76GMWFv6/FKorDh
Tkd6xJAZzOoNK/x3jzMnBrQCc7KMKdiEsx1GASSEYAj3GY1V/vGZRfKuszaheT8M36AezDVqOyIe
upwbRnfMRgJeUWnihHqPu9s3pHaEUkHdj72g+6F6Eyu1RavfSQBzXi4puzJT76niZRD4B1yZWJs8
HJ+r1hnFFJV09Re9DoPfQIMmZIt0s4mgCJlSFy3Brzn4xu/NXMmew8+SCJXdv9pFXpdpStbYH95Y
V1ABkEns6WU6zIq4nzgaDKcVraxSRxZDKUVXGjzpBQS1Fd1BZ8wGOdzqtGPVZ3g83HvVpHqPBL5A
rrM1fJfl6c6vo+z/dIqEqoAHdgZ0rL5FF2fxAvxHu8cYsOFHp44QoY1cBHIxko9oj/gX6PohVnZT
QV1LJtaKrU+uaXLVVUGRyRDAqW8F6KLkkWrDSbyjBrMK9ksP/5vr1e/uOjlToXydf76gFti8/pDA
AtouJFqrUrYyGbILnQiSqarysP8KCbHwNzhXIFo2bLYMsVQV5eeQgaXH88x4AXvAo7lAQ1Jx5ZZg
WdGXJYinOkFewgXQdi0FTqC6jEr9u7df4EI+RU0z2cBkJLOBKi3zPGxoS/P91YE+cCiryJjjsQCR
osAiwGjctZGNJekOsRrgcnfFw3TFlo3T2THovG6/GhfVRZfOmNvgd3/1lUTzP1qJs2zOO8j21Tqu
z/Yb/cIQbQVm4LlwnmXswlN/xDWC0sqrTtETwSwrIxTxHtlQrtjHNXlxqIIC1uqVZDBLtL07hOrS
cFmtm+m7CBFlfxNS2f6TJRwpppn1Ubn8YzQGp8IfxNiwlUcCLgZFS4cmY7Dydcn/DdX2GHNcX9GP
/dB+dguPgU68KM4UzkHtP0EgQlDRTHTHSaUT8ogVRyPHl22Qeauup4p1DDMgEtky5aoEitEFAHC7
OTkmJqW/AvGfrDbYnM4PTI6FKSYCiAoukTBfyotbP3Y60HMjE2unGkcXjQNKhP5v1JAql5x5MsCz
UuKtqU7EwWreIZZg2Bt/kP9fCJoHXEMUHc6uP2SxXi6WjQ56y31f1+O1+F9OQAqNORNzYSANA5Mx
a/9lzqOKzaFYh/IIsjMOPa1RQOkVw3Q2oAnK7N8moG6C0hZuZbZfSAjS6fAf2gjnHYWOp7uFj8Kh
aPF6EWeREL3tc/0caiKeRIn1BXE7qvmiY8OZ5p8Yfu+K0J2kA7s4LCF2K3DU4EyKb/CHbWeI4+zV
jmGEi/rx6iu59JL9hQcWBrdHh6//FdIpEFV07XZg7QTlQN/thF5E3ZeHLDruXE9L+M9ZBniEbkrz
2gRguRngmUvZGlTcXMOYH09ZBrnJ17jqiHnUp8H68+aKR1TIY+pPtLqwwZMjbc3m82YzEHFOFOsW
TScDCalLHGwPjPwtzXTyebdCA4eNWpUaOojhjoFpDfpqRopcWko6Ib4gjhERm+FHowtJPoSp78+I
aQwk6SOTKaFl2k1Hmmof8p74fq/C2R70y0krTo4W0Uwz98wp5Qta4kamzByFZ7VIIhPltVqUk2LQ
wpoi6PTYK33gFkyAR5kQapL/vt/SWMCUK64EI44NxxkUYiA8/SBwlfoQHOx39wgdsQoszgHOBNIY
SUjQ/9c22bc3c3wO6Lw6FPK/HmXLQQSmrIvnhZA+y2WRTaBEnDTqhz8Y4O1MIa5khNTOCTOSWYwd
w1enhTqP7v3MyDjrUP40zjHuZscO2cRejXxbaW74LZ/MWAkKGrYZ40nv2KJo3Vm7lR6QgaX0sZyC
6hNmStaoAn7JgvH27Hv5Kh/OXjTazl8THwxNiPwH+2dSrAZA0aiBdkgajySCn0sd3kMujl7shdQf
zI2nf6+HxLwwxgToNVkKvWLESUkAt8t62lCbEYCRlNiG4bV1Kl6IJTObi2VkWgEQaOz9+ZR7NxGy
lPWjNywPS/jdYcw9XYbgFQvXawf3hkivatzkJkjfr3iC6eetRzUmIzXnRElXM1aPcL4JFd4heVUK
E4BBenUrWSg0PwVR
`protect end_protected
