`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
B5oV0LSLJ3kUNUJBKeqsH2WUWt2sizysZ9Su5fuxPdZiLELaeO1lgIXkzjA0OX5BSj+jslmdq96q
D4sk3R1Zz/itlnQJcZBUg+JeDkVtiErb94w4zE/AQYCHLtV3/9zlvOtBxohEkEikIe7umVEQ+y/0
B7+e3B9OFbI2XaORc8QQrxdbtCr5yKrWAeDEDSpske6H2MkBRhBKOfBlyr9AHjtW2mqzPRC3ZFOm
72tFzqpYEs07W4IZOOI7QSWnFjY6rYXVuFKlnLTzB08rd/lQ26C4xXxOtetKbQ73AuIikn8R03MO
NmAe30OCr4Y+MrGbKTT3h9mMpdQp9y6/6OpKTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="/EVrWzwK8QplEXK/3dwbeMnH7AOPawN1QoLDWP2xKlk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
CyKTdlSp2JSTVxLZVuJ649XXf1rnnw+C+3jnmQGUPUjBPYV94Il8O55UFk4wMpPQm5AU4BuEjc2a
LDgPTwuS/ULKYpUEAvP7tjv7xhuXELCa1/LU6+qIx5wQCkYi49mMqcwYJHpMmMwZ8oMYu11ga3Vo
FJzM1I3wwYOfWL2uWkLzbzbCP7lv0uFHDSyJW9lTBUVp1yXy3Gv3GTTvXbD4YYZdN11+2OQyzOjp
urbb2jo7/KQ4J8iEHrnmZ09CMVZ96QY7LR6klVDT28GePhs3V+DQ5zsH8CZh2fY3/XGeit2mtKla
KpXBxeGBe9JRyg+SK5pbi7N08WrQI2UELAtBl2NqAZmbQJsfSkknlUQ6AxD9fOZ+fj8TarWIHMrX
y6ltRt4RlyBVSG3n3VA0ESUCZfgmZwBEbGgxsO/rxHxqRZCgYVsuinbv3pZ7aJcUcDxJi6UZ7X8c
XkB1J8leJC4iQxbZ3QopoLEeEmAwdlUqWiHUdgQceIJadqyowF23mmRldQGd/FUzg4PCsj4OIXtm
KHGo3ppt1XOOQAYzY0+5PYD05OEA7WYr+bJWc7p7ubavJVfcseontHHCBXauLiy0e1qwj2vLHfsb
X285/IUhLLTleonWF+Ao4ZZ2XkStVW0TAhEL4w515SKgvQF1Yc0XDc03bzEbR8sxU++PCyuiogx5
zXT/nu3vF2l3IFcb8bAc0mB4ZmJG9X5VN2tlTQ/RsXIimabySobwM4tGKsBwqqrhg+H0MMVhbPwX
/3a2PJkinxO5qzqy9gFR4lgiFbWSN1VX3HXUlYV3G6LSUbA5+PkUbuclAC7vS+mv93XsSgeIusPc
3xkS6hzcpaWe2+gruXwfliqiWxAsn9H4NWFqK1o6Vn7CuILr7bLz5fs9lu8jHWtILOGsscfXUUSw
85gRi9njYr3D6Lu7aK6WMxcCRsxAGsHqfJ9XVa13xeaLy45mbYc9Ky/wjS8UdSaQjHUrTMoFa/TB
QijalIrimnWjyhCbg9wieYzG9tot51tEFcoRDlvr5jY/KNIRWY9NEaQLRCkXsyqxFVSq1eL2nXab
A8gZCkj70CxrBT8CbwmlkVJYB65RPGJBXlWz90dNcLiWM07NHjeb03W6NWfqSLxOx/Fcb2BnXS3D
YxteEl5VMBjajTLqZwGRxtsrHmMbhs2nCOQII5HEgpco1ewfLVta2ufktQOIkWaZ0esOJ4Navaa+
ynWkF7n5pOOUmMuUVHiiOA==
`protect end_protected
