XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8,�^��@��U�e�QV��
�|���ǖ�QY�g����1��^*Q�I��  ����"f��'-��;:��4#�fR$8�N��K(�qh��+1�p�{%=��	l�2��Χzkf6�c��31�A��n��!:��-��bG�K����t�L��Y��d-ظ3���B�p �;XM�{���(�'�$��#�	�gY�Դ�M79��bB%�]T��,sm�n2�-@�����[~���ν�I`�Z���l#e�w�p<��t�Si����c�P�$FZ�ʨ��B!�����!���Xolͨ�nP<��O��Uj�j�r�s�eS���X�9Q�"�������~�BD`�; 奼�DR���*��	�/qY����F�^�oB�/��~"�eھ�+���'�_u{�������ڍy�֙Ǚy{k�(��N򰥼G���t�GG����p�s���LK�o��P���W�}δ̃*8���8�l*{�x�^�fFp����S��d:Ʋ������X?�L�!��[�J�
(��2c��޳���2���R���h\�j�ue�M}$t�l5�OD2LY�(�jr�d�ޗ��g�d̵�ZSb.>=j�|� �0��=��Us�e
4�b���w�_�_�8���6\�|d�`�XA/u�.���jϝ:�4�J�w=�ㅋ�g�r��y4�L�boPy�f�?�޹�h����DPiԘ�Q
͖�⯻�Pܧ�����uΪz�� X!O�}����!�@�������q�}<�UXlxVHYEB     400     220��M��pS���r<)����oq��3#$FR�r�Аz���-�?�ŏ���FS�m��z��-Ao� x��Ê��2�g�.�`[�&�O4��Ro�N��}�f�2Z�vx.WL�ScR��=.�����=N����>�8-o��*O�$���oH?<�����K����I��e����+y�G�C�_���:��"��}hK0�X�Uw�߷��w/�"e?M���	,��h~(h|������Z*QD[�ԜM��iB�:*�^��A���w�c���$����b��#��yn��2�yTR��OrV����}O�sFPc��K֣�a2���[Lc� ]�jH2C��~_��S�������yG�A�x�U3sT��p#��m�-�u[1rE�g�a���]Z�;��
ޭē�����k[E��$�:lH��	�'7+�+ZϏ�D�v�"��R
�ЉL��r�rs�����N<%�]��C��`�g�&���mqok��q˲3&v�&n��ֳ=�/
�[����0�,kXlxVHYEB     400      d0=�KQW�`-$��M�ߟ����j4̏'~�$�ρ-�I���/���ߖ��9��|Ǔ�t��z BDnƵ�<�K�Խ�	zp��1�!c���`&��%���;�]�`�GC1ϝc�b����>w���5�J�$~8����a��c򲩨L�g�]NEu���b�z���3z�<�9>�#�Pҧ ���Eh <��+0��;�kl�c�
��5~�XlxVHYEB     400      c0b>�8]�T��,4�_ڗ볒�0Ĉ�y)Q� L��b�eo97��TX�
�=�����I1��pQ<O�i���D�nM%M��')/����Z+ڌ�;l�Գ+~�*��T�S;����# )a��=C&6��@4a.�X^EƋ^]x�e�I�5>b̍���b��f͖&.�kn�����s�½�����{���XlxVHYEB     400      c0�����==8�5,q�y�Lo*[z%�b*A��[�E�^!�X��`��%��!��h����_�x3?�'�m���SH��lY��ť�G�l�}�%6�|�o` ����3��ೲ�>R@$�S�gA�_h
ϧT����	>�lv�B���V*	��3H��6���qJ�cP�&u�>~�>��z�t��G<` �XlxVHYEB     400      d0��e!��ѓ ��r�(��m�R�F�|�4H�Wd��>r꯸���C+4*8,j�I�f�F`��;��'�o�a�v�L�pu��&L%-I5�n ו�ES�I0PA'k����S�?cG��bX����>��}���sЄ��͙��zE���+g+z&��-��������g�Jl��O��Aw+�a2 �L��،j0���&+��=XlxVHYEB     400      d0�0`V�+�>N>?�G 9/[�c~��bNK$��A�����}��D�Q4ص�����&�:$Y��{��6X�j ��W;��G�S �y�U���g_�rF�~_��au{ݹNN�ۍ%���%HdE�}��[c5�25YF��ק��~�	�r�ƨ��d ~ğP��vC�آ��^�9p t<X�vW�KI�w�*UY8�߅G�;���aQ1|?fXlxVHYEB     400      d0$�g,��Fb�~ޱJ-��uB���L����0���ml��C�[H��_��3B:u��9�Y[���F��T.��yh�'�y�k�7����EZH�A3m��SDH�{Y��{�{g��];��۔,lA��ⶏ��!��m/�;�<HtK��/�D�[�'�΁eW'����]K7	J����b@=���w����Lui�'m`�y�XlxVHYEB     400     170$�O��6�~>�z�:���၀1��9j�l�102��P�	c X�i+�J�������!��[���p��~ �K��f|��e�T\�,J��J�� ̊=�k+0���>��qUf}K|!Φ����n���
F�P1O�@����ߩϙ"3��^s�W�;���D�S7�]������wbq9�х���Zη��S�u/�yY9tc��lIF%��p	oݵ��ƷC��4�E��
jX1����\���wMAj�:0F�'^3��YY�ళX\�)42^Q����/�.�*��y��fE������A�ĺ��P���'Y�'�P�Iި.����{M�<Ý��8��'7W�j ��2�sH�E3�����S�&�XlxVHYEB     400     140�ـ�BűS�XJ]���(��V*-!]�R�9n.�d4&;���9I<E=���0lD����O5e����(���a��@�ޟ�W�	M�8������k/�Y�D����bl��)�ҘB���j�HId��R�W��+/�x�}V���I��8�<�c����$�F�ni�x�q�g0�qI66�r����q��z�u�NT^J݃�&]���z8�"�xWSa�eC�!��nƕ1O�����&��D*��Uw�X���\��!#���)"���0r���!\��3���RY�~�rov�\�T��`��|ߎ��ށx�#z�uBO��W�AXlxVHYEB     400      f0m� W��[Zꏅ>(��[���gL�d}ё������_d���v�t�v�{mk�q2���Σ��)�1d�JgC�لܨ����=
q��`�H��+���|��	o�ٰ�$.>�ľuL�D3�<��ǡu!xa����W�F�n���p�_�O�2����r(��5��Y�C@�C]ȃ����g%oJ]ZS;4����F�X<;(4=]1���xT���<6�" Vȹ�o���E:�XlxVHYEB     400     100ueȍFRHʑ�����E��!O����L����~��֘�4������52���-66z�J�a���,�8��_%�*:��5�v���m�5����9���7)ܱ��|x������g8��Wg ��Æ�v{��~�f�H��LT#�Q��`��'���vSڍ3����w���}y�*V���4`:�}й�R���)vT��v��|��܀]���|P�Vˉ�C�X���k�Z��2�(�A����9���X�ռ>�����XlxVHYEB     400     110��^񬰶|��"�<�>�m��"Nkq�X�p�5\⋰D=�j�2�a`�?W�YI��h@ٔ�[RLQ7�ή1�a�E���+*}����p�c!���4/��?/�@�����})��`$R8�ﱎ�0i���\ZXvli}�����G
�k�<lP��]���)q���I��Wx̊K�?�7x 	��.�)�(
�i	�_�����"Z�Ve��=�3��V߻�\h�?�,@��.~b��eV�s1�Q��в���mNJ@3�2�`�XlxVHYEB     400     110vls��X&ꖨ����H�P����w��&$�=>d����uNu��2��N�=���GQ�sY�N�(50���]��?�!8͢<����
{��1"�Dex�c�%�<hG��aG	��*��FƇ�6w:;��UVL%�:�K�ܳĐ�R�:�~*�����J��CI�I�^�>���������X�c���+" ���9��L4�I�O�J?tؖ_�q���V*6�)?d����f �[C=�5�]�/Ǌ7?��H:��>����q®���pV�XXlxVHYEB     400     130_>r��g�j��"1M}��k�8pt?F*�G)��>�y���'���~]�ȋ	`�*eC��!!�ѷ
F�Lrs	�t�$W2�=�"�]�(OY��g����ә����u3�*�m7^����y�Жne�K_��Ft,J
���2}�l$;`N��+%��ouJ"@��Jp�jU��FT����<�$��3
��:v����N�N�muY��'��@����ך�8&gfFy;�|��C�I?���%�9�.�By�\Z��/�0�f�ж}b�&	@$���O��b���߾^�h�|��|L����=�v{+XlxVHYEB     400     1001��zf;������vbi����![K�*<�H6��nO��́p#M��4P����,�i���.:��s�88笌�[��Z`&r�Ё��F��tA���+�k�����z^�� O�43;3��߱l�iU��t��9F�5lB
eI-:*��{^��g�P@ -^$!f�	
��\RL�|y�g�������Cl%K��P@Db|h�?��ɘ�O�?��x�$e�(ƛ��0V9������ߤ���G}�3ѐ�ګXlxVHYEB     400     100  �J�Rpq.��b��Ww���٥�%���'6zr^��	�D��>Upu�������3I��)�j4Z{�|���ľ=��I��L���N���|�4�3��/<�4�a��-4RԹZ�1ֶ�(#�ǴЫ9���G�����r`!�t7���)���fT�.�5��j�D{\�>���$�V�x�pS#^Ki����mO��@^�ٖ����J���4���cM|�CTq8��:��.*gخ�%1|"!y���txXlxVHYEB     400     100�.�%�7gU����m���K��3�n~�*�o����<�_ft��RZ�XT_���.��s�{֦)���j%5>�'�LHu"��8���"$��V&jU���z��?*�b���Y�WC8���~e��*1�
�L�'VhA<�.v���^�����C���*r�_��<	繜��_�Y��$.��r�{2�j�e��uk&s���}�z���}�~T�R�&�#C@<��2D�~��9Z��Ԑ���>'����/񑚢JOGXlxVHYEB     400     100�i�][����֭�Y�B�)���=+��Q������u��8e����3dk3����l�������XW�Ǉ�zC�[���
��{�0����~�;�esG_ID��� &�e9Ս���/���ѿ�:��x��0{|�=�ŀ\^��E��J! Ȑ���t#
��_H����H��Y�����MoU*yb��\B'0�}�C�EK�,i#�澿�xZnM��a���@�Z��"%b��{�����a����(XlxVHYEB     400     100�_�F�o�bGb��S�uP�S+BlE�dG��(vX���xf�cĔ9w�6��P�Z�H�ͥ��C0��	��9y�b�zl1�� S���$�0v��ȶ���V��1��C�c�|O>������j�#xf��L�!�i�L\�� �|ȑ��yF�ţm�� �i �e���D������8��23{hya�^�K��c-�!U�u����� %<h"Q{U���9�������yvxrm�e�����Vc���3���. ��XlxVHYEB     400     100������N��u��Ŵ�p1mqV�-hl�T���v6��:2�F���i1$��V�����7ȡ����5x�P[��b#�IhH����"�K~���^�����EŸGVn�O�S���^l�ėH�]{�v�fJ��V�!@��_�\?ih�.ynZ�f��U���NR��_�XB�ЙT�{���+h�<Ѿ��i��\����r�v�!�fh��s�i#%�R��,��$ޱ��Ӷt��a?�p#C�em��b�%iظ�Ҳ4�9��XlxVHYEB     400     100[��&��uX��s�IgvO������d��G�2�t_ ���p���%q�>��]���U�;�&a��k�rV΀��"E�2&w�t�챹FPZEn���V�Y���h]]A�g���8	q1_���`֛�=�c�|�c��p0ԍ���5n*�+�L�wÄ�M
����.߫�ʢ"Hq	 ~Wa�Am��b�k�bfA<�L��!]и���m�,ת-�*tv� ���ɿRك��qM4�ݏQ�V��VگJ��XlxVHYEB     400     100�0Z�[72�P9����u�2���������K��������b;`�2��8��L�*�Hb�x%k�ԯ�\�Z����T��JF���E�臿ӣ�T��K� q�l�&7�9l,}
�A'�!~���MD�i�d��Ѵ&H��������|�gD�Ҳ��D,vV�P��������K%������P�]!���]�p2�0i�4�*d�L���N(�P��-��������3�Vh��,�w��V��5muXlxVHYEB     400     100���mp�����h�5[3u]� Z�[q�24�i�ۉ*�A�ԯ��k=�r��>b~n�b�0��������n�5�qq�f�wKXd�4������/�D������ ���{.ɠ�����u]��}W�Ͽ��Wq��$�����ȏ$�'1�}>�G�H�GWGML2:�1|ҳ�0n�uޟ�
�pxM�8�1p[t���Ё���S�?��f`'�H�yf|C��[Bz,�LPK�_�B1�xb��e5��b<`XlxVHYEB     400     100E���D��{ꚰb,�:DPT��h���'	51DY<F�7@�6�[%������Y�{N��㞀2�XN�8�F��$���|����J�t6���Ek
BGM��|�����?����z�� @�D�TiJ��
#�ER5�w#�kb]�5�2[�^n��ϟ��c���+���	�	�v�.�A�A}r��gD�b�|��8 ���U,�b�GA��)n�S�;�[?�6(d���g!�,9��$<�"�6h��P�MҤOXlxVHYEB     400     100�=�#���^R^�RwDҚ��x��!9UG�0�� ��)1��c�%'T�i�M��4Q�bq�ϜS�(H��~�!��ί��'d��
mq�Q�;�m5�(?��huA�ۏ����g���^]74����L�E��$�Z[�8t�DH3��i�6���t�*R_%�̋9zu��΀m�ÿ�<�'Z����nd�U�r�2�o�I�_�Z&����{C�D0D��Eh=/4�'^�XW���I'V��m}�:̋<ˁ�p����XlxVHYEB     400     100�`^_��F������Cw������oK:%�y�����VpoӅp�^��K�hg<���˽�R��ׁH��7�x�d��/ٺ�f��}��!��$A>P��� 0վn���
��	���(��O��3.�R�F���'`��Ip$�d��M�s���Y�+�I6::g�wK?���'(g_w�}:Dc�d��+�ʠ�3��M��J6N=]�a��Ne.�U�`6{���_\� �?��u?r��S�CE�n:>��-��$�XlxVHYEB     400     100=�����TruY�w�#���,��0gv�Q|m�"���2Hw����H����A@HyB�j��-�M�1i��c�zM-��dR�a貽�5q��*�%u��ݞ�_�{*��tٙ�7��K��v�]m�[FS�g�y�gK9���GP�����~����#E���� ����s:w��;���W544�#Ip~��ǎ�F�= Qw�$�-�:F��q�6!U�/�@"�xd|�Ʈi��ua�[�'�����XlxVHYEB     400     100p 9�N����0t�c�nG-YB�5D�|.���!x�ko�n�n�W ��	t���'�V���&N�߭��IH;qԟ{�Hˊ9n���Ϥ
h�GD������}���7��v�S��S@�+��TjErL���e?�#��ЊeC7CI#A�vdX��$�E 6N-��`�ϔ-N�%`2�-��Cx��D0���+4dR�2����̃g%���>С(�.ΐ}ð��sA:?6�y�쁒�w�J��0�aL��x��^�XlxVHYEB     400     100Sr"�c�rY^M�s�^R���f���S�)D��2�n#{���i]���Yݭ0v}ఔx��9�2{��0ǚU�gz�|��F g1��ތ��rmt���v[�c7�P�܌`*=����PC��%��e̓��jX[ltYe�۔}K�W7�N7f��z�n;hy�����"����EE$�D�-��og�A6��J������2<�x���u���ڂ�w+�l��y�G2�x�EҼ޻Y���ۧ_����J6(@XlxVHYEB     400     170�`�<T�$ջ|�2��[\������y�/o��wO~Oʳ:�XK��}q S��à�ݔ*)Hg��=`j�D�!:��	ܣvf>oى���w�j��O��D}�$s�⠀�ʁ�R�;�-b�6�$#�	�Y�fOğ�nY�q}�1��_�]���a{�zz\Ǡ�N��Q��Y��v���1p��ߧQ��'Hj2��1�[�wK���E�}�Jt	G.S������f�h��q:�K^��빽{���9�;������E���>���%v�:2�.��,�]h:r��K�����-3㓗#�?Cލ5ܮ_�l��J���~]�B7�F�����B��۽B�<x9D��C�c}B�-?�M0��52NW�XlxVHYEB     400     100Qа` m�s&a�WH#P)�/��dY�T*�9s�:��Njŋ�����i����U��|7i��ڏ�i#N�Q�88��7�g���:�"&�6��S��� �Y��N�=���bw_)R;�c]%��ߊ�h���<�&�t,�-.c;�W� 1E�tob���x�c&��ü-��˥.:o�nՍ��{iM��W�7�y"���:�@��Dluh�;����6^J��g]��܁)���迭5Ȼ�!��/,�+5�XlxVHYEB     400      c0����\W2�/�2�����\�ܱG+P��ur��{�B���	����Z��&�w���sp~�E悚yO!7�HC��,��>]p
��&�幋Cu0۹�\�Ңg�a�K���8P��Ń��>E�EW�q�l>pY�����(X�X����B���u�9�
�<��+���ڳ����C�!��[F���y?XlxVHYEB     400      b0	���ʢ"��"P�$�熭5������ a�d#+.\W�<#�b#N��!�&wy�O[����ʱ¸Y�1(ԩ�+	�/c�6f�r���5�� �њ�;��4Z<�c)�_�������ظKuz���߿�bƕ��^�ղ�s�
�+�N oȨ��^��:��>Ju�uwc{p���XlxVHYEB     400      90phP25�W9�[#`<S����@M!将�������̍�ݕɶ���̅O7�f=KhJ���ـk Ɍ��ՇIcߤ~t�#��F�A��N��q1g]ʮY�#̵���GĦ��݌�����ZQE�YKf���}��XlxVHYEB     400      90\������Ĝ��h��FNĦ�.Rȓ��l,��Z\�Gi3)]����A�O��k��a�J��;1��	iy�j.B�Mk3�������_�}	�s���/o5wO�q�>�rv��:�Ц��(��Vt���j��X �wzDP�����2XlxVHYEB     400      90}��x���l��WKu~In�1����$[yR��rUח?�D7� �j]��q��.A,Ϣ���;�Z!zY~c����B��R"uݍq[�U�:��nJu2)�SV�\T�g֪+׼�Ы.<}Q#,�C���ư��p�%�XlxVHYEB     400      90�*���np�A7��d`��j�7�,�ߥ�L;�JuB�G��r_�v������pvV0������|�X�Aaj��6���4��2�?QK��[��fj	���J�a��;f� ~Ή���68H��%��P����M��*-��XlxVHYEB     400      90����2nx��v	[9������,#0�B��?��h��0�#�AҨ�K�}?�QUKa�VTF�ȡ�9菱0Ӡ;��Ɣ�J�\=�he=@U�����S%Ý����;J�甴j1,�	� ?�/DR?ŋe��S������@�̩�XlxVHYEB     400      d0U������;1.�=��gY�Ub�3���5���p5�-�v��1��e���D�ۙz�a�mbn��,�F1_ۇw�'BtJj��f��h���xD��
9J����`�$��c.�'"�� #��kjQN�䆨�<�N�� �E|�G��WV��ޫ������~��}��D� (e�e[�ޘW��YOI�>�;�C$6��`�XlxVHYEB     400      e0�M'e���D*���6��\����W�0�~ď�XO^�TdG
�Y����%O��K^�����N�YV!c/�X�𔽗m�5)6�TQ�u�sS&9�ɢ����o[o���Ш�F`P#d�H/ـLN�R��i#���_V��T�����c��B�S�4�}�i��F<����	��~�Mۑ�|��V��u�~ʇ^�f�KC'��^�^$L��fT'�)x/XlxVHYEB     400     100>h��Z��%=tY�`�����o~���.=љ�zM:¼p}��]��������њJ��6Ƀy��"YE2��Ib;������?
�)�n��[N\�|q�T�k��zK2���cg>���,JxYK���B5V��P-,�;w���~��ɲv������Z�C�~lk�8��{��XOY��M
Z?ϓ1� d�B�3:-A%���ȧ���=����T�L{�s��?��9�2>�Q�1�Ln@���V5݁de��fX$�%XlxVHYEB     400     160���Co��5�q��|M/��Xo�^X?���\ݔ�������1�ZkP�D��"���d	+��D�*�`Pb�ڼ�����,�>�k����'ꁌ�@����b9��[]���3�r�����eY�Gy�l������^��=z4�Ԟ�4�������4/��O�Ѡ��VU
A-�%n��z}Y|�
�2/H}�*#��[�I\�}�$�`���.a"����ޮ�Ҳsu��tTS�@t��oKn��*��G��6�����t�u�� \��p���cH��ax]�[��mJ���y`�<dR�Y�]��Q1;E����DM%U���~�ؚ%x����X��`�8\��B�U�XlxVHYEB     400     160T���]�ݼ�M;u������ϊ��e�4�2��iw9D��[�Hy��fǲ�9)�����9��"?: �n��;���\Tʦ$	l��Z�S\QzۃJ�
�x�A���U�h�H
3��Z�R�HxgA�'�������f�u�N��y�:���Q��u����W��SEz�̈́M�	��UAt�P�o��I�:Q:W��K�
!�m�m���t�%���ёD�i�xK<=8�?��r�2��9_F	�d?�H�5wA���ؔ�9��߹M�F�f1��b�s�����B3/�h0{�%F�Z�V��~����N�������;t��Oe�2z�ec� *��{���)��-�XlxVHYEB     400     140��-����:��f�<��b�"q�=Jj�ͱ�~�YH�q����t>��A��1� ���@ߎt�Tx��?2,B+tJ�f|E�ߋZ�����i���0�ô�v07�%rh�F'����� C[
d�N��,ܫ�f���v\-
�fA0�������R����)MP6��k^k-��*f	`fů�n��.��<\�V�N�����P$(��c{J�ˊ3���3�Lu�����[l�����f���wn��Ѻc1�{���A��{�����M��a	ѱA���g�t'ƞ߮\�+�K�6¹D��XlxVHYEB     400     170��U��c �N��>�]Gj��8:ѓ!t���]�g%��D�b��֡��e^�y՝<.[�z����6���[`E�g%�$J��O�>��}�y��@t,�1h��Y�^�nҭ�%�cm��Ӷ5�4�����[��\oY�=�/ެ�2�"�AgByH�+B��m��S��RTN}�<b���C�p-�I$�^X�ŵ�Z�L׬�1�"�6���f:D�������ѷ��ny���B}��f��
D��kz���c���_�����t��4ک����3�ఋ�� #Z�ؤ����[Ǚ"���x�b�^ o���7�uH��F��/��Hyx�N�6z�	��y���u�G��偸�5dh~`�9z�)XlxVHYEB     400     150 ��f�ٛ �����Yۮ�6ϾMtEeBI84B^8lz��b<P�]�@R\!�{���ԭ��8�O��$)��J}9�e�_F����.�63Щ|��)�Y%^ԼRy 3�b���i�_$te޳���K��e"��Ws���o����e�������,�z�f�{I�-ѐb�/�9^p\^\�۝�K�\.�R��@��š����M�|u�(��%���Q7���\Ϳf����$+Ze��8MP���*��H�t�����qM�8���jGԊa�άb}F,�b�]�a<��C��s9�H(wbt `(e�
�5�������J歖ʵ���C�a��\�ZXlxVHYEB     400     190V)��!
��+�~�=����Ȉ���Ky��"�y�������ct�a���Fp�FL�����ɐ�]���R�̫Ż���+��7�;%�>'�*����p�Y�����?�"�T�kJ5ug�zE��A�����'r��4�)@:Yc�a���<�X�{��sYZM�쨄l9��t��Mk����bS�*5}����9[�12/@;��:w+�@�6�7�����e�|�Y|Q4=�eX�{���ö[fÅ{��EN�](獠�� /:s���I�Ne�]���n�������U|I0=&���D8��/f2i6����k��'�5G=��t����/�V@�	����0��#K�RGu�����p�W�UM�E�Z�h{_����6FH��XlxVHYEB     400     150��ʨ��ʮ���<�#ݪ�5�^7�pIRۈ��	� �[%Ƿ�δ� ă���9!��?n���\v��u�HS^����=�L;ͲUH��Λ�gpe���9v��7?�b���D��:��5S���P�(�Z��c��gg�L j4�-�:0�X��L^�iv6Y�ʌ�q�L�O�x���� K8��ET$�S����%ø�
dŪ���C�\����)��(��D���IFC�j!?���<���y8��U+�t����16�sR���wi�ӗlѥ����xW鲥��H�����i��,�������r��,$��@(��%'(�M�F�G�M' XlxVHYEB     400     100E�c��LT�κx��{/+�� �s��n�?���&����%bF7��$1~6��v���������m1�e�(���a|ԫ�o�T�E����Lm�"ַ���v>�
&��,��OHc�\`�0���G-*k�������U��jqܫ��o���� 㒕A�x\�E�j�H)���_oN[AP3�!*5��|U�L.�Sl/x�����Jё���C^~_z�`�յ�c��P1zO��:%�.������K����&AXlxVHYEB     400     190��e�\l���j�Z+q��nw�d���V9�B��0��r���th���(d��`��k���[!X�����<���2�8wVCl�:ow����	<�\L�����yp��7"I�|�s�����s%H��Ϭ3v���< v�`��tP�^��]��߲:od
o�1�^7�C���5~D�}�v�ְ���gML��)FR�Fy��H�]�]�Q�����8Ct��fO��ۍQ�
�Q������{d���u_3�(L���d�/�.%���Mq9�XiYV/Ī�S'�pX���D�4(����P�
��%������$�+�앃ߖ�Yi�@��a�*~�ڎ�q���&U)��P�AT�Q�YZ�(P�#��qcUȿ)���s6r�&��� �څ%?�O�<ݞ ��_XlxVHYEB     400     140p����%�u ���$����ʼ{y+�;QL[PqP�����_�l!9�ޜFM}�N��$��;� 6T�b��:��/�����]�o�K�+�Ey�T��Nnj>!��N%'�#վ4�B�Iӓ;r���xː��B�̃1V���N�2�HȲ�.�H�>�ԗ;�فʴn^���g��!���5�B?ih�J��2��k2�Zu�	�@9��

��a<^��(8�;d=�Q�S��+�o���(0[b4�H�u���f9�=�̧����U���i�_ 1�)U>�mE9����=X@�Uκ��BE+,Dɾ����#3XlxVHYEB     400     150q���@��'����l��ȼ��ǡ��� �C�����/ @��9�փ�_e��,7��2��U�����rV���91Bw.R=��Q��˲��"Qe�{�)!7MP;� '6Oc�ҽ�7%��{O(��Q����x&��D���\��4�R�'�ʧ,|�� QO���ދGts��q�X)ːє��of�!my �:p�}�7 ~"/���~�V�C���$:*�R�����������9�SN�X�8𤨧��X3�(j�8���W����<����JD���\�r��rU��
$yG�x,��	9�̊��2���c���XlxVHYEB     400     110����U�Lh�p\b|��W���Ѵq���$S�-�ۗ�9V�6{��X��aw͡B6GMx��F�T���@�T-��������HN��5��F��Ę���k�C� �d��]DU��� ���Cpn<��O�!@�*��<�+��O��h��r�	 ��4�}b��PP�O�����u�u�*E��D(���Uy$UD�Y\����B~�X������^�'ZTU����6%!��F˹A��57�[�*�i�2N�|`�V��r�����
XlxVHYEB     400     160�m��=��Gt���h؈��x(��õY#g>�/5g&��D�.AkVp�?�h ��@E�y����o]�;h���� 5ia���'^3`�&��R�l�t�a@����5������n�6DW10���R�ګT�u�9����?�g	�b?��A�ﮧE]��R5	)Ǩ�M�fr�8S�{yr�J
��o' ��⟓���y(v�v�}��}G>ǚru�r����¼x#yT�=�"��o,+��FX�R��4JQ
����9��;����1ߌ�u;�t�����]�V���<N^���dJiJ��I��q�M�tb��1����M�>w`ƺ�M��#!����<3S��F��p�XlxVHYEB     400     160��c�jdW�̽��AN��������g��B�6B�/��� 1���vй�X̨~�uUnZ�Z&D��^ʡ���f�n�~��4 �5�J�NC���,!C�{�ܺ�L�s�Y��9���Ch�������5�P�	2�J�+BX�_��t���q'5�Eh��M@Po09q�ӄI�FQ+���
�I�[k6!�����鶪Xp"��/@$t��2�Ea�X٧N���6~g���'$�l_�21D�kڀ*v�+����{�)<il��^b�{Qj>�Y�ߙ�Jl���e>���$R �-��wJ�$YA�\�@�v�`(�jOb��=���¼
�j�w��,b`����9X��\<�XlxVHYEB     400     150߳���r��I�̶��1��DF[����'� ��ӝ�'����Hgl����P8�^�`��(��f�i�M��8H�,�dF��b�c|"����fl#6^�vn,�o� Z\�r>���
n��Y��)��(��
8��X��7JԒ�˸?֫�⡪�^��y�G�_`d��[��R�  ��L��s���� �
�2�aJ�8�z�l���4S��\�We�����E+%��
�q����xa��.�㓢���,��ACo41�̓6|I~�W:�fPax�K�uw!���[d�	�]/q0�-e�y�O.Q�tw���\�Mq���ʹDm���'0O��!�u�XlxVHYEB     400     150TK���w�.x�탈�� #p��3�Q�VE��Ծ���,-rً�Z���Cm�/2���'�$�Kl�3ԂJ'�z���t��� ڜ����t ��U�2��Q1Sp�j��H�o����x�a��,�-�P�xd��fO�ѩ�'$� V�����|��v�
�| �x�����*J���c��T!����Z���Rg:�05&�;�|g��4�7	*�p�G�Mܼ%�᜴��ϤK|n#>�c���H���㪽p�I�%�Rf� �EG�ϔe��$m5���C��i�?_�y,PfI��%%�>���2��KF�O�bm ư�W��eA��XlxVHYEB     400      d0r�"�Oz���θ��� ��:�^b�%z%��p��B�=ȣy�o=���^)�f�g]��E+S�ŷ&�5Sd��0���V�R\���M�?���gx�P��Yv�
>��\{�SlC����pw"�v{�5��Wy�|��I[�_�<�w��x#�ny��J��KP�I#O}d��a9�s`���tO?)�'�Ԅ�p{���54���Cd6SrQXlxVHYEB     400      c0��<i�c:���� ~�{�64���
eu��{2�	RqC֚�e�*�~��g�?�� QT���Ȉ��azʉ�>�n���'����&��=��cv��n]�2��N�4�3��9������k����o��fȈ�|o^�c5g��iV��4����l�cF0ҵlpܻ&s��`��z0� '�A`�SXlxVHYEB     400      c0�/N"�8I�^�k��Z	0�Ni#����b��܁�:E1�g��D�D[y3{Y�Ex�v9������I,V:M��mE=A�H���e��r����Ժ�;H�����\o_4[�J�̖J�^��(
�Jϻ��߽�n� �]�f��d|��o��_mu5�\��z=5C6r����P��sXlxVHYEB     400      c0�^m�=X���Z�n(��0��0?L�0/���#��u�h�)�:�iW�:���Sr�ҽK���4������|�Ut���[X�cO�{Α���ڦ��2C�U��k$>���r��c�,`�r^���nPAR�U'���Mo��uV���Pj��(kk���`W�e�
�0W��%d���b�䐈�S�}�i^XlxVHYEB     400     100T41�u�<a6suݵ��~p����/o�NS�ʹH��Ch�;64J?���ﴐ�n��JmΣ�"�'F���	F��Z�U{���4��&k,A�;����K 81\�H��r-J�hw��-v�� xF�};�����f�z�t2Atz��Y���B�v1���D.��Ǆ}?Z��3�4}Vԛwf���d:` K)`07�{�Cef3Mf����H�{�؃ɰ"�1�I�_���[�y�=��ԉ��D�NWE�\LP*�+*�Α3�XlxVHYEB     400      f0�B��N�u�1�.
�r	�i*�a���2�-��.�!����l���c�1�{S���������*�⌼�Lu��66�:Ϧ�Uf�r������㊡�U�ID��%��Ʈ_�tO�gU��oz��FbFE�-_g�>���T��K���z��
h�{�uEq�v�?����Eъ�ۃ�&���x ��Y�t�K�6\��Jq^�:�y����u�Oc�ѣ�$d���cI��m�oBAuXlxVHYEB     400      f0�#YZ:Z��x����ڇ&ef�G�`�E-���RG~+ީ����d���Tf"%���e1���N9��W�.:�y�����6�_t���|����:~��/�Q�K+jZG�Л{{Ɛ�"5�����~�9`<�ᵒ�ݙ�0-I5�܎d��}�J��	x>I���q�k��ٽbū�2��r#��e�M<��[����Ǝa���G��_-�g�B T�;���J��t����B1��1�q,VXlxVHYEB     400      f0�T���������v�zK4� �c����"��x����ӵ�o1����"���"���3����@�������t�G�e����g�1g�c��I�9S!�U1�g�ZO�y���\�V�"ύb�M�,�LM8f�,Ne�NԣǛ��=��s�G~�~�	�wǸ�i\����*�M7}"�/�����h�y��7G�ϥz���H�W��A"y
i�"���g	��ԇ�1m�I�����Б9�6��W�q�XlxVHYEB     400      f0Iu6<;�h;��'DB\���9��:y����(�+J]P������|~HV���H$�5�e�6�j��}�o6S9��qt[��T��p㾻4d����ɋ��H���Cۗ���G�sƸ���u���vS�¶|i9�&鹹��T8kC�C�s*vbh�9T�k�M ]������5E�Im|!4�Kp���u6��ѕ�l3���QJ��kį��(�����d������e�o#Q&v� XlxVHYEB     400      f0�3��5��Z�%���{9	a�������o�m4���q���ѕc2ؤR޻)a�o*yN�E��iw�-f���9�& Z���[�@*�q��Ҭ��Mù+����{�Jţ�i�
t�C:���sT��!�-Y�
�)&I�v�b��w�2zk٠X��@�D��#�R(gz��A���5�v�j�@1����k&�ud����D�fh2�y9�7���d�3W�_�ܛDr��9qwh_SdS��~.�XlxVHYEB     400      e0e�5�o!�� �ϩ�C���_NqjָnT�����juo=4�S?n�%������Yሑ��r��YCfcQ#��_�p2���|�Ŏf��g'jC��c̍s�:mkd��?&�+����5IFbu��l�]��Z)�EjM]i\�2��:�g��|R��U�P�^XU{@��M����Y-תǏ� /a�B%!d��;�ny�%c��-�"`$
&�w2�t��XlxVHYEB     400      f0�G��^<�����VT8��u�M	j7+*�4ڋ4s"Y?1�TE7MM:A񩕯�= ��v���
?��^Q���|�+uq�n'��Y-s%����������{�NU���d��+~]�'O�)7���]�d~d֪�n L��uKc��4"�{��6}���E+�Y����P��dB�
P��W(~a�C�Ú`�"y��\��(X��s�އ�@H?�}B���)k^󿠮i�XlxVHYEB     400     150ͻK8fF-��3I喷��_K^ ��G.�f��_�����L���>� ~�K4/�mC�䐌KO����Y�R_����xX
o��}��Sw��2�m�*oݓ���V�C5J�l���EA\R�W��g�䓳�$=v�nWąܞ�i~!1�UWA⿝�z�9��I���L�h-�)!?{����?!�)EK�b�3���ќ�`�q2.�kK���GCW��s�r2�/��i�:�&=���g��*U�M����ǮJ�dه0��:z� �D��]p;�arV�@���v���q(ǣ����e�͘8W���w%13�s��b���_A۰#D�y���mXlxVHYEB     400     1a0G:u1'���P8 �\CO�E���3�9=MLDH�V/JJ�̩�J�����M�s0�D�'��oлW�N�cg�cT�娇�|�k XSCy�ެ�
��DH����%O�8��c��	�uY�	|��ԗ���l�ĸ�?�_��RN�mr�w�*I�\'����^��=����ozRz�RM��?�j�Gt2� ��u�R=� �B���}'*���`')V���� fU�5fFϓP��s��6��69]��CQ}�l
`�va�kd�����S@/�R��PiR�_�㿔�(���M��1��2v�B�#�������b@6���h��M�i��P[U��%�}"�Qs�>g�DB�~fv Fn�D�/y��4����fI�W����4UtYe�*��*�x�c��(F�wx��'�ڼ�{�z*x�XlxVHYEB     400     150HLt$n���;�Q����ڋ�n��p��^[���ىw%,��3
�
�	,��i�"_g�0U�FB�+h-�E]B�r)���JFH��p^��k�s2��]��r�Y<��b'(P&�l��2=��k����ޮ`���o���?!����g�`<����̶&�k�-bb|�wɝ��H � �RB}��X-�i�B��k8��=���\D-�a�qN�LƎ("�˧��u��i���+�!�.��꺇��/��V�-1i��zJ�1��kv5��,J�ל<[e�������ؚ̬AcݭBR�!2�X9Ɖ|��r�;��V���/��D�:}XlxVHYEB     227      f0��L�ŝF�x
+�����O����/��4=ȏk���_+�B�J�SW�Ae����}��r�p�i^�?��V$_���u);x�T�~(��(� 3�Ǌ�w���e?��|I�����,�~hELF����۠
�#����7�t�>30!n�P�UT�����YD��v!(��"d]�#d�6�g��	����f�3����t%�����EUwTk$����.���PS�������<�8