XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E�|Z��MZ=��4eN�FY�(r��C���{5
1�E�"���5iKK>��ɚ�>Rp�������:�ե�������1 k��Q�#�yK�T�Y�z�3H-���,�B�[��/LFU��d-&� �m~�O�J$G*���ٻ��yrmj��,�I�MT��9�y��<�Y�=/1���Fd��i�8�M;�#�5m��
�J'\.H��YŪn0^i�D�hFI�V��D�SR���ѯ��'q�ե�B���_�Sma����_���+�rL��x��ۚ��2k?��PEȢ�cl��:��4c��wU���DJ&����{*iMF��}Yu�)	V��9/������7oH�u��4(�Ey�8���6�Q�>,��_���U/��}�N^�&*��$(Ă�����%ύ�F�%�}Z/���n�t������w�2н..#�%��Q���smz�	�?Q'9������tzț4'�*���I2׹�[_�yd�&u�U6/�G���3��nR`���3�}��
{�W U!Hkn싰<`iq'�^^��I+�e
"d̓W"�2��꺐�Jٚ�=쎞�̝��M���1�C|L�rsI���ŏ�ǟZ��h���m41�Pw��]�T3~U|1xŁf�{��/[��yV��������.S�/�@���i��e�xw�PM��):{T0�Ng,����qL8�W��`![p2�H�u�A��� �_l+�p��-rz����@rP[R�����<XlxVHYEB     400     1e0BG����&�W�c�l.8�2_Wld��G�1s�܏�vԐ�2�bzF
b������ʖ��y�C�;�4F)�3��AM@w�I�\��8Ӛ�,Ug���k��/����������Vz����LN�j�2Z�~j}QK��0�9�B=�^'Hl_Z�f�A�1%P��:p�L���ڄ�d�&۩��;�#L[=����+f%���sBn�F��!� 4���}���ɿ��s��ʹ�y��`-j��[h<����kbSd�5Nۡ�}������/��*�l����s3mt�U":&ԍb��"��&����r��w�B�/Ѫ�q*Ki2:}Ֆ=�5�r��f��c=~��� �qѹ�|N���V�Z)����� �aA 4HT23J��c�7�QK��O���>/�<`v<����84//]�T]���fɊʦpz�Z����;��D�H0��;�Fu�f��ȗ{[�.8Scf7�XlxVHYEB     400     160j���
���G��Zj��Ů��)_�#Q�D�}�U�^�ݩ�f꺊���{\b��(r�
��Rg�a���'�=��E�����R�;�*$��
D���$/���P}]�ו?��]��t���m=�_�
�b9G��<��ˉ��M�|�F��砹�����7�4�D�,�s5��ׂj��Ƈ{n�P�i�ŷ�!*Bz�i`Ǉ�:��2�"6������m�����w�=��~�'�p�ޓo-=/26aFu�(����U�[�Q�MFqI#�9�f�����X�#�R�%�*?�[�P�x��#�� x1��ovRV�@eB^i�L1�q��V�9?�'���Gt����XlxVHYEB      50      50��b{�coM����Yg���XGe�M��@v=�.n{��!�50vok��)�-B�O��l(�q,/?8�G�Җc+�`k��y