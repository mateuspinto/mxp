XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)�K�Hy� �����5ݕaɘj�=G�D�8�sw��B�}mt�%�U#�eI �q��^����G����Jv|Ċ]ޡYy�u^E(��v����|If��y<���H	��W���E��,���~b	��9ͤ��N>ؚ޵�ńJ<J�1J�O�1H+9�io�u	2�����'��� 򑠜�^�s�۩MF���������`]��] ��!���;�{Y��t2�\�5�^�,��W%�!W�c
󚴱$WA\���L0�.�cL�d�+E��/�W�G�Q�1��e�[a���"4��=2��d3ZZ�VQ!��o�D�
�F�3ў��F��:'��?&��� o��2�����4js���_��E�&Y��J�1'��=ne��\d֙/�.n{�ܶAQ9��4�NxƱ�`�O�g!!^V0E>�č9��N�U���SC��T~��_��M Pw�N��ڍ��fP��
�1a�[b~�b]�C�O��S�-�¢��VX!;i7]��=����|{�h霙����e���)�}G��;y���=������Z�K��,��g^���~KVvrk�r�6/��<��v�,�26�:�����ͱ�ܰE㞳p���f}�e�i�GC���'�m<��g4���5$wd�G�>�J��w�K�I�"�=d`I�OEa��F�.$S��a�Q��7�7�.�n��B�hx������QQ��\!H^��:Y�y�_;�._l�T��a� �Šy�?��P��3f<"H�9n��o�XlxVHYEB     400     1e0��w$��+0��m5?J��i�[�TC��*3�E7J8g��$k*�DjJ��|-)>׉쪛N��e���3 Np3�'j�7�#}��4��+pX������D͂|w�]#�ٜ]��n7����NZZ�Z�"B�R\XyH/�Uˣ���Ѿ���U�Sg�,���`�gD�����F^;!�XM�M�#
}J�伹q;����بn���dӀ'�(աd<l��=�s�H�QSl.��ն~f�c�fEfy���g<�ÐB���}<O�'�G� ��w<p��*i�?�Q�t�zA�p��7}Ӂ����$@h�qcKL�� (U�u��Q�];�8�E���P�j1��Ԣ�_�6�#�'?"kw��6��9{i���W���Ïl�ڇ��4pЂ��W]l�Qx׽*����u��8���pȆ :��]"	��Z���!(:Q���T�A^�8�gq�fT%H׼v�V5߼�J&�-ms$=��~�XlxVHYEB     213      b0��F{�븜f�����ǯٳP�̜�n}!��]�n�-�.�{58��|%��U���t�I*��.�8⪗q��^���M,0W�����A-����S���c"wmS����%42s����g����="�>KR��"�+kҥ�"\�Bb��@5�<a��j�$$��/nC�o ��