`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
b77WwyPVSKqxXg2VTzfmcYqM1+03NMST7yHOXRdvfUnNf2DbkD3sYJlbzPTW6ktN0//8kTpFlktG
vIxpMQXbci7IU8uZooiu6lBrmkUHm68Euh9qzEYUZXs8GBtAEa4n+R8ZHFgMGfVDQapSVa1nTP+D
mEFR6LSFrKdd8m78VxAykhSAF2BJVukP0i/Nrqo8pGwiy8UKVcJabdihJ2Arna0iAe/58B8BO5AC
PUuZDReCJvMP0K2wzVT8TvWGjpOG2u/qqOUJNJFHbBbtVCevtOkA/au+mE6XNjw/R2kaZps3PgFm
7OYJSQ9YlOtUjtncZmDDKfdAvMGFSra6qMhzoQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="YEb0C4X6B6l4Uz6QcbQ1Eh1nhCzfUEj9pMo56kd2fDI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`protect data_block
kzo2rmbj4xCupzmQKNJhFNCbTmOdjj9DHic/6m16RNNf4sxwhIcFakIgE24kQTFMczIrZXacqVFO
N4+KLseXhYwnwd+Szxy0UrNb4//ynr3GnrPgYebqXaZip0Z4bBHxj+bCAojfFPDBOaTh5lzfzwT2
VFIhmBYW0r9UZn+cZeE4pIBw8mfYIsf4CvwQvCKLmZi5GlqPmSfp6PppSF03ieoAftpjU4tfUx1M
9k/hVuUe0q1aV2HP7tRMkc9bgMSey1n75zUSYpHSEQLR13pr+qTyCXvUTf4Ax0Yk0Eb3txY94uZP
GkHy0nCVbyv+EC9KrMjpDgK5QPmC2ESdQCMIYwoaa0Rt8+BqJNtMCwhjwM+RfoLs4kZZlXXNMIrR
SyRCKNknHFVEhhN6lmR57jrWOhpT5Ph9pHsWIiT5E3Bq01hZk5ZBrVO7KqKX39to0Vh1INwtj6GK
P/J08XrK1SqYmJRuxXaJGeR38BxaxCKtE3HBVno3bUR5phKpgdk0t0miWru66nef5z7m0FGR6UuG
WPVn6EZ+3VSe+839A5H3p4NlTNmUu4J021Z9SoOU+2XiNxhit+fuZMzBahLviDp9RVZHPTbRq2Sn
RMahLmb+OnNqkqF3/NnuoIHUJmGony1WGujH3B3X2j+UdWSuca7FCTn3gqU+NZpAb2kj2G74OrpZ
kTc17+HwdqScvfd1moRDyZUZkv5MWLvmRDNiLRolka03yZF2dZDWJQBLoR26oXhvXuHd8a228g5Q
iN8ePG5YnkkUqLvufW3JcoMqcxPkhjzAU6eQpU7LnzeebnhIu+PKSL8ZgmwInqhoVQf9kRyDk0iM
/fEh+A/eemYgPvoR5WMB6C1cYwC5ij7Xst98QIUwXhUqu/+7nwbgMkfCCFCbIjPHLF1Yl6wm5vZV
lsWDWdF9ykXoFNwssi3Z71ElDq1hyyuHsyyeNm2RQ2HcRPWq+s0xYYXuVRBt/jtpzNNGpV9il5xD
N67nAf7TtV4PcAV1gqxhzQWB/QCGWQWz6omDunx90u0oKtlSeRNx1yMODNDClKQAA8ug3tGstfYL
Ggz+j7Bn+6mQCPzQk4GbGMchdI5t464hFcvDoYDf/Cl7O5s7pg5ODyRHaNp6oWQoKHTyoakKfBt2
CMQ/tgAeBkmXjlDmGGwdo0V8oiTLqUPbZ7jwKQI1ds8vHvgaCEHIILQDRtDnxZWoS9P6+dmDGNV2
8bTttWsdbAUML/3P0zev4ksvcP79TbHqbtpNzg2F2x9GZfDkYC2FJK7/oduavvlEMESwXtIZdwRD
po2UBGOYN8224mylMjyKMD8UulQw9O+l7nKlvM87ZuxlONL96U+V6c6PtdKssZTfRCsyYyezhaB5
MGrwlBWmVXPXfyUZEqrc4SkFXBsNhyk1CgxVmChiqcQxixqpo1pDeaNrhSEnPs4/zMc8erAxDNpr
j1p/hBQWxhX7VGanoFn+cGd9W2vjgQwvOgKj6rmWDaqxblPOoG0F5QMajwP3q66mv9Cca2uzlGkK
sesOCxwfpzYf45/O7PGEeQd4rXdpx0Jz7b5MEGINaWOFWTKckWeVyXgMTWaOf3qUoIhOZdouCzti
gtwCJi4Evik3MqMbIPtEWvooPM5fjS4gBgnCp/ykygMaTcKAGDYO2dIviqk7SjeE//ynQ030vftG
fx8j+/J+lsNeqEfGm7fLvt/8ckRnNEQ4+zSDARkuNDAp44jW0kpQTXchdU1R7vNv0uwih8MXogUT
8qe4navTUFdxvcB7SDgZbj+iC/pjncBegrM/CC32L6k8AqSl5aWVocclEgnAeUrP7k4A2L6mIqr9
pa2b5LXoha6kjCW5wn/p10/aCgWbfPdNn+sUigdE6jJU2o3cielHPJSur4s1Tc35PpYyoeA7zzvJ
gS61BsD3reVSPUnVzB/8J3YRgP+wZ2iwbqy11OFrxkfw3mVvY6JZwawVbOjXsq+rJFCWwwR1ZpQA
eh104bg8jUCVQBBVZGjwJZnMGSnN89Hi83oP64uj+lYO6rJ8ClCGMHQTPd3/cut6uUqGFyiCuCDn
7APNGxM8+kvKRORF1cmM+FyV2N10nocyIq6E2TdA198TKjnIMDcD73Qr7vom7/ae3OAd73kel7IF
IcJuPMj02Har7aLFNY2XaMT+UeZxMRlZDJd3iVD3BOP9S80dz/uPKXtSh1bZgIPehi1i3+c1OG4d
Dkym4R8jlhO8sAlr5zqRzg1E8jMsKPDv0uvLPQCripDcIEmF4YBYmVsRVuC2Ue2MvZyjuqdEAOJL
gvd5a9LzPQornbSWT3Pd248yDBJButqx1AkIbiwfZIOVAUwzhZEPu69DXme74G+l5veNaGdgRSoS
5TLkRtn23fDpx7ZYzinw72oCaNVHE9TSX7nw2ZIk1FRAMll3oSO+M8P5xQsG7RmkT6yD54iBonjs
Dg3q13AsmeBF2OBjhNPLbbRq9RmySHIrpIiCK//y+2JUn9mxLYKzxWMsegYh2snij4rzmIlJEH9k
bDCPJUHdbirx6WMVTdlxgdIO4mP97KB5w8iLiE4Q5FSxmfy5MuHp2H+3ou3gX3vgcirmXSzHhHrO
j59UqO5jGI/JQ1UQ6XFBGGdybj8j8WYJuobLBHlS+KuzP0OM+o5LxifkNBxDgc/OZOgYUDkcBS5D
YvQF/n5YEbqwQw9wpW/Db9yKFkrvyr67vosFdwOZz+UPjbSyzVYO1T9s6cI54rhiW4L1VFwEuVSL
SzAypYF9ylMAqX7a9q465fjmZ3DfeCdRsLBq8yFClBp8RdZ9GRrv5EFb8Cd7p9rjlo+SFG8mFbE7
F0E+irfXxcAbLnc6lvMBqfIHQw2dMP+eGOYjTCxkLE3wysHbswcujw+AZmTCKe67Mt4sGEQbpzJc
tZGBEXN3+bH9c1SAg6x+eEHlAScEeY1mlVBO0lsCJeRcAbCqh2lmd3TbGBoKTnQW4UZNZ+bGEYPx
PpTu/UfkuuTh2GIKC+SOLc632OmnIK/cLbjH0oXETjzVe/Z8+wPhEQAU5G9rvDF01uPOF0hHjNMP
YBecaL6cC4qF23rmVyE4imc+fzCFxzpnF/X9J8ijx1D/QD9kBVIvBfaOrfwVZE+jzRShrhOnhY2I
GjVbOyrsue6Z29/UiIhcG+QrKgiVs7aoGi4DzH9ypZN/NeuZsvmctXwNBPbPnm4u97u5NeiQZBgt
47WrvnouYbCgM2oJIVvrtSyg3ysuVKC8FuNgXT6WCC8Faaqh8nxEYleHa01PEQR7PvzATIvhZ4iX
0SzsH+IIuHsuC8g1TtVOE/JcgH0W01LzdlTFCv0QE+sUabY7+NVt9JZQzQil/c62yaq39T141Wpf
oAhqG2MpVYjRe0iqVpmu9mB2TTYKhGwjVjW9LBKjJXr/slaZtuVgBIKbCeCggYI5My1HLhfBiPkw
IHGloz+eMQ3EB3zAp/tWMrL1g45WUF3zkriBw01NYF/wu8BxJVWlbw+QH6I1IUb4YO1+rbb2beWt
EqcW3+DN9wpzI48KtWUZjOg7qg4D3d+wbEvW87eJcc6M1AYty9fqmh8CQrTXMi0SE4eYDoNh9Pge
UklEOUXlUOdVFUcploiXQ2oUEf/Sd+Fy99xoD1xhxpoXqqs/azIBS1HSzRRaomdivtL87b0haR0M
KDhROEH0IhoyIvM5orNZ57qi0A92/BzbbvUjRPS/w69cNtvnf7wOQMtLN3yAv8ahSnr4zWImM3oD
3Hx67WI3OPC4xvqIC8R4mucN3ZsFYKNUz3zA8RSJG7e7XAzpkjZJ43WrZVdZnV+NctNt16VPesDo
UXH9ZycSASknsfG+M3V/eUvXE9BDsKivKRy/a618eWXnohQZOOuFJHZwRng/fr3b83Rdqe0bOLVb
KbyxGkoHDEQGT+3Ez0KRz4hLdlpNvaKGEf3RRC0OPRTsH0T2ekxwT59qMeTKdqp3vhfX1vDXr9aP
qDuSt453JUo35Bzk0reQkN1eXF6T+SQQEURYprRUTEKKt5gsTP4OZqps1M7jtBSicbKkM2p8qEwc
MY4BVtvIrt/a/1l9td0cb8gu2daYcDTbG8HJJbeamN/w9GRjWT0pWhyj0wwxAbCVlzTMy6WsBnwj
LhIJWc9gtrqkv2zFupCpeJbdjVwR1bfT9kDJc+ICIvkths4vySTYMxCFdDah4Hk0DS3NzMylaZat
rMrGJSsTZDl9NNfVjFmYYIUlLcSu1tA7zyiXFcuiPE7vzRs4yFq1sQwG6VCXkmzZRhRaETCwu4Og
Tmib96NqJWqRYgJZGIaguUSr1SUnV3muw0lrYMKOI/XxYtTieKUGT5p3xd9W6SSsQwCidMjyyOm3
3ft7+xtHC7yVUc1+ssG2lqyZJi5HhiRqO9jw9aCGv+kJTZtZVqtaA6EeG9zSp+d5u5quIffGJjhM
DVxlbu7G4RMXarvW74PFJGKp96ayc7mTYYXv66LT2hd8ltXSRY6qkmTY8CLVDZpugKHas834aWNz
aZB9bOYtvKQDAIp42WQerwXJJglBHwJFVyGIimd5ihoTaGU3+NYK/rQvUX1V0NuVIW/iWKcRDwhg
p10khje88lMbxBn7RajfMaccfsJ4Zb7w/DxEgBDJJfv3uDGLn73DX0mStvAsUtxv9SCMFDMsIkCD
UEwxKBbOoXMAkL8e+Vesn8OQiwMPHTklgOhtPMQKTabiVKKi97IlfMXAOrDBFGjpdi25oMwDD/ak
v0W59r/i028Cexm1Ri28giH5akPgNFF/BuLcje5ifDsHq917gbktqozx50koIK9S6/tkyk2sv8r6
n+Dx6o+LMmbKWZKOfBmInvTsIQ8HzCGNRBkwnVYiVmN68JBsnyQwVm47lu+Aa0aQnmqQEVriq0Jk
y2Oz154l8FXMehMyd68RwA6/a6aqJoQXMhzHItaPuyqvFM3dXhwE4AFnmBbb2PExhI1OlJ2AKxGP
BOCkuNR9XVZ9ZaNEPPBl23FoNuEy/FBW4RaLzJtARC6P+sIVnCHlWg0J9tmjqs+JNvAtrLfHqI1I
d5kgSD0Q05qtCaPKJRzDvNToOCx3tVVpVxshzGp83xy8rmkdhZet5tm6FkGY1JQku6uBHQUA+hkZ
XWZcBidDz4Re/WDwcqytwozYjlYPTQCt8Grt8yWkMcZM73+ux1R8SNzDb2dnnfAmAxl1iAByQ0kQ
hTlRzbZoV353Vsrr0A9KIhYAmBr1TFr/OsHRDC0ru1OPLGhFjIzc6EMJfQz/Fht7FbMiUZ1R7VhA
NZELAyMm2gmZqrsuwdF9zrTyS2e7sDtajO+DU0G08n5+43fVwXom+YGONE1mTOd5xp2kfaF347Lf
Uz44+/7BGtAxSQWegHnOp/HyRoVq3jLtwJd3/BTbbENzZo/sl5X5VtaMTvYM1zbQ5nN+3d76Vi0l
RiuhLT4Ei3Wi/He71S3fogUu/358DVA6CbQXT2tOxQYauP8Ws4UqfibOEeAm3PKVs2NfHZipz1YX
vnuTh88OGSzX51HyWBZdZaY2xmaC15EEpYqeCYwhkV95HQgxPtbi6QsJXb0vvIy2EQnUZc9EhL4y
wb6IP8VtMOavsUwqby5YuYbrSXzFxtg9BxXVjuRsS4DCREXhYUOZ5d7z/9NG0/AREU82oqDNEFYr
If/3MP53KNz9nhEiGhASGwm7awYUgrRY4Dy8WkVv0JdnuFQzYMMZZNf1EwjM3YvfTTNpUjsLfW8M
MPrQaShH3FtXZ1tTXMp2nPGnyR4NZMqU3fjr4//2lTaKDnEp/UnhUgUQEcWPIaSQ24ACK3EB3F2p
bEaY1NzHFTugCEspHHq0xL1tuiEeNLwo4oUL2o4KXwIHVcYiHy4/P5FXXVqUF4lOQjdLCqVGN6Sh
BkS6IHePJFDp4+M81tOn8KA5Gm1M5VPW2PSoOb8Ie6SMKOWxBfE0mrJ3gjHwj8tI1GSdBsf68RAH
2PTNqfm83IcMmrdvn85o7Jw1ajdQ5EftuLF5L89zLoVJ1GhIQbkn5ORGuT9aOLhGJ+dZO6c12YMI
azBui/JsnkC4hL3uI2VB2JycJGTpEFoLl9mcR5pK/OqSj1nYcc/K1rZtCtcea9A5K7MrOF9iVlkB
ltS/KP5gdZdcgjGpnRnXV5VGF8ZfLCQggsswFqENo/DXWAYoudXrRrRDL5XLA5+r6alKR/DB5UHx
03Uv3OVyeqCT/HPHK/jIX2DT5AaNvMQFNGix7iZomJN2KbtkFvZBUKEwBj2axxtOb6x3KAW5fwNZ
sHXwHAio2zQmCCte29b8PnuE+URRQTJbq0pjCDjCttpsM3l8lM8l2q4NelBrdVb0P03z9cKZCP6y
N8qW6PmC15+iSYMkAkr5z8sYGzQ9b7CywuA0X6qSNZouPlI4BFBRvA2Iv4Tz6qClJcGteJiZLHta
hta5+z/CGhigD/wH791sxkuqjZ4pONro2ci1zrJYw2AMyF0h2QI+/JOwBR/dmYuSiLSj7UZx/cWC
SvnNWaBh96sSLVMxvoUDg9orOC2cFR0fjqq6oEXrpIwPggCKSDqaeU+ffaxHW0ld5iSbpLZYiSdv
BLviHdOfmWkqNEMZilkBNARaU/HXrIBe/VSPVpbinwt2qiFZscSTwQBUwWLE1T69Qd66M0b1FAuW
UoAd/4a01qRj2xe54jeY7Tt2xAU+h7UI29emBzj3vIQOdOBG6LopGuVo+uAnLdR5xTmOHl/8trqB
plyHILr5oqnbdMZ8LCZ2pfja16rFA6Ly5JYVIHLRilPL4EvvUU1bqmsE7D9zfUivHPDL2W9rGJ1I
2srxKvoujxJ0PXHrlE20NHVqaM0+6IfruBzjhSWjHrnqgtOaFqb+tGyMgf5wfrd9Bjt8qzHJZYUy
8kLNRhbgHHaRLpvpD/g6A7+wzye6MSNSxh4mhOoJEk9GIUAyYAVhjRhtsaV7YNUL8Bsn/B7eH0N2
FI/FNyZ8ugqZvggk//+lvDbMf1QmhP6Hd7onKRUsjZA6a8+/Q79EHxVuPAFuoINeOqfqhjcQcDTe
4meMIDqV8gdnVO4PZr82218DRdbzVjHJ/w/8rOIn4shXvee/2Is9jsTsFdRKG4KqJe067hG/twLG
QGccsmLQHxtiGXu+YCPK7+EK60oMi3LxqOWSmfW2b5/4ZxWtELcmJOUgAJJ1IV4SVGr6n3GBsabf
eOv0kUqbQarsVJqlO/GYiFMmXWqil8l7yrY6+WpcQkd1n+yJ7k2p9qguNnjPOj5cQ2PysPp9BN8o
Mb9v7agzVToJ4eWN1gUQfU4qWCfU+irBdmnHLRUPNnzdIxFbgQEotk7FU+DSdgM9+sy5afyD3uhl
zJaWBK8sVvSkfKF2e9wXH8g21xg1DRnndYFSyJiPn4JPw9Cv1lCMYPt4H4DwkzBAiRaxJqoxwrW1
Br5e3AR2Coqi2SRMxkaxDBwTs+4Ny0+endVsXCnI6ZFDSZSVW++95Qna7LujEytKniMNGJ320PPa
5bLdac2LolmkOrHpPjxeAnp1e9lk4LR1FrVNAYgowBkLXQyDlvBpPSRt/eY3kMAuyvCBPizTa6jp
CMIKrXb8rsamZhPb/QH98zUM7QLOfA0BdemMdP3WLYc3dlni3uC97z57kfv8OBfKy4urKRD2Vxtl
jQqRvtFfchzvoaCznM5oMy/s/XAHLA79eEa0+fMnw434ksZxIef5+sVfJIwMxaVLUQBZsds0syix
LEAKdgEqLk14U9NLgjFt+40auf5z8rzdavCt3Y1KrQKfgPHl3fCW8pKQLwXU5zte3O0xGVDsfutD
paEC6tWKich/VCIut0aBTHUcjArMUwsnbWnKkdUQ1m1Wlk5mdaTujybPfupGfKu5CrqoKoWhqXJZ
77PPSnN98dKQt4PBGSwUdF5UEwRxwKcpfm9hp+SeRpAVToRNGU1Obexp9Tgd0FkMIGH3AOWntKtG
jKAC9qPGX9OlByo9ASGO2T+mAGjwMcm8jvlreb3crh3SzZ9UZ7xLgIqktyTuekR5nPtq5twIVgov
i3sqCsfSE1zdkLj5NwO3P1aVVitrwZeRFWZFjrHDvVgboM6JGJ/6fXb1WpIwzn1r83ORpA3DVzhE
b83NmYIh1XgMqiydyiyU3UGNodNgxO7xSWgZ9WmhUZonwSbEOFkgl8uYvcUrM8WWnXn4dMW6Ew1p
noHpg8S8G/aOKRrEPqaJvMAjADJPMjzXKmnBDwVfbDAf6tM7+mg5PFKm+1bVXYQ49gfwPQDm4MGf
ftxHl+GFVXKGizWc9WMiOhiAqsTLvILreu2wo08qlA+vILtdMcmcrjwnnwIU0kQQuxE+Tkvyh6bL
3t/1Icki/LuaJAkxcqtpnoHgdviQuK5F1fDQf8RONGrLSIdsKqQ3/YMAia9+ejNBoaS2dgZMgJYZ
lVUqht2R5mfafNWvlhRqMEQaVfXB6y1Td4aM+TiVWMO/M7dNPIRb2sEQ2AbbB8xJa3BAOlHGqqS0
rz/ywlZI8L2SX6dML20oVwNeW40Yb6+RphaL/c7XP7BvuUoDI4CB28QpkYEiOYmbTl+v0V7JYKQ5
4mtkizg7/yuxvEftpeOQTb3kEJhMdao00jGvwdKaeIqGpGcPuSiXMK+T3cDvnUO0efku9twb+riS
/GyiLrCYKEyDgCr2Mi95aC1WP6XCTo3kl8IyK0r2a6ETc7lw2irfjFP52gdOUpX/f9OTam7LKuXQ
rxCDv0Y9K7OAyyZoqDK3KgraKMDfMx4Eyn+/mjBfbxSvQOTMD2KYt1kLEC/tAaQfsLWq8BnkymmP
l4JBO3t8p6deiakZawtwdCK8SBfhIZGx3+VMXgPzE5zMYyBHbPHWC9voe+4N2C/zNL1TFpHC+2fx
KLP9nL6xjX42RKOZ5dPMFEYwBDjtjzZ728AGeOx8JMyAOEeBrrTKnbXLa2nwHPm9nLfqhOE4KzND
t+ukCyo9juXvOo7gSBy0SUHV8Bj4NAfGi30hwWJIRQ4QTqdanLBRylwY5jzEZXG9/mMcr1TVtUim
5hVBNWLi1knB8o8rYL5pMqzrAxpecjMvcdb9oNjdeJCzDvy7TyK3bE/oD7U+GqzM1NbO1fjSQi5X
UplTALmhW4Yw5Kpv6x6RAfVBFeRVHTR18ljlq8hP39qvV+fBrCsWxWRC/GzU7qCCI6FYOIWNu3xa
+qjYaseYGwtw8iuV4JvPFyAupETc3I/6N6jOKPUgttcAgr/ExwlrEcxPE7gg7UzCkAFLMHeIWe9l
t0559CUvt1wg7/jnsmXu/uLflkb+f9gp5sns7rb99MrPUjibciGd6gxBjSuG6DQBT7i9M/RTzwZh
4YE52v7uRyv4lRQ6Ab9V4PJlKeMEIOK91IAAiKMQVxEL5doMhTHdweLTI99kQgJazei4le/nRcBk
DuahEvQyUJ1022CnysPceuj7XfRvpHBtbUwPiFjdB0u1VBEFB4bgrbVfPqzsbTHUHKj0HEXaiu4m
VPzfO382YM8Q+31PcIxxvdZjLED0sKdj5Lb0H96AtPIyi2Tu8kpP+u7bqYEnfODWih6/lnqLsOYx
sZIZOD1SWYDYbHrRoiovGQAu2fm/ut9zljZv0zKZMLT2wo0WcknY0sqRcliNae2W0pYNs5B+taDe
0t80sd/H0XZDXZpPNMCR1Z3txVzSzW9P1ZFC0uFz2kdo+sMp7Ws/1z8sZR3XD/J2VjZFyrAeP+Kn
08igIaYXGHmDSmji2cnYHqpp4PcgTVioOo/4Bw9PeciL9hi/YLiHb+VmoP+9dq4ybG5Ss/t+URnU
rJKHmge1X8UBwJxcaCFwKy2DOtnevBaTvm3XoRBvgvNEqk/2M/X496W5f6ohT0FoLpTSmE3qz1ty
Immj0CF1XmBwr8pq5mA/M1GU63n4mc6N65wt0nSq8/3xFvhiUUk6xxlr08ApDzNx468o4MRxcsbU
wi8C/zpyodEhEqjeXPRKG/el55wSfFT5kG5Bya9BiMxlR5k9ohiQmRunqfNeB4SlXRDZGEUf4+AI
IkTxvPSuKZ0XG2m/ma1GasJ7aT3+86dhVgcJ5oa4pibD7JreVG9eQ69SrqefYgJ2Q8Htq3wX0Rs1
Hg9WJn/NpygGoGqYTG6llX4MVrAmKvjbM6+Ps39a+9u19Lo0TMTYSfOLY2hf0SYTrw5HecbJ286Q
87RjeJ+eF0z8ZJfYBjj1ob2qs+kckkR7TpoUUy/82Hqf7Z3jFPJbQ0kP5GApJNEvXJzAWxB85yL6
SNxkHOT3yUHAQlkXxaJhHfabl0vOehOIhyUG9aVpr2werixyWP0Ecem4pbNNMgJv+zrlv0azyymG
FbfJhm5Hiyst/HHhqZHbP/11795vktIledjlnsRztJjjbPdQeSqrlC8y01jarwCGiwRSIs4ZqMfy
QTCxQ5R5+zg5l+QGINXEQPag/HMDCah26PA/OkBxAUnUUaldXl0u6H6GK85MkdPaKLpokN5/pzac
+bnQyz0U8Djm6Nn5sKqHr8tpIZ+U2ZgKjxSdqvK98p9a15c7T0pQVhDaUKshtSni+wxxNsVcmhh/
ivdf2MV7zPYechJrYVcPhN7hDOFOOMbIM6Gu81JjK148v0r3Ez01GGqe6IxH1AAhh3YGZJOMG6MV
0VPEghdkLIwP+nE7gNPe9nHprR+9E6qyz5vbfvv2Rtd5YtRcMNn0gvye1gOt/86PFHBdX3dMooap
+oUYh7vlig/7vLONMLaR9ICM0DJshce6mfxNuCgy1cH0r+yhWn656p4ffaboAIe89TArZGerA0zd
UoDQEHNsh+n5WYSLr/wcIYKcW0xSxd7RqimmLMts4yrbE3DZUEgIt5z/cgmJwCTqnjR2ydVWKbYH
9EIX9777jLOs93/odj7i1nEuGpdVCu62WiOq3olwF6lnD+7rxcQ/VqtN/buIfYyPbDuf3su1vVJf
qgUfhrxtKhTQKek6woCmb6gKBe9GIFpZrtafQx7a91SZz84NPmQ4ACPrpMwGRy8RginSBqf70bl+
R/9dWfzx5U9F5AVU44yRzwKYs+BKlXgQ7HDyGE4zB7BF9mYIfEree1VDbD811Jj360+gfC5KwVVk
PlyQRgBkp9qYkilgXyJH+voOY/jOnhFgulDXxs4BHXdAtlBGnFtTJaGHkZQExyndj7I3A8M34AgZ
vKRbexGJOhmTGttygLKB0ratUEIE1Z7wVRDxrStKSKfVVKfWAwYGdgp/bslQHkujWSdqCaB1VO0b
nTx1J3ZiVY7zjOfANbB4vI1uF5vDhwfvnSoBDQaoUV1ZVuc7f6zaUDFsqScx6W+p4GINyDwkJeS/
khL2RgzEqaMdVsUn+lFR8qN8DlfSUkHNX9JgP5ujxz+9dMLSpY37Q2pzmKFHVjo8Zdof1Una47XM
gQOBqAuF4i9G3rIkiHkdNcSKCYKwuKGPAn365q2hDc00ykM8qUBf1F/soDs27dASOCDyqw5O06p2
JHJsQQIwWUiRcGuUZzgUhNByjeSG1u4oMzTUhetOJ8Ff2xnjvkLDWmodVgliqBXhl5XrRDP6gj+h
xZ6yAZzipi0+0SFr4rlE/1O40JQPr9RzBurGgpV7HNl87xd/XC92IYJjouUJXFQFNN5zgrcA4pCn
vV30Lpo7jXEtqV0PnGxpSdTfIRbhknQRdcDWaRqsZJ88kyKWdOU7oZeun4E4dtgH8hDhRK3mz+hf
25q4saxCLRMDeR2oIjgKg2wu7Fg8kvufkc5XGUpY8bq5PL0B9MjwhEmION6PKtErrfS5S64JLern
fijJnFQGru55ZfSnakOFJk3hv62T3zfXmTFq3PVhH/aCHb94LM5odYjHthI0SF7uOC3ILnG6NPIC
mabwMwcnd1i2MuxMfIj+L2JAFK7yEl0ZZfdSyNNLO3pgkUMqigo6Pazzz8E84snS5wyJhYixws2o
AvYrYzlC9xvLVa/f9ZcdPpTp+FIK7B4uwhtlmOvf+uUq/zBcP7RxvuUq7wrTUr9OM8jd/OKsC9v4
97q/Rky7bB1zu3ZrP2gVx4+Qj+tWgdbJ/H8S8AF6zcc83T+xk2awV+bggm9lSQcIcw3GyFmPWPfT
c2EEZy5SCTBz3dMFBCEGBMdC0/FKxz00+yqTwUYT4nXztdAyf+BJeG15k88NqTfDH+uo6k+NnAEP
Dmhk7M+WFkMh1LEtmfYaTyO//9QDwzOMR1A0yYbk3tV7dAXNirrTy0BjzbI/uWWuXnJxCuLHPxik
jX86K5Cyr2qQpgl7kDWLupfyEPnteLJ4AIdJ2RvIO7HH7Dj1mLUuHwsqG9H5K7bmEu5emkVtINcA
RSQyafrANRYHhGdeW/RB5P5oA1YJ6hmNzMnd/kqq1HuPtl3vDtCtDdPosdJHHX09T8T7/KlhooqW
NHxNXxIYKmv4hht4icYie9uv1sLWA6CGG7Fl9VkkW0WjlNC4wGxBxMYorjjkaAv9DCBgqbOp0pdC
QZ4PGeedGm1p+rFi+IP/FX1E12hsQZs08bgvMnkX6Wx9sttUuz3VN/XbeuH8xuwjWLuFDu6FJT51
eIjO3QiQKGD7GlvfOcu936zRYeu2NWuNMJjaDnMgZW+T5GoY9kS8eMF2sj/X3jUzWauWFMw6Znyi
dJ5hwmPWH6I9kiFXHBQQUambKM0Sob5bVSP4sfY/lXmEQcCAR9pun2kpXLHysyztV52Cx1EctbP9
N/OYZYNEDxgqVmiNB/CI+4L623hv3zDyuuQsg+KBg9L/SvKjw7h3SwoW4kjPWULtpg862n7A0eiJ
PbROehaMnAxeOCrObrjZzZeYquGpI5HqmdENiPLWpuCJOG9AAxmdCan2GAFLzsO4NOlyPcNXv/KX
tsH5eQriC2ji0ukc9oo0sEE3CYx8ztxmakjARV5sG4dAQXfS4FRN19a8aHfX/NEB7O3e1yd8gN7r
8M+OdnzAt/vbQYJ3W0G99Cd5eYNBKUXaouEXAEmPvn8BQkwRtJF1JnhR3TuBGbu9pg5mMyp7kmrc
exsix1yXqvPYCVJjdzR0BCyQM2AZ3SzkXlB00xfBDsd7ai7iMt+MiaMorZu5T/WFaRecPthDT3Ym
IKI1AJ9EV07kbyaBUn8oPt/r2hrRpCWeN5bnagzY/EmFxzAamoVT0h/Sfvbgr6JaH+d69W/fx77o
KiQbqojdfFtYwSA6xvO8VXWU8Z3TG8k5pNHHx5+EUJC8ma9ESB5XBX4um/I4EFzdG4GbxmOwhYCH
NJ50VGdGMSNxiR2LqFEvoXpiC3hkN84t5Uauzjrccs4OwPv1J1jZCYvcu8eXkFwLJXk8yUzwCXop
B/F1Z3zbJLKFCKFStGQJPqdK7MSWClbnppiu/poaMMchhVZ3qbXZiQff8jViS1R378sCRvflxe/L
GWljeCDNFFjOfbohgektBvyG4MBkMkvPmyZA/K29oPV1zkRYa8zlYkKaJMAg5cfO7gsrT8gpbFQK
QOc5T1+KmjKZq1nr7ZVOWDrvJ6ceACxOCgJBE3+QaTjLcNAgefXdlsOrr0Sf+BZBBwHfEKOMYIzb
HeWMYMmH8Sp4zZSs/yMKk3MGfP2ekY/8PfttD7jJWIkUImPkViMx+UF90ljnd5ldR7soMtsJuNms
rBge1iWwTmSidAOL3H8RxJGmNIvK8IpG1DVY/eUhlHai6bL7z5VjhPzUt6N2SeOAiblVEojsGCLv
boPCmeAmGky1XZHgbMN0ZsjpN4ptvX6B2wX5ZrHgt+C1a98tqoT5x0UeraNq+6TrWfZex90bTLne
FTxG96Clm+ESP/2FdY1z0S9xGzD7AUda7uHx6TtaHQUUsbwWYsgGSY8UDljhoQCJlIPJkletdVup
+Bf5gphMXn1ZUgXhp2iLJVXPpQGxqJ8IToxvRIxb/grKvurnaWR8PaN+U3swqJTHsVxbJGso4my9
mAImRqne4vjtTzNWxFt7rWloV4nKZGqlEAEk8fFT3/mhawJUWdFYWjuiB99fTW60G1mcs8cA4yKa
Th+Yxu52p4IrXvORSGcThdjiSeCwVooZSpSgVWd+FxXfti7kDV3lPN/0HsdxcKkaC6T3pSClB9Da
w13eFJyNZo3k0JGljGP3swefTReyrfsRid4iioXzIHlg+RcVSOxbqmorxxNnHQotwX6bLRQymVL8
V677j3gwfmc41x7iliAaPCw+Z3VRoMQVmiGcfbX5Mem1iVqET6Dd90zQpcSEK2HjuYIn0A4AowGq
tnA3h05MeD+D1KbAM4NcN5KtttLpQnXUsGH6ZJ9grqrKgldmTlKIbh+zN5CW1/7QK6F4gH5fbowo
12sS7TuyV0Cti+Gm91H2dOT9Pdrm+AbdmQdNDFlgRRdAT0Df4FgbTbGV+3BxVxPEM3UYkNdJ9sYj
b1eqp2du/Tehr148utAzfwdFgeZUEpT4rSixktFTaj2ssJcwHkpvl6PitLd74/2+3wxl05Od43Gf
dPcZyqoRMerzlMM8BEt9eHdLSOiHlPNVtWVWZ3kXlbIymwbCWsdarkg3pwiFrco2l7Wf8OmecLFb
dI1lXFn46TaV8Zdpe+JtBvEIfPoQg7v4OGSorKCoJdfKrxyIh4tpZoORRf7e+sI4CI9K/q3ydqFw
IAXN3x1ugae//AUm4d2VUxw0l+B3x3aAI8+uk+riz0PEmyWE76kkoUebdZLjP6cGLgnWSANHcSuD
bL7yqsI8UqhFaZajxGFVcC8rxdJngdYbLvMo2ZWzfl2Pcb/vdW4aV4s/qggPJIeDW6BCEEwEJU6B
yCin9nIY8ZuXaiyYaa6wsDwkcIIezkcwV6GoHjt6PfyOFpT1Z0itcr0lZniZFrXGRco3MNDwK/LW
LTg2GUFQr5rQlyclnZEhRfJeLm/CEePbbZC/Q/ns3eZlasRJGfCYZgYgrbkzf7DlsWSG0cSWX18x
Gj02tE99UaV8GR2XnfUqWVANCb9rqbdZtN/bbhk11UnsRNu6bOiIDu4fllZnUMQ9T/nJmoc/Wy53
KOkiLLzBE1pv3nVEDCg9gUeoDtlradf8aRl+QR5iwQSJqXkdL9vBDm1WjSYJie9Fr9laQYmvWjiJ
pQvMzROTodOyUeqkSS6ndkosPBVxruzTeSPZ8dYo4mdSx/+3E7LNwOfqPcxLJKGx5wEO6eaSGsa2
7qXrzR3q82eNKCzWviIu4tx6t3/egGDDCS6uRx7uhpNeiAFqLIb5TKuUbcDVmZl6fG+6HjNwwCAT
kT79zEcye7bEFxESVwIYfJPhnPV7GW1QjST9lEzxnUJ0v0BwSwq1MdngsMHcM/Y8inrsHvRiON2b
+BszmY3jTPo75Qy9Tb8uR16hWQ6pIE3M5O9tqbABXO+Z1e4NSW38GQLxXJB12Js4GtxomIEbAnrV
SNddnjNP8WrKmUYS3ExNC2CvXuW3Pjrm0hrTiZBKg/S0h0aSIpAOivFVMs02vGHzNxm/Cssyr9TA
/jrhZBdbm3RPaOGMA8aWKzwzpDG5EH40maoEUXGNiim8/3Nd3LIxTuVVn6HytMBpBoFIYBK99IXV
MMbrMqFOw+ulEo13DZJLWzbeJKxLwzpuTGXaFBCDH/+JthBg5cgUpd78hVr/2J9tY2DCueSbG63d
51fSJHBHtLFR0hfHtJII99pbhq2j2Y4DQmIRu+MXXV7xRDkOTBU/HpNT18xWRc839wv0RUBVB0Dk
YR4VK8OeXmdpy7TeggCjkb02+NrlvNeCSXabZHTdbOF/S/YYSy4g6sDi67zOYZCtCwWZJ2NZpSs2
Uw9LsXHs2fT+hqc6OPIxvYDszr5luGgyQxNXLSXxGqBXvpx5QHboyb1319o4eSWFalvpyqsIG25Z
Sa/vvUr69OJrmPn4LfTd/ggpannN2qUZV73VOCfiV2FE45A6rybladtknYZMrRfjL3c1fJWBP3g1
qhGFsT9uGzfUTVWofxmMpc9MmloZZnc4O97HUhACufW+x0XBKH+rANefiCqS0g9pYDfeU9F8a3hP
Gb+qZcN5A9XXtS4B86w9CG/kxbvXK0x+TT35vYknYHZzfwOdkA7OiXiptj3CvPRiVhNH1ZGx2xJg
5qN0Sbb1zT/GgdkVRTM=
`protect end_protected
