XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L���Uq=j% �D:�{Y]�sXM4�$��i������Ű/g���ifO��4�{�R���X#�"*�|~.xb�9-������W;�N�K�B}/ԉ�Q�Wr�m�1�G��NRĘ���zR�O�z>_:������c�U��G����TFl�@\dK�Gn�;掏�O��ux���\�������W@���g���$"�+�q�{x�^��<�3#���~ݞ��S��Do����|��j7��h��g�9�`8S*�\޶@�
1�.ܱn����k\۟6��-����z�Y"�kn9��SPE�X�{�;�%���\�@`׋6��ɳ�	;w�j�}�����튅�=��ږ:S��8��hgH@�����GG�r�b���m(뽩Ě�'��#,��,:~��6�n��#g��Z_h�7����;l���������.i�����9O2v�y��>\����wG��S��1�Cl�"�)�� ��itK�;��m�JE�e_1gQMZß���Ea��-N��bدH�5��,���Ԉ!ChO�m�QJ��̥�S�'�!{�ڼ�f�1�z)m�c~�8n�,�5����bb˥��*Z�q�Q(�ZA*3&�;���x�8?.�#I���+��l�>��,Y@z~&�w ��_��-�n`�"�a[�<�T�[=4�E!1�&uWg��x��ӵ�i���	+ܳ1���U�dM�wV�	rU*�.q{�>s~�a�
�Ak������Z��0_��ie�H���3���޹U�N~7XlxVHYEB     400     190�w�����=SǝD����4�F+�m�}�W����X,ki���MT�Ύ{���!5Mq4�91Ym@
�����7�5�����*�w�zn�r�Gw��QR)��q9�d��:�3����6�h�
;�����$\"����s�^_p�$ܶ��΍�̮_�前h���%�������C�GR��p��	���ũGg߷�`�P��2�Hg�e{fbi�KS(<���� �8dk�qR��h�^ИRS)�S�m��e c�.�aжg��|��F�����a�P�m韌7�b`�ՙw���ۤ��(t�rud�掟�ל'���`x4�EC�ltKM������jBG��I��X�� �Z��vɆ}���UN��3W ����c��6"�>���sXlxVHYEB     400     1f0�'y4w �3يU���w�j<�����R0�m��j
������4�-����Wb+�派\�[��gh�A�K%�;ί����]iV�R��L�8m���H�=���ߒ���QBVD�2���m.ʮYy��k��8"�7�Q�Ǘ�g��}}/;�K=�*=2�V�(��Eǯ̓Fê�� �v����adə�*`��@!���uH�C���}�ay��RK4�>I]Bρ�UE,,������ʬ[+�gy��U>� �r4+h�c��o�Y��-ͅ��HZ���5,��f�ϫ6W�O�SXMޭ�{��*es�G�r�>�~��g���ti����e8xE��@>ʤYa�6��!a$1��tSx~g?T�&��*>��'v� Qi�i1CKd�Bg	�%�:�lD�ED��P��ѣ#����Le������lK���H���l�w���u����&� ���ְ�j�̇�ܧ��#��{� XXlxVHYEB     400     200�ズ'�N���j���ZtaK�H�'�D�n�w��I���� !q ='�5�@~h�n����ˠ��$�ܖ#�u��4�/����l���J�Q��M�`Sf�@��>�����&��nT��Csb87��@bX�<.�&�7Z���$-h�2R�4R�9)�j�}� �٣���p�K"�(J�0�"%?��	۴��|hB�^���لy��W	8��}�x�r�Ǘ� �X�.ѣ FS�h���b]����k���~��Q��Q?�����{�WS#O�1w�=g%O�q��j|���(��6�n$�uN�\R萻t��rĻ�Q���-Th��?��xS>n��{���1\c�f�K�o�L[u��qNI�Z>�"\{�w=n��˛�yj���{�������u�K�ìp~2��/�2 X?/��)Q�foF�V�ؓ7��]i��.vg0��H�����3;h��`�<���&��FK��������*/k+��\����G�XlxVHYEB     197      f0~��zĄ��N/ʽ�~�K���_TN��Zq��_l`��_[_L+�I��A��
��*���Z��t�
�}!l̷�/.�c������YxL}�%�΁�;��M�����e@�,�������_�pu�:���Y2��Bn���r_��fGB9�3KX%��k���+�gNH^���;�t}'mcb��G����D	U
t��V�eT�U����qLx�e�somǬ��O$�u� �vP