`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Wy81LFvy2vm84nkJM4z0CwHBwIqwEsFhCtub8hKQBzo6fSbBxt03SEPyxUzsCnktLUiMvknyclio
o8VfBvPboElkWzWjQ/lbEWNvPpcnrcG5N51OiBBMdKuQQKjMr/goePf0WpSe5bBealmW7cSI/MCM
zbYhs9FngzlEiNR6bacWyIJKKWOXSEZ06qcUgxl3t35SuLqTmgB5UjzU/4U9CFX3RYtHKonOMqj9
ghv/+3wUWxMaqQyKbqUF2DaN4rzmIsA6PXqG5B89mrPMBgza4CwEsAtQV0AnVb12bJK7fAxyD/Qr
2HtIF2okWSenpCoSSSXEMcLx3FgV44GlpfM2Jw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="6+CcWj1BIcNlk/FxZ18A+oaHg3MKADuH6uclydiHbds="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11216)
`protect data_block
YSz4FrZSri0+ORlJxaJZb4//w9mtusU5YImwfq6wzEf2PCf3b0n3vZR+PeeY1AOKKsX5AcEQVncm
zwz6QuurCSpc2F3nsWHA4kUB4vOssg+LbErnAeE/7QXwCuoO3oY2/UBvAHMS2zVFhu+SdsuGjztj
bKOZLV6nHKM72Iv5C+HYH0R7KVeILwjayCW4P2u7c6dNng/niOQZt5A3VKrHsIWk/OHcZx/6VmFa
otklHkqgVHGUG8zoIyDtoeFiTApFALn2ABeY19o3GxCnAGk3D+08AckG+TuJBRGF0fO7yxY0u2Yd
rrHku4kv7ffKlGenPC+F6+4RCxxLODcegpNvsMVoFEN10NkEd4i1rh308mLaBO5g+68mK7/FU0ZV
C+LQko4mQhZhPZ3364flCm1lt5OvgRLWsSxJCVzHgQxq5yLAgrVRSh053kQKjAjgQ5z5MQP5MWhx
tEQMR/Wp0nJVOXVK/ynWVpccgowqTB9rwja9K2A0EyAuw2BecmkeHTEEuSY+/6dZHolZkaP1v0Aq
l+5d6JGbafoGN13TMAvsAWMZnPsz6EkL9yIKyjNw5/23aT2AAY5TvbD68MRq2DHDDtDxejqByKkW
248+MFL5RfG1FtiqoHURKsKJhfPdLqEEVp1u42iKJ2B2OnyxKvmL9HG94892ksRjHscmigwPOK4x
qqaXaTF02nLs9In4hRXD+oQENIifvLL/mjzwnXBMIkbU4IC/13Q4Acsx7PZ+aBaqolyZ9Ejn1RbZ
5yPpXp3zXngunj3qjr0KrPF3j7VV/RZ8KWXs2sqHXFRnyKyidfEKTKHMjHpZAVSqvqgjDTRgJ/Se
SsGw6fgqW7dGff/rigynXzdC6stql7+87OFuF9zop9UnrIiIDBjxHQLpmrXr87jo7tii9jsvG6Hg
8Az6/uj73H6MGB2CmIPIi91NoBD+mEth3CFemIgy0d5p95IEVF7SeFa0QIyH46FzCARK/Lr/eM4a
uXimuWF+dpICmi8Uj6Uu1lScr0OYpnxtw0ob1fNKIzw4RCYIzmv0TlhEsf6JHTHwm5Jn0q0YkB5k
HNQI10mHdSWPv2UspTeBvbo5bC7bgVgTCxdJFWS2MtgL2MEN9pJgDd+vxsqhBNrrcSigchRxR/H1
rxqHNCRt00MVgkx5vrYMaPA+M2/e1dp8Q3LWjUVdSGKgdsmdJO1MJ3u0ZQIap0yz4Qv78cyPftt4
tFxTdfDNuftb7UodtoZkZsJtncSEIJsoKTDtFoPQQfeiuc3QFEvzOvMpsFuRc0s9Ni5I728+230D
PR9fTo5CZQRXVY9L3rWcwsdNWSijVQiL4osoxTyBFGfjaOIuAStGswvG+wVM/ASHQ6dhsZ8xa/Do
n/SpVKaVLHxGvQbjPxBC5Yb+Z6/+6WXHTlUqd/neAGbQj9j+tpwfxcsPGn2ypxNfxx+Xi5Tn2F8r
TMeVfWPJK/pQ5tToV6jeMxI6ofRkb5/hDqFcNwgnk5lb/kgYKm70U2LMMYL7IqdTFuLE2mseK5Cs
DQ7OQIN3Nb01xCu/XFSJ82TqQkRKmnOVERbWQlaZSHjyK7/t5uo1eKrPWc3s5Ax/shiQdWfMheDA
/FVeumJIQVklbkfq8g3Jw1b792s6/sxQFY/yQwIkYBdNr8/A22yb3NZWD5EXBCpFsglbCyJ9uY/J
uwiAbnnV2zn9ygUk2lwNNZiXWiVfv3IVRxcc0+1oSVIdeWUjJC0UrOZS0DCjvziTg0UqtF7kzE+l
XGs9lvC4G63A9sau5GhZwQ6snA5dW36rmdoJlUfqnL2LCSAvY3uQmhxpqouAcNVpOiDdYoy4F1do
2M3VmERetOVoN4Nc+2l/LzVw2FnQaubiAxcM7gSK+1sxpyuiBzrCjtSK53E4sKkF1EECTHqrVSRl
CiFjQjgZxhWzQuG9FnQjX917w060meIlZJE8eR1fJ4qZiVwWrg57b4n43ycLiu7nrhquK8l991M/
aJyGQUGvrASKkRplkbVYDSSmEBPHGF4lAIlo3nYUJiBo9xGpnHGe9Ih21UIMgUTbdyuZjyD0Mj+/
WIFLPMkXFefTO/wtAARyBmwYZQ4qJ0By6WNxvd6tRNF1ytpWE1hkjPfj4QJQF/WCVzmK9KU1Bk2+
a4tTUhGvdkv+QOaMbB/BWLx0k9Rm86xhn61xhDwOrhBxiZMmKdyhcrwM0vTwSFi8oPVKgsWLQzFZ
m+o39CH8N63SK6RN+hlcjyk5F4IQRK1DagldFqeDndiyXsHMuhWJD/ciq1N8gxoYcdLQEXtvL5oS
3lQDw3U7DYF4GfOaE2kNJBUGAldkX1flLQzF/y1S6ULlRVhCi8cDp6MxNMOYjMMqMpljBjYG5ocV
kIZwpyF/kJ+LlW/r+vrFclwjGk47CzXHbkinZG7A0HM27Fi6PcKj45DiF0pF0msfWEdB3XtZpYVE
4RTbMbEsGo0PM9KDGlVqqmQ2mCIO1CUDTy8Yu6NZYMN+CQqz24CBQw++iJmpHiPq1X16Q+PeeCyR
Rqev/+cVbnHR4xH9tWmGr0G7td3K+xQYIkDDyAUkUd0RTClatn5JBObgIIGGP8sN0YpgeEuviqtG
s2qO5Xup0AUJMpmXHEYvugCzUtdERJ2T4kXKEdFSwDSpSl4HXEOzE2cG9mAImDl+vAicOobd+xaX
UKMJN4+hmQ90jPL2tdere/Mnegs6vrdM0TcTGz8c8ufCYpJOzta0uC6Fk1MKtvd3x751yzHCmRt4
qABmw1m7/N2TWfThR/oDG7R3sW/Kw0tAmTq9n1pPOXQN29edsVuQYF29WG3bl0hjHGbEjo1yEJVJ
eYSCCIoz1mIayPS19FK8fVHwXoXndb/c/9CGztASQVqbaJWs2DRdiNWFpkcD5bnrWx8S50bf88cx
L8IlJidW8m7JFcLEAc+IfYPp/iDqfurz6tzx2YQPirMTNmZuLCvZOQmNLyOC01p3KVTbIyU8WxFq
+cpuJ478Z/3Gc7kWlU0fq6Va+drfSLEafLv431drDF35//FC8uPR5a3EVEgjoVzCteBBtylGITCu
JOtTsTJCDlA3X5C8kdQ8Hh1h8Nx/K1m8ehGIRn0jW6uzw6Kt8ebhSX8DCLO0kUTo0Itir2T9Xu14
0O8mxYP6UZoGYzTuG7mB/UpB7/CAIFbZN6KhYzr+FVy4hOOrVJvrFxCUbfZ1sCsz8PdfRSQ1045H
IKdPXU0zk9YRjwgjkdMEqgxDQcBcKHOMCG2MmD+vUNhneCA/S9UB4+g3alwkeeLOQkF7Ec6fg+jo
ELBZPVUIhuCBBT2b5mVdir++UV7OhC1axGPvIlc3CvrM1mfp+vJtcd7mk7l7dGONEDXZMbOUynUE
yb2zAF83Uim79pLZHI9SDwTJDCvrDmchtXUXY9x1fVYZ4OyRRm/SBzfg+1J0cZxs+yugep6DGHjo
awome8j/UXoMFcG2nIJnCYQAT9fN7EBik05NcktysGsQaeGNpWzc691rvj3Nt/oWJ1UI7Bnb3Q05
IaFqkq9gdK7OUKO1lDGdiQNas4LiuKpujf4FqoywLOLwEgJLlhvmUdB30I2YvT0oIuFelU31Hgho
gbi6HV4EkwYV5+zMFxwTIh7dgPTsnonYaR3ImJg8WOVhCRK7aJVpOclpTp71ikbQUO9Gh8IFEeT5
8QmzxTLw5EQC+hIPp6QLmyFJ6zFEwn3ss+5o/v0825tacia8aRblemPXMTG8rmn+wHcrIQG4Yu8q
dNtTsunYqU02fxu2qQ3bltRkzN0VjXuCe/QVLt/5xq7e2BmF8lYehmUyNMCGcuvYfLht44HW3Q5O
8Uts02K5M5QXm+z04EqzlQefhey7UqXZhRu+jsxPTphcQE98awcDHu1o2WlJciy7iYIcsnoHBv9i
36A6tzUPBNnSoYggQz6/hE67hkeWtCny853IdnJqzIJnCj7y2ICKI0QQ5KOQ3vv3g+6JqbyhyhpX
rHc6FOYc54LpeVvHr7e1TOK6o97EgUWMzIlXkQpv5jL12b4cJpNYYI0y9Sr8idYSr01UW+oeH5CR
LPq5rINAcpj9XGulN69wzOzYGfvmshhWr2sHFdn8Z0GHkNHjIix3nz9o98jSepPNB6POCfrvsYps
UZ5djmDtduu5gC6TKkx4pY7F3N7hnLe1YeQZX9+5WePfXqGo96IDh1lCYjLLZnJQd1H4S+x0lErV
Tt6eW6rmrnjAFypKJ1DuX+MXK0+2R3MnqJ6Hfmso+u+T4RbfZiMtAAMOV73R+hGU9A9TDNCzkHYU
ZTQPipEZ2Oy4DqBXN1ZPRgZ3wt7Mezq5T4nwp1YMxzvpLwD6x2ZjvbvW7h8iEcjZLtuPtO369ISi
MZ0KolQ0C6LIwEjsjY0bemXzCKvAISXcswJOWqjEYsS3oufZWKwe7MJSGDZQTIVFTUiB8Tlq4QhT
6InB2JqjNTJ/1xpZjgu0MdpxLvUYC915XggBecJMUO89hxTViQXxISqBnniZxXBhfU4MY/VC2LaW
FqC+2xZ6P7pBkChEgRwv3uwwhW3c1UsxY6DPdWBsy0D7T8Rh/mx1j53IZMcxvdShZ3E+sdUzKaud
vRktxZRpI5Q76UKCkJh3Iw0p6QGOmUxgr4WByr//dNWTmXht9wYasJvf2xBqZbdXMWigZ+AfHd0b
yjP9/DT73f+BKJLprW7j8IQVp+PXj/f1aGLtIa6g2UGDGNUeQmMCUiKlP2WMIY+CXQ3+MNFJ0qxJ
pnIzY+eXrM7HSMyMTxFq0tlo4BZLjap6zEIJkMFXear1RrYggq9VdHpJOPe8uio4K/vGLa4b4miV
noNNGto1hfYWg4q0QCEhzqdgVQvj1Yl6N3HOpZLr167xbWs9ajimWHBwPZFA0ElbGKOWo5x9BUSF
gw8e87Ybj7kmCFHw3faJ0ztDgyu8QFvEDHecLkQaXdXqfuZPVkVPCKp2qguL3LGJ0WWPNwSb9Cl8
UBNilThHwVb2PnA7BloSlt/+XnkM8BIB9Tcj0OyByfUxwzIDeWOJ6w7JuwloXsqFqbj8FrxZj0D/
ovAuH6pl5DWjHl77ai156gGLOzfQR/XGlyn1CqyHZBOHXP2ZrQPmrXKD7Szpm2Rsozhnh6yfhCK3
3S5PbaiBb3pPyPfXSb2wD5XpM2oD1UwpW2PDU6rhC7pNt16sw/Qb1F8CPEyflzA0LiZ6csKXIPii
VnaZXmzEjr3Gxvbv6+mcNNZI6zicM5ePl6+S5COrilQozJ79qctaANkOFa+u7DzPAWDY4TqJ+ll1
d0XApubNAaj3I/Vjkh0DZyirO7Gte2jNFJHZvIKqq+9OuJoam54EaVj4fEUaCBTacyEWNhRH3GA9
3ZASiD7D+EYTe2Kx8KwbU5GJqhDJTyC/Yt/lZGBOvp1RquGQWL7vgCa+W42QN86eeVM7eJqeaoSZ
M+pddU8+SH4Iz4Ya6quD13r7dgOAdgNXV5me1ViCNUY8iA6IrmbxynkbhNK2us4dMFD3eumKrzTV
ddTzF8kSWXM+rCTrmHaZFknNX9N5pkiRMqMLZreF2cKhUxc6uCDB9uz5UqLlvufSjA+4LBClRpZD
DSD061Yiq9tb9fbCEfiu3Yi1F7RxyG2SPwIummhufH9Y5IqxMxdA73crOO92CstKndt0zJGF3hmX
icnBL+sBxU3RohK37rB9RWvO7Y/FhfYLg/7sl3Pvv3R32lx7bZqjaS4uTe1fWLlwHCqm8MznN6iJ
hE8wMfQysZQ8gJbOYstPbtjLSx9YEHe9uSaOhKJVRby550F3gLj0iDmkIIk1Qlr+LX5XmOpci7Pm
f0GTVqRtrSgj1Ny1vprNCjSo5D6BayERsC14aVH+rhbrO7a7G37MvO/vwGTwNL377VYjc7a+6Ecw
xJFIzyfEo3OsW97S65WQ90+V6f2nsT+AhVf+neLl14O5vsY0F2aKIf9YxPRvVCDAw2n0vwTh7Kms
90X7qbgYTzjYXtLWC3ZnkAT+kuooW9uavWiQb8vKwgXINd/l+/PWEycJdv1zz4vJc+iEkrFdJSm6
HOOJBTWYKbC+eJKbcxItbII9515nW6oBEiHrK8r+xYAENgN3DX5P0+qFE0hGT/mJMUK05VJlAWE2
XOXtQx1LzDOTo8n0KUMYbo/LlWOsfu2/rIBfWBnr2MebCYIBhqS9pCzZCs0nctdwyUhEd9MYAxuu
bq1MjB440PcxslSkbpFAucwCMBTfWuzFL3rL5G4XUTXm3S8XkSadbT3JqYnxsHAJ3hih9Z3826jk
bD4TBxY38J0dxNC57Pc4ZgkeYMy3xU69EurJsVFxXght9O9H0+BAz6YCiOQksDlutBBvxBzcr5AW
tfZvIVIIX9uH4+6Z5THoAkmuZJ9ZS+jpKOhbfFDkysBXnlyUsoPhkWEup1xmeZMQOaY4MchSqZ2w
OimUnyk7x0OHVGSRUYUiFXf0Una1if2HEga9BuIbeQECfQripCpZO0G4+plVu70vqdwl0fCMO2FS
2P6Bkn5XePI3GimCo/sUQ+4zjylaKKe/EN1JhEf7QFp4p3Q67kAFa9Z6Iid2Fu7D70XBfGynbVF2
9E+GeF3oyQsnPEFL8OKxSqxxPq9jFSobPqx1ekBykTMJtwOvxOVTg9mUZTYidNt6jsZcXtROGv/C
VZkJrflxkLH95WmWeV+dSEIUPBncw9CcNwpWG2bVCVcPoZNG8Uy24ALal4o6fOe3xg5pWCvSpRMr
HAYRuZutBH5z9Dr/v1OnQYXpVD/LntPgAZ3f9tDdsZLnCYipaPmsM/R8s30Bt5fKARgVDTJDRFdz
5RTp+4Gil9WPsKkXWNJ9W3jqeXCLnfPndekKl2d0T6ycIJBXwXOZ2w7RINKEioBnXz0TZC8KVUuH
iUUrbGv4NuohooHAeLx5wxe2VcXWoapUcQV0TR2OC04olyQZKuKmkNi1OAPEWhzK44w643AW4PDl
pvhPn8sgiLlT5JdwvsyqT5UEykZj2tRFCMFgZYgliMJAflTI5Wl9yDKgvkdfKanyEGtsJefrC15R
Mkso5rUaVn0pYdCvsLoXvqhenmN261CgPEIFZelnVu8KmoDe37KvvTWyaaulPbEAWij8cQacRH83
gC0o401ucEJztIVL44n4TC+hWu7u7nKbaYJvRYeqyDrcKXkC1nFq0NOyf82yOhBcLyTpLC15GZjx
l6vJ0408oNi8f+jQofN8QKDDdSi+8uKZBRJZEehrbEvy6rFG2mFMFkataAEmRE5KlQS8MBXDCMja
KO16u5aKuwySZHPc4Nx3ZL5vWPzz2hP7C//PNMP4KT2ryx/ShydWKnXHVpda6KhUNHBhb4CTCUZE
RSYjJIAKRfwC7eFGhJoHqhjSNLGERC0zK1QyzM1b84BAsrZmmMzIOB65MMLJh7gdI8U1QjUhINQ2
9vEmCrr0OS2gzTjtOH3KzJkNvCUgImIaJISWReG4Rd+VEMUVmYc//BwLv+9xK9m6hkGY0k8tRp/f
2hwXZAIW34HvyipyL0rx/dOvDjk2njhcYkBo330bqEH7Odum4AQ5cKJEK5nD6+1KsIZK/tEQYFfL
C4EoB4mRwhYAi3GptwvHKsNajTAncojwqsn/txPbs4ZDt3+b39o3IAouTna80uWzqHWaC3porbR0
TLr8YnvsViYQ4dSMW2AtzdSbf9QI30+Cm8e9GJgkgr/3oupgUELGhGAggkz6n9595sKSnrmyTv1i
gJprirXHSEHDf6OubshTwE8tTW3qWKHfOUxRzd3/lgsgoqSodVTAl54qJQX247KSBd531/7+PpjX
w+XfsROT8HMlOLBp8MmYCuWH0r1vqR7FzIa2ne0ZHoDIzW0s7DDbyqeLhOZp+QDg2qwf7PUCTwmE
miyHwVblLBv9wCHFzlb2JcX38jtgjx7gccT342ujEaLEoePTZNHlzthGG1WUskGqYiUi63peNamW
D7a3gk3Ei3HquLUCgc8GayBI//vRTPUTaMxePboAEaVYjNAxBQbRObkvbUP3hNH7rN7kcClnscNL
nwMJvVhn0Kb8fH8ROeIuLyXmKSHtkGgXiH4K1yCu/Vew8PZbvxa4d8AuulJQW4nZPHmfDb1WwFKZ
ugX2wR5ormIPaMXO4TPCOHle6qyeilImebnk6rHvJEusAeii27hknBeJ78KAGUc3bV7ZNNB6k1mc
I9DsONTHbWfy6lIWMs0nfUpr9ElgYlCBe55BavNES3lsk1KD9+7NwKxbZ8HTogwFOYMs1EROUv5R
qDahir8bWbha3W2/c8HEtjhrfXX6L9Wz8zuQufbCyjg4Z10icso1RQgwzLK1tptydf6iCIbpHfze
n9spf3QfqQIxddZ9LoOgeYmP/bSRQGCUMjaXXp/zA49klHsEwaAxxsELR9l7mTwW/a9Wd5TDD/Hu
yUr8ifSqngpSdRxtK65D3NyKnxc4/x3hzvIwXiqYDQpVyqWXNh67DkBr3dOtguAT54w+No6/rt2L
HZpERCrrlzjO65qlgWkIwLcvlvNKUv0CWkdbr6ZztX6eYyfvIbDxBlCRNplLqHLXCpLHYUiy6eN9
8GF+OlbRVF+92x3WHWUoIVl7PWvGhF7DwORs68GswOvHMFRlwvEJqbvKbwciR9Ac7DM5DDJan0iZ
PYy7Eh5YJnEt98nJDXLneOdd3Y0VpeYRinpaVqZ93ULwFaouh/ILitARJqotidKTL4gZm0SewhyK
29U1bG3bDCDw15QBprf+Kw66EDEUeYjh0YCq5fFlkKbV/7e+e9l8QURcXShqFOUj9nbCirRa1sE6
vqCQnDmy2iH7i3yeOfzqR90+tCiwmrpU0o8wyzKweT0J5iTDJ9Iz5d/nFZHf1d6NebWcMje6HUHd
94Fnyda8aDl5jBAdKAoSYxE3HCbUDRHEY1uRof1JERi3aXqHPis+BRmeQDphqdD4Jsqh1gC0koiQ
T89ZltYIiyAvatPdT2/vXXGFdRYF2DC2idPkb8LXcpAgnudACD4t2qJZqgqSiPkWwAIoAvlZh+8l
BsXlYYpVZeOsZ7jwdD0Zxwu31aAoAc20qnimzFOM9ZDofJ/8GsKN6MQ4atdU9LNyapEpHSR8M8kZ
0WQfwjWtT0jErQ9750eBDBVSnbgincMWliFiHvRJVfg+SmGOkc0znM5uB67coQxy0LOJuZISbCkx
W8nE/sZwsG4krFb9rNJZUq8/9yTbnwkMyGacYx7C4Qdm8DVgDde82FPrN5ZHhWAOALHSkm7kMo3d
jAMiRdZ7MvDnvPMv6znsoe8UQek6uIpcYU6Qmgo4jhXtrhl96DYCM1IYdt4QI2dwyxp7UugkgsIf
yMP4A2VIa/gzbwzdp4vscozrYQYaYOU5uN1UOtFfxlvkTj/S4Oq16N1pWedO3elxq5ACKi31PWtH
cgzNc8CTBzaiPEpeHdlhuEOrl+bEPFbKzFYNarcQj9fxLCx6PUNzDC/GJsTKtgufgtG3q/PbHo0V
v3vUBgsiJYuNd04RH6yDtvmkX8SR1hQomFCpsgj87NfRbEe9921DcOtGKN7MMtg286UoKUiCPt76
pfiwwKe/h12PwN2G1w00FEG0N4eho2NfM3ewmFBzIuiWdSSkjKylohfYOoUcZDC2dOhMC3A0eE3t
/RVO011GiEAAEo84awSTwxyxkdeM9aZyPcZLR789h2SI49W5BwjKVXKvaudWCkhT2UWUy+fGUQKV
kKDkepJ8qd7mU+zMVKfaxtZskslQmCvIqhhTuEwRIHmrBGdBO38bS2JvoaNAtNVu5qdm4s6zt4np
78Gko0Q1vJYJTFfKHDPPBdOu7ICFaoi/X4cyQdz/YMEHgP6FP+i1fh1GYAEHCaJ67xnz63nIWvee
PmUrfYOASoweSi873Gg+JF4+EGcuMP0AWTj2vE48kLUN2jJHP0IXzPd7dl7505mvLWqHekwdyRr1
PNqX/1gFOyStZk0QXYLTZp8srTChWZ1GUwO1ZeqsQtChb2GJ0r9D5t2vkk11s0TA26nGumj2ri+o
hmZMZsg5an/w8ryDce04sWrc70jAZkBM2iwi4ER0NPJcyk2TVdOlE7bc5WJGrVvqb+/0K2VNNWhV
xFRyr84tHNvPQ/JP/M0sU8mvAugYL6XCQw0VO6vLKWjA/40DTTqbA/XbpeI63vCYTBVfi6p6S7q5
FDDkGZCUaGxnXmBovc8O0+rtXBaeSUhRJcnL+O+YwVbigAP0HVehd8kaiJNPB3uAHcgnseWcKJz6
Cuy390CkVeV3SCfNxLibEcL5nGsixJjuwnRvDw+/yJuYsx+1f2Fjb6R2pt08KQaZGH+WINUP+7sA
wy+OVjc/4lE5LgVgMnHOdszG0VMZJSMDUwYrUJZ7IfRWyrQL+AMu22lewcVO2kp4lYZTKHzlhz+S
9O2EA5NeYh5FN/83Fmhk/XisdjCgd/CfGI5xT3ascFrCq0Aw/yl4Np7MgrU4GlDfcsIa1t63ORLu
/Y6n04+tqvjyAChj806q6vda74aq5lLxizGKSZCJtmiEIgHIC6vXZfDhnc7vTf/FY8kdwi3N1myI
/AgosTj1ADztCYPld7+B7yENvhJknZU41GGpj6WXsnabf2I920d4P7c3PE8EKwT3nqG2LwXezEek
Vj53UA/4pgfdtAf+8pjGD3eww9PjNeJ1VqKChUB3lIoTN2Ns3fBTbwA57B49DmOox28M1AH+F997
VGOoN8UlwEasjrGqI5ciiq3nyu1z4zgfsizvMB3+qUCDDMzvuxi3boiGzE45VcwjE9iV3ebFPptf
aPeWzexDzIwEoG+fNV7smWilMcQbGR7QfRdPH6YKspxs170WzsyXfXHHMZIJN+5LI+zdn5JxLOcF
EQsyZvKO3rixGahxTqtOnpF8GQ4ROxX4v22zOHUkyJufw24eyrSjXLlfMZ6yqW4DVPQlbQRxelQP
yN7TZAl9sOmdLfcoZyh1T/aRzT5VVhdjiiku3EfeCmNkjc1u5S2AspVjZsU1rwLtm68ThfyWv1xW
m/w27gZ/yeOEm97ikHIgbjhsKhm1Yx45d+zRh1f/y5Dtu2y+3v78drpjJQO7lsr0wQUKVYzwfv1e
dzIxYiD9Dgtxhwi719XPrLAVkJjI2ZBUbgq5t441GIWhbAxNONPvdFI36iLm2xvklbiDD1SXi3Zt
Num1FvXjH+8MRJAdbUdyC/z96xcO2ySIs5M7Xz4R+W76xDmKXl8GNQKlBkxVVRlEBArIubN8t0Bg
WDwYmzMz8kURHlI/u4rHWTNsnuyd/cbGaPVTnlVmYMSnMGN9QigGxKt6Wh8bm/RbIdIsu/TYMHlO
Qybg2kigtRogFd3UqG/0nRUWEn0k53bsye9DiHyyhK37dKeeGjZbZc4+wiQfAYG2grbhfGeVP0Tr
UTbZpIS6WtrK0alYYf6nmLhBdBoN+gXrTjkKj7c1Od9w6osLvsZb0joJ9cTETF+XZR/iboUMiRXU
H/qC3CRDvoXbh/zScLbzAB6p98TDes+4Wlz9GxERkKZXySPAj2/84YMrSQDgyZ8evxfQmOdpY4hZ
DHOj1hMKkjoYcR5xKjk3PHbojyxprb9Fm1ggTgxGQTxsXgCsLZ5DxXu8LlrVONqi/CYo7oWFMxBJ
l/5b7QTTXpek6eEVQN+4UuD5J//28/qVZhdjuA2YdCRCVTcYRsnBtU3PKE3F8PY8yQfh9xKViYTP
2+OE9ptdworUk2QVQNPTOqC91i16f/srf21krWetzI4sy7f3Uhq3FVDc08jNr6TX5L4um62pxoQJ
rNwBI11bFhweS1BsKh8QNordp0nHOd7oofgyHtT7IEHuD/tJFTllcZJh8N901suDg5O4Ha8/1LSc
7bDqWHBoBRwMrtWsNhHjwdyG9257WVCRQTFqpfN8N7zaCAMl3kN5rzgV2SaxmYMepGX4S37JJ3w4
X1NRVFEhFUKkRt+Ng2S6/ebxQO+R8QUjkF18IUk8wPTjr+VL0mbVucaRD996Lt7jOpu8017O4PRI
y79IeLBfRZq09dSDqVpYs4bU8Hcuioz3VH9iYtCe2mB+15zje0ogLVmUtfoCZHjRpCODqRysmV8L
HO/KbE9pLzoJKsupH6NTFkb/vT4V4zpnpX3aRGf9OzRzWE4rCeI0cxevPhyuEhvHS10eIwd532er
tU9gw0ZuZMjEADfbIKFbJEkB1Grh3EOfZJFVb76/625ZapP71sqEHMmukYNWxcbxufoCDEvJZuLJ
xHsFOAOxPX+ovMPBwHJ5YazS3EnElh3NG/2wNSLu2fCVfQDJdMzik+o4DM7gc6lmm21yiylsFH+X
wY2wGh1IpEihxgS1VhRqvjW2PwlJQUQD5SIlH2leh8SdcfwqZZ8+BZh27PJNrWUy6HFBzUf9iVQR
ElWgpN4BbMwKsbl84WXJqwuj3xOG94snIIuRNYIqieKAg9MG3rKC5k0bsOMjI/TcElBZt/nVodqE
adp6LVaNERAEoCpdPkGDMqLDMplpB5VOuoGwss5cFCpPpljzyg0YddZhP6a4cMceOB3eZqCPb6Uc
VrQKwJYtjpEcd47O1RK1h1VtZlscYsfXo/8jODtEes+xlqiDja9ejpKh09wevD4CK1PUVLH1/0fp
T7dmKx6NLcOkeMedQx12vg54AFVlZHkj1IVAMUFR+6Jl9+u9jwm1uIpglDBJiw5CYlvGBCcQXGcH
fTngBbMMxAvGUbnJ4vTD069AW79WnE1Mi8FY7Yi9gtEQRmvMCRJeGLYasunRaB8SkcQiryV4ACII
H7KXztlv3/tRQnveguqR4uLaFxNxbXsZWX6/ERgoBH23C+SSfXva3OiJ39b69l1VmZ3IrqqF9OLl
0OAlkn3x0DU7cwDXlgDlt0gQ4dApsDHnf6xDeKx8PAZCy27SoJrmjElo21bz+PZPgY5TNfIjpem0
M2UttJPOAAbFMiDGFlt3q5SV+50t+RaG/l2qtcm2L8hrB2HvH3gQ9xQhHwH0XMesfVKSgdACP7oy
hAB96YU6JOsUDRDrdAVJhK/tkk8Bht8a8XkmPZqBHIkDlJmOe9ZByA5kXFbnHMZkm3PB2PvKFaS6
N+u1BuuoJLyGO1jTHTc/njpCFrzdwOYxnBG7msbYFlIEjcHnI2aCHv3qnCCEvIh7nqfcJiJJju82
VYMz2p7SyfwkOcQwIdkNaeFYi7CFGYbEn+1eQfUC7UiAHVd8KgA3LrJleOxFcyHDTxPlaZmW/21U
1Xdqo6r9c+MRDGwtRByOC0Sksm2GMco/zZAQVPm20ds25Z46X2RmRGIvpJZNj1MetGwGutWDDqpW
QlKRUM0I7U27QFs/iL9+nUBtlY/nQZ4+8f7Uc5jYLGAkhQHg30HCiWhnWeNBLM0AJ1svoLGNEyoH
fLpa38PSJYtI0Ib+ig+blM37M9bltC8BHZKJ9dpUI9teejTWUCsYSgK3bfUym8cl93c/ihUP1p/J
Fj3hdbzWmZEID/rsWp3aNqnaFmmkY3+qfCj7fGOapsu+OUgSilUpAaho0+XmJos5VDvTVPwDCu9j
7W947W39Q32mtQVDvLJiS0J/GL8eKCECfS0PwtMlIM6MZPRKcX/KXI8mqZ0Knza9nUFXyINaPSrd
cqyd7Wx0QLfZPvwDaG6VCqOqHtFbWf9BVvy9NoPOpKKSt7ZX3+raSHvZ8nQPhL2M5ofnhyFAn1ew
WoNQesawKD1emkKESYAss2wf/ZzAOzHu+KRrwyu9H0208tA8Ilft6A922BvvWq0uRUX74StPg2+E
OwUO4gVSTehl+FGMLvjxYeDY6XDST6+vWS2HvTTjFoHIW3757gThaHsDZHjuNZdbOoZ94LP/Il5U
5W7763oA+FwgadUjbQgFFyPrMIsYblM7ff9E888qgyAmWIijUwylfJPbRMuJo4w/wdPlaBXFObNU
2XwpVKDfCNCQ6yD8tstwpipKlTsxlkftbr26FwcIhEZ2/5MsjDkqfQKT8QO6L8xcE5uW4WnB+nLi
XgfsDOX/JrjMGazKFBkW4Npw8owS31pIeQPM/3+z8tBLCY0TSBG3gcXFr2TlQuT9Ygn/IeEL1Joa
DZx/moXLAxZt4IObTL8BHruc+JmkvQ7qK57iZmOXVpyf+laRIZpP4vIB8OQ3iA1X7Z+ELOPMkNrP
GUqulgvkti4P/l1KgYFuw42ZoJAmZ5lxyA5g+ax/bUGCTvPdYQ/wpnIBz/Ehb/bTtNVlig3kdq3b
WYvtKAN6/ADaW5iNfV5VTK07HjFIbwyPvL5BQRkqi4oEPbtkmGWwAjRVlCz0qDVrewSProoYA8Id
YjylwViFccNh4EXC18+ylrubarVVpoNp7rHCyjbKWDfu6ihROguVvYn/PcEHYM7rJBTVgpgHN3Iq
ElOCBtwcpkBldQ0R+EvS5mJL21I4I10GlFwK2ahHkHSnFdokVWXhHfMb7ShzcTKndzz16GCZQuZq
JpuVfT2EqRnDvbP+IwUD929EcWMIClkjYMkEE/S1u4uDrT/K5JadPp92n4t6hHrLmGscRxMvI4Rg
dj8OzPe4iuGKSgW83JC081QxcmjPOfPAqsqR/3l4KHoli4rYSJ9Hiq5V5ywnXxfVBlHjn++pulFc
RoYmrG2DtQp6NUVdpuhLhVkCWguvuUW6GIj8jKgaLZTSqDctWhD6qjxix61wQanhsa5VGLdkjqZd
kHebS20z0yPpwi4NYfgjZe7OhXr3nVVSJAZ77tF+Ob5knea5mHqr5R/nTXoyo4OA6jn3oKUKQKtH
ss2vLB3/P9UNlBluyoSyLpytQjhLzdFjRzN0/2IQyuXw/0NFieRdtUyt85QjlAjebk4emsY0k9WN
gKSF6XZEeXKMD4B+x8E/dHFHw0FWhl4elbtrNYIaM1R6z7psjC2mIcSbu+ItyMom+kWWYwMBQQtH
mj+i0cQKLBAryPWuai8krn1WN4osebuglYYlnwIa8G7TygKwVBL0x3GW4mqHp7ROnglIpic9AhKG
MQyTzf3Ma0AyTdmQgIHRRAB+Wr+Aw5nKdQAg2qMAXDTpkLfng34Rc+4uRhI=
`protect end_protected
