XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y[]��a��W�lㅾ��ok��GoF�O�o���[f�2mU�I<��op�A)�V:�|���p�u]�n�E��\��O���Q��;A�1�,����P��ǥ���h�g�^��a��z �>]�ti����ֆ$gw�f�gXD}�����!��>H���g�>�"���8��r9<K���7�����(sˣ/ٌ\�3�Z}�:���� &pR��^�Ʈ��|6�A��x*�1�ĸ�V,~�|+J7u6��w�z��<½��K���$���Y��pD�$]���o�1����S��/���G����[����۹�j�<B9pk`�#h`H������ݣ*D�X�¦N̴C����,���]!�+���|˅�������7�>�1ݥ���n�sČ]߿�-��T�6/X~�Y�J���Z�6�XmK�cgI�V­r�4h)�姑�[���W���#VP�!��Η.�q��d�N��$D��a?�Zҍ��+���ڀ��̭��(1�*��֐���^l�S'�i�Q��@2-����AxW(�)с�4=37j��b"a�h�F��'&zѵ�z���OkqX�
�(�Oe	���T�m �.5�{�re����y�W��W�6�4���ɼ�>'�Gٳ��ғ�d���u���ڿ�Dmt���y󂤃*�K��K�}���|�]�H= �w�,9��bk�A�����/��He:�)�)];�AG�q���-�Twn�7>��07�%��6�.5�}�9U(m�U�XlxVHYEB     400     1e0+L��p�n���g��(�*��n�;*��	���A6�)��i#���N��/�v���1�b��uey�	{@�+�W�a�-���s�+�Ҙrx��n�3�_P����	�>�igl���n� � ����N?�������Ce��gQ���,y!-6�12[��%}�ns�2��ق��8��$sq+G3�޳��Wl#�(5q���(�&�3��~dF�B4���m+
I��~�w<�My�c������?� ���DVO��̆��HHi���2�kr��|9�908�6� s��H8A���������8����R�C��9"��vH3���R �%�0���Nw���?�#��pI ^�f�ǏK�_���K�Ch�2�y`s��V�']��%�2�4;j3���%k�a2%X��*i>�[~�8,��h��B�o����"��*ʖ ���?����ò�����{���*�,��e�R�tsR�)XlxVHYEB     400     130SX|B�B��N�u(��Mߋ�e����]�N1�)"�:x�O�E�v���H�庠�ǚB��屼f@?���M��!�[+!�,���L��d� ��,O��+�*8�Վk���!�l�h`-v@NæC <y�ރ0��&�������P���>�6���%)(&6T
�D��ڊ<�s6]�/N��{� ���Ŏ,�-{{<��_9xD��V�֔�g5ı8��	_u �&Em�f� >�iT�1��5x�&8��·���Eț��K�i ��[P=�G�7��k�X����*�^ʕM����"XlxVHYEB     400      e0�?�6L����fAs��T�<h"��pxVv^�Y)X)�1>bw<A�XBW���8�N}��F���:���u��
�Z&^9c`�����p�S�Q^_��
��LaK-4 ����>M��p<���ɞ�4�XF�'HAaJ�Z�؇�6U�><�m�r�5��:N�8�
������s�[��N
ܖ|����^�<gA �3x����aP�S{`��JN�rЌY�3_]�XlxVHYEB     400      e0������v�LP#0��n=Ocy�@.�9�:�Q��^Oe����H*�q���*_ͭ�BT;)Bk[���8=����2�O���j쀸@x|_1~���އE{��m|�uJ9ڋ�2�|�7Z��v�ɏbd�����>�ny�;��C����#�S9I����v�%f�L��� ��EZB�S���sĦ�oɽ�!�2J�1#�Y��wͣ��S�0UY�H����j��F�XlxVHYEB     400      e0��J)��s��d�W�5����@2fxY���f���N }��i���	�)<�Go��5k���4ʸ��7]9U!�G������qU�"�*�jx�4,6V��I���*��'xl�+d�:��d@��,�Fb}=/�/ߥTdt u��ҹ �D&֘�z%�y.��"��j|I��8<��K�T`�"p!��gv+4�;���,�%��Cn��U�a�k�|5y��XlxVHYEB     400      e0�T/._+}m4�r-�lRc>;<�Y��(n�|S�l�Rwlq��[��y@|�c�|��Yt&Aj;��� .`��N�%=��x�8sx"���(ں�fQ:)�=�N���;(�0�t���,�qp@ĥD����,�$�.�uV����ɶ�W[7Ly���:��2�@�ĖlB����>3�J������T�O3�#岑j���%S���C��s+Uh�	��Iy�&]�XlxVHYEB     400      e0,����_�(���+�Ûh��v��zN~eZ��5q&T��b�V�M��ή'���E��+v��i/�JU��eawiR7�����q�@���PZⷍc����쨌$3�<��.>�g�����VuPQ������Bp����/$�u�N�H��3%z�V�~u�+�e���<+��X�p�g����%*lv�F�77��/#�<6U\�WҢߨ�lT���gXlxVHYEB     400      e09���V�$�@T���y��/�r����gMJR�q���d�&�T�,��Ism� ��;��sA���#�dZ�~H��"��Ո�M�<�	�M�U?X�T�ЊCUe!��������h(�ns��]�PA��WP��LXn���5��}m�H�MƢ)	�+�8�v�`�A��Nۙ�T��d�A�~EhR-o��H��U.�# d���P(��5�X#p^|!�k����XlxVHYEB     400     1a0�g���MB3�	I��B�2�ŋ(��8[���ь���b�{�n��u��RS�j�
�zk��[#\y����_�"�%�����/-�(<Iu�5%�K��t]��U:T�i}�$&d�Q�o�;���dRB�o�x�&���rУ/
/�Э` �i�������^�\��G��ŕ�a<�O�V��Ĵya�r>�&G�&姪'��`���<PeHs_�ƀ��z�4a<��O�zy)�¥��
�ot�L�!�+N��2š����l=��]գAڔz2*1�>�B�k��6E���?��Y0�39G�-�U�=��n���0��a�����Dԡ9�P��N%p�Ȋ(_�C�2��$ϖ�t���O\:��ے���-$daj�,>�Xj7Ծ�>_a	rAצW>��u��g�a=���y4XlxVHYEB     400     110���d��_:�`u)��9M��S0.;�L����4D`�N�$�/�l<�.%�l�*ϖ��=}T����5ˌs���t|�s�#S��H��j
�-�l�qE��v��b搎�a�3����̏�Ǿ N{j��w��._�a�"��y�����e����vy�浓/�R��sᙖq��8�=6o�ڒ�r��K�i���8��X,�`?�b���Z�3�Џ�C�RQ��r�4�.���-�ߐ7�³��_:A�օ�Ӿ���W�:��XlxVHYEB     400     180m.;Lq�F_�x���]�9�����k�;����-�F�������|�J��;>��
�/�0E̹���FَL�=�`��`G�W5mnrqu�	Ť��߄ 8n��Pm�䓷��Ck�I|}5NJ(���r�U�ի�� uO1+������9�r�7����_�:��e���ƴplc�
�w�7#ǵ�>�ڦ����g��t�H4\�H�Eh���XH�EL����Eᐷ&�wK�6�W�(���e�\1In/[¯��?* 8�#�(ވh�վ�spI�����
Ό�L^�E��b9��%����j�M��l_��":}��#+ ^X�8�)�Ԫ���K[s�M��v��C���"�I����>��$W��}9U"�Uȗ7�3XlxVHYEB     400     120����q�Q��sMl`0�~1�J�%���P9�	yCM��J+"a����R,ZU8?S���hq�W��ٹW�@}Uy�.�ͷ�:�}R!�KP�Ӌ�z�咓�6~
�\��֣��~�(H�I 4v�WS7|h����B4��4�T*Z�#su�w�=u���;w����' �����CnI,Sn�FY�f^e��bF�e4�˜ouX�Y����*��MÚ���B�tCYT�dHYt�kn
���&]�^��Y�T��f���zr��-����7d�҅�]��XlxVHYEB     400     130*]�D��N��}��~my*�5νk�y��i�5�N�1���?q��.�����Ɔ�;?� %�KV1J{1z�f	U��4��%�ؒ���ao#�z_�{�@��_�T�/��7B
+�⤈�����a���g�0��S&%p|�v̺��X眘J���i�/�)er@������٘$�tR]���8[w��mt��j�����G�h���"t�d͗DS����r�+G�\��a\�?��nՕ��mb����ԗ��z`�L�ۗrXL�pH����uΜ�<��sB �BN]_"||K��T���f�M�M��6XlxVHYEB     400     120���a�+,h��
�,�h�J}���~x-�鄃�$#'����3�y�,qߏb�,)�j"����ߪ ���b�/�CvD���"�v�����+���J*]��WN�w;��¦� Cm�"g �>�҈�d��`U0���ր�~��dfb7@ v	�0�/�a���D3�#A��qG�����;h�Ʀ����r��P�\�����^�n�h�p$�� ���>L��Hib�v��?��Y	cM2��n�W��)�X���(���b-#�|f)�"��Pl�u�E��> �Gr�G�XlxVHYEB     400     140c��Ǟ�i~�Zp���>[����ۘ� oJ�'ը��F \jފ����?�~���5�_1|�V��GC��LB;L^��▬�,��n������3lb�'�2�v���w����$�-f��[i����Ơ�"e���Y���F'^�bX0��>�H���yk&���`"��I�ȣ`B3�g
���$�Dʷt�T��޶���'��nҴУ���e���(u�V��|����	.����쿡�VNe�v���˷�1/�� ��^iA�G��f�Y�Ϡ�j@������ejc�%���` [g)��I=$�%���u�x�2XlxVHYEB     400     140�7���H3.�Ő�� ���a(�RDB8��J���s�>�`x�$�������_~-�����嶰��
�AN��w����
13<Wc��+���E��p�J��6��&ϯ+AE��v>�(�m� 2I��f&R4�ark(�|��j��`�T�ѽ1��v"��V�3�J��*���TmAc���~�g�F�Au�UjY�ޒu� P��|K�j���;�m"�2�v���C�?�._���ܚ�ܔ�4}�[��r0���t���R�ﮫ�t"����ޏ�uT[���e$~:�Ky�2�K�������Te\-b3U|�� �SD�b�RXlxVHYEB     400     120~�i%�Ƕ�b�>[?�:v�	D�ĆB&l���"��;ߣ�N����g�/4��U�a��-�����Z�6!pL�o�o�=̫j���C<(��
Sb��8jp�~�Q���Z���.`�2�G��W��R*>��<���(_t[��!�uCz3�� O�r���w���4�������<	g*pp?-ӽ�a ~��ڠo6�H�ҿR%W�[�O��/�d��E>�s��cu�G�����'�_&eR����/�,���AV�m�@��y\J~z���e�ӷ �	���_XlxVHYEB     400     140���0s%��O�ma #�${�0C��[��&F����žY���%]F���[��iz!D!:J�?"ɨ4S@Z:P9W3!oH��Aߓ��R�-*�S��R7ޝ6�:�*���	�*XN���a��Vd�$j*T&�,�4���"Y��P���P���<nms��zhq��E�;��apu IF�N�~���D�fQLw�|Ey�:��n� ��A;�m0�t312d[��)�Q�5D}�!W9�vp�Z�,��v����z������
M�ǖ�����ZO��X�8�\�
�2�Ȋ�u+%�g&t�n���1�h�停a��#@�XlxVHYEB     400     120�x��hvNf�G��.v�E=<�L�$�s	-�u�~�gj;'v^*�,��Bt,G����~��������DY�,��z�wE�܍��{�Y?iE�1��5����qt���ӡ�I=&�5��{�U�9��D&1��9�p���}�>!D�1�몍r�blǵ�%��r��d:(SFD���z�yfT�gdJ�nݧ����WaU���eٛj���M���k�fۯ_�*TE��D�Wۛw$ ��'Mw���KNP��x�oa]Xk�-ġ`A��o� Z&��i��Pd���XlxVHYEB     400     130v:��dQ�G�]/K��	d�"����O7����U3��ȥ�g��>�3_�Z�Ω���9V��)\�<���)lI����1�vQ{7��D����9m����¦��>�}��O8�D��� Be��W7���`����W^i\f�Kz��l�N಑G�!�ל~�<�����"ң=F��IW�@� �+�s���1���B�;��so�3�U��j�6Ъu�����4�?�ڨ���g�����3g�Yk$�k��H�.��� cbFh��~_��s;��6�����EĜ�%�+��SQ�T�g��x������{���XlxVHYEB     400     120�8�Z�%?!,d�������%��R��n*DɩUk�����\�B��]y����;��6��[�4H%��u�~����JH���<����E���{�+#�������]v�l�\z��ಷ��H�iWX��8[Ӂ��7I���4����T.���%pR*��h��td,�#�D�F�iŁV�;T�"��H;�u��i��8���4\�!S�7�-<ɢ9FgT6���I������N�u/��f�� G:@���%��~6l�Dl}m����5��0XlxVHYEB     400     140������2wB�`F�k
u_Ql���h$�|Oi��u���6#�^�C��=�PL��WW58���S�����`u�,�����G���J�:]!� ��y{��P��������,<��Q�^�.=$͌��h���#&cf���J)e��\Y\Wm����f��*�.����׉�v���z�yt�ˢ#�Ƥ��˫��Z�ܺeu�A���!�j��a�L!��`M��ye��v��		o6K@� giBa�PoOwH�xw�*�R˽���O^�a�2hϺ��VѠ���'�r7u2��O4�в����B�h���S���Ϟ��XlxVHYEB     400     140�7���H3.�Ő��Ne_W�gE�:�kjP���Lo��wY�MK���R�Y���P<�)��?��\��/��K�S��({��c�$��A�5|�Bgћ�t��#^��RjQ���K�H$8�+8��Z-������K��~|}��)�vǞ�ݞ���9u��nBye�p-�������2�v��#����7�co�w*�K�����P� ����0A%�<{
8r��BBf����O���۞��ø�g��H�y��T������o8���l��o=���54�0�C����{/1��m���*�=�ԈXlxVHYEB     400     120��~�]�E��sL��f��C|�Z҇E	�22������Ξ�hod�(��Ҁp�-\8�sӱ4����z՞kȀ�*9W��X���U�Ε��F�Ca#c��Jf&���C��.d!�����
'۷��b$i۰>���6�elZI�~mbÃJ��Xk��8�o:�݄�`ȫ�򹺾E�s�=�%ބ�2Awn.��ʟ�\��	��3�׸�G��:c*�h0B'���@ʢ�	LRu�?�~��b�E�v�v�;3��.X�����a/țOW	�XlxVHYEB     400     140N��Ӹ9�6�ꊄ'�6�[A��|��;:��'���҉K^��([vxm��{.E�̮��*�u�
'U	�~Y1[����_��OI�H: Vo�u�S�ƨ�|L�6T�v��[��1@�D��	Q@6	N D\ � 2����v��T��j��nЧ~g�<fy�_��h#���MEZn�j�z_��n6{s
M��)��	���7"-�H@G͛˾\��aC7[O��RW�d�PQW^L}Z��Eo� ȿ���������_��<N��(���l��ą����z���B/ɑ�New�3 O�{�;����Ӣ0�#=a!&XlxVHYEB     400     120�x��hvNf�G��.vܲڷqPAad��겖�h�;E�q`Z�*���Z���Eu#��drL���* 3�&Gq�u��h�=G�X��Ԅ�)��<{�d��fO�͞�D��.�?9�BZ~g����4<�1p]�����i�O��a7���F��@�;���E�k�۵7?ء�ц�z��g�q)mx�������
���{�i��Fx��0���2�4N��)��)��N���z{tN$ށGj��2��*�~D�$�nn���}� ع9�<��_XlxVHYEB     400     130$�E�fմN�Zl�pu��VѸ�������=�M+��>f�)���Y�)W�����"u�;��u��H� ��	�_���v�P����.2��%�N�K;@�G���@e�����mH��c�%����%|ǯ�G�/�v�҈���ve
����("	쩹��U_�	i�'!�2:b.����G���#2�G��ɈZ��`e��@,.`��uS}��mLbO(�cqjӐ��v]s���jT�e�R��~�s�w��;i��?kc�#1�)��0q��g�Vn|[�jNS��F�-�q���+�^�i�؈۲hXlxVHYEB     400     130�̶��� fOSl��|U�����߷�W��a*�j�:��n����t�$�J��@�M
�_���1e��k������_?D�Y尌t*h�/I3~�i�����'a�!��{��I���eR6�KV4�v��S��ɤ	���uu�:�s<����8@(��m�`�p��$����`��K
��``<g]IM�V���7���^+(:q,fj��R<�SJ�3<I-����735ϣ �&��Ҟd�!�8�J��vδ���E,��It6��%Qט�����X��ϡ4{�����	,�_��6 9)�XlxVHYEB     400     140��QQfP)PC@HkF��Ȓ���Kf]��U[n��1��m�|Q{aW�y�t2��αu����-�ܧ��a�m�y�ZUżm�B�BV��%eF��N�Fhf�S�6��e�n�����[��׏�{�o���*ph�;�@�S�nR�]�`񈸤�,R��"
f��`�Cn�JU��Q
��:(�d�F�	p9�]���p��?7��X�H���K�/��^�#�l��$�7�<�-L����Qi�Y)�VY�{���8ǥ�� ��5'��D�u�i=�y�G�t�hM��+/0x�i݇J�ҭ*�c������Jo,�?��XlxVHYEB     400     150�7���H3.�Őlw���*�Dl�3�cY��G�͈���Z����㥣��5Xa�l�(���'>�|��5и����񂑸Z訍fu�6���uo�������(>�ȵ���r}a����d�%3�S+ұ�dMJ�Tf&IM!j���
�V�w��0~T�
E�r��S�E�� �%�=#Q����Wl	�4H��Pg�g̀	禮����4�$�~����">ڭfp鹳�(��;�s&��Y��Z�gm���N�͠��拥��'�ͮ��	!�����o��o��H��[�^�rο�5�ZKUa,0��!8� e���A|��4��~�XlxVHYEB     400     120N���ZH^�dB����ÑL{��6,�X�Q�t0�&�.��]K���n�`h�V̥��s2 �#�D������������bѬ;�4��)�2�b4>���U1��	�}X	�4zA�8��z��6���FrTJ~�nl`�#�D��B�x��[h6��d��:N�-=�횕h|0����hi�8sƝ�l�GB[>�F?,�O��8��[�xZת�1���$��A�˞F�sD���t�i�2�gM�"�3�&�>���g��a'�,h�)�{Ot��!�C�g�&�@�SD�XlxVHYEB     400     140���41-H�ܨWPR[X}��w���nm4o7�b�d@ک��6����ZT/< �<��c�Ύ���LU�(YKف0��>Az��ǘ���|�4�D5s��0�,0��)�k(��ړ���>�1dK�� U����OI��՞�n�2��6=� �;�jmjq�A����$�+BhZ%���ׄPt�.���Е�C�A�R���`����Yd#0��(���L�w�9���Bzͦ�Tku���j�;�-vMԿ9�i?�i" `��j�����*�$ ���5�P~��e+�f�Jg�ϳ�*E�����Hc�T��27fXlxVHYEB     400     120��0��J�(h��m�,Q��ɯ��NE�Zcͻ���
ƾ��`.a\����M���K?Й�M�y���I�D[_l�� �-!h��%�"��d���Ř��}��ɵO,����Sgf��Kt` �0�?����1�|��݈{���H��=x���#DBY.
㚟pzgUX����L���n��n��E,�a��C-�*Ĕ�����_GG��K���o�䧬������/Nq���[�E�P�0f���YSw<Yu-��v��nnz%���3{[/t�w���XlxVHYEB     400     130v:��dQ�G�]/K��	_H0R�rY�
�?�(���8��O�k0�p'f�k�ߏr}*D1M;�?��-m��V����A@ɿx��

�I�mv�0�ne�֓�%E�10�tC �V �((��n�^�:������,��%�-�P�|���[� �b�0�T�kf�u�t�U���V�S��2ZFH���r+Q��ȑ�k�4��?X�|�1�d����C�W�!ck��q�7�ɥ�L)|����@0���9��=������w�E�	$i��S��1����y?����d���f�m���J�XlxVHYEB     400     130�̶��� fOSl��|U��1��y�c����!�lo�kg�4J�{[�+OO���?��[P���#� _���@&�˳tIf'��*6���n�f���t�Pw�?�_1����GS���pR+�Xi���f��0�[�����&_�mP�}ͽx�Jr}J5��M��@��?nx�:ج���*�շ��$s��R;�j�P~W#H2	5�����[)�^Ip%y����V�9��b؜[a�V��1�Y�z_�;/@�rȭ��$�C�yY X2IU*�/Į/\���=��:^u�Tt����Υ1
oN(XlxVHYEB     400     140�3|���y4	���|�	�tZ��k�.(ml�F�b����Ey��
1�� +��Weu��
օ3����)��C^9u�"�*�z;��KP�L~�u���mLq:#	�Z'���<-<=�8q
�6�?`#z�7���X��3l��,�w��e�9��������78��R�I��MG�Ԭ-�3{㿢�	��C���'���e�ib;���y�4p��Is��!��W����J�)��18����I�ݼ*�
>.�QN�P�3l���ME-dz�SD�W�,�7�9+H:��="��~�mi���m�*t��GXlxVHYEB     400     150�7���H3.�Ő.0�r��	[U�%wg�žB#��D�T6%h��l�!����0�%
pBXR��F\��,��w3�*�W(����FTi�e��2Q�F<�2��~P�����뿈	����&bh�UřIFa"�e˾O�K�6�7/Or5�w@gzgӡ�x�S�`�W�߽��Н����������m���5�A��Wn����l���j]��SM�᝷�����,f.��K(Yϐ�E�����莠����=mG����' ���OSn7M�z�bc1��J�
c��θ�ߖ�-���N�l\6�DKDZb���drI B�\�	lXlxVHYEB     400     110MK�[-;�:L]�`�Z��H�Cy�iS0�iDEg����<��ӧ�!���ō�F�ĮТ%l�a�)[���^�ͬ��Vr�q���m]߀]{*2��|G*��S���t���П�"����tzI��ƶ�O$�C�_����1�L��×������(�	�gi�0l[�����a�����sR	�����\!�}Ϋ��i $�
.����2��5�]�b�U
��u��nQ_�ڸ�54���5�������@�'хζeoS��'�rgXlxVHYEB     400     1403D���i��Y;�C�d50
c�\�_�����ډ��G��ԣV�c:x�h������Y���!�4�8�����C��5y�.7R.�o�4с����n��p1j�I�������P��+�s-CE/�+q�V��^�c�jf
�Kk;�����Ɯ�J]������Fp�yl�f��P��f��w��׳%k��j�����)��,�r��G�	ӥD�2�09kQ�fZ���y�S�+\�7��
 ��]�Z-`��C��Y'�Q�ߎ�W�m0���%c�}I����r�W����Z$u��ē_̈4��aGϢ��>"XlxVHYEB     400     120�x��hvNf�G��.v�Gb"����7W&���a��<ן��5�|�c���)٦�:EZ������,�)��vLsi0޸�1�����7�T��^OZ��u�M	Sq��1��<�����L�F�y*ħ�8H>�˲U_�2�T�0���7i������@��)��qH�YB�	�Q�k)Z�\_"橔m!�2�&5$�eҮc�Τ�Β�� ���Z0�FH)���̿�$��j{���p8h����I�c��;�$�
S��)M
����V����4�1�'��UXlxVHYEB     400     130�ĥp��n8j(�#F���l̨��pf]ޥ^ �]�<��G���T&����BM���fCM�r�����Wo�a���i�}M��1�u�w��fx�M���H�l��|�>D�6nAxD\�`������#��\t�8t֤e���ͪ
�KE����>(r��+����V���Xf	z�����~[������1�ʞ_GP�'�rM�b�B�����Za�[Ҭ<�E�?b:n���ȁ�907��$N>�G��x�Ab-�R�0���}�����J���{+�5o���ФB�4@�XlxVHYEB     400     130�|��V6iYFF��c/u��
���t�F̾;�I��k�P�eb��!h>�)�r�˹�֞�^|}�"�]I(��{6C�y�Q�a�ݏ��QK�$ٚ|�%\s'�i�Ht3���/V);�F����(��0Tf�25}^\ϸ`��B2��j�aT��%�^�9�ā3�EޯO�P�����5���3�9w��w��C���N�׆� ��k����;q��v��<O+�02���~QZ"�N�9��(���`H�<p���`��%�p�zo�np�Ϝd����X�"��W�^�U���o8rY��m�XxXlxVHYEB     400     1402��G�[U�ߺC�L߽�	3�D�;�E���3

��bƽY=�/�2����Yqҫ�w`/v�))��7�H	;jnsF?vμ�T�I*}2��������ĺ�[VEeFhkZ�qfO# ��ĐU�6�Z6WQ��F�B3Ǟ�p$T��;�њ�h@�i���L��b��e�YX`�Q��~���.,b�o�o�C�\�E�ӻ
#3�q�17�j� �� 4M����KXPl�R�i(�g�/+`����6���i������(]+�HK�� ]�̂{X���C�֩�x)�$��(�=�^�k0U��XlxVHYEB     400     160dbw��q/������I�5F��U'j�o�u:*H�N*��P��E���&�m_#������m���[�u R]PS/e���$NH�Xr(0���Uu�NUZt��g��uVP���7W����B}���^����	� W_�iy{om�\��vK�H��}�>���y�#߸���v�MKhܽ;�:��(������nn�H��ɻb��X
�E~�bg�Z\��Ip�����,v�Ô� �8���eW�d j+N}�,�u{�����u�δ>��f'j�t\����`+�S�x�"@6._��~��!D��7��]���k�\���rp�s"�=$���7N!�x8x�6�KnXlxVHYEB     400     100�=^�8��>���l�;6>��%�b��݋�Od�������J�}ʮa�s�1_"N�:����-��Ѱ���h��&]��F��~q����!4c�OO�km�[��������=RI�0u��yk膓�5�mgG�޽��UN�r������\$�	t�;]|�Z0}L�O�s�ѰEw�z���#L�]�cþ�����pf^|uX`z:���7`���E&�<J~D�aR�0=��;�A�ۚQ�æS�XlxVHYEB     400     150	K Lh�M�vS�%�hC����륂��ؕM=]��J���l:��o�,\M�J��-��S�D�e�7�&�����J[΄/������΂0y��[��T�t��� ����U- k٨�m6h��F�����gl��m�7�|W���O�H��~�r���}�?|��)[w�J����D�w�]:����(JI�5���q�ы}k"Q����z�Wb6�ᙵH�V�ׅ$ �k�B�un=������$ྐྵ����xS17���ۙGm��5��iń�C���u��2����SC���M�J[d9���5�#�S�Ǯ�O���@/c���f{���e¯�XlxVHYEB     400     120!�8�'wdv���NQZw�n��Oi���u�������6�X�*�^jH�I�y�h ��w˻�4�?u3��v�'�����|��+�aT��L^~��r��c�G,���R�Z�R�~�K��W��D�FA�k�f89N;��楉�[��c�{��:л��i�
�~������n*iKu��Pƺ��W��˫DI%�1Dq�&%��V���}�����^�t�6S��>$y�*��Q��J�����	�O�(¹䉴>��[���J�K��l뤮XlxVHYEB     400     130u�<�����]l|����}2�p�ζ�F�Fy�Q���A�d���1;_�dҿT�3��g�ol��};����� ÿj#zt��K_\�1�Q$9ל9AW=�h+\���$���,��d��׶��`��.U�'�a�mYr�KS�k�1��W�_����͵m�Y�t�T�{�q�#�c1���F���Kk=b]Nc\̜��<V�L(�%��)P��H]�$,�8�	��p�.d�������´Nַ|�ڛK���1o��&�*v�<%�����KU���<1���}W�JGBhY�$������g���wXlxVHYEB     400     120cL�nZus ,�		3����:�3�y+��������E.D|�8��¦�<j���T�`Y�R�_^�岓X��)�p�7�L�)�kRk*�W
�B�+��s*N`����^ɏ�[�0�c
���aZ�=��bq����TfL��9G!�p�C(�!��	��j
�x�}�Aj��n]Fc�^����7�8ΨF��O�4dV_&���	�Q�Q	��=�A��X6�,|��
���A�����Zٽ����\�-�Jν����Uθ�5�7/�&��=�����aN]������XlxVHYEB     400     140*H.��!��A=B��-�Or?�iou�P���c;\�ܖM���V-�4G��QW�x6���%�3��"��ѬGh��
4Seqc�b.�q�L�Ä��gy�l�q�;�2D�;U7T%�;���$1�n_@��n���o��Y_�L���~��|��:>1"��m����ݦޑD�ӅE@�6'�] 6�lLs�w�
/y��y^�!Ip��[=�g�z��H1�	�KT�+$h�ʓ~��~2��jf�[�ͤE{�U'���P���'�8&� �̩q�)�wA�<H:�1�_���p����?�Tzz���ڛc���XlxVHYEB     400     140R�j���ދ����D���U��F5'�ȧS�p��`�auZ�:M�}��"�6ShO&�l55��)W�����£��9b��߼�Z��?֗f�n@m���߱vzQ��|�������/ԺHZ��AT�w�W]�M�
J���C�SW8�7��I����h�w8E��_BB�xAє�c>�O�|+�\}K�LD�3:ibUX�[�/s�A���  K��6L\U���?*��Ƌt.��Ze4z����,�_
<$ܤZU"���K��>ߣ�<p�w��g����&���S��Ä�GZ�!�Q�@XlxVHYEB     400     120gcZ��g���T`�.���|>�T�n1��3�����oF��hWjj
�ៜ�w�8��];g}�mQ�����x�Ň>�����C�h�F�V�>=
Q�kg\��Mz�ܹ��,{'4V��5.+�=�?Cݎ���"}����k�(�^��lS�Z��P�6���
eIk�u��y�����V7�8E(�춣�TC�5@"|���X�"~˞��@��6���6�a� ڂ���ζp�W@K���X��أu�O�#��Ѽ���#�)O�j�P<�
�%�ԓ��qXlxVHYEB     400     140wf�E�p?�������K�E�m�����CVv'F���N�ϗ�Ο���LɮG&���4�`E?H9�ĲX�kO�1-��~Nb��uZ�T/��]����}5�/?���>V��(�"S��4g�F��u��Г���c��pϪP���Ῑ��M@�0�� ьe����c��J;���\���u�o�ƦwK^�B�?7d]��Ɲ����@��4Nh%���̙q?�LU�tS��	$U���4ia\�g�K˗Z�����z�����E��t�C���YD��Ȭg�F7dkq�l�N�֒[d��eF�g.�ߜ�{���s��-g�U�XlxVHYEB     400     130őz�)�4�P��!C���߭rBC0����3���e� _��BYzQX���z��������$�?}�p��?(ƀ��s�zz �k�*�m�{���@v1�u<��ySW�j% ���M�O�6R˕��2ng�!DB���M`E1�*�`��o�O�3�i#�/f�{ܳ�g�KXiQf9E��v؁� �^C�6&���/�hA <�%r�!U=��x�J�$+�Oq�zè�x���4�����ʎS��c�zy�L#
��DYeq��г��#�r$���ȠB��;7Pǃ��Y��az?����XlxVHYEB     400     160���
P�S���b �4c˲�fX:�Q�
f0�p�%Q��j�H_K�ٰ���zZ���!'Vw���̺��N>��@ �A�sx�˗P*����W+�d�ĈF�|\Jl͏ PB�%��ڽ�����~vaΒ���)�7�eVU4`/ݦ�7V�4�UX�7n��sS���ިF���k�Sh,����`!��6��1�����1 w�v���}�z`%��\yW���i�2AD�-�,t;��,]U��1��2��(F+jN�Y���V��Kv�w���g�1�[�}�2V������M^�f�����>�ɞ&�s���Q��Q'O�^��Us�G^�&u�XGsq�D�"�"Z�XlxVHYEB     400      e0���mٜ[T��]��^aT����1���A�
�m�\+�o����"�7���>���T���'��y6�R���\���L۴��� �y֗0�I���3f�Ļ�Y�?�L'��YxD
#�	�+A�Gl�a��R�% e�_Z��oQ&IE{R1�f�ts�t��e���Q�aMƘk�oX0f�$�6d5T�ڠ;@�8et��bVD�6j�p��QYZ�pXlxVHYEB     400     150��M7�25��J怍T���/W��j-�7��8���-,�L����`�X�qo�7$�1Ţs��a�y-O����#��gCя�G�,5^A�5*�7���gbh	է�F����)�!�
�=��S� �W!"��ȝ.�~�`gf�R�r��|y��q�N�fS	o�в�˩�-��c'�	a���T�2�g��i�'G/���+�e�빲nm)�{䡼6t!? �h��_�Vҡ��c���p.6Os*xj�HX2҅H�������ii�ª6�G㞑X[�9�T*��AA��\Ig�$��-���d��<&8��|�H�*\$��5�d!���y'XlxVHYEB     400     160;Ro��$E�._Tv!r;B�'ߗV��"��Q�xDWeL��	
K�<����m��`]X�زÃ�����*ovv�v�hú����BsOL�
M���`"4%�5s
y� p�=�n� �v�|�|�&�Y�7n0�=����60'��$����am0�zk��'c�x<���9��8�3ν�{�WH0�=؃6�Z�
�s���(Bo!���һ��L�I�#�%�ݐ�(�(�T���nr�38�l�����k�����uX����E� ��7!���v(-���p���KOd��Kv���E룓y�JD�z�9�5�w
���V�PI�_�1����Y��@��Ī��<;�ٌgSXlxVHYEB     400     120gcZ��g���T`�.�2�jȓ�^��A�=�e�:,q�L�.��w4�T�%NY��j��|��X�Uc+J�p��7J� 8ĝ�,i8Y�1���e��h|�t5	�aS��+,�8F�'�\7�x]75����j��u	 ?:���U=����lx��T�$7yd)~�I����"�aw����}�Ih��s\�7��.����͆����vNx]�&F.�#�֟Pz"�M ["��=t�u,d>[��Eoh�e��QL�y���0Fb��)��nϬ�w-쏥�4+!d�=XlxVHYEB     400     130l��_�b��	hLS�Y�S�sL�vu��O)?A�ū���}�����i����F9�����aP�tU.�	����U�5��~
��R�WY��k6r.%m������wBk���n؀��|�B� OA�N�l�?90glZY�ƀ��4����C�cpo�j1���mLyb�_��YĪØU?�P�m����*yO���抵�����OI�T�ZMજqR5BŻl��'������>u�^�^�"y���;��W�K��B0uݼJQ4z����x�g
Mr}Q`�m{��XC
?߆M� �c��st��uHXlxVHYEB     400     140�+��;���)oQ	��Ʀ[�>鶫��Y���0��|��l�U���STm[e���V
��At�!�-F� ��.	{�O
�LP��8�E��F�ۂ�(�$��p�l 1\�1Yo���	 [C{&������~�����z���`�%�G]�{	�sf@x��p61�)Ya7 ���GQ��gm-"H�o�{��oH�5d~�R���lr���� ����5�r�v��DdS�-���V��t�GdgTc:X`Y8���Hb���x����a�H�x�S_@Up����g���m�+z(8Q`�KMz�Y�����8!�XlxVHYEB     400     160�k��dh,&̯�S���#�̀F`�$8�w�{s��<����.h�6��8zn���Ix]!:L��	�+��sODP�r���28���C�w�����f*W�H|\�,�O�&�#����};Wi�I-�4vs߄oD��anG�����Y`�sT�B)�3'�G��čV�B#g'�q�6������h����ؑ\m��yGs�F|Zc��5�s�~V�*؞T��OTf��gb��q2�aT�!Aʠ�>�&�K��!����@��F�Z˙%PW���_��8���\�`ݝ�J`�aR�d��13a�F?���յ+�?�����!����Oy�ĂuXlxVHYEB     400      e0�⧨v�gP�]A��)���#�F H�l������|h�,\�Frv�0 X=���WB#n��=�4*�	����\F�`AGqy�y�J}'�����7PO��QLWwpP�i� X��"Fn,�[h���>g����Ng�`l׾��tHc�0�9{��}{+��Zݻ��@�_���x��VT�ǻ�#&g��v�dn��;W�\�l��}�s��$�[��U�XlxVHYEB     400     170��s���dE��y��$��	�
9�Q����sl�U}h0���N�� �ޖ��v�P��_���ؚZ�= �o����@
��H![���I�@���;ٞ3�Nn�:S�8���#4DhQ�;$����cc�����)���y�>g��yĴU��a3���Z���,=����ݐ� ��>�W���t��D0�7f�l�> 3_o��ڌ�#b]G����A=_ I59i(F"��D��	(8C3�ZV�XO	��9n����C|O.S�����a޻�ןַ���h�V�4L#>��y��+��2�����;�W����S@j�&�Sئ�5�\16��_�d2^YHxOb�,nS��Z̖�����L��ۄnH�m�Ρ�XlxVHYEB     400     150���D_��vqM�2��C���#�@���ۗ����[Ye.[xS��`Ѝ3��,�ުJ[!�r���I4�.�(�cZ�5�8\���iy��ه��7�v��V�R��1�{P��r����m>�x��p���P#jZǦAO*C.I���D=���ם�������@����<smZ����3�@��0�_���p��k�9z[	�G������1�c�6�y8V�Z���՛�1j�c�{;�����vDj�b������6)c�o�(Y��� ���j�0��Y&�!��a�X�J����`�"�gϙXy�Px =)gM;{�r��2�q�*b�XlxVHYEB     400     130[d�lk>�|��љ�M��d��kP7��a�^��ߘ52�l��F*�D���*Vt������2����4ww��Z]�ONF�c&
�HK�����Ct����}��B߭�/�Eĺ�4�@.��y�C��*K���F�%/���o67[� +d� 
~��q��i�2x�kN>�7?�,��F��8���!z~�p�Z4]�)L<3x� J�CJ�K���HǑ��`�.s�3�"��TF��Nk6��Nژ�.���Z��*���2�)����޴�~�`j��"x��Y��E�T-�o�XlxVHYEB     400     130mG�h�.��Ě��V�_<��6�C�����{���Glg(̏����g��H/{B^�_�X�9�l����Zɗ����-C����dZp�5"���Ik���(V����9%B�����k=�'���%Y6���A���g��V؈8�~�{���yP�o�5�X��>�*�Z�� h���0���1-��*�z�$�\|��ZVQ��g�5{O#�S�.������wp��٦={Q���LX8��طژdY�G���Խs>��
.�z��ϐU=v<�+5�KJ�ׅ��1�u��/��Y��XlxVHYEB     1b3      e0C�D}��o�D�e��J�-&+�T2����	E�ԓ��U�� L��5{�8�m7���ڎ���[�ި�Xm�땫#i���熟�'��'Yn���Q�w�@��øO��5~({�ʡBG��d'9#3�L��(��>y�P}���P��y�_�s{x|���Z��Җ`�FÇD_��ށaP<�O8���������:��1��_U.���U�v�"R~�٢