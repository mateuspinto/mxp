XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'�E�H6R���6���p���kLG�pu'�iU8S���<xׂ��pT�S�����8���������b ���(�6B�����2�D	��&�gM4p9�h�W�鐴K���v�yŌhP=l6$���nr|�~�4���^q8W�$t�(�����fl)�`*�+&��7H5�
t��?�&�N�޷�a.�7�G�)���i�16o����^3�X�۬�N�l���yz�5�c���~r�pٔ��s�QёH�Jgh�D�BV4!c���>t�Y��T�4� /��cE�-6��L�Қ�*��^��aȓRb�L%�ufbW����Js���%��>P��Sg��U���x�?�s~�<iZ�<�~��@=�*� A�+���TN�.�v<��3#�V�61�\%�※�].�O�[3w��>��?�U�	�	$q��8!������ћhȱ,�_*6#L^Oj��LK����f�����;̋��%��PK�_�c���I�寑�T���a�v!SV������B�w1L�x%h�k�gtrP�ȅ��6^��/<�y�����K�h~N!�F����x�5V�Io�Pw�dŚi!K����ʑ�!q�q��q5��@N ����l���b'�'̎ �*˱���8���8��R�VAdG��K>Y���m��l������B�eV��,���O� ߲AhMq�4q8�PD�lc���-t�-q��V��QO;�(������|���nmw2�y���;�� j�XlxVHYEB     389     180p��Zf�����[*�
C�rj�U��G1��4 r�����:�y?��z3��=�̯��#9V�����k�L�@/�4�=��s�����5����)�D/��TJ$X��ߖ����"�=�^Bg�˧�4����Z#��J#�_ �8�o��͎���W.*Bc���c,��S�?,+Ȏ\ї�����<ַ�r��Ҡk�0�+!��D�4ы\g��W��ƽN��5�Bb��.M�����j�p��!�B�+Ѓz	&(ӬM`;��Aֹ%�`�?x�E�A�)�ҍ�񾗿��D��,�N@,�����K�S�I�#�H�N���ˇ������W��߅W��#:��&��{m`������b=��_�Dp�k��Ƹj