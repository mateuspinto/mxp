��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���Z]�� �+J�?�ɲ~}��R��C��֢��=����7�����@��Y4rA���K?����X/Kd�h��?e h�S�H,�^�J���׎�1��
4�!fQ?�Ok�f�@����Ϥ焕GUH|(��H�5
��fw?�S��js3�r_��1������htA�����ύ�&�o!�y2kH��$6��KO�峟���{paBw�%s��e�h28�A��FC������Xz����ֲqy��Xo�b�:y޴95�Ѐ������Ĭ �[���0�Y҈H�[Ũ��Z��̏�����	�/���=�Y�"���:�u� w�z��|���ѻ�Y�]g����MdWev>G^���:��Z������k��O�2��Sr�EҔ�X��8�G!X����̞;f�+��-]�[�԰>z'�1Y-���++�Z1g8���@
ݔ�MA0.���\|�!_���`���9	��.B2�	[x���v�&���"�9j�K�}�Pn��Dg p1O��e��ʡ\5�7���|BT|HC*�Ai���)��ɛ�)���5k���_�0t��J��v����j}�x�W�G' �����n��0��7�t`��*�?Xw%+�7K	V�I��S��m��)"�����}�.�Y9j�u	�X�G��q����"@<v-�E�sB.?c��OA�-�^��HS��1����Ҩ������>HA�W��%�������	Qi�Z�����}�q.�V\���繐nU���M��4��,˯1�}�櫐�
��X&B�n��SD7����
��N`�n%��,"��3�E�+O9̓T߲�!�ċy�x�x��'X�Z���V0���E���e�Pu ��o�we�^v&UPY��9L�V��2��'K������H��,P�~�]]S5Z�4Bb=�Q���+8���a����,�v���(pp���Li☆Kc>��}���ͱ�Zdn#�f��_;$:�AC�D�^�z7B���$��͞��"0�,���y�,�u�E�����g�7[>(=�b��!�X�'~@�t ��5h�R���	�����^��Tw��ì?d��S������J�h��+jY�iER�1}x�^3�@��2�_9vGE�#�>����B�`>لH.*���thD��ά	�����#�yۢ��� "��k�8�2�qh�!�&�,s*Zgӫj�sK�/���TG���7꭛��Jz�_9@-Ф߽Edȅ�;i�h6�X`q��x�����Q?5�g>�u�����X�>4	&�zS��Q5�ME��>���\}��;��~ł��?���ɿ�^���93T�v����%����b���+��%ܲ +�R
"�n�����R�|���~"���`��.�ws�7��8E`?RR�Y%�����~�R\�if�teT��E1�2cq9y��¿���LrNl�^oSvZ��R%M���0hc�r�_��5�L�=�ت�D�ܝ��5@,Q�����}V)����7a��:萕:�@����CP�G��l��	K�eI��:��%����&�}�85f�	��wB+����H�	���W���_���1s~F�S��a��q�YD��������,#��EHG�;щ��'��ƛ*��C��ׇ5���gL߭�)�,�o�8�uه��DCʑ�����5RIj�ӴE��o���~�$8<���w1����)�7R�y$�T�KcI$(���Y%��t�Z�.�F�����D����[q�v5ꃥ���'s�'P����It>�&UpU>@��v��ޗz3tbYT��#�Ɗ�'�R �<f�o��E�9t�Y!D�r�(	�`�XSF�ε�z=ȊYc���/��O$"ʞEL�Ixf�_V�įǧ��ß���\����i��ҁh�A�6��I/�@q�]9�F�D	<@�7������q����.v���C�c�ߘ�/���(�taE��8֓�o�=�qClhv\�O[,�~\��s�UU�)���9���	����W�lAH��m�� �D���"6�ѭ�Ɔ�j6�7r~t:�����.��
�R�e�8�7뮅�(����B�;cK$�/��v�+d����X�)"�B�����FE#�o�Q��BG��Z1�K��s���� TtUB�ׄ�F]�:�Բ	�������:�ہHW1%d��F��֛���jf�b &��{B>)!y2#��g�n�@N @�`��d���^��_1< �=������������G ��mE۳�h��x�qUu��g�&��DJ�����?���#�t����	y_���3"'��HrS���J�si��Wҁ�@D�2lw9���XxV�OG3���N�����qq��Q�p��
| ��>T�%HM�jxF:�z؄3��Y�5]��!�����v_�¦_�&�-�Y��"F"]7'~�"'BC`"��<�y�S��|�09¿u�b��V&�L���c�5�Sn��`���~�����'�4�Z�e.��{�t�h�̎�f3�&�^w.=\��R��N$��N�5	2Ë��KQ(�s7�4��I����Qs�N :�V��5�XIK�&=M-'����G�1�c��?� ߡ���S���&-�RU��;ԹR��(P��1����H�l��kV ���f|޹����Nǯ�\��O$(�9(Jsb�lM�	��!���,�/ηY��:��I,~�o�J� �w��%�#e�\}�<��#�F;�Oo�j~� �E]`�xAF�
TfS/�z�*l��.&�E� ��gg�4�k�#��%<�,Cm���H�
��"=/J?��k���N�^��TA-�	��RtE* j�Q|��3��	���w/Ed�k�5���(.���L)��<%�����b��,BBö��1n����ߡ�	�A����%���&����_@��@\-4�����fa܁��M�v�x��(��V�'ժ 8HH��=����Vج�ph��|��[o���|d��1��L ��su<A�a_��7QRϰuS���̃�u�uq$�6�[䰛-�<gw�_���ʪ���Z�rW��:k������A��+����+�Cт�u�h���tl)<��TF������7S�)��v�+�"��q��k���/V�gK��	����=(4 �*Ӊ�'�0�#��2���v�d����Us-a���Jh\�5��@��;�|)�|+R�o��Lqi��K�p��+�8r�xW��i�Hl����J��XI{p/�