XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� �)�HY��E�7�k�D�S��&��ǳ�~*O�C�
8����}6!5����8<�zkd~"ښ���&�K��S�ݏ�BeFV���>�YY�c�֫l����/2ڢ>�[��aR�=D�V*�:8ƿ'�==FF����T/ ��O	�5��m�#c4²��`�}�fr�nZ��Q��-�����ѪH��7,���`����a��������P�yOP�C�Г�4ѯ����Z���w=��r����?�q����k5�b��66&���%yY�YC|��p��p]"�N�/(��Ύ��^0@�$�ho���)�*���|��
�E_�:��h�M2�5G�CjJJn�%���M�uG0"�X ���B����f��z=.�F6�k~��{b��̓OP\���O]\�n&)dmP�T1�c�,>J:I ��?�GYC�	��%���ۏ��5��~�R-�<�i왞��ӊ����A{��nUg��	��D�5����
�d���2��ϔ�8:�)��Ɩ���ws�ev��d��I��u;��&�������{��tw&}�qn��0J���%��Ij�2�#�
t�U%��%WF����~O�� 2&ˮ��ώ�<b��fi+P�1����.@�_#��v�WJ�)��*�|8��=���EC@�hV�ނ<P#
�=h��5 X�gJ�s-�?��Q ��Fw�2�Se�+��#���~��]�!�OT��%�.�M�g���I���b��K�#�XlxVHYEB     400     1a0%���p�ébj�U�e�L���h���@|�M���ĭ����O�b�E_ⰸ�����h'4D5E, ��ת":��]]�N���^�\���'�D�4�)�
q)���j~&|��M6�y_[���h��VvHD]��LU[��"��ʌ������������)F�+O���~%<�
gb�o�"(�l�Z���<����O���y��T=�J�V��8��lȴ
l&߽�o�+��?�0?m��e������+�=�B�R�R��	e��1|Y��d�DkK��v!�Zm��\�,*�f{3'A׷�Nv��g�3y�Gxd�8��F(@�axn=@wYˮЇ�m�R�p�n��lF�$I��q�;*i��yZ�<R����u�_�Eҳ�]����k�U�<a��a,5���i=����A"Yo�XlxVHYEB     400      f0��"� �h`�HQ�����;�Ω���Q�Ɍ�}�Y��X����K�� �	�0N�[�;lcY.��߄+
�vP+kC:� %�r�������$R����2��ɽ/� y���~�I��V&`����%z�VP[_�_����F?:F�Y~C���^x޸`��[�D���7uu{�S���R�t�q��Ni��9�Lf�����;jR�F��#Y�l<0{-���Z����t(O��ds~C/�XlxVHYEB     400     180���6�b_1�����(2T��k/��9,d���W�1܆�5�g~��3W	� �{g���4� �� 6����ݰ��]P�J���&kv��%��-�g(��~��?XnУ�W�,�����T��m�u���~����U�+BU�������"��s��FN�o	���������f��e���HSh��K����ynD�\s(e�_�T�ҩ�9ΨW8�^R/���8�t����V�q���2���@j��9;w�'��;���𔁧��{��|G�K��Y��eGPsN���Zm���@g��浾L���N�.���dg`��%'��ܿ�����DFl����^I���&�NY�X�zx�i�i)�j���¼�X�R��-�sXlxVHYEB     400     230
����S��`��KW����LG5��7%�	`Q��������J�w�g�	r��H�)���GՎ�}t���ODC�߈f,���K� zzuޠ��ю�;���ub�捆���G�%��Ҹ�ҭ�^�bg�~�n�+b���>�J��?�E��߫3�F�`-�պ$�T��H)��JCQ���/��yE ϐ,���j�T�)���W��=I4�N�f�In
S�\�}��{�iMgQ�0� �֬xl0)J13��$�E�c���\6�6uR�
h���aF�B��Ԧ]$�J��;���(گ ��¥���k��$��p�� *��p��׻�*Z�ho��Sŗ{��XN���$��ã,3W��Ř �dK�ҋ�|�z�1�Ox�C���J�Jp�c���(m�r�IP�g,a��Hi�Z�$!�F�>�W�)���)n�����`���î�5X�o�R�� � M�ʟ��Z����t�5��4�d�-��r3-7V�)�(ErlWH�wt3q�-�x"��f�J�uD� ĭ�F��Ǌ���Q��5"Z�DXlxVHYEB     400     1c0�nT>5����4v���$��)-8�9T܇Q�L������o�?��&k{�"wz�t*Lt��DWx�[�cSUV�P`D˒�ŏf���Ej��/��CQpQz��*4��B���������.�;<��ο�ܒz�[, TK۶�y�;3�P˨�=�
-�POLv+wi`A��-^��q���9�f��Զ)C�v~�����X;o�nwe_��z
gՒC�*w�>U � JO��ڰSj�સ8�E������N4Qv}��ol�2�
�9�t�r��Y�,�l*���q �^`��,Q����g,'�x�3��S)雬���G�Mp3̌@��^�o��f��m_}��
t+���������>Ӻy_���B^yQ��������k�b�e����lc��JdtX�RU�Z�$���(@�ətj�w�ޮ��Nj"�a�!�XlxVHYEB     400     1a0N3TU���x��;�z�z��pG�1Ƞ��uB�MJ�
٩�����
U00ݲ�C��S���k�M	 ��z�P�4g~J������i��4�"��r�و��H�F �bS����oh;�G?�*��4��1�1�9T�9<�C.H�xW[�Y3jU$���(��"�]�C����X��_����TlPM��+nT8瞗�Ơ��^F<�Fۍ�Z:>jF;��'s-���)h��Y��xbU���� ��!���A�\����^�7��╆���3d-��s����F{�Jh���k�1va���9�3�1��5'{;���u��M;I�E�����Fܛ��q�}aD��v����U�����<^ǫ�K��b�E� U=B<�*x���ruH;H��3~�wC�BXlxVHYEB     400     1a0�L4]0�"Y.���.�_=Up�,}Y����h�˾t�Y�j���U�HBM�fI�)�^̄�䒌.���]Ά\3c��oC��M��2�M˺��[_o�1����H��w��G��g�5��CT�gq&"�<u7����n|���� �0��x�qp����oʶ����^���� �������詚D_w>m r��3@���+Q�*C�������Z�1��ב�,�>	,�S���O ��&=nn�XW˲��
�젫�3_�vRqT�S@BS.N���4����!��>if.�K���GL�`����^�Ǥ"��ϥC�l�!X�l(��!�R«��`�����4� ":�!5��h��t��ʞ��,m�f�$y��Y�~�Z�����T�#3G( XlxVHYEB     400     1b0�.�=�'�5&�]�,�E�3��5D�a��v#$v�9�k��kB�4jt)G���Yo�V�Đ�v�jged����HK7���	��we��R��.�j��ft�;�K��׭��׏���� 6��X�e.�N���M�������6�.e?!��D�/cn����Q�yW�����s�V@etk����_Nx��Wk�J�f4V�%��w�8��f{���s�	9`a��%G��#9�q�gD�^������FS��W)_g$�
D\���S�ÈXIB#m2u�մ-#���͇���4��k����$��`���p���X5��y_>�fUjAUŌ��So�5����v�<~�4�f"Fh���(�l�Ug"�O��_�^�!Ż~)��$��ɼ�azvhd{��\�<�W���\�L����XlxVHYEB     400     1e0OM��}U�SK��V�3��葤���i�Qy���9q!<���Ⓠ� �A��R������X߇��cvwZ?,#3�a�%��ʚ�˒!f�pL�Vy��os�(;�%� ��MlHp��Pޓ(��%����)��E?���Na+�a>�P!‌�>%�#6��Z3��fOO39�ZסE���}!i�	E�t���$�~6��:��k�����T}�{T�<г�X&1?.I�(�C%@�F>`却%��mv^�G��
���`�2c��mi��Y���D����_/Rm�)@�}�uy�d;�%�$��nKڟ���=Nj��fcPB���9����~J��'�Q�*���w4���sN<��S[�Y�	�=P̉�Y>�84��^{u��رJ)�?qH����J����Cf�6��'�?�H_�7�����UJ��ޒ.:5f�����(�4x펛�=ƿ������׼sk��eXlxVHYEB     400     170���BJVB���y�K%��v�cY�-���
��QFPn	��h�:�aͿ���rL�;l�gH��E�C�Oj>?q@�&]��+���!w���}Tw'A��TB����d+�)�8��*�S�E�S��w�3��/Y���3뒾�ʸ`�=@���70g<eu���X��߳�LdL,X3)�R�E:;� �u����-o��u9�����E��_���k≳Ma����$+'��x��\�/�~u^����KQH0�C��Q��y�sL�&3�G��+��7�s֎�����o�8���z�ѼJ�N��ǌ<z�5iA��V�Z���:��L;�����䷝�����OA�XlxVHYEB     400     140��j�g����Sob��F��QE��	H_��
���;�z��w�������{�8V�Z|��!trM@ꪄ�<H���?G����i�e�ea���T.
t]�H���R1��|]#��j$u�@U�06d�U怕���0z���pj�� �!֟�������UA*�kMnי^n���>I!w�9=${�v��i?��ʶӟ�!�|C8=YOzi���t�[ѯfnY�G�'����Z�:V�]X����H�u:�@�c>�ſS٧Jr�<�����Co�z��?�cO]�_��Ȍ@��I�?p��`m~tք��%XlxVHYEB     400     140;�qcA�(�)rƝ3QB�&��g RxU��p��9u���3	�+���:)O:O�9]��U��)�8B�_��J�b%D�'��h��g���üP�}�ي*�����Ml���=\�.�G,�]3�@3S�{}`����Y�F��w�d�������T�H�
�Sb)C Ǝ�\��x"�:`���`��Y���U~5&G���4gR���m:�m��;˱W�U���=�}qKˉ��:�$�}�z\�ƧԼ-���k���z3�^핇4)�^�=�]��JgF�@���v�� �=�яM���?F���ds4�o�T�G��߇XlxVHYEB     400     180Gi����I�nE�[Qi֑�s�z0?0��"��d-x�G��O`�}=�*F���R{��x��Z��E'���7�81T�G���鐂=�\z��B���`���<��0��9r����x��z�r/%��hb�)U��IV,zU_�X��R;M��I�"�{�����~�����D?�'��Z"W�0��X�G��S1/�u]���{Y���w@�V�O��~�ӱ[���S'��c�x�G(O�*ũ���K#/l�#4>n�)��/��>�+�xߣV�����uͲ���V�oDco�.D�6#�ޝ�̨����ъPǏ[N)p�R�ͥ����+�gK��N�	Ժ8�!9��7�w�۸w��V�x�a���:���X��V��]F��<�CyXlxVHYEB     400     180����ˑm@Gw�?�/�����V�H�?��v�ST.`�=�"���>2�����L�V��z��/�-ѫ�ar�����>I��P�V`��\�N�r��(ť�t:0f�	�&Xoh�.�U�Q��ox�z5�?�L5¹r��BЋ~YI���?6��7�U��v�(�+P�����'�  ��TΒ����@l�<ڹ�k�m�[���>�9s�=�%�z�ٵȐ��fϝ���ɔ�KxW�"M���A���hC��I�UOe�QH�[/ʐ�m��3���@ �N�*̎�B���Ԕo�Q��h� 9���Ry�������<��>��xI��+s$"��s�[C���rϏK���c�\g
�m��h��,��Un�Z@|m�XlxVHYEB     400     180_e[��R�^dF��ű��XX����F3� �t��ʲ����;{�u�:�z�4�u"@�7��2G�_�K�1셺���I%�f����� HZ�?�P8�� ��c�y�?���TU�!f`�+�N$�X��J�l�s�p~�-L��2a2�~1Z�qϴ�����ʡ�#�k�`4�U��U��}�գe�����e=���phE`��L������`��.�џ�˭ÎJ��b;�YJɓ��"� �|/ǋ�W�Ư�ֵ9FJ�����C�ЙURz%e�W��ٻ����A�ˎɔF]oFd/qx��t�H[���!��vWC֡l7s�Pb�CR��p��&����r���^�j�'Z��t�5�l�c��q}/
XlxVHYEB     400     1a0(g�_L"�̟��!.s@%fD��o�w��+���@ʺ���&ؽx��!��ɺ����ɼX)�D���u�Xq�\|�"������-H�4�4 Q@��.�L�O�⟣�t	1�q\4�͗gw�ZS�{Шoe�h�����Q���>�m+��(sfj斅ʷ�������#B��{��
V�]�;�zŀǎSr��u��Y��b��61qX��_�"Ã0�����ɫ����	ޠ�g��_���k.r�8��8�J���͖��&��e:@��K�LP[�٧%i��]
����{'Fh.bF��^;ߺ�tI_�M��Ш�&¯�#%�i]��ʶ��L�A��7��J>�i7�	��"�Bވ�=�R��������>��7d�OޚJ)e���ki�������eҴ^�o�E}ٴ��.^j����XlxVHYEB     400     1a0�$��f�T)��(ۤ3տ��qu�^��CS��l�0J�uk��
��)��,��VŞ$�����Q*u�]��l���`�gЖ�ӶN,H�Ƈ�n���,�%-��I�f�%���}R�M����u_�,�w�Pց�	ˮSBO�����A���\}�����5��GiJ6"�y�oC�n4��$�^�m�۬�ۀ��(1z:nZ<�j���M�|�Qb�Q������h�p����;�Jc�����I�yҨG�P�H�kn�p�2D�n�ð�W��=$a��7�ڥ\�`"MP�J,.R�������>��Ԃ�G��D�f�9�_]�Z�v�^(�������y���/�q�I�%���U� m���t��t�,zP�n_���6˥Ef���i� k��]?4뮎�W�m~��YܼZ��H7XlxVHYEB     22d     110`�`�`H �OV�n���R�qB�VfG����x�3bDeo�%\ǚ�fKRt�.�'킙j�*�Cn� ے�$��+�&�$;�k ��3{��0�רz�FcLp>�9p�6[W��m��*'�X.��<�ȉ��yQ|h?-�Yo gø�ǉr�E�<К׊��>ֵo��ǵT�1.xFq�E����h_��A�w�WO�ܒt˷�`+�k>�@���x��Ҡ��l˺��[��V�����˾<�AͶc����|�Y��g
�E�ʜ#78����