��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��в�{�����2��͏	�o(>���A��R!���Ϙ�.Ѱ��Ԅ�q�!MB�c�x��P)�f}B�h,��2�)y%_�/�e΀=�+Nr�]��Ċ�bВ���ļ��m�F���Q�ZB�2/e������!���t�So�g��Ĵ��U�q�:X�k��4�O�2�=�Ѱ��w�C��0L�k��U��H��b�`w�=y�Ju�pJ4��l�ub�f�>�"�L�~�E����>�(��{��rx?C�sC?�Q́�����Fd���J��<���	6}��́ �G�H�qظo�����?��i���s�D(q|5+J�](�Ɛ�g"m��(0��̛z{���j�s�Ձ��:pi��"������irO���K����5l��#,�{�L���Yr�#z�]�I;�2{�����:�!��G�T�O�G=!��'�����&bA1!����u�</`ζh���䴸�X��]@�K��I�LI)or������ FΌ�S0Q��P�� ���!�Ȣ��Q팿T�=b�&���a�c���i��i
��Ϣ�Ll��+~��������i˾�R�?eo�	���ܫ�Oq�:^*t��^��X]x�L���T6��j�~;[��w7��QS
��s:8_�m9L���ec�p���I`r�?!'cD����
פ�xM��*����+���	�%O��Q���V��{�C��=�`��c^>��Ȓ<��iH�l��?���������估$*0r8<v���s�aK>�53�q����j���AG9�~� �x�nO@E���[�(E�pH����>;���^oZ%>��s!7ٞ[5�\,93B��{)��{8�.���@�m#U]z�&�G��?��d�X�^�eo�=;B��Ii��W�YiP'����͛y�E�L'ְ4 �Q��u�g1p������&�N�+3�sV��H���d��?�7BZx�0�ְ�����f8����ˏd��8�jJƬ�h���Fx�zG��W6��2��]\Ɯ\���O�xN��'b|6�����nJm�ie�怟"��[j'}u��������Ŷv8��w��V=B�^�����έXt���H�^��Ȑ4�Fl�38�MDc�Ꭻ���_R��3dSk���\���8������/�UTHi1)G�Fk,�� L�y[���Į�MRx�,�Dg��N<M����dı4��ߖ��A������VsB�8D�(�we.�(ͨiX��R��W���҃~?��_c���V��q�Hh���w�Ӣp�B��<J�/c��ܦ#��~�g�åBr�v=��$~W�Q	�Z��2ͳt2U��̫nE������K	 ��Nyʒ��[�N\���1ƛ+� |z!��w��#�"�y��uI0�W�����.@F餂����Gn�W=,Fe:�5���-����kne��O+E-PbBl�%��ۓ��k()�ђ�i�"���n��;�IuC����?0�U7jf�N�S!@ql�>��J;��6���K��>��T���8�m�_���`⪲��1�7^H\�߬  츎܃ Ы�� L�3��"3u�HN��^����4]r��t���ɟ+�|*e
ؽ��?S�����Z�5���p��m�Y�-�Y'7NÛ0B ��ʿ<�G��*Nag/˜Ş0�:��7�G~,���U�T��An�;�@^8aM�^s2�%�>R�,PMff��`9��W�[<�ɦ���_���X�W��m�hN���dm� ��݁�uд-�*�>�ퟣ��=)Րޝ�s��1�đ���Wد�vo��bZ�X���ǆQ��k۝�ߊ���Yq����MpD�Q�t����᷸��f
$���[�Y���R��7�k���H <�V��.���>:K_
�#6��wj=UY?���lG�ʍ�lQT�1�E��$C��3x�̡�Aj�F/
k�u�W��)a5�\rAg^����أ{��L��]'�X��a9?b�1O?f���le@�r�B�Y�_,��x���+^bb �)M��KpWZ�>��:��s��w��"V嬟l�a�o����1G���ts��	�:q�サK k�~�ɹj��z�N\x�����q����	E ���F�]g�I�t�vv�{v��$�Uܔ�n���ΐ)	0D��y��etuT�ry�yF
sEm�!�a�R�F;_����'� u�o��d�..V#U�J̅P�
A	���Cqn�o|I���ɯ��ۊ�}��Mjp�����r��YK��_��Z�#�D�U��w�O!�<>�[�SMt�ZC�5���V��۳
�u?���.�`�s�ǟ��෨��(¥"��/=��r⪇�R�v��0~_=��
 ���ݨ73] �1i,@�M� 9<U������:�g�����mn��Q�'Z��7�~���k�ƴ%Fa��e ۆZ�Q��,r��8~��P���T�j��D�#|�]�c݊?��w�m��:�?7U��g�JJ�$ݼ]���t<�)Wm1�a#\R�@�:X��af(�3�@�8�l@��/�V�;X�O����QJ�ʎ,�r�lkgq϶�W��a8��i٣v����m[�dF�yR{�a�N�Nl]W�����؂p����`闂����K�1Ν��n!���r�~���dt�J9���.
�Ey�弑Y�=^Y�6�k���Q7�¯��_���`ڜo���r�|�~��y�i�"��6�T�����j��m�Xi��Kd�u��l�U絑	�z�pƙ��#)�vU���r_�r�4��Rur�����@�N���3@���nw5��tU��# G�I�yֽ���U���30$�,�M奲9�M ��W�r� �q­\������;;ؽ�h9��,�ۮ�]Jt8�Xq}n*��&��o��N3��F�!����Cq�q�����Q���R� -u�!�q6\�I�bk�l\��q���a�6�ضN���L3Ą#+�࿯x
�Ρ��O�� ��2kޯ2p���Bt��B���_���t%=) CT�[��"�|���\��~�J
_��f#Q��%�w-C� �oL�y�⋷qHau뮎�Jz�z����JL�d8kz@�v	e�<�O��P2��{Uh��'�+j2�(��C+m}���(�wtRdY�=M?�ˈ,$;Q��^Z|�����c�+�Y�#���F�x9m2H��(�Ԣ��𼧺Yk��g&�Ե��Z�_Z�e}���Z��-r���{����]B�p�qp>D-c����]������SLǅ��A��V���A�����{�Z��%h���(���:�4�E��0׷o����8��w�/��4t
�����������{�{7(E�!�mq��'o("T2�~�.�]&�!ޮV�@S�H��>Bz�s��ԺE/%7%M���D B}�wΫ%G;�h��2�~	~�Z�n�ZAFr[�����ߓҧp6?����х'�ի|�(�G���&������Dr[�ƚ46:ej��cQx0.ƕ��E���K����7���G��P�rf�&��ҫ��KK�{�����X	]��W�SX�Za�T��!�Q��;�GKی��	%o��vzۙ��������Y�)�^���U���+VV��8�X��`����*�I�]�9߰�m�CO�(���v���Z�&_�����x���,� ?M'�x.ݞ��P��L渾|�MJ�s8����ECR��(}�f��uWf3��C�W,�36ި��r]8Ugn�nؐʉWoܩ+
%��+�3�c<���w�S�b���(G��d�8����d��7�AK��y��p:�bAm�J;��;��9w�_��JD�ҋ�	�Ax?�����^�e��	v���ÐЌ�Q.;ջj^`���`bgzIP��4�{.J�#�</�	?WJ����g
�/��� ��UP�����!o`��(c�ƅ~�C&v��|�B��w���Q�Ɩ�����T�����z�(�`d7JL�1t�M"�;�s
}tbDw�E��I��kkH�eXd��a�H)�q:St�B��IW9E��\ ���:����M�zS�2?,�%�fz��tN[=�-��5Z��n�=��ˋf��w<�ݎd�dv�=ڹ��B�����!��gݢ\+��=k#��[�qNH�v}����pC�P��7]�
�u���[F`Ң���/�CmB��&g |m�cSʒEg�u&K�����VoN�>;_���w�E�F�fؔ	/]R��ZuA�Y!g,�<3�sx��St�~��j4����0�K9_��L��OF�c��t@F�Ҧn��� ���uw�&��̬�O&�� sN	���u0�*�h�B�g#vwHR$Pw��n��q�ꤡ����|����@3v������j�d鿢�'���2����g���k�ձs[�e����{��o����B�{q-kL[=�\<�⸠�fo���	���D����wW��-i葹�Ӹ\~kµZ�	���)�b.���/!|I�)�t��S�f.H���|΢%OɈpEфj�]�
�P&�%��<{{�j菄0Fc��@NBz�^wDc<�M�X��:2K �q����f�~�8��ސco������d�e�K_+;/���ԡ\!|x���u�&� ��P��=�:z�-q������VvM$��a��"ڳ��}M];l��B�"�@[��Xp9��q) ��o7��tZ��"���ŀ�=@&���6��X3'AbD��C�Z�X�p��ZK������~���]�$`S�&hb��"�C��>t�~M�桌�_��_[�{�r�!F�����:������;�x!��"�q�E�YH`��:hV����˨o�ݴr7Z��2�����yхy@��[���-�F�zi��%QƷ��ޚ0A��2M=��<��˝
���'6�� �3I�3��p��J��ga��넃J%W���U��i�:C>pA��X��}����i�<w�wޱ�s�`��oQ&U'C�Z��o�`��9�W}����	f��q�6:�y�Ȍ��W�%��y�^ ��n@�	M��x��r)@3�V� �'K�5o�i��p%���������dR�|�Qnh��r�.(mQp��N�>3��Y��D�b��$��,�%���[Lij�ym-���]%�{��@�cT�K�R^ ?���0��_��%�o���9���F���GSX\ܳ�-�O��'�rpZ��x��w�Y
�V�q��FV}u4��:�}��my-u�Dk�{��Q�|)�.�X�*��/��s�#�d���<`�s2UJ�	z��想9!�(}k�Ї>An�q��]bQ�CY�^k�3�0ή�;G�&��AT��|6�Nj9R�7�zIL��e�v��vZ��g��|�$j���fS�`�9R�`V��E+�C<��Ɯ��:u��އN�T�g%dh�J�)�0�I��Q��Jy�[m�T\Ey�^��&���G�m���t(1u�K�2�:7x�rs=���R���:5��,�w9l O�3�_�ۇ9�>���r��yʟ.���K������&u
=�� �:���[��/����t�˯7_c�����	����4����f�hGx���e��ֱL\Ȅ�������{J����lz���Z�B̕�a\  ڍQqu���ԕ�J���w���*�}i}|�!���AQ �h#��k��dܹ\�?���C��}RC6ދ��|��6l-r��[�N�C�c�e��[q�{>�K�F�>�pa��u�8�E�kD�(�����š'�߄��z���GG�Y���s*�!>C� L4�6�3�5aR�&��)�����9_�z���G��Ntۂ��e/��5D���m3�p�3���Sj�;B �+C�jP�E��k���N��`�/���9��h�Yd��V���~�?���d�RvH�7?R���*X@e���(�.���@��Dԡ�'7s!@u��^�q��f�b�|���f��|��9e�^gh�"����ZemM��f��Z�l�@V
�+���PU��T��8�bߛ��Ɖ(�U4o��|���G�Q[��&(_�p~�2B9�*"Qt�|vc���4���n�,K�m	zMo��yq��2��2X7��[ a�����p5���h1���(K"֭�$+�@'|��YXp�պl�J��R���˔���-Hd��L��$h-�Jө����+j`�y_����#8Pɂ;�-��B�����&�����q�V�%�C�V��֮5BE�at񘐈�M�Z�'���C��l
�-�E���@��&L���;Zi�0n}��C,^k��kEڤK��ǿ�:��ۆ�p�8��QT������ݿ�����M�����L�N�~Y�ݺ�l���e`� q�Ԋ�w4��9��Ρ9�J탅�V���ٚ|W\q���Ɣ3>u���Q����0�Sb��04W�"��h<*�z�<K`�*��-(ƆZD�r�([|s�Zՠ3UQ{R�����3�P�E(�����Q��cӔ^ܿ�<̑գb��Pg7 <o��
4���-��}�[Q��Ϲ��X���5�ov���m�ϢFX��>E#�>0�,fad@��>(�qX�b-���$C�m�eI���ǽhD��l���9r*^	z��y.�;��Ɣ�z�t�8�=��\ JR���Y�s�g��Ľ�3��`�������9:t������#��6�ww���� &�M����3p*N��sD�W��5����E��-�d��w���]땴'̰�2��R�[crE�h-|�KZ�зL	?'�o�xk������A�' jzb
~_M����}y�yXQk���R$�X�p��aVwǀ�7��{B�̱�|���M��L6]�n���4\Lw���7��D �(&��(�w��?7��)��,�9��χN��VІ�o^d�����_���#On�ާ�^�O���}Ptx<U$6(�e����~]�4��F��M���N���8�`B���{_�F\X����p�e
��O�C���-�58'������^�;\H4Ŗ-�J2��'��>�mmS�byp�S�h6�y
_<1:b����B�m��ۤ'�����}o�.xr�?�m�>@g�@E��TU~z��.v�fs�����!t���S�����b�!�׭���'��"�x�������QW4]����8�<��1�x��iPM߱`�W���� A �rۡN�R#���m)Bⷌ�5E2vo��`�_���QoZ�G
J%*���{��8�J���s>�v	��Ńpu�d���:��h�@(*�c��?iE �/��V�U_uw��m]��i��]�e��+4|����^7O���yyO�7Z��̡�H���J�R䶀3ڪH�O�~�M��#-�$k�����I �ĥ�/��a�M�>�$%��M��:�fG���ǭ5J�%1.t��7��I��Tc�E�V.ˢZ������(ї�gJH+^0����/i�h�>�	g�$B��O��!� ��!ۓV�|V�pe��k"Y��7�^f�N�<;��ED=�D���o �n(K	����MH���X��H��	���'����gJN�y���@��[^��4v��,�R�	���=MA�2h}G�E����鵜����b��\[�)��v|ch<�Z��_)�M�2���IUR�ּ� ��6.`L������v!��Z5�J�� =kw��BI�((��v5�l��h@��y<:V�����k�Z>!qlL��z f�}�@NL���C�i�%w�C�%��q����Z���]������B�׫5.�a�]p-)b���"Di�@Nv��L�l�K����ף�$op���Y�nb�_�G�d[�ǝkD+��F>�	M|�Ɲ���d�GOJ�y�C����廆N����͘waw�8��;��Ѓ��"-�N�
�9E�$܉~X~G�U(s�2���?�v��� �S����s��M'w;����U�R���ac?Y>խϾ&���Y�E��輌��ԟ��_���=��ɫ��VsKΘm�I�:�(�Ⱥ6�ksP%D����Ypw�W��"ߥ6al BB��gd�p�%� z���Ռ��P6?$��IO��g6�Έmk�"�fSb�\?V/[�l=t	4�L���*wDs�ڽĤ��-�0F��D0 ��=�� �`�߅s_�Hn:%��j@�h�Ѳ�(�2�3����t��<�Հd�K�Z��o<Ez�d�L�	�V�Ih���y���R��-�cJވ�7+�M��THݜ�� `[}Vv� �1<��4���uMI��KI�Z2����|g�iWXXK̲�m��������R�#���吷ӫY��9��mM��7�h���2u��1�}�2V��j��/,vg~�bB�Vx/� !�����[[%H$&`���=�>[ܠ�[CL���m���]f��n$O���|�{�+d���������	,-S/y�>*nc�0��c�^��,���rs�<F����'wϥ��I�Br���䗟�_~�Թ6��a�zo�:��P����WQ B"H��Y��A�n.�G&x-{�H�upl��l�c9���	,��J�S�Me1]!��I�g��r��r(5�S��?�Hoϒ����d�x9�y����uqW��5�L*$�/���6QY5�洚�+����S��~���w&�=7��P2Ps���QN����N^� ��-^�#�����d�lW��0�2E/Ų���Ē6J���(�YA�Е�.�� r:�e%V1(��UlQ�z?ج��{z0�fg݃���"*cB��]֞]b��r��!DH�sۼ^������6����Lע�~�~�,���E�#�T�U��fٕ66��,.�*�E*w�=(iR���Ӭ�Ox�h:*�h�{�ٖ�R�L��9vlS3S1�a"��R��{���C �+�c!�����{��k�6	��o��"Zl�~ Lc��%���;��7��f}��w�h*����y���%�8@~�4SZi���%4�[�&W�T��M�ܚ����q2�I���4l���t�0�a�rm'.�Z���><6P`u�v�^�H�'/���}m�K� ���x�-�>x'����v��?��}�@Q ?�dRcp���<yg�U�������ŉ�ԪO�|�ȝ Gtҹc><$,+�_��Yn��+��.S���24.]Ct��V$-��������(�Ҷ�t�������0A��sIjWR%����R�<S�k�ٱ+D�/V�q�Q_=�p�Ԑ�҉o��G��֙�3��4Ӈ:.��p�퟾%�;����fJ�.�}Sд��8"����Ps�����Av=���!�6���u� ���~��{����� �9$\b�-
�񺁴�K4:K���W%A	4����BR��T��q�FX>�<-��esV�8�ƬRg�އ���4�	�Q�B�����S{Е-�R4B~Y$�^3�?��0x>XX9 �lk�|�r���;v#���n�;*
U%I����>B<Ýi��J���HIz=�6�`B��G�v��W6�z,zQ���mX�G�u��ƾg��'a+��"�+?�2�ƀ��L5�g�o0��Ad�u(��հrnW%+[�mW']@�m)�[���rց445v�c?����� �m�HWb�t*�+/U�]���1|ʼ��b��9��9��0h�vߎ*( ��o�Ȣ�S��S��jA�y�������&�s��D�OM��}m�����8_���-��<'�����gs��0�͛�|]�9!k`�3=*h裁`�u��[J�����O��t$��´l��1����su�,����_��~:. \NPS'�n�r���ȭ;�2-�)���Q���v��ze����|�KO2@SR�t�t�و�Ω����f�5�$�h��V���(�3� �:s�$�µ^��·0����bc�]��'���]L�%���r�A���Z�ח��.J%�%�٭5����}2�?�V�]x|*I��1��Ia�``��"���̔�1:R;���q���(�1lkڑ���J�M/����I�!�~c���uC�"����>M/ ��X�u�Xt`��,���D�6��7o�x��(�l�Q�'�I�l��
 T+�1㉶��@Û��R��G�/�H�Ȟ���l{%˽�����+�jy[�z@t��\#�k�=#╘��kj��Mu����s�
@��l�L��w�!�(�	������B|�� ����0����%�{K���ա%�=�P�
��Lo V���F���D~�}�$���S߭��c�����,8FF�0k�2�lE㾒x�CN�ä�=A��;���f7�0_������*vW���;��t;_�]M�av��xI�c����T҂��u'<R�B�E��d���U�\�AX���~Ձ��G�����)�OM�S�gCG��G����zbְ�O0e��]����[C��N�2�	0��*�%�S~�V���F�_:��I�[���I�ݩ��,��G�>G��م���Y�Jт�	��q�~��z�Ihi�#p!��a���N!�u[������Ii����1Ȧ��Xݨ��m���ׂ3�z���X W�닪��MPh@`�'M�<G�V�V��/<a���B驍�Җ�� �v��x@脿�r�M�����!�7�e���Cm������XX��ڝ,G��K4k���੄�Ly+�E���ϰYT}�y�����4��$��BLw���]\!/�g�w���;��'����\��0�ݙ1�,W�}w�m��Y����hyH� ��<�^����]��	a:�
g���̢���U�.��U���~�S-ӕ�E^pZ72ʋ��ˍ�z���m�4��|IϘv�gy?�vF=�M�<B�mؓ*raʼ]*�e���}������&@Q�p��L�Mm�r𷲦����s�8W��f������d���|����(�c�bw*-�RC��r=Kfs�v9��S���7��=�M��g-K�9�?�P/v�{��V���):�a�A���/��ؒ%�	b�q�n����uIVF��l�
=��H��&m�$��X��uG�պ.����ؽ� ��VY�vG��7PTJ��#}V��{ӴY���2�(Q)$sQH�)��Z�=����^�.4$^��q�� �C�������Jl��� ���z�:h%�Z4+��Aq�g����M����9I�Y"���2�5���:�\J�7y^gft��rǐM]�U�!o>%n�.�Gݢ׵.3vv`�����{<�_�5^S��M��o����MwL3�]ek����[���l�:4��"�ڝ�Uݿ��r�ӣ*XlL��Lʹ+���W%w����+��9/���0�UXA��.�Uķ.y�"����W��Ay:Hb�|iߢ��˱5��Y�=KxK �w�?�A���ZB��=�G�o�>rCi�T�+M%*�&�>S"��[�n��LDpc?v�߆5���~-�#Y��M�gv�;� ��p�:��S �O:N:�[���܀�d�`�ɓ�p�M���&�G@��?Ȃtb�S^.����&L��s��r-�@4����G�c�M�j�pt\�}��^�u$���V�A"�s���P����l�2�v�R�S�E7��M 8[��<hZ;>2䷜T�K�l3���eo)��/���%'��/���b�(�c@����'��l�)�>��A��?���a�Sةp�e�`����;�H.�/����ȩDf}��G�O<��b��:�T�S�s4�k���]&�$J[����ri���H�K�C�a���,��i(�ǿ�"�/2\>��ʶ;��d�ݭ5�>��U��NW}-h�Z�^��NZ��[��IʎO�� �Mm��x��K��/D�ZU7?OM�ne�ko��Y��'�ݸ��/���+#�Ɓ���q��}E�+g�ȅI.����La4�RY+sX��i>'{�k�ߔ6��l���m����&�߹�lՀ(�|�I� RVC�ȧQ���e E����A���C�E�wh�w,[�WCg���J��`R��}0*���-���G���(����&�pؕK�e�w�g���+ZJ��.W��!d�ـ��%��_�#)|�u'@����mHtT����ۏQ�x?�`�]�6��	K��Á����n`�d��a���b C�M�*���Smݫ�Y�B�Ա�3�Z� ��C�ί1e�Oo���7��/ ,��.� ��ޣ�Y2)qW)�����\���@���Q��T�١�?�0�GY*����lq3�7ͤv��P<��y��k��i_�<�8��f��1�.w;���s2�oPN���Ɣ�e� ��|P�f��DT�@��)��y!�l� b$��o�O��,
�5s�n��g_LeGEc�~=���eҴ�,��,�I�׳N��N��Dp�
���gآt��Db�!�-M����̮�҂CR�yH:�M���9��O�U<[O`��V�5����L砄�mB����mP����)���Z{+��v���$M}�>�VL�w�*ET-���dN3�zYi��W	��b/sQN�#.���]�s�yw%KP��	�G!ь���Cz���,`$��,=)� S$���أMφ���L?z���H'�dZ�;ˎ�-�m��T.>ޏ��}�����L�_e����ג����r������:� $��F���N�5���AL)ZZ&9x��K�y��Iۂ�0���][�4���ևE��;�0ٟw�WD1�� �����ø@7T'=S�n!����� ��4 �=���n�Zr�`EU�����ˑ�{���6��yx�2/�I0M����Ь�?&mR�^�����N�
�"�0��wĠ�"�iyW�Oř�B���cJ��7��d*���������xJ�b��:?*��C�� AB�N�=��b�|�-����+n����yꪁuD���w\�b�Qd�������Pg;B��k�J�\��e���k�9z��ټD������������?qQWl�kz���bվ�h94�n.`�/A�^�_�����شk�J���W@7��0.}���zlP��"Zj�=�!ouMۄ�i��j�$2�#�x�1�ȃ�В]��oH���E�.�g�,_⵼�l.�e;���D��%����W@^�>�XX���ٻ�A⏁s"��ߦ5'������qdi�@_�\K��}������D@Gj��o�I�&�-6�/=W�-P�VA���1�(�Y2�7âG(�{A������a��Q�g�-���Gm�8z<�c������¨���	(le���&}�|�A(B�)$����!�����Sd���ב������Vb�A*���8��%����H����@�!�O�k
�&���Q�ˬz��Œ���[�_���J��3����>L?�=�-i���ݼ
)z�BPkW�O�<u�n)�,4���V?ؕn��ɣ(A��p�ȓ�W���)���z��r�s�&����Y�!l�g;�z��2��~=� ed����`���d����$Ns��aA���c:.�YbY�-	ȌW�)����ܬ]�Us�	�2�|'���,��WЍu1=n��~���-�ۮ�僡�mW�Z�R0��k0&ȹV�p����&�^�SKQ��WG��8����&�>ty���b��'��;НDi�.���4$m��2�l�������^tǄ�y�%�\�p�C�>V���Y�t.}�IЕV��qm��]���>$����Q���2e�oƑa=��<ub�J��^X�P�,���/�ϕ�8M�\�7��B77GÙ��*a�@cB.X�+����=@����[%��tb�ߘ�r�8*(j>���8(&���b��(��+�6��"CP)�
�y
J�oa�X2D�M�^{��F9і4cy��y)(�ˠ�|�|v�d;=�m�!@�Ƴ	S�X%S摘�^0�R��}�)�Y ��*�P�(�$�i�G�����������M�����`8"�ꯍ����^���<�^*���f�`-v��l���������X�7Χ��~�7�yB�=Zw�Ԃ`�_��@5����5�{���}lt�]i���t	?:{���;�ޱ���>!�=�<X���J�iBF�P���%��sQ����b j�exk���g^Y���s�0p�DعN1&V+�G�E����#�^�c��E$Gͻ��6�j�^��]j�� !��NZ��4|̩d��ǳ��cn����.`q���a�U��Q���8���F����(��nA#j+�T��Л}�"l@{��=��mK��q�}Dr�pq�cѹy1��d[�F���$�S�@��w���\x�Y��>��؎?z�����1k�V�e�+�<~�'(��E9uY0�=�2��\aj������y}���r`�֞�,&���/uΥ��7�y�~�.s, A_\u}��]*��G����f^�Lۜ�jzL�N�m�F��;!�/�<~�=|�If��?wX[�N?ں��4=!��Q����r;��,��%��t�t��f�==ݧY^� �|�nc�a�Uת�c����T���5� ��I�%o�Z�sƼIU���wUn;ZS�����(o��xG�Ѭ�5a���8�c3�T���1�>%Y��o�->��e^/>�E_�����HǷ�W=z����jL�G��,�o&�j���R����UJ�SU"Ǝ@(0C���hP�΄g���)��o��Λ[)мt����C���Tz�mþGb5ŝ<�1��>�u��7BQv��
�ۍ��4�(�ܱ���}Axr�}y}��0u�X[�꽘�o�y"�-��n�����Y=��uo�>;�4�_1����+?����V�6�y��HfA�Q�3�U(-W���_X����R�\4����&�R��)��>��i7�x��"�h���Հ�
G3��/wg�������q\��;OL��-=e�'�@��^����eZ��j9�Ԥ���Z��j���Nco�4W��R��)/���9M�}q8eG,��
c$��f˴��DW�Aa�ȥ�P��4�K�l(��ԐQ�;� ��$�dMwzW�	�q���~nK��D?�l�n7�Q|��
�%���h�s���FI8b�*_&�6�1m���@�U�a�7萩6�Hq~�'^^0ΔR�r*���MT7�Ɂ�4oW�;h��L���>�$��Y^�8!N^��� v�â��<����$����z��r :����3�\��v"�eE��s�!����h׀.I(�9�0v#3_�3g�wG�+։�7�8
l���T��W8�vvhL�'>��䉔�ª�|�\�<�ڮ��y��lV�<��):�"��YCI�����H�ʠc͍`�К�j����tL|?�А�����*���U�EaG"[0�+K�w|X�a��Bu%����t�\��X�Otnz+tqzGf�҄�����J��s�1�OPJ��r-jT\»�g���as75��s��-[X��Ξ��֧t N>!�#\_������=JȲ1,�"no�I���:1��?�^�^X�4{��<���u��݆k��\�0Ȃ}֚i�Mf�����Z�4���F�n�H�̈́��J��%�P,�u�7���+��%�(����$�}���A(=1�b����ڛ.1-�Q�l=;p���N-n�$�4<�"¡mnGYC�5�����:�y%C�K�GA�2fK	x���u���-��Q��j2&�Q��ƹ��� k����D}���>��p�C���rʧ�@N��gDa�s�]����̗^�C�����y������g�<g�d�,^�Sh�o�]{<�媏Ie�kXp&�O�p�?B7��Y䳳�z`]�z����k�C	hD�|dX�;�	Dp�*e"L��������UV�dT
�ύ�;$`�{�IL� r��U/�'���~�t�s�I��t���)	�U2��'z��?E�Oʢ��X�u�V��H�$LQL�wg����(�칻��յ��I��}��{*����l)�����r�qH��NWlv�~��g'7��s W�m�&�gef��a�zy>�2r���1＿i�����f��y������8�5fl��Δ���K������� *D�<*�:�>X*�+�k�H