XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D!*��>Sf!��{���#��L @sv�$��s9��of�!���u�0KE� /_n�:rX��`]�LC������tе�j	;��vq�H�~G�E3d3��5��Qvχ}}>T�8�iH�{���`H"�Ug�Ң}mARD�
���jK���P�]kF���<���v��t4o�u���	�� 迂yc(�Vm��Hf�P������5��=�xY�ls��3AJ�ʇ���\�s��J��v����q�=]9��%�ǰ�x�Z.�op�}�mO��a��-w�Թp����Jq'���ƻ>UuMN(�sh^t�������g�e8⡳�f�7�,�$B#g=���R��'�b���q)��XX"
��4��A��dTHM������]m"�C��b_8W��K��m�v���C@�r}�~�}��%=�s����@]0�P\�!�ڊ�s5���e�(�o26���cG�"�'�#Q�;;,ҍ6�:���1h��K����B.�9�h�d�N�nuU3�jL���Ƭi��̻�՝w̑e�:��E�~9G��&��������ʲ{�*p�ַh �6�~{�5c��ϓe�z���/��Ilx`=��l&�Q��I����:� �USK´�A6C�)Y�f�١�C�??ҭ��	֟呶]^U�(i�Z
Nh�%\/h!���Jt�Z���$��[xv�$Ӏ{j�|q�%�Oʷҏ4<�$�FT$��u�m�qb�xQ,�سXlxVHYEB     400     220h�(l+�x��u7D���^��k-�ߨ��b���0�q�aD1C����3ׅߨ�&Z.t���xq�=�-�)-�Tx�$<�h]iH�+�̯�}�30
�iJ��������[�����)������7ik\2׌YV��g)��O�n�|Y�({��i��D�lNo�e����i�uh��]W��3�rXm��"��ws=C8yی�.����N�A|x.�����$I�q-P��{PCO�w��e+��Ϻ��60ͅM����zFK�`-<�H������ëP�w��I��� 7{ٯBzk��#jIe_��D����%F2ء7h��p\�9�F?Z��}~�ML�a�tD��r�#m`��M�"���\��wD�0��Ӥ���M��dì�B���ë���!��# ��t5�Nv�w����J��?񗞀��-����l�"�e�X�A��� �P(JƏ"|\�X�=<4�^1[��Ű:o��(b�g�����(�LbG�:��2'���������1��s�$Ċd��C6*9�Ҟh`��0XlxVHYEB     400      d0��h�b(���ӊU� �t�-8*��{�v�3u�͸��'m�=Yc�O{D�>���
�"Pf0�2	�,��Ѫz�����7�k v��iB������ޏ�,��D�s$tb4(އ���j�3R������^��Q3mF\�򼶄���J��Q�z��6*�;]o��Y�R���bP;}V�+����;S
a$̇�����<�ǆ}XlxVHYEB     400      c0�vH�^�IJɃ+;�����T�%�~x�R芥��\K5Y�� ��} se��4n�ק�ń�&	r�'�%%�ˋ�g
3���U�Tns�+%�P����Y�
�	�l�y��!N�����n2����p���T@����@O�5!x�'\�S +��1��d�Q��X맲b?�1=xE�gt XlxVHYEB     400      c0��~��M�u8Ƃf	�;k���)T ��7��t@5}Js�I��ӎ�`��[r�~Mb�)���D���Mc�E��:�L)-�����m�{�J���y�K���0?Tq ��ɣt6'���B�t=Gn���wg�c�ޱ��1�P�ܼo0G�<\�c�="������/w�Thy\��C��dXo��~
�l�XlxVHYEB     400      d0�0 l��p���v5�`�;�_��)��َ�K7�w�J_�\��'x����h���&��K�`��\]�I��j9�r9��5�Ӯ��nC��sx�Nq+�UD�&!�F�{�k�()��Ӡ�ٙg�Op���p�XϭB�e1祚�d��($|�\�x�P�ӿ��ݏ��Ƌ ƈ  \uՏ*s��l�$�D��`⎽-{�'���s%XlxVHYEB     400      d0&�SΟ.o��kB������>��J
�CTgZB��f;3Eb�b�
qEˍ��n�������c�ؤN�G�aF��'.�.1/�ܥI���0Q�,M�J5���&�����k2�Kmʲ��Q�5=�v���D�Q��*�NU@�]�O����;���E�b��uh�e������Y�������1��1��+'���	��/�|~��1��<��XlxVHYEB     400      d0��P�k�c�9u�wȈ�5�z�]�i���)ő�}�#0�����c��䅢�I�gb"�_9�������B�3؈�����v��ؾ<�>-0dQ���aq�$�LX,e�@���� [W��N��Uw����W!R�]W�p7��nE���cO0�U���ߦ�"��Y�ƍ�:d)�*@�.e �<1H!��xR,����XlxVHYEB     400     170I�e1X�d[� ù��g��_�e�g�
_7|b�r�|��|zѽ��\,����EaĂ�t�<�����nl�ݚL�{��A;�'�[�^��TX£�jk ��g	�l�;(�Ws�>�Kq�8���6� �I����!ú�Z�R�i�˛����=L��L�m�1��v�6
�����uН�Z}h�&t6c�`��0+ٟ�,���Պi�OWm��U�w$�n�<��g[;O�>X-�,+����~�]6.
G��*UaDw>�N�
�2$��L����~H������\��$��K��D�T��T�%���;MTʼO*&���11�	���ڝwp��F"]mއ`!D�&���-W�.��XlxVHYEB     400     140�Ѱ9��\c7�L��
7�P�����������a������c�
��q�������@פj[ɕ��&�:�-l8��vK�����Ԁ�H���Ad��9W��`���%ӹ��-B8;UD�{�E|�W��r%V��_�t5Ll���RibsЗB�T1K�iĊ�SF��չK��y0�*gm���ӑ����y�k�}�$�d%޽x��u��->��Xt��Ն^8�}��B��Ϫ�4T�hAb%^7s�D}�拾\���pGY� cW���p�J�{_�Jp}����i��@�!�c6J,�8�q��B
����XlxVHYEB     400      f00%�&������a_�e|�s�l�ܱr� ����(�"��C�1~J촶0"'�������k_�4ȣ�/�� Ƨ�%)�&5�o����V�_�	3����ԾV!��sȧY���;��>d�> X�7�1�Q.t���5Mu�̙��NT$�s��	�fڝȐ.7���$KP�{}Ր(,[�����l�!�T��b+�`m��[�R1�q���_����x\��՗�N6f^g=���<2XlxVHYEB     400     100&#��_8�tj|� ��l�=�ߒ�-���~��7N��f�������E&z��o�D>��૷�nנ��?�pI�{�\H 3[�Q�)Cn�q���̷���j�Z��"�Rd���GBv������۬_uQP$)�	aŐ,f�o�x������1I��hǠ"���xX`i���8�΢�n>�a/0Gnܫ�2^���Ԥ/P�<�����>;��U�v׬�묽�WZ)��!�
8d���C8qqG[�B��ގ�XlxVHYEB     400     110R��㳩oIl�N���Jw���g�>e��?P����p����v�� ��-���t�ɹB�7q��ZE�QT/_��%��t@P�|���#�C+��_�uR�%���'��Wj�v1_�W��l:�Yƍ��s���t��ٌ
�>�[��@2^�-i�T��������D��VE�/վ	̪?OP�dw���j)./�z�E���./��N��W���^��n��t�����$�2��{C	��hf�6���E�v��I�ޣXlxVHYEB     400     110���k�e�g��f��a���u�/�n����j�?t9��� f.�oZ �.�%}��`F��@-���L@yK��>�Ӑ������E6d���PnA�0�d� ]}��]4N2���Hd.�N��X7��6�EDԞ	���̭lmY�/�� �����j��ua��+EJ�t���p�\50y�~RD6�CzX�^��T��vO,�������3�cRʯ�B�g+5XgS�G�6��q�ⶮ�=
O�>}���c�k�ʬ���1߹֍=(�XlxVHYEB     400     130�_�bQ�+�І����::��*H݆�j~�W+S�l,�QzWuډ�H���w�n�=���a����#�S�$?�ڀc8��ު]m�'+)\�p��C4��ՋG��M��m�@�����@S'\j���My��n�p�mEz%2�X;�Q��	:�b�D�	Ğ��X��4δ���Pk�=�Yx�N������揁6ܐ0�?�?d��G1���b�*��pz�PB�F��>"��W���6&����3��ԥ���N���$Ԗ	��n��&��h��"�<�e�XlxVHYEB     400     100�vg-ڀ���+{�$+�pY�<��oH��N��M�	���q��=UF�hi_���6��/{J���y��z(լ~���μ�N<����"�K�t��C;���W���[7�ƣ�n+r����Փ��x��sQ(��5�[�_�\I�l
�[���fe�p���_��<�I��{�b��nG����Z�g5UIe�,փ�i�����n�}��6�A��K����K���y�/�I@U�U���͵lD`Z")2L��`�\XlxVHYEB     400     100����˻gp.���*������xT~������3�@YU����ps�x4�8	=��6�,h�6�����#�����\��r�A��. =�7�7��Ͼ����q�.�x&��MO ���H�VcqI�n�7�<ty^3�L#���|��?�d:R봧�Z!���a�T\Q���h�GlV[}h��g�~��B}��0��Ƕ� �T.c�/��^�zgEԑ˄�N����
զ���|%q������Ԭ�0�h�>�9�XlxVHYEB     400     100�_?�����{�����Uq9��W�QD�q�4)>@����:	�f�D�����D��b��:)�ܺ����U+R�@z��$�����{�8���q�y@�!Q��P_������CH���w�.��u8&A��R����L���k�>b.f�3�r���@u��>un�xt���}A���'��׋33���T�E��o��K�L�b�%,�~�!s�s'��?d�K����f��ݡ�zCb%����FXlxVHYEB     400     100�6����n�Vi���Ex���ֻ�e|�G;K��ߢ�L<0�~7<-�%���䈌n֒Ͱ�N�j�\b�E:�4Y$��놌>4i[&�}���Cg��^&�]w*�J�|��d~�<������\j�M`�d��K�,U^�"5�R����,��o�Э/6E� �}�-�bCQ7(�)��zq�R)LT��m��?�C �V��z��G��:��B�n��w��#�[��ŕօ�6��������wXlxVHYEB     400     1007�*��q�|C��yf�D��:��_Zj�#} \e&����-S�R m�}$��O��+��%�O�kI<��Q�<dC�����g�b�=+5{�+{LHO��aF1�d�}����٘Z��+O��J&ԛm�6N��� [���Q����#� ��K��.�h��_ꚨ�j���~��Lx2�t|������|f���Ƈ&1 m����Pk��<���[s�����}��NUV��&7�%�#o�G>�'\̤XlxVHYEB     400     100���
UZ�,0�9O�ȣ��tYK��שm�{b��?0����(l�b3s��~)�¿�>ؽ	P'b���M�kb�5����Y�ҲY]C�R���o����@���C��@9u_iM`eA.�<��n�#z�Ɍ`��+�yҖ�po�\��:������e�Vt���3�z��!a�D� ��CA��K������d���h�y �{�vR��X�8^P
d��g� �f1`��
��{��:fiE�|�v�
a'�XlxVHYEB     400     100��v4��Hr�0�,��6v��	�j���(�p+s���b���O���2�2[f�= G�CX42�F�r0��l�=Ut0�n���v�j�8�tw�s8�B&N���"��G�}b�%������fj�b��D�*솅���Z��/{��=�1Rˬ�M]Qs $eh���� N���5���jۖ��^�A�M��	~��^�[�\���V0�(G �'n�
7�R����̺0HE�f�a�+x1�lG��W��XlxVHYEB     400     100Ϋ7T��qtQk))��bS�����%��1��7Vu��V��Rl��X����y��'��T�\��qT����|T�2�UjD���h��;�m�F�'�Ƅzu~�?T�Z�z��������8�L��Q�t�]>X�b���c5b�vG�Z����dm�������,�I�_�6c��ϳ��~�Ba^nY�y�qBZ{Ү>�A*�s�w���T�gc�,��~Xe3�k�,괻���w�2�M6�.���T��3��J�XlxVHYEB     400     100,�ǭ7���P_�\->��<�h]&�o~Y��`�o�9q[I����<�>�o�;Y"�DHo��
D��Sy�+Qq�%�b&>�+|oI�iH�e,�Ùr�20���������+��23���)o(�5��l,)�׾�����*.%�$Ӡ�ɽ��2����J�4d/�_>����ًĽJ��J9�e�֮;�8��`n�2����|����i]˒H��ū[�[�2Kab;jw�G��z�!Nm����;Wh�PXlxVHYEB     400     100�W�UO7��1b�v�Ek[��#��m��_r�wѱ�|�:43Ǖ�-�c#f��6Fi-.�xz����M�`!��������#�M�IR��1F\�8i��� �^B,��$�Y4����آ����<�ӋO��}�b��]^�����?�cK!��:�Yׅc@���z�Ll� ����i�`A��?��e�vRD|���x?�|�;f#ۖ�Y2Ĩ�§=.���x���*Q�9�as=��xj���"-��`즳_Wu��ʈXlxVHYEB     400     100{�)��o'�5�k?�d���ځ��̚(*Б`�������t&��@���@��_@�:�ũt��q�qe0M�bz1SN�8����t��Kۀ��DOM8kTQ�Y���0�+�����:V�m��:�������i�(�7�Ae~�O=Hs����-�^qN�`���V��q��4L�C%U
|����@C_ڙ�k�HrڭQ2Pu�SQ���q�z�ܲ[<Z�^��E-�M� �ڜ��Le��_���]��0�M��H�XlxVHYEB     400     100-�ޥ�lzDrk>$U>K�B���I�-+$���|_,�	�3UU��0��ή��Nn5�5%A��
�J967djz�,;b8�2������e��z��d���8�nn.!_���C�����)�L�ϣ�2��V���q}�Y� �<,���\�ݑƫ��ȅ�\�9�-�2�)��L��"/�ېѕ����*=3Dײָ廃�r��]�����ʭ�
�:����8|��������[�?.Oz��'atXlxVHYEB     400     100~X ��gi��"G�>�)�`.���b��?AbE�:���0zu��7�����}��6�0�B�w����7S�t}�0F	�s�%� 0��/�2蒛T��l���q��Ν J��U{� �FJ�����1�X���Y	�c?3�ĭ��:2���t��T�SYu�B@e���|om�Ȟ��,�9^��+&
� E^��s�i��Om��$�޼HR�/�4�k�~�΀	�E�8N��A¬��[�]��z��&4b����XlxVHYEB     400     100
,\h���d1y���������Ģ��D�}�����I���k#�< A+�,1���t;��1S����CD'��H|5�u��@�_�&Bz)����a�Q���̌�h>��SyG�E����v�~R!j���ڟ�R�-��P��-H�Փ��{,A����$T�IT���E1���zQ���8���@��)�BR��k�Ҳ:Zo|�S�{u���?q���L=o��Hv�4Dt��g�
ؒ�Dh<g���XlxVHYEB     400     100�?��f���%� <�86�?Ć�g�Q����[ ���ѳ϶i���V8+�g�M��Om�z]�fr�;S��X�Hn�I�5T���/���i.wKOo����K+;
��Ǳ��~+oV�h\,?*�Z���-Ml<�QЁ	ng��<������q�J\��ɐ&�*���;.�^J'��EQ���S�4��ժCu��=|��%�O��Cn�������0�[|�1��v������!������(�
W�C/O�	2
6�XlxVHYEB     400     170�M�(K����-iժX��dH��6y'Ȗ��)��g��]
]k N2W���j�hN���V��JU�v#"�{�+��<Zt��S�YsC�V�w|6I�pz��QRW��b��>kJ�M���m�Q|�2�c�i+C�F��D��f9�w�}�?X¶K�ap\�F�VY���K�\.W� ^��?�J-�Nn���C���AvZ�?*�%��OTh;oS�E�XUU�s�Gw�R���'W�x<�`���f��\_�5lb?���H�+]�怠zq�>�#|F��l7ٛ�g�Va�\� �D�E4��ǔ�ͭm-!9!�`Ų+��2)���x��'�W �)��5V����'�ʷw���k�"��U�#?�-SXlxVHYEB     400     100*�̟�[7��1�����І��E���[���iz�]�+�f��3��������M}�Y�!�`��<_��|=Aj��d�w
� ��;�'�s�mk&2l?Dͺ2� '��o{�.��cU5�!�8�������t�av8��̈~�X�kҐ-�Amb
�an�*G7?�Gu�2:źT^!�J��P!).jȋ>(��0��
�jQ���4�b����(���-�0�)Ԛ�����	���8�)O���p*��u%ۘXlxVHYEB     400      c0 �(og�*�����|)}ćC�Ɲd�))�a�,�O�>�T��K�������.��&�U4��-ᛐ���_*�vȲ���0 aV�v\��\��^T�E����P�Tb�Š<�B�q���f�y�]���9=#��%�S��<�����k$9��s	�Ӏ�����^�GD/����ca���l�8��b�XlxVHYEB     400      b04���mc ?�2u襟++v@G�].��$tr��:�ݙ��G�H�ѕHy�n8�F�7���Wa>2h�@.�l��b��t�����Rܐb���������S�d�,�=�bQ�ݤ�n������A�P��TMS
-��si��y�eoEF��dg�f�P��B8���ԑpr��XlxVHYEB     400      90Y~WJ rʹ����f&cݱ��q��ǧ�:�����6�Y�EN7_���f�}�pM�wE[�6�}qJd�_+ ��`�q *��6F��`�<��j���
е�HF��r:�:�Ə9��_��/���~Ųk!0��U�/��t���,�����XlxVHYEB     400      90�	�Vd���8�!9����a> o~��:V��(����u>f�?ۦ��)G�^Fgy��\̢�_���Ʉ���|F� )���Lf��v����p5�]_"���({k�u���-�����I�+h��{M�Q�h*m�'�!XlxVHYEB     400      90�G�#�1f�n�59��X�GU��\+�F���6"K�:{�O7��o���/�\�0t4���U���"B3
�iH��I^c�@��� Y�'��7=d�SK�c���2���A;nm� kӧO�j�a�n��,��o%�f%u�4X�XlxVHYEB     400      90�D�[����m\+@�>��E�j��������1��4��ԁF���jו궜�u+oU���G6���Ӹ;�V�c-LI��S�Km���m)0̗�2��z�E �~�D=-z`
���.���p8W�P����ſ��Y/B7E
A,�&�RXlxVHYEB     400      90����RFM�V4����N� Pzm���q��aK��	��_��+4j�^|��&��G�@+V��^�+��1�K�=��%����M�R� R�,�}40�p��g��x�ü$�Ge�k�ȅ��̝�g��H�5t yx���t��/	�XlxVHYEB     400      d0Gj�����UE�~5�܅����H�V���J��g���u�3�� ��~�]d���.��æA�&� <R��3�{+�1��1���
��M]nz�Y/�4����An3z�����xɣ?��V/�w��M����$9��2c]v6�G^Q�yj;�m� �l[#A*� FI�|.�<$�!��X�*	n�CW`�	����pYF��r�XlxVHYEB     400      e0}=��뀽��H2G&Y���w�vc� _f�H��"����u�|na-���`�:8W�~�
�AML�d2(X��D���֏��������X!�=�!D�>�{��usƣM���?@��7پ�)��i���rc��-�7��o�Y����k>�	!�,�v��տ��Q�1����������w��O�(�#�3U�l2X�ə�7 D�\Vz0r;��4�?��oXlxVHYEB     400     100�o�Z�I Ll疐)ϒ\1˿���F��@��kkr���Φ�O��?۝�g��$ٹVgSԹ*�b�${;�����r`,4w~�(k@B)<~��������L�cMu.�Aw0�E݄����V�kD/^�T���:PS��o�Cүck[H��G,�p��+1�u��di�YS9HgC�KxՀ3�h�we�Vn���qs'�����%7�B�KPaz�zi��"#�z�f��ʰ#�B���r\n,:�B(����� v��Ou�XlxVHYEB     400     160��\U��Z�W�;�F�z����\��w�HL���a����0#3w?�|a�6�	�x���#X9{�AR~;�(��<���Z��H�@��?��1���v���\#�l�:g�D��ht2;�`<��~�z7��H�_;��K�QpqB��r�o�e��D���1s�ê;~{���!��W�\�P���o�W�P�;(�+�U4%�|RK1���,	ݧ��,�'51ѣ<��&	¨B�����(_�tx�qi�ڥ�&��@V"!��[���;�� #��.e|���{�f$lfw��v*�'%<ǟ红����\}S��:{D{֢i�P��W�vpC�3y+,'�
uۈb>&jXlxVHYEB     400     160A��.�~ =����1 �c�p�^������iՇH��\-�^õ�� |�a<'�o��d�lJ��>���5��`]�g)�6�6��C�<$Y2X��)�������Ȍ�ۮ][�G��r���m�N)��|Mt���7�l.�b�Ci�I�qf�C�w�����x/�9��d���9n�H��N{�>�v��y��0�l���]�C6�;{}�O�k<��M;1��]rsޏ�h^	������HP�))V)`��
�Ԙ/wGAK�� OP3��c�/�i/_��܁����X��zb�L%]�e\>�ٿ��,̓�����6Ub�7N��$䷪^_A�ޜ���-�Q��XlxVHYEB     400     140˟���ޭ�X"�NgЎ4K�]�]��ܵY*؋��j�@#3넲#��������ä�}��n.O�Ƣ�]�����N��^)�"�+��ea�+�k@� (kJ˯�Q�U��$n�1���MX-<I�E�-�� *�騌���P�̺�����[ ��b�fֹ�z�z���)�&0��R�V���Tq���{y��7��t!T�Y�C���<w{]|�k�����H���|,�����s�����"�|�_�����)�0�V>��p%�S;��,Q$�ֈ��&L-O�ZoKx��x�1��˯�]g��HA9�XlxVHYEB     400     170%tv���r'�[N��_v��B�z���P
�������Ե�'K�௳�����o�(s��W���ֱd�Ze!���6Ht�����~ �1'2fm*�~1�lv�!���o�~����y؉Mn��a�����ӱV��Fm�X�f;�)]�n�[�'�7*�(���yI��w�H1M�!wΌ�*U�em��6�j�}����g=�$�f ��q��<I�`.&:3����0�1�P�����l����N���tL>Xb����C	�ȡ��-7J�B5�f=)�/�J��W�94]b��B�������j�h�c����&w������V8�c~#bܧ�rl|�'$J��Z�K�;`��G���XlxVHYEB     400     150<�ˊR��.�2�v���M�h�+�X[!�xB����q�)�+d@Z0��m�:�cDu�����M�~r=� �;[��ן8\�$�Q��纰����=E-B����D��3�@�N�B"�У��7e�oc���igK�]7UU	����"q^�6���PD�܊���ųg;�\�p�Ǆ}%��k�EU��}�� +eI���H������zUSWMxZ��#%��	����N�
��">Kơ�c��si��\�p�z׭�h�.��fq)��m9�~ڣ��Χ]��h	�k{]���'uVG�Pk��(	����	��7Kѡ�ؑ�,u:�L�uTsXlxVHYEB     400     190�-g ��%H�WCQ��h�i�U�T�R��o�g�]�5�I�2��#�VL�]��z4dfL���ޑ_/��յH'l1+FYb�Bn%�3�.J;J��놛U����O*����"�i���M▴ec�0l���ӑA�����e��p�a}B뛨:@CA��}�$7��Yb7��5l*����.ɢ��g�!Zއ�D�-��#I�+���p��*�7:H��H���-�~3��l�i}��Z���xRk�68���4���vFv���X�G�.�)������P���q����)���3�I�Uo�|��j������D��,i�B|7ǊyMK��k]拄V�x�e+�e%l�@��eK4����C/��@��^�ؾ��Ӣ�i,2�1����XlxVHYEB     400     150���������9a�n&���]z3죨ta@���&޶��a��������*��+A9d*�]�>�.�����Bdܣ�0�w(�@��<宯�1�K_c�$��0���ޕ�(���+_:;пB��d�K`"�O�7bP��DPV9�D�P\mw�Ρ'��K9�Qd�&�=LpM��С�<�W�v���[����f�f���1�(���Q�g�}��L%�\"�G�;,�_���.a�G��{��\��O$mWtC��c[�1�{@c���;�����e��(���vpp�쟰��a����Dc>�,�ѣ^Z(\3��%�xE�:��lj(�����k�XlxVHYEB     400     100|�|I��Wn�sF8|�����Z��M��lR�̋�3���/�Q�h��t������t�ĩM�H(v��y�]7�"������Kq�Y�� Ӎ�T�i 	9FDr���>I��+����U��n��*Bh,V�pN��d�4���� Mf����Q����2���8��\�P���ق:\����ٸ$��jxa�x}��U��F�F�r���[x��_V���,��E�q���I���B�9I4XlxVHYEB     400     190�e_^8�Q���#���@pUl���m�AkM��YOt �I��Dx�	� �H��J**��v�DE�aÀ,]�������	Υࠕ������'y�DC>'��s�=$o�=T���N��d�
>?���bRN���������h�_4T�+��?J �+ޫlIE�z	�h�N/��j⪞�S;�HRM��VQ�%�u�Q��`]�(*�_�4��I�S+\��#6^�������b�
mݶz�Y,�m2`*�?Q�b��9�<��f;`�-%�l&�:�$~�U�R�W���u�.����b��l"��L�g$[�����.�ͥ:�;�^~��Ա����1���O����j�x� �T-0�	�)���$jj��t�V BoQ�xݸB XlxVHYEB     400     140�9��bI���ʁ�z�s9a=�{����\$���T'��T�`�g�	.�~j��]6�,⼨`l��e�5���
�7cyD&M�be�	�����1����3BE;��@�����qU�:��c$�[�0`���������3�M��#��/�wf��%ky^�e�'4<�ņ��V�h�x��u��C� �?�#��>~�Y��#�)�3��*f��?�%FLo��K�Z�wa,���{=�V����%t�c�/�/Itu�++��))� �ƥ�HTZ��ᅴ�oX��f��A�+������T���'�A��u'b�NXlxVHYEB     400     150x�6�A�m�1�q]�XM��q�&���a�'�����?�!�`ԝ?�2�rPHK«cu����I@R~�'�1�?�5zFӪoL$���o�
�Ap��vؐ�߀��8r�gM�o.L�$iG��~��G~���Y�b�[bs���Yό~��S^��5��ӭ �,��XS#Vd9�԰4~켃'PĜc׾|D���1����^��Z� FX��X.��g������W�5����U8T���U��C:��z�b@#av�zvMa�����=��;Ն��!�w��2�_3��FX/�B��Q�1�<qw��;�g��,��&���e�
������XlxVHYEB     400     110�i�|�QgW6��۴x�hs�z����AQ��� �*aچ�[�^%9� ty�O��aa"�OXA��j˹{\64YV?cM;�hVu���	n}�Y�*g8O���ePx�4��07' �/��]�cU̔�IpSzv���_�F��t�u�t�m'z���K���u:a������K�rܠ$I����=����J,�lӜt����P�]u���ϧ(q��s[ЀQfqm�[Sp}E�d����i���\T����#����U��-�,�g�XlxVHYEB     400     160ӹ��t��PÑmYЌ���%��'����uH��ib-l8���R4O��v��q�����qD@�I$��r>�*�E�A݆S�4�=qy�\�c��{������%��lY���<d�>n��T�&=���K�?+an!��T��
�{��A�ž=�.���N	/�����u�����%��z��f]�{p>Q���O��L�_Ň�Z��������(0Ą(V��l
��AH��"{�~��f��Z��hU'$����#��� �*4+�	tW�_�Yn�M$��	��ȍt~���>ː�^Ӄ�9-�E�#I�t��	VoB��;T3p;2V���'��O� �2B(=���XlxVHYEB     400     160@H���#�����5�+j��h?�Qv��h��\v�!z#j�'!�X,G:~r7����dֵK�����Y�|���@���b˗-�g���b'1tڶ#g���P@�	�6B�⻢��$C=n��s�'�0:x4�&����^���=&Y�� �{�Z����ߨV~����K��T��sgG��h��9�@9�-_.z�Lu�	R
�	��'�x+�%d���#4�9��GpI����ӾW+gb����I�l�MG�i$�a�+�Gy���"ث�y�g�lO��������2y��K�L��#� ��.��c�2�j�Xj�������[p�Ј����Zթ���XlxVHYEB     400     150c�!bU��1��z~�ȇ_OV�[BtE��*i.U�g������(�4���t�u�J�i���s\�ۦ���=�&Lr�~�ʾ��9+���;���!�<J���O��%X��)DU�OC����g����:��4j���j��5�T�B��������y����X�/%�� �δ��^�փQ��۬Sj*�*/0��'��H��G1ٜ]��5E�\�P�����8��*��>�X�A�C�/��� m�
=�5�b��WwPa7�,�YF��q��d�۠jz�Kxd(6~�V������;��?I�� +�V/��1yl�@O�^rL�U���XlxVHYEB     400     150v<�L�o�B���� `!P 6�)1Nq���]�4�m	[�;�Z8�v�X��k7�sY>��_��M`��ǲ���$Tn��{/4��J`�ʛ���$���RI��ѭKS���K5�Z�kG��FU�,�r�������D˝�%���Beث��..GX�5L���-��;Vڡ��&�3�#!�H��Iϳ2�����*/s&vy6 Bk/V�~�fx����Y��CA	��_��x)��:Hl=����AJ`Lx6q#��I���~r�TF�P�� ��t��tRAZ��QJ�_g�kO�;$�Y��%Ǣ���.v�}�|Ll��=w5F|U����F>�RXlxVHYEB     400      d0�d���k5x ��:w��ǎ���/�kݿ�;���#�ti�>N0��CU�ͳ�fO�h6}�C�*_ć� )�����!�moA���G]\�����x!T����:�W!J�蠰��c�V��<5ʷ��&�ڔ"�9Y�%�o8k��d�Ӕ��F���綳�m*���	#�4 S���7��m��瑎��so��}Ǯ��XlxVHYEB     400      c0Y뵏��7�z��N\KDiv>l�M�
�	�N�zQ��y��D%¥..��N^{Y�~�:xvN�Th�J�	��a��W4��tߺh�K���3��Dy`;�~u��H 0{Jv�,QAl��g�&Q�K����o�tp�K���R��
'~�.�;%r��v8F�pҌ�;d*.VpL��������snh����[XlxVHYEB     400      c0n��B��!3?��&��j(.�x�`L��U���;�й�QFG52.^P�ȝ�����<L�Q���M�u����x6��
��fLV�����p5VF��r
7��xG�1��:8�'�f_��S|^�(�ς@�i��n�
��@5�R�ޜE͎��|�ކ
Q��̀z�x�˞�^��4��\��eXlxVHYEB     400      c0���@ٻcCǏ�c��q�S���bny�vǵ�S���G�N��Q�)�SfU�Hpy&c�"�Yw���x1��
�����,���J�"IϞB`Jk������=E{V�yQ(��W�����_��M;]Ͷ�e�!y�R�qd�)��r"nA��t6�+j ��l�Ϧ�����jT��[|�K�����&XlxVHYEB     400     100b�.cX�O�9Mt&b0i)ڤ���V#��Qi74�I�)fH�#'*�g,�l:�0���&C�zB-2�mΦ��L��/F���3��*�
�5���=��Su�"`�D$��&s��7��bT�l��n~�W�j3;c.H���v�Y0�`U���YJ	�T7���l��].�w_K��Q֑�����>(>`�T�8���Nd��^�5������C�V����(9&G���/�Q�j7�=ժYj�7!�L���XlxVHYEB     400      f0��V�.�K \��-�s�8J,,�>�5V�u�v9�T�T�����L��O���M�q(��E�`:wW�@��&,��V���}��Ә�1�����$u�/^.'��C�Ƹ��+��)��Ű�TlS������i���&s�[Zη��<H�2����N�*�u��N�>�E1�U1�/v���bϐ�D)��Cn�����x:��@����14��T�|:��2>Cw�ѿMm,y�z�XlxVHYEB     400      f0��:�ͮǲ9J%
*F��͝��̪���D����������\���~��)e��晢�h\��j�I7���ڙf��Jz�?@({�8Iw�,q%OZ�%�c�� #�lHu߹��sD�E�6A�|3�(�Z܄9@&[��Q���Њs����M��"�f�i`�cd'����V�X�;?'%P;�j�m���I��-&�l��͢�,b/r���m:g.ٱ��~�\.�dK6��)XlxVHYEB     400      f0wю�᷺��;�^|�y�P�:e��Fn�	nA�W/�؈{�"������,➪��T�cB4��[�����d��N��>̛�hTy�S�T����ǠW�yڄ�1vU�}��-$��k�>h�t@�V��M���z&]����UC��v��LBؘ^�ۙ��e�+�B��s�r�w9��/�8�&�W����3	�cE0��?7�����q��_Y��T�G�G��(H�ɝ��뫃�ҨXlxVHYEB     400      f0����NR�n/y���hg��P���(��^��q.�ޣ ��#�3g���n� P�'�׸�ȷ��͞���eD�g�}���m1����qY���,n�����XG�%q}@�P��k0��l�?��QȂ��� T����K��� n9�#�cCyI~���I�5��t�CƮȤ�۔e5x���
u:v�z%�h<AX��By����җ�V�����;��f����g��(��
=���XlxVHYEB     400      f0T
m�묄�#J�6�Hb�e�i0(�K.�SLe�Qdv��ݱ�~���D�(ϕ�楖���Q�.��`�.;�<��@<�h��rʸ�[I�YCG�	�@*3"%�����_�n�?��I���(}�8�Z��`�gV��O�C��.j��k�JK��%�Y�jg�}�gkS��!^�	T����� uq/����FEA�Z�����U4��Q�W26=;�_�9(6�^�S~5ዖ�>����Y��XlxVHYEB     400      e0��ı�0��LsI����F��{�h�|������ Z��"�f&?�XQ��Cb\����f����� �pɭ�x�}��~kz�ea�[�q��l����8���v��7��,����p�u;��Wap��?�n�Fbz�k�uF��򞆟.�ql���e	፜K⸁�2�lH�K�%�����C�w9J����pf��Q�WMo���� �`��v:\ ���T�$&��XlxVHYEB     400      f06���n}�<��]������b�HE�o����oÐ�3��p����*ELP2� }��ZԻܫ�UK+,.<3��zjP�p?0a�H��޿Ujd|�v'���kQ���~�}���S����9��;�8-�4_�&N�M�-�?��L��h��]�x�&7�7��3���&�mɣmk�ߤ�3{�h%l�Th����bGvf��C7��d����r8$���ϙ���]m�(C������XlxVHYEB     400     150R)�]ʽp��� ӕ�Q
=���|�1Q���T2H7l�Z��~%Hg��;���f���\�%�iud9��ک
*�$8�[�b"�>Yqȣ��>C���#T{Bf�c�(���1�<�U9h�HjS!i�3p����o�Р��?�R�H����x.��Τ@�J��'al㗎N�����G+_)�Y��<S*��#:���ׯ6rn�y������PRg4���ōokG�Q6�O,�n�{h�]��KTq	�($[gc�:t���}&�F�o�t&��=.�j��&�UX5D�gw?q��ayeJ�����W��ŏI��������XlxVHYEB     400     1a0t�lg]����ˇ!��A�w�ꝏ}�;�B�dS/�S���-~Q,�+\�g��}�(�ip�Rʔ㍌��!��6��|�4��������Է{�2Cv��k,,�Ғ(�?8`������d����
e�2��s���W�L��V��m�ٔC;G�#�3m��fw1lUaB��(x�Y�o0P�Z����4�����N��� M�5�@���q�81������e����S���W��5���g;��ç5��D%��bA�B$�lD�&بA� �5���p(^!���?\5u?��BR���� �r�p�#�о��V�2����V���H��s��^`jz8=��>�I�30h#DMNec�+�4�+�����hŻ)y���{G]gb�D���
��ڡ��|�[�y��������XlxVHYEB     400     150:�j(b��n@��,�~���<U,�����;~���W��JǗd��q�9��i�_�.L}��oP �^�%b[�1���t��weP�sb�e�XXW���Z��amE�N�|8$�-�cC�䩙R�~oa	M%<C���'o᳂+L��~�]��8����Il����X����me��p~ߘ�����{o�'#+���x��\vl:(��6Oey�TJW C��wy(D�!$�M��<\�ᵕ@�'`	sĞ�>#�V�oW���Ġ���"#E/�r�σ��{�H�5'ŲBG�p��C��mI�����~�\��T@e��8�s�Ӟ����}�
i��XlxVHYEB     227      f0k�}A��hB��0�x�7�q@}\a'���CSh����r�or��P�1ż]��Lgm�%	f�I���-��J���l�Uw���'���=4�$�_���AW��9F�ه��E1H�tlQc���"��[��8j�>S����]��v4���B�g>^��>�,��il��Iq߼�,*""v8�܁�4�y�Վ�
k�[����֠��zCm�F�;ia/�;C��{2:C
f���p:K�Ts8