XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ľ��;8��7�,�[�����N{pfY��Gȴ(#M.���)���ė��	����e�K�&`;W²����F�2�)C��AcSFѧ�Xn�@�{�C�lrִ��]��ې�~�y���J��5J@�e/lWս�{��gy��G�ސ2}�����
o6	%�t� ݾ�k�(�����&4��{@Le�bTD�q��K�9�e� |/�r�<[��_�{>�J��λ�$��vZ�Xͨ��-F�F��-�����x���@��xb'`,��:�hj�$#y��Ji�YE}Y�X~���t��)s9cD�9Kӣ0�ho�/��.(3TV���&�&0�奂e��U���$�o�d۽���M��������ݫ3_�Et�nY��g�2�B�=��q��S+g�M�DB��ԇ��_�)�_���6}�7l�Hd����>B�$֎ժx:�M���Tc!��Q�>�m��Լ/PJh���5_�-���Wtj%�3���{�������">=����&^^�1���㾆"��]��籤r��m���d�h�f[�b���e&M?�!>G��,��A�0�"B7{S������,��G��^�^s�E�ƥ>�qb���&��*{�	�ׇL,~��)\���1��8w�7()��1h��Ô�P���\��~�ж�ͦ��Vc�Z�'"�3��b�6��T������+�ˈ�t�����	-um��;��� S�qŚ�]����\��ЙK�ƥ��~�g�ecs+�XlxVHYEB     400     1b0�%������,K7������k�=Bf�����Vn�OkEނ�y
I��4�������`��V��y'p��zm�����C�D�ɧoԌ��*
�}��UVJ ��G������oV�RƦ��>�?!��aΕ G�֍�PE`�����Q���T��Ƭ�3���ZM��(����0CKJ��p]I]�y�>�� �S�@	�oDpq�'txwN�*���)�����>r�\�٭P�.���j�q4�ɡ��D��%(�����1J6�H��=���P��եw�I��A�[y?��������7�
׮,$ ���ˮ�\��C�w�_D��>�P�0֙���M���<��o�ky|?*OQ�����#IB��f3��f�u�Y�<�ׅ����2�M���%5�uU��_���xr!�XlxVHYEB     400     1b0�����`b����JE�>:]��i��ʩ ��fR�j"^�·�C�����b٪[9Ӫ��"�G8	�ϩ����Pǥ����7k^
-��*��n���6�6�X�=Z�
E��Pq	+��Ip1�|8���'�e�)h��@�%uЕ����k+(�v[�G���FH��:�5��E��'���@��X!�W`�W)3�VGzs5P����QN�Q��U�~g�q�V4��.��I�m�6�?34�;V$|JH���4�:���0�uJ?F,X]mXS���C�c�@'l���:F��	�;���[���>F#����4l����$nPYj%<.�h��ף<�qk*��:�ݒ��~s�)�!M�r:;_��-��@E�އ~P� �n/��-%d�'�d�	_tnX��]`�śm�C�XlxVHYEB     400     130yW����,f8�5���}�
��1�Z`�r)�����S����b%��~��!ADMG����l���A+{m'M?@6~�i��1l7�S��2��AE�6��AֱbO-G:���Q�V��&ߛ{=N7r�[�q��kЖ��6�û�!�3-����g1|Ya
R᛹�aݕ�-�Gz���0ι�� ]M��FZ���N�2w��$�ۚ%!{?��3��08+�E�Vp�s=������hh��&L�Ө�v���-�MM���P8��J�"�D 9� 5;����	�ͅp�����cc�J�K��JXlxVHYEB     400     190��9��
��h/����$(�_93��j�'j�q�)��H�X���(��p�������#�w���mv�X
z�|��:�Y���G���d����sI��f*����N���)�)���AԜ섙��[�$�KA�Dw�l�Vi7�C�(}H��L_dS��+�R3�3cM1	(�;h�/e����
B�����e��%��l4�cII��ywhR�t���Y�����z�ߊzñ辍�� ��re�Y�P�{�Ǟ���Y�x��r�J`���耸Sc6A�>�X�c��s��p�Z���(>�&$e���m�kM�@����@y��0��iJ�<�Y'����d�|�j$fY�¼�d��ث�1D@_n�����X�ZV�4�����iq8h!�<XlxVHYEB     400     160خ� ��Oi�ykH4��Ȃ%A��mi�!c��);�ꖼ����Ɏ��&��j�O�Y������Yn���
BG���+[P%�·5����Xf�T�9(ĭ�P;Đ��%�dS�6�f��)���%���}��}J���K��qZc}�ՇṦ���3�a�7���I��`����t-#��=�������v��T푑��m�|���t�6�!�V����%%��=�4�`�T�X��O�8]@�}�~��z��?|���@���{�����X}�_��/X��z�˄Y�X_�&Us��@@�����嶱�t8�D��M��^vܿ$�*�/�iF������)��\R)���XlxVHYEB     400     1b0�w�Zї8���i�����ʰ����]��F)m=�y>�RD��:�0�,�tS��I{�������O���*���{q��E�mb���y1W��t��ꅭ*F!5~�ͫ#أi{U�����hS�^V��h%!A���Y<�܆�/�[�9���z������ �������n��ޢV�0\=���ݞ�l�@�����ZE�'���𾻩e�a����n�K�|��	ҚZT���CR����W�3|őe�;���6��������C��������1�
"�	V%6o�x���9�Kl��Q��~���ό��.��˙q�u\�C|�
d���+b[��)�s����#����:�$��C�7��䉺��\�����;W�8 r�l	B��O���n�3��J}A_AmкXlxVHYEB     400     1608o�b�@I��U����b���aG?C��G>l��<�#�&�sM�b��#�O�iZ�q�~��HR��G�X��ߗ��R5u�MwV_��ӫ�{�m�����N{�.4�������0�1NOE��Ly���m�#��Sn�3h�|��0 �[����`ۈ�1���+�%D�	�Âн�����
j%�4:�u��V�F�Βz���CÙ��T�VZG�F�0p��AjU>n�r�z}����~d�KC�QH6mA��IP��8'E��#�4��^�鼐g�S?O��^	V>bS��˵}w�#�(t��Ffkl"E�����m7$Y����RbB3$}m�\�����f��_XlxVHYEB     400     120��"���}���g�)Qn�@����?�@�(���2"?@O�c��!�F�V_xf�����~_�����>X\]�*�t�xIk�j��}2�O�T��P�vECfC���[j���36�љ�������A�F�q]�� �/���) �H�c��@��-6�0�Y������@FR�j�rS`p�:/d��)?��.�r�~_
�W-�qY�>hD�jB.���(7�˴���4���BU�(H~J���SXED*�cK�D?Z�]���B�}xGxp�f؄���<]��@�V~��j�XlxVHYEB     400     190����oY��cC=��	��K�,=-'Wy"��q���L�U�"���ȼͬ4Ӑ��^`�vq�'��e�j0�B���J�ǁ���u�~���eh�>�n���B�飲�(��["����%�
 ���U��Z�5'~�=�*��M%Ǔ���4��4��fv�H!*fRbVɅ��?�`	�3����}�@Z�J�Q{��"d8s�Pu��k*,Y+%��4��lX|�ij�ڿ`C��k����K''Y��K�0wլ$@��\\���Y]��u�4\9_��D�*"��H��2�.�+�m;.dx6N8��M$�7�"F�<B���3T�0��j���s]�k���K#sr%C��s5�Ya�.x�-蛯1�u�v��菁�gO�9i~�`Y�}�Eȯo�XlxVHYEB     400     140]�c�)�s��
M?��Z$�.I�y��$�R��5��y�֔؉�l,�*]w��yDlu��=�$���n����MQG�Պ�`z��lŻF��H�<��<�?�`�19Q4U�5���X���]~�3�����̾u�	�9��;��$�� �a�D�	,�|�Cbh=�����x��͟�~gq��"��s�La-����eX��wlϒnV�-�� \�9@�tp;�EM�t�s��/�����Cp�]~��w��_A�\C�Q.~X-Yw��K�i��^�ɑ\�@�j#Or�Q�t�X��|��V_���T�:!��$XlxVHYEB     400     160�ɞjj'��¿�/'ū���?yY�L.Չ��:k�xyN3u�W�Uqf
7A�LVn�O0L�S�!���A���H�:QIZ�X��L�-��}qDMJ��<S��Nf#��N���P�|����G�hUx�gv�QQ���ȓ'O.���E~2����܌��sOl�A�5��Kr$T~�,���
�^Gm�K~e���|o��XA5�<�hl��}zo4�m
-�c���X6K�-ŵ�xBe�̆`����ͼ��g&��[�']%U����J�%e�{�����{S����3����zS�<
�]]+�g�H�&o����6�R��AzO?�g��-Z�Y7]c��q4SXlxVHYEB     21a     100#�pû;$�����F���9ο�c���Wo")AC����cj���� ���ݣ��+!����SGͲ��I�g�q<��O&�WC��;XW2�.�F�	uՙ�UUإz��/z�]v���='� �dS^?Z�K������őT�};=��Z�=�m��~o��M����w�UC�k7k*_�z�����/�7P����m�eTŃ�#�J/��݅��֡�9ʳ����y��#��/uQ^��U�V���_
