`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
F2VF7WCtih88I/eCTt/tOSXgiE5I3gWmqprMgwG2Yj5rtM4GPmCi5AC8TuPoDJ7nmkEJDQsMSePO
GqQ6C/fhO6Zvpcl92oqxQr106Wbf6eRS3vBYrELmvtba7t5TKe4PKicHWiRstUbJq6IUOErwxOMh
dhfVqUrqpZQe1Z08tNrQnycrXYT5vTnzSSSuH9NvNuzRlvJtP9lGIyom+ePJekhUZ9OxAo+8eKz3
nnOGvY3kz1IMN9AlEUURGKbWda7ZBuET+M/+elYTPbiw9nArS+StVKZHslqZMOEx6wUP4PnOZs49
4IoMUvS/34VbDHiuUJXNlu56+Bm2j935D52e1scYJhOggbvJwqQFYxL9sWSm6Y1JL+j5neRE9S6P
GQg1nq9x0vx1bidml/2hfKPDO14ESK8EB6mFu8LfWL9ze2Q61PrnKk12bgw+MRzA7/88IuFRqKFe
+/o7c7b6IuKoJtyMO+9/wroXm+KAFjlPM4N9A02Yc1FUqUBRNRrzAicEACFCxnw0jBPnxtXFRdjK
PfZmaOnSFo+QN0BQPK7tRSHQ0swwIR86Rkwd18jeOv1sJ38pziQw080+PkeQik6nc/a+CmH0KUiE
NVPa0aD7ddwoGHYlEmGZKH3bTZmsRvFhHtMW+CG7Mg0tBbYV4MyWhK1LfQmXWGtbyp3OjyNfm8LR
ReM2+18zIrxq5LBXQGMJdg4KYkGPVE5CcNIqQPsDTQJaRAXFRyNyJATnLQDdVLoAhk6rNRNzlwwO
UIIMRA/7ZP7gW7MOfJmh86BHKBPrjhZHq1tmkI90tjdtGHjFqVA7vjvoitzsRDWnTSZEXs3W3+QR
CHToX0E5zV0S0CkdzgncnOtNn56zuwySksj/d7rvQX6o5uwADX0md8QObefivqKCxevV+lGczE4n
0O2jfDn2BcSvfnsDCjTRNEGzLQ91u4KotwJtWmHT+Bmaow6M2u4I0J4ujA/t2JWJt/BRgsgT+QWd
4sZbMCW1k5xx9a6ASmV+5ZHk8Q/mQ74dB0Tu84SVAx2hNwfDVANAElb9bU/9Lo7gVs3SSUE9qYU/
AmM436jo07jyLsGFM8lVNCHMKpU58u+brKLq90fjidIt9vNjWxaxMxuVf2ju8yuwqW2wlPkjDtIF
76gRSE/uYwqKOOwOU3HZaB+1bcrqfQgOctUsKen/KpVvLCIZ+BzI9dq+iQ86EJa0Vy5y4WN+swoG
SAUcWQ5ljXENFoEkq0BYwkYbbKYRN11Vb9sHygeg1oqTsCDXLCdFw0gauj/ocKlHzfTSCtXcgUq2
+KC/c/Hh8Xdxo7+BpVfzfhNyI0r45TEwvufYS0rTxG2Tad5iIUSYlKP7E9Q156RFzXEhaGOERjpO
Hz/mQzUTh54NJyAjggz7Hhyb2EJNKR0ZrCC25Kp66SBY8pYRdGOy+eQzMYtz57Bm4M3SVCUZtOvJ
6bJxy5/RO8Gzb2zZJ/rujDyuPxkjSgoqw8bPcZJaxLkjAfbDFo93Ht7j9RFhTCTkMzM7AdLGg0Il
cR5Q10GeQwTXw6mzCS7Sbth/rgjKalsU3wQNCAi98NdRX8gPYpnlUXnVFPj1fhjbIDIDKZauDmy8
m7j5XNvJKeOYVWQ9NI0XPskqYKlZGMiYdrTEpxt03N5UzF7sriJWpNJUC2mv5qOVLOVRtp6Eyp5x
uIRlPtSpp8KbB4fwldlUolKHbWckhKqI6Q/Ry7CfsJ0yFON48OSizQEis/LckFYQlNO69fNOdhRz
Db6lSROiP/ja9eGvk94UbRTmiijS58h0dHrGyts1ljryvnFPcmcmobKpmMZ8IFvudZCdztlxWfEv
5kgsuF/DJRn+1vjyHuaBcyltRPNs7GMMUhCdNT9eYSSWOSRvpoqKF9moGXxUJ1Y/UB1LZuIh82BZ
Iuzc3EhC335qlako71ctriV1/jodFLFdTWA1Jkr8fzsv1YeCuYMIIfakt6FDwLTNmDfsIJOt8phk
DpRdiFNTYjPXJNRmFAHiDfhW4k8Qhh2UE3Ch+dwwg2Orr392ryRWo21+StFiCmwr/mllTgzc/j15
3xW0PZq5Ac3oEfO+Vej4xFs17c3e6AemI+Xhclk9B5p9l0opZ5FGwHeVysGDba4wV2LIiwMgRdno
1QnK3PapYQrRwC6MrETvqjHSq4R0Uk0wTklwHqbVgndipMoCSs4H6nYTGQ0FR3Sw2NVFSvh/zkVM
fu9aXk182bKohnNm1y5IxVS92VfXL9PBP8Qzq2mw/G4Ik9MK+kaCzb+VZmwdU9wv0z+0dFgYqEtP
jTwhxYobhO5e8JCWjzjJf9evnaEaCsWZt7VoEjvvHhf4CU0oKMDdb/sqPPjHM21hZ7oN373K7Pze
B+XVi4H7XRu6ZD3QRc/vv2FffGbT/lxTW5Wd0biZLh6E1U4AE9Tgzlnf44ADWoYfqqlU1bXGEsYa
uR5OxuNpVznobhTMqjH8atqJhw2Mzbo+qpYwqz3gpIc7IE+VdMp+Uwe0tlE7m8CQoAB3kALbOxgv
WJ7gz6bWbzXZ596oPlD/XodrOhAbrRiT/yOercXDXOqBJ5IyOfQrNUvZzXDTW81Ztf5N2a4wo55i
prjVZWmidfewuG/EePf8J0NXZEgw0V32FtuzKNPF2FJ9uACvkRGWGrcXooxs/GlPDudc6Qm8cNLR
ukVvr/xg2929YT+Xuqwvp5z4m9zHHEl8RrKtbwv2APvSttiwcwYfZCxphZ2hOhRBGXYKYN7Ihk5C
9d8jUpfP6inwGM/oi009m98x3KyyeMtsmsOtEW3f7MKISCIgFVGBFZCCzHZYDoQOFFlg68V1IFWN
j5o4Z7BsQxkFo9XzcBiaMC1YnkrNC+i98LWWMuSE2JWeHQZip7WkmtwcmR2o6TLyTdrApWWUGWXC
z3q9k3jLNT/nSRfpE/cJtXcDb0viU7L00hF8uXVmwKPZykw3kYnSIJd7kfiSWn0Zb8QY06k5N2vU
G7c1hwueOp2Tjbzjk/Mi/m/lnPcKX8mBi2GiPAb/W/WleGh8BHOcuqsuWdjyoLzBHK8X+Ab8OV19
yDTxhTxmqRHnpNP2kpRBPf7g0UYSYf4jAElMpP+WeZt0bHJQZIBCyrA5OiyJxlhokr/dYvqAY/bK
YeLmZ7SHIutTmjYeagtoUIH0NajICbzBBnOhyARfmoXPTW9lo6njCm7RheZXZqF3xnFxpsBoRT2A
PSIAZwI5+5d6bZA7LK6yMojWWvv6YPT7OI5nAKmhNZfw9ktomHhx2s4ur8rVxW9vgG+nDgaDH8oz
Zd4Nj73Au4MQBjERNDm3kafLxk/4emXOdoBTKWdPmK9UoSwu0/xs7bfWobD859L1bfzLm8YxRfrl
+QP6CPpE/r+uEPRdCVjbnhUNiycpk+q4CPdOEEC0tJ48cP5UTf51ZQ3zdsiljqYMGGKmPxmuqfKL
8NezCpBb5aJ1604pGRtb6G8PV92Wjw3e1AXPh4zlKiSvhQzPOaP33Usrk5hf/u6TXg1WG8PRyXJp
P/578VmK3F2ajvm5OveS3yN7NFmxxcNqNYC8X9Iw5dbqjKRIDDfrLL5Lsy2goaqHbck0CojAEfoe
PH/Fsw8cAYL1S5EcrN9zLSwQ5N7/eFmGK2j2wu1MutM90JOhWOviHhPCcU/fqvtX+nBn5wz1CPxL
kbk+s3C2brfiCwdFsmVwGBq3ycDNwOUYx8zqk2VJ1MNBEV8NdT0tFNZ17fN7CQAaOOYI0ss1YA+W
prD8gwbinWrKxI0UY53GavvbXyqOgj+rHot1Vg9hTyMkzB/+qwW8zHqnFs0wXFFDb79faCsp2j1G
Wm60VCeNiQktX5j+lbcodOWgBEIK/9Y8+YSNAwdMjkxqX4uPhy/2mm4FFJFOJc0gTDGplyXZ9+UM
h8ZK1s411HMehBZeXgkuhkLVs2jawf6J0yVu+FVuQYb7MaTKtM5C02x6EwMDWF2mFv2EVAco/zaW
U0JyzPd9oZO3dTUvumqUKdYXR7myBx0D5KzB49NYYYa+8p6FvcYQW4qGmMK2gBGZxj5uaxvS2dT1
AdB+zI3+xsk0EgqbDPfS+TNlaA0U9/c3C6iFtUk2TnvfuVSvRW09g2FPo+uQfnWit5BMb2/07duD
EZ8p9AVDKe5K8tJBzDzJaNyhad9KAmIgbIxuYb1Id0R7dVJz4B8t4bOcSl8TvrQ/nDy0HIWwaAO+
NXyOe8EeOnGTbqGhpy3pQ8QSUWA3SsOIs8gOeaEvjtLtOykQALKK3GipWS5PA4twJWdoPCgb7pI0
dBTvfi1nRL/2eqVnH0pGDQQr7rmyqeGGInaBVtK5rRgA2IezS5/h0hZS3E5+Ewsm9jVkBkJRq/Cc
1cv0Sezh8Ms+sANSCVXugHnQUK2Grfn1MnF88Pw630KJJXsnEYFwkHPaC/mpqxYSl4rHGFG3pjzk
RgiRLHj+rQixRSDUIlfUezruzDj9y/qTos77bch+B8VjdAXPK4TdjOg1LtqNUKFdxpaAsATXPzq/
J4SIj7kqGhmE4uzqn4Sj97R0JUD5V2UCYf7psv2yF8kh1XfoQ7hJLVaWn4rzNqxll+JMp22k1xoQ
uDJVUjXaF0dZ2VA1/l78SQqIunw9uAblIudEOWMQzL3hyoxpwoiRigSTXwIg05GazjLjxIdC7x9M
SCGvRKhoN2Sgzde3x5Kgo1Je00Oqg0gqWMg00YUYqRf6lRwT8UFLE3nnzIBJSKCUQJLH3m60vmxG
uPiywBT0DIEtuZgtJQ1aUERbmF5Jo88CEbC/EGWsbmDGSuWhAlbJ7w3HL8OlRYwJIxc2BtPJ7qWE
h1UjCoQ819YH1PRrs5nYq+VE0he18HH0Ng5kdhEF9V1l07eUF+/03xQJvvyEQiZkQifErEyopS7/
CedMCawW/v6tQsKehZW0ua6k1Qep3NM3GiYbakKHsvzQAoTaVLHKCqPDJScgpWek25dVf/gunwdE
GW+pfI/2qYcVX6Npc3XU+2n5A2miCKbSANzg/dswxrFOA29qxlRbg5ozdqlSLhF3R5p0uxpwuIIL
d9TqwD2livJGnEvkdQJC40el09FVjQp9lhwnW1tu3wQTdLb0htMNDYN0O3LHeLrbQpo/LpLvcdtP
anGEXvFwlok0bPL2H95J8EKmN/0wlhtDq2xP3SY/mlmVzkncr2vz3C6Ysm8QrCSmX9yEEyiRiSRb
J6ipC3YR1c6/ap8ZErJfT1nxB1UlLnxvI3RhOsMX9W23/NsIlHzAz0lwxfnm9o1H97SvMUknIDke
1PDC7Rtv7eEzFShdYgZvZFpsqKhmIikWRb3Hgd4IjIPof2w0bxbrViyugyCvWnWDfWa5Y95iM5FW
7yrwJX3kgDnMGhUc8i0Jc+5b80i+3q0PoxsRAvwVkGdnS/QdekxYxJuNrIQZVeoKAtJVcMn89TpM
Hr5RswwqdGPjO5yFbIt6BA7bhQxz8Ca+lSK+rCQNb3ZehyUxU34tMpe/u0inckjx1CSnWG84R4tW
cVWbHohVScLPCk/6p6PdsAqWkpKFYwhxhpjtxeR+NkhlFZKy0lapGYkkv4wm3/p0KIJ7BoWD9yy7
ARQipRPmCQGFnu3w/+55WoZlDCMsPHqie8b7mofmN95ifeV8TGgYXhNghCb+NzAWohcOGr0xgCvp
MPvOngNFQTIkzD1jUJgmha63InlY1XF30MowZpjiqmpZCxOOrzFGAe3lwCvUbdy2e79y8//kjLCS
990QGkbTx5WhgZmdrQNUcUp4F9y7WpEWDVI1gYzVygz03UAsP5lIgVvDjqaggHkVduy36NHvLu/a
oU4T/SuLahVDn0xi7Mw6gBbETAIN7jwNNGlPaOAOGLLEDGhIu77mO0WE2kUYToDLLPG32eodn0u8
rXZSGetQh8FjJTX+xtfxLFmTBsbe3GrzYjuAyxWwOdwTpG97qlnsvkUW5n8oAlXNTLFoWv+7qhDC
fgIaoOhfmTpvnqYAvtvTCz/pDrjeFuMAtdAhUYGBcKO82ZgG0UlgDrS6BghzU7MhMzdr573TE0u5
FTE4bmValArFEYYIl0NaosLcrUpJ8im69kRimC7mFgM6Fs/82G3fotivcw7onmFLNJedNRhC6crQ
x/yaw8b5hQG/l9N5/nU01YFlIrsuukVU3rUbtvMg/7sjz5twyoR3cIhWbJNHRRPr0yCDj9RQptV8
80FKPURbyMupcjnGmNK+dY379qChJLB5CpFbTSGj89l9YL5d3PDRkMY6OAMo6kS2wQhSo384L6Hz
yFYueyBvxCSVSXJUv0K9ONmLt41Oq4nVVVNF1sXF4jXn49EkCjxi658VeWqC4d10Bqkroca8Vfnv
5n4tGPORTygspAJX0v5YHLjn+MghHNMJZoI+JsUapBWyJenl7hL8aAWRXS1XsUggNxXhYpSPZrec
G+N6piKorj5oPcJa2oWPEwlCkdDI/5oxVR6yNIspVREfcy2DUDjl7mN4P3hdr1YPgLWObzx5U9Hk
aDwJzXYPHdECID5e/lwI2a7ct6frdaNzEQ70oMjYbdmGNjvk+2kgdtt48J6yLz9nMmSJTCMMvY1I
JYrtZYdLxxcKWb4bv3pZLCbPzznXJVOh4yVdQF1rqtNV4P+2VT1SbOJrZAGOqWBWlSqOurUBpa5o
LquNFnz3Q7aPpcWNHNX6KRNh+Pb83oqRbOJga01FjrDn7I5oaMM/5LBLroux8jgtO59Ac7IBGDbW
qyg6i27xurGpfzV+YJPbUhy5Fz2aASuWZgPfxDE04hprGlnz8V6izTulx3OaltEdU/GITPNOJitl
lYNRBr6U9itnVdqMggerkAVPbExXYtjStnEi35M4MnqKDV3pfyZW3tQWxBopqeVLSud+/ShVvXiv
6uw/1bUHFimdNsweEOkl0vV0C553FhYZF0MRHzpDO5ixOjyjsTgZyhPI6lDqWsnr6dFikKf8XTgA
iOInoSV5McipzUpajD54SpiAtlE0guO4bm56GOgSgXsT4z5l0cn4U0Kc1LTv5rW6ewxE3KZ2Idf+
yu7EkKpW8lhdI9+RTjItCa5r4Vcv92NfDKJ3iPzpQs7ohsgok2oe4xT/Xn+92CdlOhBTftvaalwK
5fxD3NN3yeRa1Zk56jvtipfo5ehqE8MEWSLB21Y1Q+ppOTY3i6jCvOlJyMiQwGkDY2f3SEJ7S72a
jNFUN8sFIU49n5Q64ziBC+FhAnOYvFcDjX6h0H9hkJ0ZGOoQU/8WifE9hdTyATBzERdd/MF/iA3Y
lDYjtqwxwnua3EoYees/CIVzz2uC+vBJz+g1fDitvZ27VvumIXTNmT3featraKZPadGHagRt3p8w
iGgUi1oV2aDill+iqc/of1H5Hokx4O8m1AM19CmjFAHmGldP127L6qtkMFXlPucxaOiYo7Qncaqi
FBscPDvq5bl6q+CBUpH2wKJXGCYS0miTYI9XHmqdRSZYeJjrr9cUFXCCGXe40WoMHAazBcIzNiUe
SWZciglpmUJ5QzSERkms8oDzT3q3oIK9oDReyH92MW9HlKWxcuZ5fgmldDeLnnHHgvPbtRj2soob
t21g2jbyXQHzqmSLz/K3tELoEwDymlcCI8ms5zCT8IkVEqaYXEEPEZeGa9Z/eY72t2zAHk16Apgg
GVeZ7ozRmSK4p2Po2q2ia3zTk8pZCs9aCerQlC69LWux3q2B3MkleZYsnnCN0zStyo/+2zojWwyT
+FDpYEE5MWDVFXzMiylxhPTxynlzKWfLg6ZU3fD9J3riVb0xSq5gfpG1CJoS5+Xu2Sa6UOIJAzKQ
vwhNxmx+qZqOKuKQ+3iFgWJPMDjD9sHU+mSqzDA8J6vV2KbguTa2ZR1Fgk4du92SQ5J9y8Y3nzkX
hQyMyfO4JUngIy6rQjJqSi/8kvMouxKDmMeCrl79SewjtFs/Peur6EQK3FvKjwScrH0IR27SGB5k
rX+iXWTiSS6AXjpriFZ2GcPvv/B0ncrIAV6pisx/WZTI0wodP/FH+y7LbJFx3878LEN9f5ofbUK3
HBEhbGaaXY1BgcaONioYJi3OIDrXzR5JWul+2rbvquJwt+UzE+EZxul7WAujBcUCYXN5B4Gxx3lN
vP3mOcZfRKaszKDJobwzywEMS3YwjKUAlNNTIsmZo8LGBMo00k+zREagg/GxuUMdEkI+iDOi+Fxa
EvxdhvBbdft0xh/79LjcpvQr24iUNmKVrrNXr0D+88IpBEklc+H4c51lsnj4pA24vbmVXCozMKpd
CsbsmQCIcq5twcWWNXSrFCaDgS1hDLIUkp1acpHchZicvlYzp4KhcChidfNmBi9BIg9Lu5iSuiGu
s7Ed/gH746AkSMZCqK3E6saK+X5vpKyLsqMhQLapYXVB8SHT/PvnolVSpOZUdlDpfui3l8+ksRch
PvjNrk6b8t810q6mSF/XLdjK4fi4SmMyoKz+upw14cofSL5Kicg1wrozjo2A1OOMtcbko8lBRCGK
UR5s6g7TQ0tVcBeuQNLtKV/irVyydV3EIOFCNIbbJ6a4len9abT3HjJYpOGkzYLyZ/HA2dPKFIHk
W6/J+ekttOsV+edxCThi8ph41ZoO//XlY3ouhtEEwmYMU+apVT/mS/FtoQWiaeet6qGknp+rFde1
+fYqXhHzxE/Lks1l22UgymF8MaFY4hPF4FnEmUYBt3wT3Ic6zcG481498o+sK9EU5Tc6OFmPzmtk
ha8ONa+95w/rbGDJBg3KzBeDuGrl9xkv+1/+CWpkPda8nIJCZ5uUsvFp2BBr2Zy/TXIV9uu7wJUK
GKaNQncDhz7r+iGb8x+ocRhM9jlYGYl5Zeju++oXaEj5dUJkiHKsBNCq+9xZ1jdMYM2h7Tt6wwyv
s7F2+IaCfU9TmRUrgvliazH/bVB0Qi26O3O5+4gs67uAtiVNzjEOE5IP1+Y5Us9cl1WXoLUMBiZe
JdNWq1LYjdfHWn/hD7AwEF3VB6Hygbhw1vmiehv3loJIPCvAuoeLkJPM+a8EmpJGgtb6hHFYAYib
wj5v7PKxmCotEELbZ4tEwG9/59ysGlBTAMIDkyH70exmNYNvs2/qlVQNEXBm9hIsD9rfwS7gqMax
0vUhp8U3dKAG3Aw3Qo9jtGDT8RIOo1dfQyKGrkYksVQgbSdEFl2JO4WaYO4zYh+Mgtq35pZds/Bl
uK2QiIONCe7bu5kE/OvVqXDXqRw6AytEYcayu11DgtwOrZOs/vHBe87Zxdx3JESgoiPW+/ADEuiC
Sp9M4PwZfp7zSdkErStqni63Qjh3ei5RsKolmDHxPJdMoXFSkjJw7jg4z/i33Fxe5dCjmjVzsikF
VgkZSGtCGfadK1+temr2A+Dm6YQxLZ+bS6xHF2ALiM/O+SCHqSfhyN5bO43O5sxNIXNV6GQOU+zZ
C5MY++ikUQWVxwf9CwdRM0coOWASA3dOH9plzS5dKDuJKNFu1Df2GCWNKOe2iAK5pX2PfQQbf8ct
cGtPl1lEXz/j8ypxWpheHrlWeq8LslvGp/Uml3nkn8jcH4ATooRs6R/bkSkM0N9FFMjVbAmbpjMy
1gZg8KjqKwpGcv3VJB8gjUhSWaciXcMundq7EH6unnIQVkv/cj68WdKaa6Ru/pYLL/UAwbf+cuL2
Y9NbNy5whygAy38qwVoVbTKPwTde48SsLHLgNqJtd6fycrRpy3I/x3FxAtu2hLxAVpEXPUJOPswG
AnYkLJv7B7kaxfIUG6MPmj0z0y4RRQ0a68ts8DDnoByp45SeLWtBDtq9oatLEs/cb05FcsGZgcDN
BsR+Rod01F9wZuCOm3MlLncxxdsaPTqx7sO1sxNmqAw3Qy5ySPQqyrH8nu5WJUgHWTe1djGlTFEt
yK1/aEwQsZ5d/OLMC2IPNdnerfSalmJtPgjEaiIsVp/9MGyRZWIg/SexYg1esUe3MMTLeoK+13sh
XMw3ygxY+ViRWPMoywmKYtYvdRBLJRhlxeD32IiYSdwrXHSEE0i82ulr73llgJSUNhK6q5ft4qU7
o6Gp5p0CrdvZHeA//JPPmuUKdWP55q4/XQImaH36TFaYvTHtuxtC7BHowDYayxcfL1k/Eb8wUr6J
GLqeCW3ZIOK5j5MY3hiJBAJR6CtvAwDaSJo93urLXGdGiTKmtey8UdAdqcML0tTZX2nCKNedP96k
OJ6GmXlr79YCddoxiP6IfsLgrk9yo1aMLw6AHOM3ytyLLYiC9QOFm3J86wKy4D7muqvcuDVmIdzw
xv9Y8MIGRgv+itKNpHHPeobF2iZ24o/SCobV4PZ7KT8TmTVXzu+TkBxK/X975drLI5nP33bOoAag
ZMh9qr09wMwPWenf4IklR9B7QiuUfSZhd/4Tc4hVOAQDaQY+/kE1W5FlUpYcC4xB4928JCMNZTY7
1IdmOt8kbR0WCMXp9POZ4UmwfNoyJl6Gf5eqNSZXPWyeznjItAkiF+Sd2bWP3Bc7wZSxVfgoOfok
tBsW+P0MaQCcqo4p4PvqIcjkOADlmje2E3ssGKl6kWCqmh0hZNb+cfZmlJTWYcMGTY923tYRd1ED
mJA8NxhRI1U9K8wcCFqEoe/QhhqSr5RnhnUeB8v3grpeeFARMoo4xY9sPMWu4xklvMbtKd4AqyWa
LR2xFhiHkdylIBRCd0tBW1fY1E1Xjr4B73gOmP50h9Jz8YaWzyv2UjXp6UCHzMtzNv9LQTRtePPu
qdnTMHT+ghKaZb+LhTxIWVT8fJjmfXNNTfnv8qnB+UqP6zr1oscdD+HldGL0Ted9VkBqOCIg/TmE
sZpwHDiaCBC15bwdF1HftETsW+waI6WpZamrLnN7NVYSh1IvgFEjaAaWZj76+/XTTY4SVXjE+TO1
uWIq36NKhxGysDtzuu/M7nPxgO+hSPCcG6qTJiFEH2Ckcemb95Q4FJ+DxqYgytmTQgv+ZzPE5oOq
4gFefwSxsdOVtnpYdJ7qt0zFpFEtlSeeeVJo170p02WFhlCPDeMEK1YTBuE8RT5U2wVAln4yPQDu
2y6RApTxaEkygttWAY8W9fyhfBPZOOGYyusPiZv7AfVPaucYRKN1bHQ0uJgNyTXEo3Y4kMH+Nh9W
8ThVr+NKmrhOpR18RQJMDM8/tjBog8g1/oe8vtN19TVXwqCcHq0ytQI9unxxSLxer00TXPFblXYd
R4iA/3h9Qfq+yR9qDATKAVDgnj1GOp7ix3U25LlrmdZE1mc+O5mCdu4xO09Z8BgdosX0aXAuIomH
dIAU1p7zaVMAjt3RX2SzLW8z2IVtSb3+ARjnGxYZb9l78Llf5X1hlyvx+67cwc2L0aooeSkCXH7a
dRdTTZKGG2JPXJq413FGzOgpA7oHISfGuPiVcmmrM5mMgEN6+dUr1hL8LnnSFT/2jlDI1sP8z/MC
7ORcJKOOtrZiqHCuLjWtvUQKROgEI//fzPXPLM9fMhNlnUfWv1Gob9J1sF7/Bx4XJ7h/KmQRSLkf
pe2MFvFLiBa+v5M9GLarrWojWEUYXgEYNM49ofj4J3hd27XSBtE42E0m/NHIR+25KY7mjPJoijMp
LxdcP2hPOCIlSHgIixHBoLqxNx+GTQOz4JTChu+/hnMUQ7wSVHuiccmNSHGrcLIXPMgt8IZhnYfT
i+218iu7kilnQoB4g0m1npM8Gzayh39ATj2U9082Q5vw7dbMFHEVH07DBlPC8FvrxzxIBc/5T7XX
zupiEFgCdzHexHz6PXCXTu4a2nqnG1zLQDmxdyBunu6NFk5x6ozjkpKNRPJ+x2ieLn9/p0I/CedY
PU5ISjUsFF928ux1KwXuvPb7UxXpvqDgdlHopPoxxijXhSowe8zOeKu+ph8l/20TsR1zg6+SR+HA
zk7zZFSmk0tzh6z6AdIguSqftp+p8SLejIaL/VPD/xDBFYlSR2v9AzhYRzCyxn9zg8+UvnzDazfE
DjZCtJuKwJ0kAZKjSzeD6WcTxBkwiUhOYp44VdoScH+ifaFFbs/zMXZ0HfGxg/lJsmLOCou3YBIm
1pYA9hWSiDmRkgq37xG5YF6g+Ccv6M/EDjwAAs3UtT0ZvX4nXUUFPa2UY+fcsGLyXXvn/sxtIAwM
7az1junbVDeGOLtM4sW2oXBYwTfa7C/a9TV4gYnhi5weCfgy3a6ewx/pu3ywUfKG3fpXEFtrl13Q
/I2Iq50iUXlalPMzD4fwP8bcIOK+R5QxDC8/IXgWqRTi2ySXtYXgjvRdYq6D6pG6P7qV5p8LQVhA
0cPdp8p2gYislCzH8BWSv38Bf4yXhz05kJuNW4MR00PhukOzBYxOy6wVXmaBsXu+dM3i5M1qy1dg
FWrY8NfQsfM+uZUVX3uvgeDWqgXrQJI2SNRnvrlLKzoS2085dpSNjUbht4YuWk9R2nEgOJ8OgQXk
NxuR/v2LiwzE4SgUt5jwFZYoMC4an6/hIr+TG/22XrWL3NAXfFSO+QUYzgApkCIuDd2Mbv1EaPMa
rYlhQqJA9pfgpwpXfY9vU5/T/HnRGrHt+KwvOKxBU1XQiUVtGRBgNM4y0XFn5347s7li26rSe24g
6dmFv9sFaJH/3mpBVArvZXz72HqwcmQOYDGc2nEeULI/ThQ+KBPWclDL4UecI/LqERfNjmIEJ/a3
OzpPt098nC1MVV5Cg8HukmnHCWZzZk7euYEzY+VU/CEH+KTi66/IzljOEeBQG5m3/2qRiMYctAzO
f6/7JEmyCiYD9nEVvn+k+2KTih9rxQH81tRc64axRrRpCSJIegPJ+MzO+lPp/dkGTkTLAbHpXxxW
LrUUQJoagqw/F0Jg+LQ6/zUwD6YuSff26kUEFQL+Ny7D0X5jhPwV5XhY+knpGFomwRPSrWeNXm4j
M/WA/wSad9dNPBGMGhiw9EvSgRh/rGe1NOSBZLA0zDedlurKs3R6fdCeqVZg16a4S8747H/sdhlJ
UOiXqCmzDKQh5jjjeWXlt1yBHG00HqG6cCdnB5y4aHIYu3XBZIwZQO3sMvbz6E26qcULk5egdl7Z
QK8hgerPUWmJ9dAl3D5HwdMyUyqDjg9Qzca2TBsGd1ehXxNVrXafQzKuiOP4fc3rZmBadkdYs2QO
ti0HfC38MvcvUXRf/pVAM+fIzaioVht3Qfuvbp+N+CbEg0aNA+CPZz1U6S1OnqOrLwcxqWd8KLA/
oS/EFJ59S+4pwyiuIqHY3p2gPGMjNfMMszGVhJpEj8kDVo1fKS8kA/+oAfN7KvOuUbLsCny86dM5
BkU8fRNY8uOglsKp9F9FJuGqevgbWZjmII3CHO4JlHV1G/ml9fjPaeChGmUqSA84v21t3+cLIk41
Y58sKOXwx7oVdpZQV2lEYpJ+HW2aLHerrWLySHNUIgn4N/U8x8N9ThAQJPKWc+ewwCkBq40iO7m1
LRLhAPs6yscFAcjlQUOgy5QSZcJ0+k5H8YjLo8ZDiylSnJhAIiAutUtp0aTbLjUs/QOkeDotC6We
hBw6TLRyH32ndhx1kn39UdYYUFW5LKSkpmyzWuZNfwnewLKX2kPvfMi78kHJt2tvbN7/99rIdYaa
M3kbN8m9IsXANe9iVfbW2Ihf7AXEijLwUZKHCKcecUPJjENH0jVav2NUkpViJRbQ7QhziL3R1rVU
Ui52CranGcgaKCBcpvk2antTxFoxu/UV2z0pCJwdzIe4VAWT5+FJg2EaN4UTwIPnv8rsAXTWZhr3
X/ckZ8Ojbw8dx4fpbGuiGpTSa76RoTLEFZBQtKhp/8W/QhVuTJKGTxCJ0Adz+nYlbHRpPfs7GVjg
fA9ncuW9hDgNcFkUxsCFzpVT7VetZQYUXjyqnW0G+z8NGT17pBSQ/0EPHoFYh7X/GXEhlwQpjz7Z
C1ySEur67iH3jIAXbSkEP7nu0tZGcdLnFelTT4YeaunpxUAR0NqPRJUfd9CVSrMEr13TB34WvJld
8wscQ1IiXqbCxW59Ji7E2iZaOBZKn3YlCjCjBe6qYBad84lg13C6koO/QIg4lKiippTh5BRZFrqb
zslmSghVqHYZte9x1HjyG5ouZsLfEr/4VkDqp9qlWCIOykEib9uGD9k1eDEIy/d/tr9dMqzscfdd
chiBdEduXR9jWmbf+yBGwKm/BeqkFKorw10o5YgkPJP5VFd+PJ1GNj+v+aTuVsdT8lUFSldh3Rlz
TjFBWlHK7eMqJka406pocX5ZxzNYahNGtyAfsL2dyHENXbqkfPBYYmg0eX8UvTiXoK9r4sLOSP5L
QfCB0Rxk/n1iLPhFekIPS/bjtXFKNH9vpYo46xvoRhjrwkTvBB8th/8t6aJVL76Yyd3zK19JVEt0
XAhbx/1KVq9t9EKGAmYE1vsOZMUp2bhHx1rBSysqokRrQFfEyvtB5V/lq3HHeRpDHRbw77S1L25d
rlIxm9LdxECwAoMdeBdt53Q566CsmPyJWXDqRUceupQxznbbx/ejuVFd5f6yb40Hsck4WXRAtq7P
2clXbfuGTIbD7E9dQwiTxWkxPIlqjYUTbCgykidUtqZ8uLrxdiT5MGqaSYwcKmBqT1+P1fG3i/Vl
/Q8XYcUgR5JJtz+WHX8SFCOkBnktX4jb6Ad4nx9in6+JHGs7fl9Sv7B9bZ85IiJQA8m8gEI67W2i
dvf7Ch2OTPE1/WAYcEe0+KUYuqZM2NreHhdnYJnSMNytTIGa8EOdSkrct+8lTz2fL+C6b8GWLaxB
Oj/CtXbOKw5mixNtq+b/SbDTnVH4uz/2Jl/4eg4hPQ8Oa0ZhkOxN6BpVqIBRvBbLdAgzrW04Z2oV
Mz+MS8UIUbcqCwaY0iZnf8v7i6yVehpgXqvwOWb1XzWt1gfxseWR3A8XSio9X3KuGhzNIZNQs/b0
7CWAlqGPtiLuKrN8JweW9Rna9VlzZXwUj4kdJ/ZAED6Wafl/LrceoxOjylc9y6xemJayLQVTX3CL
Vw+isKd0YLWDv4N2xbTzLDO/5gipE/TxScbO5GpAFKV+UljWPPStT5zJB7dDDzpy218xGQmFuqNm
Ke8qlUFYgJHm8OpPBI3+FrSFTD9Y7hOtci1H7bTJKx+XEylF5NUG2TGtViI0KqI4zZzWKvAtGYfE
Ox6Chd/+gCj3YpYJVNrFU30ioxTDigqQhsPUhZiefBWN6izTjvViESF748J1pl8Rxi7fhYvWWUCM
nShytJwX1gOJKNmIiam/OSwDW3daSN/nb6JPmFms2at8cN63LoJ5itJHyZkAI+TUu0VstvG+6onD
jSdIuQ9A29VJ/yDbCtwUzjo7c+5Ijr7IgjxiwbT2/ije+MHtlfHEAsijEnMxqtuVLVlbCjLrTsbL
JW8khnHB/0HXHCWT7i6dfBbppVQVfXNECyPPTS/RTngUucoC7FaDv7ISVPH8ec6y28W93rSqtVyq
bgvHoLWQV5KBkX87MnI6F277nKwK+lekxaTWt6BZ+xjOuYdfP3Kwi9FBogTD+FULcPDiHLRQIHK8
YnhPZgGbsips1Dh61e9ZXrLLLeEUjsBPV0xQKehNqfCf8W8vsOZnGIFAgMEfJYCg0YvlMDK55zKK
J0wjd9lYbniRpvcyUCSSbVgpNrs3349O1ccjmRBjAyq3kTV3Yf4hLMK0TwJXEqUX9DSrJ3UPOBGc
LDWrnvTUsJt41PBAQD3fMAhI929jB4Hj+RehidYMJDEarqONiZt4oGuiyIqohxfL8GUxQ6Fb/tTv
1RV5Dw+lcXUEOkWZZVYm+fj1SHiHYO+9hMEuiFKd0riWLbU9mz31b+kw4PFDqZyVulusBym7Vogu
aqXa3i7BJ9IT0Kuoq+aP8WzEDG91oeNmBb0j/EEq0iJRpwMd3MoW4jF0QmpQR/QOojxOi8WE3Eo3
zEh12+YhmsXeZgg4NKurwBltzc2z/Jr5TpHDdcX5WF2Pwk6CBYAhVo8ySTe0JOlc2MoYAHD3NVRx
rqzihpT6FTVSYjS2tVUvzXA1opBIT/EvZtNulPONfPbyU1XvIt1Mo1Hd1luW6ECzm11KKH9g1Ahg
q9EHV/ItnXsNBzkEdTmVeek+dhK0UCZE1mGudLJGnZGz8roIKSA6LmALMZhlolI1SrCciPN4gIx/
KK9ulhCV0ZQcx+oJxG9UhcVVgjYxVykqKIkG9NTgPkV09XVghOJm+yNR2hffN5O3n/zp4ePO95+n
etMd4KEbWSuYFtLrRZSWTyeY+/NDhdw6L0CZ8q8Sgpm106tbtA2sMRu2Mn03pWMZC39oVhWLeq5w
PjyyxWekwAVV/jOklCd3oDeNsmqC1suVIv5qp6d72Muwm3eFqMtSreGSe5/JEdoY9a6kN7q748vZ
meygQQF2NdERrbMR0zApoFCJxxWvF213i4O5a7BNN/PbF47yxmheGBFQTNW/QSZFa4WmlUKBp05v
Hhva3BLOYMWepbBAP/cr3l1RrpgfIZiGggAZnUKteHeJ4sjut9wlXYV3d+j6EGJCBmLDNrNDBOHk
2kamqEXvEu3Nmf6TLoQ8L4jt7eDn+66dHRsDAjqP5nO5yYZ2xO1E6rHpH9HWuGD+WKnYfB24FZRz
gBSRVNL/WON/uemumBWTiDsiMkdBwfhRCF+ZYd5ZDLU30zddyVTdCkSA5FyIOtZN3QyQsZRTq/qC
hP3C6jX+w39Xd6R54GsRAJiC0WOmFF+NmSaYTxXjqPy6ivxQnjfphTRhajRvgks2puZyDkyxl2gl
Y80Y82wbMOgAeWJCm1VkU7F545TeDclgwLXchxGpvN8uqxjo25NimVdu3ePpLeKmG+E7fKMMLtmL
mcSoegPWjKIyXVqAFFf0rjs0mfUxF2Hvzj82NxQMcKBF2XnkGUCWmOxK/6rY6lQS2jtXvm5zCUBr
5JS9072DksCbOS8nFT2npNwlUoVpbjaFWC9d3/jT9QTWgWCDVJIb9mft8XDxO8xILrC3FONYmJaN
NP9734FQTd4h8Zvvlkn51uftnOyv7DQcyJi/bBNGcVX2ldeMAFKNgcOk57mDQzb2zSAd4OXLJmQd
JZIiwPGfXCb9XFl1qxa7LpDH0Ti2UpVXyOM1f+errYr6QHlmhgsboCjv8MMfujMNzWYYqtVmaHiQ
olaRVFfiMD+QuuzQn6seBucgAB3HqUygPKl9/u0h5c3dYTPQj2W5R//8x6Wm90fOn9nF1s0iofV/
MdIwLWiPkvQWB1qw6p9XBS1TqAXL1G1EaN+2bk6uOFJna2UUujXIXALo4xxW2StiV70+WUQGS7Nj
VXi46sWi+OMQAzlkvkWrd9ZKQJH2M3b7AgZXHP6db+ejQg74P+kM0I8Dql+iCJzM8e4jsU3yluYK
BqiWKzjEdZFEn4wWvCEaqZnJwVrhuM8zy4RZgYm5zqBMesf1hEmqnqRAzA/rqAVFi43ijzENx/Hy
MaqFiwhOGCVkgfU3SpCoJgRLwuUoYf5UQv0uSnBo1UbCB2GLLVZFfP/MowsWNpggCFnXMdMhsimC
v3jhmk266zmsFuVw7VMB1raiIe4z+KNZw7aU71+QMrsQRGRaXqAfY8B9bUzp6czQyCiCIIJk/wjN
RjYMOK7F0Ct3s/9YJO8Cj4hquxPe1NRUZIIYh9Ac3EHul0TQBL/7NCyhBApEO8jqR+CLqiV7tLXI
0YzP7ehGky8hPEPqkvQEjjxLXTKPIbj1GVDhTXfX4yKKEzjEUBQENYNEcYlgi/hk18vqbe1gtcm5
SKFLs2uBRGYP28/AqAH7UtmXFEH+j1rEcotJ66fpjKczQ7iQ95Dq07+F02NZSkKpFRp/46X6j2d3
S95GXc1pRSkWViw15oFTz+C51it/6U//PDMSxo4ROVJBvxMsjG/RP971Cf+qJhzZqXS/2D6XcTZ6
fzbU0WB2JYG8a7sc2ebXGX/vbf8akeOxWtmxU9fkkvsTBkY0YqN2ti4kyCRh3OTgf+FkptP9Kbkk
lfYYBHx1uoJnhVxhpaK4D38K7wNiESgrs3pspGRD5rAOlyaieP1u09mg8yw/HDm8UtjMl72qlAMZ
QLuY+9AQwACEbR+GoWgoMbBVAnBqvUljqxuAiQNrN7upHw6XGHls/T7xgKSvmVSFbKXDPq/lrMx9
LMY4du2d4KafnPUMV/NevIgRkML+mkZMwmisadeBcJrT2r+7m9B8pvngmzyMWL+zPjxRSwXe5sIQ
ZA378m47uDRO6LPkt5RYY9ZC8hsliEVxTyTh3BZGyfaU0HYdCY5oefYO9RD1KEb/Q+PUEe7Qbiuw
QYop2adDSMUsUz063Xb0K3aNnTY9F+zfRiHCcXQ61oGgPkUnGKUI+pof+BlExiWR22zkuyVe5Td5
/sV4knAsu1HiwGlPymBoubT6yiV8RkbkNhA9G0HmeQG1k+9qVTKtzNxvKKMc0n6C4HSE0tTyz7Gg
vvbbRamZ5TfRBdm80chEAPyIE20SNdLWVAxwJROSgVNNPoD6uychHLPXweJ558fker4RY0Fnpn6w
dwNf5/8+/QU0f7HV/qqgwa4XhuZrhPfCGN7etk65Ft+XDpyLaED3KfoT19TIwdyjl4MXluY6h9d3
i9M4uDr14xTHvcjJ55nVP+itb+n9QtqqJ4WU7zY6wTn4meMc3YOPyQeIITOScyZFxCp1E2pm6owr
zw8nMH6IkdgueKcj+orzS6kFxIXwAUMz1JpCdh7nrL5NpXAQf1jqTbVDGqJxBpAIdPb7SZ0Lb682
vqi2XIpFjp7vyQyJ
`protect end_protected
