`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
JHOQf/4bgGdqvPbbwecocvhEUdNUcHx9MD98u8SGwdTbMlb6cgIvYeccOBDTFhY0uJe8S7bNwkcH
VxrlbwwCWe3PxIZCjuqDIFKxa4CWxYfb3DC0zgFjpOhZ46bdRpb2IFkgQ7OCAiJPOE0v083y6Df+
RfVyE1/c2Fj8fU2s5FQwRqQkt/M32uDmw8eRIRnstsnLqPKSzXsKAnKzjx2NU+x8up97ovPKXRnN
6t8m7W9hIm1X7BIaKohpGIBoNFTQdhnU8ou577yxcEvobLN01goKlyjHowQ2fXod/Azle3YyXOCh
0OmCAf6JgeVvfSVlamd+vAP0C4Af3PP090IZEPqQfhJ+uwdAR2gpnHofmOfUFxUY02tcy2nJM0xJ
DzFxs8uo9Ia1GSQbEhBl7Wl0lVM7HNRhqEsC8hjKjg0dJfejV24Q1antlG/opC0ciZlmzLrqg4K0
R5DfSe7jIlTCVnDvUXwurXQSwl6n7kYCLRjl4tcXHhs7m7qQLTu/U6sAAREo9mWIcJrfYYUEP6b9
/zyaHmVUiBkabzqrbVIqWGFmBxnuDp0uX0TDjt1WhAdH0EHYgFtyN7Aqxnzq6Q1xNJd4CZYSgfCY
HLdVoaeycVR0/4AtqmUAgVNevH4KBLga+qITIC66Kt1bV2+B7inzQkopR5ciVGvC2GtzaRVxzpb5
3sMV/iC0T8GzALr12ib3x24d1LwKrGf1vxhCdl/SYRdSFtSyTdbszCUW7DbnVABX/688vTt11o18
+9LhRWYhJjs4P7C+feaAzZQpzJWmGCJ6Ij5ac8L+RItm/Achou4PDnRnNbI8akdesoHGxTTzoZBX
/75Be8GYjQMMu4TeaEsCBUWaaHWudFJEN1j1c+AEBB0YaqoGTqFak95QS7DsmuZEihZuacQksohX
DpNa282HHB2D9UsAD2FuCxMZH6VtVHvpRa13zDFQ7l4G5tDbesyH5cTXy8T/OtGdjMKBYm3/iICX
igrqK/ecqBc7w0cZRdwvLeZFE0vM1/aJBa2aZG/6CG52CaOyUS5dtuqmj1jRAA3orVkeuFbUOzXm
uIOk/1ngrpqRrdZ8kKGVhGYWCqc00+UDf76UtC5BYwS9QwooE8Y5PZYzMYUuqOBa+UDGlJzOKAbQ
wB5CR7mcgiLFPpY0m6q+KWm52POpVJBONtf8YEkAlenFoQENVGIhataGyqu2igpvQDvoJV36o5Oe
mh0H/vi8QmhFoZgCMpfR6d0dkSPoD3n0PZEcATQDmtRKbjMMGi7BDQD/4Q6rqUO+aDx6Z9qpb/+Q
m7ZjsIyq0JhjrbXffZ75GG3XaxF1o80atJig6KgY5YUfsU3ct/h4THrpvVGC/kNGkTW8z0LWkCzn
RHxu24ZjabmLVx7PhHcRKGfLmBtBDrSq3Wo/enEWq9wfMMbwM1JYP3hx2vODhdWfrYN6CCZMkGDg
BxrVnTykALivSl0Pr3g22ynprU8i8JYqrDA6f/9Vk637N9hYR7B8XLqigqpOg00m9VLuq5D0owjo
k+xDH3SpWCe7xOvJZxfrNJjDxr8C1MUDry4zrzd/JZyuLC7ZYmW4S6HfVzGJt1YdU/xsXLp32vdH
TGgdM8kanWjwi/C3vQw++fsHPOlCp3sOWM5xIMR3tZuV8TZhJ6hr6QQ/V0jSS0Nflq0ueUTh5U4d
N29btfIZ2QgkNM5FGfmTGk7DC2YUR7gJH7uS/5ziaRrKGatOuPU++7JUVMzVbZQVnFvItpSKxYo1
EbDFR2lqsTk3mP3PprpiyoffXflCUXyyvk4+h/cPRSGv5Ph0SML98nUagkpzLtCBXxeP+nUaoGTe
4A7wC+saVu5Q0iRg6kqMy+8oX8slVzdB3dljo3CJ4VjbNVgfALdVP0VCuq2d4QgCHY9c5U6CbSsL
vRAkjgzJVj3hz2uCdtcnkQtI+uWMN1OAnErTQFTLpm8LBjcw/4Flm7xc4Bnl3fT8B2P6t3yXlmFW
eVPHIb4RlMRguNNG3rKHSzMUOhhpeBBufsuwJE4ZRvWkQCBRfW+4RzZWIey9e9hWJio6RNN0+tm6
Osue4grVJr5nQXGChDwnj3kDd1c6FCHac9n4BKf2YkAOxZ/qCJi4Dxkg33nYFrg1V8OUGv66+518
1AcjLud/PbvABIcVhtMki5I3IJpGcGuhjZ4Pf/EtxRckT8S3T5/XGT4rE/3byJ216IrUqjchXZLA
LYvloBuMM+x95JfW1rmIA/L/bzdA1eVWnQlSp5n45W3XhPkbIpJ9nUfwLIav3UkL/1mIt5USvAQg
/zqaGQ/aVPqya2T96BRyoYCTfmYQzHoP9dMr1wGaRHXngMIQsI31EXYjxZyM/3zhamBRbAGOXd3k
oLSDhn3bQF+2XSxu3mCha2ALWoAwQilHzzyeja/NCs4xJA4i78R3HH8etqV9V6vUTyOgtBTqaiPL
QXvjx8rWGNhWu9psd2ewkToi9nwGFBtutB/vs0gnLRgJ3pXUaw60OcgQLOT6UrKAkTxDL9bjZus7
8dFKta+rqzYHRNfoSID7jbebVlLrC6Kg2BTkuVZHSbKVJ1GhBYO/VJKjA1/vVY2ycoMDmEa0DojT
30m7TA+GsiQcOdVlg2dAgYZxBV6xuH3zjXqvC6muMOkTDcgUYeAxXToUv3f3T2GPMdU+cW+VMabz
SUjVF77Z5WCTX2LYj+izgJ39dOzHfmOQpPHFClkxIkbTSVMBW72pQ1tKcyOre09HfZoPz4cRifa4
jY5lye3zCaC9ncjsdk8KKxVcttUxc7xubnxa4u2PJUpOacG0PNpTYlhpB/rtZUic8VO2pbjrSwiP
3r6GzeSQzbBuV5Z5DBD9VJrfPSa5btyRjNvCTdp5maW3Tb9T5YsTAD5fz4Fgxxdg0tfjaKrKZhE9
ToYH88UPgOfbrhsDV1PYW3D+tcfWebt4e4yuGrTd6WXYFAKSyZBT65AJ0/edstx/Ou1YmxWraQyu
9lqZohf61ouPFDmsSlqub0jUSC8YIpHA1f4Yz45J7U6da64RpLLwJSz0RQrVUHnQfB1bIMxbzhzk
JfzL/247Bg6O5xaMC5oqxjFBx624+qCJ7gWjE9ZJRS7sG1PiSb8oBtN5QDRu/tsxYRedyS6IzhR1
r1Lj8+qURFdCWld3zp1UW3G8Ciy/R7iYKU4lfJ+lgrkEK8P38+6yDwXxMUklOX+XmmSo76LUY3l+
2CuIQV6yPf9d2SX7ru7Ss4GUrnrRQSsmuT6CP3yypuPVJv+ztHOManpqpViYNbZUL15qwNARpoxL
R2blLC5bpk/FKVGvrrXZOvi7105iAsKvUMwHGcURKEtn8S3MCnyb5JTXAYrBPGexNUfzq0RzRjFX
nPzKz+SogSm59bdfjRASOWDvHTysYgRZgBS7/KyOs31f3Dzgx4jeMD11WMREZCCfG+T5y6YItSU9
iFi/mzzI2IYEq8ehRYS1vuKgZ85O1xdukAN6G4Lw6moYX7Wto1d6UEXpL+aZKM50t9GV0ms58kx7
Xqmk1lyRuO8pVChREab3fVQGFn77iTmMxCgHyo4Q+7zHzQfoClKDB+oDnv4P2ZJQZdxVEiV/DGUI
Zbtpp/drYIW0p92MrA5vAiXfk+QFQbZAQWCYx9PuGF868Ob8Xn4PNcEIGxYf3ppBYucUboShYVSY
z8tV92MgtDJkPR9Kd3noQPLvyy35ssVspALy/BQVNAdXQd31hkgHC0xYYNBy1kQ2XDF5lxB08peQ
cPbVOMY1BwQWgsRT/sQ81JcLo7pRWKrZ1q7Sg2kbqdRwRitbe/znCfVV8iNXwbL8Tyl1m5yVEMlz
ExiLo6CADV4jHCSoj/Ruo1UF7abv2EnzR7uZQmPW8vnyqBfWYGTxszCsmbn6HxF7Q390prCTsRDv
Bc3k2Vvpq/1kbFrHSC9mr/1K51Y7jlhOx3li+MeUScX9f31cr/F652Y1P1X2Ze3gvtArXjjHpVfo
Yi5RKEW4e1cMyXVXMjaYBtp91vc7ges1mXEH40AcdTEsGwVLUfl7TsRtwcwtHsxQt0prRzFydp0O
LZ4n0TzUSJaVkH04DAVYlL8woCPrbvXW4qntiyXxMJ7zPFO02mRw6N9M/ZqbrXrwe6K6Mtyh1/9q
iwzUMDFMTDIdCd6BP96FddgfFZdLT9CYtOq8R2So70+PMA0Ytk+CBb8q1QFZssiNGXViXpdQJZP0
Ht/LXJ9xKzPY+pqDmhJqvy+vUdeqSFijUFqd9662QVEzrahlb5E9/kTSnJiAPCqehiLBfhqD6/Q0
GvX9lyrUNKvPpip9RMwS2gU3JkKZ1c7e842vGEMN6lXqR3xmika4tSHYBeRybuDp3nKHAfHjWfeq
+QKzUY9PsGDE9Wrsmk7h66o2mThY17xJ7WfXhHm3/92Aq8F84VLUlkQUZdkaCZqBvFToK9NzNJeP
xGucZbl2N6ACQ1ds5IrAdX2TD9yaqXTwPNDZ7ywsZcLywNO5ckNeVPyIWCPS1Vp+UyXNOs+138IX
WtK9/ugbb+iyrodm8Sm5W2YQIT59PrrJO+daj0NVxFGfBA+3mQrhXfqaFKI/z1ZwNKlDFhPuLW89
nOa6LaU+/FAz/xAXYxf7yorYlKIuExxVvGHqtRXGYsp/0rgQDlIuXGMGNvSDrJZU53MUbiSdCnHg
mAfvpumRXMSAQXNOlOEpOgD/KJGqn/ALy7OrSh13Bafh/vwt2qhAhTkTFLEtbNpNSql0GU9QGgR2
tWUp8TAinB1Jbs45xd/8k8nijFcRIjedAMCew4Uf3XdIxjovlP0NVmbRcOGtvn/EXzvdY5fFCT97
3pgUL74ylNquLZAVNp4Ht6pd6UK9dP/t2RDbQZfo4ChhlyllYniTWiD9W+qsLHFy/YN3PK15ymfV
LxRXTvYw11SJlU6kqQsvnQ==
`protect end_protected
