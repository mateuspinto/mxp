`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
RxVo7OJfWQaLKUAf98kuN+pd7z0ehDRMcC+101eqvbW+rBMsSNNtTm76iU5Nr8+b0akghRlieyVB
h0C+RqbtK5vpkPFcw25S9Ek+p04c2uoISdrg+9ZoPpAWB6CrEofDn/s5vHfKzc2w5onmg+5V9mEC
ILwR+BozV7bTvVcno/lMFDMMN1Rara7E1okdn5K5joZQ6MgqrXaw3O4DEcZFjTb6ppmEhV9hZeh2
X3oiaVoM9D8ADfb2IFdAa+f7FijzvnkmPHNb5Buj9OsUImizT9bX+5Ql9zdQlUYFoxpH08ARrGJO
iCnt/zcjcQODZ//rQnHw3kmMQaaF16XoR99MjA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="T7VEKJJCiesUNn36zEfH0AsdJJ60gagg4S+zX56Q0Y4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
bKEIjJm4RABBJRutrQlg437Tv9gle7dSNxmeecddTsEjq8UW+0TjQmhSyZaWmCtJXVFxXabl4vhn
9blgfv7dt+PMM0vQWBfU0tVX0o5sA4t5R7r7WpbBR1rWrrduxdXR965hAyLaNexvv5GX/lMRaK7b
1hTZVEnrRKS3WzFV28YcwPNKkWwix+DnbPAtGEu8M/koyQ7SocVCuCmxq+YBs5lrvSJSd/HSkFV9
gRfBQQolxKeCH6c/qTh1cbppHyS1oIUd4gGnlDBAUtDidPQbgKavnN48dj5AJ1k9obFtDLj+MZtx
nvkZp+5GcljyypGJPtbvkiBHn214ghJ/Cjv6eVe+l3P+ApHqJ5kPdv8NbJPIDpsOwEIia4EhzbDh
bC+xDv0TjA+bP4ZQr6dQbgnG2ha2yvG+Lp6CpsYgA104uzwxxnslMpw5UU8WvCm5nk6U9z5G+CKi
zHKWnrnQ5bVxZPNh4CBlRie7rvOuPKHuB/wnqNaZsGIzgRiNfRGsz9Wkrl94dSVQ0IMXH3FcpICz
LWxs3C4fw3ujgociZH2HzpPW420nSk+JI4VO6GZFzkXStgjUDPvp3yIzhTyWa7URVwnSEAiArfXM
UH0FM7xv9gYc4UnGC6ENPHjHUXvvB4KiOq6cbi/r7jWIZXAAirxPgeBPM5xUrggtJfK5Fzk86uTf
Oq5viIp1E6A4rN5MCVHrGtsDJxwGC1ElslXud3i5rkEPZjqlgBJRiXQuzqf8kj4UUmyfrmgdN8vo
xcPrj7p3e/8qBWJvUndpLIuXrWjhPPzkR5/TGbh31VjHK0s1LQld9Txbmvh32jUErIXl4kVqKu5s
5vGLLXddmO7N23h6wTgwIi3oumLgii9Y+0SFKKBIwRoZYA9B8VpPdteKXRQfTu4Zr4FGRJ7NkZZI
gqlsFQsmMEN2IiNsv9D5YBtft7it0c9sIxTI9Aoq+E9x5qKmjGEhuqnzt9M0yyZrGu/UgQQWuP8N
GAhyGbgEZDE0wBvvSD2JpmqK5MrfEKpiyB7qab6+AJvkKC1brbJr7mkRhaifW2UdCLJ9ZrIUP1Vj
irBTJZ9UZ66O/TiDpg5Q+sh4L3iwC2JyI2OgJo+fxlxq6wWFgZe5bJzCMC5khza3ir/WMylxDuRH
TfF+RQuZu2ARsTarq5O4PJeWPrPOLTvyOG8voaOtChAli3VdnHnkS1ftVqPD5YAjGagwKbsA0NNt
hCruFN/VMRYPeICsvhnjsxZCnfs27mXSMxv9yDmfxKx5Nm32mdfIaDtAQqOoI+/OQcX4i7zChBg1
KCOWhGeUsUVmaQ+KDuhoafUjQM0AllZngI6ORF+Mn9S+7AQbFrrjK00MkdOObmQ08rK4raP1zrCC
uur8YhUKJMmt+L9e/2fDYzRL6DEdoYCJ5C1JC8tNr9SK26eU2YpwJmBm9KVPS5Mdx2w9ROYWmq3T
ftMVSxfiVetYGwCTHYlU4GcBza5rZrW+R1tUxrEHz2gTuT80M4SqlW7qpBwwVhgEejwXd3k6BJ32
MV55oeTZTePdv1pDg7TSg6ApRI89W2ifKgyWlaA+CFHAcnnDDEiDB7Qkk0z9ySpM1yK/wyImv9Ag
FK2iGld+UgGfIV5LmdEQMpCEEIZBG9bzXrUL6EdJpChVZJr86huIcN/pD80bZ6dOJ+j8WwxirCG6
q11rRjklaDinEUV0KJJzVPKhXLGuUD7OGXUcUdXSJnaQQCVrPbh3KPRnByUY/ARh1q/TPEK3tz02
c7IUIqrApBz8wO+IEqxv2DbY/cy7BuP7OoXpy5NKCNET1CCG6y4f9nFQkGzoDIX+y2l8EnIq/FGM
rrenbobQNwDcCkkZFFO05UumKqCQVqdbDpPoHKTOn9ipJwLeQQu/1fXyq59v7Bpi0FUvL9o0RpI/
s+WtEU29Qbni1l0YgCU1UV834yS/UU5fvUCFnpF1lIznp3a7+gneNGgMFpuCs7omgdg5tMtPoIQB
svtdyAvnzeRXkfi+yRrqYgl5uxUcPMyMQlrtlW8PhYwI5hTtzHg6l9/FiW9o51LsL/ie7IHZRx8m
duMn3X9N7vby3WgTlcMwK1OsLDJNt7XAuQbo/CzYN9EqVf/XUBtxyTKHltKalTBxK4T6Lw4KpNJq
/IlFJJHpHLwrXIQYZqu+//yFXnKr9DR7SaU4IxlYSYsYzdo3mNyJM1aV5U3KeH5W051Doevi8AKZ
QPeD3i8uS7kq7JXhBjBPikuMC5ZdUU7obU2JAm9UjU7dG5fd3oa4p1bMEvw4rbcTrBaZxyaSYlru
5hlu5KOn8gjZqx0G4dLGRgauE3+aI1zNLytnQ05D6trM9q9G+iKGBzwmdf5HyfjyqYqzQgf91dz3
m0Zgma+nZeCTLTkp7RGcqTwpOm+GPoW+exqDTH7KpLl5wDBwGSWFDUt18sHoybLuJFKU2RkeI4Rb
bPupahVgkOfB1hs/LSFnmTJLBeYrHc62HFlI6QT3q4DAhSKKN/TM1w9gVss6liH3htj7Am7KOXsH
0ETlcrHvvUojtq5lg8r61O29qY2PIiaPn/ytrRObikH7JJ5ZfPe5t2t90TggP/rWegSQIjQJY1HN
ecOe8MsoFydRK8EbrQOlboHpc+p7EiwTu7hYLtujSyW5MD4LFfgjfcvXAbXHaSAaQKOkIbcXdD0x
SGZ4ljm15tlRnLUaOzk2qEuBykMOYj6bN957blVfyL2qstK+zvRRAjXwmTcUzNHpAu20l9PwWJml
mY7gwCX/O0pUYk9XMX9TUMk9HLaJI93LXlh0yzDLAP/CuD0cti0D8uVES1j6g+dkzFq1seGwC3CA
Q+P+NkQSk20641rZWSm8Z65qqRMmLwc8odYwJiDa9D2vLwEA9O4EByvu3ynej1/Lxx2Ju/v2mm1W
kJDHlniDM0bjqDOQy3tvrs+SyJ+a/L5IAv3h7yk+/TKnxC8jJvCJ/NW/+Ae6Ec6MnEbUwN3yEQLp
JOZG7DdPD0S15C6oJLdMorDPY9tnSLqoziU0aOTex4AKGdxoBi+CyKaUCrhXXM9/+ghsWIRSeh9Z
Hpx3oeAuTKBz4Y8ndDi4GwMZggYY9HmV16izRkiaHvWpdy08qX2T2dciQeS8tFyAr5eSIJpfq9zk
v89+dRanSRBgpuNzCWQwhQ9JSrMo5cMzA+S9WY/4I06Q+IQ/9GHIwTuTtx2Sct+Lu6QFTBzeQyX+
2DEpiYIzggbG58K2FQdcQx0TLnh1yVom1Un5P1yiLZtaiasLt/IBPU0nmUGxTlquipp2uGYA/EDi
5A1Q1TiCbzOCuz6tzZYqtX2HDOKT1q4GOnb4+9QiHmxTQlJhp7XtDcbtM6sN21HKPJsY4QG7Rjuu
OtCBmp2wIg4XGZ1g7lPkkhCpFPyZ3hBoDSvG4+1bXHR21481JJqoZPBUgmT9RVbxOcpCOsb9DutT
UmRbskhOLnWb4TQttHSk6hKfg5rsyXHEjOvbZseA6AogYgXvS2RdZKuCNCpY45u4qjiEMx87vPXx
0Eu5EmuSSQoMUgSC/iCn2dZjl7PO2IhDBcK/Tt/o4gb50ux/QN/idNrnBCgTYKPy6I4EGduL11xO
vJcaHBDwCftmePu5UZi3LTDUREEj1GrTlHEtImdSpo/07rNrNdacuTILZk4uBcSgOBpy4UDOe0IB
1nFRoqiF7sOtl0t2J54d7r5+KB9QIaUekgWztNbbFdceE1HU7YghgJhl34LCdieKeo0zdJHQtiNa
NKqjHInG9AxzhlDQN6pMHyc8s/TGRkXD0k8T8cSHauOs3J79176vdBpafL+O7VmO2vb7Nzt53IOa
J9w83X+uYaQDBK0tToLbYJO4lQqQnm4Z1yNAOSaMHuavKjsTs9AarB8+L6CBTjnGJOHzwVwxBEa9
a+bE5YIaSQ4fQnlA8q9H3CUAqEBaUNQPHlvO5fKCMHyJSkvaHq9Eveclt34mj4DwMseSEZtc9fo9
qmYtzRj8ZNbeWOcNQOu33eLvLd/rAtVj+jCog8p+fTlWvU/+b+hKGC0VkbRI8aCa6nNofYY8bKHy
dllDq0R2eD34O/PQSydGk7nauaicrQI/s1ZaDVtXNxp4OgQYvELcwXHnFpi4G0DfW/jsxxEvhY4F
Fm8OdeDonwbnAnOWV7ZT4RL1B6nJ2acsfZuAJdD5sZL/cyPrCRDsfNfm5knXY5bbTxxHirSK6TLC
VG/SIkuzyRggJ6q5Wf0lCzRNLedBYBUs1aoZi9eEtoenc+v0tc0l7bdCQFiGE9roR51g5zRcpQga
vHbUc0erFpRQwD0N/UtsB2EM/DYI8oOqNb9LMVAcBqun81kQuQwNqYms/+2XC4+a1ZOEwPG+79Nu
xkHa4DtZ1rxqO1YczHksuZ6tGV2hiAk11Nrwx+a+Vkh3X1+Eaw1jPjDJbk9UqzWC9iKxmSqnIDZ+
rYDprPbMKwwG1SmVrTpoiGFGFpSe18u1IIdOroX+/qI4XdyP3H8fWIcEtHDR6Fd+Fs7hUTYm31Yo
iu4G6eeNjoxEiaG5h5WpdBzUeVp7AglEEZZYZZ1iovWHshfpFUiBrAW37khBlQ3cuhIx+DNn8nmm
e1mIPBFjvzGWTB3vjSlTAB84zJi3MMrqXCDV6GQS1sKdavqNAIyYeixCwta3mVOiL4G6Nl1a55N6
SQH5vvhQWKeyz52cow8DT6s9dusYLmoaXCJF
`protect end_protected
