`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
29UEl0VH+HzloL9E6mPUfqpfs8deLvOdnc1gG3V6bulDUk2jypOvFqMA0vuUlR33aalfmn0aoFSD
629zWTAa0LWqDKq3UXRI9Ncwg/UdP3SN9OwFcAmmQABHQfvdqD38KKsS5bWg0CQB8omhmv2GEQkI
vUAJmJ7ooZNl1n2VDjfE5YH4O2H1dsmf4zu3vCLqerZmHZ6EsbLDlVWqVWVbishtc6bPyEpnXujd
LGBGWs4uBuZ91Xe+vbefnzErjBBeUMnnVkr7uEvnOohZg/teJ5RYHFdbJbeTGZ/Fw7cOv8ELypUH
cJOHKod3jzBMbeod9QfNP4+BDltbg0ZND4aKAcjWrxzyoYRK5Pd/oUXXTv+OVdwscyrIZAOKrKc8
DNWreGnHKE7wBnsjbbdrXCGEzctiljPsc/sQ5RpWg/WEycpTNwaLVe0lI6cHRNLDKWhaFDvQC1Er
JOw3SBX5ELc/pfRF7VDkk6B9xLfjeECupBAayKccnqldLvN6cyaWiwfAwpNNSpe4UOI55ceN0JMT
QcFMT9c3SdKo+754FAfTP1XDeYBUCFyfMvSpQAy2pcLDt/j6aF7YFfGNpMMYIvZWNbENJf+xHfv8
ig+P5XIzeozOBZ1ijbc2zqH/vIa4fbEj5aHCg96W1XX+pKfEn5XyRyFRzL8JL89olqopD7nRtFk1
MILFq6myV9tMeuPFmMxdft+2gyTqn66I+D3RIlF095ILxnveBYd+tPs8HNGgI16+4deiaortmqKA
jx5KgrMZT9SEO8nLzZYxNO3PIiD/EoJ4rwMedqNyHf02KqTuGjJ2Ew7fZEX62GWr3zmiXp9bl10e
K+112hpYhX0PE3PO9gGIntgF7JTSg3lwV6mEQNRKP9+8sCHRKvk2fHZOC3+7RXR50NEodMiLxvCz
r1Fiow5PrmPeYqRM/+OTIdNNXWj90cObCy53UxrPelNFjz/UOB8gsRj3RI+l0TvJosibJrtQy8mR
vGdkEz+rPhLHVyJqN2/4P8QqKQ4h5ThykGPubiq74WtGbjGgZ0f4sqHyN1xZMTsa4+luiGpw6xkL
PnospaiXA6ciQaIwiynEYFLKDkrXWjkBOkBFuMUJIRi59v36IQbzzuXNPBWnBxoZBXlss6cJVbAw
XDVy8a8bvLArF9AzjM49rcyFeuyN1TFgy5A86O2yIHWQxFaJ4mPdgRaRt1NmUdTexGfPd7icb4X1
kVyIdWZ4IImUAHeBBgbKk30Jw8zHd3/jQFVt0aGlagbPP9H93wfcmBF+isH0K5WzbwxWwnKmAf5X
w/ofawD1iZWw9Y3/MepMjnY8Tz0dinRMp0vj8LFjKw7g5paeb2tlahqL+J4abm8FPZsXlonKCzQC
AqGOb7yNqTCfEUHstbvBlJYrWsD6FcwzNgA8K7/NpeJMvdVbuPJ91nATUo8rih6Eq66oHyUl17Qq
EakCmf5R4pCHqhIosLFVDgw38QvKHJi7xefuuTE5tHiG7oVrs+t993xOAR9TlbM/yClGeCt4I8oB
kFVvDMP/nBktSvRQNK8CG8QhU481nEN6HahzB1mwJrhDKhkUXRN2/hgBGVlocgzAzQExSXMBrQLO
DNXjVO0KplpPh7s9u/FQXR/HukNJ01Q7H0ppw9g0G9O3Cx5ITQLMO2/AAANcr2iO+VPwmIeKU0l4
KVCbhfiMkgEc3017ggw8mkyA4V0ipg6oaVqEWR/jY1QKQ7j7VCXl0/9Ybk8b903oYQ17huTyvrln
+enfpI5c0WaSH4ox5xuYunrSE4Jv1/UjiItwLe+Fa7y3GRJdcjOmCkxDKUNQcUxZ0L3dueGYt6GD
qfyxDUp1rYGGBD01YuqFHJCA4XGL6hQ9iAFjC5CisC7NQbNpeN6gdCKC8G2oGkUfcro3Wa5Z7TGD
uRLtkQbnX5jjM5fRdbUNHsAWh6Tksi+S4Hys6q51/YTQJhB+H5ozXin8QxQKsL515pJMnJe2SmDG
sDymdF3apSOnFN/0ngNwBFvw/3qkSjDkwazIcWQPO4OjtIWoSWVyNJHkLIDKUrvA01BdCxCtdLWY
r3Ua6ojhEiXERGU8xjCLN8tSiwYTAVa1eel3weMme5grmsSMV8+KQJ3aqma0QAwRmhv/29sReOMI
e4gLj5Z1brmqxRwgVfyLMdQlga+s6nvplLlskv3iIPh2R6tMXDJq66BS6XICpzD1/mnBxnYWAjwA
Rsy4kMADB2Q5LF0qw5i1enkwk4DqkeV3P/xsNgpyKgi/PI+V8cV5fbk/2zt83w1yyOsuhxoRdpGO
EQxye+HBvExwJn7P17P3Aw8p1q7maDI+wAQk77W1k5zrqZtn9bBv0srVBVEhMME24rH5ycipfiPq
gYTZ5zgiWgQlAGvcAXiD+9E9dcvdvFOO0dpqyScbaX6aDMhxYIjltypWizlOXOMTQurYrgsVJwgD
ZFgTMzsPNDUtcfMyl7uSqhxUe6ZAIay1fLR5EC8pi3eRnLxgRkTtGZbuJeaIh2GShWBOrx3D62q1
Ajj4XBo1yOGqGv6gjggJzo/XEvSe7UDhdPitbzEM+jWzCRaW4mkIteQf2rt0GyqD9qNDeyH5SlX/
PFBr5a2Qhgz7PhbhtJ4JDwpk7Tv9pHhbut/MXBt6M2NzPBrcquTiEOYGpeEDyaCEtSjug3g4mq+g
1EP9oYFLnKz9pqxD1g+kWGvlKAGRApbnIJoSvZ9NfWwx4qntVsuRcjkgRvosQT5cgfEO4c/t8VhH
lD/olo7poItqpwgVp4wQGIGVS5syyY4stL/jI9TmS+LgiThpkwBy7tZyBJ392hnXP1s9nAHpO2HZ
QPmP250XVi6sEcLPfqB1y2vvKXw0zapOY4its6ao/0INpTS6SCkF/mcr5qRpVS5oBDyx0v48twAE
q2117q4Ny8YwwfS7wdN0q8n/UojTr4mZG2VnVmBcKoZhYyoScotfS9k8Y4i0HixU82BD/V0gKeoK
ux+0YoLOLqliBv+qMZIeeJwLEJEiW4t8C6TkIxaWyLr3Zvg6WU/NTYSatDVdk6zTddqMpY4FWhkT
HgAbm1ygVmGFVMGTBh+41rsV43CHFEusGEMP8bkjwlg9SYc0X4JMAe2u6QElKjJG+HzLklGfurrA
j6qHMUpoP3YNG4BHnSPpvUWqlodXCf1VrcbZSRmNt02EspGHg0YIYvIOyi/OADkBBys/XjPEvJ4f
c7HkGo0R5UbsMIgUDy2bCPokUjgONeAEPqiENHZ+SGeww2l+W8vlNty5Q6Q3sINyxAudYA7Owdgv
xyy8ZiwqT2HGkNYNlRdtKy3xuYFzsNkldUfc5jbl0cDeTzuoGBnTUtPXcQomhpzNw4KSf2qx3AU4
iP9f+nc+JW8OVEg1ItEHs3b0hMF54hlvnxFb35Qc7cT+JzMurHabMs09pRbiD2/CDgaR52FfN993
2BrEAFjKiu6qHfckV5hEU4s37LVZq6451B2rwu/mVSUUjNx5sUhWV4bVPZwoEasAGC/HAjgVHXGZ
tXr3f9YbWGT8EFPAF4NhQsjqlKi6meQ7KrHR2UecfbOdxnnixiJHtm9tB5j5kyjvp8vZ9+REYpb9
HKXZggtNI/nPifiV1wRcgOHcxSLOVelkO+9kfZKIbhv6VsJ8cB+oh1iy/3qGb0jYPopEFopqM5yq
Ibr6+500oTmaUM6i07305QoyQjHSWTMwjMcZCXKqrhBtoUJzqJ65piFhhCdD3pdZKQQeNQ+VwCwu
gA18iyV+VQU9OccSmG0IEFYHBdpDjJRrT2JMlTNCmudK0ufE+hdCWfWv8lGLidj9MEpoabh9oKfn
BRMhhK/FDu4mgw1wpDNJTX47u+wPrzIRfoqVi5onRQuBpF3sGL2KkYDon0mOCMtOTdeC0GXH8us0
TK3LRdBu59Qv7Lv8Jg9e8hJaVmLHoABzHuhuEcOsJeR2lHCDLcQe5kNPImuHq8qMSoH53zP9msap
hPAz2izrYgqxhZi9wPsUDS3rY3VYv6LSnU3nlWDQJoaeM4EH36Gy1u1q9Gx/a9CLO5KTNNxnD8iB
ecFs1Pr4j3yGYPVXfeob5GFRPey+r3MS6PlCmTJqGRZBOzXIXUghuLhHYJKqCW9Z9cltk+3oTWfG
0QD2F4DkON+31DpYdjloOMYu+VjwOu8DgD5BEN+wVyu60cAN8htEV2JWTSeJELYNjZx5rGLPfxct
FcRvlWhgTWb4Eox1QobZj37Ws1q40rxtdudT2GoF7fzhMfleADBbJhi0pdhR/GRjYrpJidtb1Hbs
8kFXZLo89sNdNcDBUS24Du/fRK4lwONhTJ2m8WKELCSaZacKxPbfsqA7EX7hleA5vKy5lRHH7j8f
F7cKSLCh1tNVQ3LL0AcaSxfnUukpMOIs5KHENwtJh5fDK5Pdr6Ls9ICYsOhikGQnyhzH+LaxHyzu
I4WiJENVe8ens470FNU9yuxBhuEHnwIddYBcV7GJV1yDz1v0rigjljzmCTihgY1aLEqE4SqFGgSt
c7IEdrrxAx3FX8PNdjrUMPd/PDtqPHsPfeEGWoMMqsLfowAMJ2oTLIrx9rn9T/4Dk9dZPnOAHXee
5Hd6geVGSBCHF4wXV3XqxvFP+V1vBigBkRtf27KBeiohN3QowQHvZpPHJauG5xBpISNYDSLuSV2w
G5FMXx1VSSKZ01U2xaw0efUC4vg8rl1aPnAo9nKM/6JsdOVmwgTPAIu2/kn+R7hVJVoKdems4FSS
j8GZc3paOsDf1fqQKGPmsa805JxLgdWJSIpOyP1NvPbKRr1720g3sTSxhMCw3QqMhc0NdrWtvi4c
j4aulvF4efewj8td61cTeYuOd23efe+Zh17mmzMc4G+bwvt4ii/Xi31KcPWPmlWtFvorxtsf+dt5
ZTqsEMaCXe/RuLS0nP0SIUKDI3vgqNyjPJv63d6HwY/ZVSbo4biQ3tBps3MScK+miPpGRn42/4wg
Qsazj7AOaPcHtwObt1lmxPqYADW4cdJi8rOT15UqqkykeJqNpCzielzJfMKVTx5YVh3AGFcMmpna
ebEnBjeWWy6oHCD0EhsiExn7lLDq05t+oS+O3+6HWECrFvdk2B2uD65Xb4Dt+Y7gLUQVoo3zoKlF
fkbQ+2y0EWIdOFs67bi+phoiLE0Dn6TkkP4rrl7vBEeU0AxPnU3wd4gwU/LrUwXzycRh7u5hZsTI
TD0VD4GD+WnMAl4jXfg1ihoyshNXePLaRH7LbrEe5QfEh7X501EFcIyHz0YlxCyUBfW1R2SxZaxu
1gXB1/OMroHqY01tkDcOz+NRDvjD7h5cg/ZfTWcR//xznm40L7bgn0+FR6ppsvReu8/IiXA8uB+b
h4ZY9OgBbFlNv3n66MMeb84Tx/UN4D2s1MfWqh0pauTKS0sz7OYxjDxauVQg9jRXFXjwAffXh8MU
0wF3YKNwrlM14Atzoj8GWqoJ5sjANrOWwr+BjTqQFBhkx0o9h1JZJhf6hQc6i630LyEo6+EofZZQ
tAS+0ZRbZa5FeM1vk04gmyrIoHJsSkBnf1F4N2V2jsts9KZsVB+4GlSx2p1PWxW1aakqZVuxOpUm
cnd0HSq1qb7iVND6IcHcxlIKFAdnsv09SRVK9GEqpN7Vx02imnnrOTJiPqdyRHXk8qvdHrOydu7/
+hFNI8BFN+7S68yIZqEBNhqNAcx8gX6b9/IPdMM7EgRMPHbeYqM7G6d3+lTYx7dq/RrIbA4Sz/6d
FBK1ZNd5ze40U1r6dfxFn/sAWDYKREFjDOELyTVxnFXhHPxhtgP8Uj4zSzhqbnzC5zh4mw3bMQf5
KjYRIJWpJsDI52wz3sCp3ThXsTMuW7e8Vcc19UOMFtbN+SzGDQeXAqqOkLR+PcuEmBMv6op3llBx
oMd/ZWMR/Ydi2TmIyx/9hxy7qwbaAdcIbbRtq0NVTpzVkG7zI93jKb+tsNH4latBnT5Ox9zUCLbU
kBoaUUYPt3kvu/aut+UvY41J8XfUWqMlNlcEOpbmuP1cb6J1/uHHtXJNf5y9p29WcR91ia1YaiE+
hnLdk/lV29BigtAioMHaoTe0/2F3V/WUzVMaYosU8w6rTEfZEaceUE0ksQQ7dMFDRxnzjAZN4CIF
cTU9Vk5Eex2GmzDBOn+i4/fchqS1pwTmUDK2q6Fl+utL8dOsFJPbhpqfTS0/yY8b9CHeKXZm2j6u
mOVjP4tnnulCTV/CRVRWnQM82Xpq22ugd4DR2gjH0SNjhQSc5/1nC16YMelnLBR+i+qTKTyt7j7u
gfsPxY3iT1oyb5O8J4WGe+Qy+UKqA9UV3E+Rrn/78XhMAJDgseZXMruXiQKA3BjaH136GmhA/+0k
C35oBULP4cYwf+fEVfNgmA8542J1wmAh5wefHF6clyTTOyZvanUaPSvxazaTJsEFO26+TjRdiuOg
NUIcq0lea8He5ZRZcybn4mepUU+LuLN4usBkx3W3lDTgOhvv9UeOvZqbjpv8roOtq9upBWCVopZ0
un8dey0RfNTxvPFjiEm0ba7kqigHjgyBlRku3kLfuvOJOG2lTk2qvTKlc/aq/MwU4fs2xKWF0unC
MigGnCiMFCQleF7VKS0HowNPkgsyZtqyQ04ITXX4/86Zch9i8+AwOoBHIN2+zcHcqNgGCG6dqDjr
JJnZb7eufjBCNVZwAInt+U1yxu1yqQlLBCrWRnRfGYzDlrh/QobSy+aNFWCcpoX3UpJAgAETuTN6
2pNcgEzpEtWdxDujUWQfqPA1slfM470iPXbQae/P5Ib9VP4f2ICa7myXywuuKzE+ZHJ1KtMF2e1Z
xsv8rIHwj2snChaJ0DZ3PlXEVD3sxCRTIUvhe16UwdcHq0uyxd9yEVZSRmkkuvcPmz/VNVO0X8NB
Il6kaKE4vTWlTNgzM3kFKhB2XETNWCKbBas/cBpESDQ3Al/HN9bmp3AZbfz38X1C60I3sfFFnHXx
/dEsFoQwqlizQeX19+pqwaCnnG1lRdQq4Zh4cvRG8SBIn8SKzIacqbTJEWSpkNB78wDb5G5+S3wF
GHlKquaUQE/2HRjZ2c+GLEgfZpDNdoLSP2Olc3GzZtkzCiwunms0P76dOtRNDMefmiRsmMyiJUAw
+dJsGIdZRQVl7/Al1LOZ9H32V48hfDovo0p3GWCvfVFjpxuxHygcjyF1NhPcGQfMOPleqgb0g/wu
4Bhj7O3ZQ3W5WRyJYe/9s54c5Yv4O2KCRXrg1kbRgxsVbPK9fo4kX+z4jxOoS8cr0vylU4+Ee7+O
BrRySgboP7AWDkqECECC3uY935sWAB4c8j2gFJrO8qjfTAntRm+kDdF7ZxVXyIzS1l52tYkpG5F+
ZavGouh0Ng8aAIl4VvwEaCmb7NB7bUnmhfNY5+xfwY3UOaCENrxjmP0DZy8QxGGXhZyhztCFVoxG
ptC9QKfQ3DmsrQC6jk66CFnS6R1c1Zg7xJ+o5WzzTbuG5l+Xpf2AvJf5RgAP5b0XfolM3/5Ep1vB
ka+vcBuVFmNPBnY+ZZ39+o4/lnWq2c3SS2ID9q79UQmcGIvt0Z17pm1bnHlL/9omJ6q9lEue54+9
ZHwOylmdAKof9OBamycPOJ3rTXkqkO1MlqTtisxfw2cQSin0n9HVWnOaEOH/5VZmrmA6gJkiaGhO
GoTxCiBgRC0ZE6E1/lthh44NW3Tz2avGll61a9XXwjMq8k07kEnRLQI2zvh+c6mza1sOwv4GkuFd
XLDUFOp7dUfl7Jp6ZE2JnTDZ9BXb6YigDlu7ERn/f769hyekWhUX2GAHqPHVKVxzac5iWlQxnCe/
2vkdeoCBIOezsgh8v7qrII+1iNbbUBWqrTTAJlxTqMqowv1ko8Snv6jwtxeTqGckMw3nxEOeZ8LP
V+9s/AWeyKxKPiu5mhf8ZcXGNpIKK3DXiP6KwplJW1FXg10MCEnMXPnTTqjvT0JKz58xCxmh+ids
QHOoMBTYLg+NodkEfBAQOdkpiGdZ2QI/BOkLQgHUbnUa7Cs7mVVGc1lq0dA7NZlRaqJ/rDuIqOyI
GlEsRQaFZ+j7Jubl+bgSYWya3x+xQ0ij0w/t1rZzIFEvwDNazmrp+jhYBMvaQqykppkdl+xuBA63
2ELzB4gWXE+DDy4KbIduzBYspyBYHUrQ4qU5HQgchi+FFutwINznjX434E0eCdDSjqqAE3eNuS04
Aq9QhVJ4m+/u2QY3LXOw8kJjDRte9CNzo/ir29HXXR+Y/OOWn9RMvthwC+rRVaiV6SSahQWv8h+X
y85bBROwEUdl66Nh+kakJ0OcUW1FrhzM1fkO+UhS8AIL4npyGj1R7KyulIHaoSTl8SQj4ynVSnxT
L7naiOGHVvY4JvxIQRVwHA/6QiO8ZEt+4/OyFca92ku5csZitzstLdi1ebipKn5QTwmLfGpdH82C
ArBhi/h6JttPY7TPv5bKFKtZ93sxzcjYP1jqPiHLUbftyMVu9nJ1f4dO9+LSXBAKFwntpMUQObKb
rYyIWQCg0oWeQal6aU2UWBRWJeLpdmXi2PX8gMQpDzdiKMI8lrVxVAdviDfD1rSxfhDk91Y5w3gT
JZ+2+HuY/BwZIoGFWJ3zoCbIEdClsc7UtmAjmkcxjfZzdnwpRtYpZBVTxUY3sYBz4N+pSmy2tZBL
hdToMQCNlzsw2srSPTZAbM2LBp/bLul2kEPHbiy5dVqMe0h7yjLxZ+zPeUSthggd8H85FTZLY4Po
ahoag6G2orKG36FCgOcnxwJPzwIgtbwm4SU6wMC60niDFMej5TglV/yKG/LcDtc36M0dPeo5KLaq
2cN/YGNXa+fN3R+YH7j1JQqO8ShM7HLOq702eoZCqjaveal5BoLfWdJwI8KTRtNuiOHhNZTZUP+H
puerwdIrrUqVfs4wxjnr6Tfm3c/nhpFZGU20uuD0qF3Lv1F1RBP7KQvhuYgqNshxcnmwlc/qldIp
92QO028q99O63MhlJCWplPGmc7aPnrBkpOswPBdpqw0gDU/oycbRwnDmNME8TRUZIPiYKBNim/hx
xECanrX1vxA4xTGvwiulEDL0qBk0likmD63cCyAZEgLdSD1I/nB/KVgdZAbXO1QsodllrvHYtccq
KpE9mTyyXpy6ax8M7wdHW+h/5pY9VX+WXvAIBCxj1GUrOcLmBMDlESPqIGc4ifa9XR8Brs/8iPyi
EACCs8/iDCbwQyTngxRRLoa+ErIKlDu4NAy92MGI4q0/LVgA6kIt1EJiGwSEtLClPlVHOWuuIZ/s
76+TV6xwqTWn/lsMwLtUbJ1bZByq89Sz6yZODblYy/Z/viLt5s1d8mH6tTx40Ls4rNlP+CDlnk7v
kADMvl4NoXzlkInyuw0poYmxuCcjZKHnMLosDTD4sTdwqMYbt343ejXfMpwst+msfOt63EHmASUy
rt5DLpyNMLuBsqSnabd9wsbbYVvq3kKklu8cjUywxitvTCdhX2CnbFws037HYiYiu1eSCiuNNBHO
U1ucdYmBNzB5ONniQgufQhILAhIakUZmAg3l4OSNpk0HifucYHmWvtD1gEnRkoL1iQBbBdWxqjiy
p7XKnYGDiqYvdP/8Byr4H2jCKOGxs7JJD5Dp3wsayMxgb7NH6OsnXlobPci7jaH8DNoJ+JDgyvml
ycz7sy1Ga9Iy7cxWLn7+y6hsH9TUqv97HsaK/c0f02DRH84u8Tzxh1hJvsoQ13pY2SKiBEGVvrBo
jrr6/q8I2Bs9ZW/XTewQKqeO8MGbiInvX0aTBDTtxbYN3oeEFdv4fiXtflhEJ24lIalMiTmNcJFY
EvWQqGuzJHqEE1khYbuJ4Qp2xSmNygDtzCHhjgsnZvu/e8+XKGrc55dVyWNMABcjPsT8WEeEltJV
duB2FTS1tieU35a3ZgXMGybRdcGgtbLbcj3RvlrT2lAN1FXZYOeP+9+690NuHQtTJwo8s2SxHM5y
Raph12yjJ+XpMU5fkMEgEwx57Ns3O7+kFzFMshKm8IpwpkxIPxB8JgOJa9psxGXHCir+SHa9iudu
zJWSU3PlbwrzZgX4dWjrPTFzfIOenC1hF0VQk8guGKCqske44ViMlyuj2UFuiHe3puA7LSd8Fat0
53DsYxyXpeT2eAfPmkCsVQ+nEVIKxUm4DcYh57WExYxVgEFTHkDfpYoJN72GD1fcUKev6gg7445g
m4PKS4kuUQ63U0CQN4Z2q/oe8TAFvScH/Myxkuq+jT5aNPDGrdqRrE6ABmoZhK1Vv7qx+Pp0v8wG
HHrr7HTizXGv4y61/6qvJAA/7vauhNY18Uc5O3v6Eh7iuP5QV2+LTeGr5sBo2tI+Xp21MfLxv8l3
GBgrafq2rdknmt4Cbch0OXd+5Jox0P2+DhYuZX/3lgOOSwCRc8jRg6frDs34KJds6hARli8M+7wT
bT+c4xt5tFJg6SHieBNZbavZu6FWVst8giuRoid5uVC4wfGii2GGD980jUoeeynwM5o+V0Y1AAHz
J8ygyHI2lL0Dc/cJlVHqGj47WaX5LgRyfxUORlMY8A6HSsbMDaYKCHmxfUuysr4POWlIketmuShF
sp+uI4nO+NC+bjMFrfA2paUOoPMb3H1R1s+SOVtkxZRVzDGi1Fvxm24L3STCbNTpA0nR8XIp6xYR
E3kUBsSV8X1NMqM8q1yDrPxios/SqLdJztfWos+xZsuS/iKjlj7HMLIkt+CMQYgh4WSOst6MScgF
3cTcHU4tv9sj5P+ZNKGKH9W4ttE/MSTtQSwmBH/guybJ1zsXYhGMOuzTXvw1wBctOljo2fbi1wiT
bWuFP3msoWIFTnEu1zYj3chynWX8G1e2x9hZxUTJfvRf+uZlfyErA94Ab5GeHof23iNT4ufN4fAt
D/yKhP5Lj286rbkbzJhfPz+AN/n/y6DLPShDPWduIIw3tpec2sbDYrutJ6eZtkfU0qGiRpEGUqly
7sSObZ8FlV2kndlu1ozJF8zJZWkjAnl6NbLDEmyboXd4sVRSLDQ9WhWiFFnmSX2baoWfq4XUXi0U
4a/KEmZO6qaKTmxn2JWd39+B/0QLgr8x7VzXxa8Nb6oJ/FAA4tX2Zweq2cvoR57NQ6xJbICu94DP
i99f30GT0tXfSLb6ITuGcKbP9OXkwRNGfH0ZP33MHv5VnCVUEM5voUuxXlyiqF+qTADl9HMezK2r
sjSRjO1VjwbTQdGNygXXAt3/7vRGjcTYIvzZhh7elfLIPsMSiH7PAIIWOn9BD0CG8Ypim+10cjfm
Mvpf2iOnDCiJRRAXzMBsb4/TbhkDQ76bLpDe8DPN/fypJkRdhY9svDdDzuiquRB+LHCnB7CeFQCG
Oqvu3753S4CuLup2rIniUx3AIDY6DMXYZMdJ4kwrthziK0gzX0NKlciSuv3Q7kgAMH0BUKnXTabB
ysC0o9p1/zO6gNHVQN+ZE7rppyVAXwxHTRtXukhz6gxSIPA/G3bDyWbSgHkNLrIRaNwjElkHKE2V
OfUQCfe/hfLgHohrYFpc8TeC3iZWR4gDnJFwsghJacSdlxNFhMbuk1HtvfRYtC7JgRbkcHirooeE
yT4PBzFxbAtXmTg4U5xMt3TXAJS3hcX6NRACiO1QkgrlGWngwSSm+5iGZD2zdgPeFDVKfzYYz6Mb
f2VUs1Tczx2L15n/i9rT34khPwQDak+qoZw+on/2gwEe5QeWmxss8Pc3kNTgkl2+8VcGp+zeAyZP
rFLLbH8iyDX8pYOOre+as0tSgKl6iOhsd/616fSu1/kbP2YtM2T/nog/FbLu32d/XclKgthOPGBa
zLf3JlZrDRKi/DGrAiJbiBWWMjksNvOiV67yW70vnsqSxC3uuWWHigJAuOiVxlFzr5KfqtiGlcgE
NKNmQO+1JMiDvwTt2nSIbw05gzwEMC+IqmZYjTDsa4llRNu/3Ja9UxuGkyiCER7HFx9VkdjQEfdQ
v8HoIK1LXZuDNe1QlE80dbB7w4TCMFbwfG6gYN5/Rv6A9VxAYosBnnxgNblGIjoAZZ9U5ERfI8D7
rx5EXVR0lLRqmEZuTE5s2FH5rkXwvBbogH/u3XqlPRbrsshU18U3IxqS6Qifd59I+WP4mJjcZ7Ee
+ZtKTri5icBSRWv8ITGz8SEdhl8AGKQSkIQg4/EsSUZjSdZYXwK2PBy3ElusscbOtFTzPKFujfjE
7A788tqVKj4zOFlFtqm6Tp/jj6hc43B12tE8lNUJPJQJwx3wYsX2KBkDrbZ81vUglegqn9G4Mzsm
UE37K0siODLb/Vt6gvgUkBmQ4UU/WNVK199TQUwsGJc=
`protect end_protected
