`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
hkBknfs2vwddoP/Qe1qxL+xwUJYjLRlvDXmvo0xfAK2fwvYiK6ftyayNrhKEwQTQl/u3GUNlzpAm
kCx8EOvK5ObbXm+OYgtG3Su5KMJ9xujIuREVDQs01JGW0MsilqEP4Xk+/mX2/MzEuvXhnUQBw3Rn
uxOCcibokezyAx+/pGtiP50U8t9wO5tbNlHNbcKVnn/usXl0y51FZ4isWbI+asrbhChTOUmdDAY6
iBbfS+jCRqKP6YaoCWMEVyDSsk+KGVCqqys/6U/bwVVfN1WRZaco+/9JJ2Wfk37546MUIjgixgbm
uJggly0bNHq4/DXR4xmnTQEBSDPw/6i8WjSL+Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="3UbguDgv+6HHA/Mk8aqIbuElqnE0U0hsuEWhgQfAttU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13808)
`protect data_block
ueBgSw977I2Yj2xL0T66zGfZaWeIienPw4xkvH+rlR3f9AymFJYrxfu9Crrti8HoQv0P2quvEHUW
7kR/9CUqodnWjXF++2KG/X1GoOaay+kgS0D23eEWu7jl8TLBMB6OTg3WjI5ec3waMgsWOKsQ/YJw
abCKi4N/aQDcBGWUQy/SwnARCkTwmEqpyzq0sXKCCRBnRxMm/mRuj7v/YwTK1euiI/igXQ3I58mQ
4mfsZIfK82WwdzIcCEwg7lbNOumDmOLReXawoUsuaa7a4igUNgek96iGe5gZCfmqLiK8HfxDOram
9qud9rAxCwVat/7fbLkRNDMW01mE7GE9ebuaML4645aO3AaJrBdptx9+lJrW3J30m8+7VDRzvcJs
RyBsHVVPeEYqXTA0YpAhuEnkqT/MP6FSXQtJF0SzNs68DS1hf0Ha0LOAWM37Hg17GY6z9KfG4dXv
pe8sQ4urkjGRYFdAHHr+CmIRFR1+UEGzPQWAs4f08RZFRBRJtDK2HhPMyQwztTxeNyKKCpB58SDq
phch4WPOBUfCDtnYwYEi2S/ye4KXEfhxUdZHVwRtxRcjQkCgYvnorm+QqNakhu0/CzR40c4oJERB
0EKmUGakpyoT9+8ZRAynrOPoE4/eeNG4ZJH9IWz/JggBzmpnx+ELW7Zfk+xaZ0vx1yIQw22DyUfc
wB1Zy21O28D9zYLQVXYCJIPFpwbYI/V3Ztdv8GIywHYm1Hn+LKSflpOldCjWqwadGlbKlt1ayA2T
fTOpi6dnTRXHU+gBTPh8jXr2VuqjQC6EyNub2s23zwXMZF88hMRepXhqyKPCFKCuyr08PTxGmy9G
mTh7rxoGAfM6XQ1UuZvTTHvYV2ljvem1bMfeRZFcK9EUOuZdAH/UJeeXAbpb2wN54h+EBv1079WZ
0fzcR7LqwM5t/VE7wsqit71O2U5Q50fTHnpRurbU0BMTKKeE/2WpzDmjLS/gfRGph2gbAIC0nkx4
9dyBBYxl+Cemdlbw2KopmwWjw2tKsSUuy2szez9VdEkY8bQijM/My2hhn7npBXVNUihgHqHNjcaQ
rE/65BORz3FxfZcdg5VGYbiQHRlxZozOHPENhh+KLi/a+nklfqE4F2PgMgLm8Ef4Sb1pecBW4yFo
/O7OOo/1sbbeYIUC7iLAsQh7h8zZDpRzmYH5ITuVa8IzypAJz+RWJiPZBqsp9y/ylwGMHP+HT6AL
NIPrb43tQLe+utkMEKlRKloqrbIy6k4FmruNidfSKalpvz428cHxcNOUYClqe5XILkYBMGeg596b
mxQeDVcrjImAkKeqSCbMMTIgq9zIWL2hRtlTGfQnFqdeymnLxCtcTkSAzFqDoK/y67RYTblnqV+O
l9x9x74InPvj7hFS2JOiQZcjeEZlHxlJLzQA6drgpdV1kDyu79G68ydXlVyj/EfAtK08zRjSGPvZ
NUNN2NMN2WopJNAsLgOVD4HVtVm9IWN+dtvk3oWyO2ne6qU+BZVvCjwT7ibmBKzc5NAXbiwDZ2nd
H+KdGPlLBhHFFnU7AMqXxI8/F/Q0MBdmNubw0MzsFoAWfHwgu4p0WMNPxOYcwA6v807corhnl5xz
zQ7q5VLFwKe8rV75C0n2ovOeXDULh5aoeLiFHU/XXcm4YN9FsEZixR/ha5iHlfJUENxP7ufg/E5c
mlzYCF9KsTknjENQ6LYGcv7FD6+YXArMj0G+80qpnI8df3NSX5+5D36IzjL9mHtp+4e8Qc5SyqEf
aNPZ4aRc12v3LiTKZNqpvrBjQGdxgk7udXP8aXbFKgbHSaGi5mD/Emp/A8hBenGrCBtudlxk81jF
EC1i3hQzLokSRqt86Sc5+gQ4D11P2hI6pGNiy2q6baaHT+GloPMKL7yBINOzuoQa8GblSwBN7Iuo
UZy7Qd+wXSLMoTqsx6wfRBIZ4ICXPsGoiIWoT9KuIbxaS4rfODxf5iiUNL85ohqzgckhCLAKwgLe
VmltP78qZ/dLON9d1A0WzsvIyqLLG6DRXaQV4n9MlWEnld0eBL9SBstEQY7DnkxoRtNEoetng5u7
IDASUMKsl6oPedlklDJsDE8D2Fo9ueRLZUmNGsvfGIbQeFAIGUU0zF/Xd/beiIg3INvSPlt8OB3G
0K6a9F7gFLFiL1OZjfdZwrqSfBBxw2jLWkyZ5R1dNzJ21/AmMf8ksv4S72lT8dY0M9O66TUZGYac
GzeIJ7TsVOcwm3ukQv5uRsytP1gXVuvqqAWZ+Wj2VkPKzqg10tgT9U/4vnJ5nmZJNclmuyx4d0ky
+YCd0kTezM5P6uBcCQAYFP06e8J5P4nKMizDp+x4voWc237gEripL0PscGJZDfNDIlzDTJ0v73rt
cYiCuDiRd0EGQy9QyM8PKfWpDNdQUm1xVqf9yfvyJnnonGFDkbfvUzhu1mJGVvUo3FF2VZTFlEmq
wtz3SGSDiERMWC8JxQ7X7s/aie0tq+etdDJ8J7rCEdhjJIslzaUA9Sb+a8pg3YJCl3W0SxuCLftI
Kzm2HBSW257xMA0DWj2liAQrlbyMUW0T5An7/HKmx2cb39OR9aQrdsYWWGho4xHhFgPLY0/PvaN2
hGr80az4eD8EQKMchJsqpA3t1kj10siOq+EM8rCiUZOqGe3o8Uzj4tSAaVOrXKVzeIpmKmPpuubv
/8CcDyAhkg55fReNG1NJ9wwhrW2gU7L4uFmGh2dIHG2nRunVgybT1rIu3vJC3A903x4aKR6JdiSw
HdIo3qfRDLOZd3taXo0fCdIW59qj8B/93Pv27JcFLX512PFBbEoBNPnkUoM4Eras37gz9fzNfN2W
/fOCKErIjWqkIdgzvXcPyG4+y2qC3WOmJUUQLdlgXQCZ3eiR1RnhaZZtXAxUjuIZc7DIHjklXjsb
KHVffBVJ8Cwk1V1zeaFxoOExP6jMh9pESHjsfYXvcOcnBqkK8rMVlvo8Qr5P0LlNxgEGP+E+cuwu
uk8uHrX/YYIHOk34ZgPA34ke31iaLK7KvUFP7L6ndqwXcKkph19/39Mv2hSroAzknJSy5M8IMiwH
ebcO8KNtHcvQwjsTXvLGbNcJxmKseOcFfwFhgqfXm40tgDg9XnjUfT7z3Q/q6np6+Ewl1FTg0u57
vLsLFi2EUj1u+FS1+svTgBiN1rNhFSpiC96ax16CAeYTtc39QBOQ5YV70uW3SISqayXC31qi2TZ4
TfyRsxrb9Deb0tSzmsQtUAMs1bgFOsJHtYQry0g9Rkl9xXjdxMIWHwXGOckzREqjsOYIFTKJg8fs
UB2isWCgO7DgqnKKfMPthMGxgmo3yF0jRh4NTY7jSowSh9itHIf9optAE+9nHhdMTpoLUF1d85tL
pj5As+0H7v2OBjdrioZZGEd83L54A/dmhrYsEHs+xjxtsXilbzUriWA72gzsPM4hkTdq2aZ31kjw
CizhIIFC7z2SSiGwNgnp9tWIFStVE64mB1TChv5d4zDMXGezhRok2YnOlQCML6l+XTYEEolMyPLK
nEpFHQ23TNL/aGT60q3wVI5W591kW4CVIjFjoqIgXK0qCN6If61KcXKi1hf7BUMyA72NA/agmQCd
CTWWeoaCYxMYVttLusLrXC51WG1cVTeBUQttNHgB9dcm9poNWj0pVIP6kpw8BUvqHuPj8JIcwKjR
NeLPLMpIluDfqVEB3D9eRfMYiBtrYelWntTVxpdHIekCbA1JvN/QDLv5rblbIIHjnVjsDFHHUSBH
T4xBGTbKh5YMjzj4NwXbKm9rvbbguafeG7LyR9QH3EspshYxP8dZbejGoUFEMsf1kmk21/z2zWt7
jtTxICYgWb0u0kprJkP648mgobqxEKsyoEw1X6xcEHN296qBFSDMluX5ho5s/Bqa+LE5Hc5IMZGQ
vyALfLpoQrsUEPWx2v0fwjy/Fd5La7azqtj7Up3WcK9Sqf1q+oga32RNv5dY2YnaB5CGYMy1EUSi
WY9HPxT01XTXestsRdGLGDs5pQTEON/uQ0QX/TNIHfw6raVvggrJLjvbDRAJX3SF2Yk6tEMF/tCg
f5P+e0J59F0DAuZA+jd1p1AabvCi7pEZBUNMyjUOcI/Jg6O8Q4tCnWxuotIR53424/TTmsHUwxeS
2PFXt02oTRaNKakGBM62yiFaQFPvDhEnppVfvn77Cu9+1kO9DEo5HRANUh0HdEGiKmkh/+m0hh46
+367qxV+ueLTVkV1bZ0Yf9evV5qM8VSvQ7JSPkBqZhYz2MzQlZmvhQNh6r5NtaynIjcruQxg8luR
Zq8mj2g+5lORid65u4Ktqdc+JcqxS4sJzHUJBYbx/x9jCZa+OeEYTNk+jjwDeOLZw4te0eO9OrEN
ehkQ3DluvGwphCqnZWgkUfRN4LdOIxc65jlYQNxKLqSRkzbkXzHIFKIPJndum+ahd7tgs/STVe6v
7SnR5VRuydj7WBisqbd23caKyWQTMXWvQcDd3atYy2pxZOFZEtibySpt+OC9kluoHEny0DL8vD9X
Bgj9IbN9B/+a4WOSmJ6UJ85mtN03VkdyxyG6ydjDgviH4qh4DOGEATRLZ3Rb2qW9zVIHFkLqSZRg
gmQXQMtNgTmnr5KGFQPJWQ3/Zr3qDSqyKNL03RVcpTMBRSuouIgkKFL06uBDKhPJ0spGk82jJ60m
0IIkMPB1H+CdCdpT/rwHXa4n0YK9HzprS5vlO3F0tBYDDqR+kNxNm2jyfoVofKwsu9d4R3ZoBogN
e3RnFqBKZQTRRwT1N4A8JAVfeHR5W3gTBLrSZXj0RuxD1uITKo7VJaor5PsNzj/AlOC85pl3ovdu
EgjTZlN/A3k6dsWA33KQtAVUXQaK55kpBSXPaUJT2arpV4lDptyuaR3GovTym1kh+eJPgbi5RRZJ
p4DYvCh8caUTkkP8AFiMB4tvMCbb0y0cvl4J9moRhQS7ZdP97dvcPD/9Y8gS3xvdohXG/K85liMi
iVhHyjQ2kHkWkZmqQS4WbirWEyPJFVWR829M6aUYmVbcHf3pZhsVjb7OHnBHj8iaRuLrYHg32emD
tYWp6TVEgiN6YeQ2oCvuX2G5W5OuZqruPE9yCRC6o7WzqJEsIXdGLZQ89fG1gHiJDUetuqe2+0nH
7DSDb1kVh9PSr2YqQP6D/wzprP62tDPKDfID/+T6vnkAj60bZXNcvxHA5wMbhQzQjPbWQ3z62eSS
gAa+Ol6+u95L6rbUq8M/GAG+IELqY7FTAHpyleUVwjGsld85rvq40x6BYwguzw85LarxbMw2IMOE
aaELRFj0McMyiPCnf59KEza5Jf8YKH//1PLfyjHIWCTF59l6cm/NK/hqoyBOcxNzh3Vahnmym2m0
8xFVmIHZ8DO8ViZVNZx8AdXEtYuUngDC/1WyKJzWxWUB3w7VegXHvgXbWoaiHRt/TCqm2/ztQOLp
BkHyCZSIg5KrxEjV1zneO6qODsgxqpqTi0IAO/+2OdlGZmOxThc0n1mrOs8W+WvFu/tGiFn9a8Uv
DtvZyDaFKTDfXs/dMywT0ROGcrWpBlmoBZmLMxRZ7SeGKJaYD6B8KI+87xMiGQP7ZlIa1QSz8GEL
iiG3W6M0Y5zdhP02nlHw+tnKeK5QKT9t5F1dU+rpKhkoJqzN4JEU8mj9nnTdTE3zLnoCRHPZqUkZ
QJDdx4SNCaNzgrMGaclW7q9D+/ruV6A/oL/uyIQTmuAEyZdq3jfV5HXh6CGH+rqGBz01T/Ds0Gp0
P5hIDCCf7O8e0uBXGzLcgisNvr5o2MGZT7cQQVfJWCfvRUJWYl6+EkZhrwh1zrI+fl2A69aUTxzk
vhUVAUAfBSAIwAsMGFeXSrEsDfrT1BjqGMQohk1+lPHP39DBQ/nmkH7+u2NJ1RAOgNJt85c2FS6e
DtV2Difoe9P9YV5SpX4ruUxZNHY+tVH55R83yAMUn0D1sEaOonsm2hFKVCCbNAa1cCKy3XPW6Aro
C0Q0EUB4rq8V1U1WNkO8c9aAVOCWtDc+UyZlhrmD/HER880fxh2jU3Feh7q46UnmV1iTV1qp2Pd+
7Po41cmiNzjakTWZ4mO2JeFgJ7f8147Y7vTO2nQ7r2T8VejBWPtKv9H0Nbfcp6bOuyGPIXtDwjfK
MR5fE+XjfplvJGlj8Pe+eRRzcmgLyQ9pJi144gHQiaK1G6RFDhENSaSWhoQMlawJm5FLl4ASc+iL
fUcGz5MwRhZyP5L6mjFPV45D33Bp5KIwDdIP5i9fhLptGG5qErOL9kOg2gw/9Ewlno88lz2EJ76v
SEiD6Z7bJ32tWFNXBfoaIOPDusCpimeOGnMoGURDzXpAxZAa9xFEWSxr7Gn87moEJDHuNS5a4286
HV7M6psURhslPOkluYwFa+HuLrCQfVdEjTwKP/GOzR6g0ZnCMZf7BE3MlxfAWS6dfVCoMdpcjSj8
gdgUe6+Lo6buAwa+fFxledGpAXYwOnQ2lIr2FJypjSGTAW1hC8vpH1YyX+/OGuFvMQ7FecxxmKxU
pdxf1MDnxfoaxZTxxWawT9sClDigFI7EOu3TY/6boj4QOWua3LCHcMeqqZT7BauWYVS5HKeyI1I9
ilclfAarxmuu+/LvGyy52671KgNlxQ0LXQotSoAn3tMYE4g83kQZLO85o7DcOKBcmkBP7MZs7tpg
yPo1poihV21N//hJBYy8Qx9KiTOPu58hyNiXOdCbMWAuiwbGX04LAf+Q4i8o/XMS2gdt1ZHFm1Nv
7tMMscgTjH7mzgwBRsDVc3tT5aKt8LTpEVqxCZGiC872EqP6iAcIFePjf0rYjg+dy4QaE3ZLeVB+
0OWVl3xDPppPghaIuLDnnK0hAnkM1Fv+7W8cKcmxKVDSiQFZAuoV/aTOPwX+62jU22TEnrRolC6w
XdeIbA+m7I+ATAWqEX53KcxVYINCa+RLQ86+bR28o3DBs1d8+70d2yh5IyP/NmhHIvzOdwyyZHkM
oRRhOiLh3HjN3lPz+WL34JSWIkAbmYc+rrBGS43Ot9teO4SNHsoTA+aD+Yj1hdYo/192TIcU0TpP
bHtUdLv4Lh5o8Z3Kt0T4VrzFgp0rBqEUUAeOen4p0J6cs9Zf2E6Js014NOKZKdKuS2FS0QmsSIml
58wkhrRPxREUDAUjVyBGpwfswRij+PnNPR86PopspODGhs2/kzDrepyG777ZYOIIpUOMRZDpFKz+
AF5xi7MOos8lyjzAkbnJAlhfLJQfQWPtM8etWBqumQsXTCa0gbYVFD3jXQBmq87E1LWImSBB/Cs9
RbnmkzyIUCtKQI7dJv0XHRbIm+TAJ+INIMHl3J4hsrgMV/PCzieBerkCm+PgXSP+BesxTgfseO9B
fiyT035uKS7eK17c7bBnTW+Kw1a8ssFgoaS9NabDe3o1PD5SwplWoZk72WEnBJk7uF22+6teoADk
7ubh+AWfr86AbcqdQisKcOPfZmxwgTdxeQoNslnKiGBjhJaBIyr0qpXZEs8zrtXkRxveiR2Rsi9c
XhUEsVcmZVltdKcgGRvQDF+JYed/Dxcr9o1qTJBi+2hopwEDNWs5gHlyC6efNbzg63sHAS2e9hPf
ybX2qv+7rGrmbbh8RxPk8jF3OvnXlrxdOctO+BbaMmT6lwbeNIsHOHE9nP1Lb3JiiJrougli/V2R
C3gH6f8D3PIAUa+L4eGPwDynAnNuAvq0TT0n2MSXYuXnVpBt40CcLr+/h73DYSxog2npMB+iM7Rb
ij2bgF1k7vSoaizaKSj7YanFH4a7r4tsMVXB4qWR4WigxCn/sxqDAEH96XZByJPxXGzeT0aK+IBF
WaZSOHFKVk8tkpaSjxlOeCwTmRrB7ohK2Div9QNKcJSEAgjylsPMwuo37BPigF7YGuvEf+otLR4Z
M/ismo9q8L8wLfaa3/rngDCfMtbQ4HjQ+jQXJLC5Vrnwex6g3PKag0EQRU1L5o+il+xi2U7JzIZK
BdslX4T3ja26g6PdPwFZBVjxRDW68/k1YRCH6cjFeV1iBCz5ZkR3JvdurPC22HmKMwlrRElxfAh9
tPpPiisisuDV2HjJcd0/a47oSyM0NXdwQoYRkZvPnDUqdct482WMdx7C8puc1EvmlBUqeTDugFr9
28A+j+XfqnITwMBIYrc0fObNJVCYjOUaDP4opInHNKSoH2a0+9bwHUqG48o5+E74Ni+xT8gmrhcu
joVv6fxDlBNQAhL1e28S5h0z0cOgFI4tdV15Mg/sU+CrEgwqspJoNQL1J8r80+6uGGyUe3V2YVm5
7knlf581wyOzk1EoTj+oT3VSoV3q9VORPzBR5YWEI5HaB9QmaPVsGN44Rv6exnzOmVqhr5Xdbynp
creUlXSvK4npTFwhhTl+RUehgnlDD2sRoKR9bI7JgH4dGXWP5FpD5knVyaXQIlon4GvIulOAanSy
JXyB6YSJ+tnGt0/4PXYalHrxob2NUEFFDxmiZMsE+ABaMZn+i+jqtA6NQ1k3ir9YmtgSuK+qD7xi
eSbJCNgKEcZI3YpiCrgsKjixmBCSoT4pM5O/8Jex7ToEiALa7kmsHW1U/V6VLaTv8ONY++To15IZ
FETEVFBTb+TeZ4bOgYaandGEm16pPhayQmnDvEp6W9URMqalTcQ4NMuj940N/CJBqpfIX8/xRdOh
aQLZL/EdEmrSlWz6n2O/TEK5YRSjDmNkKo8S0Fy6IZg5Skoecyg32A3gzwClAlzrG22BZk02Ygsn
zlaVE2SA2rmRQtlL9fkSUB63yVmZAYr7rNgdkqebzR1/Ex9SAhFOTcRYjPx7dkCVUyYNsLUwFdbT
P1cm6xrO1TdtUhUC7O1c565ScVLq40N2r685PQfAlSjLxCWqUXYzaEN0RLuSUJhDtW58JI58KiOg
Byt5cQUfKyCTvLTwp/0pPPVWyDIUBcPwybAvDN+KS5BvoVV0iIxNWh3s3pfe7i5xBfms/Z4BOFA0
MDFgjfLyRHhObUEw7w4NWa2TCi6VIEwLZQnYsWP7FIrKZ4JR7gP+d8icLCHe4GwQWppbfLsRJm6J
4CjSZVnJN5py559693b77ciyiJtjt8c9UsczC0MQ+qxVvKMzc0uCgeHbs+L8wyCdQL9Ro9ZzGFhL
4mAk2/RWCbL/Tbo4WaVIbhRMznFKNWOk/vuuWzgKIqPGJ0q64m1HVVTKWz6lBxl4gKTUes7dYFcn
L/81FLBuAOiAMuzWRrVKIKgQAwk/FtYkP2vI707pzCDV7IB8PNRmjUxFidRfFjgSHkD2A6BEIyVW
VJRi7+p87Crs2cCCaeIgXN3Pnf/VLVIFOqIGb/KXxndLLJyJ6BrhYemasxclb8sVDgUm61YmkSPt
62oThO1Ao0EolbOy+JmV2Vv5H3lqa2NJrFYKDHhhk+2ZUSXG6WLHjsdEdaWUDOn5ADlfgddz6nfl
qyLZOP3Vy77pnXhbByUSjfNnbiKUKBwcYdgIm1GcSXMhf2haV43cymekyqKdlCx4rlHDgnG6mMvS
4pAUqtsDlvHY89Nlqo7Cv+Bv8D+vCXwVADTbsGN/AlwrQjJ/iLFAgj8ymscMzsyxAEYlXJKeHfhZ
bJ2PhHNozJtV5e5xLgWoXYZW3KHTo3QoRZHMDokxv/tdrxp31dmqSgGc4auOydhE3Fs82AwRj+AT
G9Fjz5ypCU8bSRNvYmjt4GC8fMXhF6nDFoBfU1RaxobMAxBf3hZBxnvwxT0xJvtn2exNnJXx1u5y
eNWgYmbrUI/Owf1LBgXpaXuRGvo1w0oXpHQ3F1X3crElllWE5t0blPVanQW0pV1PGlEghQjbOmKW
y2tdCQgrdgORX5pELv6CiYb0R/f9xEDhkQe3aGa4q8mmQxMa8/oLzPMZJhPqf0cimpBuOy+pvXlp
/iOxI6QkLRc4t8c7nJgyMaQUKUhUX+6Rueee4ci8yjqbfLkgpj4oOxMjoYkDd1y1/1jgDubU758n
ktWFb2EEhPBJEgiZ9mgiGrnCbRavKd+Qn5EJIC7RapjDAOjbP1YqEu0dqkAgAxzE5oe+zc7Q453X
ks6OBf49aAOs8Em3vecb2tep1OXmRo5ijth57CS5J2S4X+OmwoGeDbz6VaxGIF5uw4azG8jVRfW6
yX2IQT55Z6a5dJVrth6hoSatbVnA2seSbqMW2C2cqkYCiU/Av8Xso5baFixJ4welCXG0l07eukga
wBar0f0rObJ6bStokJAioqIxHciy/DgEwVMHUO8o0JtNUAT11udRESZONFYftMWj9MUTNlD7vvtn
mTPLYGIgD0jwxQVhhgSuPT6RmUrShcLQxgy0EIjGYUyPaQwxvLb0GT2YSG+QNfyxdUOArxxpiuCt
nA954uJPAJVAchMqeK2jlfpV+dVIT7cHZiJfyrkpCZqJ43+mqK8k8UJ73wLazYTqTzf0O5ohfOmG
ezMhVtiMKwM3AOmlDyym8Bj3HUR9GP/VHAWCpAKUIZCBdz50cwx8DC0wDsFasur9RPlgV9TUoFxM
C6xhxoPPxiXri4+Al0T5i63SV2dsC09fjhRXmIi34UqDHAuN2jIfpmXjwlHgiEAAV4dOJxcO/ZGh
4SSHWD4I7QLHiMDzgWDapXiTs5139un2OT1V5xFIHQFGczFwwAPnHfP5osrQhkbCH+eVir75t91j
r/fJ3/aQOuR9QTtPYUU/rJ0ZyX1NmNqqAC1u4gJ4+Q9r/UdZ0EkuZ+g5sqx3lMxq/lK+Q0Wp4Cdx
mphHFy1b2MaLKW0RHhRXGLAQB5FUJOdCZR8FuPDAdqpRoQoz2MoXuPA5AKsYgoNur7hFxU0BJ1PF
jcUU/XxixjT/1guB9TuCavdi0GZAfmZEsH4Wcew8yKqiF9zSiB2V8f/iXomLDYyFbHWQuv6svl9a
2cyuHRZoBrnlYSElX/+GJXrvf/SFtVsxp+ubFyUj3KPGvRn+rL+6T0g/ce9LWl7J1uYm5W2ntoge
57sWpg5hBNYD/K64KJCrg91anxUWcYQ2Swn5rHGcQ5vOZhqbHj0upeNWKRx9/KiCqx5aQWiKsIDr
JaEcf8pMnMI1GUnQaF608GMLXtf0NXJOLync8uUYqxtKTIs0xMYxmlTVVE9eyBpKLogWqWSKVqsm
bO5/61TriyoAMMyVkatH6he7OXMNrAr4Fkq4hVmBE/P557stLWqlRPqigrqUdaECHbD4zK0hhtE4
oFFYdt3NVe0jtc2pYbNGzKIs0Jc6DnCiQjpkMTe0f0/zK59U94yH8FurzfrWSZ4b8X+jJ3OI1v41
oM5WOJSOLl/IAwWLpmHkVlcm2WIQ7ya8xRzPetssYX25qq3uA2jK0xaw+FHwocLyV7JnFbjpPxap
Fz9FmuB+Fcz8wwpwNTIAuVKLyQRbJiZm4TGNcl+SOujHlaTdfNYnRwUZ+JgZ0oLZ+69X0QsMMXhH
5vV+6kMiEh7uyuHwjpMW8QD+CYTcRcJ8smf5lsD+saSlUyueUwK9bNFNfT90Y32V9q5QK/BRRx0j
AwfccU/DDnNE7vk/+Kgc0znKneQnS3GfyjIvO/RzZfk2OeQ5f1cvlGOPxcPlT0Vwu9ucn8J+EVfY
ftmKWNdD0Q+KHejlCcMuEDh0s2DcQk2XPWqdM7EaVUdGSBTLO6qinOaXZlQmT66DebPa1XW18epb
pNXSsgQi0JKDgyLFei28RW5O5r3/H7MIUiCm/AOMO4GqZJoUMx9t/YkrMYsOsu95qIyyoUztNKW+
SlPtn/JSdsoI5SfjcvK9XLQgY/qc+VIS9ztosfHCqdZk9R+9oZs5bGduBwWhMVvqL2MoT7nnCkJx
uInYFAmd8qvw9hTjtbJt4OVlnWEizoEB4oAgdGCFeAGqCWLk8c46Mj0cP13Bkf3HJR7xGgKDFepK
8nbZhpIZ7ASx++qXIJVdW+u/Ol5RrnU1ldwYmz3ac9aGHxBpg/st3fTvsgYV42KEhKuyC4cueBOG
jToLQ9+/OLRv5Gengl+kxNbqjwBUb+jwwqAon9fNnaemTJRvwbDjZx5wLMJxCFtKuNiKT9Zc2Wk9
9Pxg1Y+nYeWc6FqyABBJpKfbBtpGrU33jh20VcQS44n1pYXSQswWk/mpma8eqq32O06CcYZdbvHm
qL+QLVehrUAk2RTx6OB6cGjlbTEYux6i0rPwD3VsSKh533S8IVZrOGNlSE0ehV7erWerTqitP2sh
VVYLYGn9dZX9vyTAHcVEoHME2OWbFcnJfw6fdEF5U+NVCYmvgEK/87C/unvQho3khbDGVmyfVyyx
amMKwRVj9LxNaG28uwjkboKt2RKQ78VRjtFGkvqhg4mDSHp/yVwL/GwDo1UGl5ZlnbZH8DlRCxxx
W/3/wckteYVLBiXkg/wsUWaCGTACc0GxJPBdqshvJV2S2TnE5I4V8333kCJg2qqjtrkgglswfnSG
sknfmyAi174BL8nEJtkXx+Xy2YaUn0DD77a0XSsdNHkEzYPmlZpyYy7+NYVIPrjya3CBFtWNHl1q
qGo7McKIGDUFMuaMk8lCCPxl02rBS/Jy1KTwwLRPzK34W7XGDzJtyZ8GE+XHD3cbXXKssaCTtiFd
7Z3/wE1/WCotG9OuTkhrJNgjpUmqrkE5BCrTivLj9TtOdnUA0TyELSD9mooMn2HwKktwlQo6Aqtz
RG858zQeadFHnmp9LhwUm22rHmqhofXK2vom7th54f0I2Ja9LmfS9l10mQgHapvkp8cmwPQgIB0u
HU5mCawBG2+psJxao65ebdHKvVE+68T0bSaWbeuokCVK16EUYfpCqONldfy63D5gJbQ9pmayP360
c1IXAZNM8E6xgdV11oGqyEhFx+FzfHuiD6Zs0rP/Mvvmd2NfxLl7SfcGZunvjIEkGlNI1Mnsutug
iYGSxgX3pfamlCLG8Gtbjn3Aq8GqC+pH1f/S+Lwqofzrbom4PQhPwTgGKeC30H21HjnPCcQHZY3s
BTOo4ffPDdLQXDbxVJLCxb4eYVs4px/bbGGJ/02jpEitMX6qLg2T/bJP0aGvd+jgnFqgs4fCFwnl
mF8JmqHFmoLtPLl504W/jiAunPckO3GPVsNQapWwGJjKHYNLe6U18eP+H2ZWjluW3j2msK2hGSYk
swIfzHNaQNQXhu5UdYYrdvQR7oaKk00aBkqIxzrxjKlQNh6qPToJLw4Mzc4S/yizskbB4nM1eTmK
hGVExOYcx+Zz66MegiTWEUC27Tw3T9uZC3sS8WaD2tEuT0OzcscFGwyHEl7kxLy0rV3gzjO/nP0c
9HBsR0NYnDShL+eTmbeIMgFA2cYuehBiFhMk3ZL+HTANY+rGDSNZ5+osc2RST+b3qD/byQ27JJ/M
KRNwid8UJfN4hu9WcAtIeYvQsXYjGqgoC9QfGYSAYFJC/TkrmTVk1VsvOuwps44meU4QK273/EAj
D8ffiNuNijEnKkGAuRjUJAfLjZfj0p5Y+W6rKsdMVxhcHFhH6PTj4q5KnffBVF0PRVpgLG7d+7Ka
lyKFxZqcD6JCoyJhLa0mJrZdgsEw8gZ+w/8zrBL9RiYG3Ju4fPzj4eO/26YfXF27Ukhgq8UNiNm6
+Hnyhk+QO1xl03o1tAT2QvVeCPDnYYFRrRFwAAn7ac0PmtGy+ckIvXjFaluf6Qjc2Cb10B5CbRXa
tHcThjc41QR7bwdZHwlIXyTSL+aM2ZFca9MulKBdUfP0eOsayxGZeKZsuESXy06qCUuJik8hifqX
1DlaNg/4vLrIy2jlsITvVsFj2sPSeT/aRNmZPjDK9UJLM2kCDKxA0gBU4qogyyQZFhIkBUJ97Bd1
YQxXfcAl4VuCRj7Y7hVZThZxUIRvS1K8ROj3mgroNbwGSRHqsTeDYUgQp0DWPx1jSK+rqE52Mc/z
Jyabsfk6C7rsIQaNIlStsvibxCzyqHnvVgG9dVpyTbVlOqeD+T/1iwsudNV1Fs3Nrfbl+as/6rZM
4a+nGN+Gh53iXjur5BCfgA30JVfR1HPMPLTUT7+MaXV2cf6DOyu/e3LI1NP6EJ6iecrLnuWE2ZaM
rBUvxM7S8xMioqQYdWHUsLHb79RnGUclDBm1Ft5RTICYAPz4Br31WbqXuuqLwr5klISoZR02bQ8p
mOueO9iJYj7N3z6YJtdZUQYmr2/daN7jx6ZX5DIG1nDdI668frNpE2D4uGzPvdLMDVYmmh0lDd/U
sDbqzU1Q09hqscbUMrwXOt1j5rao887IJ8yW1ncUliJk9F+YFQpAF4srPkw0V8NIBVk0cgK5z+xw
ki9Jykf4AR/BjJ8XgEfLK/diR0WDwPNWIFMDsjoHpa621+7QZenDQrO4BbOAooyFb4JXTuYl/7UK
FPLEtVSQnzKZxh4EThyqgWOAKXR4AZbENant8vJwz5/kTdTimcCz3fX+yzvNHobdHPVTf+Qg1gdx
DfX/5La7Poct0PzG6Hy0a3RScbfYANz/ykXVutIfvehs75yGKUBDG5HwI5nl+6uYTVqgpN0rNBAA
asczGWLOXbxvmV/JofrvUouvHqAJqLR4BGwlotRTiM3qGeBSvk6h4AJJwGiaCO/tU7jZ5U43ZoK8
RXfJ9nH7d69MjCEYRvSYAPuw0av6dd+YTO8Ac9P5QVg4jEiYnNle20Z1GuY/oULIGKEOVnnO1yyG
N15gb/BkxW54re4nENASgnLxDLhFRQVH1GlKP1P0ULboWFXl3VZpFNqMzNNT0r34b5PW4sIAeuCH
yaDQ26Tua2Xs92mkNGl4878aaRPb5GarrT1y9MPuysOc3AGoKjVfp+Vs/M+4W2Oz/rdmbrIXuc1a
1/qoQa2BhAIqdfXQPrdP2Pr+x+K1TyqPbvibCXDFfcEVWx3I9somIFMmBbHHi+UtYr44UXuRg/Ka
tPXJKDazd4VrJ7JUNfL00Po/tXk5UaQ8Y85YZS5hR/wHt+NcAVpQend6dnoNSM11fWDTM+VANQtX
a2mZuvqU8F0hBISqgB/R0X0ZKBOIeQ8co3adlPv22wKYEKnQwCa2E3Ms3gphiWqzzaRXyx9drufj
6cZeLDRHi3qXuoakS1uQ1QAMEU+Qu1dCvQhmN3jQFePF91oYLGdxzZRACf/netqd3oATq2qESNS1
k0Xed+EX54zOh4gLBU4GQKRNaRnssXgAaiGZjrmhy6ukF3GKEQv+t/g62vrHCwOCmzDGCbZY9+ZX
kili+D+J7lXbFDPkvW4sKWHvadKkpnJGRX6EhX0p+VbCTRvea113/yzYRxcQtBaiA6/ZXMcES6qn
J5iLrOs2vxh4pG2YJ/CtY1DzhviUmeP6Yt+sZRHMXW/bXr2GTa1xtGPwppq/TzhVMB94s5BTThRt
IW97m1HeD2Si06iPXg+pQS4mnBKihMGKNYlNZwujT3Wvi8rCvFkh2PbUUKtOBq+j67M4BN6RN5av
wrAzE4jsMhHUpXO8u/9D5D9ExOnnIziUoFsN1cdOl/rEMDx5+STbNWIR3j5fwTiktNFj73woZngk
aUANapgPAQ7OUvRIAmpuS8jbnIeh/JZASAWCJSPYEziDTDI+BFXkSMAsVuBNAgfYSoGYxeADNSUz
A8pYFbz0+CTtjW1HpayxBfYJWiN6NX+/XVuZnOfZkau1BquflO9S4wKOns3Fs2AFVl3S67CpfOXX
6rjVMn6Rq6kaYsDpb2hH1WPtdpvCMwel+6veUqCelaSXYSjQPifdn/KYAmbOaLzfjGJsKOmIa2nf
iFkXdVR5FfnHKheb0fWoLSWE4Q24siHImSVK93/NiIb9VkMPqBXDNdWxg0Uxc8QKdiH9N05m74+d
6BDbDy9H0ggW8HM0cqD4ImfhTeksMMAdIgcQzlMV2np4NX0kFGru1DGTA/wnqI4LEmG0AevU9csr
Y78CRt7B7tjki1YN+a26QubkUCyAKxjp1c8y1XsB5paJu+bYVnpQBXiXywuyX0FfVOIQ8FLtZxN9
T1Jz38ZM3oFnceeu7CinnXuwQ7NMXWV0391pRYj5l+pK23596RrqlVNxxMt3/6eqDiAPyL9zWVkw
EjY48hff8G5T6Qo091UsGhC4ICC4I6kaSERilJGNYdl0g92sVAALxj32oWQc8s0tEMCJKhPTYUJX
uCpnAumjzPPdEcIzDTFNZJs2m13AXYPpJTTTDoeheRy61oLh54neIJWLpKW9lLkyyibwGU2WP/yd
KpCb7oJ0j6+io0OVg1soSjHi6nbiV42OTqMOeoDls+3Xx0M5sIAlfB+OS6GQvP2KdXzzJy2qgG0b
p6+l79F+nXtTgiAMiTeyv1QUTipzxgmqDPa123meUZ3td/Eh8RA7aK6KrbHLfYSrsfL6mPTD5qSq
aOx/j6x2UgVxC9t9hTBiIq2wmQ9HAknITq8ihwh1U6dqa9htj7/QwOkU4QfC0bjOAeDj+c6BnhBC
ugq4tKSEvYi7naqoC+Or2xONYWTF8oa66ND2nj9HjN62dgJSUkKYjKTIyWF2gFphxBG9SdKPCqgR
a/A35rf8JBso8WNiLmrOMau+/8vrlTyDjmw0WVcDlErCGVN0MiRoi4vDaVC600fLBZqViG6WeePr
+WOqQoQGJAepzOqYlh1AHUO67sC/x6psekfKTrGjAM7yeSg2dFT8qJ33Su5gutfcA1JXJ4semaHE
0fw5iEpIWZWnNWMmbGVwdmP/YyzlkFYgU95CYE3gdREzEhIHO/jxfl2GBW5+GlHeoq/5IeQib31v
JmGeJtIBRcfQ3QQYHaKl+m85zUx2n8vzpz8fvnkNjeWxO4+SpnF/IMGbuyemNppBKitw9Kh3vjRa
pwuQBOZK/RQHbfl8zaRkELFPD2LGbKPCMRZ102C9M8Tzc0CDukEno9v3zKKmJcTq5K8MtZgVpzTq
DUUM5N5XxAQGHKGg+7xhZxYYlsTgi6JiSJe+1/gD+gH3//+JQxn3ISuLNgYA/9CM5THCshlasI14
xUAyiJYoN9gq4dALd+DTfmXIxLlYylSisfK7KQpg8CxBR3ZKSFAa/Hmk66tXSsj3uSJXngTV3m12
nXYC7zCSpDu1gJvGRiYldf5Ar2hO0FJWNR/VZ4AzfLzuIKFWLGWJnN4ZorIKVmck0xZi6SGnuzmq
sLMqyX0LhNG21WvC6jw+FvFFXIJ5BrLQUjYTq29iFubh/U7fciLA/TWS3M3UlNkGV6CvWtH6B1lm
Lpr0eFC+Ops6lhHFkAmY7fPXBEnRSbX0u7dgQjhShsUe1SnSFFqZEY0NGbi0CDGi8e/xzN9MumVu
nSQfgX7FfjnIpn/ZM18feMWRJNj2EPAclrlDlxhdHrXkn1lIdRAYCLiNeVq7PEmzUa/J/4G9V9SZ
kDLC6ozDxmiLbvIyMEcUk7iTVDs6gm79fwzT/MhxBT0lwt2UNNLSm7zzm7Fam5IWiw7QNxa05yeM
z9vnm/0H133AzSmxrBMESpeMOwb4vtEjhwdrlmdEqBI/3PCflSd6g02w9yX8MQr4/EPyzhUW63rd
CHU+ObW9or9EpKcptpR5Mc82gW4QtuPPHSc45hVBRq8sppnMdGhqHNr92b6woW81ckGC7PjzWxmB
c1pgpNprImq9ink7v8gRf+DcV56LiT+XGedghJpIQllMz6R+Buu2GfmWC3ScyCcDdyRGyYbqnJgp
LK3FtxXWwNb/3QX/ZjhYm/9014xUlsSFoZpWTwZREKUhivHqL4YbnNUrJGYNwTxlJvea85bCarLK
EBoMNRuocKySWRDirLsIl9W8HWRI08jFFC7Gzyv2uGzscRJioCgnIGIT0rLYc7ArAvDCwYfmQrtb
8zBsHITKeOe/bP6UxwvZQvEL+gpcSC1Q1xACSacPMhtyksEXbTVoBEu5ApUQphBquTPIbAmDhTSc
E+xbaIUnYdy9Cgu4e+iuIAOZjzKQJdj2o6/tzkK0JWQtoFir/KxaM7OJZLzH5C1lV/6S+zdfoDUS
cFlUrBqAh6MOa+ECE0AsiwC4nU6EY1dzuTjeBI3sxL3uXmvZvAssmzIRUNJaCyXo/7b10hV6DuIb
rOavvlhBzlMBSnqsZAn0/8m6IwdXCR+erAG4dbeeJqzB2yx/B38hAodgSbP/8cUSYnND69TeVALk
syfME054VK7iIaAwv7j1q5P4xwTGdkc93S55k0NXO2IHsRWn7ONGq4vCZXYMScIWXBOE5aScBHmF
y1YUd1g+pAP0aZ3wHu98Ug+pcBKvscubgAAOZvA/dFFYlHaMiouafYl5V4AtX/OaKBh14VLOPJoE
xOuqtB1CEYv4ONTbftpGKGq2MTz9V3IvruWzt9O0K470YyKddopPPFNJtrGnmmeuUA+rGYVzqSTZ
UilM64Y1bLTUR8/+ZsXSqRUlCRYp4e7SHTtEfxysDRJBmwdQX+9pRm6Xiu4pgfvN787eBypbCTUf
dtGpDWRYGCsdAjEoiZMmGTx5jcylOwFdZF5NHaPitqB84UzrccrNCHi9p0AzjzPJ2S2+YZCz6WTU
NJdE1PJWFoPHnlMSyKTc3gq3xGCtQPPp+yudMnuds4lD9G7JGEqY49d6/x0t8B4aacb3JVLVbfV5
jCVdZBB3JR93kzajdAg=
`protect end_protected
