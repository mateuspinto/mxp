`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
Wu2HJK7PxxLGtzwgnG0YRsfXFjC5fUGJcdgld0J8BKOUiRJLN/z41UrRQpprcWecWI70uLyaL4AX
doILZdkYl8IbVvO9p8Pse0s3WLsWBjPavR9QQ9JKUc1g1RpgqGIxDzQ9Env71kqnhPyCN8YIpuQP
cQJZcSehuBFo80n/YNU3MZmYAjoV6IiXct4NqHXW1lWPTbMDHxW1F5jtlcUnafDR9uqJmh4PKqUC
tqTv1hI4BPIvmw8wMoOfBRBkmCjkxqC5/KF+aHdmwZ79jFxzjRMPE0Y+HnwDi+VQ3Fxvc08LsgaP
T2vFe4HmDFwRWnWwmyxlI/BwRObDRPLJsacaIaKU4Wo/1ZJo5FMYIcKe3GVhc+cKOlt9S2BBCMoc
pYcax9ATBQPhuoEgeHLh2Zfv1l2gjtEEcvC9/tmMniEJjo4qR5F1aCCi+UElcl2uVnnQAdmWgNNV
DDEY7CFnNC4t8h1VT8f4ZCJpRnmG4z41D82YLqV80SNF+ZU64bhr4BsIJJ9Dk30ru7bwKIDXnbT0
1mO+IinPA3Me9pu+SMeODuLJJmlr/JHngHvE3Elv8GGqVvJUG7L5v4O3bY8tumvbi+O5Sk2QI+ZJ
UpXpbYHE11gzOmEL2+/vOpegm2SBysPhKN6VRMnDCfZytjj8faI9Ivl/zKZmoYrfi3lHfio4FVDd
c3zh3xYizOAhmyFVaRbVqy6OjUGZ8NPW6Y0BbkQvDX6M+x3QnBDzswAYW3Uf994+MoETcPlo/mgR
aUUs3ZC9hmGkgNDRbiPQkPcjZVNq6CTXspfgNcYu1mSCXDoiT0SUZ9PcrxQsDM/aPwZwcpm4S4Gx
oeazGimBnurDbz60qEGSGPFqauGbBnxGe+tRS8aZYcGd00maOFn3AYMVyKtnZC62Xlwy25Cno/LJ
Q7HYr0pr+sYtHbuFzPGNqRsXqrUPkMd9Hoer7L/kqdgQhMl8p9q+jEUJrs9bsv8q4s21e9yUqRTu
PyyiMqNMzV7qbUH9oUIQxTNzwoaYeZu6bJ5e2YkS8/w189i9hzO5DIJtNNRIt8+DrNVBdgjpm1WM
fThjr8y9/FsYLdSMOsYu7uBSAGSzen7JL/o8P6pG+/ZTzUvXSW/efCExSUV6gn0vzVrngW1Fgrrd
aHQ8VbfCd4oqgCnLJhTKJKEwP8YdIiI4ACBA7Iom1Z+xFaxP0cTjCjcIU5IGr4GUmGyjfHaxa0lI
uPh5GCT62PKuDMLnUKdA8Iad8DPxwzeMTYWuPC7iGF5c9i4L7+UgWuszjxsTDz+hOyxrXaabM/3M
fgbiIS9sy8skjjut+K7gWKj3dGv5QZ5UmBg5x4v6kDf6kLSfSQb9Fjm/To5zP18hnezXvjLeLGHg
kQ56pmTKBv+WN8M6jubaeQlSUYs/iQ5ZMBr1hOH5AVqDwsKfa9uKZPKcVtIV/EHX6j4fiMAMCGGZ
lq9UCLSjL1rvE+XNNYluBeaqxAfD2E+EcV6T5ijZuHHs8iczxqqFiQntjTGUS9eLoO7eWDScQQWz
mYCCDrIUwOmC8D5uU+ilUVBzcspgGQTxL83XhxpsgIIZ6BqV3qI4VvyoMhuAaAaKcVzRO0Tf2Mpr
HRuNFXgDQra1Teo0LOFEr3TkP6Cmwae1RoPOFyyt/4+xY/R1TsGY3RCMuc5K2J4yxid4bY4puSlR
dJFteE8XJvldVXJWIZmJ/YDW+YwEw3AJ5tcaK/xeH4sEekGF4h+Fg1//CpYUXGw827+Z0DthO7Iz
N0Fr0nsDie0aukdio5icnoNd+r+IwaJ35hMpFDIzfxaJgcXx10AUxTBTeD8ehXmD++c7aAYiHbU6
xfFn2r4dUvuziyXwIRkmBERFM+noRab6jrnyBt3wuZKs9hCDBcI4ElgGuUlX4y5/sMt70h4DRj0q
+O8GlDJ01o2JYWe7niri8FxmHMtKEFS5qCL2SBwqc4yBNAXWZKZqMM+IJWf+06OmlIrGn53P687D
DOWiX6IDyxZKB3rp2fBrKWFH5bpJAcuoT/On0Zzykd9nwwo3r8PcVV8kJ2adYT/j5whE8gl3aQXD
+8RVLxNWuCw+TxFDozT57Imm0+jHq1rHCfFu1olqfjXXs2HTIq7A6lfNY3myx8kzlF33WrpxY516
7GW2khwl65nCIhtLa4hv52/fWBEkCN4xWZ/tF95jLfLELtTFqM3JFuYUQNhVilcfRCl6cYa+/uD4
S7r9TmG2weJM1ME2qvfvpvLcvjDEmp66ub1R9yBgc7CdbAhlDzULjD9TwuvDxiwumCt0A9y/iBUO
H28R8L0vZZ5patOg/3y84Yq71LpvCm7Y6tNrT+/t5igwfmPztJO9M588xJ/NqiWDXDmgjzRZAV1u
gusNk8VMN9aMH8pS/bYzpsUeZWV6o08VhTHKISRSC+aAQD0m6D8UF9JItSunXwEJwVTVxuX+1hF9
Wna3DBKmRgv1RwQ6zL3Hkq0gXTbLJzo9Ur7C9Y6l7DjldR32RDmoPrrIHlqzwabUfwou2RXHw+s1
N8fTbd370VPWWJ9g8Mh6wLQdnq3D16pEUxpoDW0qZCK0MfIc61Cb44HtmLR3agyVyLajHQo17YSA
sAQvL9NhB9eGS7OPtAXUvN/9x56gB9m8SPYZuUgYB97BY4ETeWSwh2eInG2OvFJI+1k9vqCh3fa1
pwixHRFOMX7Fz9LZcAkhoPyeVhwQw/J59Knopp/Cp4MN8+63Ige6Ykz4tXb+IuGPs1pXM/he09FH
b9rDcn7yURgxhCfo7h2RV2lb+mg24xgux2xAJn4dhF8IECYXEgS0V+IWUG/Km1s9yY+bR4bfMrPb
G131gfBcSILRPjqIHqOxjjJhkexaoey3yNkgiIexzO8pbZjBiigMebebtu3g34YVdLopKYSS17fT
lg213oRNtY65wIYyjsHIWTzOF5goI304xcW9dAsX+g6ycJD1DHDoSfchdo9R6Un4rYy7OzYFN/rV
kroT+SifG0qLAiIG2139jpS5UwqwUz808Awjye/LKfZN9CmnWepxINDIEcQBqj2L5tm/GpAaUYiH
JGroNj26G948e3q0gcv+fuSPXO5hRkNUxBJxSHhpVoblyqmPzYOjTA4oWbETqEOWHQSgGlYZ8NVU
YFaZ4buqEhOY0q/0tW3LI7XkKhLcb5PMOFZ7xJPcqKUHbEoWbmHnJQkMY0oaihbWZ8qAz68NI3hu
OUcixw7e5QpvZuopcJgrAWDCdLUJd/SA172fHInkJ/0xxT1Xj/iJhMESREmXZEEw3ZDa5QMJzprx
6UNTHNGUoAcQM7YEHwK9Cy2bghxialyKMrGsKliq+0fDJNV9/dNGrd9AFAcvJdyGK2WTjKI987/E
snIudaJBsrGQQ5tGIomEKTU0heybKnUmbC9ho2myZrSLDDlC2sLvCn9LGh7uicILhN5wYVvRBJab
uRrA7LtpIwJjhOHwrqi6ZOcKLOfOh9wro1YYGGPradIBuQcE3iDKjv8VagCRgASGpIFB5z9xErHv
VvHXFEdesECp4xDLmy2YDKJEhz2rVP5UHJwr6AZiAcnuIpq3tnkYBub6fTK3s0fwefBDl+Aq/8z6
5QGdlnTKxGeqve4cgI20IReyiA5g5NBrqaIoCDeNahE/JFtfKtkQouQxxhUB5kUgh1Fwcq9MTJug
EKHiOARAt33SaSuBe/6LBv+OSrdlX4jG419y9PRT6Td77Vt0WSOqguZHFaXnulP7RyFVBGxEpt4T
lEegZHD1LeIRQ+thS3hxX+OTkJU7JOPPHOqv7rLqEdc9enkq0f7vAsmbVgqlK3ocUXRHaukTo+vb
pey7a85PuXf772YNOa1i5/zS08oy59WY0v89buBvWObOFx00V/6mqVtk/01GF18OoP2xEGsyDkO6
2WBOynLN3zEzw7fcu08mWjBd6DygQmgq298y6MGOySyScFpLhKJuyF9ffkjVKVYAmaA0ncX1WMea
9otorFqR/txAKjzPGQ1jkN21U1jbmhks0gyHyZox1Ttblf5UhjB6Uvi7l8Yvh1PSWuLF9Hl+a60n
lnnaVtS2Aqco7K08nDS2cOLPNBX7OZ1vxDjYjhezB2BOIfsZzfrdut24Euux2YocgN8SVKO/PtnK
nID7C6RSEneD7kr3YT+Onj0Ilr5C8Dnd9co+wWHLnaCBI/ZAxtkTvPDuqW2nkFVom+ZRfthG9DZQ
ZYxauHBJCS4kJVmnrUJGC7HuvQSRnThb2gR4gZpp456Pe59vA8gY6Api9ND1ShCEGbAQH30jqHHb
gC+8/rdcWqQjeAkMEZLG4VMHCPEPQgtwCtd1ASVHyeCY7gMHvvMeQDa1fwIrOo0X84P2AACsqkl5
6BkRPly8m9IWv1FexwT30aFNxIFkAGWyAOIAVybtLK/76rh9XkA5h42nShqH8nv46+iSAv7JSo8s
2mbCxVPjgEP4ZFp2y4lMAhLtabWOCWLDbNIrorGKB3ThXQpMGSpi3l0uzwFudbZftyViSvuE3SVT
23zGKVXPwPdmqwxZlZZq9cvjspUfnFnXDGoldV1xa02/fLpXykSwT+/91/p6R9MOt2LEf+Or8xAv
6Q9mjnrRPEXpSWzkAynX9Z40Trz1PUNkNJBycd5wzY5gW5e364g3S9Nu4mHhQ0xOxnXgKVI3k2pz
S2evXnqlp3vNDa8G+Xd16YkMhtXEiLfveZHiHUzny6n/+DcAmsMAV5tstSjgo+Wlmx9r0loDxv82
zlXfBMyoeLJXcQxDo1bm1zgGI0Z9XJ6Q4LJtWCsh5PzWC1WrWEsMxR/yHODZe2OdGcAQcGXNT5zF
5pCryO6rjjhsCn8uIaPNPB1LajbNof5x3MS7jYWIcbhoysMe0omEKrf5nMb+30RipFL+pjCtQFRx
IYi8uzsS2w1ZVly24wkgMQ1uk6Nn6MENvALxhZBRmG05z5nBimgzhYBlnudBUiUrkMbC2M3NpkP+
muTfY34BHnvhBHW+3dRy183iX1HZL2ajIUoUnO9eAaMYxFtTWkquSsfUxtulxM6eO594SIZLUH22
gTVScuKanKMaw9iWMdYqeYi9xT1ODYPy+e+TtOYWTRuRr5P/legQdSRM/csDPvLK0zErp810nzEh
fkFg2mQMAn9J8P00aTmKiuX52+p+taabpXsNIvSdpuLuPh4FTnVu+r9f4akp12Y7VrQsJwjU5t3k
b1Y2EDpDG8O9KGZ8OXzyOnZJ2OQBRt28oIJPfLj1ZEz2XAyuhkkABBmAvwYjHE51DSiNss6yH1MF
HVPAimae971zn8tBSJr0Q9x5Vnq3em84TvMxcBQrkmoWhXMdUEKU2H78XZn9ykTNqYmQS3BSwEw+
245Hv6pVVxkhEQuLFD+rcQYk2dbnGo22G3ZHf7aE7zbvZZRIfAEZDnl9BRcJpzEU1yVlxz30kEix
2aXg6iSK1AkvB/LJQlf/olYl2ScFbEpusc+sC07VtoUfkUftwkonPK4waOgYIaETFhu24c0iCkWS
sgfc7OMNplAFJlG1Bo+COk0p3Wk52ll9IN/lPvB/G6q27VMly5jkVejaIj+EYb0LaTxV5l8fcBTJ
NT8i4GvEXEBzyM1qqGYz7rJgTYn8gZESf7ssTqWXYHy5XuW8bO3EL3ClKEH6SWuIITME9POh5xX6
BFLsxU9Djd0fWtnOpC+4Rg5uYRbEHccm3YGEZaN5Prci8JXPmnsXCxdo51huu8O/TD+49PYaCynb
qhbJSlmLzLWjTC70mpB1Cn2+ja928F20daGLvPKUQUpP7oFPr5bfsh8GkHGODAJT1f332nNKzq1t
sjdta18sg5ihb5xpf3mPYMZTLOhdRqXlVokUW2Xzmh5q42aTOty1nF7sH2U5ZNRzvwje4pPbwe+l
+U7NdXpK5UYueNotXn0YdKrJP+LWd7UBPz+nrgzJBMptNKwYIh92BwHdmTBd72LZyRp68eJusGBz
LWNNaVH0Qih9aCn+I3AoCa+QHGDxz9XAvdnEdRN8KTo9OvDZFswDRqWu+X889/qLCqgcNlpe4L7Z
s6lt5n9atpXaJtk1ZDZ6n4xruJQ3Y0DWY3vDgpzTRzvq04a6hA6o8aPYqw47X1DmgqkyA7A9cHHM
fBvdQdTVDLUcLIX+tqI1j2IXRh2xXxzVzgTm7Wp3FJdHJSHJDk6SCue3vw4cT45TZUpL1+ixiI5n
xSwqxNO63WlnkHIq5Mi4SH8GJ9PqvhbgnuG+IYDYqqduXPWdAn3ZR6qxENOsAuuR7GPnbHuT/C52
g37PfHpOwiVGVB5opbCrFuHdNtix9Kxt+J3B9TIF6QJhvU+LsoMTshHCovaoXc65VQ57b47jlhTg
M8uDgdg2Svr8jFnEoj82f6xD66GL+92SejjAnZ2+MK2mu5pGxbdYpdj3Ebn7J9fMqK9C+VrFgfGP
LUtIdezN0OtxzNs4JjvTSZfQ5KwDDNqlAZ+K7DcgtI5bJcSVECC2e6TLYUBp/pOYpUOj0uq51RED
ZQAE6N+Vm437jYaCXPoWrZcRQw26cX9FuRwfYt90QSXYzZWPn5vDWfg+KeJXl6yJTX+pafcnViuW
Y6hNQQofQ7zq+VAmijjKnYUlIlVTsK9BSgiu1trF1ljnR/tB49lA5ojSj477nSPBQvnnYy7y/aN/
IYjH/k4TQdjkndbTaUxRBlP0yfJB1VsQPG0imhhUkbn11LPiClf8AcCp/xKxO9DE5SNlVg33ItTZ
WKBcvzCvi/14DgSi8n6B71XTnnNZvW8slm+zacBwUrYq1WF8DHzX+FnbaM364R05pEZ6y7UStj9A
7/17uy1/SceUHdF/oeqUSm8LuOo2OaCrAt+mh4Yw7cDb0aeI28e5mKsEuWwEsBZO5iNK7nSnN+wD
bwASUbeuTRy1idFCyqZOdR5bmI8tNhplkNud8TDu4qj+vJIL7G4FQwnYRH62xUSQvWjm5PdnWrL+
UR1c21nfATHCsHG5iTfGvuqp9V7c0U4wsCkqdAlMCB9OqMyv+2biBe67aFYlWiaRF+N1UjT073Cc
OFVR8aqKH7ymyPeS/M1e3BE43ZjH7ylYbsfDe4BoOfU+V2Y60g+oYY5urT+f6b17OVrkpvKdmYWJ
/tLEmBM6QDoZK3Bg7N+CLlKebsQh06Sn4OIUmJRWP1HHUNhD1rN++KcXeOW4cOxnKIvHV3LRQ50l
xkPGKzu4dE3zD+3kRwC/QAxstxDNd7O57GNdXA6qlViY4+aXlN9EkfLgRW7828XcHHPYqLMwkvdX
h1S6b9BC3H89UXyuuGewSlk0gXGRNXjlnBjFSsRwJGi1x/yTVW42ULa1wp7Bb1g6Nnv2Yk9y4jJn
cAjAqtZSadLp2JtUsx6V/XISgE72nP4lIlO6/wooKGSyVnUb6eoGz8x3comz7XfSjL/LtpARDEHY
lN1W388g/dl4VslEYdaR1y7IKoxWlw3EmkH+eAtTbfdiLpaIS5/rQa1/CJdOgSG4NPSqFAVoh3HQ
1w3vP9nu0MgWq2o76lyN4qKSVeXC8RfYypBljwH4UYznI5QM+3UG9InIUbbAjL/hcVXwQ6V1J2nD
zSyy3OZNdB+aUvGS27+6Y9IXIy8rD5JDKOevJi5yuGiO2IUbLfpmOtvW0IZYPA+nAWtbCvGgmRRv
4mfD94WEVQOQbbakKKOsd7dYYZdQImQlPAZuVYjxEV1Zb6q+X8pefi+5ds5/JI66SMybz9SJCfk0
EjeC5gm++1PoYQwcn95/FEGS3I9KFYRQGE43wO8iBSupEDefZeHhYGvwXayYtc4yRHknZ7ticwPQ
0a4RdnP7YtjDHYN8EyQSuVmvDJaiGpRGIsefHtvYMATiOwvVncBFHzlj/pOIlS/0lA81U5Bhkr46
A957hwsxv4vKjiuajIo/8hXAjTlt1OC5RTEa64vJ01RxToQabLTIIlaN4sLwLgwfhwen9K2QLLGh
BYR5cYhikagxPlqn/IwtEEGIsrM/rjxiY1Gf7iAKPTK7hLTEYIVVGwKbM9P3UcuquObYSwmPjUsX
crfRXY1bWBHmXch92CC7nvQDWbgi5k/UzgNfawEV9rrf3ol1gHdl5T0mhl54s6CRhnXIun4GrV/K
01duWy+m4rWAKyJjfvz5IRXRVYU+aD8rM9bnTlBIVt3WFJKKQ83ibM16ueqbzm0Eo7J0IC6sH4Dn
1fDuyScIEZC4poBKef4iX3DpavOWxdjgY1YDl4HsqvKvYKbmEkb6W6eNY+VrHPHIaWOmmQ9L2M82
1v4X1eWzX+fqSQu4MSfAm3Ea97YHrBXJR8SokjRLokP9EgFRkncpSFlaTt3u998HmSeqD8Za6kBO
XSTe6I1ky4sLiYFOJXIw7D2HfotXRUiSpzzRJkKG30NfW1FnzkEnWVFNQOEvAXAr4UbcwQ7lpl6t
N1XyfrTpEcsYElvbBLvjCivTiP9KuovD3grRnH+3ZBeg1czjtV/6FjagoucYhDiKba+Qe8GiJPgm
OxIcOcxbexeQ0i08aXCqM9We3K52f13Ld/qiorQDvk5KhbQeCDIEIkeff9mTo6d5TUeBiIE1KC9I
F3bREeV883CdKHacKjD9Jm0VwWO/D13ppleiuw2WW0JzUCe3p3Pqb9yISr4+i37amiz8vR8+Mdyj
Zu0XGjOuc8idNtNNsZSpvcdkzXSgo/8shvTd2u4EwiFv9Sy/w/jjwUL/t5nedpfkJLR4m/fsH04b
6p0a3+8G1ad+YfZ/nygmKU66j0zRMMpyhqoJ1in72xYePLDj2JhgqTYsJx5dyheNExD9zzJ+ZZPg
RDCLB8gfw1Moia4IxHbrdgy/y2y5tVCEs35UwiL8z9Ox614kAe4pzYB1CsyDOOtpim/cb0mSEAXE
7N8SNtMHf+0nrHEZSU3NUXi/KgzbrWIXy1+9nEEfz5WxZCugVa8bbVLknA2zBX8JMYhivFa2osRg
GO0WILvyEKNzibrMvLRV9rsCaQrnlnztIYQm4Onzpjdgu5oDYi0i/SmF1HM1fLc4798Aroo/ZQB2
pyxPlYarERaqai50gzlN5Ml6yVFmZJCmETlpL4DTue2zzNpRt9qZm52/60smPqyUV01U2ioXkAlM
faL5Qy5V46Nez7wzOSrCbQLtH/9NYBXeefAo23XGodneyGAoQdtt8FoU6j8Yjknwux5pBptn9oWC
o2y6UlW6InIORbVyFRf2VJmmDtHRD0jXoWMd+N4ehHBKD4s8APThfOgju5Ih0/GBNgdy7fvw+I9w
pa68fnJ0s6TCRBL6m6ygMeW1hhYxoZU0hWz7rkT1LUC1zkuMUf9NQlBKfWY3H/7SvkT+B+Yu053b
ofTwMVEcZJxqFAEt3vT96HhW/i9qDE5N6TxsmgoG6GwN7EJlXAmB8R8Tqlikb7Dts0mmUEbmCKek
HEwelFAd8FXyxBl6YMQfio04d8qzT13soJUWChLND45e92XoBaUDZkLjn4HWpfcia0CDVNx7VDry
Ae+0MA1iK/lnI7w+KxH3AIVSVl5O/z4wQuvaKU09rZ0B4X/tug6nye6MfVXDI8u4+SOM/I190uuE
0oQbYnwCVIaNEqC0s/xpKffTKb8Qcxz5LzDTC2yUyga6xXpHxKOUCNpk5+xDPA0oiEgLjYuDKUbi
Pk4ap9SqKM7bhM9LPHjZbschH7krVHQWGNdpmXCYa7lMEt9Wc8BXpSaNG+kN1G0FrvApv3vSSBj6
MlwgRFCEMAjQOV0zy57kZIN8uDtw5J+AAErBRcEb5dChzrqYhsZy8v2JweGzQDkNe2fjCR9FS0hb
rMfhzyfJz+Nicy4UKjBZQu/DzMAN6Aypigf7llYo7TzjW3ioiHBnCIE9E0LReEQX7KhNVujLp+FC
FOdmpysBH+TcSn8Ynzfn1CKB6OfVOKRhp9eUyl7ThHN+YUT51hfhyrd1+zPMSrr5TenZISVlLubd
Y0WagsYCd3mN7OKBmXVro/61SQ1iBl/NsCw4jyVXq7JQ6zBcBbnyFO6XVg4e0freYQi+DjtSM9m1
CA3oMkEKwNXIWzWvLj6Vyf1xqpy92rFHFtSZQFHkAnPcBGf6oX/Xa05Hv2HekAlJsWmgq5iThOHY
xu+TRmYcOIRwEqYbV4UG20t1wzO9fLKcsYOEgaxecpA4nJSR5XUIk7W0u9nKyuvbgEY2AJZZyeeQ
YKYosh5ocuMchmMR/MBLHrK7s0sfJtxbjmDKCibFg1a61FbyAUUcuO2qxAKQoUez4TTR7nncbfuD
+Unp0emVCGOG3t1+Y0UYai7CfjzKv1nJr0z7vk/B1dYcXmcUtnnLpaWUn855zck8u5a/GGBeF6Op
974TFS7b1UcBHn6V77opPYATQjRs8tRkK24FPwPJb8KhsDa0Ia2tO9B6XzTu6RcQ5PQWLtQGZFPf
ExtajOKm2ym1MdQMXfAo5qUzZdckcsK54JXg9IylLF/Cvojz1WMouv2D6MTaANulkY9AfyRi3c93
RZ1aOVsiIUEyUc5XjcczJF2mxyCJYQpMdUo+zuOzFbWN17v22xMcEwV/Tx3xEYI5jut/uvfVDkZQ
iWWodETT96KflfH5VjAMPpOfUmgka/5L2FY4LuwRuiEXuO+b+cWDR+lRUMQiNfNvAkA/fZ1EJFNW
G4/GvTWfg+PnPrwGePk+SbMc9N1AxhLTfJN2RnWe8eS5G7oWzSNI+dP0L2ZwYjnW9IR3rB7INUGK
HcJ887TuiAgJ3M+jM4Vfn8P7ddAw2vhpf0i2UZdffpQQ+kTTEHeJ47FZ4O89SngIJP1go3+u5s6C
CpOY58dEhc0PBLBKx9w3E8eJSmC5d2lRFqQK7/ZkxB+WaAPF/j4Mk0EAtyr6soW11BJNiNEzoks/
4Xdp1wWZDFIZOwMSyw/egONBPABwIS4k3zKGJSOd/qCRcuw6L5Hhm3YWdJIx4VooVfuHRqLB9CHS
R1uxRPXwWewzbfOXJ7cxYuArs7e+bbiX+4CrsnMmhPgG3gM06EtBx3UffIJDfT5o+kGaA91MiDER
aQpKZFpK/c+zKhDnDfSRA4/oFmLPMEa4hiCjUDMb4e0gTThIvPFkl33QB3IGrO8EfJO3ykoI6e0q
RECHHMFBoDz5dtgVt4lpGkVb9XIFL4Ea6yjmeqmuyfKDADYBt/CD8nLWwaBYtr25Crrzmi54F8BJ
r5y4hxRW+gwk84NmM6LSdlQKhMvg6pqfPhxkEhvZHHxvJOl910lFoNZ4YXG/9+lBz4v/rUufKesM
h45nBqtVw8yQCL1bJ6FZNztjuzXu+LQ+HXlPDalyEl9GtaNVfmHLcIhk2Y0zkr4JhnHGJl7aKufJ
zUG65Nv+Y9Ta9vesQDPqEEZIXgOG3nqgQzbWHF+os8f5xVDbVjF5szsp1FqabDC0ctwwSKY9eWJn
zqhGX2PHXf1dmP3ct+ujEDrPRuT9j4SlY4KJnYdbwh7Ub6n4DYqtr2KlAYKnfb8fS33kyE1kcTw8
736BoJ1rosviCmT50EWUhKMAQD97elcJdF5XjqtPbm7JWABddYpUIbNhPTDtmmbFBUOE+Hg1Jfg/
4GqO2eTKgQ36IK7rD8a9b1bOWwvlUAegk0jPC9NBweKH/CS1JwzaOmXLKiIhHaHynnO5KkHEB/Gq
LrIbnsrIHPwDjD5lxgCUeH8H4C08Cx0hzVDR0BEsgbK8ttLP1Bo2eS8vI7po88kwoYxSO0FR7fai
HXyKBSgK7Oj/ZCFaHNYRYbevLLL2VFalfQK6brQnaKZzmRpOMbRm6RiqPGfYKlNNSbDbsCMUP/T5
Q81asORN0Mi/INRgHgNjqM7n9ig76UzX2c0RR2b+JAFb8fLumUtCPGacrpijcuNOU4mZxJyBQ/W/
rrKN2Mus7Y653HUGLLbO7iAT/GgPDIGSd8zZYulU+wre+MOVM8QiK73CCFArrwYmx6ewSAQnUCfM
uopEzAYG5FO2VZ3w3FyUb1yPEU5aYAwFrn99XmG+r/u7253IHpoA8HXHzYUfKfFYTyaZbT1PPSko
vglVpp2DLD41GpChfoPOmFdrqdt+cSGHD3YFvnDNO12k657gDkHAxiaIGn8sSusUNuHEvbe+30XL
/kANwL+ilb67mrn0eJJEpS/tDPmHxya9uAHpJuHPfb2DAOS65cq3nC5QoUfcjFvP7QsCB3YjYokX
HK8phIjTiWHOWD5TOgHq6F7k67AxYH27gmXUtNtJrFDYsOsx/VYYer5ZC8nwmJCprtYqjiA8jd83
OMM6NmJaZjr7uD/mbesh+mkxoZwImLFUjb0s+9ehwVUUVtT/Z7R16rV1LkwN2gv0dN3vCsVXDxgh
m/egeInhtXClHMw0D+EDvp4n0wHORwXrxUHhry6vkx0PbQDMkaxCrLtmYVLdLZA83A5/YKoZgYvF
+4fBZ/OYSaE3KywHKYMVgX7YPT0aULIAG2/eSSjoBGcl2w9lw7fdCSUFD2PABDuhAeNFXPQkw28d
Uq9OARPaoqxX2GocYxcWRUuvVFe6oWCzOP5z836B+vJgfrgIQCzNP+TvQ5zmf/+pkC5uvzqSRiUC
gycx4dOhjMPO4cTk0K/Z71uX4JD63A1T2e0IgMMDpXliMgdEMGOtGpMTVBX75EPv6+NkeV4kDwBl
Z4gp1N0o9Z05/+zem0aOG3i5pAlHMWR4MXuVptQe055cOGZNV8SGJOL07jeVPw1SNnzMS08YwJpn
QEKvGklZPHR7t6yYS55xwvSX7D1NWMH86IYT3ArsnnNpn/sMLmtpr4Mh2zTEWvqZZJsrqhWImsTW
bSMkc1LmNz/Ap1rPWeCwCgerRLLdvF6uIZ/LPFCgJcQL7hKOwzRdplt8X0vWrFwPmt9XU1ZVp6ZE
gco6eDcc0sa2sep87pUW2f1Namfat6i3m9B7+JD81R9ks+B4C9kEhWZbBi9OEyw6olE0Iil9bDvD
Ni+PfzzOSe35X0Ejg7to02s3qz8BcbVMzOd/P9vj2juDp1yxatpgm3Qi9a571otBh6l/x9QBYZaJ
c/du/AD/G8j5NNaDm5fQNrl+Ypt+umua7oWLvo20qcjKzxCVKXz9gyjvcvaAvEkeYwcquzWZzaxR
NJJPBIEzAiiN9Y+9rNnTqsaMVC+uknJUcWo58U+I5i+0SY0bl2tFHcx7CyaLGcUFj4qxjOM/ZbbN
dFHzlfyaiS+mFNxDP7vWUdEhkj4j+Zhe8Pj6Y6B+eEtB+k2Dlxn46BcCG+hX+JPwZYLiud1IL/Sl
PX1hBz5pQgOhTimibiitb7sayA/tnp9fkuDVyfQtw9nuWOAhdU2i91LJN5QTaz1mtJ53j866o6Jq
3OTpJS0dY6bvUUwrA25dUCdJJ0wrCBoEkbIDYi92PtwiiBUGAhlzY2cnbVEUeOMtqECRsGEfZ/ec
DSh+MItl9W66XDzjkjwauLCRGXulGvSj2wFiXxUGcvi58NqKC02s4lmSI6fVTDzUBdutZvwwgzDO
2QOqo/n8ntTB9ye89dE02L6QoR1//5n6MeCrfY/2igWKAL1q+ZOvaXilt3EI8PDLXnZyzgx4cKp2
pJaY0kzBzcYZuqtAjey8BXYs0UxWX7jVPHHpDchcM7ECpydmg2hNczwIvJGQp0MG4R7pZUUz9Yxn
kurcaBXYjlvw+1o4HFPCca+WCcP4vtmoNtsg2mMkAP5nb+9E3OpezgfxjEUou6LO5itqMxyEuaZS
EK0LLHPML1PInJlMhfpyaoW5O0JYz29SoOJkerw02uNHS8fLAlvdG4+h1Dtd3XDzCqvdkM/4UTLV
n0vd7YomJekrcC8gjWrG0pI+Vd5f7RLVkJHvIjK35eBKE2XJ2uruXbsWdZ0yKKwz2A/lqXeTgdYB
2bCuMBzdPU3vsCyB4ZJ/r9Z66Pj7KzH4sL9tZapDyqVcxB3hfE1C28JyDCTHNWFf+5I/uluqFZRO
PpUVp8rfreem/F9cPtpvP+gglatCu16YEiSfOuN8BviT+cAcP+giYI1zOD9LyQgP4SF79vEHAQCG
JbWk79MFKXDT2cMaRCbREE4jXuAOsNOLiV/6iIrEiUBVpMiuE4tEcayCvnciE1LLk1u75s8sJ1qz
civEN5iKpuIIVU4kud0D4JuEc/pTv+QRgXMY2wSAE1sOMaUE04EBknKMW3zrgrS9Su4+uMwHICA4
E/WX1D7eNMEvigUzkAvqDr5cYBq/BzaYI9/Gxvb7Bn9bNFVCn+9k/iN83KSizMdqzmQP+GlkX5g6
SvmxVQtskNJek0wVW1rfiLdRn/ifA60e7PG3QWSxhLrs9WdY3mwjWKPErQYV+tRPMizqN45QAXd8
QJQHKXMwIBzMOk1FounoCQo2ClxNY4CFbfREuodlaklvfI/Gvjj/RDk6hynjBeJxE3MhrAk/ktMW
Wn+vTEEQl1KN/izRiQWBMSKTXkoEH+ic7BWJruwoeGNZ1BFs8DHqU6nCtmMh45jHhNeRF/O9wArH
jIQZo4cLbOHp1sXBEW55ZCxV3XrcAsoz9ksosI6hmhviGT2jUQtyOWJWtf3a5dFr8WFaByuCAxpR
f0G5cX1Y8OozxKSAe+hjJXMVG7J0yAALja7kFeeUXB7KTeSYLLkbBljUQyIchAEHtgdUEGr94jyI
8A97h68tPky7cAyYWbbjDPyRHRjYPigGtu6WIXgfZ3jdZGYUGhLI3TDxiM+vS+hJ2YVwYQYj0UlE
vWLPbNkfWf11FPBd5pYwIAZQbrUBtt7YQquvj47TCOCRRRxPviYeVQ/8V+NDEGN++7MhZoVxmOCz
Wucypv2cDGMCH4o2UqXeN9Lxi9UMc7Thgv5e2tRTYmLM4owzmLceEm9Yn2leW2g5n9UdJFo/jnUN
vwiQ+b4EHwkcytmyScFPZHivfZkxDslA7p0Gr8u2sRzMXtZgPHmLALBjnp269AcZ9b/Gce3Q0zvu
PKfFxlbMF/TqTlyYtHPbgaO6X0B/tr++O2olgd0UALQd0LwWRq1b6Cue/9Mji7CaD5YGzjlLVZLO
iy9rmYpt8y0CZrYxX3VQhTjie6Ca1+Tm/vRLCzy4Cd7wi6NAVkBezxaPu8vhssL5Y8831TWDC2fb
o4Ma23xU5VJDIhte9Kn9tr8nngZeBzt4Ue0aJOcJjKkam9s4rOQGD1OpTyfxjro723fyusL1DDRk
gHaxb/9GTaGmaMh+k2/hR5iAZR5kc1I+lDBGHi7RfQorQZ1QeYU/F4y/I4Q9D8LmKgPotDPo1ydP
sk96Gidg9Gjxxw9Tmx6AG5AF4uQ/w3BZ5bYyOs8mZHVx0OmdL8VSBbXno+uiZuzCZmbFwzehBv4H
yc2NoUiJbTC7zLEl6M/Yw/1Hv/Z1cwCeGGcD2fE2VC/1OEWySc0WxmsZxHjFbN2FRJYp3CMSqGrN
VHnlyEwxCr3ZWIUj+SDmUXZctOoDgTqMZQufKLtDP2SG8pMKc+uhbeurdf29Tj+6mGWM8S/6XgYF
/EXm0pCqdoBjNi0F8IkSneBBdSot0IogpOvS3iy+Gf0wkZ3JCO//gEUAgeFqJG+I+yxUn162npNp
XLfPfx5ONQPJkzN8pm0L6luBljUrGCu5Jt59x54I+gvtmIHDES8lL4/WwESQldf7IG8y0meJTrIs
mQke7J3d2z1C686dROXK/Om0SyNg4bKkBVgXd2qB1OLBuCMrA1WFjvfkwQXhitCmmiIphYL5JZjV
D66/IqB3/Duno9ZgzwSjJWVRUQviy4hZ7EYNIdj5hjK70wRCg5e6kwzluGHtFiQVs2jko+IEkOET
o+jKRCO/gzWBCkZwxqKoRqK+MG2HvPRMsXDde5r5vA4FRkJeQ+nI+CCTxtw2epwQB98TbaCcEIIG
eHwGp6kTQqFZTzaCnd926Vil71N0QI6P/5pXwpZwBY0PpN3mPKtMH/bzYXnPTkwRkijDAZq47uSK
UnK5UEIoWJgxGXKUJfWR6L5vqDorv0F5W/orEun63BkLhS+RgvdiosQo1Cues7uBwl74gilpJLM8
JhN3DzDNiJZqqwZM/T0AA4aBudkx8a+wYfjApEft/ERbyY31BVLeHwe/kj69FSJlIr30Q2Bye00m
SqjbrJPu6C+Wtu0bCD+0jv1FG6paU5dd6gJ24O99e3CoOjLgrSUFqsZkN1qua+hrHDP4368zMtVv
I+ULP3farm8xJemrFaDkhfHbEZ+q1/80n6nU/jbdegS3PtmhsaWcjrBP0NhtS9GUDFgHi7mwox0V
pnva2gd7bBx8s5LHSn8G+z+u5Q93yV7EBuJWy913s/MwNWQnSXgf+f3RHy2cOOQSd9F/lI+Voy6l
R+jlST7KbwfKxwaPmfP/gLwe+WxaXO4p/K3JOQzaMcsJpNl5HaAXf6fNlLyP8A0jKnURit2Ge7sy
EDK8YVmZj40z9gvGY5DhI5Pg6pB3C/8WT549GKGbsawZw+Wx/wAMOlYB2HB7bqUHmc1iF/eXbf5C
I+F94XRajihJZcMYHj+qRT4L1MQadplhTE7MVK5Fj6BQI3vgotepLK5nIbIKq37zXaxBypFQ0auU
+RiTb7IINcsaBMGPD+cjV6gss1HEdTWGVu2cNmIE/tNRxa3URgRS+L9rvv86d7Yo927Fi4AAauLR
NNkDyPo544BUPmnzuBz7+edXNj9joT9K9yl/7RgM0cRzO+jxwvfPSccw6byl+R1kkLUDwDip5qe9
VRlAzvCnRNziXaoQwJNCeiMVYZt/7hhbreqM/WgiuWmGI7/at7k/ZMPzCpNLZ2gdZWOlDAoRlTqg
uFKMOrQBGg3Bu/CZMDo74trUn1Ojsk5ViW9es4R+r7yBRxv8Zgr/8N4UdWiWZ4kPUQJCd6lpGy4o
3u2MBHPPag9c0QQlMtpwY3VNoG1NDIUQt/4qtEiPXfyL6VxomJG/NeMVwqM/IcaOyvZzqeesnoB2
V6e83+mboqbNSa1E9NN62o9azAdmpFj8mXx8V5I5rJp1yhKkUoASzAVamG0YQoGIyZP1C6KtqxZ5
PCXHuO7mgGPShy4QSwANkkbKejIMtwUwnYXWoUSbTyxXKh0eufHVWZQJc6eJJnXtEzHnbndqtDOX
Dng53+0S13HR3uylOxTgZU58mDap8SLbAcP3pX2crooIOzdFxeKzYnUKSA2djIidlekXDbekiNze
u8ZVOhsIE5W1KdSpb2VTeu1M9+m1L7DRO9+f3eKiPcuenpgmsQudk2FdrqGyjs3sJ6QYBumeWb4m
2LXfUGkRZiX9jKiil7oy3VN4w6CihsSbRPWh5sfW/qjYrBjaJq3zuwT2wPZ6M1izZGwJizvblKUb
AflweriVf8Kuh3gtdAmc9zf8pMg2HQcZ4TUP6jRgP1liaJq8/pzrurJbLDJ4X0DEil7aa1MidlYW
ctgxZ+L6+Jt7qmCRAff9l2sHYqE4jxpwHPa25xba41NyTtQhdKEwLLQoZ5mRYPmhsgIohJ+Ir3xV
4ybLr4hu9znoKmj0ETtptSisXfDRUOuYV1zyBPTr+1SHc6lP0kUewO4CWuzj17u0ekj+aLhBe4L/
F3C7RQAVonH/Eha5SnNnetSyFCinE4IeGI8k8uI3zvZIpDabK+9xjDXgwyeDi55xa8Qng35rD/W0
/vaKya3ldCLaQctoH2HDceFG08oYkzG/QTze3CSvUy03c/M1HTbnPyCiOypifTBa6xOmYyzvd3qP
UvNuGlSSEWMzKNnVuTHiu9b83P6c2Vjb+fsIm4A6eEuURIvbQLWFNi03OgXl0KhBjUgKqpuJAzMr
7/50gqxB6f5AXo8S1bOEyJ6EcR0r1tEkNwM3dlBzkNqZJsOSwm1l2vJN1EX2W31QJRm2sDFbz1eU
s9IxYEg0Ix3dIpFXRubx+DOx6Ka4+tJHI2cPHUrtxRB9SIbIJ9ki+LK3mk7FVz6SHMI9H/27wg0/
V5PQkV0xIyV8qTDWfrkGPvQWIJxPXmJiK/Ro8ljSJTPreitNye2+pNuO4FZ0owCdhw+M74N21BAg
//XfCkrJZ1nvctRVUMhvaU//DRfesVOe1XJOlG3sr/lbuEko7AgaaoUj66iARiRtUTrzfQsj/hP5
i22UXo3bymF188fT/f17Q6Kel4w0icmfJuHvQXIfW8kt0410Inz4MOAxhKmwScvdfSnxa32QPTv8
pbXzoq3Q8fEpJqNR0D1bsswvjBFy8k+XASzadkljzxEHsl1YIbv4TiIF/5I7wG0wanl9QT7gAXL/
U2qjpXZByrRIpVk35A8k+05g3K94Pea4glvwfEiEoWhfcOo/I/ZVn5rV8aug5CEeR3uakM3dGIce
a34+vEaH6nxWvMg2buCbyTgkvvcjUSmlnXtpboD2DNPnjBEzmJUELXh/VZI4WTuWZWQi+wmpeZew
nXLPWxhBZ3+03Z+WUSL8+9jLqN5/Qpt7Pc3ICvgcSr6EZOVyiBDH2vZHeZHGkvQdTSD/6oeRNdYJ
BdWaEhEPyqJOR2v8gjtjHh4yQupc4+7INNpSzFMSh29imGOAKuFRH9BRH3rzsf2lhPq7k5A6VWAo
KXxmyp5EUTKjQDsdM5iV4gsuJnK+neJZgSIaDfjsIV0Wi06hARJnSEklbFmB3GTNckV7jPrHhayU
p0aSQhxJdgldkNzQpV0+WlmnUnS7uc8P6QQknJerZCBmsW6YvqWQv/A+t8rc+3WDKHCEZfSNE5iB
nNExwt6xH9t+LC6l
`protect end_protected
