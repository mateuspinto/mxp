`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
Yx8+Rp94WXVIcs9YqQ9KkEtU59dZkxQrqFihSdpAugq0XW/NqdyogOtYa5+heC1L5MlosC4d7lKQ
Vj7cTBqbQ5kiP0k1gT5nwkQyJLf9dGfmMws63G/Dg1mQ4C9LoTo8TQCrOLx+p6fxD+a2FSq2WB1/
4jRLzOvakUo1+yd+kJ0QwWI2CketHi34B9aCsPIiGDgLHo84J+2xrHalShHU+V+UlxLQT3biTY5X
zBkt7dJsPFVQGyjAjH0Q5eL+sGtgvx0PSQjCo4EYqAVmZrv4v+V0qYpXxG85iTS2/3CZpJDSNxrM
GUk+xqBcjF2Cj61/CmJ0EYPLsH37+hrS2R04LI1ZKXQGwjCtLtc3rRaE8xwszFcf+RDEM+zWaeiv
4B3YfrjCwj+lr/WM2+ihOrhU1AlgrnPDJpCYM1AKg02CrP5/xumS8L/c4c/JEE2HNXKCrybpYU0j
mDBwk1Q3Hh+duKIX65XGL9Ag5Z4DAI0fYi3qZ4NxGEAOqoRGo1Ztz2Ah4SsTvZKrQ8nAijBKIjN3
WvdyqQcYShh4A6zgotI5zbgHTbfKv7814L01tFeGz1EMTtXAS+WpO+tZ3efcm4eQvsQqn59hw9rO
WHbM/DSozU93vqZO0N/RVJXK3DaIbPHCAbLxtYiD88bv6BNjyacTO72Cj+g2nFTtydv0JHC1xdWW
vsrwxDVKEz+T/qkXWZAN9n8N6gP9C1mQ0fMKJV6T3Meek8bzCg0VxnDQRpDbEYoNnY80xv7oz1Oc
6HyxwpKMrdJJ2TkNiEypo0YemxpiS/zsKLHnWQ/dvYevF8eF/ZTWoRr9SzSJyBOUhLAl4j82Nu8c
Xh7cO6nrDgJCQiwbbVjlY4SyLjs0qboiqvvbqwiaxRBka8h1AcmMTlikyd+zYP0JYTGJVTjJPLf5
0GtB10+JeB1jcDKtJSa4b5EKF+uFH0KKSenuB9QmPsp8RfgSlncXFLLBKfaoRe7Qmf2Q0q3kmI2v
onALhq2OWLgmOo6EvHnCYMXbln4EEnuxyzPYU5VC4e+ZrWRTH985KR2+HgUKxvcftqyt1gUztKb4
c/CAwCtJ6lqDSbo2orY6hk1cv5uhQ645rrFliWGvMxlUOCxiliouaM6Ejl3xGbGMX/rjG7PPtQry
Dz8hhg8rZ65ZXrpuriaz+8rjG6JPaULoOR94IMlFiK4frzCkv3+1c0uSENR3G4I6PxwXinDIhzUZ
JWlzGLVLnytJsGKbxmbXl8smg97p49K0SdKe08uW54Pb0MF9B+3Ba6tnkWOJn8+lBVegI6RH5kbp
/7EG+WFapAoY1Vw/QhtTK8TWEzJHOGykKnj0x+undNfLrbf4q7RfbWnZQIOlGOgja9upUQQY9tmy
3ad9bGr2DwGjm5Fp6kBtA6YggRKcxl/JYf8kSSzt5lWGuFANn62JVHBFnZCv4x8gBXWoSnqAKdWn
HOZYWdIdggKjQLzBNO5gB4uErOsjDyr0hYl2pxlDa5fPdc16WO29DlMGUzydHLlLRN0qw40idgic
mmJih9imrVGYzEejGN/QktEOcv8XM8XIQhQ+fosAxqs3gML85Ms2dei0JPOetIIjUl0ZcL99+zhe
w9g8e8EXgJtUnbew0CtoixRoSUs1XA1CtbPPWJeE98ByrdyJWWq8alqcpq68e9dWDupYaruznUSh
Ow/sw7oc14JPcl7DvHF8DoGaBDfm0FF1NcPPSvpdeR5L//v3rrqzz9G5lWt56g6zVezYV1+83u6t
MHIuYCHj5Ut6aGzdn5mJN6LHtAXNM+qBWfJeN7e/csrRFH3toLYDpK43FzokHOmNTcKBZeZH9gll
R1wRcf2+GjRXpA7jM+B1aOZsSBUDtY0NywJwf07LZDwEw9XrcaekD/7SpsGHeprYHZlQGCuolL1T
Fps+ClWE23s+Xr7dprkMGJB9UCqX90FIfHgsJOGEoDmGprzogAsQEXw3I0CBal47r2kQGPsqL/Ul
M4+2sLBM/lvV3jgGWWuaomu9xqOdRSXfQwtEFIBZ41W0ARylwiaXVyUZg37fiqCjzRxgj0pXr7jn
BEifoAB6mt4dD2JvZgtLQpwOdTYv65V0v1MXNIuuqET++6BlGzwEaoFJF6GDHM5pMJZJ9JqZBAbk
37Sa4yJKzyJs86g4Kx9MAG6MurXIvekqUxxLSO14MNnWPCFq8tVg3jkMSrg8qG4GhRu0DL6LEMgT
pfw4YYcPb86nHmHEIF5M6RZT3umhL/ioFzDnCsnPXdoeXrrjpbWg5yPPOJ8nJbGgSXYGy9sy/5oc
fntv9pRZeEhbbukCCkijgIDyYi3H8wZyROHZRjQTjbnOE7s4+Xiq35J30HjENary/9OsvVXTBXKO
PyXZunz0iZYBlse+4q+/h8daws2U4wS6f6Ca6+SjEjyMeOCaI8xdHtKG11Fe/It/ZU7BPTflgk1p
vgfoBaJBVAxf/KSb9+gMXCVUriabTw8avy7nuSuy4keACaNNm2dTw6iaX2ZdV+lwboJAdll/GbCn
IUHzveHrdPtnHeoj8pBzCyWkQ97hzU4FQFCxZ8AJCc6VI6IcNh/JOVoN/gkPooQ6yrUhus32cS2B
+kUobAgcUtErKnFFQcYJQPJeuWHPsNzMWsGzrJxsLsp1+FXTfuCalq/JIs+K/sRdoubQ3b8ksBf0
w1HHFFDbupg6ZTD3DyV4fzOwDBknogiqv0yMeB0SsINxE43irNLOvTe2CiWoH06umq4dpBe607gu
Z+wapaEq/ImXXXL0BQ4oOFoirkoZ8aCCxhyGMJixjqjGret502LzwMkxBOtgnmEJJT70OfD3jwUb
POe5/HpU139PIAKzQR4CbbZ/zYcGZUj0ETd21j09NDdnGyALls4muVAS6y4xZfHGA0Fqj/3a72m2
7uZNxa26iBHPh35FsRRfW6wwX8iGRvcGu1Vi9kgE0F38CXHlJnmMrIEZEKlAtoOBccsicQdGTdEh
YzF3SsSiYhmOxbhP1dToWgC4+Mv1TxYLZ1zTn/la/MwppI96oueLplmtwUmtmWptALgQHPryMA+1
eTYHsxJV5hnt79aJ6QWGSzltpIlZIuECUyJ/2WObnb/wDosY818Boo5I/pXbKMWVGpwMikUFw0XL
3S/HfTe46ZZiwiIEcSZV5+zYagHYzvum37hLEwFre0biJAOPkPpcKmXzXDv3p7Ke6GTucQvXzHEo
80s7eUpkp1qW2GWxw131piyZzoF1uuz4krjP4yAPwoYbE8x6pYd8fQxcVIf2af+sYlzaQo4C34j/
bMxXWLNzFzJG6P28RULQpH2m54Oq6Tat/c6ZOV6vHgDJ1pHrYZU+rKgzEPVPM/FQ0ElyYVrSMWPy
msTiNe2M6J4CvWEu9CdN2rKnho60THxxtgNqFR2l1lIOP7s/YsRnMOHdvdLqVdJxyixkkFrrxir2
RLQL9Jpgeab4GSIEiK8TcdK/gjzopIlSUeBzs7qquBiE0DVPbie1lbxxwkiYFGlNikVxlKtDvkYE
dFl1nNe2A8wrfUgVRGcT1eW88YviYnUg1VfCFDFEX/3ejqIJXUvPjG8KEMmgAc8uzrpj29XUBHMT
Z/k1/smgHDDN8zVGggGvAbIXVk7Iyk8DnC1xryGs82VlKHofkbwsSMR1MYEcmbh6GgT+rRmnrnn+
rfVnmfbIfjQ1g3bUnr2SS3LS8+h+yM/spUpKH7EBmu8hZ0kRR8F8tAyjhxUhlZMh7x1yMztzMDk8
Ise8yp1vIXNY8+mojTjKbhjJHPa+oLxl0p+WLK3xFEqU0qWGjyKLXO5vDDd1ig87J871vxt7msEC
SYNXaTW81RgV+XGSgekPUa4MAblGuTgOLyRTfoqeyH2xmkZ2g1YEAZqJ1AHPEHcLQ6WUY6lXn7pT
BkGyxxWlPmyQyx+4CU0EoHXxExTWwq2onN8JOkM1jsDDJrxBy/8UBMbvfXYGUXCMdXcb9xHcFZyB
YGwkhUopMAScbA3CJahUqBhBWBYk0Wx2yf0+EoWh8DAF7mYhN/Yqd5LgH4rBoOhvsbFWNj/d+7EW
boN50FC7ZD9VYbUwxtJAbnHBgyBWBMWryDg+pPx0g2w/epQknCxvon3l5WN0U/OCBa7p6FScYwQa
Gu/gJIQ9fKNgX0NSn00YpH8NPSPHS7KTRkYVFqEUenNxxbRmmxpTpMSZrVJ+4p5pecg+xkn3yKBb
qUDm49Iq5wrRITWp8YpHQW61N8iBBrTn/iHPm7byLEskhe8F9Z9Ydq6pw3mD46HvzLhFvvRn6URR
c8Yjw0MsNMEuavytM2wZZYPT0OSAD9CfP0qfr+24lxwo9SEDM6kRA3dKSRA92TYs9rjsxKumFKdS
DoNUFxHggDsb9tLdmk6hzG2Aah6a5pRxyBwBpb85lxYx1Yc5eIUBttoFBUFOx6UPC+RqxG7GavNp
xLBtZ8n7IkZITBgCM3HKpamuvPqsjc5VlSfZPPxYJG4VRzZGDvm+Io+x0a9NDLxQurI5Huo4JH12
u0F4thy+l2LczOiLIpkurjLntxMoUDHsUoAoEAj91fTGzPF2QAKuEFnyW5Tu8vDv2V5GaoL6D3hM
omtwBQpe7W+R8elqn42bPM9D9IFjH7jOG5zc91qpkgtDEBu2zXAgBCjFCzmwwPmLyeCX8JTTmZ/1
23K0qR+0dhYQtqcGxlCeVePKWc25lIEEbHDECim/02q/yxy0qE2iaEv1Ew6I0oCYBXk+U6Si7jlP
p8hwV1Dhn4gCkc5tWcI+shOELgOuLTkv2DASx3V75H8fTmTafO4VI5Qz3erxx5+qFLkTyVOvczKK
ULVUkMD26jvL9lKy6WE8Htk+6A88f3IhJoUBFUyFdVnF5sMJSdI1AcdUAsClLPeca4hRc7SGI9Q+
eRQTjPYtmitlHDQlXxXqw77Bw/jA+Z8t6i35KteFZpiDzUVgfnt4nd1xnwlEc+Unog08Cx3j7T4W
rpZXRv/tanRrd6staFCc5p/3XAOAgK/ndiSfduZxmJiQi4oVhjUClkCbonHKsb2nQUmn6cAyb845
Tv2mpxfkuvGYBNiPbDXIcttChGrjuyyDRcOqxc1uGO8uy9qLc3WnZFlpEfdmBMnvrIziSmMwEjk8
5hFlaBke2JLvLvCwLQbNo+FuP23lcu8UdxLRaoQ5EY4jFfyEq9LZxPPfNCBgnwMgOyVs2ubJWjx0
6xhECjWRAQzOgkOKNEIlRh5swzhoh6hIVS2RXDF7T5pzbzp41BANbrMMs6m+RvE7ptnGXmn8du1C
LXqoT2X9Ze+cKVsM36pVP30Frww+MSVhox4PDnoaFnGFA2fVelOnb12WfBCaxvxD8FKpm7PNvoEa
4QgcYyxHYCuN7AXhRxUoykzTpENQLm9MUTL5x6dJsyH9GxzEGdPxwbtEPUN6r8F8Lv/0EqThL7Wy
onUQFjQ1rd6FTpjfJ2TrvYFMktSK5riXileXXXZPztcxWG9apm7ueMs0K5w+fwCbIrOtK8VAm5Fr
kAf9skZWFwTUH0OwWdICi8SpfgjljAS88dAcmZPCMnRnNEz7ULZ4aL72NuG6NHo2yjnVQYk9ZhPK
AstQa4jSEB2ppFinBNMDXx2IAvd+EhUNrr+GcvddN1P3pqre5xck7lFff6lNc1fVv0RLORy+Hx/d
iUQ05CVF6wa0DFFnny2kxzqs/npY5zf8XfzC0onbAT6jtgqMm5J3D4Q+/BrGaWXutcmKK2fsS5Vp
7Thrsv981XUu/gu5BdKjzdVbs936pZkn+XZzHT9/9qsfR5qxVjA7QS7w5p316Ukj7ZAr+mnTubPy
xjlvcAxUktQmAQRMHJn9B6bHxCh34oAjUkmsEsslaW+4lmeNvBMTdbu2uTtZLbKinraA8q9Bq3Es
lxmXYKMuK3/sElZMTQJoSP56bgS44f5BCm//d6rdaHheF8VnXgDmcF9QowZrvk7jNkb6jhDyi/2g
GddC96k/KnpDO8EFGhyUkC71KI62hNE7c6+l4CbuHhXahxSLjvWEG3Qt62sRMrRH6RckAYa8r5T+
aLboHE/s+8XJT8e3vPW7BzocrI/etheC9S0qRacmPq8nf8hA3trhE1HvAx2w7kXbsaNbFLkMUTHF
G4+cpvprMjewZq1+6kTlWe/s9h7M8R6dDsN9AaPgZH8gftgAlqXQLQAWm8dOfObf9vjj2ekaLqvy
c3Q9PfpPPOyITT7d3vSS0cXbmP6xePIB7gvTjamrL3jwebaGpvbvkEQoJY50Nyd2mTAjAQ8jlmU6
58B18IwPbFIhvfo4weQtulWKVVvrT3Fn2L3aWIhUXuQIYadW6LXJjiSAZIHUgkz48sxnM9Borwvy
r0AdF9IcpRnRZvjSXCpHS20NtfJXYdFuKnOjWjtCa9GwdCVtVmf4MFF0+yAW2LdQymroxW08ap84
l2msU80SDX4422nttT59I/IUu9UcYZgipaPn/NqqcYbSC3iGkdX+MyiAU4rpioMt/qk6rfXRXFpA
Gw3MFyYWJgpU/Dxb+vz+/Apt6rCajw01kQC1lKphiI9GtrMPiULn1xT5dq682AwWqDnb3svOAOJF
fNlvdOcaNDD5hcXDhIVGXuU/qS9q3PDxsoD7uBm6xzjaD1Bb+ZU5FFHvPitbs9sE4GbT56KbRkBs
9tABhIQ+RPjj6Gxni70aYtxK/CBmM6KGRn8U47X8EEh2FcVBwKne+R2ofjw6OO+Jdx7eEHHdBUfR
pRqQGcESluJOyGAC5pH6stweshb0VWGLyTPCdPvld4j1iff1mNWezShUVDhr/qoQyoijfywobCkv
eVkgiPAfA0NHKU4eQMeiGVO+i4duCWBnUvmQARSC4L7Nw31z+IigjwleX7yMEfRvFQbVzLxBI3MC
BbUUthSwUL104B3KQje5xcN+RbXlXZeLbRVfjDSD2WgcSMWIe86cGly0C8qfOAopME2biiXLNU76
t+YPd1xkiUfMPTSASxXS1BiwBjPgoinuuYIDLnFbH0jxl+Kw9EmoRG8p8FMR5ytv+6pWiTf3894F
Tyd+ziYLtWtubCkC6AjJN/AlPb04s42ayw10ZrVAmdthFXc8htlSEIuQReL7PpFwNzHJprxu1PTW
Aoq4DGxTp8EHnlHdZQG/6AQZ3FmbvhldHU9bThwGGSa00zv498ZrQFGzA1RNKgZqHGB/rxO8TWAT
flaA18NGGPDvW4Ya89LZCQCiSSM9J/wOchhk5Wq6T6010zwiZG8kL/n2hgwpwZXWRT04jhqDMJmS
ExEqCVyWgn/dMVWJv9scyFkaKoL/h2XxCphvGlBgDq2RxEmkvKJmP+13ngr7l1H0DE0XwlUBTZy3
V4iURdF4pI6PnxfELJbqS/VeEiJLWAkheS5RIrzNfbN/zD0pBKgmptXauqEtTcd/ikbwCG1jDjJu
KoL9WJ4N4BcqAtxYFrzOB0n9j/4ExlRY99JR6zy34b+jFcFkw+QtqUPHmb8XeFCbG8rQ02trGY85
PKo7JNWbnDbDX7ry5yPQp1FjxP1ZjBsgMn2B1vrsGTvmDmZhj7cav5lQqz5VE5ateAqPOgq1I9YY
f15gAJoEIreoC1w++abdkBc/diTPz1vlNCOpxaiYldvX4HjllC0MGC8drqCyq4fZhQebZg/V1H3U
ISeDt4T9APAjfNyOwQsHZKmvQnQ4UyF780XJPa6JWPQCwLpFndqbYHWOadrUHHZ+nZRoO+rkAdAU
W9/io8qymqMs4H1EDV17wzoZMWG/XfZT9yxYccU71xn4x1oxpvOAmMuRYIKgvecaqoYfNXEXERAA
GQImU9HC250aoOywn5MWHQiNiFRYMZzm4ClUBzV2g0fHWPUbGN+BoezV6DASTD97GJeSom08yBlH
qrW7r7lBvhmit52Fbx6Ffe2lie6YgnUIvlP/eqHokMoUN4iXv24HFWQiq/xJCnFUjw80GhwJWsDm
1Rv/PlJ23WS8QKGFS+JZyF+TgxK+vWQyBA2uWqhK10SDE9/a7wrCLmqlDzUGd9Ek2NjhGjo+VMal
K/2gA6CNaaeeaXMn6FCS7ZQOuJgnMYk2hKq1D0qLCVcnsSfb/u7uatqHqAGf9gni6IFClle8+fLj
AioTw2/iFEv8rvJtLP+mww4JqxILswVU4rqS65D2RQ3g3JJrUx1xTSgYF2wou4W85gsHJLwqE9hN
SI/R6G0dlArSVijIySjlD42hDQ2D7sM2T+b5KC3RV7nrnlSU4fgz/IJ7WyHXz1euN2SS+SKPEcjs
A1L8VcDYaI2+KfsdfmH+4vyw5oZOR3UIRvWBVLb+6Zisr2EOvD4znQs0h6gRKRkktkV+QoIRlin7
GmbsBvhSGIqmF9S5vXU/fLHmomLqopFP6TjzYUHaxkcZxBdV7kZpk28YDt/mXcsWVF7/91BN01LQ
QVMWazr0BtF9J9NkwPjFPHrK7Mxu1zCiysuoy6rvzDreyNToqANeqaWTscgFh1R+ec41pkIDEl1H
iUs1UwgCpHYdf+8ejKSJSZ+UL9odJAY3RdlqCKqTxRgWmgjOEt1MVt+aDQZPLE3M9axfuwWUhpxs
WD5qPiHsrv6BlaQEM2+ZHEC4NX87d/AzENd6cwUZZ9PSXuKvoEgOfReBoUpAzUQtF0nmf2L3eDkN
Nov+I/jUM/WHkIwuzsOWr+KuBCoic659+Bo82yNUFZcL3KWkkg+5J4pDVngOZkJS4n2fpdVL28mx
AIBXsefSiAM+jidMDZriiqZbD9wuLk9UP5oL3Fpwb6D9j3+/vlPwAQAjSVQ61geuaaVTFy29wN9r
uQoySTLAjj8z16QzTHcSDat9ynDMU4ittO158nZMC4GhYmn4yJ6E0g4DIgsdBwIS/HNLaYutqEAH
rpYaTWEkMx2eCH71d3U1cCBZ/Vjy+G/uo7EU70peNpwn++naMq02NIvgtnEi4n+7a4JOYH3T3kci
BR5Go4e0hZGRqHVjc7LwPA9n1j20tVWpJaDUL1w+8gwACIEy78hxyD0nhekMrny6j3XxsWQVy3Ed
e7Vn5XHz4999QDFyi55EGH6Ks9BdHl41xG1Pua08JOY7yoy+k7MbMaXZdW0cfLI/u1djasTykrkx
M/AqJxGEfy46RnjVvcxa0DzCRaD9gJo+P9Y/3l44nhJ7qhuoulizOp5X2HUeXLhvdJ8fKFULfyJP
o4dg7ZIDt9xFlUA0C9h0xcP5nSd0hEW+F3/l/KjwEJPTmMW3SQhWFLpeVaKr2NXCFEDdK1sW3N6m
L0DrLOUdFETOKgaQ4Sy1MggV4yQxxdv1YDsXmyLH3w5iVRCrHv8LbEmtXDDRMl8cNGG8WJDxXAXK
O1GLOjh/FpCzEGTL6pkviW5cS/lAsBk06j4ryniZkgH4PShNolg9425pC2LWhAE/hckK8f3g9hiL
L2WYnjKs1c4tHgWbYlATPdqbMDfruFCHUaK2DeL4oRmdQiMHOaAjJaXBGJRK7AHSll/FjxwkoEwO
pfVOslgYjmfCQl+hZOG5smuG+p9q4uKENvj+joxFEnroTMBq
`protect end_protected
