`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
aF+vyFT9BoQNXIut1cySL26fm9avwzs/s9FDNCvL/Lc3MlrUDP7RR4jF2pUSaJBBzz/0e2MItg+9
DIGUAM5ZKl+FQVkiKnTOKLih9bwmVUxM0H3AL0q5mJuyksMbXng6uGqXI28cTz4xdNjOOe/IvqlB
esxLQFvmwXUCYxhBs0GHRJnD7UcjBbOrvqZX2doR6Eyu1NBL2sNxbDkjoctutC/e2wWznMi4H7w5
VHoBJS4bF5B1gnLDAsIToa7Ez837UlrW2Taier6eH70HnHjsJyap17hkYpreknBcGUmUlmNPYYq/
JzSYhCUJ4/Mufq8c/tAYLghLQNLzTxqdejAasI5BH1qcZ7g48/Q5RHAlDcQMMwo6jOR494sQQ+og
i4FA2s5SMh2tK71hbY4R4fdLyE8s4HEm+ohVAVVYG+cRyEgh3M/+YWwQ/oADZYAT1ydTqGVT+w73
QhdDeWdXkEUhZSJHeitC8ZSvE6Q1VPbOBT84oOGHpQRQ5uEhfyCqvzRL9O+YksTcfaXZMOKgwSom
5ljdaULHtLVwtHt0tUd4L+7I+/GwiKkQuJLcMSN+gUllIQTHZiMy8stcS+D2keKDs7Ma2TuXKRvC
IiaAVbGl1zr5M9711Iz5sxCEbuMtRJWYYyla6Q1uq0rSGIpcR6DjFxaXP46ixErfRPTmqh5Czm/q
oEWh9zCJobKfC0kcu4+hxZOyCgpV5nA937BpDJoEOpBTEjxDF8o2XeTuey3VlNeydD+RVW8NpRqo
wW8qDyXUEv8iUV9awnnA8SPBHy9VzP3xU8Iu+Pm8h4BdMCU77OBB+OApSygvcqNsmvBUu4X1wBpr
6T08TQXcscI1f/2YoYo7zPIGk7WV4Yo1IyxggITvFHDP5VOLv/1t6GCEbVu+IHBJm+DBeJPt9snz
r/P8/VAEO//5M/2E45yHcSUkezO2tDjDo6m4Gche+SiwEwicfRnhBD9ZmSciC/35hxZxXn48nXHN
12mhgxWh8RielPOPyrWu++Ncv3HRXFwEb7gLXHlZ7BnDdStryycBWWpgBxHxWpnbekK/K/uNevDQ
HHMFkAC1tZi25IhbdT0Z1/FBjngCc3mdZwy3I9Se3Yqq+PgbaGKNEEP/t4s9lhlmqN+eEWSFxHiL
ElnatKmJQiKSL/d5/SkM7i9BsNjSJqzU4/w5EzgnwH/GZKmsliFxLspgIbIDnvdBzDRBEW7ZZ2VK
4islbPL+g9JS3m8rb7fik6WVSo+eZEvMx28f0xdgHOZl2eCOzjeRSKp9WsMdNTHBSt7o3iDMLhI3
IPNmPG/nhABGc5f4URPcPV+aPHsooltN5g4avMDkFJ1RoSLcWCYLg4FieE2Jklty16lrNKP7OYsG
kOCI2NAqH7Ly3W5jVJSiRCBJX9K1pQA/emr3T3cbee3asNK2p6arnfZoR1hARu/4O6cTAlxSBDPq
onysVRMIvYmcs3eXoNTPtcz9mAJdbspjQEkUjiiqQsyOMxNDMQmtOTEgfJpxCJDYQGxCBENZRq0G
6k9kUpKaDECbz1VClmXun+StHAcj1yGucwTgcc6ZZxZt3xCnHYCCEpQxXptf5WXrCf+CcC1413kU
r1zBW3dgcxQGci6b1yL2YbOsNZeWJ0wea5OnoAX1x3ga1TA0+1b8n+I1tNepNZvP50QEqmOzazrZ
EOHISqoDskIrqhJPUuiE7n3EJXyteOvI6X2GuiOfWNC+ipmTIEkwrEVnhmbPkU0pfKH/8phigqcS
2wh2ZSp99OiAqksemte9c/W+NagfosI6O8ZcDop1XyekxONBwulKJgZyaCaoaPvaUMujAhvY50Px
rJ737/vJ2GqVzrNQnFiRtlSPISUbaOFdSOYZ9N6OLuSvo/jW3kJN9Le9VscW+4MjnSp4tK3Y4rOV
403Zj7KmdMfUB/h5jmkUVYItawTCKVZH3Il7z+aY1Ek/l/I/0/mmQVVDxK6OFtzuQP5ez51A/M4X
d+E4ZSpd7YTcsEl3hpTQHIXxVcd4ikXPNu9IOLMh4ATwMWspgF5iiTujeJ1y/JYAuKjVEQnTDn5j
J1wLkl+zPrktUVP7wlpShrVLEUA+y0ThqkcIqVQ2OJKHVFfIMxFMfMsWAid177OsF8Fy0YBQe9iU
xQOsK7STce8K7xqE5NWSfjtbP4VR/wFyao2/up84ei+M6IGEXou48mDIf7fgpu3f/HaRq4m7QUCU
+CAi54dRObJ2fMlZlAWl5oTDIEqGASJwwk4by5LkpY4cJVdWbnBeBOQ7ahsaOI0gdlxXfWH9ISEw
X86wQWzK54t0OqeLADWs9ZPgHXN0jnfGZwouw9oCBWHjERahdTsGAOigd7fRK5dyapRpRY5C7Ev8
U2b3VU2x/IX9OFt/z9/vhsOObh/ScDX/yNbDXrk4/MjxMPSMrMRJfNyOa6WGFsdqUt3bLqEyfcDE
hs0JtYo9Na6Z7i5WLodsw104ItYUqxyxWqC8FX7pP4Bh+RnIej53K3a9Jh1MeQEhp0JG6hbMyeqt
qEdwh2OWfK0CzyFqogRZFcSd/cJuD4SDz/Em9XgeDs2GIDFUnz137bGtIOPkMhmn4tgFPMPqnbHA
aejVlspSbujgqBnIFedzmYahGM6En/MaMi4+upXmCm24zZ7mKrH7Ra3PAqWGVHkwFrQQRuQOS30y
WFqkSJMmONGDIMnjiGtbdwakPUCRAUZoTsTuEt1iNLJSyBUh+1jXdXXPtKtfqx+3Lw6k88FUOgxy
VTtcqHrf9MzkVfhkQ9aOjT3QBDU1DWxhql+OUrThoY2AwOMJ2U4ftavaQ6+WKadnR5Dksd2ieLTl
iRTqXqHdhw8fbwAiO4Qf+Gsom5kW/CSf7Ujzz1gNyR9QO2DcHal4lLjyQqynuA6MGaQkCPm80Mf9
+tjxnN1kFXR8EB6sTuFvMkvyt1Z+fxPMQL7JT5nrcyTBHUGD9Ldqh8u+cpbMXWnc8+pMhQ2Q4PrL
HVFWrU1SMdwJ6IFhJSU421shjXkjW7iuCVG6MFg7OZ5D0eojuRY77tVhZVjkuj5p+B1KVG28A2GP
UFOkjF9Wxsz2tFbBeIX1/artwl5kVXa0Ye0Fwju0SXFNK8n83yfbAHcpe2bl8SWBfxpcANLEpofx
Z9NRmz3x6hDYDkZI90dUESq2baM5z9hDyUcu+mQRBpBTXoGpmsrGsY5w3JEYQv8Y0pcz4JFGun27
bjhw9odkVWvTDE2XKVyh+ZSxw8aDnqE8/eTlRMDvmsqoKF/AVG8/WVaHSN8jJM52Y/wlzTbfKU+W
y8AZlN4zDQ4NQDniTJfUygZUqHbmSmQQEWEYMtl3uJHj8JqoBxtKB0gsEBDNvop8SyPhjf9k2t5h
GhZCLkGJtDMUVTBlrIcl48gI1i5kyiv6OjpHtUa3xpTqeH0kfeZcfY8q7sQmMeiAn+FC8RyVtQWw
hxJ7qcrkUIZUQs3RvrkL4ahnwCQ2gS8tWcI1fhoYVUezjHO/Kjq8LupVHy5y1bTmxkoKjnYO+lN3
rOpBe8KK6ZCwSKURz32OQnu2MmgFqWMQ1u6Yek9fzxmbNnW0chdvKrylRpKBuMgHshF32MaYa15L
B1H1a//2NhgkQ/oa+1vJ2fF/B8L4L357AW3Si/xupvgHGgaYhXYJ5VEM10HFxxnVjVRUUDadVPc+
O/iXkSg28Q1MuSgAYm7qM0Kr3envfPxj13TourV4JvXup3mv12ApVGbRMPSQeQcfIrI+VpD5Uxlq
+/QsacQe5/NM2QFIy+tkML5AxDAfxRYBfhGb2DhxRdMRzcXQvmHxuhRfT8rWcFM1o3n6+kpbDIov
5HeKoE2RIq6ya41BHT2h/Oz2ylYuyuxV0IXejt3mwoSwChw1cadWVjMC/tf0FO8Ws1l7u0Rkhs4m
Kfnp8AMkilfDoy8wYmaESJqZGhJIMarZFStH2NTrypLsN3CNbNiCLOIgJKZaBwo2G+sLsMwomeE1
3mwjO986Gcum4fti4PZdLdUnJ+LJHWd4IldIKhedf6X6eOGuc3dlx2xjDf9dCCg2IEOAS82GumbJ
5z2DljZNO68EMlJqcQvi2BHhC8Zn1kxG8VjlZrHEJgIo9F5FEJYQnRRwz/KND0PV3Cl79WzB3/d3
pD24lFCyH9ctRSZdPzgvfKfojA/IXZCxh09s9f4tqxcaMWm1RcTIOc3w3g6g3ULiPz8qs6gVRt6V
tKTanS34e61Z/pojjI0NQTlQwToaEtkjoKy+21jnTmnYk9BhE9CEDehPua6mmqgtNqMJ28V2YMYq
kNmmfTq89fO07xDHLnzZHX1q7CdK1FCDY4owZrAJGtB5TIsI2HUW/hPu5fkqtAsLQvwybPXxAOSc
wgL6mONtJk/FRyd16M0yNBCuNGlZoAHbRrb6jgq7P9rAihoUlraStJQCULCOzXWGIsmRd7c9g/1Q
g2RVy9hwbG8R8GoQ7LdjrKvgQ55odhprr/LZi3syMMcOMm7UvG26ECbC44u9vazxxARhs91rGdJN
yv+RYXAP1H1eihZzdCPI4j3CYgaPreLeeSuPEzXDT97PkO8lu2LxsyJxqS8fFLR+cWiNyeJauQDB
eE5Em3gpEX+Klg3cF8RA9Uv04HJja1/loBMbOegeb0zvjhz3+ts/zqA78CPVUWJFuhWUvN4+f+Vp
Zye/GRzpqBYSr7pddulvXEFKu/Msw/53vYwmGxYaQNU9hjmyX03LEEjbsRjwdvoAtF+rZ2MyMSIT
ZB9ksikwbP2zf8Gwj5BAMDeaOpH9qKgCLevOkrXgYYNOFi+pF8vtUVcoNlzCLfm9HtmoWMcN94cB
cKbkZB98BTyRwU/wftxGvoCetlJf3cNHOFrwOBEBC5QFgX017rUrmG/l6p6t3wxayBeJhiCt06Sd
pturdafNSd20gYBlDuHwVVmJuDWpRXPCtXNW74WTtlD2HUFSPwIQ7lDQ7rCvSCNnmJIfikIKAVG1
ng35cOYtISN9eiv5GOL+obUuOUUUT8ZmI4CWr7aiARlAVOSg2VtJXH5NyjO9tImBPmZt9gCGXX2G
XhuWqDZ+qCaCCTbr/TwA1FWqz0lD++V9dTXbiESVLjSlY624o+de/hNi28/w+O8F/Kp3+2gDVcO1
wMHVMjrFRjsp8moVk//lBarbVtfrl7A0d6mlkMUTVOdxu64/OG5VsHcC1CQ0bqJ3VXhlsRu1E09S
Zcwrg+xzff2tICP0gvnuZWlpCwFBjYuSaa8rhE/RFm9IG2rP0MpSNmCN42luf+QQXPIvmDFRJe4A
A0bAS5uW3kdX6xzHjy1Ejl8RjqBcL7VSf0Gw4IqZKp9WduQSRtmE7TrMtlGiXZDwQ2eu7/0YUF2D
dwYAqjfPSMmH4KbNO/4HXTBkzapXBnekc1llbj7USuC6QxPqXixoYnuZvSbmKoQElryLWGAeXsny
YFdBfTLwDc8WdRVRAdVh0uMmnzvV7HRH4cc/6k+xh8s8gdPQM9IWz174TqN4kvwMtoaQY8NAcM+j
zH9/6HOx9seId2hr0PUoTEUp/ItPrEZQ2XK4GO1Jbqkjz9912YLUNBpHr4BZoiQAeLWJJHpRLyk9
wOqGlyPX0+eEuB93xZOC9LtpeZDLQPQSVc24ZVJ8fmeuwRNdzz3POZMr1OoadnNtd2LfQarBrQg+
QiGLXF0nWfIian8NhRHigX/0y8t0FHC+28Q2v9+CtCnnyMIt0zW2UXnbtgvufL+VlAoagTCHuMNJ
JI4ACA8bjkMxscewx8PLHiC1Ph0rr9O1HvXP/7ZZU0CWFDsKWA9rkefhcZnsHPWknreFKxG+rOe9
7qysw+uxdDhT2ukVXNa5E3vbKdewQVlu+HnDAyy6KFAgF4+1hCOOixWg54GDzymcfyIxzNSFansi
GkdAZplqqx/Fts28/4iXnAqzH1lt3Xee+gDVjhbNap+mX/40y6gddo2lcc4tv8+8suV6KRSZcKDK
gUMLwKCzBQ0RW+c06gymEhkyyrgzJo4qcB/827PD5Bty+2ZBxbWk35DjXbkjFV3SLBrD7Kkusmwc
9BMZ+y2obxzur4/QFSXJtX3JDFGNjKz4Mzi0t3H2A+RLkcdLc5609ZeM/fqCSgo0io07Uy1cm1PX
q3uqVA2N5YfJjItLq9gWwht4ra8Pqc/nei2Lp6FNqJJty6QG4oa1b84r9skoXhT1lPsXz7jRKhKV
dSwa+z/Xj1VlQIH1txaf6M3GftN0tU4uE9tjZuExNwhV60j0JFUJV6+dPM/6R3rGivfjSS6d6wGV
mAgM0cONZ1CJrrWq8IEk2EQR1tlY55Fn8vhQdVL46kuARJoXlL3BcnTqkAVA0Rg1WUI4HmAhUq31
E+4n1IuBmtm+rHg+cKxd42aq55o9IxrVjV+OlwYUO4eAd851IzBFLdWg9mk5BBeLhhCIHxeXVbD1
1WK0GLulLNACQR8vS67mbQodt8Q65VprrAL4E1G+zbWwuccOE4x3e1mUY4dbWyH9LD30oHt9vYWf
BmiNh8SLQ5/AkEC8BQwZsqzT5nYp8S/E2bmzfO/67EShp02TbGqw+JDZKf/GYp3b0mjLzseZ66Ib
3DBcbtzm4c06hpf/ynCgoJcwBpFv/kvU78HRNsMKJ7cgcNPASRKZXaEC2fv617qBqVlLJErgp994
p7qk63nhc7DHJ5e13c93/5MqyrKqf4jlJ6gh0824CkeqqT9woMxv6TQE3/aibUgLG15Dvy2Fgouf
B0aW+T/CJfASSkeDjHtA2VdrVWsyPBegz6O30aojUyiaLeDIDWhEVuq12a6RdHDG6ADoAIvY4jCV
U8iERrFIafKi5LgkcAYl9XTnY4Qa4wPhFTSECdXTtopBkPKV6B8lNYGLvCtsT/xAEDV5yId1qGep
5CFRRfyWyjJ7isY2a5Q4yMFpRUrDn4NBz8RsKAlR2R5horOL2Lw7I8WG0zv8nvWfFmWdCTGxmeAo
w0KV98Ro+DTOAu8+Z5WWpz0BydUMcEbAsPzCcVEs1MDADsv0fUI0BjlYIOTaxN8QS7hW6h1U6sGF
0OYmyOHQDYTc8hRb7Lxi7kfMsp+swC4/dgFsfqDCKRA1QGAceFTg7Olg0lGHOTEZxpOXqJ7+oKBA
nmEI0+Kz17axF14hLws7ytrB/Aul5KsBv2Du8FHEp3rlnJOl4N3WlW8j4FJhwTJxmgvDBEMXUSY7
9A7YsBaWy+KrrZMwlbrN2Z27dD9avYpC0o9fqtQ0KP5wq3J75Jz+NVagQnwbB45T3mmIeUAy3XAn
YUYDIBDij6m/ZaxEoZTU203e2EFvIxSHdDH3lvZc/tM3Ix5O0gXisfzLG5BXNkBHePEtJDkzD3Aw
woNmwh1fiAd5VQFFxbFcjnt1utEuNur+uU80DlLomhuJIFoCV5bXRFOug/OIlzsy0gxl9eNyF5sY
czYpSVriS1JEuQ/qoSBd+BT7KurVbsqlgxOGbBCN5jZKSTQDPGb4HPfDgmmBtS71Hj2fiCIVy8uL
lx0BH2MWhdUsoglYXnRCNKe/Iswnuh9vvNOKmrmKUdAZUuu7wsutGjMIn6w0X3ip1IX3xgRF0E4T
hRuQdx0lP1lb3fwOdr4p5Jxuidlb5CpALNPFJ0hwerfpXxTQOeUfXbNiFn7XdfCD0/J9gmwIqhsv
lgVFbfOBtAPy21SWYadLbPk2tmuI7H6Ix3/NaM4lYCFJ/LV8WW4yZpjeY99vjlXDvASTKx1hbMH3
vireSN5TWhrsoM7dNgBxOsIYisL5v0AiSaHFMMThBRXbJaD/Lud/ERZQCnNVY1oreRALtIXqj3Tx
5ADE7dANlw5PEhTVRuABnA6+EqNGb5qCzlrgEOtRPYSMgh6KD/eh3SPcDnxitsZirRrk4gn2C8dF
Rub1tLATih2ZpK+6HDu4f4c28T2xZCHACj42I6m3W1XUNQ+/mdNnOhiaWxGUULp30iDkFSUYBQLD
iRVQV7A4MWaWzlgnfhXMXCHgb/liJ8HP0dX4R40TVl2xPMcT/jLgohH+ET2xCgjOeV8yso9+kazK
AuGRbWIQSsjM5xwsZFKWbH5Uoc4CcA+qEZbwuE0g8ZppIdHO0ILUm5JC4EVUGfItyVYJy51ccW3i
SmVWmNkw6RfupZVnXe+79Hq5+0Rr4vEwa7OadQ5yyODN2sNBUeZUmZ1XXInobocQGMUCrhZvSxY9
IxV7R+bS9wSBmhsPm7lUznLwvi7/nmGhWS3DUtyhxNZyrxszue/wjuZOeJfu3EbEY9yROO2Beajn
33NfHfo5pWHarHlr38gE67a9qsqZyEVtKN+65rVdEBgXeCYISyZVM7cfe8vzdX9fp2aDr49Asm0o
F6pWYSuzOMPiKLlXyb1kKrSLkJAXOcru8Ppbqn0q2NX6b62/hMHHerhT6hUEPS+4f13YI9gVI1+k
A9qQvzJtBmln3M3zsKBnrG8HN8m0cJgmgBZmcWr28lZvALD7yCif1NfMVFFBYkJb1EgPDJrixhrs
IZT497k21VIAC10rbq+2t3yIexs71568hrfaCprsHxWkKKZJzLxbM86PictjbIBKqnFTa5WccdYc
lAbYGSpXWL/kMpiEQNLgG6uQrBx4uRLJyhJydmGsqwEtV0nz2Zmxo019GtK38C3D57DTyvoTp14X
UppvHw1bM0GD/aXcz+lP692tMhmwdK2nBng5uT8J7oY1diJxHba8PUVf3TCxb/NvrJIdClkWnDyE
ALZte8XB88ykWK+ddzs0QEe1cr2Z2MOHLojv27OXd1sac85hlgem0HM3PbG7ZaIewYsYnIPExVXg
jcsUQiJhkxdFukE5ANV3rWmAeAMDV0qRae7E/ZNnGjE4a+CluCyXCm7qlV8ON52A3w91KerZAiDh
HtzbHVLR9SAzNa0TpIh44D19j8oUYfys2kK4K1FBQYr70e25mPaahjRmKCZh+ipiSKz4et7ex9VT
3SCR0jdgcm9oZOfPXFyAW1+tFaR+f/XYN6SqA9WwBjEw4XowLe9B5Ywl4AfoOqFV9TcC8WgWACv9
bngmriZvOA29jiMB+3dTkGt5mf+Es4oVPi9cC/Vmflv4aTDz9m7EbC14QV3Ls3jagSQ979SNvxp3
n50LdbI/CL9sS5NDRFcQcAjO8Zq6dOXU5jmZ4eKbc0YnHrcMv3KxmD3h8Qb3V4nLdEThwXED0Q8Z
lsAl1zGTQyki7kD5ch5N8MAua7+9XbYcy0COSoK+AM3R3+JgRppMZ9z6T1vpfN3AZ86H7T8D05rr
GAyaOrvKtXo4QDFJi7tzm8vqzTbXHqldlDgAiuVFAjC56cAVy+zTTfnipM3CCX3mxsJzCikwnLqA
mTkfLBqkl4dQsva01HlVUfbr59TacPEtpqCIAa0+SPOJeK6YfuDIiEJtT/rO8qocpc596/U7zBhk
OkPj7pp0Fu7O9ZMB/mcxMvEITvxrJqOJTD0kMA/PQf/HFDG7Q+z3Oqin08OIu/TP0rLJB2AtmBP8
cgkfWfCiQQYF4TlbSNKFSXaYoD21HIpRSeq/jgrI7lfv7l5IvsmRbcLiXf7rSx8k0Tm0CZ9alSjk
XzOec9okCSBZzfRO9v1P8ElYFvYsUDVZ5xin6NCd2TVSyVspzG4WED5feCVMOjZaH24xe7odsW0q
zPMLPqkMdh/EmmrQeC8jPA1WGVBZpXjlFOdscMtiitn6EVudFavpqsylVjRRSMrCICLIsWi2qtcC
s0+ZFat7n5Azg4ItFAf9E8AMyvBesF9exLZ14R4+gEmq5O264gTnE4syMIvttEJFuykN80rnfJ//
N9PjxnYT+q+YsUUbPkjNEskZOCXo3Ks0arnwjXZ4Pt+hqa5hg4ZwxkbwsyuqhRYXeZtyFzNeU+XY
eeqnRGOyphZ5diQwjnBMYLJ5mkFYh2BH8O04of2xhlFHXoH42yVdHRJV6P0SuqJNkvB4z6PWmyy6
FY+kJeDFNquL811ja2Y3roYJlZrFf9Gx+JRzKCtq7/DSZjLFnhq/YJ5MP52JuOnrOqApw2OHnHxF
pGS8RliGcTKkImGesijpxlksZNoUsD/As2tTOOdGAoA1bCpTqDuyh/tSHcCFnNejuqkizm6ZnruS
pRd36nfZzSOX8Ix3ej8biu/Fps25Jrizu9rp+TG8z5Bg31mJn7WrU0u64SUqTfR0g5ul9GRURu0N
sZIyU6LMXCkn+RVAQOYHK1NrqunO2P+niARv48bDI7gpJdy1Y5oXDhtDAGubkZJdcKQ69r/I/IOz
u+5Cacc9Or9gDcTfVeisE5szNZ0PK2Tlh+JqLFuPc7GG0D+6jamMGT7Ll256dwybOk6nywX+iyTj
vO5+gth7mP1FejE2K/zOvDHCAsTG3AVlS1EWjX/6XGMlFQNgqnLwJIunOqmC/ks7NwpkrWaxowKj
/CgxBdMR+8EVGgkj0zqHkPyEahGbHB3LIh7FUiNclTA1D3DQHps1LX9Z+M61n3B5Cqvrlnl7eH5I
eJPiBBrOozEiAX1X8p0bVgX4tNOtvgmKAWba+7dm+3Env1SQsqiw+REmehwoNYld7ombXC1m0EaJ
cX+QYgrO0oA/XVruaCdAvbmZE4KbLib1+PlDyf/u84woq53nN88N83+gwa5g23tmRXLZGCzJ3jhS
UHhsGZsBqMPEanrdwa/5JtmLydXu1k0cue9I1heaJwDAzkIjDjzZphm/zlvTz5IVOaJl8lzf/XoN
QiUIIrlj1Fwncr7WNgtq520RIC3eCs1HOJFqdxqQ8Lge3T6gKofWoSN94KdAcfCpMYSpmscmRa25
XSuJoAoG2nDh2x6uy7yngnK9qm+np7F5OXVp4utoXxx56R4wGE+EacWksDhRXsZ2snXF0s/T2jGz
WDrOiz6ilgv4D7hzza+HwladsI8mRyAP8krNU/T7ejJgFQbtPEI1JyUyVogWd6Za4A8uKRkhZQlq
8agOtXW/qLUTeaq9x4nMYR+hpJ6BP8wEz116eR6i3eqjI/r3oMYa7D+xR2Xp3itYtFUbO+C4H0uX
7UA9dBpZIZYbOS+5aCN5bwtvp+AYbYL6F5BBn+O4Gy1z/cKBDEYWPvH43Dx9ca16Bc8nXTxPW/uz
8Eg5vHk9a9HnbVBTwB6K3pT90g7yJsB83z+G4nK5nygvvm1libmSaKCOpAL5rzKoQWqkXFxbYskU
fQihPe5ferQIPNyxbQHl2qlPF7kgBVpO2qTz+afhxnBEBiSzhqYf887pUFyhaVpmQiZav0uEbrcz
ngbpl4Kyh1GvCRJlGeGqwfw+Yxc8LMNtY4NCtQuHSYcNZPv1CsbQhBByUBsVhkx70Jse5fL9LaGv
m08vvKNTpYr9J1ACnocXsOAj8cPU2hzzbwGGqqVDENeC3mZ0+EK14npKDHUkMmZ74/lAjXWkYmWx
Of/ejYwcyhoZThZxq1n1nY9s0kpNh2cuEg6GWQ/IWye30o7P9aNf1ka0omBmJMtnrEzn07bopxjS
sLOn9DDxx6KOqocTJYbuKnYJfpqxAZSve4Frj97KSDFn1RY/393k8C6mu8DfGPM6ObscKWMp4pK4
XnzVgiONsUP5CddHmKRJhGibVJGrwrbU8buXNIsgwczf4/DyXmdMlSEgaS2bcB4Mj+Y9BtuR284H
k9qBSIipTg9/PK1+JUKO6gDKSPphcPTsAxgnrrFVgXsVa6lOauA8iP/Y2+8U4OPehI29n0e7cHSb
StpQYlmlzMke3+DPD5XipRlykrrDRziTGbHZhB042Pu4qFyTzh/Be39mwJRhLUKL3yCyLl8u/tzt
NHasOEDUg1BLOANyBaX2Ao+nzdMO8jhI0vwZOi7YNY9VPOIIuRKjIL0RV+JXbunqIIeJVQg7gvgy
4F6aF78YkcJSrlk5Lx7zgjoC7cOE7WAyZp1hpYze1GY/bw6o3XF1/Krlog7ULOACT2JtOn+GrE7w
iBcE+kRwi6h3fvecL9Fw1tU4OLH5kTV/20ngiHruEwNoTwp/EIPfXA5WsecZrtTcKi1Vy7O6Jw2y
8XoQFqeum1pQqxLJJJtS5EH5hM22b1suGBA/XzCe8wJfJvw/6+z23VwnMUgesER3+wDgjeJiSHcy
pTiWO6pMQdm37Z/edHrxs+AvuGp4mfLKc648LYOHIK9Xxr3BQt5JOfZpN4IqGBMluQYL6gmgz8Lh
C2xfQLsphRKiHu5IG+KLRXRb0s2ffSdJ8rU1pPLj1SvYtfI2cMmIdY6TCkLlKrwvbgH0BOnuGQJQ
BxVRHyoCKX5D5EqGnEw4zmCheRWJr79YWgLUgT1R6HF7gd5bJso500FnWgpfK8xIx6J/31Mwy0MG
R8N72T+Clc91VNtB1mzbln7hiLjWdd7sh/6kC++GdjIq7uPSENgnQA8XavJQCYw1uWLjtAJ+C2ij
gHP8Ex/cs1s+LTnoa4neafqrT4lZO4e2zpjpK+coPf6phSdfyl/bblPgI6SrNgjN33euIKrR6j74
o8mbPSqPfGXSDJBTjlFMKDrkt40oKmuV8VUXJX13kmSYXfZ0zPUnO+AA3+ppF2kbx47/xFK9p/pi
llhqv/9c5vDdAQbXgVtJKNo8hCuqs5NqmnSSDjnrynZGLW+jr8Ms2gQ0fz9tMN+hlLtCJXh0JxYE
OjdvnhtIYQos8isUzTo/rDiv/XVXQBuCoZ4xFua8KmJlclOBUgQLSAWYdGwslzfixKQHw74GSJNH
SI2cuPXgFO4WxVP1D/DQHx7pB0eBAlwpn3bW4uu75Jw1L3pjmdrhEoxFp8dwu0en/g8fFBWjQeGc
69USAuOWOD/XXZ0B0ULgoQHPtaGW5syTRKzNS56KZEdV/fKRkElujj5Ql07uXeq5Os3kdM+GfYnU
JVXR8bZvkVGvtCgg+6oqwJR/uMqPoJicA7ZreiqfqgVoT6selo06yDvTs9nQjiukTwL6P6acKkZJ
KgFe+fwjUfbSLam49CNpptN9fcX4chKRb+mbtsXwE4orJEl1PvOXvokjN4R/h+v5uNPT3YOXxxwD
gjbiZhKToDfiyohrS9LvEQssiqJxlG78hedA4Eq8Q8ZUVwjsoQypJsg6g9A20iphwKAULVP1ww+b
KZey86CiPB+sRfv3f2q7GHWH/Y3jdItYzfSAdHxVMl7JCRkKmT19G4HDW3ywSPICeMirAjptV5m7
gG7EOfm0IyjEcSVCYdhlTZYbl4Rhy4KfyZlrWmjTExuQ2EIxo7rHLBfon7fUj0k/UPTIaI/KFf0s
zsugSGFBhi9oP0to0bu7zCaPYCON27pvYhYGchdK+W9vQ3ezBjrrZIqux4cLJqXIhdgtKYKXkCeu
bmL4uFn/3FOQ88pKAboevrCjz2YZ9nhIBdSPyA8OjybwvNMvTgaHXGV2jyxd+dr6TVNkBVJ3Iv70
PfRCAFJhI9OV24EZwelR9Pr8fgcbPhXwcw==
`protect end_protected
