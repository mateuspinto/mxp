XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|ӡWh(ICϕ\���6�,�>m��e�{�c����Z�y�"���N8�=���1`K�-آ�ʣ�\���N�kJ%���M' <5���[��!�������)В������A����)�Q��FCN�aѨ�_���0F�Jy(�L'wd�t�f�͐��Y@ӑi� Y� (�WM�r(oi�ϥ)[�����[�$�5{���Sqf���~9��6.���xr��M"Q�t}�K8�G=�9|����^<.����VA?�*����6m�/~�WFᓕ�րI�E�Uz)s�'i2O�LM�w�phb;!��tXB�L}��=�Q���?X^�{�	��(6���
������_8i��Ƈ��FYb$c�F��������V-%¼�w�:�gJ�u�0\P��J����HX![%�kf�2`�8�����=L�*t!1I���1<%�u��j)(���W�Ȑ|w�֎��AM��g��2��$��TPNG���d�S8AԄ�O\)�Ǖt���e��Iz��4��mu��l�$7Y�3����ɲ4=��ϭ$-bs��k��*��ڛo:^O[Y-Y'"���6��(�K����X%�E�.�7����\s|���o���v"I�*A:_;-�"�| ��L�V~Q��)�@v�/2��6ȕ؏V��-�8�����BoA-��2/�}f�_9��d2�l5�L��,���� K��'9�^Jv3f^⯨�8�K�v�{f��yR͍n3/�A���D�.9��M-�h�~��?�~bXlxVHYEB     400     1c0e��BMћk��#W�B\>����rĨ�����(Tj��A�NFh`��Dڄr���f]�e���[����'%%F`�]�y��?MQr�Yn9Z���~�D���tgo�S�P����z�+���r8Lp�]�F~5m��-bd�@�^c�[@gS0�"y"���Ш�d���	`~�H��}\��5�O��ە��z;����^����u(������c�F7�85���BUM*��q����I�fD5n��9<�	��t��0īL֣0I�ֱ��_k�5��Λj�S��5�3���G��hp���ԧe����K��Q�Ԝ��Je�`{b�QEp3`&�n{[@X[�X�y�l�:�R$���Т����|2ޟzr�=�q��������V���:�,�VƣBą��'@Q�/����}f1K�j<�o	����<���[`��H!����?XlxVHYEB     400     180(�0Rw��������M�Ǻ�,�ʐ�2pOQ�g4�J��?�1#(`�n��_����&乥ۏ;׳9xG�SW�Q��W�.���ǬIBś������Y�z���l�IL��/C��R������D��G=�&/�����oca�`�<a)>	�JZ���
ĉ�JZ�	)1-�|�klHĆ(����|�l0�W�&��J�G�s˺^'K<�MA�:�Z��Iÿf�H��MoG�N\7I/�3�D�R��S姯c�W{�s��r��^�qؖ]0*��2��GQ��Fx��U�Gu~4r��3���`] ���u�/u"�|x!uF�A<����f$]VX��)	�s*�PW���a^5%W�x��q�`!$�����Q�z XlxVHYEB     400     150t[Ow6e >ͫ�i�8���P�%�*[a��Q����_x��ʪe©=FZ�z�Z��>ԋ���Ї�p��!&�K\Z,�Q5W�[��8�D�w~��Rl�D�:�E��#l	�X�6���;S�~�xG���4��@1�_�=��,ɡ��J���Ǚ�J��l��X�ǜ+'m/Khw[G<�V��qU�r��D����~,�Z����h������ d�lB��?N���;�Y��;�xif/D�ɲ&���w�`P��k���.��c���P���^.�8{���=͹��"'x"����P|�<�����<uǖ�>s/|3��fm�\�IX��s�5nXlxVHYEB     400     1b0�J!S9��Y��Su7��j�G@Toip_���(��"j=[��`ޓiU���;�]�/�vOuV׀@��+v��bN�ێRM��nUL�W�����Ff�}�^4��p�y�ɨ9���f��h��`S�� S�T�(B;�M�}�J���������:����/��:X���w�;(�C�m�t��|����3EY�v+႘^���n6�e�J�W�굎��Y���g(�n�/vOP�19�R�����BNQ@��y�*�Tz��IG8z��u�#?�wx��C}��<���\����]W��M��x�y�<ߝ��=��zoN�覈�# k�; f"��qr���
���.[�GcZ��LŁW��p��F����C�����a�V�L~(����YRw��x8Yf��Ź�g�y�6�k�PY�p��WXlxVHYEB     400     100�^�.�`׽J�hz�$�i⥧.�HXw,~���:�G& �ǹ��=e�.>�a-&��OŤ�y+�Qf����W�m��F���G��D/mώŮ&�<�3���=��m�4��rx�N)�z���#�[�0�R� M�eB���­9O;��`gǻ�o�F�7^�`JF��V�n&�AS��ҫ��*X��U���������I�y�u�wL���ĺw�G������=ZV|O&p�qiQ��M�Vxs�'�;�XlxVHYEB     400     120�1�YQ����'�s)���TxL�a��y��3��n�ax;���o@]M���OE�� �d6=+��G��[JÜ��f����&��@ �u�M݈�}�R�Q#{�
�v'�8[ʑe�6Y�����W��G��2C}:�(��P��Y�C����(j�nG�ӏ�=���K"�� j�BMWB���R]�m���?���3G㢯��,K1Ŝ1�K��U�Iم�n���
ѱ���;B݌��/񺨊�m��״3-�� ���{lVm�[�0��o_�,ge�#�o��̷�`�4XlxVHYEB     400     160�R�}�F~��M��ỡ��̂{��V���d�p�ۚbB�MN���$�V��p�u�aK�t��'��)S�4b����� ��8}���h9�|i����z������5>��0�^�]e;TCWA�C�-���Rg+0%wp����@_��](c�&�-'�o{�حe�LȞ@Ə�Rp�t鮢5q��Ԧ~��O�o��X���@�0
��I���#3e/^��C��fi�)o��XaN����a,*`�th��zGl�C;��gI�Z��yЧ��D;�<�m�ĩ,���El�� �o��`����L��;WX��Q@��0�d����	o?�Sd�|Y kǭ�W�N,%XlxVHYEB     400     110*zjRugG���y,<�I�ǷUCH�MԆE�d2* y��o������'��m�f����>#$[�cn���}����i���0��?ɲ�3P�#���Rײ��|�`�p�xހt��ul�5p���R@�/�8aS�I�w6[���M�^k-�d۱/�
���򱏃WN��f��5�Uᑃ�� �,�/!33H�wf���d���`��E��̑�rbMy���"�̼����8s�>��i�>F�k��9�����n�+3{�n���\e�ӀW&h�|.�XlxVHYEB     400     100��+4��c��(	���a�J�F���a��x�ƥj��7M���{�L2[�o�z��*��l�����ߺY{����y���E,�:�u=Kk�l<�� ��s�����&�O�`��o�e[*M�7XLa�W]e�"���F�_��Թ�Q3i'�{�;��vmC؁��n�?�"mAt�E�x���%�g�/xg��f,I�� �K�~B'�:s�fk�\�n{e��	���/�;�a�9�
G�Y8̑�3��.<ׯXlxVHYEB     400      d0S�S��i_�.?�Z6��w#x�"I<�E�[X<��˧	�QJ|��;���{Ƽ ����/z�Z/d�S:�^G��+h�zN�	�G�/�� �?!��*�[>2��׭7?���K��ix���2�A>9�b�~�A�r�H��_{t�~������?b��F��p�8�$���h���`d�P�"[��e{Ƒ�3B��	𕲙C�"�aXlxVHYEB     400      d0|8z���.T8!�S��N���.�^z))�OXiZg@���)������֢I�j�>����f���� 9I�&�b�G���n��C��4��U�r�#.2i���΃"����'�����-n�r��/j��?#���?z�����sk%���!'Z���@sQ��e0���7-ՐN�|̝H�}dj.q�e��Ԟ�r�9��JHy�XlxVHYEB     400     130*�z���l�/�D�u�`Ûc�
��<yQmj�(�. F�������f #���y����?�8�v|����_.,��(�m�% �Fh�q	)цy�,��w���p�?6/vb�u̢�*�f����p�����
��2.��8I	�O�P�Q�&j�^�փ�_�zp�0��+WY�VC���5��"E�ƽ��Qi�F��c���x�[��Dw��x4I�`���>)*�e���s �'���l{�#{��X�|1�G�LQ��S�{�Vq9�3s�z|� X;�UX��ݻF�|GTɝ]Q�>A�ke��-�~XlxVHYEB     400     150�m$>$�D��a8C�D��#}��US� �C��X-�905���a
��/
A�T�hٰ��a�>�+D֦���.2��.8�ڱ����-�gWw�T]&�dI�>�ֹ���bL��6y�#���n��~|o@t���?L�oqw<��9�]����{����s<zb����uP���Fyh��XA��Z*����W���w��`	Xҋ?�rώM�6=��ݔ����C��Q9:����&��G�FH�����#���g��6�M�`/&�C��.���u�>�q�J���ؾdl8��,d��20 ��v!9��9V�"A��ޢ�F���'��h�}-{��~�XlxVHYEB     400     1701��������>��1zv��L8���1CP�nr�Q��)_�׏�t-ï-Iˌ�O�[���)Q�Y��r�lJ��A��ߕ����Ou�d��x��6�(�`M�h^�P�_jA�;�a�T�c���6�;2U�y���{8��xL��U�Ә���r����i8x��5P��H��G̭��1)�f PȘ�8"fu��I��j��%}���9j�5.D�Ⅼ�Ly�|YC�G��	Ch���s�&ikzR�1��}�$yvb���TZ�>@s���x�<��@�%�E��g��, #}�l1�U����!t�b���'��s�ֳ�E�4�yu������xi����K,2��(P�+�q>KXlxVHYEB     400     190�C����Z�P�4�K��~�\��
Vsl9�!_��@̖�><��o�P�-����oy�yV�6f6#�5Q���֯g�nK��63.rO���p�p�Е���Ta�sS�ޯ�D|��u�%D�]H&�������!3��a� �uoq��;��|p`3�PL���$'��E��#�T�����K~<�z2�\-{5�إ��|���'ͦ�T����+zD���M�NŶ���p�.r�qjv\�	��y�Sz��������G�^~��nA��qo=�O4Axr�k꩑/���?��DG����YoB�rĄ~wݗ�>��W���Iz|R�xi5/_�W���]'*"�q1qS�b�;N���8�m9��"m�*oN��t��,#��fk(��Q�XlxVHYEB     400     180�>����ǔK�^�
��~�o�����B�Z�x"�£8��S���뗻ˀ��4�-R����84�oaNl/A���<m(�����%���.�
�%��E�A���=�.^�]��*����|u�$@�AQի�]�K���ܻ`�������#寠���h�Pa��L���Cs�}L����kLYF{^}��8�˪.�;E\� ��I�Qc+Ln��B��3��5��������@�z��
!��X���#��ے1���Y�$74�{�}��ߪ&��m���R�H�h�ȵ��&�Qs!���:�?�Ƚ��%]Ck0�u>+�S��\T)k��� �t�3g��qW����?K@a��t�Y÷��b{SWr/XlxVHYEB     400     140]��ψ�"����lP�.��2���	��/�����SIW�@��O�T[0w��\5[-�;d�sr�%2�`C]қh�	�3>B�
��7i��Oܐ�f{w�4j��\��PI�߫��x{��ua���i�_��b2K�.ֲ�!9.�sЃ��ʌ~p�i5|�YXRs��"bW�}b�2��&�*rf#��}��w)���R��زK[W�ot�Iqj����^�h�<�i�H�u�<�=�hh��j r{���-��&��8�w��1��3_�@�1f�����N�B$��S�Y����֢d�� ����7'�q���yM����&XlxVHYEB     400     130����mӨ跡�ډ��r�g80���m52���ƺ"�a�v�hi���mNW	��z.�+���Թ�෶ҥ�_���Gxb�{�ۯp��к����&N�Q��y=�h�1�?r�{A�^ȄJ�~��m����恮��Cx:g-gќ�������5��l}���cw"5�|�>M�W�/�sr�9��+���\�葢�<�#ʽ�8v�'F�0��/��[[�W��{Rc�-ߘA�������X��F�(Vv��w����,���*�7r3*ªk�hvՊQ u����G�4G����N�r6fXlxVHYEB     400     170� [� ��x���W0��nZNP��D�|S�\>�����86[Y�o"[o�)D?�3���vZ�4��������SQ��)O���1��x�&ƓHU�����񨶘�$��d�*�6E[؀,Z��e���n� a�0�i��nH����<�*�P>�}s%���s��6��R���v<=*�"�Pb�t�)a�;t�:�1?�3��_�Vcll��y���v~%�;D_�O|�`+Yݔ?G}������:��e��sbB����s �������T�{�߿im���i^�.w{�f�]%}@���l���Č��Pj�{����kT���Zd�Jf{I�9k�Q�>]�|N�XlxVHYEB     400     120�K�Z���H��BKC� iw��K��Uӟ˩RL�*���&���~�eV|H�,a��DRLz��{�2}��:*��$�x�o/��6eˀd��$�3�#m�;���E@a�k�fkhA��I���Ug6*�Z�����UaC�����������C-���U���$�N��F4�VP�T���#ʊO�×� TH����i#8#�Lc��il��i�i!|pd�.�����7N`���H��$ <|�d���x9B��G����V�����e���<�g3!l��vӹ�s�|~��ٹ=2�.XlxVHYEB     400     130#���?�0�%� p�@���tq�^�I��H����i�G����w�5z��y<0ef9�	E�U��/b�\��]l�ۀ���E����� R��l�y�խ��BiP���b0ę4x��;щ�^�i��P@6�A|�vu4�[*�Nۭ�VgD|f,��Y��Lh��d���ٕ�)�]���x�,a����F�:#�Y���M��K�4��g��b��[<�$����8��k�Q�Ь3Q�+J���N$�6�����&j�?`'̼5�6����^�:���i��[�&2s2�-��$_|P'XlxVHYEB     400     140��ŧ��):O��ϼ��Z�κE!�}s�.���\�[M��3�9T��m��n/a{+���,����Ȧ��w�g�����'I�r1p� J ��s��J��!�5��%¹��8ƪ�qQ_��B�d��M�c-VMS����u̝�b��xa;���¬�=�r(�I֯�a%[�j�m���;sĴ��������L�;*��$#e<�o�۰���J�5h��rf��Uӂ�'���9q�E�|���T�BI* ObE���a��F�&a�b$�����slf�a�n�x.Nm�%d#%Qm̦NG�$�&������h�4/̚2���͒XlxVHYEB     400     1a0����Aޣ5ԋ�SF��j�d�s�+d���??��������jאS��k:�sƌ��JgR�|����{�g1k�"X�O����<�s��o-�<TU��pSܿ��N�����*}����BN\�98��Sm7�GJ<@�1����O��@�!x\��F�h8��^���� ��A�7U�=T��5ٵG�V^;r~���3��!�_��s6��*�ĝ	!���U+�V�����R�(���@}��>2��d|7z��w�|T�;���b1\�r7"nk5|IY��� e�����o� ���f�5p(EA�U��G�j;�4�X����3����ZgV}{Ǚ
:�ѱ�����5DV�_
�V�8Ykj����_L3�5��r��R��_h�i^�T���r��5?�����e)XlxVHYEB     400     180ձ���ڷ(�a(�Ә+�\g��a�Yӧtz��e�:v�SW'#hd��R�i����"(W}���7�VJ����l�a�n�t�q#Y�<�[�}o��n�L�79ơ��f	���m�*�l�,?l~����3�W!�'F엹�jj�X
�C��c�%����*�L�'t��!b�5��>Q̲��5\cx�bQL���*�h����ւ�W^��[�P�������l9L*��(Q� B3a'������d����m/\��(7qH���#�U. "��[{�4��G;�Ρ4�H�����ػ�:�45p��Uܜ�cU�NwJ������L�2|�mpoQ����[��(�����2��(�6U�����2�XlxVHYEB     400     170F��N�əB^?/�+��WI��P���P6��FE�=P[�?& -|V���\?��K�Y� �U#�Z��|��iܞ� x�~��������T� �)��[��"R7���3�xZ�A�$�S��q)����k�K>�~m;��٩Ȕ�<F-i�N���Yp`S�ѮG1�Ld�8��D�soQ�/,��Z���2�0p��;J-hK�Ԧ�QY����i��*��	����`��#���j�g���پ���w�1i*ˌ�����}"e���/%��j;A��Og{�BFE�s`yk\o.��yD3�|u�1+�L[�Z�^~ux��A\�)���^�~�|�'�y5;�O8S(��~֪�,�U��O����=���XlxVHYEB     400     1e0�S��z#�+}�te�4J�$����L�@y����ڧ��-���Lj>�¼��J���ɋ`	�G��#KV����\����\c;��x��4u���9d�1E�Y��j�i���ŷ�������_�y��~�<�M�]
��헭�,a�P4�u���tP� �c|�<,�-`��8$A�ͤ�ŵ9ݤJ�t���#�6^��6�: Ff���P�#�������f��z�8�V ���j��b��a�����E�{t)s��E�}WI肎�+����������R��,�؋��I��\��O
����B���v�?퉯g ��9��iWv@ZݏBO�߸��KR�(S����@��*!uD�c!�p�G<[� Y��*�`�/N	KI�^�l%VOp������s8���"ܮ ��l�x�v���w������|�3��KN@᥷E:y�5��g�'� ����c@���XlxVHYEB     400     1b0������T��c�9��Z�h�x�n�O�Gj�Ga�R�.�5A=��E��p�=�r��Rm�L`�N �5�k����t�/�:�n������ָP��ڔ��dn�9��b�w^Y"�[|������H`�
n�%)e0×�H�V+��d�V�M�u\M.�h�����K7vX��8�xp��'&���@��V�c<�/������K��H��9��T F�j~��;z-(D,R��baHX����d���Z(��)�Lr7Cs\'yXKt����9(K���<m#t'ع/ԕZ0���_mhxG�2��0%(�x�4F��A�M+�:�q*Î|Ibr��D�91���.���J}Rz��z����=�@P	�U����3k��y�_����y�τYQ�rN�2e ���0F��D��%՘��1N1�XlxVHYEB     400     160󵢄I��������I�XX��##e�z�gl\��	�2wV��N��I�?��Kiz�2�+1�?d�魒�|~�#
w�̟���������nF Z�<n%�N�:��{}�W��:�D�\�-��`�Ѣ���D3ҷ���K�{5��?�n�����{A1���)�h�0Lp7"L�,,����%p���)u �<[�3�#���*"@����p�!�0����v:u���
�W=�T\5pok��%ә���ي�ތ����`HR����i?Sz��u �ˊs���������� .���Y�ĸe�h���p�M�e�.�o�H�R��H�y�ꪞ?wy���t����`w��XlxVHYEB     400     150�@�K�_?29h���^�s@q��=]��ٳ��@ /��['�����AI!QUbF|�����$�� ��ӝ���̌��88i�=mP�t�<���+zT�!�"��2��������KW��
|&����d��Mۄk[���#���ڐ�Y�',�����TJ��4*������T��c��%rL�ɫi6�t�U���rY�Ҵ�����-�;n[��� X.C�(O�.#AT��?4�c+��L�?v��Qcy��c��`��M2I�W?�S�����Σ���d���h��4iD�O�!A��-,��/YU�[���.Z<�|�����g��ReXlxVHYEB     400     1a0(Pz��>�k�i��60c������Y�t�k�Z<�C�F�ꋁ�P"���Y]9�5�%qM�D�]ez�yj�(�C�~O����i�ն2:���1r����B=�C�����ZYz2�'�V��L��$@�諐�7�:5T�i�`�X������B�ޅ?��{��bG�Ϣ������>[!�a7�:M���?��z-h|4�dΕ�n+���s%��cGmT)u�Xi!���mS�Gߏ���Vi�o�����v�3���&>V��s���e~Z�N����O>u����O�������,�7_Ce��k��Q�	v3�	YwK���W��ʹ�8�q$/r�Sn<d���E�1+t��},076{b>���a~�8�m��_��ܭw�����B��?�u��1�:�OW��\���50��XlxVHYEB     400     150 �a���f_"@7�Mʣ4�S��Wq� �͕;Op���y]Vk��K�p@c'�"LIS�*:UK��F�Y�	�`�..��9F��7��_�[
?kg)6���F9в4�����[c�x�Y�� ��V�X��Y(lj�^�(w�/甎�c�:���l�I\�����~	� m20�߲�]#�::�΁A�I��)��-*V�W5̎&(
%bE�%Hu�+�ȑ������ ku����T�W�d��L(u�AI�qy�Ƕ�.�S�����C/E���.�#S�՚�h�|+��&�p���$�MS�9Sfo̴(r�����03BE���������-XlxVHYEB     400      e0��d"O��V+ �U�`��2٤�C�����Ň�n��_���ʯ$���_S���>�
>޷=R�K�fŸƫ���p����E�g�4^�1d#6%Als��j�F�����3�������O�19eևk�����83���I잘�g륜L���1:SKF@�}�Rg����&Ba�]�V0�R~7,pu)�h���`�����u*���XlxVHYEB     400      e0WTi�W�Z�W�J�Ξ@,�j�nn��-~��l�ͬ'��Ɨe!������7��:��f�3�t��"{4�kĲ��n�.�;�C�M�";�}�uf����Z�Vzs;N�5���%o̔�n���� ��|�\�H"��2�!M�SU�"&h�/���`�����KVR�t�Z���ļ�Q�X4�E A��}3 Z���SmL���y�Aۮhd��5%�ʊ��[}�H�XlxVHYEB     400      f0�y��߄���=oK���(½�����]x��۸L�X�⟼�D�u~�/X�����-��(�X[�%Q��3=�-�8Z���Ƿ�B1}��
���;S��h�P7���Ab�􃬓��O�5!��M���c'���L�����-�t��_`���7='3�	r�\�#��� ��r;H�%�b�-����<Fm��E�*����s��v,�����O��8����t�V��`��@^�o�ͱ�I�f�XlxVHYEB     400      f0 b͑��r:�89u����`��C���ªw}D1��<�Q>N�����ƭҮMulpB>������m�- �	%���v��I�,ڞ���WA�0q�Y�9z}�"+!U�Bad����X�q�W�D6~�4>�f7�0��bǭ�CD������V��L�[}���L�D�*���)���؎%�ڼ��z\ ~N)���u@*��-�Hf��vAP� T�	Wl�?�2˔NoUC���DXlxVHYEB     400     110~��ɩB�˵�S���J6p}]�GX�'ђ�;��W�3�ڪj��z�B+�z
��t���4�!)$*v7��WbI�>���Y��V�{Y�k�$+����8�Tk�5M�,�V�a_� �J:G��YyBY�UW�^L�c��5��Cb�x���l�u�l������W9"M�K�7������h$�Gj�o�u�`��{�-��Sb���|6������W�T��g&��5y1FR�a���(6����&z�I?�gx���;�@o̩p��%�XlxVHYEB     400     1b0����k`��Ŏ�$  �3c��F�8z�\�[ �q> �)wr}���x2"�������6�D����5��q������e���/0�W��H�Y�]u�q^��q� )`�}�:,��[	r�gFT��/�^ĘS���Ӥa<�0����p��U��H)d�֭(&�`�dE�F�Hμ�v��M�պO�:T�"q���_�{���Y��\ۿ�&XAy��.v4�������!,�A\��1��6Ez��O"C+�μ-~�	��������h�Q�z�$���B����Ҍ?�X�gg5���%��B���'�Yu�׎��e�T�T�B+��5n�H+�]m�k�ʷ8�6�/f�����k.�4��{�ݞ��&��e`Och�W��<�~+�nP�����ӈi�4��M]���-�;�^�/��(w���*�zXlxVHYEB     400     140��>�4�.�n!J?D��7����Y��S�Y�]�ŵ����+��-�#K̔��K�Yq�l��Һ�0��~<:���S��䔕�4��&�WO�>:Ռ+��y��i�^4��v��<���d;���I�
��_�U*?*.t�쾐���g��˪��K�qZQ�J��a;��v˵%b�D�*�J���d��:���'��\b�Fu�Z��	��V�\�s�]�߽:kY)�D|�q_��$�7�H�GH��M�G�*�f�a��Q��<v9�ƨ�Ļz�y�Z!�T	����P?�P��A�IJ�L�Z��.�W�XlxVHYEB     400     160�a�H��������F�kKtz�I/v�N]�C{V�̨e+��z�]p]����q�24���$.$������ �i?�~�U�DaT������4Jo2��8�rI�&�� �Pɬ���H�P�b����{�^�n6(��E�7�u���^z�%S<�]�"��K�r7����F��B�cX2X��;��t�X�Z�7w@h��e
���և�0��>���؅�/�>~C/�mR������}�U�0�����3�J��x��xr ����L���I��&�� �MK�"��H6*"b�#�����P�ɔ��Nk��J<����|K=� ��~L`p* *���6�:�WU�l���XlxVHYEB     400     140ѵjO���f�*���u���\j�;��&�D�.f�p���+�6��M�ƛ�Ge�����a�^P^�tq���2�ךb$��ZXP�2�@vх~t��4u��o�K^#���Ŋ�l6Q͉�JcV07m�I�*��l>d���y3�Q�&7I�U��A\�� O`�IajS�-����F�������,=nǵ�a�4%kے ��Ha�C��c�' �;�Y�C�M`�m��n!�W�x�[�΋����8媎$%S��Y��'�\I���N�X�/
�ܐ���DxmgE�Ry(@�[m�m%�n��;0�p�fO�M�)XlxVHYEB     400     180Ӑ���!�z�������q�C�8�M̉2ff�~�1t �E�o����t?� J�s$l����Hd� *Q��5q��`�SݤME��&c��i���,:��@��i�K�<m�M�U�pIه��L��4CG�X�QL��R�O�SW�p��^PD?rm���%'�1Y#RiBr��"���Y`���zk���P��d	g�R�8E���E�H$}�=��G�:�U,P�O����{�����{صؼwӡ}w=��r��'�G�j�FHp�������]H�-���r�y�h�d�Rp.Q,V��� �.���b�Sx�2O�/E]`]����z�HPqg���=�g>k3$���bY�3-ƨ8�ulKH=�6�KXlxVHYEB     400     190N�%?F_�7�
��1^v�E�pu�o$ÈSJlA��ϧw\�W'i0���t޹`[:��孍8��f��?2����k興ǀ�� �s���׈lM��[Vq���ug���ܤ�jZ�;fE�rI�%f�h_�hy)�;���	ҕ[!*�P��HZT���@��>��'�5l�!�������N�ީ�(hn>=r,�{�����)3��W�[&���q����ff�52J�<����l����?w�2�Ǩo>e�����Y3y�FM�K����Q�uE�<YL>�*T'�!7��`����\�s�z�h֪4Y���D�Q9�F��!?�.W8x��P� ��k��%W@m��C��W�g�8���+�ۣ��Ò���d(z$� A�\�^鼶�`��XlxVHYEB     400     1507h����hՍb�:I�1�ƦH�-�{���6����?��t3j����l	�e�إQs�Ds�3��,�m_��vܲ	�Cw��8'�2�ߘ� U�� (&t��Ӷz���^uױ��f{7qd�Z��w��_�)����
C*zKMM��0܇Zi�o�ڑ=��x�r{L'��5h?D�i�z����j�«/�H6k���_�k��2�FI���7�~���f`���^�����f��E}dx�z�ph#v����}^��15X/cW?s>�tH�T��w5R}��܌^1����(?��\���F��ջz D˻��XlxVHYEB     400     1a0�EY�i�T�$a���z�� _�|����hC�zo��Ʋ��w�8��&��G�Z&�Q�-���J=[�{o���蘘��o�^<gt��G�A6����t�7�ĕ�����~e�r��G����P�.�9�U,�9���}�	��L�S�D�29)�~�Զ��6��m�>k��"(��_1�zClv�)>*��L�'$�m�v�_��KP(�����`�<,?l�_���-�r�}K�,��))(v�X�ǟ��6Iϕ�b�+ݕ�|��KOR��X#�.|hZō �����	d��`��������q5�H�E�?'�&�3B��(G��k���]@�%�.��z��mK[Ѫs��e�7�:Q�S#��@�y�x��	��:����q�,��ZaxC+,g����C{nGoD�HXlxVHYEB     400      f0�`S�.}��ڦ����
*�`#�T�
�@�R�K���y)�$�18w�"{�&?�E0?~ޡ��ʣt�e��[��6@y-F��|�Azhڤ8_x������
�&�p4��~�)�Pl�����@F����i�3�e.�k��n!�����)������F�3�9oPP�F$���������֟�j�+�����h�ߵ�8fFd�b
g�Qߌ����?H���BV���0e̖L�XlxVHYEB     400     100bQ�1�l�r��J`�CV��	�8��ȃpbUz�r���AF
���@=�2�,S��Ϛ���^c0�z<{M��q�}0x;�l�a��w��~��
���GA�*H��"D�tOu��:ʭٺ��h�Z�/�����	:�R7��bR���ވ�σ�Hn�*g�M��[\y�;���_?@�D���c�;�b�0�=7"��M�6u��o����g�_x��$�q��Y@J2��g�H2+�3�8j�+��t=�_���XlxVHYEB     400      f0���t��d��F����@��:�F�c1P`��iHD��=%����j2���$��$R&�lO%��~Tlz��i$�L�& /�����DWk��!u$D}F��k=	�@|x!�;Ru����X�1�C�8���b38�)�\�1ݹ��7�v |O��J![^}rh�jd��;�PD��WާZ���b2����'�=p�R�A�i{z���ꬬB��e��D ��[��Ų�4F!.�oXlxVHYEB     400     12002С�F�Nۺ��sA6@���1_n?V#h]6W-\0Xq���r�S��
�%	81��C�^��`�LQ��յ�ab��<7M^L��1l����N�G�ySk�+?f��q/�j
Zȡ�|0Ʊ7>���w�<6���j\�(C���f`}�m����]Q�!F���[��yc�@�m�`��u�7��.C���(���*z���Լ�0��\6+�[.��9#W�7��-K��cz�fm�m��S��	����m]ͱ^��˸���x��S���t@ ����XlxVHYEB     400      c0>��ƽĨ�<J�TT���+T��a˿��ݬ&<�썴��j
ӑ�(�㯺�-�����zN^-�l��^hXyI��_}S��ȼ}Xg7+e�:@�-��r�F�X�}Z���*�)��=`q<�d\&��g�Dq�
���4y�km�AS�!i���W�]Ɓ������fJ�c���E��HϾ�5������<�4�5XlxVHYEB     400     150Adr�����|��a�f#~�_���7�1�k�@�C,�<�$��k��j��SI�y����k��q��h?N~B�S�1���j�����l�;��rfk;�F���r�\�M�����z�ѡ���N������h�N�λ ����M�!>��3�U"�GE��ׁ�q�����IT�,��LWT�\����&��8>=A��0܆�F��¢r�A��p\υU�����p��<I�񬔃A%u��&eÁ��H۝�ʩ��Ҽ��&՞�z��~��rx��F�H^��v�9���Jg���p���*�jMzL�\b����`��#ity�_}|�XlxVHYEB     400     130Æd6��m�e'�c�D������y`@��
(��qj=��'�	��0QڼZe��o�0�ʧT�<	^���&�(]U5��lr�����	�á�*Eܷj�HVפ��8�cO��w�W�<'�T4\��N��퇩��W�*�q[�L�q2���7�p�X��g� ��2���䑃Q) �����f%�������XD��o�A?��9�an|6�(���vy7���x��]�~ϴù��q�s���{�:#�Z/����('�6)�2b� KF3Xok|FiR۰G�,���ݯi���U���XlxVHYEB     353     160���a�ܹm��-mB$D�Y�'_/�~�trk�
��Vq�y 1$��_������\�����Ҕ|�����כc\�Z�wE�kT�+dĚ��_!+�h�ٝ�S^r� �4
�ubn�A����)=��>s���5T�K��YzE
4��qXj>W���5�'J g5���E�-e��$.�e��L���9����9�:q�)0�T�mМ��nX7��g/����nF����nN��]lB���9K@z/���\���|Dr>����!�%��lt���͑밸ͤƵ����b� �\#��������X�6��HG|v���g{�8] �s���AY����V>F�