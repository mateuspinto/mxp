`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
A/S2IBTXOtlIGTMOJW+/QR4c3y0saDie8YXWdvp+oLNhyltbhbRfT8qvoAYO7nmi08qQ/StbhDZi
imsnltNsyMwHgbQaRnALRqKEjkNJxAlExviGhnmNNWDfYJzeqp26nURBbhOcabHpKXjkRPTlEs2l
k52KYOTHvfm6EkEp8lHGH57YyYipptP2AXLnVvjaP8BWzB3qpFhXA3DOyg4HcZdBTEr89eYl8hHy
qf3t3nUHURO1HCHsWsd6RXCrO7HmAyY/3mHNROCLFN9+tLCVCbfoHlYrr4SANKm0ydirz4iCp+G9
1q08BfDSKJFURYvKguwENDlSEd3HDif45BazLA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="rsVbdfaqXVOJjzxClQNEu/J6QDfuqEJtw+mxpECFxhs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6912)
`protect data_block
9RJ0Wp9pp6u1VrXSVQUO1zuCjRi2tMvLNfd5FdqHySnsb+QSaIVnfLfezYGKSCYOOzRDn9sGS2g/
Ca7wXpR15gLXssjVhr/icxLFOYIV8bOKArog7B4E2BWf3m6gDqwiKjXxXMOG8EMZJckJ48PApF8Q
tJiahVZOi4ddJFbmn04Gxl2mPpNg0vFLjxk3Nv7/gXq5NuKw+Eh/5HLTbYQy1/y1+1raGfhmkzOB
37YjI2+KwT1QFrUME3nvN1uoD3aZZZhy7mYhWeU8nU1HUUlnasuasb8G2xAQXXC/OdDRuuQqzlr0
kw6EQvSxKbwRvxRsQ4swjTo27qRO6SxajVWtExoofonWWx90we+Axg+ksf/fGQeUDtgL6nqWFTLx
rQKUOGHn1jp9TNQ+/OzfmMGBeTCWIuEpKWhm/yNQanOKNcx71tF+PR7Dd5FX72GAqF/W+CXvxv9B
2zjcBqPJ8NwUON5PsIUsfkbTR93yOCaG4AJxOCeDohCnoLG0NQA5avYE2anVmZ83MYdUHChKZIla
+mJBQn1EQ/aq1Te7l9WxSg0KrH4Uv7IOUIjFVnXCyCClzkLhmDE4h1E+y9WeeWTjlzojbBMuOamr
mahGvUbzMjX66WoGsjEtQxVWbut6x4aQ32LqC5vJd0N9Z9WAZ70O97fyME+v59GiFzsz2PgTOokU
ebLLuaR9Em5NFYS2XQQ1gBr54tlpXjgE2eNN7kOKccKVdkCaos4CB/dnpkVlAfN+ERayJw4y1qzp
2AfiAIBF6hUSUNz/dSGIWrOX48qJc+vEuJqXZshpayoQSPT+KLk8WSh6tnZH9eNAalc7CpnQ7tN3
JmJG10izlHTsFoA/xlMvku4R23Jalth/PRZon/itgoYSEmA8ZlLUOeMWWUbXYzYKKPt6LsY3PMia
q7KU61QkeUZKYVLcF5HpHcsHVCc+0go8nep6farA1GYEs+Ew6RtPsq/0aNfDiPSVU/MeqCPHW44E
eLzEBJPiH4VKgAwhqexcWkrn9iixbW/aoSMgUCD8ImxRxKzS7JkzcjSE9//wCr1+GiGKiEQrH9r6
D77tV1uC87kWiv6lD3LGraesXpPIpbsMSAY92AtOAajXyhlC0KgGCyiU/EijCsfT18wKyBtrBLLa
2csGqUEh80TUaUe054Lq+myxM6H2/YYB/3XLRN1DhcqresBa4kAeielNqpSWX1DgMaNjGKcS2Gjn
2wMOo0UBTOVAbckCknRklXTnfXR1QNAI96gMG/jkPaFGh0N9DM7DlAFi12hCjBOvgi5s5yxhteVc
Bz7Fp0nwyzGUlFLdFEPsE7KbLCnUtUcW/le8WD6QqqG0ptiTtzRWepbbsMLxpua+5RMFPdxUo9Cx
LzcMS5gSosPbgqnSOArSZsDi0W94503yLqkaTR3utLAa9B1Bxr9Ba5ms3Ai459HL2coQMql15D1O
SNBdx+Gbc1koA9ELEUFd25Fy/dC32NxI3PJBnCfwiZEESXG3fVry9QjnJkfOvuPFHuyLZ5MvfX5W
ccUE8tH+r5ZgN3HQhCpmYZEf9KYB1EOu3ACEpDVlgiAy7yMHAypghi2tXGif8O1yZ3J33Vnknvwr
Rl2NS/1b4oPR6HleX/nr3mxMlYkuMGiXNbwRBTGvGaz5zCH7KKTd0emCCW7M8c8++9s/4K2jvOxg
76Sgx1Z4Esp6HnLzwgOkVgE72Xkd6dAIeCUI/dBXejoyxB1iZ4dqonrgVhabvM7yiRTKo+z/ZWqs
O9HKuaP966aDDyRJ9Uq9jXgw0L0QfjaEy4XxGNthi23J7PW/7FdAboG44Jotxuya5959WqLZXQDn
wLo2idEJxrZY7MeMHqJ4XoPGPpI2I/uZuDPjbnHzwPQY6bA1wVD2MeSHh2eslXvb+hYKlQAkBJ2C
CpYoswm6M+ZwIdSubEvsWMRDW5D4VMAo27WxsYS++L99j5FmRdHFuagQg7xDl4ylYCDjpfPatrdV
AhwTVWg8WxfcVR2du6W/v0Gelcw9UkVbMrgf2n9oqMMOM1RgeNVQKqpr6TTgArsev3/SiXzjw7JO
Ckwc9A/y9hjuoq6gK9uFDa5J/y19C2Y0miX2x5HKONEkNLDJr+I4xW0R5kxKy5esrpzMVaw7jJOK
vGMI1+5lCvyNEBBpB61LQ5FpXmlalrZJwqY2b0WbkiCA1UlRk2VtAXI/TZJSHPtdSnSk0Ov6Wqag
f8XOjBMDO549LKr2SVSYZ52O5N3CuTBTz+2Og53fWlWPzQUIKtbHKt9O+DGoCyZq+WgEzARNFqAH
7ion2/to0EOW6Ethnwykivb/hDJxIaao2iNB9Ek94f0g0J2X/rg/hJuZu/RTEVpMmV3nYZFN4M4K
ZyNl2+rpA8RVkeWkDlJiTmI+YHVX5Mb7yTSRs3/hCfeyYcmpLgIIoK+q7DYw3PKvVPuU4RDbQk0d
9DDjT5GlKMGwfnpKnw17GYn5k84Hsj2lXG8Ny7dkVMmJDTteIFCo0tWRN8DW8JpJzn0pMcJ3exjp
11wdmdZn581ijvEsOlsfu8q/fdlgf/8tg8qAjuWOgoDwZ1wo0C8NajMrW383PVL1uhiwrm8TNF5y
CtJSKQv/jpLgQVA74BrmoM+7oXXnB7twt2iNTecIBJR/N5sNZ1go7mJu7nlPNLNhvPB9ZYR7TaEQ
/SKtqm0yiVureAvCmpZv3m/V8ZRMfFyP8+npVJ85YLsBhl1MpSuS/wQBRoi0jeJa+gevx8BoJQzY
OTk0eEwvUp/pm4zTEao+xeR+9ENEkJS1atWRoxWq2cA5NtwCiU7HOAuw3ISXZZyUeXVSXZyPzugq
OJSYPomJoqqSLU0EWnGbD9yCSo6uHiePG/UsxSFHPK2PejepOz1jHnkGauUSLbXcN9vgIpf2joJq
V/bsVsHYrUPTWRn9UoBnAA+jHbKh6G3w/qpQcs64Em9djAlPYpRuXGsLXBqvBCybfmknruUtqcVi
v2Dfrkf5mmdkcwub0kYpUPluzUIEpaH9het/vUQpEv4sUIuKg5Od84yO2WojRoOPdqckFNedJPMZ
wpKV2iDzkbkGzB4ONvkNkjOHYd0MZxhbqQTQH4S8HOMyVDEi4nsmfylb/ujSBLSCye8RiAXlCxsw
t7WqTssInjyFugXYUb8yr2m4NUCPAwYC3xt2oIwh583O4uisQ+aD06M/IengEeYJ6Duc+ZiN6EnE
mDH0fIzH2OK65saKG5JkGelTDCLCqG+CUPy1NUDZFN2rYN5w1j0ecNejnbYJr/2PrrAJL1o0Bmgl
+Sgqgh02l9c6Xvm+yKhq2YLuzi6MZsm5DGCk399DP2s079c4OTCqGl5Kff6ttN+eklN1st2pcbQc
iyoqfsrJrJTLtw5OjY80/d+6uzJat9TnGvdgUUKuxFWepeMnQzTiIL440R+VJ2a1Sw8yJqt0fBo9
M+cg0H98lKw+Z39yDcwVeGSSwjYhhc2sVkVX/ssSsx8VyNFFTQ/D0OGFeCySgXVrmFpDHm+5uPKe
lZEkYORAiR1gmk3Dc4izsWjayJxMzjeNQrwqFUADlHhOoI8cRrxCbC3SrnfoHBa5JU+LBH4D+56B
8hw8KON30TgBlrObnHtAKUWfFibx0PIgPfiWZU8ZFBXuqoyNG49VOIpn340mApr1kXt9qcb1l3ax
Blhq0CsKg6Izf7K5Wg2bU9JASaI2MiF5Gyb7lsMXNNVKf387qp69Gaua/eQ2HWMH+/SRKzcnJXVW
A/0VA1wsUgB2VXonMB/H7bMC0HSb8h7IvxbomXa7y8OcJftrxBApMwrL0ZRi3rXvi1oJe7ZWNsYJ
G4iaUSVW6HWKNGG95DawmGVVJ/9xPF1+PbVLayGPmY2vOLi3l2sz+ytR+DiTct25hBe+NsMEzN+b
W8WTQ0GFi9bvAnVgtBtmp9YmsLv3rYt3l8rC+gTyaIDo0nNrcobmtVNwanGing1/EbpKOOq4wDke
cMcOczPc8X3RjrkmmQutIr+FSI61fshe1Q9w9UMq+kAGO2Rqy1jcuuLRk1RQoZzuaBQK8FZu2KMh
VUgO+txhNndebZpLVtMjNw6YcKo7M2SUt146bVF0lsZFYjn/rdyYdW2tP5GWCbLc8vdUtgUqSNzv
q0DHaJQzz1aiwEiBtsqPlX/aj6zeTsHm6aIEIA4J9UGhF7qAAPSkuRX+W8aDCeavm3/8ZsaUNFDM
cJ8dK+NQ6f7kMadoyAYxbWJsaNgiDax/yl2c9kt08HxLFl62E7xC6mPicDQRlrVl2h87Qvqwslr0
hOvM7nmAEt81hUFRGgarT0rprBi/Izh7aFtoS/2bC6TGctgnimU1fE0u5ZUqb9SeX5YSudAqAR0L
H/xgDI/QBE1ZCg9lzG77fyZu4vpkZJRU79gWupTgeClIe98VH4LCzue19f2/nadZPZPWd9mGEDSG
tYtG0F8aRVrVBrKHcszaz1Gbu5x1bXVselq7zR6wWCHf8mpprGlKxe9eP+VV1mTVL2SZXXwKgzRl
x6Mz7YJ8YTeWeJbPOUYi0SM/pKJsddRy4354iM8hwly62CitO+f/BBA/H5CH9CNr1inPJzF3NldF
RcLnvKLnGts1VyplniEZ64oT3PA9gnSam/vFkE+8F1vMDuYw4zY7jtbXH/mmmoGtMKrEq7E7sb0K
5lMy67yn4kR0pUtNKw2OAEtTp5RtXpb+nSOD0piWbGu/ClUQNrZTJF/urMvupO+TYwmWanf5Jyk7
6YxxA5HJ9ks6c21F/j71Ph3TnBFviV7x11DNSrZVxNK+86P63DVLAHL11TlrpF8iec1LveVkUKS7
7mvYi05lLyEHnU4H0fjRBQpglrlP528g+Fjvh4RHMSvCw61CK5eA76bLL+Th1llSzfH+Naldmup/
QkNLaXrkWhDToqHQLhWUT/9NBfWEK57dX+tSD8jo8ZK5cYRx6UEp2obOCJKBe1SKXMe2K5LR1CLs
r0PTXT8H97IZyEndgynfWMhHh7ZBOJHFnEchk8AinPZdQopAa4RQk7w3HZeg/pdtn1bLsp4sigIx
Q/QSSuCDHVyXghPlVRU3dy1U1En2ODTCM13sU9UAmPRcd7+BtJAonLHKy0xFzVJ0AcMx/J0ciQ/i
mPQFMTEXYi9Tr03jVmS57/iTBWLL/Xy56mBwl1AsHyXMr1qsACpyOZXNFDRHugb3Wd+vFjcj1Uvg
V1RxRQaXA0avU94WFiOKASW9Y4nMZ3gL9r1i07An2CSQ7NMNF1ifviIxR9Y7gAUBbKteEyR6H0ra
8SOqscggcqh9ho6HrtYjtjdKpFXn8r8uLqC3bY6IvBF3tKlJ2iBhBy+Dpna+MD+NHXjX9SQ2efEg
c3yLJgChMwwgpJETX38iOWk3orPoBHnV3iLqNyCWPP03pCzAG+CoxuSnMntJvjcR7cCabSv+P+vn
X9toy0P+RDXJl4bM+moy5LoI2EilmpFAIyS9gBhojtHb61fwK2F4lkZ2NevjKYZgAt04eHKbz8Xq
YAuM5JqcLdet8MMnNuvZyGVoUwwSZd7tATohXp6CUtXPKFMWfEQmhxZTun1ihiYzjtlgHREUnaeG
Jp/nqlgV8AWftW21aSZCv4qcJCQGZdGKSLTAClhB1zd+zWvaQkavxCq3MHQw34yYY5we6W+ERAWM
Ze15JEum5Yc8uusozkfw97p3EqEZHhJK3qzOaKD5hkcwkjBwFPIog2EAG1NkGfVG7+gW3QwgVKiB
xrU8ipaD+a/09cNWwDPSzDcoyLNP7jg+Zv7sfXbWMx/AgWT7p+7j2X9FJEWE5WTclBmyCw4bD+oI
5j48ouf//4HWwbVt5qZYpdq8S1VDoYTEPotFbeO/t6iVzHSwyBOZS1n3pl2tn9dJAbUj9KBrGfGV
RxpdGl0+v5Uo0IxTU64JvFoSmgtkpyizfRyJe6f3bUzXZO5P05bam2xClcMLKTo0L0H3cfmg4PZW
ziqKy4snXGK4ywyLInd+WZCmQ1Gw4DCQEIcNxg2+t64VjO2Hxyqvwxj40lfFCHE7YqlWtlUSFmz1
fmFXUBF6dHls+EdhkLIigU1OBcUeyX2Ik+V08dExxicHSajrJmaVosrOgaQmsalUagufiCyx2ke2
7o236iENuLkcIhLNdNM+vtZYHwEhVqnN/kVyOkkSEklMqQJsndwT97pt8VG2rrUj/5Qa+eObW4Oy
Uj9BcFoaOFXsN+47Xi0UCoBR0J/BSqg1oLSTHuLnhNdThAeEoks2HOTRXiNxJ5IX1eiVhfnOYh3z
Vcc6JMwxwDWIcMIFnFnbzUXW7KCeUPrT6qbMcdH5iD8z+j+T1SNlTm0Bz1LvnfJKE7l+3hVXSCTI
mXSttOUAwHxnxLI9JvcewAQdfyLYyn372kbRT/bXeb0PNskBo0u30XCPj/h5N0JKCfP+V3lLiFOj
pqHcegAM+K8yA63DFPRnO67JlQLrpomkOFdfFJlDEDODzkQOPU8abOlFAFqmG7VI/lo8t/4t1iN4
rPmXN5yyvZ3CV4Ib4pH1E6dVCNnJkELd7qPufYCxZEunfCWp1qX5mqxQOsmhOYvVAglCrbNf8Xq8
5FXFbB3hor5RC/ETVqSozEJSGIjwmZpd9Is8StHX07N0BCyXh+v1lE0uhZll093qt4/HEZQwsWe+
ktE0zF0ruhZqRWl/VEsjqcieUJ+BoaLCN2BPCbFnwcVDXCko3coAjFqv0aBLSAR6LAqjO1jpFMpe
V75kPC5muEw5OU2u3lwPrc6d6MdFtzEQZ8fXNChyRphIFYlw/GgTBKoB1sFesUO8Qa++Qt8X/lzb
1zD1cAto0nS3QEjXqZXzyYMjm3YqWfilFIBnfzHlIaeLiiK7WLoMwp2BYkQmQI7km9XhNhw2eSBt
LFSmQV7VWHiKU5aUa40Q7iSqSQutBMZ2zvCGHgL3iTBCircZrk9zeovUjxnXP1i3+sNNOmxF/mhy
jHYpMyrIOBX2P3S9wEN+ZXvAo9zuOVs0btbxTJK0+QBU0GYMdWSAUaVnA6jjkV1tra8JqnkmGxF3
G+GdpX7Gc16jQ08CMNsgYCRqV+97fth5lPrpVt0dVDvUXjsw/siF+uk91a7QKWdLDtJ1ITxxxNa4
stOSe7Lt5RKwk3Bki2aNgO+e2HDh33bW82clGngLGXHqSibh73Kf2/in2fkK3MSREa7ozpiE0eo9
0wgXD8K1CxwCvw8RG2+hTYTV53DBPPG9RVlKMpH82IZ2wovPp9EgKSJz32EV5/cN6Xf69l8TECpt
ueLG+M3slT0PnEpZWMdMmIzpR0uqiTnM/c9Fi5Z2sQZYGKvJNyz5glXdGQ9qnty/Uq69YYtmRqo+
b+CkrGldQD1XX365u1hbHDn2Utbk9kjsjQ4aYhA7GDcPthBxBKtUh54IbD+NFEsTYj3mKliqAzAQ
6IgKAd8jDgPJLCClrdwLR7JIqypT4l5S0L4oWEcejHFRZ3D3CREKD3u+aVlhkMwblOXbYMAfDZu+
sM8nU62qKTXD9wqPgmCZ+1rhJK2wOWemvGvlwnp5zhwgumGQvzow8MBFPLBNZs5nD3faTCZZbIm3
N+efswI47WRNUJGKJYDAEKvqg+f2XiGkGSqGOa6mgSgBErWQD+R0R8PqCVkRKzho1PoI86kpbXjd
va7WBibjPxr27UPlLhEJJujQW15a606PFcC2KiSnBN8esaZXNV5G3OFpmdqTPa2sQihg6ty4BtjE
fQxUyZQB/1FCZcfEsQXuRDG5gkgFIl+mJ6YSyfdSMJBPybzDKc0DraLS0/nl6xVbYiU7VYJJypMr
c7FJmmou2V7/X8mEJ9oaShOA/t9AGw2GTO5gHuTDNz4m4B/AsUZ8mPNiC10g+uoQGDNujsWUDtyC
yTom1E29tM1bLyoHRE930WK1iWbK4lV2iG6/QdRvKnZ5idGTuK9bxh1UKfpqIl4oU5qr38lt3J/S
Nw1VD9uuXlyfrxJa/uk8S0R/dYL71BsSJICklQWOLSPxmgrnVY3x59DxFoFgXxIrsvLj6K58Ug8u
9oR7d9sOrdP+Lw98eOxwhlRjMkGpp7g/GireT2id7vASUoMyetFIx3ngWxHqHwEP1/pLW80nW7Om
JH/9z73Kc0iUgD8l1gYaO5TlLk1LSolZCa/2bXMt01wUnXtv6Q2ae4HVj3ykhJvywKOf8350Q59R
7mTi53SDC0/p1fkc68kyumpsKFG0z4RPWgMMRf/9osRsVjZLgyEHXRW/OSEe6wxpaRzlxu+UOYg5
3zHjqwOZ6euiblgDnsB1MX2b3ZKmhnsIodjGMuym4DGKuyYSeX8oI5c+GWkSsttUdpCjLcAUHqa0
pEWQcJqReSG68yHsQNMtUqvvh0pnTmUkdCHh1XLSTsUYMMptSZ6dXz60TNZKa4drxNIiJjZ9zgbf
RJrSoMIqh+9biUgf6zzJx/qw73J480VkRrUfnvVTh+ilsZrK1OX27DHL5mYsmBp4QxCWiFWJ4s0F
982RydShp5TfwjTQAvLr1ebL5dd2tJU/W6tCIAaDmrv2he7atFM5zj/kUfdl5RcaUObYbKg2HtB+
cyFCn+7NO7fIDAYF6XmC7AmCCG3NfHNR8jnpn3YZFsB07Cff4sizauyFsSi+5U/8UfP2rSI3L8YG
3sa/rjkDtov8by0wlnAXzWjphcqi25kqhEcPiKWIBcvwEWzTymRuwiMhGuzZxCeB4px/K60/JUMD
IeEhkpVFG3DBOx/qWEImtgSi92Ku3batFUk9dcjtUMb2A+lvapOKPcybz+j/mLlpj3bRmZV1DvLa
/PWfGbIzB9WgKklA52NsxqRE7wGVxTEVqi8r+h8g7x/TGEVaGhXJauIA5W+XLOHEmASirOolZxyY
px6AbZVtivZ7Ar5m6YfuXPOOb9rgtueUUou3ok/vKOxcNfx7Xjb1WvNYWDgDVXN1xpbQR2tkiKve
qZg9XfXCxIG4y07xj/mVtDAxZ9sIcFXyHxVDDk79BDYRAvcxOOyweS11GbMw8/Q4Cqf63RQljxMc
3CjkMRBtY3qFwfrMqnElNJ38YyrjH32nVnbTpTeHk/SCVabEMJwnvZLt98M2GZp6SfCBFBLctuzP
tEHVc2QGWYnkLU1sd9+9TLpKFfqkXrLRZ074N83OfqJBJ3BY1dgPP2ljwfIyZla67x4e6hXFCRA2
LsVI0KDaYKveE6JIhqNnd68fPqFLg8ZBCh8sZt5dDMIXyMvT5T8lOX02cyUE6ORFeDinHHAQzbRB
J06ivk+vKvaDv6ZFkpc0
`protect end_protected
