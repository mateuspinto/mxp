��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ЦT��q�e����6m/��p1��(����F��'��1b���gJE�E[�i��=Ue�eR}.l�(&�����
�fYk���X<�!�=�F�o�1b���nZ���K�ɰ�9�O�Hcu����lb3�[N���{�����]�2[�/���{�h��A�x'�"�?�ֺX�7iv=�0F+÷Lq�+N�6�.��0Qr~�w�����V'�^�2@��67q���`�|�R� C^,|Z�rv��|F�Ԧ��S�^ȵgYh�������%��dV㧷?�)�����uxV��" ��5�\�o�u���`6C��ޠ���"g�y�B/pK�����7������b�mߙ	52c�k��x^���H(G,�-�f��.D?�
Λ����+-��-̉��ވ�[�&�����X_*���=�ףT�<��H���c+`F��no�H�Y�0�D�Ύܛ�i���&:��ֻ�ѸZߋy;6��
܂�=R�]?z(��-���:��>7>&��ȸ=�k"��r������I_����R8�֮����E���u�N$RJt�4S}_8��n��N��Ѱ�s����c$k�F��Hk�FTZVO�`� L}�� cgO��DhU�FϞh�ŧD<�h?�Tþ�/����;m�
?����ֲ���䊨K��]��Ga-�ܪTn*����ǋZ�Ƒ�I�w��ܤ�� ���D]p|[��<W��.�&�Y�/���on�q�����0����Y��Xyv��/3Yt�;�IQy�:�|�@@'l�5a�1 ���3h�2yO5n,��N]P=ś���V��<`��^TG4wX��NUi������.g#c�HI���e
�i�B}�I ������S��&��d=�e�Ѻ�EQW%��|�%���ǡ���i�19�E���K��&���r{�ݏ�M��5UKQ��z�Y[��s!� DW�!�2��8�x�oDv�?d�&�Un=���*�Z5ږ},���ᵍ,�ܼ֓�[̕����a^onLd ��&0�o^�e�{L��9���.�@a��z�9��h�͙�ѐL�D9;HX2=��+��Y�/OH�����b�6���c���</(�Hv6�~W�c�h߼�^xX#��5YU��Nմ��y�P3+Q�����"L\J��%� ƪ���5�)���i��p�	��R�'^Q��Oʩ-op�!�J�v��gD�C������&�N �J,_��s�	S�R���{qq�?g.���\p]�遟�������JX�t`����^�`�91e;��A^޴d�į���×E	`%�/o�܁�9e�>�G͛N��5�e�(b+�KV24Ғ](����C��G)�����ߟ$�6���*Q��l�#>g�b��ζIx#��(�J���
ͣhu�u�.�d!8�w\�_/_�7w�D��m�������9�D������ׁBpi7�	U����>zT����c�p,H(����76�aZ�b��m��?
i�ag�W<K׶A
�:�s����4ᏥP�Qf�)�x�/r��Sm�e��!H��"�:����@'X�0[�4Bݷ����RԈ؞��e?�Iࢦ�lA���b�xgD���S�b�.p7��>W)U��S��L��Y �W63�1���g�=@��M�2�`�+z�4*���E���*�bI���h�ZM��ww̮i^�Ν���O"�>����lq�hz�����0DP%�^]��N9yFgr�ɟlX�n���%����Ht��-&[:s� 7؛��4x/}��}I�w�F��ܢ�I�T�=�vv��]������'E��
���5�`x1���u��D��wJJ�?��T�d�4!
˘s:�����3J�¤
�c����6�+���c�5�Q$*B��y�p�t���HBF�ɉ�yUůs��w:���
����ܒ�B���8<�pض��mP.3����>Ҹ9��b���[ Y�øK��+�E�;�R�PO����)؇$�=�����0Ԁ�?�;)�m}zW�B2��Zm@��GH�Wc�a�kH�${JX��S<@v7�_"xEc�
���5Hߗ0���@���c��Qvj�W
�_�]TXM�ԟ�O��JiS|�"`��rRK���1S�>��w�ewI�^������<�����)������2��N�I�W��(1K��CҦ�Z�/ֳA��������Yab��G��&�6:�7�;�/��Y|�E���iT�hiR4���*ս�jw.��"m�,�`�o`�	�a�76 �@ H�UF�O+���� 0/AXV�4�G�nex_����=T�ؖ΋4��4�z�m?N��$�� X(y�AI�xH���}s]�>�l��S��[O���������"M�V`�F�b��'~a��ԓK��Z��T�x�&*�Ij�r��q���~��I��N
s��W�T�@D[sMW��27߽k!�݄�N��JT7I-���9��A �����{a1I�R�99\s�.������ؒf_t�u�P�!\*od���Tf�d~ǭf����P�c�!%�:��	�`�?�����`H>�[�y��Jߙ_I�G�T�aiq�E�a�d�
��Yd�Ja�x��h"eZ��gK�8`�W������Pk��z��m�c���77��W�OK�d���i��#�?��}���㙭k˱eʈ�'�}ǻ�<7� �ό*j�e�nU�jtZ�9J`�&s@1��a����I_:3�zy����(oQ����16��F�aX'&��$M��̗P�al�F&L��'Ͻ�ʻ_��n�;���n	�Y)P��c[����g�I�	�|�:�p�"�&�+ڂ��5o����»7���y���Ar'�{���=��ՠ�1\4bo����9P`PO���/7��:��W���uq�1�FkX?�V�k��r�.�n�Z�����\�a��a'&�l�if��_�q5g?�Wulj�*h�䨯�^4�����df��GIdA6�c<k]���5[���RИ"��3�Z�Q�s����f�����H��%_����K2Tt7�LS_l�j��<���ZR�[�1�AQ��B�hmen����%�ӗ)�"�q��ԕ����������(}ڤ�9'��X�a�"���'�?ۣ˜�*L&i�;��?������c�7!	���|"m�㺗����-�c��j*�LR1Zo�+"�qڵO�t�^#�H�!WfB���٨�"B.�a3Ԟ��lބ�K�K�oaU��뒫 �v t��ކ�l-�0N��e�A�hH+�jWVP��P�^IU�Q�Ϭ���2)��*� ��_��[(����yʾ6�����?�%vf��5l,ɂL�ȥ�ar�Q.�<~�#���|�ZO���Ҷ'����>��.�o^��I�m/��Dxo�D���rC� �A$�.K/��Kq
�V]��_�'�+*Rx��)�ce^��KӬC�&6�^|ѤM~i��	/ �&Z_�~���<�]���EV���pW�"���j�)�С�k��Ӝܗ�5�T,�b�����p�4�/
.���<a�{F��Z�<��x� Ƨ~=��q�Q���9$�b$Z.�jйhC�F˾�Ǿ:.�,�����V�;m��?0��ɣ��,U�D��I�����J5$�.���'�j3_#Ǟ�h���u��������+��َ�;�-Z��VxZ���6s�� ��U�N""�?�E�:���Ɏ9���h{�/z/*�+*��-&���{Ν����/?:�E�e�r�C���E�B�=/���2_ P���8�5o3gz,�O/b��`aR����4��(%j��|�_t;�c�8���X��s���&�^�0l�</��y�rI���įQ2�����Gk��(=�� ��SiL����tZ�[x��'{ϓx����#��3|��S'ud�.�T����F��)���L�EK5�<�^�_
�I4J����[�w�l�!In����WK5�V�G<��L����{�u85�)�5 VR.)��[���؈���W�QQ÷c��� )��o,�V�g^��v�[�Z�+��^ Qӄ"�0㈚�a�ҩ/l�O�Cl1CY�b�gGg��b��� ��~��qؖÁʝ�\y=�Տ�]��
���D�TІ��恳͘F0?f�V#N��Z�rf|L}���1+�-ӭ|�<��F>�MbI#c��%�S��R�RC�ݑ��?
�l���:»���r:?�Ѳq��ң���6G��f�(p, ���^1'���4�jD:'9m�-P����m�N��cj��$�g��)�k��y\	��_M#خ�zS�fi���|y��0�T�f�ӓ<�T�Z��p���e���u+Di����7�4�4����l׊�2d)������w�������bc�/ޗ�=o�Ϣ*]T�i��y��R~X϶�q�C����X�����)��M��/�8`&��+֕�Z��UOۇ��B"���^8E9V"X��p	@jm��FY�k\58�����c+�L�&���^��K�F�;���h�Ykl��@�SoH'F�QD��de��B=o����(m�#�9�T�r��Ejz%��_��$���gʣX��qE���'�<=�K�m3��Q��%�6!�>J��a&�4���kD��_��O��ٞ��(�:��՟���[�̭��<�ud�|WN1uD-l#����t�y#d0W�<�z� �\ ���B�	��I��������������T�Z>x�0%�윀�|ћ�5n��nW��mJwtf�Bk���y���Y���i(��.��2dif޳��w���|�1�/R�А8��2�&<�O��8t��U�ki�� {�ʿk=-��^���Z��U����s��VWKs�;�T*w�Y���V{���P#ȱ�-T3�Jhay�"qi�ؕ�=8QQ��|�5��u��ir����\���)����܄$���K���9��^���b�)���¹FU�GU�DE0'�G$��n=�z:/MZ���|�"���>�l��z�'{	xf���2ȑ�(	rZ&�ۨ+�C����Y�.�i����K�������[�RH
D�_97�C|]@1��|���~-�V�L�C��2ޮ8��4��u�oG�_���8ʒ�)�����=V}k���k�'�^��Sی�*1@v��6�4Y��&ؚ{:zҰ���x^��Cv��I��4�-3!�)k�������}����/�6p�ͱk�?��a�6VEm��-�-�`S�?蠋.6��5�1�IH�i�g1=+��+0 u�=��NΏңG-7�y`ߗ�q;4r�Fa.7�i��2-Grr��\�s���_��i�ީ3�ќ��$q��:��F��g&��-�nc�h��$\����-ۃ?� ��b��mKP{��֖�я��=6��/ot�7�]�诐7���l���.�q��*�MWs,C)���)���YH3:"�?=.�n��6��vz�X�v�ar�=���w/�ٚէ#X��Y�7|���8�:��F ��@��O$����j�;dn��{
�����s`�уP7aH����'�NzAK���[&$�?5��h��4"��8��U&R�h�߯O��Q�����	kG���o'ͨ�ƣ=)�g��J�yh�k ?��6��:K�y������kx*hC&Сe��D.?���O�7q�6����|��Oo��K p2^�Ȱ ��t����zX���$Ȳ���.�����0l��a+ޮ���h�bM�ט�;mg��7�.:=�/��2з�|������B�CAJz�oZBE@�n��+!�7�4�L���8�Ý=��R@�������2
zK��x7.~0�	��Df�>=(�	)2 ��(��d� ��A-�6�{y�}oĻR��-��������8������pM��\$�,>s����X|7̗^^g���je�-ȓc$�%������VNg�m�ݍW�d!,����P�&).�o���o/�s���	� �N�F֩|D'�Z�dXO��u�Y�5ru��+NdӁ��{T�Ɖ*�a���iZ���	�ɏ���S{��,�l���Gv���_>��
��q� 6ma���p1	o�ǜ}��-)=z ������:�K!�vQ�o2EN���-4˻��qw>tx|}/�/�S~��O]��;mv��$�;��?Z�Yx�xE��00�d���kM�w`�t�fٓ������=��M�*P?��V��ʱz2�zz�̼Swh��OMm���HN������]�%���J�T��v{ȁ eO"9FC�nwEO�J��х7+.�G�WBN�r�ε� �ϑ7�3�)��Tdw[�E���������Ck�UMF���r&��Z��ϠPd�3-n���cV���m��X�Ic:
����� ��¡>ѫS�y�U����pL��-;Y,��0���O�.xb��Y�v��ڻ��eL�c�GƯE�H汎��W��a��������'