��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���"�}��c��}1�k��Ϲqk^����%ʺ����N�h�M%�Bx[�ۥ�Mj���9��Q<��=�B�0�&NF����b#���0F[!���1L�*�F�J6J7�hn�6�i܁.��tB�����F���:��_:�@���˽�O��JIt�dC��Ba�:k�R`;ٳ�v�:qf��;����b�<r�+�׿i�Q<0�c����Ա�M6\p�L��ЀMl/����2I���(�}b��N���>������.�ެ�0G�8�C6 ��^*�F����^��]��GæDة�������f/9��;�f��4:�1��Q�CI])g�RU�cy~@�[K��;�i�;Q����!5 �_Ī�J}zŃ��E�BVQN𺹦!\z�SY�~�]�'���!�[��
w�R�Ӱ8:����2NSd����~모$�Mu ��(0�"����'�X9����úq�+������,��ˣu�������|^�<m�2��(F��q\�X�����`�n��R)h�J���0���G#6�f���Z}n�~��(�v���L����(~�oT�`�^������J�O�Fڎ4���Yn��]X���:/���?$
2��?���Q9�p�';�Y���E�c^z�BQ�,,r��z�^|��,�Pi定�a~�d�c*Y����,���N��~����`m�"M��Y�v�nl+P�`�@ |�h����0aZd7H�I��3�W�R��z�t`��k�ӱܥ4��y6��D�ƀ�fW��%��sB��ㆴ� �B7R4��O�AȧĎ�lJ����[��!�z�$)�f�6�;�]�z�()��U�%8�3mĞ(�Ry} �MEZ1�����rQ��*�cЕ��dp�'�-؏Mp�{�!��\^��� �C�i�~H:!}�Q�T�C�[�L`��c�U�C�1�w��D��NPs������{�]n<q���������v}]ZUWc�+ĈF�J9}�c=8���*�n6����{�#�-wt�ڣ���4grں����-_,@ "���y����7�:��B�,��!;D�L���'u̴�Xb>�E︌}��^��i7*��"���MS˄�b?J+ %���3����Ǫ z!�-�͞�g&��-hx��e���������G�e��v0�f�㸥����Tl+��5y�˒���T�����_i��^H�Ĕ��d&�Â���s�B
���B�{�ʳ`�c��T����\���Dr�!��Q����V��hVڿ�"d����KK��9�����v�R��.r�~�؏t����`�"�O�(`����X ;j#J��3�h7�����(,��+�Y^�w�]����@aT�TZ� VW��j�gfD�vtu�ad�𢈻}�sɮ��W���s
�f�����D���2$$Ә�(6Ԍ�W�RAk�|���a<x�*�nX�E~��%��)`L?\�l���/�����#��/Ig��*��ubm�"4G5%��g�C+c���T����	M3 <0��;�/�y��K���tK���1Rl��.�����%c�!����������^�[�8����m/� ;A$A��r����a4��0�B+��=X7n[�*�k�V�k����\�������4?U�t�]��.^�ҳ�E�+�Y��Z��@�8Y�t�iXE
x�n�vA4����G&��=�#� ��q�u$��/�,�+.�^ө���O�Mǎ��C���9���͊��0/�p��£t'�?)]+v��>���ԥ�`���qm�W�F�wz'L��ç��$��W�:
����걙n�Z����&>�
�4z��'�k"E���hd%��X��Z8y9~��D�v�^Q���0e=Q's��\�+'ϫ��5�l�t@��\%�>w��.��TR�|�^���?��_�?���ʆ�3��z���fcE�#C�7���wB�q�����fw������p�"���hD�+ؙԲ�=��C���}g)�J2?J�p�������e��=�Id�2�N<�'���\w��ͣ��&��b�ՙ�/3K��@�SETY		v�x�xX�vh��,��3Ti���6z�}��q))����%q�F�d���D��F|^�ѝ���:Z�и�F��5��Ԕ
�˟��C���ԣ��TfH�5��.
�e��.$A��2-�����"������KzJ��A$����#��������І4���)��2�~\3��+X�+�N�����bR��O;3ǌ�C�ʻ�٨���0��08�5�"ȩ8�2$�f)�WSk���V��Ž�<r
\:�{�֒�HMy-�N	�Ԡ������|��ذ�+&5��C�ҙ�k6x�x�T��D�,x%������}�qIE�Ȯ��M��3��M�^�H;E��x!א�!b��R!+�h���CJ��<��
j�GeA2�n%נ\� '��!��s<jt�k��� 6���!��u����>�����'�lOk���H<�0y��p��;D`?����S[�oq��D?<*:�R<э�Fl!�� ��R�';��G���������!v7�%��Rmc\ f�ndJ�4��V�:Y�ΰ��?e)�z7%5�o�a�vL������ٲd�BH�������Z�.�	��|���!\Qt勧�����mj�����+���1��"�h�<�����K�^�~;����@��<�ъ�W����J"��`c�x��g�������{�d�6r�s$�O�M�G�7��*dH?�{H�O\[�d�U����K����qӉ*6}�on�_ ��I��d�k\Z��3���`��90� +(ض��&@�����F��,0ꎪ-U{'f8ed��&��`�ԥz�vN���K*�'�6�рr���@�~�u��]Z~C<@;͈��$�LBh����� 2�}��X1��B�B��j��߅�3>��ʸ�<Z�\���Њ�8�@"h�jp{�W�u�e0�=�1�Zҧ~��k�1OQ�I,��M�ƫ��-*�_��!8�#���J��M��d/*F��*��т(��$���+�/� ��?� nw�_@� �E�����υ�xܨο�C�<��M�R%���.��)�X:*�7�X
{�*�*ǲ�#.����Ϟ'�^L�o ��gU��A�3�p�-\�`}�]W��;�
N�$������'�r=q����+�f)u�l"�����ߛM���K�۬x֭�T���02���}��mcM�G�m]1��IF.?�bu��q4����<O�F4��u=Ώ{4Ҡ�Ӱ=+�U��z�bR�^Ì~�7Ѝq�
�m�OB�O8X�����+r��o��X��sc���2"�q�:m�?�׊qK:�JBԋ	媍,v����^�!je�Ev�gR6����U���mP*ا�e�+s'b�$E�Ѕ4�Tz��S$[�s�)�S_H�i��Y�N�  ��s��pQb��Z_��}y�ģy�T�g���g&�B��)�V�&ܳQȦ���e�?�>���wP�i;��(���+���b�����dF0�K�/�4�
��i~�}�*Ԣ��Gwg�k�辩˯�����k՚�dW߭��ocɄ��K�+Y:P�o3�I"CoQ8<�"�R��QV��`�"�,D]aE�}ZLg���8���5��m��+s;=��m���U�Z��~ǩ�eAc�(7�A;�5�h�J*Lx-Z���?��栤z.��ŪK=嶃�Wډ3e�]p��t��ڞ���$��{|o?�Y�"#������V���)[���ǘ���(]7B��f�}�p��2V��;8�ݟVџ��Q���o�_C.�^θa��,�<�L{����}��U�G����x�}��N�S?'~*�-@��%���!l`3�� *�>�ѐR1��]����ϙ��=�C[dX�m��߰v�%XW�<:�6Su��:}�Py�Yȼ�6�'�G[]�����|���e ]��<��s�}Ι�赭���2?a�O�$h�aS�]��X���r��[
mh���W���hp�W���Tu�)MC�?ou9ӟ�n/��i�[Q���/�]F~���mRfF��vd��KT��07���bN'9���"HrH翉�i2'����1
���Pr��q�=P�-KM��ÕAJ2U��Q�]	4�ꟛwv�^��g����߂kV|�xI�R���W,B��=*v���C�#n؆�|x�*���f�Z��N]�%� �)����j�5+�$1:A�q� ����Q�m�A���d��Ȝ#�!��(���(��Dw�.M��3v�>�6��4�mzC�"�Y U�e��3*ͮ��Q��Nl��z���1��$6m����Sh�Q�a>4E��'�z��]��T�:<\�JfC!7��]�w��F��.�T�1�N�Of�JSm�������~�Fш�~���J�[��tc��Ӿ��	(;����e���V��gaXv�����o돳��▯7�b��Z嫎��\�{�N��=��+vK�3�79��)U�^ވi�[��7�%��͈�K�N�!�[��Z���s'���)w6jV��PR%#��#=&f` v`��bp�`f��
�Ql_�)��� �W>���#t{;�YJ*t|t��uj���t<��E3�*�$��XG�%�X�l$�*]0rJ�[վ���Z�}�G����$�[m���T�s��0FfG�a[�V�<*t,xw���г}Mˑ��z��	���&�����>��Q�!W�O�PN������ɍBs��;Y�2m��R~Z<J%��Kh��e��z�D<�\�p���H�'��c#�B��C@�k����%CE����>)q*&"n�|Hеt�Zpٍ��T��FTQ���s�l ���rd#��^YC���?����M�.�
��J��U+�\-}������,M*�A�Ɲ�_��Ŋ�9���	m_��r�B���ax�a��LUڋW�r��̓YѼ��+4�-��I�RE4"W�x2#~M$(�����;�W�11���6.���~�$h��c�L��N�W�Z�MО�H����U�����A���kr�%�&a���g#�|z��t���yi�G�7�?�#�24�lF}ُ≃�^�FA�w_)1!��3#���n�C�����X᭎$Y�:�X�ەhP��rGbύ���ҭ�7h<����6�u���%Ǘ_��,�[F,Oӄ���6�H_�D!�����؏�:�Є��"�8����1�v&�Z, ������=��WW�LFumB���7��*k9��u�(8�5܎�lY�1�b?K�5e`=�	�+��uɬN^�Mf�
|�Z��D�ⅆw��[Q/7���V5r����|�����s@/"�_TǴ-�9~�d�(��=\J�ѹ�ϖ�v�c�i�w}=?I�������p� kd<�=�.����1U+���m���BD���*���q��d&N��[>mu�$�_	�	}0�MZ����݆%��.�э��E ������Q6� 2Z|�A���R״<��}����w�X�'�s��Q5��l2rKg���L���&����;���ֶz�躁���vXK'_��ͽ���g��Oj����_�aD�'��*�2�kh2u�7��iRK�c37i��Y��
��T��o���޴�9]:YF��<T�PX��Ɛ��A鐄m�Ydmt�����Gs�hod��z�9���״_r0��B��N���YZH�����Z��.yC����O+��p�ԝ�YݫM�<�;�;,��NY��"	�5�9͑Ʃ��g�pi�҈�D�yO�H;��##
i׭2y�5u!Q
�Kq�Q�}{^��-��U��L�:ǅx����4sR���C�y�z�"~�'p.yox�HI��]��-��!ITDF(��&�W���8v�h��cL����D�ۥ"~GK�tsC