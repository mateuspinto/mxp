`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
0USWSUGxovGsyBJteYpEob+Dc4IxHQ8ioNIK/qJSt0iynPxXszTShiqJeEjFuMAW7SVK9JTQbzJP
8GGzV2ygRIDTrBf33/X3bGoxglMvlUmndy909EB4jy62X/1/FdQyrENyT5kVw6NqIrC2Hx7TKIZs
YCetfE9YYU84qN//8nfIqlaOQvySEAI2TmLyHfDaqQl6NZCzBEL5hU1zCJfZfEzBsc1VmuXc99Zv
K1YeznBw0fDevM5zCCYQXxGTgH1gtBOyikeG8nXWRA+0Ch2gyWZuIfV897QWiwfvd1b1cu2ScqrS
rXqM70L3xwC7V5mj1+XLDN2FXV6pTiuE2HalSASPppiZxlYi0+sGXTzg8XjynL20Mog/uh9Idn3K
QTm75Zaw4yCOuJnT+udBt1w9NWH7bBKxFvWUpz7sgyN5ozYdbf7kUbiR8ZVqZVI2RdDYPSLl+6rL
LVwefsLwYaCwycDjC9TBVqjr8wIuCgak/Nw9fTutfgbE6gja31p2643Nr79P+VQFltwKaI3/MSAQ
8Zcgd9VwLzlu9cGQ+Oevcu7CFd6VrRFiKjEkZkIEUEYYT0/2vU0RazJSD8DNLhDoUDT8R0njSXad
pxAd8hJ7PcP+yg19VmFFuqBYn+wuhknbHA4yMlKCMpBuDPXxPHBEBTILQSl8P3OZl6OXbb6+A3Ky
mShNieJQMuphcSty442gTcd+2TSdk+/SzamYbobcadoOYzYJP2sAgjD8QoA/cznk5A346hY/VFde
7KpAvhOAm+5XNhexSdmkcEw7+7UsaTGnMQ5kgHe9YT6JHbyic6L052Mc6yME4hOF9RZdWM1VISXc
kyDu0+QGZIppr2CGgI2tEqc+CdFWKQTlfUQQGssiE2Frk8Ga2M7k1c3U8e8A1RiciXdBGYK8rHTZ
4WT41nCmD84ck1UNvlRESgNDmMELRWZOWRmOo65MriOhl1qApJhMalafseKIbd6V+1/LQLnmFBro
0pd2k5G9Xj50D29dv3IQhVFfXu1vTqeyFFPn9BuLlxyoiS7Nx73oFsKHI5AQlIZ14f7a6vm6X/4m
NkCafpASqLe/goZN9rZepmTMTBFO5eh70VMB+wAp9MmXr531tuRScClYdHoiyMTti3X5VnD8Sm89
qovd3+MzBI2Dfw6MJW4rTcvtIzjPyouTQN+/jz50s04JcIxfU9fy6zf9vXAv13kGYqoWbKhAFTAo
eq+8QvTk7waBb6aRHqMcu0qU3f6frHCgB1QQ38C7Xa8ESZOBxUb7Q5Sk/w5J5ww9uZAqgDDJy2/a
mHV7iVMpSwJM+N3S7vjt5x+BiNc6GaQzHYtZstbrNkNYUOPiLHxxXyNIutRNjuNFTW+Hq84arX5r
HFL7IruoHShG3sjq5I4tL7FFVUQLSgkdvTUg5eUkasl5mnW5XG2qTqsLFDDjjbCxhODe3n7i2FXu
Mf2XVv2COqNLO3oeSglhzAx5O/L7CRk5n/CDThaL44u+fjl7vlgtSBXJLTtoj+KzftHhFsqo2qh+
39XyTEG/Pc55b13gSn+I/bquu5tdLqgyU/Wapjo05itjLriaM3aCcmyVtNxrLVRaladhc4Gj/uBU
q47cbrFrdi4eu3GyFNkRFqd6YH3SCsjc0WufvCMk3PI3gAsRdd46ZKadcdXPRD5tIi68XiJLqETa
EvyCx836Imj/j3E5ZkjrjMAJWbQBGkG/rsRaYzWMbxhqvsH3cWV6RAStmsDr0erYRzWqQSFiaYxd
HZEBmgRXwLJODFPABs8GYm0j9i7mjDd26oNPlosMdZZREuVOP8KVUzdfuO5xp6RJ67Ckfmpk7J9W
dwzOZM1gbV2fnkXQ7iRy78QnNjfAM33f5hq2C7nv4vy2EaQ9QK8VB+AO58he16OUAKqvgYKq6KWL
JRc4bVVKFg+c5G5FAeZwRaHQNrSphlZfnBaHIw5ZeFfRbJy+I79LvtLDfPbXw22j628mLKxuC3lh
2Lne+yRQlt0cUH1C/FvAUwExKDC2d27krrwuCLvipdpeOK7FpIu2f9yumvDt2nx7SuEPWDNvPxlJ
diKBTfXl5Bou+6mrLU3A7HbM/g79awo4sTCmt/xP0c6oL9q1+CstDSOCiGgL0MqARz3FUFXptR+o
QRwoR25PdpTv5GuowoqcwssQWaAUDC7LIrViG5XTPJjMQtpdTBPmpuv/SkduprQJrJ2Rs6z8u4gH
JV0Fa7SO4YW48Lk+Pzxp17VdOuTF+Vz4M/Rc8usyjARNoR/VIDg3VZ5w8IJeGwavDpLrfsrfmxD+
flG7Asl1aIwATjRQZ7+4RomN/Ehj0WkIeCn7JkMQm8uX3UgKYnjNkSQuos0S+q6CJdhAV52V6n2d
4s1KGZeZ2Dh14k2uVKcvAr8nursxCVotpUNgzHPb1t44lTHGkbcuRW07oBGPw9/NHgFornKUFAaK
eGYVzhAX3KnWLw74V9znoZIVU5Z47ETrYoeF2I0quJUemRDlU6qkti6rrb9bmiddWXt92aTj5ISS
Pp1wcfbpEbP8yS4bqDkF0vsxhc2DEu8RP/btfGYr3u4/TgUQkZRL1U8ZfctQhqSEK+VhGFQSOCyG
14eILyI3zefFmhS4hPqPWGTHULEPbkA8HxBT3KN8d8rbUZ66iaGixB9vD2g2NQBHF5GEuOg1zbFE
iJmqojIkiNeW6fjH6D05TR2hsH0oS8v+WdKamVmt6IKAAURAWLbv2af1Bg6c68FZx7H2+HHS6B59
m3NUn3j4WQVsLbM7ZfaNajNavpi89MPiKHhqAxDCeMO+ADNdIWlwy2fKs4V0qqVx0i2lndo5/vyZ
1k4dPO0kvDml2qIc3nTteFtNAb/xXFi7YT6xSwSiOzpOL1Qo+RsK5jHgE6f7vJxkNKthMNDo1LXq
7i7AEprx9ywdx0PkzaAjdmXRAze0wX51PWH97bnqIq3sCVJ4pjlpCCOY+w8cL+nCxaT6WHp2dRGx
Sv/aJm7IKkIfKY1QuNllejkmDszepXI52Qy8fSizqo9bbxUK1SGvDD1+ZBj8JtngWTkgSBMJMOeG
1/o9McLOCxiqb7XiYYW9e69NDjke8tUpMT+nabwkX+xICiUXL/XgphuQtk0DX5gTS70pEo5gtdFr
UisiAlF1Jew+hBzrGMU/mK4d16FyBWBn72E40zO6HT7O0Bck76SIgU3jPJSJNmTH25RyKaUNJBLw
2UmRJHyWJr3VclmYz9odT9axQSdkBWxa7MxvQIhh0s8jdVVI7tkd59chRquqi30ebcqZF9QLISFS
CqgtnxIFSE8BqPbsduMMBCesMK0yOcxM6w3blxy+pw1Vg/xfVZnqNZGOG7vJAf8Wl71powDICV//
ok5XL3/22vo3tHudKiX4ciFpa+pOQPBWgTl7jawjZsxZ5M8KcejvV/IbsrIGubtLVHWHZYeA1VTC
rhWtta4EVbCFbLAPw/OujmbOi7+AKQGUAVrRR4mCIYJPFVYGVZbiEp0HsyvPvJsqIl+bBozorQbu
JRe/Q4YV3wSLD+ycSpTh2p4qPKq1f5QCz/mnLTovDIp6OcbblvMnYLmVU9UPMYBIUMBuemwZjxMw
twKp1Na1pX4hZuLp5e31lU2RY5W283o2WBJjdY4Ftxs2YQxUA91o+0Eh+UN3+PVQpDifCDyLYoXW
br1YAqZskIn0bD++6hm3vAe/zoLbLxtq77smVlCoZSRSIJd89Up0Ou34VJ5Ns6pM4876uNm6Arx2
kSoYuU+IZRITeS+saVaUtGwedkdsC6yWsJUJxb0TzP9cVqW/wa4SeeJJqTI3awdPW0bdM1Mqk0ty
acleXjsDo7kaW46d1+6QBKIYeEdKUZfR4ZTglubvVNZkiFYOuKiKqmlfCtybmi3f+xXW42rlyxrf
YmfLX+dnsTU4gjSsNRl4CyY57ubWBuRaNqVPRS80k/DOasXMctFTlzddxSO+I3IhzKLtKK6MCQE5
7pa7NLebAeOuJRqXUR5DLpIVCXx8/1pz527VsjEvY9baHKDKB0Fj5w/eYhvqHpcnesD32LXd5Arw
EgxsLChS6UloAmM1sVoW9YqsN/ZqfZJjD/Pyon9CNk7uSbqzMlvZaMjEErlk+2FK5EI0i+T9ORyC
MzFZQfZQAaQVoQ0yn7lzIuHEOV/wFreYpiKKyTNyFO98yVZBdgZAigVI2ayIoI5sFawveQ3/79C+
bRgI63fw1lBu5qDSA6COk/mcOu2a5LbQpAKVzAqLW9Ma90X9En4H/45BuO6kCYLtGut0U5xb5cPn
MuDnqb2i/zv/44ANN4/fEmChgiCTp0yLODc3tG1NYNnY4tnO42cFlN7+Qa3jBtQbWhX981CmNdLa
FJP9J72iMPdWk0reUkyA1hYud+IcVPBnkba10SEkZADRULLj+9KSzFiBXvN+CMYSMZjrtA9zLrca
ST2rTV9ZJ0I5O13/PVaUaILVqQ0gAE9UGyw3jpwlratPr0NFMl/+9zrkFJ6E+LGzWxh41PKjq+TO
V4ujnYGFzJcoqBxIyyplW6tUWHVjEvwWBNaLQbS7WB9YCpSAm/xzwlj+cQJ+wDCRGENPVOvja69C
4q2fomP0KvPJafhwVhhreA9JNSE5UUQmNpWPBz0quVBBnTdHnfGmSurh3wjyRVemSNpzjqin2jrM
zFFuz2rkhpkNsKMqhA5l4e34GZqrEseu3CalKyd7Iq38XMcREJG7cmVgxH9geKVdF2QHVtT67zRX
iFsGQ9atxFKZhpyRJHH8IfGHz6SrBE6IocwSic+L55yVVobEtwDtEJLWv8zKIO7y6hOLG2IeFEGE
zuDwX2Bo8SGWdcnyzV16nt1IBwJgG+dZOOEkMlIX1cQ+6aCB2XSwPdfncosaOdzr9oF/dwAk7oHS
gzXgvwzIFUIi/HrkAiXJfF61yvohKaRIRyaARM1KYTh7uzDymWW9BxmSU/dS/e9C8YPWmu9gdRn1
ijxjOtQdErAJ1/ZgaAHcmQBSe5vQjMHZx9WXjWHvtSjnkxa8A8vXT5DNsleU/0+o7VyHuBuqY6H7
zeBMcHV+btXryPgTPKup+Vli9sKhpLSFEtrKJhUfzTu3UvcUXJCzSVqqSFvH6qYi0XBZF3iKGlWa
bgrMuswlX8aIAw0Wwq0kiX8qsPZYg7aVvmoap9Itvto1TZ6qjt1Mk9+GBLDMkjL1t51zYOcqITiA
Xcwn6i58nq7CR5Nhn4HhLXs9ppAV82/BCb5FSmRTMUjmxg/SUtRYaOELhIJKCzqMmogcBEZU3Exl
wHiGeL64NFKQVtCpVa+s4SOmWa+rdw4KSxGubP9U8UunLEa+7SRpj6gl9ppyRgb5STPTaYDaqWJE
JBqMrAYGU12a7MgXVNgCIqTuF6mzx3pPnzk12h4SN2hb1JGctsl2mHEe6pFdf/8EzZaGiSJEXVDD
Uw53ZBjK1eXy+M0rj+fNKD5bIUudH7LGfLIAI1pB0JXnRmby3o9nl8CT82S9gGxxzDGgYpC/6x0V
xsA9iBFmctj9Iqbr9sOdZFN25+CrVvn8QckMZdJi8cf68icRiaqawVFyU84mb2RJFrvH24P0DA6m
O9ue9GfS1BV50KMV9IQWBcZRucMo3/5bt4Jil+fy8YGAdDy2RRw65VwXdID9nAZiDaZl/nWVCd7+
0kxOu7IBn1IdgOWNjHQkpldW6GzFGfXsP0oZwciCTA9fC51wT9ARpIKVHFxeGXVBZeLhyFb8jezc
d78rx+L+y0Kjgy/jESt2QYY5cqymGz/Lp4Ny5Azk5q5mWaq4eOT3+m1sx/aW21cLPxNByIwqUwbT
FaIpcrVDb8SeVAJiYa4qwPEWIflccQazsCGpJFT4L3H1Y7jXSF0hytuffnVwbE1NH414/kuWjVX4
OrLs4FjQj1HW5IElpweSwUjYnsgnNViNttUaeIHkek+grbfIWdrSJViDXl+6vDZs6NAFHOiRlokl
L+q4PKRTKeiEwy6stwhXC1Dn1txUwuJTkZVaDRQrAPe5xqzsEGdhZhpSn8/8FiQWDIe67h0KsCmJ
i7VWhTCFBY8f2kvXfVewxTgEnVvmrC2dqaBRHaNjVohMzoWQVgIqyJxluxzxsQ4cfZKTtIe2SkCP
TXPv0jirqjDXtw/vrg8sw7Uvv/IsNYdx5z5HEz8bV6WFMOUDXG+V7lnid1lnNTQVbrGXao0aagSN
ih+xSNQ5emuH5ygAH6puKANFdIC0q3VmJcX7R3ep3MSJl/WMsruO/4TPPNuGM96A+AJ2ZNyGL8W/
gw4QBr3o7+nrvUfcT3H6/YO7wTzUsdxIg8P+VF1AwkwiUDo3IStRR0yzj5Itct3lYcCfB11pur1P
7YYxMv2DK7m4twAPBVZ3XyymPK9Jz/czuBHwRxC++teqzEcggfRCb8Nd4zgXynmbqhzSkv+6rMIQ
zlCEHDK8TM7Fy3Mo32F/50P3dfUYadPX3lNIvslJPuGO0zF1+RXrHgv6MqOiBHcLBcziOwq1oTox
sJzLhx7mo+AvxEb8bQ3hVIH2+HHVeSmy1WqKWxGxofFU0dYaRY3kO7jv2TNt2pe1ZhCaHyGQFqaP
IlIn38gyZZE8eOxyuqHfBXxLGiW68vOjsBTRCrlDmpie01lbXtInuuY2BCGz7l3ufdLet8zkoaYL
HsOiEzVb3O5yElRN6715ZwJIrdvE5I9aIWNY6NIOPjqoxkqvdpX95ojFVziSPNRav3nOG8ahmveH
roGFIasG+k+XhGmsIIcUOIWzZWpwj5L7ermONgn0EdWCY3XwstR2Uq+gEKJ/gSnIHKG3xXJS8CLW
IW6JbobImHuvNwIXge9fudsJ7qIBsBhwPsO0k8/mp1d2rZLbbgXTwGEQuSOOpyMZAOxJkvY3fKh6
29KxOTIjokUJqCslLqF4SAhMX0YjQeewLy1eOqgtkDxk5qNGqIroa0CUs8H20jLheGBeMmv7ujv8
nJPlTswKsrJrVMlZs3M1dQNgnjZ7aTKJ6mNtgzQIsshgFLLLbuIQXm8kivwGPN87cRHWE5jl8a/1
X1vChwovc/yldD7okwRPssVTrWkXHLuXByxtXTpmcF64BFCcu1NLyFIo3ewYrursYJi2fov+B+gh
uHT3hTvR1IQaO2kUYsbRCkZQYbdqhD0dL5nlUKcT2IVtfmlSDtSIxueqpWAYYOS605AsS8HzxZ/H
0nkbRmDJrzfiluL6Az+1pyMr0SUCMjqZ9rDfEOr7htFxlHk+vAj0BRC1nsFAc+KqkEwo6TKVtJR1
pB7klhAAawlMsTeZkr7+vYKnq8T+FIhCatUe08SoRZmQn2snwIMEbBnaEDhT30Dq5f/LNzogXQmE
4vbR7Tte594MajnJxZg8LLLlJkx5fwag6kcTpkc4ivhF191zuJgoHg7u0OOJ6PniBd8Cpk7NmRth
91umaKlGKEgn0bd4Aj346mhIKmZrJ+Qen2wQmAu6/Ohdyl+k4y1zukpQ/T5x11r/O49kF6BKSfAN
LQY+/O0i5jcrO3dCimByAcAdbmZe+tfhAzENH+mLHJBDsgnGkSmxD9OhFyDWP62hW9qZYNYeHt80
K90ZYf/NaBJDo/xljvK8JNA7v5+Z4ZqKVT9lgRS1XKNjVFZTxNfuMM3qYHvu4qrcBpjw/uLJWGOv
StafAoyHLHEH+OiVe4s5qjUgeIL13M3bvsSSXktBG0XZfp9XMg7DxnmPczgzfOpfs1n6fIpJKcIB
MzTJBsgteMXCK/kCJoPaIL9MV8iItD81U2h6ECCcm/kI8pQb5h4LvAiN6oh27WquW8FDOX5F0lZ8
Q9dprS/p+7kZJPM2UgNnyFQ7R9IJLJsWwjR/LDJ5L5fOOMey0466DTIODy/8ZX6r9AzWkdxrpnDL
qte+reYBp4NsjyHwAtAUNbfFS0ZGXFfkwn4MdYfAS5CZDBz+qeX+8NNXeNEZN+WVUiGOyCQ08h67
t1QUhQ4eGkwZVtPnb72hXPQ/exNKf7LLkaaz0DQKul8/X7Rr7zH+7MZXCuvg9gy1jmmWNnpJuXxQ
US0WJsdqOYxqT3tGweVQ+jG/a5+mSq2wKSEiaSAE/WQYc4p+o6yitTSpbMr48IVYanWGrw07zwHa
74Fv/QUlM/ytRuqaG9hbxsKVeNVdK/dq9XoOxptleh1f1AR5t+ibaGRK0vL8G6Vy7/JanXweLWGA
YG0o8a2TBj/ONqxaGpLp/V+UyIaMs3aNXQhqNbjIl8kXBbCropHi0TptMNdZ6sJjtThhFdE3nHG/
Ld1ISTLNaNhN7AfsE2JOTonjp5qGDQZPsGePzOv+5v6Gmu3SCgIvlL23tggjebqkCGLYbAxqjKPW
4rCrm5s1E6iqZwXCXGcPXQHxraTW47T/rmZmpq3q/+SiVR+99hBufLG0fLBxcg0ABkZ7f+Pxzo2D
9y8H2gT5qeX0AbcsHF34KnZb2+Lxe6Fkqa2araswbZ/mgs6K5/9bArrpWH7bQ0ebZuawzQNNCsar
vkTpCdTXgahLF6I6XxC9/wIHumkBC5sc4nEabYM+LTbl6u6V8U3XuvjskLxlUMWMn0maOJ/1KHQt
ze1+2TiKnOUdn4DwYL3fJ2ZwKfCpYAsaT6Wg1h4x9HsJg+LZoRXolwkYeKxxMN2/3a4F2EM4LNNg
6KYB1pSbtJUXoqIq6c4VXiuaiRbCiiC0y3Kd33xSFTbtoJg6gfEAA1vgoQAUE3+dg/UwlXREtI0e
rNfVH6BNMa39z5xJynrubPy1GbKk2Gs6L+1XiOZ8IaBG+JQE+ZSFVMS/m1iqmXHInYNYSK+cau4O
NvQ48wousAJbjfUz4Y0olaCqSaVeq5znXYvQyeQT6SQdc0u8GCu2+A9vQioRssaD4wtF6++VvMiV
0/weJVc++1/wAiEBR7hcVE/uArT4J70EWT64CF9+NC3huf87tLSqCuIAa1X7ZB6pKO/21K9vRDib
bVFr8htyj5IP1s8zbx+rtWAs5TOIGgeoRej4TJ8E1buVnEKH2BmfG5ipDv0mP15tZDN9a2soU0s3
qNjm3MhOikYqy0cBgrLU6G3Vf21jOVkvMypeCMBSIFEm0vuSdtbueJe4rmkuDnjSIQ419QG8GvAg
DcY3a6p1gfY7jCcOM4ulvJ+0lSGUjxJPsPtzzX8CNamiwZG5icZF05ITcTuNfb081XfkFdhsoUwH
8hdCTsR8uhIYTLuUJMVcZkLtzCCBcppmFRTyJXti0egcnbCLk8e5tjhTtH4W4znagc1SRdYgpKuA
ZAdiQ15PCCHkPkGI5P9pDUEM5a7SXnd/iLyt9yjW7qJzqtsRpE4MGECJ4trp+YUcKj2ge2rT5PbC
t4fsICFyL8rN+k94FRm2MziVr/A/IGLiMnitzztpJjtNi2c45TT0A2ZuqNGfylP8JymnxUBLkX3G
N35LxkvYij69/F0bfZBTsGmq4hrGVh2JXZoxoFfbVAqb0LeYXLY8Weg0Fhe8WJDLpRcXSRRbD837
/K8nJh8dYEJNygo+vjHoqCU0tu+EeQLRtPxE4Gs4AqNEyLpeCEW1odBT90gknxRRFF0lGbSRdMPI
xWz8IskS6O2rMPHIG+Um9Lqzgk310ybWrUv4t2qKl+Eyk1UqzfmRHyqlZj47ob+nwWJhxK4Hhsa/
OwOgUQ1WeXElAjKtX7Xb41LLj+rC3kQGyTeWsrLpIrkcyubJ/JhL+DtkKDuuKaA9KslOcaArpMQJ
9folm6JjpwkhOKedpn/0Mhxgp+9ZNU7uUrYWfDRyaiPE9u/9fc9+oIvfD4M/gLPQOi8SjbMg5Bpg
NmDwAbp94STTMjWVlu4qmuPbmiXf4H0Smwzr32cms8u/xB1caKr26wxFv8pCF+elxctcJC4Weo8T
zNGY7+Mw22DplUvU59xM4HKI8Hf3v6QFb5P89t7qp88b1O//+rIw2OFowPh+gAlxEcoTV3dNwLQJ
sGL0AWS0Cbombt1SsDk3Ms3DXaZ5iU9DjAJJNdT1uL7V/VRTElVybrFzVGTrtjXugY7ue/l9XcdQ
dyPPxn6FDyUeGJPeRbb08A+TZUN/2YhEtdOMuxEmJhR9rRLFkAP/IiB+OLisSuVCFYJNS4TlPyj6
ggLAqw463WC1KFjbuW4wvg0N76EyS0YGVGHAFCQR5Wacglf3O8wtecrjLQu1iLulY2/o/nqobCDe
qJqQvKojBsiwYHDFXnKEWOKUlt9kFPeXExbA9p5lhPX4FCKNzRNkd/chzAVRw5VIcwfpJTcyay29
7RTisvLu5UsURgozA+OT7Ov0FWovGPmrAxM2DfZIk0eA2JRoRviBVWA4Wh9U3SQ7ruEJCl6zGX4N
Z4dFb0Kn+CzCnX2GSyKfSIxXp5VVSHlMs2wB7xMp/oczZ2ajoo7eim9WHLQIw9TqBeZe367q7toF
stcLKlUCPSs9uMkxoHxSeJhtNT/i3wMzFZhoQq3jhVmg3vRhWmN2+rUytiujrLMR/Q8WZmFwLD8P
EgHtz+V743Vmiexi/U/2Qq8zqpTs+vEMiA7Ul9ahFrUsrfZ5t2AxupxbOoi8GUHzT8Ycffe/wTNB
ZpmCyUgrqec+LIbeth/Y+T/jmqJoSSDn28Wfea6Nb7uwWpQu+tSsL/L0AlSQhdDkJlujkT7hduE4
/eOkUb8c0jA5d9nNRJ1c6CxT0J6lWnwIp7XyCrs0zqiHNtNOVKTRqQ4xb72aDkmPH/3k9puDJagi
nNxRZHeEn6UmHBTUUSlqDTJwF4UwwBN6ZHF/81fWZj2X3i0vFPD5BNs9yANu1dTUvo+zqihvSIKb
1YZbKFGOBaUZjadSAg1yI6otnhKA4La+igGmFlua2hhyiWPBIOrAAPajN/4abEEIe6qiSg3KhuTe
OuXOTFzSh/pspwDamLCO0yiSEgm/5L68b+jeQfkDok44rp2YM0xEcOrn/IyHLl+zTi+gGj3BK6NY
XmGs5z1gXV34WLd/V2U72L48YqMHCziLztQA/wxdQM5psseJlo72WsGQWBphfDsYC9plDICe/jwI
P+HB5/Ns7ljMtwkniTvrNeN+KeJbNarBMofyAwNJ6Nad1610XiskcctR2aTrqTB1a27jj8HnY5kg
U2V/M5sXBOOV6A8uIQfuRl+DPul+z6AXQPcKabZA5rLL4HcRhihKt2VgtCyeAaURUXM8ZSbQI/Tc
0K6K4gyBAp0xzEE0CHqIobPO4mIMAbxCg2NSw/bC/y2O32o/WMcuVkmlB4Bhj9kmll9sVs5dVtH4
Hk+9yzT5+erkQuUxvuMVEXehpLxfL4BJWAD0+PUPnrdNqkUFVTcDoTSiyOu09Z05D4xqMasHYIgI
JNb6phtWQE2yxBiBRTeY4b49lazzOpZ8thMIWw5vijzndOXlqa8Z09uQ/P8U7JaDavNKCR4YNTpj
zrvbu7Fg+Ih74hjcb7Tv4937+AOKkKklMNko0Czmk3mJsra3e7rPddFV2d/80xG+U3k0v8U0vaxO
AxrzX3FhQns6zi33rpRqmYShI+iWK9nEPA9GHdaJplaa1otIoolHueNVZVpFCb++/fXZ2l2MVaCy
uEAAAk9IZV6FMxGBiiWftP1FWdLKEqbEIdmx0RQRlqF5kGki8QfcGsxjwuStAQ5V3O0+XOj7EQfO
4s8U4vzR+cbO6EuMOzSnj/UYWBy5Dy9N8Gz3id2tJbrI5c3q90Q9IpYEsg/NUbFEITdSGeRRq9x9
jbKQweuH2k884qrT2T10rIPdrKe1MFGzKIn0c1GGRm1zu8gK6501I7Cl9fWyaqqBrR3Vc+V/5tCp
BdecdW6HBCjfsi0lTh1gMObrIR4tiLgJt56gxCTCiIM95Lo+Uz/Hg1cyrxqjt4plihmzeFLsXlIb
nr0OrLMLMlC5x7N/AwsCDyXr0AxDvtwwhrdimOlAgkccSOt5cRjS80LaN+Wn0rlgMDVJXuS1ilxV
Xv6ZImhv5EwroM8C8IJukFZNP6sN7mBYP3msWYK/2w68K0uDnBN63jxT3kA4r2On/bSEiaeweWrO
yj+8NA0Uq15xnO9DiOpUSTDr7Ygx/zTrYUY7JzDsQMT8HqlIawCJQL3tlaooi+HZOfMPRYMM3lh3
ufxN2VmLvQFWYl+UvUss9RPTAR/EEVIHr6xNMVpZ6Ln4yp+fXfDX2G7KkJ2EgEzzOKKFIsFHNaHB
RYImWrTfy/+J1JQlYcKbs8wmd1OTeo5gjxegia7RrKKz/nUkZobQkZjuDBl2r2/yrV6n9bspMWVn
C3fMxq39aOQxst8qLtTYgJb8GxXeBmbmJo3loHvwCb0vjUXYW9TACKj7u1kDlx7//Q2bxB59ILmK
bn5yVmPjCPLmVmdQBSI33sYAPk7TfElAYFh3APVfIQuiwCYIG4kn8mODpllCa9CxblThLmYNA7+r
E4vLGbTPA78+FahEyjtePbInuTYzrdHZ2j7qgM0/zhWnEEPQNEF7OTeZPDoHEczxOJ5jMrG9/DyW
fbUf1hyt5/SpPXUyrnbWvujgyUanEqwEuxbgOmEvzIS8wyYZfWaJbvBAcIzq+4HtqKDmoLsq46ev
H6HeySNDlN56NTM7Tb3qQEvPcu6WRGIDdvHwk9LDLjOcFsBufLWYe6sTD2HJV7/rQvrhj1MHDJPl
VTfNso99SObSCxMNWlfBTlkvA3sft/DTRMv8FxqPCxS/HE7uR30efOe7NwIszlOZ8Z5DF2OCmuz/
gmev4GrmWyPTG4fksLSLGbzCoAJCRq9pGGqGA2or+sXLjuzeU8YxCXXLoyaZNm3Oz1Rp5ymzJFFd
lAX3AFYid4aiabaWVA7l+n7Nnuj/TVHotRujcgsbe+a9Fj1Pa1eUeZVcAS7gaoA3PgLDVF8yYd30
7FMH7sRvGx7DNvv061TKa6KnAy7bM8r6TlpoV0bx/2KDb3ru5nRZ/DuYKnyy6SX4TTMXQqqmqNGc
DwUBWXoK24fL1XuLq5ok4TFRHEDg+wqX8o3FrlMxlkAAd8vh2vwWFs490VxkEHYotatz0YvaDqk+
/ZTOWoJP3bpOpBdxe25fKH7qtLD53864yUL/Vpg8maAbazIM31MhACdZgYCUsF8oC1eqicviQGTb
B5pZSDltyrmqvCvXD24LUrxijxG6CrwgWyGy7wulM8mtJ0vvPx5Sul29mBTqgeLOjt36kbF1TraM
aiuM9TGnRAcMvHsF9kC0kTpUk2BSg4qEKOeMDLKhIlHJdD3ssDXAFKLZnaDo+DlrwsvvRz3AEpTJ
fH3I4zJGKSeJ53IyKtMGHecszY+j5qmzzL+UdeabYGJwQNhYFMw+PGuR7qXNS6vTdAdR2wsGCjLf
p7FwIuS0UXzXwXPE9ejfS8UbvsGI03lEsxyTT4ZY2vM97p/4CH1YCgV9RRPFfO8v8ODnaBahdRU4
MVKWPAJNLioSTwRnW4Cqx2KoLdt3rQQHINQEhoUVhZJKMeXZAY+hRJthsUjLANTa6VLsHvfx9tT3
fdJaSt3CBPSUXTtYmJuvAEZEwIPldrvHp1Iblw0gUL9i3mNN9P265ICf1cIV0UNNn6gapup1OlD5
V/QMqsi8j6tUM/dEe0bVhxV7Z7wNJKon8vYX0j/RWbQyJckWQM+wCJ9h4l/TDxy+HGzUyuUiio3B
/DDL8FRGoqlFWqumqIVJA5zgV9RE3a5XCg9+498lNwlS+2jabWoAJHlFyT8LSgp00RM3OfXnlsPJ
QsHyiCcQyo2mNtQRNg76WBScIbRdtyi/djv+H1dgkA12KaAUJc/DKb4nMr1bLIMej8Ibe8TJcJ4s
8AXlqg6Q0nLXDJgXhpBVMAfK85tGsaQvOFRFL31zPHbDu06z49O17II1ILQSzE/Bz/hm7YshkqSP
f0VYOMFBKrHhrQvsxjgSGzuzZ/HXpR0jr3YPqYef+x8wZqKvNlk4a3oEoX8KztnGOxSJZZGp1U8g
iK6Xm3ph5UmVZ2dc6Y+J874RO2BcV9qnja5Or0X7lkUBz1G+D5iNy2IRfeJ6qXsDVGkWnbR+SucN
rRjPlgzyzfGLpL/LtGK0J2xGOrq8tfpmaro+aiHAn5ICGmxT+Zu0awLUrvuj/pfiTiiBiW3j+4b3
xCFxJb9K6aO60GTGylelaKOqg7QRzyX/ycCSjCev5J+Ch3ePeAuP9sprFarR+tZzOOtvNf/TQD4n
m4oDgu/8mLlunRquuwDiYIkvfidsk7/yWhgy9s7R+Wg6wAI/jBdosn26ELz0AuQXi4jZhKKsnV5P
ikjGXHBZNZX8MyOIYY8fVgej18g1fdBB+SaS2QeKYuKS3nS8Bgg/N71PmpMQJnAgWURxGfzaYvx7
FF6mo8guzH8yi2w5xegrOgXHqzhGcRze3U2/xZN8tkpH0aBlxhlACz8YwCBu9duZ7xANKmKg7gy2
Xcbaj4oPwqrJ+bBWadszet/BAB9fHj4jeOVM/a5UYO7PUIf/68Nz8z2iyZrGJMwVqK7BVMlaopQI
/KejHzaJVL/xhDCVsE17XV4HS/JYEMSpnVuwTKfjcsovwkYJjf7Z7bkbjL/xasOU9MlKDtfdc5yR
2A5LLvv8euTcEOJbhLoJ+rRwQo+m8PCHjGLIq8gg4U+IK9jggG9yJsuByot4lM7Gu4Y6xsnvLP4N
KU8GshG8Kd7E1Wb2HWqpLHmm12mMuv9kdLSEcENl3/pDw0KyxUsf+xIyUoHK19jSsCUsMPShaHWh
0yP2j5C0/iw1ecBpgCf8UYZjoQDQCiYAVdA+rFSHWtscojfay9CQEJP1g22eE5BwrPG7dKybxerx
7OmgN1BOIym9RV6INNuwJ70WQ2xfP78Ms9DIfxadeNi7N6+KDoooUKU0+isl5585Boli1aJWQ4X6
2ioLguwzOLJ9elMj+KuY9ZTPf3eWUYUIBP2xuMEl7hB4aAT9tBkKeegMdCElHSGjoM92mOKvx1C1
1dya73dU2ppC2efZWU+77im0urT7ho1a+iI4DF30WoioJxXspMsN6EtXFUJ1BdoSmKrc3XFZ1QCP
oloBvoMQuTbEEB1+tIxBm7jVkE/dwie2I80mq703BFeLAt3tw+tFfrsemhRYLRdE5pdP+0NyZXFk
p+hVFvaGWVu3Z0aD1Xz8VcB2suT4L0u6qkpc/HM/8ujYu7HNX7dhl2Wzx0UsFRtPjEM2/G0h2fwZ
Ihp+12J0rAmozmlR4zx5+cCnFgAzTGAR6b4XrgE3/ZLr3j5QosV1IRn8/b6zbcPSzxOBkLVH2PZS
jd5yQ9NydDEoQfCz65EmvbDLqTODFvdq8a7ok/brW6GGae6kF3jWsFkh8lFUgBULdSsQiI7PmNpP
vLIHPmZT9GrXi63uEviJ4fpXuByfh+Jhycjtuaz2neiFjTonoDjbIYEQEIJeGKKUR8ejEzezk5Bp
cjZ+OCg1kHtXO6qsswR5z1RwdJE2/JXRcK5jzEYsIhShXezPEm7CnaABfbn64SYGp4hQpSz9xBkI
FALwyJdKsjfQwNMNFTZg8PZxqQVOmVxSDROj5Ls6KtrozrR/A3GutY2PZg5aW36Sc2K5WdARwl4S
fs2ZeQdEu30bu0K1pV2HqmdwjvH77/ONP5q2vTP2Hhno+s14z4x72STWC3AvTbdbXOVAq5+B47ZS
MCrl69Ev858mjddANDH9JbEBIIqCnH9kCdOS5wvoaGn+HEvtK4J6+I0H6EG8Qe2UCwtpTBfR0y3C
FoXz7Haj6/krfLeJBNsNujs+Ecq1UAVSIAYRoCrbj3KDdGmhadgRSk26NveXAeiChURSQNvVXhee
LiaS8GOvXsTCddvgKU8v/4B3aeQZOZG69Y9uv2YlidPmEkArqvlUa57CCg3mbs8HQWi5WrhpSHVA
LTtxLmPoXQaoFhHLpb6etozH5P8wRPSz6bY796/Ccn2/Ub1ueYdyXGXRTP+eZuQhTRY4yuw3+PKf
/bC6XmfpqygbHck/r+ZQT4SX20VxKIVAhwreZIt7ksLH3fDtdSMG8DkdQazxoM1M8/x0DnC3/i0P
MXGM8WtZgXrjLyUwl2usx618RegNi6gCr/224Nh4+U2bmd6pLOSoNSERMs/slnLr2CED+TYKwfKx
n7iU10f1yfWNye+r1E+suLH7XIkTaYgO6EE19BMGVcp0PI0iOymm7+GslE+gJ8+fmGOdYEOJhgbF
cHXVTJS9sTi8SjwxxyLQpYxcnHloe6sDMMpqYE/gfu7mLHYs7wD0fzK56w450fsZTfstSuplVv0s
prvgoAZDrC8ck6SOIFIiocbTwnybTwSahndhExe/yN/ahk3Hw5TlJQJt6CG/TRSLeNmuptgld5Bh
VxO2GIkDPbYsmOXQGrkBj6bx6Kx0eAjXlkuM1cWK+8uqbR3TYHR2Fet5Go74rtfJ8rWuNliCnqTd
wDHAFVVmQQtLdvjPOHgDZVYMF7/0nDiAFv5Wbirp+d81QmVnHBOYKchdxgXuoxAKSz4mc5McZ4UY
gDFb5teuH78Bs4AcI1t8tZDj6hgtToxV823JI2WEcM8EFnCYNlF0IRxmzdtb9WMMd1pln8C793Mn
TcTkGpn85EXQ6xS29tKsU7aBBt8QdgY6XRAIb4S/X7naacG2LtKtWkJGNiReKcYv0AXbY7lbyBzp
/4CRf1gnVlKSz/HMXGrJiEBzs5s/8dB+ZunErUTUMHfyFIMkpGKsqXyhchRRVCHw8KtjLu66usBs
YMX9KGXItbWAelKLe8BlahRHlhzu0WJCn8mvHHMgQq/jrt+dD3CNgiXHg0QebG45dbTE02pGky44
7zW1rPggXFjL9m0jixa6FE3KOii8A+k64P7Kk3nysT26+NHzi6A5S3kWPhzR9d3or7VaABTaNcOh
6zvIL8VwhbnLhP9ySLjKsUfMIK17KFtVwzEDf2k4kKhsDaN9L2NRSqfsUmrYElGjwWEWPlua/7HV
jkh2gZqEtcZvg82kukXcaaEiJOimXa+jhmJjAl3i27OgBHr8p+aKUijeaLzMB4Th20hJCBTZBjz7
/jDZZ5YOJc2cCR0EGYRWdZARXCB5mz3tlorNp1O4riZP+F4iHrRLJeStg+MbVbpSp8orXVuVi205
zErcNklT9Hp6o6YBO30TX8SWRc+kHa0RFsEw7jKY0ychgxy8WQBDayBqYPMiLMBq/LrP8SWVYjJI
YHtdQRQOM0S5PJE0y6LOnsM0ycvLdpfmRBqVl/Bc8TteCt4g+RWJSsPdJbHxo6/aZ/7f1N7loqLp
AOZh4ivCJkY8elHEi04EzD+ffkLctGqZTzG9YSENQJdnvvxVpDixboR8mE0B7pit5hZ0zH4h0CkZ
U4CIqnlk11MOVEY2Riv9LHz57FmV6xeAcaNHs+aWLNMFnPOk899a3q5c+Dp7VXm1ld7wM51dG3td
K3bMSoPLpyP61D4QL0uB7qH8sh6NXVPIbIb/eLs5eGYOsr2CbI08AQ0xuJexAvpkXZnqdMIp5LoW
FEjRckuBqKN8vIpDLrNu3b2jKvlW2qsQ/lwu/VCXv5XJljPaFjyofjNTAI1Rz2qiHTwp6rvH570O
zNdXkY2LL+3y/Yjp2EKU9LBR0krTgRLasY8RBrtB6zaclsT8TeLVBJFoFgBWNLxoAKsDAT0MXxhG
5sZrxZHQAg6zY1sAwulHt05CsZ3RBLiZ4oX0oC/jCRsV2h2iAhYGUkR7EQDfDR51BXWBALb8jI2e
f5qAezksjUpYqnkiOzQOpFORxCEe1sG4o1/STFolezIDIZRgoYKkPafs8k39is0RPgqbT6GSrvuJ
61n+4gDytP4PYfnkHr/4G4PvqVPVwHfn8LCtdYsG5ZAFW9yGyhbVubSV0vago8xZtYN7OmntPhW0
5PfO6A/PMDMSPD65iSPrGuh9vysvRjj3RfX2rOlS/pjblVjC0BrVLrVLfZ4zK6G/zeUTCyiE/nxX
4D0rkd4dbKRUhMiUDCEATKD6PSNJD7qxFj7O2eGZteJVJNf+cmd8EPlW38q0i7+IDN7IU31F0P49
AJBp9yRijArivHLzwm4LeVGvDJXe1fsWeJ0fXly0SP/J1w0/P0BfQn93rE5pVbjvi/phq7RnpPn2
E7BcqsCnfXMCv1eeuLPyHthjVY/vfhiTfx5eC1eQi3+1fwyBUXSNemLBjrmFrR4SZxSlwpmngzBg
7kWJNY9r5MAyp/MfvMKw1jiQmE8K/bwy7N031JH1PXJGjuEOWjXWcBwyEY+7b5dtAMpCxEirzec2
3DNSWSMOtVSNUPBUzEjPiQclccMu0ej+Lod04rLQ0/SG93cX+qmpPlM5MRdNmUKoOQ+MS9nzZoi0
1ubCvhF0RxW2cWygHC4a1jVEgc2A0LrCPkT4XoHIGkYCieCz7WHcZI6PcRYydhWdm/39YawW5c/5
DCbn+uAEfzVKUDJbc47qFH8lhpfyO9BGjsAMkbBSV80dSQlgxoWtFkOwevO3vKePie4UudDKISmd
pxqQzF7FrzOi6wxk3I2BNZrt6UXew6BKu/PZbQa63snvmJ7N8pRZ1HiO5RnPr8k1xLsyBLZImjNB
tH6YzJN8kjVQxZ5XPkcYYRu47pvquNfg7X5gr1hAPhExuOVA4/1H9hzJun+NaddaQu579n/z2fhQ
P8svhZ5ppTkMotdeMweDFrbzSHo9pWRj07riovDKMShXfPMQNQz3pgei2FU7P0tBbRXGxp0jzkde
i6+QikQSaGBwDXsPqSJl3wF+kXxfW/WytjcMMB1WZcSrttnbecYpKgWfd5vYj3NzBNN4Hu5w946K
Fdtd5xxFmlpDZLLdVNx74MQNtulIKwXsfE9neXFG1WR0ei8mTuz+O6LxklhOGnOfJwjp6ctLTAAG
wtOWJKsDVdCcs/Ur1yVHbljMLkeJoiXEnzVrcMbf8mucqkYz9lIyDrrkFuNgZbUMsp/fCEr7VGD1
+7waEQgnwMcy/Om2VbWNXPv3F/qrFsJh2kI5sx0y20VTfFM+JvJmtOoJpa1+4HZnBLbe7ZIKbcgc
JrhBw74n2/y0qo5AGpHNGJAKtrmD9s/jFqOiEdQnN02q37RNsaFlmNe2gJJ7He/NPIg/EkjhcvHO
9Ga2/b2gOw5RbTOoGk0CMfa3/XPxTr7Iyk+rB9Wc11TTQz4GDuv/EUSEUzkbCRbUWNeRMa/1icpb
7vnu575Mu4w64Bs1Krst0vyVHcH2Aaog8DWYzVmRu9s6dDy7zKOPjMszxtuaoNrLiT5hCgxUfbUO
zEf6VtWN5aWpE8FRtJtpyCueFr/FBBxTo4hIC8HO8OdTFqkRLlfpS9b61PX+/Ah5LpJ0aykTa7G3
mQzefbUy0+lDdkkypAr+pQ1hbWrhNvWIaPuymd7mxYko/l+X6T/xLdGeWHM6Kho9Wwn9GLNG+NlU
WhIoxvHZyU5RfJ3gEgv0apRuGN1r4s/KHB5IB7r9FhJYfr+VQOjhBRMBNpZcgg1kzuXjLjSpJftE
JzPgi4BkvrnWWjzfIhod2/v8wUWg721FMRnzdvuPHYMoOQyOXFAcQplHJGRVIEtd9EPxwdwqA3FT
pFlxBZBD/2/MLY/TQNCEW8mM0NzDJWE+Nxfi/jh4J8ecCxU9ltRBe+uyXddg0PNSEIMabybmjFwG
n5jr6qMu74EC7RXm4ARwuaDmdeD5D6Bv2Zxshruyj5c3iFihWrescnF3Iu32lVNmT7An6nDttIo7
ZHRU2g3EHY4lsgNlitdblo/qxTJwFfUqBls7N7qd+jkZYRQ+upeeaSsXB5PEyfp72aYXkAZkvo1e
tmDt+am2xaPnOkfOGuYIjSBWEGcKpxDmmuvjsiUXV+RVPH6ZzAi6vOo2KIa85+B7sfxElFeVLHCc
G5BFvnCWylLhTVqo7gLGp/PkyDfNLuDF0+rw4J3ki8kZT67Z8/L8sWLmyjP0xQfBuIEEzEH2ekCx
i5xjaQS4ZVMGqgd8wliCI6beqXQO+lenlzzxFaO5OIm6lwJ9XsBaHNdiCnZUccSvnXqrxJEg4+me
qqFAtcfeBkTO7bVCrB1A0yLrb5SGuFbZJpReXGxTfKGR57ybP4gG1mJoWhzfiWj6L4rhDjVarNPB
UE0g6S+uLW9ZnS39NDZ+s4oBvdjpeh7xLBnf8xyX9wiRFZPHt1vWw9DRcqPc/SaAMK1KU1IuOhzw
cGf1VM0k9pot7GokkH/ijLMb3odSa9sT516lPYwLMH0V4AACgjafi5vEEtwFnHbBQkaZQh2fm+Su
eBQr3dTCekWPH22/dLSCVqWV4usZyYWZnaW2MlSttP8D8l8bHbRCC6zF5NZdBBZNSUYvBBXr8psA
nG7e+q3f8pJE2vbOiFkUQOYq8ETPt5N5XYXX4vyHHCwt74/y/0ZrShbI+2kTFYF5/atsh4pZ7Vqd
alziCdOGs+E0kwoQ3nTYTJgS+vKOA6DHMpV5ycw3REqupCmJP9Z4OcHOhlImNLCVOwWrfLlCupgi
IhCnTEfVGwxbDqBE0w0bTDO0qt1YZKb3XdnzGhv8kV3di+Wu2dOyVZjlFz+8GXMOjXKBfudGvRxR
U094LmLDVB+N8P0W62UI1Zv3vBVHm/n5f+8ZAoNCVpsz5Kv26cVGF7Oy2rlOysbGfNmQcYduf3H6
W8OT94K3mLkUsFMzSoKjlTU+/Dbj0qF/YK2o6VrEVKPSR6/5TLbL3PjTUvT3Mwwh74ZkZeH/K3RM
Jxh73LEY/vsL1gyqIZlXqDSdx0AXcdRrXfFsks3H78Jy+K8v2eioIJTCTZCafO7eiBr4oWy75i9m
lWoenQGGdfOBd5YGNt194b6zd4G0VmSelXd1ZUU/ltk6GpHKywV0OCQeNsMEuod7iJBzsmDeqJF3
795sU8wwrkjdaOfEu+WYkook25uOfVmWFwV/1YuA6np2sOBCCoDF2pQ0uYNG6Z187/tHsEU4Nm+N
FrxEXBpRffDd9Ca6sP+qeBcuPpOKbsRrKQJDNDfTGbtP0XlJ//D8Lr/g4aplrctReIphUb0pHyQY
WDolcbiTc56yAXesowQjiS4IF3lxl2r89Uhz5RyXjW4BrHWmZuYxXK/w3z/Mgj8Ixp0dWPW7bqKJ
WjFc9JmOYCpDWNDU3UXzIRhCZfgE6uf/U1wju910o8WHE6pTvLQH04DGhgiU2J/N5F/tFJ6vlTTM
L97tcObk7UYjZDuY6/qFeqTKCs4qlr4nwK3hELsp5NFYmRs6vvbPkY4zlLsMh6Xb/ADn2dztsPqF
UJAbYiLmtd3h1W3ugwSTW6FleMawIeFQm/Tl3tgPCq6ecJtdNDW8aZAAjV9F2kFDjgy1NeLYuyF0
7/3ui98qXQjmgjxuvLEKyit/u5MIi1jdRY2dXB2FQiZxyYu6P1W/H21e0mpJAjBvFLrsJOXonmHL
Q2KAQqfLG0eKMHR2NLynG7EUJELPJIhjp4+dE9dcoAxO47wnsN/Sre0Mjumzbx76TULmFerygk/O
51QC/Dxe52ZX+JBdSycreeOswSPtr21Oxgw5ZYZ14vHInrTEHCa9ACmfj7qfc4+zoD8G+sjH7SKy
k8LTzb9um4/5rt6nIfAVmBsrVGn3xBKI3+1Eu2kf2TJXnDMytzk9JIuxe9LuCSV/KmOyTwFbYKMi
C6KZUucHQZ95A05EOM5Hg1vjkjRamtztYzKYupiWzMeR80cMysj4LzJsddLhOGqZtb0g+s9fmYkD
t4tjXxzifE57exOi0Qbsi+PlGuXIPeTJyhZEW8CYszpAF9LbuSapOCiBTOl8kRgpyzuZ76s3b+YH
GHh2rOCuu2V5STKsftTtGRjImnV370xJ7bU/KG0kzHJQyYgEbTuz6kYWXtGDZ4ZhQMqyWrsLyXDe
3QCuwiF3egYLL0OixRfoEkaDgOHkhMayqBsILPJys9qd/DhlmXW7y1DghytVWw01idKk7afhpxie
SQ1KL7LMQyjkdkNiGHQPUDhuusrkr+OU/HEn9AwQtF1IvQV0tG++jeDbAebCDKwAYsU54624Cs3o
QMCw8w1MD2z0osaTBRCzgO23LF2bq4L17nsDiFyUliy6CjzQO/cnuMFJW3gkisJ2I/eJD3DqeJ6r
VYuziA6PouKvW30T9OiAV5LB4mRJeka+4MTe6ASX5dj1QoNYqXIHiwAdmPmNlCNg8wcOjf7F2tEw
u8Wj0hWdBdJfP5/mP18JSWH37DYqR+SguJt9ZTtt24xgnOfLTOZr2kmVpSKyPr1SJd4gW5Al4J+L
OLTxVLhZwxSSNCDctfybqB2hWfIrLWM5EAKI4HRQCbSmxmpTY163ej0dD7aC5j/vMcqfKyXEiVX2
ElwmRHxs8zee8LhGs5BAlHxAyTgk2NvYz2f8i3jLRAumSK/aT8VqNMTSB7h4/3pby1uQU6OZdVJ8
M3rjyNxtfY9LEgTquuZnm9hbYDh+9bdl+i2uoFl3whaBRuSY0hbj6l2Sid8K2zBr/NjAxLaF3/BK
/NBL6S6bnjqs4wMJVjAEX6RaXjvZyDT5d3IiJUoew5ttZZ/OJIIeox7ZPeo1PT4mZ0zvrpNdmIUT
Put+zI87XiPWcwNVEoPOGkLv4nolgBAskQgU0CDXVvNPhmgS0xE/0t7Y1MRGcxDHZ50ITEkaM66T
yx/2ypjxsgfSnrz04OMMxAUr6yRg2fYxMwG9jdY3gbBiZRUzhRPg175o/tGABwRbB4XUGsOPbemy
wKrrxscEp+VnCLcdPMHQ4Vb5du3fFPl3uUEhM/1kCRFoD+FIKI3y0Vt1vvn5Gk4Ql5hEk8yWT+KX
cvT+vMcE93UKyI4ai1ri7d//wvoOS9lCR5g4aUjJL/4WOLPqiLKnWh+hWZuiZizZoXh4GaQ9l6rh
DcKd1i0kHEnNcd8rQ5+DXocqY7qYdNQoF+FfwSiIePwk/fV+R+qSU9ZThUdbt3MiyIJujjWIwgO6
Z0B0wZi/MMn+3WhTO31Ek/S8MxV/l1G53ctnFubQQoqLK8wNS9Kz5Lrgzsj8nlgeuzPqLN1Z5GjL
aGM5Zfy9LY9kfSjny8iW1weOP4oO8KxCwBu3HNR7UZE685VtpQ3nT9mpjwXDGeGYvQZ0HNdAFigz
jMpAxSKC/THdF9siLv7rFT1aZWvG2H3k/Sv7wHYMzfG3hdor3iXaKKaCdlfNcyY7Q/Pjm1Le+Tly
K0r+7HMZHpztaBhBACwnnoMC+21sAw9L9Ow9HEnGNaXYLM201WlE681ErrXG3LzZUVzEI06VtneN
tGd0RyNXCo0otjK7jLCCoLGRFAVhR35xphFG/+5bvcdpYLPa9B0yVCSIMd5xLsVrpiWbO3mzB3bU
q45Zvr3NAXgAnAkycEqjBhEJUCcSPtvFZPMwcf0VQ7aZEbTmnOv9o7JR1N6/IdeaUZllHKTS+qdK
n4es2pNTsLejbooCAq0+qhopUlqbx8j48gfpg5vBo9LFZlcquHJIlr3adaofr82/ke6iHKeQ7S/N
hpSu4Rk+q7XOPEjIDkSav9xVwFjqcoEGKE2xT4xAR1ccIUc+C+wLUv1B96zbxYJIYB6Z99ubZm0Y
i2b5CZ3sssz2QhA7ZmpuEXXUK9NFTd6TAWBCEegoyZQghCUcKzDvQvtM4pcI6LnKW1lVm+pP0C0L
Sxb7b1zhodKH4AUGQtpnDvMv4DGD1C+AKzGRD5aAF6hjzHFcT2kKqFg1esTfd+9moE1CC3rCy9n2
A4goJ5cErpoG8iIGi5b16oZk/GS1SbwZTTgtLF6JHjYgleWAa9f+1r7845qLvzHqueaiBvQdwy8+
O2Oux/09E/Ni5nFt4zP93U2WlHiHUH6OS2nAfoRdby+zj8e39TIqQ5nhx2+49ffaFwmYWn/kgu8W
NfROMnCgqQj3Xn9MLvWMqPxiPNJxLop9jtX0VvkwAErxDdet35Qc8Ni6BFbUYx21qdhEzvvXOEc2
VQ5ogWCocJsi19v/BnmJ7yMdKW05ycfQBfdwm1VXeVpTXenTR/Q45EFlfUpTdGNm7eV6DKKB9x+d
TaAACgW2eMfa1iH21t2pNm2GYT/9nRCcHbx62ctni6FsgbyyYAoGX0EGZW7H5PkdO7FDyavnNN1G
4/eWrQN00D+jwReUhCtQsnfjrPlIBQtPptIaUgXWbmYVpmvJcwaEzW4onV5m2bQAxbO7hiO7/Owc
yOluwk6lMO+EZC/+dnmhRpK3e67rAB96f6OqkFQgMjgmZBR5bDYKp3UbTM0UgDJ2W4ZzoOPJTHuO
CZxPalZl0me74IP3e7/Cr9h6Zm24+G0xgyloW5acfvms1Qyu9SlYmhIt3rYVRffD6K5RQJScI6OK
nqkW5uIwj3r/gCXwAa35edbaL0frVs96X0y2TVenKGjYO/fHLumDc1NH4iZ1PFPKByG3/2I4Fxfy
+Ey2sW2UNbqOoLa7W1wghlcHYKEBdvaGedsIdK9cTfVw55HM7oAe8mL7b188UXv8NDGrAExpkhku
aQPZ9lVC7NmVbZ0f3KCbBAwt9m3hUl23pJVNMUja9h0CM1WS38TaEP9CbXkDNmKjmpHYY+mAEqdz
pYxFc+Rysm8yiAbot9N0VdyJCLS3cIURNotLY8pJLdwt7ApAeTliG2wNYeBunI4JBdBM4FbyH90/
0TMPwUqRjAQK1G2aYOXj/jViTmul+hhMbMm5kvD7wNtuZA5h3dtVXoN3cV1h17aLuGbEbhrOiQYH
u6ZGX3d7fLnBptIuK2PTyf7EY5gJbvAvDxygpXZlsYYW2xqV2kXSxrO9VxWimXjPPtDNFuCbtY8a
Amx316l9QEHVYHuVAmsCGB5iZAwCb97NBWHghZiM3WNHvrDKaBWu4FRwrvxpKUOCSfhmpzsWfOEb
fTf8yxPwQKdh89PRikq3EMCNCpyb2AwKf5tkX0PQZt2vvIivK5jPnRBlkCHsvpCEQLjd9ffpgZOC
F9jEPwZb53Q7W1hTqb1i/IOp21eld8Nr4dokKWqo2Z9vlMAx+EnTl7Gb4RAFcfc9oOYwBhpcpNfT
9nQw++BeYQvdMb/hQ3jiM6N+fnUCJgAMLIS1/SSzALO5NOQqxytF/ow7oN3il1ZYqFUsXbYDRRPg
wZyzpgv0aItRmn5dFjFWPjl7zjevtPCAbNKAcGXdXm39vdS4bp2GJzoq3vk2W0Ax1eN2zjs1PeN+
quH8YLQa9A2VX0xVUGEeLF/quWjvtBwK5jDMKMVvqFFSjw/7vfm0Lj8+kpy+M4ZYhvQPO8nrO+06
cqVCcOW37Q7tPwwV9jqJkZtRbhVYVXjqwt28bRasqm/vCaz2oGFOhtbvH47PyuJ6+LHXQFMW5AcE
OBEWn033zmiVqXwNyixDKi0BFqKoktFizbrbIf/fjo7iAwXA2SVi3abLYmBYLK4DcCeTiXSpOwHQ
ZudyZcTFJKOGkuksQCrCMIVwU8xJZfYWUggRmCp0p+qmYbRFrX9Hb0J1apPQsOAN8F6y7B49wWdL
r6JHsaWXgjiGdRcRJZEuOhKvIHS8WiDM4cumPFuvRgxw3Aco3venpFwi+1JeN+ps1v6hZlAKmSWr
MVMYETPv06G+d3HsnuyQN5fri/2oeR2ZoxVzYV4SJNTN/vj3is72+AzEDOm/8wflPI0/BMbcZ7D8
GxNLwMDh88ZCuZ3vkc9uECIY6G2FNfAFuMWVWgCZeEqYbSmnei4pOyCHI8ddGP030d+HahQGgCu7
MiXQU8SFOYgglhr5m96BblgTxjf2Dojwc+cEzun5VBPZUFfUqH0FRMTzVZ+rWkkjOtrjG15DmJSB
Kr3BJNTnYQbClYI56UDGUf7YroHYYW+FLR1/KmAyLGdkZMeB/BQynrzH+TAnYdUL3XzzcmaJDH95
RqwkExkwtWcV3TntlhMlKM7MHH+hL+zO/fMdO8gzf9k8nn8iQVwcaLBgzNPwdcHDqSnjojTPprSp
1+4n1FjH+J0EmRFsBf1VSKHWHKcqmuVjqTbZEGGqwTMb+d4lwf+nEMhV/5657FjP/uqz5oENMh2o
GwAj59iSHDxEEov1liu4dMCKS5Tfr4Onqniw3F4amq9DZUx/u+VOXOoYz+qp3sSyr3B8IMGAOl3/
CB+hlBPwrD2OqoTsuVeuiZbGnXHnYF46dvg7XfQho5MaZ0jVFnrE0AxHcXS+dCbdifc5jcfP9uiT
NQSP4EaYqmlF0/TJ+gXr/G7zpX6TgSlkYK70Qz5AXzI+Dv+texd8QImymG9FzwsHCZos0AJHKYQH
7QLjHnsV5D6uJ0VFVZg+/9F935+HY7FtVA+qXmLIIOaoz9L24wswKt/DM95jEUwkmOvS5vLgB3ey
BX8wfGXDaIXVlx4cxGmI73snAg62JI4AIxfwvl5o9aJeLkvgPsbQLbjDO+cjG1wnmtSUWWA6FLyY
LqrVYr8wf9mCZiW0CzW/GDGcksjwZ0gSB9llBGwj2L0A1YR/P+FTAw9pLyJwhuUYtyJ4BY4fRGju
8en/zdKtChtSZo4+cmk/dqP+fBIyWp6AESNQ2cGhiMU8ZCAn1fzROJ2Cn71wLIyLqo/rr+NfmPRX
kWYkuZdrporvA7TV2cnCBJ7bgPVfRLMn00ECgaIJKCOG59K9GMeLO5VPdRZ5sXu26CvsdpMIq/u6
YMTQCiDBwW2EgTXbOxGyROz78fl9ugDiJnHrb9V5oknbaGAiThJuscEzSO6G1Tjp2FVgc+wY3vf2
9xH/q7o9C9kLEdQVD8i1lSjqBqqkCU+vuuzC3ZcUOvfF7qyilgg9hexs4DDH8zDg5LH7PI5oylG3
7XzX1Peovm3AErkoNvC11cCGAsr2P5R+7KmdMPJS6+0xLPR9GFZ7P7CkMN79JkWeOgPa4UxgZ2Yw
DNZZPrH2MhUUWx2pEiHybtVSOUvv43cqodj5UBQ7UQA1GHCgdRno+qPjMkAVEhZbmR3dmYIISLou
DMNe8yHm5mKHCmrcfor/3T8jNJHKV83AyuuEUICnfQmThP1EqdawO5lcE5RvaV/KZxtT1uOMcrOm
EiWUOj4SXYDJpHK1iPkZtyYP6XhEW/na9aC/ElPRjJqExLZ5JilVoJCkcw+Ywc26u3biGf4v0JDZ
7TdW/Kjy3gnwWSbr/TGJze/2XEdNoTg6HxB+JbwldVJwk+kUWdW/HR7jbxFFM3bYazaXFY19gqXV
OL+uYOQFXOCzdIQTWHFQS53OnPmWdIC1ruwYYA0CYqV1do9THjYkid15s4hibr+62fNw4C2KrgHG
6OIw1vLpW8AysqbxTlKUxny4HmRd7HjWPkbXs61NPzbUZpXa7nk2pImFwbFVd9fLKPqAdBg/0kIa
Az78OZM9LDmC2yGq+Msk+QmSemf46IjnhesXuI71vkfncN+MXcjv6dzuu4ePxpVB9QNxaKJe9ydI
XjSGGowSpmPxwYIpBESp6gsD4+VpvF6lQrTY28pNYWb2xQ/scDybpx2Qsb0ndLZ+A2FwJ8PW0P2v
2Sibo+ivmWtrSEtQnMxVKPCbl5qNql7A6ci4ZUDfKdL7JAgENVr11RzXjil71pnWqbaCzsaJr+1b
xw04ki+T4RCFylxf0WUnKEwCSysb/fmKvvzvQa4Sa/NR2mmK0+2tEruUX+6STAUp0Zutj3eDj9I2
DazXPr7YD+rUxbEmYhHwaQyd4amLUJUDRRNKQ4/jx8UNQSbssxgEpib87hjcgTwBLLG2rxDoozG9
KFdA/dBw+WZuctacPu7mkx+r2TLLk3GhdwDUEqW19RdfrHYTNnzswJIrECCJYMpfgyQMxL7u3b/h
4Xdkwfj92VDnPCO7ZqvdeABE32u+8iT8e69KEYmXWrJnBxH/ILI7aUKB6RhvdcY6tFPDfck66lXc
ZK+YJIiyMDeebo5wD81AryzS+h9Ml5roLFH+cRiICiSOzb63d6PW7gwcjfB1UKNXt7vJd9DaV2fU
HD495P+qJcUoerOiNtzzpuck7Lqe4sJlf8lX0EZ2ZE0p6jHASNobMADm2VH2yUy4KK47kRWjHutK
BvKFS8VbTgqmPXyqgqhT2s+655aQb3yvZ+PeD+WxKqfuZmOD9vjHVI6SWIV9jrzo/5zdlMV6WRTB
tajnIRcbixhurWUgeHLCjsDv6C/nLNlXDGLptJFaMWlT4MunhlhDoIt08kkkA8Q+YDBhEQM6/aIA
uB9t8sq+8sylO2arklzVd74dM6LFV33w3LP/xcd9NWQZ2r001akuKFC5HXCRa6D18MSqvzkYcbJq
FEdxRAWjBGG/hLuD2t8sx4lS/NDWL6xZWJpkyYs13NPKwt2R/SUGXA439GTdm+KERBef8TgUIcr4
ocL3YddD5/f2H+IbboIovtLFPaQifgvgIDQHggLmx3aYsULH0DuYwXZFSwM99qvUJARXDy4wIkzf
Xrimt+pkfJ/bGvv80VhgpsVbyETyQ9uBrChpt2X6VjQUxg/CQ91ivIwUv2uPYpdJXm1FCTXJDMdr
ypDcFfYjk5V/hH+o/831V7N4e9GF6QcFRqc6rDlhQyfilgVgATIXVttk0YBHkopljfZOdDWsIU2o
mZ1ROp4Nz2BqI11mFL9/9wTlewFPtCn3ZzBaUZS11Fx8+aaMa1EMJVM/riFXnPzH6JoCpP27n7tx
WdFbrfMtvi1no/h+aaukxgFZiG6UxFEs+ydAM8wICqajmEXXJDXOvIRhZNxgfCJoetngDusmJMMK
l3RyfNzAuQ+ugakA28btOX1rDdwdejhe7DCq8Bwjy3/RmMmFeqtjVMi6WaULi8b+SHzsiUIjCKjC
iv4tZxp/+hb5F08OwTIftcURsOLOoIfc7efwRyUuLLFtR8QjUZkLuX2PbRJj2Dh7/2WRf9CN3sCC
DxUnoNXBmo6SkWj82hB8ZN4ocLVarvPaAX4476XQU9/R47KJ2FBHSS23I0e9feV6RKWMvezMrK4a
IwohuhqpwqiaaTBSLJctvHTLY9+cRELxvrjgAtDPoC3VozdUsM+aMVcCXEHmd8OHkjaRiPfefaVa
rVihO5xIxQT8MU0LRf+Jd1S1BQBxUBf8dlhBKB9xkx1L4DAjUFzSCI9GCjkFlDRlrPt3+CtgeHdt
j6rldGRBQTHGWlOggQlB+kyRIhYKqmwHmcmwrbwjeUfoh0U7cEKTl10oDIC/mctVpQCpGkTCxbY8
nGJF6vUNhyHmZd+6+pU5RgRvw5xz+93oGmzaksYap/wQfJsDxcC9FIQFiOqz9azJB+2bht2UmI9V
9cFZLa1URkmZ/zQElhztXSfSFh2QFwJC9dpQyrIUpJEZ2HRSWVVOJnatIHfZouEcrtnD/yhFHoWV
c4nknlu3/+YmMtZDqCkVjj4Zh4S5oCAy+P/P2wf/gU6FzKRXzKl3XaDw8GIMSEbsI6bwdtzP9rI2
QIBWAT0Cb1jIyizY3k/YnGw1sLz8iV79MMr0F99/N2vN8wJkZkNxTKPqzDSpvfvWneYyZ89EqC22
Jw8vs9uKV73FhtyJ1oHQ1DMoMN8eaXYpg2JtPU5v95F1llBj43QMj9dv4lovTG9EmkcPDXmLxDM7
ODeG/J2Jk7tB6POCUT1QyXVoKG+EDBH8R+swz/HbJnbT1jFXa7lfCcs5NXi8kn0Xv3cJUKelPQR9
obnBswJ3E1tY6Abzmxaq0a6kxtN7EO6PcElTGFN6TkkrA7Kah97Hf63jp7qXhwKRm0QzLX1gBxiv
Wns36rEkwJUVNjgBZH+75A/EjmiyyC3tvQDLeZ8dIoWN4gUZIxjx8En/YrIizH5Rrm3lixnG4gVe
6blWXvMEkBIig+7K8gMkOTh3xNv143EfvhUu45dMWg6ac9fYg4bCuupW3WCW+jOG+Cyn8A/zZz8p
LRAHKyB/OAk+n6f9wzzKyXLxGaITTHntMExSC/eqikkG3gDdL0usaoBKnzs/Ik4fYToqDy9sQEDu
0Cvmngq9c10Vek4ZJzViOrbUezJOm5FNg8GyMw093Vp4d2n8iBE+MbYcVJSQI5gAi4I2fjlMTLbt
71q7uA8/MsLBXWeHWhwCnakP4bB61+bBFoFiHyc6Sedsq5Vz0izar/L4myYSN63PyIXO6Dsyqx2Q
Y8F1hKK72P0zlTjDnzfHBnvdUevLbhPILKb+Qrn+2qFlEAlyy5fmgV/S52iijo1Vp/aSPGxdA0QP
0KLBcm62nntvEyIPJeMAmSzVvD5aCCKV+STucaXEmkUJS4tLdWsjfxGohSVmF2MIli0svo7iKZVS
LT2d5wuqSBcyoeK7ttxxpd0YqH4pGMFK5pudByozohoHb7SfDaWmCCzDeyDXn5qqoiN3a0+58tn/
seq4abh+s4a/v4Bx1pKMN39p4ZVgB1iYP1czEH1+0oV+HghV2e0ly3+uFouglvMX/qUQsAjJ4/kY
Z7VwPhRezHoKvdjvkrD8E96bSi3wDYQXlcLvIQEqN8B21QIT+iHpT8sER2EwjfdfE3iCi5TmK3wi
7sf4fIHVvqY4eiPqSbSCUgm64Z1OXOewiE9PMxhm+Gjq6RKAWLhWcuiTItgiqzsNIwJut9vZ+BoU
XlT2c1q9XA1af88OKKT4drtz/YwgfQVmLKYt/ajhKz9sMTpEQ+Nwnm31pYakDMWDmOqkjZ49yvFy
fpe7GUyD5zZzFV02/ymUc1cht6oU503Gb0hGLuv2kaeRFLb8qsFJk7+8T8aglyB/CWTQ3nYHx65h
UhzU9grP6H6FDyfIY6wXyqvZmTJoi9maAmsXoltA8D0IAu4ciy22hk8q/K9YDwL1NObJ6QgeWHw8
C1ziIySHtApXONtnsTa6/adRYNwZ9GG4CBzzUm+2Ys0wa5I0/MRIZPSHBYzng8Ky5zc7Q6sZ/lkP
FTdX2pGcbzu3aPzfm9RdJnSRSgncxLnU1hWUB9WUVGFRuyAivGghh7ZwdrZdNJVyxg7ZYjQC148N
QymjTmthM4Pevg0Ad2TncGlStoa19PzWTlpxHemQfkRYlK9nOjuv7SnetFY44ItGFtl+YsRA+Jb8
A0lmP/ZlOy+ieGRcBPLM2aRnnMSplA/nJ3pF0X6dN7oHmz/UQkZTIHXKW8hVmfqEHR4PYHutl+LC
NWGxaayXOVZ+n11/KU8FRGGtnV5gB3+jDun071Wkyrvhil2jiPewkQun7Mdvrjo7Zi5dfupxxpJm
Oe+1SOQtcq3A3wVr9exHcvUUQxYU7f9JWs1kUJAz8H2r04a87pP+zLKGxlRTWEkq0mOb5uVY5K5+
5ZWfeRCfRyvBSWgSO+vO71hHwBrayIt5L06VXu3W9gyz6dWkPXZn1iPfxrdnWLixj4HGZVWYumct
MXA+PscqlPKASYzlWN1AW6mzafZxNxU4Z2DA0mVgS9B4XW+Vd256nWFyeulGacKejFF67MwMaoAN
bbID7dNBVY/OszRg2ebMe/Dk6SoIOQVRL2s+W+iIxm7qG0hz4drtpv3jdZtbHSBmW0IpIMktrQMq
Ynn6dZ4HUbjJvAmuSuh/ZvbqCJgQIWKNKLQ4awb5r/q80ytckyot3HF0uVAmpM3qTMMMs0SjtA8k
k5D3A8ci7cG0r9xF1O3kgOpg6xl50ogi0KisgjqeDSCEjTsOrctwsxflAjnn3/pBBKLK959Hh8Ts
3+eXdBMOvdO6trCvK+AwRQYg8fB1XOIhJf2iqTsMHuR4bAabOPw+yGGEUN2MumjsFmuY3Gu2kVma
eQeq/Us160L4/gRxbienaq8YU2qnUgP7jJmMgu5Xc3zEUaggeVRpgUNow/+aSJJrmNiln+UkiGKM
JJUD36GLM7ZR0McObb8Ncjltlqj131AR6mUQBPV4yTgymx/+7A7JLUJwFLtLHPYkqRozT6iCmugd
RMl+vBVP8idb3Fv/jZeB3Z325lLME5RMq9T49uVKiu7G08n+5GOd1RVDWEVO6mV/Lb87zVeGCe02
E/HbFFzbKDTxq5I7VhHSqjmkMluftppKU5c0lox2syeZ0m4r3ohO3Wjcr22Fwp+rxgZPtUKlMw+S
8xqO29wJPBaGGhZs/5NOdmMPHAbYxY+1GF1yc/eZDPyu7PhTD6Hcsc2LC7WasODgot8OQJ154EgU
zp1gprJ+nIStcMR+od5iWrEm/Aqjt0Y5muAIdjEbsJJuFwuDQ+Cw1OBcYGEkZgTMm0DDxYxXNvoA
CL/8VOehTtd1gXiyBnqA/EW8D/lr+9dU4W9cws0yvy78+d1GsTdCilsRzZxdeADYqDW/LpralA9C
EQLQTeyQrUdIyRaJiUrRqueZz042WS8FVgxPJpgAfl7SALBqqzlpCHMN7s6FlcPmdRw3b73F7ePK
uY0Uv5MLb22656TQPdM3rMx9ccteoQQrxXp/6rUal5cBJ06f0WaFRVrCAlBxPwuReauhwqcxaMFp
smk9SBt0tI5s2MoRD7b/4V42M/tmaGo+oOM5XUWcVwRzCRXQTWHywv8x5K/m1WdkfASdsKRgD9he
2p8F1/mXvDctnqU2ry4jaoWY34dLoECtnNslltSdOQVLsC2NLGeXpS3uk7hSkoKDY8TmVu94EYaL
ME+6XBGDAS7JvzoLuHibl/J9fLA3709gX9GMdIrkXGYRp5n+SsrZ3rtxzuSWwSKZlhwAVNPc1/cZ
2mRuqDv8xVFBZphwc23Z8hYOrMp7J88fZY+/tycy2OnWB5SxR6ZKN8gDwCjCkzeT/4dcqb2jeB3z
kNJB43qrR++xWvxugubF6yC0oVchIcRE+hh7pI+B/0PdpUNg6SEK4cgGTE9xvi1iDnN1VwjVZaNB
9IGaR0omYMx4ZGki1n2cC+KpbR0EV2ObgTlw5dqEImZWJuSQ+1tN/rQS7KP/wA/SEHBCzCDn0V9d
RYT7yRzhNYVM+A0nKxKFK1rR/PsiMPgnd2GyIjProdYCDfI+w5WSdwG/8DDbDxb6vd2h1/Y0KRw/
eQD8u9gzIZyhFlePSzksa7EYYqtA56h1uaClLdY3PPZ8/zXd6Hg8jzltoj94/xeUIgK4sNBpI6Vd
KzLXXh6IPcDkBQI0evaIRWRHimmjJurkhlqlibZAS7a9+K0r7tP45RRHY8vZdn+OYsPiEMt8cIVQ
hvBTVPV9HAScvS8tciaRQfjPVa2I0fHJ0mo3/QlJOXpkM/L8ZQC2PPxrnMR99yZkQ1+3jCC1BKc3
rrsgTurY6gJq9aHgJFPQQIE/t0x0KUKc+WU5IgoN0gYvn3Xs/hOOOn4HbIsKhxoKt7gBwC+oBkt1
UEr1WqrIs4zo9EgkLUt0OeIu628o2aMlvP8ZHCBw2EcHomnoPfa3W6pRh+JpulB/PlHHTKSlAwaf
EKzOqiS0teG6fQWXMv7wzTljdQfNfATsUSjTKr4DgbqGAPzmyKaBx2IrA3siI1mj6e0JK6p6onHv
bFE0OopbBQ9dAXG+4sGkPrg1z28OshiAb1ZhM6492CZUksa7jmOK1ATijIQMyMxOswmM8PlBzJic
WOQaFk/NQr7+XaPdMpBkpFo6ijr1uwGe9jutNHY5Z9de6BfhUoCo0LlK/OtFrD60/6v76nlwGhPS
j7vtiw28fwr/i+WfziXC/o0+DJn20eGFOawDA3qsKPyzlQYk+Gg6TzaVLmcPTEXuHfA3cXWo44TL
VODvkQHVpWNqKj6ONxOf9GMDqlidwE+zMINpxZK36cLfuhv0zfAwiWJ+/EbDHv64gnaT06pAQTpW
p+GIlnBOWqvZHnJT+C0q49Hev4UpckUj1h7BG5jnja1MRimRMtoM9qX4d5MNmzB6mGlOD4v7ElFU
CqMFIAiBVmGQIY8Ih4vyryVdOgJB+wFFw0wk9/16Sv6VVqQgUcENE6dviv7Rc/S6Sbx5sTbpmFZc
8GcdQ3WUsR7PksDwHmzjp0y897+5LGBeJvV/V08RHnP4BU/v6lc9ZZA+FuE1Vrk=
`protect end_protected
