`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
/s4smwdsOw1A9c2QWhMhhTiEaUri9DgzebkTsEGTJer5MOb8+3eUnNB0efSWURUnjnyT+uxSMVvh
MTjBNtAwEQv1fNL5BvgmoQOd2k3PNZ1OKztf5wW8nq/oyNY5P+QZX2hfPBlaB12o4XZM11xnX+if
jxmlrz5sKWn3tmjxAIbJA5rOjQ+5cDKQJYhSh5CsVJ72WseXjklNY3JEpnqIleoqHwn15lwKhqjn
U5pchs1FR9OI/97nR9v3Gw/mZgzc5jifbxUb7f7+gtttxJP72Yo/kSDF0surie5XDdC2tzNW4uJh
Kzb1g7rTm20BKJxpM24WayfTVdHEhC0MXIhj1y2vO2PhIhqBU2TrYkwCMTcVPYkeFY2pXSnsCSo2
fGD41wI0jPIzH8rh+3cQviEuJTXMWKffLj9fE0+nOQxL3v7uUNk7XDr8iAlygMtAc5wpZyEuSljJ
nq8LLACZOAI2iQkByJ2EgyjuG66K5bmEbEmKzVE5vC6YeDhGfvi/tsEA4K7D4+2gkQFFgKK2EENP
CQl2gheiiQG7GlipD0/N8zceNYF7vOTfkE4BbwLgJFF5AWRbLDcYEH+C0fCtOH7USX5d58ypVPnx
yvuTv28mr7uhP5JqoAg+ZMBUt17gzz1evoBA4ij/jRBMV+ngfiP7CRejzOzOmUIxpa+chdmfIGei
jde0A/FpI3QiMokT0oh/aHKVeZVuBIE3GLS/Bw1Sm29Op5n7WxiLvFvU0THGZBQlGvOxz6WxHh9W
DyqNL6ahgNlLmpl5lDMsK26SX6NCPz6bK+BQIP2JAiobRNFD4fPolHHP0C1O5lFFllFiI4RZSjCG
lxUr0dVOBNw66LwZFi0XuHOXK06IE/+LZkx+V62r+AVuKkXPNVc8V25sheNchcGR+5+ocx4qnmIH
8GaiS3+L0Ba9xnKTU5EMKqcecJm/QCvA/IZClqSMaA4MXN3he8tD7wI5Oit8clmcnhCzvS6FN8gN
bBDEzkwdUrTF9hTIZ8j8BvH3sIqKAPwBp4lnXq9+lXeiZorA3LLSMd1M1oj8tK8pJ8bVjhWxp9n7
EGbwUgGRhAGveANx4f/U9lArgfPNkDM3eWbXim6plgSAN9FoufZJZZYL81kriuKNb7yREu/Jf4SY
nF76aBl3Q4MwPYo5sQrszi2PHNxid84Ndf882/JQQVkx0Z23nijs5Kn6ld9ZLQfy3khLx0zjnVQO
9QAx98MmQeQssFtIIArKnA==
`protect end_protected
