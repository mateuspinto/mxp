XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���BȻ�M]{�!��d����.u���eg���rn������d�������U�t`�;����WB�
�%|�A��ua)#�O������i�5�\�š��W���!��E+G��'{�/��x�M&��}S�.����u�|�@c���qW�'�I��u,�N)/����`y�/�n2��O-�:��}ܣ���Ҫ��Ǉ�:Ra��ڥȸ#2�S!z#�2�w+��*�P�m"��P�J E���C����>3�8M�J����"���a���N���$�15WS�R��n��Ȑ�"�,�6U]ɫ_�D#V9b���lxkEn^�QU:�^����4J���CZ�Z@��˖�y1ˡ�X��&�W�i�%1w�-��=�{������7� �m��csN�,��3�G��G�;UA@��>l�>gJ�u��)]tm�n������.,H�3I1����a;P�|X�к�N��w�������u��ɝD<�̾��a�s4ɷLyq8��25f������0q
�q�E�s\V��Sm��	 u*�q�b��9>�j����Ui��h�3\��3��?eBޛ�*�q�z#��Bή�B��~��*k�QR��i:",��8GQ����<�q	Si��n�%ɶ����JMsG�����q1B���j�jkȡ��]]�M�~Dk?%��=���u�a"����W��͋7��,�y�͡L6��p�����f"���ۨ e+2���ĩ[j�U�3�w?N�4LWQa����-XlxVHYEB     400     190��w����5�4��G�p���\�7�Ӛ�{ɤdD��J�Q�F��A�*)F���4{����"Y�c4;���߆�U�;�50ʦ������$�P�hz�`i�rj�k���%K���me��b�m�wM�H�q8W�^��]Eu�ʡ��l�q���B
DrϺ�b�d�E�A8��.d�,}��s�OH-Ȫ���h\
��Z[܏vu��m��A����Ypf˾��C߅{u�k7�j+yKy1x1�\��'
a���lDI��=�|��A������8����+�lX���\-���C�ܒ�1����q�f��T���f;Ŭ��C�!�ýω$�eV�F�^q�%��g@�˲{�d��$(�\�u�m�%c�qO���zh�Z|���2�� ���4�z)����3��TXlxVHYEB     400     1a0�ǈ�Du�LA/�R#r
/�}����;���3&9t����cV�^���E�ړ�k��h[`3����?|c�
MSr��k�r,�r�;����M%��%���D|���� :��s�}p��h�[y�~�2xt�5�?=�.��?���3'�z��ߵ�#��㠨�%6,ݐ_�� D�Д3�կ�d�*wO����5́�x+���� ���<n*��0w��J ���P�<��!�����'hh���־�>.F�}Z/�X����o(��_/N���@-H�ɋM="������u�|��a
*~q��P�K$|?���Y�/+G��[挕��xs�$�Ȫ��ƥ�8!9NiT �1ɩ���T��OB(���gR��@�R���X�Z&2�(T��������x����#XlxVHYEB     400     1301؀�2�B8�m�y�`uF`"�-��Iy?��*��k̳H�8\%l	��]���G=U������{1)̧�|�B�k��.��x�+��,u �E��A��W�t}��e}���p�Ӱ����?�-��Ժ����BF���WG��~�@���,�O�ՙ�
�����J��2�L D"�������κ�휭�."�<�n}��*{}H��v��R88�H��CAysN�0a`-��4s���]/�ak�F~ 4��g���2Z�1e8��!.�>��u�R�; l2:���;���䅚�TZ�,*�%l\�XlxVHYEB     400     160^����z�Sa?���F��y��k'�Z�'�U	�K!)��&vߓ�4����;i����}��x���2W= �9Y�Ik���:�{m6���Fs��x�8EXw��P�h�O��{�vN	u��Er��b��ĉ�"Q������/�F;D)�#'�]��q{��'�#�)��A���{�i�PT�N�PZ~ϡ�s�"�a���A�����6v�
:1K�RPX,U����[�����L	�����6�xoG���*	?Q�6T���Ң +�?x����*����A0c�*߹{�����Mc/�H�����e
x/��OύAPS�#�8!�+�\mXXlxVHYEB      3a      40��?s��(�``͞����~�?���^���kFm���R�#5�MA2J�Td_��t�R��/�C���