XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t2	�<������vO�$���@$������H�d�0H_�+��J'l���	��Ȗ*X�}9�	<$�uF�'���4[h9 à��y�ɷy�^f��8�BOlNR��0�z-c�Y�&R1-�tѝ.��F�L0�#�C�ec�{ľ~�G��bi����b��i A�%�p�vMg�"�cB���N!�ص?�bپ	N�7��"�L�7=�O�	��v���)1C�Y{�uRY�g�.A�R�4m���+�W�ъ�ˊ�Vy�3�Q=�sޜ�G`��Ӧ�j�Mk�Q�ڎ��Z6{c5�x�e�I���	�+v� ���y��-0������e�&w��h{�I���8/-Y��}�7�B��Ae*�������@�1U a4\.Y���E�A�:Ȃ((/*�2��Kw6���7R�i��D�:���Ӟ����s�f];�7!�)�T�(�.���Ň�v��IЭ��CN^�����	Z0a�N+�r��9i���$:���o���EM9ď'��7���Nj�9	��0��`�\|1'`
�����c?+ߠ��'�"2sa[��(����6Jz�cڍ�UU��|!��2�I�#v���6x�<�o�D��P�E��L��߱�A՜#/�]HK�of�G.��#
�ɐ�
�+�:�;�lB�Lk��g��[N&�n��g��C�Oֵ:���`��I_�'���{؂�x�����j#���c�je�@YL�s���U��B9#�m��NhE��L�U�� ��<z�c���aEM�g�&��
����XlxVHYEB     400     180��fCtsy��ױG�D�� ���|Z|6�؆x��i�N��~&�)6�v[ɕ�(�	�C�����v�s�CQK�EH��'����<n�L|}�o�֫��.ѧ�Q{�מ	����fh�2�r=�Fj�>;�8��O��K��ߺ�Yt�;���|�ۓ�v6��E��\�@�i�����!^�����|v$�u�U/����fJ��&z��!ܮ�d��)�=a��sn�L�*9�/��+��P�N��C�Ry&�,�?X|�y���r���4��v�>,9n�m�܃֞��bE��,:JXG����>��|�*��b��7T3����Nc�ђ�Ѯ�D�����4�,c�_��\����ע���"��~��v���XlxVHYEB     400     1801���|�L��{Vs�kq����dY����Ǵ�����X0���Yf{n��hd�~~��,r�c���C�@)�Hn ���X������{cBIzhn�<l�*� Rd���I����7�dF�^P�b3 ��@k��c�H�E�y9��a<$V�j��b����m����YUlqBj�g��l����|�k+!���n�P+#	��Uth�qx_o�G=*l�����(u�b����G>P� �[����J`xK�(��Z1i���9�&�M�Tl7��UxX}7k�B	u��L�I=�:��'�T%X������һ,Tp�c��x�,W��8��{Vr?�8�΍r�ڊ7�N��Nm.�)�\l���R��U8,,���U ����>/�?mkXlxVHYEB     400     170��"�����|����hV�s�ZFjy�Z��oe^��jk؟�KZ(�N3�Q��;`��6dp]4k�sX/B��OC�`��o��sCf� r*:��|�p��]�?�UE� � ���
R��ިǤ12L��F���9ڿ�j��Ns����Y�ǪD�L 9�w��"S1,N N���ت��W@5��{>�A�d��}~�5�9� W&��`��`j��9ӏ	���hFT���"�G�"k�N�]t���b2��� &�:8;<��)���ۖ"�����`�����	#eE-d�����kK��ƷJ�A��+���N��^�x���ˉK+�� ߑ���;9Kt�:�Xs{�T��Е��XlxVHYEB     2e8     120[�f�4G�sY�/h�"K��7n0�!�9�@ G�	NA��$2��G+�-�щQ7���Q������*��i�)�@�M��C�J�9lB�^��rl��O�g�������ɤ�Ύ��fq�3�ż��k!e"'!�����3�Vs��3��`�w�Ƿ?�)blV�	�؁r�	T�+����I�:�Y9%#��%�gU�Uk�����'���j�� ���s�Ю�L;a��vN:Bb�0Jƙ�\�YjE`�|���U��͆z�!��A�a�*k&R��������b��%�