`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
qoEz1cIEaVnI9afJ4bcwjlodk3JilWZy8YBEI57ZFf3NqSM2qeBemnCIEaAoAKgOXO4ER5HYefOt
x5m25AqcHvEO5m/OWUREihNszhBYSLrHxdY/HGIhMPgOasOU1wJEoHycOzyOPsKFhhBQ4eLVXW8G
/ZfM2aN2G4pRCpH8I1VC5NanXM9ok4K+QJuL5+uPXdJi3XumRak9O0Ivoy/OkM3/JMtgka+xrV2L
fzqSGccbBlPA39pSbzi0bYF9+TzNWnNePfY9eyRF+NFbvoVOnDJhpe5+t+8Qh/wWh5wkE095oiTd
3LdwrKGa+292xpNb8DEA9deVGRS9dXlwvn8p7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="q3mjuMWV/Pu9HvAmeAjh0pj0rdhoxfshUnVjXN1aNOQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49760)
`protect data_block
Co2ZhFWXwwuCcYp7Gv7ynkG+cg9BAJ2OOv34V3OaHkWIYL/6AokATGNoBsHgBqevILmOUchAMpZN
M/IBByKCbjfnvlPqH1Iry+67p+NGV3bs72pjFJFgX/I2SdYiC/00nWjNfWtcDwoYY2hoUqFodILP
dzsql3csG2tgqfZqbggh22lNpVjcwKBSzMMgA1j+aGwQlSTUyxtafRCt8/euFcGSNsLToWTYMye+
f9y+6Af48lO1D/hvIGLc84Nyqr92Ss141HlaMLTinN2vPc6RHc6xjDU8noBwt8bihqHvNd7lFIfn
RogJrDQmcRhMs6hTsUNjFBd9xY46yxc+NnYANf/8JOJYYofJKjHLgbmSsQRxK2k5hbqpyzGO1nCH
GwG1oi5W2h3e5VWJEK9MARhuhKmIvYeD+RFbphqjwWcoJ/djfmC28ZuxP7od4RO3HapSV/H5o+Rr
0UVpDzWj+ANs7U0qlpfOshr0YAA8e2wncEIrTlOPhmhBLCH88l28t9hMGsEIuaPmnmetauLmqNFV
m9/YTjjqDAwih6e5Lc/HWZVFedjhuI3QYeiyIBjR3DRFNgLTzKg2ewqzOiW4jbirrGfVLStzlV51
1YgE3s23CN28FHiurmkY7eMSFa6ks1Ynaz5DVaMI1fC55H0PY4XMG1Pgpv+6Y+WRutcRg/P1NvEw
R/4XLqqz278kxD6oTX5Xyt3EKvo60zAk4zPfFPJfGNbQesHLaGTPIGT9HYiOpcVoaFuOINGOIKV2
WcBA/vgfZH31oIEUrucIfZDYQHlq4w4WMwE9GaeRXDWwmV9oY4MCfYM26vxAYRW25zZuDQIOEsLQ
tvbWiYuiYc4d4+r9YZmszaEU7FIclEFMgDe2M7fEwzT/05e4G7CYUESNEpoaISVU50SqBY/F58et
5efh9wJZWWvh/6rGJX4kVodQ4KLNl78gmODLvICY2daWeH2l7EMriZiTqySwNl96A9qsv77DeKBm
Z8s6haGsUn9kmUgC2Gk//4o8MlzysPRe59iC7zq9yVvU2omOCYr7N/VYpzZJmuQlQoAWfty3BLfc
i4+gcdsFXbO9SiKRF1fXZloD537IYX5SonAnN+0D5Rj9ip3+5KxnkN5eDL5hyYmk4IzvS3ti8/Ei
+TxVN66EXcyZ19Cw04xP0sMQM+s2K1g6FD/TRvZZOjwb6VUKSkFmTuBJ3T0Mx2Xj3WFDeXkLBojs
ulDDneYN7msm6whOAK+okXIJlUrh8WgC4+HFRJ+0KOAy66atuzdklksS3J7e3dxot0L4Dl4gcgAg
cx/0IFNzoC/tjoX3PWi+FyCFBjYDMktx5PzhkYnz8/051g44uvw0QLhw/mx8GIsbiV9SGnVckWuC
wChEBuo8u9wRmSz/VXzHhdMRmIV98E0Bip2DRa/71VqDux/qkMK6aE7ha5fgakeVsvZUoic9i+Qo
iOBv7W8OaRaqxFib3H1nXjdjBn6kXJfGJEJWnLNZ2P9n5K0nPRP1r7s75C9dPCKth42y2ozqQtSi
b069nLSzVsARh78M6wbY9PtJ8p0lig/AZFwjfgYIjuUC0vxG5LMYUYYIQpDPzJa+7kluEEefTsll
6D+f0myiE71eKInLB4kTU1MDnAaXxyzvuAjqgUBzo7Da1Uueyez8LB0s8hnTsl10UKm2bRCx5b6C
L3w/bp4x0WRlFRErCIknl9wCGNuniz6n1UbeDjaKRTFeq5OKu0Yqf6hdxI32SVVHaYbveqUyhFVc
ZL7hZaRH3iJtBhmCBVCWdvm+Pod13EVbyyWBZjT9HwQTh6pJzB9ZYu1R63nidR5OG4GR+pSXluVf
3f59oJ4iIRKnswCnqN6vaPVXzf6MOxO6hQdbUH1lA3BtcYAxLNUDpKitXTRXp7gybi3EBxdQz4zz
6nlwPGcdXYR0AqGZY1zJkWF/EUXsngTrrZvI+s7UrYcYTZFquJsX34Osv7Hlgd+OLAtlfN96qh7E
8FdnglT6bekOqcE2VneI2Mw9nks8n4O+dqfjK/IyF5T+QlVpHwQoxLDC/iiHGytfgmeQVg9rR9JT
LwXu8CuG0tFpG9UMd/nkiYdY+hKUDaxy82349H1y1OC1fd+KLFiE1njoOy7hK4jT+k9XGVkMUvCQ
ofHeQkkGE/Jf6Qa6KSVxgaf9ohcMQ5wFKOhrNVyJUYaNjT2w66MT50lugXAInE6cCxzg/xfUTJYj
HL22HH6NWtM9zg3jBxgX6Vc8fEpYpAnNzAiptorldV72gzPElQLasllK37eMShHjbCAQNoBXlUtS
B2gNvuDjZVqBmHIM+gU4RukibDHQjWXI2S1ZRqK4SazQonAmJnaB0T4rOgGG/qZ77Q4S1sp0XuI0
GFtNKbDoToFU9+dfdiS7yjoJcvBOFjO84El/tRuFp7NeZZzcrfmbILq0vRT2OqkLyvLk8f0DERdY
9030n/OsP7jVJ89dHz7OUmdV2a+B4xB4zRPYr8VbiziJSJDRReqO0k6+UPQZl9SLeoqvefTMYqi2
Amclg9MGmwK0RkZVZsSb+muVa6bYSqEsO4/2ERAcIiyr3cVxdYwtoiKcyOtDYkaa5eOE3Syiptrl
7wy9rzedcD2lDu0Gqm1s9vNqT35Zk96vkxKaQk2YO+UNLHzAXyzGbDSotp1A0M2BHyiGxXYPC6Uo
SmWVU7M40kAu/1l4cXsncEu4rrEdMJBKM4XObtEzUJknlIo+9vN4GrpJNZyzCR1njE1S7OXWqWYd
516+FJIgTQbMfL+Y3/VSBAuF8uY7Os5moeZ7cAa12miV3sMmC5ai8rB8/WTVfIs35zfhp9nrAGl4
iRJhzHLFH+8WcISOsftqy+bDy5nc6kyb7VNjQs27NctQD1Ri8AG2JSGOMrOoDV+9hnYJ3VS4zhJ4
QSi/waDyHtvdI37QeP1DuvgEPkUme7ajL8eVEa5sQ57f2AZH3wAzwkpHmllm1XpQei6Oz2x/DnyA
hBMYelJNHKRhN2+ZDsF9tvO+J9lYqGxwh7MzdIizWRfR4+c0y2IEyT3vQHHLb0W/rOEmsgTcvKkQ
YFLop0rZSsp893bPsBnFEx00HjNImGPPDeiaxHS6UNa6YcYwkOEwNihYGmwUsGUgSupW7BVZc/AQ
Ga3yiKSiVV7nzotV4UnxnnzMBs/v384TZzAT7DsXyNg3AVSRfsnrvd7PAMEAB/BEPjShgbLNFPa+
P84wg0wv/JS7tkDVeTgWohgPuNH2vYjgcoMWaUhRirCEc9MVDzhcgfwGQd61SPfuqPEShv2h2WSS
WmjN26VcRMSlJb3qI1WBt/RyVCtX/FJYkvAUywhqY0X+Lx9jMEXUzpSYCUB0kK0YE5Y5qv3ckJpk
NRwB6NqUYf3xh1FZY6LasYsDyafcml3dbsnUol0TNLLjMz2NfJhcGXl3Tbe4thw9kM7mlFZZoTZ0
cLq4ErMJtNshqLcst5OKOV6f8H/5+siKlO7Afht4R9AonRstOKVWRm8OS/4popN5LJkq8DHw/mHQ
3Av/H38tQcT5SEzMUYU5bKy/eJPYPmbZ8k/tTmGJXZhr/hckmoMTp/lemkSpyyC9KqmtvbrhR+CZ
ZZkAIZy52JE/lkO3SwtcXcKcfnaa/GF1THRAcxof2Mg3E37yBZJjFnQLId/vAFvHAcx7dO3zXJ2z
AYEESTDotTdncn07QyGnNOYKmE8mpaZCKL3z0jnqd5E+A2xbydBC/owqKVu5ZotVl/6QthNm3VUe
5s3MQvJW/M0aCUDryE2MZtb9dpim7BBLY0K0uSGC0tZ5BMNNE2NAImppOiDplM36IyKeAOMt58r/
ehpLQ4uH56XXqaYd1l6pUhfZppgoS8bWhQPlP+afHKGtnPjrCYn7hqtWU1HhayBiAUZND+i74aTC
6A2U5cSSh4PUJ22rFmrhK5dAGNcSqukhFUFvrGrQiOgKxBrqUUrRUbaAYyf7Wgf+ROOnpOExecWi
Xxh+fVNVhtQL6Yn98gYGQTnuQkkur1RVwnGenFQZWqApsCW/p77E2De/0BSUsQnAmueMeNCAATPr
Twzu/IpA56lUxHsH4Ang/7NiePhcrcUN1KtzODDUC+WOXVOjpPfQchAwdqRnDSefysTET4Ija342
FF0Gl186iCFvY7BrJzEr1FSIV8WGtDr4PISUb3c3yjWiHn5rp92csAEnFMt/ncqDDcvbbr59y8wj
P5jEM2LX1ym44sMzk3MxP334xAJ4JvuUKiLmy32RjKvNs0ya4xUllu3dLwWiTw2pjDCVWIjxq1qX
/DDqnPBdz5TAzLqth95E6KnaLH6OQTQTuiSnQGQO+J2WaLxdWUiWUltVFjZgQcRajq5DLcR//c9a
PFOe1LZk4dpT1RE1aHv+CrPmccHaU+wYaijY2sPWNTBH1A2L3xnAlJZAI8FchifPfwDtXIS43koW
XzNqCheK7+DdJRfaFhkJhzKMUQ2tiLF7jsZm0W7lpnsPmi6r2mjXy7vUwsj0oSlfAnrsjfv7JpCa
WO0rFjEkNqjRCnpKUHeBE0uZM9dKZbiEa6U6XU8Ow1WD83RuumYoJSx88t/hDpx4L+dN8DDNMA/X
Seph1r1xyQju03aPJEBDAg7FkTLVA3r0pS1IYmPKt7KZNbKHr9yl7/5Fq4BgE6S+B15YEff6FLi1
A/mCEFteMnHFDyYIFQZxeSCQ66bssLEJRSqNBcO4LyxLYS1kRw+9wMVb6tZDl/Uq9rhOe7ufSgPi
dN29V+kqomKHfG5nxfBeXTR1nJLcixB7N0LqBzRpSozL78KNKBtpKLIGH6k4TBvEOQ0BDq7k8Lww
y4ZXWoonmk0t9DDB1ChOEpmYBVGiTfKg835c9E2FZTa01vopftY43dVFar4xAfYlqZyrBErwPuXA
hf9WyxEUCY74i25Rjq+kkXVdJ4SrIRpvcHXLda14zvAwNZUtDqvR3ZXvImuLMbnqIwr/PcDm8CL4
2fFrlG/OhzVHGWVsYmFvb7BRvl5I1muV4Zw1ToEt3cr72LpIi0LRCbfpvnYHEcdlnbS/T0WV48Mg
s+n9BN7z793tcU4/G5J9Y7IWXWdOYajmxLyvM40lVONuFnLN0XW5LyIyS3xDNJvzKDKnTZnksnl7
hGjkPI/ylbm+g2T3Nlp/9LWkRYdbBatI4bw/XudzECMLbvz5MAaGqxAGbpOIZ6sJY5emSL0ShD1q
skBrxgvDpCdw17GB5dALQCeQ8HoBS7Jeb/Rbtd03dsl3mfSuBYCMAm0htMdy4e4ohNh1fuP4cS7a
r81vVmqAwRCYb2S/Rvbs3+/WryvyrrZbehoRvRkze1Ml4btCXUBb3Zg8WswcdOODZkhDGboRH3qZ
1F7mFIJjMnnclGGEBVglG5cAtO4n04hqQpR+GjTnTSxgclBYvDxFYX/4de5ZnzQ6OabJlqB84dR/
6MAADlj0ly0KbKsWE9mx1kyHc3XO+z7DEDAYOYQGN2UEm+fBxo8QaSiC0/LT9HkXCWa1CdQ9I57n
SFBhEdpE2fJ3bmU90A5aWaSAdaPjHxXa+61sOzE95zJ+p/SpPq1tgGLPKv2vZdeSO5aSzk0CS7lW
+aRpaz0Yo/Nkxj5pi55VOsn+3/QyOiEc4MSmcOhdVXn04biXCqxCCiaSlZdhw3nrShOkR3+fjRtp
l8tpWmJRbbmWRbIN/HWJUQG3c8zno48HkV4RxFuLg5EIGqIDRLP09VEKiBHt5NT1Mgo+FiktFMzx
4cuzMA8vdWsccLSQvMrRs7TpYZzLRyq5doe2gzdISBJ5OGphUeyczUKUlosTlS+2Ek0ZomhAc6Rb
XqbL/Is6IcZUDkZWYwAhXAPIwoNIujNEvU0XIIEdSq11RNIWOsYx3nP+gzY/JRNCnh4+OrElXGmM
FzctwCCRfkir3hFERJdeSepox+LxOE730Qsk7Zt3+aUA3XujmejYR3S4yyuhRT4UFr9hPDgmdvTM
2bXLE46WK3jT4noLrIiOu3PIYy8N9BE5e9o6QPKRAA/0qXAVlUE73DwYX00kl2WZYiMDkeV/0ayI
Ai6+AnHBxuMtAhdFI0Eio/MslrobDY7Oj6bcDiegozszLCO9jU9CvyBDbbYupKvD/i8LFZsiC/S7
cbIYduGpP1TqhqTWrHOeRQ09VGXfO3ME5JGY4ZgoiA1Wx7f+4mRsHSLkbvln9YIzQzLgba6R+8za
Umn7M1hi2zIXXa7VRsPsoPWt3KZ3bpVXOthcYt12EoGIwbpiZNelwHgStg6udylPSLeVMZZo4Plc
Kn9znGp2+Dz0rxcbky8hhEt0qkH002vLSfGTXMyR+3IzThQ1EuR3+0KdAfgXJp1bIwCa/U1CZQbk
aWd7oRg5oIusVQ3f99s6YqIVO7K7ZDuY2sdHOz+Txmd5qffrwono+XgoR6P3rzT6p78OR5NzoGBk
kN9hbnljQBnIRSayez670un64YeXxcNnVBr4WDYt1QocMVmOUmOXkl27oXHO3xZLVH3Qmo0aGD/b
6w9ge7Zrxidnd2/A/4mr3BZnQ1Spi6RWtIc8BfpB4uFjgYwG1TlWsWnVJBMr+ACIV6+02b8iENHc
oGiCXvBtINCfhyicRfGFzxY+elTIlcw1HI/G0M8y6ye5WLUFH6qMYCkfFLLQghO7PVrhh1JxAJe4
K2VEtz6bRjSRXMN0veEl7s7G5PGcgYgCLetF4omAAoq2qDdPT0rCrqLExLPQLbz+99Ot+umjbeG8
aPLH2OtICQS+luue7tpz3LL9O54spLbL+xaXn+aS6ONBwy06jrkq1o66g/KZ9tJfR6uaeEabcN1m
XDfahJMH2uHDPHsG7iAQFaO7VS0FeHh6q1m4gWsJitHJfNTqRoiEb3oJwlsboOvADhRv0omyIBez
ZG5SX9HvGO1nX15kshYZkMq4OfaGvzk5Yu2rK2ccp0oXmHaNLO3UHgbEGaQTF608KItYvZnkIdM1
lOgPPzH9C8HNUKgw6Bnw5v12FJEeY6DvNovvZiDWoqBeCnjOFNGcvHniT7TX0AhjUHsYZF40f0qm
7WZXzd5aumx+tSboA+UjiTpNdlHz3mV48ml3eK6B5ZmAiv6E3iBkLgEBfrRh6K4uoi0KhmFoEoqs
vYmb/iY2Km5/96oS5dXozm8b7XGaaA7slJJ8baz7Sj8C0E2tX8sU4E+DAbbsyNVHHmyJ+KPZT74G
1UCtXQwbVhjZ+JSzNxVqh9xOHHOs7vDGds8vajZCouxZedCBXmUXCLiA8H21o70HMIoRzusMVcbt
qDsiGB59zq+0ydH7ZfdvGJR14OMFUN2ndpoA7VHbTmzbZz2PXabYLQ0Bnn7mobFi1zmisJ1ykPyM
tEmH1KDuyCYNjrAPTq5CitNobc7lczrezNMs7trMsS8B7odAU8s2rvrkezfmDc0at4YPnQ44bbZD
Po24bfWa3qQmOoVDgeQ3fYYki6cVVUmBx6D7mgj6Ts5cMeTD7a8XCmIIXokbP+534Nh6alhuuTsr
uOEV2WjPW+s3F45340DvIHSivPAYleUu95ISFPrqVOachtR5/u99d6qZlmFUH1WbPKtIZg5rkFUT
Ik3b7yHtzgCdOu1vMd297D4GBBjjwVdowqhluJrLd49VuB5DZkzLS0+/e94gIfFDzuK64sIyCt7z
oLLgtJEQ5dAzyW6wrYk/sPw0wb1WSwwJcrgw3z5X2bAeMb/btI63y0QQS1tj83/u5xZImYsPL0yw
71Yb8v0z3h1NxSP2AgnFOB+dYhEVUcP6+1HE4mAbGLezDrBUyJLUskR77mcVj2stlJhjRC5EIgzQ
8z79lEbXkZdjqigveQ5KstAAltJz6+tBGiElfAFoRwo7pSi7bZdULiMFS/sQvrkhDqn1b7zgCs2C
AvuazI45iONVAioDwoIqnP7giVuEMPOuqVLiHA1xBmGDOXzmeZFUewVtM88BI45gcoObF6HgD7tD
bsXJXotAod6cQqwQYLKwhQuhOLRdPBEwLAf/ykpddHB+BDRroHGtHMA3DyxEc9VO79IJSjI4jJol
Dc/a8LzLRnrNjN4f6mpVOvNDEYbUIqbWbkuY8IiLgnj035JJSlOerFhW5SQgwegU0p5EsKizfu2b
m19KmPUam2DfVwivONFBkcInY7fDjrtJazhNu4JLen8zTox3tybkok70t9nmmMlXcfRPlAhsHAAJ
Papc/9/UcYYMfZR8rJMI/kkKM/lxJICnpYX1vWOADbVoOsW++ywij3pTS5yOCXAXjMfKlTwVHk4/
YtlplDJySyGzyiHLURCDO9Ys8+7zeNezbNT4gijMhG/QjXJJKTTf95jEjcLlzCLE6a8jahcizLbk
SP1CABFW7zKHRrET/WBqYcVH2YQoKxi70Ht9wEMQ2+DF6z0I5LbsgdNq7RGkNajruPrnLVlw5+JZ
cvUOQq3P/2M7iMomOnCYnpzbHe1eWc0L/8y8iyvPTHGnSouD+JR6qfsIMBNliyj9/HVfMoM4/FYF
MyVDb3qd6my3wpRO4njO5mEKKwn7fz7EyQ23KsJGrKANwEiu+BzoWwAewDmlKDcCAhSSgeDIAcKe
BOjNbBpp4yHQsysVs0zqbY/GZ0wGvcCN0q3KYsCg0gNHQecl5i+AwhAQkAjkZbyx4frQ5RP7UvBG
fnWhxjXAZfAlHnmcgElSrh/o3I0uttJ+jOgX4iTvOdGQurHYl+raIH7tktBb3tdwAcRR1wWqKUOv
3+beX0Xbw1ytYzZ5PfvYBUBilw6dNo1ckBEMeIgah1gXt3gCk6up0xtJ6fBKV1GSdyIig6HLUToZ
uEK/+i+P2gMk4GOqGZEEwE7fN7k4O5L8FfK8LtOmrtEREnduQD6JNR6ll4n+/LiwKaDyD3/K6ouq
6NxznrcteDL4wkeQqbo4HzSid1mrMOmLeYVruJMM5qqpYFETvZTEb0dW1gB5E7DfRfTWm1kWclZ7
BpI4ZDEnuYUQ+cCrfP8y8vLNUEoafOkCzgCZPdjWcH5187RWS7xc8sv6iRf4qq2vPR0Uh1ko88nf
p9/FoISkXpmxp9l0H5znWOcBknqyN4+hkqVwG8OUIoNUHUKTKom1hlmou8NT72XhKYUiC+smr1yz
9iMQpuZqN8djCcARIhQk718eBWp6NSveJN2XnKq8cDPRMqWjZHsw1B/uvpEISO03n3peZjXNfnEj
hwpChBTO9VO/QJ5HqohYIjQsHADFzywEDwXUSbQhDAD+yS1po3FFz4W0Mhv/kxitvG2T4S8MHyfw
Fby10DrPgI11PW90bMPYGW6+IsBJ55RmpI+bTs3hDOWAutaF7HBN1UZNwX3D7tUg/pPKZ76ITyMl
MexB5332Ay1DNM3MgmkdmPpPqVehZfn0/RQZaNACgt+XhCZE0JsemVgdh5JldNLNHPjixq0ti0yc
9Dj4BKQXfbeMcS5yrvjjn9pNMy4Ia4hIp/Yg3s9yVai72cFX1llbbCcsyT9yVTIWt3Cu8St86vf4
qKYuN0NW8sapabQnL9zcXp7zqZTXRCBzTTjgEbs8xD2LX534y+Y7/eDog/oOBA9WTunVDlKMAB4S
IpnYGAi3aNbgESwZRoKLAkB+0sWH9YJvoU1nliJrRgPSKJ89qrbGiAS+ZT6nMtpIuwEBu3E4F9mr
xnEnt0hqcZOUqfvMDKYKAXB4A+T5Z6M5CsW9pWvHK4DPmBop5Izrh85XFdjsvaDPtJlCa03BvltS
8m2ivrVUtZ/C1k1j6boOkvfQUTQ2fk7ULIv61axz18ffHtyNwqM5qWx3p2eKBFBLDMmTNIX7rT24
FLbRC9nYMi72yA1UxRBKwioOftLT4+sufoSQqqE7eeYX7RV324fKYyLtvsjrvg7QKIzMGnvbVpGw
Q3cUXJBj581bnc5KFZ2BowPaB7+hmtUWXN88Mjnxc2F4CHKjLe7XtLws3hwJttiwQiooGSR0zeIN
xtbXKHzYL9lOeCkjkmJbrARoYWQ4xtbRQ5ANxN4upqnRM3qUjDas2Q2hnEBOJyd4jwbLGrpP4ihu
Nkhe3rIT3+Dgl9lNrZ0LjHcO3CGv7JR8DfHoTpNFQBl6G+g7h6L2nUAijk1XpAkXoFEEJTNq6sBZ
ppeV+vWF+FhiwEPul+7zKj692U+kHsY0XUeRmJpPuiju05bpYOOSgUhYPiVsQKM5QFCN5H3EzLIQ
KRq/H9vRSWESktsW359725lPxLjtQFgTv22V7wuB+5HzrQTYIbu8juL1zo7D0BFcBhUcA+g0EXx5
PQHANZ+lR46RE9Vwoc2MX12TvjGYSfpJILAOESuFDOhld36KHOROcLLsVJVyNzLO6YmYUS4zqvLy
0JW9T6jbOb7t2Wqwk6+AuVgJ0ePDbt95duZ2XgOF7nvyue9z9fRkOim2iwmJXbRvPaSvAHBL1RQ3
S4tFlqRxKNYoDoSMASwDbLy7f5NH4J9S96rrVZTfFQ6QfbP1MtsgHtHEyXagzC+vJdQGoOUkFwVx
54GDnAqIWlWUBfA1s2Sp/lFrXQL416IOEHUH4+yxJtpq42zQCG751VeWLfHssVphfmLEZj64v/js
qyXl5MUUVdtKUtqc9nMLwEqQwiWAdkf6I6nEwue9gpFeMnJy4yGafVxZ+OddnJ0vN1qisAJN0UBe
Vx4K4DCRiYYwzklDyi3GQfnl85mWBgSDLkGwpnHcJicGbaK97eNzBXy21kwIiZgfPVyF89AUitkg
Uh2NSS61qUr3/w4m75rCqgX8QorRkfq1BJ78rxmW4m1xgByBGpal9cpJqwEkokenkFtukEeS0sLR
ZempcowIpvKNxyuu9GN+wtHOSI+CD3OviIV1rns+q7+C3BCWYDmOzDQhSDxFdTDK7hAvmHKnNUsZ
m9CFnwcf06ul6TKCFfmop37oVYCRAGWHDFw1nTAv5EXeZquQv3DgnyZVNG4shWFsGc38lFtBbzFX
TCFVkWnMgipQA8/PsZfAyPBqYEh51d7l75H/qYt8RDIxXb5SlvMAkcKiu38+uztnJoeecJKPTvu2
JPGuuf3xU4x+Z5VEzG+Av10Y1kSVz56hUztY45x/iHv3qoBYhdRUywiKG7ucnxBcRNJAQ3frbzM5
2h3fVwRByumS8dS3RFeMKJRcHX5gQmHcF+1wE0NPpEUOtOI4SWjx5p6gxAM8sxF1/nmv2s/usxL0
zrRZBo/Y6tfFqsKXaZ37vDWVuU62ib8pcuEXO3kIfmfOHwcWmKjLcFVz78NqS1s/vzKlxh9nd6I+
0JtMNqGbOkl8W79CMzPfORxFmhWitEnUd/iTTavuXdzS31HWlnbc/vQXgIM6tLPVYtfBDMuzW5ay
Dn2dDqYwVI/irdPBFfHQbO64GStVIS+3eOeuT7emZcmETnJPZcqg8qK4wIU2+lrMbxG10aLKKu/3
vy7Y5E7xD5LdWE76bwBNjcKgJIbegil3WoO3AzE+tvY9PoN4jjpr9iGm2ayFMBE1RcbCRS+rSWzS
U6bNovS0yOOSnifIx1t4IBGN5WwatCZZCQ0osOiPrk/oCq4row9Z4qBsZkJG6rGMKnQkXuksJKF3
8JVW7wp+mvoFTxnYuw6i3qG+XJLMbKC4sq54h/Bmtyi/qHJ5UPqrmK988XCNFnGR6HFT75wP3DPS
gv/+m3g7b6359iBPx3oxXoBeEDXLqez2TvBfwk2jFbj6mBLG8T7Waq+GalLN+djhWuXAmOlQ0K34
YyDMRhf4lb6vCT+Isp3Pa2WUFVv7m4RJCVxqIxG33HZ0HYv163xzr3mT8ViwlRhSkoDiE3/bQIzj
ZfQnqK4ZqaDVBg3qyIq+bNHJ/p+Lh/QGLK9Zg5E2RhihizU2jAMyl946tuoJ7pGYUYRz6xhXT+MO
ZJGB9cdWdtOQVPmxK5kCt7qNAJks8oJxcI345Ljeuol9dvmp29b7Yq8kuspAGuBi+PTaYzH8MuvE
nEBkQiFrgZIfl3C9Ckfylxb5SG6hPC/N3IgC/RNA4yowklbA+Es1xOKLEs9J8IPuxTl8Wgt2ZdGP
2rNmv3YXW+x5C8FtJCxZVt3UnfOTFfWVOAdhpckbHXNtoOQkvQeD9DLC+RRdlXYF/tT5thWzd4Rr
cm8j3kK29r+EmjntyqzrjYdul9r42EGLMGGbLt3/262NVsUIq5pR2GkmaSAmTnUjfEnqirU/98jS
7fw+n+OloAn2hPMRE32gX402sPuGvPszxoqs1UTn/bFCWC9HrTC6AA6KStYFdq1rqn5ykDqJiO1J
rSiPuqxryf62VoOQ4SJ6/pAluZWhH55sTHQCJRZMqdH2M1Pytmwuo5zfoeLofDJFWuuBXE8kuDsJ
xjAxf8YySK0JvJKf/XnyDV/LEyFZHSHkV+PWaUHQo7opMZ7p4KpmZDb7VJKhwxUyi9p5bXo7fJx5
HiMgesNUPO68o8lq6nT8RX76QCLeahirSRP7WOJtymtg3DYHEEz4/RU8GyIymMuh3IDljFd0PFeb
h/dGkhtehFeV6rfvy9ckxrcjHLXuPrBMMVpVC1s6IYDseIL1rCc+cJJ1g0hJ66XvlW38pnKnAzx4
IdqKyrwOTRVPtfSg3DqGcFRvEjoUlv6tsaX6q+a9gSxhbZVLbDahNpomv+dFqrqhb5OG5iE6KfHr
NaVWmjmmeQC1rkw1f/geSnPR3SDV895axbNjx6OarNcte5MSoTW+0BYYT5n+eYC5+7Q3ja6z1mse
tSOMVbUCLnPk/zEh8gwP/GVa9epGvwX0gATh057s0fSaZ4d6q6z9zjTK8Iq5QNq01FNH8sGPo5u1
Fdo9zAmw1tKI1ETrdr4M88QeWEwYNKVjkFP1WqyNFf7j8JPqCKJUSbCO29NigYUdFMB2X8krzEyy
gcZlTGlpy8Pj3mqqVQurDXCLs6w2Oh9nfgCpOuIfZ5Brjxahw7nQLgdRCDsuKKE68IURWLyblYLj
V6RtYpyQdqtOme2kNSeEufCPGzRPQIpku+RLHeoM5g2ygUXLFqJGFUBnXjOoX84yaHEe07yu8Dj4
BHeYQ8LDCdyaWfS3BrHP8HsvT+cbz9J734NGSpoTDzx4vKl9AuJdaQg3crbJnP0BjG90r1MD1iUA
J1KLKATKayW1eoB4VzvjKhgKzaJ5F2sSHtUJUquSEmRZjp0ndIzIyf6+fTZLP6VlFnl4j9Mi3Yug
1adkS6W8IE4kENg/ZL5g/nxV5VcLrBIO3by8WLTnkJcx6mrX6affKeTqp0vwzI9jbD/rnctt39EL
xpIBleZy5IvYdtzl56GzEDvPqp+vvRYnx12OpA98N/uNkybTHl3ISTHwQcaGMwSm1gUGn8ulmkna
V5Cg0Q1cKWTs7COdyhGxPtBW0YOhi7pPl7x6FW3PAjEhWkrvSDRG4b8cwVYBr5IzFfRtpHgb3C4d
hC3ti9NoHKBLr46rruB0VhDK//4Rfa52fSlTmhFbUjNd8UIpbL5maBQzUykHykpK+6QsDOOD66ns
/8gFgMRwAt5W9oPTv0fwWaFNCj1yJGf/aCGT5xgWEa2e/C7GgkIcRBgewQXpcesg1h0EyA9iGlI2
6ATQ+HysEi81oXwrOoPHEGN2PBx7q5nxK9y8poJcLXmlv9rzU7OurbWRrZ/k1jLzkFW796UZxaa5
Mn0mkSzbxNn0uTyX9VHn595PcJ7zy+dxA+21kHmG49vLkJsa/WFUU4mzD/v7ZGnwOc24nlUCQSZT
Gx7zj8CtxwjgwmsTYs+m3eqznRypbM/hhfst1R80tsB3z2hrgrrvEypg+pOwIlfKnapgB+AB9MPS
TwJosTi6RegO6urVXuWDS2HITEaKM13e0a6ByNW8cRp7r3KGVZv/sCTCvyHhbPf9xzK7/ho/UI9J
UeRC/MgBXrIGHIDusR6UDvT5eW0b8FUknnwlNU3Nx38QdQHKKMRNweYI9uzsUFeeWlxYqWVtn2gJ
+3ppoT68mNHGXuGZjeLKtDDVFtr/puZO56itynU1pvfs6lq/MWVgHS/Rw7vg9UxvCJAYkYySnCyE
3vUZjJJNKhcybMmZuZXaCQwIDl+EXatZCRFVuxCtRS1K3ScLv/CUSXDD5R9+m32pK3CSgxlmjkg6
tl81jEvLG/0TKZBHaXYCPHarAIgGlY4fazxhuMR6P9COY27s0cgPl9vuHabvYZZyB1wHx0DTgaBU
Nar0iMgncB4fDvfg3dm5393XnCE+oUHRC2fpt0jt0liBaGY+AsFG3FJisk5obk3j1EcpU3NfreYx
zD+lTNl+9tnQaYHaDG4vv9gCVL+GC4BYBpy+lINs+Bh8m6reHkXtzTpUrw+ufY6UVC6JSywqngXm
aNOKLwzG91/waUBvKoUtF49phD5cHbtDxMuf7Xlfoaqouv/bnCSsZKtDju1yJlpBsg6auAaLwX38
UcDb54KoyrXVdVLAvEuEUaA8mpWlsv0kJ2LaVHw7w7q3j8Wj7qsU46i04UFv9Tcf8DrbpSeRuPv3
0dmBU9wuHgn72bfKqqHESVdQ/RnFFDM9VSw3QD59IE1943apQwjk8Pt43qIWfbk3zcj1VgydbEwP
6miGmYY8kBx3vPHXQHS2AtpXfLPiZ6svEI6hnPKsPUYBv3IQiCkgmIZFgY3vsiaVd4vxO11Rh0ca
hsFMOQMkdpb7czQp62QqPVNFM+FOE3Mwi44hBnbBpEebYGQC6kzZ8GO/FmoDtzvmYx8sBBybqWUy
YNJFnN7fs6HfBhpSvfxw6bn1kWXGI6Fa9QMKoZN1ii1wIDxAXiu8/xiTY46fW1/V96leFyuA1JAO
3Xondj05Ul5hQXvZYBSVUHCGMJHD4KGm3dzpHwi29k1lcbfW16+zh6wtKWaQ2Xmpa+KiAtB1LDgk
sEG+aBTZ2OwTkCULL1SKTvnmu5utB/ObZAEP8gKNqB/ToRrApdFyGXAbH8nNEamzOGzV6COWaJYi
3ak74C47q/qNvgjxFVr6ARM6DXqpUvOEGjt2zLXvZvwkrK7dBJ0msAgOSrNMhGsneqtvyv69juC0
War5C0QV9m7fpfqi6XJ5NTilj++P8isIo+J0RPdTdAfzT1xmALgZBb5ja5I+0XaHOeJqXH4QEcLn
RZnLkRvhWxvqCSrKzJkjvHK3ccgCPHw2F6Vsk0YahvviGVPbD+ChpG7JuHJYUOYuU8wJntj8PZFZ
RlnFPh8IuSeS3C0hN8g2nuJGXX+aRYs8p54CDdSLloxekpIRlC7TLQWhHA5qlZk+K1Ofo3i+1LBs
x6cRa5fte/cW0yf65tYsjFmWCpHo/IHxhdanoDaQZEpDajl66v51Uqov5mp1VtSPcoq+V8Hjv50e
aQK2sZzn89WC2b2ORoKkKtLCx6I0AZDNUsIKAca1ZRk0PdU61wHZLIxOCMu4mZw8VOuyHsNSo+XW
nd5W9qEsNk44r1UYLdbTZx+ZS2PlqRR+YMrg9ybiD4Cps0X3JX65W7y70lcSUBxkX+wt1LcRjpMn
RPqPPvYw1D7ZmMmwMVnA9fKFIlFpNxGn1mUjNXzz6sW50fMEM8R5BrDUjD6/TlcxMyCFaOMBPpIR
8cGlioMiWIYGvVwYqOmXaxV0ZfgICaEcpPRyLdUgCXaeabyygH7qgTzOlNGpOo/VUpUuHh4uRy1h
ebhAgulSSsCj1hzBj03k9tgDjJa9QrdJDWm7lwrOx6eNYF7d9lueCL3x+piV1VnNhvrdezgVtBSV
ZqPkfDJyTFg1IMXtzbs02vkR6tJo1BJqNV11Ck6e6Yg5XJ8O4BcWfr5Zs9yqGWu2wr2JLwpV6zIL
XPbvn80dBuuqu7z5X+PGtOXCZsgYi69YGoubbsqb1GEY46V5ww6vwpKVwS9J3b7cjWvMGFk5Jt1q
Fz/sTfa4qO6vjstOneWF/vOwTvh3IPtHXFY0itLyURj/j3YfMAuzb5Wal3d/o/xBY1GynTpmU21j
oPf/sAPC67LJ3gkIruT4F/+NBTeAzJjUGnuDfJXIykfdfZuGUpIxB92ZeuheNervaCk28pDJPLO7
FBT++B4lJktU+N19/fW06OxEM6QP4VyXO1D5GW9H3wC/gmBe9W98RNZv3V+x3Wl/p06BP3ypMaoZ
+9vKGRiLxW4IvJc7xp1okwOO45yxw38rZ10JNMcmASMSReJCreGTWmgRCYH729FicBv3aXCKJ7cT
soLko5oU6BjQs9tiPb+kW2bdQZ095czE2O5RutY8Ri+SUym7Tc+QMvr6lukNZzpBs4BGOVqiZMtp
iWRTFTZSm4hp7si4+4kV2uF+Yw6Rx6a6LB1Sx1BeZPUPzxMRF6abUnHiVXFaaKbk9yNXPyPAO1cn
IrPS/nqbRXKnNxGYSRxXH0Vp5vNEhRmBZgQqIIU3EMIVyjr/5dB35VVkwPzaAZxmupfc8SjMpQaq
aOGF4ocGBwkNFbdp+JSweoIOJagdN6dJyAr9OIh2LNBv1tX+L80g4IfQANssc4/Ky85VzMwhDrfc
2RM1Wc6WRVY5EAekkzg0y+SHdd+IVjaMcyDoPPdU7B37wbF8/QDd7RirT1zlh5MHXbAu9f/VDbcT
Ne94dteFi0FEc7BXVreP1mlvfCgapogpBAD+p3e0CPgufwW/+YdWn0j9GbkaCRyC3stdVaAk2UNO
mrpMZPfe5aSL24HjfkZHUIMy0dPsiUideRj/wl2W+vgsghSic8fhPvWf7YRKlxAuermAxm3akEKj
DmMgxhNbbAvTERQRMlBz2lIHDT7pCc2YXoTuL+8RV2IyZfCXy0ab1+rT1Sp+mcV+NctBQJht4ut5
iib4qONyfVwqyruvefux5qHdo/7vagENejY0MZT5CWijgLlnXzs/D+QAlLaGn/jIS3S3tLpjbsEf
4hJwI1Uh9T4isn09V3cbhzn5wgrMx4rplVI8IuiW+mgjZQP4Ow5L7phuEM9QfGJ7VoJuLDTq6iie
7JcVrQW5gZ3SoxDppjghmm0EYdcAnGTADdPAxpWi+vcGqVhKG2A/ZkWicyMnnWngJ+WGhY2/UPHs
oC+9ClNzIx9uwr9IJKu9c9t86qkaxNvlFAEzno5avrWTiCABVq7HxVK7if9f2ADmSkcmOivufLIB
w8MjQtUjOKHwWncqnqmV9qgGrQ/nln1T4M4eh28n/tLpGZJbMtQ/OHRCp5Llm/1/rTZMdYpwwd07
AaRJSeJLVNNfGL5YsdViTxrPotPDqdE79ea7EO1Uie6FUTKzYtiYara7gGE7xEN8os07WdvRX7db
HekBU0fY+o6bfXAHc96Rgv1giz41TKmq96/TP3dmMhpYx5JYXQvy/nLNMAnIXM6uDf5hXVuclTeJ
JUKjXl3TWtcSyU+OyesiiBgts4avwez1ObV4schmxxV8257F74xY622cjVRUmDEl9Haq9SLUjbvD
99YbCo4yDcO63s5iBMYa2dOtvnOteS1ZAoTjysQBxgAPUod7e59Ang5ljzZJKP4V21jSgO+tO1W5
hISx7mH6fP6FO5zT0kDIcFZq0nMQXglyeOFshGO7LI6YxLqaRww2CK/02vSoe9wGcTxPyl4HNmme
hizBtBLRdMe/t/kaYx69OoOsHC74zHJOXpPqC/fYGpWcZzLdUNYo7uthWn71K02dQk3CZzjJGVHn
jYfGfjohOBuT01Ro0awk6DfHjuDiK2ZebZ6ypJIKTN39biRbE7MCA5hXnpdW/6pVdxbsTg82G81C
od8btg0/koZWpb7vPbVd3MqfS84OIbZT45txgpLAyVWxEZl4yI7eLxgplYQ2d5tJBbNWDQzOVrYC
5s5Zv5dDYcfHlwCwMvEJvx/7Oa9IW2p+ZDGYy1iyYn8Zl0Nmop5skB2XlbDzTGBCdBwrq6v2mN9C
KBM3jqDeMldRzdvmKHvAEZ+wL9hSFqMkfIey60F4bjwqJuf8B2r3kgVFffzLinO0eB6q3MEWicDr
UHIV/W0d5Grf9xtbropuLp5IKm2xQznU72TrNcHNMDP37czoQglYRcKb23AR77A7FNYT1Oo2scFq
E/Uq74SMh1s5wl/zJOsuvF1zY22WCHUQklK4xDvNBBRX6jC2W1z0K4A+EMDptt5tL3wH/PW+Ur8M
0l5KBvqEr6heSZvITte/okpAod4XbtuOxJvr5W1UKxtiUDR+89+UcvAOigTTBd7Ibae0VvT0t87f
pdZyCmfpQ779eOJ/R2S1BsBLMRPQjIxEDEMHRFknVz0qCYdQbmVlPAjhfuUGl63q1TRb/BxHVtRN
8dK8xOXTJwozWAUrm2BtmMQV1b677YRkrSH0L240W8rlj7pki/DgptGztNMafAnQbB9+dWlyuobD
zGtKLu75pXk16vyy5xyESrrz/gNdM65eCpdXk3+ef4dvwSoQy1yS41J+mAZkZYqIhSLfbLNlCjjx
2EWVIDsSxeGm+ax0UkBBnlEcfxw6pSWjl39y2A4dbaJnH4stKWnVWH/bwJzUHpbTAFw6InsiJa8F
Dy7cFS55LpKh/h7qyOlzvW7z/7c6lrD/WFRTm5aD0VZ8bfwR7XGcWqmo3mj00WN+ozdHC0D2soW8
Ucp4mRtDx/jWprpSUldG5GwwNC9gn4Z4mWg57zf9EnkeaEgQtMVSy5GDO/nAR7bM/E0qg3q8nJ8I
qfZo+Ju2zD7CK4zZYPtpKXrr0y9DtSkdf3Ieo3dIttu5S+nsOGY0ejTDEpj0hBL289lg+r+Jc9Ss
hTU1VIYDa4fh0j7uOun2TqmVYrz9w5Od0NZIIRIPhiKIoIXlf8GNhO8zdiiYjPePdks7etY2M9x0
iCQHxKTXka+pEHfID8rEYXAbM01TFl4UTckrFIzWPXNrsRFhUJku8EexeetApbmJ5AtqQ9Ah5Qn2
rESOzDJ2O3F0ZWrfmPPiQ0l/6RhbWM7dxOV9dRvAXyPoHflVspZR1qlgOY7Lm09y9e55Ra2s3jQi
7yRb3v+uzY9ZkIdVOp6U1IubveWCVIDVNjelWRlqpBoE2EfkQSvMhH3pCf2dnij/deh7y850hzxb
Ndw1UukkptXzziHv8WXM8fv44IUxlNhIL58/LcsYkQxAp8LoWg7re1j/D2TuaE41JM41XMaSzqTL
croGbAQYzQPLHppr/gG1DvqevyLuXGu6ba6U8GczH6W5UTSmVr97gbjqlZmdF4OhHGiCmC/06nT3
ff/knRtmOtNIwNc4ARuX66ec7jBoReQ4BMZfV20ST67dcspC9Sbt+ni/vIo/0YaD+ak7Hk1YCpSp
lE1qKSa5/4j3850dpq1ryXIfu2+7arGlXZTBl/zH35ZZRwUShM8iEiZRsLbF8niCnluT+Ep5CIcN
zkhXL2zN3VfXoE59Cc0lmYbJdd08d8bEJQpJv4EsZKFLZ5LgzlMuiW4HcWIQnBPJa/QpOUUWEyZd
uYmkzSBCv+rTtKj0DXESJOhi6DHP+ZSJuXu2EhvQiiKuiUSIFXNOB9CljBpF1diKx5sEpmW6p0oo
5X0A0s/Iri563cZVBAEv2EpNRv8qtgz4kxsSfgkI0RPCQahWjBZK0Ay7s8rgJDQH3UOjgJWh0O+T
fdcByJeQieZK1HzchTYStbyyhMfiu1sca3x1k/6QfrHdUEjHI4ucvoRanJjZJSz1esuUfXB6eADs
4x+nIOkjjNEdxe+heMQL7qf1eSDZSu7drKruY8g5hilF2zzkswESHp/SaKKim/Sgw0kaMXdjhEfr
wu+Ei4S4uKvZWxZHogOojM7ISHeFUaHLLsobIYc9ou9+pzB073MxKC+Cf6+6KpQZOntPWnCo6GBg
RCSg6SjHFabZ8WvRxjEEsy5+wbi3VDXKwY39JiLE5OKRtGGix+Nlv/0fRC09gI+oVZlo+j3nMC5a
8xOiiKK0qGbURf7KQBR4mLEQNGQAkBvw+5h7irJGiOKx7Yqr0g0oOF/HZoskpcfBTWo0vLTxMlxX
GJX293cmO+3mZN49tpsny9oEOryd5t824us7sp6UuB/xYIYsFz8ipdsnrJE/oGgL6voIky8M16Aa
KlRjW7yucjeuzIYTQSAG21J67/3yFHF31d/3C1frxflbPuRdgsXa9sCaNlnCgsgNggtc+HRhUmH1
+0dgQuOC5az3uKGK12s17YKI4af5DCZqZGa6I6jtZs/3mHnMxHAlpnYOnED7B/hBLnWlhBOlpNg+
MMUxKatI8ZaeEKsQgeVxBzancbv3Hm5v9Vm6qBiVPEaIkUXeO41XvZortiXPvnmgrsHAzYIrBWaL
C4dMLGxZnt88slu1BRG63B+M6d9mfLZ0ZQuq3JvNkBzzaSlcyfAITO9XnLZXqE5opg2OtGfplpPU
EOewrj/KANZH4jAZbe71IFlzvJL3JqE+SwJYE7b5N9TsFPMyYkrFRlcvCzwA1G+gISQnOYYXehoo
7ueR6zQTqmjMNMCWQwiSLYGarizsOFAA2BD58xYv/hG1LRiSX3dW/339N2Q+VVdcd0Y/u2dLjPTB
WJSwhbxE4Y24Oa4fOJk6Fcd6ab2qXcP4YndZCw9d4P5fM/yb72c8+j/VOsDIicdLDB3EBKXwc+0i
cwUs6Ez7Z+JXkl8WkJJ3Gp7WsgGcvSFV4Dl3XgtTa+YUVRtk2R77SxpBXFUa10meKd5xin244xUZ
rhXeR2OLYfLpM91WZt2npKFaI3Bhrof59BCegVjm27/KmchyCNCGt0RtgiwgqNAAsnC64o8mAe9o
j0HiAAm6fXV3VzU3ayFNKbyyQgkk6N/JbmSahtPsoRzJSIIZO6h7WN6zOhAH0vpsRCeeZDdyl5Xj
EeFaf7TXFCBudNgjVcLDuS/DRDPOqhUGvHbjqUW8Gy+AFHlVL6ICwvEaml3pqyAbvy/B1mN9AABg
YBEQIYEg9I8Pt64GitHBg5I0c1m2OkWsduL6TNXQ2ZLP3aHNIBxzNmtyT2MZxYsX7JWvEyBvSd7t
PuZdegu7vrM4j+Jnszz8QZ0ipiItELzaEYt///2EPIvLLALiiegMgx8DvP5dQZ+DBzRHZx79JG6U
z/nyMq3rmHbN9LpPNlwezXfnd1g8N2jqsHhJGcJ7lkTaX2a4MKdUc0eKP4bJ8dBPEGQ4U6DB5ytT
vsr2aB5SCyPI3qXiegmmNCE7bek3IcfHcwfAlWjynvF08wunVBzMOW8nVxFfBej7thAHtE51crUN
pnojMx9PF4QO+q0zU46y/As2NDCTLSZBVKayySZfGf9DYuc5wBkz7xKTPynLD4sCNXXQ9VGrwnmE
l/Zb6pLxp7kx1RTIOVqfjz98tNlMCNFM1KXrIFrbg4BSDagQVScrdo6SE+22IugOSHAqIixVB5pz
Z6E8+YIxwwc4sJ8FhL1ZC/Eb8fHW8oDe8+aDVffz3OT8DFQoO0+FpvGktewF7TrL5ZxKJ7PDBzuB
vNtbj7xzmXxW+ThoGkO0rKOGkrAFUZdV6peiADdxGaQhm6ee5/8e4+Sz0FvyIj5lAy0U0HgAJsPl
k+z/J02CL80r/otEXLLOTjiBGP5nzHJLsgxTHMSYDlEq0G2yk6RQ2qtrpwDPEkbdm5p5pCgL6jic
eE8rReXe75/R9j4HxqKvYt+7sMQgnSxqJ6GZXA9eangFaHC5gcC7s8PIzqocLFCYOSng2ybez1EX
1NPNgKMmsI7GtGVnhaajkoedJ+cODrIKJcMqu/ByJ3e0xfeMJCvuefBnJyG4qKcMZS09Krjq+jgf
0lzQ9wVpv+Rox2akYbRGhynZvOFMpXGnD9i1dQRS3wTijET9SdlSpnyY86SgxrXtKudLPz2RWmN0
pKIWXLrNzgziZNCUXcL9lHtNJASGMQI4ufHXxP4lROTmHxWVBkUl2f0aPes6+xcHa0qOmtRHvavL
SPGmV1gCAvRK9puXPuqoeVud6zeGUEasID1UN5Pfru3Q9QukdBWBUVKt7XxCwsii+b5aIj6DJTr1
90sR5W6stXlKp8RFXBtsVBIHyOU4P/PaAONwkh0nIFcHa5qi0+0BrGMwyrnWNfmTi21FuCtyWLFv
jbdwfZtpHZMFpMq8/m/W+B/hPtiocpi0UAs9B5eJnigAptK4iJMD9OUGGnefj4q/Hft103ML49Nq
N1AJX1PbuPV7ZOpDw/FdOS3QiAbSWFR2KSdeqTJADMsJYwH4W1PaWEfTlEf7qzGs7/5XWYg5SFdg
P+q+SiQ5/YFtbNo3kX2QuWRhfU2+RCo21DyIResKYUeM8LCBuchoWxPtoc+do/Z7DQw26vU0alwK
FDIq7lb9l5boNL/NRt6qs6oFrBoZm2t9DDYUKWtN8ae6/gOyMMDK04XW/b4FRiQzQA87gl8VujrM
ZaVYf2KF7XHi/twZdZzBhvpZQQczuYssDeDCpCgLyVBr07R6rK3yO+TNbVyrrnmQQz+WeJeQ3X9K
VShU1aw9goiFuI2SWBPGKA0o/l5Y4PkrzorIMxdQHQeCig8ibtcPELOhcZ59sByMaVkFb0T1ux3C
3NxxgA2G22sbHHsUtXr+DK/zAKoMd4NOtcpa51JSb4/C+C+R+ttmQ667RErQ4NSJOJUUn6D6KLcy
1rRzRNR27AjdIp6B5D/b/X+pVTLGnkesT1+l8/W7Jtxt4cOJ12WWrLHurSw3t0kJx91xzPyAfRCx
JER1zUqv68Seb+YIH4SUnuoj+cqU0WNyN0x+c21eXjYcIv01DsYIQHHBxmLjH31Xeyrsia6iLqJR
Zk25hx/dbokVUqFolaecfZwI0UmdE460SE3nBksFvJ1j0wmam8nggcNJvXqUfPtdOkiqblQ2HO/I
88ORYzhwB/R5p682w9sujotxeCFsEB6xtb/s59EGHeHbZ0mPVlnrTQpc8SXYRLi9I63pRkwGQ+EI
MzkUIwrGBCaYAWjqtMpRgUFbMkpoC/ZoowNqSjZHjUFe02GPMgbKfcbHUBL925W0kYUYgxRqOsBy
kUWEFNLuF/EK3SRAw1FdOwLCcF0y0h1vlUf3MdWny8gCg/SW9twvKcix/uXJAOFNbOAdG4IrDz3p
8Utg8mnNCRD/hnHJ+XrhG2GL/5Ns0TqbtNK9VM5CxMg5mvDgDfQcN0/8KMyiyT/k30ds7kqvVpNc
o38KO4benWiG4bmfupprIsIKUiGDyCzZzw/AVn/PGZBiXM2B/7kIEfvMGoranHHYd6fQtV8ecGmT
gZbgkiVaXP85Nl9Ml7tKmQRw1FjLu/yZ1t58Tpq5D6kMcjMq5unhm2q0h67kBp90mhAk/f6yFySR
T5Lb+0GAw+d9n8lggEyhuyDU/KFmkggEOW1Lj3nK81TPKuc1b15cBuNjOOmn3tolFA3SFNmfs+uf
Xzsik+QHO3hzdedJ1Hi4S6wzkLlaBOCF2jLSNs3maijtEarWWk49XhX2QWBtaU5AwgHhTtwDMuMY
oiUcuRTtE2hC6DAumfMCit6HwEmHL7pxg/KN9Xo6873wE4tDRpQxGAFJkz29oB7cAxGZhw6VX2gW
tRuXDkNx5dCJTYyJqtGkfynkbAIErIbHJiQ5LsiqSO5VJ/3ZE8kiuv51iP9NznMfbYmebf4K2oSK
C0uXdiVHntxPnu3xzmuqhoYGWLNJNSLlwzk5hZ1PB5cXsIlyl2xYsbGTY+5Pml+RLtQFwqUr+JH/
79WUmc6gtIOd8Bw+sXOObtRNm5YoRMwAsSdRR/3C0q8MqMr5gt626gEHaFnvuJup+LlERnfIOsha
T+EXq+q37fbgM27bYtdc6V1WQYJUgVsawzKt02U1U3TsdO5ghphM7gdnRMdnzBeVw1/USUrXcYP3
q7H5WBZn7HnWN7XRAQOgzESaZHJT552UUmM4GXlzCkIxFgYbme5+UGgpRY1V4A4w6E+VcHM9FvZ9
/ukC+j8ITpF3NN76nBlBZhsWvPzEyJJbpI1/S1OcHg0VGblA47eOG3tykc2NRvDggvcFX0WXtvW6
n7sGqP+G8Bn7zztmS7/28UZazX56/k9xowHreKIORmN4JIi4lBRuG9GpR2HXLw/wnJITAYMLHlNg
EFQGh18/iNmdoPeiWfvqzpqiy11fSufoX+odwRm5/Q4IXG4j1gVoz31salaRNSLjbjeOmzai5vTI
ow4qrG+LytkHtjUPbnitLAYszcNbVg65orG6sZJ87q+rgXgIG2iGddb0VTYYyFNsOWjaYam3NMTH
CbjSMylcznZmxwO2nUJd6aGHnWIFp+8/x3HEceUnemNxY8zRkNyu1kwN+NChdbCz1zRSZgtviq5B
9Km7ZT4YpEojx3AfSBRUgKNWTCDbuHjwptVNV7ykghIeqc8YlmVNkJ+/8+eARqAry7DIQiZVQpiG
/rT4WIHtgDGR8/9zNv8au3TUscDknwJOqGZKId5SjVmHZQnDmX6pMk+PyxDZYradq5yxXCynlfqS
RlG+j26wwJSJpBHsbDBMtD+Y+kNuOZwEpUIMaPtDBX1DV1ppvvfUz+wGga4aeLHr3HCi4B065tGC
ThNKzRND3QMpyJaYTFBi6zYhu4kNkHt807kWnAQyaaCsUbSsvUQUlr52bv9nkVnG9CaJeuEIfK8y
fUkfNsroMmblvmSBLAmjef4MS1LORngznm0Yauz1jIsb3JVSMB1vFgjlC6Ezp9AJu1le85XLpa8v
RVeORDeptbj2Z3jDduoTWQMjZyGOtXEOZHRm6FfnBCCt48t86gpfLKsvG+cJ+mqF2tY6rx8DPBwt
B3TP1KY4X30/Pz9vFTM2ksbmJEP4QvpqU109xpb3CJgxntDDToNJxbt7PEk5964iiQy3PERv6nHy
Xslq/G80fZraNU0w9ruroCO3NBfYkkSrbWx0C7Od5gVV5tLnZM7ogJz750WWeZsOJxRnHJUKdkNQ
4xv68jIUQomKzqX1awweW8dl+OKmosRn46gU0iQ8QzAs10Y8fxFXRw9fV00UhsjyGhoPQVzY9DOO
5oU2xc4Daxo4Dlt7tO6PlDZpkA65m5LDrTQKGN+2Y+/Q8rPks/KRAVQ0Hj6nFjzBzE3cRedylE3c
DaJPZ6UmQsM7T8Q66FwiR3WathqZB/JToherujidoS+aVz+RLO4MYqC8bZHYPoh1FWKJTFDgZIds
KXxOver89Bi75DvtULMbzVRjZ1AjtwPJqM1aAb/UYVlNhwrfj3SvKPnJ7xqahxPlOtMkoB5dbXFv
WE1fDVhto6HlbV3ZWrTcssYGNiT2OC/Vf9UqgboI4azcfet3DrbXPBqmv39hIGlgyoxEAZZ+HzA7
ExMMh4pzXFLo9w6pHpd5J9HEQ8af6k6VzfrPH/PK4cEH4oHSpaLUpu+WCqBvYRW/XRxGpIpVPzvC
Nc/mwDgBJxdjdMslLxiqT9lxZTcrVsNe3uc81d0/c9xCFFePdEkIFmdhU8cBQcHIuK+rww6+SxcD
OxiycAhr//Kr6YF7K9H0vaZxL5i8Gc6hqaT2OCaSz+uJQ3CEHosPVN4FRydg9XmZS+h4H2UtNNjs
UMWw+OW/OCfhGzcG33nFcYUaKoJZI1Kl1WzpFwKyfUf6JU9QGCLz7SowbCl8Fy9FI2gcMsyTYDSn
ZdKJ0Va1Pu6fTsDpJcl5avF21Bnv1Wf4r6SD5X6RxtUW4eFVaXw/gdL4ZDItbHGJR+r6dOUyQQAs
AR1UVrr43vrQDKLXFB+gOxjwtXYMMcub5IFQkLZ1oWSLVSyFmP/RJkRx3eQTZsWlA2DBSD2KCcUT
iajgoCQDghUyzXiDPz4swUJ58c8G7CjKKk4HT3t+tacUJXUldP2nPGGE4kir5OZQT1mULI3SOjqe
p1kOheNeihV31lDCu75wmzgzs2FpafWT34pyvhJ01a1yJfKzwHyxhK629JsDseOSepcYzJ0HhVv9
sGAaRpeQAl5cwWrmsLpterKdqCJiHFWwEA36or+ccU/JxTaWOjpUHrs8rhdNis+E/t+OMxaaPSgZ
dhpvR7dOOWWudcP1AxJNfc8JRn03VASVYiA4dERQbuLb+Ts7Ar1LPzuRWJO3FgCqvoVKciFXiB8N
bgoXlkK6IrOhIo2XBqDDmfsv+AbQ6ZzTGjpV1TaEoUteIe2k9CdyAaGfG5Kt0QRTyUpio8xefKIf
FnaHuPyYue+TVDc9SbIfjOU9my+nCdB5lrl/txkj5KVCz12J7W2y2o7h88+XyzNpltf7gVTfP+kt
Bg+xM4dlUWRX/Ip181f4rF4wHdJ+QBC7/8qV8kFTiAkxPrr+4ru0Z88V1wKAYGZtcLKylLhSInbS
ONEHSYHAZQKMytGDrhsMqDu1BDnv0a5PKectf04QOqb1SLn9nr8kzcu+gVmNGjL3h/LLkKrvdTBV
0e3VBTvxoluMqT8toY/Ww3h8EnNKpNtLhxgrSYf0VFPnjooDE7eSTJgyQ0kFoN1H7iU+PxBivIVV
rqS9BwWZsO2+ua6ulrXCNW7GDihwa4MiFL1xbLs1GOAcin6W8HBzPj13LtuzCuIRaroRCY1PfxFA
xQhSuEYjV1R9Y8HpXM6+zlHT31zneYmaqWh2iyYOddBkkjIhKX1RFSQyZM4ipNTm9VdOHTq7VNRv
TKiNH5nPC3CllzFbBCysvwD2qAIwc8Rwys5qbt7J6WovvwO/Ugvjbk4cc9kJ/k8BvPclFWAfLGC5
4Nk9OGxoqbiQlnBAyIQZSblRSVCdS1+4IUw4cNav1IYZ5rXf34XsSxpNSXdI9qgL8GDcuF1xxeBl
D9o2arBqiSqLm/ggRvcm3/RJ+g+qAm8Ydum/THSappvX6UXhrOEpvSVEtRYzf74TEJvM8UEohFci
cefZBxoPe5292NqdqjzQZWY7865hh1qU30s7MUs6be1jg9xsL3Ycxdeh1btc/wk8cm8NjqDUQEEb
Oh/LfT+2qmKvuWzVbXCmHk+x8khVodpC5Vm2V5BVhobkcWRUOO7WSUXgfgHQHRn1iGY9skjlKfYE
XrFsf+hDf3bmoVT4AzBGJOpqVeziZNujCM7/sPm/qOnSU1OX9GDdm4OFi/U9O5medvbbsyGDHuGr
sDvuFgYJit5gBM4p4eCKX/bQnLKTI3yZlJFohXTemGyKU6AT0olQ+CmCUMXkANjsGn91SIi7jdUn
yczXcUWJazKeuksSIiMJS9xAt5KbsrfA9JRPszKyNTUB2o/nL3656RFs6z7kAklWI8Dz/+wfvyvK
c0j1bN6z43S9bLoe9P5i5Sori0F/QJkwwU0qjteDBIjWftAZdaQJdRMwTuFJCjTkIrDCUiQf2Fts
t3DiAeIlf0cpgejrECOU6wfRQC/ZS2lhBrdM+fe7rs/IijEDzAcn5o3hOZKjriQ2YDHPBAClTkcg
qH39VMjvbQypry/PsDxjShQFT03LGRG7mTVGpQLTlOaOtEW/uICNQwz18AP5S7JYphzjscnEZ+8a
e41CAiForF3F9haATn2HC0jfpRL0k9PUhzBqFr4uSMZTzMN6X8EYa94BRSJXw7mPxi3eZyLE1owJ
8jy5gdyXKo1bHeAjvxtwRfC2nd6rmK8DffknoSHuVO9+fUABWrykoSmy88w/eZ4vkCp9+TYzI0fZ
3/mmOJx1se37ns2imcHIfOh37SYEtfxE0kJ9YEX5n/FruwEThKJSgeo9cicXKZftRE0t2htW+IPx
QS2WHX0websosoXRrPvRzui6xajS4FDcA/DwjSCAES1mr1Rp2VansfBTkzUfa+Q7gMV20vhdzeH0
+5nCGrlEse3X6amFG/F96s5kX6Uv8t7aecTeVUKjNrAu5E+i3/05VPaOgH27Z1YneeHa3LcI3Dnt
7YHyvU+n5wfsHNx9luENq0/MVkC5RA5d1f7MYe2GblnEQkjdVCQ0X7SBhITODyFAiGUVgj3SULXw
SiaGILja1l8Ta/A9dQ8jBhdLEBl4zMupwXD8kGC9B6R3sHkHgf4+ELQj5uzIDbZA/dA9QJ2i+tQb
2Wm41LPD77hBRU3fSKgfzo325kCC2KGkS1lrenO2va8sEL3xXDFBiN376ITQ7F5p6VvqBV8OsSU3
I+/iDmIP9qwDDnep1udOxPjesrNxQFrcR6CT6fteQ5C9cY2lwtgW2XzE0fx0BNB/IOdBZX+PJcna
mvzjq/ykJsnWRr7VeWLS1aoBLXoyAzZv40rqDq3m6Y+OD8K+C3IOYClw48aJf7kdDCLtJpFizK5P
2CO6sT3C36+cY9ThbC3HgjPqRoHP5tURfgoCcXd3e6eia44p/KC0xIO+eO0eumLD8EWFYUiUkpKz
YuKV0T0uYaX0sJFqz7PHGbIgdtG41bVXJNJzwLUic4ofGQT3zn/cSrC7ty1t1XMFSKYsJ5whcs2W
nl3a8kM+L6bKAOgelMbcyhuVf2HgpRmg+xP0YTy3p+LDez2JIHSr2M64q8YHmbNyJ2+Ok5ghCqZY
CjRruVsnkZvUJXwSbAwrOjwho0rJ0lPKCbbU+NG9LNUZWVYo2hIDy2jGkGWkgfbVzpAgaL8ccCxV
qYvjUKvcDJ2gd4T1Y8yASJyEYUmZKBKlF7AJrcBrrWIZXVHpAA8Yf65ezwQVKdkDNB/A81rXHPuF
VWTrFpKHbkFAnfZH4XYhyVtZFLuF4j7P1AFFIfS5W9xbP7keXyjAjsjF1M2Vh26e3QGBJSNAhCbj
h+lH+ZLrhSHrHgK5pOgcOmLi8iK+9+PCy4Zmc0pYBej0g7AIcogxUx7rWsLuB6HSHbr+O/v0sQ4I
h0TgnVyzOwrVAhcEt50883k94hqbH6J8ibZhfXylW4IFdQlhMY7Rc5ildVZGyBKHQKlgmi1QCQuR
xu5LuKaFUuiWkBq5mvA+qWgFJE9OUkQea3D1qMunjuYMg5B8ZQUebVSKH2DmOCSVGJR7p1l4lsTa
ubAw4l82SGs300P+BXSXzaOO8Z5FXnhltcErLaikn3fOSVG8035P6gQx5zbt1Rhp9/QQNJsFBYeA
WDvHIGJ/x37fPv3YagnPNcbGcEVfb5oxk8q94rJYWJZb2xCpIvWLyrVhmnccW75Osz6SBYUmnM96
zoYpCkeIlXDfKVXbZ87cwEK59szr2FeEdUuTix49hUAsnzLIStEIUCnWYasVaoNvTdovMvj8FeJI
a9FCWzJgKsm6W9NqaMGngJnLl2dmd1KCFGZpIoY78sj9ZDEYnnY0le1XXaItgv9jo3ws5Ku2emJN
r0J9L1BecFWElzU9jBrT1VUJy6QFnMf/3jLbt9t55CeqWL5+OV7pdyJRjt7ppGMNPx/4MTfLQk0g
YWUIPKKaE3eb1EtDtxgGNSnq7ldTYocWNxXP4kJHPB/zUWONN7PKZvSg7LHbAEV/NMvaswbIKEUo
M6uQ7mbyQ/ER/Kxdl/5svdTDA9VjJwF0ZABKvrnuKaj1RKduVI4RkUfYvaiVTTzGb49RxRscmSzz
yiZSDJVkNAwSJzsRv+BOHjcnibRbrboQ4XhF3WQAbEB+QqHu1owMNi9o3uTae9JCIlshPl+DgVFc
43JVj1ET/9ZlbqtWJYq/qA53nIpbG/N5vr5pu78eLSPbx2rjqumafOGAA6IUZ7KQ/dTmK5iFKF4q
aknOg/L57gsHN6uFbsJSTpTPzVekMBTOefjoLeSSfOK+UdGEldno6n5igU0csy1pFFqBanil3aWc
IHY8Ui4/phFxC9ZJwp/EqSUI5lUaYDJvIb3bBRrqBE8V0CoO7LVPMyvnyuI+7kO3r61n4e1W9+wv
rs0PfDybyH1rvGGfqwknZx4FDMuFmvvnv/Tna8gVpdAZO+KnJgeR2k29oJkm6Cy99xcnVCjqBeS9
Rf1K0qdFIU3N+Tktv5eQRrU2ZDwkNEfVfwxW1TLg/vTCWmbm0ZgGYESV9PRaxk6QMtkUKkMiphyr
RozS1FBATMRIpuJW47XpgK2FHXTUUhL6h1Ozb2tm32FLItx8YkNoVjGY8Kzazfmzug5m7qLZr3SB
NNog3nvM7xqwqmWSpoVkqTBnm5ftnmPbL03Z+z05oiJVC1OD9k3yNE75YvBVCq6EYTC3qsH+/2Lv
Ft7p7BkQ/+OEd8VxaQckHmBTuJTJpBIVkrmsQgAHYqhCFuir3xhYnBEHCh2RW6i5efedH3t6LavV
i2J7+SH3tXpCE217yIIA7E+jinh8JSyVwLT3do5j+wzVu5gD15i1PuW5f5WryCMPytGyV44jTCQc
oYB9ZOjdAXh0s14m1Leoa8GLm5megRaWHDsAbS+TwynEA+U6TfvPmI9vIyMQyUfh2Mgzxy+DOyFp
Q7IQCbjok7CrofoQ3o/YrkT/xdUaM7qbB527iLVvGeR3drAxaErExzBaWhPNdKpLJog2FfDqqgpN
PXNpBGfWKpUsvLoQs8EV8plu87+pm0SutG2SkOruE8lK3eRRfxPzJWg5osUKxZM2lHmcO2ZZWDSp
cdyLvV3tqoPPi//pVOTku1tvgl2VPk3C9uOQMNOV9In4QBYlXvOi9hXM3vl++ncmqTp890jLkpKc
vtiLEC2ROKtnYA6kQA71YQBHqpwnvsHTsMWcGlb2Z1wGcU/aFUqyZSskM0jqPoIq5/kCg/sK1KmZ
TU/LsAQwgt4h7Kq6qKP4S6iW5xbobkhbemwtNrdPPzG9xgK2CUGlUjePdpCEoq5EjWfPC8zfz3YF
aP3afr+pyvznZq1xjDNNcFaBqv+02PYmiT2jN+8hrKf+/NjxXb5YTpWCCpKsQVrBAOz879RNE2gs
4JIJRMTpr3S2KYyDjTcZJ0rfDttm+1URLuMYmQWvTPX7/QIaZaunlbp8dvIpX1Yc+Qb4oWsDcUgo
ndd23rxWtgYIrzBAUezu66Gz/NYv6kJx7MJcBU4j+XZ9IT4xQs7Nc61r67rxGyM7aPNTbwRw120X
q+KT+BWPh3oIAzGXsmo0faljwdgXzxl1or7uAh9IjvrVc9UV22IWdxT2DQK9otaI1M1VteP0hg49
isXHfWuQPMRi7VH5ooNKtRNsJuddrXYfYEmHBxRd6FZ9jq4jptrpnZAMEHbxVQrrmOM3P1Hlweto
I2ed7Gc9Mix1+g4mRuHa+llN8on78p+Fu+upLYYl7+aX2DaupWxw/W+hD/+ud0Exl2dgqSthUeoA
4qwp+1LibvX4tGJ7UYXYwNSysfsijRQY7oxYauxlNJqV2dMO2zk57XVnJVyFVFIkEvfcehyOZpc6
Qceg1PUvQAM5gB6+FfUf1ZWR9XRRO7TJS9dwtu0YLOPdSrEMhsc4uqO1dtkvzn/gpwqetRiwLSIH
GFhyiwvlKvs02FuhnezkXMf091xAgWCVfpDsbYy5Tnqbd4YXt84ce+20Pvs3PA5dO2ajB5nd5pkc
Q6T/o3V2C85hlHfyWhnY2n7okXfERAFfyFTsRRiG0iwAfIfMBhT2HbjvCBgNl5X0x7XA2CFspX7V
8y6M8LsgsGmIzR8L+UVf/WKYnI8h8rA8WJB3UqXP9tYc4xRjH0jKkuQlMejJDCx3YapZLJkUs22S
rHaCKBmWO6b9nZA9IC2xdYAtMft6iRlPhbwOtwLRgdRBL8a8kt61mUH1oZH3N+YXKMStqLFm9n0A
U9OFMpLvrbF7O2v3StYth90jbuHFviZ5ncKqQXO3Kl45BwFoXPtgdOYwM2tQNXellsI+RnqlgEje
s7EZGqDbwlXNI624HRvLj44hRFgCscdV95z2HVNhpCpSIhTi5V9+21w3F4yUUZjQakbNOuqrUpbk
ygov6C2Y55J0oAlv8MK1TI7FloDhtRWcBbQuY9SbvAKC6jfJqoBV8jqCOXiNVSb6fldnXNaVNHul
VrX2r2fLTBhquuHv+RQlkD4SEvqj7E5MjhC+by3YPRtU5hVg3fAdr/FbVZd5lRWAo1LlKmLlJVTn
w01W8D5gjFNu5DwzZrtT4PVFqSsObf0+gjm8mCjzG2e1yTIExGT+oyX8MJbGicZS05AgL5zSmQ3v
cqxyLflHiK8L78kEsmuQBKi0YF3Im1fP+rU9w2MSjR1oxWlFfCkPIKtqAOcgUv6VuvzMKUZ9L7ms
oYgp/HzNaXPpPPddzfnbG8riNCW5SXQwbV8FvCVFKEKx/PyUses5h0zohAEZJwWgcwSsaJqC4N+T
4TkpLt7OnjZ1+EYm2i9T5X/Sp5cKYf/qDACYQZJCYijyY2RdF6fZZzFcw3SOggojBXUFzkeoZSz4
GO9w0EQ19+J9pPck4LH1CDsizW0EXFOiVTCE88VNK1aYBcE557FsnmUrfSZ6KueyuhUIdhcg8ywq
Xb6WLiuCiiilUic7A2EJp8yKgRu9UACzuzqkkdPW156Iln+4tbQWcH4rVVXZ1sYUpWn0x3dCHKaP
3L9DAHnqJ+A4Eq0KCgd0B2z9pR305edA+GSWmA8q0ve5zY2zX/PGtHFNx5wT7hB309E5AV+wv3eP
mX+SihGP7/v4tH0nVJXiJV0DRINJ8WJWdiqzeCfcPYTqK21bSE775RP6NcMVJEKOy5YcLfPw2dWx
2dgwQHiokRWC/pVd/QDcFRWpq8PhaI+dCFWZWszsPmgSONOogbPuW8VTqWgBNbL8aR1pq4GhaW0K
DMx8naloIdsXQNSpK/Ohwn8h3EW5IjqmZsLcaieWF8L42sKujg2Yb5eyLE4oGtNIWxx0tBBjtHw2
ndZisUurXZcaD/4nuZ/LQUL7rBvYXpiNoXKYoNGvcX177vhzTmM6c/lKK312xE9sxZiEg1Ywlekz
UEg43E+mxq5BDDFh1PwtSHdMb1BvJCGvg7m3CKwpLco6h1C8D/MI4V2IsUp95fpFFD0txLerGoId
qwwzVQ79gvS9ZIH6CxASqb4OvgbyqxbtmcZc+MArpCuau9e2o7pz0uMcy1mIK6/IR5N+iZhxSX++
Q2PMOlg0ooEl/UDJFWxglJrF29hPGoAQ6EWBBw+YH59QNowp95wWORDXzVHtM+HRGojBoFDK7OQo
CYJPIitY13WkTpUv/+ryKVRJtxP3Ut6a7TehqXelc3mThnZKTlWcJml58htS4/YHynwZzA8nRbkl
7OzymMk16O4kc8z61zd79O34SPvw7WLIu+wedfdQUS4egMP2WVPk5BQh7uhb716bJWLNmNHTFIA+
Pc7smvjRWvVJY1c1CEPk4+Tjn5/+aYiVkqZsCjF489TRZEhC/SnsM86AqeiJtAXQDj+peF0QVlHL
/deteXOaNCQMjoBTGuIivwSWvro0yemM2cpHJHFQpUabN0tdoVBstl8tQHNgqGGz/aKzJjpo86A1
K8i7wJxPx+nQhGP6q1DJobLe2V6mIxi+WZ0PRLmrVNCKPSu61b/qLojSXADBzqFKodIgBmp1IOgW
Ap4h/ebMwcFhVuyiV/+g2nwUXTVV5UACMeMBvHdtFOXbuHQlR2nClYKD0YSRxcfdMAiBLvTNBtGA
k6BdrPpLsZwhL6yiBtQphCqi6jWGTkLIYax1qtaEHXwbTA4vE1+TjPIIBWHqzvpI6cZs4bTtH98J
9KKmkfhOiHd5Ozjamf1ZYD0hn/xO3BXu7X3Xinqy3beoTMFAH+oBSwHppe7DbHpxQEb7iJTAdDn5
0J2Es/XpuJhQFBIJQg8aXzv0vY+Q/D5g7Ok4M8iB/oYLBRPzOa/GPMnIx7KyYgXrzHYYtY42HG/E
1TxZKyDevxFj2HvUSavw972fEo3MKZoTBZ+OETn40veqRZ4QVCF9FnYBBoqt5NljpP81izX4Ei6B
+IRCzjs1PKHLYKiQH5B2exeuv/Q6v627Ew0lc6VrRgmxZuVICyB9FpDPOqLH60BrX3Qy9X/rPhjn
0YFzABplrt8RTpHBsJO8HIcXVeePZVCHECkhNz4BgIpMmA37XlFVo1immK09T99UBdMB3yacDmhK
0icAMLfPbcGJ3UAEXbRRT3szd9ja1sbNhCvYyvbk8t8T+eDKjEG1f0C5o1ndPbYCRUZC5TP6wuzE
EVa96giBP46tIW02ol8/4IeG69MP1DBq0deCPzf4qt0ARBgJ0mtcoZ5uMV4x9zBenEOJzHCZ2f6R
8m+7abWfO79OVZ39K66idcWkLXdiP646N7lg8CZm6iRol0f/Tg0mWp+mMsfGLK2tysm0wnzHqclP
GnJYheU8/cHCtBfdEopy+fuykEWUQKzVGndPXV018VvQbrmge/XWsK2kH6LTpiHhQzvN+yEc7XQ0
DmiK9NlhvTK+iYfOJTcfFqAgAA2c8pHelZPWw354Xb0jZ/eLQJ46SNY4atn4Z7HiguHyPFmJ1tEJ
A8rrKEiLC1BJ2e5n9il/EORkejbC9JZRjFfl5YmtypKhwmh27YtFQPhg9SFEX/iJOMBuI7cK5e+8
mejOsTLGADcoke7XMzm7eao1neV6DJdsJrz0tAlpM2X4JTWil4cGzxBlWCblsiLCzou+nuQlKxLx
Uc5OWUC0UcettqOYBMSYFcoV4ZbDrhYKvArNGhUXQ19soZAtmQNpsgsXRKaaKn5L2yKuZ7IfUUf8
RzOpEXGDCtBgzP+JnRFuZn3P8WEffsGHTC6dxNsZ0uVhssd+cj7Q0b1li8OLXSAzyZQHYz7NthDB
r3YllH4WjJQAWVo2L5zL5HE5v0OnCmzsTObh16PNKYVUhW7YP3PTx5wNqI6xH+VX750Suur5du2B
5FEeStBkxVAYXVYaoQjXAZhHYwelxtkQqjCpZ0pVxSwqJOXCSszbX+61aj6xNC1EfSDeQ9Iw0e5H
EUK5BgeXuOfnWdxBGHbYwo67nhHaJpUz50MzYNVHbQDcKyyVPKNRdatKdvk4yb4oblq7XsGi9c3l
tZU3uUFFfqM6xA3HrciamL9cVielVWAP3MzlT/eiyXvv9nNVPzZofwmFchTznep2ERtTphF75d07
FaNbQ68BFGlS0YYYmi0u8e5/klc1Wz1tkNPKmIJfEeDSGlI/rhRXPO4BmkHytPCnufQ6I++L/o4c
9Wr9SEdJqiwSLbj5l2Wvf3da4Fu1sipEMDY3wkma34ElPzflVUwAxaS5idqPGR0t4XxXieVWJ26h
oQ5FQFXN8IGnCgF7lOK9+HR16jwS+LYjPOrUCJNFnCwYDchRVIRf78D8fph/wWb3OMiacprUTmXI
6wq+eWa/QyWNnvshOIiJjbZCP2oLMJAxymsN6dCow0hGzH11++XZsLLAVTNzjoV7/MYqsr9gqPXN
FyfuX4Oh5Z/cZCE66sujqTQVdi79afIrewdVxd1QaecFTsXVDkdMnHfMPwgG9qofLn7S6n/m9q9f
S7Rss5+G9h+jQYUQw49OPDgmli+b6fBQsJmQ5WtUZxqjec6X6OrzOIRfVUVlGafERFw9Kg+v3DHA
3djr3J59Zx37RHUR8CLrd//CSv6DIAlsEcmE93Nyycb/brFV70/rGA9RBpvhUDhVs+kBakKX8xxc
QKE+UhleQ+BQgLPaqrjjKNc+Dw+wxGNw2ric+4e986qivgVYDoacSo3ntJ13ovq6QxMy7zzJil+W
3v8nVI6iZzUYYJma4+y1D4u5BvfAG1+5epth7Y2RlajA6RYUP6y/GGzN7ESAmFlwSWoF1jRyvPnf
dDNAHGXDjtXfJO2BNAL4YAKTQXnUMKjKqlyjgzNRHj14LbQkwqMpeNqXe5ja0WNl7pajteo4IoXF
865MpGkuDUCLSATUWcDMYzjfn+uLpEanXoORASw7+JAfeHQmmGKPgsZSxlTPBbEHaICyyyJlJo4s
o8kaczw14DFIkds/9wKvhPwE1SBCpYv+cLRFFaG+mSt+glb96DFMoowUYedSB5GFznyslRMd+9/U
OUPCPBc1Va1uDbv3Et5M5vL5+FfQGVJ04lyHYmmUnPQGDMM9AeXlUrRFRFZ1xAq2/CYlF0nMj986
hFd6Xxiwsb6MAaOSMFg6rEnyqHQclgyKBTIXjlPhO3mLzOdGPC/lHhfKyGFjq3AyuO6TK80nQBI2
GID9xHHNQGtxMyjtu1wXsBERmW+zyVrRQm83/EEoYqsRdd3VE0BZqU4gkpeiKGXT920ex7xgjG3V
77HaD+C5pA0TkOtocKzr2CgyS/m7Y7fvbBfbsljL8seXXBt3nzkUjXSGUv1TwfshknIq86x9JCPh
nD/IN2mHgU3lBzvfiPCJHKRGepV8aZLT3x54qir50H/Qo2JWxvIQvSs4fIZ5vLmJXBopY2VNnasg
K75+8XNtuwXlSGRMA/onZHHAr5ZafAqhYwaCofAVgb6B12wn9xIphR2pkqyd4lF/n2BwaFvV9K2h
84fbDOgUpNharMhASsO8xHA0uA6SKcq+Sq+zrL5kdPq/JykfxgSknbavjdfqVMR+Sdd5QtBFWB0+
w5LDKtnMYW13jFUTnInISdqp7UgNmY1jLY3oX+NdrIFQAQpA9xjKMZ1Kti4G4JYdwoQGO2yJIs2v
o+Io/P7QQ1WrHxk2lzZ0j0cL6vDGEXpVNQUqJCTdyP5TpTC1MI1U2NlsfkxS78HrdvwV3EdCTIYp
FwCiXlqFik411FaBcgS0h443gT3MyvWTy/Sc0ZRk8nFBuILD9Ps9LuziglyqoBBBcrQoXmYq4bNf
gz5O1TfT/Xbqe6DKBQcQgbPT35qMFMpi8MeA9hZRWWW7KL3pzW7SvWyCgT5e1+o8xTNjqLkYm+3f
dFd8b6KRgJ33RraLwcBpg+htlmlr50lZ2Z2e8AoC4p16/QFSQZSpW/dLjJ8mbwLdjvJUPZLaBMHr
z/Q9ExZdS7p6r9SeZQAmmwls+/+AeS/gitekrBEI0W+mB5vWQFC0BXHfEla4oCWbRbt+fJa17T0v
RD5TyrQ1tNo1aUHlulQtIzu/Dq0pVL8QLam2ZHqR4c07ekWgWz3JU5Dq5JwifmXaX3syisbq7dJl
bkTcvW79j57zlOAFlLLsRqEJgBwB7geCVT0QWf49eRE2cvqB1YaDjoXBZvz6rQryh+SoEYtqua3K
h1dJJ7MyWudqrdV0yCQMVO2zWQb2tDbXgIj48XM0zKAgpsP/UvpYd0gtOT4n4FwyQxp9o57lN1pe
xlj7As7b6q4ZLMb1B+vcBwoxeUKpTZUafa+z3oHijM3ukQ8R2f9NwMpZb8bB93STiJiKMCzgkcVG
xvKNrR5Mvf2+jcE8pnGzC54cLQdcgSuV2yffurAdCD4pqaZPGm2+FNTQqxGnHTH5/MZhdjr4KDYR
xIhTWacMSGCnFudXLZ9qe/d40OIcrJLXnPOSiSQaid6LpthRdc7TjGgZr44Q7qJZg6lIQczXuTkz
kjDWe2qJ9CY6aoOXN3DTp3uR9unyeZ4eOcggQmRdIMIchJdKfcVq1sNqwx+IgZ4m3bUyXDzfS7ZJ
soBYZkhDYs7yKrK4GR1lXLJ8oqjMjqhWZkPGptTgEwaQHS/pncfgazNINYGzWvutySqkSUmO7zEn
XiPUkBouV54Uz5bNMRR1KywZDhSBYp3i7umsNCSgu5+N3F/nJfIGtGj5QhW9dImMJftf48t1eAXb
ETght5celY+hOyR8IS9sc2gDKYlbbNxUNih4YSAYgTHWbD6XP+N4k7XbQM9VT4VOSd7R9NXjC4/L
tt7fM+TXhggsvqAZgFpgQ/bk6+m0udKRmCMu061nj65T5J4RHw/E69OqwsIu8m1/rn9vIXHKM/BR
JaMaQOzlKb3/4ZYEqTofCJUySj8qhbQiY3vHxkLF+GYZgTzneey3zfrHj/PHgKhG09/5/oK82LoX
4wiTTvXOPUtJwd+zatCzJzmGJSy4s18PKa+X2JhkpEq0q7KT0ueuUsMGB3HCIGVk/326s221XQ9R
t1eV12pZFHJsSR2VLgq7jx8GPKv0ae7Yhx1DziYAMxNsxzQRa5mM31Cd5/lZEjSyynPUi/EKg6Us
RR1cT3A52h4A6wxix6qmWaCVNLFowUG0L0cS6tXUIruLyxBI3KwLYN3VufRyGL6USLQzy1zb5QEx
zFNCEsJq8SbjV520XeeNlROhSReCFXrQ8PZncOboFR3ds7+N8CwSkwlN5ET6p0jtByuXeMG8keO8
DJgxuvdvMEgcwMwxt+fKmlVBYMJanI7UBb884ohwusgBiGI9+yZCypegu/IXjGPxhwRfGaShZzZK
FROKaaVUc6+1dTZCs+hFIZTvkKs0laA6XdMmXeJ2xvHAW80NlH+9ZNTdVXmZfTrzyKBjPRJx9DJX
STWO5LwkUL/gLZkgt4yycukGLkpu2aS3/wwBdFzQje6Vjkl1dKz+lZ/X12leN5wLqNIXzgps87Vj
ghqajgJwonWT6ob9V1QqOwGYgH5/MPtQseHeFNGnJKEcyYMqbLG+Gj/EtRDoSgAH2TPzU2BMBFPI
lWcebWnntRQKZA9RCu+IDSnJHcXpA+MeFLmZ0jbdkHhMYSDpLgzXtroEBUAlg93BqBnNxg539Zcj
KYhanpnOZdvCc66tPiW0YSO91SacNsHHu44Oxqp+IOeNFW+aA/Sa9LSS/H2o7Vk0lUO27N8SUcnv
QIWen2X1pT1tTtAjXwyuU7guvUhfBqmDwoC87WTeuO9OsbkqWgVyZTUZdBFkLK49j0q38BjzPFbr
Ok39O6czWHL0T9YwEMOv/CU94FQsmcqoTuZX4pdpzlOzrpu5fJA62kEtc3Y8kcN9Z0QYJWfrN2++
XR6kLmzx3sQBFvZYFFTzZqrTftN/zjjMdYPGtntg2iahkghrhPGNeQurn7LCBu0/bIDyDL1R2RYZ
nz+Q31xKdJiWu29R2xTA3DpciFwKtVw6v7/oJAd0WFiHZsFHh+WjzsVGkvNkL65iRq18/9sPjL+/
AjpWNE1rfflNFMYqo2QZvtUoHulQ63lO6PWidXFTmSAGOKXCg5ksxl6ngWY5Jt7hAdPZNqtQeyLz
8WiCjqmgV2MEOwz2K0a/PlPnAYSeF4QS5bad8m2fKeEoEf1hmD3j8up23UcG4SuqcCGBnz0ovDTP
fVRKefpniOAnTZESRI8krJrzqQxTZYsVahB6hfD0uISE3JgrV1YxCIVmsDNGj5AMw8W/NwvKPbiq
9k9YGfccXUd0/6YWawGJ5kNJIFiTBclHO8TVJ+edMTxadSUXhaYi0RZflrBxK9MYcY81sYPVuQv/
OmFUGaSf3W1Y9d2uZtZwlvgF+2EYTSTzhzUUnXAMlS8fRWLzYmhneRRE99ytJhG7EEVn/tNlaVYf
3Edah7DuQ6qniSYuKCSOBw6wNRCe4l5XmZ5Q2FUNB9Bu03IBWZAuFONggmRo6qgOc9ajWhR+U8Ba
9mvSJG8wMo4ZufQeqcxm58+faL2ZWhNi7jmL8CLNUGpHx9UGhoIpqOExm/5mZXdLvFocvrALmSm1
HRjbAJj3AxyOJmZTqg9ZNttbRcr0po+QoJiU38k0GSWDZRzTVQmGZlsAZsIwam0StWD1d9D9ueWy
wJmroOh71icFKu6QKXhryhKGIc7F1eg4S4tMn+TRBzV7kiLlY8vsHztnC4mQzMrr6aAxwqyQh+fX
4o34D6Xys0F1rVXVt3f+UHK6FzEp5qqG/lh9xC3DGsg/JPqZbEtniiTQH+eabosVTMlCDJq5EEoz
JB0/N2BxY/+pN4TfMMbKVtWEJRimffD4SEc/yrW6JpYsAaiSa4mUZ5zE9SI8KS/Mujm+TF9Zp5/9
Yvc7qcb8BLAY8JemGNmZutFB2N5BReXzjJ26JJL5eVuMrOqHUBcW5KxisuJ9TCBwKonmvJ/rd5vy
ZHp/mUxso7MfLdXKUhlpd5/nUVd1t3Ydr7eJY/8wQysm6Jk9HSz53fPPILEk+jJVPODL6tN7vYqK
5wbijdVLn/Lvm+BvqypyEy9GsANGGCuKp8iueERKOKPFoWOKr+3cLAJJxy4gAWjI8B40oU7UQWMJ
vaF4hi3ybSfHgUR9+R15P3JzSmyIPksRj4Tmvek8e3VLSpd5h3PP0jlhPKRN3lhpFmT9nQdy1rpk
a1lY5r0KIMhJ1FtyJ5xuy9VewY6HXd6o2cFHCVCRL8UCtremmsDtvfAEK2AQpVljV0xtNhCmroKx
VLgx5oelUNHMGUygKYFMn5DQLaUEq0NiBteK8riLYAItlBlHkIFX7hqd7DiDKXRHVmcjlSnUibqr
PqoUwwkdg789rbNedoep562ypzRfpA0yQ5/HA8QboEb7Zoiz9AQ+tQp6Fqtum/4ba0K7dz61WPbI
OZVmyWptQXzRHm8Wu4ek4ndVm+FTKmRxwmE/2v6yZdeKRKQF/m118enP0bhGvODSopRnMhI1Ry8L
rK8GzrXd4awjHeP1So5ctyAAzjlMVKYxTGRRGrpYPIeQFG+D3nvsVB5ZaQr5xuU9AjfnOIZbsa3H
/gu1UVkl7+RkqXBPPlRCi4R/jKTK/6rlh6ogikQJ9ELgR/YtOEjHftVQP02xUrDxKK3N0DibgiN3
FTH79295Whl8PWF1TmR/Oh3xCdV82vAyijuXvrxXV2NRv8vZvvbZLOI8lE5BtvibwcVqssn9XUr9
d5Rb2rVTJfWwszwj+hzy8byljhor7qggEuYSAW8BiNh8KhnkaIK/uDaQEHQV3gv3F/U4z612LW2D
RciaA2Pk+AGaaGCysWxwKa19amPravjR+WEZHb1qa7+ypiY/e4y6MJmIlQCpu99WPylnzN9STwO2
Ltu2YFSe32OJa5LPc7PhTWwo7nXxNx78nY4eo2M2teVGoIZDbcmYAdUNa9rtMOA+eDZZsdA88cWW
zzsrDUv7tWcH0P9wb0xEorULZZkzVhT7IZ3PBegirIA3Q2jT9TDUJreHiyqN+Vnha9Cbr6Qe2185
B7yISj+zqkQ7D3g/4Q/bmTM5WXy9UWOaCfw49vXMvPCn7pntXmTGUSys1RTMsX9++yHsbga9Gbmh
IR9CFx9gWTRXgYYJ/NqIdEC4wsQKCZrtsWqSXBqCpOZJiDEctOVNS8JavxTc5jQLKAp/N1smOJIP
mRphhny+g/WoqzJt1zIzKcBBBb3TUFoYd7uyaW5yrDwm/j4HZb4ndxxInAbkDG48Q0rgtYCymaZn
3Wx0ySZe/IowU8qZvfs5q3mCynYs7yI5mejbTWTj9pBw9O/yjEVMiMCecs/+KsJcZcUBiRDrFKqG
oPExEmdTgoP7SlN0SzeETfEFeqh9rEFfdTxtvqAUpfGopFhR9IXJcuXzfF31pkjCo69NBo8aX8zj
4/QYMrKN3LGfe+uCORvU8FY2Ueo3su6jH5CXJSxPzgvrhGfchRUpdpjlmZZVXR+waLSWAAQH1pM8
mRYkKxK5jwK6jhBSHp8FgqqkxrtfJ+LiOha5wvqzkMd0A+HCavvC5zRX9VNSKkDfNulYT5zwgIvZ
tQ4qMqyF0PVY+O6VuJFu2j3qTIt+PLqdhng8AFor65ovXHP6TLziBJZmVqFY5dkO1v3tACoGjKJJ
uR/YbdjesnGQEDVFPd7AwK2dzXVXp7mGmBoieym1R3CN9hYB3TqbWwWDpvTcc7/fU9Ap+Ma/ENQJ
A3VRrTF8342tuuKt8PKwdpLJ3DatabF5+Sl/O5SirKY+Jcif1paQZ/TbIyjeFBIdtw4rx9LSWKri
3D+1m2ar6zUq3QeunkTNLuqNql0nhCkJ23XjFeQNRFsS4Z+gpbSVHnDDB34slsRSWAtHCfMPeOlk
g1MqwtxIwyWqt0mJ4nYD+say21NYDzZLkQE3vouvq13x7yEnZq66rGRhdaveQbFqko6GyhyAt8BA
LgTWB4nz+U9sK85xFUzHs/QqoXfXlyI6ElzKVNNJd/jdHOlEl79ofdLlyg8q1K0+BbE1CKdnd0Ne
08QMuPd8g25pjHfiYwyj38gpY8DHS4e+D5ZyCANvN9uf9eWHMnULfvc24aThr5Fe4mhSwuIwZ4U/
DOUi9/0wvWdYnCce3pHvCIkUI2EcfEs4icx/JNQZsehz3ffSVh3TRvKzz2Sq/nBxH7ObtQsBHHR3
2A5PV8O+qMgWuN/CyERWZqwgVbkwIWgN3JfP2fDYwj1cbgiKXxun82123+gtjwIXJYeVmqydw+Y4
G7UqCi/Xr+khzUICym/Q2ihL49h1GfhOHCzy6/J4bbgaUPtE9EYgsV7+SKELhy58Y+qsm5PafFvA
pcEM2pjGBQqS60g69ejZ52cvS1n5hUZznVBrWMcYWQLWXJrRduFz+4AvwFllLme8tb39E+95e98q
S7jOETxifCG+dYKCAswQwTTpcWmK3V3oQURZO9bmGWNtQ6viWL1ETlnWebeE/+gVpXrp9X6MSR2p
1KMNJCzDhZ98jdQNRrhnOgVg/caX1uuukmvK5PKWRHq9yxmBtfJ+a83gGwv2WRpM6dC+wPcbPJ7g
GIx3W243rzj34OH6lKnInQf2OHeMsSS7A0M38buo2OsQw2cBOVjItaYABz0BzlszGtNGt3KKU51T
cw4h/RxYeI+VTZwlA4OP0eeyRAr2qaX7ncgITjLduSPWNYROCLeTDLdh96Mryi1FiB12XKuuBoMH
8+FFJiytOt8S+PfOGlFNWRLVRzEiNIDIR5UemaT3Im/QKwKKji/4lIykC9Rfxf0COovGtX9IPHpi
KRY+DJwmat0x29DYvHh2OJMzpFAbJoxQ3gxxOAdq8FZtbXdMlGBpm1FlT5OBbYaARO1g2P/8xE5v
mxld0VL3wY7AACsGy3XOFvbOGlInawMYcDeg2g263eGwr4zmCNumWl/ZNDnEDm3Kjagqgnbr61Dj
+7SjPHh/pA1I13S8i+ee5NsW6ca0sGCQAIkZCn+8DhJRBc/0kYejUXvNddbxOBJiqH/sftoYZaFf
BvH/tB2U+TqIbbpoD7ZQmiO6+w1A2E10CRRTRGF7DYNrSYH+79CJtsnqqA2oI7EqdYi5bsRFYkB5
7WWPLgSx8hG3Jpm2GYm7QerHQNMKa5b872F31dxHLSnTyGYH10k7MFgxB8Po4Tju8ZBYe+D7HodD
RtcoGTdiPGtURLjDuGpT9nANT9lXlIokaGhYiTXJXJ9lvh+/yLWkKL+Tv2yGp59ZX/nQpteQoZmZ
7sGsqd9pybdmS/9EnNM6xSOO3HPMCdEifLiqI7dn94uiH/zIuWiXNEkyMQOi3X+x+BFIHxUtSuru
xlXi1fwDe5zZUSZgLnr64SU08wr98KCYaTzqx91CEfzyF1Ms0cq2go1CoOG+0PAE8JjSRBgl+luc
4aXrEsDTk96Ex7RPpTuokpFXetMllmD6XD4gRGJ0Ut8dMJUJwCTObHfH26G16zF4e2nREnWzJlMg
kJNi3Qb0wSoQNob4Lwm60vtOkf8e/IXfZ+fYO4/260Dplo7STZMFgjUILJwz9Cc5GjuS8XMv2SZ5
hQ4EnmqOJKNTbMCMzkprb9MobB/dkIuK7C4fFJiVwwZ/6btDBTS9q9LZ+7in//TF2M8RfUDV6Uak
aQ2qRBlLxpLeHTy7fyqzg6HnpLUA6pXvutaXHMgq7TYWOQT97dJcYelZKYaNzwQSeE9K3p4axJo4
1zkNIBvsyny1XyVyv/Y7DgVHADLjzcGW0vhstINWHsO1lANLZ6YmvvtpSHaztrITAr5dby+flx+W
M81TpSb3+2kA1hu8njsiiUGJdoZttoIyGRkXRuFk7bzuNwY/bTkhkDoeJ+EeaUvjRU6iVM+SfktF
eYmE8d5w/nrUHCoQlfPtgkwcwMOZrnhpTU9t7t7y0eDgx1i/R0vs8zKmmMPtWMAzGZTb307imAhH
aZPHljxyz7k3f5cgA7PyqkHRRAcimnz8aleZHK/Im/h62cBAveIz+M0XyMIMdiK9ml/Ij56f9TYE
G2hgpm+wqHRph4msIznsyLMSvUG96+a7AWFJ0/dSSgdHP3xZHFmkxPVXayQK093NUdPaLMUYZWTJ
cxF/siOw9Wb2m28G1Z7/+9cCuVxCmMmVvL0j8UVSz51k38IaIudiAWXo3G+C21m3rUwEPsKoaX8z
rXYOX3zPevlvlHJFb08PWMKNkP/tf4M/vjjJ9K63zbjieySHo+sQ0qSmYgI+SKjXP82FBWfIi2xV
k9PfGXY0JZYGGrPidlFNLbbk3zSE4QVvjdIGBAw3Dn9qQDVuuIpwBZ19SeBpdI5N/o4a50UXgW1v
w+BPLXdMRmWdJoWJv8+foR+s0X4DSWPFKtwDBAbAO2cyD17I4BR1xV3TJrQ83gRj6Kx5XWBWlFfA
ePk34/4RuPZfyLYRR7zoLa2gIdj9bsPlSh7UUJLBV5FPyT9AXWNHN2skjZkiKPrLkInBs/UKgxl2
QCKvpaJD0VPL8yMAza7zc7j+oI091hvhuExGt8lSDR9ovR8Q9b3KnPFhpZyuQcFg9CDrT9+M0lSq
f/PzY0P4OFHPdsHP6kRO5+m/87Xvmxt2sOI9EK30YFZAMj1DCBGN5LI7JBGTMGVNp/TO02RYtt96
IK2ESclzqeyJohXooztd1kW6uiUB0LrUd06j2Nq4i6+Z4M95kcyNL4Ia1Bt2cCmVGjJg76zaTBKF
3PIxQG6bF7CZeNf5gzGKiDn64lht4a78cmZj1H7OA83+JLIsU6j5wEm225VzS2PsQGCDvkmaqQfc
Hfq4VA1PxMdaJssgmNFcxRmfXsqKhnPmEIdYG5Jy+viLPTgtaxPET2RSPrpmTFeTc6jZx8R4Tgly
TGVGKgt0M2q4ENSccdOJlpvPW15L3333VwTxG7SpFnvNWTBFnvUYwTU/Ua7uYUCWZ8D2e25oVZTM
RQLDA6zu7CUb7yFakVQX1HaKRUkwKaTgrJsOvfzcdL/6nTAuVLshB4AwXe7VY/ScdP/jaU2Mf04+
WZYt1Q1iuR93myMzQLeWedT97ZHjjxyKuXFGqFs82SA50pKlk+iQf2rxmvNFXPtBsjYYmqaMJN1S
tMNl3TiT76zkI1WkS5hIkcexTlmoH0iDgm+7jKtWI5T4O9+eKoqPYcrGJfbG0DhPliKTcCs865AZ
Su30WRKPFcQ2EOVg330G859E9UTDMgSIhxdQgSJpdBSvVUiQUrz3XHEwirXeqSAGWmxaVtVMWfdf
r9ZbUh+xHz3yaNiNCe68Az3Y+1a4A/EHTtdQiGQtjhEus2AjfMkjPDBQSGI70/wO3jDwtwxbvrGA
/+C0+8uVIXNVrcY7vY93Owdtp5BTqoEqUVc+Afgt5nk3PM0KTmh1KUSxIlgJwn++mwimHQVAst21
+DAGrp963v7zgjpZQpnUZumKTpG2Q/i8B9Qm+CkFx/r3ubuygzIt5zgMYjg1b7M6plhSAr+MbDou
yIWu6hw2iCHNdZpMbsdFo+crkfg/hLT62Y89E08g/RFqTkQV5l6R7wsf25jBls0SGVY7TFUZ64KJ
LD4KMI8helRYwVSFcR+s0M5Ls7lh8mRCimnb6zx8A5j2HN42qmVRKznOT7war8ocmudZh9A05seG
eWn7HK1n8Q+rcheosJbZgonYI++KzXuxWvwCzLEaKpxBa3PkqNUwd7ePrHOlaKPIACZ7XnPER3+F
2tMqTqNViKP9jnw7HC3vXByPD2flOtwCDRaoy54xDubnmvFe/eWWq6pYrfzShnaaarf7egL0oUVM
vqTTW7OqGFDF2AF3TV3t7i3w8SAvnHaeLH2ZwlkGaEgECXP8vASbn/pG/P+XAoFr+jAbgPvLNGYL
cbLOUpDtkqtk9E29Q14W+PHaxzj0JCt79ErDotHT7cWCZh6ic5ye7dDzMlHLw+06+Qk/1qJNuiUB
42y6q+aq69yMO9LBlOhp9Fabz4d2BzOGxFkCmVKeRfSTi5uKdSZ8GtWWrHjvxBQeY4hruC79bYzP
qi5E8ZG9L7BEZWb4vUJht070h2ihL8cmoW9DqJbW9kW5eF9YaWyhO1Dbk8lFynviL9oU3j0T+u2d
NteiSp8Ezen925jHpAGcczNhTrCTHb5pzC6lDc6FLY9cRoLA4qYoUxXsCUnbm+eys+pSSOSZ2uHf
87GHZSpAM5vZuQpB4lUJfKdVGcfHVSyK5UFMvYh2m1ekvAr7YuChvYrOb3VXE8PJEeIoe39sJ/Ok
ExftNNv2WWTZnCPZldbQLK14zmk2PMTLRSivw1SOmxv9OX6zddx6CTxbE+GGisxkoYLS/evuLY5u
jG1B3JHwS1JhKq6ZcmAjPHUCI5VMFb4An+Zt7ac4Y21tAXyPfmQZ1B7ELsn7Kog6eoZ/lZEq7PXy
6/5o+FO/Fglb/2lXHPXs5Gn3HpMkYVTlhxAYp8ndJ1Q43B72Wf38Dg0ZAJuTa3Y/huWFkcUSKGZX
rsefUXhU2jGIYitSl13cmekJIZ3d0qQytKLKd8eCRs9SB5Y/4TwZ31YUKzLFLysTxke2Qbh4xKPT
P1WCU2KCyyoqDmG0t3e8lfssWMmjxytPO/Zee4cjUQR7Mu6Zx8y7hUFxqDFqJzko4RMnepYAeMF6
WcPNuPVacIbtM+nmHWniAx1XVkyFat32UuMrm/UHEgx4h16KYjCM4e1lE5TOeDRGKQf0Vmzilyal
tspL2mAtPneltlSHKMDdY26r66cAklXEtS8SGIhTORfamu1MFJOlWYNdpruTGqquBiriqQtjlMtV
W1i7LPVIQ09GEcJSIDi7gGxmt7yOLs2YvMmsGZUb8VbmCBGA/MrxuvC4x7RYhFDHOcI2i3YG3o71
U0gxJEJcnZyfeDoutXICTY+ZV5pVHDQX0qM20emMfvBtFHn/LjN5cpwuwm+dNXwaniURpgacYsS/
wOwDLj+Hlq8l+OhOuh2sG2jETcSe9VNZW28j36aPqwIWcNvej2AK2Ay6CjNZ4OzzjyzcSsi//9KI
Rkuwqolwm5PCFWynS7jb2OfaqB3gvL1Y08vfiP4uRiBxiX2m0SuY+V8xUPNWiMtwlDJ0aksXrIKf
ET6vvnW0VFJ8SAkSNZiuo4+SGQRLhcnSkPoTJh4GDPv69mBksdxby1fKZN4RpNW1Iq59+fxXJ/9Z
0A9hRPJYYNoy/4SG+FxgoX7pKtpe/EMFj6I4SrGTuwl5x9IaNMYOmNwWmZaIz0rIoR1p8AIP/+cO
Yf7crEPna0oV8eejQt8vutK10QqNJ90mEyC1KyY7cgD0UHBoNmOWF1XmONLL8AKMiEhys08cXBrP
UDDbh5ekPBl/C5XdUPmg/fB7qeR56ylcUgazU/ZbeNSsrDFxvrvhmKg7EZ/wLhsWvX0BPoQ3sE/r
xA5k/9d2LkVEsXHaStUhw6YfrmpcFy09PfLMex/1xlUHmCmZclZaRwnf1BFWEt1zSkcsjGZIjA7q
pcdFCWtiEb3qZcwL9KSu2Bbf4Vmi8QExss0eh1+rx83xF56+qB+U3XmSIRnpuHbPouHqNklAhn6j
BuREaJhj0TlghVv/TLS7NErleXJIsOb+zKi7B714YXP83DQuoB/CUp0Kzz27cTrIM1nwvDmy21yU
0mIR8tIHe6kPDSUt0/+N99PGOLDxHhI6FpMsET0dJKfpONrprBdnr5PXaK3TWaAteHORVYPSyZos
DaTrBBnYiLdXIJw0mFu8RgCed74n4izwrZROpgVy0PKCqpeCJW5jbTP7+3jRjLp6RtFyQnOIEzmI
796NCPR9wc4hLqeJdxABA0GWqU+tOW7CioKv9/gwY7GmBkUjOEDPHwR/YDwqJkfekZxUouHf8Zoz
6EVq39Cx9FfyQpurxd4IdH9LMD0r/GznWWnU22sqotXa46s+Q9G6YPQgOLeeby1RWiGr7geIqOXD
r/KVF6tBTSklmSJq3ABJ+YIIMNgoL5k9wT/ltqIFRVhS7Nuo13ss2czcXRL3rBmFcKrMZDZykZR5
6IXGAmYCPVXnNic043y5YpcETlPmAAwdp3IyB8Vt+7CsQyrIBA3D5SK0CLWzcCnGI4wZKZ6Tt/wq
a44X1zP7Vc97yYOxM9ov8f1Udk9ANSBcVDoxXPQwpfHcz94t4EDciVZ7KXGN4NCX+P7Od/o31Hex
h+j/xsFsInMC31R9L6gHdDHndoVJ4VtR+8oJTHFesKDlJxxSAy5nrZ5a77XKLfHTRcWesxnjv0XE
kyq481vURYFjBEptk5eegiB6elwdAmuU9b5XKwXC053af5ly/d7li0G5TvHR7wIyc4aJHujLMhHg
Zs4xeM86nCCP1ZTUby31v/FpNB32VE1oIQEBE7XL6rXu8sqtQtKpIhj6TVmxF5fimPY1JH2dSrel
eSTK/FitC2rGwh3rEtxAjrHmOO7k2fB/wTp18zWMnK/+Aqa8rhjkDUBoyrTXYQb63AcerwpeGx3y
T7zgmayxUrxqYLBmsHjYnMUJ+noWCM7C53Ns0lcN7zVymynEqRh1f6EQJLUPdy03JbgjJYZRPtkm
TXiXHSxRo+3EEup2VbPAhOyE+CQCALwvpfpKc2H2PaCJwDD9HuilXs8W/wLyaHPKZLetzI9xUFJI
5DDMdGBesw2Dd0Lojjv3lFMrOrGlspUm55YmNWXzbDmww+DxfR6y8SVrPVCwbsVXD2QYuEoCG3Z1
FbJCALg20k3rGsVggvarCq54Ugx5jwo7eoSRxAGiI17M+jl0RR1n5Bpao1HXiSGrpgCjrOWBz6l7
J6x5YL174atqJMBapd5Zy+Ug6QnuhkJ1uWT7qfjKzM6JssIglTOtLDcuHIwrsa8yAeXgqcYmLa4j
RGuhsGcoJJ/O3QlH0PEpQkaCzRxbAkTiGXyNZh9IrO7d3YJtr6vMn/vIpSIGSC8pVIxuHaffemHU
BOzodKL/hhjzhw+u765YtI9ALEvjPyGbhWj8Q9q6fxk7J26TzMTBsgF2GJ9FNFH1rwFdSQnoaXEF
1Dzy6m3z/l/qCoeIdpMnBqUFJyoMycwDl4EBuz+ObppPpnEmOIAcHZvpPKsW/8Aw7TbYtHLMzhvB
wMH5OixMyWsosMiebIACLpDqRrqlqMrj+4eNCgPrOGwVxi5BmGTMcT+rFMIB6P4qSLXHCBg585+a
rn/W+Gj9vfsD/CTeQOOgHlmuPVI4dSJW/dIlKjZDjfIPZCjyTk/GYjFkrlEHhh0PwwypBdfKKPaM
NrdN28bE3iHLXRjeEitStzV7IOcQTYdGWXhS8/jGIX9ThbtEwFi9DxSzOn+t0Juog2pvMwF1v8/9
qfuiA6i5x16BhXkGxNYqPFG6IJtWIlmBTVOK8QlQee7dl79pLn0tK+2oCd9lSIBhawy3rlkKOfEq
vdongwCu+aVJKfJ68jjaxrg+G5YkHpBcJgRPQW57xa9h0DDx1gfiuV1NwVt4bQZQMeNz5QZmsqui
lGH/wldp0A2RyAsO1pdnd+PcXwzAz6+HJh6hSqLkSnDCLJk13B7RvyPAQqXEdXmFM7MbazNEdjUP
FgfdDHgeRWvbjlwcVz1fWH4ce5bjK2S2saNAEFqSGxQ2m7UvijFc/lCxxylwjm56Ec3QcPXO0B4u
rx21GlrmdCEgUlVPoprMXwdukFCKhdH0USMEhiGrA5Q+1pgzwAKi3O4JquHo+xaneUd3Zrrtjhuo
IGigb+jrEyRFyQTTjPJdabuXWIlAIyXgvpbLWzwwskfUWJdomyw6jdBihAn3Mu+yncuZ+Jciw5TH
hKHpzqc9fJznKt/BipQ5uhkRDXkxdaHx2gi8iwp3qyQeMC9m8Y4UZRQlZ420pl6ts+BQFv+lCDYQ
8J56aBocwY0rLGOv6BPYXCrChxWNUqTcJlYusWxx1foQ6Bq1RvMWaQur4gkd68iQm562Vg8KvW4I
ti8ckRVOCmAnt8O/2m8Y7R1wGewsh6D3CrP0PYdc0hyoI9uK4e+LI8MpXr3bXTQwGjvVqQAX7Ou2
lSmdIOk0Jkb4cv9gfjw2lme+f4tSIveijoFV/L9SyqxGSsnIMKDDxLepKkgOcWl5I7NDy+0KbdCR
ohulzHUxZSDKiyRhIfttY1vbqrAaPqfJw8ZTvO8aCutSmn5Jfw2SJ5n08Npbdg3uPGqavm0KX+s0
mINZ6nSb/tYS3BAWPTwAN/FOxbtQv7yXtT8WY6b4hepHieBUqu3etfwJbwodwdPOUpDW8DQYi2yM
KATOS++vnoTz/tlg/rMsfeXON7JfITOrGM5LjF5Ehh3clCCPuhtQUFxVpjpAjw1zCWc+uBeGTkXe
cUx7k9ElAmi1ve7gVIMzqnaLOtAxD7NKxK6bjqfrqaI1NO/BePDwnBTKxCkzVu/bxLtHmM8HbTvG
5DZxH8gxzj7VzPzWgZrC6Pdh2cqdH5vUbsybLMAqKp1wvi7bSMroPkaxPKJIkB/1zOFC6i/ozGD9
FwPT1iZWyzL2j88JqQmEmFpbCy45aPK1xs+X9G1j4U4YPMV1m5UpvrVNivodaBEns1QPMcxH/cB/
A1Qy+1xlUT1xt2poTYq30oOj5HBJZP+KCp9OLwJmeGPURVVU2k56Lfmc7udVLNy83NtyWiLGqqkZ
mmlcX5UaUkiRsp56ytZZxEdXPF65cYT/DI5+xq9hDRFgkDOAbOuT6gp6Os58zporQ78uzo35wLO1
oKgv/f5awsp8w110t8k32GqdPEzHuxwYcyrkyfR5NFOobfhrUQ2y/HqqQoqp5eVrfBvu02eNxCOy
QqHsWgxVqRB/9AJKuoGS6K/qdNrrqTjqd8EIXp2KRRifkgXDHpAjlN2LIHj8LcMXFnfqAhNYgnl3
Ez5MUs2rPwU+MyKhzOjkNWp7IJCCkYh756DGt/2eE8SgeeHPV1VgksbqkAgxJE+bWxdGGw/2oCJP
UAaDueRmuhliuOjbe9QzRLYtQX3PsxuZ2TyaamZdsjj9XfBSa7Zt3Es8WQMREe6oAbc5ivSmnWZR
dDAUheoy2WSdHxCgKeAaYm/13ssvn4oxHvjm8h0cir+3AZbBnU7iQ9wAjuWaK4BnTv7r7W0k7LR2
ZZKRZ20Ms5N/LyAyYRTKxW8zvggBiIXdNhxupOKctmQix1e+S9Y2twCUxs/yrK8k/4fc9XqccjxC
VGTqTLQFdZbcPiZUWmZOzTkkWuAKJHDZOpfEP9vs1uUHaEjMUp8tVUMN6dYc3A4f4lh4n6TJX9eo
grKJkNQsqjGL2ag3TKkc/YBq96NzXb2mVpY9Ik24ebFZLJVoh0lKQ5kuND01GHPJ1pknt9pjIRno
pIDoe7CAERFm4OAWMJEBdDSo9IuUTKJMctNJYUIy9LOnLpky4e8LtEWlC1VNNumxUvl024j+Zuih
myAIeJ3mmodrIBYA23H72ASFjciVvhIzRH8AO8JkC7I+ok0ekqRTTynDIIjj79n1ROYhkvQO3yfx
BqXjcyscyeVTFguZNtT3AV2bP8nWceP7Ny+2O1tRbULDmGAYKaeBWwHx03l7xHRo9seRdi69VToN
H/06MttL7+av1TfTiF0b6o3mPfNmKibdrFYZKWEpQQgiM9pawu9iwp+Dm1A1rW8IsPr4fKEUjvtd
P28owBHSV4kQzVZXGD81H4GpwCwI9m8fIVLsTAkFsU49Eo3vM6cT1uzsI16LuEdxbqz7E9pZe9wK
94zcc+kcYLXXox446mKhJUfFeTfYvZ4jzjGQpWC68CRK3qOwBJ6/BoEZnWe0yhqabpn/esLXATa9
Bdks/GkS0M0izam+bput0f9kn+hNJYBB6ojZIIKcwR1EwQMgvrQ08SV6i5vnScquhul/Prj2NMW0
C2x4T5DrOqijh0/fTNavdJgS2LaYdydUxjtCtLdTsZiP5Qrf9P/IuX6CTJKe8RBVOrzjBe+JAaM/
Ldd81v5w0SN5E27tWOw3M8BZwNgygBn5TklMjg7ttMNCc/wPjCdBm3FICuOx5+le/KQ3d9vr0mXD
+wx/oLLkz5HmEl5q9KgZieGZo6f/vEx98PNX/oJnVcUYD+gBf4AReHY7fD2KsStKGr0kD/rftFm4
KRarweWv8d7tqshhXzvGWfK1Gh6/aTyra7p0HjLZX5hopOWGfHuuVzTOBKE222Be1XSs261z7bnA
UFwJdQzBszJxYQ+Of0uvvu2W0siQDpELjA/Mwt24tN0dYM/6PT/Zx3+a1ApYt8TcqXqFzS6DO3ER
V8GjoUX+tMGHXvLoVofwglcesdfNHMX8cii0tSrXq7Azam8Gb7dIozIhQAV7NkqVLEtrV2X1hWry
BUqSBRDbT7EqQWUrlQyb2pXCW/iwjhRKwKRmws/MbUppzNj5cE2PMwYwLi4tqEx5V7DK4TGwDhDa
fa2CTHxGEtQlbkvrmXTRJaypZaiyG7vSQxe6SsN/7Q/d94qswnzVh8adO3bPlTORvZtQu/ifhH8L
XRWQmyT7R3Av+W3qEYToBpkBHeA+Kel6PzyVQ579U8AGwQYJQp+LVelJz+gRnu06vjjUslP2rnDS
6OYnTkkiOdu7dw0KmjvqnqTIU3dsD1+MTtw+FFAB927eW0woJE334WkI15vdAO/pwHKvKfPAzGiG
EFucZQ6iO63BxfqVagImzdFFUBUspjT2FD44nU3ICJBos24NPAJwENlACt3lAquAQ2LHwwpJdDMq
z8eTRgpvMynVt3ZYFma0cQwjGERDQWqipWSi4zl1fj1L0kQP12WCxfI9dSfi0LTWwsda/FJ7HFB7
w5o5/+fmaFklv5gZG/10wvZWAaeMdGXn2H1w4iP6nwYovIYY8gwMPjQY57kKcW+OVxrnxT4y/SYH
dMdpEfmZBxCmV5cLgBVvGL2yQ4BNXBOLZQzuWe3A3/3yckT9gBNB/FoctmGNlexgS6HjByMkcsbG
Fpv+oGY8+wBcyCpzK559L2GJmkQWhOuCs7FD/XcccCll0V9aEk68jPiUWLNOD+BScy5zWuYJrsdv
uZtfnXh1AUL4uvtaHjkIdHUefWlGo0qoahya1OGp6aD63L/jFUGBV2RtLP/pkQHlXzgmYK4bZ2Xl
S4bEJPc9QIsmzoUXS34ISnD0RYwlfCJxrHcqnSXljrBczvGZR/J5DikD4sqMJmEmJKMyDi12wqn7
4KST7aorZpPTDwbzurOfIWxX06/o6kRHhvEmgItGddpWFPEnRvG8RULRFuLbC90ocL6rRRIqgNn4
vBIvkRw3pO+oKobNiFCOxJvo1XYIg10n8HwGcehgw9jAmies5v9Or3QXettovgG6onEbJ7pGGGrv
TTjan/QGyGhsEuyeO+5nmE+bygZ0O6pDBE+TXy8EobggLIjfVunv6swww23ZSNZC+ZLNDCroF2Rv
vEFkz0CJc6Qh+VZ9MZQWWunvcn5UmPwdn0izXO1a+AuSA+ar0SANMB9Wt0MRITY4yK7o0qVMxl59
C1icMrYYLrDA9afWRvOZreqBpyxE/W50YEsoqzJMX6w5DXxXqVeCZ0efT2xxZK0iWCW1Z4F6FNCt
bJj7X/rPXpOWjvR3SsA5NOwi8spUVDzYxDS2sjKmchX7MW0DugNxyoWaS/P5Hycaqj9CxvsJUVa0
WlIfXVrSGDNxOp4SYFP1wv5IBzeMPYouM2afEi2y0tkEH5M7dXv7A1Bl0k2nUMlc0SHuB2G3vtVY
K71Xpgk4DxM9S2NSqo/FnL5Oc3mp4wnJ8bEENqiYZjuRrvf/OI9yDOGGR3ulkiiPkO8GG/fjN1mz
XZ6moQIwQt13SnA43O2sCHPiKgte/YUJv1byfv8BkmkjSCv+ZFUjYrkbAEeSTwdGTzHW1OfJF2ni
lQ5xS7u92vO+2J2zR705LB+dKAfumipCVP0M7wUTmpf4eWKL49NIxJg17lEIRifdGe349CCcLoTc
z35YbujZx+UZj68eF4QQ2BszcpiCTlVhTc0actHVOy5yIejJfufHu7iJ21y+Sw4FN1r5z1Bf8ETV
kiBk0fviWGnHRuG+vSH0e2op3rArcO/PK23xvsfARuAf4eQgpu/8QE82wsYqnlzSZ5f+9R329zUw
CVg/kAfYuzgYZRp+7YY7TS/CBb0rc0i/CzCH4cZumXjza7AnJHY4PWrHX2l17haX0h4sIuPf6XB3
rJc529YPjLUAGMRKnd/MDTZSe+fvDCNLHWfijZiCvbHtsy88Sj2LGomuDOYQH4Udkslo5TXv+v5V
Kx0xkRDOQI5z0c0KwCBEwbwl7h544Wvs7/0hEhm578MwVXxw2uQQwy5hPpRvF1QerSXoEeVvKpWR
qQQfltJs30ZRM0etbzSmLfTJh0BRUcRFAS8JHl68/nQLRT8ffh+6MXdmYRS01TlD+ZlOy26vs/C+
Qmyr76grmsRtKK8/trzVgVMNAQD+tZiFy5ZaUIsuiIWwQ5G4CUyFOj0tgCtqR6ARViBv3sWBCTh0
1u1VMIYSC5OpxFWQzMit9U6Hof0y1dMaz5POSmLR/+3KIgIS3mYv1rbizb+SAznQgAwor5hV3FtO
2kDz76tDRC2n/ULvqAiOVSjPZy+GHR2MrKmOLhEjXc23Tkd/MBh9mm8KWws44dLUDpIlNuCJ8C+1
NkXzYrF2uBP/1MhYjEJTTUTEEk2MOqZw++EOauLEbJ90Jxs+/3PMD975f922GQX81elDxRHGosl2
KkGAFU/Vuw6v1wfRDwA3lXKwKbv6VIBeMVgx33/VfLWJkOV7eZyjUmK7EHY00Bszw5doGCo3TnBr
dBvDLUDcJMlAy+LXTN1WV+2Xm22V7Cq0fI6wW7/qjmLQ+UUe+iAun3ZAYj99+pPs5LYXndIABiRC
rA37kv42AhiTOAHXYF5+toIxvG7i9+vEZn/49Iduefadwzo29A763mkTk7TFnM5PslKoOvKSYKOq
yIxDLJlq25posSrWhn/BXixlTD1kggpJ/YKwY38IEctdJmU7RdDWzlS0q36GwFLpkfAHfnB25s2J
+MeYpjNJkiWL4SUfwyS3B1siXGkMksQq9a6kNKnqy5OAaWA0I9twU4/3LscjzgNOnHbaVCyAT8Fp
1PlfRB2hN6Hiz3DlGAvTtlao6jyZcE003k/4VkKAnwO+/rqaVjaLO2sIIX76W1mzK7pDLSv1Ujfr
UlMhFHNNSm3j37S+cgPjRhbw+5VbDfHN8VkyI2bfj3xHTsjcJId191eH5Q0nSQWuftRSqoVfwjNu
TSS75XtCZPC4n825aLWgeueDvTZ4ef6EOiK1UgYcxRftb1n2h8Gc2dE10xWdA79ktFw2wrCCro4o
DESPLvdzJPP5KdaJ9m0cUGEotL3DmopeRfEpZcqM5824dNWZlM4a6rUrHjExkYzv5tMkJJWVGc56
NaZagoELcX7HtbkbZc8rR3PI8D6P3DZfcfezULx/hNdR0QCgBNLiTdYecUT1DfE3ygMqh4+8/xbq
92fiBRsEmObq7xRLvYCowY6GAt5cUC4k856/mVC5JtkNDcthiIKPa3PpAwwhC5h2zSMudOT2mb4o
HOEGJ1TvsaeHfCJrsPZg4HY3uBT2eaXx0YlgclAlFuq7udufV45H8W0aRXWM0Yw+Ga9yr/8wfDb3
V19GsVinMzsXULwiswZ5aetb2v4F2CqXOQ8W4kaN7R1EsTsw4vEGvojlY1+1DIPksLw/RFZC57Tx
fzEPe79ZX/iWZWLlxTRpQpXFqmiu9V+gs7WTeo+PQAuMviyDMW2a7REdNb1wU0Rkif4NUtQLAyow
zDVFI8qVVMrcZXzZZQ+KxFta+CxaAfnehIvbL36KlwnJronVL2G4LC5TMp8mLJxPRW0N99dd188s
ea+3C/S2/k5L9ONzP+7FUQPb4TEcjgr3AQ5m06fotQeR74B7YvfN1zW/sBFshwPhWDB6hfLbS2SR
uQNEIcC2VnlvOgRLZrarmBbpj0ThxYM4IOc9hykfGMmN0VSJclkREV4/x4TEEIRN0oDhqs+86sWs
Vb2ZtUZCgDQ4qe75f1kykS7EQCoXefI/C3RDBbM82GREdxqS7qqWt8Sxcu3+sUqg5c1A70INaPLx
2bcnl+5kQ8V7A9ApAZBFTGwITgPu1UKKmhktzetZfqQXFTnEHoXkQSp/IqehmSmEEaZWaNYsnY4N
qkjcT5UNg+vUlnwdhmFas9zXWxTddNk+Uvj8bxD4HvTa1H1iz2bnRXesSpjEOjI4FEx3bopGMr+H
WXYqifC4dq33CAkMGUJGrjsYh1PWh6M7n4vRAac8N4CNjoah74n7c6yZDJN6I0oSOM1O7ZkIDlxt
lJzW+rIHeQUc/4o1b428TQHvaThn90MGFhRoYVAN51y82Qsr4FgnPlwdC25tdaM8IaEdZkMfsYsK
8hOFa0OLRnjK7tf8Xkjak1DDYHOv2pn7l7hlqLtTKxH6TZJyIStPHg7qFiNI3FeTqHjOBKrG3XQp
6cUh5+khfPBaJl++TkWGzdAr2+ssgnnREplkQemtIKSwIcgturu6l20LsBOarTIZkBvI1G+RBUXN
LoImEKEvs+eGysVN4A1dpULtw0UNOONuIY95NebmUkcCj4+i4FQrm1mpLnay1yDx7/8Qhrn3O/Hm
InNSqY+Lb4soy+X5YkZsQ9NFJoxMqNK0XyBkVVRLVJnJYxFvjaYHo5O5Rcxm5a6ZQ3IAoD/nhlMq
+PvGlkTKA+nqQOl48UZh+2IDlY83/GgySbfzNEc1iD+pmCHGfGHZH6ypiti7ywORFrBwKGYP5a/U
VtOuJ4HEB11cheoibunMKGHf0J2YKmZI0w7CIKNu7z1kyWFu0SKveTxkBMNej3q+WAA/NI6Lr5+/
UdaaoSEngQ7bdbAZTkVDKkk+DkfuanMp7uZb2lQtTA8jQOlos+ni9UJ1hHXUgFSKc2eCD8BXzfIE
u9q0HZJSnuDenfoss9S01vRmNPVFMmzNESCJABwW/ltUHU5kR46Du2Ug1aDGcnITyyPevelgzbBK
bYK9KgyCc8eDJNxf3bwO/AuMnaD9JPtUotaA2KgCCTJG+Nsz1leU+UUEIEx/HTEVm5j0QsfLfvFk
HIqi7ZLErfYAAyKWWWbe0vdP6MbV8CtnEdCLObROTk9kuMGrmqw5QBsiB0LO3giCnK2UMCi8PrwW
x7MfMbHFYoKiKrOfylMPjFsYmVt5geP9DzQ0/ZObSQNHzUI2+dAKsOeNm4AvkJaWF/gpXCsMaOo+
RkUmRYdE1mbZqTrchOrdZbFpMlQvQ7kM0qgJNhr1dXA1iDT8lixY6qLRjw22zhiVdgzylzoz56Zf
XAwdzyg+bKtcMzDi5opL+V8wIJxMCTkbKq4vSBy1VeP/d2/FKKSPL7NMyWMyf/PSrPBEkQsKU5sZ
OHzsIlnGlu2z9wnSVGCRbPt1asVvacsi9SkxYC7MatAGYnLWoG+tpmKbjkXCed4DdmnDdEhDvHkk
xpCoD8IIis9+Sa+wrbzba0PWiCAEptVlJW//FNuKmSiBL6FEE24+xly0b/gPO/Pehk6NikouyZdf
rDom8duSiDjv0HK3A3vI4ozU8Tg4Ukz7tMqchHh3fSwapDzT7nruaDU2fp2l+BPO5b/yj//SKE6W
Zglx5QSkczszDAw+3GuYkejcHNGSlT4MQQpbABb3ed8seX+/+o82W3S5RIDAyLmmysPo+UGYEZTj
lt2dU2SwEuXl/WHK6tjMtA3hKFuBOEAk6LQ1Gl1agpvasvejE+MsKD9CuQbRPEifEl3UaxCz+eyi
lyiNvMhzj7o8jx/7e46QZdfYIXfi+X54njDSiKfcXfxE0hULMKntzSjeDRMxDAIP7ee8WbMi52CT
XCVqrKMsqPkh3IBj6yEZoNvtiywoN2lgOpwNQOv3HMHptZHolw2Po6tjoSgHtL0jhXFPXK58VPS3
haHFKfKdJ74Un8E6RjGW1p2agLEUIrBq0iBzf479vvWTyLRNSfbQKWJCTs+U50ngpCQgtmDsRViw
e0V3gaTORH2hQLPokHHRYdwoY04qOpVbk6Qt6MIAbTVcgK4O6i6TmXnXkl8sjy5ZrSyjqDZMVLaf
l5Q/p6yxBawmF8NULJI0o8p2W5wfBDjK/zf4MjNjGQdHHJv/QMchFh3KzZAfDkd0gQluvGJtlhYU
bzhY0YT9LiwSn+BC+8atuPumRxoiHSnYYdqL696N2BTxQLe237lk1gYG+N4lrwNDvt5AagQ4Shdk
gUD4Z4ehOBNFmxW1ReKko8oT0gpRVCe8bhMYeAoF5ew3tW3rshBqOM5yJ+BkKOurrPLJk8r5atOC
l1LdOgEWJIBiNEeihU9L02QCmxEAbnBl+1HJ8O07q267/aCk5bMjaBVkNN/uSvKv5h3WRfMD5s95
GC3yMhbWPN0nLOwq+6tIr30qXx2FG8Uih+He1QIOEpIJ3xSwKrkwLFj+ArW3DjONS4qGT7/2VY81
XoAluLiK6zsOFxkyg1wWTwdjPbPyIxX2AoLu4768zPNMyXWHAFzyFFWTxUh9cTMLx3heIddhvC4k
lQIdYCvSBaiQopEnE853qHQ2aVOqla17ImfjfrnwIypPQ+BVgvhfr+2ealIF3IAqmQ9+cCO6aeyc
6Kk6dqkKhbjrPxk6ZKSgDnpKKrf7Cgd5Hp5Nc3hKC5TbYb4YpXJXg54pOP+M05RjXnto2f8sG7JU
Br2//vvY66M+dc4zJKatngHQXXerqGzFOj2qLq1gg4+Oyf0bYmuzaGvJTXLcEdAiRPBBoN8KxznA
yKhHd97BwHKJzsDGCtfP0ND+aY6VfbNFOyUuqhxFk0aa/q6uGSHx3f5UlikWuhnmZY4/PywUNGuK
s4w1GKm5kPBc4WRRkR2Z8Q9NBgHaAruCj+zSo6uJu4koxMWdRL2IMN6IqA8liXNppOmoM4/Aw/s2
HoLD3BmxIfdXmPUr6rJhtbGMNjn522nzI1gdC8M60V6yKpqEZGgNkAlL8TUQQprWXkX5bbUspGiI
mbyKRI9QVFNYXSTiSWCrBFL7LSoK1x6uB9E9GnbN+thskKqbBwFiD3iMVwDDOaqbpNOe4wivhpv/
FPVskXe6TTrVtSXEQMlGy4wBebEHvNFg+1Ej7jp3KGrmsCRX0Sjn/Qx7YIikLW9nj+6U6jGE8ysc
xfpIamiR5CbbaIwDkdWoG2EaZ58rVR0Vwwk85xCzM5ry3xOb9S0OYj0oPqXkxtfSKDXy2/A2qh/M
Yc2mKNNBtamqRbVVSqHDJgqV0Dbh3F4stU2wGvqscgXx8Qm3itXatqPudNOpz3k4ZmAS5kL36wPW
52ddkVFiyalNuEIevAiL1KJEXc6Uvy/29CM527qOpZG38EwyaJZqEYBseLPUkoVZwFxm8fNQ9OqD
mQU2K5cAqsWoPAZiduL2ZB1iUmW9yDkyX7HD6xkaHd4iP7t4y0pPdF0QnTV2z/CfKEH4fkRT++0j
Dk7DYmfpUVOuZmQfbwTe2u//qcBIsIMPJZRL0gzWI9yVIyg1+d9w6CA8oaUmcarq5CmiDKKrqZDz
JGB7fGY31Ewkeckr7wDlUqdQBgICClZztRlNVAzRqqOdzY/5ENYboA3QdK+JVN0ENjJVm3njSaRU
nvEX5Ieyvpz8zO+FDnwzbY3rW5xTIbK5jwBp25LKW3Qq2vKIEGtKreWyJKycSyujTNH3W2rqbAPI
1V6thFClU84wjCs5u3MdisSc2bV1RDlZ0G0RiwKWsTF0b0x4BAjXdVJrtjg0MLsSWA3ijGGWWOiv
WgvNpxB4ZFpzCEYWHhpvqCA7jD34Em13xfFsyz4PNS5rGcfw/Fy3ZXrLZIlEznLJPbEzRjyTUsJ1
uJK4V5y7K/oXCQu7rQfrHNUmL+w26GLEnr76EXooXG1TFuRZKI8pyw1gR5fwolM6jxirB0A4/EsK
jDfTqSOWCq1zG5LC/kg238THQAoEL0kz/bfNtf7mLXUvLgLwFsbhvAiWXqG/96u9pZTGUGQafE3p
uMzQCO5YzW/M0m7J/rATJHA73BscYLGRLxhBkgODJ209+G31NHJmUlEdfq9hVx5qFZDOICbDLw5m
Dpo+CnGCy4r2TxoCG08OwUV5A1bbO9pRJ92DKLQT9o+zCRGDvOv6yOCkReq1CuzLzaGJGsoTBX86
ewLC9f+1wIAwrzvhzCJ2Id2tpbOTJsScBjqolzuQvs6RH9m4UT6g+lH2ljKSsizbdu9X/ZHt2hs/
5wpocetWlxKbHKvDdE0KWMPwXZczNRalBMGA6IZdk6/Mx62EbqgOenu7ltdYDVdpdUqYZdC5C3do
Df72jyMxojU38uim7hvwJ8divkhMyWUx4R96oavR1x5UfOwSbH8X7xrpZu9xXNP8J1sbtDOv0XJQ
8/VSs6KDuFOBJp27Rq95AWsbg9reNqrZmsK5g0umAl5XjIKJRdxhIJOL94mwIHje/LjzQmK1YDfw
3cOLxVkLLvQHA+27CwuBBv2yrkxQCzP810tNhagmMIqGkUqRizPCOIHxtEXhfOAFtD9FsPaAAII/
6ue3CADum3Bme/WfvEmq6k0ce8/O62MCzvjQqD87Kf/lrm3HheoguvxfZ0CouQB1J+SQxLFzeFDx
gxbGgzdftq7sjjKPFhc4kMnT4jDYTgnNW6Bm6IpIZwqJLRL5PEYOTppz/lNCOscK4xL73n9Jxxjv
4n9HaF5uIvRDAVocaCofdcjNaFyU2GzXH7o61Ll1UDV1/MsQsMlkcnpDxCz9ACk56E2dD+fVhmkp
xU/KM4F79No1aEybClyrH3nelJIHwmlF0EmSsevD4xMk7qeShOtj3a0pIDNCHg3lYpzImTQ43PlY
/qOTnqKPDm8E67tQGD+WAHob+csjx3Iq7no+5UFNO8xDXDLHEE1OB7woKkws7MT00V13vgNCr6d4
TXwnmNw8iQh12pirbddKGR+P2actJEatySSiXgsEhhbiVpvVIyDehBuTn11QzteOclLwdgQgWk0y
RkVAWeXWZt685AVNG8VrHnXyQ1qSILFjRje28jsRGLa73o04MAsx+qv9enT2gGbKtSol0OUMsNaB
dNOgMHx4fHSNhJNTI8cfoM+Eyh2FjKr4c7R+qL+ZP1n1DclHtUvST7SfpoZGVJo/jJHd3tQBSHN7
hUxzarH50GelCWuOu3xte38GidA34BvXwqzSJZEPfePXSKTu+ZmXjYT5ktPMyGwJkTJ8wi9buSet
XMqa0PC1tg0oQPERsMr75OwmmtxzeTr7G4UCYtJ2myDXG2feeWh533tnGIdAwLGMBfOn63T6QqSt
ImbqoiDMQnBonlJXNweXsZuxu4yVVsePPfhPAhGx0orwFl/Xc9QOJXL6e9Vsnb1aknbEnQ8XpZPw
PY1tqu1exK2o+ti6y97IlUJf/idC+8nOZQ25Xrgr3TwBy8TDG4vJ31LxOO/KzMJ4Dwj0CGQu9B13
eiBGh/Dbq2Ae0FJxIT7jMOK/wC4rzzbRTDcrD4Jfre8n7f3H8mHiYOWuqPW4iLZS+IU8aMe4QXul
u+AcrmHFYHqatZlMusC0sL+sxmWsKIUYi8KfyIfJv1GiBRmWxZlXKxkQtg68KfEJs2eAHLqNHSHv
kswqHCyyoze7AcvukYboBzK2Ec7s+YX4QACa/KkDL2fHGZZRjhaTG+orEPjSavQOT0JqamKD59mg
B0l9gyJcnTZzCAroRj9EuAYg3kGD1rEcktXgpE20FGeRzUEzGbsj8OHOQo589GAIOxhDCsq4FXje
020ix+VZwQJd6iuWhcedSawzYHA9fCwGMliqeiVroDdkudS/0j5XuZNIa/2K0CWVtKDy7ZYEg+Sd
5YNOeXVbwNrIeg0X6GStZBmfu52TSQscGhHp5reUDehIu1nA/9G9pjvcOIUqbq5qkwuXCrBPVUxJ
MxW3l8bD8B9Me/67b3wObiF0fWoqY1Cxl+vF8Iklv0FpBff6WDB0+ElcjJw4i3M9b7j/B8QFPzqI
KdR2YPf7d5eQwH1xXIfwYxQiwXAgkYLE5c0i0FCQZnv6tp7XTm/dtw0LhcFkWwfKAyo9WyiNMF39
KfLp+n9khFHxTfRC/MAOY0g85NonFSeSrdkdce6XG/lVn5zbLIDz2mLa4fNSImSYVeX41usXSwRP
xWXSeY2fPy8UzUzV1LQgnmOzGHwqreTUrV+cir6uCI/9VibiLXk2ZCSgyU6cGEMZbOkKOjC7v5H6
YQjLcwFz/K+KLkI9cYrHVC1kHMMW+ZUH6GVvX8zF7F2opduD4FvVl8ERJvc1GSgA/l56kK8Fkc/7
GQ9zoxEntnDuzqhakx0ld7F1As8GnCRY1tlZoGByjxmu7CMDqIszSN7yJxmjFj7H5SNr2BQ2rCml
hS71bn3nuLh1YU9a/bl9e/bor4BMOL+uj0RG+hkpydZB56W17QxkVF88JhW3bGonrVX/Zf/oMPUZ
xYRxqaAH/LWp66mfO2shqxYGIG3hHiLBWFbcaGRGli5kAVzQLdXctVa0iODdp/iIPUgBmlUCSJ0L
IVkWZQm5myjXRSHiBoR/Y0TDDd5fGbXQbOcbQ1Z7v1ro2LWWqxVJGS5x94y0veypzCUkU33mzgwx
8LEGDfZzvL2cRFkzpysKAzdpgLsD/pbFTNj28I74Gsd5rh9KoBO3vO4vXaOhfAqnjZN8KsuItNNn
HBsoTgQfJXey5BZL6D86BAGA/S0+re09bMMo3l+ZNDpw1uf821sCO0+THl7vC2cO6GM94s7qQ6zL
VIEwiKuDnPD1mKE+hkRjp9c2JBL4qZ8Iah8YUCbuG6zTean6DKxPWjgs7pD8qBrMlnWnJ/KZVOOq
PXU/SOYBQB1RzZ8kZg1lOmLzO4haxFrWtNFyumUUb+J9r8LKum7tmV7S5i5z92cC7A5klonzfGUB
yM7xPl17EQVL6w4azEy2MQ67F5D37Lm9BkEpt/4Yo2cuCScNu/hT4ij6VEDrN4Zq0JZpvif2G5cr
jHoDVptzdr+C3fxv3zRaoab3kclYZkFUTb8RegJ9x5tezWQ4RP4U9BT/aD/dyoodKGY90Sh47XBr
KyOSrITTdgqsXotEZmEiqLB9Ai1u3f0mIM/xj5TwK+9Jkf8OKddtMyYFLMIAbOq7q+1NATWx0Kd7
70T5a3ILReuRCoXva06DUJ8RUkUfioVFaKUHfFngXDdK9TIqOJQsIOM882zMk/5TfwPusNf40sGq
sAWUzI/XhXKz0TOf9qzErEvXS4w2A+g/M1Tpqwf2td+YY4CjK0yJhn1DTWL8cEtyOiT/NUn/a4lw
NU4eOHtXxlz8LhZXh/HHoXAQ3JamxMs+0OyJJMElew/tbxo8YoJIawXdOQVmiSTlrSzrcVl8hz82
+XAUrLtjXwn42V6l737akPHc3u146J4r/z398wIDeD5Us4GhwqaAeD0P7m0UNYgyzWA4GAI1H8z6
gZHCNatlnEVwbvnQCs60rxfjOxqFGKyOI46u4NUfi/e469lMr1wP8+fNp4HOZCuHxkohUawt6YbY
woog5bPjaYuYdSibeNUlkqfbXNzs0337b58YIyetEWoR6U9xEPbPWAmf6c0/Ryodb7vpGmnJr+vk
qgWx1XrEpMfIVMcEtN8/wssw0BrMfJteQwTVx1Y9WdPMgNzINtXINJqe1h+ELi1NoBR6jB+LQ3EK
URKH35RkPrPfntaSfKH9rseCo/cnLwdvpG8zYxwy5mtIpt/waXZTKdNWCp66D+EGBOgXsUH6A3q3
kpsxqtUJt2UvI/1gJo2Mb/VveUxm+eKxVlicvoV4dftB48t2jsbHGPn01Ixe5pcB6wGJ04kuAuT+
7soIoODyZIE19uvhRIJGj56NxjwW53lbNtN4tvN02EAe8vC1JP1fqXpntLvO3pDGjNud4dTQAXXy
kx9NnCWsP5GbuBdJYDJzog7KqS349s5voRxNXTwSZNr++nUuzUGhHXU3nGB2xyfDZ087m2XnYTpB
wdzeF+jnrno6BDtrr3/k6NTf37IJZLp33pWVmQullkqHBsUSImdVw4giXDQGs/ENzS3MhGceGm9i
iNjWsZYwviRzP5aGy6WuLQoP4VvXPKKlJYf+mwUqkfHD2cgBg7W08NWOMhqWEY/yA0NW6Qq4/VvI
rMReQJf0ng5BHS7u37YC548Wft8cIDoFHipePKVBb4tqchvM1H0+DQ2Mwp0vyZ15idoPTd6vxZXB
p0fkKn87HNHpOhaPeTffdjoQ1W2zOS/IPcDOzMH+X0D8L2SCjGEoEi7y8Kw9Pq+Xw0hB7qKF+Ovs
AFlrgT8mZ/3QP9lq4c6m6c6Oltj87tDWiQqdtYu5lU+qQU8oryM4qkf7D0T1JJPOI+hSVll0IJr9
1CiJHrHkebqfR5GWVD/qjYLYnkyq+hVGuZzd5VeragrcSv7x38/MHZMAiRoIGcthPuGYMFTv2Xkw
QO5V0VmjdWsLO5FVEBLawqh6auHN6WZVflb00Kt/dQ5yQtuziKI9Vp0JWzz/mVG1L1e42nc1sPUC
hQmxn3Tod+12eUCdy7R+Pjoc0R+zk6qJAaHZH7l/vw1KwxfD2z3cSLh36Wh9k36zPaRUK8Zvoni0
4J3AkMbql99wQIGJobqzIn7sU1J54qgAkz+L9BA/qVypn+kDsYfNg4EXCGAloCvkAGS8gZM/YsqV
4Llm9PyN+YTrWltCp117lSHnRaZVtnpth1p/LvSfIA5Lcyws6MBqMSIM+RmjdvYrVm70hLymnTZw
bcz2RmANWe8LyWBDKUEr2h6y9KyteTHtCKkbXIEB7ehiy/oMLUI3/H7KIlXV5+hB2daVzVAX1aTm
jJRKg7AU77TGegargcRR8SZwpAL6Bf86bc0wM/FLUBb3p3++3y8KWHNj3UIdFks0vEOapswx9I+r
NeYu12g6gu5tk7kjjIlmFS/p4M1diMgEldG++Q9ZleNkQrhpil5gnB/JmN9J9R21I9ptMfI4oHYh
hl10LcpcKIAFp71Cq7JrE/aTFfiRGLqLTHOJAi4tKxceXjY40iwNiQnIlsrvpqjZbSE9pDScG5Ae
i2779TKBJ/jW0F0NUb080jxo2ljnu2RChkoefNah6uFIEOZj9i6M7WklbCKgHw2XWYo6O2h8Co1I
E1h7nZqNouKylj1JSXPs6dnFX6t8o/GWUrXK24dVfkSQwHK8fEm6z/IaUMGT1VEBK1rNSYjRQBAZ
BQySpp2WxG8lj9IzK96vAYWgs01mpaoyQu8B1/UTTQwBYDW+SFxH32R/lXwE6LUH5ZabC0PQGHnc
8Xlc+It2o9YzBjrulbZVd+mraKZHKDTCoGwMR0Z9RXA0se+GXRsoQ+PZKeiF534HcHkt9UH+Vto1
Bnvsa8OZ8B5QxiUezxuyiUHfbbv5viu9Ol8oGvAM6NJV3a/Ff9cNECI8N9nTFglgLysovghD1Fhf
/Vr0URsp0ZW55Fd+M0jybYCb5OioQvv6IgH9/+z8vyqkVJwGxJCORiPHXbOPHRE3y9TRE1xpOpjH
QafNs8uA2+dpATLcimzGY6H4qtiKBRXBaJssesNVsmka+QPilJNcBOPsX1pQBedjFNp6qOBeKoGq
wxJ3RLeSJKWe/qTvV7Csn7ykQRE/JeMGbJOvdjUPDXgCJNEKUX1O46BxK5FIArSGgjxE1XyP4Y0A
4OY2ID/cMODOyWKelSvnzy/5uTABzUqSzqw9i24cLMk2clxftwBId53AznYiGGchkK9jz5XMkXhn
LJ7Eny78129gvUbwK9kd3dYXarAa/uwZEJvT62AW7vzxpjbDN0AZL93eicW//GDVO1e3imKS2TXf
/ZMArANzZbMIKA/fk0jqfjU3S461BLhnZELn4S8PctX8hCeGYgRFc8tVecdeRNif0vlOTyjszP1P
QKdnQcGtfS1uyoBJY7Pjh6Do6pcnHbyUJSn/J0cnNOwaNodNEMHexvKN9RWTH82patDpRRCg112E
pKKQOKmF+K6CPfUaAoXpvMj7fK8q9WFYjue3aS8dk1OyfQAqPs9PFE/W7EtlRLZFVZu6y3RuvoMK
5LPYsx+8bBPJGdl2YzwQi+0HpBDZ7WdjAcugN3uks+zcN9HZK+lBIObxQaSXsTyIRifJmswd8YHa
ls1Xu+3dMEIguI78iJRmj5eYfaC2ICdw8nJwKcPWOLn5j1ovLJ+k0LapbOX8hql0z1I7KThWQzQa
iHTP1FXhB6JlCRar6Qq1g+Wi7QGm6GPyQYrTrQYxM3yUpshfo/KXj3pLnJ/2hdImhsobFc8sxGsE
VRO8svbLoMod9UZzyGx+Lcn6DMp9sexx0MpzhdreJyXC5pOsilc9vy8kRV6vWNWC+hYJbF/i0euZ
CpjDHhtwOvw4P9Wg2qvKJL6kLJf1+uQi78P1wcDWzS/pw86qMvfkxA//aogrVEObJXV+A26tjiqK
qFFz/pklKVDfGpAxk81KAgKfThhp30kEOtDd4vyMwrYqknvpGmq1ENiJiINIlTnzuvaunuaWC8S9
s9/DSzXIphm+Aue1qWatEDMcO3VpuqjyKhq0AT+Br966KryXs6vYJWbDwbvBjlM0FfPsG+MVqcsE
GbzTW4ZBoNVw9gHbE3tPVQicckgXam5pgpRfPMBriSO/kETlwxOGt2W7r6WomhBQJOX+J5S5wxOL
7/eZZuH2NR9ZWVtcH26TBqOd2DMpMlaJ2E8AcPy9UBueIoGrn1s7EGjW9B/QEKW6VZMoE5S5SLeN
5J1fyXSwH0qONV/T6eAK0sB3RSAg0I0Kt8iSuxWdtCBZcNNL+8IGubUmHb4DN93bAZoDIn3Ws8K4
MBSG69Bu3vInP8pswIqGgXz4zPNHWZW9KAK4z4n+V8QJABcU2S6f+1OcSkcEwi6MgfUsi5flPjuv
8N91fdkpwTYs0BRqDbv9V5TM5W7lGA6DLtfixDiJbR8prPBZQb4s2qovBlER7b4U3qiR5oQX99sh
SgjgHvO8TnuuBNF+aFbW5v6+lCLkE8n879/DKja3hqCY0xyiPWITxMYHdD/xmBVmDDNc+mxLubt7
uTsmrLVNmKmALVHH6eXx9WLIMhDx7nW+4DA5Je/mEBLUjuU2GSHqHdcZPFGnrR8JH731ZkX5bDyu
0xQrA2chpNlOARMTewbqawNyVGAid8mGsh8ILQPyFWfmPjlUr8v1mz7oA081+mEF+q/OPLTGCYbQ
rJNhzNEhbh41lkbpKTFCizbg6OtKbmEzd59NaEVWZoC8epqlXI7OA9w+zwXPrhPy1DMAZeHbmp8=
`protect end_protected
