XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S����a_xw�=����u���pϥ<�n��߲(:)�3���<��l6v��]>�M�l�i��s[o5O,vI��x��,k���0Yu&�@� �h�'A��B[��TKg$���j='�W���T��B�g��H��p�݉E�z�ڏ�js����rj�,����'q��G�o�������|�t�f����^{!�$���qr�.���7|K�����#�Q	�5(��Oy"!ED{�C�-��b4v��T��4s�4����V��G�U�d��v�<Y� �J�#6ґ�;������C1��a���r�O�n^	5}0Ss���Y!�:�K�*�<6�H�G�e��U�g�^�˗��X׳��q^��]�~%�6_���\�2��OC�#
��ق�5��TV,Exh�k���GjV����
�ho��M��F<� �އ�c-�)�hP����<� &��ٮ�1NU�72������\`�����=�Y��5��%�r�S�h�*�|���Q�dZ� [Z�Y����A~�.��sG!�bi+<C<Z�!Ƿ�d\�yly5�,vj��n�[g��09y�����KEz�SC���X��Ra�;H�T�>�'&<��8��D���W I��0�QW�QxX��82���q)�􁏛��bXe�J7�`�n����H�hUC��D}%P�IQ1�@TV��KX)#,,���o9Q��T���R���T����`vqQ�m��K�e:|O��)�Fo^*��5��`�'qF1��-���g�D�XlxVHYEB     400     1b0��ׅ��������fJa�Z�$WL�WH�w��c�KC�5fi���DH&*��e#�^|׆�hNj˼D#"�����c�b�� ���>�r���z�K�8����6t��_4�!B�kQ�a����}���.#�#�Jkv�Vi|L �U����jЬ��4�sQ�A�~�U��\��) l�"�ة]�
��@+.�֭Zf�H�����֜m����xQ3	J5���3W*IO�$⪍�%���W
Ԕ~��rh��Af��=k� 	|=S��������+�>ITX�k�׷%�"�S��jE�Lʆs(~�k���@=U����B���{�貓&�@����A`�_g�������ҳ.��[��*�utM{#�c�۶5��m�*Ç��{�os�~;7��f�Zg�u�߀^�|_����XlxVHYEB     400      c0R���n��rF�NG��g#�����5�A�ҙ&��İ��ᄫ�ڕ������dHCV�:X^;Y�j�\��������y��(�\�a������)l��X���JZ�sԮ�h���c���2=<(m�0� 8DZy��yZ�w+�$ɸ��)�f�D.4�����kf�_6��s�����{Wg ����� P��XlxVHYEB     400     1c0�� ����{�����NB�W �ަe)M��DF�l����P^��&;'�#`i����1��;{�ꃴ����g�e\�i�����F~M|�k�>�xҧV�mur�4�����0��Q_�/*����_5���7��}�����8�ֵ�r$��;�v��c �l������7�az-���>j���>��c���fҺ��c�C�̔��N'�2"��K�-�����&�~7��X��W5���q�|E\mo�Um�w?re� u�"��Ǿ������nҡ�R�ތ@�7NƫX�"���D���m���d˖�DW%���G2�?�a�ub�H�%0=7�!Y�TVC��%vx��Q�S9��3O���wW1�{-.���8�B͏+�榸c�f�	�t�(������)��h�ӌ%��t�K ���S.#lMb���69>����� �1\��ѳXlxVHYEB     400     180�z,VL������3Rf�
O���[�[���B��d��]��j3�b/���C���v�U��[���G�U�q�L��=��'8joY��	�!���l��(�}IjY鵘Ϩ��P#C΁���,�Tג�&eS�
�}��fG:׼��6IU���m�+|u�	�ΘȲ5���!��� ���rU5�"��Gwxw��b�[-n�7X�yp����^���G�c)>�zwa͛�s�qʉ�qR����]o@������kmH�>>�vLL j&�6~�Z��\ֻ`
���3|������L9�G6���a�(�(i&��Q%\��� ~�����؋�D���&\z�MNS������rQ��1M�Y����KAE�XlxVHYEB     400     160�Y'ц	&��N咦���}�8�_�a�f��Zb�����W��E5 jM{HM��s��#D�#�s�E���TS}�"}sk�0�w�J]�5�ѭ�9���p����'2,xvA�P�D`q"��/������Hy�DD3i�N����걅���-S)"s�|>��$�n,�8$V#����#��Sn8%J���B����u�h*԰���YU�z{�zb=����S3�	�-�[�clYӟ$���ib����D�*���;�����i�Zz���i ����RZ8���`n ^0��%�>e,�*���>���`�W>k�F�S6$���9x๫�( od�2Ǎ����Ѓ�	�A�XlxVHYEB     400     140ktehԅ�NM}#e�������p_"^�Fĕ�gr.sō�^��zp�δm��Mj��zk�����D`��c��6~�S�7����2�F�V�*�j�R�u�w!<��f�uݴ)�'��=9���/֍9Ao9b�w����_���9����	���mP)������#t�ǧ���+]Z��*10I�.�S��	D�n6�R���h��>�n��>�4�BU��"�&�����Y���U�X��2�zk5.x3Q��{%MȦpw��u��CQZ���Xb�U��#�E֦3��ٰe�q��6IF� x�t��JR �y��vp�$�XlxVHYEB     400      d0�!�ڍ�b�Z�C���q� �¾�I�@��t��ǎ�*T2��.��E?:�=���i\���y��T�6����Γ�R%�]��5�O��1�ꃢ�>�%��1�3�6��9t������ϰ�Cd���@Z�E�VQ����F�N�՚�7:q�GCs�ȇ�`�;��
����A��7�Oxr��Rp0�\V ����!w���yhO��	XlxVHYEB     400     110c+��e&��g���%c������X�I9}�;[��Krm:�Ov���N�8�r�K��
�D�6Ǘ�F��e�߬3&��&-8��7}�.F�M2�} ����_������q//<��Ml��6c��NV��q�b*�W���sm��D(coj~�\��Ξ�6���tu��* ��2�;Eǖs_�q�����||��0\�#��N�Q�˵4~�٬h�ǭ��m�{����!��@]%��)Lя_	>�"}�5w:_jm:�b��@BK���H�:�[�"ف
�^XlxVHYEB     400      f0�=�BE��Z/��./�Ԕ�K�Rn�&�xO��@��n�-D�~h��A�!.�q� Fne���:dt��N�D����(���e����2l��}���*z��g�f����>lTY�,%��#�~K���6z���A>��Q�@#ѕ���O{�i�!v����zͼF�.u�d�/���f~�ߣv@U�{?��}g��&952��1@�zE�����ڠ�XlxVHYEB      3f      50�3��[@�$3Tq�P˩�ĜI��5�6��d,by��9�4k۳��c5�����z=��� 
����i�GG��c�����