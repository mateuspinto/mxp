`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
DG7NdwdAMEp3xMoQoBKDHoYN8uSIVQNs6pFVBANyL8OT8QVgibWIXu/P7PyPFViurcTJ1lL9yKyW
GzIIyzzDxxM95fYiX3wktV+utuJGlN14GiXsYosJKRK1k2zTuHAZiK8xcNG/qzMP/UPIsBOqgDBb
FX+q6DlK5PofOLNT4l/td3IDWHvVQo5fMs71irFVP3ozZHm/CTbfa42U+eexEpRML3tpPzRV76cE
Ih/QfVfwGYlvz/kWgQjEGtu9WP+IF31QHDWDIa5qdOq+tGwUF/WCdRMw/yUihYWfB9Qybvyh3FP7
wr4NSEu8YCL+ADXJqYIHEkNfZt1TliXgSRWmP51Q3oHn0pEBFUeW21HvTHORa8ZmTKpPyLU4ZMEM
Blz8K/Lw9Jfs7J8+cu/hoUlUFoeuBTc3NyNycWguLV5iS31gJdE/jA2TARu8eIooMdrCKX797VeF
LMcqEOwo0kVO5BOjrcu52AXdLQFD8S9Ler+ou8qxHFJspOPNCsdNw5aKwsI10jHg11P5Z8iWMEZB
BMj+dsALbtxEvgxGOX12HEU2eMn3hLVSbLjP8GzrKryFRSzJq2oPGflNg/OUOjYhCEvFO3Mx0w2G
g53jZQX/byKKagECYaCNDKXjFxC3keJEB9HzwSNq+x5IBjEaO1gAESefr1D8BBgOhZZmiCJHZrOG
CXQ9WHW029yYdOZ6TytuFjXxZOLgUNbtmmy/4zqnbLvsCU4nTAFKyGh1xOD4Li2M643aJP+kNt+o
Yy6W7TyQMLanoMoiwdBywz6JWrKFRFgULnG3q8LX0PkEnCLVT21IFyWyMrBw59TIrfcE3togQ2dD
akmxGVllMcHBy8zw9Yj9Nk47QvYAPGz+INRo3jF3kfrpoG7w/9AsBELn98ihNwlD8/2+REJX7SWI
sCJAO9k+VeWLgQ4SjfF+Y6zcFuE3SWjcP+XB1Ifdel8NlF4+Jcy/Re6zcVg77NqmQlthdOfyxbk9
jWBzbnFc5vtpXbbAyvrijrD+IC2fHrjBzl9T/BsB64ykqMNyAWsZjUiiarxLIKbypEJdZbglf2AH
IoLK5yrTriTyVMhc+r9cZ88nnIa9tsvdC+HHOKqMM2pxRk0vCZd8X1HRr/v7NehBGdTAIUc5iBZt
ohqwyYyH2Ac3989NJNmLPqIoC6iu73Q1Jz9RGsiV/vvqMhrKbUrO/wprFNicb4hxkKlQK+8IBJUV
RmJsgr5zCold+rkRhzYWg3igYml7edwZ+uIvoyzzW8XZMi+pXlkM/vrl2ZZniKxJlI2+eipmPoXe
t929qsJ85dQo3V51w4v4hOSOGI1gVvaFHqxCn6kVhd+q3nGEq3Hc4HhXSLHonBUnxKCDZZk6sQZp
gh324WSH75z0k8JnTJahHGxcWmNmw5S+UQBcFgS1SP/Yv/z8tQ7nRhYFM9EONnP23/Q1phlxyoLj
WRGO/vjl4jjsr9EvA9g6Nf6kbuyI8EOPwpVuQCsmXKyh/zYMae5xauVt9BiXCAqdbRXj0sIljlqx
PwALWJgjnWUunVVIFmvu9EhxKVPj7XEbbVIrX+cA0fmqGyDUt/DAFFHT7oOXJRat/OANXez9oJre
kolOwke89bLIZVDeIR3mTyT2SRP2C/Bn+7KyFdkw0XPUpso9GBbUX81B7W90/EV2z/JlvEX90WKN
EcZ20UNWblNmn/M0ZolAtvTumRJd2usQRDiiYXfsuoVUJ0MYXJvzQxltGL6D5FtI0to/FGEPKNNc
TYuev6DPdQpn+AyEY/YK37JIv2ZHLTQi/2wssgqw5J40yIwWQ8rlruZkIRDtNCtorki7wN5Eehx4
3Nx/oyOkcCNzC9WLrCEJyeBIP6xlcrT5QZcNnP0yzcfflqHfi5eQ3Rp03YMBtGY/azSeV8MRxF6X
P+YJtiLYDSUiIJNZkEzirBusy88b44MPbnk+2NoQwHqrmk0824hRHPt+oDzx/JpvgHkkCKXq86NO
TwV7q+tCrNwYcwb9cJXCsBe3kKxY4MUzg9cPGYuC3+ds267aIcSecpk3LY2j4xJR6Fh3CW7nS9We
0NGPA2MRuvR4LQRgGtiA5Bnz6OSOYrizJwPE5hxjfNmmqX6im7zTjZNeM2ST
`protect end_protected
