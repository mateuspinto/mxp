`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rrl0N8SABb1PmUP5CAbpT/IG5k0mfRd6/Q0l3ge7U50HiYhFrUmaqN0z0Th39I0q+rS+LXgahwqC
m5ldiD02Fu2j7P+cudmN3/6x6AVTWRxgGRUOIE1klObbljE74OWvcmi0fwAMsfnxHjYPgzm3ERIz
QGQrmmimrXpiCXW6j0eJxWsGpY9qRP3Toqv7/0gtjmdBC/Z4eWNXm3zEYh9ugjTYascKbd8f72ox
CUNQX+VjH/4pyWtkGHmxP/zOl+xH5yXcp7y0U43EW97pabkawnh4uFIxjMpgEAt0I8DCy6Y8Q0bR
/RLDAM/PLKLjVHyKWOm5TyDA9XIThOlbt74Wyg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="U4tzVde1Far4k+wkes4XtsAK/nylMoo5+4CbRgenH2I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54608)
`protect data_block
rVHscGbxeL3HluhxbWLAGUu3WdjFZqQr/PTREtRog3hcvpBwj+abWgmHe1v3ydnUoFPRvynnq+Bn
agfQR6ueF5e1QdjvnyUQLgXQyKvR9d1V8su1ozaRT0A9mjYJ19U7x84X5d5c4juTT8VQRgCxjdLC
i6i5wvhAtbIDdNNq4lwWPgqH2n922U3ECT1ZnrfgS/hp/ZqQA3i3WmmLNtWLXR1+i6C4wEynfjMA
ro0un3DF9a5KXPLvZvp5yfledVzqvXYWDTSrASDmCY+mRMGlw9DMd2mO37EJRTcw/lCHI0qPPRV1
ZjJ8jp9wVC7OS/8ga15RlJPU7lu+Yt5AdaDbD6Y6DPgjqYnLeatod9XH3ycXDGQKmCL/vqtFVlzE
j3devKBvrzpn3HP+o+wNeZr9MrrD/O1Mju/nH+fkINqa2o+WRC9Ha3PXtRUbLaW6TWhsLTcsV519
SDfjI6rpDCjxjkrf2xelVLmDqicgLvu6/KMFJPWMqvVBJ74UPzOsXm4OcNpSPyw8TB0gUgJSTHya
do33zu09aakRdRJTjSFLNIJpCGf64BQqrXtcCjcDgun9NOPKgUfNHUjNTtw7U296Q2r0Y0SLh1A7
GxIALzur4eZ4q+lKpjpiwr1b7SwnCzWbE9YVUduUXEdslL9U38+HXDuYNAgGWs1czPqC6Ab1skRc
wi0jBEUmOFifXbnSGp/GCP+xF4W2igwgfZmJ46QL3dl2/xvcUP+ITEwV00ZE4Bq+Ii2tYPmfHFMP
YA2q7OIbtZDoa5MmQWnDT+DkdR2oFOS9kw9ur4k0acC1esbxpzLHJJe4gwxx1R1Nh2/TK/1WWNnK
mYzxqj0W4zEBCkCqPBT1psl1fQ28ztiLXdHX/tflZyS5hEppNpW75LcbMY+X0lru9vcQv/G2E2ro
XbDvLOOj1hY4mzc0IPqfu0A59sxYffRw47a6EtUDBUT2Q7b62kgabimlU/+F+AffLCaM/0P3Ered
9IAhwjVNwdrgom2DA7Pf7cVizBo7pVhbMBYoTE2VeHEgTsz94UzzUhPB+aa2+jKtJLvuYuSvQg/X
Gkrgi7XbIhmiGxS/kvW6B/sOANnU/DrVtIw4416ElSGBTGHdW0YRRWNvcJDd7oT2yowTk7gX73K/
1FQA68jy51qjCbTzg/g7LyCG0zJPCNH4bxCrThUde0ihiA/q+vK7PVtn8CnjYkLHq3wEeLfw0V6B
CC3iDFFat7MWOcHUmqiVUC7nzHhLsKopRG9MHo4RbfPtHof1XJcDZ1AaN5TBbPJ7N/TkJ/muB/mv
/IJYII6xU21fsmYWP89U/noXz1gCJ0UzArDXXLn5oUFKzyWNtaxMlKjVJH9ivQ9PTDwSQ9xFvB3p
LbOWkTK2PiuLgNgSEHxKXLZ4zbu3SD7GIEb70NmfwSjkssKudYjRj7b+aPsX/waSguddnDVoyJb/
72auj9geUI7+aDo90XKaMlBtTugX/biCRU/qxmb6sVdtkNnRyN9dPFI7TRe88cZVtrB3Pd9Sjwd3
wX9pDBFXbOJ5dus6Vken0bWkFZP7XIda+s+9vJMSBd3M6RbddWzVVk5YhIF3mX52B4Blbo21O0GM
x6hXbYIHUVqJ3kxasYq/ZlkBnKfOWeOs6y3AZPQS5CLPpD3R6EBblZMa40JMu7kN8EfMxj8lIWNg
8b9IavYyjdiHgYKci2P2QnpuSeGXhg0vB7jydP22g4zzVv2xAZ+tLH9m2QxwhstPaGLteKUxLgm6
pdTETssqmnpnWKdahkjoJbZ77x+Iz/sQheafe1yCWZsCApufj6xtCbwD+pGbM2aXKUmnHT5DQvyH
tgiwJvbsQ33VADyqgube2MW+hCwq+bQyaXAPCDCbzEO53Xk12i7RcI+ckWHKZdCmLpeX+VOrHp2e
uebUPE8SWG03pW/xCtfor44F64FvrXNhGKmBUdDWkvuG8gJURu+uem2N9EDPHUDeVrqn4oxvIDwE
44ESQ0BFsjmZoI6Bpki2mgIAFHQChxWsttI8LOzPhr1UC+bU4X7gKNlCycv1AtymaPoMIXKMrDbS
DEvEBtox3S2hAoz9KaChQkVwwbeWk4jrUHLOy4JISoFqiw8j+HGK0nq5V2PDRevq73HNtdVT0Cwl
o9WfAJK8X5l2NONPzXAbL6Oj1e+ycoVI7Of91CWk3e5eXy+/COJo5X776YNAxJRv8LeJlUKJrQmY
+wOwhwwOU4iw9jtBAeFukRop7qIKTPcIMlf4pU/SO3pl0NHs1oL4wHtl1V4AiD05VhZCkJAZ2ljo
EmVn7nYTTQWXhvMaNo0+z2Y5X8LHPUrNgtjmVyEFkJMn7f/E7IVUUMFHHTJPxlpjtuKx/PuEOrx7
pFkJ7csQ6gviFVD2dacGkB/rrFyXC7ePZroZTsjsWf5317Uca7OmB2eh1XmD0o2ip81G0CibJ21d
ndzjpYxyUDPPWlvnd2NQNbDhyV9S2DmAa7I5HsQwLf2C9H+TSggqXKu60YhAKknPXQ3LJyyLC/a2
znrRFTulw51AFg0ozyjzK6FfG5ynk4WitIUcrn7c4vCeEnQJ61ZgiSmGkgeB3e7gGRJedRvLHLVE
wb7DXE5Z4nLPl7hRIr2pFajSFMNyZOuvS7h16EyF8aCqi8j80u2FJ2AD4wUdnvqhtWzP2y7g+wAV
5Z8sKtfsaA9LH5gCI0jmc5caC9DlwS9fe+useJDa3+EGt/mk5ZskbnESVGsEpZ3S6jkFzuwCey7e
B+8PxuuDgO2XEIhGa7faGVSvQ2cKjHVE2DyAmf/RMyZgw4ZMlPq3qRa7YhaiEPvQ9Yyhw+Ew5yh+
aiiAJmecFspV/PhNRqp60SgKLFyzMFF22fhcCkWu3szCFydRJGLKEOJMOv33x5DJDWzdenrQ5n0N
Hkm3KV0J8Y1CUNMQyQaKSjL1PaWUUrMA0NYJDNpnBP/88BtKfttcdkWz8Gtt0+06DYza2P7MHi2G
YAa/uCYuSbUOOf8nbPsTP69c32otLoJfvWL1Al6Cy5i64/P3ElAgTqtVGigA4fM4xV7OK7FLQQuB
5MUZJsBaUVEnhefOHWQ6D/oTIiJu7UX2NvSnEXbzbQ7LN0oE1Cjlq3ZZ6lmhEQheq7pPTxS9ec3C
ccJCYtgs9HK8R4FoasoLBLyUrKfDYPU47BNJ+UbktPHopzSs77bvwvM8MZUD9g72fSTyde/SvYY/
vO2LJKxQpP4nZ1Ro6scXXBG7A49lhhs8KIGYTYag1DLi6nV/2LexgzklW425XAdMnydTsc4UELbC
hOgoIuF4H7B5CiYp5C0WamXHnkmxWsrjB4McuFt14XmPMWQQhOHRqzq7u7wSqoEVBn40bMTwp5wu
/MZPq6DlT2GxfkkeehTTIGObNhckKN2SOLQueiVDj+u0abNtXYc3W4ArzKhRUU4GGroprkDQhwYL
jb5kGdV78/X6tz4Tcb3FmdDeStvNoU89xpNMynJFOtRu1dlO8xNiWTQyaU4x+zjKAtmegL09xmMr
NuATPs8g14FG7G6L3UZYoHBedyuG9utjwQdXIRfxstPWBZSb4mpAl6uDXnSBJAcOpBjYWeBD6ncY
WTbzsyJI0yld7D/xdOqrsBAm9OWyN4EjmI94JhUid51csxvRX3ttk/f0MYVLgKwN5etb5XwgZsd3
dztLIEdPvL3s6mVwhPAgbfzQj8tC3rm4pohNdRngWc9cud1ez0DqOxQD052tfVsaq6h2PEmT12qB
AniD9SKEB8ProunhE5u/t08pNldZc2hpzbId53+F4Y9dPovwa9NxL1EurfeBeQ20KlsQVf6bmUvt
f/1daNuLqYCeNCXPw+DMPqCOIa8oBfNsdajWVCYFl+bqudB2DCfOieh4Qw0F+5wgl4Cp0pv6KvmJ
ev/XI8Ndb8lSo1oEc+aetU4cdYNp11AXkPt8rqMh6NGMe7YS0waYu+JLTB+7HRYTf53eQZISNj9C
pdILDOtyPS/DtA2A4Q7ldIA2rLbbVplqtlHGC+vKwZuUhaCs9AdoKaHy8IBNgxbjuegRSRzkwBWP
HgCOa6YOcfnD4JREBriOqNoARSN/zY5/zMA0lzLDtp7qhOGYnKpmIuAUT1ZkDcTA73jzPsFm7cBs
/Z4vKHIaxrsudIOxc9YdVyRObZTJBWCx94Ix6Bbhcg66ke3rmT2QRUAtD5kSSc6ZpvppYnB/N7rG
3Q1MeJ7BG9yKa+IVIL142MZNZjBFWgPXPCxPM3lwy5rQcMtBJj/1oas1e4JOx9RXjzp80nJs3jMV
tMeQmUVGq5d69I7cBdMyVCCitTwoG3nAdl1NKScy5T4OHxPUoJmNAuTYtiG92Hhe0ATZGPiHfQ4h
sOK9UWBAk9DxKW/6szikGZ/zxkLr+Kxb4EzYKan6m8AZVwLZDSpki6xQFMtcq/yyNTy6QudjkqIn
8/NuNj5J6THU4IYEAb0NpF0eR6Pa9MBMOZ6TV5Vk9SPGn5nFTJKPmHfKkqqmfqLCqHmranEmEisX
N37P9FkxMT3pLIpxkSTBkB72ZV/7fkH1toxs0D2BkXSXGW5Y9VxAi9BYj29SzE5eAPJPkEQ6NrOQ
8vPfcCiEZhdzuO7yl08dhCGR1YJLrFQPhbbIjAOgjOc/BP4NvaHp8lwODjzn498sKhpt95MdJ3Sb
9zuRH+ynD4pItxXTCbJRuMRAUVx7fawQRSv80q/XsLl2Mfaxzvptmeq7aEH0Nt5twiB0SZqjNVH8
PcQlaFtovQEAtNGjPcKtGM6bsglJQGIl3GNOKWZmaz6Cl/ykgKmqRTOfQZ1aNNdqq4hOK4urWZ/u
q/w6ImaSqrhjPApnHVVi1GCjSbL75XHgFFbr5N5nKDVpfL7ro3aHt2DicXf3DUABpibzAUPDdGjT
raBEJ2wChHSCOadiyN1BFjSiSIV3yfXn+v2YC06RlEc4+5QJtrAHc+Xw9J7UlqECvkn6oKqPCWG0
3zbdDD1IjUaC/ihBh0jf0z2VI9I5X1a7kSTgpXBrDj+WfOxRofdiccRhJuhMXxztbWeeGLRtKfK0
noE/+OHf0tBugAdwo3YN+RLFJmjLebjwI3FDwfNwMX8JUOVe1FzF7rBBbANlEm5PV6hT86bPEHuV
dk2eFPbmvD9RvFXp+rq/kcNT2cc6oOQKHSB04jqdZQ9kjNEDb1MyEDXOtM3qLFjB9/NXkErAM4tU
8QVFO6fYryuyNB/POIOmQfpKmRRNt7Q1fXHXMGmsf7xxQqaTXVu9q+YaSuvw8iV7uSKcFH4zfByH
hEEKlsdfuJNyJZcHlb4XbcoaOyZu0Ao43aJ0yHyz2r+1SIo78YAZiyq2jYUtQwLkbUfsoKNZT8S4
XkwabsLGVeG7aVYVbS0eHfRRlrC3rU4Bok3mg8KE2yn6Rq2+W8Wk/x204N8rjfyPf6Jhjia4NSjL
c74G1+mG1Gs5yVv5vVK8bqMbtL3b6l8nIH+nThaImnAURAc9uDdlQuphtpycFjCD0rC2w4dnHIwR
6/4tb+NKzg1J4qFAuP05XGfEmZTBZacM7cycUEEgWLHskv1hVYYeN13uWvYwGS1TaNttSp9CR3Xz
SLdpSJj+rZNiQ86zl318ksjqaK1ufKWuXS+8wKlJYbDpKrgrcYVRb3lPPq+8LqAVDeRE4k2IOKaB
GP8iP7kSGILc3qHH7nZ8G2sV3Kv46r7mSeXmvhZjQmcHHzPuXsRbsM3G8xPRRJyBi8glK4ep5KzM
hr4Z6fcn60ac9M0T/ZVaKSNvYtvU/fOtVIpRizBMFNu6tYxWOpsFV3aj/xCJMlkOrGfoTyUu+9Tl
Q/EEF6NyIjIGEqSIlaYlW0dbVgeIvoiGq8F8ovg8WeKGzISrO3Rr7KyIxiI9nyd51DXBOgfa/7Ru
23W164+AGGLTcKsUZBcXTkPwWjvoXzcAt0zLeTibJAI80Wy/U6PgX8PZVGdp0DxVvfoIX77YTzEo
KKMROihZBB7jZB7lPfDiWlukY82Q3U4l/aaY9LPefDEruxjTVS593t1G7yzZFk63nfaYbJe/bbVH
U4RQPElW9YvFIrMwmww8f9JoMfWm8vEX3m4uEMdXBPz2x1hMLvD3tQ0ukyZW+Gh+0m7pyI6vALb5
6BMsy7t+5exiVZ292ZJ9UbbzpgW9sX9l8I4JU4pvP+hySCc3NgRSmNOPpUbLPEOzx0bbmkbxqLmi
hi8GvIEQXif//yaQyx3Z/i+eFCKJ25jz5M7InpDE3oEWb41EL7gI3JC5ZkrFQ1B+2yrlZNxuruMS
9iQjBKpy28pq9lQuX4zJ0JSF4w++2d+lnnOyGaXZt4AIa6VWtSDfIFoqJ5GV/WBjiVd6LysI9Q/f
LLEneH15sCTKryh7dPIm8LB25uY3MH7cDpnywe5SJAA0h+q+cuJamtMPGnS656yXXxm8xT7AWu9h
qEjodGl6UOlnrt+wjMMeZlz7UOs9xGFRDsQ0L04/Lk5q78pWnjFhlEVoJ5nbBplJBn1XTEAp/iGG
lpP8+PWFiNy4+9Kc5PU9FOYZS7+pZlauq5zMdXd+ViuNSBSnjxJha86Uk+heIpRHMFxYTUqs6E73
sDFEry8K03Yub5Xe3PRBeWJBFZY4JUJRlKnTJnuvB+NloPn1Gfgh80ueDaM6mzWn1n4Jaw9ioWyi
XiAoD6Lc7P3YF9Dv4iHMsSrf2rvlG9JMRd971tefBJn52yAW8YGwFVxFNmWEB3XYm2ffjYsJUTsL
ZCy3/nvD1G0N78pN1KC1l0JxtRi25mT9xsSFCZ6yT9Cd1kb0pYp0Zfuqy7gqThrwRKwX8za+St20
lBSw51vH8el8PyLoTalpZY2pd6ZcZmozxnaL46NYOjupUY9ssAG+iatAjgYSkEEqrMf4XawN6+g3
8Y9Y1fr2E4C0JLWka1qR4CWD3HCrqZwji1UVJ3mFxWC8gBzI/XNV7UkzvQS+omRkVwii5gZnbBNj
2m8JlI5konksfEqLp0/STiWo3dGzXaB5R44VN2wyDsq7ysc41r8J8f+dRhfFg3v47ZecHPsyK6uE
mjsdPDOkL3MvvfM7Qa0T4QVoQSmM5C2mkWVP5M96c+u1jiwJVXkwEo2/gD0SJZZQFsdy8YvtYlWx
qaljj6cJgwTGGfiHc6vts9e652lPNj0nVcQAxjrrXH/dlYu78okbKLKoi3x0DMeD/l0QTDLvJ64b
zhgOGhdYcVEB86lWm4okuNH1wU66a6gYIQ3FEyUEPIOzIKJgRXgcJ97eg4vPedokPXwYztmlelV1
A5gzYgDtafrAyRM0b61eqanF8DOPYpbhBIrHDOfjzYL9Z1PpyMYIgohjyiePZuo6LHcrmY1erVGa
FcO5IxQ9x4QFO1yzmVZY/jrlbwDMWE6oXeFMjaNikgbYnG/4qrmxWEj7bok+ypnJLpvSOvi81MTY
AeTdAwhwLMVmomA1zTQzFoybingWBy4jYD3Y7H7l47k0R0v7A2ggTbY08n5iZo6qwpt0F7R6jt3n
1zh3q4wVWOaV24AKkdjE15k/YWioGCILySb/HSPi52/QN5ZA61HTXNeKOD3SwoYBQtQRK/H0ZfCN
8CoIYMLiYxdWBYIRtsd3Ed6UkqJbg3IvdxClGWg9zECVt68Fzx6kB2Z/pTFpjgiXcH93EM9G9ida
UEkogW+Gl2eSg/GTHgVNaWmEEX/Cln+KQkKmbFw7nbYR6AgA5LBAzNONLC1mr9L9inJWk9VQeRuM
QXUpHdMazzMD/RRvusf1yE/+bKURwRC6+YWYFw710Yk10UYZCalV/vxWodgdwMNTLx9mubdetvLi
RoIOcc7C7LZpeKyZHIbmDkLsBo+oqm9dhDFppdPoR61HXlH64686M612aGIYhGkVuJGk5FGTZBP7
I5LD81W0pmjz6+dlawIuaYZRkJ20hfQTcSyH+cgQLz/6X/uovf+s1oDbUxqUVYO0LNElw1o9JYoZ
MBwUbntVCXsr7Z5vAj2YeOKAaOK/2k8z6MnkpTc8dSrqjNvtzsx1L4u6GYOENCBZbVG2CobkWDIo
+8vZGKCzrKrrGuEV3J/W8EsrUQnRr/JV4otJ3Lgv4SeLBZ624O7TV0bhM8YHMaSFKg33pea4ydHG
WGBU4qNl8gMZqqZSAycfS7y5e0YWS6/i++LivjehDkcwvvaIQ20HqY5iw2Tl/NS/yIxCC456WYcy
Nfcnywt7TrJnfLWCRkoeHXRg9S5HyxYXjD3N8ODJUSXm0vs9OGnMImkE7K/e7EeBb9iTp777jqsi
eHUlFqq/h/69mYiEk5NEgp5EA4J8Aqixq6zz0+fD2e0S9D2z4+Wrsj8n8J1DYRO1stibP87hQvYW
OcWwD7mohsVmK+5NyHMFjAc40RCo7bOJYkYk1qUNLGp0z/LpaBvMYKNWySQd3lO/S4mAHuIbWJWP
lPlYwDrmkzlSDHCN2fNNyrMW5wSaxSaWCp9YdCiztR5ARx1W+25t5fWYrNd7jxIoITchfI4k6A5D
AChs3RZ+taqdwG+jqG0Ls2ng0AzE4jjKcYo5JsWAtDHBHtr1qw0bhQvjDqPofMaoAsi4ccvLUIHC
SwWRMwDHd9wQpLgOBX5UQHdFthzSiXgIkLIDaO7UKNWiMrqdFWNtG9mT1dPyU1tH38GblMBc7r9s
0FID1k4HYoaGgnS+t/fYTHCQXVaKOFAWFa4ctaL91mFsp2ExqVv2Jkj3w1esIiHPXje8l5CL/2fo
AwVT/6v41g0CiUwfXWOt46V/cO3r/CeWQtgQYpNbpHLPJfVlco3CwKRsQlM2v6j4/JrlJRANIQKj
UhADTwUCp39UXQmejo7P58XSu4GHMPRf/F8eat7nPvdkG+UTC/CV2PkvFomgKUoSIJfOqobBUAx7
Z80vQ1C0oMYRiHA6uNReemDOIjYyGf8fvvOdeqabatIizWYHYcCmkj7NIwvK+4F9sn9AzfCgCLIu
TdDha9BH75caqgW9c1YfF3msbsaK7i/opNWTaILQFQWA68mAdCh+z3VJJR5q0BHwPZcJKw11qqsF
5nILWnc5HD9ayahpDqWxJdZYwcgfdwg2clGiRu5rlebq1geXC9l6ijAUPOTsJksHy+5Q9JgLr9Du
TuuEMXeJ2HeXlTkW0x3qgdlbodHNkjAo7MOLf1UbW4sGVzyxocCdj70miqK4VQyBh/+z/gFGnnUQ
hyuV4h0RqWoe1rPiyTWDqLAhUTFnVeUvc/oB13Ybt7c+xLaRzVax+ARRgiCKgCs9IwyflTvDwMmE
LPJOJtjjjo3dQxv/jLtMDxDXqSRCBJJuUmDVjxaFfj04qwd8RvIl6SB3eRNptDg+5+dUesNsvN2t
652PEGcgx6xPUhyB96ub7OKfeaIpaPTDcNZBWbLrG7mCYNOICA6yPHz6M5Pu+pbCEDvsyxII7Y2B
M+azKK2VlUQ55TBPQCcbnx7Sr3MLKMTdN/9v5wfqLcjKEnj5bNHHSaOAJseFNFejmH+33qywKb9T
zrel5yZX0PJ7t2zNZw8//0VTJ5Y80H9YjjokO32w0CdPOzsFdgOWDBeC/CeT+3gqEKYqFAEb73u5
65uAPD8jA1UPF7kZojVHgEdqrXFAZmDkBqLbY94tUX3chlwhNF8w44xGUw0latt94h8+IoyafHSO
zn/1E2/EivCwXX5bKM+yY8i3Q6KdkRNUYpAOMoZicjcGxhA0XmY7z5p+e77javjbwGyyj9GRKbkR
+bT+xDCgXS1aknqw1hEgKGnkOO8BLmkO/84s7gh6x2r3FEa5H+ll2zlYkL2PnSKvTVvraEcYtMti
FpLODQt1vmkdee/yi2lxbklktUYa2u/6lkOx26gKpixtTzrb4P8xwDwM7EWMMUA/Gi4ig585/0eq
5d/frqgGaVC3O5AwQaRfjECc1W8RAOPkkeURSE7/tIy9GzHLDXQkvcWYU7/lrUOMK4LyOnXMy4iH
bbIJlRYrRIn3wBA6pyXidEpFFRTDPqw/7ep5Sc+4ZoLt7pcfIF7aLypWIqsC6JU0T5r8HclQ3oYS
GGAqz5E6UGRMrXOqvoGeuauNNW6QCMYZGCIKBTXNEz4qT7N7YEo0G5F4YaMLd3HmHksHtuMbfvrZ
+Wb6ZVbJXKO+9kSet7AXxEhJzsMxSjqYonM0Bk7+t4PJHSthZtgfJUanoJPATdQCdpWM03SzoO0Z
o81XxMuJtgd5cjvoQHN5wreikFoaILfzwin3W7XZzspTOykXS//HR6LZt6tiw86mIYVLyZe4WEqZ
P38eMs8qRBnLMVbcBzlQ2sXO8BXOULrg51MsBPlP38fogMpzjzFUSEcJB8ZsfQ8y6L6gMaNIvddb
h7BIcRo2Jb9PqWBmOLGc8aMug1ERoD+aTBF7Kqhtzhf8n52dCLcLEA6HfDFlX4XAaJhKD7EMtS18
3q0hI+NLbM++mZPXFDmnO22ARvJaR8Saf0HxHTKK43hfbXUv3prnmkG9Jf+VGN2qHJkrw0zUKHk2
xdWX7i4gpuAHfqXLbGIFdpYzfVVCTc1LJgHcyUk1G2wKngnTWNNoZbpMqODIAmKZJe9fjU/dCb6p
hBRpbdDcveG/Kg0wuLzKa9k2OfdBUbShh4t3i+O3UW2JuNwyfO2wmtl++4Obetxhmz+/0O2893l1
pCCue9Moi/o2+/t8eyt8ajkT4eeRNtgMh5Y1TwBB7Kno+sjZxH59LUZIbAt7a+Op+nWbYnx3hBcQ
+XO11p2sfleJID6AerPLdQGgR8NMrbHUb8wvDLiJBE27nDxw5shKDEQ9cQOxKbHXvPt1x6u5u3xT
5pnESVF6Lr5bi0HbNdABTNjsgWKi5Y7UAiIE3n4OcslJVpl0JkwUKzBtwSLWRmDxaLvpnQhRQCBq
TgQzyhggC0DSzH61xLSHvDMw9SXDpf/gGWFIUzETBUeB1V5sfJXNP6x6K+fy2Qxhuo0E5kbCP6tc
a3FB4xeh3VgG/KMYZUV7ei1hSLBpeQva86m9PUaNonkqlsnoMauPfoCL15fJlnzZyW7kWxztW1XD
9rIWhAcavrxW+TEl3xJdcGBeY54DhcO7SYkgiGZ2jfDfWMV6ymcOpun/Q2DZBrTlYiAbAd/P0tY3
SeMSzzIz599ib8H+lxHUKXN1xRQeSnkto6wSSxiuHMaTEO3Pmk08wDlL6Rl7Dq7dETFaPBBqo0XC
NzrKk6DxATnIt1UOW6TH0tu+dMeRerRcrv8xNbPu/GlVt12SKG4ZJC4F0McRbarOCQ7vxkz7x85J
0z6+gyqWPRxbuxICdgyezMbN1oE8L7rP5OE6feLrTzorYePUpYgfSgn16WWH8ppDpFP0FNOUlSHj
sySV7bWL8I/OXKdoIMCrqkoO06xAY4Gts2T6WlPW+D0Sw62yweNMPOLwtOBq7aT4fzhHoZpzOTmT
9RaQg0+TtTydANP2/SLmFovfptOk0m20gmbLKoIb+WyUXEo9SH1+cR5wW2T85SP1iNNys+s7LEnc
e7FDJp1vXkH0l74LkIOQfNa+x51Tzvbms45eFtblLH/6HWaZPjDQTAaER+Dw0f49SLNuP9TVVXib
O7/Ly/Q7Jumhb48BQ94rSDELw6eHv03XGbg32Pms6U1mMdaYsHH1Sm3zc5lnMKHAhYYfGtq8qnke
3PhW1e+qhtnEjBs91BNDsd3uec+HmmU8NiAJunMUVmP+kRBJez+rxhzQzK39Xk2ugXB/nVZ/b1a1
68BJLUAcXR/srIgRrCoErwH7qgvVJaPyGOZN0g1KJAiAamiWWHCBhWf4lESHpDrXkdxGfniXQBZc
ZfZi6Wtsn++FeuzwIy1jIBW2KjTdUzOGqoKANLD/mrTmgzxzpiqvcLcwu6r9/JoPsz71cK8gtVV8
M0NYZkGh1JW5oTyRKHbHqH+mtcha5H6dkZ2X9WF2+RjiyfH+Z5IT5V8owe0FcjfG7Qsdfk+V9nCC
okPEFsZ4hZ8ZV4zHXEQUAYyqVMxnlcXZCBKGrEoRjmjjWTna/jJmUiOGAUkTLiEl5JkCB3PMRgBQ
npZVtbWOY/YAZVYW9F97OayBoXMqPwXT8UCM9V4Gdp5ZD9HioujYPIosnnwU4hP/eE8BHUErlNfd
ZXl2lQqexrBsU5rk/FbQZyTAdiHCAopw8OKW7YF9m7XJBHeveST1wVc1MB9V9yZpZPwYQl1CPK53
/J9jBiNcNciwFN6rDPw504dMw0v9D1+HHv4UxzpymumL/QcjykdnvlQrTiyoppgtS157GuT61MuM
Ji5oCARR+hA6lPV6kZcuPyGMUm+PAFGOARbc4DIZnmFwy6cZXQELNAe/eO9trceG909cB+6Sd9YE
eBAcRgqUB0ahSyKu/f/aZvwWpZMbthaHqsg/IfjguXX63i5FGY33Tuq1jaMVEMUgp2wNfc73FAQj
K+OEyzDIjQjvEe08P3rCXxM05NxP8OqHS8Al2XB2dX02iFJfZ065ww67gKa649Cnzknz87t9ZqKT
Vw0M3gp1FatZAfSPIA4W3lRfk7x+wW8rrWQ4410dOo804fDdZLvn1OuSITtchOMLA9J5jA0IZF+g
TrjPPoF+2NwJJXXpvwefx0Tf+cEVZqhExtymM5XgfV+D9ObjVMQFZpXXUp/vXKsAciaBf8uWvjnV
BRAH3bhZ1mfuQORVMbByBpUvUvz2ePtmZ2nhpEXF0ruW8vTrEV6lgPDMABodVm4PmUj6VH+IqkLU
EAHZBhpUjgQV19/4dQkQWPOp559vkL9aeVDuYxrd/LSJjb5JWynbRJeZRsJcF4Mm06lTL5rMqdUA
I+/N6PBFctwNudrA2UVDE12pHu9H6jRDI/jP0wyC4A9wt0Yb5AcXtZnuMpTCLxsZqdFNtwx60SLT
RH9kyxgWFbPg7vigOnJcGGtxhKDeCEKTLMHuQztOoVyw/V98rOBwoO/kJBM6nzDeuyg3sPZYTeLR
TZY8Y0NwVGkFHR769cwORPPMWKHT/eQB7exAgZHhmiOEpRD6TfnOWO4DeUdEau8yULCOoWKEzj8C
rtJpTLgJk14xk40H6L9byYx6bx/2Y/l4LU3+ZTo/X6jdamL3p3d+G6EK8Tm/KUAdl6ZiEn+O1FDl
l5c6udEsHOES13c0tLiISlQajgFjbq4PWhZRP6+aJM4udH/m9IUDf39IWdpphmEU7AXN7dSC8PL/
cxF22RUNLQIx+KvGY60NAJxwBk004EwE0pFxwUvuxEHX3UMoGPXA6sC8DKaLVJK6odCZMAY2lgSj
tbsk5JvtboPV3WjGmMuuiH6IvTl+YINS0AIyF9b9nrax026NObBeFf5tBwULetIB5DYuzhypCaBe
hLBa3CRjQrLeCwReU+uDv6oCjjRLXHZUzz/vnB+SwRiDIp6K+BvcD2aQqcQlMUfZIbAIPXDx/sw/
dU1ObARc1RixwbctvWkxGnk+SqRTzTalgNClEl0vGxW70eskqmBl5HcEGoJZnkRL2/eXKl78iPsZ
AizNwR5VARh52FXJ1ViftgkfBWBUE/98cWy4ZJJPksbc8hsfNgYV2w4I2PQsOqi17Z5D4jhTfj/z
jQpjlzp0mK6AS48ESB4arVgZXm1IQLgDx6ecCO6e0Y5mKW/hpvl7JdhXM48tDLqBV+T5P54JuJlQ
gz53XQ3JUtqSd0LnupQnU3VrPRO7wWKMKlIurgL94LcVVK6auaREf9R3Yye0RhihNvPh+zhtdSCA
eahIN+/+T/LnEdzZ/Y8gvAluyb9JjaGzre9MGAfPW7Brhq8bWC1jQj2oV/zlad0rMb+GtubtkOAb
c34I5eWOCTfgKBXwig0oeDttEghHhynLwtMnyDQji+fKCrSqjZa9mniH6rUnuwX5eq51/onHaqU9
0ffIWcgWWMiFAY3RKisbrAgxJOVQGGqtcB11VFsM+bQ3SHNU0bNezIpuMZMpUkmpzR0RVQnkdfVB
fiNjbpkvdmhoJUiset6V0wJUBMp6ky0/IVqgtLw2gmWEf1A1KiI6FI64uS+AFhzGBUmgxgoi0mPr
LEN0vojSrsxxwdzUw7MzyyV+FowhRX78b4LqsVJyLSq2v7+5U9UBi14osP/+ay9gfLAQI57cZYXr
wesv/xafocbYRCkMgDJ11nEKQWXO5j9tznjOIJ2RdyPJIRbg0jjKcQlJ2QCZlNYLh1vjfsqDTZJN
Q7eL2gsgJrCGaKfnCqnzp5JhCSkSDBgM1BX2Ia6fTe38W4Au6RLmBJc0d0fktvcX4xGpGUaI5Pci
Rr50cGPr8Y7c+reqQWuo11pM8zSgmWhV2/Sma6LRl9EKaBXgL5clUkBuHexsDaPn44j9xiTB9fz6
vNHyz4GuKugJ3R+RwPbUsjGZr1B8GCf7VMKqRLrBGOAJ4JEvq/7pya96WGKVAG6fk8786eUSzWAH
hWyc3z3XQuOg+zbT91WAMoZR8LWQxOkJ/OqBaS/z1Xh0nolB8XV6hTllWrIod1HHYbIqkg4QLqVb
C3r74s5dYhQuIHeMHNfNTS69TVJQnABxKCNQJ1CfTpnKLCEiS1lKmrI1fOcG0SO7TsOeM3R0ebCB
mf70L2+w3uwKWvs7FgKsv2P5kFZX8nTc4SYLPxCEGfSKEY2WckCnIxLfJqZzUKIP1D4ih9Sx12TE
kxkBYQzwdH18d5Pk6GDae1jMxypBH73LH17+97vNRQfcitCMG/JJkTRcRfk22IARq1JeTsSWb1E3
AcODiZ+xck+6HCBb6B/Y9Ffsj1e6WqMrm5fFqXGye0AMTS2ESGWc/q38rZlkCAyupg+lbMUSrWoK
oYCZcp2Z0wvGx6ev3oM8I9PXoiihV0FiLXRO20bvD+KE/rDVEDpzPbuHr08WHXt0FD0q8CcefJQW
S/Zv1vBzg65ZzPJiktp7pRHUYwn3KpNbUVu4Dg+tteMuYhbiBcdYpJtphIyYUKDoExNXLH7hbpkw
z7CtJH0oJk0OrO9hUh57pMb4hEwkJeOP5k1xP9R2hELBHIbU9KEs7ulpYt8ggajlbcSCS7az3qJW
Lcx9TJvBXGgcMi3t3tuZIRsTv7dYpz2t5wBtR+GoGnvXRED+BBK0YEa58yh6v8aN5CmN9aC98l+F
h6X8AIDJ6vikYQIBAsiM6Ng6L0CDhmNWDqh9JbDTEec7q6HOn1chwIFbcZwifYdSVLxvV0iCgtMN
dBQHlFcwwnOXN2yzCdn+IPV/hUTaOee/ZyNeHpfZCjI7lfAGhDNnRZum3VwB7f6v5zbK02oKWWEA
Lm150EZpvm9zFCEm7T/QlItQO5xNYaAWgghreJAZQV4horQSC6rTAcmImU/5aT1SXcjM8JouOLj9
0KB43FN+KF+VTgkn1T7TZqeZvDVv+1wtID67KqBSUJQ0HFBkQTdkNQi0zCFHlSqStfA3PMqjAiyH
AlStT9wIZu1S/fnuxEO75JH7xYU73aTEPiH2JNWhn6pZlhe5LbD8Bfj0lebmCqNhogDcCPt8luCp
lcGcpSuP2NUyBbR6MpDbQlp4u8ofRybV+gCcdp3+0LNk9u0fDpOr+hK19p2VYv1ZehdyrVQN4gan
260u3B6Olz/lK8pC8hYSgQpiZ9COYp2gFEhHb165bUkskKw0xMY362iqG++Qx+Npn2UBwL3DchTn
oKOW9ejpTNpQLpePEygqU1cAvVjgFq/jj4q158gYdGjPkmPPVD3ma4V45Y3SKJTADlOLJB8hKnRN
y5g4en3o+hWKotMrPOY/HK0u5MPCcDVdCpFDT5FD0gZLGZbVNMQg6a0qbiOlh4/MzVHV5ielVeRu
L97VlW6XjxV7WwPdL4Io5u/N/E2TBMISighACXocf5nQihm0N/8C43JfKCsQupcS+riAejGorOrD
c/SKsS/lx+xH76AnKFdmKWWTJaelRDO3RZNP6DQOVfccC6SLWLjVMxLQpypSLlYM2VNwPTLZHhoK
MyKglgwFbR83RFObxMN9bSFs8+bwzAwxNHcT9xg8ya9R+eu4QCfhr/gwZvHUXrqQYqRMHPSuZTea
eeVVPAEvr+BeWabKbhfoQpKc2Sr2kG6cUb3VPo0xo6QpeqBPsa+6USK9z0i8VxirRgqmszA42nM8
L0kY9cr0qKZdoY1k8pqhkPNRnf3UqqS1YuWZHtWMAwZzWEq7ZJjc99bx0jvdXQb1fWjwdlPOalnR
WXrcWt2VOx8xJ93Ie+WmYRm9nuyTV0NJ5Jp27ca1MAHUsUvWsN9kYn+Qb6h31Y0jOAjXd6J+JKrF
pyh+kWQX6GUNlGFSGXcssDds0zzT2bzmT/gRKDMxEuZmtEjoIw96Nm2qGpROwStcD1YK0jKT90uO
FF/zGuvnJsEAwAIzOtWe6IV8EhV4ofwPj91lIQPleOfHsnUhnMubesDWk1fHNvyyN529djmWlJpB
YkGvbGsQsN7l95M3uPoTGf1BlLXjy3RfPAELAwT7St7TdAEL+KjUcSCelmNaKjIme54zeikakHo9
SOk8s0PhAxjrI0Bcl3P2FjK2eQOzv8BXn+pWYMEMKoEiY97TRgW7M6foA+08ZdUG9cjK7LXVbuei
MfZa76UKwj5VyUg/+c+jKM3pYow4LWHvbZLaxc2T2iesc6RXUnk6Wp1F15VcKbyXVE7w07H+hvH8
6+atTr6YxNtQeORsETwwmp6wj4uBL6qhl8gzLEyBqMuH1OmD7x2+wHZC12ZpmFvClj666DAYIuZU
34lMvIf4A6QmqljtqM0mv9PehVS1wvxGIjYcboHi2k07qUjXLjzYrk2bqwRHZW/kTgULHrvjxoIM
oxvJxApSnKRcFXUlhGKppxjmM+4JiCpkYljZTiB88ix91HtRt0OremIazjCTiIunxzjmAHw3fxJY
Fiu2IUQvKlrg8yAHzZmWRGyh6h38v9CZIq9R99Q34F6Ep3rZwPFKiDfJcpRQOVCBOloqJ8Prh6A0
owvug774RISacnggUmAq6jUlXgH+A5u9mJU6qtKqTrLSyltKtjj1RvJwJSkYNP7liWUxEBZbcbIf
RrnylNrftI/FY6otWjgROdqkVf6EKBG7jXyCPck85wlB9O5dZtRCcgaFjXgektCH/Kd6qHCINLkC
uGKLwGF6qRKaTVwa75wFXm8fv2xCPRexkE3nfwmpyg19D6rhmWNpnFy4gSFzGDeu+bvPeNnzzzvA
vMYdhFJTb59rsn0oMh6RweEbRN5IECrOOIKJGlXRq6ehHzZvtp7h/u9a/igWbP0Q+aSWOQCCcq1A
JVCae0SLVoM0dUwFGM1VsyjpFFun/kUM2MWr7FS0EYpS9wTX+ZQM85A8sySE1KGsfQmmCtr3dW9S
vQAJzWuI4wF+8OFj7Ok+cHTdv61yGHTJkJYWn+E6cHAHdt6PY1y1Nh0y1EENo+pQHXYrcPVJ7eM8
u+U9Fp0C1AAaOsUgyMSXb0KnbeaZPUxP813zFJJp///547oMbt0fOUwgOVySCt8XjbeLMAQb3gz1
8SOypK8bLs2Y0nxnrtbyR49jDtd5VDENJJ5qitVTFhS6ieCGETII6WJe5lIOdxL6GL85pg3kgvvl
aSjTlnoNWu8HgXCqYCU+LXU7+8RnwumlNIgz1680qtIX+wxbWIkLXO7bbnrPRHSucbLpnptiMVOj
FuE1mZ9Ks53D12fRHsnqVioj+Sb0NOXFn8o35xPwCEQI8DgFygKWOAOlRMjVNPbwJ2pHHpRQ0rI7
HgrwziJz9NadRAHMryZ2hJ4NMbU7JYAHvPI3lT1nZEeUp5RQb7O4j9VDxZfTsrF1+n7ph55IEuVq
dhhdxSW2hCZRVENXdValuq/LrOeYUHfeYdUEdn1an8HEbM/AnMd3mBbiU0ycUIiyLPB18rcdUVFE
dtW5UU3+/Df6zLIa0HsxHtQwgPqd4+GS3PnPzPOtU73AwDYFgmj7sK4YgCwaIRM8ouvx+vV84tBZ
/v98YL6UfQLxn4saqO127APGwxH+IHw+NZ8mcfAET4wmjbhLesCP8XKltfi2X+WVUV8jrNNqyHul
uepBRoOLvakPkMdv9bYz3EWARVBTbxWhevhPSMrCdQneUuP5RweFA0ofk9yfBKQ58pk4vEkX1OV+
ZBWnf/tu4dmBf64uH3FfEl5z8QBvB6rPSYjSAxh+6EeTBIUddNXzYU1Etw1s3fSwgCfRGMwva4A7
KC0+b2/giCj2A2vUwmT2sqG+3pgw9McsAVYZ9dsJ1cqHHe05cBU+pMN0EJOCRt7K1kIRE6iPLiiW
cgHkm04TUZofHUk1XBViQK/iYwpooSM9nbG3vtxWWQln/ROuWNmnI/DxLf04QIT6T4ZzuhJfh8J4
egURUj4utPOgTmbxrhForzEpv8lQS4u9SyipAPvpCn6wdYhaylUqIEx9M1tUG7THZmSl/FtvWOMu
+OASV9f5d8Wz2bURlf7PhpwTyRyKsG2sMcPwNQso693WxqyCSdj0rk2sUiiS6paLAZtRzEi3P+Iz
ojyiVfMZz7yZMN4HPtg7TsJHafr6hiLgS+cnYDjAhN9qZdfsz5N1QgI5Oso+kj1/la9YSA43sz1V
q8OA42oSqHH0sFGlHReO5V2crOz+OwSsLGSRp/GdPBAnRqD62axiWOj1MTSYILisB/7Jsj5G3wVw
nmuCBP573CCe8gcxWVC0Y+7WYHF95NWsMV48auHimYDuXMDBz6O3H13UKSdine2bc25BjGvVWNNg
3LRrJIBkt+0HrS2pNFDmSQtRG3zTL7TL+MV9CjFTlgqviYq1LR4VtAr9hRtDlOl2JXduZjFRDxlh
ivuG5Z9Lxf4z7vSaEzOZEtgen0wo4kLcIcWzARIYQ/4rbY8Nr4nTaI1T5SwLUmbFPZpZ0YT24iYJ
GUfk9YeisNVQTh9OYbcrOxWMEqSzGYwR02HbB/70IJDKTpI8WAz5fsl0wQ1ELReswJ+VLDnpeffo
mWwmozLQKZf7yA+gREbm+pNrycqJSgd3RAmxYgfAdEzQl5ztMj3cGUgKf3wmddYB8iEElo2BlWQG
hIzOoiXQ/3irvrt8PvfsJ4jixpQdVAbgV3d7en2lnDeEqLt2uq+56Ika8xgZ2jXoIkYD3zVlEY5e
7fFOoor6pyql5zazWbBa2js194MbCi5LKNUJynqgmx4CT/n5xavk2FLk+hC77z3sF5ISEzqykIgU
PL0wn6TaLWg4x6K3W/C36CWwN2UZpxIPFxkHd3+yhHK4ZwUJqNVT7ES2hN2IAsctv9JfYugfiXjT
KTE2oUFwX5cfbm/lkqmm6x7ykP88zJ61HX2hNmfHXtsVC1X5PNtCirAgTWmB/VNxylXWMoVd4tq+
5qbQKMotKtYVHwImIGGoUXViesE6eCC1nSnO2Art5ABAE7Ui66U6whH3YG+EF7jCVLZfQehWt/7J
Tc+WGKJYgDQEVNaWEyJsugjDYjqJ3U8qS/l/I+2ttokAZ7h7LDXSb1XlVm0KFSq2cT8leVE+1m98
KzNWzc+2+7l3RCcThdcOfM58gDBo0apQuvmsXyYIuGgctb6wGEXBlpQlYap+gn57NLq0IFeu4QjV
O0qrZyT8nrglAqemNUwh07OSx9ordDJyzy7f1he8/dvOByK88J4115i1+4MeOdTEK6EuIlaBj97E
tvAGTC41swFat9WRafqPeVbPYHjBOlNayBPvmRZj2gegdOMw8Oe6SnjV22sPofiULg6E62/I2Cxs
gr+I5EoiGEIM2oF1V4wV6UA6S333bik4rgOL71g5H69w0qdsN09cIAYwqowv092ZFl4AYiKt8cqE
v0BfjWwYOFGjiumQkj+oViwJYFMCifTkCzjy/vtbnZu6g5AiKHaQnqGV8Ta5R/Ruu+4oO27tDLO+
khyJq8z7Zi54a4kd2gj22Xg0Eag5avlbLTXz/d2Zh9sL4TgPjIK4Ovq237apoOUdMCDw/9VPbJ9/
M9UzKuqB8xVfKSEHB227fAUjlEA8PG2qiPRPfR6/HpLwIN7u/L545CrXUEqhZfhgA4KVHxGu38K2
nEWjjO4QPckBtkhFwPPxfL13M645cNjhs8rd4gqgkbTIPefEOwAIhriK8Q9SEIy3A0PxZ+cTFSfM
sq8cPYvmhVST3js2ETHNM678iHMafmRcerLVGyE8fDcyf79OtPybYJKIdnBaYqgwhmSZv6H/mKmU
ovt8HqrpI+lYufbZfUpDkwoU1PmybqdArWzLcDOMhJDchYKOEax92HEhL2AcQ+BkEd3mRv0mdZQC
urinu6Z3C7xZcNCYkr0q//IA3gyd2pmmkBd4EO+EvaSC84o7vfDAR3z1k3tkWDUle/aCExZLFZ02
nUWxZFNPn1XH8wVcyFTgi5ZuyjV4nGTnTOa/SWNswg8nWEbj9m1R7MUQ7SoGHLwwBjPgB9Iw02qV
E5L239pactmgZmrxItjGfaIwNtsqcj8G23aa8ViTWADn3m21zq4dG3UyHFOBa5/o95HgKRkBN5SY
NCg/FIB8StO4hDq055t01A1uClHOjrU0sBxR9NSCu55x1hBM5NHy6eAQvVwpp9AXO4KS+Uns1Cy5
ecE2YKQrEUK4uOPPZu1rCOGXM23QQyN0V+vkPBemhvKg5I00FJdu5Esy/RZ2Fpf7YU9mEtNA4tSl
dG9HaYaDKt9mxeO7agmZ/UGvkwjDTQvoyQBJRyfx28q6jbyZAWkYHNou59S+EH73HAd+2x69RiPT
vInEmcrtWz9xU0YfrL0Mi+IfqrvY0xv/BWHBZLCITJC5nhNyNNxGOqjEynmbMk/NPXVAtI4VmEda
YJuITjPijdjOuK3/zSyna+eItope/vsWAivEWEzOWP+XqqryTNCf6NFF1P5NlNWMLMg9w0cn0Bd7
omJUlAuKwgRenk2YNKPQvYH1DFn2AEA0KX3CbciG4tkbLTH49wiw9sXuXwa9VLhI4Oci2t0qKhSe
GwclqpT01mQTwbcBxzFbjb5N9k7w/2AkC7Q6wAp/oou7oT92xCMDiN5klL9vUOlht253CmRVJKTg
/TD1CsotmIyI+tOIQBzeqpVZiAHuYqBwKvT+zCUvkMxwOV9TQtDkeDMOs8J1tOSpsR76UrtaQ+LL
AP0NI51MGQGAlFJ9GM7l6sVQoR/oM3iuF6S0hwDB2eldc6gxhGTZUxciUTmgBncPYgjY3YYDBGhK
WTQp2dq6f2mp9bJbIzFZ22sxFm4vFZQVpZ0KmriukX6EALgDDS3NzHeM7n/f3Fb7XlQYGlRiIJGC
Uaky3IoWDPiz4OacGfFcLXTGQoJ71FCfrU+HOj2auHCzQiJayprLV6PA2rUQBs1S+kw1VA/rY1M4
GCcqUhNpw2cayOSJln86dhL+J1QW7034PQo3YgSCFYF8mO0DOEa0vZ5MaCFJe1LMWDMfFUIn2IQL
+/fRuCR2dnMIEX1yRVE8JKHeQag3ZTC8L9qLCwNu/iJhJDbnkfXHglQQz+nIlDayFU/5YtDlJ2jg
UIy3TRLkGPrcWJzrlgJQ9oQm6qGTbDFPL36TLGKcxAchR0lbwx8YAZwzHHORqu6LXngXHd4OccTC
teQ8sfUmB1hDMc2+kfZqQwNdw8YhWeYOPsnnP261XpzjKhGRsa6hacbIeptCdstdPCKI4OVJhsiJ
Vk9XUTBGjjAHIZfdCsf4DgXhxezhH4lmNCRjNbSIMY6aEZ53Shn+XsQCFfIQ+urIKxDCeItXYSlJ
mJAN3wt5RDQG+/C1bZD0ipRHhD/v5yyTV0XHgDEchlZuujZI6YJbvpHKNP9rNzseN7AkvbNbQ/6w
alHcsjqtBik++8qBP+xanuel63jCImcXm05Z5s663VJ1/I7vZeLYbw1cxWbH9K14Oh7UBjgQEeAn
zq0XNqBni9zDZ+Y8E0dc0LGnnD07wlujDvGAl+9+lnYfPywTpQlHUYLzE5Xrwxgke3vHO4YRV3II
9cbZSVsXMH7OzAK+xZBAuhuMHQ5lOpRn2F0DQIV16lh8+LF5+asTYw79KJkP3ea9zIqIlWGS/wtg
V+ReidktezwoB2UkCKjQ5trNsy7X4siSCfnoVnS2Ok7x8sHZbDLXrdnpK2UprFOZYQGR122wwdxo
0f3DLgeBMynrqNDJsPxRjIN1gUZ73X8aq6XuMNR6mDTU3voAPWx9fxb0iHxnVuvtx03wdVsVle+v
q8qHMpbShUCZAb5LtzqgMBuRg1ZI/B02kEnZ39Jc64Qdh6bqpq92dAM//qgYVyX4ko1E6TK1kpmP
gQ/a5GkA6+Nn/FsDo/iZF0mvrZhBtejet3Sv7mRIocUK5UsIuZIvlgZ/fYWZ3QYjYv4VeA/UW83b
KCte63woA/h3ZJhv9Y4GnCUCZikXYVWlt1ZESM7DBtAZzRzSFU/unSSz9m0QJ1CRJEeg/rwMY8sf
SGBhZNXrerHzvGr4ccjKeZFjYLT90pwHmEP23hlrJC/DVKbV52IKSYrisgKnsfz0+EdrSB4hl4KT
FfOl/9o6IfrCgmmd5a02g2eivKh41yC13314mhsCcwRUjjm6Ndf6ytr9/2oSb5X2+e9enxL5wYsi
+buvg9Cxuj62caxaj/l3oxjaWGQyWIFBL9Yo1aeKRhzqhfXrfiC6b+59x+CyCnGI82NECl7DFgfe
SxggNbOIp4CoyAW6iIyIV3TMBpZmynx+amqOIlmVc0lsAkuMA7rUbfj79eWOHs7ACmTMXodrV8Oa
rdCCahtD2mWXxaPyB8a4Io5ncV6gzxTVfXqgj0Ly9i62M0Tfe7/BRKCs3mDK7SWgzY2FNwq9Mf4R
CXxi0T0uL3KvcpMcSkdaEEUeyV/Q+HNHuHdyt9DASLnP3vGnuHgT+LIOl1KtRQoCpF5/TZAvXgV9
Y6uxj+XdbFCvxxBZkowDTRHvwVRhwuXRc4bIQit1YZnUjXPmjdk5aPbUXF+Ct9DxPuUCveFir09e
3mvxbEQmqQfIthN0A0LzMA+xD3UvzMNnqUSBEAjn6jywOMzbi9PzUh6cK99WOCTIUkfRvGiO16yd
ID4/uJ0chgl5GhWYMItEFkjnt1EU8JVdgar2mb1E3A2VegTjNTSsNo2Bg4LbClhD6gpNuPMji8ZH
1EdKDYN/MEbmws89QyofebTmfpQMVN16sGVYptLg8SZFzqrXZk/n/mQ10GWp7P8QlWgbMbGgjhvi
0ZlkDj6pDvRYobx6nshXGgAcB9fV38W5eaSBlEvouOL7e2c1RidVLheMRN07iT/OSmF4wg6cT4NC
5NR8Bl2Fy8a5PnrLwLQruZv5au+S5mLBm2wXoBLZG71QOCIGCqCrD8h1MoYAbepBwHwKhyfHqPPz
F/LX2PeASHEsza7azWKVadeJYLgDwdzm9tkf0VWWhr3XphslxedMJ2U0jkskVfFa8enLRVZrVjZQ
1L+IWgzNpOnyjLJWVx2Kzma3QcBj4yvNbfSjDE4qJ+T3QFXp2SeqT3aYfplbWMMQ43kmU929qUFX
ZmJxSNMmbLf0qkkxPeoDaiWk9lay6gk74j64AvMHHc1uaszFB9QUervYXqW6EpavA7664+bRZ4gL
sFIwdKRnhMfRCxRkg9CE19vwXiRy45hWkS+xy/CXHn4YcNRmCqzQt/oYSQudNRxb30oKPgP6Niai
Een2rszeWXZullLGGo8139tL+NKUbDZW5roMUCOZvm1tmZcHpV35gQPbXb3Kkh2DD/HVcVfx2qm6
h4Nj576zr7dvxP7v/dayYmnzwJ3Is05GS9WSiK6lfBAbRldE/CLibs6QyQluivd2giFDbrUkQrrA
myz2PRgPys6ZdThf6MvjV2WBQqn9rGLmR8YVyHkD0yvr5jEWJZOZlHEntijDL5+zIRBTEG2qWkhO
zLHpZegG95k6zVEv27LDID6xnme0eAV1UA4RkkJ2IUxmiw8ie+ldXdNk40zSb+tTH/H2+jYcKJkh
spc3gKJf42gjhoBXLMuP3bhpItmsCO/MECr1Ld24Jg9vZ46hcNP1NkL0yukVHSrAUz3oo/STvpvd
80i03zOp8KN8kBjZDIZds4afYarMZVRUxZHgEHXjXEDgi5LPGt/saGTFWvh7qDraV71c/dwroAwy
TvhO4IQJp3Lgc2qjSpsAF2qD7YQzQm1EgUJJeQs975DUwTs5kK4AZvPCy/MK8umDi0TSy0Cz+fpa
7uhxihJ1InL+8xgKyuDIZtz9RSTiFZ2CTKX0Z1XrPx3Hv8XBhH+piALUMzuPvl8jWGSRvQEmmxdZ
svkiMGldfKjqenmLND8pJqYp2lt09U/WDhLTgYJb5Sctz+3zSo5BdKdmrThW4OWw70FQJrIW6L+r
XzOCuclmV6tDr5fj0qDrMNm5F1VlrivawyQs5xBcQ0pf8z/yY/aKYwMyL+nCmY7gFbEDCxLlumfa
2Q64E92Q7mp9OKWctAqkU6BAgidOEACfKjxrlINQVVo2u7QoU2qVKW2EN5tveOKQK9DRDVHTyjsq
GqKTT9IZZKf6n0znSfwF4p+Y9ZWB2zQhjsSSBP2oLUD/91e523yVF0BCcc68/2ygj8xUzcM3WNMp
U9nSexJKSt8vWJONjscqfWioZ5cRaSl24n079CG0e7/AGMss+2BqTQJnkB0CKDaVsWO+JnRSTnIZ
JMdiNUXV8yqnS29n+GeOnSWFWSwEhYyW0o+bDVAEj5OAh8LmKNeqji3HAI1bdKxaynejLSD8j9Cr
mAcvmdy3JugQ9tJ6XtE4A46ob8Fw2+b0NA7Y4F2Z1ZrJUmLm000xTQlyRIHS8Tzhm9b5wd29XJCw
nckr9m1PohZUwhfYPX815Yu7TlJrJxeqyLh8DNMQVHVJtZ/ROuwy5r8bW4uqQZRUT03Y2udcDDt5
0TMJfyL4U2wUICHRyvY5ABc/3B1+T5lreAJEqFuPUAVHmSAazK1cdJUEZSdGpZB+q1L6j7QU+WVo
tEU0NIXDH8rHMlZcEGU0qf0l0PMhhc8OQJfyZLvDye2Egn85R5kEjRnjF/IoK1QzYhbLtdVMeO8a
rmzeWisKGemyuoeYT+P4Fm8Kod5jnm3n7KDgTeM064oZVPqYyVqzlNaxs0fdjhzxwxoW8USph9yh
nrbVIcmt1n5H5cjbmcUaN8BVIpqckJ1feOb198NaHme8Fu58vS/6OlyVEKoZuqUxLGbwqbCwhJdE
Bf18RT4DiZD5vAcXayAcv6QSwhXVyRuRPU+bCPR6VSQ6TcunqZK9PREsZTePJHhFM67atx/JNi9O
zMzaMYLnXGn5IMjhI2uZEq7upznPX8dox1BQ6PfmyOjl/Mv76j3i5tTE0KMZS806p2rP0LDEErxd
sLQ9eBLwxMWBbOVEpA9hhz51BZW60wDM7q2r6GM1DhXfml6TiyRdssP0nth7qAre/Z8H/aagwmGF
fHNNyjxae9kbWPemg59RhucUS1psTSgeyV0hSC9V9j337XHoCNkTnGJcLN7eHzoTo3h35a3/O032
PFcZ+3J1KgeIBaobKD5JiSYzOpn8gHueFGAWk/LS5+QyscLXkkyyiLHT1ipNrBXBKLzckaT4atq0
Q+mTdiaKEzs8VQxhxX6kCLiZI7j638KBhHIxxFGM3pzgRqEWwAienGw7nkyL7S9AbvJfmrWEvkGa
fWQ4kMyhLV2kgk2BqZ1rrvonYE+xPqh4J7JtooPbcb3e7NMVu7qlIzyN08090aodzn3RmYYT3NHE
4u05g3mLj7fJUQq9t6D9MQnDfQThMS8kSS1zNDO5WCQfTMI6jHqZS1NQw+IeRRdbYzJnyf94xTl9
U0mMPfO4U0OfpQZPesLLxYO/C4sFrvBuEiahhsvaRP9RNG6GBXrflONM6b5p90DvxWz08PX1JeDw
LGHiN7TY4KTc5Fuvh0W1W5Z4RsZtJt6DR/nXVfm4NXT2yVJ8vOxk8j93gPXzB4qpE3o9BkSLoFvK
QtKIidzJ2msF8jOvhmezndRTd2paTK8vtHl6tlX7jNviXiv36NsQRW/fH+qL/WpjkyH40Vod2B16
R3J9diSAkGBZA1ogRsHCyunMqEP9TjCz58urCyRAyuKewXX/8knGSuR7mvxfhABM2sno9uQUMSCa
P59nHr7D+cVJecYVWvYPvzZhnfuJM/uFvHeePy3JyqAS+dBOFirK39Z7syJvuQU7CpiU21UiniHg
8WIuHm8PMZexqm8MyzzRo7P1CxWQkWybE0ZLjlvrOANf/JKgJL+Kp7Pb4TQeiamlAn0CRmIxBSgs
KyOFbW9M7QoXwxB0aQUB11nYY+wRilzzHpIzQCJdu/Rsx65MhlLKT1EaiyKWxlGo27E7raId2YxN
CMPL6tk2KUE90OhCrHVKZU3o/f9MZC8lNAG55xMfXnZy/cM8Q851kJXF0GoUboz80WYCcBiLmwu4
Wal317n53kGPWpGS6kjrwiuuHXZ9BDFZsjdPbkBRfwuw99UbyLcR16V94hJtZ/UnqbhqLPn6de4r
1v2ycAmzxdMuIxTJMH+XWA0Ho4MsxVOPEQzZ8jUKF++G6/EVXgB5BBUjDXl0jNdM6AJcI/e+Kw3v
Rq+OsJVsjTeM0fI0rrcLJR4ZM2e6jpd3IkXrWDw22qee7GFFgfMdjZtJsX8FccPCCZHzCaaN+EiC
hFiAta4q59V1fJwG/WzPJmm+qXVyW9r3ZPxxzBxt2nIpgEm9wKyxFC+ECZwdD+iKYMdc6FELmUoS
nUqBMZkc3Ky+OOQkUBE+Sj1hCbJ32gx2tyGeVcLFvfrxqhCDFCxDBuMMgKx1/qqEQpp14AtNf+8X
4iK0s2HnR04s9Gs8qa6EIHSdAvzUWQnKCOrfB3Mnl2TIUY/yZMW3qwie67m4lm2RtbQPvM6ryiBW
1OWMNcEOGQld5loeaWm/0Z7Okl4KrnD8I4J3m2dgUvs9NjSQPDFHCYrZSjVwCliEjzt6rMK0OwQx
Fmfa/dRj6nuaRumK1PyekWLjB3tGf9D/RoAjTIMvvn36fZqabkECycgl3f0StAaM7G54ETaZXstE
adQ2ScgpYgneCew1vq70Ze2hFSk4ZcAt8u9DHbSa7IYFBTu9OSe5sgCgvOx4EuUIUgAeZ9eXKIVn
kGOB6GXRq3V2XXDwoI322PFrhc6QG968Bl0H367BWlXIldow+je5RA1W5gPL6HwbjtNJIaLFrHU5
TNSVxhNzYKPKqgR69/tIUX2Bw9lTInPzcEe/nIFlAbvt041mMVvEsr3pIkrVqA0J6fZU5Z83OT5r
eMD4uvqs/bVvvB3EKCYjgeKluHRzes2qZ/0X07bDTznMcapeyQimqse9V/xJelJuSkT8rSTGL1Mn
LsFcWQKM4AArMztVHIwxu7ZKSTjVeeL1DbU8S05WeqJEUVQFHivPylWvDjPUristjAvn8Pu9WKHF
twVGdDjNvM2OMHF7EQrKEJ9VdM61uEIpNvBKW+Si5m/gppA+Zz+i7pgEXt/Z2DD8FjjmtmzReSo/
I3NDUFXsRgPqdtcKcuNddLL49vAzbbtaGCqBxTpawJMXhEGvvzDta3RlpbUxzbFo7iX1zhHR3vfE
njcqO6Q95prF49YkxbTudPSebdHzaz72kI4L1A7MD82Piu+Nlm/DCKRRDBQxSruphOoUo/W2dMrT
rkLgKxow+F2KHmpSrT4/qH9jUoHtZXZmWu0LXluqOMt0+vS26v+Z6MIgZIwDFcYanMoCV/VSdbOX
Tn4imNwU3AL8KxHtodbbDgl6zeElZAoiUrWxFV8Zx+Dw0pJc1vykpUTTbrfPGc9+FDl4GM/j98/7
Qtt0LBMe4guAH7Pk1SkpvGqekIDMPapDU1QIulOKdO8Nd3NcXx6Yy6EIpltIWbVqf9h/oft3q0vB
Pw7xN3YzB75pOaxhtyNA9oX1TKl2iGKdFP4x9rpcp99eT/oCDKXdqGI/Vf205Uhi6DWqRSwxU32C
xvv5NGZGeDghOWcc+gmfSPFKteNS19RiEhpU3fQV4Y5R3rvEKBtBbU/J8aO6B4HP1H+CqSQjhV5H
2jsZs2alhZQxE29szrjz4p3hKngFP470/2zt37CRq0IPjvA6CsqoS0qTuGgWZDAEhwTIuhjhQip3
W6pCl8wi/yH1u8PpFqkycWmYIH7ZJSOY0SdG3z7sUJQZj6d+hR8qeM3Z9PCnbOHLwvbBLUkhKs0T
2Iu/nv3w6D0emkL/i0WMBt5s/3qC4iD93C8eANaYL/n7NsXRK3yv9o6ut6J2xePQCpeegrJ5K9dv
JEOdoGghroZlFs3DdWBntPP1hQ4/pY7OB0IWEpztjltV3VN3yRop3FuJWzqwdPEavQznn2YoE51F
+ql8Yv8eR4YEGKeJAhnlAOfwTTmFmsYTBwquhZxB8UEO+ILtBtuiB0VYAZoG5n/ixLTrvG/sdGMY
17CZlk5ToPB5lebbeU2c2X9iSg0J6QPMdxCSYCmlqF3IP52qks8dgyilQz2UV1BmJa7AqO5c1Apw
no5V39ikoA8bWROu8jyXWPJXOCVvrYISD1iwHMLEgroZMp26t1RQwjzQrZeVNSlu1ssjr39gE27X
5a6a/1cDmYaSTMY13zrcvfQLvb3UBesYDGwcfaFwx43lkgMsDXab49l7QGgE0stuVAduwG5cci3L
R4/yNv4hgwF1v7jFrpbHg6vLxVWSnE180HkKNmYy3yuWfofStpbEOh/UbvhjDWt5DlogVUZgcSrj
0LKhVmbZnUUcpmZ3l5pPTsyGxKRnTM3IfSH0V+FUy/AQ5egL3o8svPCLyAzr2voSuVmOmiwpVIDF
q13zLPBCZ4cntNpUTroJGGUCBB0CBu/kyO0rDEtxv8ElGfObB1R+z89V4Itj6t/5Yo8dCgJFgMnO
ywPGvuvG/Wna6anyye0RMh4vPU5IN41W/2Ofmpmc+GdkFH6Tb0ycwlM9oEHQmlsQUr8CS/3g103R
11tMocs3oW0eo94rTGOZTLa6o8jzLsq5ZEOvzfIwAkcVo4FA5slBJafdvyN4tXXjoZZMHGV1opWB
SrSkKKzyS16UgajcinBwOJyiJPnwVN6OBgeKKIsFlPPYARgMPkqMp6jokpTfEgqcYfkt8/8N1QRz
xfsAMwbZbphE5ZMguPjjVQhgQFHJE1wg5L866venv8tDtvoYr5f9rpPUEG6PPGtBIa+mxnGvZqpF
TMteWNwF51JQ2iBaYntZ0LhXFcCOYpY51WqA3IxstjIYnTjFn/uXbEFlkm8Jh2cOg+WU4J/SHYk3
zYG4ddY0Gtu6/BtIT9bzWWjdvrV36P0v4zv5LMvBVqEAgZK9ZtuCvblG2aeGviDtcXZGs4h335HN
pjinWzYnlJ5Zf3ZYin1R0gX6uQSGCqUBB8kXFf/gIQQbn+O4ZbxoPs78vzrYpB3cuhCjsOsTSCxy
awVgp1WspLFZe5W7JnZqqw+Md3rmJNKh80wb5tAld/Ty54kJExZ+swoXLBXIO+vY5wCMLtEC1qP0
IKEDL5o+Clsj+d0mwpvL/N63hHaaW7rmF2yBVNUjj+M7Q6/sp2PCxJc4T7cPNO3hOam1A5XDQLfg
MG4lw1QWyIagvBNKsc2aUZ8UGLDH9YWxP+rMP3bHiiLUCtiyJChDE90XzCQWMCOPyIgIzRkIjSUM
/32ZNhMTc3NyOru1WdVG4h8VGVIxixyfO/BQkKMumUf6UCIMDVGs6DPgKbgfrQlBSwi+75A8VJUc
oeqQoPDUdHWfZu7oQijBZpW5jVBXoaooQa/dULbb2hsWL9Lk+HzWTeCEPt05rMKhanbSu1UIDuiI
0FImlfkOuD/2l0ySW64f3/C/zeKT2gZY6ytLjSsT1L6WwbwJDoBQTdvSQMURYsvy3Ig/nlwIPTTy
BceH+gugfiHeH6Qh0VSbSu6EMbxXY7ow6f03htFDgn3MCAuuJrZ2Tl0KWQJNvHOMJosZ9k5Qz1TA
zA5V4QIAyR2D8YRkaMj2C7HE80xagBBHQLl6xhAnfajRu828HPwZhffxTcZgPQjcP09Oc3wjDF9l
SagQQki314H5sKcoqoj7QALqrQ9IuvFMhKPsPhKXqk2Z5I3kXMAILXwe5WcP/MsEMN65H78jOT2o
G+UhTyk9ktscYITrphPTNuxQln5zaG7ByzhcEfsPONXZi6wLRROsBhaYzc1R9gdSbPqkHrgt06TA
rv85FbwMC2+D0wUPoYEcpznhrZujgYpSJCguUx6Tgb70nTPonwAiVFXNcOSCR83kduYvIhgKvbTt
ROnH0Rxt2ThAt9C7nbURvUt10RTYP0DOOXjkRzZzK6qUOSV8wdUzHIehOTZUxaPlzOBN6qFFdlbK
BNgNH+oCwrtqQ12yrIJCGFqw0t/9NecHPVe1OpKBiaeK3u4+8fHL8mOXLV2Ghc6LzcK6xYbDUsUo
sgNgL00xkYyWosgKySSkCERyfQ7aLLq8M+gxBFB2NSO6OFaENRtmc6oKrT707a1+Ee5VjLOeJ/SF
0tMTEj68Udpn/zBdEZ1jZSQ2o+vKW6EB/kF0QozOPA4GpX+GcSX49T1tIoT/ltTreXCtomRzqNui
YHYiVPv/hnc4gPvqIj8mgtkRq91u20toBqAngizhQn2s4kYt45dE7nogiWwu1cvj6LBMHfeEa7OG
WWXfyLEQdDAsg/7heKQ/v5bCqs9KRYMuDP1tGoJhRLljB5OBbo/Qtz2DlOG3phfZx38nmINhPysG
L/Qw2ZB4i/C1DjbXoFpPlrhLJuzwaZ5AUyA5+HgWNudVfBunG2mQzt1/ekVm5KtT4n4N3DeNvE2n
ErkjIcIOZRoCz1GPlCrJyuqp0tDeHRJqYzjDwroY9qXoGV6FbK5IWe22O8DO7sCTmmYHz/KZVCGe
TE+Y/HToQ8Nfaak7ZmvIbVrP2iXwS0QibPonb6EnbFSpPlgEd3TMtAT+l49RNc26azi3ZGYG5uFc
MG+f9HLvwJrbWPnekA8kKx2qMp18xddO80WctLy+GJg+53Ptkv9dXDQQu49NQscAhVPJ3ddb5Cmo
FI5JUTTr4pPgF14SAogjGRjM3LTzl9nxn7usmoeerxfRkkmN44rpQs4CMoR776Q9QTe9SCEUx93p
OafigDj8fh9HFGyYdvQVZH3UEgHH1Qu835xJ3Ru+CZoagvAf2ga4UGlsKNzWI7Is9YuK/eqzlfOd
52YVajWO3i3YOEBiVzFXxwDTsq+XbC91nuFY2ayWjPZ4Il9zLy/LxNxydh6IiRNqOgfCaJGAmeKM
uGs1vhe/JcrpXhFgF+ElsNPLguzNA35wWFjf8X3gIwIsGW+JBw5B23UQr1Z5aRCGfCzhlYkDgdCi
Alcwg2PknNNV5GAuNjMTTRRVXXRR3KQCZNOaqTEs3JkEdHlKx5qQNpVV5sK6ruOGd9YZkeRn/V26
EK8+f0wRk0YfhK8/jJx3rf8Aj0JSKrK/sV3nyRn3UbL8eOPE/TGvrrM936pXldhIAlV4afI5/7Oh
jmDYXm5nQDAE5u36BbCniWbWZ/PNJmkHi27hEZzNu/sTO2T63fHHchLBpfY8VJlcn7wg2ABO4fo5
EF1vjBUtchMPtvG/4tXCCJic4FycNACgi0iXSe+mTcp1nfw+1LrzkYt6AsXPJ5B55xMttnngx7ME
0frsF7vs1BwC4dPruGj/UgxD1t43JlfdsSlObEg9STzo3O8kM6+R98SNoKhg4qIWWE7fq5uirMVE
ygM9SuuZsUnJOo5pjBAPqgMVNyLVbcKTzEoGSg2NVZrZA9EFEZB/veaMWX5jb/NlQmdeCzmR8VMp
eM3Z5n55qe0Ym2O9asI6H+Da2acGBcWTM+YVrpKtCII51p3+fxLS+bknElGUPhvZp3GSaDOZPQxE
efJcpj4MqmxdtPw784E4Zo4OLoM2kNBIQV5w3uwdNsAlSchPX+MHkkirk78syaBHYaxQTRHeIufx
Vy0NpKzHziJWXXyYg1JZPhJ3vRm1aKiAapVIDqtgwFpi4lHHqUU1jEZQXe80e8nb6FSkdxCHhqk2
p+AWsloDCes5XWlUzPi0I9m49UqKQcx6UmXy+puLeqETtU11kBHpmAgnB0dPWcik/uVf+IOKehHc
MfYE9pHyMos8uBDpO36yJxNzsQPbNE4+KUw3SOxRlMJEU2xARQvyrAUA5VlbEaFFrZru4f5wr1W0
SfrGAsgu+F1joywjNgBCm9Jtns6JfZPcDBB0yVs7WcMMd2CuLEj/Ow8Ije2uNSKJteVklCy16fbr
wokzhGYNSpShDVbtlRQP5oeQ2y6LL6QvXNZ5jUEPE5buVIb5r2FksCch4Y2lFPot5is8/zMOVCUk
rXFKcDKWKrizVmSuQ4cpzPq3ONnRo1VsEIeYJfPCzrDvYUqWHP8eIBJhn0OIhHtp/Rw2wVsjTSBB
eBVpKccW/KX4Ck8sJAvPeFUp4jG/jaOQLjMtrpHe4Io/qxik5bxTBPr5DvE71qSAR5CaoW2/OYRs
2OdRl+D87W72u5uhDkFeI8MmAWQrENsbPnJ7ksvfwCaPCz34gXajbf1t8Vnf6YMh1Ei4iLnpGb82
JxnEezyFeFWwsXrPs+VFcZIroyMSCoch5EcQhNPLOVF70dQhN2E8XWq3vZuN6khJxQgXqV0Imtqn
rOcxcXGRJXRBzzlDyzfXLWUiIDNb+QWlaIF7AhSwivjdXwgDO9LQUdyFgi8nRjgwAJ0Vk+W2k/HK
TQYU9UoZAQmkAKlGfRX+lwqnu2UDtkS6bTnCgo/v1IfXvqxnt9oXeIreoVYdYlsDg1XJeGKcHHzG
Spq/Vf/2Pe6pvGvIPf1uOo2TF5GbALCXPx0GPslsZaeHJ8W79VjE4CXfta8h+0LDnp3gYCuJPYxF
epnWqDLLH4qkFmr0k6zljqOPxC675tzdfJRInxVbrxp/EZxYRpe8b4YOZ37SinALXlqDg3snz+4Z
EL9vJ4ArTgOlWDmo1RHy3HuLjioiiJdgQZCJ3aPtzivqQRb+pinvejhVSzNUtdBe0Pj0nmDah0GL
We8CO2KVcB6196/V+51YOIf+MOkMsVANVQYQ+oDYmSh+lJFJ95QyV0EAyNZ83K5THOECg9pqSgTo
j1vG5z9E7ES1Ik9xv5CWYkHEB17FRhl9ps+eIlCQPYgkoLtebzT5tjy/IX0ftlOZO3Wr+n1rXYfd
1GRqbVg0H2hgAIemW94cWMyutB0ax/Jv3RewL0umxMpA1OugYwtxyMmk6xxCB4s0akpwKlubOIAU
CY8uNQT7QVrbPYT6ivyPsvN1+lEEgI0R41U9ivaP1+B7bGYL4ecohUIo/YSCTpymKpTXCJx/HVS2
qAETHbQd3rfP0dYe+xXPTHFXN0ZHyBG4j4NWN7V6jYcNFSJUWL3BABJg/n3fVfp4RkcLvJbTL69y
/JX1DbQL6Swy4QhiiSp/9iftJYK1/VFFRf9QC5cQut6EEX/KekyjULOXp/wNJNj8MH7rh/ATw4+O
ylRZysFKFORMkW9pTuRG5Uz2wjkHpTa+AqJjSQmGLJAmx/dHizXdXKnDoJtbbPRd4KzOUbEMJ5MI
mmCnv7ypcSkSTDZTQlT8zfql10+tTjhcy7BSEMDZIzlaBmsQhO46ctSpus0dVK3Kit9rrtwdYvbU
Xz+eD7Yq7N4177llHBUrR5HpMFa4d2yYnMzeTxqMBO7mk3EX8T5i45DTTqcJzFr7sli3qS3mzxZe
TVTzkB70InFb3/9b1R1c63bAsedmf/CYEM/2n5L1nYMzCJf8Hrz+CNZFf81uv4yON+72dzlZEvoA
SCH9e2KtWvUVj50fxiju1gQQPGDMLyja8Vw20J1uYMOJl5oVnooFL0nAg5ZsUdYoQUQTit8a8PDi
0tFkCanWYHWLk5AitEIL7fUo0zYbUO1wNzhBUazp37h5T6+Xo5ie69RTBlP2k2MIww9FKSVy4KHn
MNTXiw/wRCk/T1iLD03IuaMLF8uk+uSr5ltFmaKGZ8YNBASFJ/dtNcIT1W1cql5jJrAAZanBg4yo
b8582gCBTknwHQhIwC7ixIOsAc3I0CkWfAZB5Wm6GBdKxxUIxJFB6XFxM80h+0e2cuE2AB9fvrPB
jaf6GeAiZ/KUlje0x261gf+2Lu1gKtp+oq6TzE5QaIH3AqWjcslPFcPoKzMILS5Me2naFqXipIz8
BpZHWni42UYG/tWrtYfpYEfj578CrZAQUitBczqYswLfg3j/aye6ClBICCDLKrTRdYM9h0sO0kdH
KQ+MpjTW2dqirFdHkGRGm1WGXADBFD06gT/PWQbWPC/atpSoQL2ZDcpOwLZiLkmIhrLmz9EQ5Akf
DEic+KduaibULV+BI/7Z0kEYOjBf5+jms3YYBZXCrTE9TXfQCLlmvU/KKhUV89rrpeSC2kj0OORg
jUfa84sN3JoA4H6jIwK40THNQAGWYuHv4Nc4Vw69TnxUujPWCAZXeX+ZnwYUIs4YJ1LYHLNp8WGe
uq8n7SN4zEsOvXzOYI+KpXvaJXSgjeKsYXbxkSH84SviGsyO12GMm+vrxzBMr3Y3nXshNabiyayL
dlymTTXDCDQG7mtPrAdMj+O4xJtbPTSz+XfnKlZG4doq1f8kQjqn/p0eMGdVbd2oQMgkaGamP1We
DOdAfEHbvb7a8OqhLrLKRxMOI3dhpc0ITuQBq5/O3sDiPQl0ldawg1FpISXS1uU1NwPdNV5YVxAC
I0XsRxH8Q5qPYiiXAtl7s/AAdjE3U138RpSkVr8jt6Qr+yFJ9iD1VM5M8TqKA/5xba+yhWmNSWWn
3iHjUPAxPcTNhZgEvjkbOCEjLLcoISrePJ+nGsNbk9IGYsIaZidyfsgk7f5Gcf4g1FeRZJoQYMCR
XmzB5MKtGyU5CnoEdTD1564iakrCLnd9frgGa5B+8l26q9BmPenQAx6MZRK3MqGpabMq6UERRd1C
vBY+SajoYraJvSOUe93n//PQFeu12BW5O0Tngd5g7WkNPFQR0U6pzn+/xr+KNbWMx71dsmxbau1m
ROAdbPeCUIrq8vCrWi0PhHu8uuVb2lZirAqotTYAbwV+mdVkijPNEnEwYVbHNrCpRoXc9dbMiCz2
x8yW5YB/ZskflDnRMi8MlgvWVE27EI3coIuw1R4L7ohLQ50rz0IyRGBAX7L98J/iZbR4U3p5JtYi
dwx1m5CW9hPfmpL5w19ZCrKrol80ZpUhsS5U0z/nnxmCU95OrtW4QeDT9n/U+O7gPpyQ4W/XdS52
6D1Hn677xyuUpRySPePl12VVQOtBV0i0WCs5RQeV41cMVp9jfvP27z75jINRmXqrpfdyz90yt0mf
GPiyMepsyCQj0tnbC1ugtCsqWn0/zad7eofZ6bbfuFOhTFJ82TCn9GdIWtmymWqaK21rWld4cNOV
BNZEk43NyKs4Cr72uzYmtvEKNBs5FNTQjKhMi8CNN9JWQqSyr55bRJ+dsSTrSb/m89UVgyAOO9ZN
zjl/ZoNgvLrlai5xR6NHQ0JxAx+cQ/DQ0pjRZkXJicXKa5grUd3wPtU8x1/6TBwZDkuRUYa7dviY
6Z9CstbaEdKNP+jTpAy7dS+Wey4KpqJUB7yfYFQo8vr+q7QPPP7/CquwwvpePRMivTYrrvtf4P3b
NuFLf3XHVvdoiCqrSrgguE0QTcrQ3o442teCqjrX/MezvVQw9ELaDwnvMGvP1cJkRzowozGCUBqM
rO4ENprExsocOJ6mpy5onAXSLldNaSGimgUhJUGsdNPrcNRmfkv3xZrmxj5J/ItLCh96NXo19ZDL
ctACYa3wVMoo4nSMgwGfzIK9+SfHBwmadGIgPfHXZuzHyAG/rStnuEZMkJ3ubA1ilcUsrTYtskhG
jcBdmaSprwRhPnVPJH6QbFZjZ1SrlkJk5z04jMiX3ayZInbVW0JerQYgr291rKFvIVniNYSagB/R
k9Jna3nd435rQgLHaepwHR2ZpEPyOSSsfHA5PUhOxEAx19mSN+Aix5u7gA3il/AioSJJeHy8mdAJ
axQCvoaPMVtpoRR+HI/pQWmxtaYu/hyU2sa0Ere6h8DomaYjX5HRzRiuXU4iqcP1XT32v5A3W1Hg
8vtSXFW0pYeA7Cr3WL07/gb3ZOzIBtx2HtBBDPFjldhb0DYiWXbxXCX3GOe/lKVBa40JS2ehDgLO
+9r0NhUi2Ao6m9vnn/+T5COPhKjmO6eUjY5TUNGnt31TDpNps4cUpdNuBGetXn6nb/4CKRpYqR5a
G90kAO2ZpG+1jq3Ct23kw8zaXRXyUPKjAOqSnUOSAuCE0gvY8L5ASaBbskVbeBpiC5sp4ZKa+bx8
pS9fz1ip/TQyyR0n6Fi+hnS2AYTwpuzlbTC7B/f7MA6qyQyiV3f1j9/tvAMFd8pOYsjxYQychKuj
caFCscIUc190LGN4frTr+ZS97jjPgVPbf3G2QIixDpkAmiaxYTiyjcxKcuauTE0/wYjxaEWX4wpx
OuHo1OqNjNKoFu00UkibGRn6BTIGD19nVEy0c5SjYIudy2DgQrChJH8/pC+fliY5D2IYZO2FFnQ4
2tveYsLrNwwSvISDHWqpqTcKvHATFDshpwhYwJTt7eAcQPaXZEBjGOW6I5l1U0guVs4IWzk9PgfG
AzduADB2nFle9t8uxmYdSGZUNdCx5D70T5PN57b8mKZ8P/6VdHNHmXAgpKbTt6jjp7tnI03ODX+4
TVA/YbeLQBx4pqylZvrc3gpX0D4+K3ET4f0+pzLrUm5JwqIxcU9PTUqd7tcuOZ0KPG8q5KoUogw4
Jmo0Os12AP2LGuzH/mtjQRI15UVIVLXlRtW/Iuxhd7j9VJeIaXrqc5JR7NVbaVS6e3DnPtUjDh0C
7qbpajBfPYCAxl/LvkdcGpGv1Lnwn3vB0kUHdNY6TfOxTj4gbksU2Ntybmmgt2li4hsNuITsk2lJ
PZiM/NvDH3XGWrcsZPNMsugIN+NtqjLTcj2KIRqsSeg/DujLr0d8tw2Zn9kP0fEMANJquIe0Gpp3
UaTPlL/OtT6mp6esbrG+l0momZ/5ou+5wUNSIA1pa0i/UtJDmv5FBdG3FVpba3yfR98l2cSZo8z2
nL9qk/J8jkB0pviBnoW3ifWlNFGg17kwTNXngl5XKAk8BHueaJyDM/KzAsx+nrk9ulFpbhC7ijhi
j1v0H+AvKyNXBa6HAzacnETXNTIKed4KVTz+3Pg5JqbePUN7yDevkPNm+6Praa+4PeySTcPfr+5r
PDNHh4HWVIC+eb9njM+VsMhaZE6qNOp8hCA5/7wkcviThRg5/zzetBCS6IYIiXByxlslc99V3ARX
Dn6+/NXm3Ep2es4DfrnkIpzepBc+L6pr3+2cyWGjzTao7hL0oxEBhWW8CcOvLQsaPbFiiA0NDe4i
oc2z8g8y6FB5P5ScqqF7WdFx12/toGJiROza7GGhYC4Q3OePIt0WDxgMTpawhckH+GboZ1sPrSdM
GUMiH6XyHrl2hoqZIL4QYHv/CCGRa1Bxq0IviqwPxtYyRK42DQx1ctevBRCO0M6cvVG7mEl+IAcW
1hxyEcUesJKu+PF8dooetfs28DzluBjfBtiT1GPgsHGN1kKnh5FLijTmfWRrDkkr1uZ2CrOFTUvc
vgl3M4auJRP0RbTgf1R7Shi1jl6iJNJk3/UIOqP+i86/kU/is6oErDByoSoJ1VigUesf7zyx9Pl0
jAHslIEIhuwVFN9yh8A8sY+Q6fmeWIvkR/UO5Qbj9Bid4TZpM4tK3NUGKCD7HT4x1kRNldaVDyHB
f5voeWQvcA4ejhFp9CvlJmUBPKo84cAvkmZb++PKQpcO3hYuzzfcUj06rN9rWXejNwz1egwVYJvW
+7XkAnOyzcr/alB4cPqQVarvtBckK+QqS9H3wZ5otGS3n818FXH6iaiANlYN2KDU6qNWROxZkWik
G0wjt1jDevyafrjuD6mZCV0TPri36xXcMSkZMAvc9Uayen8KWfe/Uxm9pV79i+9bfoyEALZ/sVLd
1j06xnPIk+jBmQyScbtuaFM3oxlVyMH9pTHLQLMRZZH8R2NrvzxAqXtpOveEhqdN6kwlYe0SI4VV
l0vg/ubdUUBSekcaCqqAEqZxToZlIjrkfvGslC4kh2BgYwOgLZEXtrQm1gua598bowz3N2ck7bvT
GU5oegpaMu50WqczRC6SLsjzC3Tov67XROWf0O/nh/aMNMAGNEh3uMq8JJPxbOrMM7kZM3ronSRQ
OLCiK6RqihKq0FT2rlUwVikAVfpSS5ij2ec6YGa3OR0fCBj7h2+pjKSq1QNKu1exjByIEijm54kX
wvsHLEA/m+LqI8cF+7nOgVN0DVau39cMRbVdNf8C5hiFp7CUBzY9hY+wNCpCUovkpqaFceqtOfjR
4mpCIccQn0YbFgCCsKFKGYw2LlWp8VLYcJ1/eVKtHhvQ7Hf5yfKeuJRVMpL6c9EaFy7r+i8ugCek
lo0ULWuefZ34gGD5yS0kykDEQEK4GfmzDf+hSOKKSYKsA31v/6mwkbA7q18G6kOXIpLFFYFIHxWZ
p7ylkxSSaOv9YWS2oqbvshBSxB8bsCm6FwYgY/Yirg4+xXXIE+68tFMn7MWNOsEDBt5It1QvfQy6
FD7fYlgK7V7l2X+dUOiczfKwiNXECWb5qfV4L+OmN4yCKyIqiup2sKKm4lJWtM/JRwlq8fXD7+iS
KmSnK6GVZKBqB6xwYX7UY3eXW9bFpywwYi0RihQ2qrJNMjdiCPB1EX0hMP0UPXKcwKRACiZ9zjcM
k9RRawYK36AlBq2WeiXaTnJrrpLstyNGKEc8n5cdh9upWC9xEb9RphcfgnQ0IAyBAO7ocx69pMAG
XssXCW5PlrAzksTgFOA//Sil/yMTh4DMG/o0NT5XYRtnBJ6jaXAJgsQggmv+z1+c5DZq+7VqDAky
OjHvQ9oRsons+TWs51FG0Pynho7szs6PAKbNivaNSBP0DZEHnM9eXu6bijRx9LzwXZ4oRzyOVtNX
0w1MgGsbPzht6kFza9UxfYDhDev2AAy3xHsXojVPyZUq75w/BacUEQcswK9hLw+7pogGu/5do2aR
3SQAK+u4on/uai+LXMwNqCTRrZDEwAl60ZncP7Y5HmbJ+MDlkp0C2M/FTz53Hq0/z2rriOcHwAvB
SdCw8HsroCZsZJYC0me1QsEwJKtFfFsz5Q/1J9BdeX3GdvY7w/Ff8WbbnHq1h9foiw/ORx4iaBsE
n9u/stru6mjXOzdr6Nlx2RNLETm/XR6/sfxvVS/hmDp9YOg/o4zYZ30SoXlzOyfe2voC7Lq3s0yr
+Gqsw3Q/9e6OdFNkdV6WfEZf11Wy6RvmGmxVEXQw3vS1oK5H40mfuFTCRRbEfje1MJBNKh4Q54bT
pDRe1t6vqpTm8psKFLSbmlqrQSdDgaSIGtfO2XmpopsbwdcNUvfIs+1f9Qi2HFFjzM3wV/jDeS3s
2uhooCnfOuXZKN9R91G6FnwD6AnLIVyXtNN19KN4zXtSSUC9SfYLdVPmJ/afjBhXWkKZ3eIdVicp
otsS1TbW2G2H6tBiwdqRwl5nY99AWGGiaV70gBRlnQrHwUgujsTDLjnHAnynCOk0N8jXFXirZGsw
lOR8lD3nXxaLKcdKS4W/F/AAB3mzg/Zpuw1bWNbeip62B37Pp9oK0I3zA0FBwVQFQMRIZHEh1miV
uQthb/yxJ4TE7XA20mNy7XYelHosdyBvmRlWoqlqLrqEKHe08NOcqRz0NBx2cY0I9e5XXFSDXJXQ
/vV9QAv7zsTZAfYZJYNHWJSKFKBweD9pnftfgtlbb/ZQ7oKqEcjIXeXs7J0mZF5VrZjU0AYuNMRE
7JqC5y89M0Uu0EGCxr4epCRDOk5jC1YjNj/QSG5alArufnslufa7Jvfx8BtgRvWb23rKf1z2pqCn
1lbPJjqEoJVu+ivddS5uZuq9atGXrWmfKIgSjqMxcU/TtCv4I1ULpfj02mNpyLpry2fpHArG3g8P
QggefTnliG1hx+lolY6ge6BnIil4PymiqB2wuPx10Ibcf09af//zsWZNdWDhQMYhsciWAgnpbecJ
8wlYwtWgdPz7jsOdKl9rwAGzGZIEP74i09AhUfRPLqAFV/wLlbrGcd5dy76stMISODuLyl7um+mz
Gz+r/p4nA9wLN6/NbVqM1iyyjrTf8MRLdHXafRhbnHn0KAdivw9iFpDy64p3csLXS/EW/V7SJ9IR
1sIuXm0uEjl4NNpqLqctIFE1HN0iJ1mATaZ8Gv4TOHM7uCxjQq6DMgRvNck5qcw9Oz6lzCbC5ISj
RYse/4y/YMWmJOBLtcsOXfj/fL58xFLwsqLzB/ji4G7KDe2XRsFlmYYnSUxCDXYhUsNZGrtBDsky
uRwGtOxcOEwiTOuB8+qIiT0os1YJqhIiNNAnkAty44OK6QUjWSzUQ180XAxPgYrhFOLgWzLrnAsO
uiZd+bgehTmyTQmS10S7jfUa8c5Ffhgy4fzANZPccpqp3plWXW5gJ5KfoNyW7K90ee6GuNZtlXe7
hGaSSTTbojBEWMdtuE+C8i1IyhTpYQTb+ZI/vww34hgfDKpuJ3NwyD60UAKIumAogRtChNxeoup3
Fb8HdyrIoGNHFzU2vPekHSD5qj9NxrKUfkNErSbRWJD3a370DNz4UAFZFYhmizHdmAxZJc0iAm6a
QNJtMu2jNHgYQmUtfdUFJvR2lVhKywE/44mgMGHXYAvUbrvnPlkIGzSf7rqGsvY3UTB4nrKBVm3k
AFD9jo19e/2Z13kiC16oktbSo/Ks7Ck13fAaILmosbiyq8/j9fIsQpahJUcVMVKb2ZSRkusvlpMe
TN5mV+tgDCBQ35uknzaG/Qahhs8hX/M74T5NJAH3kryQVxr76hI+CMH7CImRT7xGtM97BxJ/Stkf
OLOetZ1Z5wnTQhqSv74Suw+YBhoy4n0c/Yo6aeScII1yBxePVktidq4ZBTpayKvcYtSl3DzXQOHi
KG2JYQYDrpqp4H0Pwb4UWwgKED6QqJ4D+BoU/3kykGRVYmb3i7OkyvVp0KvYTMtVE19s2hW08hgc
4cdPN8G7Dkquv0Qng2Thf5M8aO0xsAqMCXW1f1LRT7X357UcPeCvM0KLMzHYFm4rLjYsSCG66qjo
iw+xEFiirM82dFY/UBQZIgiAHIejtP6QBjiXccFCpSGigdfge3Iy0oi/q4tHekEffCdT/qT7OGoS
Iio17F1uTn6Le8VlVVsx4GruvzxqkU1dWptUUWVcuaQaAsfXjY/gMW2PFXswVXssON15NHEpEBJU
wcW1ZYjVY6sKd4RcwitiJ3RJRSbgHqtLRANDfjQibAZwT2kNkjg2FJF3yxPKP8Bldr3fXs6EMW1e
zAHhOQFH2SgHm7RiCXzmMKt5yF5eQI8pfcnddrtfPRDjAApQrY7CsXCQ3dyuUmOhZj+k5mjWOKEP
8UmX6322aJ+wDedM3MxdiQj8JhZrwclmL97SgVxDXWVe8L/HNieJoaKSkk1mrKQW6yMdYNGSOnLR
R9VlMloFkymRsj8CR7Siv1I5f2P3MTg/XNJ0PRNVowDkdUkgvYTfFe70OZ05fP6A6I84gRAjA7R6
cOxl21UHyRfw6rXn33KNAKlwLBf7k4IYQ52BI5F9W6AN7ZWQG42opOcZHK+a07T1OcriwDRiLpKt
7RQ5hL+Y7yjJCqbLnVCwNg4M1CMQP/YEVeSHjMJypmDZpi69YTNzXXDXxKezNyTZydbkytgBlvFI
uMuJAYNvDgbQlLLceRGYYI0SbVtp38Wgsg1Tu+MXOfDfLXgSi53ES8gVJGUIlmocStfUxmqwp4np
+znFCf6RmpwPRa9XtHNnUzxfBoId00W17pK7CsgzaHVFXymv/VKEVDFEvBGnJnY5O1obJvjC4/rv
JKCqS3bpXEUD6udtEEGTSIxWo/GNzrCAoyu3rVnqcFyem7o52PPv0Lh1A99BljgDe76f+alFX1nv
yPusBi4aC6F+O/BZVccsAf/s0ISwAjJeY63r98MQUluk84YkGKfZYawnZcKOJokuLVUFJfDdwUz6
+GMejloTmX24EGs133FbTbUwfcFkinp4zxbbmTaqoBgs0nTVzQtRMA2Dw9VcEzxFeqokgNJv7Sar
mAMeiINl+5VgJ8KbMkGQwofO3WZLfCjoC0aqZ7YgkLE02Fp8E84OyilT1+gSXWKxFn44qfo58yLp
XR8Eirgl0+7jnMagrGzw95wpuisnDkhF5oph9l6fq8QadvNVgEgJA3qILwhBuhcf6/yr4EDqfU1d
Qgx84adJ25fpYhOKmVFw3EGn/1mg8EVSImy1jteWiRZG4MPzfU+kZRy5gjCYCieVtTgxvPlCHi1h
7R1egonTlhZIZ441bypqbGqEz+Vjy8Ehd2tbkA/ok4C0Ev2ox+lG2N47Ohw/4gaEpPyiuYT3+6zf
2HsiJXViri7U6RuICDK/8nwi6e8Vl2RknH93CtAYmadLpd7T5lAvdyglHCPsVwDS1UwXU+moomZA
gexv8wo13QgGJOm1iY27bY2SQe2T7yEtBrsQRfDBXEu53v6AJWXKltQ59klOmxYJjfKKcPY4GGFM
0dfQJhe468coq6JV2LSBbs7X3NCA/mawZz5hp22ZxBEjsjZerHB12NlhvifVL6rm+DQGXK2OUJJj
Y8c4CussDzoj7T/1KnwWmcrRfQ+q7M2jzhCOPy6/K4SuJgoMQWClGRnStTxJnFuxhY5Ho7leycOT
UF0wX2LdOY2v5YN+eWB25Ez6tJktIY0IrCxnzCFU62cBjzWhGMPd3Ss70LOMcyIlwmFryM46Om2A
tYnWzmPEAazrdYcO5ns3pXmZyf+3F56XLrwxinTbKbmbnq3fjXVGNWmpZzJl0lqHCN8y8hoSpWBk
qsG0LVHqYDCZz30jauC1ZgaN6W7h5nJ0qxLR4O3M5056TCakmszFIa4KE38ZNV4XxoONc+6pSzGC
nOcx2U3ak10UG2UcSDCfNEqySqDvjvQsawKMqPcJ3xugCk+7KRpHLO2faitl5SffAwcOP8gdjJz0
XfCv/+qiv1ya3Y7Rv6r6t3ONpFt4/lZdCyONdrO+yit2nS8J+5KknvbwbLhZskWIB/6QLaDjEDlA
VxkPwH57bY+LEUToOwu8xliIQPP1bkhzli/ifjW2yPWu0nfRnrUerwtaD53hMfBHsoaEzeIS+yeA
B6Q0Il2+QBv5iG/sEOXpMvvGBkwnANVxxokloV1yIpSPDVQxuO3sZdL6tY4Dp/9ng7bUYAUqiVii
ul2WWPUhQO36dVkyV8vg6V2Eyv7pwQDq1EuvFvVfjerudFhfK6I4Tr6qK7zRnnEywD8M3ziMoMfU
DZLS+OJnQZUKtjcuv+RJip+pswSGnKXWEpIEppvM8/7gKndoG8vylglFlVd7+yq7hnI42nqI7CHb
nL6P5GeleOhHWgB9vhAOB0vo79szzX05ixzFlix4KMa8GC/S9hqD6dySEJNrvFjw2sUNd57T/Yd3
H/TjmvQUuUyrA0Smv+o9quFmtXrB1ObN/fz/9D25rMhQomNb0VKheCDcOP/LOHSSwPLHvfVRj747
zL522Tn1rky2oJjnKF/zf8yNkIOvlHVWSwLC9lnGEOYyMJA6siu8HX7kPxHX9zLbtq+Fagg5l4bn
t59/Waf3BohxFVpAHgxwftuUJ9NdPrk21AAS8C3vmgG08ngryeuht02yEtxy1Z1fth5IfUHK4DDt
wybnXY/iGUnZXj8vtygEbbnCcQwlb3ieBtQ4drPKGZQ1uWV2R2DwTMJ/dwItPb/HY+074cTDX84P
k2z2Sb1J7Nenu8kLX4K5vXpuXVJ5lm6u5ppxd0SK/WE4acRXfaGuYmrE1XBq2cUZvkEiz1Be2Dc9
1mjw5XBDlG2xfwDHyOx/Uzw2ggSglEp+p5TN6sYd0Hp9sK18BU27FTkr+JYa6r9io/EufmZNqNjK
NkaB5BswdBKMKEtbiDXFIZ+GtwZ5CLz5dflCtYwYa3qJoPEkzmZGUE9fi/9kF0REbpLVFSdhNIlT
Z/t3T9AJR98Oycqiwg745f3P5b+gFW6jnDF+3+/3+jH4v5keEZneocNZKTVgirb68muARiezYXdc
jVk8cMbHiN4BL736lzE+Vm6ivxxVcrX2D0AnsZRPvZUpMzEDc5rCQFaBnJYOwof/v9IZPRhF5MVe
stRr8vJSKg4mM+WmXKpocCWfHLfstE4U1dEb6jS7y48TE1XrRRbuXP3+g6wzARYc7rbHR9yd1wdE
vwgHOcOdLmBU4aUJK4I2Nvr6KBNyaPUOrW2hrjGmFWoUnvLXNSE6hPTNvgqtPG/mv0zThXEQpJLL
Y92SUb/xGHDw2p37AQ3CSMJWkADRVTNdWeF2TqrUah0+BlnbUAK3Xbn9JlF3HItfdSq2ZCzibFqw
hbTR6A5ti6KapzhKyITIPOpxcFt+hrzS/ItHv5kAMa6QbAEjg13i0TerCv+Sm6yVT4VaDB6oqDBf
jzpgz83dTjYG4Mpr9HHb8mEOfkcRhFzfUpo5MYpChk2WkjmT8yuDuSXSRravPMaBCE4ZWM0DAPNt
NnAZXlBZgzBZodob2AWXag7W/ipbvvsvZ48PhJaOxdR18Zo/VgaN1Zg8yzhomM7Y5dy3QFwpbrln
Qw/rB8DwK36GKt5LkqXW+pFzU6l518YkXmxoVD4ntb5RRaRgOIWtNL9q7u+YCuSl8wlE4uDnw6TZ
A0eMGgaPfaWjxqecT7uoYN7JbBx4kJVLaovBt8jKeE7fGFdVYtukVUtu0+1QoqzRSFwKcEBzySde
ytULvEgvW858BxjjwF/OByaSjXayESUfLP0mqdhyC644B+ZT6wmjfKeJQTK3MjNjxdyzvXw5vbsS
4BiLH/3P3qf93Y8l4ZepVF7sgWgc8DcQ0+XRxs7g8zEIjNRQtGDne/2ctA93AC9YJrKXc5tyU7XL
LBMB2Tq4pvR30nv6sU62sd2WHq3rhuZASB7A7Dj9xgnWKDrnoAt95md+f68t8eyyZS+6WDA+t3PE
8L4/ywhteCFiT3lR0qklA7OodtiTPNHVRklmaXR1/LUtMjK0kuVa8KFkORJh3JClmCwp0vb/mTgl
LqstD5+Yn0CG9DiAHy70Qzd905otFUFWVRaFxZ1gE2rCW1Go74NhjoKAR+UFr8aoA6tWk2KbO4E1
Nv6PGz6R4YjR3eZ8pT2PjzeaoPpBchiU3YSx9n+P81RyfKmG46N8tuaqARFKGrnuHVOpe1+ltYQC
Y+lmNy/de1DjlFAwG8r5gA+D6luMAXw3zvu8T37AkCisVx6kzM3XcksceFM03rRzE+CVAnlv57LP
ZqhZj3ZOgUAqfAjIZrT0oXuc99ZbdjoDOS22kq++lYC1n0O/waDSdaRmuLA8CCaZZbJxUQuVGpn6
ngkeX9rSoGvL6CLLDT+bPJ9NjNbKZRDvpXcUhNDPZ89sfYzGNKYTssXI8vyuSb8I1j83rBQsqIW2
lqrDb9O3Tmtp+8DQuuQ4nqpmsSUowZf2zXpXmOwDTBuQq4qXtup6uKw4RHe5kBGBYO8DZPKv3Dxe
iyiq7zldO0ipy5nteVy0F/WHm/tI4bmxM6lzJqgnaZRYV77mkX0sRDkl1ms/B4g/CO1QgVX99VCF
Z7qMwXb0LY0LfMV1M48lu5USvb5zjkQZuJhJUQwT29v5+c2GaBP5e3usRDtoDM6UvOVLYhqp2d8V
NVs9vqd3WvdvL2AeEWB/Wiybl+UHvEvAcYI+WNYh+oWxrCBpokSIsvv0JMfBbx+Mvsl0sxvFw5lu
bzWKaw2i4/Yfb0s91izMpdXJpmVdvcdXCkq9fBcHqZM0tvTnkr+aXe85NiCAA7Xvgxl39z3FV30w
wVPb9BETASmU1EmEgkfpEIujSeo6sG4NmviUTv8xYpDy0FmpnG/7FpzT4PDFWB7J194GyBDC4YhQ
SsWXxZiFYQvWPfVdn5Y0D9Ij3Hdg4g+5P56lAbY8i1r+5bI/Nw03oFnCcZL2K6rDNb69Txcn6PM4
TjHDbCeCMie48fpL//2oe4SwZh3kcbx6n9IoDS+K4yEVrfP+ZwkU5BjXHnNQeiGfyg9ict+FvDq7
RRiEQYfRIRiPTo0EQBCVfYA7CkItD8QrG86/hUWk5rqFoY+uuzrGbApR0fcbQHmutKyA6K1pNWrr
/qG27WbfeCeUOadIyUjC0fVvJidPYmXaAZ4EgpWndZwSPFSF4nseAc15uUCxv8RWr7laiylirJwi
3YbRDnkac7jvHRGm8qVImQH2cpKyhq7xv9A/g9JNfemersWMFMPUY28NpELEWHnK6y1EV6VLEHiq
MPrboG0Zufgok4oTf4G550jqqWncKDBnZ7kAESWvsiaUzbdKiuGkVpgR1CqRoQSau8D2bxibNU/J
FJicQDHub7Z14iMLnqOaHrl4dwndPj0QjcWGP47uJtafbaJS1lJKdd+dNWZ2zc674zmYl/qtJ6H5
MWG7Olq3kcUx8jOsUPE+SBqg74EsnnmcSlEuc2AfiidEGmsIrOsV2j5GJRZ4/82wzhEz+ki9XEGp
/usO7U7ZBVI3AlgsXH2NKf5vz9Q+cQXysLYOiT3wWgJrMzsjEKyEB8izSOAiQoCy185JbfjxHCRX
W0CBAfG67Y8KHKU+jkaNs/UF0EYQBDgI2N9yibsKrU9scTss24/hdH2FYvVwto5gA3jqfmr//+Wd
huqYLH0oS/7JbiacuhZekYcbhoKc9oOef7xgjd1KNA8yOVITdCNYcJz8iS7dNt93MgIqflfBv4Ba
y4BeWp3l08mBL5fzOnpwmWBNr+/5GHejOLxW0HFRTAdlPaRHkPI92ntD2TVeiHMS8f7FabiaImzX
YdO7aZGfxPuzJiPoLzjNRY0wE/YmmcdY7ru3FqkiZ1TlVcf/tNbBcaspF9kncUilnXxqe1v/sWmS
LhwYuA309uyNQEYyQ64QAkWRswv3UinssMdAwRu0770qiZg5NGTcnUVF4SRcAecxZdwpuht9yUC3
UG7CeDhjbaVyTsDQ1nBjL8IyY9zVpaiggnX/etl81JDsHV9+QnHQDRUsqVTL+ajmYlFpqP9EtdYb
Y5nstVIutZBeJKNPGnDM15hJq+3TsU8uO4DfWE6wseA1v5ICJZbtIUo7nRbw/xDSdxOi2C6MGWYW
SMa6rqs8StnY6uA2sOqYWuN8oy4e+Y+COSKBx7+dkrHPRteq3bl3yoxV7+8Z3YrLcWd7xjeNnYZW
ULWFcboUHS6CuY6G169y38r6eLNBJIHIhfyLHpXhWkBUQW/6SQLS4OdZo8Q8sgpYspuJ0MSmUabG
UdW2DmBvzo6oT/yqEMQGr0VvCa8TXbtNySEiN3A96YUj3UEITT0cyqlWrWWMEwSl2RKjeT2UsQnY
wmnEKeTEGw0oXc7qrQdffh7v7HenOwKYUfSJm6LdzX1ZJRmwezwYyOZetFKkrk203hE4u9xlEc48
unkFG5ZFwqHWgW6N/G2Eofu+UYtgFvT8MNQ1AYF7ike+k5Dkz25CpjLCsu15f+fCY2G0Q/DHGnHk
Wm2ET3RheWvAZGL3428sctns0GGvvKjDr5WLo1x7lkH4792Dc6PEgGFStH+iLXK3W0vKMMI1bbTH
IjSIfh0GweuUk61iJvvB01pxFMzDd057WtnsQ0tRKMfBkM/BKqrZXre4Ailh+/pefPQIgCcpPsjk
6+Llmh4hv6IZFdsSgTiz4iaDTHolba1SG+cuJNDNOX2RSd9TPLMdRWDZPqoUwmnnE2pmg3iyoak9
M4DG8jwch+sGyXa7DGqKoeXcIO4sJpQKWEeIsaZhGbYCMD1GHV1UpFFL/85OjD7F6gg6AlcknjVQ
WLT66aelfeL7KY4IiEw3+dNzHhdhXDayw7DBdFnr+OqEGmSDFI5pOdUFJtkB9eXUTX+hXdTVjV8L
+ht5dQFLyZ3R5fcVH7Lc0Zb4K5MWjH5DBKe4Z98gREFoG4bnhuJBncHU0x6hkN9fdCMUTc5/iyD9
ukiZmGVKU6y0DJx5l2u/IyhgjrMP7CxFLs4fQPfzTVn5lLjp82bX5BPrvEyKBFAUVVWs3ABbfMo+
g5QAmY8uuYuYAtCjFNLSXvAXenwqMq8d8HasMPLUyhscQyC3+RpZWMXGOw7Q/VXWsjqH7gQ8/Jej
+gUeJhjDy47oFIROtIZfJdCTaQ5bm4RTNYhGFEtFhd9sFqP3pQieAujsEah67j0+60BOD6ey4Hwo
J6a+OqqL+p9uBGRBd363A7y5n50AZvACTZ3wfweZtp0dSpGqvP7aAHhOrszSfQJWzzHt/yH7XKcX
0GNuBsFPqxPCQY1GGG9ahmnljlWCcf6fPDbuZ7045GhXcV4C8UTMOPhy41aJEvb3epwb04ee5Ubr
sPFYJJHw6f8B6zHnfgJpCfj6O9+EmOaeAgdtzq+439AiYVqVXMB/dqYTBgsCyrnTtUR3SoFgqObI
Rage0hYsJfcftYUGtpLBBkZI2yrKKEUk1f/uBn4XoW7YJQVIXjtKWWhT6D0GOOfFSn9P2UioiU4A
kM2Ub/2omOX3mNWJAQWN7ribKhWZfdhPpFIbFzHYDWWarCD2SNz+JT/8/LOi5+zj3Kv5q+BKcTus
GTn4pdGPlXhkL6IU2dK5DQBFeUFe3L64M1UUv+w1ZxDraDqf9b9u3IVWgQI4+cAD1IssGaJ+gAbl
uszfsdJqZNv9TvqlREWD3wBtl2lirxxmii758RTypsj1OASQlGKMpPaT2d9mPpLC/0j6DGsNlelT
KDRRo6UDIj0wEsSPjZMu2CDDAQJI6MlVo4OAJKIg6/0UaEwc84rIwVB5thH29AiljCqt05MCV8ql
2ExDdWMntsfPLfiGALHu+ypuyQmK/6m19FToE0cK/4sOv/zoYaNMbw6t2PQqby9zO8rHLXy73PQ3
G8ScUvQFU0Qx8nnhGMzTlT/MhthfvT03eK/+nwWdrOW0zYiJQEwFj/lPCjrARo4eETz0IN2ObETw
J8xNSRE2wXhJgPmpqDeVQ9ik7cR/efrgWhRIW19+uqX9UDb2LS82XBXbQD769wdXufJVAlPu1Jx3
4jYzFknw6pf+YSh/K1+zuVIxhIzRNxZa1Uqgwfi1yGnrocIfJH+YQWriewqytAcngk4cplQUP54K
2L4WYWmkd7Vocc5HPODloY3CKP25gOX6keBfCj4NGH0o2LWHV/UE8DJhLUVMW1Pde93b+8R8ct24
RHiSt+4Tk2yMRfQ+iuksQwunwkBsHGUCF2tqb6UG/4gS6M14t7aRaFqBkEDmhEGakS1u6hBUS8wB
toAufIBP2AfWykiCdR0q5L00VYrdK5eKhFDcQzVzC5gdrne1KvlX+FMD0YEc3ihBbeATgq9enC8N
quhCczUlRBwTfLfXpWxUL4E2uHs51rxELw2uKtyZvx57IatelHpiKcsXhLO7dIg32pAPQUFGtSlF
qTjcbvL8zANoYzmJBsyEliW/3otGRr1T9sbhHxXXHs0qeH7WQiARG63jBqcf+/YQ4ZEQynbTUvSI
nwf7I/LN5jgmND+3nEqjbZBFbqnGhOcqd3ZpK99pQ8UXJLnYwJWf6RSYOaodiSpnmE4qWU+lY5sC
h10Z4O+wtX3uctWFHlXIBJS2m52M8Zm6SMm/jzU1BAjgFruPO8ACUIhk6rRSYa8iYjsNIqbUCTGu
8uoTGm2E4SYYhKT15YECme/+IlP/bx4DKAVL9wUqI7yjr+/qIZHeiS4WHEMV0Eu7uFvlfKJgRWFt
hNXSS1UeRcZVLVh0v+BUaigVg35zRPnUHwjU+WhFX8/vnptGmw0gQi8cipypJcrGZVlYaRNW/7uK
eDp4ZhtkPx1Rzz2u3pxfKrShq3sNYbCGY9lKjKJRc9sldUj7YC715PCiUOWytE11ELtmSlu30wvW
fwMM4wAEHoHXpsasLpXjlJy1AGGV2HTiD0VrQatshKFB+MmQrkR0c8hEYv6FsKDHtpYDQJXdEzJF
MrtZ3Q/PutvQDFfjDqeA7tbq2FTR5eNw2cJ8n8gINx6tdrW7ewXZ1AaV+w6GHjq12aS97MrV5ScO
MAN1JRIgkSd3Z6c1dYdk0/ndQyjrzlQQIPTGn5+Ae86ucMvZ4TNQMKHN3PWlG4FxAKPVicx9SgJW
ODtGW4ItBz5ZUMofVDGsuZUQIh2SiS6by5J7WIlU2yfyzIYuOltlrnXx3R3Jc34elVbtJ9DV9SWO
pn7IVBaW6JBw0oHLFtAXDiX+HKoQE8tUEfpqciPqB12fTof8Z/vqAx75628r1B0y5b5jhOcHeqBt
IYxiocOEYkXkOCCEu57IwYM6jgLdmG72B4bFkAJBhFD/A3uJmOw0J7k/c9n7yBFlrwen2QC9l+iB
d2rngfqEc6E8tkyAWjYonQyVQNS0Jt0OVFuAounF6dn1PKYqJ3ZiEjgrAmf5vRoD+foan4Ww4Uts
GmyFhov4u2iLBt/ztTtwmmfng7WgwklFiSbzMGCivh4KgdU9gEpyh6UsHWRy5nCZt7SHQGLzpaIb
beY3j4hwEUIrGKJdUs3JaaaKFf4H2sTxUt2EUN7kbZYtgMMncm7IZ9s2cFC5jKv8KD1xAyXztGA2
TWd8RP/jkxZ/vYRd3kVVTeYOtfT24gjrMdvQvwiFyo41BtTf0vmdPdcF/xbs3nPh4utxwWlAKwOm
J/dMKAFYba30XwInvfgvAbXqu+WzYh1fSTMtBUUH/zdSRr+k5c6/EJNGcV1KPtkqyu0c5YbV3CM0
b1yYw4e1bsOyapb7vNUHhb6dApP0M6Y2Ff7kTO7kq5i6YMdlhgATdQuB4wvFJiWN/EK9FJu+hK0K
tBtVU+1PlF0lK0NEtxFyv+wTNvwUW7Wmjaz8yMTpOldqkRSy1ivVqJw0L1O4mm4j0Et3Zf1UP9lx
tCPEB8SJdnvvnY4U1F2FLc9SqfUyAGhpAdsgdtQIGkBr8T+0gVfZ3iKc2XpqRqGWV9yX1hEclFT8
Wyj5p6vW+NPlhx4pcOL8GOwyk7V8NvJxmqAxeneWg9/7lI5oWAY1GMa5VewSwc1RclrwaCY35Ri5
/eClvju3gHPJC2yBz8RJnN1EumFVOdkuX4lybVYJSL2ZFgCKb8sqnixzdMOrPpjq3VSChxPlWNBz
NFXFV7VmJNCoK76Vt3gY1w5Za+1cp60MX1Du0f62qal8FeAEJnJuJKhPGkWZpZ5XUoxyWKdwgR5Q
iN2FA3tcuFXeG52Q8/GCIP75ejiG211xrQeYMZMCq9s6MyQXRtAOqyk9e4gZO+Oq/uC7eMwjjN+8
F/QDsOE3BYPjaGWQ4snf61H2X4I9NimVt2IIvM3YsQa704IWooPv2kgcF57OskPxAZH+JgE9lXyR
RAy/ssgNAVN9fz3YzNSvQuSLx+RWQZsQcxhxDehuKcIH6SYw6vrh+BuJKH49e53PpY/2SD5XGt1U
iDd/zuaoatCbKe3jvRBlXy9XVkCtxP/xuCLrnFgQBtg6LxfrNXtkwpUERLoV6tUsmxbyA4ShXCsC
jw65udbKDp+C8o2XfCeruXaQAFOUYlxirmCSQUWFIaJJTV7Kh44uNN7d28vILBEuai1zUEUNUx7F
kNOxJf06Y1w5SR8goJD5xtP7q4K5NNZfkq7OaPpo4uysY/oUNv9veGkfJI5buBGY2KXX6QCd9p2+
1h3lJ4ZU8OU9ggFmlqxpm8hr0khD6uR+4ZSLVnSxzkE2sDOC5GDsNKNkCnNKUWylI3baDtWAMPJi
WF56uedHjCg7P0t30IeDYm+2sYzlD4Y11ymBaKGEcHOPmjTmnZwzfxQCqYSwyQzsQcNah60dEVcN
H5+FndbZUbQ/35DK8/2vLiaaz2YYpv+xzy4syMH435Euma6LKB2YlJAHi3JAToz4im1rPEqa4z9p
5CiJxA5xt4C6XXMCwBTdhpH507xAtC8mRRqEUADAMzyK8qQ++miFOzGSvnjL3zZRWm+yOGaeComV
9lmH0h407H79cMxijB7pW8FHh9RGrucpYFLm8v0sgcdp2Xx+1t4/GzYjsrfkeiroMDEnF/dryXdm
qLvtCf5+QOC7MeiC3fYHui2fWxoyDr4zj5lfhZMikEM+wzaF97JTyN1t9VxJcVXCM4oQ5iHKkN8h
080VjytBRqfAD5VkHL4qyBNsCb9O7VqKBXxoPqCoeSU6UJMeTus9pSSDp9nXMFgzg49GhXNThQBx
UowQTduxF/Cny85u7pMU984idTsmHa2fNMqBkhZItptsdKCVpC47FNPVWn48NqM0O4oSNVFZ/Mm6
6Oqop6TCEe7ad5ds0Iv3vzkzHm+bu7lUw5LG1BAIkRlnEmi2gpX7/XodZtQmaRFP8xLPxztAiagY
/hTTNCAvTpep6DbUpTdhb3PmU2Jv8bZAA98RFljg8oIYj6NNnOs4tsgcNGrjtQ4/1BEAU4sO2xzV
TZ6gVTqiP3hRhfFNaDPXaQc7kLFItiRf2rKqdj2rFIF2Nj7vJN9ZA2553h1iDKxISGyWqU30tUTq
Mx8/9MP/ZPBzBNw3SeuDVq4buQBtEidIXHWGqwfyV1Rb4lfu5O05l71Xw4PY1E0eLKcRfxh4WyAv
3CqvTg1WPDQ8cPomFl3daRbPVopVe9Z59ACXW4hwe5yZtxbeChsJenAXLdCMC4aknELfCXboUuls
LFdMQGPeqP4vzUhnfF8Y39B/Cfie/mlTsWKA0s9zMS7hkw/9DdlQ3EWtQYe+wdPHJ7b3I6G6+a+v
6OoD0eC6F7S1PdSgh1SZWmZdL2u+FxYNyYRiEJ3b/Yu7GySAMhW3WzfLbEbbOlLiozFOmV70T9PK
WPRsae2QXmg/M3+bBo/9lxyBVhG58Pk7r1Q4TNhwbqjImE2kE/JGiMCZB2gpY5nOiQA/FEUk5LAk
t52wMiGq2P6OoGSOCyS3PIxgWp3oI+Qj79LbauHmV2Bssno4FfIAPI8jIfM/UGnIs5p9PyUzsKJg
lIvdknAZtQm5Vmp+UgrfGA1HZ3YfoU/7hcgcKEUsXf/km/eklpf5Z1U3pGGmOvmtho0Vl6kUsXkq
+E+RhGE8Vgm4P6mV16SIAuqwZUWLQ5wMyW9ChvhRvUZda+WpL0cjENpfmxyE0Ix0DvL3IOUFATFj
ahrXODxktfowjjkXpt+3WyhqmoLiLZ/Kaz72Pv08eEBG0b0UYn38gleFtAVOJI+0GBOIRRoBJpn8
WEfcxqJ6u0U4n8/yXJ2Os/S9PfMaAvuXdPDfReD3gjsqDgRbX1pOrfouLBCJ9DgOA/DrUFb45TkP
HANY+LtkxWqiLwFq0lNOXLci/PvKzpFRqJJuAIW03Jb9i57QU+Y3l1YqgFLxJvzZy382yvW0DFJq
emg9y4SAm6M9eBo9p50MXgjnTiU3v526ZHPH053+U/xJRH7T711iLLfudJNSf2241DuOO7VdzxDt
kJl8rrhL0tkoxMuYyEnbhcHDeuZrDT5/BHT0KrxW7gPla5Mppdu94kEzhH4nZJjXGQ4X5nAV6eXh
DXyh5pP0IJZ+aikoSI769ytn3RmCgTpMKJqvK8n14ms/4ohTHI1bteK6MEM0YzCKWRFsA5BY+tHS
4QZXScBfX9ZYypMmCN6N9iTcaKIzdgkgIT8pfdBVr4WUP4rhNqXCHWfHrWNghMRHRIMPMrPCGEVn
lhyG8COlgce4mizWDmJVHIk84ldXciWhFWVMfZR13n3FW1EAEMl22dg2GxFqFr7+mOJ36Z26ji+t
qfpw3KXTjKhsdwK8T/reNphw5BbEfg+g2IL0bYaes2kpYb5Y3HB6EGy4u1dI8uPUtH6lplbZJRbZ
1l6xo94FRbxvD4RpGa/2QxV4CjAOkZ4vNd06UMB2f9PM6C/nG+oFlCxg0OYBn4+Jm38FHXIU9fY8
NkBY2kuZNm1fHbj0kMUYsjoko2SrTb5jnwXyTdQIAwn9T6lOnI9NjaLHF3xqJbiSaIUf35v7J4t5
P2Z8Plmu5BmRk3B7JCC/QWOO504/BjErRolK93XR/nzVV0XybQzwUPHYbqGqNjlSMEJ/n97/Qog3
Xv21EiyT/wmJj205s2FAob+GWoRrry4oPA+lmW/+fDl8YJPILv0owfN9WfWc/nKFMKy9kNRTGdGy
4FU/QKulfhA1fLL1aPmLwsmd6Ns9l0ToyBWh9cN1lIYbnAPfax7Pj1Xfy+Yx+NtZttVUG6uvAqgJ
q+9UH9KpmM07MjfWXkgKVQQ/S+WcPmMr6LFYPXecE+vHBe/40luvE/mxD9WW3b2f5tzC0gorQIZq
5r5TYsj7unLvD2V+WMLlui0+uozpmsZ54n5V2aOIlCtxlIU7cqUpAv1hZ7aGATddlPdJ7KPJwVcf
jZCVsRTyLGL5jMhBl0vxIG68oWU8IRvPFPr0OlJMkIbhsxLoiRs+PQf1SDz3NEfsWKTnOGbktDq9
2d0TSOO6xDcDUgm/l9N8p8pXJ3ymrn2maz+KqwWdDhcc9JZX8srSBny+KLWvO68zmcxyV6PWmIfX
LW5blrGp+w4axs07PzPgUQHqa6VAjMIZ4HvHkjpVt6E3ssouWrpIv/e6qhMp3N7RdxCPcu3I/7j6
9P/z4Skb7/8ycQOfJuUHlTDGcTLssNWqKJETWMSxixi+lEKqjdN321TyVI4hFQk5HJwPzpdj3YE2
fScjFmFy9G0K5mSo8ugGjOcMzZ2zMe8z9mn6m+R5N1uaqRnXtlOKMSf8FzX4YgdMPNipggnu6aES
dQveYYWHzkVKI3aUj1rhf50UuWZXgBt0vBocIEgF3DayN1q+lnW7VDt9irXcicq8cqRFDOgFTYUi
y2kw19Ns4NCRdvYxVh3nTJgMqMkkR4lrdmJYYCzIApUu7PlzihY/vzfW4R0LTHoI2y2ydCW8S6dm
TBm15DXZFz3lGXxMU82+T8zNCXI8OqRlGr9DsaeHQS4OCS+qRKuLbvQuoyJim9bXsZT2Vscpsj9P
HXiVh+fVBgl7SYVt27yFqm7cFKhDn3dMc4UCo2QWpGITFh/FUbU7/9n+nDCvyMko56AcsI7RPeNd
Dpce2tduB9cMfuYo6BnSDxxYZ+mlDpoCexQT/151Xu1wAQxMlk8dC7IdmYuctzdgDwPy/kz5LU+H
0WbrMefbDDnfC7N0Y1jn2r4cbBnAouF0qpFpiceQcAc5G1u/i5R57hn8yN5zejjL2jpEDrlH2nKa
wjyFDjA8dITdV5ANTTamG2PpmtA11A/xVCzgLmNMVEZSiijJf35ibllMpntwGl1JXd9Hj30QT1lc
Im0wJ5zqRJ4kz21XbzACKhFQCowLYkiI8UUzTWu9oE0CbetmdGrcE/N0FEfjgnQrSy2GwpG+RN4f
ndy26KmaR6Eu+TeUhiuYSN59aO5UAr8vlkPXynPIRDc6IbzJO8v6p3uVRVXKiLNl8tTBWf3UEPL0
nSxC0EZAw7LhHp7Ozxz76arV/kRlAyNCi56E1ioLt4QRwqHwo1lzZFw2JlBI8LZyOkHllBap1sFL
Rh4rSf6NPT2309hNHqr31EITAnSNvILJd+P3sOEcogGM40fVEcDOz+HdvOc117S5soracvI7hbe9
1PzFYS/mi6SKHBnMoq2qNWuhJFWJxoKDZKatZyn+tBZtpCKtdiWD9Wd/mHf373AsT+M5S2XTDx2m
omBc2FmEwJpl0AwxnkvXsSW6/+/ehAGkTw4HzHSSBH7/AeP52eFBsnxi1uugQ4A6XxlU+3nBB69g
qldSnTW84x9sRKefABVw53hcBcpwuhY9HJ0i1JhG6PeComDTZ4FZ/StPGt4ogAq8O1eaCcjY5oiy
cCDpc7XX39JCJnO5GCEOrmnYlsUkVktKhAFZu2t8ATnVDzXa2KkBDmhvVPPAEwRfTUke2qNHQYMF
WVt22i/oSvtuCTICVOdzd4aUDYKjolQtdWUN2oP9yMkdZ0PFDjai9eAOtAeHxJvmU2bM1K7LtGys
nJCKRrLfwdCRFxnd4QoTktxdtBZtyDMYlZrupsF6RoktZ5pGMibqmr1iowJJZ2hiJYtyIber+k0D
Hts7t/MYuKeh4TkmGXrnqcGMdkfvGfbJBZqAYKfO8AWweMqMh+t2nRroesUCAHJ1z5ycm3mmOMaS
yosoUC/uXoj812Zx2TpokbVI/mfwJKoHavfjVz5daQezXuqiwQQGpi2pDBKFswcUjf18bGjc9TIl
2GrvbMv1CONkXTm+RVzNQr7dC48rTe/vMZrvB+/o/5gVZ/9p6H+d6I3msnX8ZgEjnBaC53gHE/33
ltPHqZkULC+BTBwNTm/rTV+WcHqLlJIFwuI7flUCCy1xOwt06ANtyHnn3FYzaM4c4osgA/d6+iSq
5AfJW9FxtHirdTSOAe5EOachpChyROBL6VCGJeEe3ax+g2l3QTPEQHg8wZPEKAf8lcZnnkMOal9A
WiGzf0qqjXUC+eGzUbs5HeumuaY8CDqoYU6EY0c0KSE/vduxBpRbPznUM+Wj9VL2v1sVCAj8a0pg
y1Bm0Wpj6PT2J3y4hSVVWDoOsTD7xelDCb14B3xAIoPiSQYHGHbOs4COVghkNThPX6IQBSnGs+Eq
cI6nKpDAppUbgIFd8TylZa6A6HOpVRe396yE8T40wFgZp89jBXBh1QXZLFT2n5nNbfAexJI3pI4J
dp2BrRgxqeitp6M8lCc4RwrhyR9MkM+N33fv+mraZPlmxf/2B7J6GZV/lBsLPnlmPYCpJ9PJFgpk
AVczVdEoujsUjN0xg8YgOL3w86yLasK7urOhHncerVPIXxouwHmWWDq5lar4JSVzS11lqz+X/KZy
sAYwh7XhLjDRR1SGA0q1fiMm/a/CFV3/df1FJlZwThn8G90APvGKuc/z+5hL8YGm+1/ygVR9bzGA
ypvb0yMXr6oRkyfKI/5EMa1M3FUMjT6QScKMpYA3tgdodfsk3+e7hiuKyJf+UqxGNYLjV6LGlRM3
JSu2l6WHfNe1UhivlbN7mSOitKhBY8XiSLhw0mABKvnzjJ8TDnTxB4q3GQHUDANA8EVtOQsAiv4g
ACwt2UvJHxNawZmCeU/CLLf3L7hWHGewEb2XY7P65y3YlQ2K2W6j44PlqdpPkuZMgEfPol4O7iom
7eYI63SbTdfwc7/QnwHy+aViMnVva3KgaRFzfEkaG9XzCIi0VvpRJsdCbLpXt5AkLXzN1wrM6Xv/
Giup2lguSnQYiqOjx/wm5p2+yWNmX6dQfes6vXywsIgALPjJ74KubN67AQ2sTxMeb/dPPtvqXF42
oCR4HUeIxjCYxNVtvh5R+fjV5LFCeQXnS/VJXTrdZUddYp7L7JzQWpU+c02zuEsuQQ5w46b4UNEi
l1j2NglCmvYKBxdMEX3S6pqf+HqunkbejY03wnSQ5gFCy8de1tPVWYVFI8zV/S6yJ/VqLiPVqsso
F7nPAC9UNl9TPnvqJt30jbDX2q+bkioXoxgwo4yIbryvhYKRdFpOH2MPKh6JrTGZRf1vymZGBJKc
VSu5Q7ji/ftqjKHX8sNHwtPWkImdR+8CVvFkSJGaqxIjSUXOU6Fj0DKe3Z/qIItvlMVBU6lA1Ef0
/FtJxUInZwawfubfMP1TvCAkrfQpd5fb2lSZ94DIx0EkfJjzIKGfnSOdsegsIuQci1h6c6sgFHev
cqPqOBM+bmLbJupNdrHSMzBK7xvllz0pMhGjKe4GdXJAsy2Ml0icNORvBVigkOo0DIrGaaDZ/j8K
nRI5v00Y0D47PmlwWa8Pw+IX2H5XCElt2cMQ6ea4z7/QK/aeYGh5Lio603wQe3K80b/Pjnowa7un
BnLBt4XWKDixzmkHDY3yg1WZ+dqLi6xFvHddDSktnBNvJT5JdqNnu5byP8/sHkHgJMuQuSnvkF6Z
drGyCVoF5MVllJqCpY7zS0u128KcynwjmOa1vja+lP6396ML45RK0TXuaBDIgFNaDTfaOdVZ23n1
biNQUncVbmRW1QZtPfk/4LrHF3cy8S1ZjeaojOt/GB/RaHTYJr24TH8QNqbGeDflEYP7XsB0tHfC
xBng/wXd0K4JeTwTJGHMZPm4wYGgNLMkEe9U0MbZV69JsHj4hP4LqqZT6SlPa9KmLW3vbBK2bI62
2oj2uONOyI3Wkv9GjNTLg7LYugbqW8s1esK0s4iaVAzdaBSfIOKBSeR/ni4Cx9cNTxrrAe907we1
18eESS46h6BUHgt1GXu6oyyGr6KSjPTwLtsI0jRvsaVXENwmcYX2lPS2RhvlSl5A6TcemA1yrock
vFYLqeEB5UBRfQY9KVSyLKV8AYMcl2yxLFSG+Y7pV8k7veVqa05PRO1qVlpJp1UlPm+emOtQK/el
O5cbv/udrCenAPHpkWmXyyDEayMcIjGj6I7JZThwutuqLMVHsfekEP67xU4T29i3br2+wc14sLiz
BYcrU95rGGPziEmc9dv2INcGydjPh7wxtNhJQxnFedewp40efl6jJu4WfdZUi66EVoi0EKgcF/uk
G+jycESkJIztpPOlOf+l3EUn2pvwfDIbRCtTI5jOBDW4NLPxZQN0HYwtsDHLc7Xj6Ph6zVVNC7Uk
KJPwT/VU14hul8udAvZeyzRgskfvuQ1GvQk82zV/JOztLqFSEw9vyWsxPoChTyAfX9w5tw58DzKk
hJ0WpPTlvmE+gUJL8MfA8IR8Vozom3Sp+igt2Pt6pa5ZeyZl9A0xYb4aRKWBFP0J5+eDMLpVVkIY
I+8TAN8g6+sbtQPgABHZ0CNiJkJUWY6afqCHypoUC68UiqFZDtwd9BB7h7ScqzZIAEVVJb19T01X
soqwHgFoEi1jFq5upuT1uBfxv0jJpjzFBs34kYdNAzIpEAcaiTJgut1Iptm6hUW8u0aUz/pN0un7
2rG9OgqFpswZCTIwDGN/zc7E2fWHGjeLNyLuqzApoKkE1rTbQjv1YVml9rEcIAc9Ja/KW/re8pGb
ULgQJQAyu6soZaMkiXXr1JUb7Nhw0hUT1VJiJADSKFaskjV9jEO1BDaBkBj/1qt2C+f93LpKgMet
aYZgZxdt4292JoM35FGXQGl8rycP81mQIXQ8P60sfQBfnmKwYBWkNhvqFgwi6IAriEBSEL0FaQUq
vVcJnVPkLAIZKW/UyXPp1wy39hi/lXSWdbbOuZ2Q0Ry4RdmacvMo6XyqMiBxa1vSGVss7b/XiQaL
vzI6XudImN7TYRwe/JaxHDV8WIHFeu7GS9UUJUPGzKex+WZN/40a6t2HrqRLU5WJ/o7ezhCdCU+0
Bq8BsMUGn+I+GyBKJjP95pkVeUxwzzuXvJibZJS+Pcr+VJJ07EsPb/0v2GtT//ZJ7ydHxM+OxVZF
muJCT+yMKtG9H4AWS+rRaoO4xLrYEP64Nvfy/mGMFXbjaoIZFlM/oe4HsPkmANTzFcBQNrQ2P6Rz
n9wX+fhxP499E57m4uTbkvafbZI9sxuvHsGkW2bAu/sXi4ualrIi6l0FXw0xbcSguARLai9sEYYn
Fq0j3zhfY2nCIU9tvrbeQFmO/M5vqdvKf7sjfgr0+/6SncBQC5PDAtfw65+OUFmiWUliVc2ydOYi
nJSeOH5dQjoDko7Y5quzEbLJvNpg7jW+bvtCdRfLTZIuklKXfxqAmqXu0fcnS1ft/CB3ydBKqEHU
Uc7PwzMM/rEz/5k5BGLOTQsUtxd1kpfqdJWEXPQ4yp1LtclfNYts3bDxWj/7sDji5r2l92McFBhG
wL8SAtUTWOzlAJXYeuLdYNd+diDMaKxYEK5ZU7jvUd703BKYc9sudP9MkBjJni33x6Qyz4+L9hic
aTItLZRmz+FKuW5Jp8vFWOszUoi2DL1ufw8SbFJosGnWiK/RVmtX7u74X0ir38V0hxwFlIN3P7PN
uA1DBgENXlAWMbeIz1+UnZHFuHj3p7ZeQOEPUOsEu90UxQwXKYPFAr6PGXbWQnzmsM5UR4XkucWv
tAzQxIIynGgyQJTTnAJm7KWmaleI6t9kbAth5lQ0Q4zmJ9GwZIWUqGb+Iu61Q0IYPanTWx9owrgi
gL5nPu9si0Br0h/GewPM/JSUwRDCi4KyAGXP0iDxVdBHTsl0oh/uaTLuIoWisrIpUxgrEPH1Q0A5
d2xgmvnovw24+dUDA+XljnfZ3ttoCLpIlV0KGftasatv9WsMXwQhgfgIokpZ6zI4UNhZ17AR9hkp
Hg5n0pNkdBctUaV0pb19cmwU2HbCrZHGEWlD1pnMzaja7BW2bHkKWBeYUzGAGYnAKnCH4/nrEClR
roJgXvFi7+p+SW5JBCRvocbUjcu2ICBLpsWK/S4SImCKsoOQfOx+cTo3ldYuoFO9ar9U+TDIz2tk
K86ubsD0vSBsyiGgWu++NuoX1qd8DgdkzG5gGZkrr7UISbd6riMg7OiMlgG+SyZpkBSDmo4jdaF8
tDO5Ydw0QrPsXFpNFb2uEDKQAz8EesZuwGHZ0wTL55l3a9YJtwznwtN3Tl+x0QbHSTd/MqlSMA7e
fyr3XEWw8jl8k+ikUNr+t4Ey5IZ0oTkva4gLRMyCdR1aJ/5gnFQaOdtv2N/YbZF0dB2zmr9wEyfa
ZjJYbRfvpQh8Rxku0DP2iU5LzHrA0qsTOq78xf6/QIvtcHRBYrw0kj3Y2nJqXNcJ7iSb0LQba37c
FeDIvdS+Y7KqIFtIjOjvXDvZxCuZ9JL8pYlidBP0eXp7Qn09fmb5cKjrrukPcIVo/eqJBCedpTJo
xB+WoFLEtx+f9ImUioG7sUyWR0Mnev23HhLVj7+H1Rs957dOiAyzfEWOz8aJKkH4ccaNfq2mcYq4
GMeX+46K3JPz/Qw9mUMtq9Jby0BhGmBtGI9cZfT1EofFsQoGy5hDiydgmL3aPjXq5RRc19iYzhE0
BNd5dQvuwfL9bqtvFFkrPIFUyYxpWej9ixSbetOld50oiwV6Qf6ld8++t8U1pFBlcBCkAFnoBOuk
O+mHbybhVX/r7lgX07hUuTlpVHmti0u7oqKVW+vxz8TIoajVyPk/WOEEDueMWGmI5Oi5nMh0EvqD
3yLg8B2plJa5uMNjwfZ45gsAjsX2o5UveBaEzldmQe1z1C12pNZEnrCmcQCtDlrCnqHy1csoi8tw
h7MIp1MBNY5AmQ/nILQd1hqN++olI8vDEALZ79tOTeB5XqUFo+Bg3xWLbwOFZo0BGkqlG/fxJ7O9
K/f8/u784wcOJeydh4cA5QQMjnyWQI6ugiUu5NSYu+5SXHrUJxxzDtmq60QnT8WRQ4/4KqPmyrgM
86+8X+zcwBmUFsY68+uFcJiA8lNmuZdxnbKyTNnckK2c6fKPwaH40OemScQmg2mcI0n3ZSIYVyfJ
QTVeb0wZbiKeBDnqPjn+wPdItH+Y6F7gz2JG/tj20i1XW8XBKf3Xs23ammKxSeHJtctAOP8RtNf0
ft8wRHWVLF6X93UrN+3MoKSyKFhWGYThuvNNsD1gLGOyatJ+e8UvbP2/rlD8HeVKwKEraKf1M5Bj
rk3fPG761jcXUyKRGskc7AzR6o5Cuhl9xr4UC5264iQ7PzE31S5W8LZO8rJkl9R8xV9HaM2S49MP
cwloFm4OxowYtVkq9T1ROP53ow6eC5G5wYuFQ7UlR4n4K7z9vGQaZ+bUxI0mK7tO7+QtP8ztEAdu
0XtmucW2YmonmaSDvZaJQXKW+XrkpayAT073ud0ZV1l8qZoPmIw6SzPUaEWrlURZsfwa3h+qalLn
zM0vyOoSzOf+1u8VngcSaSmNZjmVrrlD/lPXKkvVDQUyyMkywkqMUG/AooyksqLb6hzih5bPUNYn
5M9PoG0lx8uZWeOlRokzQwjwMtacwBI3g5eITqcKD7oU3Y5BpqEbwJhlBjEPuNnthMzOZBwPwHQm
r8VHTAoOwXXYdXgTy4GezlDmLuQv3OOx7jBhTSGgfZ7C3qci1QOS8lJlOsFDilOwdLv1+TDC+6h9
nh9RqSjFwiKjIm1p9Ycx8glgMju64rTV1Yep6cAKxSpwf5HqSbhDRjx04Nde0543aXzqtoMVhosc
ZDVQD8aplJC2xGpNqJquF+7jC5owFmiTdUCTOCYLRhRUTICZVWvb8MKtFQFedSmEkd+V/QE86qt0
ViD1kGBL6/fST0heryJKoBFUqXlSZGlvabRk3+EmcZk0eti4jdAYuTC5BTWTZQMgPfaX+N7I8bjQ
lk6LSHZzGk5OKlWCtCZAapKxRXt8Z22YtECgj/x3Q+5dgBne1s/+giRsJ1nVsupYHnF574A7QHcn
v16weJPMy1rZFUtkhXDoG/IJ/OR25S9IPzWx8LoFXMg07gwBmoRXFol89+KTXiVNmnRHcgLFZlgv
7V4G4IyusP+WSM1my5+SGZJd2BqiMJQ1wL1LlW8t019ijKpKttaVo6Mf7kBPBF+DOPZaphrcydDz
vtXwYRFCpyX9+0Y+fIfCLKPIWRAkFm0jlJyyIIHGHyHBUTUJaHae78qza/GMAz23j1li7yyKnEh6
qwUt/Hge44QZ4YKKGWxmjloLq64Grumhi9W6xk8UOxa23FrkpFiKLOPRz+IFNhdIcxbBJQDrHA8V
BGoYlMq0vtdZCbOer63OV0vNiSNpI1QyWd5rQ3b7sfTq2lzGgwhuIjvZYe69EHsBpufSICoPbFk1
QTGXQAQX0ffYFRRzuOCtJBoSup2X9y4x3IBm9Eql9UbFVgjLBRQ+lI5tsgXDyM54xqSF6jccb8WR
lQYYBoohjBH3S5gCR0kzj2XYWqmu3NEUP2uPnpqVbRzaH2TnJgQA/bs6uW44l4bIAFZfTwPknUTh
W+zWySd0g32pHyie0IOUJweMH543367GLiCXU8dCFyVgbnRwUy+Rl1YclvbivCWAQit/dROehx2y
IABv2SDe2yvUs6liXrUrgDmMbaFGTWvcmREofb6mquD8E8ZLwS8fIEz/DRVqT+4Elvmlvsb+zrun
8uAuwuQH1kR1rGc1oMreuxr+fqX3j4WaNl59BdhorOtNdEslPFSziV8IVi0mKYetIefd1UmgTCI4
6lcFfOWhsygKIgtG8xpF/31ZsTvXWrieyHRphmLK0/n3H9v5UiNz4RashBTeLdvQCcn0JO8KD4RN
lO5FrbD93g5BZpyYq3q94HWxmLXXavbRVRyxx5p9rem+Wz+chbZl5+KSNWCZMsWWlBryrRlAKCPV
5vyXrA63POYurdKvgRkKndFUJmar00uDBAcG6VrzLjZobAGfTpSsu3Pyej2UsaMjv2qpzzveEGRo
JrQE29bbRvuDfpDg2uUUHrxJei56cCiEAvvLqIme0fmZQKxMUM6NlgGR12wobTFqfs36v+xmj2y9
CsUK83ae7EXMpSRkqtKEBCtphQlGFfpK2hb08gmD11YrdMwYO3nL3nWQ5A4mRB1DDZqluDf8oQ/l
4dW71j8hsNV0OMUBrIxtJuqFq6r5sK4pjOz2xOJoZt6HuhDJLZQ5o7T0StEWzAnEzXEjQxby4gtb
pVCILeg8ZIn6Uw6Nk6O8TzUgKCg0OrEVP+I/sceK0oW3vfl7ZX5VinuTc6hjuLIPzeeTx5HpwYWC
g8KFAcBc8xjOpMYmpD2hsK5Zw+jSB1PCARfSaPwhD5W2RSK/TpOXOrYRlFAaC6gfBFLD5TDjsHOu
bjb7ABnCr4O3vCRxch0KfRCD6M+0FM+sRfoMmysL7C8wjeHTt8loefHWPDqrCQwu+fOHJgCGjB66
zmNULggi3q+/TEOnKgImU1SUEppZ2Vh0KPY+wTwBNWDj838Sx8pbvmQDM29VvGNXvyF2aw7XLviN
vPvM6mv8s7+nkq0FjAlUDguGY1IgNUClWNfSM/+eiCstTWHDaHuFENeobd1ZS1um8K5R4hZm7Yh7
jZS0+YSUuDwsUzzXqiHxNOh9xqX4SCUzkUZlcgomot50m4QJc9H7AHhkcaLmuTSOFtOJLsJA7M8V
AoahogQUIpx7HkXY2j114olNsNrm0WjDOAlInr9ARY1zdXKarwsqcTndF/uGJtokPOFsoAGe6Qw7
xDajtwWvB3Mtogp/RTjYOrRIWpqKt+rFPvaogTfPyZWRxPITQWixeIVj4ZhGkSz1WHiVnTDj02C4
UWAhHiY08WRyTnneHM1iQRKuWxqd8NsssgutWb7KFAEnBYkuK3rajdehjyxVLkopIkEyCxKKRhd7
2Q3iVqwdW9tsZhAXo4A4nHAXaRjfIGM+J88jlIm1GzUdDjkZecS9HTHWlfZprsZ/XbPcaI2djspH
Af8mSI89UW+t70bf1TnD47VfE7CcYhSQGP22mI+dJt2LCm1YWbhirDlNUAxTvY34m3SOSBhZK5bJ
7/Tr+vd9jkTHQnfj/M0N1eJqfs657rb6kU5tuNF2O8XYgKJeEuWvGhH2boIpS0FKe6BB0uqZUPW9
nLEN5iRMnOGFVeoVuu3DrOizPAIvmVMvLxSc4x6oHD4g3vq6NEp71AUeA+85p0aKY0fX+ATsMcbI
bwoJMRwpwpofUP/1w4X09btpviWv8h7oeXaOWXcYnrXXmiK3dhuP8U20kwxdSFf9iq6gBtajtpKq
3vKmQb/Xw6639m8fphXu1x6F6LG1Oy9nyC9LWVUC4ewEZ/Wt/izfz/SjHSpfQm5X22tJnziZNeev
hkY114+9oFFZ70pi17zzjbk98LQiQnxnWc9YsLOAgzHRSJ3VDfWF9aOgbm1DQUCK5kkMDi4VztHa
MFT19SCKbq+ZTATjKLI/M8nfUdtNRAYF9WGtxkzQ1NMOpSlmebBrwQP9dYbaRJLfRhkbE87f+Jij
wiMHgvELU+LaXbmR/cd2ZDJI9B0kvIWQdbhYLNcVASmv/ey9cKsv02fn+B0GBsQYtMs88HWpikpt
5oaMO77CJEflaxdzjPI7enIBgxMx/mI4a97J/57doxnoufV1/+gi2S+TzM21vMvIYvMzTiah2BQ5
+q7jgsIw2fR040OCddkrlcM7JA2muaNv0aoN5kvf4a+aDSuk5eCQ3e4I5cg/70LgFFyB5oUDLVPU
rpXDKHnUyLhvFIUGn8jUsyWP/2e+7BvdCP9h0e17UK8ugbpBm3mG2GWf+B9XaWF2hsD0sk5LOQRa
FPKm99apaO0HL+uiTD2gOmZHdayqHtO/0nptfoI1JC8UyFVk1az8mAYJC1xCquns4UTFzdQfSr+f
NB6R9G83YwK3V9ZjO5SDfnaUDt0P/exh1Hj9zWA90xDpcivf8dizIwcDjx3EwLwGyr+98wB9HL/W
Y193Kn+jyiaxchD7LFYjKzl1HAvNXsVPVhM74bbBpkOFISFcsRzGPmBAAsZ+dSmKQNt1GJ4k3/2m
nl9IWFau+Q2AOb7Eu/TRp3qRFJDI6/VJtAVh4dMUaJVDGSODaPLN0SX99qjb3i6x3u3XdIIIGeyS
tVG1pLucNpyvTrT4au6wpqlonhck3vA/5Ko9R4ulO3t0jhup6dqZnetixNGy8iS5MqhMTTBxB+Md
VzvGTutgwFM3LS52XQJeF37NAzrfYsQ/RAv39eHywkwWCn7XmAW+VNWTEyacL1r+T3LaZyXUQaX6
It7ptc64iX+YiE1eDrCy0+IGIdJe6Psie0dCOOTvf292qJulqrCXg7zk3myuZBapjVz2OgPrdNyc
1emGUporr4pTvL3FcdCKE4Y0oAxTnY/q6mBcn6icvRTnOiLqCk860UR5HAtpPsW+EXIlFmk5Ium7
T9fIQAbX6Ibk+Ks/ioZFjX3t0nxzNpdRObfpcB1Yth5LJxegiORH6DgDPLEzEIcyQbpIWvADRbn1
kAet4/FwB4STr6vPXMEzG2V/RPUifJKMXk24Yo3UOfjD3jDq7OApQxjf+fFdxPAuEAOsr9+pTMPP
eeA3k7fUsHKpNa2P16Tl/j3oSgCpT0GIawSYz0gZN0Z8z+ot87Dqs+IlQ+gfEngd81H8tdwVZgW3
2nerXh3EVUYrIB9ZH5eyBBmhRs3ujjYbIFOZ63J5zwCz1zOh441uG63ZYA69WaepgRlRLqo1I9z0
/HwRyz52QaCCokiPpCSFcJWM93sfSRAPLBYFqTO3VLQ/sXJhLTdqhVYIF+lUS2h62TKKDuFvRMVc
y2GF0ni5SqQynlQjWsMN2FcR1MRwGFp1QKMqnN56eW1nommA5XrPaSke2l6gQAdiFlcS2Acv//dN
KZ7FnYnIEZbACBail8nnk/FrFKGecj3R3WJ504ap5kwgC38k0FSOg0se6Ia09YvNEtlXdoJ8fgJz
LCz4DYnmdPx7vS21yDVIUQfXRs5EjecvjuYmKNuUswoz5n/8HWGje6SVkJCqSBbbKy8tjbYunJE6
jj1RjlBnKfgOGLjxMVKXSsD10AkIt/ePMx14FEdD77E9zMnIQfqyz6iF/S3UUubrcCXBzU5MruOr
OqW9hgI2Ve0PIigecFfQyOtLG84oGKBF0+txoAVCj2hRsDbL3LzIvuXe2zZvepUgUEcAdjX/4adK
kW6tS9jvdClgoLIeZ9eOMQs9w71fSrDSedpobgs4SUVK/4rJx0ibIJl0LDwZMieP7efB4y5RdbIs
0f9Z7gC6L2zooGt4EiBdHgUuZZA+4ra0RWVhTJ+KMe//FoDpibUnMbH6lD6jhsNC68ar4hkBkXDe
aA8d2BaLxuKZnBGjiMvsQnRmskC7wuetSC/ReqTNi998z8afr9+JF6FnZ5X84t0FUsrG/HvdaKxk
4egUwghd83JBjbZxsU6jg4GQPGf8TW5hkiac6KtXp88XenSPWmzSmmOjktopQeSsfc2LxBXrYywI
QwbKTA9T99w3rjxOfO1HIxxZdMlVQJlXLoiHBag33/znQOWW1KWgGb/vfx8A1jfBvCnjBXXBhIbb
KgTClm70YpbaUEtSixGdGXF2cB4c9AZ7kJdYyR/lRYbDh4ZH1EJ6MVzBznPliHv7PS65gvEkZsMm
toU6flJoutlh8MWo4GT6fFOrGeDEoS6egLt8si03hDJStNGV4lpHrYqjqMeYmE5g1WeTS011Y5u8
fXFuFewBd7RmPimVAf89bfDfW8uDY/OMw295egbzdEc+5pL+84cdMNRZ93lLsX/Z9H96rT3XYsNP
ZJP4RSz2dVq/5sMzmtXBnlkoAO8gvO0rFmGeR66EzD4SLwOurFJ6hZ49YknXGc0woGZ+QEWCaZSF
M5c3oVSlSlneHwjgk+ex1s4OlN6koQ0wBqFaEXmv9O/+KJNo1K+ZCDlkEC52F8rrQNOyoyqSITe6
uglCKf4kNZSeGhy7k5gGqs9lIQFoTXeqVI52HpilXaPNzCim9WW3nGZQOyhBEWst7bnVHt7K/N/d
38+trUGvdQ/gWiZdh48qCNeAhaVJRQvvrl0OyJ0ShIcGPXtSYgRXze7/h/vE+XvK7XYjd3K7uPgA
LXZkCwVgnCBnEUk+ArUTpToK/v3QTzwKFq/pSlhPiU0ec/2a1e0iY9shSG9F6m3mY5IESOCk7/n5
1TKjoBBqtp4D64/UR+x0/fjCwKJgtKC7mmhcIFqZS3mMFQwGYoZCO+3Cs0ePcwaLDnrHZjmg8Jmp
U3M61dxPO3aus9wS0h00ndNCCPcIDZeHQoJUiuuHSILcWgQ9OGt3RE1u6w/T1rHP5W/kiJzyLEUT
/2j8DlXpcS06I2HD7jzDgmXCHj1/C9HYeFU+LDoWfQvcKZA+Jow0dJ/OYvkLC0DB0h2imS0xaIeR
9Ae66A2x55VGy2rvo/Np9hyHNwzgmP7b4UImAkkiMFJYMlyVpWDoc8Xqd3633fw57Wbjm/rqVT9u
IJzzVUV20aT16q+8bdx/oK9B53tFbWvTJHwLSf2qSAmUzpgOgLWoalsweIKeHYBsbatqtcqmdXOi
korvloUFzaioTYovG6O/yZxVAjRVfKFCRmLwzTEUyRuILSqVAy1JLBUcIt3yo49ATO7PYaD1+HnW
PeAzzhOwuJUT03+H2ukDFJOUu5XKFl3c8A+v34ENYMpUxk+xPf+yVL2l1r1iGz9Jmlpuw34CCyDs
a8YgrDJ848FsZInfk5fXjao5m/xtL2XT4U/EIPQXoXZzoeiqmEvu4UcLkGT6OxopWEXNlvv+X8WS
y9608QtnzgWkBNBYu6EvgJe9MvZciXkQm71RBEcvzOKwK8FmoBMIdRknp1Nc5B/r6EBtqYyQt/o5
x/tJTEReYFSXnN6fx2S4+AumQVsuEDRvwwwUBHgx+UiDFH/jw/4rt+JjTZ1rrkddOq+Mgabt8FqB
d8f69Y/na1fKk+OSsBKEfOkknXcw2GQSPjx9iR7C8I7BAU5iPCQNwnuffaHrxAA9766zQnlVqaVB
BLE4YBzrfu1Wm1arQiPCFspvdd70GiT/w0M2LH0PVFhe6BNeOMJ100RGWuY1QCfoY04FudQfvKJD
2yiiF90Fo28ybITC0oBRLtY7wmuZtgWl5Zc2dvrEC1GuTeEs3+jgJqecDwqEFe2tKSinZ0u5TLjy
cQPi+D8naI9mQmEIQ99Zji7XGYiOmZrx2+6kf6APk773VWyQW0ra/NB0SDNSktgQvSLKFfvKqy6y
Jl0dBrUkn3R5Arsz+wtGAtZcGcyF/xBX3ATrGUIZ1xKk+5cbhrFVPvU3n2cdE0PvtDSAbqcdT8oZ
8USXB8iN6MAqJI1Ava3R+X5qvFwGPCGlxYILDSFX7+enY5iwI86D7jFDo5DFc/qMNgrxvO4YMvKa
3crn/Vk4IYYPxhxC65V1IK3eyJk/K87IdBKx62AO9PLw1CL6ZrV80wmPx+Jp086PT3lBPHGKRsJ2
T/hEFOngLhxl2nrm6rhx4ovqSxwTvNl6odG4B4JfHcd24MObGnrUyawbnEP0a4CDsz5UX2+PbthF
IJnIDkuHt/TpdXxOHlgK7/9FrzjiASUZG9LMp4R7SHr13+MC/OBv2FiMmRY+kN2PwHxRbpVREXW9
8LDBTTRsrdwP1P3v5v4Q4wqJnImjXx5HMUiV6kZmyXH7dBdP57a3vSrc0qoKU3ARGCzuVBL5jbwl
y1YaUiPHzwIKsra/7xXwZ2eJ+Wtcfp52jFDjhvrSrd+cE2z1A0mmjghDXF2hk1OrzrM42mH+S8n7
hihGZMQSVnc8Ky6zfEbwrLYhy/ow3qQPGkGtoXn1+bQ8o4aaYjRVACEJTxHmANwuXB7TnwKFVrLn
Ehk7LYsuIasljPrIPrbljUzSWhT2A/6cL3uyfFQxWTESuf8RrIgp0VTOwXkLYdwaJmRf+qsKE3Mp
BDDI2yGg0MvqwDD/JOesHLaCmClFfQ7hzFt2N5b0ZX1LFPtr8buf26VC3avoLcRcJlmw0hTXDu8p
ApoKBpk87vpDCoRE86esaFBz0EPkMBtklDypSmfVJinlaYfvhpBtcbK+/dgYJsukhEa/PbED0gS9
KkSXpxOrg6Vq9eSUVSsD6klb9vJz9GAPSZPW3fu/uzHWOh1uw38+rJWQFt1vYgL67k0yl2QbI2hv
oSsLZEp0RFVu4nyp1TpqwV9KDlOkalB/WOnZTbygrw2JxqwB3FByKV/bAlAl5S36J8n6ldTVsV2o
OrxAOFipPTu+Ralh30Pi4BV90zgzrSAtNteJKPspl5LMmxdcnjdqbpmnjVTf/w8gnp8AjHshPh8o
QnLAlRfMw+VkaS7v4tADm1oQYfkUxAcanrv/iO7tz2z7StuR7ZOCmGxtMzgk9CIZethZMg13oRIe
hyl4jTG+StFCAQ2eCPicIB+8GUtbf5EHHEfBCx6vUbbz/UB81L7lerbzSOgEMyPONNFQCl7OiVUz
7UK5JHDtjOHCe3rxDCYHF15SI+Vwx0+pae9c6o6+2VMugM3nfnyMUiiw4lDPxrv1Zgy+H6tMcoKf
Ufu5oz3DxVZE0UtFvx4145O8HQFZAjusnkY3QBUTEsaOAqHTmF2IlgPy2zf2Q9/09a8xQ+6sGa3g
794K9K3jmSkPG/7p/Ae/e2PIFCmxFpZs3XcErqknKKaujIq+SlAbaVcbQEzZdxLJn4YIdz3tyg4c
AtnnbS7WAZFIR6x9And/maSB1X+HpoG0A/R0B5Tc8h47En8DUhxHc5UB/Bg0fhvc9K4hVLxemuNl
D1dHkrqZrIqVVp9si67KhqJLzKA0RGb8tZG4lz5E/Wj7RCU0hoKCpRkrRFTCI5hpx4P/rLAZ4O1H
qbh02C1r+BSQBQVFK7K5Xd3Un5e7Eu2K+EsvPM9Te0uCou3Lwpe2aOs9hiWu1y+bk2iSdpmAMPg0
s0+X4Nz3Pk5UpLqRe6mBthATvHx76HBSexknmft3ACw36rFospqw3pjzUMJ64kMNz39Huq97z3uO
uJSCjXNm6iMQgVaXpZuS7ATAAnQ9RTxWSNYpHybpLtJiqQeTjcZgrY/jkz6xynrgcMF1RhlZ1UHy
qJW3r6ztyrTO5H7K2DtWksjKPjNa8ai5kPahgLy4cle4ZYwKO8ErhxJEqA35R1dbXbspUwoBXe5E
j5DvTvba/HSiVxzKn4abw6uGwCwjfWdkuSOrxlUG1oVpW4mDokPAhxu5q1YdSrmUyQ6cUoAdSwVc
YM/DY03+pbmSfg+MAvSXnsyGvfWeggfSnhNAlJ7BbST3VHzXJFCpnqaNPILOFCx/UQreB/rsXChy
gl+SO8UcM6BHMYWzpCNFVH0jHx2isCYzZyysFCn5FTONbYmNsWP0/gscaT/jcPqAoa9a+jgq8Tzp
yO/ngXmlq2xE2GfRjp3x4mf1nDqEmnE8NU6Qo0Tu785X1/mQdf+h72THhzMhv9QTnC3ZxTiExDju
owYXLIGrkmc22drMdlRCJ3Ii4Y3nMfEQlL2xYh1Y+ap6hH4PAvwiT5FNJrRjYBLRzS+hS0HKEzz8
g7n+H7/fdSaJPOY6rHFl9n7PCiLBzn1Dk77lb6Pn2IWveXL074dHcKqWgGBc16cRjVsyCau2sUGw
307req1HQxwEgCjzRBD00SKfyNOKdSCf5aOB9s+0XRCOta8DQ6hY8bVuGIOBGrkYVpi9BDWqggqc
SWwkE22XPSj8JJcuybCwFf8VZRR7KzeG/qoMICaYDFi3cDVBb9uy78hVZd3CKnqVEtkaJSV7YB9q
2Zrv5mzQKmphF0IZEpyg6fNAvK2sHZe1xqJQZQa/uS7IgGQwU81+aixlAvGRWhnLEE4eOgwKEGZC
nkV9xx6snK8YY2QDYO3wT0N/mRdevRu3UWZcVJKdC0ZjSgfgBEDqDfSXXlRxkLGqaVH4CoaEgayK
9zTBv8Zjbsb2EPW7h/PHGp61S4qlFtckYTehl6APqzfZ00gWmZAbj6mjF0MA9MRsyBkFXO5DhNt5
8aR91aGM8H0LQp3fMe7aWXTnppHUdZX9SwkPY2ARyvXtZViDfC6LuWUYD0GWcW8SbtgGfv5ylB40
d92T/aK0hKidC4XEBGgLLWzmKHLHjWQYQiiRjAyUUU5hMSZMkDG7bxmo55EE8yyX182ep5OB4HJr
LtCBLF5ZM2UVi3+w+e5IDTJ1HRmaqDegqixKJpI1pm/iNhvWOqtncc4HOw+XkehK6nPOIp+bIZiw
0rUHfsfQkpfgjWnN7i/6BRMrktQnylrsjgdfno9prcPtvudDZ5dNP39cYN3mX0d/aAoDsiGGtjyy
9gi+YzrFXMfEN/P4ve0JXeAwdlri/fwA3Pd2PrjC3b8vht76VKIIL26+4HqlZTaKqs7ehtpK3CZa
YsnW5kyNZG5h5n8beFqfSdpvdOzUvGS5nVS8KdL05eFeGC/dX9/dXheyZOGhoUCGnQWl44Ost8FV
TH6Dlzc8WKk6OJ0HhSjQdGbEbEl5/Njlo5Cme/y6yJ8sIjcQHK4Ca2WmkvSG7OA+0/GNKQubSWpT
T2oFVKncnspDzDwyYg9POGAjhEqzYKEjXTBPOgJiPl1hHxNhuxZIR35MI+aveAbOEfTN/PgkIdfl
DXuOld5KCizCWyXKV2iMn7eQXo2ELavxZGjfc6eBtwQDSQ2M34JXzaRHeMyU/WiTXVJM54NSbu3y
5aH4qtOMSZHviUKchrZ4emK1nlKP7z2SC3nF6Gi/smUQsyywLHZyeF9SWjvhptmrE/m2lgs0SXxo
P471S0rknMb4CibBNrMnG2oItc4My6DI8ZtUh4kNS/6IgAI41HeXubTBRYp0DzdvsFwET5W8Y0Uo
7zDUQwT6aBFUOPmsNpRbZVDXIOhe/fwzq/AABqv+A+PXuVg7LFWS+X6p5cA6GnRvdfLwoVFPPI6i
I4B7Fn7Xezu8vQCOZBPVSESm9xu7IpwCSdtWwBbJiY6yl2cLAUY2O7Q2SahzZW5zeJCiU8NeeLxU
iz4PNRFVJ2y7hrG1kVWdkWD4p3I1A6unCElU+DiPVKI6FT8JTnn+96N7pyjH0ei616HpVsX0K52p
Hf6nekfejSiDJISQLWcyV//d+g7VpekrZzmJ1WKBoPHL7K0YfTxP3xQPAyHXvNBC/yFH5pu2yRIc
1jdjkr+Ph/mFvFj+yYQdYjSATrJoPw5A3kJkhnAPpcs8l5QRR4xtCPtlurhm8/ohvG1oO6l76Lpg
TKa00ZJKKo1Y3ABBbhIl5qiSzYbQRFEUNKJ7uSpz9K61Vz4EykgkS5+7h711DIwuBSrCzU7vH82r
Y4m3jFtNtf8AjKA+QKeV4Ujnmfng6tOctqljLMiNWiGbG54SxO7OlJVfzbFYpqhio/JpAGrTyXeQ
rf9rV4lwrykO/cEL3u9YnJ8A8Pp6St3U7JMc2nFyNYDJ7AvhoQEYat0JxU1ilpHvEwUWW+48pbF8
Tbn89rbL31Y+MFhjyasAZAZ1Lfxql2hjSxvP8TtC5fbaq+fm6dmsJi/8oNMG0pxQ/lcNYH4jxgAH
EHSlAVT0tLXEuHPvsRRFdNgnDPJq7jMUw1KR/AQgECJF7FC0knMXJ57oe9prKOU2q5CDWWQU1i7j
PLm8YnjB7BEEfdzS7+xgqXhjhvvkLyhpnSfXPTNgriZxJclWoWG5wc4T5rsrj0kIEUz2oV7WztAD
x8NYw7wZJyCxQFyVP2J7PI3SzH7RkIp2Nci2uAenuGrh7YYRL+q7G1Hhphg2LyFDEqEdQ7nkwZTt
bdLQ8PWeokn/bnky2c09ra+X6WphaQygeMnSWGYZa9bxO6HgDR1z6/ScWoFoqPxbLAWLMHKsC/WB
PqKSXi5tCdJqDhaW9LlsuW/UfOjhEc9aU3TEyIMWCWzQzAULT+W4AcVRwgKe9PkaxU/Pg9bacblF
R74QyFjW6jM0MQpLfCP00zVA7i0/g+ZRYM/SL/ePzkh5WaebN/BrC1H7g9cUX4ginvxnutuoVDUm
4A+9e3Y54LOvTR5+1HxEubrFRIho9/r7rVWtf3YEA/PXEMTQvr7c3Wk8U+BRIUC6d2ZeVuIhBy/F
xNDMORcuFuQJgTf7+J7TY1MLXtMFUH4YbK4PmqUhm1OWbcGpSsDS5pdVj6FzmJJIvcNNtxgMGfL0
G7A=
`protect end_protected
