XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y��Q�5:��i?�A��jz�iv���nM�'~,$5ӥ+��sͰ&�h�j��B8B���h�5F�[I��z� G#�G0��v-�oM�_��<��^5p������@i`mѹ��Ǚ�	�wϺ��mA�#���Ht�T���n̏}R:�)�YJ ���ޞҀV�Rv��!�#�����e;W�Yt��G�=�I;B�#ȣ��ⶥG�4n�Y�k�E�+bz�kk��N�*���bg>�^�����#;� v��^ӳԯg�8ȯP�%�V�8��I|~���@R�3��d���
���=�Q�2KP��8yh6��w�N1��-��	4�Vr��$4��޳_�L�n��E���N�� �b����ߩD��M,�'�� ]"�o$Uq��tߴm�um�����3��R�
+,<@�ȭ򟆈c�l�+̮�/o�����J��6��%�\6;�>���GueU����
fۂ��ُ���HU�Մ�S�*��!#�@�:��h��*�����a���gH�Ȋz@�,��|*$-���1��G��f�g��F|���� !�9w;�C���-�@���1�#���m.�]��T�~l�h)��Q?ªc���;�b�'xaՃN��dE?��(͔p����Q�,؏��E�����Rk���tL�?Ɨ�J脴:z�=���4���p�S
��ѧ6��sMT�_=�&P���\�2Iw��x�)�e���׍4����!Z��'z� '�x���;c� �8��H:?_�\�xq�XlxVHYEB     400     190P��K��K����X ��xR)�9�w�|}�	D��ў����#�����,��2��>�v�5��%��ۚ��=6]%��[��&]&�+"�T
�3�������(��� V����|yx�9X�PWq�o~��锋6
=�YR�Ŷi�ns������x�bP gBD`]��[?��[�G��>6��A�F�
WUz/7���g��3�I�O�Kt���!LBE� �)��M��0n~u׭q}ب�Y`w��~�MS�듟z2a�/�A��3i�ǘ�PV[J&zz�F��O�v�od��6󚶃�6��z�z!n��^b�qk��B�n;#e�s>͝��D����Ȋd:�%|���}�f�8yʮ:F�:��0)lR�=�*q���0�uXlxVHYEB     400     180���>�O�Xi��q�]{��q1ǉ-' Y�Gi���So �(>��N�. �0��#T�l��0*�۵�I��2Z��c$�~>�ALL�g�6�55�O�2׌F�zH���-��OV�(�l[�M:��"%v�ʒ�51)�K�Č\����a;��@���������lu�����sp�x�x�7��~w���=��[X�`�^�r:�b#�B�����Bl�~�C�pq�x=Z�OK�L��CN�K�h	e'�J�����ڑi���ըm�QNY�潜��.IO�	ճ���~z��:gN�����eW���lkO����^���Qwg8d��װu�����8���w���K����o/��%�����9� �ON���`]��� r8qXlxVHYEB     400      b0Бӟ�T\��!Q6�6���Z�;�~:����>��y
���.֏�O/_V��@+�]#��!v�+���'u��+τx���nzX7�Q�����)�����R�j��r���%6��]�O�0?�"=�$b5�4�MC��u�n���<V.3��x��̌�xpZ���CRg��M'�XlxVHYEB     400     1705[������-��5�b:���`Ρ�t��C�������?��H��[ʴU��?G�mt��V���>8�$^A���N��^��A�F'	.�_��z�u��b�C?�.W�,D[�;��D���v�L��r~JX(��Wz�'HĴ֭С-�.=Ω�r!~��j)1鏻�y�*�gp(�T!���0����U�^�;0�Fn�/M%r
1�ر�Me�@5�W��U� �̇}��M�3�=�ACR�s�G_@s����Ɵ樮������G˒ '����)Lr)(�!�e�ӯ�6�0,~�e �۳Lj�#|�kyN`L�����^3ق*ٌ.���8e�9AEUёx�������\�1��XlxVHYEB     400      90�.g��1x��ò��-`(�K�c-
!�Z�]�>g���@�T8d��V�~�}*�����R?��!� _?D"���-��rI1���2��X��34���a>Opә5�g�K�V�x'����������!b���S�����oVm��XlxVHYEB     400      90r!4���Հ������p������1�YSS�����ہ�V拰�L[�b��Jb��2Ēdj�mEuK`ɠ�1&��B�#�����j}3gw��|��K�����l9k�u>eŎ䙎�8ɯ@s4ݸ댰��� '����4XlxVHYEB     400      90��1T���>
�s��M0uu�+��j�"�O�5� 1�ڏ�1���a������!0R���?.��\,8�k��{˭��s}_��0�X��|/�'�z-#�5�R2� �Ճ]����W����h����~���F[$jXlxVHYEB     11d      50&���a{�nO��Vz����ȳпM�I�N� IKa�<|u�>To��ŵ�Q�mt��%C6�P]��RǤ��PZ0 �#�o�