`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
aBkTzut/ru/gHzvVLS9J7dpRmLCM2CECNoAHJqqwTNxF+eCYkcAU0ih3wKvUdadZG5hCj+X4ulNj
FWsCSERhQVr7FEuQxwGGLontAsfMi9vYFCqfus0BK43rY19+BnG+KAH1MDvmdcPKobqFdXHB1/2R
D+bgT3pSjYV+cAHOcbbW7hS6nDza/cSrZhiVJDuuB19XBjYRTQHxo2+hfO/JvCf2B3o78mdib2La
QPWmG7o5XyuLcam3CNvQRtZFUJxsNOq4AsWtyy4f9KRRjzTArezWVHtTGaDupRsnUStkhCmVFv6v
X8nC0SQzAIyFQ3FZnWPePtFy9H4uU9OyEO9ea3M+XmKmTAUmzAw98fuDc9qLsQLRO18gAxhfZp0L
Mswc5wc1ZqBs8SiSqe+wSBhqEFhegb7xaVVsERZAYXgPBb33p0bxX74E2IK9Y8pKS7G2i60Lr7SF
/wQ/sz5MuecvzZ23DhuVhFYZvHK7Wiiiw/o4QkwqFODwrPKZ0qU9I/3CenXABzGmkHlZMe9uL72x
yK9KedHhFyFbme3lzb7nzHIMDs1HIwHRsM2Xx92/jg4hHe+Vr8AT3yncx9c4deXhIX51+d8Mazm0
oBgj7lNR1xSjjU6zkD5ZyAGwmSbbLUOYN5sDemFAqpqhK2uqW1AWF455SN8qDqGYXJvbXRxddZ/c
zAAZPnllmJ+MmgVG7LPbth0qrVvVxNfL8Pb8rAlFXAaRCGUsDTQZLtFmu6vJ0/v60ietPNlKttCC
9WjUsqZEvqK8IjT/T9NK0Bze+EmTthCtZLMT0FGDBxPHuZO0FBgcsh0WjPy1oUfO0rxvf/5BsNyP
s0YBW++pGmlnvt5mstWRYTgik+5I5QUw2sAXks5Dv1TIqqUUkFmElxE72M4eNYkijAfpcnuqLLFv
+amqwraweR4E1GLPQWkrGdwyBjImpDbH4cG+Jnw9EhNRfBVIOO/SCb5YcDsBC96Z182t9G5rKDbj
/P1gHmnMQulki2SBhrhiLvAMyvngX18XNq8htSNRFIOyKSVdMEN/I7Y9lcpNE46b+5dNW1lxdBPe
d75nedsNpowlD9u3xDArMe+pm7PTd4TOFzBJNAyGJDIH75xFntBoNUzIvLGapRXBo67V5c/9D0Yq
IgXpb+SOOKJ2uMw4XWUTNurTuzb1fYJUePv+jlhXnIc1inqtFN7XVwgrKFNmGCuNpDJ8wvO/Y0pS
RZ+b545B8hdXh2SuC8fonxzhYoJwnJiIMMIxq5PMS71qG5/SH+MNc8C8nUazhq/QHS0WyYNv3UkZ
013JQOe5t4F80p9/MruYRZBF/sEDOF3E8KXTVaBWUTH8GGC+0X4DMHHgPd4ey/668VNjujB8t27m
1GycMSjhozmyZPlbyvRLQJNN71Y0sx1kMcH5EqpSCWh/3dYNg+9uUnDEtxkJr0qzl4oCVzEgFmK8
8HFGCqXSSz713dyU1vSTIM8qQxKpTpbPAp7n7jzRYYes67iK4dpp/cyKmZs+FMd0h+V8+Vn0M0/t
KikHzCe/SgQ+KIel/Y/0SlPtLPYcG/pK2e3rnkKx1HNoown2jv8w+4uIFkND1CRgaAZvwvIZR1Ky
K4ALd3M1/QhwtRJNo0Bxptk2/H4s+Gz0Jc1uTrs1QYFeo+ZtdFs7YBwALfBaqewK+cf3/dPwcpbg
JBjXSVkTdR4W8k/HRhz0tq0ogZuL9O9LVAL8f2i+QJQSqbnmGpjQwvM/gNsmhzcgsoOTPu61hXQf
t39h8NtbsKZgAtpSK4gbbLdUFAM/p1jtjl4QsBY/TDq/kzbm24JtSzToaw1xRh42RV3NI/zdiKqR
f8OczXQaKEr90l05l5Q6vx649GBBJPYvRR9r9dFgq70HZhWree1JDUhEVCv3Pk0PAjSwDoCeul1G
8zsjKc998ekKXMv66oCeEsMaodX6gtvoQCeIPeUG+A49G5del3J1Gdvbpk9nEr3KAdVLbPMzGnSV
HlIi+qGx473zJANwouS4mZAObEG4HpUGAJ64Z00FZUJryeTQ8rIbNdjvi1Mgg7ZSdW+1qdOCuzDM
L3jKhcfkDdyxtJP3JRVuKKS7pm/Nz2TjTiD/XeQoYv+f+p+bgtH396Asjq55yGmjCWfiB24wAtVb
U+5AmtXqLS3s1nnkuqjkQDgJHVNbGFVQM76BYp9kP5M6gReztDSkri2BcvNe6oizDqseTL1PLepX
naQIqu13tfZqrfI/meAN7UwuZGIJdKxb4w3uZwFNrV7Vj6FQyVIeosXuc7JvoCZMpfKjhlH4ENys
qc/hn8OzCr5grYZgsA6U+goClyYjnfeG2vBtM28g1ykyNzgbB24fmFYC83iKyAUKKggH4cu6/RAA
iRf2WaM9QTS3FFEmFBUIta9UZVg/Tyxy3kWkAShA9431/5sbps7GsxQHahE9Bt4ohd6EC6x+3EN1
+I+RZ215yzuU4PLLQmDXa6ugKsES043t1xNJzRB8hV5mgqNTb+60FBKP6aCo9iwY6mCkRzb5s7Cm
c9+oAw4Yc+txQCQ4JffYoEuN3PuNqec55v+z27a8sHyOjZW1whXrpb5WL3T6MtCMEwo4XOvgpgsc
PdYkilMOd+LXEKIbORNDZkJmuYd//T3nvIqf345fdrqT+re6RTD1CYYleTZ2hCLMpu4T6dqCRb9u
AdsszYn2HTGQX8UYaM0YVcO+7IgKiMkvSM2U5MYaeFmr6RWYzOz38CcgFCkaa0Ch9v8uJWkebcPz
G54bcGI5oH/uZkrIFoKOBrqxC2oKuVWRd1jz3eUKr5dGPThm9JrGgHEUtuLJij22hsAqMYru4VIF
mPPkQ2/Gx0wXRJXwRfC24Q3sEgL4U6KE6jOBIuFkx7yL2HEYUseFYOc9QNG3WZewt+K6//GLpkvp
WzmU0zmfBlwZHqcVrYxuR+pTesnsQAFO1bCYbKu4tfnqfuBj8LZNKMVfW1d/0w7B3ouHkgr9oyfV
uxNE3+lY0nTFSci3QnNR6Vl2pYeSjKhxqE6YSnoivsh7xwhXH7MRlCpbw+ODrAXy9BbLsF24v8DG
NSrgEtkW22BQa82PLvinItwf5GseRlgsDXd//KzJcZHxgsdSnfbap+X0kYPyW2U2PH0nfizweMj0
kAkUP2TeewXOaVjywQ72xcqmTe7wMInWmmOn9SAePxVlIsbBUBOQp6YOaVdFLIi+LdO3wvTmF/T+
kisiRxsF6rBYxQy1OFXwnSZN0XvnNCV7g0LX74vHXGebZdga1GYOah8bsJVf3sH1P5cigQstw2Am
SIopDezrYgHKl2tVSmU12GMbk/dxYqJdRUUd7OsJpPT/e63ygFxqQMzimKwPvRQOOvBAOCI6LyQo
KqwVa0MflJmQ/+L5EotFzya87ukgZ38gAgVnXdIU6VUhuuypio6wE2OtQ24ggwtjpOoieD2BCYvR
o1T/+PF1ZJlqWcsPlNJkY93FAA7eiU38Amq/4sY6XQR8Kr5WAHywIlZWQGKEifzVMAttRYwE/QbN
jNdOBpUkz/61brmqwHd8xT9mB1y2LFDbaxvEFRctNoD7RPw1TJsSPFSBzClPbCi/IBaSVQGydwVc
46XN+r82V1+RJ2Yfg/jyQPY6h6sLt3T4+kTbQArwOIcqUp88fqO40d4EiPv94XlRBv0KZ+dPo7I7
fct6crjulIHdJuVv/n7b7aqHrkCfPtBYB1tDYk2xjVxQnrQ+XEp4U4InFWzaVxi0ChWBmBMpV+vv
ptgygH1vvFA2BE6DkKKvcPQvDUqx6dIjzOZpZtRusnit63LsuDmjBqrXgHQksFT/fbwPT21wlOMV
oxBPaa/gtIaeKcJ4Ylu+o5nr4asdPv2nnNq6prG1EeF75TeI1qr1bN+DP1D4LNZp9Cs4Qyi61WbN
7bQgTxqCDUj9nmGwLQD68B6lBqS4ZMozNWzXtIlqBb0PSURUi2wiuo1+A2x/3EmlC97s0lSrX4oW
okFEnpBJlODz1hqBdIJh0z/AgheCwoUZugAv7sb3fM7bluNafbmR5+DY9OUHEIH96Ml90xu5vJdE
J0QDaUcLXjlLgf0XSGDjS89UE3b06NO6F/NbIxa+f24hKREl6UcpdYB1kDEDgn+8Z48ZgPZuHZKT
wspL2MtEdQiGnSHvJjDbhnsFd+mzMGe6CLx0vBYdrILjlgVm0T+Hk1JZSR2JO3WcYAJFbPcQ6HWR
XHziL3DzkDRTvXS4fCa1EJihTe1G0hbKGh5vsydydbj4z2Y78DZgFt4Ts0hX835NRYIJRxCmDQJD
HxNdCaiycxTvI94+aUrAXXGRZkYNK+2uzw2Sv38G16hYB2Kpq4AtFhtBWhacNfKw1pp7mMPIzMw3
sQevMo76QnZ/um8VDcuCYor5+JK/9N2DF9s4BXd0D6WJs1eV3CTAWOYezXFX1nnwoYIuMZqjcp5N
tEmyqjzlz0xwO0CfTjSyQuAJu76yvwWwQJmAhqgpxMipTqYx3FGhmwjAvKjTCKZwkACn7+LjCvMV
LXfTe6/mGvMbs7DaJbvXxScEutjSeQ3qWxCgRnWO25avT+PEct+9Q0JxA9HjtTc9q7C2C44J4106
eqT5Q1ijsnDi5oHUnodcw+O5gH8b5FDnoB0f0ss12AGln5w6jOfSQ9qSx1ns3HbmpWePGxDd5E/G
g9PZXwLSfQZFgVyFuPobEs1gRBkL3I2LonE6tNjtGiZwRHPzJkWqFIYNTvMDqe6i//gOzNZL9Xoc
uvWAwmdsIA86kupM6/t73nJMKj3qTMV6FZrsGqa/EUuLx41fibP60YMPue/1CEgbaNf395UWUQai
8PMRxyHn3oFV7c58KJodPuooKucEznUEKCITCuZzi7HM92bOGZ+52k2XDb5X5apHqEICRcc6ubMo
2OiogfeROB72i8cKviLVO0rT4rVafCg6u6AO+JoZnPF2w+Z6iTZrjU0Lm/TayudaCHe83DiL/GwV
3+jK9OS++li3rpw6KuxxLTFvG38y78kS1FSWYPm81A7PLtnDZJIQbcCOeXusQF4Yotrjibm4s47p
kkH/Uj84LLn1OW3ewiCAQcyRUE56SjBkqOsz0XBuY8pNXIfyxpy0IBXBvw0xZnKgrvuyH7YDadKW
ojkMFwkx8WJfD1mTIqDHM0D8iBpJJIbedvZ1uzkGEdMzudq8VsX8W9LwjM7hd1GIcxPI4n9aRI+o
dfMnCDFtTQ/BDTGnWFnRnzrFVGrbvX5BH83SZw8+ER3Afv9m9/9Q3COpfzP34DoF/cZVjEinNkp3
xY/7A5DIfWeGLzotzsOvq05VkUQCWFb4bkSzPgMejVeE6KexRsH+54Fym2EMOPlOP7w3jXf9DxI4
Vr6tkluYtjBkpLAjaSmJkjn7+VmWHsb/hwiZ/JpLWKrTnZuwSUgM5L3Csr36GIhd2EONfm+efPLn
XnlJP6gGVxG+3oL68yGCnFlqDzPcePwyN3Rn1c3AiByrjFlAnYv8TzVIS2uVLm+ecqKTtUmWsb84
7OyNceQyqByyQBUp+zeDjrbZ/toAUMOG6mPOVuzVMpVWOhQ0wVBQ57g2y753ljVzJdtUVKF0kn8k
z8BbTLJgTz9V9+Y7BJlYZdKeO48b5H6EVEfB7rg9qitGi1m71Qna+Y2LXM+DZVd1/Nr9Imc763JG
PbyKmQuRRpoibsfyxBB4H1uQ8ehwnVAThdx+5mkfKyuPqyhiw/UIPHfUvfyh8dzBSZDw8oCEV3Zq
2/wvW4SY/eFatlB25ZNG4LujVp2QkP6i7JEdkfmOA5TB1BFDZvY8qOdCJs4AGoXFL56gGOKSIkmq
EWZhkt6fX1bkgwHayjqdrMwpmQnZL7QhcXuZDvnvq68XQE381vMuE8j4+6UjoYF9f9B6GOzEql9u
bFv53+FijVsUy//yQ2Bg1SpuRyIT5SYzyoxZLL17jsfyHqUTz4kBvSCUbf1Hmzdq3U3UEUICwf70
uDSH3KSw6PO7owmXx0XZsgsITesK+S+HqNvgs9rEWBEgokcG6QPXwjnkj8w27S6WqpxceG2BrHpG
M4kr20+3aOfVrGbUwwwc7LqFkDiGYMtNUglGp17RIFYouQ+wZnnR3t5PdPo4EwQrR0Ryx8Dtl2GI
f82DzGmT59gNXo76+4ZxzYYNX06zmi4HQYDwK3ukk9TTo8onNG+0gF7dBn45EJ5Ik3otclNwEKv5
CMHLO7oHBrVvpigDrgPSJOT0WPoHazkqnI6ls+QDOxQZtVZ7fJOnqwvJn5nkq8ZCEDFWEza0OGBE
jzx4mv7Kj7wYg58LwEvEM+hQWL9nV19lhCRUKkpXpyfBnJkDfOvDPeTZduct7UJ8Ljkk8bk7sQn4
4quLUzvE3RwcNqV4iNu7NrBwruErKXv4LcJojdyHaXELzc5e9mFs5qX6Y+aiqqRh3gyuHHmpf54V
ndUDvpkOYIN6ql/uN2yhL8q0KrQwz8BoJ4ihiYNVYK1o2WnFqN0OmXtUkFDQG3fKfkj8SbtS+UKM
7x8Bl/1oQIuQLycqycn45fXcQuEAD0BV1paOBgwRLF8c0hpFfOG3Hjbx/B9S1Qslp8oU8sSz8c32
0G+rupAT/T90sBgGrqu7YywB/qvFFRURyvapiYwyErKpqmk27IP1TLmDIrz8clKSTf61oIlVppnk
vum8ahKlWFcsm8Yn5LPcnkaJSkVcy/QEA8jIQFByGy24M/v8eHM2OiSQVdXuFBgXcR19te8K0Ufb
ekrOHJcjTeUNjIY/f1rnXTxG77xOedz9fPlJ6n5PtDQg6+13/QqgGE+e8L9DB6LKAmsPYErJVtsY
kBUvuQU1SP1XMMv3Q4Y4zjZH8D7rrqK+lFbynzYfHl5my2qXoffSy6E6mUCe4xqHCGyc9cF6NwUc
Jb4jLqE0+nXImskUK34A7YcAcdqV8d9O9eg9qc85nFjG9lRZzzZc/choBmTtKmboVBfvwGjw9V/N
+0h9SP8UtopmkwRQ3hHKWynvr/S7N/6w187HTTVefwJcBARkQ+id86IG9jUQJYy7N5Ju+H+3cRwv
hRpHGZtPP8uCo1gJ8ARZYxpd3C3X9XMFlxt8HNb/PKgn91gru50Zs9OdmLYhAbxGJxf/5sZfVOJr
cyQGJ4VjIFuRIcDYQfQ0yxdZQ34PWRx2/vFSsEzlRCxwXKROtkNrvIdd7Xur5Gg7CawmNVXjiYBh
p1fW4UDT1G1vK9lU02LXu6Nkij1bUZ7yEFpLhL1P5LYUlROPiJ2BB0gTGet7OnHoZlN/jAm7DOz1
NBwNZZexaU2lAvDBYWFgJe1iUFxET8ONbpQVhhAAB7iiZ3p7WOza/gHQGh2kYcQpNXmn3HFPeFf6
w6LnDexr/SNdgW8S6fiKG2GpWVkXhlwFWBtZCsAmSDVupWoBJmo8cUzD2a8jKBnlkf4YymyIq169
OFL1jNGQ5KQ51zOFGJzsAbD5+3xfFL8vmB1kkHavx6oP+nWwa6ghbPgij2rJk9eIGIi6TWyUJlon
TErsagpUVLWuaOKEwOvltS1ZXdLY3AwCe+F1lSK/ged5VLDJPePPYvMk/J4PYWn3twbneXYeps+Z
VignefD2xnJzHp0cv2DSexiMcW+vwTpvBdhM2cN7RApcj1ACwKEonSSTKzZb89FtoiaMK5dzDqaS
i2zLpUdvWD3YZRqCJWdXxKVxauGgvR+wBHfpzCCjdNv1CTajjgSLpw7DNckv8LNQuW3y+2tZT2f8
sU3E9n882QrO/VHodKc4pStC05iUNh4cH6U0c4UIgHiItRjUBOOJghYGkGaa6hl27oBlIRuKPUXG
PH/FUE3r8Ch8nNflXgDwpCulxLPBLaeJw3g4YG8GvS8zjV9iZ575FTumu66k9qkWZARcz3scUlV6
QY3j4TKRHUjIcaiyFI0QLdyo68SU2zP2DEeLbpJGCZQGCw7ByC3U3EXnkpf/JwNiA8rO7XEc7roZ
Y2EWC8d/PsLFmlik3pluwsQE/wmjH7DvIk9ftZQ1CC6M9LZGwpMCs9luYJ4c/lPVJuhYCZbVU07+
Chm0A5ORb0gZGKIFn2g7DXiPFhgeX+axunhwGNi1c3ihWElE8SZJ8JZ7Axm7z1d7fumLQeOC/exs
cIZLRsAuZr0CL02+5IbXN1ETT2rvnAVBGZGfMiOExPcoASk5HGldZ1PmSBCZPD4siB4ZHTS8WM2G
Sa360qAPFS2N69Z4nHUPeYe++XW9ShVQqnhKYgeO1fI4SnA6lWPQ1p0A0KkbHwLO3QT5ZTQBhUnj
STTivpFwtGXDKwzVeeDPryWeHbvWUDKCqCYQhpktHaj5tYownt2/gf9FfXb190EHc3hnBqKxY+Zg
Yy1vOxSk7XuH1umIK968k6x7ZryfK11fnSMqII5WyuGYcdqJzWImI5+pUO3zEFQWF8ySFJUMXu8v
V2WzAhemU8eTgCzlx4dL8yW8s9FaURGHkjM6owU3TXO+t57NYglXkDcVTYPtCU3Uxm43dU/kjALd
8YDFzkov5M4D5rNWSRVV5SM4MxIeB97AF5bYRADF/5AkPh4fhAfn2ewLokZ/5i9nos6uPh618QQ3
058rtAbhaKeHA33Et+LcRUL7SJT3xWOvWtXr8/bkaGAu4w10I9naOe3+vc2z10wMvMXU6ZPYY8QA
hj5Z0TCr64/YSPEeyHRUWEC4GRd57sGFgV1nVKit7upoMymtw6ir3xmJWXzePDQ6b4HeHrewgxRO
5rl1wUGFBetVPA+nreWFLuchf1zk1jj0uspUIx0KNoKvR7AOdKaStGIBw25m5wDpWNqXUaQ2MHrP
xDNV2AkJy7ZJDl6HqDJcliOyX2D//ym3TtKMQjDtv6/CoKte+dfVfv5tpQQKIUPKD+MMH7QEa3Zu
Agtd/AfolqkWRs1JEIoqF3CsqvsGBXPPseSDpGZfkXqqIxuuXbOhVaGZCt7FWnpieuJaaNDtcTEL
n/wRni1XkvMEi4M9hwQ2YfRcaElAl96J0sgCiGruSDMnvLKfFdkeU0YiNSDdAzurL5pigRe/dXrr
4W/6GjOOgT81iBE9t8N9ESsw9ZBrFYvBUx2kmCmC44BgySQsqiXiquYw9+efu8NxN7Lm5na8b+9d
ONtEjysZIKxx4Vb0B/puz7mE3a0CPbcB8luIqNAgrvBtNTx1Ks3IvLQueptwpacUhxAk2dtkXGfn
HxzB0OTts2Q+NxXY77ZRWGz6aGw/L4hHoAlxeaczfD0KBUAgqy3xRTBw9p4Yl3dYGjbvtphAcF5o
LdhekYDX7bmIn1ef59at29tG4gVbYM7rsvNzIGZVO6iq/wYfDNN2CVsux0G9DV+tZ7FdAaqgZ2v2
v7m/Rteh7cTaCiStOWndZUqWOcrlhHmvNrtjvzINFTLqvA5ezSaAEWW3EI3XxT3eUpSuaGKjXOhv
OVg9OP55P6NsqJcGpH4A2R6ClxLNoT0FOuIOVkW+vtJg6GiHWDwlV/rtUqHpd9N6Lr8ohIPcGPqs
HFJmNPs5oDap5shL2OFDDSz5Qze+njJIMeFHx63YTi6hlUIs7R4QwfPfBWgRiuR6j8xb0qyPFPfz
LBsFCqoL8z/zJOS5OmbWJZ7PHUhYMVgyUp9oQjySgmbKuGZG7hphuXbo5gWPwLv1QbRaAR0tRSRi
jsHnRwhM+d5vY2XPoyPx7ayDs96I3ao6quku51MxtEtvDSUq+74n8yrWyD/849WeiwyspsezOZOD
a8nu/pDMRpg/8cg8dZX/+h6eTvWbiO14euPlWPwyxvYFP+bl45DfG7RMezc9jTaztfn4v1neyFxq
V0EIqrGcpbzuL5Y6137tmK7b3D3TXOshIs3+c84YV+ilIlM0aMilRUaBuRTXQfjHLcAXDBIcy2AO
P8tWKEg40D3X17rfJQf0Dm8uLCX6FUr8Vpp3k6UekD9uVrGSDMkEtzuQRw1cV6xlzl1wxnlX/BF2
zTEaIlJS8fcF8w6gzCQwv1GjpqVJxnnjO38aARTeSluaX/NztTE0tlARHq7xGt3oeJb68N/v73DE
gXjb1iExDwpWJF6XcKb7J/CPKdOE4sSAlpWfDaUxvt0gk4z+yKqpyOJ1AgOKbttbzo9VIp55zYZu
K5ButGDi7oEVkYU4ZcdwSXbWy5EIZnva4bzYyQPlJ2ry8B8JCUwirTtrlivS4lV/EaFYH8GwBPvq
ZKoWjrcqxCj1tc+0QWO8mIGihMaRN528z3QRe/6kzleuw6GXIVKRVh6HcHcoGKx2W1oxtyJ4UX1c
61MIjn7ymWVBrMbc8L7k/NupwlzRmc6VV87Rn3/163pcroqiWEHkfOaL2AmKu2MsoZGDGZ1JV5kx
AaKHuoSYPMLVTUz+Xy9dxktz55mmUMHUYM+Hnnbe7sR8ybnv6TEe+7xE+tBx7lB8bsRv8yfyV0Al
blPBRinLZhEz8bLUqIREzkYb68mHEf8yuHY7Y8Y5Jur3QnQgHLIRlCiSdE3PNSu+8wDF/wknr9sE
ixYmHb6f+WW+sGuZTeQJKTtK/EqcqjTMcSuo6fJQNwZrA72j/oadZY0rYXiYOoYlKUkwPwtxN2fl
0xgVbo+CmC/dOFIQeZ6gceVUyNEByuKkIWeZr2ATN3Ikg/qHpkPOfL1oh8rMzdgJSEFDfNF5OUe2
9wJbFh1Zg3ZpCmIOpHNdQ28Vf6CzCkv40Ed+R8ld+KuEIrr2s4fHKHdvRH9/Ia5V0QMi450gdGB3
cOStTZOr7MxBvM+BtHn1W1/XVmq1r3aa3E+bcQLj4BGveI4cdxoNdMjk4HOUKRa42XTmUjmj3LQm
ipZCYiMclLvYp/JmGJxA2SQLDNMyWBqVd38Xyy/sZxulOz1zABMAMKO+pJNrXlLj5uD0/oFW9BRK
DR7m7xn57SBHO0kUP3UDeRFOaVUvlAyiLxX+sQmD1LVeMPocUl1nL86O1ops06zcVx4izeGeOejm
hpFmFfdC9Ut6t8w/Q9COkaisX7EUJ320pcTFQ7bv0kz32gzEKqHoN7JuC74X/sh6fN8RmBOs1D+x
jCSub1sWJMnXFXObS+4ake538NVxxDbZYu94+v01yDPwnyxUo8ZMuFp7jxIum/m49wynq8aoTXQI
BpxZXGFuKfSMKORH0pyjRd6gfNsXJQicKA0aShkMyiV44WJQ0h9702u4NCsebokrmot2EU5WT8kn
gWqHmsvlAbUOuC3nXj2pQkACEeor/goW+cjnmkXqUcnxCrb3BkjOyQgywcooDoS8XdbbY6IojtgR
8AYcbLrDyuXelDQzNnZAS+cITb3ArPBVTTDhAbUwho2QaVWASrMHqQcAcflA6jqwRgsaLYg1pHPW
71T3GJU/y6Qf6/hq+CvwNpKRyirkCK3l03c16dv45N4/2LuAa3jvKiSjQnVhj6aOLmGOnHeo2Fp7
iv7hRn0pjp1OkrhMsAg2/eg4Xo+UXHSMFBMH6QU5SQeSxuqeNoXeTEWGS0xjBOJxXX4RlkD2avIO
BYfUeYa95KymSW9wu4StuLdCr84ANtiEAnE77TCyOs0dxsptXVVcTD2OUpKAjSBXUnnlgq3zyrMr
XP9jdZxrPHe28NAZcb+ogHgPZOsg7zNsNYVJ1V7lm1jgK98VzPjZDJ+pzhjMum/2O/NztrAoB8gb
9Bh7FjBfljjFqbGKI0L01Cd/Xg97/MqAAaZiMQ8FLa8IgSHGbR/RHeppCw4ZWDiM2UuBL6tTxsm3
KGAdTcj1ryFTY8UclWqSO1LrbAJZud1hvrzNjRz0IiXC+0VYV7VFCb8Yd7202ZF5xxNOYYGNTkUR
DUgmGSppn4oVxL8Zc6MFfemz0ufofR75xINewe5kmvwPWhKSeoaWIN0WHeObwYCMmu2WjwHJXV6m
YgcyxoXWTr6JxIdNx8LCdGC0KynVF0hheqBFqNg92EVdd389eF5ieWA9ZaWZQgwc4GYWSc6QQnns
QB2/3EZXIsGGxqI14s1GeTBensQzbp3PSNRZSMbnQgZe2x+1Ryq9lGZnU/9TeFocaxS9+OKyOsBE
KE7fY6JbLWNwsmGez66gBUuqs21J6aOmfaCpRf+yJytFX+QJD7TbJrlNsTRZrY2MDSKx4WuaVnk1
YTgZzyEf3mjGLJlgxGtmsYY6s7e+TtNIirJrkK3Qm1LYbqyC7RTQTkNVFTu+AM0AieY12vUTUt/5
DI81yhKBcJhJsdL/4gcSMIJv4MVlF/KanFFlQiKXLI/kFGfqsCN+fWiUfGi4KTE6AAgUx+vqfgt2
9sNnj9lUr8gY0HEWDtl43iUMGfHAgiZMx9E230gKwj+oAO1LtqUo0YG5pDN96wh/hVQNBZCun/dc
p+iv6Iu58RG7+gFdzWFWjz/jo4IFmzA4HwYE1W66DQ0QdoroiFLF5gCvQEm8nO+E/LMX3fLl97+o
6YSVtQV0/+MYV9S7WiBsuICmo4KXL+u8acp+5ZDh2PIwxGc3ebtEcOJM+BLkAI1uwsu+AFq4cYe5
mmLh9qdKu99jLR07SP3Gsg/NGwMG4CwP81KkuNqVYeAbimsmPvFjI9f3sppU/JZ1jrhxGOvcEomn
3asfEx53E4SIcXNrEIBy0Ziyi8t2D6Qi84sSp0pKxhP99PZkKGdq+QhKko16vqhd3Dy6SxIN+Udk
JcIRISDVke4wA1X/AoKJ8ba0s6FsNPENUfJ0lBc7zBUxiU3tvnkgQ9HZUYsfdGlOLADgdcRZ+xVk
MxnJOPshC9Rzs+jKicIl9zAev7f4rrQWpDwVHVvWD3dZSS/wNaA/XYPsmwnL4jpFRib+gkDbJ9JN
odcOKEOTaSn5kEj+SLHWbj6tOCwcFdrS0evah03lGg/aFqJLQIvUl0X6AFz07VIx9O858LKdS7hc
AoYvAbu2swrOi0EBluyWxHtfaJz+7WSeSer+dItNacNz5c+Wr4JLeHfUEq0V9aRE4M7rUvFhhmpX
3VVZrZGrTLCSqUA5aJD7rVCpFNTJxCysaX7S/VpntqWPz4NyFVVjaI9d2XssWdddYtrxDZsd+siG
rZwO1Ia+hSjHOxHxomXGrG66R6evo5cWRkmbFhmMcUMsYiCASYRutbTGcI9JhhDfoFYW4FaqQhe/
N6LZEBV5YbdS0GWRjN9ox0SIol4TmEkinceeTFGHrPO4TSjZq0lrltuMHAnTM70kLJoz1DBx2TSV
Hm1WsQkJw+RNMbZ5si8fw+nCgBrSut4J62TSbLSs5rGeb5jYvrBstp26fjjhuIPpYiMdw5f2uLR9
kb5oFjNztb5YJpRbmc0SethRjT2o0r3EY3iJslstLUgSVdeRAyS5Ie1qBqz8pDNahKSUM6qsQnvy
V3nwAbYMXflMzZpxIpFsNeny0YILRHrhKoarbyTVgHAvZtjb51UM+e/UUllmXj3pNo/5hWL1hX27
PPiWOJAe23KaNhuLARnwYML5eryi3JYNzntmga+wqTv2I/RahBePaOa89/WYWYgwgSX7giiX71io
whdg5G/rmILJxJ9ajdndmXzlal0miKzqY3KoCpPi04Ola47A9hkxFgbht9Yp4D8aQznlB+hYhv0+
olRwqvvWilAS9+pxAVG3fDz50bFh0CQBTlnd0w8HWfe2pno9HbYBBjq+resUmTEeUDYRM1XD8YUg
DTQkqmpun7ocOfNzOB1XLEFQ9VdgqQLHKHZLcQBgIwDv8+9sl7DXekUDcvla4u5U8TyyShReqnPa
C3aN2ite2IT1WR83lGgrSheWPcZnOkb8ZdfI4IQ8LsZU5zij/0+t2RGeZJjOJV98cWf9TN+DDi0Q
fEq+Und3acLWRse/4i7CRiUCn6YB25KUky1CGzYmGuCP6LSYimeeaZ6eEc/sA6/J3wRUl2T3/++N
LI30C3+XXCEQV9k2lY6VMgBIXEo36C593uLGUoW0n3ZCKKbotlAWhmUk/REGdanV6aWmBPMYByHt
haCOMdzFqlym4ouzvIZ7J/vKtMindLnOpM3UzXx9gvjqDn6X1bHFZZJR3f9UQQKrCTq4t2Gs4aY+
MJMDrfHAY6NL6nqeGXs9JNXNftkvm1Mn+OF1gWCet+kGTXim7ElQck3l/8LXnaqTy0mcYppFT+wY
DL6nk8P39Zn2MlT8unq5jlWOKyWoNyeV+oqifkoxOF3593yAxDh6gxOJCVyvzzVfG37hjAJAACgx
WkUVYinCWpPzoElA0HFhgaPYFVY+eEv10BLlpH3YFKjhxmoE2ww28t9RbTnZP/18HTNpEROHZQb5
2IX84GH/7/d6nta2iuIEF3lXDh1jyyIewSJ1pjvDHInRK5tWyn8=
`protect end_protected
