`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mrN+aHPwqESxkcnK8FrjncfmS30fhz+nVCjZviDRtCfUijIQ0b9bHuGiKvyA1+64lc9Xt0d5oIN8
ylrBkN8+DOKHyibe477U8m/lfxaWrGWUrVNTnvDIa423C4M49Zg0SMrGtoEyw9BaFc1nnC72Emnh
YPDl6EV11azFBhK/Xn7U2Fl7AdhGxRwP5Pk2UXv8x/6BL6gAtpS9nM9q63cpDDhqquFL2SeYpv1R
9LyKv7qxRE+X/AoEokMs874Je/81ghoPr6GtmQEJBPmy3/Eg1BTZOpJIC/4pUESl6waYu+HCP5Ar
Up/WSuGMdprA7ANf7om23jXBzKOXeZOTgdk5wg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="e/6uccpDube+uqyfXStoy04QjBWHBidltXIE1ttyAPE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 75616)
`protect data_block
r4gqLRzh5EnZXkW4vg6cQwibv+wvGonAglpa5Na5r0JGKJjbu/doNC9tjtc/WkoWzd60jKRHcQpj
Vd6z9AgZoUvGQ8OB63/3jsbDaYrpxDEZ8K6XfRJhutBZGg3+H3nt0WMfJ+lDdBlmbfLFJ0TMQAcL
Ddou6n1B3OILt2qHn39pfweQEudbOIZIO8UW7FAhlt4pPEbL3LVpcaF5HMStS1RbKl7wH2huGNlV
ZG2oVsbfMLgrswkUDpZlEo+22i9hmM0bWvKu1qqlaFO0dZv9Ey+OvdnEqAjlpgyPWnSJs/UWhWoQ
o2xhj1VM26wT3zXrMvQ3OWYYbyAmddTHOUuek0LZEK3Dp7zWRHe3jrzempd5KSlL6vCLhkPqiLxI
eI9ajwbsb03XpTjBNDuSX+asP/aBpiQR1Bk1iCIxR/dKnKhJ6Goq5oEouOmTjjkYUZ22IrByFx4A
K56Wx6gAOJCVmGP2ze5WI+4BhdDyoJTGnAUubbybnIwZm50IYcxTVG3+HUcFJJ0NznbZq+423aqU
qkJC90W8+6ipocLrKZFnQGgcVETrbO55P3tEyf5exhevVGVJKbE/hZUkpi7iHaZqpPpfwMOMav9W
d5MiOFIHh/P7XM7Rd1Y3SNCWdrkAAPqs6z5Od1lfPwzahVwkOI9CyZ5FmCUt19JiTE0NGO+kjmT/
+EXiRFfzYz5oGVQChp+sgmeHLsFMSkv7/iZwxfWC0WNpFypi1yiqnA/eFlLR7MPoPmiOr9hDVZd0
JzQa2tL/TfvReP6daKurQy6yWhh02uEf2lxPeKO+dkB/3BMe1FoGEmUVGUQy07AjheosP9Rg72OM
gQG8sQiBz4SALuYqYd1Gqf+h1sJ8tSBlID1Q3brwfwhL4H9f7F6Z69u8OpyHHtSRqeKmSdoYw5t5
hHUEdZHMqQ+bVvHFoNa3RD43MxRcBJmW7uSvCHf7PDcKgcOb7FcYP3ZA+II4qtu0jYHEBsOein2V
Be9qO0ko8UPVY6oLOhOzWZor4gXzJ+Ldf6NVwri/qz9nquK40NuLL9chOvgsLO5tR2+YdWL3U7NH
hMfIYR5spJyE1cYGl4cIiU5ineS7HSie/KDl+cEuYEWMKCjlrkAIv4H6pnRkAsmliPZ/ztKlwIYW
7bn6lPeNohxBc+iZMXyC7Pi6XO1wz6oit6/cKN9hVQVMpzU5wRsc5haYm65BuqPM8+xFdwvZlgHT
jwN0F1rzEzE0ts+wJtOp6+aCoi0ahHcAPQr1b+Y4QSRhZsD5dUNwhTeSZjiEYTGzJLVNywrwm5Nu
/p8wUhWOLNAige/HkpkLttYNtrMZSMmB9KZoavwQmJ48+0uBxvawLLc75UbbdGa56WUy1dgyLVBF
rTmVF817dZmC+F5EJ/StbfrG8JlPs+S7liTOJKAUrolVp30rALsQQ59XROtIs/YgtswZ80nMZixu
OLhA9kjxLBE77miSPfLQKsRE/K4tZrIC44OF79vMinfwU0pbWvjozW83uQGCJXIaSwHu13pwr4pF
rbGWnYv2bMMDDNYWjbLMJIbWk588Hl+6uMgr+LPkJswEwhfsQPKOfqQmylTkh3Gkz6U4JiSeE9M0
cSp2B3ubJ9YPpT3AQoivOYnvKGqNQ/ZLMVuxz11vhwM2cY7ahiJ1HlYGekeWWcQ3tktdLNPbjKj4
LU5qcM7SxgfrmHdjgRO55jAO4taAGJDrX6zP9yPHfGnuejDZHXLX2G0yUcBiJ14LKUhaXnQLnjnA
KWNewyqnU4ZsrfeGgtDIKNfoA9MlZS3KYOV7ija6XL/C0LX+hCJ5v5hFECs3cfStMJRL2pP6BlCD
kqLsDee58KzNicLGUcewVEqcuIeXHxmKfUN6Es5F7zDayGSj5MVinmudw9fo+0pEzxqLdIOIis6z
39bSrCS5WWWUwWH7ZIfXA2o14jbC7DdB79yZwk8VJMInoGLlofrWhgyzr3U4eEovWONUc8hy3I8l
kHs69Kici+CgwiFonJeyQ8L33GFuXNN6JqqXyl6QRa+G3niQ4kO5qbDS6WG+AZo6GdrWM8O+1VX6
AysELboil3Aa6V5xsTtQFyIue3MLNlUEgYfLAPtbml01MbynQyxoYjF0rSHJOJ5hU6dQq96RE7iU
D5H7npdlxu6aydMJ0IGuicWw4cxnrKj7BAB8hUNUApLL23QmVjkFmaF/Kb6wh5UBKZ/wdZrAKYPD
VRoS9VDnM6DWuJd0cf51l/rhIz5+tH47brRlhltGx9xcNQxtCs5o+u2rf5GQiF71Xkf5wHfBDu6v
+C/xAB9NLNKZp91S9hUwpEVRvJKC9EJJD2wPKFyX3nn/5BRY7WbIOpgEfiakusrJI/c2Bi9NO9Cw
StJRElwA3Vn1g8a2yFb+cgJ9JSej+SrFggfw5F4scAlKQLch1AqIf8MvQRkaV6q+fc+JOBrO72gI
qfG5lLmMhO+p0PboCN6a76zFeif3KPLwaLvDZQ6u5tgeURvt/QuOAvhoF7XszXBA0pG67+5WD9PJ
av6sPpXVddcRe6wLViA9NqDNqQX7E0qGRKsWiC6iIJ+OgIv6iUglUOxLK8d5bwDQD8T5Je8CUyib
T/8Eb5bNo5LCLZ7Avs/9iq1XJfCgRsztU5wOfPbdbUb2O16kv7kMcqd1T7eRdeiFfFRS+3p7ldm5
e5XN3iHGt583wAQS7hTizgpQxg4VwANJSMU681WNOWxnIQZmYa6xR2BSa2qn0dxm4TbTQDdtQJQr
dZupfNVxUFqxWKMQXXavEuZ+9Iv+skhJ5LSDw9HFKq3P70vrGQCVGq9WE1LuxyWhlNctylaOAr4o
F3KhoS7l3AjGQUUGGOkraZskBimq17Tngtv60reOe2dnZKBF1s8PMX4wxsc1z970XLRgc+3xtDMs
dykSw/vvvhm2VQPw2/thG/Cde6s4xz89gB0kfFJvVEwwJY4njZGQMjy3wPgEzt339Ve1PTe51sMH
MqSeWRuH+fOJaso1XYIYDgkpAbBRxnxEGc9jtJDr3A0GcNNnDmBDGvZkSO8dWn+TrEHP+MlJnQGM
Av6WRDAEPqE09NlRg0dl/VwQa1YjGYRFpKIb9VlzDH+9lLAGyWK7/s5tjPS8oMJi83wPPYkCB5wD
RfWh9QuyNqQoTq7FYMK20BH67mEsID7ROzQH+NSsQT8woVESo0LXnbAbg0uEsORUtas2q739ay49
VyaEuzLZqRkpngQtzni2ByZ6Efcir2TwgpCRCm8wzrdBHlCSPb58CnLYc0cpv10bhfJhAkiXrPDZ
ntFXJetZUXMwJEsDCCktqZjOlaMn3dzrsbbghXnnNVIuE4wQUVl8i5/1SLNs/xjk/PGWuNd2zhOc
sU60YB2MnT5Ov05uNsqDFyhJs2UPokcf1nL4IwIr5GJT6RH9BMaRme3A3u/QcsazSvMGt1vgwN7m
lqc3iPskgJh4ZuDTC6DvihrUyXDd5m/5vtsjKcYs80daNYrO+v5ZF1aJnB6M+21IeN1DLFEnV3u3
JS7mQMeqS3BNH6BuXtKI/ZUtkk8f6kdFFREoXLcM/fL7fuVNaYJ9BoaZsH49Q3S62+nm+9qgvwtm
LB9BvosJACPvF6R7LZ75+uHGMFemZuG9xWE5mkdB8FrqWzSZQ/J1pHquuoy98MfDpJqAvUld7B+v
p5LtUoIOsek7OtdZcv5oSzTSd76pfOw9Xrpnge2V2pHQdp0eYpRAYpxbBm0F2ND4F24FFC+3xyXG
i0hrOPz9k37HGoHMQbAkebNHNXV7e/4sAphfBvU7iW/wGFoeypetWVV8rjWielv7SfHJmxBGawm8
UYszc0CuBtk6n9G/MEYWdfBIuOreIi0lzTFngvaJHg2vvRfPg4d4nyRr+UOXHxdN2eoswh88fYkO
zsv/gP83Q2wrzUUAVAy2LUdsp5knhbwX1hSonZmgeuAPBbALZCaXyQQ5HI07MWnricbhkDwaekxM
Q7pswAJnPF6iEWFzD1+/W6+aIPrfJbxWq2K5fgqDvyK0nEewb9I774N7FUvjWbrWq9hpvWrWp5aU
WBdk+UadfYbjqtnVKRrmRWOiCc9TnWV5XpTEIQJtk3jmXrbnjnyukH7AaYEeKhx9rJnI/i4fUuc0
cQynca3J6PGKuspw6JpVCdLWJ9fUWH7ul5y0UJ3F+Jf5QOEU01mpCHd5kwmHmq4r/U8Otkq0GzAg
BAugiq9of55uOKJGapVKc6psTvyfW2vZxOq+VtU+96iJL/F7xllNL7nWPGALnKES5qMRx1lMdbw0
+6eKQzKVO1S3KIPpVzUd38dRoWSyj2reyQtd13Yupc8geZJPY3B+52fF9NwQNU17mt5C3XgzkV+Y
apT4x+m+Lke0pSKOsT5NTpOy/40/7OdbK2KxVlXHULmp/WVmYD9xhPKfS4pO1v8uRYX/5DdPJrWY
UI1l4FHDZrct+chtOCIO4XiQihTX4oPBpmNCQUWX/dNavm7ZE0YZPd9WM8JsGjse1WY8a4DyLudw
M8Ptr471P+2D+w56LEcWg0TzTcl3fULGYyNkueu1o88FfORCUObkG0Z2q4aZEPNVaMiy3asI0vWa
BDpLXSsmbJkau6V+q3edE5HraZbNBaH8Ntf00XEkeMX22x0/uPwAGOFxtzkz70VOQJwqY3+/LkIy
CUQzt0SHOHWdSd/UikoXG+OtMYs0Thu6xQV2Wo3HwCXkH2esL/rR0m1KMQfgleaLckND/wz1hV8b
p3vXwC0jQ2E5dld1zgVdLdTfqpOsO0Bvg3J5+UtfnarxNsc9Sh1qtpi5dIyIxNaSO85X01sPFVEv
MQVB8+zrgKqDHxXDyDEKGrpdsHzwwojq0u2UXakrH60XvnHP3hzgrinQSj+3H9FIYP7k8cme1evf
I6sIk9TTkTKGffzN3cZLmmtTN2ANFTtmkBLKrnBM1iYPI+GsKWZZfzxnBvai3K8EMocxVX2a9z2f
y7TOoz3AqQjz1KxfHlG6tV9TzFkwmwl4klDSJ5SvubQ3sEoU5X68wIcoGZW85hrOIPXhrid5kWdj
JzoN/x0jO6o/TAKoqgriOmycO+N4aB+vhqRX6hwJggYPrjHFlyvAQhDa8aiKymbgwLVcJg17wWlk
VIwDNGm42RIufQnNAJC8Lj5gYxh9sB123DTPR9QNh+PnNoGl5ODg6S6o+VOsXrIE51b/2Fmhuwm6
enLWGJvC4stwOi94a0x3ek1OuelFVRxMjvP0A3btZtmW9a412irzA9tC71t98W9WY1g9hJg9cv/Z
gyB7wBu7l8yTEE+mCRVci7PUmDIe9DDd8DcOVP7tU82GCuovKZzJ/5jBYTwjZ1+woCSrghS3ZO3s
AL3Ia8OhzTt43ARUgZFrB+Yojftc7W7j/RR1s2G2xzhFsakjN7CCEnnrR4nhycQItLvOR2lOBq7v
xVEw1YclCYePltHxAQX8tIlWdYBpZWJK7uyLjH1EssXGrfK2obuRmzdQb7sIbp/T+n6GNtdbAVWc
AOGxaAG1dVf2dJXpP+2hKEAnONyWXfkaMhT53Et2GcQB7JP+03c/2ARdeCfqj4rC5F6wxBfO9lVe
QTABPmsr0y4b75foCKTnAoCWjEqPwxiv407VUolRZ47STheDcpG8AJTrxYXT6AgV9ZBlS+sabPAD
/9IRN3Hy3l2Q6G06rbkPn4wQUw+QMRIuSODnlAgitcGSYpz2IhqSImzYUoykqrMCkTRG8jc30+d3
H2+B5dVVXingkyduLIErgIEzNeWdSehNWGaxNMRQnvqoKY74uflIiifmu9r5DFlK3MTewi17qIqz
+yK5xcnkI+K0durD+Vh6oEzxVISQq3jmBJFvEXLcqRk9TrzzI05em7sSVUto5BAgTHssn2G2IFIo
ZCAFR4tLYCibMwSjmeJ/Rvt9sfqcnWF+EDnCEVEu4fb0weCxVAYbRcZNIgw8Lw8qd43wXUkcJrAx
Z7LR9JJdYnPyvETg009ybvqeFXpdGmiDbqb0dNUtq17blayZ0P6ZpoMp82ac3ygNHdKcAc8bZktF
VT5WOqi3tCWp2H4LGgjlGX3w+PQhM75fYoQUnTSBY2jFV4MczkucoSHynMABYt2X/09KQ8CBjnKG
Mvga3h9mF0H6VyopPnJKzwdOrut6qHaJgiqGtmaxNcJZyXXF7ps17pDut1etEdRy1OEb5IhpU5Jq
A5GCh0FSD5qi9ZkWINn7apfWlmBLYeRkrGWu59xpUWOJC9qCQTQtdZVTn65q4z4CvcQZMZ/QEmuB
xa5tzwOOoiEMhHj8n+CG/ZqkGAlMkkFKsygIgG3hRKa3AxOwrD3ZIxJPRJTR4mEZ9oxs3e2DovYt
db+YmtTpaMnf40o+LQ5SVpyJjseGmhERur68hm4nlnmiQDsxiebzl4OMEmsprzXBoRHSjZOnp1/I
uH21EovoF4/iToZ+Oj+3GsUN/oxfJ62vjoz5WRtRlP5cnVM60xmEActOUnrIA5FFWXBaGF6/ZdGU
fQYM3/QlKR93L1QFIHYddH2D+1DyTnObQHaRbpzc4rzlIrDubr25g0dGOxpmX341cxOB2wBH0hI6
qkf9hD+U+iIBc2wExc8K+NKmfL33uWg9wLL6MNEBgtklUrBenKCMyO4RDkhgQfxd9oF2D6gaX7K9
4kXC51T0tDr2m7LEEnwwOijbFQY1zsLO9M1p0WdKZ6y4b9CySiPtR5BWEuLBU8oxITJhtVleVKF3
atMrede336Cts04n3jv9sbR6ObkiyZ1/nAjiF9a5NyP+8kwMRNzk/k/vqKzCFVD5S0wtVt2YJJj1
w/wbspmYxYmyBRpny6yhGF6PiEi72oOAJPl+OLcru5AJSfEbN62eepLg6cuEqBM7gZg/1NGequrI
FM5tc0baTv+9HfkzVKiaBQa+XI5Vrm+K5OFME/NlAY696JRI5bfHPtvLh4p3uqeLlc64fPeVFwxC
j9QEpg4o0WDXPXdEuaeO8FZYu64E5OeLbd2h3M5Y5E7kaA9Zv0iB62pIRa0dXRTmL7cb8GZMEaxu
k05iVFLBxRKYbwMjcN51bppQuYg9Dd+hoWitdnLWb2KUiXe7zfUpeCj3RtyeXqru3SZTIchhYLJL
6wv4M0gt+jHVs7JG+T/g+38MOx5znUfOu2UkiBvEPxCUKsA7toIuQ95Hf1rmo6ScEYEkeamLpZ75
Zz92Y1lyoyZ6t63uCUezqa5xJZljlCltrMbdDEnrWCIIJOAsAnFdJAOi3baUgOOhCxlrtDlLlkM5
ZQC1MTY9QaOg4Asfv+GpLMq8iPMea5TaAVayixxYL03+MV/0xc2CknKUajRzDxAJyFx6w+oCrIDd
/gcxKNdZSlHuhc9MwGyZrbJWlgE3lC7+psDDk1s/38biRJATkaNS3IKADIQ2z3IJBTW+ZVA3C10q
tYG1q5Vc0kM+E2LKxYo/uRNOOUQG0lkhRxp+01avNJ5E81viWtOVKf0OATCGPoFJviLAdM6W5mxe
w41y3XBlyoG2qswVyv5zh59fSZ+0M+YKFW96mZ7MFC/ts5zQsuLRCdkmX1zkOUNpJqRqBv3tzrhV
O8Wem4UibUMn0fhOufrziA4nRx7nLNr9ABQXvyHFVh8RuHv4kRWuYWTveUVOfUiGqR+8bqH1Tvqb
DglCJglL7RYtm6AWnMvIOEEk9LZfMBt/V2uc77JSrI3vq99sc9o8mUYELDT/MPb+Cj/uk7CsTFrk
sF7PokDRHrN7wbSH25qYHLH1D0umJX2L1iul/5ROSxpGgJdUKQQp11nChpTPhmURosYSnt65i8RN
Yamikhe6E7l/dT/IVndnDz4mHJkg8DZfbmsSLabBkluK3+KIjjLVYMrMKjLWnfjpFceafEXl0pCG
iBxtbSMcrqS5HCAxpoNyxFJEytGzd/ZNW+pON+qOcFRkY+QYsxJyPmIeVXOu6Ro2Uh/cTl2a4FCK
XK9wQjuCNTJlvSWoojilB9J7rqgso5UcC0NZqxCYmdvE8bQZkNSv09q9e3+ERvIp/Rnl6VHE6TVq
uUx01lpXv5zrKnQDveZJwPoz/tfWUtOrZge1Yy+0NL4m1CGvv0F/iscj4bU3J9LorFYWib+VaBGH
DdW8li36S5wSXSf2S/IEDSEXYOTqTOb9Gaasb/UdiQD91WW5r9kuebh95yt4TMAaLwXpMEfi9d+q
ZLaLL19awd1mRnIyZA72pSA1yEFXioMLLzgJYLgWIbcCn8DnbypImV5kU0UWt3dLoIan8NSyRSpp
f+9fFz7SmLEUmkJMm4lxYQJRbDhYWppdJevvtBM0izGdFS+X0JNGNH+093Z6Vfv50TrD8bj0204I
V3zz2tfDaDJXlHDiW4o67YMlp5doTpTduz0kXzgRBKGiMgE9tZFGJG/mN+dPRz22dCXBd1Gdbbyr
gktdiZMFNGZskLVmSnG/BULihx6sOdOFhU4koPcsLMIZ8QISrPvLstgOi7wSNhQz/8R7vLRKFJfo
PwiOo7r6M3Lq2EsV+JjBesZQKdr9h2eh9JhSZuhnLco8Agdy7yPFjYtWpRqn3dMoXZXfsn7tUf4y
sCfqSbStf1rLgGnI2k6z2BUt61Fan/5/BvTQedVTVLozBic2QpKTR/InzStr3zMNQGTegpmUpZSZ
AaP163Ukj+6Evldmq2eeVEqSMhFivqBBH5/TiJycbjtVI97WifuEvJwR4mbhHOC9NzBF1nTWQSab
DUfF8Z9lvD5cUhH+On/AuVfk405jcda78lmIkmc99IoyEKwZet2EQbE5ZUZbFINgTfstqnxJoEN7
Qetwwqk40J9AqDiZCt+iGT0k1WmerYJgh2iK+lyignyg7OQxEnZx8nYyge4ImhjJdyfrhH0R2nsG
DInsEo/AcB3HzLXn9z1QyMp4h58mV6CFBtcj1EkToY6SQfyl/dKy6Yykit0fHS3xwRCCZNjxmy/6
PEct+Zp1PZkaGnRioqE3RbhDYXvzHYpzpsAyDYA+1zYxGnT63ERqyfb82t9pItrsi8pavEkEiqLu
6qpFHkzCkvg5cYgOfU8gkI9p09SmdtuPVMQ8qlDQR/kfM20ktR2wHMxd2f2R4Uig8P5DTJFGABrE
7SJWXcRVTHsyjmH4YUeZoY0MzM3vrSwXTcN9barKvB/s0xksJxo0gifn5cftQbZb74InyPXAg2lB
UguKxRnkDtSkVLN21FNBa0uDSg1t8HW+sJdUQHRAlEo7OgmP/8KTz06bt7yjy84JrcbdPdklFhce
cXuwcr2tB+qKMGOs1ytRVk+cgFeoJHlhh5p3oUxS+Z27qpYAUHklg1hi0+DUPKzhDKXaHqf4ItVQ
4Bb3fhOEmbv+cGgxLKjgxeZ7lNEOMGz0WyuP2Ip4RdK5ION8nr0/dHBgjQlW5UOqtt8Sk7K5Stot
xyUS4+SPq7Ij9Dc/iT1AfN88vmH55RMJtWKPqrnmDzeC8jg4ng3GclUUXVXtZ4XGULmgLS7a+kj7
+D4+5esmjnIpMgWQ5H1nQMPmHSGPBS8LdHxyNg378vnTu1NmyvtcuRiIJmDsDgeSCBKyX0pWASph
zZd47nH947KRMNlH+xC0KqeNIZkbyY63WNBpyd1LYm2X1fdKEWVDG75RBH4KFLi/mjcC4y0U9+R+
UzB0w+ogRgACZ6bXt0sqjxPfDjEB/4DFO2n9gfTO83OUv4GCbHpWB6eDEqnVu2iFRLYKdQE6ipcs
bR3YAxaiChvzC24OgtLOepgRESoflIEvVL+vHcHlTbgVO7lpbgmYL5B4oOjH2BqGVhuTiVyhl0px
ZyejF6yb9GoXHwOCFBIlyscCTVInxgVPDjNKjFS2bugsakhDd0WlsowWPLAaGzH3r5Zol3Jgl+Ew
MIzBdLSLMELgaCqPiS21WOaaueoqUnDWMqZSEI5/Xh1kV1fC71mJ0HmQuLmoEoLqT/Tq2Mniby4q
VWsIXIgs3Icrs977M7suy22k1koq3aWKpa2Owg4QZ5PQ7btbb95bai7yfD+HXVqRlQfnXWtoS2dN
D+YdkBN24/EUnlhVuQKR6ZBVp2C/0KNiGwgpHr8Av5rLdahgSUTRvWCp044ynyZ4102RvCxN/vmv
7er2AvEKINElbze5MEvQvrrrGfGXduQfQGz/aj9Z4ZUXzdxX4nlCvHf/wnH76L0UV5sfT9iFnvC6
aSXtDjj4pJUXkDdFcoS8sI4lNYvIkGswB33KUJOWEvdXeDuclJX+hxRCKrSzIwvtCYrruPTn5qQq
Jjn/vNNZtUMtpJfy1PBMUVjTp7ufiTr2D9HB+tBd46z06+fqgLDmjr4Y7WaBucDM2FzF4BOjdWlL
7ZgLg9BgoTOBF1+i2d4eaabJbJ+KZ4ORHmAbq1mccaaDOMOM0Wv/e8SLVm0xZaRLH7OETznDi0tU
wdm3Lubi4380pTjEeBN+ZeLQMkHlnHRWLLYVeiYVDku8yc7zVDEzGfIikEYwHRd7Eb1M4LaZLP7q
BqfaNuypYy3figo3yUgSQRdlEoBlQ/CfzLE6+wRcaBIUS+goDamOwIGh5U+6CMkTE+xteqzyvdgL
U+9qCbcBIn+AXrVeeNOQ4J2pTdRApFzFBn6S+4rICS5MdIQEOggP7cuRgLlScjSb6LK3FCnVzhM+
ICWqqf7tutk82C6RCcuWI9U+52L9pdE7JnNpJMrJkEfKadO1yClNDnj1EfqQNd4TcUPAyHITbawJ
d5YumSNCzAdl/39J70S/OqxN7qLi8lXxob35Aa8eb0d827iRVmJyADwCu00rrYbrG3MOuoRihRD9
Bw70Lpgb31Q4JdGFezpIYONvkn6Gcp3qk5/dVPrM2vAWMhJ6k4ErlWycyEGIzKfdbQcx64/wkxdp
RylkjYpS4N/9yTxRvnRX2GTbslOu1hJ/2Za/gLnxXy0zZhCY+doS5oVtnvbKrnG1YqrjpcJWsk/P
pE+sxEvSGQWUNULZXDwe+FPcsYlPxTACPwFVfphKi43hjcBZakO+J0XW4S+FzJvPoNgCs3gdEZ4S
FXXShLjNMCDBaOO0MTn7EDy1njU9CTeiM892ODXHGZzknUgZM9L5PsTHJun6ywWiufESmAaek+7A
scRxrpYmqgKtz3ia5k806dKQjD+kBiYSWP3RS/hhjNN/BrjqWOlvtNAkP/zZaQe6aAGsx9zqCX9t
nT2uHfQym8wMXUgBMXExOwePRZa8LzFcwJBPKvLFVmI5Q6GfZvc3CQGBdx5K8olyPW6vpooZ4X1S
2OxObvWslCLY6lVvMAA1YFUx+jzN5fHVVsdbwKhVUX+YAGVcxKveZosysUu0xKgunQpDkNBm73dA
M3ELhPFvawC9axC8mclKm9EyXHEIPL88To/1865Hozr/zdr9qidmPtEKC3kIXFp/0f4S0O4D5Roq
BKV6tp6azF2dUldPiY1FKZ10WoAzi132PCI8IuCV3ar7Odelq35wcyJ0M0BOx8nBeKBm9anWw7PU
Y/FWFF4A/sZCRqLQB20rm2RFKmwMxoYeodlf3OczEkdBVXR+tl2axs+JiglKAJxzutBlDacEbg78
R7h3Zm3g1HnX4Lgpw8tMkt9bJ21kivIgR2+LC2L3SPyiOPhkLqZjBHLS4s9k2vQw62SOnthmFuJk
eLXxJlr4mYqvyFjU0kDsUNOCxS3wM/p8HGtRqA900CFmq2hSwIywnFK4SIgJUrpWdsYvKbNajQZc
RHKyooUwUyMC2d4BjNrOWsQfEbTTsbUH/fzwL7XJtSNAQoJJ7EULcBqnzHUmo3aNobsns5TKr82f
mnYIV9J4dWI3OfypCXqNV+QCUVuDlY+TIZApVwBXDnIlFii76DIZInZA8KShgEwXEuga0W/pv9TO
cSa5KzdeEQ4KilWRDJEeDdxEc39s62Bb26yhGHnnzVMBPi/U5oaxQeGLltIAlERIaIZ89LlsWELG
llZwfmWQSVJKWXDo7cp9Cxffq5NS03rZ/9HUp+aJ2IU8Vm0kBsi9ubwZVRSWJBZQqqgtSGug8Oqg
ZTEEJsrSHJxRRd56VCnX56lF0Ybj62Zjv6/x2NzC7UrpZPavYuOjnal9neDqaGmYF2EYmdB245Wu
AKqjTVl1/cMYq5MElY5BB5fuuCKFvb6l95ShGO0oRqZj/tjbTO//4THzTxW+ijl8oyj7c/xDm9z+
as2kDM5D+FhdU0CB5Fd+zCRV5A1dgHfjSoiSAfn9Duhz1CuSFVa8ct2snE545G5kOQsAlxaa5wTI
q/yopyMuAPcRvjBBw64hW4LDnSyI39CyFLPnv5LVpqfvi/tlsQP7mbLHy0OS85waT/aHmT3uIb8A
GeP/OIZ+tOjwlT73L6lQihOLZX8X9NC3BTgbBTuctUe1GTUVSV4it7A8pqCtzFE7cH/eMzJVTq0U
24XLaJDgdB+ML+icMK0cLIkyDR0KW8OZNrTYgxbeshdTx1sBJOjqqwd/fXDHYKLqRVYkYBYpDSbn
ebi4O8TXaYYHbTq+Dk+7sYZaqOXcdH6mkuK7adKhNrvzRZ6fVudxGYXtz5E6kULjC4GWkDTf6A2l
H5RAqYAkHu0gsafCT1o/NyXZ6KTX9hRi05y4DyBHhkv9mLg+/N0RGVQOv8dMbQe4y3Szk8ELDt+K
8iebiuiip8uNlAIW3u/NQMdXqgue2MnVOd6vgGJSrJRgucEK8eto0hoGMPJKapToNlLiOroe2bDH
tYzeWUL6jibuQOSf3mbiS5R0SFCAuibOUrQVKYFl1W5kqYKnNHbMQGlu3jdbPR0/0l7ha26m43dc
wkSC2zM5vhbZDCfg6AmHEmaWE4cyGfqHe2VMdRN8ZiIgaFgLp7Da12Iy0yIRQDkC5EXtuw6Ryyr3
jwe6JFoDWncdFQKEcc1a7NzjQf8XRQunb22ClsoQ1xVKGAcsGzlQnpD8K2b99wPVeSlWPvzV1u+S
/4uH4mTG/MxDJ+KPi7d0/ZHTEfkrB+UxJyt1VQiYx04TnKY9bh73JxPOG18MeimWUA5QGtFYotV8
MQ3JZ5MJbXA1uuXPbkYelsWMunsgfkcFQ68mzsAx0kqBKOIGpd6L6LplGN7EX2mOrzjjY5Bet9LJ
bSRV5fzLmc3cHJBU564wbggf0dHblnyJtoJP2gfQjZRWrG+BGXK5GpaS6U/xr86P75ctDl42svSc
Jthx0MFVy0WJR0EIrEHpGmVB94y9ytbBLf/z3Mm5qp9CULIVDg8Fefl5THTnOyNHdCwridV/dsTI
fNdKMvu/X5gPBPTZlzU13t+piJRKOe/P30Rqup4j6eihNbWmb6FmfmA6jm+XrKy23O/GVrLumEaz
PF5MJM2lc17pf7QuuVK4PH3CvQ5bZa5bwZrLIOxMo86EblOfz0HljeUKmtVCybqZyVUxz7B1bQ1W
vbES+ZV4ckmAEYtDNaSEU37GARmtOWcoDPLlAJMFnVOVNZSAPgBMemqHcN/IiHpsN7xq2bLWkKP+
/tXaeF7TbQuNS7pTLUSBQeT9iXYNyDWo+nid6M7/MCJbno9RRA6RQ5NE+bgf1IFhataARtkaodwq
ZiS60rEDNcEDXsMCO/HKkbocCYTHnbvJR+NiEb0XxmnZvHBVqZQRdjqx8e3XV3rEMrYdT8ba/PEv
8U/Xqza3uqJUYjzIhz5BzzC5DKZuchhi4y2DwbO6hgQ1GHSxpaLV0AJ9AWOvkSVsrwH1EL90wM87
4PB0NncvNuOrmIr3W3/uFrd2qIAvGwMzoj7e8XvU9haWRKQ2on0mSQx/UYcw5HY42Wd65FOpeNOW
wwi2Z3OSArSONVdV51dhSrY4UN92lH+M6nqr6CuL9yJigcHAk5F+ddUOvu1HGXlD4DTh8fT57IQ7
vMOnyg+KUquZkE9vGsALpEyIX9EA7j4MbvzM4xDp0CG01zeUNApsJ4b2mLQsjhZwHctCYpKr86bT
I9otHIFoQ7OkyTG7xNUSJEZvzWgszzMrfpTmC2brKEipLgTcEKiSFM2o9WX4LEhWSpb/YNyaW3Sp
GN7UURPRTn8aeuX3Y839yx6+nDQYSXSWx0AQwjOCzg4gvCcb2AjLeARHZiBdH97WD1hFAsaY3Bk8
0iyfIapRnntVw+Cj04LjaFKBkdnzK4yJLJhu2orwWlvs+FHU55T4oIgZaX7fZ6w+s1aQj3/P+Gbt
MsIpmFb9A+EUptmzQ4zHTMBXbIBoqH5Ub5J5+Pxj0xPzj7W8OzH1XwYeJQbfx0nDIqAco3ORv8nu
jkGrVxfiy3r6cxuyqApmWIBd/PzZWaZy/dYTjyYQuoNwA7nWGu2Muzv5voYkA2QqoGNfptfSsIyw
2/XjXkkMpWUvbpN/zEowrkJz2AS+StG7vsqO67/OROGwzp2l+pr56jO/brm+CmWLstcW1RmZ7mNo
0Zxh9JpWgPLT6zr0EeQlJccscJfoTHTLN+4qf3FkKsusdM5QY3pyY5wLtSNDF+ceP2ibZH28btu4
K98oNZFTN6Ty3HSdNOiyqlXSBAvZg0K9E3syJSFErWxsbg91CopbAbjGVBKyenIcZnXT9ElVRoEu
tGO2H0KtlmtLDX0ObKOszUMxKNxCSVI65jWdYhbD8F3w+Vt6r4BuxZfa5ySZTZQLvABgPlsxm10I
rQPRH+eHoYpB5FGrMb2DlGaA7Z2YNwU9EwyUuQgbugNH3oQJSvFtQ/Ukzu231gKjyJsoi6Q4Vwp8
pJoU7f8s7w0Yh+Ie0dciYdxjkh0mAsZd/c4giahn4HIbyJGBEsz0LTaUKy4ai65jHEjE3I/4Dnlc
Z0C3mFXFzKtiJOO2AqqDNIWlRK97IxKPh4WRE2TKWx2NV86Ufa5LfLuABXgPQ1CWICWHvrYOcYOC
bIaHJqXxyIK1RNca2RYnuB08xSL2g4Tw417QmeHl5UDlSsDn4uhCph5ym2Jw3ueCp9BJ7Us+zWyp
cBqfE+ONIDpNIXecJb2TE3/4YfitRqCAHsrL5c4sfu/SWomipJdPvdWc54uBYmdXbJm1zbwygjFE
K+XVCUZVg67FgypucM0dZTlIzAA99KbIFHKQG3269c+aieDtweTF8nR+dgoxAPIJJNGWKa2xXkvn
TZYUvfOiiowHlhExEyILcMRoS+jOfkYt3T+2p2IFfB42EvRn6kH1lI9TmZHXSi/wnaszTb9GOknv
ccpYizaijYYEM4toahPVy0spcjc2wGnnxB/dkHdqUSy1qZ2DUnvWZZuDBdW8p4OcWuKYbTlw0+Xk
QeuMC+1k3lL5qJJqDJ9qXvuWU4hgbsGHoBW0aGAjOzMHtUvBgZMvNlvEi+LfnDCCKSkSDRr7zI3Q
xyDxk1Osp4XaTwl+0ujF8uT/Kvlt3kX0MCOmaQNo+rKkvfqzUw9e9oVyrnMuB+G95pVsh1tskD54
KpkchghOY4Ur7q9lMaLCvhCtN9FRvMed/IZN8xcBB7Zl0/rFSxUImeieSwCwseWsswSOOar+8I1w
Yy2OIvgLAhlYzrd6nOKzgP6InaMtystoCpFWDiLkQBLEdAoKld8QfwEnqroxuAMoyGWTalCLBQDG
5jYu1kU615I+c1LJpZiMW6146lKMTXoOvrgcmhI853wbJhlPv+X1ZfD6bRSo5Pr6WXOEeVjf6KLj
tL3JRqJAcrVsmAjJlXwx3eYHvJ1gTpBBve+Y3PYytbcHGZdH+R2xBvnO5YCcduhDLzm5e+gd+BAp
FfGD+kFzGV9zH25vF/Db7eTFtfCdW0/zTY90dRX2gicubyCQPBtXJZ83FIbkq7b66RnPoJAuHPQD
WINvgynmpcoLURCRf4lrPo9kFYeZxdsrk6B/IXRtrvrFMIPeyrVOlpPuhn/tTR3WcU7/4b4FuRNo
EuJPRl0xbf6+E+vZwEM7VMOjwJSulwDaK2q6nrOsMq2oXyRduuTyFgurdo10G4WbJWJl767iQQvg
LSNvRv+aPBvyEPueJq3kDc15bWf7uMjuf8/F9BSLaRGh9P8KMCOoa4g/lcfSQqVCW1v/vMgLcswm
HvRejaSsoXJrycvEG+UvqPpsluUkE9PJyo1PrIHydYqVeHmeeZU9fhUVoJa2yxmCbkQ/SC7N2Lw9
msypOUmNE9BSUjsG/rVdmn81Ne9tQq4SWZ0BRNp3GR+meV8ydNMyPZbKUjCDFd26J1viiqdCYBHG
or1M/fa93OD33JQsbrYoNPXfEIX0By1v0NpYeKr9eRGIq28xv/Mj5tjFjrfs+B58BjKo8gYDxKrD
biAg43GTHYQRif7gPniO3aoYIPUn05f5jExJ8upnnor6e9zcRdAOXpsCTaq3/mQlXUkr7CAYkDQI
Y17Prwv+CLCGUIPPdWtn6sbW1qFUj6BvzDnvGmSkunajNx+EVzUufVCuigsBGADZrct/XA8xIY9F
1RpRqWMcXLHvk0uEF2HRIz/7a7ItUUF7YVlsBZkn3PlouGbTZ3fdfCu4kJgoYikpMRQS+aSL6zWN
curiU8R74GgI774BTaubodvrf6qijPQGv4qqt31yhGQ4mAaSGJKnFwkVVnBfwtM3FbvpluzG94KS
OKqQQGrIm1AZe7w3o2VqXJv/XpkG5yXxqqIVoqOSMhFKjQK4iq2k4aCevd03RQuIhya+XE1Q3uqm
8YmcSJ6/fHmpsCIUWZMJTUZQAmk3A5GWRL6MwpW/aTluU0NAMGL0KY9QzJreAibOT6rrwUHHU+eC
zlVgL+gjxs3YevNsGyM/I6Gv6WnS9LIJ6AF2NetXq7ri09aKuz3DlvXhGQ+c/yACOVoe4yt9m+5v
LMbxqKVP1pTyRgtOCquL+vvHVQbEyWAuTkp5q4A4GVrkPk3BevVOIbIqFMMCWAVTOKP9KxmU31cA
tHSu9yXHWniq0SGyMl8YzXmpuX7J75yTHsbDZR9xweofamkIKJHl1xrU9S9GKNpOHrUwVMOEqbTi
hEINY8m1o3hAo3FPRsmHcHS9vq9KWF+XN5vOUGnP9X5C1mguUbypoVDZSirhECJI1ViAkD7n7qYP
YxXDT1lHYi0FkmtWegZ+f1elDHNeMPL1zkS4k1KQVA+YDIvrj5VKOUR4Lr/hxXM3ZFb3r0954yYh
KUrBynOB5xPniEqdm8lKUKkAscQTCL4XPeUy8SKPAI86dgbU5NGWBLQT3TO0VOgRT77zCdWo+d4k
MfgmfE+cJil/WQRtM3mu8cIveUzvWgiZ5hqvi07sqtxhnjJlpriEs08ozxSYFsR8vuUZ2UJ1Yk/D
zjUV7TNOsvK+ghMwVC2UHHm3L37gRMAFRWKDoEshpBDiSEaVA+I9Raju4M7LSFOlEM0j+BFZgOPh
0v9Fifgo167sanOkUn8yBEs70kCa+c00EsYSYkDfphUa13WcGlgpPy17qIj9Yq98PzpnmTo+hqyt
7ttdVeGxbWyBk1jGW0vZSzgQmnc8aZf2W+rn30kxCTsmc9zMSsdGzDTAYOJEU17s1/hJhTGRQSjk
sHrlVlcHgdJpRUcRQpNAgnYpki/+04f2uNBN7RAm0ckV8SnfBNpG9oAYe7KM7j9BzCjA9I8Zv52N
TIFqydM0cqvLg4eDIZqdB96/9zdH4JHn1slw2N/GicuPmgLt3m3rfkXddeLVea4btdQlZQ1gXoVf
1C+r5c2JS0/FYeyjkvqLW5RHtSCv0pvg9QFuiA9wNYElxUDM0mF+wNKmzH0PnEbciK67ifWTF75W
Et4JyHTP5/7OmI3tE/uNPL0vzo4LrL4ihsmBXyp/N0tuvKMDrnHNYbyOG3MA/+Qq0EHP1f5sBAMM
378iUVjRQfb3WPtdbeoT6tVbf1VFh02edehkGsOk5lCG46u5igVe20WMcVNCbwlJQkvJK78Hwi0c
bOO/v2MIzM4dJWwf5kFjCbw1P6pf8v5TXI4uZFSF93tljJZ7iA5BVgMP2MfXHewu5FbejNfspQ9A
FCjlssVQdIvZBYZlZWIBvUDRi5l1tWAR599rfWIjMro5AA5cP0tx82DqJp1V/HAQTlQGg4hhJKm8
aoykQ09wA8kUYebRM8l0XOOwpCIs1Z/psFYqqS+jCwdxtZDUy6chb6u1nm4L6Cgzru0n/8YG8xhl
Kcv2k08+XBRpVZEJuMIPSKBTSR4B/sF4+iostNcmVckdkV7ASrtJzu7Bc+wXwHM0hEeL7l9fPS5C
7pt9XhqQmif7VhXG6Ye2gJHFqasMPIBR4JMItxNhMu65THtEyELSfu65PcxBNf+zRNlkKFu5FEJJ
ypYF3GiWnKZABm1IZFDC5obN3/tDZghDUG45OkHfM3eCZXFndxGEKGVc87Vtm76M4CRkq2l2ne/Q
xeYPshNRk6Div8xR959NoTh6JsS61G73elqlwCtaka7koIizdi0dqLK9EqyJpxHVMDaclyueslCv
+LjtdgjA+3ioTTUkY0vFk2EgODYULp2ZubJnWDHBF/qlAxUxRWoGfUOfCXhhNLubLMyi0y7aG+Aa
Urj+3RqNdzLC6dYpun3dT1L7HdKbVQ12xdyoLj401nWuC2bu/35snc6xjNmqmsF6orLPy4s0v1Ma
yfp3T+waBjEQEaiasjqUNx5k0ts+B/xvIxchaAn/czIntGvkludthPVEUYQ8sH4y14eS6/6OV026
VJOgdb7fAR9vQOvhnjqdJq+BBtMVCdMSlnZ5BYNMKAC7voUi3JxwoFiHYsu5Zrpc6Z5NsN9PIHGG
0KnDylG5N3FSoj0hDZJxTlDdBgJMigxJp724pjDIBZm+uKjevR9P0ziyuupg6v0jOoO+YXoe9IiZ
S+7gC0PKKxXlIJwMlNfhROMwjDOUkgBmjN3bi3nDgnSc9hMUkGWC6ioXjk4vBFynn7uyQvP3H/hR
nkKqcca00qW7nzdOxY26DB3cHeOyDdCtm519chpRX6s51Zt3inWTI9xRHadV6nIEx3Y82vwqJ+bU
8BNPBrj+l/z3CIw8xpYwzdpIIF8NdjmVXzkkNRjHjUUubNzkHjpjw4zpEZ8szPgbuNdCQqKINDq1
Hz1KJvbqinWC1ktuHq3t1XDc2W42dIiX7NIQnVskgAcuzMB80qzCV2+fDI0YdM/e+vXTWdGQHGTL
4CJL9E8o32oPcnF6eAS9DqSgopEF8woWUD2S393sPhHTMS3uFUEABAZFTcdY5L51oQeHJXxwev9Z
ovFnnhFu1l22Ph/I5VncZJ2qnPMco4gY4niiegZmctUr2iOSkMda989e7UiCSTzxrDk1oDoHz7y9
5Ks9cgsWM2alx02NA8vEsE7s6LHdDZzbC5N+yZI4loZNYAcr0AKblZpKEKKmVq0nwWGhGCh0JI3n
H/jwtbBHDwol45vqNADalQI6Do4ARmkjDPL0vpMNl4RTzKEszgmIRxmxd1yqLx1NSwDiqxvdeMdh
Bmw6vrLJVQ/phKpqcqlcW04yGL16bA93tBUXF60fN/9L9AmtttHcb5ostboFSn4fKxIDFPXldr2b
ety1Ht8cUuGwVWiKXgpiIDL8NZ/W/uSke1s9sKQEtKlzqge4wzXnceioBy25ka4gGQpmWSLY7xOD
qBq9xT7idBQjVWAJ/g+LDzYm2+WApafnqKOprYIQP1aaeFbbcEU4HNzMJk3xtVwQGRINfF4o06zZ
jq79HZj0eH1r2/F7cmEUHINyHuUfMWTIyyUsPztCCqky4oU5+heKhy6nC9lX3Y1//3PQ9rfT7ckv
ZvFYs+zT6+3PS2gO2hkepY+RcCt/3uRzDR4rPSNfNxi8ZdgvtglGqDloBXt1UhEwWVvT+Mo/0/u4
nQYDi3/EEuPyEg7QQy0GBekCnOF2HyWRFfQxATAeWBJRoLqehdBg4t3vLDToDijtJWRThWFaYw1F
LZH2d6x1alJ181boTD3b7/KDDAfVmsCWTL7ZmiOa1NgQatFoztak8GzjGcVoWvSK/MKSqjWIrnrl
aAL3fwbo0gE/TR2twyBkdmgiJnjCms4EbUiRGfQNiQuGpNAnZysCKGPamj+E4FIy9Ia3roJMUQwK
LnNeufPlLSiE49o4IRELxjM3XmbwJs93oNgqP/wUB1I0u/rs/SMT0Aak3VtrEWYg/9hTP+Ec8CwV
XlJ+j8HW89okC5nTQYWKDSADTxAZEX0SSD1K6lewt9u65x2C8Lt5ydfjhAGT99JlG3M6V7330I6N
6kRlE5NE9aVG2E8oeeywXSTqio2AhkEg81iVR4tUjNyaH2hhQrND+yStI0ebJbDFSR9Zj/7pZ92c
sfULopWKmiskYAXynragNSVkBVf5LL4qdgPX6mitj7HpSB4bM5i63k9zbUKUVTMuYikjBxv5L1K6
qCabI+/cYISOxS/gUvrCCE/I0OY27bfNz4tLV1yFEHUQLa8RFzEb+iud8AE/Gc6sOQWKLfAX6oV5
XWmiI7wvulYxd/paqbfr9npDMLm3wfGvecRrfrISsRJ4rWAjkHu9nnG/1Y44ZelBVFlv8YzT7lnG
c1Zx9V1arnfbA3gpjzaJGwod/6WH6/1dElNUWGD3pYPMte1o+T19aBBGimhGGc5Lg1THgB4z4LKW
PVDWGmOgRDgUWzFTIUR1f2/QHpsGxapmlufqdjFX2UE5IXAowVrd+PGUcPqKM6lhHCHl98snj1Av
6THC1KMe2QjE5If5nMg0NtHOAP1ML9yWllwq1+idkFSf7kTPooEK9sz6lLY7/kfScvmqAxMZvrDu
XNjAvxrEttdjte0ntPKqGCljtgsdKaH8sTSFjjFz7cNmSnId2jcbaMZX8pENaCJ2tmVT3MoqNjUY
xyYsgQnEDboZt5Q4lVYp52TdxooVnazdhh6hGe9WeXD6mKZbfPlkITELoow72Fg11qusibDz3U4m
cvzVALsRwzSDT81pr0G5K+J/1PH8RtO+p6UfEZBRhdB/O9YCMfTkIpUVQODt1spBJ7IjfwsEHUBi
MbUzIoUmw+b73nvzHT4QGD5IE97IdlzuZUG+niEQu6VZF2HCqWMBhUxxYxogFivvZks5Pfo56XXH
v8+y+Gyhs1BWZ15ZFcEILhPAngTWW88rdw+clUyrL0Gl1C8sBL0vh3vXgSelnzf0cOCj5CXZRhBW
NYYL0x04RS9/LnpMeq+9n6EXRAcRhI4p3EooPtRY4laIxoo8oDvx3DPwe8U9+zI5kLPHkipp+b1l
rtK2Q5aBVLOwFeuqulChDR5mjgfk9QvS1QcEogeG3fOmUqJ9LPa8XUb6VBrsTSWeIwZsQ3T+7Uvs
TgigwD8qvm1BxRcK260FFuE1Vp03bshaibCtt+pyV75cfwG8bw6dDWEHlxj/iM2Ovv6CvnLi9O0H
Vts12bCefgVfQJPitZN4+Hj3PWMkEKI8PMj6xcWYivfIfDvDuEXS7l7eg1tnhRYXEmhmSFdL92NP
kW3JdFdAo/nbSXSHh+hmtzny8farLhFkyzVhQL46nuhhN2MrBW5Pyyr73lohOkzaTTbrJXrypI5Y
T8YGuyXv/CjcPxv/NGXwBdLfzPIcMDbQh4O9/oy9Tp7RgH1a10O08QoO9mGDyJ+pY/V+GkVit/Ry
Hkf4StnKuzf9H3F3PazkPokdFl2g4MRm5fpDVv9lEbdkmueEVTwlcqHavkT6YBfjLn12p/9wE3b/
HIay2KHfBRli2W8mDzjbAWAFZDk8UnUqrB0LcHUAFpotUNx/Vozq+wM7iG8GW3GwuFNfI77J+2CB
rmdaDj3tV9l/nUbdIJtIeGOQv87GbIyVTR531TZ5Vy3Sh3pri7+7I8jjeHT/DhIVbIVWfkXvaab7
PnU0Fkk5S2tHL0wAVswaW5I6L7nQkupr66zZrNwKSo2OrqNoIQWM4N2+JIwaJvYCAvsXFR691KDQ
YaGG1k/U3E+J1cDKq4QtyYi6vBGfk8aDTUXQcZ9CtL8NPbygCmo/ypQ7TX1b2BZqvSzGzzYxISB9
fzM5Mv1L3JosMj0NTxJEsPwxXjxMmnAuZ5RqfdM0rwuZ19VZWEuDrW67xI9yFUdHjtdtTUds1Eyn
9xqUo0bJpYy6nG6MHSgj0HYChFq58Dim3G0D2yQQNlfbLP0kC2z6XzN62SodH/00czN7naRQWD/+
VV1k/oeJld9cM9JybGHR0YMEZw15/W2sdRZ4YMzVsEIsOFJq6wpG0D6ktlsqZqDBMgP/zhPw5dsY
jEnjFMeYh8bp5aZawDZQUqf0AlnI0PXKix2/hagMSDSIUQwdOWk8cc27HKpVxZ0eQV01ql57kKbh
4UB4SXyqyX+2bO0IIpk4WDxePobpJGLHYP6M+1gO4TKbotsma3Uz8mtyBqrEAVifPQHwP/VTziyt
Dziw15fRMLK9ImpCM0JqGuZ9YfHLQNitBmiqpjvG0wqCYNyCR56fyMlgeW5xh2x+QLxBLVSgyxey
TGcqYU9/XXLp3UfnSWI5GV2VtcU9pdhiN29XAwWhZBxjqpN7fxOGk4uq+6XXgNoSUk7YbCBcnk5U
QlYyd3Q+gXsShiEcK/go28P6uOU9s89+j3qdg5t6/de9Nyd0FlXNmDA4u/f0zyp8x9wdAfQphUUg
p8wfKBHTCIwRh5Cw8vUqLSTNDX2Gf2JIYdEPQJTbSjH6KGhR6MWNa0IbgwqmxynHKwSkE2E27g/A
nBe0o+iyFvGYQBlIDCJnO9XYz5F5nFmR+t6END1nSbD7IfUFd2fcHeXHjCOwgIynjSLGjaFEzUsM
SDdcGQuTBUPCUJJjpjXXvSKy2Y5OnpZTLVmb0phzMuEKGtc1pPqg5UrtistCciqJqg/4y9P2HhO2
j28MkI44hJUsJWtbUVFgeCLjEi6YxL1ogm8IKA0V1lDi4XBtALABPnS7H5nfZKVQIwt4gHlEUPKG
mnRr5zO4XoskPPz4006nFuFk2sILaN3g5/mDiA1Avv8CCe3cR6dtC/H4VpEw5VCrdo1UGI4NOcMN
I2E61PULypiL5veDA/AVMEbUSjZbIe15zPyrrBBOooUCXk/qaOLaCHb8KJ+Oqr3hSAAsPrM56SqI
4zOzYYWRsmUKgzbhFffTJoX2+UNGWybBI9okeeRbC8DB/tVLeEtVU6UHFTxNp52yZT7CVWGlGCaO
FNgOi9Kbloma4FD5AlFfb0eyNsj4XrKKvjYNms0SdYiHMNSlX+51Yh2REkgZrk+gqr4+w0gYUCy9
gGqWhIV4qufZ3gIRid4tZVWgjFa6J5IgQRfGw9dyp2vmME56/Llja+JwCQ3kllpEUPn2hQQWV9wR
+RyrQTuDPXa5USZbUCMBN5H2j42I+F5FcL1CHGJwEGinR4x9/Cfn68t1/Z/8rJ2ASVqvX10Bhn+L
vdQpap0EQdB4yPAbfMPrZ2x3oqXVcY8cu9uJ8Ed1nwwR/UanTMR8oVqY0PM6Qbv8rsEvOsXNjNh/
RgnSz74dixPEQUVj/Nbo1zn5AMjhoa2SdX0fOO24L2ikDTmwop9zB+czvEWi81QNwV/vSsjiTnHl
C83v2ipwNq8uc5ObZ5hjypdSRlTJdmIjb2hyhhL2WCGF2CQRKnEsmsDSMA0E2urQbzrnaJjQ9hFQ
G4gCehd2SMdaQ8Z2Ck3j4L8T7IUntATYVfsTaOBypU2UqBNxYrXuGJKjUQbF8XwhHDCfudoPdnSE
g3IoqEApQUDTMxsjUjGoXchWQIqpt4WKhIF+k2U+qJfB5igBt6xluK+IaStVM/Cem0q3V/hFXRb4
JIzM2ak5RnAremPqvcW8N8k0GbyYiITKkvSSGbIw2rPxevUGB5JQmF1BTcKRVpqPuuIT1oUfo8wS
aNbEis5evGGzeaC+0myryEK9w5GcysiE8sUxE2IH06JE0oThspDuSrancdhc1uQxEwxGqz8J/DId
uRdU1x2Q1agNM+dHyfz50bQbHmOZDYRsEidaMzBAZr5B+noYqAN3AZNpqJpobT1KY/9jlh9+ZnCY
MY+Qd8wF/qiRTDzY3xaM5mgvTheChu2TtH33kpDKjhDs1nSLnmHFUsDbpohbO98C2mEY7b1kLU3B
JctRzfduvXIzPj8wmXw2hcNTeqPmZpUZBx6Hfo/XtFVQATLUuoiE5WZhjFUeS3/UMd2uE3CwAjMI
YD8pdPyeyuGsAA0I3O5Rmx84xqMUoMYgwkKAd4JL0J34Nxg88NDiEp43jafC/W6E7W4eOejpF+bm
zQMLs6eGg6oJD/pDR9qMJHVClCWSlnlt/Twnwf3hkVHkk2Eh4Od3BbZjyVgVtxg6j0Orx4Pyd2Ml
wz19PmzEUrGHOp+SzqeyVbBpgcnl//yK+PskkqYLiXx6zdXmRZwCtKgNDZ4pflFCjiwCS0UwDJBX
sZ5kGdnHWfPd3qyBCGiYBxYzWyw0/WAqHWjbShYSL+QNO+6kXlgWZTEjtY8SeB5OKCiPIVZqDJgI
Wx3dKAugAyupPsOARriCYQ2cS7RCPf1iZoECusa0s4WYMvLugVktl4x5ysH6TZ39uEW6S75EKqNh
fHKrlNC9pPpMl0SlWIH7t3x64fSqiOGpOdoUjw6Rzq4uY3umaa31k9enVfy3+D+3LLOSheKbAQX7
MSd68YIEgQNepBlz8GsH9GwX9fURIKw/8+O6xYw9MRQv05JE9rTa2E1zKl2iHiX1S6oTN6AVqR3Z
wywtOASsVG9tzrHCfb+a2yLR9hzZAs9aeye8mHL56NiOM86TbhtS+Bly23jB64NPmUmQugjqIHGt
ln9gX21SbyPnRt5ipnqWsupWRJw+PqSaMIwbUaSll2pmLYhNlRilw1Ky9qTttkWx1B7Dl4mdr9Dy
qYBZwL0UJ3ZcFZGAf58UUkKWhPBTkjoBcrQxrxXhFkjYr5JqGI1lSxbJvR24t6/VmI26VIIPMcW/
lIJDhmHBqv+VWm8+Km/wF100Uej3Ciz7M+sqDF2H+uoTkZ4V+FOzGLXtqHZLPK8SNbA8qO2e7EoG
y2x0FBdcYHaC2W6n36ced9RtCSiMZjxTapbJkDapV7iN1dOVHRvzEtBHW+nXwbCGQRtbreY+BHnm
OSEsQfNl/VPJYHxu/Tb3PkWQn+6QEA4PQyc7DQmZDkp7pyXYI3Esou02HhanRA0NiXxBwaR/pXDR
WQgHy/3z6ilsRcFKrHnC42UqO6jsgwZAq8yM+LBibzWFqEYZy9rE7NhIgqwgDMu9Mlyq7+XMvqEC
OM8u66quvHFntT65RGUuGBooyWMW11q/LyoC7UdoVEuk0CxVFAQ4RcF7cLB1g6/Phg5KQzWlQfS0
XRUP21t2otMmbhKp3c/LFlDPfu4CLoDUo4nrBwSDSAPrZATOZJtJDMo4QwcUlKcNGKfgzJ6xu/R1
s58fAMMkWq/xGUqQFl+dmrERredGAx3FTK/mmW42l80JBBVkCFKWGI/24ZoZuVn19pScTmo6LXGM
3yRSgfgYr6XP+/jvO+FYGA2OMVN4xUgjKPXEprLNV9CSFqkDDBq0VGXGW3gBo2iMI7Eh2f8vNttU
Zw/XhCLN59hw8Fpt6tXby0RQKIfs3Jc4eeK+b+eIgw/5ztOuZuNO/0M8XsUG6GW4GaXYq1PE5rgr
zydAKcrFCidsJfnZqNE8eV1pwJ0A9PTZ7m7Zb7JLrpBeiEyRXoJzVrBk/7sgsbxe8SWTROg1uehI
Mbkb/rUx/aQYbuVQ7IqVSEdrJ7HN+yFD1HIMaxWVPEauSMwMBkJ2txKMC8KDTflOudGyh9ikXFtR
iKBOuG835U5318VQtMZAiFhJ2hOpByCEz+KukFYUcJVC/NwYyu+5CMmurwzzjRVRdKTbKKoDzjwt
E+NPHHxHrGYWZSEMlOvrqwCG69QL09yOTqEaugGxXFdwDFKwtoRn6PHrlZ/vYS6ZqL5H2eu9sIWQ
dLxfYoiRveMi4rRmbvhkwhDVB1RsWfS84Ru+WXa4dQyq27erP8kvWRk/Ju6WdcqJA0Re0PD9RcH5
qKkK2RFeaGvbyyxQ0ylKoz/E7RF/hIbYJvGrLQ5Uenbkkk/dRESaivHOPACPnsSTbcyqhafklDR0
DoKGhCk/5KzqR22yNwAGwdaaXp1ZAXMO9UeIz+ufkyhEvlFOhSFU2l5TwEqeAPIjdxSLVovkbDEu
oYLLmqn7shH4Eyrdrd6blh5Yo0RhwGCAIVjg3xDAKbsKU/Z862X01GpMZ9Lt1zjC9S3ixrgSHin+
+lDX9Xz6gjlB3v523hxod7EM4Oi9s+e7O6xBKm/RZLddQSjvliwHlVinGNzsHLNbL/pu7r2Gk/AO
jmZZaYgwDJR4ESJ+l09nJZKdSzQHNKe/jwqztQXyQCO2E2xem5kqsKhAdoK/UE/vrlWOyT1DKhJM
NLFTi7894FLjkqIxG6ykCugeeUF32zCfHF2YHxlL4eiyssXCnf+NHZVZ1NTQDhEwNv5lkP5rfLC7
hDt5XdbwZOrdr4NznGQW8iaREYAhB0beMFXXh3eTitOyDVYOHs0S60eM8rE/AAcISPWcPV3Ozxve
bIwK8/dVBiKWuCC1SkUXTyYrNs0Bx2tkPO8d34jwBcqDw4lzbNJkIPMxMTMjas/yWeAe+YJAxlZc
a5B9vDedteTxW0IZh8dW1tmnQXks6dThGQrcthU6G454RgYV3UiBSaiHK8SCOgjWojiq+r6mFSPi
/UwT7QeIr4d0dM0xS68d9vz0z0cv1N5dOC2GEnF2Y6GT7i9P/g+XmSrLAhZ9v+VWvNeBZmDcAAei
2FCeLdQKXis6Tf7OVvJIh3N2id83cZZabJgMzsMAT3VzgZ6dK6PlvwxW3xaVGrxKQFIuYF9zpfNQ
ervoCaH2sBVrRBQiyi1rlgcNIsVzrBmhqOXq1fXF/XQh3L2yWfDunoMqFu/W7DRBFAcJPX/gjT/S
D2jWV/W3AufK3aAj7qL0OgLNPWIVQGEiOqoWnOx9pf+LfZsl9YcmSNpL0OpUupDQOU9evubzmdqT
hGK0/vJZPk4AHYJTIDyEuwHoQGklRR5W8JSMldeHpHnDq56d6yf31DBrmdIVlIkOGJs1+hbppgLa
mxOE3CShWVG0miPT7ct9okEj1zr0zjlcBA2qGYTbmgMDFbmiAkukK5kyrAXWt9nTtvMC8Bd+QOKe
ojxv7LEe0wvfsBUOQnH6hkxCsIrQEFyyyx8vZdYMBw8TOyXElobRB3BLdh6khmGXe7jr6qVlQj1g
/80+gzfEIzaVjgbj1hwU2rFgXj1xOAcLHv+DL/ml776dI6X4Rkom7nKUDyUBeT7hUwpfTLT52oxh
2pVI8DP6iZMI5rCOMaK4bJsGnpYvTgDqsO3Rn0OqqiDR/26eBhj/O4I5FsURYd2myugrBLKIVotA
uZCFM3QMWkV52xmigjIyA+uqW+6+XfOuUMRKK2oI+MyM4VFIAl4NK0cUH542E3t4q+6bcEFgBmdq
1W1d0nwar0xqQIz5H4pujx5IXh8Q7/SQjQmoR40m9kXGu35UYN7+JnLminjn7qHevkYJXhXu3ZD0
ZUXFBqjc0Y1M2HJN06M/MDZQlY/FQZoa5X/N8mvrfc2cYmzdU0DkCovQvpZLvOyV7o07XvbDMcoV
UIFLDqFF2WiiX5RAmBcpOCPReEU45d7KNtHUNf1zRkkSQhd2k5f+Do07rpQFz3soWTa28Jb1bEhJ
ms/N58V4A1i/XZMcNnCixv1RW/1K35OKh/mSAbg2+jWtOtxc3VctUs6UvKe+dHi5DdYIrYm7PeII
NJC02DFRkX5T2U0LFyuPHYClpoAE5gF/Nx4btZn201FPv38j1i7AlgUobA9lA0PW0AmoXSEXU/fT
tyrQAIL/gAr4AdkuRoYL3+IVb4P/3E1I6iAyovYZHFcwd0dsg6BXI5oLnxcaXWFkmZYxbRzxmLBS
Sl60upvux2ajnHrcI5Ps8Y7A1BKnNAErLmsG9dwusGT/1eG9KthMJ2dpJ2qzbSBOlYW56AYmnRrk
e11Lrw95Vsyr/MVk6uHn0IhAPIh1UFk3fBkAdw2Yt8EzH+7VXUt07FFSXhLEeoQ75STexJsBd1DE
XUZtpIZVUNMxDvqk4lVc76Hb4GbgCYac2DLCSfqcGkznCwRQ0XhOm3V3GglGFlCiJJF7jj8Zeu0l
iq5cCfDpMhMvCJuFMNysGnRvL0MUj8lxDZq46rJuI4Heh7Cy460MQ10PF2xyKlQNck5KB/YuJ0BA
AK7tUTJ3O9ibJUfURxhRUX7l0lC6WmimSeTW6RQRauP4lVkldMvqAyQ2LPMV1un6APXJnl/xNBuE
QiGlHXKx/BYqs82HJk9iWYvkwl8G4yyF2Z/u/H27kc3xXbqkQn5fZvCIPhd67ZTRiwRVo31qxfN8
yhD1mc8fKBA+B8EgfEQm4woucIkbgx1Q2yH0BBRjjtXw58RiAwY2DE67N+dvQtyvK/49VgzDlIpZ
CNrtMk+RF6FCicUTGX6NZ0DNo8WJu8AHQadwv6T1Fo8j4tkVOHFeumUWKudNxyY/CNQOPxyp3fvR
zTOZm0xKYP4qG2zwKlWN2e58oMTzbkTOC91d8r7StY66hYS/odRhDQUwAuH2kkLzk3Vil/eLS1F1
gIjwuvrtNMHbuGQFiZ+jcCJYaf4uhoPmsyHAB/ldxeS5x60oDFMy9S+x87prBEsfXyvUDSEwnM+F
f3RBFYP2RqW/7zLGLOQkCFIY3HOy7q9gDtG+TqRrhYH2ON6tbBz0OGI6UNAKIhE1En1xintRuAkv
C4cBTDpzf07tpF70Ed55hrE+4W/96BuR7t78WAj/UZTXtDrEqxwsJP4P4g9YenYltOYrvOc9fxGd
x5Ae1O2rV3EUxDyw/Trh5siIPARsV2FXjZvJh4fwdCUQ8jByY0uPwr8ISfVa4Zs1NtEVd+c8DPZV
qkMFrNle4F8iPWPLjilR+36MzjRNRNCsek9CcSSDjpyfXGjjmtcSgGFKi6iCMvIlCrNSDjoD1SRJ
Jdk03W4tshQCSJVu0t65rUXQrbFJbcQ+6FpknCHAQoJURMMkRKqF4bZNDMCG6qrnRSq2hDK+1jCO
GOqkt0q5dkjqg7x/26Q20HkLZjjwEFfm1kzdUHGWhx5Syk73y5ho2+dP3MeVNMGYdulr6Uc7xt1a
Y0QjEeoI3ER7MPeGm2tSYA1bzL97Ozn4Upgk1EER4SyV1f3OF8va8JFn6Ec1YL84SqrAiyE05c8a
0hozmseZlit8u3now+gLAKdDJQ9DQT21Xrmq7Ho5Us6c/LwTrQYGUkVv54O0kF/0COXsYSHjN0jJ
v8ClLUKQcjylG6mGcyXBKgfYy00o39uKsypjVZa/OQy7TIDWyI/F0L30sfBYNdlp7g8hHxmlaHuj
6RmMsbarzGe/WLFwU8F7z82V9cf/3G7jmIN5/154d4Zd2ZNNNm5OPbBma61LUdVGfY+tIyaYr9En
+xJDPM0wU/3eHw/UzlMJ56tl9fF632K2qKXG5QSxLzUoRee38FcoBupFm2sw+8DD0hO9akBu9xk0
aH6tTnBXqaPZul+mnETEV15JTnOpIMu9PmnF0Jl1IA5OWXSvzrm23NcjhNoosjTjw9fpGjo1VDRr
UTK5qGm/HAr+N7kDKLwSzViMnOvo5se2pT4uSMb/PdsvdW4K3UO1TibX97otrAKFxexsqGA6F8Kr
Cm1d7x1FMxZbYQo5obwL8XFPYBpQUIYh3qVV6A2SwskWQ52mTNk6V0R6WsCVwMttlUORQ0rnxXSx
kIRERgh/1qRbaQeDV1VVjqWPFPnaoK7ptKw6qKmrhWNOE86ESjup8ib3+rN4U5ByyHVk7CsSj66I
+olAOG1+k1fDkeHVqQ/ldwjz3bB8/MZFA92ldRfK+tlfR63nNGTI+LvxgX1cHZOwYnqsMpWG6Xtz
qLhzwm7NSP4yvXe38OkhIpdYIeVfpM8JaOPOsFmGvWprgsQuyyQqQWagnEzWLCtFC1Wo76H+5/Mq
S0equPRYs1Jbi1VZaTXYxBPZ1gX9pkdoTTEKlVINIxdfZMHQVzi+EezKT02M5bBpiANh4X68AUEE
IR5z9ReqCcKOK4eT3Wel/4WDGA+xgNtVdicEHTw6ZoRgWXgzVyWg7V3Hga6UMJdiQO+D7P2mGDof
Ytms1y3r5bwJ7YzOf6mKwh7JrSpxk7MGzLpcK6McACTZj27HdTae6RRE51NzrL+9qQ6EM3i/T/wp
hTfbUq7YPiD64XM9ACNDDPIIhUPOVjLs+u59zAMRfFnv95OyW1VZNjYEyqWZpFhDIQNmJZy2q8tj
dM9T26qtM9/e/2/6eg7HvEG+mtkvuafhyMqk08ouCz/6xpeCb/Zn+MowQ/PH1U2opPd9QuVT4lP+
gxmBEeLTjTNthCCWt4dWdGzqN9CkNhTpsqWYT0FW8x29z4lusj8q0KWgd1v3iSCMQAHV3ZQLnOZc
NWf+28Nmw0KBgWZEmEOI6L11W15RgGwLoHa3CWbNAnZ7DSt1SgXbh2k96rgNC+1PM0Rz3yyFVWgO
fwEOVY9fjrvJQ5eCVyIC5l5rscZojrInOY9x4k0AC3AparWUk7M16rRBP+xSCoR6ntCjWizuay04
+DvR2gx8Jprpr6Edj3KMNrP+TDblOA57H9UkVr13y/TZUf8kEAJJ4IXUBBEGcagNFWpFAiIfZ8Uq
GGHSVodfuBYS9ORBNz6EDBV7xArBWO0AcVWBITrNQHI0XZGy9WDRUAQeGFGyUOvSKrg1bHNUziNB
q1zxlk+1cl/UK00By6pn0AyP78T7UWNTo/JcjMDIaarqqWV+o3i1PYeWeamx3yR4y6Yzh9/PrYGM
96giIjX4tTQ8YC4IUcmdreacqETeMqG7PG96VyNrM1NVT+squ42hCRYMMuBfPvSnq+fRUQhGcbJo
HCQoXTbBWlDcWbJk2p+umFqgn9gLUfk1OFn3QWWIIL91lYvRP1Brq3ehMUX8orzZtlEckkQzjkSx
JzqJ9vlETpvBjF6tnfZMe114bcpxKQmFZmmd8ryBX9wDgbHNm8V8zSAdTFDztCcpa2xk54uY9MBI
Z89o5SIoGmJVap4HUxw7oMPa1LFBk6CuMGEoBwekmziOHQztDKbRq8Gq20fgmJH1PTDrhcfLjnUk
b2gHHvYVFc+dvWOFkNRytArKKTagPdcHNwPFcm7ENlCeUiL/rM/QEGZ8bkl2HP3Xo1vn240SY+Q8
hW195jS5hsLW2QMSV1JTgNuKLgJ3+1uOHIaJ/eg75eO90OTnv7JUDwAbOesA64Fy99BwBf6ty9at
kFE7/KVowyVxACMXj75Hd7EP4V77duuARJ2Td9OyXc5d5PFcLqVKlI6C56lAAmxjbhD93fF7lS0g
5k3kE2MZJHJ4EvqgZta2aVnyYW6uJkG3mu7iUVi0aNw9PIF+se2gr24XIvYfcZDVaxIlfBYSnOlD
ReMqEWNCgOovamjunXUk79ujCT4vQkj11qMD+zMjtkLI5NdXa6wQaTvoew3vZtSVEy9w4FzCi/D6
/zq00XGDTJCmgzKeDuZL3N4QWbBliE3Azwf/neWuBCVFGo4YEkfi9US+HQODMWyEt+ozwHK5889v
ojfZKe1hU46ZWIWQtMgAsN2sFFY4VA3p9Ba1FPB1N6Y8F9PPiez882IYVjyZ31jMno+I+p1po1tL
oVZX3OrBgPpUTJ1HUTOOrRLLECavexNHMBC3dRWl/tlhuGtjvoP4FI3nAEacTDSdxFR99rUFlQtL
xqfoIQIgPdVwhFO6UOG4wQQjZm0s70qfQp6QaaxgmuAp44bQQtWOccD8B8MnvT7WuPAxmTrs6sUZ
sFA3uungq/FJ78qQeMRkdZYlZVm9RyxSk6RtCzV/Ixpk404StdS8piEkhj8xjccOh0ujNPWxNEKR
54RXhoE4wXGvUUEo2MPyFNMioS+xFvN38tvzXtihzQl3vwwnlIbX0fAt3Yhki+C/0J+1fU1r6+MU
EZsT3KMeGoz8QVoWRBnIJNKikYrMOExy0plCNFOF23SxNSV4rcNGBrBXn5fxVgCXz0+9FAX53R/z
yMYHUeK4IFR7tSZqTfZjenxe3+vFJ1QwUs+EqsDh+xUTwdx/0FdQ+YiNd02gdglGr0CNJdHl1OSh
MFhuSTe5P4kXmY91J3zTWnhSWWLnV6+AuVAhRDEwtiiGT72rbkKr6Og7x5UeFo3n0ZhbADT5Esz+
SN7fHo0eI1fpFkCdfEJuNTfdnrM/SIOQ1cAZo0q5YFeT+ouRIlOwGL2HUM/CtNy2GG2QR8MrCCgb
imcOewJMdZ5L0+N0nHphFw/L6TlZOOHoL7eZ6B7RjFZJeMyULsyLJ6PzRiHZz9+RxhkCAW5jG7TC
kctZDHv4ULSvMfBfgFB1BZSov3DO6BCMy3gCNTEOK9vO+Rjq2J3u8W3aPcEMnbkx7fwWzHLErk2q
wD3jRxL+kOmvNjKtxwvqYn1cgPmitgyV4B2+d3f52Yq7uED0oLMKUmWgNakwxzg6O2XWaliqFd0r
roeYn+NSQITLXlhVrhBw3uemxsPLbYgZB8Pdb7Z13io7QBkirHZzZklfjfBUXKtM+UbySy675jwS
3JjNYLNirrev7zRkuJYDfmRMfWPUyRYRJ8MSdy0ujeQ4xs1Tvm9uUlXc026wZHoo8mOLRzBNuZDr
7ynkpCRXo6xgc2xz3LiRj70MqgrgMOYn9fELCB89XboH3uUPGiQQziVctFpAakuoOC7353NJ+f93
nP8bJGE+RF2rd3xJAwOUNyKswsGaY/rQoKfpQvcS4NJyFk5cUGMT5dcSrMeKYGW59cGBoJinAKb6
8LADFWD0wTY8x+xT98YMR8U0KUOQB5zuLgWRtJXXkyiukK3lEMw72ul1zRxVvnNpL7DIrnXkqMFm
3YQf+98MyjoSPiMUuIpHpG+1g4lRmscYZspN2l6pzxifEbiarf+pXknusIBXLmFrZzUdPcvyQNFr
dS7F/IwxxoqQ9oWsmpXGlDjNf8fniYsg9cMBfIQQ/jbsSQBXoz5qOpTpaD/0E1cd/hiFW25uWTTf
Hxl02B+wga4XxxqDhlb7vL46pbhMNgMNIVfrrrlXDQPGw+OlHViwgRxGgifsqcv8bWSkW0xlVHia
kAUoYqdMafL1jn2qO+dbaebW+Bh147DlWtYxY59Rqg6hDrpcYbW7q1yNZz6GSQo9O/F/njPV/AxB
xK7ilDranyFeFMk/ePVmL1WY01L+WRSW2b2sEz4civwU7QqKPr9uH5JwktuTQ0X2mdDoduTDllF5
5twu8V/t8RBJijwi1UaDJVTj8/yxaRYQqJdJE9ZqBUKHF2Y4J4agba4kqld2a8U3+2/aL8hcZINe
HrRJkV7u2dPUj0EZgFt0WzJAwneid6+x+1wK8+VUgU7tDqIju6pNyw4c69C4k+gwbdwLtAkYYnfY
j/uiZ2TmTnuXa0SCIQJiGoiSNXOMcH+G4ZS8ufyhWqGbj5Idt12JcPJ+PRwVWWSdf4uNdiNBnRnF
Kr/EVFtJQyCqbif+CwkenGd2c0AdNAV8HeDg7fc/7OBIn68Rlf5nzzJ5T26HEvMLNUKLoHTT64I/
GffYXd/5q2HdCDMToO3NVdykVm76pCJROhcRr1OmyUksCniYABOVdNl5lGEswt6gqz3TbP/uwPn9
BKC8wtlsbLkEwHMzPEcmABi6PUWJ7jEeW+8uZGcuhoA/v3/qnZbJmAAGNgWWleIk2KIqBBKFlzqk
OIbynLHsEim9zC/HQylI7qdZd5UcZPAL0N1+Gz45BFqqkZxu7Zcr3Za4MW501aWcBkhSTGyz1wPF
EQzo8/GmcBC9hQhwk5dvyes8gRHvcOIMV+bFUc59wpzHBFszjYz6EmFBUZ5UZRpfPY2a8fxQboq4
Mf/RKVYXTxqqtZDcDDlDDZN9+T/AVrPSnkrU9Q+Tj9W+vC4FT2bpGC0/AD8fE908wUMZli205nzL
Nv/LgYnb6bGcnLvG/F4ZuO9Df4bvDPMO2ge9mjXz6d10690QZ5OVQZst3akt1WMbvdlPp+bFFZDl
pKlNXyPaHRi8i8XZj7XAmt94jzLLiVRqClKhsKDgLe5nidOS9rch2QmRFLrGYw/3HKDgTKxvkyVe
7hqUB7CeaoCShNFj5lv6NFZ5Ivu/ZL/39T66Ka0Pyj8vLeiRoY8ULEAEql/L944nJbovQ7ZBQE6S
XXJE/ito5ltyx6rijhagYgxeF6cXAT6C+dyAqes28dZs+6b1rXOHa0bWBsEvxOJE+b8T9VE2u6CY
Kxy0eHgNDV66giQT5eL6DnF39Pjvu11G/S4u6coAU+D7TzYf0diFV1fppDdPO4UGXw51+f4nVyvD
cx7siTVc4fTWNQwEx3nR6IJopkZcnkACgGryOp4bLVg3+VRKcQ5tI9LAGyktM6reF0Cobts0JBVm
KEFmlJu3Ccmoaw1WQ9xX6SVLO3dgbDiGledKRY1EvBr3n/US4xFWmwSSUpjVT+KdzqNa40vaVWl1
r6V+3ir7OscBwOkv8TOmmPnPHY2UOsKRh57SQ233ST253St6Z3a+t3/3wTVFQBTpxsNcfLmACK4f
yLxjpbxJrBWoOWGKRb5hWZZHKyuKERZkE8vgNaHm+c9Fj2QLScqLJ9Sl26+OhyjdBlIkgbXhBrUc
I+FEdEbbZraWYXovjDPsT9yw+JQG8dPwk8AhaUsPrsLLrl6l1leI31F7eYv/803LzKsztyk0Ucx6
Sb6jh6vEzaKS4Lf7NEx9J6gue0WvApHxLjvEmWL2Xq9OrDNxiQdsfkz/9APTDRZWfOQrI+E82+Do
llk6pyhk5uMc40OFoIjNzeJjc2A29N2y6jg/ZhOq4yJHWFrL++IFQ2mMpbX8H+jHLTSF3HhYPi/r
ZC4lUDOB8MO3pnuzW4m/N37vfQ7ZE3z4LjqlLPBDsaXe2YDDeSNncDSQvik09qYe8vOLWi/mR8oU
roW6CDN24+R6NPl3GwwoUvKhrE4IApnujUmBbVd2T7PpH39kaH36hP8Obs3tjxIthfOO2M0DU4b1
sG4uO66WGaloIdcwPDjSFWpUwrQPu1RW1PEONx6mxCigpEil0o+j3WALrC8dOvDIan15G2vhfHdO
gQfRafy72gigxhnh3kBsD+AcUqNZIovRaa8aLUm4XXAMD19w3gD8krci7LQTQDliytq9UOVCFJYL
+pYtYoVrnkR+A2li+xvLWVhme/kOkIj3LqQDZVo0U8oOLjxgtLz8yZdcv6UhlRHzoxZBVFm80ajA
1xArku8mGM9bA2I9gKVilaSNL0YZvL9GrbASlQeT3ZPj59HtQmHQulSpIauZoNstA2xsPdIJiEg7
XoH7CtAXFvyMz2AucAtzpXpa+ST/Y80rZ364RuSj57qPdOVa3E0qnolGmGcAbcOY4dkzfz/oyfDb
3dRepa1+B8sImyR5M8yPTOCAtWon+wG1ASyAL6dVFtjhlun5fCdWIOsVb7xKWyA/IKTjTkbR1irA
tqaqh6PFvFLYTInZbfAdTNJ039QBOXi3ZzQaTtFEZaRKLWBJd/01cymE8YdU98s/Ffoe1GCsfYX5
StN4YK1VxRqitsfqUfTSJFqgDZgEnG99xaG+CJ7PZKDmge3CKV79txscGRNoDb6v1MFZ6XiIaHeR
1jxEK6fyiauAuWnKC773X+Dw9ew3m6KCadHOgqGkAugXlnieOeJmEX9TaMCex/et00BSig6/tjTO
7X4IXD4z2PMktbmngfBdmsjKy3dE74nJkztRXY0J5dfKJi8Sm8Th1K1CGZPNLkmfxhEbzOm6adS3
qW4ri6yO2yh2+7DJ8MFhY4Bg22o3toFZzEtWXVhuVLJqLjvs+K7FTC9n08F+8sFP4qAKp4BFsMGB
5rFxyv/pGHdbU8LPio5D295oLoLZZwRCmFNz39USud8Qlw7cDMoWlVmHhBDtZ83iY5p152FNVFvu
yfmTjDUKF3LuvkyiC+5XghzXexaEuOabAdriuUJMar3YtdnTxdMNBpr6lga/dge+nTso/CWiER4J
fdNVbOvKZBVmxNIc8WfpauHf3ej21Md8184YT3IUg6avzl2npmnzCY0DcEmeCHc2EjC4r+d3kOsJ
dXlXYBnv1jtqsAl6gYQ2iu1V3P0R4CuBhvJLd+pq1x5mHijI6nTne6Fne/RdZdzXxSXueSY/XAZC
DqY3onjwSrRJuZ/mTQwUV7FnHT+rnMw+q8YGqVIgdkWRxwgPpg7KxMWsNGzSJ5H1WCnq3ztKDX0c
giylB3FWtNbwBL8DlEf4s3xaZPAhg305thzrtOFxYOi3BYfBPFC5CxtsdI0T7x+0ChsV+Ou+VIwO
D1E9kKk0Du3LtCrqukhZnO7LA/n8Bhj+7Rq4NpSy0lbrGp4I7bamBy+7QwbhU9CrD5rASgGQNgv/
GElZVB0XAXkbeqXtlXgTXPu+3cj9SHoPrivAJ6dVPAS41Eiins2fEvkIxN5jedSs8XDaCdVkgab0
FZIhlu4MdmwJRD+fJO3VXssjEvE4Te5VebLy+XC34X2rYH3qlG2IXNNmhBZKl0Ea5w6vEY4NqDVo
8fgMS4olCUMiUDCt91ePMnN6ZmE33YacAZdPRE+XCzgefWHHsLWcALIT4TfMF5/z+OUI47V649de
qHXZwZLTr/WItUBytT6cSR7mGajZ7SCWs56ZYLFNrctGZkUgKDCMfcXQnDg0gsCVCnosmHP50CvQ
BhwSdRQTTQv7LGf0nutKowGkI5UHN12xH9T5VoFmxivoXA653GoyRgj/UhrudCXbhi3xKxUy2fZA
m5RCGeCyVPqOqnMzYZvyRFenXOflg/KfEjxOz8qgc4o7qr4D/LIXSfgv+ouBIcZOi25e6xV4UN1H
jU/7sZyphLOmq9J4p78TVbbVoLkszWKWMRdKrblF77iyq2FcKrsfgrjoeh5xbZcm1GnUyT+vzSW/
pVOzrU3XFUJ1be1NOEauDV86mROldsL4hUbJUBPKS6tEPTlWYjby6q7BGsjQ9OcaE7ykMUL+ymhw
iio8jjvKPVrU70OsRoBjm2hi61tm0Y6tpof0IGcFilC0AfYnPlTLhGptHszcgU80+IfSh3kDp5k6
ni5eqoA4ozFClbalKB9rqXXxwZWyf7lPXE+571hMH5zhy21hcsBIMsjSwIgc3e4O10pWBmDJ5TU+
Ckki48PzHGeDorje4QCMTWmu48/xigVlqxszL7j9c3B+Q8lJ7Eozm5bddvLi+auBdDyB7Pli9LaM
agNonKLZVjvoVN5ja77OQqGjK6Wk17cgnVhfVU27xGxjr7u4PKjZMCJCgxRAH4sEd5bmrENLk/xS
D3YiSWlRfh5RhU0l4LMHrEQ6DD2p4+ui1WN4E3+50Nr5d38Jb5WSG7ONUgkcQOjs2xnh58/+77Fv
feWEqGktznGMVSnB9Z6Ug4kJZOpqxLBicLocieMsFUhYfFcVEGXCBu4KjC+uh5ZbWDd2XOXY6FAG
WD0V3ZWO649mOll14ZBTDu8Y+BKi7OygwtiTloOrrkQ9FLEYHyy3srg10VqPRD2KhF5dCah8badJ
xmwAG8qH8RBekLTzQjrrTsibDMWBcFKbcBqPih8oQboPHgPh9Athw2kYTpjvcbp5LZRCqIQlzXIb
nyHA52NFOUDb/fAxxrY6wXGStS6JnPXscboaFUO5J9Aa47+Px8fxpNhhRZ8Eq5XLr3Cns2fqgrCi
D3dVjpPGIPePY1okic4QWjK3du/Lnw3edz3HhSwBugNO8m/ve1T0q6ePkZNp0UELj07plU9dHwp5
sTz+u/MrGKPWTyHoDjj1RVjkoVA1c1Wh7jFIAG22G32rHvuf/1icnP6YxyVZ/TI0GzNvSdY0Sy8U
AWf1hbSaUnRJcA2YNhkmcvtw3Sid12z7eC7l6ygh0ZBnn4B6FUWn4M+6cVJttdmAlYI+3PGMlEkw
34+LyUZj2qxbZ1pTEdLpjF7VhoicaWzYiQWE0ToTkqo5YAOCk0lEOzgPl7cCQ9CslvCtyfoV+ZlN
+8NSFdTvrAW2fTMtev+9/dRFd2/Gzb/IOgTgZJGb7BHoxB6nQz5RpbMmI9InxIfV1f0ZRktDZAAO
pA/KBHTLx8Uom32Z21d/cPEcpavlKT4vIbJEPXRiSqf/9IWE7WSgTUmJcDDYwfCsONWZMhX6CGB2
CqW5dOugQ3TJl7T3O1pRtCwvG01IiRT6f1YZrqhDZQLw10TiAk/xHAtG2v0I2hdesRelRX3hMAMR
8d8Q29UBpzTpVJfzpN1NG78vP/1iCe6ZkyN/HYU9Cql+JpSc6TnN2IUlVyQAiQ1DLDXteiLHfaKl
2q7oQIM+iQyC5x30rh7u5U0fPagjVyya0MyGhZIO24TN4Z1qNChmcNoCg5odfs+ZQYFsgXM5Hg9P
YYmhfEUm/UiU2XBMgu3PGo0mBZ8AZtaQeeHzf/Ld/IBeecrKlNMIQhdpy5Y3sO+OG82YHsmGLQbg
QVgET/K37Jqzb+dKzIo1KKzrwPiPRMFNunHom22+v2L+WCrjXMqL2hqVhtw6DM8wgkkNf1C093j1
dM5vE6Pl5efqYcbAaJU/cVS1FWelupthq91TnSMOT2kPFNH/R9QDPGQohLOLqXMFkMiUOQaDVaAE
yzeDxNeBmVsq1rq/g1arUL4c8d8QV5q9F4qZ1VU6lYe/YMW5twDdXSqdQoybHR7Hds81x9OgIc2R
/sKGfvlNtLqqRawawFA4VxCPVIL0pDPYohLR5ga0IP3vBxMvCPMKyu6FthbOjki4IuJxWyvCTfBZ
udCGh4jMvrUIvFnieoBpt3tq3kv+pqyJRAjI2PcZx+RmhOzpr+nlzyx/wBCP6lWWNG4oJT4htWWy
jIc4IIFv8gFBewLfStBoxrYatRAHwt8RPYtkCMcXKRNm2Ozk/8yv6b7lZ53QJ5fQLZCl6zLHH4tn
glvisCDEp19e+o7mvdb2mm+iUyf9El87D+qft5nHfzdq8yAC1jqUBfHfE1GgCuzeXuFu8JTaM3k0
D1d1w55EtiYCsMobgEesRB0smzMBSGa9yR/PFZfQwQ1yFcZlL5vdbkfAdivEmdYdbGXttoOfErO1
dIqPV4/Zbw78Q9l59/T2dOayKZyKnUDzqBt83FKtFS9CXNBN8vdtTj2hxE8JQDcP8Y1eLbnOJv3+
DmXe/rnUmvZg749FKeN3KwNGIlStMYwoFNPENVYgGbK6lVgM0yLf8fhaBTBbpKx0I0qt8w7vrzbY
W4hDHyiKKvBCBJ7JLYkjael77UsgLdv7xuhfMfoHeKkiWXastSMeojh+Vv6DecpWO/bzLLaf+e5V
lh61hlQh9YRA4sM18wjzhuEg7x20tndI6YAxpboAt8TPcoyrYkFNak5e25mMDpQpcb0hvwk81kt0
gQl+49fKd81bdWQcdbVMHNu0cMoyjKTwL9Cc/54x4ot/mN94vu0Ww1ZnZ+RrrPYVP0GsuXx8hyum
F9tDsBgTi+H3rdEIN/uoR/48gIDbLXgTYAWYvJHPoHbZ+vvf22xcV7dh4HG1nxAeuF1p5USXAdUx
/eTA/NxuzaZnAvGCPM86ww22fWaPEoVmeMaqQUsgIK7T8FeqIiEq8/UFgjdFX/pugBy4ywPKtmKW
oHULNMyyezhmYEASwvuXj41cUvl/QJFNCh0/qdQAk0FSfhm6YrY7Y31mQhzrsS1qH8U/RpM6op88
eAVFKUcUqcF7y7f+IbF1bc9DUQFJkwm4AeadhwbCDpsaqBZjSUDaoMPZ0CGgY/MUCRejVetdAm2+
B9QINef2GofHvI5sdRv/gHjWhti389WhrS9RSeQNJvc1YzcAJEQ5O1uGP6BKBuCpvDuaGc/bZpnt
Cjtj+kYE3GJ6UadxtX71NKlpk8DZCtBS6+/BR5ZnSRhb3LqBTJKnT7H8aKwOuUsWUtiXR5uaamF9
+n5CJRDESmchzSR1l5jng3B7KpfhINDD9Y3ucIJpJQUlDvuBp2sXaB/OIqzSBj/UZoNWR9NQhn0S
ZDnBFKGsvhXF+jdibAQ2T4K6OLpB64gSe9JcNcTT9BOfiUvhoxrpz8MkGepSI1Evxz5yX2NopZTT
vsQ0hfyYKBMqceVrozplmLWuroj4Bn11I53zdBiUp2MhbzMYLMJ2MsblVk5Hq0ldrADL8fw1ppNm
VGCfuXaIwmORf11aLchl9jOxAUAdtvbUEw6qrEe3l2C08Nkphy40ZhG3K+CYIEkvC5EAcXHy8pE5
HR6GGp/bfNmRfDTpa0AXQUse6Nyf4QV6YYky6liJa21ciEDyuagH+huvCEPZ3ifQdIrGqENzuSDb
qFBd9rCWWFvxBvD44CkaS63IUvM2seovb8sDefqpIp9BJOhLbLjVD/tn8LR1l0IuYnhxetu5vafa
83py0G8vfdfGSi5jXoMrkY+dpmh9Llu939GeRp6KwAhBeqiP+KACr5izCIZeBJMGF3Ckar3Te9Kj
4ndOOxprs/GuREgxxdehJ5kNzicnOVs7JBtRMURWAqPX0TahrVdncmUA+aZBdDvYK5e5Rt6pZZ1a
9yI5o3/MG5fNq93r+wZ+Fd98ywdBLdZTw2qep011gAF/xuUSwJYcm/VcRn0DsIs7wXBO3rciNcMK
RklCj0O1FWuGFXvnn0ge7cfCTiubDWNKL5n34+h2BNjhKtQMjePwGFrEVwPpaReNkLrC2o07itrG
qaZIbhiGjPayD88mDEoVDQoOjtrMWFXQvBufOTxyDFYdEYeBPOpJEj75XiAFKvSCoSNtR/VTDRta
owhWsLgCrINy/y5I5q62iSaTlXsJXj44u6Lbbfav+wKzhkNJGq9YtEAFBknsDSgl8m8ic3AigT4X
C7S+BZ40Qo3Qj+2eJ41WEauSjtTqu5N3jyF5L47835ggRecjm1b2x1Dh1veOeNYOuG6XPXFfTd3G
q/z8Ey9GiLBq5QIz9XFaKYsxEO6yLVw1cXxFRug09CrJyK9m+1z85+U2ls+oVQ9G141Z0R5ehQ9b
5liuqb10xiDtI4HtFT9pvRFvW0BBuwV8wifIxrmsAVTkPwrMQm4CH8HuiZLWrYQGKfe/LicjSU9/
bsibHBmKXGZmi87UjeB+SdJGT6WFwhTN8bGJzupCOUCxu2YJV3gCDZ4BBwnjDje4DAz2SvCwRB96
rCNC9k1ybaq1Udv6+o5RvY8g1+fTuK0BIbXlSJAJRWQuRgKLm8avz1dNrpHPPKRvCRhaCfxEQ0Vy
GeshrGhv2tolGF8OpW/SP+Pz543awgVLwl0WzSBTmbWFxeWP0fW49vOIxX0M2T8N6mpqfFxwQ3LW
3BvTodbBQTfY+g0jChvgtWbfJ3alJ3bnMslv1aVIBlXcqjtYAx+Mrbz1aNuMhkyhmu42QfV1xJL8
Ladyrsv/Egt+oLSe+LNzjhpw4lV2Om4bDLhR+bMFF/mkvGEXy+rkLUhwIkhjYB0EbgZv6QYBC7zv
6Ji+L2mispgefAw8Owp3kxneg8i4T8PPMPLJyejdDvZV7srdBDbww9+FEIFyb76pjeiRol2dL8Js
QakCgq5RatNP5v2EoQytpDc7dQabt8XBYymyg9ywDLIjghsmnbZs3h/VVkaa13YWKG93J6JxFE9k
D/x5htwp/RpKRtdhL+wTGwGz5U+Yu9UskHhxJMggitWnjTYdMRgkUS71LdPfiBwf9ukc12ss7tuB
YB9KirJHRbCypyfp/kuZeTqTQEI1tMQCoTJEzkjD50Xa7apujajHixafIxjnHl2wEsoVb2ZKENJ5
6uJlu8qpmwwSmHPY/eRb0KH7sYxHt48gjZ7Acv8H5ZYS0ammsXmGUStz5t0M7D7DoUfEmHiKcswt
uNRopkewaCsgJf0nPUIpMrOLheMrSxO491kw1YjJ5zdM2rUitirTolUF+SmRIhVnUCod7GmFYlbd
/C4Rvoz4Aduo68CfvNpWxg3eU9Z9iyxvFBknrn5uVTcmHgxdaUBGM3AF+EjH23KYQM5KcbK+6FnW
uy4ZmbWjBLLHj6S9w1k4gcYEPn+QujvcUrf9xr8hqqW7a+T5+emX/0gR7WZQB5F0HpFB5gH8XuEt
t6M835KGimkjhtzlv/B5bmzewM1sifQxBh0v8u7gtijv/lz9JabHoE28437w8qsmauPq7Gk+hnZp
5mPN+hAvD99ZY6+pdE9H9SfeCilNMCYxIstSK0ToVGAyob5nUHWfXroSdtn75dZUBvvlnRg0kHvk
44vUc1blJ5rJRruhXa9T2rzIm+heElqLImGej2PDH6QRKrtpAtC1Yy1aFs3vermjNmkCkcTnJXZ1
RhUM70/wUgsdasH34aMBgGJ6OuG+LuwlRzn8pxgxUYzJ3QlsQVHAb+np367vt2Xv6b0GMotUs9ws
DbyfW53esd7gam5ikmfpzeoYQfyrJl27vCKRqSjPcG7D0CmTUsQ7heva4jrFvzj5flw2csjuGoyM
5zdBuaB+2VT+rFreXrFFGzzzsSglBaZ80assLuHIXlIkPDcvioXezaJHI9Krqv3+RVOIfvn0Kytj
CdA7/5weLJQQWrvwHTxcSeysHBURufZdQZARf+kny0pxurlq867FEsuq3jZA5g+1V83j7rD4TP6+
H7bO1ORv6QjCXrfRP8bfVJr3T32HNc3gn7GCSGd80kfcH+qk4cfsKFMQd4WfOwn+ph14g97CB6lo
HL8u7jpwe0yWxPMfs1nYShlMAdg6a8Ex9KhOxY2SxGon2rw05zHZSsAyf8G6AISYv1GKMqwmqdYu
3sGKf19QfMgV9tdEroh+hK5yGU4X7d8AlDS5Akj6FbSOkfZNzl9jDiW7qQraNRmoRlc/hyOQmqjB
B/UKn3vMaljdrCerMpOwkMcG8qlYLBw/OYozNjASfQTwMKvhRt4I/r5LmZLimedVCobUHPK8BQTn
uOBUzE54+HZEyfECQ8T//JYKA5Ktow8ROZvP36Gqd75f96o+jMtmSg24j2LTSaCtiDEdESlyq4f2
jDrtM32xffgO9BLqIbmuA09GHu2UgK93ZxY4QqAcpIpmFkjVIRqsBn/yKt8CwKInsl14A73mUseO
YsatyOWpsh5vCdzalnH8+caO16el0V73UoKdYHLTWH5uru04xyMuHmX/lt4ZbofBMHta5j+cg1O8
HaT+zmvDyvl4Sq6hFU9mxVfuw0jzndsvnAOeJ+hn6U1XhcPrEZR/JRSkBsezNmef4qG9xce5lyHA
/JZzxArGv0eTpUEPdgOARdOrB9Nt7ABCd0NemRQh5XtPOJ4NpfDZ0SvxXSEokoiK/He+asj0gOzg
HYdjX4OhfNlQziXDr4emh/fYO61bfUf/RdcerdQoFnMoDMNMk+piBxJOZer/9qRTF7uxurqUVnYR
omnK5sy1s9Rf2GguOT/fszPV46q474/YoeiCBW3SFHD5K2eskbIiqYY7D+3biJhL0lytktoAxTfW
BN0BV3W7wwdLEW+prDiBo0TG1KtchunLzP+jERfiD3JoZ3vgJ++owzwDPpszAupDtwt3JHpi+sY4
R1p7P6U7Ly57PIQtPfM09K+ZpHFs7Qwd31lCBrNgA1l3KIQK8hIFnoKx+bfkKxkHW+FUBKs7UD6i
Illd744BHCFlm+zadDEj6EMGj9F0Y1dbSQGKPxClP5F0NpBUHMRiwFW4gmBGXAap/vL0tN1wVhxu
iFUgulE/aXEJkpeNa0j/C5XedTr2dPMeNaUECAX/xZEHrGhBrWeop+6QkpUPMTJdNG5Tt0rROkL2
DrLrU1Jj6v8vDCLMrKkK0S5J/PczxkqEFemvazkEJ81bcba1NfHcBs44MTMElgLYO+vkywCTAqp+
9qBHoLgrBb0RHVxkO1UVC06Gwzyyb2/kKS1q3RW0H2azCadnWPCYzXUPJTSh1UrQFKODEg6BXfc6
3urenN35cuK+1evuXVWZH7jgSIneevmKZKC4WEotwJiurXszemAovm5Pz00dOEfs4oBWbAXpgwNh
XJRExZJr7H2z6c8ElAhqvC5rS2MTKA+1eHyq7Fkl+0jZliYhyWco2LQ/VUulcTgubRIyuGMlH0mQ
02MIERZTm0F9sGmvleghmZhjgZzYGoxuAg2kwS4SHlkGCcEtJ67FvbOet1saSEbmSH6dWRi/O+oX
lAEsmU2U0qY+4bWszgpeL+qsiZ+cPpDT8gOPSxp/KCSo13B/04rWn9ZPTEPw2RZcuv8hAKnhRjC8
BPxjBB6ACLZRhNk4JJfgMgLPbUm5YvaUxj+3N8HLLQ8IA7xBCmtwuArzyMnCjyCRZfFKwtaOLQQ7
0UCjpLrU7nIw3kVqx4QTvpm7YODNbZla9hGXxQg22AlejiOFFsr1cKVvULkJxFmuUw9e6et6ZNcg
fLebsc2QDiDw+ukbsVIDaHvMPQR1/cWpSmwv3HU2jpoura8kFae40d+wY0eNzBKPohiB8Jw+TaeD
AmClEk3jRZfkAaaqP24OFTGe0qEJC1d5tmBNZThoVQ9Fns5E7qtVJrRire8BzLWiEFOrf5uconP2
7YOg8yRK+R8SIAwKVwE7mKdudZleE4asN9bJQ4ucfz1KSbGAFGv0jkjqv55oB5XZrEgK/tBzsQ25
VS3lcTsCi7fqm/W69VWH7yST2jREVcRXk+kNnrFVzel+3SN2nZLfhbAb9fsrLuEBpglB0SUhLYvL
65ysILnhR6/ITT5ENOnu4R00UjT6g49kWJtmAKIM8ilL7YWrtPlxp5Ty1MhotoDzyt5lkuGnra3O
ptWeXXGwRm+uVrc0MFH867oPCffrKaad4p8Pffz8ACTh6iTrUDqJmT/cp0ngy8W0KLcUuxJesCkx
ScxXYZS8f5af/Xq8HpozfE23DH0vA56EPX18cSiJZGJBRBaxkBSPWEh5vidEYg3UjOxkuq/owaX2
p9B2mo2x7Zl+QfMWq15WyH2xu5iCVK7MzXW4rcFHsMuIG4UuYRVDD17PWRLxdc6ZxNnxlwquXzWg
ltmnFVcvwZUWSIu3DVUZpT2khRFSR7aDBlaZM36hFhbXie/0lNXOpQGWevlqBOw78eehV9OOo7pC
SigpiNS9badWe9wLQa3kT66fcxwHOdjibuZnAvmWuJ3d1+5YR6XYNkh0Y6efbG/gtLSCxrXc0tyk
3M9o2CqMKpbTIAHihp55rqIyQvR2gxUglhSL62ijxDEOcdPxhWYL4uFBDFcIznH5FfOv+uwz8A1Y
qwgcPYX+FniIMxa3Apng3ps3doOd4puttYMpgE+/nUxnDfkJha7Am8vJxBqXZooz2P9byNoZFfwL
gX731hHuMCgLIHJei9g1EIag2NsQpWYZaKGpnWmfYKWwNX2xlrHZ/wIU2/YUgIWUWV6UhIjluxDt
0hs7gE1sHiKSH4mabU5OhBNfr4aSTWPgCFL2O9HbohebM5SPYvudbrlz5pXyldynkRGw/Aszxn8t
XYCdI/JUq+ZwgU69/7gAsDrg0yOreTU1Gn67b+kS4wMmI3LY2QKwSNq6mBJ9zm1r94m2KrdP6wXB
ihbUqB4In7JEf1RTmeTzoUWRN36jSdsXSEswZTTWeWImze1terwBYIK5CW8A1qHCklWRmlcWmBsM
feBCc4UwM/bneRzmMhH55qqQNn0IO2kYNeWqCNys9id0niwDt//CYJ330ToW0S09C6eBZMCBl8GB
t98OuSR+CdGwYzh0idy8Os4MWEzZEVNSWmhGqj4XIHS7p/DtJeyOXLhrirH7Z09R2lXUsVkI99JG
8hLTx9+lGbILF9XOBk6inwwgrTAUvUjZJSgz+/v76k7dlVNyTyfq9J6d37Q6MMRnGSarrhmaB9cK
v3E6v+rUC3JEjElv9ywFc6Q9qYW8JE1ESvhOUwvN8lCbeVuzCv0xxO158nfPBM/WqZkTbWVxRMQY
eDTMVMy2MEZOgv8Hw9HDyILgevYlzTIIC/1Y/JrvQ6z9GxFRSsE73MpJVO8rp0suHuR6h7D/rxwo
0JuBKYGcdceZbNG/5koVRAIfZ+O3HRLcpTjrDCEUIu+hUOLXSM+hVq7Nv5Gb1zspHC0JPXlEFVOZ
25qiu5CswBsuYEVFMIajahwHWt+JKxYfm98v3NgoHTj1D52LmRvDsRj+uKAgZ6+uBmJwCwFhBfkX
W6+j+aoKXVWZ/KKyjalNljUqmoXx3smgRNleUnXuHiOV5PmoOLwEPfTxHwVvj+2NZ+3yJFpSJjEd
Nec7xQI3jcTlfhJmnyB0xvxULgVeBhJsszjeFKawd7zTIWfiE1znB85z3EEjG87iELD7wtyUuk0J
+oWgKiIFiZhLylHT2JHyrXJwCE0g5FFHMXPchgTGrn1vfUbCg16Oo2hId0Pqvn3JdcVitBcBnqsQ
hOI3OEW9+15TT6VEClouC7gfwOpZe/PClmwGH4quSY3Tuzgmy5Xr7ZXQBB8FewWfzFb1yZpSxw1F
h9T4tlHLBPrYVr7V5x+lyjaN0VUDMovH1m4lbjNCrvTMdIS10foYMZ1NCXtJJJWYuFmyBW/eEUtK
W01OYmaRI/bPwoE8Z4JU0jdG2Gjd1WLxSRMhf0Z857kB56zo/5atOi33D+wDknqPy4N5+9h3stg2
LV3Y1Nv2GmkITDQAMbrJ5GkCjb0bfv7k+quc2xxDhUfX2auo2WcD7xW/ok6f5DEmSzGTOUpKrqNk
b2d81qb3dabMMmRLlFjFcP84i5TYdb62I8Z5mAkBvHGV3UFP7GFJf6eDn3otr6cFpwubWLWuqqY5
w7qtmGAYKdhbuFdTDMetDVvLXE56KMXED8PRxDxb0S1/CLVi/GtjTPA1eWyfz5nKp5T6Rs9FpacI
9gzh0N38IkzehcM6FC0W6Jx02p4CaOVQjIFyuKrcWHn/k7oufB9a2PBzqoBdtWEGwG1WhdZ+aY1R
GTqsG8dwqN6SrdBtuZB8j7Nqyz8teds7oQhEmfOgO8Xvisv8I61oXIMrdsTBpITyaspLwpTkqxXA
vfSkeji1aqnF86LC1nbeE4bGwlcfLoldWNblnHsllFgoqzppv4Cr3Ca5v2lbreSfTOEkiRXqlsr6
bH3fv4euf8RW70mV0MXNwV3xXrdL0aBXJSjp+eZg9IjxS5xxKQ2Qtp0BIB+HNT5iOhQXhQIvkmQ4
kSG8kR+z0/xn+akLfMfqHWd+xElj4Rhi39SThOqDDv6W/BMiH/XEUffXVJNl7bPLhXCYEvlHp7Im
7m3WW/macRcPR0BDmQhK1SQBd9lmuvhCS97SM4gznW75TQds9yRKmFkbI2wbtlEKXGAYt2mtYI5I
1Z40d3nDqltcP/vsWy9tCIb2CZ1PZ4JhfAqI4EuabTjBK1KYHOI7wCk0XzZxVDTI8YcB4XAP0SbD
u4DDYOFHlgsX3WpFPnkyklBTkCjMIk+ymoMT8XrFdZhPPe/7KrD4E/TmlwMj1p0pmFxmg5N2hOEF
rpnyDBIbW25B//WwIjsu8dh2pGMIXGEytr3yWBhIqNsO5wJOKjez+RY3eFeQe5I832RiKY+zZHTH
HqBlIr1LR+gUvtDdDz+FEy16BA6cqdRfEIRcTXv9DVkyu/NVqAsTKqIVCAFAoZeVaoA9Tp9FDU1i
Is5j4B5RtfgaIlsnimRgEnvjqri2a3XbNrDsLRYLDgnTNvHGxaxuy78IjVlGFoYCeWTq/ki8o9J2
RtuLuJdTG0OvxpxfZLmW29KOD5CFoLvGSQJdQJZSvL7evT+/rSNC110h8rU3+1Xd8vN6Yscu4ea5
U9ryj2PHO1jdKC4zAwUI4Jg9nHzzVvGF0mXRxw0M75mcYTE9LyYEVPSNsTyqCOYRI7tNVz5JwT66
DOiza/LzcFsaDjHTL6UX8O+B5JB05bKim6KxD91QdoTgDZ5aVHm7G1Tv8CjXdYk/Q42vw0DkewOD
Q52LVupwjr86xzZc9M3nua5y+m9Av+EJQac+5lC7MYfRbrb/27vizxlQ6FbGcbKtOxsu0OSBPcfX
R+9k1/L4FtYYSRPywou55y9g3Nru0+knjRujGLK/pCNOuwMzMUvC98e9wRhRDjtEbf6xstGvc401
qA6CRffnPhtKw25tkQMYlDhB1HQ7s2R1JecU1uK2Dy3EtX8Lm8KfpYr5IprGRe76AOtgNdnqfs5V
tMueOkOYTgMCtBNE4ZviKGNG47b4aE1MNrlb21XhYJ4oyKByBMFZFVvLkWIKI00tZtNPxHrFBaTS
u9n/dM29RJCLbqqbUIuYYf5lgiQ3pxcWA7B58FCxUttx+14rROPJGnk/JRta74QxkYXcQxaZyCMU
lOAjueHSJb4z5KxWP7+Ssnsi4TPjBmcT5bo7ohVlBveow7ck5R2kzaqXEqabAenCX0U0v4eK91L7
hSDTroo8FvMokNnWaqGs2VNyhB75rHXuWdV08DwsB8JUmBEIonHxLpjLnJH3V1JpIoL27tUQBrno
TIIhZIWCzkbiS2NR/9drqulOW3tvmDfPMRZHpGnk4wDJYRQiuasuPnL3c2FVi9Wvh6X5ag7gKymo
xaSqjXcIrtvzsjJ1po0FmBR7pIOkG2UnqMDPX6ef6LTpM4ViZJqcdmhDfrJEKp4TUCa+BIIQyX5G
z56lGe3TsSNdoB9S+5hQvnL/ZUjIi2iEUCgDLI5dP35cA0k6Ely7nPRaT2rBUvEASfR/dPF8HPlu
0MkAv8Hbn7oYvEMhsFpDy8ViWVrZYtc42zCOZNiay0HvOTOPURX/F2PN7eOdTmm++8A/lX3ubbt6
mcMD/q+Qn0yoxCF7r/lmIpzq3jgCuovlwj0COqAB6NT7lYKFI/MsrNO5g8lDKhPRsijG8rUub7w/
wcKMiiz55tT481TKk4MtN8/tUnN5l2hDug7NVI5RtLKztxbs0rMbyIks3R1l674bv7RL+QsDBZAz
RQSsIIhbBC/7NKjd7O7suSNa/6Sta7fS2+v69JC8uVHt8nNZ1P1MWMjL+KnPqJEBJgHTQjPlsVu0
EbPtgSZmfoZBCiywllwV/bR+wKP+wv8X+jFPn7NcVnNouaUVCBJVqKjKwGFoKD/+Bu+eNrItxS+1
Z8lZ1tXkYaciJlc+OhSmtTNvSeXcWNtYb42pNXjya3bShdBaI1VMqkZ4qQM4ttkqlHy54to8lBob
JjsoPlRJD3RaYOT+fnQxaO/YbGaYcK3X0R09cUmo9G/s8th8gwT/towjV19Y2I7jK9f/8dst6DkW
+LWRdeFW7xoFGsTh6lxVfve4Wbdte0h/+oVX4/+JdgMwlmmu/MzVUuj5x5VaTB447K3sfIRppe2E
equXeIFiSddQxTiCffkMeFwdFvQRFu0qWBI4WuEJq9G4vLjoUqafq8pnWCylu7jJDtkcafVVDQ66
l1mxij1+a0aIiJdIAEkS2AJN8nQrNXUloVDCcykIFqnALMhVHoYSvWbuwHhCkMvn9vX4kiwWq7Hg
s7AZ1NVkiDMXeXPYfj3NMNdQq4dBl5P0hcZrNe0+bQxAh8pZXhIeKLI4YGo30jmnSpgbVzOXvxAt
bkjiMPlqqzmB/2maiNVhhqUtS63A0if6NepxxoyE82I2gvKVEd4CBnhZ14sDE8kfiRxNxo8puU7h
RPOl3ZFNh3rgjhcnjpZrALcC8HN3uPEbL7jK+d/T1RqUEhSFxMQh3vl3hmsRgmXwiCJ8RNDXQWOs
zLFFxy/82k6USjMlxdPt9kirHoSaSZlr7Bx2+XhjSrpZkdxenPJIbxZOuPSQciN9qLcrHYWWuQ0z
VupCLVNjaTYdiZwNs+qO0drz7kOTTAf2JepmOUYWdiypEjyUOTitG7/fgbUJtch6Z3M1lZON//CI
5ag37a5MHNV2zLw8n1gB3uNO+HvuRoxLQkMjt76vEaa3hjvkrhNYALRIAf7TQ9w7Mk/b9AzPmiE8
GMdDq42XHfOdmZcj1IEsMZjj3PosO43tcwuvFce3EBBEq/mOB0S4f+f5ANUnUx1kvxSRoUG4xEzM
CMLTLQvhlANDD9HInMY3A8+EjKhU4rTjNLkfQGEtRI52ojVvAUqwkztoXqzWX868nNPZb0BHcIOF
lQQPF+FLW/SDT/iMABL6KHSZ1wFOKYpLcLcU0/Hxv2UP0coqhyP/HfZM3e1e+gWXfXcJQMgvUJ3d
8/ilddoP/czJK3+FdPdZ2GjJ7uSY892IN4JMjuVi63c7c6LuyYpOTpBI7iPWpFwIgqjczndRWW2h
AsTEXWru92ASOxI/202uXgLG8QjGF2Ltx3Hcvq4HqkKID7q8TCafOexpNVRmZmxlZnCCDaCy+8b+
w3W1bTfd9tBt0XUhTRSI0JNsl7YOHF9bk67tHm+xrsXHrMq7fXHhr0Sm6sjLH9e8uGQDIebgTFOP
qYibM7fdTY/7NS5f0Da48US7Qa9Z6qa6U6w2YUy9z/UM02sr1ZnEIYnt512I7E2U1p9LfQpn4FGY
0IF3Y3y8Yf7H6g8VtRh0L43mMqFdSITE5tVv3+jkSQbANWABSneISAVbC+h7BcbK5ULax0JNbpZ1
rRnPuVnMst7hSGb82KkV4HiyX7FMkTG+YU5seGhlkJmo1siBXmJ5FQnjfb0A3vy/fkoAF0EmKcPk
RQhCm3o+ZxDCvZ+97j1paa361KOMYBxhuJWV0/6mQMKTJsPfyqg0tN+yjxyt3tk4EX3rCHo4o8B7
bhO/XHFBlKyB3l1j4Vcf2NNG945eFqGE3KOHvLXxG+cekKZLReCPFKtKl8Yi7otKaK6513BHcNbO
t0OncVzLndCB+clT24NqQVUbWkCl8Tq5R5MSmDD13BRRz5iU9PkkQne1RPP7SdzN0zgFpWqpYnzW
0Ktm7k9JwAqBhanniDtyjYBW7MBfzww36a9u8aOI8NCtdWDwzfEFSLD/tFveW7EyjKFKY14pptYl
czbjaaT4GJzSZd/Uc+s/p+jZRGwpgScOKYgQb0+2fRVxtqu1EI8bYNWtITUtEex7lqC4x0LE9LIA
3fY9qA+vAAwxNaaHjQxfIT5SudHogVaFFLJS0/aBFBydRhHjHALn2SG5aNWuH0Pm1U+VlPljCfRj
bwPbhTLd4uGCXqSfnnm0Xw9a8TUNXVAs7t2zAd5w7KQli3hU8MC/x4mi9njF+r/WPnbvKShwuBH2
uPfUQYZyKIWxXESBYP0eyXRRYYLXelVfVn4O41mR24Q1Xhy/rhpRvZswfaZh7dwaeD+i00l09ip0
VI+QztvokXHRf8a0p3C9xIrj71LZSSSZ88AaZ7MQKvztq61VeR14+mFuwgaTuY77FRKKmC8FxaTU
P769QqHqzGEeytyZZIyfN4DqalJitkX3RJO3qX1LlFgABKUD9wvJGK7oYnN5pssajoLjCCDdt2KB
335BymlPNRiOTjSpEZIzg7r79AA+KO0V08B2303Kg+1AAi7uBiE6iE7XBZqBVrOHWepqwvNxM5fp
xhVkrsq/kc1YcKTXNYwtU5D4gV82vKh0d5r5h96g4/zO23ntsx7pT2KhGKbn6Fy+0nRYtnzYs9VL
RCiOoXEQQwETWZ5+ML+uUtR8GAKIVrrI1Hcy2a+JwSRweo01NrtoR8KYGZXxuSuH4Z+rfIMGEPel
YdjlDHoycy6EXkUx0+/EC9TetkD0c7equ/WYTnokoWhT+wiy6g8QnTiMUFaJmso5uNG37NzFaZfL
XhrtgEg9cfAqd8kfV3C10rnWgL1nx6TTEUCpT4nqps0JHigstgxZJTOlnQ9CqKiYqLMf3VwNQnsl
GTNQOwkOBU2ZTAn5/GkcHWwr5pXA0o+EBnWCNsl0wcQSneBUcnv1mSIK3iiAqkFeGF3Hibatv8pn
6xRm9wyoUgX6kPpmzDbWlgZkmLEwSnlPK+qcUmJxgl0ROaMPMIvijt8T3LeH7eoRUpsK5LwrddFE
H7L7UlUWyn1nUtSW6C74DxZe4rx/7wLDD7kxcEeoWFKPFrXFA5UVjkrg6ybd451TeHFrg0p2Idyl
7JaHM5woVt7WRem5sy+POF/L+6Ki6d9dBfmnZhkAT1gb+tBAu1pkK2OMlT6RFXPWPgHYsRZG6ozk
0iXGscsBpSeAY07js9Wx7GuSad3tK4+X8owDScuOgmAF30DMF/n+8MQBHi/n/786XL4pNVgJ2qgM
UxRJ90RKfE9WCSVZn7jN+4hcnzjma3hlfbVqco62X/7vKwoEG8FbVoVxTxIfQvT0Q0NBOm6C5yI7
i0uHTlS0Xbchqxpr0b6YttwPafiY+lEHlhVNUO0tyiXYYrAeRjPNC7/mgBSGozDPTT8n4yAAfny/
RtNkqTr2A+vYiKyqVA/tC026aFk5QTS2XCCd+D2MzzuAB6GwztW8YKYhO+e7VYxUQbxHPLr5FvXx
iP4Ue937Xxl/Zmr01SyO31T4B6cpvZNjOfCWw50jyxRZxpZA4S7muxV1dlXldYCq50rMvUAq9zrZ
O26UF4aQxZeWcLw7yCDIOewaaTL3TnCKaptwcPNUiILbwruXJtxAqeEndF8c5P3IRlXCmuPV459O
E4fJKe2nyefIpTl02KcEzdmMSNXTmC0Ychc7hNMfadTUdUlWN4sYhryf80KDwArOCPbbVOQtaz+5
jg0oHmrGuO0grbgUBD1xZ2IjHCfSrprRdnTXDn+cNEwNRcp/YTWLQ1V8zva5+xZD9vFDD+bxgs/0
1KxuJOuHBoFvbnPCkTsj4FhE+ai3OwGTxWToekz+DWnHozIZ/LxV4FEhYaQR7aa6JeetrojC3SO1
6mf/KGrapAWv8nEJ3yAaJfRYkAWTbl/A8Dan8gxw36efgqlKw3BZYh+33PepacJ+tDVhz/gmem+N
h3SRdHoa1AYR92Q+93IZwTsXeuuF90cLiAmlBXAWcBLieDnsXWsNxXw6WCsxNMl6eLJj2W5piz3t
sFeRh+vUgTNrTbABUuvF11ltCcXslD6aXX3dXKW3LvrURKe9SVXjDRNLvw6cZLNqivaNDDYJhcfV
LsawsxilYB5qGbyakZhzC5cKJ91143e8osl1dAppFfR4/zOabhjL0JOvm4aF+VmYepISsSFyErdE
f6uIi9wuTYVKISaM1TzJ9cNGUYg1Zm7HyMJbfW+p6N0BbB3T8ZSwdL5r1e4LcrD5SPU9b9T+w/e4
u/4VGEH0cXyYue1VtcepVQ7jtud+BkwilMqUQuC239q/Q9g8L8Wrf8Vj0R0WeiR4yV0+S78BVnZC
Cx4pNylY1+wATnF9dssAz9mSugWAIxKkiXIJNK4yOSXYQQ85bDJckHJWW1J+Y80MwIMtORqI4GQW
Yruo3fHo3z/qxpZ7OmgC+B121TiyQDw6dp+/HLuFTYvj3IBaoucI7SCUB4q4jUDZni+n/5ZLa6i4
YxlPOI9L+46MM8i5RoNetNFnrY357WRf32k6UL+M7xiifg/Ia6My54Vb7w0YZ2ClmwTaztpN7Ufj
CD66/k03Sc0Tg+uCW5g4OyBnc9Gxk8j6+bsfPXuygJzi4FrowOaFtiCCT6IiOnYTHU8fkrTbtCLB
fEo9OzAsEVogzifCjIPtYZ59zXh3Ngk0LFYcB1XiqiEnsY2e9GWmL04XXwJG7anyFB6TS5mwpIr9
HH1LnturU+395RV7jRrBz15QQn+2RJTrn7z6R/DJu5QIw8L0he03/EhFFfDVwx1bS/u3nfCH6AxS
tO4bUzDSyfn5JANZkVtqXtotOYYpUXGfX8oz+F4LLO4x1K4n7d8zaq+XusLdDDKvryL+/sHV5QNi
RHAkOPtJp6kqhtg78p01ME/AqCvQvIbK1TdjSy5AvPueXFdPqJrhkERk9nl1LUzVGqvi2LEwmHnL
YvSQqtBczAtYovN43QZOM5iXI+UuBixMjkU9Vf9l9ftMNFuuY8Cql1Bs1Zf5wwbIOnifGGmB8buJ
gs2GDSyTLuztZenlqtYJaFgejeCPQrelGnAalFwChRJQfmnSEhBFErCgGZ90L/+rFz4/uIOKoa8B
4hCxj7baWH3/3kyB6RzNW3NcyP1AW+6InG88EFcuHKs62X6FLBxqzwa9Mq2q9f/OW5ZaKFz64CuQ
GOuPKnQlsXRn8Qe3ZKMLxiHUm72ik7R+7/VQ46n3Rq/NhAAInh3ZjdvXvP1twl1Q+Qa+2hpUc9dP
CTu+4RoYM4KUcYvbiEQCGOoM1aENtViRoJd/YugfpocoHaQVWWC4K1WFw7rZTc5d6nEwLC5P5Cfc
1wyzBQftBMJtY8vWTCv7Hi42F49bF0DG4m9hkwM4xG9nanMRKEi5HIKDSCWSV3FN3HFbEasdmXjG
9yxJHhO/RCpUn3lUXYBWzd/XfR+Std3mCPOSXsZYknY1deUhP3SGYWwfyqrPRZZ4d0S2cE5hS2qY
aTChvPnA2eLd1l9q1hgXhKQfkwe+2IBuQ5cLoBBRszqo7vyLQkUHOamQity3I0gAT7r4ggFwzfuv
TnPZVaAkCgLiyIV3n1lI1e2ZDLda84TJhC70xSzBa+0K0m3evk6dNxGctWK6yd9HO2HOW7XmFF2i
C1oSVey2eb3h4xEkpy0NNOsdpC5pqrb9rx6i0pBk7x/GCtHDTbCbMdfXcHC9ctg3deDqwiV4Dt+w
N8s8pIYykhMk0YSXBioYTlUzGTFXGBe7WiHN4rBATul8uSlfqNeUUmBHpGfAaIlZo+ei4UnyzeZq
8v+HjbWlua3gOGYWtYi4wuguOfvsT1c3j1ScV7va0ruRAMLnqcTflhZAleRWqTTh0Fv/z0AgzWwL
uDIhWBAV7eVAJoyhhtp5UxXXDj6udhtPxxJkBAWmi+73id+pkIHu8f1qNgxPlZGOZE/RozMOehua
+5nX2AUwBzCImeMKgbnnVRatpr0geDsmT0sYbM79n4/EmdPnPtBJPp+7zSSnM3YRwIXs1WSseFfq
kfoZqP0XrZ/Xhv1QoVAqlyQkCI2v+RyOeb0s1WDQDq7DUs/+PujlnRQrjZjd0dvigwL9+6PTEN+T
NYCRzkii/nJwgKfz46cTyyJQqW++Q5uUvHIfJ4OVWr+USZyZT5e8xg9buJpRLVOLCpAnUy68wYDF
d9HibEPUmlBI8SGw5zw2VGfd0kXjm8jLl7ax6+KdzdWrOQTd3d+zFW7N2QwTPh4hw6juVr85S6BQ
hy6uoT8/bZpktj8xChgpfGM2uhDyZl9Irdk9LpQ367JZHTWr/MONvSXfPbOMAB1RdKmpxIWhOutJ
RKkIVS73aDJgn/BVNXCXXhMb2Kjb0SMryghz+1Z5+6CjOEpKjpso/uhga8ODbV2d+ZJmt7J/DFHI
emlAZR512uue3ejngxoKtk0w/248zDY4XZINulZpYm/cozFSmx0l9T4HKiVZWlKOIZwo7Rk5aX0M
KFAdlOUAyXELOSPB7S6ZUWBAi7J0RxTYxPU1OkhvFlhG0l7q29hlo6UTMEHJZzS+B5KY1EcphENG
78IobI2FTSEYA6qtb6alFJHG2MGZY9SNe06W/OT8hO8VgNAAcALIzPJYNpokuyyWW5OFufbE9G4E
Dyo9p1r+1mV0SKg3HVz2PqzkdywxQTUE6ndzfu9WpNz+9G4/SI/RVUCdGIORTpOOiG7sujs5VYPW
trQi82Q5j4GOml0NSqjTA3jY1sb2syq0uqz9+wnZHxVM4GQWSXiDYGon6UG0/3IjyuopygHByNVB
sM6uN+GXrukQm3Fkgj+XbEw9sfxom8QIr/RG8QbOPm+tnlO/BUe9wRkhp6XFOrGtSlWo7UHJAnBN
TS7nK3KLrXwJHApJAgW5kjB9mI4yClPjstyUrI7MvbC4mGQAuKqay/XtYhU7xhPylvfLaqWWXW/X
N5ZD2kkEYEVL3lnty4KYSNA07rQNbExF5u8B58An3kgOYFyqOG8/Au/hC8lthCvWiDWX8N/4EO+k
CEnz+hiN/63ZWsrEh8fHA5TRTGBJ0/FoD9PGQJ+bULNAIL5vle/n6MALPdLG1IWje5dmvcWNS/A9
cWcaEXvJBFqNR3LEEUGyjjay2uM0TMRy8wVI3FdBjBuvX6OnBcEahhRYXqpS2D7n4ze3n1agdO5q
2mYHkcmRejlmwGWgtCkMox+Cz9qfMYFhgYIerTmTnqOREqZmwvdqyGobwqbm39zXicNmWlP5PM2o
VL3RAdrHVWotEI8ZWwF9IHv3+B6IWOqGQMq+SOoxWZrOXKRluONZym7Jl+AI87h7DRKYI00XiFYk
d4mjvP1GlpGsnN1iFrhzk2dCe7ynbUVAIJgn3EVRteoEkWh6mLM7W5Y7gbgbSTZtDbfKDBKgpapk
RIk6v23HGN0MTVBQ5Z4ubtZQsjqS8hGpUwuQibbjy29qJnwflAY0Fn4eWDmdqTHvVRfwcn3yVkfO
O+hpIbJFomWojbCKZbPDM1k+fRxpCWSGq34NqJj6CgDdyuIsdc2YSjCugd62NM2hlJfWKUwAdEMz
h0t1VpAHsiyDH467pvc2IgeJORZVIdugCM4TxYpwnTzqbQdEkz1s3DyBTcxiBoV0GlWabilYZ90M
uywg3+tKpMhc+DuJvQBHquUdMlPYJcCjW9LHlsxs6ev1ZI6c1tyQq2P8o8gnejr46oiBPw9XJR05
jMWVno1bwox9hjAkF+RhfeYwcSSLsKAAowp6J3dJTzhfdxU6JiaygRUNxsFaL/VYXWnaNZy+d1DK
cBwZRoj2D0I/yGqTE56g0Z7GGHrUrOaSl1Y1krYevFZVQW/GnS0vi+Beu8We6DVBnvsy7wrm+Uoy
C03dvfrUP00oq7fuL6VSXNwyFajN74fts7/YnSP5EW5xiKxhpDtcby2yMa/uQzCMJxTaIf6U7EoJ
3TKr85ffTaJaFSm12/Kr98txBuSq2BYtR8ywJm5VnPynS/JKD02DubaPszGCnDqAKT0TB9F8zmfc
fbcRAoPDeFEy+lUWV8c+ll98r8njoVICe+HD3mamr8+i/CyWtJ2KnvhhvynO5dgjsxoliG5gEAdQ
XI6qWG4G3QUUJO72aAot4KPAllcGQHv6dT41cFKGOMNVqiTLeSlsnrpu7qXpgsbOVfiRwAIi57+p
JASXT89RphcTKMS3e6BQiK7wucuWV/D9T6mkINkOQqdBELfpUaSgaPMfaGTbY8ZADOuJYklegVSF
06Lii3z2m6wECdarlR0uUI4WvuLFr8f7TYoh4sn2qOmWT2bfH/pO5r7Fi6vBp1HL/qTufOu9640k
ShGGFJRPox8doNPwDDyJAMHMDwxK0SyaExGXeyu993fmTmnPHxIX+hCMWB/FjIk5AT/ZnvDN29dq
bESooP96xhmssd26VTuC0h/NUXhbVUL5Kq19Dl0VvRLp31OW4HGBHUzi/ZRIyvnaZ5qr3uqXwI6n
wem+919M2tW73HtYL6g2WLZBOSpMxpx9oITsTM7k0DarXP4dPl+jMvwWseaMBVh8MBvSog0f77Xu
szZy8KfrjgKcSRhUU2jeFkwe/mtA8sDryi9LM5R65+G81ZC07gmEsNRK2aD1604ykI9sljiDEhD8
N/edBglLT8P/8+Oai+1Hh1Vc9TBLOGEvZirpeOQ/05KzuFsuFlTRIPRM1bfLTIf7eYVTD/jp9exu
Eclq4odpEn19jSPvqldmKgmobCmXBaRp1PWjR3mvv/EajhO/BubZ+8dkuCVY7+TBirqv7DkkKz2P
whMbSADYbklmgRm3pecm2pEdzUFyLJRYKvIyhfg9da1/rHHF+YthQPCBLXbPFban+tC5PJk2NZ5l
WEnWEyLMQr6154hrkcG7IEkDIw3m/tuQwtAzonlS7hLR/piqRasbRPsUKtvGF53Avca16uMca4AL
gKRyYnUy67h2e/ga59ohaxcu7KLQypDFLVA78ccxrJL5V63rbcxSAsBbsFdTLaM4JAZiolFgBTT9
8uJgIzzHeXtYsYfVm8B7uWK28PjFGZcTQ07TwGXoPiEogwkzf/U/TgeUPBNRuBnYuE1Q1NvoPQmh
l8ukdWmVsGBlecUTHI9/0TWb3K5dNvBNyg/wyrrldG9XpAXqPyMLstyzPEbZtOuDFDrWT8EhOTY7
ZSwaS7Nvpax/Q3pqoVzWjKteLTs7+DrbRpCXc+7wSvUUpMBtSeqF9cjUFkWkesRLfENjs1iSRu+2
7qBtfcMPDkhox7aWeGs5Oz50RTwbrpdcsTrjiM/7iEExdBU3ujvgAR/SFOujEPnb6HZGOGnjWNa7
7MJvnK6WXq73xzpY1R+lmLxAIfNmduO/1N08HuOwAqRFkE8r/1+lFrzTI7sSVNEbQBYsUfP0Nl8J
vRHTJ5jxQvGeoIGB4Wv9oab5yPbjj9oZMK/IKFyrE3ScuKaKFfICuKNo3U6PgJtzfNDdjD6UaeIn
kzoXsR65lOR/gYGKlc+9moVuRxQyCd0I6ALKczdEe+jzZ45yhu6dnMtEZg+AjOsaPDGrCm4v2r/X
aggO9ngdDoTJcMSH54Kn3ff0/ZJiD6v9BfH0BEu2CnwpKzAhqHNoP3P1ZcGD1pl26Nqcos/3ih+Z
42tQ5pJ9olpwTe7Q+fsOnXVrG97ESSXsHwC1zG7RuGYd2EDhIeAeMzuJ3+J2y0ehldTeyIOmzSO7
UaGk4VI+yLmpJOJLuwQecE9lGbbUdXpZtIzX6Fs/gZnZGEDMSmE69NaQtKQG3nXgq2jAwpt9Bs3l
eKvex1nQwsdeWbw05OkwKFadm4PeGnA1M4ONkYtjnPinK4m02RlN0spaHFitWpXHpPVVPDwRyDl3
CyGKuTn2bChAQfsfN9Aihp+JEXyXyHHN0RMljpEm2MlwjwlQThJcPgxmsUAY+en0fXs9jeCBIyW8
EZWsN8kVlRdsOF1vnab0ZdkCofyWStMHuoeItsMK+WsZVAejZZqNRkSWz+z9ittdCtN/X/T3ApBw
H3/p3Y4dXBo9kGhCPRB+oqD7POwOXbIKGaXSu95cMNzynSDR6HK13W93eoynxLZJFZEKfZstSMAm
SyqbLnI1BVBJgbtw7Tiy2XjIfJUjoPk+wgwfw4XaA8/Yk6BJDJs6tEbqGvC2JeIMwAetx7Efz2MB
TTZ/+//DlSjNNjyz58GsgNAw++V/dAoBKZwEGeobGvMX7cbzQT42EKrBA9sGQJKh1Wq4oa6l81N1
1RTczBoS0cCiuYO9H07Vhrf9E9OCIBoWTovdSoQ3N4IgmnkO3ZC6BkIagRx9xoiREz7HTeiork6r
/Wyll7NAyJvxYt75JBcywditdw4xHOUJ+pMZ56H+kkgkWwoCT3D5p9cN+KdthGWcNDS/KrYDXwz8
Ux1J2zLnBSBYCDbEkALfiLi/fvg9s+hazIPLG0WQHra+q/e+7EHGn3RlvZSyNamTlSAHYtqkN9wY
1hVZr45AMG9zXfI9AcDvkwnsCMAqk4O/YF8W4kWC9FtAVnWYu1L2IWkUN9hZPUWSvitATTI+4Mgr
V3lMD2GeK0KoNslGO3/kre4nbFLTbu1W3SYESxc4qSkTEnWSd6otfNUBmlpF2qQfNJN297ywJuyl
dEbJNJS1bJzdzb62SCbopUt2zX9GCzRby/7A3KMv9CAnbXcW4Ymia4o7+jl6TDk6LhAaDL/rzr52
8vMFD1cqpy7vZWm4FRsu0HogRU1m0XiwReN8VgOxDugTmu7rFRs2aORqzmkR3qWdVMq561wo4ioL
phXZSdbl7h9kxyt9rGKrgosN3ZOsWSwXU/JwRSQ2VV8wvMSIkCO1ArOWh6zWEdWSSuEupJog7Ktk
ZvmjEYnx5UhQRLPleOGBQA037FMAxV6nv+S76GH0c8taN4CTGWCOpre+vrVYjO51Jf+Oxdwz+X4K
nQ9dx9efurj5Ghi0hwikOXqvowFV5IeYfr304mARE0kzB+yrUC8eC57QhApuMunHELwGMQxCbpcf
2605vks0sH1IZQRJa9Gxm9q6jRPjrYLlBFaaprkmZvvOZAN4tazD/BT5OqwBlvvedxfCZVGekGq7
1jeiYpnXo7ugKHSV6f+V4tlyMr8zyr9Svbzt06dT7U9RTQhCgmScleFG4wvOXCw5Zb5d060Zdshg
4RW1KCSTfoYQ+2+iBF/37KSyJqqLkh+EwWol2Ml35jmrrZ1iEt0zbShK42LM1Mh35GHvRCzhKeOo
XxZ18jVVuPo/UIRpQ+RJbYbivnz67a2uKIolMcsJKFRV2ljDeadcS+0yUIyLVCECKAg0nho1evPM
aV6XeQoRxotWROmDVu8t1Bi8HlN9JBKg5JlP3I6NBemXiUrLP+ObsF5RNjtLY7GbXGXxjMK8mYy0
7QJteASawgQm5Mr2SAHo7p537k9sVLoHh+qygQiFiNoJX8skFm4WjCir6Ta0HqU57k9CzFu12KkL
nZrqvy3OGEIhQ2dlQDTbhQq7/ZYgMeIjiRejjVIePARw25cnoe0JQENF5VKju9HUcPJI6PxKcbU0
eOn/68OZS5cJ21/qgv8t2hlYZb2A/bQ1oZiKAPDVfzO5wnuM+Wdu382Wvsvvq9qOChZ/jeTpBU6k
P7BI05R4yRTBoAPmWWcV5JSmMhzsLyaYcFMcGS4fQ8KgHfxSoxeylww6ubjdLUCB5iFWSVdsBOBx
/HNAiLU25FAGKqRN06X/+/PYjAFMtAVotlBIL3/UHgXvZ3i+fV/OR+14g09CU9qDozeqSc1Rb7Iy
S7+hjWB9Xl9XVZXt7ST6Th1NW6crkm/jics1yg55LggcsTgzI64Xfz3vf/RtZ6jFMT+1MPP3Bnwh
Ny9f8K7VAGASE8nGGiTNJiTSDaEYh34YpYqxp4SIj4df8qdZQ3fvLe6hwqpyfx5S/bd+FD/hdb9B
jYnwnozyoJmjjWgk4FgyEZMAgmFrlny6iAzGtPqELC0g01ARK0MnmUdf+hPut8zb/T08l5GgULpt
XcTHqC/K1Jye823gAQRCOxZBzBzZVDbLEFdQenFB1dUaQRhFIF89Ceoeqp01DJXxpz25FLJHyD+Z
nW5s9iOVONIfDggsWAdodJmlfd1ISTxfhphKsSLrp6pSwHu58XDpcDyu1KrwuE59nLiQWGB+zPHh
WbiaPBkek8VdzBNoOFap6m8SXw98NFoOl3VDwm8F/mQ/f2hVSLtTLl1EH1p7EkrlnK1c+Z3Pqjz1
AhSCgv9xvfQQ5kin4bY3uNqg2nkMgqOetyRvic+CM4J7ZKRxm8qp1GIyG2UyqUNid1hYytPzU0Qv
v+W39CDXsMMy5GdVaqS73PGs8hSXbbSb44otT+z96VDYxECQsrMrqT/Jvv5I6xY215qluI3n9HrR
iX0ylMLRqQRHt1+Sas721rfI8IffYQ366+uYTVGLcUQ/aBjkjWudLTHWD8MsaCeltFb/nIw7UdPW
U9t8mr2f8w+snAWHx6ijPIJ1898F+SAQQNUyHCRFSPAWJxq/WrkhvAmkwbKmNp56+9RLbTEkB0FM
BmzJAla8GQDsJgYL5gwGq0n8J61nUr6N8zHes0K2grYVBCN3oV94thInwem/ajQ+aqb+B7PUyqcC
OovIDNz4x4Fv+Ffgul6NwWy/ZJXZx/VFoU4he4F10F4G1bMW/t+IzeOBV+QJLS57V0j9mcJyplhD
ahUTSlOl9pWkIBLqFXKQextqCV71n7UfdGIQF1iqjMjdRIYvbD8h6R4q6nXSmBw7+tgeuIMkJSGN
19NMsS+wa9ZwlUjLYytVu0i4aO4z19lJi1zzfcoI0ya5ZH1W3sOrNVeu3gbI5GxHvQTvhnTH9Gop
y0b76FqKbIP2TNMW3G2kiPmE2uvPdUUeGjCl9dIqaK5blTqTXDkK85knl5T4MxPT67pyHrKC5g9l
MoLl3/RB76NGQYTbP+CHEd448nxia9hpMDob+plvpsTHhbca8M/WVD8EDm3b+Lw/d7vCT0cz4nKx
wM4AZg7lpiWB1vr6Cy2HoWLeq/z1qdZ6yFq5HSopaKhNIyrQJ8a6W5zIwVv475JOM9/1M0sFszLd
GCMY2Ss+YX+Rqn6X3ylfMAr2ggXPAkumOjlVqDfqTsln5rn/P24VQS5y85wMleiKwNLwX5X9eVoJ
l+145QorU9bhAG0p0DR2fBQFMt7VIlVrls/ATpHml6s2hQNAZ3dUqVQFTHTiMfYvyOcWwvzqV69N
CB/b9F5+cakZ8C69EtHjiEBXEpOMqD7751QAwi1/pnkQRCKuTFjqh9oYWTsILpLRJEPeXLWKmQtv
t65+6UwV4b6cb6q+IwXdbnauTkmOJTE6Zx5tZw92zdg88C/RG2h0/7XIwSyBbDq0uuz9e6G7JiEw
mSYOEtQOSNg0j+zcr+AkH4A7pJ50wXqi1KO5M0WU1/NAqKyeHisiZP4x+RClFPxZXmXcufNjSoqh
WHXAuf3Ky2Yjo/Iv3TQUvtP7zRs1/TJXTcXsOgXaofO9KerZ4td9NU6/5GI9f3IaD3lENDEiCS6z
La/uWDXyALWbbDDqJ/zg02notaZBR+2oC5kZSic5m7Kv9Tv5kgLiqPcQBBap0CUdeF9hLse00cjA
X3Uc8OoyaZYYxveamUkd779FJmFlGL0GMniPC6Hdwrk0fnyN62lC6steyKHMS9ys6lbWbr26etdb
6buNSQZBikeVpY8Sy+zheyaGXYtgvr3BRHdMRWaea6y3tWZfu58sGVUBLIVhr5wZv5Rk/oCFA0Ro
uI8rF7DnG8IrqafhWNpsBnrZc8a+b3RntMnN7X5uKYEjGwpIqPD9xKp538MTjjEGZ6Ea50GQpp1F
mMxUdmF/p/uP9NqE5JCRokYMYn24IhpireOJSlWh0X6Sl7XnmNtLAr5fI7BDkyao/DQxbpUFA79v
N38uvoJFuIXsGiAt0tJ8O9bQE0vFADW6npbZ3syJWyhqzxeAMlkMBe9dt5R1YXwMYgaBmwjPooR7
TTPcOfI7WXluhd/Q6DccN+F67hYwLMmBL2g5zwJvUrckzVqJIxBNkrLGjBGgQ1GeV91LZ06pp9Bg
HF5j85jBf/Pl32CtYCzPThQUvxjaxJruqPR2GVnIgTzL3YsIUYz5RhHv41mmLfjOgojvoCz+cRaH
d8rlOhZPlaWOrSTaZB0p1dBdAEZXs1akXJC03NdRpOZIBnkKS/SDdon3kjL/C5NhfUzoo/e4jYI1
lwQLcG68mAtfAIuvRJwpwxMQS9IWQJmhE/bSvakc9G2AwijUNTJPe3NDHB5lYdxEl44lnWMLuoT+
0J8cBk+fpM0QVxJx0mrKMB8lcegpcCyKW7/g6Culyk9ZSAu3fGme2cjElysEdVcXCFk8KtnlfxJ0
exsudsYiRqwweWx8bcHiseCpy7vlsnVUFdV6fa+QKKcWBcFmppfA53PHaufIxy3xWVHloiMbNlMg
LqiiewUD9xUXxkIwrP0RDPBSCk4OTFtFqDiBcp5q2Yo1j6vLgRVBXnX8Gim6ncILRfnLQC/Oh2Vo
NWmv1Fn/LoIr5zvD1H676Z4F1N2o6m9GAAMqJbjqyZWHicEVuVRvWBSPXj7oO0ryeMIT1BUzTOsu
TK3HPpGr5M/fdWSkRMt37S4wDkv34/+33Q2B1EVdmc9oKFKIcEl3IyYxaCn8xOoKETOxZtN+I0jH
Bwf8yCBFcdr1iOOFS0zI+AviDyKVKMu5IEQ3E8bGSIxn0tQ6XOI1WShNIRcwapG0wer5LmoKOOdJ
zyuhlMOoB/Kh5/orxu+9/CCb+8D9MnLN/lutRy/JWOZlxf2gi8tSkjtAChvsM9XHhdCpcPBS8TRE
w68Wg6/f2ucGNFpys7kMDZsabnUmRfB8NdwMMxMwP0nMlR48Avh/12EWk6GyhVbTn+JfqCB6QNqo
xPilngu8BbdoYAvCz3K7NUs4zUjk0Tas4s0a4dNstNUKdgHuqBFi7v7kpK/dwp8qvXuXB5LxZjO3
xFVTjb3UxRBPE9M9vrA+1g+kAjFxVbEZx8uQImglzGVWxmayefmavQIFkJF2rYKkNhAQJtjTJUiP
0Zlg/PeLcHM5sfaTMBxD2iOVNdpuXhQvj71uH1PAx4WfZ8f3xYcZBmcvEiQemIrtpkhGdMWkLfHJ
k10VLODl1nJ8aDprNbDseFxVkSyz6nu5gDp/ZHNIHYUOGQCF9BvDEnJJwf9ybL8WmVBkjopR0Sm3
LWepc2jrTQBJ2vTkAmLtr1jfq8RQAibJ1NZYtlcLp2YW/1eIaqJyqH67hRA0mFlsCVzC2ubbFhap
2zweDXcObAqvt+wtvg4FS+0sMtF3NOFBCPqLHVitvkPoUkO2o5qlN4RbYyPuZmxP08oIFSfh9yCr
OFTZhtj6doCfy2QVQJiUc5YqxDgGhE3vg36YpSqaZMxhOhjWCOhGYyIBH00TPR37Xj6UwKEse05i
RJdZ0WJjn2qRypg3+fPXejlorS+VHIzm1ibFwjVTvBHe2sglJ1qubaK2xys+ToesH0P3uJvfA1SP
MmKLQ+9KLHfsdRPtSMCHgvbzhnyQi7c8Fl32cupQY2t87on5MBkphqtbmy6DjHVPdGUNjvsQHVT1
eLRJZz8OQCJDGbmSPkmUCf1+lxg7HIcZlWIFe5lME5tzXqv1QYXv1MUe/j0KiX3msjdYpR2j6u3s
y2FKg4RnkSSP78qx3WOVAIrGcAZMadsBhtoBilmzFxcWwRPpG6+bUg4fFvTHa4+gkxK8khFX9TWB
bxQ2SKW3eRTfLv7DpnV7jsz1pDrCM42fv0rKZdj+xVaHahyWi87/GLHRYEnIuyRMeezssRq39ehv
MI/eKm3cENpNrkqkSIZrgZGmXjTAhh3S6wlBdf5wENZYoDctN3UeC1HS338urgQiz6/XBKgU0UKt
GAZZ5+VbX3ZsvrVOjn7E5uxE4xs2bI3HPGs2pmzvUbj2wbUBO3rvK8QbEMgRRTjWqSOVHvD2CKjg
FuqsMOh+JByuqLoLQHS7Z1YsprxbKUQIQE/3Ccv51hN8dn6g4dKMeVDj1OEmPG3pgfYvRwIosyQh
ZUx2xbL1Kj2gYRVFI6p9Yokr5edNso2B7B4e2MaM8Dw+R4LN80+snUrRIIV7dqADiwp5hOVS4ayy
2odA5yrWv3aPQSL2/HW7kS6gjexOFFflMA6TPP3XFE84tauXmhlj8T9n215Ge69YhlPXLHn6uxR6
P/2XKfx0a31xGddEKlN2iU1KRH9AmMTvSsx1HKEjT/6im2/F3CsBPKsQJAsVi7ccpa1GKl4xaJFH
7BxKBGkHxHcdgouMob+DCidCWQJUCgXEyJh5WsBgcYneQTAU86KcxTNhrwg6VLxysc3xnfLUsJX+
tkCrVP9QYPdaa5sNc5+PwUroImVgjbiKzL1LKNdPK3KJ1gyjyP/GaQ/G9UilHo0fbx0L9My1Kt8t
gsCPMj5O97OVqwnsYDESzH+0rAAZhy/UqzIfCarRq2mLQmgxJ0sl0Tpr6kkdtGUTKJR7j2c+WsTR
wk3yQDGEmwGAusp3Cyb5SEdVqqzhiIKvD98DTJU5rmOvCt8KCl3mWlGf1EP6iXajQmb1DRloItjl
dlV8hkuPW4fKtnoZSrdbJ6rFNcATaDQhMJzfv6r05qcrZRUQA2oagb/CDNzRo7myxW+aFLZ/ttch
i6tnyULk2gAqD7wkhyPXOYqh3G/KWX3sXSfwhzpFPQmidAt/KnjgyUOE6kBlb8SoEXqgc//7aZtF
nLl0DSXHHrL1LIgdrcKBlfSTxKStLze64UvB4wIOobejFhJmIdQzuhedjIJEP4lnmhoDdq5jRVNi
3jAhM72SjnwP09ihB+QmRwjfOtkiL8nGlRdqFepy6lqRJV6EgggnJs2kqNUXKHcTWVgkBXqxe6Wx
zaKrzFdYwY6PhombghDeVaXgWnUmr8vA0Mkyb1iNi5f0ZmOf4ixafSexgeEq8IO6IWuJhbJw3B8D
DlYtm+vOIybYWbqc9/s+QNM9WZ7QRDj28S+1H4DwQlOZ0G2LEMUo15GH/mbxcaS180XckAm0uUba
fP6givWcs2smNjP8Yk2hVoFq7H5OsWK1NYAcDSBEygIz8WK8laqVkym5zYgesqugTwWlBetM1EXp
BspI4hPltMkD9Pl+dmlXsSxULC3GMo5Os5QhCZDy4vpgJPrLZuufSSH2WEZGDcKxiwx+iVVf5Xc3
vy9vlaAfNaz/7EvpuOSCdzJbk6Fye4RTgCodkCtVj8tc+saRvTJX+hDQdAzSec/E1qk+5NSZTEiw
/rMiy+JnFJQb8fq4A6aT90/B+f++nO1BBQ82QHjcYigjHQ6k6iR7KFL6PQwxLk4NPSkLtsiT304t
P3C7NTcKcwjY2eDqqtwmPUl9UlBACrBfSpd3myySLoHiadxqQaaH22XcTJedh2RimIeUFWqs5oDZ
qOOIFEuinsxbeMsLT7MoglpctYjSwMYorPfN+gVskYhcdXfkfHxk87lQ9alvbr3As17j3UW/xDpz
yU87ZLlz2xozNCLBQp3loEl9fA2GRw9V+MXmRZNs5oGakSzwsmZ/K7doA7NniF9LeZyJQQjVAhHP
+tOoitMyNR6iY/tDcjYEA5jO2U0uJoFE/Liz3pp98nuFzM3QqbnXaPAWPlWwnMn3lFmKgSayPrv9
0Lndy7X3ZysPCn0jUU8oEqsGux1MP8K86LXF9rCwgo/fkOm/7wy7tU7EmPElBtc0Bd4Lp1HwQI+j
yObbKGXj28PPivkRVPq/AqwApN7n+lp3I8+2ZoRbiCB96QXVQuwabJSyCZdNXkHzoRFCcxQV+uqX
iVy11GcgPtfe3DCPdOlKe25iLyezX7/2wWRKcOYL8Ygb0+yL4hHbwdhHV6lr+G/Gd6R92xOBZLfB
5rzkIht+IOZAnE/NeioCzB5pVKnCCMBf+TvQ5vTWZijIdYLHs6JWzkiGaOQlZ/cJ8WGqCamWwr4t
tiyum7mWdQW9sYkz8EOEV8yXVLVUoZunbxT3uzM9JFRl2sjQJr73G2zQ3Ze0AoCFM1HPjrGdoOeY
FBnLPdSQ5LpWfndqer/abAz+FacQC6UIJertyixxj/XrqLTRSB5SsRoS8y+/k5dUPILrGicBVM+4
c2ZttzxKuSRCdOXMLu0MoaxOIu3s0TtYumgIeB6mBtDklVz5Y2o3nIcmvoEV8kQfgXmXHEkjo2Sc
AGUvg6grwRIShZKrRK1kr2YWOkCddYAFCMljB9wov1WerRChjIIJRh06UWuDElrjK5MfMEX3VtRn
zEHL3o3xasrMjanhWwy4LPw/zVf1zMHkKigmMiF7dqUOvRK+wV2Lt2rRdGqsQWg9zExntQwiZESw
BG2tdUg+qup3HJ7dDah+a0vQ0gljeOeU5xeSvaI+CHbrSV6NryAdW4UEow+iyE/k5ZcZwQd5zTqi
1OhRTOsPLzm6Kj+TFp/Mf4QJrX9XIgqDft4rH68ReE/olQ7kYeWDTS+XX0tz8E7i203AVTMcXiNP
btbrRl1JHJBzymKHrO0Sb/ed0PZxz6vs9/sfTL6x7oAvEMFcr3NcY7/IH7iabRfAaNMtvFE270zT
QZ2+vK6EqfI8d+hXhFIFudNwgVL71ACvax+RZamY0ACp3EdemHMmM5k83w8zKVkQj2r4tTueb8iH
ov1/2NcTnj6Pr/6feZgx4TM5uWWjiB0P8KayWFwAb6NSjrtFO5cMQQI9sC+jRqERB7zNIzc4sSJQ
bXdin2fE5H+0h7AmiYIlOVj8ZRCdt3mn0R0CBGzjIMfTF2UtRwyzeFZulED25zRShKQhYDT69FHX
8mricuHNy5q5F5oI9wJodQeuABiAkYzWGasL0OhwXxyJDpXRFKBjZHnrSIPdGKK+yCXtPCWiRdKn
IK3WFtKJrdR4HT6jCH5Xw4/bLGejVnSPaEnWpIMwB5WHf0FW5G4b8TcTXB9+ERHNI+CJq+Cu/qXH
zU0/ChIn3akl/uTK5206eNoix6mcmnPh/Ff/Ii7orlVPc0OvTWU5pZNzIAa3QKPNdoY3CTtgC9Mn
9EN0Tz1IIKfYjC/0FQS2ONAj6g4hGWO+3LPYe8hfI8ATLqtlSlxi6PXEUz1tHUOfWuC87SgQFPDi
5tqisoLmb49aeO64qV/cQOg9XCfhKxzaLWO5u2UtD+C3SjseFYebd6LP6rNsF+XpYO339gyCyp0k
aFUd4g/CENbLUZAdF3Jda/l+lfXuB15VZ6uBBQXasOzni2buagEMJ7o99qr7cMzCFaKkuUMr2x46
SUYiUcUdtGMULbEgvKeWY5b7dUPo9UetW3r0Dp9IpapHTaBVdkaPmLjJZNmik/QvkgPf699SV7+p
ZD7peODUN+f0mHNI2h4NtUvNQzbdRJFn1wTNNbp3MDkIGLuq2iUhIlFU6v2LCtKzJLf+ZKhmQUXR
ZRJk3Gi6P3mpgevy8QdpWjq0XWsJucVq5yAamKsx5ODYjtk9UYPlsdVp/LB+RgNr5W17V4s0vnpx
j6ERIAsx2qbPNqnKQnwVD4u5c/FLNhDBle04NoXW8sflcmTaKLFAk+rM43N6bQsjaEfgHiLRMg6q
GRvJ5Dpplan0KUzY2dlnqmctHM/JkwzX2+0HnH5QvR9ozkKSzqINEshDNgVqachP+LuP1cQRH2I3
62NJ9wRwQuHYnVYiNMBkAZF//4rxQ4mMdcrZuMZn0OMvCN4/UOBYfAFjiD3rDSIauNmGbhfQzVEL
4TeKkFXlWuDlVS4gXiWh8zJuEA2phEZXsQihoTOSX7+qxUhfRXK6iFEGT1lggnnulwezoYFHUgwA
asfVECaN7cMCtUEmw1m40tRpOdR7PwNEE+0/s+YmUTNxBBJbt6gQ0qZ14L6Aflb7FgwvBHVTAxwg
/7NUuU5V40D7seG/zBK3vVvrBdyD3+k8EfNeoqmABMSjyOq/Mwn5KvwmNscXGw/G7XxyODJsZgGD
nVUccFsh8YAqSB/dkE7S9LkcJ72qdLxDewXcwP5vs0pB1F0MDLDHKdAIeUmwSHhpPSsmtfdd/yvr
DVeFe5psagrlWEGRkDcWnLoQcah7CcB2OyWpRTFINQuTeV1SSXxR2rE0y5EW0lDm0THku9RTqPCL
EMxdGGybywcRj0T7V560XQBDRPPRVPdNV6tkJMG1x3G4evgKoUIoyYzsd/VMTa2sQJIDeJIKCe8n
KxOoVhMHbK+rJ65hJgsoNaXjP3ElZaawn1mrrnh9shK3Kc6Ie75gV20o+7cB2W5TE2683uWDcNa7
fVhkv+e4SNbWP7Ix59Vb4gnnRDb2fED7ism/sVbvsWKR4BeJXDuzdLnBWCfJAJNlrosmwuV9PTlG
N8auL2eHMk35vvDDH8wqXgKIL4/E3yQ96uiGzpQfC6BqA6VDn0nlBq2LjDfiv2yqrVF3SUDZ1SG1
q99ac3DdiugOMAYsF0RzcSSSyPUJ5LY02WG9xJlPAaUCK7i3/MGAr6Fqp2hrsM0Gsm/haAR3xMW0
ZlDCIfBPYX/Twz5MpdeeYH/LeiiJwVlhZNjw/KFDfjpP/qXAfYHuYdd4AC+rM2Z0SyE1OGy3dLjw
9Lw5zyYYAoH7lSv4zsauOQWe/6oEWmIi7Zda6WSu4dkW1M3uZIJ0YNsJCSJjUj8qU9Dajn4Vd0f7
oYbn7uP/NNEYyEhlAwj5WPKgGnxk6WAWAXMlPLbBjoMRzR13unvjAbMCBYPmSFigwU7DCr+arPx/
uPGLc59GqrfGwDaYHi6RrB27toLH6S+SFH8zQLOD3jEjLnjV1ZySVb6GlicVimOWg8A5xTz9YX9J
PSOv53/p7i3WPzwVr1sDbi1VNaGUZFQpYJ4d80Bp+9mSuK0ZJzDFL9pFgpe7WH4e3Z99sHqXoBwy
WCnhTEQPSBoco6lkPXkDHWnQ9AUCgt9pgI+oEj9S9PeILtfQ3715ucwN9iYkI0ZXm8VZwBEDuDNa
XFyAMM0ohTKIIFx+Zz0+kD9iBGsY0SssIlfSE5N0lw1k7SJk9kyR4/4LNoKKpdZ8NeuJ84nJxi6C
7bc4KeBSVYADJU7YjcpBe05UdvxL/suTAGyD8NZ5WRBNzW9cJdvSgcWhry+5VxE07lkvGACbfKh0
p3VNTApX8TO32KH9eX57XpBWFwHUiarxqO//ZmRP3wxXpGeoGeburK9Yg5odCoCntlyIGxYLYrB7
uuFqj6pEh9YOQ1IZ79eSzxou2ulDkIH5Sg68d4AypBxKJkeirWqZWo+bunrOtkGzToJfILL8c8+U
XD3OEp3pqOnSQyDBBV5ah15T0Xe7s51qaVFxtupXgPBOUJ4MOW15rwKwMiKeTQeAX+7JycWDAdsf
bYbNNYA1DPotLqvwjZDPLzugI2EPL5733iJey5q6rKiPdecMmZv7U6NSgXff0Tq6sag35GZ0CcMo
SyFV5EtQph/G//TBoZnSdIXKRR/OG8+ZBTpuIsn/8Mo0L8LdHnLUuhj4lxvPiSUqgZ+dVvqPddZu
O/m6BGKVyuoT1TO55sfpp93l6smra4jtIENMOTKTmSplzkQF0UNZtgf4mTrkiYBPoall9oPzl9LN
lT/Vy/e3iuPGZ8eM7nKCs3o5P4hs2T/JP8tecPn5kObN9D8QJ28NzUuyclrg+pAxqS9nPw3STORQ
ETmQ/fIOvmWGsybk3Eq70ysBiHRdKJ55tBmVRzFsDnKKUtVJEoPbGHhjVQlfdVnGVkLjHL4KnIHF
rQXLbnKT3g9pI7IXVApPGPnhHuAKmH+OYuI9lxXUfyldAtP2dguOlH0/aeRmVZT9y9zLTAvH//qd
6IV43/kzCb+Bb0LffHgkVIHO05BE5Z0mkssfltEDD5HfbnpHmBrh0jSiahxIAPjggkcfWk5WV1DM
Nyoig+dMcPG+z+/1/P5rMhCMY8p5jzmj4B1Y04xNREHFvdcwH4SYMhBvg98QLH/3udmAkZZE05Z8
+hbxO8TRsKMJDk/kEbbDcfwEpv54QroirvLHMHToU4AhCcmgR+wjY4zQPXzmGTOBrYeA5AouVi+t
6RBIlAV/9MtnGp2Nn3WkRmT3ybbacbdVN9wMOMQPIuOKTgOIqyLidcmFWodnA6vYnQCKj5I3LciK
g8MfpyWSK2YBDYA2af8qAM9Qny2dfj/DV/EgL0kTyiqxS1xHj8cjlv/XfyP/Xn4NJ8qmnZzplq4g
zzrN+TYmbOt0qq0xmDrJAeU79rOAMjLV5fQCq4d5KKTUURd+wazuXseDlMvmmDsdOJQgGjJUm2Tk
YKc7W5xxJKWFsINg+A71csr+BrdpwNUaPsyqABrH0DGtFPQRMZ7NuEv7bz1d+Aukwhmw12K5jMyp
I7Ct31/TlMGNomiuceEezwWNswJ4j5gHQm/L+8w7Fak962/46AHGbaagBmo7mnMUqJAwwZ82geZK
j5HMQZQfqDOtEbbTt+9mexMawPbL78WW/QrV51KQyrYEHpSgMkBtwJsJnGb/FnpkmUsJgntx/78J
5xykcr7vR7TUMLAabtdJr3RLdlVgrMe56V7D7G/5AvjpOP1v/kFdX9IgkQRIEdPmeePuULRknIeA
vImOZNNz6PgxD/NVjEvcCHDFYsVImkGJcOU45BRwzKKpuWju7/QJeIgxVtDi/YYmMX1Cw0tdW+bG
o026HyArNaYsWEvLraWO6+hR1e2Kf+82mmZREw/LRy9aFSaWPTZZP8GyPflhjwCypMoopXLPI5CN
ALk7zzVDnfNm3bldVzTbGkdgag/3X17aHJewxuWtFxoes2SJfVE4J7lx8Txw+F7tZHJa7/z8RJHu
gYsQl8WKl5fq8eNEmAMvJuoLWMriTkdpXk/R2tfgjVNCtnW6QDSvhbMp1W1fG0b7cCOhGqipCKDp
KrsIbzkaG6TH1injRuM+mlcxPtcq3zhi76FF0wo2vjNq6GNYbkTzJQ7AqLwTpS1PGA3dT3PAgMsj
WpaIklfe58R2/nltgB9BjX2jhNZrx3oD7IkzGy6DHnNRkX9vmHnFiqbBU84Qjo64Kui43kGKc/Jt
/Fq5Eirv9jse94fBRBRWrY4JWSk251Ea5M+Gq0LeNjlVHswP4FrZrSH3SPwe8LFaJizxEIUPQ+33
PSAuEL/oFEnpfLG5tHxRYs/Ne3qYiCtuhC/bcTqfjrlYVAYfHNS6UZ1FCU1VVuhvDmuLKEFvJ4Re
DPANmtmhuv2zzqNNZy2xL3kh/bCB3z1czcUJS84rbs7XBrsLxjf5ssodZCXd85IzjqeD108MFfGu
DhXwgAVHAJyUinlfzhCeuulxw/RIL5hvGN5Jw5yy8mMdaOA7U3o9HlOhLZpmW6RWAcBBTpPwPq36
3ssGyW32taLMUyzhFFGSQt2v1jZ51Dwz/GVd4R9P6VUaoKgM2fv8LeSDPW0bm0hrYxcY7aYsOdbq
ME80th4eEezH0Navni5WeX6Du5pEKmzkL74Jz3+4vYuiQ0YO+HD1lqNlWhgspZpoEPwP2hUUvqbD
pZy5slOUl/szzuo9o6BOyYTvcFryVS4KRa4RutM6EAPVuHyvuWwc8h4t+v5GUTg8LKNRcNtY3+Gk
Mg68AdEsfbpqtYkKDs7gQENo0O9991GubsYLGkb0Lrh9CupfQoP0NA6yWwpeAWkJCAd8UkI9U5GQ
RxHKPx8E8CnLL9/YB9mcMWoialRlaEPITRCWa8NsiI/xPtXv9dUsqA2qCucVHLwLJDeXJwT4Stnd
v5aSHgprDWuJqN/5mzWMES+EFhqYoN+/xAvSzdLS8JpP15fZcTiXvmXBFKbqoZYo9KRET/Boh3xS
8W2USdMboIdHe+0tCYPxXWDoNIIF3GBqLUkNWwQHDoIuVljnUdAA4My+aVivDGXLYSB22EQS9rBa
zmVGPACSYn6FgMCfA7ptoCSOua7UwlhutF9en2Wna59QRVz6n6Fl3GyMZjOP/huD1iLw+VcS4I7x
NukK8bbBIYltDFGYyrXyT8dN/oNZx+bOEtFPyKZ6iJYh5q8U/1WOiWD+FbLDF2o8sXk0X+Au5EX/
R8ZeJOZGoBa+l+otkp5ap4Hx2bq027gnsLCglTj5tO/J90sIe8w/pkK5edF6BSVVa7jSc5RJM2dV
WgYwIm7wscV7Wd4tOcI79XXvKXp9vMmmWgnN8R01Nb5LPMHBZpky4Gt19UB6uiLg6M8oRzA69lj0
CeuheIBUOqXJHRtw4wqwgRc+73xGx9Ofk1P9nuh1/5KGW1/rEDszHPAUBo11wb/E1S5c+Ba2DBQn
eddilPZORuq1tSAJR1fNGzq45Vgd/twkNja7/keCTIZyUW1p8ft08+sRVgpbv/BCJYYzinlShZR5
dT67hlnuJ3EL24jDYTBUChlpKsJjPwDabbQIW2wobxZ5QMV0ohuMNvQ4uJzNxn/N3QFe3+MoZMqd
Pd4uzBHMOWN4Li0xFhqZsbgp21Uy9qENckoVgnxhCJD8NjQim9tq+7sU0rQ/dVNvHo4JL2psLvFN
4q0qcKnU6RG5IRKv7UgDtnBmQ1KaLUNegV7jfD7ZBJWcXYP/cglfEcDo6/jSdaLp1i7/JcaoBaTP
dfvvHidY1vSskM9L1e/Xoh+Bb2odma7HIru5oYVfFRJ1cnZeb7RX2Etmxhvski/oIdmoSlCoDmHv
gYy+G5NLMvorx5IZZr/K7k7eQkTkuxHOgH5xT7sKhWnwoKUOwiP8piV7/lWeE6W4Kb10Nd75yk+m
IT5I4Pj+Ea5xo9WkdZ+qfJ0vOGfbGsic6/2w0Ou08oVo9ZXJKC5eyMFVuc+y4nEjdymx4fwlAiC+
igMPEDwN3hX3txV0qeO3eKVrl0WYo/2LxzzBbtWVAbzqagm0qlhX+ajpG+Opznye3Q7Xj18/UYA+
tW5ta7O71zSHMCZTsnAFcxoH0HWI1tAPbM2Vwx1z8iLof2k9W8GuwlTR6ZPtLJfxG4hWd888NKSp
zRykPA7xcu5Yp0u2YP3PRUvim96heH08nvsmeLigFxMBk1fb49kbkUCZZSl8EVLP48mnO6kwHGVJ
VMVs67pRGCUwtu0ZFGK/dJ3XvLl8DuN9oIUFy5nVkED1Y1s0T7XcG/RFGWGxWvDY+p+N+ZI/W4ri
L58V3MedFrM35fjf4Fgg/UE223bbQQTg5hJvxPQ78eR8e9r2npf8Q1OiqD7P3ZcSG0xqRqdfLzsI
Bn0mE0onkUBtPVA/KNs0raeO7l+I5Z+ZZ6MZVgrOdwwl96b9xHDQ6jLss/0zgvpDJmJmKCyZMdXN
lkSSKZu+YKcBsYzpLZ4hDik0zlZaWsm7Ag73qi6q0heda8G/DED4gG/YBpFQvfAhhb/1y0WuPkbY
MZ/1QZqMc/Wm9fInhvIOyQIRMbuVVWMYFcLl1mRhO80DXo/yIDmOOmlPqOPHZ6EFJ2xLzOfKBlEN
6qpdMz309Qd8UEN3pdNlSfS9LM44mWPftgVmvSehoGSV1/N6IA4ZG5Ihkp2ytlxjluTxFrs219g/
kZNnZqOm8+YQYfT+mcRizzM3y+ZQoLXPUPfOmaSX8/FWjOmJC/L7dx8au437cngPN7wm4eukVU/5
j4RwZtvNRH8+Kn4CNzTi64P3m89kVLgg4RUyii4CEhIKJ0dHq1N0RS7Qj0t8Gxu9Ak+DFj9+KBUV
4ot5zuLEnWpcCoOviikralvP0tDwbr9H/62th7ZGIXlJ8vgePKg/s8wson6vvLmJRzVoaJmQS2KE
D8628GKfqmG1k5EnoU6PJZp/lf2sG1fKlIp4Xk46bXGkxFcTEPck0p3BGcmOj0JiyYwFXSYgLHbz
Zow0x5LJneU1c5+QE/tIlkZuJ3I3heXwd2ig29RmO6wlya0ZYddCRTUUYxFYSynGMU0y1pCuK6Y2
2qIQjD3aFp/haUtObazetyqGuTxzGVtZwR0+d8kqVVh+xydTJnT6qtBhQDx9K5GlyhOJulkE+n3g
mix1kelX/61xVPK1ieqMtvGUddbcpgvFuab3AjFbegCgBy4SNrAxSg5Totfmz7oMDcNR25b/mrPZ
MENR9WDzPRlKc5e7ALq115gNvGl9sFTdfylkVAMf5qPpoOdkHlul3XEoAgtRv+fNefO2sQJgjacF
RK4mtom/bS4IGuixM6rMQ+XaaOTfS4By2Z614JIw4cn0re7TdFpmtOgbXhJHkzrjB/NLze7N8Ra8
eZGV0hdKGGsM/3cPtfB19LJZzPQhP4O7zKnRPPPiMY+u7n8NoOXdpzG/DazfD+FEAAeg2sO+mGbG
IEn/flznzhznIdV7DZsIhcXaaaNcE0q8AVQr5vo7Sy0kP7BcToedupRg+xmz0/0+KUJ5DVXrIuxC
v15o0nTSjcOgPmDA4xMKWg+FP21Jn1diQuz/pp0QAQBAbEh9u85CeqFqvaHMPn/8v8rPUOrTBW9C
nA1nxDmpvjJwcpkaN9hFU8IiU9NkJW3S4Uzsl9gzwnksS3ZUeNBb31tFivbUI4mosJXR8leCJKlv
n+ktHZ4crP7SCbrKdouPu+gxyxQuxKa4x1WUxO1KpzI+KApRzy6caqM7Lv4hl4lJQtZaWH0xz1c1
AU0m7hMO84wcQ6/ktwgTW1tni8OEqIJPuJRx182/anyuSC2lYbAvqLib5HIVyjOAOWtd0+sUH/uY
lk4NFaeTCTobq69CRUHQ9399HCd72p1drjU4UfIuSsueO+BLSRqQuaDeSMXjIVH5wCa+cHje2+Z6
dVqRs91tj3RDwjhtGh7ckReWqM0NrnzdbRuKOIWgqMu3KtRBjLSW9gbfKZWPQH6xsnrztoMFcIDi
25JU9qr4NtT46lTgGet/0q6Rh1tiOOWyLykHYf+Kz1OfC1YBroPUpcefpjWwcNd6qmCOfshfDOy6
uDBcEFzSLe8kBEVKZn3q/qS2t/Ae4ZNkws+KajEjxgluavJZszVvpEkNWtclrnoot035u+vkpE79
YM05P+oJFE/4jYJQWpFkjQ7ThjreuiNypPvo8S+SYAFK7s8zqwtkZGFmOlgBLB151cZ/kFlbwoCV
6gYWyGXBMYPiKwrbAHUZUfyIxTJ3qB9+FGhigFS98mzLW5Ys5Uon65N3+INq00xrvP7AUKtVPtk7
qKvLtacvsqk/nKLTyRWhi31UQTr7WKqMACDIgaUYdLUQFd1DnWdjUJAfkHW2adh3P4Y/eaxYuOv2
C0tGGrkdxUL0b4O9L283pRnETmggcjkcayfZti41Z8hwiDDPozx5fCCfLSfMk7hrDeWvwspo/42k
QcQ2/D3G+g9xe1VnIE48IqTB0l9BBdhhpEOUttCvNYDC9wnlxGzN71d5EPvgDrmwwppTuocV2eKq
vMiJcn7No298Jaf3pofP9sZeBHoo+pBQvkwJ8v0NJffK797rTi9mzboiU83Z7lrbU5h6ArNdqRpp
FamDvA/6VizCveB2Bfm/ns+7hnEEn03wupTcpdwyxP22IRwQWMMq8ObWDZ8k5iOW2fNgL1pmg4FQ
0ieLdzbxQISMpVTuItfJvjTJ2dSHHMTEeJ+eyQeg1xNIvlL+Bro9iauV9Qa0vcsYH80zTXZa0cYo
aQa/NSMApTzR5E6SktL7A4zsX7kj5Xd+jgNQdjz7BSpRFyv11Z1TIkgZuYWEekrFhbd53+HHTRg6
XZKK9FjXL/MiaA8bSDx2d9MgqwaYc9+8VnWI6L9/kMo+rb3SrGqaQ1Th0tkG+vo1sbFni0xZoPlH
pvG7eFm8kW6nwiLFT3+S/er0B0XAfT09cotf2MBNgPXIXDQmbzo/HD1wixxQ8xiORX3GQjSMp/Qd
Cy3hisFJIen02HgYTqxFDrLDkFh/lg8u7b5CYaaq+ipcR8GebwPgF4weKuo+cOQh0bQsLUm534+i
nIOGYRuVZsiFwSv4zmy/2GdaeAugrtYBWRuEqsxr6gASUnZ5zKCnF3k6jn5kGU+plN48D9kNAMJw
3YNgLV4kE9JLk5vJHPAtCouQ5NLIwxnpxjky6PZuysd4jvbFD1Y/NsfSOKlgYoxC68NLCzLtBQpa
AjbohTvUsI4k2CHCyUhAlyoJh3j7XSZgyEHuFxxLMxd/tPwVYkZsmKh7zAJMr38ER86rzL4g9L7Q
kkSBa6Bs3snASQ10huHBBSieHKp8onj5qGZgN6CkjkmRuajnv4zLDssKDv8D0WlHn7U42M/rTk2C
LlqJeHxUj131IncD85gDEguvVm7l5gUFf+29rQhDALA0FTAbpZKYRK+xloYSPfkvdAeJsAqSCo3V
X62joZv8iuzV8Pm1ju6gpYeGvJvI0a+uI2ioHoCh+urHyyZRL9L+/eaJ8EnuVBBY+n2iToLCKDaW
Z6+1m+qedwXJi9gp1ZCmd/kzvR8o2keJNFRaC4VUZin+PoNDBoE4DDGasa+7TLKAjN1IhkBmmr0v
v+2pCWzC9Hg+ABRjnhNvmovS+3ah0Zv7qK8RSQPMVb1UGwuFmOgdUdKPVooN/lIq0RqqQTsI7buC
skgiNx0vgv566xorzXjzJ7V8+Sd/I+zibWWQVjeCS+1lKPDq4JEsA4HvG+V51Z8DxqkXuyIq5kim
Fe18M5g6zfWjeYgzPxSoALl8tXBRG56sTa6DkJ8kOX4o9+58GhVo+xxqO1vy03bTuZpS8KP9r1Ng
bN9jjyV0bJWzrSvhaxpcfk4knc/HsGM4vi7RzriT6zEtIn/If2bJFIwtqwg6ZXIrDkRJJMGY2c+o
7Rv3aYU1L+xMoAoLuAV5JUjcBq43o1oOKSaMlBrxZCR64KLci1XWH1lMWHE9q1PvXbudi2he0xZi
H9dJivMozsDq01iajkcAN1Gx4AxO9L0Wh1hZ6cbCwAeio9s6i7cDopwuqDlc6i2hCOfKJc+6+lfu
VovPoIlhByOKILUiv38AQiAx/X1MAk1D/qaDaZ/HZghuOShqEhFQsi9WlasvCXHwTgtNRANJf1ls
MzXitpRYb949KjcbbvKlUMN0BWCsoi0K3vI5RX5hZ4ZSgXqqmGZjHOgFBjUKIAQ7WN6uw3VS+VuC
iDO5zdVkXhgRWg0wpAFgD6TJYQ+BapjuZ7QMImpvrpoLNE+3KPzPyRhMUBkxDPp9AeEz8sz5Xmpk
KXsBjykZpRfhruDjubVounJOJZ4rh0pEkMuegqN1pSEovxzzcGLWEOTa0/XHXuuyLoqGkRib39CB
DQPkCfvLphvu0pA8eKX3/5aD4juJfBulS8cpGCiwbzbnaFoe9pKnmcp0XsKq87dZh3eMCfVGLhMn
+NmR/GoPsd/6Q0pWgTIhdXgr4S1FA5mlo1Lf+8evjW3Bqt2u+CB3IHREmPqQgGpumipw0+fJk/WA
GP28IaIe6Sg6MubVJHf5HFNG0BL8AjLP7kK1o40KFAcbz/hijJz9TK3LbN8Hm07RUX9BjY/LjgbD
Lfmhr65oaRZokB+6wSbhNBO7TjcEm7Gc8p1ml270Rrk1F8pTjZPY10TLuTi7lW82SEgmlITYSAW9
NsLCq+44jr+tK2l1sDwVlPJy6GpTRYjRJOaHlWJZMk6FdWCkbq5guQdEHjWMipxZBd4OcQnCahYY
CdlZFAiL7wqbh3uCRn+GE4NMO3LzZWcRK065We1TifVg3L4CEVixrNTxbIBuM9ZhfkeEpm/6houL
X6C0GPTkVBLPux59z8I7Pr806u1VpsRubqchfkHmWpbtCCogaxe9KMVC04lr6AGBAcaw4iKn67fK
PunD3LA3yqdwmYDYVSX7+F0rMmFq+wbVAiDUtxYnRf4wpGoR4N2GOrNypZIbNwPsjH3qPF8FJv53
MWbluAcUi7kDE9aUrUa61MSjId927aPLDPAr5WkHcBQxpUGd2OPXG5S8FdVKhJmzsU7GjFLft+ar
qjNnuB54FojQncP7cOZwezTwZj2vrWGsvVQ+ULr6YPHuBAWXY4Vkchxc7yWFs0LNT0QvYmTvvC+u
FYyj7I4q0OEeeiVSqQBgMOosrcMOYwfSyqAMSX/JvYRWgPZlLYs3J6GFVoZUCS/eHgHbODeL17JW
urkVEtNC8XgecbX0twBcNgnFqpz1fbt+N1EJGN9uOgZWWhSAt3ZR3MmVm0aLP2cyAVSMttuFiBFz
uAHoqTJvRVGltB2hXKrjeRrHQom3x3td1lXgNRhkawU/6iKaopByfyVut7gmsF3JOGCHSseNDraX
wgf/kLTHphMavA9KJmrJY4JrnWufo90qFx1ylS2TxTqCeJEKZLbI5/hfhrsyqi+n0CtFND8u5c27
mVnxmtaY/0zynsyzwYzQyfElHTiB4J+wO/jaCE0lg+r4hiG8Z2oLYatEBqye7FV1PGbnfHCKpiWG
ZdBHSwiHaadxSMLItgNiGP13aFlDetzRqji8WwXY1/OM+t+LoeAmYSnAWmZmkBA2gL+PNi8Rpw7x
C+YfaKxutILK4AhdiMoDN7+Zvhg7va2ONA4vP9II/8nQoAVkYhUNT7yRieDCQF6qeoC2h1ygaYUd
Rz6xE9ob6y09AOSZpTXxwXP+HBlle8pjoecFPFozM6+xY0XqAeqrNyJ8RemP+HtNegpEHcT0Ikhb
Te7oxyO2f/LLXKzsDRhAAflhsIZMAUuJh7U0S/ejOPSaKhLOJffqO8KZW7/NxwmsLkQcrd3tDd76
Li6b7YQsXxb7EJFirbO7Rb0lgleGyHNzj0FQPtpWdcMZfg/rkkJinLh3Y+KAel66vdhClun4T6NZ
Z8UHUeWLflvPIukFe1wWk2wyEitszAv3fW0YgE/nCD3z3ZkzWovGhDcQNlw2x0w/7eJe5dXuMgGr
7CVB26dhBDtdXNsc/Hr2U4Nxl0D/f1FodwMu5J3qVPxVKm42a76RqLZGXZE3d4qMRY85Dv0+4l3C
qeMfeJIeblrPEY6HQm+qanp1VFBNkg1RH7DEo8QkjGz7jaQ1JIXJ/pm8elgUCp4AXplex0o3010f
6QEseNKkE+kPhS/eDWUgeRakTy6hzLUyJczV8fgVugmbNAq6PyUVdF+K7QYSUq31RygB/kkBGmc6
StlYWqUmm7H2r5/xfLM8C1B90R2qPhgFx1v83+5DAPAQXJ+pdB6zlZIiTymEPrPjx+nspL6tTPkD
v0t3WoSR6pVRlNKnmhsaUrRS70uwA4Egh5S4ud6NXpiyB3iABdv6G0orTT2L2PErnZywOcGt0WF9
t9rAMYgkqmGwlpOVA3o2Z0XmonyQ7ZYqxQz/5AoK7k0LPmsP8xOuCUUdIFkAZRvsOtMNYw45xj+l
fcsqdjzqch0fFD7+2iaZLxubcoNxFBpY/gAUa8xP58PhaBIr6z0oY+7jPLOyBCq6oGmE0XKMu8c+
w6bioqWhj6erbUvkgpU+Y261p42UjzoaiPI6h2OJNpPft+VnlSfnClzrgjzvmBKYPs20hPq2TooD
e2gp5ZImuFerGzI3O4kT46+bJe+itCMSX9NO7ulydCoxzzVNy2ZXqUoBJY3aYmVsjoncyC/FYR1r
psFpCmu/qhX/QMju7wKte/fYxcZvMMgn3u9kpjuBDhjtlMKMFeVrNLm3GyoZpnes7WENZ4ZQBspe
XmfeVC+j2lU20cT44LoXKJVNf636+7hRGQTfL1SIgsL1r0kMAx7MJsEgbdc8/4jCTpITMDEauIPn
FsYZ8R/VSZFUtNc2gC4CMdpqItCSRH/vw3NHptX4XstT4iDJHQuHQVbqodv1bkgyWUGC9J+k6y1A
pXAGYkrgrokX7GwwjtaL/cBCKUL4IUxRSAqQw2Ai94u4O4hJqGwqUDqZSzfFCRtOAntFTH6PegWe
7RkzzX1iXE3dehOBCbBm5295i0K4WOFut0NPkQ2JmN0vuyuDLiAnAogagTHtKCsdO5jWPXDOFQ+e
yDSal8rMScFR8N5FMrcKqY2yaZ/djJ56+RdiVdJuwyFHni+EnOQYsjCZb6fM7jkytU4ATXsZuaHw
XO2OkI29+hfPGWsbb4XOazGT36syF5zVPWp7qukKmwaU2te6dMT9hJPJs1PT6wp2SIHxmQYDpwCY
ZtkCXxUDY0xjH/314Og77gFczvWTRbR4eImHQ+Xh+S5g9+ldaaf1YTnXMiZ/oFdZxVUL2TSKFBuO
bfxSFRUYeku3OyULFVV54x51qTwqSpN6XUA/FNjuWfM8OdgOBsHjGeo/+12IwekZ2zU0HdrFZsws
ZfjhdneazwDTm9s7EaszMO6iCZC+Offavpz0dvCUqrze1zERGBbP4jUTKJexZQ0hFSQ5KVkkHzt4
I88C86Az7jVLeVakIZCJ5lV/C8NR3KZ/P6WCO9CzQabc7ujtkp0t4IAd+ci/gDZeKk9JQvUqJyZw
4pl2v9vhRKqjSnhMsmsLDwri5/OdgHaOQbfkBb4IsAWJJAoUAPOv1VQGuBGPgssIRfwShrg9GnMt
S7jYdzhUU0d+OsJkfv8ntazZsdK7tjmmZucgMmZEnzw958aNmUqJASoZfSHkqM9et3/yOL3vC6k9
CgIdF1c6MkNfVhZpNLsk3Ann908G449cwZJhtBnmk+/VcWHkmPiR6h4paqy28nMwzrXmx1ndzXek
VtTD3+x4Kfe5zzN4XKVhWlmPeCEtOWCM4r9tW/gAEye1g0kkkZ0B0rlS5lx2DgJBpSL98F04WpY/
AFUiYSAAV888k3X7XKlXnr2bHOwqDF/A4fDc3p5NzPy5PN0Ptw+0mU5bNJDBpi06xjanqPU59eo4
NUXiM6QQQ7f/5rsOpw1WdTLSpPM1aiQ5mYxizzoLEUCxPobziUaIJNOQE+h5yta/RDJxrXP9YbJY
TjcyVPxrKNYJHdMtxRy1tRIKD3zzWEzdj/aslNKEQ0xwRb0L7HGEAUkLWOGmbb9i9u4RLwUXnE7e
OQcMYpcO/HLu45SAjCzONONDCTZOdmgxMIhEgSUziryU9n4/1bdxFmgpc+vFuL6lEs9whu0J4ur6
aDxoMoc8lh2k+D7iLMfYh4il7CrC3U+qKsr4gJ43vtt/TNaKFcHYxdw1Y8N8gX0h/KmH25sMTQVo
wvjDiTxsCkcGZ5qUSE7ofsMXmL+tcEzIxJaQBudaJtIyaG/8To5ZDgFMRGUiGRItHcTUQh4kD4F8
AZ9+63vfnONR1z9mfkKPWZ47X0toV7fERVjHj6sgDjeZJVDrpwvrvKOrYYToJuN5HsDDS7tFPkj4
j2dyBsMwKksQFwA45pmNVAlYbBtQLgRjrrDbmfkHj7wEl3gyqwwURFRBj1UTKzwjBSy8E3H0HRdG
T5HXVjlKrVeuVGuIXxNIYlBpVEbznWU2SYY/i/nqPVFMqGw9oZIWkRJN4JspEWYwakI9jEvxOVj/
nYU0TOrcpysVGqVCpT13mJvvGraJLKD3HMXFIp2V/Z0NIpvoqsEsaSAC39xmtX6ahY/9QfWjZwnM
9ntOhZXJ2XwCIDlHLCT1hsJPD1u1L+RIK27SzYERFVqWZVeuj0X2JrWiC7+6SJi3F0RfeMvPdjkp
N/oJBSOlttj6uwUTItw8cv3vhP0GCiwos1hBeROfTtVUhcoQWdSlrE4UZGOM8TJNkiV3mujUeI1Q
2Jcc/NOPO5SJg2QxDBjq0lYslJZFUacqShiM+4HttFxcs2jdgyLKgiLjwcMUg77oUT+s4YyUb5J9
aGWf59bBFo+peKim+TlwJGoBjKLXmnKi8584XAsn1rlh4OwG759a+iXQo5Q7ihFmbps6B2tgJvLb
QvRJqmpW1EgVuivjz+VkR3fR3uhUU2jmT8B6ooK+j44yilKZWc3GanZy6mCl4ygTivVVD+vOTu9h
wJnat1J6TloSTCk2cBNQ28TryWYOf30DhF9icX49BXQlhNvXbqbYJd21REjGZg5omHNBahirpO4B
7bG86+YAWKRZQtAtfB+rfL4ILhBm7sypelulKXpqay6HooES154zZ6XdLJsUS+H4xoGPO6H7ALFB
wQkYNBdWhqhfGRRnSZraKj3udDSrKIU/EjsqlWlV8xW1j578rM1/HQdhFC0dqBeliLM+guAlmuu+
r+iLOdJMePw9SXWzoba6xYKi5kJwHBics2HMNgxfrFKmsy22SfBYJdOgy6VO9QWbX0k7YpirmhdJ
eeS2Iqh02P60A2TD+6o/FLv4IPj6E+c5iMjYb+c8OqORYyWVK7zpkq3ryR5KI6M1lQJ2rSjkpaIu
6c7aXRbuUDIKCbHI45THpiCmK2Wf4xRaly8SIKsOlk5ONkC6VG6TM7t5cTMz+hle+kmI0Kp0qBsO
ERinCuufTfLgIC5IhR0C/pX+PjUx47wuTrwzPnfcaeSoCJiViNtey06yTtf0C824ng4yLLfbMUXM
G8/sfEqNMTcN0ocJA1XeT0+hFQ72tixRqIvAfZ4fRdO0oID3tctnEXLiVmDwavzHPhOC26c3XEBa
TlezXF1WxpeyaDtDqJX3v1of9LlsanAq1wCCNsIE/NytUnJJ1gZ+sjXLQNCVx9H1pRaVY+Z97Ddd
Qkk47hXBbCbdK8KW8oqdwhPfwJM2fGvthqU0qfRCdg8jEqQuDbizA6uDMCunGf6MZ9BxKGg7vQmG
tHKJ9Mkr4CjwnGI/svy4Sd0dPbKyZqEgCYq7oJX5tnaftD8SUWB4musK1tTXQZcNKPihuTJiyXYh
B7mAiR8Z6myaCsPD4M6e5WhPu+ZbLJOT0tHCo3QvBswlaWIjotgC3uLUxzygIiHdgzc5fVBbzZlU
0P8XPXoomeHDVggRBcQC2WfjztB3j9KBuIMUh4upbTzmbr1SP4Ha6U0AZhiHZKb2Gu6NqvtqFdmN
2VVi9gh0HrFJuCns/eaonHG+Q5OyV0VZdr8TtIjqh+4PRWNyAkLsDn9WAvhLXI1QIdYZZPuZ15el
H5cbGZQ0Z8FU3irRZy6JfZCXLsKkuOS60jTz52eW02IIKQ0jbNuGWiEUgPaPpa/bwW9lwGhnS9kb
G0eUkN3mMlBRcX7/okNaxSGIzHBELRstYwuXdw7sGJd5BVrlZ6ES6Hk3WS+byqIXr6Rj+aqWh1Z0
GZf5hydyoIdOtvAYjswR4bUcAyUPS7qVhpvHbxhifVpgwU01SzYT/Cl1e7Xjzl1lBKmmUgL6imX9
vU8IgUx1mNe2s9Kb3CD2JFrx3IgD6bc5aGbRQXWA3Yop19fSjhybN1aFXLnJnlFUIoLaa3Jb1YnS
tZRJ408u6qs1hh11Ijpb3VhpxcKU/rbXYl8YBMoFzpxuHp4RRIHrwjXYXIbK8LMDN+PPvrLGmsFo
I7GXgtOMrRP6rLL+sPNQI/qYnDTOdqr6aEotlfEixOTXSr17IiPT8YEIeypP0nNOyfgpXQiTSiLB
0yVyWoOIebK9UFTxmSkEtRAfgVfAR86xbG2E0N/HoBmk0m8kyLf4efRFpFSgTRWXdtbtHQoUAhEC
NpBUr0Ysoy8VWLC1E/kT3bg+X7EhDzbtY99PSUk6+UnVy2EDijUeIXop1jpLdk1HLml+NUdVQQ4y
rIL9W8Avk2EClqdwsj2PU5dneWtNVkvp0T72nNK7tXD+hEqWhsGhDrhPIsU5eYsbCEDoC9zGEDTC
ijRVmkfDnLtFPhbtcivuzs9FNMkxxCUeuQZ0Ia8YhKf4l/kIBdUJ6Cr54NY/NRXROre0Fnmg90oN
zEoeOiddpC6SbSr6kGihKFOz1KVZDl40378n/Rcf1IPs4u7GJUXvN0JLUt9kJGG+/psYBENJ09iR
QCvmGkmZj0HZYMfdDrpTJGxivLueAWa24sAPrB8rwFeHh1oLJqiHKEGwd8dreoA+GmVP9ArnEG5Q
vvHI4C1b6+Y1A/xzyT99bYSGbRvUV7EanDusQ/qj5M+Pr8lFBa5BS5ZiepUr6m2v0dVAnkr/YbDZ
aU+Shbb6EKNk1Qaa5kBQJlip1CdGa9Jjd/w/KR3k950LZ8o1qGfvwB5J/VSbU1uZ5Bvtlbz9tROi
U7Oa0/N7lyJda6jdrHzxc1rjDL4VtsHfHRJCFOZtjVW3+dIfZtHqBRWatGyaCp2jroWwO8wf1uwN
R3+WDKtMh0fylSJTufOmy1j0fExG59d5Lnco0z8YryscYkdMPPEwPFOG39hvTFOo+JFKebRxm2OF
vf+UJiasdHxe0KSFkjx86wF/Nraa+RgS+lknK1WaB4Bnjfq7Eq96pVw2OtOA3dix/7jEfF2VJIQQ
m0Y6KwnYM3MobjUt+L2HM/kAiJ01dUhTyV90B/SZMP79i9Jcijy6D5eK47Yd+B+PvwguRM0Ax90H
AYNuB/upJXMXlgw2VvpEOqfhF5Uta3s+5LqtaafN3TgFeTcR/Mt7cInD+SU0wDkUepN/ubtr+nK+
mFnU1f8OMPUEVuRzlWdRrbL+lt0sIX3BgbC6Y9uuNEVESO3OlfWEbxj5yLfMNIBpoi4MTlagAuYj
2y3AHSAa7tukD/EXvUSpqxzLihh0BjfvBgYXo3fVaQeRdsElhL+SRSpqE7vD0RfuoK8c7KJH1w0J
/3pkf5HkZv/WkmTmrXtD55q4jrfYRU1TgQosvWrn0gOqvBaXjumYsUFlIdukfy+X46OhPBheUYvy
7Wmhqc8Mg5JlR72xp/opZMkNaOG4HwV2K4urmmIyfAfhitnbd/wvTztHDgFJUvxX0aRoDiVnzUhi
7BkHZDsk2afmQNN0X8R/WeAKGOD3AAIYfnKgshpI2NTUI2L/pu86V2fTlRkwuwcR2r7Nr6Kqmg3E
eyF2WwIc6kHkKYnwtEbC0NTPgDfnrjcCaGZGW+TNaT7Dk3PrtRS6E52bV0ExlO2dZRLl6rHRkmJF
4JVnD2gAHp3mPHFsDDLNF+Lp8nrUnOYjZh8rRN0RS66y/XUmrIo4uvPmhBuhHHonHP+J2Cxqw8Nw
nDcKtsoEPYxildEC2Hvk1Hu9Yyk6Z1iirMHRTx9vym1w3Wdm4QQtBLUHnAkzPHHU+mHC2pCDgDu5
KM5CENNYTnQpFGFrxBXhGDITFtTgHVGz5dj13F0yzKIOpXseWtvBuMTRY5zH/R+p//hbauSFpoYo
+FEjCq6h2kY+Tz4Z3T5s+L3Ip97/Cr2DWvxJYJApVQMY/N2DuLYxb504tbRcr8dY+BwWezTWZ9Tg
UcVF26rUeDDySu3M3FCTCGvQ2CL9Q0fBEBv6Vk54/AoEGKf6lGtYyZDfKZjyyFvhQxypkKSMNJun
x0GGXuR2DbGdAImTmgQ0jLCd+zyZNKO0WxyuvFgFwgl5tRhp823qrFNi0Q2M1uQgcVDixf4lGCXQ
fOXqDPH7hcKEwiSF/6jmZwsFvk6czVw+6ok9AEQ5Qm2vCd8abq7I0Johm4eOIOmmcLW9uo3kuF5+
RDTK0KrJWo9KmpUMFHCLRHR92I2nOkiacgpcLMMncjuhWm9c/W3Lko5XYrbQwQRujXuyj/BrwSwW
bvDAhyfAJnAbXZ5TzH4jcL4iyxx2HcET8efJFTYYTx/41m1ACke2RC6zBAQfqblPdqojs7Ilb2Cb
h7+B6nPdNHAVuhueWrxiHsZcn89veHaWTn+Bke+zddu8dGERdTtwSCFTqQVQXelaZ/iPKqj6kWJK
CUaSPoPxAkfdi94sAcfRRtDwHoiNaPYItfH45VqAtSCvSJaEueJGV54QGe8IsetPqhdWqdvsSKGw
9KpcJ6uC+51YZpCxO4aBwm3vcO/LRd06i9aIOYohfQEkp86fSC98mM1hMvhit1Yz4nC8HhKnHLDu
VFURLvZnTXjiXYUD8LT0xtJ9ky+Mdtt4+belsLZGa53m31b7T7+FbOYSCnpq2TdtJju8MfZu8SHw
OoEbdCmz5ZAavfu+lEBv/0XLr174B2/wLgx8ik0kwBI1c1Nxc2w+QIXKdsPctcVWvKThb8LFd/j2
uo9LwpGAXYAsQgmMthTlUeFMZs4iYbVnCJEa0JMARMQnDTGF9nSq6A5hPp6j708mIOx90nI8RzJu
9jv49F/G5cm4rKshUb1eOjUOgRo/mgG2meXD82yAxqcU28gHJNEHH3r2xSCqt/sG1DxUbdiVhCYg
9qfQyqeQ6AiATavZDA2PG7slLwMe35A9pa5W5iYGZNh6p0BjoxJCwxSIFdUWZ6K2gmet/6tluJjt
oCfmcafHiDVNRGwnxJBZ9yVrRIUdj42A/A7DJmylMogT2CKc7NnEqeXcE/fIFHuQ/8NXiqxtgXB5
oF518q7u0g3v+2IDI8naioKSM23sdXL7juKYCvbcoEmrriOfoqyZVWQaJ4HFKC29/FvKExgAQw+u
tigdK3mjH/91l58J2r0ucTEMUqn75/nyFvZLODKANYyKXuY7qvksjkpLcfLOkkCiF/prE/1BNDPt
ct3Y2O6jOM4l6b3WKIKNZ3tVZ/491ZX4UQavURu1otfCj65NYHFbaz6pvdEzYDN8OtVXaatOjJhE
H1uDvJ3l7R6lWEfMax2boy0HA/Y6ImZUHJ00ZW/m2rlMMI2EUXBNremdLzZzvKONJ1B/Vv8ppzOG
4Exynq/eS6xaROqNsdBfbGNusc4k1hNDdeoO9cbtiZqA9rQbempMIVIdR/LB7cdLemkpAVpMmuo3
exj0u85YSI2gzQ1JuQvOpvHHESc2vP0+e7lx8omQoupfRE7uDjIMgDsf0DlDLkI+QcZfzXkTlNHs
l8rIswTOkdfG8/8YTYdijC9b/iHpMALrOPj9IdKr4kAxNxi3niOPq2gt68kXplE1NKr/A3lM33eg
jo0otzRZczz+jOdELl4GmN3bdHeqXQR+QqLtTCq7UT3HnBGPSC5JE96OXZjo2MjAbfoeGDQSV+vc
yY6qxIdkOKwL+JiN32vUJS8s4DXNylF2XbRtJjmvTomIBjtCPxevWjaVcj1/rQ97R13xiY/0pCNc
vPa+3N2aaKcWubJm35EQJjbbxSK3no3/MJ7ENwE9U8FQ+Bj4tMZKdM8ulUDPqdGmE34P+z+9MvzK
Axx+dyEWqluhAzGd8W1VVONMM+eLbMxMS9g/5IY6VUz7bQDHK6CFNSY5H10egorKhfgmx+21sQW2
rr7fx5R4DhRq5IkJYALbV26X2n8Dh8OUWb8heoNvTKSyWReVBm17mSLftLobvR4ek6zF/swCzRuR
lM8eCFs+yOug/8WzBurNfjWWwoaxYSnNCMH9aFOkveJjP50P3CwnCTOgO9kDL9mYwQoIDGJ3WCgG
URkwwFcEaIcMV2LOx8U0RfQC3a4lj6DjqFkMCIGLDe9nnHo4GPgHnwICZDiAzSWpf/rZx3bBuwsO
14LPt23UlSW3uILnTblq97sjm3y2hWeHzYPuoP1UmFZ5IG2Kcb3oqTnepuwWyP5vKD88RYhbnVGo
F0d6oyT5oT8FF8eFPFSqvBR797pDU15H+rUBK8YostnL9ABCGNni6oENdQB6O6GVEfCYRBJDIUNO
7oI2LbPhhjQaPh2enCM3x+X4V8afWcmFAd1+XwtW/ESF4/8+qww1ZpWQeAsT+HpY4CrFZMO87FMO
w/SFlXywv1ZS972IhRKtm4Wbh4v5SeStDg9pIJuOXiTSkQJxEUY+apSFBS09FxnK0Buh6MOo3aS8
o1hVzrYpFPPFgaoOOcNCSzSgcnETyxyn5BKDJbt7pQUBfB8AnPOB//BKtq2+y7rzYM6dACyhWX4T
l4a2JQ3jZ+Es2mh8i4Ne35przsqhat/zRB4n2OHqm87Bx7E3fMYnKkFowYInfltKwf8f1YEp/swi
3iu0hD6IjrDEFcpI0jhdpOKc7xOds/xzbACZRUNkooqQvnb5AddcFhBCdg+3f63onXOb68qxIKDq
EcKgjs6E5VK0bSjFe+rPVfPWh0WE3xf+MnKFkesoV5TKgM4+KPZE6dfWf/KBL7halhwJgYD9xqdM
JIxM70sypv0o4j32du5qyqgdX4F6TTQKnnPq4SCeZAr2dxjREuxOndEHFRfSXyoC5yjkeKdkqFAU
svOM8jViE+oAJS6U7hPGVx2+AKnv9SR080TgThGVbdJhHvnMXsjm/pdTByw2EO8MuqRSnVyAMI/Y
TkM59wRAOjTC/dALZcb+Y/9LSvwNuTn3EHwsTNnBUn07qZuEEfrm5ehwpomlHQIHBxBRiLDPKaMW
B/EeyJJHIX1sO5ds6dnO37cfSGonCYjypAg8iVplxwv9XnRAUWcah712K0UCaOlhEUlLQs/U+Zt2
ucVK3b7tY2qeFPciI5Fc7RRLQqo3eKt5TePxMr8NU4topTa0OvTLk8jhYvByE7MWqMlgVV8tVJhr
yb+wmlmcKv2c5TSzAg0inpt/jPQd1KG5yjCHNM6+KsZ4GTCu0fpV+6okkaA7zzd3U/G8Dz9Q9pTQ
KGepGwYHt/UqYRrOMaG4iTELFgCbyNNmDj7Nad1MMN9Vea7lbVeG8BMLHb66hHty7y/6rLs2C+DW
lxLmMFWf5zxUzil60rtt0Ft8VelRUOWqMWSOj4yrQW5qT16eAxOoPbbQo1Rl9beZeV4OPLCdGI8Q
ARgwm5FqHYhhKDKD8GM1YAHfLlJQHiaVgvBsYZdD+yizCa5Ik6FP248fhe48C0m1XT5EVh0N8uC7
Lc4yizXFCDEPhZcu8vrvfeWonJ/P9HVDrgwl7NkEH5TIaS8VQSfnj64ddLQv9zmWj1NNUA8tfgWA
oMQwAUsjZk8gmLCNjv3kzTT4npUEHvLPv00h77S1qQup+V5SRH5P3DEc/ETkAch07Ehh6fKRFJvY
iwsWEXWbwrYNM0wF+eogusB3DRk/6++0ppUUC/yMyqRAHIQ6ZvMDUTmaGGoE7TFtnRmMcEah0gH+
JAQCU+2Xk4laB0ve+9+E8t2ikCatqpgFg6Fnv2FNK2DhfkYPXX210MDVlrczrEyl+CgC6/nPlVhx
3BmJgyNP+tGU5Gvp3ZSLQSPjnSo/c1QxxEE0poSb6ds00xN0OL9YmtgTsElTiYuqfbpQqB2bHmxH
Zt6nrfLaK8ZImm6JPp19F7zJBrh42yT46KH5Op9YFKGhG0hsFvWJX8eC4ODML9OvlmLBpkNHM4kL
KrBQfjdjJAaslWJQDSOW+rlesNuPznkt+bIMOYXamnXC3BAvjtf1bZFqOEk73rfs7kQaSRdPxo/3
2C6RjuU6gRGoiJA9kgCmkjADA2QFZCKqg+a8HSQL4a3+gO2qSRXdA004Xpy0JDD+ZzvbeVTdKW7W
hmVWIkaNf2ix2R3/MmEMnVEUuERlGe+4XHicU+90PIsG09zan8XU/4T3HAJoYVCfqr5a6iV9S6I5
jY962Q9YFEdex9h1c+lo0Oe+bMi0TRuW8wU9LUFGOk33FzcFEBAnBytgGVsz8BOoDQAtJTJSc5Bd
lkMKLx0Pjp2SBBoLEMytS2opxqlwYLVPSqbuqK2B5bgzGRlJc4Pwke9NHYE8DTo381flIMT9Lb4a
a1dhkVE1wgE0WbbiWRKbYHTpfyCqVDZ/qKlhnspHO1DFsBRKJfTTC3fFlndPPEd3j8FHCwF3jy5C
eCzPUx9Z6DvVR/fEsR+GEbhO2aCo50dDWh2NQ4tZLe0ABm0ws9YstvE8x6RIhDVA+YFVsnqGa0t3
DvmYQUV+dIZtO0xLeZRBn7FQI8G4PAjDpHRfh2DQsAABP59ltjR+DQsoqxQkdmuyxBqJaKODnpud
aKaFILaVwcD/9H7z7z7mScjOKiJvXSfcDFcxT5ZHw0sZXb/yKHI8msyPHc+hmr9DcQVlumKPPOVD
rCb/GAmpt0uPx3HvvrAH1A9CHLR6V/duNxGvgMrpV6xm98iOoEp5FgSOrXJ7TDspD61M66RILQmb
4jwzIyt93CV+En+u4yqV7OJbGX7GnDbD8nM9JXZFV7bh6nZ+W3mZQbMpdkYjcbdu9f0FWnTpP0RO
mVw1fntMN0cAyUOWOiiuza7fFL0ohr8RD1udWxU/7rBfi7nQB5ubfolqWzzeVz8PnIF34yc6glG0
lqIQb2/4Za7i02vDtzpGhRQASgM7zG6Uwd0OTH/NwJ+RV7bvkPooaUArqTI4uMk7ob3IxTvJVa1y
D0RriZ4OlenkE0ClffIPb3ZA7MuTgnWsfKcH7XiJiExpTeZ9+JydVA1Bz6i9JX+dwvDrunDqE3kq
BswMw6r2WDHB5eNl0oWM8CKwd7XPtb3D93Xdp4LYzbF7G9KVo0SUVwrthVYR+4yRTteisnVmGzZE
G92bRcawyQa9rQZpinoFREr1h2KzyDoexlzVMpmpzmRCYPl4adjnOgCntpoNzenikvi5yKUH0f+E
sIAAlVp1YBZ7YE+VlTQnRkdV/Ev9Vq8AoB1akfSZaE90TnJHAUtuu8ZWrG/vR5qmc6z+i5NW2S3+
dB0lfMevOGpAkmf85wMrBC1bhB18xFO08punEV3GVvPEXJzCKAYQ49qFepmH3qMQrwDFI2x8MSU2
t3JIMAUCkZf0zGs1wndJSLvhekPuwKDJLRjhZIIvNVMQ0NBagEFTJ2bmYDcSdXP48Bbb3pnALdWH
nXTegmcoQ/taAoH8oMExmr8jb8w9FRaGun0fDR5mr95k0l6/6IpcJNazjt7HGKInCygV7SnSMFfd
l2rMfw6NPzLANepJj11ZoQQhxttr2MchzbaL86WgmfGJq8jtGYoTveJDaix0Ge2nkvIOB9t7yMs6
Ehp4Vh8+3AMXg3OF66T3uX4F93RLhoD7wwWaVuNWqsu5LbqV0SmZNPja0AYAOx5arvDlVcjJpQ1i
sBdiPSZNpXo8Pg3VwyIGgcDKwAhYtkQQ1LuyG9NP5lwf/AvRqZaF1mSJ3wyvSkDOnQ4BcDSsVHT4
s0hs6Wg95yyuqdZXGBikV05HoT6BTpqgWM7wT21R2K7pvnSH3NFXGCNVgf/yewLAXybqjNixV8Yj
2UWqTB5EuLX3PcTHKSr3S5AkVeHqMIe/WlY4wam1l7RyMLxLivBOexM5Qa6F2TLURkAHDD5hu7N0
mw1xR2HF9JdrZjs4yNuIZBJoIYfESTv9WhJrM22IN4gDNzO4BKYpg0EdlAQZuTcjaJJU9VX8e7rb
GWBEfLMW9GrMtPshRtHVFD7yEofHssFEqE2OaFzWroW9BBcKKRdmVNxlgrZdNEfpqyCawG7IKY2/
jAVc6IwvYYdnBpIIcNRwosZNSFkt1NrOBfb15lPrSNGswhj20udFOjidOBes16ZcTDLFPe58RLNo
wV6f2vO5YFr5+fh+cGUiw2cGU64gI8yfLq22aTLy/u8XfogqOGv6luy5IYmztO1ZJryIK3Wqgos0
bqMlHtX7evj//EOds9g0TetY9s8ndKV9Z3FST6wzgBY+K7k7Xe3aKTOcT4N49nKYHzMpViVIOsEW
3dbn+QUPoBFg83ushInb4F9LDKIRIIqU1q06b9ov1IhgYqigYTbRdcBuLzC7hg0kV3w0WQolSr7Q
ihPRMOmMgarFCI121/cyQtLsscpEIC6R6vAYtgNM5WOsmfT5wgPwXPQfL5smJBK8fPHX8KCdqigM
VTrZvacK6tq8D/UuYWrqVs0iSe1/Ian9Xuc0p6jAY8hYhKOPAjQsK+ksfXBJNRoQKxyJQys1knZg
gqg7qYFEjGvSjQ7KPakLcF6fdIw2KCQU8Ohylnk5NTEda8dh6+HcVi5ylpz/gzMELH8kfkxoiTMd
lGVstOnGeA0pFUZp7tSMoRy1EOBAofYA59Tkfidmjr6r/bvmGt2D86121y0RivJntvSzZNCf96VX
QWP9A6UsPx2qp4z3Y2YVo6azxS1DhDvjCwXtDsC09r7orvw3oasIOQgZikm9wlicardfmIYLjROt
jIXnw0SjX4ddxyLe8tTCHuI3N7lE4PDToaxlFAw4v/W/RCZt2H8t67z+2tyh63IfpBJ5VIh1OPXj
kwghQJjpUbOs4t+ES9VgvXLuPk+BMpCCCtjg9ZOEAdG1C//Q7myD+X2qBkPT3TA8vQ/aBhnzORWT
HFMcvbJt7RYZfMRnGkojW0Klcr6T453uq8YK5VJ36YBSHctDsIQjThXgMsShwCm7JNaHRnZNIEP4
P0OzXf4GkvMDrDrJtx8gbu44ArdFanLavW4cfAGD0O7aCzmUZQc9oyJCi0soN5Je53T37BmQ60EK
W3Veu0ZqljcX54vrNxRV/XWoBwfC63GLXRj7q95xXd+xV9KQ2Rlrm3IRPHtOUdkE+Zy1F5TwMqi8
Iw3d7nnRhxGyZJTJXBPvU3mIMa4YXCAyn1P9TOBsDm3ved/FmUk7kDVSWtrI+cCkbD9g6erb3ss/
m7U6AaqCGtgORR4nCo9vESb6CSabzzkk097OuWPp9e/qHwciy/H5tLuKO5JDa6rvnB+tJsSJKrPB
xFaq/aN3tvDyahPWPzd5uRzXwfZ0qDGsVcstKMPdYerFg91MFHEXPWtuyLJYiP6cNN6hqoyzdreU
x0gLxe4CjVOg21U02ax3VSMzphvnPKOtzdbQU2PnJJP5DOVDDkbrlRD5zEFvniH4runoY8KtU5cx
jiR9t+96ngYvgo6lBopO6MSuIGuXq9yDAt/L4708DJlU7allpLeoD4EUFkRNzEAAnN7BiVCDe4us
j8AM/A8tVfE625lvhW8uzQpNchDRL4wi0qyLW1wad1AWzI8WyJ5AwPPKcg4+wPUADSSgmqC4BfKr
TlnXhN3PhxGX87hbaJ42XWH7n+eQaOA5/QuYx6x3uo1qr68b47iNiOb+2UOzisxijRKqbPqiTlYt
GNaKwLLwDNoRoAoxqP7LVaS0UenwfoHZOWEdroWh2auWV0G6foTmbLd1wP3Ztm5Stlm//C0E03CF
YXn7XXBUehD2UwDZLHsEXIb6OtBPkqaCJwRQ6qeIm9a5B9BfQgSQW97ZYulmU8TZGC0H+GmkVJP3
zMpqpIes++KjT4hhldyzcQTu+IzGdmSmo4FkFkBX6OUEbCAizwBQPbZYcXhs1YAZ2rPl6MCDiTfq
fj1fLnosAzYJbo8mHIX58OGj7Q/EzjbSVY6i7fPj2Qc8N0C82qe6yXhKvPj3VERlaJnUtMZWHqij
8L/IPAGwNiuLo3/Y8jKXutD/q5NHfByuHJdzZyhOEGADELoXY0i5QWtMPtJk9D9HzKgGIPWylKqJ
wXGwOU5b9PjdPCvHR42BjgLrQ4/Qp9FkTNGfchuVuBrKWvWVl0Yz30ID4ThNEJ6fVsWh13vPr0fZ
jDzQ52sxtHB9go73HI9YSIKUm1Ith/w2D1zsrqhheP4ayjT7qgZ+CzhocspQwM8kSVhC1PrkbXZe
I08yiOt5v0wR15NwvELCHeX4syrYYiwRfMYGd0NvQJ8KzuyqIJ9fxg2m4ULBT8DIXBWgYWPVvq8h
GSKKEHG6YsQZPP7pZGy/Cis8rMERfwRviS5TEDfBbAfi+MiJv7v5pOkMAHQRLU5kCkqXm7cCInQI
nU1CBioS+CAPuSJEFn9H5hOYHefDGyyMnTE/AzAjrkqiKLkrZ1cUgphzQqRM3pdiEpeCOsPClkvE
6sj4Zv6EICt5X9a7bmCJ5RCFiDQ9gekE0nrek5xdgpGVFiWD4Zw9IuMOas20fZ42q5vuS59i9dej
oFeoBuxMkZSivaIO9a6HfyrKJcH93xtyj2FfLmQZy0RsL9U0s8SdppVA/8Zb/DDJt/bY9QFWqvm3
xREuow2x2oOPPjoCoxrYHaRSo1E5IsE1VNDVc8NQuF+FqX+6k2gmd+9SWT8O6jrw8eKnaA196A/k
9HwgM3SVJU2Z+qnxHaKOeuyjyRbzOmMIavr0iAPyeOYSOmwXlNl1wgyLsqlp8VjvjcwUDyliU3/6
Vq9YIJ+AcSjiN8G0uU33injJsE3vgceXiJYt/HyzQ7hr0k7bu51pE+qkPBRj5/TsalY7SSCL/TcN
4cqeQtBB14lpT6LmMYH/U4b4+syqdTpiSXDaYnoY0r3ArwZpsjtkntbGl3uG5ZX3y/60LRiD55ed
lc4GPh5nE00XW4NURi/M/yYbrh+KLaGXkpsYEkrwidvjjkOt/YEnhtHx6XkoCXkApV8ZEQjC9gb1
mzLH3wsRLZciYI2zd3ahbxf0vKCH5Zp5/SKqY6eYgoa8AOX6CmxNbXu5Qrplxhp43QHudA/w/vaj
CrlSpo9LgX11C9/K4tQBnF6tLZzM/nRqZixXW4Ebdu5Rvn/Yz/dok5QIhmki63k40EuWaZNoJzo1
A8WsphFEIZJs58mKdOxe6HVMHfxdHiNG+yX9TpWBbbLtOk/LylEuzSY0T3I0G2VhygkrbiBr+4B8
kxbQYz0ZiIJw+ehjHdWjCbexA1IQuvoii1IXDR2Ya3feNPUelvB7+W5WWq1LLD+C2PkiW9Sp3KO7
1Erv5dsKEino+O7gPHbWTC+shddW6jOiN0ZxnfFGaY/18cmli3S+vNwoghGlkaCnXr5RUSCT9sxl
k0rbchHEtelTfCpCtoCpIo+Uxp4Zfo28cUwuZpCiK2FI1fXyxcSiJBQu88+afRzf/LbI0urlJYVf
Fxf3Db4HgHZzIGmx382qaoH8OrIkNi++SUzcOzXhXtzbdj5bamDHfGydWenmjUd7oydl9hzgQRJl
PCi1yDiHKueXbAhYX5soqjxe2Sh1+krOOzgcf4A7/q7rX/zpPLYVO7R7Cs2rwjn+pZSOvBwele3V
WTdMK0DBhCIs4WCRVoDRoBO7eSKiFh6dO7m9YoCfD15kn2ZgksGaKapXu2QD9Wriz8km3R+6yKb7
ngOUVbb4FdXeCB7Pvh5WYakAj6IYFObyWzBYPMSUzjR7oW1NNUICapBD4xM/mI/GqeXrLVP0nX2a
RUn1j3nMMAToI2hmUJRNiq4+JQOoCn864mBv5ExAkgpq1WQO+FwehZ5LuuLFTd/evmaSvAikHOoH
X8xLa/kS7wCMV18BNkrUhG858SKhlKtspzx1Adp4UWglx4U3uuoF8vFT8M5Jfirs1G5MxWLDBnZL
2l+2LoIfvAa0jWZ6vxhal5QT/KRNzspU8Qs87RUoYcjWtQS76lA1Z+R9zxkhxy7V+VglkqrmVrUH
0plJfDv1Nx/ERHOH1lQy1mSuH/3j6hiF5Rj9ViZubxzDGc9Y3A4nm3Isx/YPsEJvJjEA6ZFlLano
FU/bYs9n1CIhUc4hTnCKvQyAlNvMcN8fArI3Iz2Cc/JpOA4+q9bdi5UY/F1HMgssEo414Ypf+DuV
FrrjKGE1y7RnxZCbk/zMewmCKOzTMLY+p/+DChgxt/KsD0+ZUBVj42vqrlp7AcXYt6Oe44N2fxgR
TOg9YiFevqksQ2s4G+UmO2crqtCJzxlY1UP96KX1/nSb7sKAdPS8IQu2H7yhztRaYli2w2bd696O
EPQpNQEGhsZFale73818T+3NFyB60gyvvYGPqknXylZ+LBYin6L6dXqNVdSOBnFcCUIqvf+ZWbGq
/QhiVzMW1cizyjzh0VQs6Drt87DhYJ88g17pA2vwUnxl2SYnsBynJtn8jmMXuFX1FXbG3kJacBUj
r8Zdba20aZzvtFsebNnpKGZmvO3C3fUCeOHr10s7IoWDgliCMZcOpgZsWMhk4V5DXeryGJRMs2Q4
voWQIlWd6Xygvgabm0jGoe1GzCd+eI2y6k3yuxVhCJ8wc8TnHH3HZdaSn0pNz4c8WHoSrT9oT3z2
9KvAMWLApc0DBsvIA0IrG2Ft/8JkMe2aYMGKKJbTRkem118xfo3l6NUea8Pt/ofhFfSkXVYx2F7m
LhAe0xkWAqYpCeLndvVS6IWbhzTg1qMhWewgTfM8Zjn3cMRArw+Auypj9wDfcTMHlCt2TdPKr0sV
SayeDK0nr2h2np+xNVOAnyKU1uW8GvgzZ14aLTwM//RQO/+fQ32Nit86FFNRN6GNQy3dAtuk14iH
QK9n6Rn+86U5CRTQNhToNuBogmYCXxefZwPq0wj+ionjeUmmAmDaEBoa4pYjd+YY4isnERheyUJC
HJLolQKcSFxCDL0ENxggjNm6bYNmJ1jfxv8UJA5vihTvpcnD0NugFY8/MdGF+hUIYYlFO9gIkNN2
NpkFJR++NXBwPIGBAxiQFnVZHDsgFhUevHSK/QIuUYt4tH57zfRDFz9oWYGetOE7mw+nifalLJsq
ae/A3edULALID2WtJcrVoyvK+VidxdW/QWRySyRADXqffAYodELogSY41F9XxdlWoWBfITwWgIvw
D2CDu+eDk3YHqRI38OMHyMjrdvJjj8u0lr3SCO3eMDZtt192LeAaL0gLTZYmdiuY5kS58GVbazHw
e4WCFZ7D7hSRAL4Lut3unvcHlYPGyzMH6rF/dX/YwUedE3QKuQ/fFj680/km1Rw+gv0TZfboSqOA
+q/7D5kIUc6Hu04Pxbs9Sv+iUc2eu4yDIYWbIRwUiYHBNnzhDNHKiOgoVW0R0pbiFnG2sX8Md3/B
ZMjcskbfIbUB+fwfxAGTbBZs8MtlzDqRV8/VTChNyB9qkHVMqyCs9X6pqdnfuVAO/7e6ruCp2sD4
ESSCqpeK6wpeGzD6vH+t/ct/tVBYwbv5Bn1enjpMG6fzbGdFJCTxa7i289g9h/Dwya9ie1SPia6n
QtCeW/+yOOp2i77MmRkvIR/jPO4fPTx24JvG3jeMHf5SP+FGAIRIjiGW0ZzoCSJXNzRXfq9cTpYh
s8D9HqLzKoEj6ZZTBR1YGVT47x1Jmt/y1z2CF4plyr8WvB4qZbpQ8+NKjbap2/CN3o0cGeT6J3Y8
OVEaiwsqe5OR00VWofdRkXCIOEsKDHJGx6KJCaFyHcYj1jk8TcCO90QZhkGzzziJBJs9hJaQ4VYt
WyIUxwYMX5CGW6TgaXxQcSk3LsgPebqeD+9ccWWtPdjkKlzn7pdn+IATMKQIyElh2KiYgKVhCzSy
p4u412A78sPdUhkpjpNO/DHZ0yka2gD0ERUYQ05Jv1ZZ1fe8iHzOgpEz6IBxkaNLGRYZwKMOdjZ9
MOh05Dg0fQx2nJj5VQpDEkl01gWCqvs2yN6UawRBKIu3TO86lXecHy+E6bUXFKEu2xrDQT4kPkOK
4hxe3icjjRDPQcvp9onYjrTAAML4/d/92qB0S7xkpisFEGQCysC4FbgT3Esi3dt1oJ2ZmmaU2sZs
hgK/fghjOFcuv4P+2Yv6e3IQm4Ufwva1PpiteAEpLVBMROQCUz8dkQ0ZxHdXCnsasQC6tqR7pFel
9HF3gBIe+JKzXRpGhwFeGa7qTtG9Bd6vt4i7/YuSj9Cv4/tp7stwem2LHF7VAZSttu+YH2hBB8Gn
i6WYLpDZUgtzs1eUeQY4HwdXUBuB0ZdNv8ee16Pcr+J1FNIBB2Y0hXtueNrPoquRHY9XH9q5eh2r
YKNCwgX+fWGtskgRPNzLq5Lm32tKUV5ag3HyZzZR1vbg3ATcVJwuxESVbuD/kymUtjSQ/8uPJ8Ac
RXcDXwVSMf5tqydiMhLaxwhgml6ccRDbsQDsGdWKKPIK8ChDiaRegfxyrV2dD1JvWlusZXIv7eqB
SULEnn48Qs+0xK40vtHHLcbb6mYYd+fM8l64oI1jj3SzK24lMRWZixqCKiDJc7BDOuqgCOV3iSye
FjzydoPe6GUSsjbe2GrLPYoFmSdgvt3X3REQLjxGuzrwsdtMUBi2FCyjp6VJc7lW6CWAGulGoitN
z7OIvsRbhhTqs7QEtXANWt3EjVdvVZOoDuUAp+KtURDFbAsTQj/L4OdcYbcnfThqvEXkMWSP5eg9
QhR7UIHoXm08FaIrL/9UFOyyrzZ3s1fjRuY4kVEKoZuzCR8bGYVBuf+eOXq108wZvV8FHYhwID0U
9JwDtds3zxru3wIKVGyH2z+BrCCcVM+HGB7hGB2sfk1jIJ0LWAcX9JVvt+kBKBBescyMUSvbQseL
MCLyWHwDiQRrsBAW/lp6UTz78V5rWv8tz+xZwGkniN44N/1AfOk0rmatCysmNgzLPDAsuICx2gjd
8pfsI4oHh9J5nTHFw4ErxV51KFPfA6F0jib4TaE47lYY5ClVTIDKH4eP6EDb7WzL3073zALuqJPZ
ywIwlpwJodQ/e5pfBaDU6geHTc+hp6tmSqx/+kMgYOSDu3zW9X9lDSqos2e6WU04PHj0vH/uOHQa
UifIRh6re8ezItzRTiE3cZG52KfqjHvx6Z3oR+NMtnst9LUffKjXxS2B2nKVUj8ZCJD4eJcn9hLF
GZF687UpnuyAYd4IOG/yZDdS47H25M88hjNYQR27HPwPhDdawDUT7fNVbJOKG0dMIvtvbGp42un9
WEnUM6WQcMaTMU2RkygUIxjhxGNp1SKTOf4fs+FCrrrGXndybAUgmyyA0abYaVuSK0RalN5fUu3x
vMeXCNV3z7xqwXqz+dPQQXTURHtfT1maikvH/YVPtT04Km2f0isHMFITMMw3CjR5thHZK4xLWF5o
s8l+PruNfMDtpedyW9qva2mSssEB4BEUpB2KE3ZMORSXJqi/l28QCjqlRUjkQkCs+WKz6S6IKtB9
M14moOgyihgTo9MzLIH5KBpvOfxzPnGEtEIFqjyqmXvJCihdZ9CE3hh+FPsL3nNgnggvFr490NBH
p3G5FAwPN1J9G0fm3atFd+P5muGtslHSKshL461M0emUzQQPe3WqDP65+I9MHrP/OT8ySvhOByYK
V9r/EIODTebZ0AP6LLIVvtvxFRCeEPHNSu9/IoPFT9YZfUff5kqy7+blIvNvWQRToc0tPr7pgMbI
QZGpHd2iyRf3fNvxkrtFhHdf7ikxT41zgPK0rHnxEaW1iX3Eye5ly08YPutMAFGrONK9IVhIo96y
ECVv8MJKaV+HW25FO5zOSSwN8eAoX5W0e5ASId+vUPDtUsVPlZsQ1grnBPiaxQ9tdx3ygP4SK5Oc
GVURp+8pVAp2Z4yJ9BWxeVpWa7L2vpQxNExZRIjKzMQETTJF+uzgFxbBi7b6KJNADSEUD5S3R7EF
UBjTsXiKZt1JGShGGPnrZH8O3R6r1aPXIcAtWl8TG3KhXVxKMNJKdLtsfl5P3eE1l1KRR8ZjsgNf
ORwntaIAnplPbzpjf/VFMEjidurzB5Bd+Xkjy0XEDSqhVh9KXnlYEhs1u3H9olh7HqGUq7uqTOWF
icsDaKhdoGobdaEEmFbx5Em+pA2wDuUSh1eLERTx3OEhXhXWDvUZX9klXc1Kx27CYZjzg2LzARBz
g3JPcZFrdEo818E5XA/0PGZvtZogxuEcPimF/jTp8e/G+rMFwul+po1v4FPOv7swQC8yjiXAIiKX
4iB51hIdIA1MRhdDxACpkALLMuyUM8KsolSi+YN2E96beiV5nWKHIAY8yPsU326C7nU/wzsHRrqG
T9bTm4iBevJW3LodmBYvfPfbp8cgKt8Yn3h7xOC0KNrCliTbxOIPbGFcYDtcSrqq80iX274tt7nZ
M428LCFbupgAw6h/upa0n0H3L0Gwmb60/3JWNUW7/g1pSS3Z7mG5RIhRR8/SCfulf88bZl6ulZLG
AVyigHRS+7eb/fugW+3qRVB9PhcTmH3PY6es6NpTl1TjVCPB70VntPz/h/t2fz16lih6LK9VyOHE
D8bHVhMXt7ickI/HXiLwrSKZOfJWdbucNXNZ3FPFxqbeYoKIgfg6nEyiOhli9tWzlibo8caJqz5z
zvCYjdKJmjud6U7KN4G5/fgxXLaMIVH57g3TGEGFsEud5NhEWdVU865ztVpd/yh3IU413iQNEg+3
vxKoL0p6XxtX++rqbKXn2z5NdaMjUWwSH1JQiMYzdvVtJXhPNIUrBcK1SkUVLPMomMm1fcexMplE
08lx+dk+w2EtXwi+BaOAZBguhrtPG/i5M1YOVbKju78PMHSsUdtbDRPmhPaFx1k0gUp5Z8ivlCzY
Gq+7090KUeJhiLYZhoGz0Kiir+oLTl0yePxjV2IuAWdnhyt/sLhZsOQkHR1VyPwIT03FcuLqRAoW
TwTQpH8Zv644HY/sgyijCanPVcuTdeB/MyAWuUnxXbl7tLR32A+45ODQqfz7Pr2obV8YfPINOEA2
9t1UzNS11eWsTFKC9gXsiNGu1ZrNCdjbtboMJc1iODcSyBD0rjB8a6dc0Ik+HPG2goT3l1ca73DX
HHbl0GT8Zh2t9Rb7rqA0o6RHBt1sMlo/+lmKKuv9IllQwdwQNl6FSn5dfnnuYh7xl4h/URLf8jGW
ozKbxsNBQ3hcr1Zg22c041XX1atbAK2TJg0EhqIVZ4L7cCaaftrpDsZamryx/EBS6N64XqYC0x7J
s5vwE2jkL9eQXMx2EivVANBiqLsRnrxlKMEzqS26n3C/0DlbY34rj1pCjzufMdyShYcIvOMd1Sxb
u3PjegRO6TzqN4Rirc2MiEbQcNzskUrGH3Km0SqQJkZeOgbNa/hCi+K7zfCOB/rWR+UnS7J9IFGQ
F9E4dX6XBf0h9p/DPaGKwEO9/ZaRxssuc38A8u5kcjf3YG3KDiAZpYODw0uhtHWKoEjm8zQZx1/m
9bc+DdxaCiN8SFqKuJEmHFeg/vcO9JRr3/TgPa6AcAZdNEiKImecK8FngJ7wbSrlR6C5zXBBAlHY
TAi7GMkpjaD7/Urxbsos5Nblp8/83b1JpXfW3L/GlIleqeH/CNN/PImEF7+eUqLjJyb0jC1zZ6xv
FiEMpLN0NOG0hYY4DnzNvzeS8KnT/6FwVDhEEUGbGUjXdFReXF04C2BG6pCkhLL09PkjHPjAg5Ef
yrMR77dQR/trMeKAjK3EQ1cdJGg56r4DmQC7W67UGZOI2bva/JTCTnxKctu8aK45CKuqQmxw80sy
4GCfA27hQAfqr3PYgZEr4KHoU/Lo9i7ieaqlL+1LpJgxkdEseAwNomCg3WFb+VBvq0woTTrRzkH9
nT+7ZiEz9171oi3WUweBaUBr0ThQZ5EaYg9I+hqqXw+niqV8r/DOVGdGw6+yGqljT7nC8Z4p5UYm
dcJscQ0wg7MyPj+r3S6qLth8zyNy/SV1rpbiGuG5YuRDwA==
`protect end_protected
