`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
agkIpTKiEkn6Vg7jMxvODNll0722vEvnLaHOVLhPNMerkHUe52uwESqtfMcCMhDybWJt6BkiBMSu
EryWyeQzNbmc3RzwZsOXOYjzSTo3QLxNJkzgZhedgms1evyC5xrzhMd98dzClN/msiqKbFZc+fJJ
ZXhQqmEgBXjusVrmaauibYaipHqi0ckBba0qIo+o4uBxk+hVN81xRAj7DdNsqDokx/6Kw0r0kEGy
1iLxUM/R0deOiht4Kxto1TszbFNv8/Oowdu8x9llpFH+07xTzieKbM1gLhO8CKUKX5f8cptbVRLj
57fro6s67nwOH/oTXZQDD5zB1UrTzpREcqMLpw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="ehSzIFP3EuFfMPMwGx7ISHQe0qXgbzPJTsf4gHrfhOM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3600)
`protect data_block
7uL5LDO59u02Hv/PBqphb+SNCta0HC1EkVcQiv7hcH4t1hdVTilKHKqItoTa2U1i8kfgh9ziI9It
IOkfQqZzmBblRyKC6dNnkuT/nphG+bjKerQh5b9vbqN54u4CSBt0js800chI/cjWpr7jje3scy9Z
wvrLYmCzdyk2wCDLybdUcFDd9EJn6aDEUN9t5VCLAOWeerLNIsskFZ6XEs5Ggqqp1kxHdmAHJsnU
duhOXACFQruUnnmDs5EZEzcX9aA4dOmMsOVy0XsjKQ8Rf5iUq/anqBp1Iwgr48e4mbHH7vSqWda/
vHYXmxHYMDVJ4KBpsXMq6zohdDnvem5zEiH/r2qKnBEfFDnmXFpBACxhebpgtrR9IcQegY9GVKDZ
HqTGPQw/XtzibTErXr9OR4tB6ksC6A1SodCaEZFVaLo4WETPYyrr7vFWn/1D2sx4ej0c3E5TeCYF
diVEw6/JT8+qbDN5DXhiac+5Z9v8H/xHkd49oXL9L5JQ9zQI9gtFFYxHZUG8PyufSNdJ3RJuMRCU
/pWlpIs8etEo9yBY0F+OAAtbmaUnx33j/rnm0L93u0o3dt6Jwl1hjq/5iRspvCjHwyf03OH+XZC5
mW+zmUlE4sMY2F+dfmzs31WfTto8hGV32BVUa602a8DUaiDAm1j9P01Vqg/RDYJQDZaUUzCZpgP/
hrqCOESJSh1l2RpAQTQQT+ruYixdrj6aqwMcg5puD46kgYe+lU5c2ARU5WvXlnebwE7Yb/YwWEDy
luTgChdVm5JOnk1RBTNk0cw8XAgxl3K7DoDOV5LMsfDJY5HE3DsLXnz8ze3cCTjMwKNmKQ544THk
t8Do/qIdKEBcUX+oWeJrtgYvuMN8/wczSfkkR3LP8hjuZMRy/IlqBKBC5B5Yt5LTyu52Sw7YpX9g
Stjc2WspVNzc9uYlbKOwYRKKwyOcp95/SYw07NGDgCoyXbyM8A+wuzr+D2QIwPp806MLZ1NyAlNk
badPbwiO0bVknAirpaEehpHrXPERsRIwn0Jh9qCNDy8XjaoRworMB1sSmgwypWBUWTlWUcs5EHRQ
nBCxhz/51SBVowL96HdRDhb4za8KNDVcD+z9c0ckJ1BSh+O259NrrLFAbCq6i8e0nbNprKWQNj1W
8qH2okudI8CCWNuzWv4DK6JMLWkI+jT/kJJodCnC9uAhDNyt5pIqyI0+V7CTg41iZU8GsOSgnR07
p5GPC8wDrgo2qgO6WwDve+D1lLNnkSTVLBp0OHDo8fGCay4sXz8/0S/km24W7FcnjB0MpGeZaYKt
PfqC4ekj4NrUcmADt979r6WX7MCQx0IaC90+UzCpLZKmNsmucmginOmvnx6kLrsa1LMEguzK+I7I
V82Dp/BizgOhPiSHq1G5Q+KQnmkD7lJr1Bck5phzf4ks6ZyHsZ0p+J7pif2Gl1A6yyL+MpSATNVG
JwT+m/qKYvghyVOa+VDO8wvUhnYCS1NB/9H8D7HScYyl3nygHIBhIkZquxvaDvqEnw+QmEpamHBd
Inrv/Gnn2VGuAQUVgNiaOKA6dAwtjfJDwQpf9Z2dhksaM09plljSQejaSOa1q520dPLvapkZf/yK
MZAcz+6++vlDum3yLu/J3vigFRM/+4e0Ph+90JQuZ2Cw2pqJ2MXTk48Szdyc6owaVXtJPVzrM6D9
M6JuwTUf08rU5vsI28Bx1K3Z0/HU14wXa5Y+ZRJnCgbkKoYZX7doBpcrbIfpNwlWrz9MRwvk6c8v
LrTdb+dAAc5fWDhiVoUh5tFZxGX36fNZdhsZTCYEO9bEIFwGIMIDTKRV6Oaq74oXRO31xirEvxFs
DCu29VO4Pqaw1EZEwtRFzZL8h08r60n28aRE4zviTcjRYF8W97+di8XcFhxVm96Dp2u36G6nK3y5
b4LzZdX+/MMzMnf0LOSBmtFapps43GZgOHotI3ZfyXP35M1wilw7PIdapTwi3ULHftN+7YSP8WFC
Lq1SjQfsM1VGh+w6penmE2fF0lbnmYoSP3QB14FGeuREDxj1JXSQL6KCFFl0ry/cn/8r4gLyC+kI
JPk78ZUM8TJwj9Kj7GHwhSSokelHooTdIlx3jfqYJZDXaxF1XGsI7xqKx0z46EoMJFH6PkALlv9f
WpaXloK8TrSZvXF/RiLK0cUZjIogwkvIdMErr446hMTLfLDEzB+1yBXH5WlSaRgLFUYR+v08IC0K
czCaMlxEKpaLPo6OFmuXfRXeIPhe9kYOzdtJlfa2xbxQgFA9aL1xmtLjwt+FyOwAVmR2+E/lH80p
3K+T1Sy5mpSxS1MH3Pq0Zvu361Wv3izJrHvxmHPF398im+2nkQTRH6VRp+CxIq24289BPtnnDDo8
4YOh1vpu1iJCnroW0UdkJPN4IDiELmGUPpjZSFT2CJeex8Komv4e6ovyofw710eL9ao9CBjP8LTs
hjhO4LolYTrIdHOoO77y4abOY95reM8oEAG2eMOgs2K4PmtEMysdD5IOmcj/M0cM5oZeHpyBPS1Z
rDhWv5nhVWmsxCgXFtHLG+7M0n82A+56Dk4pswW0wANTWGbeSCaw6TcfofF/bGHRteQqsXzHXz0x
cbl11ias5dkuyxWvRnJmfY5Tg5Z61Jqswm8hRLnWt/XY07JZyoRiFwNKRay/BMTm+gV6v1hp2c9k
GpI3E7lc8ckZFO45MzX+BXx1DmZx6LnGSUDYyDXTCdwJT8MBL2zwjwXlsFZanyIjxSi+KT3h8DXn
SdGXi6v9ECtLf5VvwBNmuqZ61nVKagAdwRuXa12h+3GY39XTG24oUnRGGYVqMVnCRVeRIcwWRPEx
1C4ji6y/W93GSDsmII+U71XEJ74dFQabUN2wFvgmiD7Kzs3VStR7x2y9uiVhZKyZyc4qM5wBhATP
7QPsSopIwlKdJ1efYY8xLnuMuenTMCWz/0J2Y64nu7fJlYBqhquT7bawzkUA9kRVn7ECYT8s8sHZ
g2+mX20zrsl8aRz6mPSyt22UoFFCU70ErTJ81tc9Y15Adr9BXBR+j6KeIRjM6R0nH3p3YH4PYfc6
m2Vq1AOpPEc7q1A51tqQXIzHKSCwm9332sn7wPuflt/a+/AtHN9h/q06crg1I4DFOo1bVfBuWxwl
uXHRmSjcBqZArDWbWeS/gtHAsj2TO22wy7y7LgNAhSuLGh4at0yDNFVsHWM6NBZ9N3ZLAZxW8Cp0
OSVwv89EcszBHX5/WCUAjf+9oaDfFJJ/rTaPJFOz6EaHScHcmyh4b7YQyXqT633tkFL5wKpcx9V2
l8BbIJIU0F4GgU+s+KdHAUzfUuUFDswJPeLBZ6f9J2b/0vqoNI4RaCQIMdMgFo9fFAtXyLYvuqXM
uVyVZf2H4zjgdPIlKMEXcbEXAYnXro9BtO9JdhonEWwOM9x4FdRRwxkCB2Nchur/Z70QM7L9XM0j
l5Zzh6g63CKjf+IwlMNheqY7sC5BpkVTnNpxsMZN++fTnpVfYGhdLsVKgfKK7xRCF6Smrwb8HnBu
CUpKzyllhltEmRUtPyeHnHEE097YJRrnrcWAg9FqjBhhJ4FE4qhu95RFL8CoaBzdC+zov9LFPG0Z
UZwfHmClJ/MF7j/WL2ZlN6vMFbYRd0halDUCNBBqns6azJCJn22HJTUMnhtCXiEDPmXOYEmxIqzD
cu2xfZdP+4+Uxgu+hGIvNdEOuhvHw6BsaMVphBrmfPue5W9ZAD497PuhN3gvosIo4RugBn8bmoMn
mEdhcAn4m6oq7H/d1iikx0dliX/ia0efH1vdqPF8SHl1h7Lvf7BVWL77OhQ8MTiHVKQH988Fxw0Z
8Oz1yI1nGuOU5kPlLzWEKOnTXRDysKzyHyrG0qMF7Sf1mJMh/Rk0AkIN/hbCKv+FEctRDf58NpfR
1uQ70AZbRkOySLSA1EI+HD+zG924begHWFDzYIYQtjR5Cc2MPMRPpqkOc6sHrGC9g/hU3tcnKq9c
CJ4Z/6UMZbVeKy2sU6K1Sh3bAd+mNWNLZJP2hc1XjFh4rvrWtg6lD/+0azBOwrvBrKkGSuoWL785
pkroqXzknxbQLbbNbgAuILMC2OMefjpp31KhdSRJNu4xaxoDp5HL6ezEqBn0qk7ZQqp633N2kQxr
3RR53MBBMFMk+kvp11MiNogL0tg6LAZ5g/reNAc8EGz4xpYtPtd9NnUUO+rRl67KC6wp50FM8yEM
1JXMEbc1lz3fOd9AoSVj6rVFL7a7ajt8KjyU2FiPov9pPAX8p7TsrsJnBlnyiQ05cmsDAkgmFE5R
cQZv9MujvsJjypQdiYGkTivCuYPmi5QWDbPnU7LPGl/f00hXoz1enEKpm2JtdKkb/9z4Ti6CGh16
quKJLdW8Gu07NoY9oCDpQnkWvktWNXE0vknwN+AbNwzKFacSX/uPK8DWPidBT8vGQvnK6eq4jdxd
tifo6nlKYut58+sTpDQy4OeXIFYkldvt0tTcib3vdKi+6991rH8gJwWlZpHJY1p6GwWJn0bNRUGO
ApJ9r07TKcqGZolRXHqtOuUztMGou17nOfTGFchRzIF3BOZj9wgUTT68JBvtbnj2oHkSX28XqdY6
2mxAlIT4E3zfoMQ4PZvb+T+ZVYtgMcCFvm2f527tEQ2cxzOO6/AleP1VtPsk6fqAgpTfp8sdHY5l
aUCBTZSJrIyZyrG/YqCUfB70d7vCSUVyyIRwPGGVfnuqHFEpi00QFE6hDoEAGelGHUZijKNg1Ugi
b4Jhjza3oqBe47vi3TXaKrPEgOcF0TUWD6ClKt6wiiISMpqDygmsuiCy4zqnxrYJoCytnyBoEQu5
Hypft9cycJR+
`protect end_protected
