`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
Hus2xY1miDCUMy99QNdE8H795bnEX3b4PkzCJ28oVw8xJoriQg4ds2YMU+caykHOkN023f3O06dC
e2BxdQq/4oQ9XgZa97S3FUNzMHMlGJxQJgO5L2SHbh7UEDwFhfTmrsAHSk73DtHN+489USpKEKyI
Vs+jQB4wE7AaQcn+m+GOEhxp4pzzxe+NjHipy3GqiU5ShPtFySC22Hs0PvVne0R++/dBKTvnl/Bk
CVwPL9OGA9MlMw67lL/2lv3aF3NITPwB7vadXaaocVkcSs4Bvu5srS8aRgsZMZz7tyO2l+Ap/QIV
OXENzNOxjY/whrOMeAhpQ4m5U9WAE6dcT+yLGA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="V03EO9fPDxVlQiQc4PqTCmPiPQOgDr8SCoSduYPb49I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
vo7OX25xUNAxxGzlrW8szKJ4Ajm58oB6MqvPdN2XOLJ1/aom8gT0h2NPoEFz+VCj32CXkFl+Za6C
GObywGk81IePJut4/a1JJKr/RmlXpb95TeX5+JY6X+9SaewDKc9jkkvIW0zQAOBW+5EN+tOZD4tN
bwI4XHKiaE0W972YdSD/wub2gCn1NX+bSiOsu6KTFCvxKNC/qIEQmI8oUhbfZ9VogyQtrAqjzkrH
8A2PkYykNlsWfvPjM//PA7DfGR6+InAu/l/41URq1TcfGmAFQrFEqXj+lgG6YH+K/P5rxiUTzpUq
sq836DIcRMEEABMmncA3i995nHR0Ckv9IaacRsrhXyPyqukPRFf2qDBu+Lp6fc2wnSAunUZGhn7W
3FWoPcxZHAIkSBNJg3smwKN53tqUM+x5Iu3E3quJpO7xUgpXBJKl3VRa3touzwy/S8JpjChLAGWA
23fyPABopI1wwBL/fyug6PzDe7A1prpWAB9HGZJtFh6EynrWRY6aVvQuvYe0LEqEfNLitmIcRmkR
HZ3dYxW9DAS/Mbt2SFaG2ifn5qT0b4NPhcnniyeCk1sQ/zWTyhlcuyCL07fF1CiR25L2Gu+wVVxj
xmonKbl3geiGFWwsLPMFbWxy4cxgjsxSWpQMJ5TxTfSqN7Xdcgh6cZXIxn3s6chWybFPvrDla9kE
OC6J5NZTLfABkHP6gdvJlGDR/Lp9hfnlzS9NNg8Ovgqmoy/1wEzdLpkXROzun5IaVMoC5ECsAKY9
C2MP8SngegNVPJk6PCjDn0M19vYdaCOwCLvSxsT3raXRCMqciH+3qIsK4uesDM5CduxsZRAbSpuL
PV9SMn0cSAYhgcpe+poOt/Px++/sSs0RaVKwExBfMVMtaOSdpV9JzimeorMmVnj/8aVcQ/MiB09Q
WfTpvXMOpIijhKca/q6zuuiJWmdGQnBYBBw3QsyF+2S9sJlTJv/hYDXmmyYBQCtS8QAJmnH2ULlk
KcsDK+beAPSYPgz29pdoLj1NviiJ3qcEoX5QL8N5+jAch+0ryMyBd8lsVLHXVCnYwlm8GwUTxckH
Jhju8ZnlZ+N8n4eIrI7PHhsvm9xW0Y4CHYRdfRsElkoCL4cjNAkOnYVitWpq9Vvm5SBBJ6dDXS5x
zLqOZMleySYiN4JmPyVvaoJrF8hwZdAy0Qc7ZVYvnFUN0RCyNmpbFj8LIkuqhAzKf4WxzQ1+4EoD
STfbb8pei6cv9GAlC5dxL6tN+bWXrsx1uW8w/Tx/JTQuatdqNmErThtNbhm/WWq9WTix1y715bFW
YjzgAhX9Joj/sxRVaKY5bPAK+tCtqfoZ6d1id8IRzxbX9hQs7eO5u/y+zbdazYLBOh5syXG6a9ac
1p2QojKF5fNc0mK6eu2u7MyYl1VLioWX5cR8NHHdtz060/14i+0yGEsm9c1GfzL39l/PclmFpVqC
rtJ8o86ma4H76xuUBnd8hP2pgRakB63O5jJp8pbJlAgWvfZjJwBf/0hVxqWGDYRPs8jS6wqmPlKH
v06ImECOSd2/qsuJnpmvG8tBbd8Xt2nxYyd66rqMsk2tj0RwUQcK9b4YTX9nbQ0+6zsUA9+uZRNL
ip12AVm2IRo8mzy900wMEn4wgG8mk1qbmd3uRhPfVTDTcj0ORGFDe6jZsi5bW8vt6wMuUrQnQ6K0
nL1nbaX5MyaoT5a0wKTQpjdxRp+BG2uy5Vsk0Iz3Z1X7cRq3ImRmqD0fx6Hz8T73A7T9QEDRCNkX
hHY+IFVIvKAd8RQkrjLCO+fEEx1qrZNBObV5fk9wHhnqkHfecSfdoFYq2yhn2PBf3hhSjaQoVCwW
+cVDwY0FWIAJXnBN7meiNDWi6Ue+FZl3j/nMFVHC9JL+Jw01IkWgabd70m/mI6dEirlUUo0I+QDp
fRePxyjnNgST2S9ps/6vQ4xoqyPKG42YogRmvDMKfcQXpofpUa8vl6MhG1LmFKkyCVhIQFejrMZS
Grm+6QWi+q1qPsPWsHyrTScyMGMH09wWaY/BvyFI51IUcKrvOgXKuzPdGkDROrW6c++KrjagnWAj
Y00kENK87/WYpNkj9C3DcB3cOzzAtjUDxlZ+QvyWxfO78Bp9m4NLA9cu+9Sh
`protect end_protected
