`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
U7kcAd6i/G44+X5bUvJr10ulJu2AhuIWXdrKiQhQej2p6/zlMMGulo0Smb4DpAow2IkxBTsb5r3g
FoBWaqwMP38B7PQaP/S0nps/pKYsbeP6fu7+3QW0DDDbnfwY3RV4vjBD3Fr7qkzzBirLV+5iXZtr
05/ax2aX0xgS2NJ9ybM+at2txY7IbdW2WSAFV+j4xDo1BV82XflOuXx8hJtJM0e1gfHcccHdXZwO
BEDE3vLeuiQVOxkFvrVm91gBbra0VopLNq8qmSRwR4hw7RPmFSi2+g1/Mf0roWdfM2NM4MwyKbft
VHtSyHknWxROLtz+p28E+khgUglaPLUdJdGjkfoyJgv+IS9+fAzq6TRqQcPCIckdstTt2izAKuoi
/7tNo6JmxWsdX0H5N7nVoDEpmF1e94N80ZjSWs18EyI4DAxCtXA4WNH09Rx1ZNrkk3fZ6U7t1An+
qyKsSSIK6N/UIfP04h/kRTyYob2HTkRtotMHJhRUBShwlbVZFRMznFWkwlVUZIU68mgngsUGoL9T
Juf+I7Lt+anHRkdGfPJ4RoHLzYIOph8aqGkHCdMZr7kkFEEchFLQ7GdP1/DvfrovTlh7wiV2ixCc
kMrbNT/XikFGCz6U6MG9A/oVUYEQcQVS3akTv43zs9E+DTHQIry+9gg+c7K7Po5n+a1nB9pcIZIh
9U2hIbv+niUJkfB4Iaj5MGw5zkZ8Y3SER5yd+suNbhzhAhRNrpz9LZA7DXrvk7feOkcFI2oJicje
B/MNYYqM3ypuwdUEf/r2XcypEnE2lnpP/Q7qxKM7XU62jYNh0MqxMBcTPVTFrecZw812qgW8+66U
oZjv+If7G4vrxfh2V/ZFxmCpwb/hWPxpNaks+zMyH2cfhkCU4tmEi/UpbhnWT16xcogxqxPm6LpE
rY1ENu2qy3ZUFf5CzXUvjB1deN0zti+Se3MAXeQ0fY1oEXvWrGOp4IFu51foqa9A00uChsQ2wFp5
URTbuHeFMsByAxSv+GUWz27bGruBbqHj37rba9aBw83NhGESyX72UmVWD4fZwNAxbrOaSZtSzSwt
Av9gu2aF5bpLyBJjTc5K2shUo8qsg/tT8ikrBEtwVTqfi5KRg20PZl+xfQBebpA4zV1nRFIiZnCd
753WB8FJoHI++5TnfiuqPR9o/0qPiMJOfO9z2R4PbG0DD7X41Kw9U0ogrbvg3iyKegF5X42tkqxY
k/AJalwmJ26MyLPhGoZOwXrZBso4G7rScGXwHj4nWOcDofZUqMIh9aw38mZhxqUCNqTGaQr6edwc
sI7XIIS4hDNKqn2b1sA4unWJ4SKy8E+voavHmMbMzp+DrjSB/QE7U6aYMfi6w4Pv3IPt0QXkqnHn
nWKD0fUvhCB6m0GdpC6K0aHUyzLVWEbs8hIS4HTHx4NsfPCCiXSvidC7o0c8SGhFbTnRptkn4wv7
wx+V4ismkKVSiw+EQ5qUl3THvu6FePZBcyUG4d1ihM435I43O6yzrov15UZZdVdmegeNrnJr3URB
BiyqY1VQfTzw4ZJ94zdlJstJore0ZQMUomg9bo16iVpV4lSh7Omq62cffZDpc9xZW+V2eOD9AmTl
l4tlXOaj954qk55+mwxw131EekmtBz3px8x1GpVwMsXu//CEjt/AJVgTT22YYfpB7hpKW722TGD+
VGj5TTuVCj1MHI0wMo1BRPZxMEqfw9/xvUsP5qHhO63AtCdhC0eIcdcqxAJBo9+V1lvvR9u3qHm+
TCLmAKVpxVvcbTcKuJKFgYf+vmIRmM1mOIcwGqr/6zshg035ae6sh3OuaGNrsfoUtrSO6XfpRVaw
+GRCRIy+uLex8cGoZQ9Tg3oCCV3S2I/oAeuIKQSjCPphTVARgKLrGrNYERydBrZ0k0Cuw5Pc37Vu
7udbsWgjRj6mCqwp5hMVxmYQ3PK47SHCWCGgIDfoTQorPduOz8bCa49kQu7Qyjd22Ijzl85wC3Ml
B8MUFFNa9V7Bq+DgUSuEmciviWqI69hWcwTa4FwShTkZvkleiiikrfMDueyFVhKw3227VGUQW0aa
7WNSf7lXVzDvWzaOO3qCdtXvQjT1mkRZikFH4eHwgbvhBuv2Ufhim8jZIesJroTaHYjJTChWIzzs
tPg1vyYp8uiCUdRXWbvze8OZOMbNnB/3Dp/McjspchCGwirXGWk86anOt+2cRMD/yprViZ53h9X2
Wmw3U857RwQ4SilEMuPi9foiTaKRPjQYYOKLjsiCruvHdrcrQc93Of+UO8OziL2jSFltC0mFncr0
07U1uJn3V63bcqglGbYG5EGeYo1yOMJkJArN4iCIpbPlYC618bnF8XtEkqQsVPqGodEuWXsX8Eo7
9V3aQyXWNDefhHLwSZM8xz8xUkpRblV1uRUklxhOJnKYWDHcX3r7x5dCEaI1rUkakjrhc1syUJ0t
EbiacHywtOY0gqyl/lob9aHLPWr20kEDg2g6KDNkxLvDIfPA2k0qZS7hFvgcY1a9ZsvVT0ZbOvN4
b7R47lJhFzak/w4poZMBW+osetWNBjQ3kTMlrBEYcqpjr6apJdUoSRYKZdAclky5wrmntO7mj+6O
JH8LXWYumBiE8JQY9lBhRO7bAtgQ9fVv8kCEikim3KB/YHK2A5wSw+2aRoUR9qSVDKBDvMoTpXDY
NO5q//Fn1/lRtpMlzGl4gbeGmW3y5JcZw0skvcuiOfw71XdqFu6cIWqjEE4HjX+ID0gqL7MRPFHM
sI7TIj4zWxZeVrfsEAbaiUAgJTf2KeVDcL54LR4vXmpVHHO+SigZpJjZULHtYk0c6u6ixibnj2LV
rVHKwSyR2UvSuiYGr/Fc4wnmubucdjVp5+aYkHb+/XP8/EkwRpKBOf5y8TFB0wspeqXC
`protect end_protected
