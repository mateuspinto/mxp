`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ifwsmkJP+qTcsqITCNKEHEKfUx3jUu6PaJQoquSxu3BmRgA3DhFJvtcWd6Wy47QHqjWWF3dLksgZ
l/GCRDCQTOEOXan8Am6uwT48JEk5bO7yQxMg++mjtcZQCnwWXama6rfYZvYzamnBr9RFVUg59qY2
CQkaxqJaNjod5Oakewbkut+zDmc4ohjpGZKSPHXtoEsaKbpVtn1hrT+OFzpfmiOq+/Zc4IMwj/bg
JXIOvhjXEtr7u4VUGeVMyxKfHasgAsOvScARMNX092/OgznfewFNnzSpCDRuEol7T7e5JZ/xmmxQ
vZ80iCJWDOHyHM5g+UmZ+YBsXR0/tsnGTc0zSQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="/5n+IkzdeZOjyX3Hmoy6Yg8rUQqn5k3vM6SxilqfrZ4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2896)
`protect data_block
1B1HSy4VeDloSTTiFjijLzikChcmFgu+c5FbLaI6BwQdgRAHvTutDfau1yIAgqi7oblaDcsVrkOE
J+XNwOq+SARNqBNUF61GM5cRN7Vqr54hD6ZLJNYma5l+oOxgh2jXZblhMk6wZ4PQmnyMIDKKxyXh
ELoMjtYtj+8gaHcNz5gkGNx1+cbY1j52GNYqCYHsRBJAZpeuqHrjNk9b5dgoCrryqVTsEpWxgOdR
R7sf+2lft+Keh3cy48HdESDCfTzFM05gmd5SXWXkWAtZkZa0w+F86vNmnAhVD9v7d7euWXerGQTK
FxmNQohjSrl3AXr23wf5g1EDgfN51gAmrcVNYL1IIWCd0hyK5LTiIc9alKFAoWo4+mWZPdko8+em
M9BC07g5K1Es5Unun1GvEFOJUu76emzw8okPeTskiewUqSq8Oj77KZFOimTob+qgPDeRqtsxF2J1
luq0hSfZ46Az61ULsr8yWdrf2yAoniBh1cSzfI6KM+UeCd/oX23XRuPJ59JuMN7pn5C89H3oKS3s
m9lHx/QbbynmX1pWb2Hx7lpSkBgn52kn1f8nQ4XBPDWX6xsOtB6ptgeRwVmATRcsiFSxVlGAGmW+
pL3BlFj7enycEfWbncswVXsdnaCtkk4ELi02HiC7bqiW5yGt0uVD4rSbUrV5KRUyfz/F705PVLzt
3S6b2oykV8hTiguYrZg/MuG5htLvP7+alPrEId9Z2JUxTfS72BZuoKRIdqj74rjbB9F4hbVOkhzd
89yQJHVBefG0CeyyhTohzpTskG5eFytyDgEBJvp7+S9+WGPDyRACmykDTN/mNAgRoQhuNQiFAMeU
f5VUt2Wv6cyauDIUivuaDdwgF5nNH9iWM58La1f3Oq+WmgJuiIzOaNZyudbJCxgI0mQ69JO5BnTx
frxXHJPF11OAJdJgLjubIkd3lNvAzdPo/vcifGD3CUN3Zxl1N19VW34dEnKd1j+GnXoWpQ2mRhtG
5dzITxX9uONgddPDV33L8XLy9zvgZFhdTOvaJDeaCl1cguHAAtGptlBsjvNNWr5Mx81+X3PpQqdd
o3AoDRtHBmN/CXe36RjyB91Q2qE8fbcqpUwgzF9ETVBFX6sOQRkMA9C3pEVLB/pmlH+0oimn4aDB
Io+TGdTLK5EYcskGcSYkYnxTluZvgsA2/V1WG5sONitjSeRAFAZib1Iv4+VoxwaW3S8rsoT8BLSK
spb+jfxSGaUP+fN/iNCNpZQIdO7M0K9TqUmek458RRi/n25yf2OKrPq5wIV7kJ+daWOGRt/81GGj
A24tMo6SuH7/F4KjUbds3F5euI4oX8ktxKcV2gHsQAl2ivcn/m2Z6gqIbu/vyxWh1hfFThqsoZB5
FdlnXyCpMW100E82JHYWAVh/a6oTbfcOPU3R0ujucoyJYY/8Rsc2B9D7qU6sBMqF0s3nC43G45u2
Yx34kqhWEqiWpzH1+hrFM4LqBxrtvuD1ODAMCOVX/0BSpbTNgVI07/0CWM1ky2SlFO8pSqBc0KWc
18uQ6jM37SG1ks1JY+7dYm1dMFFWU/Dj2deBDPXpOHy5txEvqQwCfQWUFf6NVDrFp4RTd4CeYtjq
vNHQFhMmckFfqBM4rkHcgSjJjwQ2G5uqvdOMUPDBfNQ3YalUuQgFbOa1vysUJTIywakw0GmN0WhP
E/MdSFRLjB2Y16UGRUemjrv0tpXq+LBHILyRk4x7J/07SvwjAPV9H7EPOV3vxBBBg5bcVmuqwju7
tzT46NHCiuMb/pJqsgl6KTqr+BOXgcx7GgoSQHwGz8xINYTBgPIJez3q1pZ8YqXAoJVtHxcjgUi3
KDxjOO3wEJOw2RZ+z7y1ltztO+0Mm8AZB94nuNkzRMfS7V91aSFcMbmMOFzsKU8vJa5G2bzUnW4l
kbMAR00dOjTn8Z1fGe2lkwFvgyd1bLHLlwx1UPWcisyzsgXSu6G/d0BceyxmBvwma6MMhbLJt71u
1JTh0homvXcMW54qB6U+KrLEhXvUYCbLJaafUQwc68+9lFdBUICotfe1xjiVLkziJ9aa4jVkp77R
G6HbuLOmoeE3vRXpi9NGY90NPsslwefGgz4xNb55oqbfEFDjz6TgP5ReUzJGnBKukcIpmVdLm6ji
Frv+XkbGkmkY+TnTQn3wfMT2EBoPNISfXrnq1bKUBMuxPmU1SKHD3qH/hkiNPnZqlzO0qE3DhD1Y
iIUPs9oFib9o6Ppb3EPq+y4xZ0DehiaL0bNYJyr1lw5A5Gp+LC/nhzCmeAT0w1blDt+sgEaI4qWD
w5gnF7OYJovI9zk5Df3AQxUKnLgoM707cXpHOmB+OjIMiFMzIoBeFK4llz3yAQQLtp/pgqZbEQcG
WfbRQyYQtEkEXflyWRtv+Abs9OKK6AEmH4lq3hfaKMFHq/+72zBq5GSdtUc/XKN0rBEzqyfY0Jdm
KPrR7XXi++qJaZ+7vMz5WGMHwvQnVtMAuE2sowlCjzuzfQaBvYqmw/3y5gc20JHDyqKOsTpgHtq8
Vt3+dHHq5a6fYhQvDNz1DfZfI7XuFgJiTMlnOfv7y0BRx54cCyo9sNEHflsKma3mMhmeztxhJKkF
yxiZFrFobLLkY8FGvqvF5Cp+dMsyRcb5bV7yzAaZ0mkie7yUwEFjbC14dO5EesRoYos86dhocqQA
85g2NLQ89Fkitc6oNSg1NZp2mQQPFZEuiG6nNhZShWlAyYyhsxP35MDDNP3zV3ls/Txts/7Nfrzc
njewiWAPJcOr99W3ucbRnZuAUZM+sdWld/MwV0bp2AajVISSOwi/3GMZrw5UuEOWl0f0R5vbQgKL
Zh2utNuLYflrJM88V8u8IvWK0jS13BRPCvtYZM7wOzwCMKg0tU3sDCVVAFIYyftodwcCrUk5m1I0
3THTc/wA6hwP67dadiZvM6OJz7v1gUuB7F5dE8gFoZrW0pCYtKMPRV0xhiSLVojmyRq46T0y6NJg
sf0w+xW/q9hbfIXbmBsrhYQDWU3dKx6kLBrVOLVfE7S34fv20+2LqR+WvlDG9N/xzS3XaJYFbjvG
K/4qYZnMzONfogaabA3Nd3hgOex6j5Czhi3QJhyWuY2KUpUcgANd4EL8yg8SS3lQpTXMkCtgJUIE
7eL2AFNZePCphKD5NNBzYmP1gXsuo3giDWzNgMWa0UH+MiL2EdIeRvKweDmyGhAi0sb9xSqHE6u4
8GHNDv+mWpePdcby8xmPSJH4VIBfRp3pSyBrYMnhegwTYcdZb3xIJoyaWHopxKrrNuwX2Nfe+ENh
1O50adwZToUGrDVrrQDeFiUVg6gAwt0xhS0V33jeU1c8se9zSZev01sEunyL/7jUiHjoF5A/6e6G
Ktm5I/jAuGRQU6yCRvKKmCg0vMj0VdMxBHLX4eVhfJrqzUiNeWf7QyQ1Pha/+4XoGWMQPEPlTFcN
yuStB//5+ljzadVKJ1/wiFgxohZteUKkshVVWGra25WA5rBZgLE5Ac5Q95cJOHKzCR5CoW0cgj0I
6VghTP7Tz9rBX0m4tfFHEccONBJe8+np0ISkQiFYZ7ZCZU1lRADmBabH/dZOtgm3+kg8fqBUvdug
6GI8vs8Fz+yB+pAhKb2A/RhzEBJVDdKxftRTaXQj8k3qeDtP3vt8Qk2StRuSPWN3kt/YcgkeB3RP
j/xUH7jxii/uqznarA74KUJw9mmv0RD4bnXJYXvVDX7kefiZZYMrTbMbacoWZHUy6Va3rPJLnBAX
RKRuohe9spU9tq5GbLP69gWs4qQnKDucacY/EFtBk+bptLHDd7ez3QUVA+Ua4opSDuGY6ZHCshNZ
n2Kd0yv0mjmZHpcz5kKcH73xus6GxilFfb9CBXurZaXC2snlsSou/ufJITHYlA==
`protect end_protected
