XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������\���l�������v��n��ɕ���H�Q�M�5��.6"�ɩI��ঝ���-�1��$�o�1&��O�j��ى�ic��nSr~H,pmғ��и�1�D#��I1�ڑцIȖ|Zb�x�||C��RJz��TAs<��t^a�� l=� $���T��Aw���T�w[n#1A�`FY��%�}�`������f%��5mF�vN;2 H�������+�U���r�]��Z�#�Ny���J�y�y} ��π���
k>�@�<@pkyd���XW�&./X��퀊o}&�BD>+�A:�=$]A�S�(�_�@�A�d,(_μ9˭5U�iE��8Qϼ�L|fB
�y�5��f�(Ӥ�(���i!+��|- V�'����)�2cc����$-�$���m�g)a)��?��ȼ�/9������_���vD����p'�Px���}�pɻ��Au�et��8t�� Ȇ�X����t�O@r���QLr/�S�gB:��6i�IƇ���ed�<�Ն��>��� 7-�������d�bh؀�|9���$k��>+�
N���H���_�J��%�L=��_`�=�ơ-�H�߬�6j���w�.]�'Y�4fI��2%�篍8�q^in��c��Z�������2�߼��#%]�U���ȕ�/���Zs�Ns��iޕb����9��ɹ �)L���-8�9�L0!�j?���j4���ҷ[e��_�Ї�8)<Up�&� ��=mm��5XlxVHYEB     400     1b0%��O��." @��r����ƥN�m`�~�0�3�c��7�v݇�Nm�z���ϵ؈�5����N?���~Q�a�/_g�ɔ�<FKV^R�S���)˯����St�����V3�+�-�_��xL4fSOy\4J�	$a�Kf��ӻg;�� �ĵ�k��쮐�1y����)��}.B@|M�aWu��3�5���3�З_\��٘�l�4�#�,?;������6���_� ����d�z��z�"����5}�z�)+�N��J;�Df_�ܸ��h�o�������\�΋0�������Hւ�����Աxx|�K"鐵���Gku7��g�H��ϳ�5W	���0[s?�� .�+��]e�<��eȒ����
��T{���:P���+�8���I�β.f�����K��E��]V�V�x�MC��+�XlxVHYEB     400     160l������`�>4�����
 %�EQ���g9��[H��k��%ѕbf.�x2���d��x��I5���:g�g��A��^�
;Y�0�����F����e�C�E�=ߛ�+��J��'j9Q�{����7�V�Gh:�O��=��`��Po4pe�k����#����Ů��_7�J�/�v4z��5u���X����w�l+\;�ܥ,r�ƣ�gwX��+�'o!��/���ֹ�Α��|������i5s��\7�T�
��(](āv��#���<5AH��-��}"�[��!�=�A�� yR���έ�l�{��z?�.�SP|]�]2�(nY�J�-�����L��ݬ�[XlxVHYEB     400     110h��\j�.>X$���P{�Zٽ @�g���E�!Z�f�y�o�u�Q�v��r��ωN�~��}��h��ŵ�4�E<�}ؿDutf�*�������9P�~���qN	���ܗ��cu���[�Ai��F��i<~o�����aG�K�E^R���B���7L�/8�fR�_�$L}�#����[4=Z̢oF���s����������1K��:�gd�
q´ʹ�$Q�x}k����a��8D甮*�H<�{0��x�N9�XlxVHYEB      42      50E�|�X�u��}x�L�e��t�B^�0���4�PH��ppE>ӏ�\BAIo�Ī��ws�C��5�EB��#�=U)�;9�W