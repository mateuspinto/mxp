XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}�\��_z�g�?�m��Q��b�H�j ��D+:g�_ܫZ����%64[�	I��R��t޽������5�uT���s ����e~d@0���:��6��9��>U�'A�&U]QƩ�L'�A{s$&��e���U�~t?���T����!0j#�4H�'$���XG�$�UP	�6#��T���Gl�b9�8����Em45�,��m��"��\;fc{�����
��|5\a.�6U�P����"~�\���5'���D��F"x_���Ԃ�����_x��x�1�i��~gJy�����skW�\�g�.�.D�=j�z���@���*�*Uh�mW��D�Aw�ꆈ�I�{|��z_��Ď5[ �<���?��jJ���DJF:��$D��7i��	G~e&{ $��kN��>�D��U !���p�; uВ�����ɡr�Ѡ����{D��WGRMe�A�fh�u�f0��/�*6M�kI2����Ϗ��V��U���x67o*E�>� �K�1��{��Gyc��W���8�6%�=�}֡a-�Y���Bc��t�N��<���3�(?F9Q~�i��_����=z�_�oc��1�.��D��08�ɧ��FM�"���4��s{^��ɷ��, �QX�֝�tr��
�2�Z/E�B�������Ɋav��֞�r�
�(O/M�f��D�o�ps���Dc���gv��*�P�؞SQ�����6i��M� ��jm�=NK̰k�^��1���4�|łXlxVHYEB     400     190��XYO�����86����2�js�}.�����M���ه����4N`u�����ht
[QNbg��9�\�/�L�T�'*�p/���i�Fݤ������׻�'V�_��DIg�-������=Bm�e�L��8��<W�bǼ{5����wg/��0�h�]�	�O-�E�N*ѐ��Mf��7��,�w��o�����s�u�R�����cɛ��p ��~߰�3IB��OE����kX��dfQ��nӏ���\K�����G��H#J�%���sN�с�*�%��[r�)4��Z-'�L���h^cT*�0�}r��p���&N��$l4�Fg�	�cL�r֬&��.�o��U7wi���!i͕(*��$%���a��G5.cwy�XlxVHYEB     400      b0f���WG?���~�tܵH��ࡽa��/�(�d�@sx�V`�ˌ�{�۝� 臥$�ҵj�}i�E8P%����X/�m�l~�V�Hj�k�9L�J�'g:`[�" �al"Da{R�-pK���?SG,�'ޟ����Z�Yn����bC���M�@�'�fy_x�Nk&qQiXlxVHYEB     400      f0'
��6�Zl��C��o�o҆zJO�҇�O�:��:V ��k�:<����\ɸ��)D���1�b����f�Y�A?"A�����ه�Y=��4�i�޽��த��vẕ�w�Bq�d�����z1�3�Q3�#D��Ŏ�r�0�B����]JθX�>�ۋ8��!i��?�H�fc�Ϝ�Vx�|��z�\�/�U�d���F&�s�뷎�Ù�c�1;�HIM��M�`%�Nr>�XlxVHYEB     400     150��g�@ȴ�-�����5(�%)��Z��a�ƣ4�����́��"��`Hl��o��>�g��7W����5G�OkH����P��[U�&{bH����k�W��qP�n���)O ��f����}@��[l�#���/a7��3�E�@�ړam���x����h�+�SI�9�����N���
j�l'W�.��8���!�]I
e��lf���߿�Q����8�=��N�N��5w@qb�H�P���P5�ŕI�����c}���1������vDQ�	ocf�kޘi�2_��Q��mj�f+��]z�+?ʞ<h$8�h}��w� ��6*�XlxVHYEB     400     160�{���RMJ��B���͝��)�x�����hB�d͚nn(`��2q1��
����&���%�t����%�ie�6��t�Zj���t=Ab`h�o�Bk���4��S�0�{{E����~9ȉ�_�X���Ci8&	ߵ[�a�W�29���ɨ�;#:C�Ʋ��s�����z�`5��M�� s��?��x�@�>>��gZWVlP�u��FnR:6������U���)"�:V]�2�b�8���B�4ҥ��5>�����%�{5y-�ʘ��7�L��P ��!Z��_=',W��U*�!�d{�{�:4��`ДU��F-�����.��kZE x��f2�ȡ-� ����kXlxVHYEB     400     120�*�(�?���+��FWN���/�[I\�tN�n��=��6� ���.���ǂa������C|�o�����	zQ���?����:�{��+C�{�m(�|Q�BXaߓ��R�,�Hz���:]ܩqVa��A��@��@8
���)5r�9R�������;>�c���8��S=D��O�SGc:�U!�B��1�8��I�ve�V?5���*�MYMg8o���Y�t;��R���� O ��]��|�S1�ut%{�7��L��?�(�@%��A8j����b�1������3XlxVHYEB     400     110�����m��eS�NP���d���	�t�].�&���mU�+<��0-�]��0�l��u�l��>���j&wq� �?�1��c�nxo�~���������)��C��A,�ɭx��v���F'By�q"���8R���Q����������X5��E���baq��s��ksu����NX�t<#&����&�m���b�MS-W�����86)@pF����710��W�O�'bp"~:�̐2]�p���n�}%]�p�)��-� �3XlxVHYEB     400     110��ߔ�ok_��� �*JHr_��cj����s�1��ު��X�2�Wp �gy)>>z=c�EG�ʛ�*D����@=��W�.���0\B�56|g1���b�nfy�@qW�!��y�S�N"S���@�U�U�>:5y(���O���2Je���W��@G��I��Or�nWv&�����WJ� �s��[3��8s�0*%d�0�ɫ�J�"w3��������~�,R8�_
���� ����׫>ۿ.�Q���-/��
^�X=����Ə������XlxVHYEB     400     130xa�%x7l�fHǌu�.Hn�&�Ű�tu�{��S��,wB�s�dj��˗��oI���j�>��l�f�*����ǜ�������w�z�~��$��r`� oմZ����nW���?�~���J;�]�'�����23C���ްbu%���g��>�VU��/���@���ٗ�+(7ÔI"w��%l˚Gc�q�>S�!9X(L֌3I2 ~��B�B���ߚ6�_��2B&Lr�N�;�Z�ٓ8��Qh�(�����P�/�Q.��9ղ��i���m1��)��^�r�U��L�#�XlxVHYEB     400     140��h�u9$��4z�,����drA��lN�Y}�S�?�V�y�!�$%�{(���[ѩ�#6Kp�J�|8��h6#YN��Ӽũa��|��y�M����J�º��_>�� L��8U�_��~`H5x���\ʲ��4�M
�;��]
̰l�M�����.����R0�Zힸ����D�sΡKn\��c�»��@fx�)�u[�K����Z��K�Ö�Ȼ}�~A���S�T��n���쨭���7s�boW<��L�EȪg�w�]K������J����I&	�T�� �X�q�!���~B�oݥBJvY��
�Ȓt�$�IvXlxVHYEB     400     100\�$�L�ӂ�},+�}�͙l�5c,I����?faG� �9!���ۊ>.����8}L���{.�k	����a-����Q�L��"7�V��8�2���~�g�㚲��BU�\?w��SN(��}�SɆCa�(D����#H��~��������ZL���t��g��zC��]��,���M�`?�gmq�o ;cLR9����>�;vx>� �%�����A,�8���2�*�#� �cp������ψPO�XlxVHYEB     37b     140�������|<���MO?�9&ǈ�� r���f�Y��2��	~��_FJ��T1�".����z��J'�DJ����>l�N$�WF��y32?q�<���7Eȫ�(��+��� n-�N�v	�	��D=����Ԓ�1�#
f�r����~H�C;(�!��˞$x%�(ĕ}=b�1kĈZq�D�O�k�q���_��-�W��M�0.���%>S��q���Ȳ-�{E}����BRQ��w����aAe�&�xR�ǱM�=�	���!N>*'2�g/g̢Eֳ�f�t�lz��		4ԆM�
�LIH6O�`