`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
oZBjLoZvoZWEnnzRtIAHbhVCTxma2UW77EoY98FmYzJV5ZY5Xm9x1JFIeUmbRIVyKnWO/Ek4ZyAd
NmdTxjRWRL1/2XTF/1pPRG5gMrJuI/W1EWyOuq8yrmAOobT0FLD+QEfZm+juf0gPtbIWfqXnDttj
ClPU+IXby3jLu6UYw1Y29mmOZZM5RjdQQmA6LU4HwIngxHqEEqulj47tCCJcPZsqwCtgIehBs6KS
ARDXxzACSFByWFcEmh5pfHOCT/5UOrtdhtdrwyubySH8MsH3E0fHuEyh7pIwFPEavmNzf9sNn8N5
zdTHNBzsD36RsnD8Jy63ap5ZRCVld7bmnKomkA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="QLWAjgDNz/gCvXtv+t63BnHPjXRA6aIjiUnWkLmTtOA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
02PhJ8iaoXJ16aq2jtHh9l5AphbAuQ0w15ipXXizlCLd4BMV4yYy92hEM2jDdMeP76zdBu9PPHGQ
lK7osxXyFoGVNDvIfcvLq+mxlVbn1l/Zo3j3dFGC/C8a0gTeidHxKvHvY1+8KlwTcRypHlCaJ2CP
E2CAh1OuObfHJ22O/Qs0vYlrWPQmT5uUVkpzGyyKuqILqPn//z0eZb+HpMnBF/hUYVDdXpnQy9rG
gxrTLaCY2SgyalhTUvB2xXMoqyO73QqZzFevXmWL2tHi9q1XKIOhLLqdj1+UihFFmlgvlGWNW7jt
Wy9ExTq086fSZbuz0oYhu/EaF44elRvvZdzWIxEQ0GMcOuhlpZBikL5ECt1o/csn7zzZPxuBt0gm
0fh6iu5ubBVdHPODC+/6LAt81bqPHhL5p2K7IBGGmtMetab9ZN6rakKaGOHn1LBJkP2X/V9bW5DI
qlngGY/eKc0lfSoZXWJhBcJOs160kiEPG+e8z6DoI4Ew1TF5RIKp1MWju1cqIXZK743plfKEXOaA
jpjWwBpYQB1ZFDdixHoD4HktqSWGH3/XclvpKBxXmYUkd3YZSzNOFAFbBL7zE64K9IOXi2D9cszF
/v66VcSrLJD4zEvpKIKOnMRwMQUUE/qIYIQcS1U0aRH9rS9TINhpD0foC7YRhzmJh5fUCMNRW2TM
0XXGTEnVg4MhHadG9LIs4+qaQYFkyyXzcmuDRMtkMfLCc5nCydge0gEZdRuV0Lj9sK0B2xFyoRyy
ogfEpm/SrrK6TVNt0s9T4jaDZ3YXe5s1YHfOgiFLkR2yvyWjm5ZMUL/V1TULG1dj92ZXZ+GQhewQ
muSF3UPBp3aNIS/vLLhVNfD7dJoYqM1bCyUPJJbx7fXt25xLOy42BaIx7OhnZ2kIu27AQBD0muaa
5Lt6cVZ4jKYj90Z6fm4u9tyY3cIZ4uIG+IlxQt+HVQta16BPDjW0wKhiVS9hdiiOvCibE2wI0OtS
w1E6SCnRxd1UrhncywSaRAS94TAeAYWGjlkUYIZR9s5vkPG8STqKcvp1KxsSVSw5McTZE/wqBfny
JJf/6KrWQ9j4URp/zMJ42ZkMWszYVBxZPt5pK00WZw8PKH/mOfvsja7e49GcFzoB0eOw6r8Mp7kw
vHWrsmwptmS+pEd8oROmUFl99HCpjMXxjVOl257sXMMDFd6CXiS1rCfqZcJjOxbxzusv0rXvuW5B
McfFkuiHyBcgeq7TviaOcdQx6oSr4YdbJtQptHTVkA0bMbknBBXHvveT6f9ZLGLWqGq8Bn3/KKTZ
NYRFlbhTdPCKWEJisQfjyJtBTmemoJK4U0WIiTteD9F6ObegZEzGxACXC3ZxedGBtWyKmQfwQgMH
nXi4k9DlQTpoi0eAo70+0XP/bi0tnLb89VBCdH5UGE1qpzT/pqkoPhrS7Gl8qtySBI32NAecpVUX
YRj5b3L1gpYYDlnl4Vl/GzVKLq6NrAfveyY0ZvSGB7FKwIdFhg==
`protect end_protected
