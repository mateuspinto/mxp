XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��5S�O(�F�|A�}�ē�O�ɝ�\<h���t�#~�Rk@����s�g��<�H�n�n�@N����OvXw�vMߤKQD08K������i�kԀ�8���R2r��|���Ǯi�Y�i->9�h�U7dp��A�RC5��cF��иt�^��S-i�� �����lc���h�%m�Z6"I�T1&�<���:���l^�ˠ�^��;�,�s�j?��W��$N��	w�*Rm�����MI�-G<�m42w�:ޅfYWԻ�"JVR�̀aE�F��}����n�<����]I�?Mf#2d�C`CQ��Dw�U+U�-�^�;+���xJ�"���.59�qc4����}5%�a��-q����X('���_�ak���;a�Ov(ψ4%wk9�+}Z���e�9@D��ʦ(}�6Ȳ�=�o坮X�xt/5j�����}��|�E
�qMEa�N< ����������m��JE^dwi���N�9h�?�~��%_���sАK�NZ�y��4���v��!ӭ�^KPEg�rB	�nɄul,�2a�;�B��e�RV�°���4^.[�{�>>�f����w���VB3C�G�g1�&9$�4� ����^a�v���������]�p7�O�9E���L�����wQ �$׈qZ
l����?�R1��](w&Y����E^k�7h�����QE������:��P�ME��}dm�?�;G`�I�/&Ǖ���S����@��_����`��[;XlxVHYEB     400     180��0�BY݅�
s��o�{S
��qط��;o��x7�g#O�s$����3F�&a0GLYT1HJۊ#�8~[� haz@���Ԑ�������{��b����	� �M�������Jv���wײ��8��Ўv�9Ep���p<p����X/ls$±��?rhY�tU�c�T�Q����1�7R��$��:�1��L�����os�*��5�|�g�3���H�a-�6�(�L�Y�)�D��E�I� 0��!�p��׺^|by�������mp�4�����]Gٲ<���Nowq�^�W2���m����u�8�hkO��ZH��4h�Ϣ��VV��Ar$8T�i� i,'{1�ܪ�LY���C�1�rXYÕXlxVHYEB     400     160�k�K?[]��F�����@śtyu�}�U��YDt]��;��w�;	V� D�t���������B���ϐ��zt�w��&\Q(���zf9�e:R���G,N�\��P4T*�A�92(kU%�<�4"�eLDҀ������i�#X&|���Q�=�v3)E4jB/-�y����{ݍDkz�L�I�(,I����[�Lg4�D7�WrxH�M���$���w^�혌U�W5{����c���'Ş)z����}��V�b�qV�l�p82�ӊ���r�,�O����$�}?��������C��������$θ*+̫�)-עinw��iϠOP(��
A�e�+��9XlxVHYEB     400      a0��t�*'��,�J���Q>�9NKC�n�I3�<E�`��'ňĄ��3*^ ,���øC	K���^�HH0�,H6������� d2eU݀��dJ�@���i����+�8r��^n{�|�6'� ��^uS;dr�T�r
��㠣k�\$r�XlxVHYEB     400     120�J��C#[�d�M?%p'�"~���Ù�kAb���x[�@ ��\e�$��|8���~�D��@������ZRY&�:��N���%��;4Zg�[D���C_���Ǧ��XM����PW�o7��Ria����*BR����-|� �Zd\�3�XT��Ij��s��Z	�|�k�ـ������dK3mhɠ� �>5'�2��p*����a)��?.�k�6 i@��j@IX����A�PB�g�ƪߴ��;A���t���������*��d$��g��!�>��XlxVHYEB     400     110:�xG��&�˸�Q҆r�ϲ)Җi���� ��w0�q�����+�=O��qLB��*��Iw��/l�'��2��M{��H[/!X��H�yY=L����H�� 9j�%��8�DP��}s_V"E#l�gu7���	2���ʼ)`3&�9�4q��𗕁.1�?��!	��ٌ��s�A� R��{[��)�%���T��=��
�!7��^�}�M^�!g9Q���irhΓ��t>5���OO�qK�g��"B|�ݾ�z=Qݴ�����5��XlxVHYEB     400     130�X3%y���@��i�ߗ�Y6��W�>!^ ��[�����cY;>̪��j0�3@�	��Ob��Q�]6���`�c��N7Dl&�7�52�ґ���!�@��l��/��"����wS��{�;�$׍�.���&��1�IW�(���m��
�]u#���_'��s2ԣjv����
01)����������`�[M�˖=xh�.�"޲�ٖnM3ܤ|{{���5ҿ�)���C0����L�9�I4v����kǻ+�t������L�8�['C���6(	�p�Π���,���ɸ��XlxVHYEB     400     130��?�f&;%���Vr�~O9���8y�f��ٍ�6kK-4)NF�E�!�g��)�j!�p����?k���f�B��sX�?�9hG��y��(��mO�nAlE�@��Y���^0�/���� ��a����K�.m%ԃ&��	���c��?x`�nڎ�۸f�ݒ00R9������~�/����A���bM�Ե�hK`7�����Ygl��,"�0y>�!��(���O�m�Uu��'�^;[6�h�8X�0�P3_����5�d�SR6�-=�[����JrGd��"d�����l0�XlxVHYEB     400     1206��_��� ��)�Cfq�4�E���_S�����Da���^2���̂v�)ɐ0.��Ա�"qD��&~l��?�l:�C^���
��q7`��ˮ��K՞�>Y裍�����l����42ԡ��1M�ފZy;-i�Ć�I�<g��ѮRYL��ߍ�q<x��K�������v%�)2�V<�����8��u� A�����Aai����M�yM��.^��������!`���LJJyS�<L��<D,��dN��V.�R�$[�!*P����XlxVHYEB     3a6     180�*��ua!T�$��	�rЩ̎5��ȩu.P�������0cQ�-O�e�3���2�0����C9c	�2���K���ϙ�jQ�ԣ��;���3��uv=r�"��ɷ5���K���6�\١Z
ٰi�+�>��+��3�[y�dm�,h�@�wb*(M��F��"���–��O�(�1Q��X���B�����:��HI��p�+Э�k��(���ʡ�@�a�$u�.-��5�"�Г�Xh�Ѕ�`��׃��� k��r�0ݸT��a�1��蕱�Q{�&����<Bw�-��Q�������e�h]FCϝ�� �v���H�y$c�vW�/�9���"�l{�D[s�P�����ʯ��