`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
ivzMfffugnj/1MRi7KGgZhgHYrTb/y5osuuxyj4YAEcHwLtOWj1c78O+p5xK3La98a+ayURlyFQh
z1FmAWryctWybhkfg51zp4+rmlvW9amR56kXl3P1WAtz+EFt83C8UcqIYCEWyJEcBl/yI4inNYAS
eqWAI2QvKi7VUgh62exjkuPU5zD3kzQ0FX0NjDBfJmo/Y98jXl34JyktUA2K58ijg0xRadD9g0bs
COW8TxnHFygmKG991H31glmsZ9HKso8TzSPcW2W14PQAvaZ2EohYpdzxsvQ9DbSqjXh7+/euFdkY
vSoY+ER6SRRH3OcWupnRvAciauQ+eDqISjInb2PKVAMntaJf0gRXqvXgcZg2ADp04ewBQHprBZXS
UnE5/OFTZI0KhWxrBfiDjNPY6Y/NLI/TX0bJ59LvtczKQxT2CVR05BwHFyG7JQjSBLa3k1F9O9BF
utzC20peh54C7PQrIpgGhyOZBVqvZDFx0C10e35pH6Fn+DMfKQN8SUnQyDeoSfZFbg7xM9thZYSp
TVrMDRhTb54vD4hIdorXW+5RH31bQ5KvlU1e8qDdwQ2lKcPXhOBHHEBoBEjrNF9KzTw/gijCaZbb
A48q5Dkt4K5jdTKIGwXq35/T0nj+jYNHZQ0FfR/Hp3Ek6n+8/Nurdakmj2S3f0WZKYFzs276Jhc7
zv+phnF7ukWialuAOVltNHAKSyKzDdGvKPwyko7cymFgmwORsIadHuJOTpi7IFdMpGvrI6OatVoL
E+NiCKVMO5zxrvukuStVj7hRJBzWQev5R1lhq5LdD8VddES7h8abKykCnxIUV6HQs1Idw2Am4j+V
j+J+LkOo3GdaGMex90EnPfrPif064azEb1XyrxNDQoFJ+tn1LFWXw+3PC9MMDNVv3KU6yrhc65Gk
kYqQNHK4XUR2lYUtFTr8YZJoBzsNavXQHyuYZe0/dOh3GLzeCTVRQCP5GjZLAR1sTOHxGndvFrF5
Rh4QcSOLXoSjIEzVabHeteplPuFB6PYJiMlfaasL4Tq6f2iR5eL9I/K00emj3jlpiKqK0HmPmez0
mj89Vu1ckMY/iRs7xQ7zGAoSKMKNuQHVhb06W8puje/jfYiYVEXQUUzRl/lTF9EzHx3/jWlMkCnK
d2SXG1xQAQAXIWyuczNdRN93iMibRDvCxGJ5ygsGzS5IRhDCHoj/73McudbIlJ5oKM7XzNUacvlT
nq9rUHEQBCIyFjmbwUhsEAKT9cNhOjFqmH4jgudJZD1biwsKE20lhc8pKR/ae6+XlZE0RI/2qtki
E0bWtYm9nAWOTJXXvg4OXmt6eA0/rsnkY545e1oLoYOUdn5K3nYsR/bwpIp+WdVxUSZpYCI1Q/Nw
WJDYWpZVApe+JUGpqR4xLnMtWa2lGQ7K6wljbhm9J72E8ywXOiQ/276pVlZ4XuOI6NporYWdnNaY
2jquNfkiVv5kqjuL3awz0+yNCXJNZ/O2jIklA0U6gO1+/RnSBYxdculwHBm3tFTz2Vjp8QWVpDT7
xXptCTGDASMAIzR3sAq6hBoWIuev1hHcRkT0E5Hm+fGB2V+zuTX0idnhY6VHOW0pSeuDgFD+67lV
05SLXdoWQJXNGxj9LIW0TFYarPdeUPjrhVP9LrmC/XUxTXNAnYZZOD4/PG2aEgHcXy092SsS6IYm
GuFXQydz/ijEhKbJb8WIcUbDtyIsYKTY+rWxUUvx/94XNk8/P0VXkPnTfioZc0ud4L6xBAmxa8Co
2GiqGkCHxhHZS/ItPl5YhcRyiUNm011q3ZC1tPtO9y8GHeUOsxKObtBs1etN3PPjDCZFwL40QbrN
Jr/KSQ/2csr6cmYxZlacQHF+KeSQ3hl0afdd0X02YStn1kofvCliM/kl3D4nuwgJ0dM4hHS6//AE
t3W+nUFWcr4oHr6Cs8fOWaEw3najjVcShtw/cNtG6nqujV/d8rCt72MiZEPd8WP5pK29JUEJoajQ
AITpm7oOFXkwDKzEkqsP4RQdG6dSRn0+ltGpP6SybpwNbPKnI0jQFiihtcnJprgKnkuult1Vf02G
Z2c3J1mzsa0GcJyAOzZ/+1poAEffi1IzC/8e+3PP/JB+lGPVSNf+XfXsrb46
`protect end_protected
