`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
64nFa6JqMrquFxqO6Sa8EYUH+QucvSKWXrv1KIyNxEVJwxo5ZX6X6v+4UYbTzr828ZQP6EbbpR8/
QUebryGzm4/5AeUn21GG7DoASjma288jujuUKRqXmAIMVQ6AEuEdhXdvywRNjvTJclYlaWOhJeo/
NwmAVSj8sdG0hxf79M1KIdkMCjWL7g/0gBNNgXoLaqFUHeMYwlsB4W/Ggb+H7b7gm6PJNqygjOi5
Kl9ubJv2UMJEKl1v8ju8h0kpyxUxFKJo2yD3cAxE98a8XHObojnA/lHiUiuRYag4A5aGSuFZiYc3
GP7xwcH9SvhsfC+B/0OVSwRH0nAdCP2VPfSB0STml/hBD6WYG00WjZiEx2Cs7CS6ZwsZhixcVUcy
86LCp7LGc1C6aIR562FpSIDHxhApy4tthb+1K+42awhOyuHwG+yi38U+HtDgZYhILHBoEM14aYfl
4H4yqzqB9MCRXzQxbW9ZWMErr+fL8IRrqGMnPjuhuIQsN2z1DfARasTDw+JzIov4N/s3vVF3yrnI
Xw6Qzh/AGaAKARzikm+XRITO8PtWi7R/FBJURVsy3K2SuKc9lSoS97weIKR+c0HvEkC4ZdLB5Z5V
q0HNyuDyUUhL1gfdRMPJK+PdwT8sSpaqe09lTXsDeyTq0EduDBYO/xA8qwRmVOgq61VRqlNtx7fR
qM9I9OZHnkJEx9u9TWFPiGsD3W2OxjAbRSIsKEF4GOmUERitUp9vIXV9gB2ANM6Ka1aryXofzKaM
pHXyfaserocekswstLB0ZGJ0+FH6lsyLybK4KY1P0gORISUSQgnCPPGf3Vl5eTspeGwgp+L2c83d
kHVnkfhEQUhiNLvdNhztUhdFlwEHFeUuhsCKeVQYOUslOYjCF+HlvlVYpVMonpezqQ3p9q95Toxa
H0AhSf3CoGeC5IFaQzGCONvEVaBtIfhB2+FzVvxszeRVvHE/FFhoLYSSPTBa3oHZ3PgdB7ESPyGh
Ec8l6wqBwMfju9m0WaOdm3nsgo+KzmNa4NSMSaCflWFSqf7mgXm0UJT4xjIHsmIpKUiqIyrOQT4l
ub7mmsxxXWe0kA/JlonJCAYqlGGoX88JSowf2GCcj5EtF48yBFZAgXk4V1yWLTQnxLyNmVmyh/p+
/W23H4XcAkC3BKJ0Mj4Ez3/V55JRmhwN7ZiO9QnfSTP2iPdAa/8CY69U0vw/gNqF2zW5O9cjAhJm
1sRBuntVU9NP9pZmjFVPh9DoiyCHSk+v0Q7ko6cD+F1AkIkmaCBqmQbTyErp+x713wW3u3kW5/g3
B65FhOBTIr1ByLX/0wgj29yFbKmob9t9gg73xuKZjASahXxqRwMJGD50AuWYt69ltkZPGPpT8vq9
8avKGbo3GHsXic++50cgWQoGC9+gmZlydZYjb+2tjxmgqWaQMJULpYkf42L4fF9GCU97ku7MrRqi
QKBKbC9pnfFCXiGUy/u3JE57DJPrgTCeUwqyCMcWppHWoxVMWqik2dmmHldck/vA5Px8+egwzCyw
ERff6PddtcWswHCnu2QhwPeII63vazQW5XlLC7eqE8wxwBf3KEA7TJV2/DlNQ8pyjZOEpH06sqiT
OUaRHCaQa6OnUeh5OU7fPDHNYvGyVLbIkYZAXYENzxeXzq9RFzmf8HmsBGwxN9IEesYBvQPfA/cm
CqBY6dAdVWxZuIYZ+oJajaHukB83k3QsqUjZQmyZGWO9bUKQB5EYbmU6v0HGfwn3dbszSdcQ+5an
/UmozLjwHgLT77BEs9/aE0jWTM2+hMfjtKSuYHyNcyJWIEaFsiMtwaIqMzenRH+v2KDtG6WG0HNO
5k7PjYvAZEp/t6g1nBGRs5/fXw4o3IqLZdV+kXIh8IerrP1wPO1dvMRGak45u7SG+BTtFDUiDBrr
PkZ7vvpyMkvQOG6GIReLNn3hZu6uZONj2coN5SnMzgkR2kbV0WyAwYXCBjB3j/vcln26ve3SC5ZD
Hk5jGBrA0THUm/Jydvt/RWSyVg8/zLEp+E2pSvp0Bx51b3X4Hz/YMkFJl7V8o3X2xYwPsQV1H4Jd
1aINN0UAb1ArjowKSuq0nmDZJ8L4EoWczIDeR1ik3uU52KFflnZ8aT7KXvVHJxezHnyOw4MbCYeU
A6alwjSD+jlufz/9XDCX2k+j9cJY9p6hGqU/RTA03Oar29NVqsHOiM6S7dAM9wlMVsiuq7Jy/SIt
ChqwxpvbWUWIWGpQOsRAA4ZJR+fQ4S+cY/LP0gwxbdGpz2l38yPqDj4b/8NHV1DeMDPrAvhfX/n6
c3zvZ6jpsOKgwAIvfxNbZwhTIHEH53kwjgg2aa4xwsiemMxPR6bW1qnrpKk+Ms21+6OYcISgtj4n
Tvm04PN/I5i6CVYIatV0vEclo+Q30GS3xrL9tonJOtGm2bH3kkRjFwTPT6soJgUb0YtxQfxfyfLh
2keIWi9maq+Bm6VY//seonnLJQWbGvQElmpaw7LnlIdKlxb/y9vGT0vEvULMSTGkv6lKtOnjZjIV
Qa7c6ReLxyT40IvHZP/ixujINW67SKvmBs8R6t7alpAhtJM++r5wf5rhAacDkpsWIXbAY3rDaHqs
gbTIpP6ITPww0ZCK7RGssldUbtYB1r+YjJA9W0adTZPbpFu6UQ/mQPS5GeX1CLOTFaimYpN3oP40
rteOl0CXma9HURcH2OSRM9HdRTEtqasOMBuQEyOwtF2B0Ohk20f3C3gUMTzSWqKypWEV7O0ML7qT
D6d2pccmwKsta4LP4KWuqbwtyrSUBjSTpcfLGohIAkNN0XkrkQwhm7mMQRLhaAOOTxskGaIjDKN7
/SvoBZBlQGsl3qJuda2XvSJKGPTJPtdhbSEWJ75xTOD1NnM8iHfL8ahekfIGrckqNjiV02/KPapS
MKsHoU8IV9e/RZ6hCi8N06+Ujvs26XN5U7/N7fVnRIbWJ6lnc1zK2Vvf0jXNWkvKPicMthpRQJvm
lmXUsbFHWOCG/eVZEM9iSR08rRkgimh+XF6c0VuFVj8a5QEXV1fVp4Xpe5IbheDdYhtJFIVpEppB
1FOdCE0ICYw7iCe4sKAhRj1eSzaWrLZXLHbJYUhhR0mQ5mQxjZ8yxD4XstMlEA3aRGn5Yg5p2SZe
P6XuuB+J1Fd8NpyMeMc0VrxmRW3JHV57hfGEDWYj4PE8HIr9nDs1PLpuaErYgU3s0K7rAuaxR7A+
OwkOPatg2aq0saxiOTaQHj8T/FT2mT1sU8wAz0Il6S8ll9OEeSfh7iQHF5dM6VG2CcFg7HKCFYdN
jLAjQOlSTSykdEQRsntPCvi0w9MSO92Ht7INAh9m2PPwhwP+oUNPiDpS/2OWPDHLstZ48HjHv8wd
oIwEk50ky4KrAxNt6XfomSMYR2/SvByEPfGsjbTBK6dogVDut6l1LtPQ0NHiKw88jTxEAltZJBDf
hyeh7Z0BhO2bFyxnjJm3Umd0rMzFcCfF8Vy4cMnv8IaNI4nXSbL1JSC4fjgg+5yXYtFmupkw2V5w
F373PnGznF5t27BwkyhMVQmtkiXlFO1RZ25gPeYY/O+oM8jLkj1oc7gHehXlgQO1Y87ZqguyYXb+
3JK+gSrJIl69f74z1I02OFp6je8cVZcf1WmnkVEKDadAPL/AeM5OPqtBjpOz5a0iX0561VFQmAUo
FSmANDCS3xl5jBaidn2H9dwDp+b69ipjrUwbdojPsUFS4bTWM57VTChxYnZionfZX8wdls3LfqE0
2gk5lgxFOmNRmaC63HQ2Nq+VzEdRrL49RHTqO7yiOYQKanPn9YUCeJc+WVNVg6xVGMm6tc3+enO7
b1Yn8FGHAbsujThSVS+Eke98b6LgbCLKa1rt05i1K/9EUVA7LhRpCZmGU7vl0VfKwCv88MPmQFu7
nrS1CSMlBXU80pJz/ZgglekQYJ1Wh5gJRDmWeEP49RMH1pZrMYIUh6nbzq1roFSW4Jxu5fdN35VN
fLW2wKmfn94FvqdP8WzV7JnYQ0k1VNaS4s9Sv4kdIrEspflxTV8sWJNayZGhtf/bCla9qiJ7VEYg
Gx8UOl/aMuEdMkN46XqXom7DzDnh+nR6jSfPYBDB+YdgCMVdr+YGMxV+ZAPlfTwsenIkxENFPD0P
T0n75yK0qMD6dcBrLKlTrBaMppzqWDmXieNkNAlcMJtXkxBPiZEF+Hm1zO2oqOOnWaFXlHS2xsTZ
y38trd2UOPiiIKKTDyLxzNFRmqrm1l0XFZCyGeTpM69laZzY6dyW4PeQPBCXWiyeA5Q7PBeBokg/
mxp4V8MCo7b87coju/uluUCk4lZe62IJrWbyjFRc/FIUj9E1M6yMihdNfUjKz4IJXVLFuAII1x7n
TA7lUZ2q0LsMY50g4dtxIIxRyh6G0NXdCQvVIkLQPvOf/a4swQMSAUsyTHGnumIxyAu5fidhaWQa
ycr3qrSC/E0NmCgjwyLeLFol7zgs2sQrAg46a8hc9/k7jSj6dpxHVQTkynObCVjUQNTO6p+1uf1A
PdonQAlVIHGeVaFJuVR7EcGTqvmaBGJORbbKWye5Jhrrl+m894/uTvH3Weh94tPdggg5R9jfZWCM
U2ycp2yEbZVfGPTLiTKjXws0JhliDVx47cNTfYZU3KL4ZkJ3YkdWwDJhQLZNK+7VMK+MgMKw9XUr
xgYe18KmqhxuWzeoTPRrkJZWN2yfWaMzVZw4XZZj2+OEZRZPEqe4/LlC307sT7n9+fBzKm7GVb8v
xJjUYQopTYvRG5dx4KNHdhwzHvZk54a2snBJLenOtLk6PpRvnsk4a3CTzYxYpPuX6YFcgGluFeRB
imdF3vK/GtktZ4LNuufHs6DbXHe+okVNTChUDRdNEemFiiOjoPI2u3dMRCpJPhsJvf2RKZyWTdN4
VU+KKXLVWVeocFuFnIV6yo0auN4owgi8eogn0VFVNjWdIWWPv2zWqtoA2VSdAKS00lSI2EaKvhnJ
EH30i3yHGYaC5T3JSM/mNhWf7SJqs3cdIahjsI48HvMRzWzqd2fNtc35hXehwBAEZoyJwv4IRPIv
5vTuREv5QydrgoLknq0HltBWMnfm2y6EhKuIE48zxxpQwm7ua2fOUNdKwO3Co/1VyYvSNIWb78LX
AS1J0jvc52WEXOgBBRMmC0cU3LBxwS50dwqQEh5AwpKRoZcUZW9pKqB4fDM29NxUtubE8d8nW0pQ
iD3u2ZvMxtAOEL20g8ILqiLKCbAI3vj/Fd6Z4i8dkKiyvZ0Xq+FD5eaFicl59F8WxEhR2afwbdCr
/mo+Uk1lC48bpMTCI2VTb2ufD/6m7W8qav/w0toaHtdDC0R0yVePn56E+X0BBrXV9nYpM8joXtzJ
QhIC+/UnoPLbIPPRgaavUWwKmW7BDR9sYzEjTUyXJpD3ZzQiwYhrKE0hl6+IJlT5XKTV5BObOPwH
w4sSDNPdK2q6cSaetm/50VgFAC76qM5AjB/L7EyVyooZvJ6B9BpTFekTYgyI9WA0sE8IHyqzWYw0
rK1VPU7RHA6piRsxDR4b8R7exKgUXX2aVIVvOZIWu26q6IpIdSgnDJOiHaafoqFi8Y1E34US1DJR
3igaJTujDZomgB09n49IizyZVMvLR9ICESYPC/bu5J8HZJdjlWq/05vlnxihy0Fw/SREgGjFX2IG
bqEW4opoBx3S2ZFAUpNtsU6ZnQOBcrIJt5KVfc6fkZeLZ2w9lUiABjv6jp+py2c+kwjnd21fV8Pq
Ex+OGghHKHYMidrqypODaIpdiVcXBr2WS/U6A5n1bxEala3b2jYnmmO5Z1CVy0rV2GbBhB4Ze4sA
fqx4drRLFOZVFYil2VFs7dMPd/EjpBBd/zH0jCjo0VaNBa7z8puIsb/zJePFHaLHZ287Vf/439oa
n88X1uJ3NwZkXAY3hnp/dT8YA3+Dam9Ayqyr38FPHI0BNcRwS4Eo7iqC8cvLJ3d7PNG1jLkE9E7E
Hgn4gj61HLzIDwKXwG1UZsqOPNpQRb/1iZ+NCuy18O8kRipNKhBsK61WaeNSjj152ndy2aC25yIn
6ydoq0rcifP02mP+/08b0oTlWy/+3F0WJQWeaUUhEzwqSc7aqxb9klZ1+pOzx3AVj+JyfrfvJIPt
CLnZ/9bfcchaldArY/XLg0z5IVnUzRkNl4BKAaTAdn02UxgH7m0vXyHf5MmIEL9z8+s+WkQ6riXy
/cKY6+CRXCkH81rtQjbvYA/8Z5U1fU8f80JtKoL0BexBv8b51v6c2Ve5HW5EcfPwrarpbnTXpV/W
RDXGZzhko2l5j+lMzXzXGRT7mfml+fxsuH5fwnLkZLk7w6Yw0Q1rUzx3kYW3UwOTwev4/h1L+d43
50ETgh2WzvSKHxUI5SQ0XEx4xapYmr1Y8/KPBzJyL5sLroJuCXORrQNLDI/l0NMoyFHvGAWN11Wa
FVULuGwCPLPmOJqUSBHKb5zH3Ta1ZkZXQae7Es2Smj5zmVwp2LWLbSJn+BZYkmGicOGd5LW/iLjl
B37ce6m5wVGHWN8ieGohD7Rf3jLmxYmMNFBasnW0B8oGmUGKFLmz+4vVTCE0Z1U0+1w0aYwXKN76
/MHaqV1EQi1D+2hGrXWJczs5E0kbVlhaUXWliuYJv6a9gRLx4ygMWQLPPyFvOjbFNPOSZmld2J/E
ZuwXZ7LSapQWEmN3mdVk8e4+8+HzYhBC5m8qgkuQZjh6VSM80ys1EoOKsEnPVku2HaE61TUrBW2C
wOlbQWdN+ox1WKdxFXPG9pbjHOK2gFyFnZl0GQZ/Z2K24rJRGQ6+SUHiosYy/qmLAjyFtkwwwhps
J1LQECAtYHSqJcucF/ETI+ZDXRDDrT/NUJqorwmwJy9Z26NzdLNv5/BBMZr7x7PZeXjJoj3mRj66
7RvWidR+x0z5wOE+/t+Uk/Pzkv35dE54cW3fv3opvjMgtP9EMf1Gv87GNcrerc9F5eHHpwk1fC1a
iSSmPGBwC8VFgEYsn0bqUYQJXbBIEjbwFTLiat+FfGMEdraHkHNq4EfaJaSz9PhTeIP6r5vxNydB
cyYrdOUE722fo+GEWE8Jw1xkvqVsoPv1zdiCO7TAPi+xdxwgAtiFPa4muR2EJwUKmqSGT9wnLe5G
z87Wm3RIWiULqryCB0RS+KZfbuf+ftMCammHjVA1n/5zUpyk3SxzpbUyGXWbe8MILYKfedLm52QM
CQ990l8tPKDmcRPdduzYtHP3fXNsyx0VcfhzZcxB8mnxfVNGLPihRU1lt22++WT1TCQP0HqZYXFx
NDgzPRb21lXFeXZpQtkV9zLW5GP1He0nZpZKzvlO8xrZlPowC1IOMv56uXE/hv5amrGlN3RfDD9G
QMe5iVj4qUupxhficMPvRNDPtIU2y5htXliDbA2V/iKWho4uDZa5mZoBahwspXfHrdqqYOyH7IQy
0YkHClYvmigzLqsIJ6SWsEY2KnZ+crhK2TIwj7kv8mBSt6J4Bpyn/vQHBDIxOppzZTQqbrp48ndi
r8la9p3lZvnmE16uhwuVS/Y3ydDEi7D4eiPeHq+CeAdo2mtPwP8MdU9NTFLuslS5wuiX92a7ZhnL
SZtIBwBignuein69ckR39TJQOkCx8ekaF67MRUirX8WV5oHXMf5NYtrtN3UPx/g5Cr4ETDHEhAbe
Ei4raoRWTDo+rR8hX8c6fRUR+g40kQ7NtuFDze8+iSGkXz5KHmTVp7kgl9hnDq4C2tE9VGkZ+KCj
gJM/SC6Wm0+TtsNj7xXMgg9IUSdiWHmYPOxO38sVqXC2HGTMIM6Xbp/lQkro+beT6bLOxhCBZBzu
IinQw08dKlfCcV0OYL9wIaNcSbGIYVju9GPpKNKAImy1wfrhFJ/JGeHY40qRvjCTu2quRWphq+Rk
HTfIjh51X9oY0RmfwZa8LGqXDELZwldmkAle+0YG4cBXGblSBXZ4q9V/ZkiLxHtaDCg7u9Y8DfkB
Vr+JeH8GEBU08h50iswtoT8ekfbGyiuWOrXq8F5GQqtIZ1GzTlsdHEVB4lzsYg19FeJ9fogU9SPx
/mgtsu/u4G8VBKXYcIG+oneZrKtwa7ty2Ul6uhVUG6HwWuevr2dk73UbS8gZojWczoUqQcWbKF2J
NFqkPwcS0VKSBlqdff+11dI9Aoj2CZZUwBDPiMx7aeurBxfH1Di/IFPKv7WWXAw5KhO5w4QbNPbu
TGiUpSj+9+KDOiHVs1Ax4UeBl0ofWu2FGV/8qYnZXHaTpvKmxX2PHubvqNwSwgi0LpVLFN2581fg
54HvdITIMNrPJwfWCcOdET+L5Pvf+jkWAre8+8DgCw7vitPOB8QsTPaUQwfhWNbRqTuPo4pWGSAW
Zy7nyhsQPgVx4whOZl6xhNBzMzQ/NXqWunUurZlqyMAKMakWmq3CrGXmoX8cqOLBZ2XfL3rmwvch
1IGDO5D8hCvv93uJbx7fabZA5hCgHewfRdSfCdyucRFUX68SIWdPVEWVEYOl7wxAbFw6okOMJK4X
K3L/BpOndyI0NyJhtV0C/5U3SqTG21xesdSrXNQhG+9suVmmxcRn2dC9SBW002wSbkcThyHJGkjq
moOGAGXMlSuQYmXxi0nWOYXZp7ueR5XpOXwBIHxzTiSNb83Df63r1qp+2eFwFrUkcrPgFbQIZrpx
yMMm1aO6HRgD/5xrlRrw52BkgtZ+dvbDjaOuyCwBtydyG0pdA2i/tgXxkgzET90miDHjTQQiJgqb
N1XP9TY408X0nCT3AyBCN/gb1EFeFQrWmEQ6u9yr0UZze7+epFIBGto+8a5AhLh9rcDNHJ1OY1rk
lu1ZXrUp3g4ltYGmf3UKwVcll8u4wQL2QF5ouzMwKOwH6noiW4E30aUE7FY3PmqIK9C2NOHG9jP2
XleGgJN8PtAaANxjoo6X8DpUHXqkaXWwP3Ye1c1Tsujai7Dk2dkmfw+qp9tdS+U69V1g8SrwZFK8
EkxVwAk8YX/dZTqnz2V+qho3hZQKR5pFRKqUfYYFAXCq1+qDHAcDMnKU+nShTSAOMC0Zm2zMsTCM
eRg04ZirlRdovAa2sneBq02zp0zrz/VPcD1UklNh6wPwjx/X/mKZuOlAOrnTZLaGrLXVqnVnrhe8
n6F4pI2EvLKsN8r4DIORLNuIgO5nvNjsPrQMTM9qi6O/JeC4XMvsQuWM2WpBCeHiZ1DBiDK9UsrY
8/8oOWlXUIfGzRhntEo95azgA9pmxreLuk/BLMPc9LXl6xkoCyNmIoQzna9jAZjz1ZIGrBpoz/1R
n/qfoRXgBKWdWBsiHm+YOLLIcGhTVZVgC0ULqeJIW+7eSPpv530EewHgR5dYXV0JsdI/sXRStS1h
f+00l0OHVuxX6woqRJPrLbkR31wINQRZL1sOnaQVXOcCM+q4I0UqCZVSdEvki/l+x0eIAWKuM9jd
lAirjaj9Ehp3MeiZ8/dbcBSdJJQwh+LkZVeH9pZ0KYCaiF73Y8OkiRz9uaFHPelv5p8QFrn/Jo2F
4fiOGUVZw87smF/cvnBuah3YW92I6eXXWbaey1UvwqodR+AFb/QO8g+JpaUI0V8iam311kWYc4en
stTSJJrVoVKa2RahNbJrNQfqNKeLk9jIXi2XLxoBEOT+jNqhPtTDkuePO33Q1dirLu3/stnFLCqm
JTzgXwtiqcr+fKZdiF223rMuMUUPSjPeBUzanEWbnl3ndgDMcDOft0ey4rcUsV0fB+Gj5F+Ve3dI
Ke8iXBVLkQgE8GSG+0jXtrxdwmmSaL0Hz3C+sR4TF4O8DWV42Qp2GldlxBShl0vy6/+u/bDP2Rh0
f966qJR5iSfRT/Dmi2xfqKxRq1vbLbdlB9K7OaL+KSWVq4CPHdqf/uWyL4YZMeodR1DfGH3aCNgS
pz1frHH5ioKLNv7XX7x+vfYR3IBUNWCMyPZq2/C4Fl/W7rTzaLRUke0b4UMvORVVq6yEKLzOvHi6
jtOvLlUWe0tG1U1auaVxUIKNYsVFQr9wxzKk+mLYuksjomDIAruyH3vX/7PtnGtcowUOs21bNkLP
iPQRvoWqfp1CnixyLESLe45141ZVetQHoWh5oIA8Cvfay46JdOP40FwuUJe6GTjX2iVTbHsIyQo8
CBEa1NqRVRtr5KdoJ4JF9PI5LYOgFuYMb+SegnVdJH7ZIck8lOtz9ybgdDh+rlfEzSEsQVf24jJ0
Tc76eTC4jsVr1uABbCD7/5ONeebZ1jDWGxctFOqvrUeu64ThhueZ0TvoPi5cu8JiNhfQhhMgsVjV
ofCl01n2mOi21/PUh/vMnsh92AUYYk16R5v6o0khsXX3zUuJRARSDRmLmf8XrvNA+25Q9qg7Cjfs
s/PsPeQ0huOezrTD86bx2aS1gt92/hMoCKHldYEqb5LHzG1CwVUyPas99dGAwBbtYIfQW7B6TZyD
JUVno1wotzM6nRlN+UB8cdlM6oRTvuFzlr8AUA2blTIe9ivPR2WejYlitDu7IuT17M+Knz8RXNfk
eRU4zHcMD6D7EVc6qtFMzYzk7otnAKyGLAO1qRgpy5HxBB+CPeJwen93w8HJAR8iZDrahqDpLMHH
5FsOTNnaxkvdC6CGQPLEJKGxjB/0JPbSOLWneWerbr6n666swJYLDJltaN5RcdwtuWK6hcJ7rdww
CcK8rJ3EPMBrovLtsz+LB8qUhTritJeVRwrfcegT02jBLxKd3WI7quStLfHEPfaFVs5qhLJkxnFd
7xpu6I31epQtL41/BYjMbFIIWR4PQS+033N7uhViP8tR/twsZlzuz/dku6ELA1gnfV0et9eRmdnw
Kp6QGB99TORvTZwVl28GJGfuGIsaIr/YI2E4rsCIorikm1tvVeOifmMB6LLjgdRgwvTJR2/rK6Hd
D1LfXYe937Ezc0NsYHC6ez1Bko9R2NcMbto0mR/t2SzgeCdNmUbZE/EcEAcwJ03+7GwQgVWsTgBi
g0q62seS+rjVbNp9Kpi5Y2IYYi6W5RWrklOc1Vea0tceEG2Lh4KDC3p6RkAmEG8XPZho0ktv5aUu
eq58cOGDtsTubOicUFNppZD7FotYBpwduUt6qlcBLMASzPGBKG8klbYPn+M9H3NCjqhdIquy2A6I
GEnY+wfqDnhmIYGqKGXqWL2Z/QeuV/BOyqo7+3vkunvNQ3f00+TIve7ndiX+9uoqBAMhmZYLQmBA
SpJSx10/NOXnfc2lSLtnmn9k7RwKl8CuuDcQgt7YFi8ydHqxHL4dybGznFi9NSJiQx6colw7GUpC
mjLicp8kGM+a6SeAz+7Vi74wTUXnXmlRNDBZGIfZDGwTq4rD4qTcqZkW1q2UXJwLCyRAg8yU8PrO
N7425QPkMEPoqzkXaw7/pSi3/0xhJgHLLQ9PollEWMIKv4Kc6bGkNHA0f/D8AshJplD6Ct4lihzk
TNidPNZuBIU49QMzb3IpG8CK1EkOyHQ3yNgcX9ZKlgdayiRm591Ls02ReM7H9cqO0bXjBDRhbF5t
gqLbOBEDVAM7DuBk7gTABbOHvGlgSEIQ3fTBhsFgNNw7INuiPyHGPHAApiuk0cz3CmCEoQ++8NNb
S6WwlhcuEmDmkMJSBfqO0CDZac475E0wezZ68fefFkW/QKj9SksRpd/4h3dhKxeVWSiJ44iwQQz3
Zz1NXw5B7eYlpqjwTubWmtThFuDd9a0pXmCJ4HRArqqJHL8V4bUh4kDqxzXX6eJCPFmMU2x2/Muf
sheQfHeSENYDulKzg3hp1dEEhR+DUQeFYY+vLz+oPSgBKIcsVqVhj5DUk3TpDKQygvnsFZYSdK4U
DtNGk+nUFsjH5QLpv/CWtS15aM/h9cb2Eid2zbj2x7YHfTiwZXW/zwTAEcT4qN6qkyw06f0CdGKY
48AGG/XRHA0wu2//Knh45i+xuwkWxJNcqwMcII7nyLi0WuIF6xWPDwX/sx4VhoE3a8VHmr5zQDZN
3+Gh1w/v/r4BHCzsJ8Sn3V0WaA5EIcKOb+pRoQ1dlUJ9oyFpqG98mXp2Zc7xuPhy5oHNN0hefHYS
78oUD9dRs+oLTPOdsQmSh6/AYhTBzyMPdhjHGL9pd6lE2eX++FS30Dm/MtSvMgHQrm9VmoQJre1A
93ZqJ9UEcAzzQhUCPCygKTTW8A6s25aF1qlmesXQ0FwXDkwlC0fGkpXQD8aAVXFuKbrHxCAZkb7h
fUBrGBuIfffS3NxzBIzQSrIy4xU422f6EFvBuk+49NxuhOpbgOrJQySDU77iCZbLmzy0eeyyGdrF
+HNuMqTc5MR8CZCXe4edMlNRGhU8KLtNzt0yJcCRfmmJ6qfNgatu/NOUyelGWFMWmqbzhfs7CWQG
FI9IG39s+HZiWVF7UnBB2ujXz46QmZ88KE83pHbkdT97SAL7JW5OTHaN1kboM6xpAgKpeHvVFy/H
PgL0lBZzUOxVhSoGCAJIx6YbvweBfPlIs1wFN2hp4tq01PQsfy6MtqP6eOEYYVZa7E7VVQx2DP65
ewcHOo1KTwcVQzg8AEPqabH28RTYdAQ590dX62WQ/seGI0gP/Cz6f3lNLCQKAmrd5pBl59GGReCu
3VLqf6zCn/+RULdbQpMBRBF3BF3fSXfmIagOuFMTghZKCPT/t3jd2fon3WmTrj7+5ph1Bz97ATQr
yg+vPpaW2wujOhvIffna1H+KmONF6is3Iwkho3v+GrUUDmxVmoDNxgXwhEhhODQvWu/1hVPN8BbU
R+hOnZA80UAXrup6kAPdEfQiB6cDtxo3gOGQ/hLOGeyg2vreiiwxdhY9Zz4FUeBNgb3Cys3MyOX0
EHyjKVnwiwMXbdxLj2vDjGE7gK6/PH9YJ3fHygE0MV/5BNC9t3Jm4YIIQzxXhE9LVI6SW9yl50B/
xy9vAaBcfA6yyXsMs1ztiS9qAZzl3PoEneKzuC2Lj5aQR6cbBtL8stHTyZZZBapJeQrT27ofHQBU
MXo0ynS22xNyP6xNO9bHe9x4dGqusL+ci8I9aq5ldeq/XEdOtGwqJi9p/mUZvKyeSl+SC1/Xqwcr
V6/ApFZUtOpArBzZVpX2GwQPQg8uDkqefH+PntChB+TEq3nG9Bgqa9Srk15vSWfQ/G1mku7vufjX
XAv27ASgsNP/qfduuTHy+FdSHvdX2UM/Xz3spu4yMwju2ETeaybl1FzH7D3HdfP91QWViaE4xEF5
6VRyh2yoc2XUWaHbrY16SBfc38QGXfkcR8vLX/E0ruJ8/P5MFBVr2OqRYmkx5QDNdy0reN5XlxyQ
W18MVJAP0MDoVPi6qBxg1YFYE/SZfKyDhMC6l+7cXCL7mx8oQXyhx5UZ9O3zww2ULnNd6agfa197
9b+h8hS2EtZwFvVOGCqi5OxclS7kyRlZduIrlIc5jgw9pZ37Zn8Id2MiEtTgU+1B65dS6ogvQ0gL
tcpdLUrubsCz5o6Vpt4A4edyIXemrQ5CWy5PSzxxAVEIJlRR4L96lckdS4bRKqVHM6nu2DBW695Q
UBIq1oFdC99+UBz6jqCi1omMbG9ZXBsOj2TeVFL4Uf6EI2xDOm2j1Jq8zJZHrvkiu2aXXl90BFys
5HsRMf9It4stctmGSy1uxL+zu8szYKDjX1MnGplyUyy/6BMLQLowDNOPvjNxarokVxj/6MzmSm2p
b/i/CAmNiCHPuz6oYU9EEyKB2cXsjzSzgcC9hFNXOZew27U3XY2Bi5bKhHyCkMpliYrrjz7D68N1
cTtBBP0IymNiWbM0/GCS88aiJrJBHNEJHUH8fGW0feqzby7KlppNcGJDoZfr2JZPeqLXwnszdqTh
okOK1blQN7M85lvGqhg63reYUZYQ4s+6JxkLzhMYud7cJu/rzogNSVfVBTmAH3OdKT/fi4igIBeA
Czt6XeY/8qExPp3Ir0VIjhgrbIQBspNdYQIaWiyIqtvXipXcZ303ZtlWuHWPG28la2iCYbDVmlkn
cSkaLvFT7LLPEZFJCvzsJ8IS3NaEfYQLhGH86fGSwoUBYD3vNKu41uTqbu1/13ZcEzwvnW+aXdJS
+s48jhZNSmuYhVrf9gdfZ4kArV0YzMvapu/3SQHqoKfdSdeBmqqd8GkXVyF96ZgP67wI3WA0g4TU
Tn+hKFlgzwxv4kcLeH/KtreSx3JOrbmXB1MU6LXyF/8dPhPYznc9S39nW3A2PnUpmoNPbE/aM+30
y/XVycWfIf8ykIE4Qht2o9NhyFJWF3ZJrpIOzQLoGC3tKLoASnXFV5GLW8ESNYFTHPc+W1mrWWHw
3RWMmaXkmH4TPMNv0Wb4b/CFXxDRBKlgynTfY9VZBtzE5EJph7V6CouFoGBeWHOZq+0Alc+732sB
XmbA22DfMxAwZF0fQC/mytp245svRswezatQvTsi/ZrvBOPUjpVwMZwx53Jx1Duy64WM9CSqkemD
TOVy5eo3z7Jf6Ggxy5+MaYhF6z/ySz3kKK0T75IEPR16aegJSG18/x/ZIubuWzZnJkfL7SenT4Or
jmNG9XL3QT0D3KGE1AGJltAbfUn4Y6JEHyVKv2oUAI/Sa5/s4UWzHo68Nqj8qbWYzSBQeNZIDUf9
XzbymDHwsjpgayMVJZ/YSr8MuBOtGSEyRUD1JxCtEa0zuBN2kNViYdubSGHgB+X7PUgI5YM69Rzd
1z9TPcUhEO/AiQ7tL5vS5hko3m21mK5UqLqSedOjyOo2SoRvNlEpfOxvQmMLDFwk/NCdAmmikxmL
kjER9n6+gMClLAfi9sKa4b7D0bVpsmzeFVfIQS8KnA1PQxdo6ZYDzGAmp+dGB2sNnaOwOiwiYLzm
AnmCUVuyFBpJUIfJU1JjNSzy2hDU/OX9McxbZk+I+S+nY/KcrJIH4FA4KfVCMzlVrVs1QTThzAln
5JZNiU14b4x1pav61+cBwegwW+uksgIiuHHnq6Nx11vHdMRvyBWqEZ5WAQQm2QWYd3S4i0KbtYJD
sM5CzJe0p72iJcr/fCm3j8Z28/vMZ4zlIMsyNB1xYqVKsDob2jLgnGqP8LLqU+ezBaEEDY+BPKmT
w1MeOgRdkihkWX1Apgk944iZVdbVTc7Jee7sLGqbC+ZjgMkAOEzTDcTFLyOPvwe2N/TETgZEPH2o
ijRY8rOz+7zIaBmb0W2WEVkp8snt472KHiJwSD/HehqyXHPjUwspfaJZV31fl1GEuUEjQ/dpJoiM
+XgvsCBKVRCzFFZDp5NkaNtVb6a+dzbH1JX4iQ0nzlcg0EHMhkLbuwyBp9nFZ36ccgCx+NE45wrU
W61FdFN4a2tRwXMc3J4GCjWADd83C2v0fLNAGLkn8U653HJlVvxBV3eD9/QAmTgV/nTA2TDVnbxS
zYio7cD444FNTogUOg6cSm0rkIMZlP4F7+usrQ437hEgQQ3u6WRYXEpL6o/T/BLAm7iEG4AoIf7V
nZ0jUknscX1cUeFvW200GuOgZihuKW8P8SWWiBLh52VuTsd5aa7ytbWtcFTqT9mpIghDQXq7jRT9
CV4N5wrGRiQloOn22XnxfrC6aGAdQyzPGppGV638dWIpHHWqUzSCoepBQDTB0iMBOmVzcS5lmSwa
Y3Z+6+T/2U34nfAZgCiolhJnGyndAWBWxVCytA1degT8g4s07dkEgxfPLGFPbzdWWGF9IUFHbGjC
OjIYBTjlQOvRCJy20dthMa4zcy0JntHo5cieNzWa24Y+8vU4OERMszpNGMYdvxnYlBVHyqMr4v2R
Zep+jYs+k9rARr/sobrH8MHPNzHEJ4MoQa7DIoBq3V6f2Jx1UK4u+xTAV/Tvt0gfsNPNQDqzSwSb
I3ExrAgaFS50UsvLRVOkRrmUra3OxonvX8pAJmvM4yiKVpi9bWjbvvg1JIB2ggwhA45MaNXZCObr
qRcgxxzRy1RUWpzBgyMKb2pJtULWbUmgZihel0v+dpBYYfvZZA3e/JUGWJoc3eqYTFGlyabDJAqI
kCjsxdVUcZNNzw2S9vBf7a7PqLD+4vv+oVAaBy4woKoZAxpXwQXrn2Rqt3ufAKn32kyjcNxwhkM8
kQWEbPTsVOmJ9ymsrB2cwineMGEKNxQnpPpqrWVtBk3BWiDhyVvrl1UzPRaMjRijzROsr6c0m7vj
6+gM1eH/cLnHd4iJf8MWxcHHqC1dSzz3K/dakxsX7+IjcUnmaXcBJsRGrw8rE7kfwZZAUUt3iuhf
11KW+g9GD30+w0Mk/bACgtqQLcW0OvS3TYxSgOVwBjfkXSWhvrWM26vUKfrlyd793yQlnsfhYXt/
iY8b1u0FudtQGo2v/xWJSyTwUVfsogwKcCcSIqVdxSdQKyUO8a4pGzSGCYfVJgem2gnDhWzZuRt4
GfOYbVXGbwyZRxZdzTUQZYIhS0n5aAt/YFAvICXu/QJ9OOfsH/V/uYOvf1BYlrwksuA4l8wi6lxl
CizVVN0drRB5rBIT1XQ+a97XOdNrTY0voPQvX1n1yhY2beE8poIxJJUKKM6geAypz3aeSpRIjiEm
tgIZo8+GgSXn7plECpA+bhumiLB1ekUN4dX8DNZXNxezMUbH+TJa0Q7APsq5IZWoBHb21fvCwhUB
5fScT2slJMiBCtMh8KWP25Cg5xOGtVqN3LTjK4mn6cC3Cr8jykmfTqPCDdOqScwl+RIBD7kbA++4
mrmEhaB6mgUEODWujId1pcfwq60L10z0QSDcxCXglJ16Pz9vByNSL5Z/55uj4t86sUXnTSFXf5tp
trkOei2/0ZtCAsmR5Zj3Wdi5NgMNOvVvg+mjV8uagkVPVBfKHpmJMKQuNW2MRTG20zjtEDSzfg35
ibalyNyymfOGbllmefp8f7NAgQlGtH37a7GLo4F6jb++mH+slTSpG0a2GtzaNryR2ffW2HpbOeWn
QLsZWsxdLKjsZUtSAOzae3mcCrwiwnqw53jhMadcjTUUoWgmCj6UB/p+AYLsKFpBw91iyN+Z2DLz
eNAlgL8TIE3c7S3R+uoqhXyE11F6uTSJVuVfEctXVy8pJed1lzdkNqFVvuYe6n506MaB8nF1OYln
rNToD19t4Nzrha453iLj3b6FoF93I+gc66b8erpa+k3sCQLolRjVABwaO0Cuni8ijYaUmaW2l6aP
bxcVo5CTgkzks6dOWq3bU5rvRnqCLOEJf01H2aHtYxr8LgUbHr8hc3srkrgX4yqK5F+iNGx5lOXU
B/ONx+WYvMmDTl/2KI8uOkeGTe6N2r4BjkApyn+v0EJdHmGzqRDpUrFz36fvBSlHInVJCtTvgljx
1uDHAQ93ZOODNZOkjYm1eX5nKQcAPMJLt0Yd8fdWPzLuGve45bTFkA6ESM8QvM8B0nm1z7nrk7F9
X4AHqiqKSHzxsgt3Zil+Xe3BHYOZoJW07w0VURMnNandFgzsBm/IxDVDUMnsaERtWjd1wjJUThmL
FwdrxvCOlrRQ6D1Qu1qF1/VbFbQnuj/iTyOTbII3UCx1yCS1OH+C9nrXlvr02vheMxndBhv6opJQ
lQaLjERwBGiR+5ebU72EH0qKalxQjaAuqF72TNNPHuhQps1G24GYipUChdiDrW3z5crxrlLoZy8W
H/w1ezdkDiivSSudia/a8uAFNV48hS6GnbkJGxt3A4mmuX8G2cIX1hhVKO27d95/NmMP1VIY8g81
BT9KxBkovEFxYDI87bvkNlbZV2u7gBs8zUKV22lJ+jqvnnO4Yyrv/FR8wkOJT1wk7Gg7kOpCY9Va
D4Ziz8ivPUHWe+0FFP85Tf4roScIh+kFWU5rh7UqgUnh4tnoEeg03+ERMyMCaeXKbOUMQSc4up0M
5nf+KKmn8L2SnDN6cQkXWlyHZCeiy1+uFh+ApA067tG1L5Izj6N4vejRfp8L7tSKSxqmwW6iySM+
roRgNwdS30A7HjYLS9Aw721KQJMYSrRL0SAgGnH3QHEWZ3pKCm1RlkVuOGPdGGIQYI4CZxsMJmn6
TvKrRtLmo0sGXnOzkPDb8ABPYW54jqsPLW0+yagnWsBAP6mSOxksZHvIJXky810Z/Id1Ly52nxaJ
e1B9/4ASPnl5upwSlpJ7piSf6Qazw6fUxE7Rajnk9EA86Te+3E3S0kX1lWBEVfciWW0kPh5MNYWX
pN+EKmSMihYgBt9j9oznKC1LfNQ2JSw1HZtVE2B13An7Kv4QXO/kxB8MSWBRxgbro6NJuqZihfqH
ZJZSQi7F+w3Ayw2rQ7xOYtkJh9b8+m2+1NVoQ1ysb9e9MBmc8DvOoxi713aq8KSmmV2F/QAxoVun
09sQ0bxCT9swC7QgjIwO2wDex3YosamSHVThe4cvKhkJkqS5wuLl71T/Hs4WrUJqh93SBECh2FhT
D7uqWErZgtfjpOWRj3PFsEH+mpL1hB2SS58imslGYcFDLi7F11BzEHkUAJoMN8L78WeEMusWqwpd
nu7Uyf3Nmf++oWe34kClIh1mJs+sMz8JzR7ch6rG1r35GIKfUQNHa5DT9PIc/Dvz7fgeFebePyFj
MhusA/9XSIzTbU67Ecvpm4aEDEC8U//tAPPVx3CfjRg5EoqUnyUqa0Ghmt4GHlHnraN9Js4Bo+vE
ZbW+/GFlZthNfZVQUx2eNUejevBHec4IH+TIgje3D4zY/C/8+3bUuE49UGEO1pM1jbvJfC1Rsuj1
u2pWji9U4JYMjAvS+wJBaW1OYDf6Hg64drwi0cxznmEebGjJ8Q34PAN4n+DZfWj6vXZGfeQARkYG
shw8NpWgj1GpN+7x9peZ3P81ctY6HxTwVN1CZ27ix7Bv4sWlm2NqUAhhbLAPNyJ0Yz5AWRgukn4u
sA9wazrXpy9Z1hBYgRqOqVsqSHr5Oo5reo8tTHjUrLU/jUXEd1D/Od0z0FvsVhqjji/qDfXGcjQr
K3D3nDf47aIZFv0CJ0UOOkaTisFPQ3gtDXdJxLqPOstkVfKHrV69w/ik6iBDFfJxknEN8Qq0FLWM
QE0jqFByclx7d8BSdXCH8/LOxHl2l+HYGpxZbtn5jUmvaAwvqczXNGjSbR3u4xj2NgvAq+YKuepr
73zc7cvfA02lQoiGUWlqHOZlbhO3NYs0Aof2Q5SOqyL1/mcQVGR5KizHr1KeOH6oXu8nFYIXGvej
Pf1Dd+9gQQu1AOK0XZcGex/THd7/ama2a+URzZXH5S0LdshuiKwIC21Zud8/jCFw2ko4kRvd07yA
o+lJ2GfItOGHnsINpq1e6a0UXiozYbi0tNkClg9s+fLN0Y2l2zBbDMoKzrHigg9EOpATD7bDAoIr
7xDbneQGkrYYTND6XwdT+HTIfQ34Z6IOSu4ZkkHMSQ0XK6AXN1+wRoVkgfCWI7vKvKTrkc/shIOE
RpSlJrhz8szo4y04JwATu+2Aohj9WRtUhe29q67x6exeL19TdY6CLi7LoBv3Qk9lx3N7CSzG8sYh
B2j3EiTA5yWKkm7H55ibR0vHbDrzwkyVxNZ7kydOGGWx6nAExrVoJT6EDNE63O0KvX6GHbp/wuCs
Eh1DlZYAAOTY3dUkTKOjHiwJu3FJNYw1ysVaQB+ndJvIKk/Px53MuPhfacy0T5RrnUhkem41neAi
NDKOGoGn6yBQX5x4DJyynrEJmha8FaBunQtHloYagqcn4P9g5aBh7BAh8IDOmILfzPYcRB/WNlJj
oRzXd+fTmVZl5QIhi1X/5+eIN8pQagaGaAv2oDPISjemOB50Zh1THSYdvNICIRs2szY6xwWyj0lx
6/uazRC6hnJbPsq5BCloE01rOrrygxiyOrLBdTJIOUQS7NPOkAbV8srs1zc0G7QPIxFCGbK+ymMm
4KCz3OOl14mvhmzAYWEYIHgWvSX9S4ml0K+qEDlPHrdZXtarSVRwlnjtLZSpKrAvHKROHEAtpOzI
gente6C0ao1c5V6Wmja3naKAWWzhs+0CK8GTpUHBZ1fqhk+smw5jPCU9TgbOkxDueTkA51IHgP4l
LMwqOVyYnMZ/iO1dL7g/jfeTgZF/6hrKI2xnAGjgB1NdYs3TUpDNtStDpHeP6OUud7ulydcFWHMh
RhN55eucSOawysQenovBKdYIGQsV5eK6CtHFJYAq/hl26JsxoXLhxbr5P7/1hchXgJMGC0NOb2uz
j9vujbnMl2uCkf57EShE1Ff0iZE/MtutLHfmND1Sun4WiprUxazA3goHrWvKFdlhPbDc+Ut5HgNG
yuXSIe7/OqjSj+VFCJMbOEBuVDRsgZACQ6UPmbpPMvb7mOky5p4xIpUkxnB40i5LF8C+VFQvBSd1
12rJr+xFbtmCbFABkysQX9FJqC462hs9M+9WJ7VTh3dRm/VPZuEFZvG3hNI3+TTEn3xGVC3Z1drU
LkcMzVcNq7fLtO1lZ8SFN3HD/1uxdAmUYq7/i2tJlhY590eTScYVvpZi+7QR9U9MsR5BZNUO5nkI
AU4DP4/yTOBFlJyZs0Xbx0EIaw7ZdPBNupi8NzxxpKQ8XVzQUgbRalMyFr8j1AuNEvs3RFsoCM+7
/9n7K4p11nX4unEz8jckYJjVuhjMosJcb2yW8pbhDE4Pf8qQkFAv2m+SofRXYbq5bu3FIzIRGgKF
fZfEqu6v3pxwDfKyQ18XQyYuFhdjjvoXUBqR7tP4nMQKqTgtShw//+ypNA+0rfznkKiQ1iGDAlW6
L1xxQMEsQv2WfOXG4IXmxi7++qoSxCyTmaFj6xnxKUaJXpnh76iv5cyL13vsen6D+dHkpCD4KF++
r+yKKsJTool/ugHaVKvieei/mZCeyPVS/PWkHL+A3HTMUGLoljLN4wDOS6DmHJkbaV9beCc4ibNh
F6TDR2IBi59ZixmdGJuft5dCpCGfp3vVRUI0JxJtffbPF4EIsZKEqQwHm06Baboe3aTwMnjsXWJ6
KGX5Ui/YN9qtecvRnhyZsmU7MFtJE0o3nEaVPwmJH17+rLYBGhXsygrwPAIkzZ4FjS9gsy3jXgVK
bxAT/A9bmJMPIlLi8GubsvWGSUJbMBIA4AhNejcKEXC0beCqsT/0f+Z14x5dVWavts5XyQWCFZ8i
83VGI+lc4dLtEbfQq/lrTuyLDKaHJ4HfzC0mp1OCOKzM0Zj890ld7h/EVDXmank3Ehf8zmWwhffH
3MJ6PZ907OnBUHcCcCfgT4XMeNxnifB6noJIylAGOrAylbMeiJ00oPuz4S3RblOm6QNt9H24awNu
DcHL2Qhx4otPV0doSLr/LPPlK5x0hQs10omYudFsSEUAdtmj/NO63gQgpN8AhrxwviqUDAEs0/7C
usJ8EKuXBGkUVaWZqy4Hhs9o3JWYONUdNISb0/eWQmIr3OeWI9vh+R2vrkl6VJaxouMMfb34EcpT
wWOVKbfw/JYYC0g/pSxspbxa1VdCBJVeyjc11P5mynM1JgYgijXARSUNYW1zwp8RJq+gJw+mXr90
LsNmahF/3cc1uAJ8V4ym7TOXucfLOhp+JaOzhFvxdRO3krz0hpFq34dZd25+HBDlp8Utjey4gnPX
02GX72i6qqNYWe+/P8xjTNt0BnlSnUpVyJXtN6ntIch/brsl35VsNhaPl7fPUxOULlLTVVQ2NCHR
SQZTtx3ewWSfBIysiBrsgBFbxAga5RjICZDP3uzPVOHxxXKEJWB8ESns/twKSsoHFe8Okj4O+xv0
LRyAzBCT16+SBVlmXJJzrJJ9pbNXsCtUh39TdPvwdqP766A3n9CAVdDY6mmjoG/zj6IBd0fTT7X3
9tdSFo3Snz7Qkg08eHD0hGunV03I0CBqELIZ5oqdV0nAWADY41zyfUMhTOTTe4QE+jBmeSBP91ms
FRi7sA0WxjUu7gdu5rmGqlMWz81s8bLyV1OTtDRLp1DTXM7AHJmcJfQPfziWklawsXg/SZ10kbNZ
ld4e/iFbt9sH/ty84l2Y0YKJ9JGfscfjnLiTZj9yFrhn7EZZ8ktt/ZgIL6mzHb5RQJbQ8DSmLlrk
4yxnAIl8JW+NuFfOlxANgKNFzqQ8skiJns+syykfhDKpZ6K41Xd6CP0bGvqVSz4s07dmjouc0jL0
WwcIb+QflCL/IS7JsGpvan1BKbowDI9Z4z8eO0ycuPw2wWFJ+/IMo3AHNkNHXUNEEjdqkD8pQCPq
5zDgtRVfEaZEdXnyoFCEAsFceap9LvMZM/IscF6vtN6Z3+FYFcpHr4Q2AwuzVNUBBN0g3yAWtxGZ
Sj16MwY81878Kh+pvVSwIgqdVtr93uFTgWoNEa0IAhSonNuetSAJzhxRg90YA/+Yiw7fEyalXVYq
C8bLYD1/V+0qTocoh8+g31zIc2DbMmDJGhwGpqUQyo2Pn3EG3UEXBA09gCO6JjACLKpTo3URdOEt
61qOU/ocXh/ZbpjR0J4a61uu30NuQYX3L8/W+s1BzJqmvv4XbZGyImbFWfzd+NQMtiKn0Y/awR+f
dOVP4pQUmFWRB9wqlNe4CrRXnW98NzEUZskBrtoP4v0BJ8RLUMbWJ0dfleYzbtx7OTDd7SDjHpe9
BBCtaul8Upq6o2f6wuY2v4uS5VSQBJGfBHUpkjax9214TOqJpVO2cZyeo9R/S7cm4gLweRwSbJOy
Xyn7OnE3/c6F8PdOexp5A3gJd66gPLSb6hx1rnQVxVAoExNKxMeCSmyodfkUUvtY7IzlqBCtq/U+
2DjG6b+WYtXEmyYHzf+Sm6+G4WDZh+w7RiiEDKo/jr4eKuP56+wXC/K9JKDUbxx73Gp4DWRKcnen
kYmBoZvYshWqyaQ/9BfHib0AS41BRSaEWquzdWZBeDA1tZf08OzLg7MEPDXblydlsEHGFfaqogHh
VdOcgbgNNtCtWgi4/QjTaxqkQUINGxIyAhE5XENgrq6Bj+rdZHAbmv16ea3lYDNHJ/6s9wxydQ3n
5W/IDNixDfgDHnLF/2vXYsTkjzdBYc4ntIW1j240/UaXJo3aKpIgPnxmHBrXKI2ZQtza0zSKKhAV
min3xZiGDyEuOOPEteDqYXgvYU5g40aJboir30kJuH/ZHbxqFxUi8oo4Olz8gXYt/fMC5rs7DSry
1zJ3Z5gUNVvWs7Q9XFcW8AtdePCB7WsbvygcVBwYLC3T8Cs2YggGOvm5DOGz1qARnR2xVj9q22m5
yjKOTQEwDvtiMA8gqz4EvoJ+4qOo1B/cGgz4BnSeV8zEJRgLpImiX1lSk6Imnl0jkUTlUXi6CBfE
txdPQ1uofZ74aHFO08cleSFsjefsFF9To8WUSJbedX/6S6khgR7QX/j9/VpaiRDMMDmJVWvQi0OR
34MkFKFS0PV/3RqakT5SmwvJnvGtQTncR8P154OjUEmAs8N185LIv3+PpN+wOEofhAawvA/1z+UW
oYOCuOjCIn/mQVXH3vAq00Ku8hM+NsNGddNyQHSI6MU7eD3A7Z/DqdC2FR2aftREKtIOtugtS1Dt
hk7ss7m4mdkD4roeNCOc8gBGh8DE7PPJUGCIzNYPxSxYWL/7Zo2/A13fuek2fgk8V044tJi7rOxU
29IxuDaowXDnH6EN6D5xgTyDy5mlBvd2Fi5bG45Fybv+fJ+BH3TTub0D339e3wH5X9dY0qdNITQP
aPpHrClaUbO1DG+dffn+qgm3fXDJYpJX7ID202kZqz+HLqZsUKk+QQui5CF7aPm7p91cHGFvLOgA
wFj7eYAHg2iKS1aPYIJn/MbHA8faBjUVz//bH3JVbaPX8b49g9l7hMAYcvDEclrDs8/Mom4INzaS
ZwJ2StqmcfPfs9Qo261dWdR5qgqxC6RYJJeOgeSx/PtYo7VzsBneV/H6dquabmEaj8rY8Ger37hS
Yt15pj8xXbCHkeYJmHqyk8Ny0hNysfrj0bQHXFgqygYLuL4u3AQup0Pf25LhX/WejY/frNLtLsGH
WPz4CiqH8qiynvPhMBHhJf6+g8yEeB8HYhIW/0EXifgYKNVOnCdyhysvggvm/qWjVrrEYhQqV6AV
igq1zIM7TpYHyP/lxRcCFQshdFVFneJkSStpybrABXTa7RpiiJLLsk716b3sEnNALQeKnSW3XZHW
DPxAuGfHoe+yFILIESpL/N+Ze8ukU8e3W6zqq/muQ4LMw/Cm/ArSZLZ9sOkxN2L085yCu+KsICWu
4E1QXx305+QuJhYs4hbj+I6taWWtAvI4HzbdnB0KWEkioEDs2ugvPXqlFYwvNsA2LObhaCDrl4/R
fNACW46UbIUpp5wGuEkWCRVDvx7nz1dHl/PNgMrGz0FQtRYEQVjC7fTtZJ0oqQd7o8Mqk6bUsnWH
7dsIJmy46gYx1lF9ylFxzh4QsLq2ZXpV6aXH3aW4okt/gYtLyjEgb62pLCGplUCm20exzurUge4s
7svkXFMSrgghNUDM9Ed/Bm3Oo2Y4I8vSCj5hOKWfNNRChuq6qBlKoV9hxvdLMV63WZRCybP1op27
rW784CqplfpdBBh9O3n1itXCJwoNgYKXJv6kvhBpVCwINiy8bcxIQMN6WdErrYZUE1FxHZmJ3fqJ
2OOcjMIZfgmZsKxnO9GLeimE2rToad++GUJidODXhrRLqM5A5QH4hxfpnFTUb2XyCDb8QuT4EtmS
aS7iDMzTD1JpNCe8sAxPBPjaaVZp4aD6vOo1wXVH1De1W7VNeYKYtNdUrGNmmzsFM9tfkXAJ0u3M
XFM6qQXmvWIFILfMEKvtI0MCVqIjWroABReD8J75AoWjzObgJnajZNMrzzs699awBO77+oPNISo0
igTjq1mHCkf1fTb1AxJuzYnPPAdC4yQDspY+zUDsQSScHYkp7kNuJB1+mnw2q49j5xNJ0dSajDdZ
nfgv27PLwb0oO1WB8jWNjw0B6NM6gkKjYNJFUXOexxlDj0ImmFZyYWN68bG+FtYG8IDi1HfRwlfY
PP8kpZlao02+cJJAK0PEX8NViZWDHqqQQh1JyEC2UF6RxmpizF2ozYB4nnwWSmlDTjFR+pgyBSgu
Gk9zBgNVFTJhc+irsgUh8qVwlVmXJfdJoPXDYbH/7RvCqUI3Ef8HSl70QWtCInFXALlrfefufPiI
HnC2mz0TuXM33lXqCzIEHeF7crjvnv330FM4H4A56mk/g+fRuOjl4YX4VYbUC5OT52ty/MYUc920
5yOyAPs+M7ys49UNu8nng83N/7jucqqhhZc8Z1AvWvxkKImSypLsiAK1zfxv4SYzyH+K/e0PvMAN
MnLS/mexw9+BBQFGe5eaMXafczLmA7fmlJDMOljrqGvQ/l3Bfq/THqhot/n4lxSilq4xBH4hi8Kx
oOf02MgF2v5LeHAx0XgnfAXGuRj7PdZ0nD4RTHMXOJWTxuA4JH2kXlFg6jDLsgujMG+aPYkoMlLg
31OGbGa8mamu72Zom8o+Rqrzt2Qee3AmOn5wfBR9OQDraDVaTlX6PXIecmxOjLRhVlJXakq7EJ47
BY59GUW9EikjIfDZHSG6cz5pRzjIivwghl/rCGRakeUY0sWLAF+Cc3JoXXYcIFPTugHkkrPsmgyC
feaBI0O5zvkyekX0/LQYxxG+XfS1t99XPu8IYPEMO8RA5UHXwhx6o3YoF8bUNi8VzPuJNHf8fZ4P
BE4pdlYDX8l2hRcZ6CzeDAP8Cf2NthVBAxk6YUJFbOhKJNK3HuwIljWnAdJ4jzF1wnZjgcs9leJ2
Vjx3ai4JgdbCsi4qoENfFZqtOKm1fbmjKcP5+hf4t7B/Vter/k8P02MwX3Bd5h/OVIEdI3XLYXcK
PZzc57NDPNcCHP1xpuTKRxrIXzrV9uF/UaXpS/C1f0hEa9IyPaupuwbbO/ykBTLDwd4p//WRn6/g
HmDCfEcJNegKrarqQlxCo72Rer/clsMcuvxfRNu8q3PBpj7n9CcljQmDZibjrnOgwkyLeP/m9I8d
lRVwph1h9nDOi86hbzOIrgDKwUJ4igzwp13aBb5WZ2PYug45a5DMFQGR0LznTiD7HTdRXhnbBXC7
+04lirQa0IZ6X3q1gteWD0hTfWO5QzZ5d0/STCzA490I3SsBXAwCL7uh9QEQWpdUdMbIuWWoQYUA
L9nu9TkrOa8OkiiqX00xgAm3VQqysn3iAJhD8AnChT7k3P7fr27PbC7QR9SGAbXiSYURHVROQTc+
z4mfkEOJfp+JDpqgCuDtY4qtZeGLrmv+Vg//5nE1QF0zdFOgr2ewJX1WR+G0fs9jwEyTyhZlINB3
u/OzuCpQa6wQrOOJnS+ZuN9m9ZDiPgmflGQLOE7N2AaisKwTM3SNf8lvywWNVCAujB1007F9cum8
QKGuAfgcJvOEa0lP1Z+ohRU0UMrQM9jvWzUzAMReymEoDfIEpwNFKq5xN/wQJwE/e1vL+3VqYGPm
fxGnxwfgoSyH32Iy/Ib41iJDAT8MBEadhMlJt62H4F0IENAuGXvpPYCVDiP/UPeuCNWCY56z3RgW
xCIagE3/Z+Q1cs7/U4qWdu/J4tYcDGbPd+SkEws5uSPe/yLIyz4IyiMhfXLlS9iqkDp75n394698
IcPyIUs+QdHSNUpWOoZD07aXOdoomWdnpOBnH47GWjl7JQ2EHe6K7wdzHejupGkpmtMh57yglmgt
zn9fsRPrbAGr7gLspQdC3OUr8I0B91W0Bmd48bFbXnu1MCIBXJLFbnM4akt8wCieyHcOp8ardnrk
dxQtqPIUfxfwmwaIrmLOatkcUqQNF7jilv+ZXAMNuamsEZAAOWgHjhGtzynXGv8BC5TMFmcMCDDJ
YNdRUYoHA4rftz/Os9WyW9qO3HQlqAFPEtPDHgSsUHKbU5A0e4lc0CllCFW/2CpDXK81AERonYrP
fdbijLvdu5E5qeOzaqdQ2gQfqhNLdnAEd04Tq/umo5T1+2HzFveJbpPySOYhg9dftHLasefWSIuk
jvD6IYzk4VLkekEUWsW4CjLDMX8LOZgeGkjdWHeW6jg22KHj/gtz6v/c4RmyMPZD6pwI5S0JrU8R
rl70qn/PIjKopvGBVH7eXqvOOTP8V9f+1vcBeCjye2tiUMdexvqGwC7coRucka3xTg11m7dxewNK
qSixZedNv8npz6PRAHV9/mvN/H3TZHQSgaNQA6OKBc3HkGTA39I3vJjGlyW0vtS6bvsAkZv3WCYx
6Lc8I8A5oaTlO56fnPzSM/GwG070Qqdx8/+FvuWWmpRH0SO2TiqMYUcVPxfpq+S193SLNwVKxqni
IXvcYEh4bZUcPxCuvUsKCGDeAR1WNl1JHTi6LaFAjfV3KB+TpJgNu508s/zHmlNdhhBCxmx5YYmH
WyYp0bdMV4k+eRjsFsKnmOY+l/MDf9q4lpgGzIsYkSqg+EjpZ5NG7zEuKWk7K5S3SXrdmvGzX9Nk
aKVuHEl1JoGL+SumfyTkhki7TXM1RRQQ92sI5YeZDptg8SnAZejUlceRIw40sEmmN0hCBG5fvhJR
KA/PlkOJRp9wj6wY+/qp+PlrPdsX0xp16+dzfMkT0j+7PQlOv6URB6/EmVXAo6VFGm2oxFIxPDEX
b1GK1dfVW1UMeEpoVd0NTTzyEjmPUaqbhulbLiX6vb4IVDovb/1koW2P3P4BWeF2Ogwxx2mn1gk8
M+TV4lpa2193CP9BT4yD/C9pLyZBZONpUoQ3+Y0b/+AvlzYW/rAjxU2Z6pD7ZTjNOFrgqeTpGEq8
tEzksTQ/LULzzDLhu+Zhg6rpkQDS3/cjb097X9XHCX+7qEX9vW+z5VK6CSbxe/UzCzR391fbppDL
CAojG7dEjG6xFBxg/Aw1Jc0rvP30y4JjGWiYi0IkTZycCFI5Y2MBz5ENoW1RjelDyaOWLphQeStK
raHDNG8kjsPuUHduHHYoHFQsbj7HiKGOuTIDAsqBIFkH58Hmx1ARqTKBQk0leRmxLMWPD4YA1QpF
zoyeW4NiNTug0IOEpUrh2UrM964zBeMfeU4k0g1oS34zPooY5yDs05dX4GPtbNWv/WwE56n0OIhr
0vaH7uJkaCaeKHefNMwtG6BDZ7bWPefQabhQVx+wVYKm2IIjz/ieOmpn++YhpMHGyO4UYIk5jma1
e5DriAfC7+A+6JWMR08ehQj/bAMopYRtv7k0axH0UgaK4jzlypRu4URxqe1xxswbz2I2NaldX1fv
sdnxxMwscbUUcstg8ibMB7ShIT0cL6wfnVBs/qWjnGZcsV4w2CujRTwnQhDDsISHXx09t+zHOLiZ
fit3nM5+woL58OIDSF9ZH1VGI5ZBq9xZxPT0aKCuJxpit+qTE8/K9zpPTAa+5PYRUb46X6KoYIDQ
I/3o9CVg9e4n7QaLe3wENQ+pu8jYCvR4l6TV5tFWDMQyjjAZW7AojT1M5/JLqLF+3JTGJYWx6Ov/
7qHGd0sP8zG0H3Lwgt7wQk2Jfh1sQUAjpdDrEjiHySwb53CrwFqKJbiMh6sBG4WvNDNBA+s37PYM
NzBPzwqkoFyICuXclt94NsWYtyx5/dj1uaYT4EgChUZ9Y5n9rKspLLpCxzuo/uWtVeOwDzSTTGzy
My0yXIcpuhtUb6DMdViBpq6u31r6AaGIyitqrGj+1L+5PEquPVVQkFlSr8d9GKCnKYLdcgHAYLUR
yXbn2TywBid9Fa0Qih8Zh6S8sS7kQeSszwaDdsbpyjfArHk3IxRxx6RS0RYgGSgdrCVPkLxyD4Li
O6FnYXCdxs6pGenNh71p79Lv+MFa/2nE9MWa0+IiwhbKent8Vfe9xmPVESlW/FHRkniE/vVh8zOp
BnvDiw19v0JWeItcpq+itsQLMQ/e5Wpas9VH0MTC4sHwZwf67Fo5zqlHgtYwqmjg5isJUKsPEpvv
A55BOuTEPoFvZ3sxBPeb0sP97QnY8yjIaTFrWjTOZvOH4hL1uu9EuDaxDQ1ecpgD2pttOfLro7Cw
Q1kHBdRAxRH73IDVHiJ/PMz/7iw8yt/LdxEWRnxeV1UeX11rQTTf0rWeLyHTaIcvlFMJcteAtrCz
GaR1NCQDozXWs2x8iMrX2LbiDlL6PYZ0qMuw0uYMalbmaQUgb27KXqmclyhuYtGO6My88khXmTY5
fq84X71RRZxVMuP24tFXLtby2TsOmp35u1+0GMCbzAjFDGDafMP02Ss4deMvAqIkh/8ecVviEVNT
Ng2xAj7GFCrNfenRQVp8ZScZDVXWAXg0zwpi2HV5+jlKDHnCGFfdc29P1VWkYOrlKlCo3GwO8vBL
gUeKhvvWWuHW4rsWxT+24dBKCVeIBnjkCvQM/TwV7pRjp2/QZo5eG0IxfUU0mP8UmDN8IIJG5B7v
VVjtHAHSvQSGq7cQYl4RXok/C3wR8wyRh4g5yg5Ul4UctkzX/O8CX37q6QCj2Q6EPI2OTFsZlNPX
tTQ5MvajRBa0jyQh/aGQms/sSNneE0PfANICwYmwwa3m+Q8VJqI/WDGuYckNziqV2S0Dq8RcSFXA
cuwhD7ku4JBvkyEj8PWjTUWc8M5OJo8xT9PBjWi0NEVHKtaFKI3fzmtj8OzVjYL30fwMg6sMC56B
9b3DpHQFwAJkeRQEXsdnGDlcQhOiIWHxWXPm/WBocWs0TWCTVL2JLxzsXF9ulPBd+K6ZQGvD7ZbO
eXZ5pcHQ8O5bgigCENL05+X/YLNZuqKaa6d8Se0pz6ISU6lkUBRzy4kfKdnaZbLdwsqbN7HSB83m
nX57/aldT7KLewuG2dI7nRCAwqD12S6vxMbJrWKWvPh4FeCHwDlYxRSrqbiIgWnL1grCcEZrrJm7
d7ftaJuXcuAssCapyJvHqSUe7czcTOmB/pM2uIvEQXOzx5ys3mxYu4IZrP8tafiznVw0HzzrQpaQ
CXTqUMrjBwfn9lLYR0NwdPxgQC8K18329MBB3S2qLkwMCzfusRLHYMx1w4wUk8tBRGMU7+fuIq8L
nm6Td8gHmauI+noMvxF4PMTeSUtyXHKDWqzAVHe5Maw7xcuTTn1Mc2eQfpQ2JMHreZKfS+GKv2mZ
vI6q03QMiTDmGkCsrfBGRRIGvpdc4vCkSK0BDOxKcADSkaVubgEYRNRDew8a+FYHfhEYL4N71+B/
GPcPxO0SaKIo+Fo39z8Y6+yA8vmelpqfepgvF454yo46op3QZCbYxr9vkfSB5WTo63+kxSbhsOt9
VFdZVnlXSlwzS9iFtCQBugg0OC9QsZSfCrP96U1C5hKOLFL7eiwFPc/Wos4JcHnRixCAUPVL8WjW
Wa8/Fd2dDIW7m/hfw5MA47DkGlGO4M30vIr97Oqgc9jmC+KixyL4R+KyI0FFwWFhfLzEE0JuQcuk
xj3Rs151zRkSPF5TeQL3fXjLkcmZcvyKQJ1EkCqnLEalrGembxuMUTavFaSeDcCM4qjAmfD1mMW2
AnRq/+Jr32SOQ48ICiui3HsL1efMPtK0WQFDQqXZSRc3Td07wxXBWk328SpN45lvTSrXw5t3s8Yb
Q5CH0nVc+RkkX/HNV0HnydBM/jrcXrRgAr3lf4BZFAyJkpWqt3C4EguEE2naQ/g9mKpkdHsV0rYR
EOh8vGzwxGLA10ONEKAfUB8LY5aBljL27ivgPNisWQi9kjz812Ob1sCOrxUQYuv/dTWAkY0DoF1I
52WGfmPrPUyvWAsneHBNl9tv3AsKtZNVZ2It2Wz33g5Z8791STi7nwpJPSoMUH2+8ttuis5J74fs
/T4WbsxU72qjBaJhs3YLngNkwtZGK42zJRANUIE+eP+P+S+OTzD6tyMv3eP81e1TGBPgNvs1Tqyx
0hH15KK4ZDptfOB36yHIvs4DxobG+HN6epdmeZn+Csg38y9j+SY9lnBOOtVGXSckYQkgf6wj+mfc
DQMBYPVrVSIcSDsZHPWQoS1ZU/xydc5PJfHllMhLVbJBig31nnbBWRYin9raey1Y/F2KHmPq8RGt
8cl5X0QjhPY14d1PfGVh3zh4kTXC2LWyFWBN0Od5wfpsOERU/nWLrDfeJvTR3HDojBiJGOZkQlmt
mzlBfGFLQ722ydbwwdGOQsTl5dnrQGeQ2uKQAsNTGD8nVPcSbn84ZX4QyVgB+V3PFGDIUAV2PNgz
NBSObAnGy0GJKgqZ5pCM99swVI3whyHzmwc0U9uxSX4uApk/y/Zst+nLOeTlTQ6d++nosnU4ty6i
xbsuX7JfojNFVOOF8RmzUdQvf3PbwnlSOEgcq0pp5uPo8h3me4JM66jsNvnhhQpalQQF5ep81Ocn
VxaXg1xZo7dFOzKQ2ICTRMQUEyKci0URAzcIkC1EhlcL2b/qgsTcACkT7j2ydCbGPWfPzOwagXUL
UKPoa81KuG+RJwx1sio6Xx72qy4oS07Cr/gYUe05+bohst/pQmFTN09ysiK+HKceWcTrMweG7d5c
DI4PBRMZSkc8dI+e7U8Dw5H2vmnCTjD0B6KVB3DDaE3YDcD5hrazkqbBHqAfCRgZlCo2YVzQpRk+
s0vsxgxOyymHYr5ScLPTwPhl0pU1SqymmG02JZlBqBWpVFLz5JELZ37Z9kFx4UOzB8z1vbRiCbO5
W7IMrfSLRirSJNZqOpcNkZ7UIjpheFx2Jfmca+l4RXZR4hRcMTwSGczCreJ9ETxDN6/KhA3BGlyG
xVCnAMmW8CGINzopHbWXhvosuYqk00Pyif3hwgg86G9NryQO2d5c9uU1gQErLxnmdDYcWs9d0TdJ
8GUsTvd/4MchiUq+UNQfYQbnk8wmkZHmJsmfgRNqGdAaRM7N4qQSx2kxy/hu4jetg0YbLUTt50dj
Znmv518iEdTwIKp2dSWGUeBWPD5WEq+mB5m43hPUOht+rdZUqcsG4klWfKmWUT9eGZWuw+oD091U
WhIaa9HPGUIjM77s9I3nBIXT4I/RFkPNpf55aADCMqa1b0yCO4nsttEGu8gLIXgTm+pbH+wGF71U
4Gb2sq5WdVdmbIVETb01lajbTH0Kv1KoHtrsOOHXqpr5MtpCPPOaYkVGQybq2dDYLLRs55L8HDSL
0TV0uEzG1dE7TDRQKNPF1FIZtfSOlGPuaCNHkTkJveOM/0iulS0wUE/8lsVAzTAEOVT2RFroO8sf
Qst+WnatF/jCXRXLZhvdTrm1ROevs9RoKyvfZz+n8lhuDZVsmpFy1UBgcYQMTMth3GKYGVsYBu1Q
vMSybKC8v8V/tKknRWU081WiQcRHarm5bU835MYucMmx+iCb4xAqh6yZ6Yu+HZ3xFQRueibD5wWj
HC/uKEZTTjD0g04xWvN17dQj9eXTOhoS6d3D2Z8GPjJxarv7pI1G4DfcQ0wJKSfKkj+xibrut3M/
NQzHxBYbvlcYpwERgK621fgK1hp9LwXJkwR8K3YFpxZQ5oofQwtLl4BFyCI6+IUcUXBaHVow0nh+
F9vS2cJmUV+U/RmvoavxduJk1kVM2Qoe5adSr99BBnZpMn9IpW+4maXZs3huS5JFqvYhRUOzGMmq
KbZ7sUtjhLjF6fDmWyQi1c6z4Np49FhqtW2ECN/DtqdiAMOjVGE8Vddw5Rz6uQernFt8NeYpbaHk
373z2o/oVlHc7NWv5qqL/G1CzQU2UPjca1CLxuTXqXKXOxiRt7MFAFabBC2qPDocpfprYHmPtxdC
jfG3NgQ1LsaC8w7COd41ic5hMty0uyrH6C/7lL90okgxJZlyac8q2qa3/t8uSs/+dKkCQ+Gcrsms
8yVXO6seElTbIcxO+8SGD3HoS7mv7UuoP0A/Wp2nO9imnENgqcMe2jcQqU+HI7knb/8jkz042eBD
ThqKwbQcXHCmrC9kvaX2kEH+XfaTYtfZ6hl3aWQFk64x+rULZrqgaZFjImUQE6hTzbrUqf2MSBkn
fc0aYltxF8/fjDk3dJ1A878kTtj7cu27jDb4abRurItP8YLvp115keWQ1ku86YbEgnEgq71J5Z9j
tR8zDSduYsmlc+IgXPb8B43uOr9ye4KkYLrMYA3bIsKExN+uTO4yaScevCmIh67lED/dKLkJSN3P
YxetKazUKy8ZEx+iJF2XLm3AEL1v4X7K+wj6vpWH60Aeh/IJJ3bb9aq/DTGAblENFytafZVex45e
J+p/R20MJS7OrEUNKR4NOTRqIEqPkfIsb7vE4KdbslMvat/zExWWIsNT5Ig7knTiaTXaSAuuyBj8
cljnktbzJeKLKvNoax6cP4SL3GZhZjpQPURib8bcMPJtl+C4AELkr+f9yDtO4kVOFGvvIVXor3mZ
K0+7B8o94g1a+2ejFY31ghUtc1G34qH4RzBfxCjua3wJoI3nfcmWWHgdYzE4bj5vUGra42XJX9a3
eGhZoYHb9F0VGnkNjUX5Raucpw54mLYqFaqfhSbllkAoL9TYPrjilZsZLmCLKR3dE3XLc+y3DU6r
+N+mxEEbqu2reZHNhutO4vCtQ4VLQMhWxN1VMMVVd+FsThPRZLJlxCwYjB2WEL99t3QllsD/cYPd
OcXfurT2Fh7WO+CTCGCo+g/0jMciwxFpc3BtqlW3bkGQez8o12TD4Ipwrky26Rm+KSH5PLQi2P5H
JMVkPYN/dkD1QaOHy2qFYZg+4bj0Xe0xfKCjZxDNl4Z5PPI3m/yTGtc5PgkKAvXz2PlABpmw1ds6
o8PJydLzvTXIisViI/Oe/QX7tpGbsSBYmPv80BUdq+0CbBhpxAsj4ElvH5SGa+WgC+bwFNnyygXV
YH7YZs1aHKpi3Hc9pMrhCArBUznrCZ5tAIhrAzeNMWuDilXR1SRT85YQg2UlCf64ay7VVbq5PFNd
KmA5Y0x4bQA6C98QXhCNwh8Zp90DAI71HkTbEED58KJoHLoEWf7UhgR42tLT3ZpUgUAOhFcbuP5R
sD1yGSoSZW7YlLoB+waycnhhR9LAAvVR3d1godY+iFuFIBD/cJOiUjUoL1UWYk76RvMvPf++yeQY
hyMA/QPBHXx26VJH9yZDyjd50874PCW+WrrhvbP7YxQ6HxiJ4Q1lNU5WSIcX8LN6jvTAev2n7OZZ
YjaaGb/ZIxtwmrXVKbkbHaHlkXQ+3s4YU7O6HzDto3a28jEBMcCfwCJr+G2e/ueT8gtERllXvebq
quCLV7qVewxJZtknXuh4CnFYE95/N2AEjW3RYKnPoBgxzPzgaYAjz0uuaL/H/y87osyC0KZRcYNm
fq74FpoDjllmv6ALsm9Wc58ZlAfYd4V9Dr6Xy+U335hgnflGT0Kb4CD6CM1L5gPrvk39YixfZ8pM
FTs3/LPK9noxF5o0Zun3M4qD8M6vz34zQosi/bqKtOdinoLejbTsF90oQGyrwX8OYqn1TgZdHXBF
W/t4vdY86s49JGDffx8+c13nc0puSipa5G8tW9EA6b7tAyVkDBpfEPueDyPyELtv9CG65Dwyzwg9
GvVV55KZWPQpU7NXb/fV9JTGhS/CHj0LsFv5FfHuG6p5btbeFW8TkpKmj8FfjsuA2qAZYVbBYrWB
JtSVyl6BGl4HAhR5gBtNi1pLuxR38Ctg/vqR1UVTs2G4Waf0oo1s7V0R/GPFvo/T1T3FTAOs5TFT
Pci0VsDKazfgb8r2ENzr9+yWwiEBsvK/ep3CiIzFXXnwHLIj0LHh6LmaP12S2CaAYnKc9Xl1FXOZ
5yUttr0E6Dwt3SFI77e95KnAgOXJO+FRJbs/h5Jh0CbByC40cxS0/UkEFTZwtw==
`protect end_protected
