`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
fIqNO2NIgSzvZbay15b2YuHOkehqwOXYH/j9PWOqzH/rdWiGewzKuRZh/LbQzgEhmETGgmfvUMK8
IEXZNWrC1Yejzi91P8D/LpALCbtl9Hl75TLFL1CwkKDrV2eNS1pR48a65r0k/TxqCg1ASUyXkMoF
dEY4Wg2EtMHrYERDYl2l2FKGjlwas2J/BUrQXMWqZApHDvZJEsXIKSSIzFDWjs4Q369vOyMF1Ksx
twEfEs1USkkeW0BshkrUmTcfnTfwrMkkUFX+ear68ePcpZxmtqryMKx+rafRt3uFib4E4cTkU851
ZqAqr429hCqhAwPY17C++jteID/O88ac2iqx1w47eJawg4DEAcq6ceIm/wdVO1YoocmBlVONqi2t
NfE5/YjixyM1DoRcV+Js6I8R4k6+m2SDvoUEEAmKPQsFDKUtpng4MN8URCg7x8DDINhl3/iZwGtJ
xpSjQqskO8EzHXe3l1ITyBAKpgcsLBHYFeAxq8IGt8UU03O1aKR5w8LjBlmeX2aIAyXYQ5gqps4W
VJM1tENtARXws8iNJGii+4Yo6BDcKXWzqnkqmtfeFGPUkDNy6HQ/ZlrVRWBs5C6aWsYK7vfpYiNg
lrarBdwf/oAImRWo1rByft43Qr5HqoXvTNO4SfYqV6bs1PKQZAxv6b0vPU0oEkKqLfyH8M5Taoup
FUPPSo7o13JMBIMZGq4BzIGRhEgDQpD3eNMz43Ykv95sORObT9hrUtkVIxcQNftwL3tMKJ8CxVPb
WlKaxnWgH+v8Ht0341Sf6k59z2iM9n9LwNJHoZC9mKPb8RO44XIUkBRbHEx7bWxSQiR4+1sWE1jp
Dh8gsSPn8+NnuGbhuCCZzVsUmP9frpF4PVln8frjqAJf7o5p+icl/tiKi0+sWBh+zvAiVUMKdDz8
Q1s9AIIAFOAofl14OQVzQKiuerUSSJgFxqSHX/3yuIscy46ePEoUtbz5BbjFuSD0fCPH7UaHb5Pn
QjUne9aMBziQoyqOiY0xp67mR/VF7txP+NkXWHXRbt09TXM0M1xQj/INcbna7rq/oSwBwQpt1AJb
UYui4pj7u8vZwlFkx4hHiJ40QLFSOZS8ExCzHwPEtXtGRxT7R0UvWKXup6Am83Nr04Fs8jD0Tzg4
EOi7iGneX/ptH76kPYQVo5fNhoPL9bJrnxajrOPajVbJ8KdNfsjJe3JtXIe664jGPRv5GTmu6Wkm
YfAaL32Fg/fUZDdqCVSJztt3R/EmxX+/jQcoPUBvhqwQufuZaXlxrpAgD3pcm+F68irri1iMKi7p
uhOFKVHUUZUyAd1nXjF54pnTHy0rbZ87C0XOuv0u6M93EWWMNs/FxlDGlnBiehJScv23ftbjAtDv
3DnX/k5zu2HpyE39BVLDvWeE0ePTXDzCTMv5aCbOQNalP69Mc1Azzri66EwZXY6ROHFhRgaQtrI4
P90uN1uin0z9Vj/Y+4Fi0x4xR6jAX2My4AZtAWCvaRSPBra9Ajo7AGcjGpHWFDUIF/asLNRWSeVc
N0uCH7SaoC2LvB2680iOnOwjJSPNrwGogN7Ptn5G29gzOGP+TltUB8GWkYY1PtMbyB7pzxssaVqE
ZtNjK3Lgp3vi4uwOE6VzI2ElVjK/nGTi2+YciJ69I626XmW2yMDNyt9EiY9taucnL5Lkf6ldP3pE
3U0hz1LxoiKZrfgFuhC4s/80STaRDT0/BEmjtyDB009mhn2ZwbeUBpx/d+Nxc9VkYdaGZqmjlyQi
9RYrzyfSdOdT2uthu+KlJFJKAd3x/nL3chJoaboulNJ//AmzbvKGOMJaAAabOUCANrDWr/N3mS7y
f0R0L6+QO/uuJxwcXP7nQt9Ry4xb7vpcnokFclxiuPZ6QQRs3LikzAbiagSfJ740/hDYBUdw6kzV
PkBvfSjU6Hqyh19wtIZlf43bE9gtEHW2LVtMDVS7MJ8Gd49j4gOtfnbB02PBvCH/pq7mhGLhr6Ls
yQaBepv3M3Kn/IGrXpixv4ip4umH2TG1F1htYIPA4SyzJm+cjDrymhC96bLyKcbnIoYOCPYCaVvZ
CoQ00HfSsSkqBIr6biABBcOeP6oC6IlaD0mN3otqIifz4r6mrsLxHhKAnD2F
`protect end_protected
