`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
i6fJlyrt1OGG9qNLnMVUk+6GOU0ceijDxNnrq7Q1V0DvVQgsBtbkBoQhj2ep6dQ+EZ6xdic0CPbM
hW8EXmEgvdYzJT64ZQ5apFa6Yzrz0abeLfQQD3psEi4ArDpz3HZWlYi54BdCvB3SCbEq1Aa61K0z
7pkJ2LDO064fiq2mrbCFCZiIJAwCC2B3NKBZxgSwReTJQG78YHWjQtY/qdwBmYKVc0m/hG3/TaHZ
/sqncyQHXh2oU0LvJ/ro/K4Wu0c1EOrLUF9BUCqaLkdWLIJavVr9hCQTGNINe21SPNqy4i4wvFHb
6I0C+LCooByGhBv0/88X8WB9T4C5SLUT5IzxQw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="X7mFmfYh2TunRWEjzJVOazbaeZf7hz+6ecXhnAZKdG0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
Cp4/AK9pibK1gXY6JvEJZDDCwMLKhVFrHlEXGoqS9GhJQ8QTGArzOAnmL5fQhlXLYgByipqZcO03
t5Wlh5RkchKxeR/38+MRWjcm6BbRbKsMFahqBbqrTBoQcuSMB2HoEL1LW0fLtlcE/YKg7kiIjWo8
q1pBSPELpK2Xgx4lPHtj1iKHNSmm8I1DAHAbmNYxPTJib8ky0jXm97ltvZq7jSG3sG+HxcicQk87
/FxMnqzTvwVyiRJU3E4aZ6jaPhrPCjjCBnR3J/1K8FqEeEOM6aW67BhJytAycuJ6ZbBgzRnBOW6m
UtUZzB5OoowX56VOZBWNudbOPpSEucwuTyzgbqkhYHMi0PFFE9VaZkyKVacAf1jSRmMpcW0nR/XK
TVjLqyF/nagspfk/muGqjG8DdtmwnNOxVqGnzryOJRpxlSa0/uymgorZQF9aVreDgWlOrTVOyePi
LS3iXahGy7ATdM0pHq65msyOyZh+hhm2B5/Tj7CPFdAMnlNoIe2HLLFlhgV7K2IoYFWYrJ91HvfX
zFwLnAYbGuaNqQcaoiNgdY8B6mrb/mdemwVO3ECLd0hUVp3XtzSSM1dn+oSMid+NyHCWNKuF2pI0
sqLqx2yghEMyLSx31OpxJ8KUP6SXvGL8ci97jcz+mu8C35E08XDG0ineXcNS152nWgcovz8eQFBp
zFGSHD51DiiIoC5lqR3AagXEokqz713/eDI+nrLZozX4CvDzrRi8YVrYGkQ/e/YG25isgs1xXgZJ
IOlecXxn0/MaHYKHnPjaHymNkRct319Umv2sGOhdE7wC48cimB/kKcg8FlAzE7ycgISKpSVT/sPf
x+lBrWsUsVZtoEx8i/evylARdHaOhZKiBpR8kBPsx3rjDCCp9aVBzkGz9Gs1ldp0SgwqYU4Fa4i2
2g7kECwopcvS5IU04ZXEGG0s8C6tK/bUYD/l8V9wQpcOwkeP2PLyXtP2qaoYoeBQwICoiFGmal4t
aa7ii3gjJrnt7IvARjoLC9QvznxzRNmRO5JPGb47DbedJ+PY9X4Zybt1te6pNZvmdjptX6rDAhSy
5n05K8+ux7ENsacLml3p7VoHUtF636lUQrje653lPcfqY5j4pu1WaIdF25H7aTFqCOElJNhNKoHE
PQDXynmNPZ44bNZ29QPLRp+oLfvSD4XllgFzXO1bfZJXBT/YBgFxV0d5On6h1yt15ZsQFqhZIYHm
7HrKT/GgeYQ7MY1onRTdnOLrEVY9R3dY0Tr0ji2mE6tfOd6F+Z9XT8iVrhctR0ggIEdeOIQHayCt
MxdZ7NG/cw0Kq+wFoC+Q6LFXDYcmloRmlgXEWuS/Zy5pmZoUQrdAOp25Mul3z0Y71cuW9VwNuas4
7ArBoOlpCSHHAB0OHNrJAkP7HZfzyQHiLxyhiSUSEnV4mldyFQYkuVR8XG4quV6/KEx1SZpjgLFw
Fersrgc81NhQz73+Bnbb67s4CYc1FDYox984uSrt+XiZbpXGEfQ26OiXlwZGabxq5AFIDvr32mqB
emHagqGlW/jMhjpJ08S34IH0yvunscYI6iTpHB9auuvLr1GxtCR3/oa0moBLAgZVn2oagaji7UiZ
YXSN+/q0bI+hyGTa14yeE8MbcXUwnVkwEw1rDL1AOCS3eRhZ0/mUk0SyP1R9CUFQPcJtky5nV8rZ
keVmj2+CMIJBk/CYkrEEa5wg8FhgDrfqNnLYfoJoAUP+vqrwOdk0V3pltXHRe+KfsY+7B9B9Qgf7
tBAlsK3gSlE3u9WR1HqzsdoVFwzq2RPoRFkL0zZZfkpevmtQQw+yC7DYBljWiMPor8qZIdRfvYbM
hJCUePyeC2jxyg0q21F5SY48kPDGsIRtlAoOHJUW+KxKkPC59V4Hwr8cNSTQBcUOryKUrNzxSWF7
vFY2piU8zSNswgdSvqzpQ98D+hABq3lsgOEY2DSn+uKuf2mL9vEZuW7GVtl1SJaoSkgVUTxN11wf
iAyWupmiaebKjJBbc6JtjX9UUn48ZMlPLhQv9OZCK5EettpUnDYcjwX6YkEnL+H7n7dkkSdBQSE9
HxSo+1kXoOVy0EN6Qi5akntXOBpsvSQ5klx4vCfNFDDMYW3LTbHr4WThFh+xdO1Kw9WtB3NDjhU6
7aLi4ef2LI0ibOS8he4DpzuAlO7aXFocdfBFhU0+M9Y2eFpseVldLsrD6oH7Z6FNr6eplzY0hNCa
j9EFeDAZy66htAp/JB0SbAq01E6h+S2Wvoxq1NL4qIfzn5YQxkBwWy4V1KfoC8ZJmQ1AGhYDvZPR
bVjjqj3XKSjgdHJxXAFEaB/MScWSASZP+g+QBnJ/kUoHkF7azHVEQgeVmw9T6NEvEDIm3cH5sNA6
GJzCrWoYkZW0SGf0pFctBZbeTzmK32S9HMiWqRajT6zSMGjXKBl1TPtnyW5QbU5qA1wDl25nACaR
/D240uZjHirC6FxUIwp96L190tKzNpfu6JcxAafTuW2uERF00RRinM3xcrjsd8PabP2pN4g9He6a
JPjKQrOqeVeYwIdqK/oWFG/zJJ8HXhpcxV956NtrWEldO6XY32KYyHGQroc4grikJhdbGCFNgc+Q
azavvGtsuohcBTlnvKw5P1bgaP0XvkyQWzhDuJEskJVc+2leRBgMgM0cWS2mljep6kThdy5ZcaRs
hDG56MGZuaPdwkXP0Y7hH1doZxaweornBgsMZe9Gv6JdDZPIuEFSYb+D0ZQr1AwRoyg12Tjss7Uj
8UELIPVYgC0yP6aMs4zpmL4pCCInT2+BhpBRoQT0avWqK5FhlROgrJHeCXZ7phMOZbHLFi03zEmh
GTyUTEnX9IgN2cperC80zaNUxegktE776til/ghe/faiNPgFq1VC3U8fIBBRF52eJ8IU181D7bam
+38UYiLBwIDqLWDSH5uG9rbRJ3YXlL2UOR4CTBwWeJObmJRJ1c/6KBc1lO9bsS1FUGMBxKtERGqq
hK/f+cP8ySkyegGrGy+oW6k5uHtBJA08qtqVsaLAm2ZZzJdpDX/PfrcGcIVzAiFFFHxSBJTUpTX2
kH2NgC6j/UeI9iNEQ/6ihxmLYQud/2nnsNy6hjavE0ddB4Ie0oz/mKeVRALMnw6/rjCSYawXlIrH
Y4EbKsw0TvmlN2qMb8lFNMIYBD3b+trNSh4G3LHDY+OqyCDxAO6bXBlgZPqHibBakw+ZkpCHlo57
WBYlonMJTmClciNXo6U9nQ1OyuY5GECQ/XuLn4UNW4ngQyXi1hAhX6BUuy3godRo/1+mlXKJUqb/
FYnBkruS14SWS6PgY1MZWhpx3Ihw7J8m3U1AsEcsXkxS+0CRtFYAEGJNCjkkgn0mCPH8+kJwe/G0
sbCi/YRP2PTq0ICWFBOp+KhTyN6uLLPKu0aFxTQ8rdC3mLY3sGAWSf/CJAFPSZFaNVqD7adhTffG
6cy/AiE9XcCRG81X5jzwiL33jxPtm9B2MIbN8TyKEFTQkz+g517Gmxnpu1LdD0V7U997gRkM4IG8
SNmupRMrZfr2PK7jxfXuXIh6INDNnUKRhswxlQnLxJzq1EjRWwadDQtscyMCkhuLwF4nWSNYP/CE
FEh1p57KwgRPDHRkW06muzISWVxjKDO6BKtTcaJ8Yw4oXhyG75rAdskmFUpKkfjiKV4lYtGscUpk
y2smGWibXuYbcTLJj+sx+JiaB7ANHxt8T1whQ5LoQkgNOouQ4Hbaa/7GHkD8pk80oUWOBvTBfyRa
6pcsJ4/vCmixja2KVkbCQn/iwNCqVDZCTyEDHRrvtrZWdH0l/cTpwVvEywE9mYaC4kDqMKnU2qY3
hpSEWoYBQbpY6ixIBFnN+R/Htpjzt92ihZ3dBTPPThaQQ707kQEviEF6nwFMF5CkyQ1B2UjUsotT
3p+nCFTZlfdTqd65sAe6tObgr566m+y51XthZyt9ykfg7NiaD0VAndN/pp/wDbq09Rr7VYPqHSQH
nW1A71OykQGbcgz4ikjtv0mTSfPCnkTSG8pxXigot4n6Jarkdx6j6cemMKSx3o/Wssszz0jlwfGy
A/rSDrJ2ZsDNkwZBWo6DN2v+9Qq0JDCSMZKkXHeIT0ib4Qrhs3YK+kRIgiajlp40zXmxDxjCEWAI
d8IRfy7y2287T1TtEXNUg/FNijmCp6BtU65slJ03UuP9OIg1zmQtDkfiHZo/s5DrWvpkr3dx7K0y
9221dpykxdgwNBk6yDaxfvant6/RxxHB2haAneytFT4/NKlfCwLt9xUbAugSg9g1iKKYy1+IHahZ
MvCq3qqdWcpOrq2rEg3xcE5372E6g9e/fS7lN6ryDejB+RgVWoNCziek+oCvG1IUF+0L2xihNjXr
JFawgt3mwzlX/ALk48GuB/cdM8Nu41mv2HTtPtOIc2uuqkna4NmZnaXYt1N8NVtg6T5qohvx/iNU
bcXPkz75+74pOI9DMWa+cpyO4KuQTcYZHtRYWCmTg+AQIUiyVKKBsrkoM7XdVr6Py3VAnm435yx+
7Xq1kUG3i7jCn6PqRi+gz8dhtW1x31tSZlFJf1lna/PnYa6JIaqtktXubui8yHTPCZJoo3hIaEGe
MBx3wRXC8cIX9+pdbW50lbmxTodYtaIEukOk8sbN0CZ5ZwIMW34ssyGM4+W1ZoawfLtUSXIgivKw
dir8usLQYVCYX1LM/TkbhiCWunLJW2CvydUcbqo+/UC9YZHDQk8C6scW0dTaaP7EuFDqU1P6xgnV
l3N3A0VlbYn1yNKz7klPMzSad+NJW87H3ZgCRSgZa9uhC+sxy5SFQAALQdsj3gEQWf5R4jY75LOn
60Q78cNiQwIGQ+HJ+yzR+7d996yU9ucslwR3u+vvcCt8Q2c6blqMMdPdorIRaLlQO2lahKbT2Xqh
nO4a9OjvI+Exjd1mYEVGhmhpx0xPNqH+j6tnoAzArIiQr3i1TQYdm0Hih5lhvkWG3maCBba5lKyp
Yap8Un+x9Rvz6TILNJyEcAMax5krhdjRiTlV+VXGOGAC8YK/f1uQoGZ+PTo2NQKCvGG1cc033iDI
yOsd4vW25fRaEVbnkI2eAyTdv2XckcbR7KsNuOK+7t9AkF512l4WC2iy6mq2keS6BIgz/aNaAwUB
G+CJCD+jSV7VPLQiS9vO1GDOQPuMObycCWUjYEPbKbnb4wH03lOdVm7OA9Y6LfIa+IuWE4QTAB4I
oxjQ89/c1ax00kXe7Hwosvon9D1jHxXoQQvVV+n8mPkN+uiYk7vaLFoYPx7M18mzDqb2DSPcI1Pk
lYKURkZGhficq+qBc2haiDRGrzMLKZSE/gJJwGKdKHiY/vH+a4TZUWgWY0W7IdUItcINnb4nY21f
NOOEliAwCYXnZA8FkBpkU7KwqUji6ou1G1xGHFMNJswll9KVmIe92GgzfV5rn3k3WiGOnvT86x9Q
V7IKjPOMOZTT+uKwQgtUe9qLtEso/9XGZ3SCRqYkWho25wGU0adenHHTMRt8xMXXDc7Xj6S9wnxT
m/jbdav+VODK/1ZWWpHdgmE+sG59Q058mi/W+uLhXkd9hl7g7N+d6/jsYKrnjfg2bQuspCO4GG0z
Ek7EwWqnav0Mg7QOwqvW9t3Jp6Ecc5jUW8x86jr2s3Ml2+FUs3I4LdOw9nEoEHSaAZWqaCw4tT3g
234mrNeFidyi7xdFoNz6fNtiPiIB5oitdQ8lt4scdUp6rbiU/zoJk/2ckFxP4VtuRLfDljcWtWy0
LZhy0/+aDNw/3mwXmg5e5Yx9KevnOCjdL2ns7rW2WJ4bty8N7ingJxdUL5ujWpAyRe2pbJadaijd
ux4H5QfFivKgla4Fx4efGUZywQkMGgNbk1yvlmAfjlSC/tQD0I/vSQLe0HCON0lWRbt5/FHFPxA5
LdDyBHo4Y7pTp1+P5aRZAkIWauZdpvV2qnDH8NjXGKzlEJV6gCxP1lpb5EA+GxzlpVbb2VhTskxV
1YyiG1oFBsSuSsYhS9fDYLk3fe/VqDvNaT1BwBF7bsJX1mqm5iDwyA/EEiwrKtgotHnl2yejDEo+
Njk/NOMC87i0tnkTVrvzaVcVCrb/Qh9IybT38kbcXvKP8S+4wh6hECgc34DA65PWLR2tzXnIFfMf
4NsF8Xy00gfZEUlNvmkLEz9ruWSdQtO9cA4tuPa3AH6q6+xwa1O9T+a5MoR4ovwcdfuc9P79xhuN
EKiF+Jlrxa1bNz/47CpyT9I9jT1U8Ylnbcxc8tL/02N7JfThr02EfopbJQBA8EJC/s0cItf8kZYY
mc2NZPVLS+kYqvBd17DMbg7JoWKOZ643sTFrr/ANs3HeAlsXIc3mInscLsF1tkvGdY1M7k9sLhqh
8qxQJayU4926nc7VPbW/N4623duw4//gCEOJs3Q9OU6eO5VOiwFDFSM3vCMlm8ec7tsJ4ew2T9tI
78I1DeWXaCMgKbDqigniX+TGWqSoO6PIBwRK8Z4PNbTKhs1wfveuNhjtA5iUDlFQM4Cn/elU6hui
AC9KNCMBKCssUBRSmhdmu0q+UI+Uy3qxmyqkm2cT7eNpQ3sIpK2geEDzk+Dl8FU3itoDuqU8tv+Y
mLpO1Eb8xzGVdw5xDrOeCilcEi1s37syvg5gDPefFNVyaazDZ/CwFrCIKNEyjtJfMnNFvA+WBjyE
vmuNoLuQdE1g+1+kMUg2oQiykfwzCb4WvlZ48WElZ6iOM1CaBKeZudEwwKMy5kJ/gLbNz22fQGy7
rA8XSgquBa97UbLn1z4ieZ1bTjHeiReDWCYU5uGAbxH8sU1EA2Q5MH8bPPVFf3L4xXIosiEmHDSd
jdOPSTDGMu2Nj/pMbctYNWX9vgHPUUVhx4xqHlloamovhsZTNdCsffZITaZ6PeBmI4XF5xpiGnBY
sw9zx9aE+NNte15e/zVU3vNdBbCJsXy6UtPyECMFBXDX0UKyL4fsDjqW+jQy7LxL2HDbeaUSCnpq
aLnR8AhxQE+DFD8H91swpirv+F/StBi80QBsDMS6qrtGPen2fXtaHUn8EKFiNTqFly4Q+mCXQrjA
qr2CtOftIdkf0a8J60NHOZL2paiueCKCAgUfiRJcxkdvL47FQEXRd9iY7q7DYUYL6Qc/6+yyzpjA
3Dv/cVPHr/ZdkozeYcr7TEFl6GvZAc5d2X9SDsPq8xd+0wakVB8Tfns0qYtKozJAFP88U+K/wAjb
1kw7sDxef011e75/cGN1iDkgbYCR2SpQvzTphOsC+XzZRbkuTF0WQ2aktn8tm5OnppnpN5ALwwJW
CtRXA4aR6YKqGd0T7+4UXZA+TUahQlzCF53vRkuFTb4+WGPRwLfCz6yznuQ8sFKdxiVzPFwIFa6x
Y2m2fv8ffqHrqfa0t7RzJahSbuf5+SdC5XdCuvsTfxTjprgFbbbiHe5PFwe5hbpeEX5zERqqKL5q
wkDuokNiZ4YtJR6RpJL2xlD0EXCwhYEKkOleAX/P4gStaNok8kMbKxHzfUoLPJU6lw29B7mbLDMS
zC0sfkP1i5AO2kPm3MDYx4eBvmX7zcJIjeVar8RMUV++uV0X1wqX0v2ZSB1p6s2wdkp3a26aGe2P
Kw7rClMMoFwiol4qUvAFXB2OpkrJOGyxUOLNh9swpKycO8gLuWVjOOSuaLn8+SwO2322PZzfCaEY
bMnMDJ7AATsMAk+b1XooVdnJaEQC4mCMVzli0EVq4t5e+JoQS4KhqBYdalQCVcMbET4otNMNTVdu
+6RhKazXXdnW/3mmZHdYS/n+tMGy/g4w736SI6OR6OPr5WdPuiE/ngxWSfhXATOpaDdk14zwJIvE
CN+4DPNM3eiETe6dnGM3g9/3rHhu0wCyToSJGg21xyEq3XuKcpNuNMxTUCM2MjWVbnTqqktFERgm
ue6rImXsRffz9azJmV5MJsW1oeOVFa3Hda5RDPbVOvAhCU9Krx2k/01Sm78mA3JpS6VAZhD45WWv
9W0FFTqMn64whYYwxQvxMY8vfWPuzXiuTm9cl4TZGlvS83KCKQQTKJSSGGUKyc1bWOHYESzoZQHs
SKLAFSykOHK63/xCjCCSnSNTndDgXVMZGgsLZK3lK3F/5D2Gl5u8C8ExbWMPH4nuESxTwg/drp3+
lMC9pf8j9F5iYkzS/Jm3qk003iwR5XiJvblVaE1Ayfop4mEiUHU8IPoJJX7XDlDR2pDkQjHjiC/f
XQaYleDCXyuV5zMHlEYdvfy80SaLu2uGZqqg9AYxtDTzLh3FYHPp8GPZyAW6TEmzrUUl2EjyhF2E
ejJQDCg7Crmd8Ofg8tl+yRtZ261Y6ycSFiUMRfxRUjxhqlBEjX4uFNBs++hcQOWPWJf+2rvgGPtZ
T+mBrHomwsnfatOhAIuVa9t7ZJjF78Veu319KXw9Aa41ShX0osvdBGzfAx6dP14qQHaDH25ujoGi
RIAVFrLEmRHDRT3POy6kwuwhsd814L6M/ZztVwGfawwZWZ4ZyAm3dbhWRfUnKX5OtwknpKBCvfA2
qnVtUa1uq8To6BSY1c9uEhc+RCO0UE3hCwZ5OZkkXqYrEKZEC+AcuvpoIWjPSU8/y8cFBnDcuaAr
B0/YlmyA1y390FC0D6RGFWmtBl8T0bseeNC/cqcfImaYxlLUBEKRZb4Ubas9cOtJM4iSUPsDz73F
Z2kSKMVg1+4yjFFG4z3m7pO0MIL0UGFDL01f/gptM/J+bceGGydpjtolUIyo5vgedT7A2Td1ieRR
5DVxo7AnVjpGm+Ijg0L4HQjj/7v9aZfyp/no0aCVjaqxR3Qq1LO/rnOeYdvyzFTeiLU8RGsacS+r
3qxefJJqignsl1sOHj3ywW/TcbSAAt4uaNhde7YG2Fw4qMMvBGiBCKxfZc88TJf6Y6LUFbPelRqb
89O13stWStuWlI07rXGTa+yuHRa7zLBxqlq42RZZoSzlbeGW7YiCI+N5Wx3NSonUcLxQ7WF1kbdC
vN0GzeiN8s4h4vnexeCLQGkxBLln3+d1WqpJlU/TBMp/26sirOW9naV8uio8pVwEEbYg89p9YB5J
KnOuuq0MDd0xvNmcQudsDuJ7PLYGP17Lh30RnuzczuDwS0Cot3szVG2EUGkjR/hqme24Iw9fdOWu
fkDvMFwv3vnBPEnAi8h6dpoXUlvnPh0U8Z9JjNkCD9jGJ8un4p/Jb55CPAIeoRQPnhUuWuku0gtg
pNvD7H+ZJFhDx5nj65v9iSmUXUwkOhsNBNOPVeh095Su4aI43MtrKhKspCtgW1uM2OaUh6jFvVLx
+L4o8JX4U6Q2g3tGnX2HdePpKXWjqf6FOIyGDxHuhwlOMVVZ6LzAkvZidf+FJr/mO/hIFyMOJRPj
dtCxS0o5XfOi6/SmsQlLEI/eZe35oFerT9jYCS/VmsFml8Gz81PZ4gWUUVl3WXfzPLsppgM9xTb8
npngXSuRj2B/IT59U/vvLu/zFSuEVbWY/k1u4cwW26eKGaQ1nQfVG91inN/kui69/znUA6GHpcnH
lVOYipC9woXuKVwABXwRdT6Qejq42BpZBRTiNBa7PobciDvaZK1z5SBlhgCREZbf2Xf1+4812wqG
DF+oylyM1xHoxWnkFYJoQ7+G1CH7VmY603Hp5wGRZ9Hfvp2aeEaMGHWW5G2RR751X5EK/DdGgZzt
gB/B+aFXoMWBngFuu9KrRxO73vvnEXkhhusF32Mw9Qv6NBG4dwfDXgZ/T41zH5nUQpCwxEPNTg5l
IuWqZEUMxT08rnpezyP/rPDq4/UTEOku7yxt9WEK3zq1k5V7UKDAWgRI1Fye5EKaacsDn8ZV6M27
MrealiXn/AMTf95kfCGX5z9sBBr4Vi+TnTZs8Pz7W00vZ+INA/E1cr/KG8vQ0gXqEhXi/FDttUAf
/z32zP8uHvb7UPKYH4CbZBKtFLg54HuL/IE3XgZ3hNJoCJlAgTz/nHC5Mx6HYQOgsR4iSitdKqNl
5je8canTu5yU64gBpTiAjhjTCZoCirM2ezQsMkyL65zWOBGaoCA2/s+gDqz8dBzXGmsghWVc2rqw
VR/E7pCushUq1pdcL/QRQGCd5YeyUJBuKiVy/MkKJZkgbnN+HA2WwhqZeLwsM3T5zvnIWY9p+O+O
rMcESBmIWBFz4kdZwT+anoxkmbsqWKCHfnGWpE5+Q3MZ2R01Mzm/2M86pkVWMxzSLxkpI46w0OC9
Jknhomp7qJXdAbLhy6l/vTgANFznYmKwPyrM8HopJIst/8Sdv8sJnF/ICHBAJ5WG0Tpx/+WcG1kS
5Ro2VLDk4sQ2v31uc/6Jm+C72g60Jzg5gASD5592KPIePKvQVEhULuSW/YcH7XD6PHrin54cY8lh
AJPjMh1vNZRYaht3ZyP7XHVuADrEIG4XZNlze9R40yQUZwrGR2PkgBMzbeneJOm/o5xU2QaJbrbU
2WaxG9hjj0BAZy6tll8MJlOq++pKrRxd05oZkcmMkBKLeKgI9mqGUaKhNyRxufxufsqDy0ZBMwBo
Vt74QaORSpb3P/GXHbr6K8jcsvwqCIRZrVBNk/bzIK6boDNaapDLqCiK6NNo24wP/C3+l4cwtsZc
2dmSBlYxt1QD4y+r0geUf9jp5iQvf2nTwmZtN60jNE4sHlka6D5aWtM0yNPFPbPVfY7/Ypi7wyop
6/JT1FFGND41MkbmyRbN+0wm6Acx8ezC1+g7/X6Gis6My3kuy9avLk9TZBx8tWwP9puax6DvhSZZ
1lLjq4L7OVs8668at7Yvcst53jyd4L2Ut/REP1195bL33qurBKAbLnR7tDgrn1ara5+zi9tAsGI9
ZIDcJZu4ay7Ha4Z3dZIp9YFT0xLGUeHjkPdEYc6dkaTlvwEFpVJez+YCw5f/t94CFJ+AnExtF33j
Mgo4qVn4AxQ9RqLtvCfAk1n8/VPpT0DHAk0xrWGHSyrRpipQe/paCToINUsoFFkbnvhmgqzqdO/9
9SN8U3Pqcou5XOzXPtAaiJm5kWnI/aFlJiG4HrNu8yKCT4Zxlc65GNci7OgXrC+lzyryrX9EbYnt
uFbXnmuo4ll5pH5AuXkDx8BwrES+HUAI7kg/79xygQyPkUHN3Ar1x1WWPCDP5iplZX8vdd8ka7xE
Em+DdO1ZicQwJSpWSz3NgXT/qtYr9/JMLUwLk0gi6L9Ho30Baw00Kqhvx+3uBJYOYy5NlBdMvkMW
Lg8cXdCz6VG2IHHvlmVzMHL/g+1lCu9VZFD7kfPh6Qgv92ZeKGxYpkLmqdluS4e5YCCfFW3OGu/A
pC2Lw1+bVI/ajC0gILOylIGPwisYQhD+nBk2W8bFnv4K4tefCB1ZTzeAEOxYlGhazWVtiCosss7p
DzWSbhqNnsm/o68BsFGwbr1wfxfrlRmLX9Oaaj1LnkLfhCfej9qd5HjvF2T4rAcTDn5kkvho6FWk
7wqrMrkIyU6ndHKzufd9qzgqrmRarbzcnuz3/Cl9ea7b6unftgjzLITa3+IkU1PPJQp3zDEdWrdU
dXj7QoEHyPM876HgfcuiWxd74GqVhRpErcay5oA1OkLa7P3RYPAFBUE5RFXaJ2+YPILVt0JmMH55
FSBLSvzru5OLJqhFUHRnmlZT4mil/qFwdcOUgY0KuRB0/5IXtbWLX0N06BTfXwybLog6VLo+jKa2
qxaOOLdZZ1EPHP5zElwOffPSmVPtHMQfyF/aaQCCu/HolxZVI/dsRFhoFhs0iub7LlbU/su75ObM
VT9wuDI51iWWWeAXajqU+VB4llU6B5eluq1QmypKX9G7qH35pFUgUAluQ5zXwcpnNNJJMMNsyRwV
IzD+3cmgaEyUFSjEYsv9mdiMDJ4zZ3KW13GLGKvLC5JMJjvVWRQb36zP4x3baGOaRzp0jniuCPdt
Nbjm7IAGHEbthQcTE0maCL0zq/q8BHQifdO4ZZNBrmd4SycckW6bfgKoc78JWXFrYoEiT326FOr8
2PIZv+WFu2cIhRp5tokInGjOKrRZLpcrqFwPaGVCry14qYEOziSg6hof0eHte0XrMDppm2XyzBFQ
uRMejLTTA2JeHl1EAt0kNHWkryZywucvTxqUnu9Ubcl9N7Le2OC7V9c55EaChOWYeXloq6tgQA5D
nUVNl/P7FMfyR8ZJnIPDy2aX3FSPDzTrzki35Y8LL7CEvbyVai3lg6dHhu6dEoejWpS7ipdjzeWo
LO/invIPyGH8tI5YJnxI4gClDqim1CaeEcsfoueJcwwa7tEi2OLySWU1Y2vPbImbuJh4X/Iwk9fi
hWgNE3Wjbic/q6d7ezCAm0Eek5iAVwAwRATI8TCsCxldfecs9Sq5MslS2N/0BQTJgzuyPxTnbc7B
dCTqrU881tlWc6OtEQIDn+yAtsEYlPx0H2Kmp+R8um5PRR7HKElPbd/ccgl/pfnwG/GXix2LodVa
imICT1CqG3yKRrrgC+uWclcg1B4MrCWs8kpxKsSZDps5XZZecnijGDE8AxZw2AzCs3Y9PmXOnKZb
NpJIJYT1ZlLVZnZvwg47PIl9/yqupgrMoaIqfEUM0hX03aZFhuBYnT1SB5zYwyrKVRf8wYPM6Ten
5GTTDaxbyY+Wbx8DNSuYoz7ogojraWrCOwa9PjhoEnBXSY5wYFarImCuKEbvfWKI48gf7OYVlGdT
1aXrriRrEoAk9ljGax/tIrRbchSEfm17LNaqaZxCz7TzEpDHvG8juklaCi7AxyZHUyTQAzjPRCnv
nqKhsfqkjcEfuhKKiDEfkkrYzpdgFJ2b8SzuZcodJO1nOzG7c03AOaULJngZkA7hemA7cDzpd92k
viyKYXQOKHqQybqWV6gka2pI+5PKATXpHSH8NPjrwOzGVuM6BtpZZfqe/pyKP9Yqn0gQehJ6pTyJ
mveHXus9kvm4JWGaVSZjan0wuNz58NxuFo1axfP4twHCv/52FKDxYEnuGqgDgYhXbv1+PLVVbmk5
qyv8Qc2MUGvFLOmbBusOQY/Tjc+7oMsQ33KvymmDT/o9dYtoOKpJlnPhm6atQjPCBFOWPtKfm5Y/
tVtLLWfK8U9320JKpS2asiPZNogNLNMvuQc61Dy0QOzTsPA8iRkyt0m0c6+f3Crjnj+gbf+fyeY9
eFilNi8Tv2kpv6dkACQvRf00ZUMRMUSlBu9q9Jr9n4ibo1agPucFEHg+raYowvHe1HHQAle1cSS+
Y9S4Rx0OJe9+RTb//+AfgRpAE4UIpmy+xRf3cHwXT5R449Cr0dJduSI+Cea2ZsNI/s0qWVtbHycb
Wd6A8B7yI3nRUyLDfGZ5ECwb8FlSd2SfWVEcFjoLcf9G2cVOD2Imtbzw2gookCVGL1Xwwq+kdt1z
P2FpxUT8xd48OU8yYMoof65NEKcwgzws9W2pmYAk4voKfM4LpyCNZdfNueXK6inhexHpJq1ivNsL
qp5eOibHQJP8ni8aJo3d1Yk47501hGoPShhrQimAFDXaPTkKRT+faJ+HUi2IUebUJIoeFVnNKPZC
Y17dv85rcZfyrjFQGgVQr/XErFl4s6Lx9QhzIaAgUMpyvEB8Pkou5cb6aKvpYX/2RRk3IYEMmV8g
UMuts4Q/t07+gQtSKoS4epvbrhFK6VBxrsIwhVPnck/dotWJtVVODno8vi7VB0IVtMeTYbIpFIoA
hoRjCZ6GdCHI4HdXJ6SN8T//+vA/IsDJhEBwDvSuCvnH5juFgiWnCK3lMLrdV784EDS+PwghgMEn
I/a9fb5YOGLbWAtLdlRB7zzjbWVQC1Hk7n9eH7m1JOhzizEMCLgPbuDHoCSI3eL30CftZFoG797y
JJOz9CkrAYSzDKDvgeHkpYgXxJrq9uLxobya2lQtexid+vFAiFYOUJTMyJhFBX3SNHypNBjCu8JQ
vtNlL4TalCXD9HRU8JCalkW4Y41VG0pK/FNs5VtjzU8Gu5fFPDnCEEmS2o59JDoqbHUJV8aWbRvg
qZEY48GbMt3hrqgJbxEmok5z8avUDiXnyJNrBwJcdpq9o+9zADRX6ycF5KJ7HFUpQW1lGy9kQzJf
d9sGSQo5OzHg5sex4gwBzrMxutqv4LQWCPAM8/QvNzisLAxaRNbGzWxZEzFwK9nIIEHQLKbWEHw3
SbJuO41Th8WnahJQUYD/30PHQqRbwOttNVVP451WInn1Eb1qOEqZnjDbyqk6llNn9CC+D1IoJb3j
cKdOy7lydED4oEQ00s2FXQ/6qmaCVx+4ZRd3NmZVxwyrZfWPBL+zz3uaL72v0DVhfiOusMQoCRfu
aTD2sQ3I0GQ2G33XxN8QF2EKSUrMk18cGVIGeBWJwd1pSNhbAFhdyeOGhZUuuPojUIDM364s8D56
+OsaipE06wAnojUIvfc9QZDdEhr/gtggwnAZW8lWDNoNfPH8Ojg8skmCU0U1AdtN6Uo4LlaJEKtW
GCae6oPSv1gYUHD1Dqobl7nAa44265k15C6V9KVg0uUywW7gbHiVhPTJoJWl4tN+EIs1jLCU32vn
O0/72zKlhPIh1pqsoEca2YW0r4PoGPl3kgwQNQ+MbPQn+H9PXMUZ+F2sExBcLWTapFazlNkJZOwA
N51OEpazMfs3f+tKl0uts0sHY4icw2sqoeHpbnr2BG2C+ia/jcvEkBhEAVA75r6T8jCVNaEHci1y
rsSDcCLoNJS5HP/lloudALOH5TehigX3PLTd/OVQJDgZg5iYJTIf6oIqRb05Xj3OikyuQT4f5ONI
at+1FGjNRY5Lrs9zYKw3mtTfLN3A9OCpWmmzVbuxXEzaAL7NezuF/0Dv0c0LIWrz4Lkuk9GNw3kB
qXuUXrqUwGkjhj431tDmdfarEr5U9jTZDQPGGGGAbazc+lC97poL4fPLn/4APPVLSU9069awTXwQ
dPrUcKW3nSirBGQV/yKotn1Wzmo/BwYT6iun4TJGiPzJ9Mrm68V7lFbkyvAxYmdh+AWN53AGfMxK
3iTk7XLNDRWCrD2sXVVgpJZYnyvE5KA4Ln3kuQqQSK6iwFsxRLjG1zcFiPxj+6i1o9Q/jbC0VR59
r1301UTX2jwpg+W1/RDYXx65wZCF0OP70dDpJyukDg2AtlkeNHaRR6WVS3Kn8m9hB6Qxg1Hb+VY1
byWcgR0ZSs+L95fuGd/KD8QXd/WdCzWtntAf2VWj72743FHZuhq/6YFcW+ac9Z87PtTS1qBW1r4P
j4bia8Rrd0tAnuBOXaqTlS+PcWUevvw1HlULHYESFZ6dWFMX9DwltZXK6um4a51U3fJOX884SdH3
fmGIROAYLpDoqkZSkX5GRpnXO6IkYK+sc2f2adgQaEipl3p5UT4Siv7mNzodS/vkPMUGgGiFa5G3
/Tsd0uRII0dKPmJQSP/cE/zscp6QMjJ2OatUlCRyv1exZmK2wZ1a8h2dqQhXXrPzsq4Py4dEaLvh
L8ivI3r91gNQTzNB/ofZs02ThJmy47G7Rz00Q2BsYdhy2jglM8l354fPuib3sb7vw0vR+5EU6mYh
cxe6PQ1Nfc6XL2eCYwCYMcdLxKNqgniM/Py9igNgM9QueB/5Wq4/q8IClvl/7VK7cDq4ONuT94Rm
fqTfA7alN8wRVw2hwvURdCj09V3b2CX/7wMJraO7GEMPNNIxGfRo/O3WTxWkL7Rzl+X5m4FsVDBq
D0KPv3Gqsf+j8LHXyHBlyhdrxHcrPqkSZZZfm8vAVqiIzTIhOGVIlTT7qnlVW26QOtlzCEMuEpX2
X8wiXT2bF6ZG/s74CpvXVK/h6asi+cdGr3HXafhlryjUFaMvCTakz1pkAqD4G0Ia6OlF1gV9HI6n
d7uAMxsinkXLRBLnHNbqEEpTdK3+sfpMXG5A0qUFyp3AdtKleufm36wBYdfA6WFH5vpO0brQqA4R
oKqVFSx4G4cfezhJy/UF7sMJtq0BpIv8n9vHBt1vTX3vkSIfos9SbrCnxFZz2Zj0oN8klXLd36v+
FvjpdAq9pV7SeZK+kBBqzaIvhVZ9ql4V2enPiB1+AN+asEVuBq7MMm+f/LkmACwgFVwRd2VtAZXx
Bim/ZE+E4QbQ9rvbHciJSb8MpyRDuvFajr/7q4oBTBAzP4db11Luoh6zHHtXlHHQ/P88kmhPTCPV
TV+R+pG7hRujm63pQY8d4VOro29/00ZfTFC5JjYWTarNgPZOVtIUwET6oa/n6yWwlWXQdabETfki
pxfSzDN30Wtsk9iZZkG142IlSCtsLjgkTl/LIwhisXljon6Mi8p0Z00QJVrPi7GIeZsCgzhAmuPt
w/ozJprZkFTb26ZIQXYQDaDq61snKuYhNyqWeCQ6kz98tgg5djj7Ikk++T/gDedXClbs8WW6O4eq
auoQRhfyT4XRxRKP6IbMqjklEEbG+S+gQYlg/cYA/t6lDNw/m2vhAfJ1F+pvn+ErUpH5mrOrRAGX
XMNp+DfdBKbEJ+6XVjIHtlcxaI5NqzgoZLNpO87SgyT9oAq6IsTXTp2GYg4MobSwode6rOVEsDa3
MMjUARTJQuXHMJaOQF8Lgnggp71fNsSF+5d4skf3MWDBorutpPNDw0DqVdHH8AUHSi5hjUC8J02r
vXpttC+6yazS+vsYW0DufuPhcYE/n5t0rr90+vhwvZaObuEhC6VUXGxjEoM2b/Q1SGtWPD6csw/g
CINSxxljA/OGXOMC3f7q2CoRvFxACvHgsYt2kuLM1/LZf+2Gnc1pjpf5n1lJcov5ANZET+R0pgXN
hpZ3uixPYKAlRG9eLSKPZPsNwesMrbdGffHiV23bQMncXrDExLvgd00QXfUhPq8yj9vXH1vAVy/2
qY2H30m1UAGp2ahvDnVDY8Kri4ryxHoSmMNU2fBYcOlFNV4a+UozfHYaJR7eTVynWx66xLcVS/NR
xBz0bO7mJwU0a0e6KJZH/x6VPr2letFzGhrHWf0rm2/P777Cr1Q5Jf5O7GYIA9Q5sieWgBW+UzHd
tb0wZthCUGfBm/NS+SFnEEl7gbzUVCvlx2SrRzMP+gewNQo134LgR0ONQumex42nEQVulY/Lzwp1
1SAT90Kg0C5UNJeWQgg5HdihctN42ewR/QNK4ILjinfvMvF6qvuYvStYHf28PS8/zeAsHtcHNvYS
CiWeP8HYWucuFS4GJ4Rq8K4oIWP7dPpP+H6izxymZ/jI+cJfncaqlNDtgzKFk5jSXp3GIJ2Gyte7
MThDme7HwOClScDPjOPBMsdG67/2K8WXOGibbOkYFx2wsEIbHSMcZOj/GRSBrRzR37WjzpUEJpdt
eCWPynvgZM1DuwqBJsv1UY1ZpD/3VS/AJX76tbohEDDZiYuByJ5/ZptE5CxhDsWdKgBkmBF2d81N
d+DoCwWK73ZRkq9wm/L4YPyQjmCoQhpLrSM8yEDuf1U9R2XACQdmXGfrFKNeS3hlcqLKVE/QQrnO
BqDxlKcALs2qx/Zwlkou/lUli/Rc/2d9NWNNBdMNlp17/OFdcTrGh6j9b8FxB3XMWnzlBI3uwzMs
3fSxxiRtF6R0yIXFtzN8kZY0blTmT63jCnUL+pkTG6+ll8vxLSPkTgputpPRe33pDAkcZMdRHVWR
d0QVkZ7au0Gx776qEZyXzQz0s4tSc5xOPgAbMLd5om8encgHVEsXR1L3aNCH7wQ4sCpG6j9GSKPN
DBiAI+0zE3hdAHyBjJ7BhIpkxBkvhbi3NVJypgO8FmwUKL9M0XYnhLCDqdyocmr194qWl5yJ7aoY
jDXONMJXl2dwj8Nq4tTci8ArenGFW9jDhjQgtUw6nsYGMdo28Cdl1jIX7M6iF6pac9/rhWyTLFms
c/z1eyIAXDbLAxOSv+JXv1v3YC+zD2lwQ+j4C3AiIrbd048EtkvSj4+HAEZMZ93W/TMzD0RW1cmd
Ari/Bo2fEjQE4l6OX+Z/sXAEhrf1Nrm48krIt1mS+g9ikHxRdjizualowSMzo8BqNViYUeQ7rr6W
QB0DsNucPJW9NTHgIMIlMCMy1MHxlqjdpOVCXbBwlbJlRiM4i3zpbKkk8me0rkMOWG1p4YKTLc6l
HY3CXyqbe6XELU2VW827ZLOGqY5P6mF+UPfc0Eb4UPDaO8m5C+0dRHFlfUYSJSnCdJ6wwc2QtISn
SsHgkNyHURNIeHzntifV389WmTlNojyfNKR9JV4Ro/w6GGQmbp9YiMt5dxTKY8ltr2NDE9fOngPR
OUpAk+Z8mqIJAIotZe/VxgeVUqs4OjKU3LMKBkdMwkT6u+DtPgINVY59MGJsYCK8WraliGi3sQNX
rD487JqVZwrVbVk+bKoO2n81Rl5QjKDMQjqeBkri0kaqv0ytt7ssz9lsD7O3vdHwlfgEzUXNQmFb
QVvYv0kTkivbjgvNjLNCVCmWOJhylVf8CHaDGLC4tyoHZxrgHrraVsxz4phhHCDXKW9H8+Ait0pl
ipASGueGwbTKcHJbuPuzKmTqUqB36qp0zkNK6rhM3fYgJSyosodrmMQUeD3KFMa2kufEF3sSjZ2u
U/eFIqYkItt0aDxm/TdxdXLh0TJxhkKtxGwBXAZUYP/mkgIL7MIsqTaYDN8666MFQh0nMlDROO06
MkfHL8SO3Vmv3WrREAjhWWQ7nd62sOXSkuBsBQJJlZGI7sxLfrBCPXrZdH7Wd3OVNMZ17hgFLTuH
BRADMgC+kVslF4yTHB+QcwIVB8KDpciD17DzA2T8tcg0EJkdMxilA83nxIc2Ige0kOqLmRqY5TPz
XUHjKiJKABDwEjKwK6wsqFsr/arTz/7qIH1sE54hfUy0nKmOC0wj21/1oKJ6UyhxLYElMeoHwRhW
FQm+Ubzu3qHbk+w3E5ODKQ3PYusvA9MBSicyC8r2bwnUrdiFTy9+D/YWvOcOAi6+SQ9Xp/Og7M7g
USaz6vQX469Z8PPs4r+1YE7YwiFWjIocAPWireIWwiqmmVtDz/ovxKcjY2x9ay4zyBbZD3FWmKdE
CioD/GBrm2Tw1x9C19VnZ3Mr3lWes4Sqor1JErSe8aItkxQCmIehI4YPSQW/uU9ivrzKCGXPHxOy
YIB8J+362z1vw9w5sS9kVmwYcivrZ8+fWBBuE+YhnUuKSTDvGwN9Ni/SixS5EXAPdTaqaUcE8exq
Blt9f7xi/jSaRie/aMP8jShjyFvv1jbu3kQjzVO2scPflShKFR4+5ZoBkbUBeWCFAp6XQ4kOpCff
z2iab7cTnpdMRu+t3I1SQ6rJnEjWNQsWY7KBOvV4JLvRp7XN+e2msex5nEn99EIcafCgmkWdFNRi
p93ARGAUHyusr333fWjxawXyRTbmGdj5/wVoRmhjNw3ZFNgpMhA4Z+a/qgtOk7eExEX4Q9YrTsqm
TjdUEvFz3E5nLF0kbnJ28Jv6QPYTJ34eec2sy+KQobs0kMWrpLPnO0wSdUK7/G4GoaTnNp/z0TIh
kebt4LUNOpAFlT37z3QH50lONmXVn8l8zUIYvybWe+1wztqurACxZg6ErwBwfULx2FBlTm9JIXa1
oMpUVOfLqg21SfKnFB+cNCqbmoCrzf+jBjrPK4cKy69piOR1nZbqzxSpCZRVhaDvqf8IgEKrArPq
5SBOoSd04tkRQXMWhKXQowtNrCW/rWYC8myeFDczD5Pi4l2tJB3zjeL/lt4O0iDdoByEvz8roeU7
dQndtfr7KCAVsbP52UzxuS8XNpdEWtMGbeg8xTKfbcH0yMpsM8zsLgzEQ6lZsQnW+TrP6i6TOKfu
jJNCYQTkWOlK0JDrQs9XBNapmUL1i8FXvUNEcnm39JOxKwrH04b6M/OpdhA+IJelVTorMmqY5RC2
XbTEKUvqVzrRJ0OBY9lbmpofkeqsoD0GmyawT87unqIE5fCr4yHPRBHZIUJds7LQ3R9TQHdQ1nNg
HA5eiycLtkeTHFMt22v+bKr9RwoPCaJVbHWSQimEGsJ5VE+TitSY98UX4WpzK7+xLmzoHfdvFyKX
zqy90Tcdg5s83rOzRsyKssqdESKwo5Su2p2FhFHZ9nhPCdUt5Vr2cELOSiaMDNOlz9Q+WXERZ7sG
MTOreYG9+8Sovgl9YPe5Z8E1cJwKbqCJU7wkGrnbnORVS36KU4tcpY5kUOSryuVYdmInVuZQMHvI
RgGGRWlN2hm6E+2grkALtMDUOTZW6gN/jpQk2n9gpq1E9F3rcOifPrp/lhrhbNP647ZtlDl5mOLf
No2JPFcSb0L/psyuZoFW8ZIjTvh0KEMM1kScVn2t3wHFMzIAKod5jeIoizKaPUu4HR6PhYSXd8xl
SVVF6lAvGVJr9/ElNoRhsRj2ehq/7ItSgA4oFMYqvdkvs72ONwoKU9hiPKzs7pQw8MogDO3FFU8H
cdrK/4iCXYPN9X17fv/DugLf89FyQODIrqjcd3BJpr8mJ/qkiuZN2g+pznBhtg6CRufny5tWvDiv
BWQW688EZ2LfqEc/heSifblbno8cG4+UONHXyvSzOYb/IRBl041TrOLyd/WSDoIyIeSpmG6kAK6a
g8AeA11qDCKaQkj6+SJlkhBHeHz1AYNjx6quPyX6mvxph5otxeVEYra4/Fv4Fo8NWHWCwWDmFEKA
hew5NkAhndHOki/DsW9BX2xXLArzQ5EXVWMDkrXAXZkqinDYZfvfITgxtdJulQjyUbg4NcCQT1Gu
fWWhRsPn9U6vnR+u2mOkT2jVbwuJ+sTiNnnOp5NbXjQPzTGiO6mHelq6LQpncGuzvCNdfaaIp2n9
XrC9sMfh4veD3dR3V23y+xH4rRoYXSuSwh82VUBJezHiu4lRAZONCVU3MrO6zxpVhckJ+nTT86WE
WGIjmQOY2Pkqu622kkrQMGmz9RreNnDbGrEC93gthWG+UGC2EmmE70c9Ln9GY05soy5wDuhpRXT+
BZVhh98VMu1/BGArlUyD/IyGQ3Yh4btDHbPjlQt7HBrmBnCsGohOf9pKDE3n51tIGwKYj2U5HHc5
p6iyYfi+0/VWApqh2Fd8Aqdk/73vxY9l8UwHp9jr2i0r2DN2o99cjQ9Z30BExHT8M3aVHLdPLg2g
jemfZAgxFjH5A0qlsnd7OPicIxMrMEYz7cExXPc1pEDdUc+a8kHdqXsYp6BSdtIsIiq28ddYmGtp
CANdj5w28c5qCTrJiSKUvVWYETnT0KnTYK9UH4prE5eXkwTJ3+dVIc9gmWpDC0hXG2fQyKkiRhYI
AZLooScJAB92uthwhMENiwp7P7mXpD0g8RpY382c2pq1A9TkSCzSqDVh8nvaTj5OXVHh5RAJuaqZ
J7cjduiPJh4tQN4GihPIj9tNUKit0p/a4rjXKcybTrk+um3TVb5GGa1Ko571w4/Bq7Q2N2lnoIrr
D7BTyTFUU/tOLiRBjgiMwCEH8oc+whSvN+Tyoubt4ziXENDQcsbgw3pE12IpJhb9XsIOUbpr3k/e
ic/67VSqS7sgCU2fC/hqt9XxoWUKHbE+ulkst9UTSn1Qx71NTp4M+no0riDAvll5FI9cEcGOPhoG
uec5i407UYA/Ijfwj+gtPTgHx7TGwSivkOH8V7VA4iBcueCuk4sq6RUo6cDvEgoDecA/nO/HsPf8
g19YAltdQ7t9L/ZgPAOp6nUc1UfWrrp28yh9XtH+qBI6v6CLZwY9ctj9FbDUcvW/63LEdEdy+Uuc
QdDuho7kclhVdQRCfcIkKeZ/6q71Du+roMAt0GSsmChwXxbpd7EWPaq+KkOt3AQcpan9BF5zBl7y
9TmQl1Ae3wUXN5CBaNMP2mfzQ2VB7qWovUb+rdCtmpOdriw83aZ356C+huivYW+zkeGGpouwAMRm
LgmSPLAq+8GsdbrrlrUeN3UnanjwqB4mMp2Iuwnq/FbljOrO3Iar2rqAPbguZL7yHQIY7109vVyf
GHnlgj2gw1/U//G5JbQtCWG+4GVaut3NsEOSk2sk/+FJr672/tmD2aHVNb7sZqnV9TK0J8eX4OCx
xV0eNe43YH3wkMZe1NswSDAUPeQYAX1LA5v5nEdRMD5iq4oDpF3jlV/7qYp99DZrrMMc3RDo7YfM
WaEmFXGq0cPNJ52kLOEu0L6viBQ/TT4tLXwGDUsksCO5hxFsfNmU0ZfQgCGd/6trM9WOTyx+NYFV
Ckpj1Z86D8Nia2HKU92wzXvIPu4TYWF8B8zyyKKKMt2dvSJLUdnVmeGqUzdGOyrUQBrNn9aW8bqY
TS/I/kpN7kzPzWT7Q6i6qj1OOz1KzeMHRSGBQ4LwLZKPD/ps96Zb2uKPkHJ7QQQE8xGPv1B6r2uY
Oj2QrxWOSOrZj4MDhvIt1qYrXDPuvIF+pJLEUFab9bUsniHxFxQIdlQ3kVg+4Ya+pgjijv19gzCf
oMl3YbR/wcmt7H0TwMqIjl0UseEl+y6Ilqpdcf9ydV6OiOla2y3aczPky5BRDnkCe4V5Thamg4/8
GbwHmO7R79FHoVN5BcejaFXtHwHYSygWPqtiItkPFNMzSBVbL8cpH6wJYz50V7hRcI+Agtrrzg8/
y1WzcqAniBJa08ZB4BTvRqRevlUvBD2R2Luh+qv+mmT+CZqu/smUCPNlyKFcRPNjs2FaIzV6DvwI
cS1KjR9zrQEyh9G4Dpt568Q4/NSopH9rsyRytAniCqwY1odM2EQBMHk0CKrLd/Kz8RXKqg7+hTy9
wXY3gcxXXu9p0acRJf36AboO0bwgJwyvSpm2ApCyQxuOO6O5UHIU+acPRkl1XQb/Dyyfm0wFoxhb
KBsAxeJ1M6f/g7eFpcxAMfZMjhihsFBfkoPlUw8iQkR/VzOj/mBNkVVdGH4MmYlcDbIJkcXqgnb/
rNMKUZmOEXeKnjCwj9CKgZarINYduoEy2xKV9C9Eao+4TzsJ48T8Zsk/sZmLJQc+MMJ0yxrAZ+PX
9yanrFmwLd4jpgl261EvbIZj8pOFzZP5gnDFcmypVKIq/+Z7bbgaGLPI988iTtqkypgmypXZSNKj
FuCOCWLleaoLj0zCo7hHHg9tULPQj4AcvTkqnoZ9XxHdkXgJvyzejttwAXlx0qwztkLf4L4cfiw1
QI06f/WgMuVup79t2zi78gxUBPwncNF5PZjPUSPTabk3F0Mka/ZpAt7wQl25Z4yQRj931eYz24Z7
7aQPowdMyzFLeiRFg2X28+Myoyt/47Zo/Cx2n8+4ZKlNQe88IwBz43gUquOqMtyhnZKtw1g/ixup
sp+M3QdnbjCo6edT1zxon/C77bAQ6idybUvpkRpCGsFfjPtjzFnkWFR0K6/Vx9PdpDUX/V0OS3Wk
f3zLSQ54boyKovCT1fGd4TZ77S63FO9qUR+i/PfgCLU9X8oDFrC98Sh9mgRy2a49VKSHKfuogTCH
9d5qHRvc+e3XG+yyi/3/iMkoL7+4vQFh6ItnOCUsg+SkXI1iAd3+wLbWGlcc/ukeCj/Zs9+SjAXx
drM8SIWgPzAxEdSccVjb0ewaQcXETJvZ0q8Gs2tIB08QkMY0a9lZkjFUicX0T21n/uj9p5P+5OA+
FU1d06I9DRT1Xas/WoL3SfgcsN/gwieOyzWUUfV3yJGDTIcdyqDovovoMs6mnQInm7iazi72Wnz7
ieCZ4pJ2EKCdqtnJAe1VADj/0LsMmkHo4UdvS5bRG9LUC5mgRJcsGxfT+iVPDQ19cMpslWBSjVjI
iSRdtpfML59Loj7jQWfUSneAVWm7RyiR2bwF5wcmJlFURVLD+0c6qE4RVKFipI2FCkVHxEsm2X2c
8qHYDMSksC4OQKLz2cr319azBsE8/M9XNl0BoGMJHzXdca8Sl9FqFdXwwmfw7BSTvyetUvdXwV+g
Mm9Vs0L6mGVWfjDF4it+uJ6ZT23B0j5tpgqwUH7AvPLVnIAwJwfgYjeOY001i5ZEKF6F0YciUok7
6X6arcHvnx7otHknwk9axChPWQ9pHGVdK9KMOpCpj3VrLfug0WXjuuWJNcBcjcKlocqTEKXjb7JM
4lMxLRuBLizevlmvx+ngjMORrWhGGGX7eOnnueJIkIhY175ta5rvdN/g9w+zeMl7GrtBVtI8fW1q
BFDZ+wnHgYozBtHrw5eSRojyXJu0DJPOxvsAM+6/A6TkNSGsa6TDnbKtT89GKsYlIF/jJWnO5WCS
8pjqATGyzJnRl0WooU/oba3aSHcDtftVS55UWvy7CkVmGC2sN9W+0LhBoRpzY6qee8SfakDhi9cw
seSrUWtKQLwnI5ujHVLZGdNiHId41xMm6knUpkHQyO4xdcgyhU7AI5FBLs3NTKmv3TvJ0r6O3S/2
whC87GC55h2wSIpY3STB3PcCkL5ZzHbfCJU5tyPZ5TWOxl0AxDQ9xgfzHErk5D6LUR9fVCqOpZec
k3IxxCpb0kT/sL0t5JvCFtMv0PSltDAweOEq3bwS/sDHYBXsLQ8up9UKYOMPj60TLv9A1tpTxC3D
HewbgUttqgkMLDqn7nGpLfW/ulfew8CssKNmuD9Mg0Md5NSigPU46V89dDOpwflPrC/NLlKhNXOT
CVxziAHE447vmNKhuWTMKXken+ojyPLBjBEn+6tH0jhvA3XJc6uqvADiADmyzv3/2lI71vg0P9W1
3c9m+W4Opy4xM3jtdev9BiFtoRQq2KUQkFf25MvP3pbdedA6xuH9geO17Jb0B6t9Z8vT1xdgf/wu
WcdaDQTPTcQ0QikvZUj4Bbyq4q333OJJH3eOcvmnJ8CJP6uoJWz86OgwbL17vf7Fi4U6otCVnAqR
1KBGpiEoYoDiVcQ5pZZMPgtrkrItIlrGHk3t72Pi5s7pkXSLKOjOMf9q+tyn+Oivaf4jdYmtLUW1
bbSbywfZ+1jyKsXlq9f45LXwoT/s3pE6L9zu6ZN8s7EOQFFJt423fUl5J4scMiDoGcVZQLILV6nq
Tq0myzJ6MzPw0gUAXxLSqpzQO9oBDUGq/dcjdQIYra7jf2xVaouwRLjzUO7TSsS7gCdjrUyr1fUd
rB8Qzn9aFadVMaD9VNsYkfvvKMokL+LemsdegIia85lrfdu5c244vjXaq/t8StH5Df2j0JtttDi9
6opoWvsRH+qst1QYpXxinB2q04kTGXZ7kzJq+YfojqhfcxEBxsz1OEZOTVKhmw2n9TCfhinmL7z0
MuzofwFvlHAKsd+LPADSgfB0fcKDzi6vThdqrF3/Xw7alW8tWfUtO67PlYds8HnoM5tTpgnxUKqW
ozG+cSzzc1I5HippdocoT+/xR+Et91MUSagv6JM2fc+1hId+X/K675uFr5DR4mrQbNjRAH8VTb9h
oRJ9c4/ksQ7fcTOGqFrpr55rgdWulgAMvDxGTd4BzsDvB9mU2V+nftTGe+evvy2shpeJ3QA9JNVZ
cR0+apIB0iO3lPRJACclRSc0RZAJRYUUIirBZijCeE/Wjr7SKmtdY6vpxCYkB52o1ZJq+Mk7+Rt7
7Vmw4wprlAdW/Z0RQHaigf5oqtq+rDpdRP3p7Sij5W4Uufv89shAaDnAY5d9Ig33PuPKFS8v09Id
GSHfBM17SzGaSKTMYgWBBttPwA9pvJHApoDzVP7K9mKCgzEGU5FSvuu6XsX81OotipYqeOzjgzzw
g9RLodUVRZ2vwhvhS4JHP35YDtb2DfjwLVwba8M17O0dwzsx0jm9cnFPdlWcx6ArRXA7PeY7Uy5Y
MHuthTYnE3cK/thT6vjk7192+TtwpTrl0MEthoi6IGSj3+qOG1CdmE6cbdMc1nG0kZ5jEEKFo4fj
TJn28GZthPukYsnlK4jeW5oBDIqTavzNiFcY2HI+K4GRlmTsKKDW8T3kyFMd6wP8TI4oiDFR5AwQ
z73I/rfk8qATojyUnsJ6cAJGiWeASb+9eVyPMy30kAWwECESTE7vQI0lZkKQaU+NpeeZNPtGjhuY
v2pxpzJ7LuN11MN06D6ZE+h1YudGcFZJNtl6uArTbopLdKwoQN5BlIvjbGJI2FBpOFxLtPEiIqkE
tdOkBGY+hQi6FVEzWb6+M/fkxj+lw604BFfcTMtFok/qqjlzyqklFjitGQqkEyd/DPwiNWCPspKa
lMTrT1L9KuFgmkndulnWycSL2BChttrfg4aSFIJ1X7i9kFj9GrWzvTijRvvNNOwMiAW5nABG1Grp
AspkW8bs6auOHi+eP0/+i8an/J+igRqXT1Sm08K10+5L3Lf8SmwhvzUzjc80InVGp7TaoFtAPpI0
1vP6ZeDwru+hcPSQ7YgGOWKDh2NRBxOkRiE76MNlniv11RZlgQz+btyH8qWRyxd2eaBEsO7PbJ6G
VZK7pOIXtftB9qA8xWDBOitPI7b43iqwH3+aMTSRsIzby1ShanXGjMfALS/s8/ehJ3Kzhmq0kzkS
5oOV3BMwgIi82BMeiWW8X83BmQNHlIcOmVZpiuLeXBloMTdw2mnsdFF7iRgs6q9f41tCDFJVHABe
f5VgalkHXGbgFnXRFjFfg+g3Mux1W4qfnMv+qRabSJ5m0tlxEcObDleHUNQSllo9cRrTeC0kFKnu
EWIq/jlOt4Vb3mGbohIBGgIXZoDGUxdccxdmhe7k9sCQVLOVta0i9Qe/7M6MO9qKwNJ9t1btSstI
WliOTAJgsk5SKL2PfhMYuWj5yhVZ0KiEkFfBs/R08JwjTpbxVb+yRdnzkEuS5dy7OPvVBCBmpusQ
rTVk7fKjQIdN5eXkyJV8yh6pBTyx+IlhRMRt+rx0WTCK6FYpfw8DnT2YNsZP4y9Su7vQ6ClQTZnP
SDJxphX6UjihLEgieT2QtdN8i7MI4vNZgcnWFrhsQiSlR0BLlESkwsYbTtaQ6Nlu3mDEqDIWO+1F
ha7/4VbE4Z0l7sVj4o9Jjodsmtr8sz31XqUgdxa5SK0emwMAnxfrV5bQKFQhrNNICH2iKws5ABVF
q6KKMmktjWvG6iFtZ1lDjDjXuAufH3WuHYtEGUac750xkcnsGwNz21e0fXgCeTO9CMjnpjXm6qp5
ZxYCbxDFD4BXid8PgpEdSc29Sn8jZI/mtitmsvmtieSvJn017FfdEELDxNW60EiRMrjMEd90WXEm
HS+wxn/onqURwCryWyGTUQuoM1US2qQfEK1pwlhM7UrjBYrWCrEjloid2c4cUe/lHcGXSBloALta
XUsf2b+/YnjbmmTiSmhv7gDmFkOiiC1djj4OjYmwWmYpOcu4kirs65zFb4n5XvdwUwq22AJQcMwf
8go44aXWG5dTnF4zgEjSDuVcuCr6yxN/6hQ9p8pnYlGMSKsfGCSB+vKB2xDXIVSfs3bs08x2uVAv
qWKmclgC4ZUX7yfYbWEKqkKXBlFki6yJ54SVPW6iEzULYTgE8PjDMT3rtu/itWKai3JLwQKxjI8V
m/0g6wynlpCUKLbED8cD4UCU9ix+IcOJfb75+rRRRP4qpiNXcqUd2hvw83Obo8zJz6e5knS73vBh
iFcqm7K/AkQs6OjDJC/zdyKz80DALcDiRzJxebe13b19jMKzU1cJUojwR4EPWcjTijsYT/THM1XU
FkRB1uG6yM3ryPddxkgdu+wWidlwdDZETR7+0CnkS5hY5tXNijzcW63R8jeN4d7tf/hOqYo78cIz
f2WOVYUN0CvhbKrijJDClAQBcdXPXxWgDwUe85Ctyb7uZI2WZ2ojEMSkGKq2WNpHMWk8sObOi78/
WJX4paDnTX5Hf7gNgnphFuoOhonQhQa8Q7sUNJ577g0hKCccip/R2HZe4AOc9Rt7HxxkGO0+39LV
EUyHaoasygsiAuJ9/OijCQWzywm0qmZLn34qeH2afj6XLSN2wtMuV0dAgW1chvtyHmQEPe2K/NqW
OWqpskl37PzBOyYPS8ddC7OatY+UgNm77XAlSP0/yldJrM3elyrTFrDdZsQUkTDRBQaUmvWK52fd
pjE1hE45wxLu70RkoKAe3LLMCtPKHJvKvx4qc1WrUWO82PzLc9mn3wFqVeX/Ui2tJqJ3+TgeVTWJ
R3n7KGBC1+UiteFbn41cu7vRGb8udnhBr2KH98sSk9tjCR3LtdlQwU7Vn9olo1lmoTPUSOiUO6gU
wOahohPZFCxIPUyfhHJing4NVSAHe/6J3vH9FS8YNoOr7sFMgYFdqkOFqQL1Qy2/I/zRi1GAD5Rw
jBo/n+S7HsV9tltZI39jpvKQbuldSkF/FUFCUnidvweInlaYdP4o3TAuRKpfc4gkSeNAeDCzw4Us
hWZociVnnQ7xswG9RTzh3/B+JD8E21KJgxrEexlkYU5HBo/03w1Lr3GDeq61lsex8ORtPt1eAoa1
j2vRD2Glf/ZU5DilCOb/kRZNgpmTWQdQzWWG11RtOCXi/+lerqA3jIrc/KgB1gd1Fu8ToO7m+Pzk
jGabAwHAj7tGesWBfS0NDJrx9tgfjdITkCeHVe25+fFJEW4kwzFHcJ9KzHxPUkrTlsGpX8nd+8q/
o5249KveJKMRixeQPuqWdFjuVQgx0TNHa0Hn/dOd1PuthLJGuPm6qUROp4EUca/wojF7ILQYPtRz
RP8D1+hYrnTtURx5+EKtaKwXzj0fAkv+Tl+DdIaDETq4anVLGjk3PRIuzNhuc5KKo3sJwNjxiEvR
YuUVBtuNJwswlW8YAxSOw0jMpQeqO5UulnG/s/9KV1lawUcgukfLCMyo+TRGW+B+MEuJmbV3YaX9
OUucYj7dg4IizEpld5/4E2Lou/hHkGpl4khG7xOIyMZe9jwjitVMMpafNXGn6JJMyh/1uP5/nAHO
EzF1zDpXg9HxmMlXlX5MTfKcrfw+7B9uXF5zOroyDaKOq6ROHmJWbBX0958eqIszK8yatFJW5FBP
UhDthPvMMvd+EBb4QgWv7mRQtmKwEufddEjsa2B8gQQkXhG5jd8ZhHO8hkdjbdgY09v2SA3DEQ/W
OzlhTXH5uDPdd9NdH9/2VIW2HPO1VSKsmEixomkMfjbmYPAoT8TgTAiAXoNfgeuabvgm6Lsb2TVl
T37HJSyI9zEa9ii2pWwkAbvFg6S6pt1DCkrZiNiTe/RHTi3/+k9RI66pHjGu3kwpRQxKSDDHWGQA
JJd76Ia/eqv7HljFjPhrLIfIuZmzFkqIP8SSqS53n6cVbm1f5G5aIQqaXIR6oCFi4p7FtQH8Zniv
wUCkJh0EbjtfvEvU5fM2VUwxERsN/eWMiI2WxMhoT4eFGd/M7rKg4vLFswIOQ12wBgSfaqjCT5Yt
ox6ZjhUoLg6XKTro5dsQDIaaWp2KpfCVffuE4P1fbinzefS2ycHsNAcGGzkEZBR6URFI79I1TZbR
Ekn2F/3Rh/6P9OUl4HC2JhOQxGOM61bO0bxbB8I0osqzsuL4YfYQe3M9vHWtsBW3U2GqnQEeh4rD
Kglss4qtVwK4x3Yb7EXZ7a1wuUecLrvalf9hkk0lD3SDBd8mpMRA1iohQDRiBKPBGcLKIONZN515
SmNhkbJWyJPk9IEd47COGVT/8g2vKgoUDv3DKrTYioyYPpv4STJyaHiKKRzabhYj1eBUypCqEg6q
4xcbkc6OdiI9PFINtEKJIfvpBGcuHWnSbteGaLTBa61y8mWUKXCL++VUbrF0apVcrOZS7z46HwU8
btsi5Ydq+LdQtWYkFyxThBMNMSPjQLVgto7e9OSW9UiiMoIH8Yh0PVIRu2qplxC88GG247zXng4K
ZokaaKCa8ZtPlH/bcyLmoWJanFprucfkE100U44ARdMB7GGLsAuFVOLL5MZF6L7yDSdDt5cq5xmR
r1LnV+qUMjGlN0XbwuItLYPyFTP75FKvKyenicaaNQXyKP/S3C035LNhkEXfZ8/ECJD3OILaBQ3f
Jh0O1IFK1aagosVZgKM3Jzk50VIoU2GRAa40847tBUL9NeyoCLbVZTYKUX3M0Xk2sf/71HL94g0t
PX0kk/vjN4coeZH/ccii0aJY/yaFvkIbwDJlHKEDrJmU8b5g6OBtvrPZfAsRCEn5hpYYF/s08Ea2
rRqSPBGYVZj3BSF5ApZ+oHwLP4argqeFcpQoOkNCfh3S+gi8Ntumj/7U7SLMoCgS+WLGYoGSisB/
803kK/FhfNC/SoinQz6TWrLP3cdBE8zmVooPUS+6h+8jjDEdBp1FjFpCs8cGbUBJ2851g/iHAB73
gj619oKVNceza5KDesRepfRKsfBY2foQpvYYQ6Idn6bLS/MffCfaQBiqGMQqEoYm9oyTYPgQ2a7r
YDtX01Cok0N/mW6SsVRt2ujrqnAHE3/DaszaOjQCPy6b0aMdb2fb9P2vhFv/WgjpDu1Va2rhwehb
FDzXFAI82nIv9J3qebMBsb5+jlMl+YcRtzmkOSlhPJmPhlhbkmkLQemIcvf6JX9RvZoJ26NSStBv
aizEe3sCCmH8BVoUU15UlY2vXRwjjZ9bp8pxYkmu1CpIRSXHfzR0N94eDMKbCOoyNim+//fEVTiO
+4FPJB7yrn1OEFvl4cqOWBlW+ub+ZVGmtp4dtiDWZujfwmGARFs8AcgrpYNctn8bzQ6VC/sv4Q1o
JMyy+Ftc1F0gnBYYGKNGiXCvy8XHenPO/xLrUnYnKB8ZCZYXvpRSQHJ8gMArhtVsoa0PI8mnRSvG
5N7DAAyVukepdKCeFBya/0dh6Yt1EuOnrsqHtBABFcuTrusMIPan7/1wdkwToIp6KgJbr76uc9+x
4TXnQFoJOjdptWtrR6Rd0m0Vuc/rAvVgBJkTGNk0p8CCSU6BBMeRpKEkVjGCyOfOmtPscdVH5DbY
vsQ38bLpAm7XvlYqSXrrsWLTJekf9SzYol/bMCvGBagpozUfyulq+cA2yI2SMNe0ds8EzkJ6ul9I
xrKhqOjHxyM7GURzB7IaT3tfK5HSlYZ5cxEkskrZ7PC9jfGs0WiBGia7ES7IqwzDhMfuIw2iA10k
TtpZ7rQG5I4QEh1m5BZ/pbTNpuQnhI3XpFbOU9EUi2OuA2TZcRoxJyE9y8wRVW5N9tzj9sHyy4RJ
zxL1V/B/4rek5IVe0UYRpq9EAZlddU31J0kTLWQyO1qoFtMTxpHi1vqp5fC3ne6vMtOlmNHdzGEI
DI/XFpH/ybPwLaGGadh75li8z9fYBDZKquKyal5uXq2M0Y/O9gw1FaNgZ3n7mJJkWqXor3aJi8PP
siDCmEvvY4B22G2U7Wsz1G2tOPjtopXA5VKRFKg7lws0TzWsXyZ5nx3xNNXyomX69BaQNUc9dXFC
S7EiQ3tGdE2TUT8YnG7+0crCqGyRrmOPVgJLxvdN5VQ3MBQPKG/0kLF03KDJp6rASY74WEPvYb9X
yGmCGUvHMykz+/dJqmV5sXcnDLuNbX87Nx4WAg/HKSr2ROt6d9u5NrAoX8J6mpdUCggusKEqO7e5
COTHiXmiT/2Q7Ks87ldVSk2FBSv+kyzwg4r4C4dUOCmM80cmNkz99FOIq79vx1vw8vcG6V3to9gH
GpUQym/skN6ukPOgoNRZnxrwL8XYW4Nk1JAGKiu74YxXb214r4BPY1jAWjTFECdLujLDeWsSL4sF
lkb98ZhdHz0J2YCatEAknoU7VYXvWoA1aNjVPmFak5lv1ijdRBkjQbknhorcJdeUIg3NSlAEBB6u
ElZDVGJG3CqVvgInWqMOWGk68EiYUURmVoMwLdH5t8JE7qd6kzOC2IRRfPEdTZAor+MY9nJx0oPq
82YmkV6z3GqsoIMeGLU7RUj5IS4t8cwVyB1B13dPEyyZ/h/pzCgzdF70/6X3T8r4I8HB4tMP49Wl
gmsLpzmTM4GFFqYwz7myVOq5RQS6ARHM1WUrIBFcigAsux0MdhsBXqEQ9LOWusGEXHAS/2gIlKIx
gy14XUHuqUM0SwBTVdbgnL1cD5Mv4Oc++mLp6HYX8jb77W5S0Vy7briT7rr/ZoHx6LXnL9r8QLkn
A+HagSq8id0GNvhVN1MumWig824LZitGrcg7z9lt8+IFldLcbW+7aon9T7+7iluMsgCtJwH0yk90
509qI68+A5gjnzwlwqwT5CWqHegiabXo0ihZJi6fNVuecDJIunwO5CXP2D0nE0kNftCg+XJYoPRL
roKU8w5GtOfq2SKq0g4BMW0rKjmjp7XgXp8HexW7ATilQyyuHLYHxv/kQyF1WyYeMz8miI2e4xqU
CkABCC+p4KhFsFosyF+WMM5qzcyMvWWQVA9hW1N/66UnmMm2YJbW/2V/bugpFB45S1rvzD+B+T+U
r61wzhXhAzFtiLD+qi8+s1GEjo8zFBzRO0AuIGb5Lj2fPPpBggIP1Tgo7ySwFi1/GxHOHNWq/iP8
lFDCtzzsyBY48cUnns2Kcx5yjADIWF6Tq/GbtDxIcUFAyr6I784QUku6vQJLe4bXRt6Xs1OqfVsg
qGazOEeNQ4SoFUCi7c21cKb4+4EGeIXVw9MEVy+QIBq9ckI38kg7nrrV6hPQsVF/NV10Pdmi9WGt
AusdRO+NamE3Y+Hp0nwWDiAgSGxCHgxpjxeAegzzuSHuesKCSIdphIhMkvKkBaER88JXhRr7BsQx
Jz+EbQi1VL1porEixfUZZFZmP5K0wntp4rESA68sv8vNo0tVLgdRj5rG+IwdjftihubqKKhGJJKn
CphLCauUDhjijznQBv+KRTSNnODDv7Lqwh0mIjlpfTOWnBSbDnMdYUX6tM/TzogPzhEFGOdXyj/A
EKblluEBbxu5A1fI8GdIb+ZR0FYAhxpURnzJemEsWmP2EewpQlhSfoNDsbvCtmbUkAlW82qCo/1D
g+SQfWEYB1IJ6amPFEFyJozpuKAXmwkvhiVmdMGOVwCMId6mv+CNXrJuL16IUspI0CCmkNSzGB3o
FT5CD8/DOHBKer86cGq8k4dgzjLGHhSxtmJsae4qkRAnuWC+gn1pd5XVvv3FiJvCgz/sxB4BrNfz
vifRrAKdKQdowoZkRMKHnHX8jylb9iLF7na6wZ/LtH70EVrz0gAuWfn5r8dtMSDuI0jT3JWO66lm
IR/L1Em0TlpbhgBAvYGN+fGd13vd3CIG+5H6EZando9hoVCVLH2uLvdanpINP/SOMVSYAntRPcPJ
tSlvhbTe+HEqFSo8Lk8AVzcQMrSZSYLG0N5Lp9TYQxki6GwMh5CiVRSmJWl4bXVQsPSJNNdQZqDw
qF5Y18ixUdSsabK+uYWVx3d5zQPSZegJffcaDjo9cYYSs7xPVSD7ciyFpt6n/seqqBmP9JmivDTW
mjxRRF/aaN94joBwiiv2EYYNieqJRZEkqCU6I1AJq7c/IdlQFUgkZ1HYifIS1NB1R1JPSVCoCymL
N17aGyznyJ3Q565ZOJviW7SDpq2delwoWL5scvoYABGJaxL7AuNe/QYEucTCZj8OrdpKhaeVJdke
GT1HPGWe0WmaLvVy8A3/dpzlzx1+H+xIDV2PO+G0TIEYQtOJ/Y0XibuIPZDYOszPJPdncX5d2eTw
fmThab455gOM3w7DoTEIj7jS6z9mXwqq79/Y3RHdzMu9cwIUi+Q65O7AdIZgDFzXDHlPH4/nZiJb
C1FPA3PaVgWdypljeYnpJiVulcX3dQV3c1VYm+vqoYIhTWvpN8vuY+yo+W9X+zwHTCQW64IooTH3
Nsz33TPA8OcNQug+JlSuQ6ckVX0kTY1q/wu+wDXRwQsCW5MqXa3iqtykIB/WlblCDKJJz08pauWk
S6g9w5HqXJxfjCLnCfziMn8s9Kcbv1UF/v6Fd06T2Y+Lx3GJMPXY3fmJF8EttTHGKPJdgNZC5T80
t6VjJZtMVfK+oVqqhm6OeWcvFjCUAC0bRz9d0lpoK6ejZ0u7B4NOUGlrEoBcNpLUluNG/VfJK29c
NlgcP/SzR9WINHoSqGq5WB+I4sHE7FArtFNTOsb1pFxwdnlvAWS5Ctmy3oBeOCi78Ns+PBkOvlLC
562WDxyzqIXsiW3qQk4/joUiXBqNQXPhG8MK6yObYkFaomV5KHZMPhMmYFW1R7I02pf6ShY1BEQy
RFxj+qQQDg1suz6KwSa+uIVMX9rUeuGEe9fMwEKoc3JZWfrj1F7WGn+wuWOOJyeh74lW5OSxJBO4
CpZ6UljmgOWpQAh0ZinzTyvXc0f1GIt9HIPDwhQyZhc1wtfoDinNoICcCyde8cHXd0RWiM3gycZY
G4QQc0s6c/wlEHf38LEUUIcVjkCnwxdF62STuaTzSQYfIrjPkrxBSYnda9O8mw/gqC4rYqAdDQCG
n8JCViw2l/pfkWBCllS0TrVHFDOOT3X0f+MmhCZOlz97sjZd8st8XZc9IzlzmptW/8bvBb8LPC+o
SQEM/xCLRvZdPpgqY/U6pCYL3RqkhrwmAwoBOUTgtcYm3jh23ye4lwDVNq25OTifYPvLf75YGuyN
kCWpzUkt/1YgIhTEa/Y37lgt4cJXb79rp8jkdWNVMAyjW8BmahwW5oaqd4NXeGRBCPVqZ0QqHvYU
YVaOATIkBKYpC/IEhqO0hRGCOFbUVOqo3fdcHS/ZU+GqxmDRYuuAT1XXyLKK89/jaJCzRBS6+TdX
s4r320p+emPqYmabuYWAx2xuGkUaK1jve1F/FIOrHVtrEH9eXI2Fa0+n7C0Ki1mNmpom1RL8Q+TJ
gKOaeewbcgsLs2WW5VmTe0rhZVqNzEz9Jb7nHtHTx029yGxo1ueVEXQ8Y7GyhBhHl7+NpYOMQ2if
m1OKhfmy0XKLVAEux34looG545kCi7szIDSm/qR+v//d/Bk6tvsVUa56gF4a7CaYHYRJIxV3cf1w
Ub3EPGiFtzBY8oyoQhmAmWnVTUr/k1SsOjB45EqlOK3u6I2Q2hKPjWFUDq5s6aIS7aRm3O6kXGVR
xc+jqmTSgl8E84q5K+Fad/mdSe4rpG8ZVySLsjpYsOq6w9OD4KG10/bYXP8LLR+lrLOok1mmTJtx
HrLiVVHWQIuQ5kZWX5kDX3Ss+1Dhztb024kEL0AoToxgqB4htOPwMYmkgr6h+gVj0ZAXm48Qm5Kl
c7iySSvgZuPzSU8xVNt4jL5Bis1Nu6b3mri2ZfJE8ZK6A5uhkKWbZC6rQLoCwZeA5xFCdWq/Mln0
QBwQ7PGMiFjKjDYA5cqicDP7K1/c/XO6f9MxA0qLeI7dTUKskl/VNjeM84S/LeHgWPnbbB3OGb87
zhSaekoMJFCwR1/UIcnWT1ss9IvZsDYWXZaDqax6w4f9EKUTS1sfwCEVEajWwdEz4OZzWfCZnLk6
HE0lh7rktaPCD0uVGW73FTCPt4regK8r+tnWJ0lYF7nMnGzW73nE7rWp+HT8Qk6hWT2ArNvzeIro
05gd/eE5LPn+pz+5gQXAwLy/phuXsVw5ua2v/ij9Uor650FvTW2SSwczD5BiTnpvSfWktp4LZGTH
Dp5EqdQdJMDv7xP7trlrk8p7RZ2JX8+gXUjT3eRHJ3+P1OcsNmU93k+QChu7+jotqKDf4XNIIip3
OKqYt8CM44TAKJDoFissNjGNmQfZgYhfkXe/Cqv9d28SRmFeJfigcexo5bOK6WrcFSuwDpHGdHrK
/xcRF9VNGsgx5qJShJYP8oGr+aA/mX5NW4xVG2WDk+fkDTMPAfvMUktLY1PdMoUTkkujIx0VN2Uu
uLuZHLt8Xp8rbFClvmGxGj08+jhO33Hmumxf8Tf5qKhylqzdB7EylLm/9dyH+o6uMZMZGt1sr0U0
aS6YeT+IBpGxmMOIo9PgQ7ltxZS304bwnPWMAiX0cud51TFGD0xoj4HzLh4Y3YH7fDUoenyC1Ag+
bjrUHsIM9ljxbukRsc303wZUO541+fBBeHj8ovqthVkTvw4DxvyhVDt/QDjogYdaDcFhsU/nENTK
rWwP0+88uD5qhyA9+5hql2+aFftE6vZjYG5QLlrE9slfWo11dmfqR8wgCP7Siu00BewEu8qyUqAI
socwlZSoCH9lAx+MTlbsKvEyUMYNqdHrRM3EMyUA5KPdZ7RGnmau5Emb3xeSpTi8b046+bBNH9B8
H3lmU2VbPtdJT0kGFH/MMPeusiW6Y2IcfqtR4ZhYjFDZoXkUlYRwOYg57FV8I49RzcWsadqI4tJt
gSw28RkGDPIKT9uSqdub1vWAsqVTNov6wwCW9QwCJDcXU5QVHy2Vgu/NbGGlu2sUEKxDMp+0hBho
Z9e2862+JjtQtqhad1E/aK3eQ4cLjrNJjLJn2i/F6Xm7+67DM5lw87tH0oV7vF06M8mlS7uaKrTf
D66FKK3thTW0n+kNC3clwIjIvjsOe3VT6nvLUQ0eL+IXMHY4NdVcEDm3ZdRma0L20kVLDmHBf1tX
GWGASS9pbe6VppuRW3r9fgJt07bXN8ORvIPSARcCGsYFfylbzykz6EFt29e0oGyvtfW/E+PSM4Hm
ji9YmX/yANiWeOqcTBQ2PJpHO2GWRt2v0kE1mCYsbrRCDtXAcm2i0OfK8MjHV+DmdxhdUq7NuB3m
Zxfh7owOV1NrW+HppwVUsOmd7zojlHI8L7wu7R6Spi31T28gvAcj0AmDZ0z+x5h4+6ef0fn6X/Tj
ly9ak15/su7frptMMARMnV78IPKKW253Xm0uE/ow3l1R8E2iX3jgiGirido75ptPM15mPtRD6pE+
rPJH+suRGY21ezh3IC/Q37nAcF4UxT0YUcymFLvBXf9XYdfqnCgn+mzu7P1x/9Oqqo+gMe4hkbA5
2WbTpBqipRW5mGAc0vofdJ8cbVDPphymDf1a1mXorU78gR5hRo/QcxN33+pG4ssetVqYONGEL1JT
1I3zesjqJFpvDDmJmHX6DLa4VF45mR175WtNNMD4FX42W4cRlSgrSaxl76HrwYmqnncSH/xp2rI4
LTF+SdNzQUZDa6V7+y6WQh9Q9HGD6bRmBYdE38FIPKg3Vn7bQa/+IQIgcGOMTMjZTGdQy2bTWLXi
eghT1DZOLeEBBYl6wQWjYpxmd5nTVEO6jsqJbzNToiaaX8IoHGCLBHmpQW2GioLP2S46If3OVm11
7gzA5nZzZpTXhowtT3kVGKLrtI22Dj72fO742/toTu0cARBV4QBMyS43bcagTDN1DFSmDVLOggz9
gTme7RuJD+2eBDgpPTKnVzuDnSOyk6DWp8sHtOibQ5lOL2G7xCwVStSGemrgn60pAOmd9H1QUk6Q
Wqf7+bsn+s6/SIMxPMSoQh66BQ0CdTq/AwJopmIjGaIJ89mI9PmBiw/fR00RC8vkTcMx0IBq9Dmx
KHJuxWXKdit/LKlEmvm7jHvBgXtGBNri6tMajjid4vaAD2KKtBucmbpQYpR7Q+3dDS5WBjhNzieO
2dZo1B2seRCzItm2CxEVSJR4OcuN2MtIDJnglLATteTjoAauTf+rA31pF+3F2y8ViW6IkonXwFCJ
Rt5wfXKfq/IsNpwnbbQvfKbNMU4B0xnNUva+KGDPtF3EQpvVn7TsbCW1FcA0dNdqSRJHf8IHmxZz
JTbA59vCCAW6v+ZhPQRR3TFoMaYm7J6Z49oKOwxXIi9jhyv5Cde+5McSfWMXaJgyGTpucu8JTOUW
1KrzrAI6Y34Ep0e4Z83C/5LrOCWS/fr94kUiDaKbz9ad4anqU7rT3IWOwsJb5Ud0WaquyC20xgWJ
g321YLl4QrxCxFM8SthPVVw/dwdFDzWuE85YzYLoNyTmnIugErAYJGN8KB7xMDYiabkzLR8Jlf3y
vpadT22QjVXhUmxjwGYWo/MhtbjXJF78B9ilKLT7f3YwNMDsFzDRYdrFuXcjGp61knmFTjrIluex
0slIJQJu2rdnLbFrKvDaZZb3RUqwV1LKWYOSDED9gqyJEgVdv6qgWm+syiCeZz5AwQCODiYuU/22
qxrjlp0erXT6XAejjF93+1D+XVo+MRyYEHe4hO1lONc5qROPH0g4uOJxx8u3+FeNjt3tCUVP0z5d
CKS8j1VFRN4fw/fvY/EeSHIJO7SfEABGlJwjxiah6M5XmZ3PhKXw0P3Isyw9wEfQT39V53QYaPLa
8mWTk48qPCIwOSNEqUeY5c1eZWlefCMXiIsqn7YPDXTZBDIH1MNjw0zALPsyL356W/yJzys+MTET
3F3GK3ORS+JsW+bXDrfCxQ/BK10w1Uue9RLTNUbDv0zzsYYVWY3zPNuo+8ep7CAFFKm09+rEHrXH
H3cALW9GjV3kZEmQxcaYx3V8KGKb+c7mpwDNOxZZhL7fUqhBJw5gsQ7s4cjR7rm7nj9AqDoo2Qvz
QQ2O2BIoOSe6lcnvZopFcrYoc6EqpRRIzkvOWajTlZ3e7bIGI1BcmxoHP9/nfSDGcVdGv0rJVIcn
0eJcxhIC2aFgpufJInpS20NEMpor4XmsK49pADzO0BsfjDEc36YMkRAYFxA5gw89GrRPUR+DRi68
UpwRa6o1i68cgyL8cPo2iXMGeOIzDRJdjFU5G5mhjyqKkQfJ0urzpRkMAVRgA7hxWtX9a22QNIXQ
eMI7xF2ZTGVqNdYSL6gQXHh8Uk3kM4ie11qK5SNasqm0QeZR1JRzNYCFFx40UjbbTtmX6w7H6hfW
12GjQQDJUtp10CRCk3PdqXhNAk3sgSoGNBYO5xG+aK8RLlJHEv8ERax57uY7SwyI9FMOKXBAxmTJ
7B33rylitD93vzek7eKE9LfBxwiDw5uGxEkwGnJcdWkR8Mjf+yNDVwteFBh0plaoDvjNKPZvexEo
6qr2+N2Lc6FhupmghhFXnjs03Wj4ESJyEv1tgH3+vof5tJksevYyqcwvx0PWLeok+wDwfJ0c0qR3
tqxUUcM6qI6MZ0vlgP6ipqLgumMxn1up6UsSu1HtnrGpYbVcNYs0iIhGpWCv05jhBYZSfBwFE3a7
SFmd8Cvozo7DYxHbhz/D0rafqLC56vpg4Hn/JU/ZortDYCyRE4E95fRyIEYJlRqxTfVZBD8M7ykz
Sc9xF2jm3u+Yfwu3+j/nX/2vjIWQgtK01UOs28bU4j1IL/hOUrF3THf5d2qahvVnGfuBoTOmXV1p
aHRQUt13T/2mUvMsg8HWW2b69EDN8jFUKNmJNH1YYg0uuKL1X6cSes/oj9znW+oMLjeXjUimw02b
2E0QZLQ5UTXz8Rimv08CzSlyKFkVzIPswhwmLNtvA3WpbVXrFKyz8qy0Pi1pu4a2OpnEPFM5bMnR
8mEW5XoJRV9lJ4iRXM+ACNckWF+iXCVWCaBkdUT4nbWMrxptH0dCeAH/djCJsnVVU6Z2muk4WYwI
9pFzCZRfquwQEcCt3YJKdixBtS/VkkDjeM41ZaD6QPeyNLqjfWvJ5cWNWYApH1U+TZJ1OlZt5qYS
vst6gs/BkvOy44j2yV+sp0WjPDjXgR7EpsYRthk8xKgrfns5cGnGrCmcYlZn03v5tMSOJ4ENocl3
s1U7O0w3FFfigqcYRkrwD6NxPAOPgJFpn6vz4ZCYczcNC8hCt2GuRPxWIJVLYKJz2kCnNrv7ow2E
1uPBH5bKyzxK4OnJxfuz6jjDRWX3SfjsfJfTKMgG5vZXRr2EwcpT7eo+gk8kPmrCgVm2FdGXQuKP
K+Zx2YKu75K+UHlXfzsTmRSUCn/flwOtHqehZcxnrM4I9iXDUWR7GJk7khwmJkO/JvSLYebhom6T
RTNstHbSJngpnCX8oHAwp9K1tnQX/a4S6bVrkWhzaEu4Bc/6zHTTcJrblY5lfAvitxoOecYWcG5O
7UX/RtoqdCDcXk92fE09o3j1056688TDUZ6QD7Ms2w7MbXtNK2nfpeXtFL9Xy0E4Y9oIw6XEFSzg
BRWxyqJNVAnxOtztUMjPyhOuwxctQaKpZW5RyJzVMZXWuBhX6V9RhmColNTEh6M5+TIGIyrDJ9iP
hrz9lsXacV/39Q/McohmHei/XeXFgK2EmkHRM0hwCDu3L1MWQoxCCh+A9lncPPKxq7+fRxcK9MOq
6SzbBvccvANHZZb6yVjRfrXPo+0ytQnvJt0kQqmYOPHX5z8chO1wqcogf16K97kq+VKMTeoHqgFS
Ajk+0GXrVHg0V/wC96l7vlpAA4e+Q25AP27dx7XAKrPjE+YGmrje5e9pmPxbewRRIefoXxa5ptbh
TDRmOQNa7H3M1ULkPmO5WI/jT9Hj7tbq2f5qtb502rkI8DoM+sGYHV4dBK2b0x28zHkUD14wbpI/
S2pcmSn4MxPyC0PDBnlxUFQ5Fje7AA5rNfr2zpuZ3/IZXOU7RgX6dW9ExBAn/cH9HoM1BE3JPZkt
TFsjbngnB/OvqkzxpiuBOIUoKcPVpL6scteRID7W0Srn1v1OCZyXPS+tOy97gLtB7ldf6jgkMjiu
JbfsPWZplIGiiIbiQeZPhwR925xSpZcLfzyc0ESw6qtZqlGQTHh/scu5mpwGF8X0C+W2DpNwlMvw
DjTJmXCcaljPTpr/VWmnUjYbsHYeOVw2EIWLvTxiiZfoiwTx2FGUxLH2HZ9ad/d1s+6lMM1gtvLf
d+FE1JgPto+3I5GyJG//s10XxvRmlt7kBAUZlVMpyXo5OaaVUn4qbKUGo98bHIDTwJFi2JCG/f44
rkm3XTO0ccUHjt+dzXY03ujpdHbW2Z5tQjfnRNCaQlgN25/aC8vMu0YdlCPPeTbaodt5mHk3xLJZ
c3SiWkTyjHDHfWFeHxO60MfPz3TI9o4RtHEpYh95YNM9oPJ4U6hYhIvso7Qpt5ABG0/yPs7mGIm0
mEKluzsIdTljoSbJYp5S/k6YIQ3S8WFAAKlZL66AKtjgrIu4zwFr2NcvzkuJ0h/BWUGNn12p3XLE
GphmZpxgRYN08XTI9bkLCljB59hNMEOYxDTRPgtREIAQXUu4iGIkw0pIcEowBF+nqmJL2HKhByfo
8iYCNCG4gazxj3o/R2tJK2hZ35fNyc667J6uLjTeTk2K7wsai8Bk7bP0WbFWb02s58oUtao0ehxR
VON6dwMMnW4IiYT/ku1Y5TdGhzkZO9uhDKl6JbKQAxabQ2/bFe7DPfZOlvumKuiMC+IUwTA2DqJI
wr74qmqN9PKT9zHtJirMsJlujLFL+z9HrU/CcwZi6FCyRA/InCIuwhkU6rKWqTwOcVDkWFyGu4NA
gW8o72f+4g2Oe+U8uOMpF6rrBuMNaxK2y8TkAYCf387NrcA/36BoT/S+mwPb8g8PZFy7yfRtxPvT
HKioaM6/qa96av2hOJA7HwhvTN+P9YzURjdpo1Tk0C84TV3JD3wXwSQEPH4QLp9TBuKiiL+MdhT4
UoKGD6wdfa4LIcqphcXsEp3X7WJ/L6PMwzkeIEknDEUhiZFbm4eqhdWaQrVG38YRL8S+nohrbkiL
uIr4Y4+HHL0zWWjhoiho1ag1fAsE8Ld0invr20mZeNkqjmDHNpGIgaXr+R8lA79OEuR0U367hp2X
p3MXQPotk5KR4FsnWn9YzSmJ08HjP8PgpysLYpmOSqZvoBem23sPrbUFf0EavLdFd2Dv2WXlWkPB
Z/P/jmj8DOvLqvEq9c1sNIU+SU+vNS0k3tM1gYC7npCgEstAWiwIWLUSDo6um1aa72cYv0JBUEHh
O8KpRIKOYx+WjanO/HQxc0qyoSlyAzXrizwDS/3u7Uygluccm2zXDypRt/k68ypRUfr+7nbf6XgU
fq5uvHtJT17WFs+SxqsbMRo6l/PCOjvr1xXHzNU5wwg3u5B0zMLr4JT8duHR59BvYeD0v94Roy9p
4GINBjtaXIz8z5lm3fmolqHFaelm5n+iYPGBW4x5feWsOnW8hlBafHkB0r0w/1TS5cfLcYhmJopO
ZVEy1mUjZoBSo/H8IBF3OEjJdd+tI5Wpf4+ePCVAgTIRqaA3yZPkR+olIcEoTRx2HRs1UT9BFlI3
Ew6mqF20S48mIw+FS3gtZ6s0V7xp/uSEKbNcgUggEdxEAF8gfuf5uRsa1IRqe7X37Y7s6GN7AgKu
gtontkjgoGqI5CKIbH2loLt+ZmATllze13gthFU5vNF0q65z4d4fF7yhbg0AdKiKBq5DmO3J7GO8
84X/HoCN0uzI17WOix2u/ldFDTnXbgZDlJHEzrZsc2PlUW3Y3GBI6rC2bm4rqQ0ocGL8/V0cWkVN
I1uEDBNl9Z5W1tTO1R7QorhwUZI5ayfs6Hzjo4BAuav7EPrEa+iOP5/7myuadQKBVUAy6p27sOlu
Z2MZzbpit2DswGwwXlDVPa+wOLwVoc6hyV3F2l1gzIm0UqKBUGKbi1EKsn9VVxXj3y/df1oRSjZH
xdHkTKh9F6KYQfjVhMcNyHYHRaRDXZZa7hfgYynawc/FOJCTkyL7jT+YUzLyE13uJsbKZqvL22P+
AdBp4wJ+CTZdQ890WuQWhGsNYUE/pJr1yvvcIFWh3JYOL121c4iE3M7tO62KA1xed86N+CC+EFNP
3OAOkDwUc/scgvb5CPwx/kqMg+ra9/qfybUeX6ybqP52Dp+CeUdMsuxwyXDEVQZyINWydO8fMUAy
KMeoc/sQiW+ETlFXjwLUwkYAlP9WxtiJ6ayu+fzpQejd0vJvJrP+oexf+WPsb2naugFlsK4NhKg9
kOPbDJJ1qXA2q9MgKxWk8sV7rAgLRjlNURJf2Rh0LbMUKCiQlrY/3n1eB+Lz4Su7zN4rFOuULdEk
aWiKyrFsKykd4URefaO3UK4ib4pMzWCppspieFV48tgOmeczILAXtZYBPEd/owfxMIQ72eNfeuqs
2OZMP65rti1j9lO/V7NtNS82amiJWSxZEtA81eGGBiX2Scf/8NXM+OIDyfU5jGWSO0LPQlzqCC1e
NqSLSLpAPY0AFS9WzC2fo5ZY4dz8iXLSfj3hIG1bf6slAbxOxuLqPY/Srq0vMUlN/wwNe57FQNyd
8Ty1NkTDv783sL3BLLWielPNj7lPMqzr5SDZgmQXX4fGGIYwVFQEat9QY7tNfOJ4EtXSKv3QQ0yG
UwSVqW5PJfdYHj6ipg3icoaV2Ie2ao/tyP0gYt0PTyefT75b+irBYzanjXlII3pTKS4XF6qEYl7J
nc0wAIpeCfPY7cq1JaoG88Xif2TE2xdif2Vzf7vmSAfZArTIegh84Dn5cCt/fs4K97wS69hpSz16
cBk4jeWW8wSWUIT6YopARE8aix3tDE8ovbli5WWZloVscTTM710aDmFX9LEehk782BUjXU3qkl+F
WHoDRCelK5M1Z+h+cVjcU3yGefVG45YAy/N15JNk9qOipeQjdY6IXW1pmEdnIe7DUnD//H9LCofx
RQpY8FDHIlKf1KgaCZVzEWhg5Z0qa1NwyvS+CDaQQ9HL5Yh88V9QF2KIeoxz/aSSmKT0itfy7Gil
hGq8VDJimA+/mE5dGsG+OTVCY1wYYF+nbi64rXXIDZo15eP7hUTZlcke3eXnmIIK9LDR5tmoNEWV
OpgcBEI/ZwLev9GdoNE/HEHVzU1WHRyP0uQfBmLdK87enDzDTenJNCdambTnqME+IP2FJNQzsf3g
1GCbIhvJHAhHXzg2mBk3jLJPlxjXHB9mmXuJ+UEjUls3b8+X+5jp0HcqDFVYW/+wRSWDIwawdA0M
06idp4GilT1zwCxi5sKQVsz44ttGfFbeFJcKMYhx0qIOVLl8KTW4px3f5kw4PxpkfFEZ3SB6LLbv
9eVuCnbMduGCZ2dizP8+FeO7uulB3C1TO9Tfh7jamLPSpJtErEXfUtXMYJqqeACb93pFk2vlfVWS
1qnGAbCGIBnFJytiCgCVjXshw4b0Uz4kqqcUuXgGV/ngturUBnQ7ZjK2UF2Ktg8oBPg1LxVxLLr7
y80HPSOdy51fiIEUS6WkKTGvtynCFqHBpNfOuu7a2+gqnPpVIa0S5uMThBwmBfzN786uZ/LW64Dh
Bby1shwtx6wIEoeGpSpZdpUaEbfQyyq/EuF0OZYBl8eRH8CWuM74eiNcWFh87dSnAKxKQkskDCTS
bp7+e1+q8/dh4/l2N1dr+vlKu8I7sjIJtm4bb8HH6F0bYzWXGBe+pb1klh0hDmgOOUTha7vo5VYI
ds/lNlq75nJu20mOFwL5J4Cfs3fvNJ+JRw1LqGfBCWIySWTa7jmg/0inimkwPiw/gT0PKVf8l76M
AJXH7ft4rlUL8vLyLIvRLGiA7NvFq9ZM83CtoifqH11OZ5rHNIxxY9u/QntO8tfpe9l4vNC8cPW/
A7mDQ/n6vunmDUivow/NPQiM2KgSF2neeM0DhrH4lj2fknS4DRSumLj6+K+IQ1n05XblWlQiHZvu
cbCaA97awYQcxgtSbKeloI+9JNsHlGBQmEMy3XdswM52l6aEJPEa1+RK67PhLgDALuGKq/o/PKnf
XwUH/GWIlzdZt89yISXcGH1hAYdXdSlmL5qXK/BieTCqbj0rtqk0VQgWzlFeURY99v9RoHC2UeTF
3IeOgHOxGAP+gaNU/zknBKV4vyqBoSyxRaKSyRzTPd2NQ28g7z0NJMeI7fsVX3I9Oyzna3O/ZR7l
acvJf9oYfaIKZL+BeeSNTXq4vonT1NI3wmvZBwRHkqCKnF9ZBDoJMJCHwHj4DWo0BeayToxw51+x
Sq13ojuHJnovQrXj9j7+5q3BnzRwytWLDLNV1iXDAZO+5VZ9fcGMfVkblrVjnghi43cw6uPsZz0X
fRaFXlM5jNr2GDwKcjc8phswLXW5I8WBwpyToCHVJ8RtOaoT6gtw3aInhmoi8cNM5u0jeYBwppug
2/4QzIDtXjKVHBMGQHHWutgiTdMy9xguE+NiMaoeFlwOywBy1zNw2kpgnQhSkEsRwV+xkrkRmw4j
fUweFh16sWdVOMGpeo8qwt/mruVhFXIL/D5yN0C5X2BcABzB8qSYWn6cxzErV77iVDi7nhaioyJQ
PnvK4Q6MjAMbD6q42h3bZgFPI4qznmVnyLkF59xbIkNiD4Qh9MJ3eMxqlZLM6PGiVQduviAqYMAS
pw2+JdL6C9k8MOxUPCVhz3lyP4exMSONOInG/SIQHuc4a9JM584VrWwUinA7LYkXLtkQKccGOYq9
gpRCIupPc0MYn3rJX7iCjFkj09n8NskMn1sr2UnOew8X5dBvNxijjERym+Rbx51Q6PoLh+oBIv8Y
0ithVil1smRolHkZjbXI3S7mHJA4WNmO1PTduSwE7zTAowJihfoJGLySISus4zFJPpsYXZYC9Lzm
ts1ENdRnwg/Sz1AkQvwgSMq4d/24so3N8RGIkZie1m36IF5omAR1Y1G1B84T3I0qf6MA2i1vlNZ5
uccbNHvBHxIcAeFWtnJCn8br+uwEipMW/2DtTOMUGS7Oc927zfS1z3NvnqMRykOxe/eC8tavh3hd
dYvp78kSGIteGKk1kgk+rnQYQje+HzjY+4mPDono12HpCgs8dFwsYrrXz5vmWQPFvEeUFrjhxLTp
R5TVgy3XAbTYjHsdutyCCZCh//WkzYXAA/cb41CmRwm+oxnIgmyZw+jpSreiRb0xBEpa1S6eK5tR
1WEHN6AfCA2UwScr1Aumi6SWTN3gaPSJ525FYMRcyJMCatIJoBfXYjxi75pYo1jjIlJ99tQnnFLG
CPhu8W5K9oJ8TVtIExkuoNQRUy2xopHEvD5IYovtc0UNeaXGQgwtfde9RPfDmLmRy79UhxvbW1Vk
3CEo78n1ImkvEzbneq5oMhKqA9ICCCUAFWJcDQpS1WCSQMSHRxTiKfjXyrLnssDOof2XkoVNC9wD
3j3xtnw8MbIi35KTmsAiptKXiDVX7gukyLtiAxl8NEflvEXzErZlYYU2nE2rdLbxyMPrpDRPYkth
ZyR4d+WBJZYPuu0L86NNyFe+pNc1sLRDO5SF5qnZOylOhclO6ADrBGJRRUpWtWKhGXmT8cV2LTL6
sYQ4fANIFjWcTGN/HsgoY0NDYGXEbo8fNjU1tB3IgZvpgQq/ajsrXav84NmWLtXg+ZM6d/EM5hv8
60pf3e4maXlPLpo3ZB/ORjDdivrjqSC+AwkITRrGOzOAIHSk4njdQpkWVnhWpRjZ8uQYzetJxP8q
HoT52aOeuwUv+3Xxu9J7wEZ6QbyRacBHP2bRhDVC7ERtTfOKJd+sd/IBoaGCv2jbFVuA1gSY0rGn
zcMDK2Yw/ezk5gKaKYzizJ1S+1Pf6YRphwnT56g55S7ADlIzUO9B7ABtcBnyFZehl/mKJGC45lCP
cTtruxigMemXjhWIQTq9xx7EHcp8XJ5+ryBJpbbNLwbyq0v5r1WtdIhiZQYSor3nAHiFBbxMPAOB
Ry1eHokxFviHZa209pav3493l3PCuOvkW9rDFX7QMwjATvJDJKHAZyQl9VlzwdQgOqgeqtXAeNRm
Wp7LRkk3FB36WcfJiV+dl7JPrm79hVXZIWkfIH8lUHZLcIuA4SEN1z7sUeelfUp6A9oKXU1o0DVr
TYqgSEQgRaoBOCq6T5FMikwcoqcDM3WG2YkS3W3nMRS5Lsor5SQa2C37jHR1ep1HLdP3zrbUjFaE
igNkXeP2n80Fu5JsbFjIJeZxoqwH1ylY+fuQbreLeww17LuacmFFQva4xw/lxiShJwUaYZzgQgaH
WVAno8kh7Oyv1XUmwQZu9f5o9dpuwYjSz9RgSzvPOGdQmzcOyujm2gseWL1pfJhb+sNTwjSiVaUv
SvSvqaDZbycxay3JnpfKAnJSRku+4uhEWwnliGDEBgq1rnvasNZeA88z1vREKMK8xJnL0LF3B1YQ
sl3/HZyuh7t9LdtE1luelfFI6oe5vU0xnp8f2AF+WphAIzPnmXjla537dN83ojuv8BFBSGQxas4a
X7RRyDM0/7fHX5ElZDfrUrmlbAa08B5/HvPztJwPYeOYiNEifM7X+whHnVKSDbKx6hB2yj3F/ub+
PGIWGsNWXbRCE6FhgrLmDSXaM3/4ZIAAkLTMFOPYPe5MCqIA0MkRbhf0nZ8WXpCtTJcKTC+xlOyQ
fLuavOJAniK1d1W01NkyZi/QsS9Gv8qw38F7apZrcSz/hNzxg/Nuuinmp5VVlsFjjB8+Ize6N6om
XL0eGj8hgn0toRJR93ed6BULUNoXWnXhVZVj1XxK/lvFf9/Ih1DScZs9CEVeBh2hp8wEWO3cbWO5
5FgUVD19g9gTf5dmrakfBa6L1DcABu1/CRSOyPT9KFen6ptFb24gVQD0zT8JBb8rJ2CoMvNawn1x
tYE8WvAYdBqFN7fYAdb3UvQs4VzlIko32T2/jxlSomM+EPmMbtB3h+ieqQO2q7F6rFtJlyaBOqBE
sRMBPBzIMkzUNOs6WOjOjivSFhwZba2RUtvamn9A+Lrzesf8vpXuFH3GIxlnlCkQELgIb22gQ7fN
6dMW7/3+FSnSr7orwEiIbbmNBndXQyOlBds1LO9STS9ESAMse22G84uQHiFBOerfXGhf3VdpicsZ
gA2pJD3eMzPAqTowbJ3HIopQxmydeK0quhzqNbSlSirWdWtFqKu8noIZKhFI4mUGhgLD48pm9GCf
FcQ7VVBJpifI94Fb80CcazX1G/TeofnM2y6MO2xtCOLPq9v+0nx3m0HnPBRSyK31N0V/+fRU8vwt
IV/0QUyu/TMCTfn2b2lFufnlofL0Z3I3ADXTFOwEBQgFP0syGkgb2YiQbl7Id0s1y7484a7Q4ycZ
wJRbBCOk6XcBK23LxXdqehNr5wYvjbIhC3rLKYR5nnraRAsItlZc+AzMwA/3y/KOjNtBSHzoeQss
luur/n5uO2z5uwuqVR5YGqy3r/hBKlElfob+kNemqAX/eCgU9s8dncBeyLfRiNioDF13O+ReA7FS
ZQvdVmjhHG6LSU/fwOydnU1yjbSKmsh4gWdtFLQ3NHwW6WOqAufYu0DDffyHzF7QTUdw2Jow00lC
hbgOhvRJ/eBmfYsd4Hulz6heb1F4LDFQKtBS24nt54yS7dHO3/4ZQIGeD9JnY7Cr2G8AXW4lrbIP
q+s9c+zC8giiuvQ/uac3e+pF9DV30qEQ0jOM6lU/qEpwYuOZ3fGCSsd1G1S4VKmQvrwG4JxxLe0J
p/x4Dt8KJZCJbeM5zXBlUpz1zr5rPUBDJZyk37tS+/XpkZrZ00yzcdhXWR6id5zSVLege1r0Lq05
+xWvoWS/ePUo/MKL58xRVcxppOwawtxssw5K9sPYRDjvnIAyRFQEJ5sst/kzUZJJMfFsjiFA7yrG
FT8xYlZnYxUyIb2gfiYMqyy/D3OnUd6V5zPiztn/rBtBDinn6H6ysJVwnvQnHn/pgcPkygvPfMeW
NrUmLfKwlasAxcB6N6K710r7jkMnxWiQUuYFLttSP+0emCiIzKfwJ9vOxut330sp7cdXfbbNIh5p
ttQO+qaW0xUZrMeQdTEasuP/6lpJXXS7sUf/gCf73lep3kOTjfSs71xRaeydurXsQCULG0aPJDRY
YT2E9KYaWslqhxHpmYscJjQbyeQcdMJnbv+DsiRflYtuNE6lHBfk+1qQvEijKeoYD1lKdBXi0oq5
SVKqcNdQqX5TSuqOqLnHYLFcJcco4M40Q3rz19N77ZBvEdhDQOUB2XFivjqtxAtXDUoyjwL1Uc6k
FPdZ1xBlIC3jFBjhQRj/GTwZw3e1+kegzvmokRTsq8VJiJfDDXnKplDq7mTjfj9nEWcsaP26WvDj
l4uV3xuNKWYU95zCMmu6z4ITtwRjelbEf4mtiiV1iEdTb3dgrD4FGbTMQWlXdM4DMmaDxUmeyWE5
H5pfWYYrXlk+ogBq5jJolc5gvqyAmM3lbsZ7YjP2RuaDQLCJREq7S3rTP8sBtVWWGIvdQj2wSiwC
GIRCRqEMzsrIBwh1/CZPKqy/jYKcia1j3UJk6x2IuPlt+zWKUOXrdJrZTTfXbpxnIWgef+5ou+CZ
3vrtKQndS8NEnUq/tqKuhjdlQojdndttpAaZbk3f89jQi76hN9HPqQnBIGq3Bcw3TOZgO4uaH9g6
xEv/S0G2aWlLrmT3kOK48tEbOuep8nZApBb4oAQcGMyk950xzZ532QkcXX9Age3j2MMdCszATsyc
Va3ha9QNYctT3A37lqlpOkQyhQSTyoTnC8NGMri/I4lWXKxXaGRh44AynB0bEvfv4rVCvLWLVIr3
cdmELFOwfsn75jmTLWgv/SSsLV1zlfLxwXn/jqD7/BcSKf3o7rp5Qb1XlwJHNjUVEIUBdSsCJd1d
zA/gIVpzneehl5Zhr9m9Jr3hFZ9fH0jeGfeSdzHTD962CDy0+c/+Pq+E4EyK8QvdU6/CC7wl0Cd0
lWkrhJo+9uIKzdDjrGDT5+e96NnlQrj3TQQOrM+y6jZxAPmta7yhqzEI87mzqT1xHrIcSmLyMNar
I6qtjE63PdDeSiHyOvbAYJU+lwWQNmNWXQ0CwHvYO8gjwO8kPnvdEzf2E5SQSYU9Rzo3WLlxoS3n
N37Grp2Z1gidlRdOAP3usaHwb4R0QDcOJ4H+fPkVu66kFBFCof2TOvgy3s3wKC2Loj6Zh7P46TZU
UpK5gV7PgB8da/ukOgkj6nX9a6omlGzG1OCW1dKaim3GxbW9l3BN+kA3fDm4H+INF2vuBvJt2ang
GKQhNJKz6mxYhUFwduSW4yGmoQ+r4+OY9ak7bsNLVWH7joThAaPI+qZfv5K5hAqYhRVtMJFaEquZ
rdGdqOWCvroGFFNvJaIMXSeo/LzY684PBrajLDZ4juy/6bHrX6bwPnAsh2YljYkKpQVdGKhCU4Wz
tynroBh6kNCACT6dFlPKG7ErOpxsEg1B44gI40Nebl5kzR0MO5ZOrrKi5cy96u/OVUNAPYwQNuJQ
b1T4tVu4qPKVgagopMMikfIqYs/rPwC4AIY1qW5WM8KOs68ZxM3Ahwy7LbupW4Ar7/BZV8jlgVp/
CLYrshKIZGBYU52YX40mMx3CgIq7LwQEZefD4hoRiXUvSuulOrwA5ShFN44t73nNT/FFTnKbZ/Tz
4LEjVjXFZBMtuTxT/e96+aEPOLmEyJDD6ihsur3jQIn/ZExaoBfXLa0GfBEqc0tL6zUXs/6qYTSh
n4Xw9J3s43q5SHy4Gr1acvbVc0agGoVHKGbzUme6PcIGOELcRVWiNp/4J5KkLDqbfpU1Bkrh3X0C
zLmzDNAqB01DZ+BfsUJvgqZwCFPLuCVhkLtOzufh0SH39Z1Sxwq+/Q3+l4dNH+gHCx6mFDWKj6rS
87rxFN7Yz9XsRNTNFP/mv41paU2malsHgijbt9p90gExzMswlw3hPCIcz+OOBlvAH0HqMbdTU/ug
sLY3uRkH9bJeqy7k+4ycNyGE+svY9LVqVKG3ZZEwWaAMArV6nZR0WK2soCHTFD1od48YSeP8rH3w
RkmOTg5Fk+voNE3pY26j6GSK4iKo9aU0DEwiqgXlHX0LCI/0rOifcRXoHNWYxXVUN9R6sAaDfJ3s
KyBNf4t4Tu9fMuI9yZtHlLbxrmL0SWG1oKYlCBHPaOIVEUZ1/vuKhiUs8eqitDIF0KcUFZRiePA1
AJ5qej/Ie4aHPcMlt79niBAImSeRgYavkUtfDf5yqz5UgKggf0yvXkUzWvZvMsSXJ7gsETm2ByoK
DQB1bGyIScHXw4QqSqenBrFZaXO+KVNxqna8Q/+bisu9IWqFU/KZo8RiKxGSHji5n9cT64bOjnAW
GfTwYsviHfxoUg6ysJx/r1ibRhKYZ3AJekgemmpavPN9F5vi9aP25gHNVEEfQte9Kr6I+rbajaYv
7A1Rjv+v9uBRlcQiDdBUUL9E3/cgIFV/+cH4CaHCJgUL6z63sYFHxKSA52FGgKNWJpx6GMP5oQst
fz7p3wfdcKl86jRaxXfMYB7fXq0iAuqvfGhC5mBxAft1DXSj9Uoy3UuBNbUiATnkai/CMgfot4PF
220YKS1ftJEw3uQB8DkqUjrAHO3BLKw5FWLmHIBTXO5nnbsfgXWahi12pRlXkcTxkTJpiKLg4zId
P147QfkumuyuDuY4W5kU5k9K3KIgV5RcnqVLj5av9K3yvQKylzra36IE/gZeL9lo6zM7AJS2rAUo
WACMcwCFuzWiXysOqiq13hBPsKf8x8ep+TiCS4dq7E5E2GS352x2/rAVQjdtDC1m8GNixgdwfPK9
tvnypxVEpXBoPSQJGGYM9u2/Tm6Le0tN7ne5wZ18PogQ6a3p1tAi+HZDiCpaHjfyk6NlRMAKH9EH
rbnYdu2KLd0qz7oSqucqzGYI/8GoeDwy0EL+u3kLDQTTyEat7ixqsqAesJDPJh6t8lrcWLp5pkxu
6XOc0E9rl0fX8ijNL0csC7HhJ1sn7c0RK0LryaBSlpDuk1mb/nnu10dKHa/fmuRtWpBw/p2VKqqr
3gmyTAVZzHSOdCR1hWyw62X3ubkCdiVle83fWE2NcvEvKPpqmeVEOSO3PdMgsQ6NNocNGuvxZrS+
YYudAGXbBrTLchq8wFmBpqfYwY9wLWpk/rrHO1wLvI4k+oIS1+fWIRD+hu7wmkYgzmtslTlAPboc
xyuRFrJOXh6KxuttH2lE8ILzVQz0AhrNErb47oh7wo6Gb/SyObZJVdQnJ8hi+c8dOQJpt0PIuB5S
PPOPC8j/9L+Qq8BkUIEnY9GlXaIjs8XOGUJkvOdcHoOG73V6DAo7SRVutxLJQ2+TFUmLIXh8MZ8p
mgdZXt9xDV25xZfgzaT6Q4dX27PknZ9sH69sh89BgQbWG4Gy5iPByG5adHPw3QkYFmpvfJEWJClu
Ki0V/ktxu+U2KZVfX43FYAfb0S9NTXdMXFuZuW2YSpQ3xCQgyOmxzTC4wbHT2Dt2UFGvaJfBQnwu
86XwsWxyQkFFnBKaLme2zNMYKhHTMup+RbM7c+71PSF/ooucn8htwonZhADEJceJV0993PrAXxTE
hVN/QJztY6oOXz0x7yQx8TDW6d7oADqiPWyBeRMbbjZgtvrqsMSLSHVna2KMaxNWY45pBH5E9XXR
OoEX7EgnAY5A0py5IWmziB5NOW0/VleXS1fRXMj8tdoCCP01p2J+a/LG2RPNryoRhY9cOf8onuGF
znMlWATIamf8N2xu8xNx2Wl9GEgquD9801sZpAPu28Ob66KKki+QeWk01r6OUzOeM4R7EUwwWtdn
Wew6IeRoCb1FJasXMyM3j16CxiezsL0mr74gx7WmOjSrF+7nI70rkmtXBRCFVM1w06X+Kq4NLSH7
QhxmxpHnR7YNvWG2b0Y/6NxX2/MEvDIV1OHw5GFlAEcPNujQD8bZMHDfQEax3Ckv6FDyoBxWxrjB
TZe7rO7BkO6cULXrCBoYdvNwOd+JNm9/YQiO1DxoD2y6DbgqAnyl897602cT//p++2l0zalG53h7
zvKbTYWTtjpCaRnIEg5uB8PuFSuvoJ51XCtIfbh80GSk+ZAr0Q6zBBmq8YlJl8QnJciHQFrBg2h1
vfGdlNLZlVo/dHnGdG/esLhY6NybY17L/Es//pn9YGoGFiJIci8het37W8DW7I4ydCs2+0Shv+A9
rph84UihEwHIL1EdRMfndD1MW8ENXMER3k5KiBe6677t2+Odr9r1OaUTRPa4iIlpQNiOLFob8qV1
gN96M69d1Ii31rPvGseep03ZPMgLwoCU5fZrqizYHNu8ZBrmdun0XjkMdNIdqQk5KjV3HXrZ0JGa
OyOzblPv7d32WW8oxerteN7DBofGM6f5MNvxTt4Aiydgal1ZrN8DBh5WH1yxmxkePC9bJVoCsXqS
FBphe/geUGq8ndTwerywJfDkg25r/61RshsY/uMDle55VRJWFSElxwoVVIGn7g4ts3fbxUOSC0Fn
fFLZ8/dn6bZmDGxHc6jgmj6mosq1evalHBmGX6Z8YA52B8m/oFX+tuM5vp23qXuUGH6KBiVlqliX
EkQsFAREm6tDgpcHrN1/6OXQkD1cs12xHixIMNtdh7i2r5j1cGCd8370hjiPr58OCaBfum3hhDpV
Fsz0pBobahrg1X0UhvPTK1TMsFiSPWenWhIRb8ukx1wAH/dKJgs6FhS/OhLJXS7E8ieYBE82oBO9
W8vURCOpigwUO4xyTzYNYywxTB8MET0Ng9dapGGXe03P8SoetGvpS+RUraABKQbF+BG3nqjG+g2p
vhw2MmQxeIoEVOB+LNP+zBQviGFHh6aWWWi2dde1Kb094DU7LvCaAMqA5eABYuqozi9d8ee3uM9n
P97FgqChEWyoLoO/uIOoAKey56FAyNBQgP4h+TL/Yg2JseQ4Iw8FTNfoUWvtbA5sargFV00Pgr1Q
iu7zU49S7lQE+9ndmiYegVsyHxBJnjLHEiKAPOARHmJQg4FN7wJRwNTmod1W++63zD+JxtV3cO2U
msOMuPhGmt7akmimu4W+1hTIMnVtgRRuKY3MBmzt+TUaMtTKBljM/faM+0ZMewPO+7X7sSlh2IsC
LavHp+lkmDgPKbSrLSa9ae05tly61b0CLUD5L+i52mJ2tFFpNn0wImyTAa1ENR8abPvyeKO+HnT7
zAt/eck0v7vcjLwifBuDv6iY0s22wS4QcocibbdSBd1Eb7Vwduh1uNUcmFCg7olrNc/9rrHDWPaa
DKjjWQ0EEX+Yef2JP5C2P5C6WI+Za3OoRHxzV9REmAQOpOvpLwT9kMdRmR3P9ap4SrHFVaipknYE
2AP2AYgY1LgXWc5/UOLrIYtJWIQjkUx4fBMXPow96RNEysACGEPlzySY0rHzeZVaoUrxEmXnQZUZ
taIBtTfaCbNv0RUgnoosjq070SD/7HqjgIKCjCmYrajik2n+SCZO72+R/DRC5RvzgYsyuMu+XWpe
cu01cJc0mTKINzMSJN4WS+Z+RW7E5IB8PbQ6ZE7wqM2h7P6mAxs+vm6zSWw/aq8uwDFYfKtpPqdp
0q7yhd1cMv3LifSqdrG25Qo0iFVxdaEA9DEKsBtUxu23GSjXI8cXUeNiW+y64AimHCUJ5P5EUite
p1NwVTXvv5IPbBn+zVzNgpJdLlpfAIhkJHDZ4USkH3TOMTwMyTdXYtuE6pwuWJfawydtvE+5Pgz8
Lv8R6XlFcZuPmjqevC3ybA2vX6RQp83bN4xAy2nmEBnkaH4icVGbFH1rbNVvEt0pxmqnLiLD3cej
CcpD22kkHHDbRve5gZ+RBqo9Qej4wvRx+af5T7lpahnm1AJLJYnIIz+M+iQ5HSs1h0AjV/b7/nTQ
FMMg1mIDFXqPBfhnU1yxD/Hp265EFGDv4VT5jNUeVWT+sccGzwfsy+wqfm0XOLWRLpEL89MgnoW9
eNhyKQcdIoWWZ2uuFU/TKReYVjYwDJrqmLrBrWIBxpzIYXOAbnMpgx0CmvDvEneCb2MfJFc4vH7x
gqf9Fhb5lb++YgOYFuTn1k7drfGV6nuvkqDFbcs6ynGzcciFmexpUgquUntuXRkibjPzK5Q8FC51
Pb5gDr8DezZmhjVrrF/AJwKc1iLyBKjPkH/Fq0ZdCFO1mLK6ytiebjIOZIZHEzsQ6Iy9J/ECTDzS
Q/z/ogoYWfKnb9JrzKhjO/B8GjrR11WetT9qP1syQkv01HmERRGJBC0NQUShwLBib291280dMxra
6IHjHWBUA45Mvy5z+CdqEUJQB5xpu2nC77yqBFQBBXdyLjitEzKhTsj5IB816BsFs4m9RM9UKvlG
08g9RwJnvRHIepUDG5GkgOSfaN8kD2qL0ZGEzEsJNaYdzukT6+Zy/OIlIebiW4GoD+oaMxRLIktC
FiwPONuXl7QZOAhTwkcmlRt+G3p1ZuZXj7py5IFerrc1EV6+0KJbgktPps74x6avNJIoot2IyFpP
hGNJawrBAqLt7bk9tZ7frxxk9C6wBX6y1VrOZhDOwzy2PBcgwLk9UUjA6bSQxFoKjR23mTzJ2UJ8
akYH79RZN4iVeHE9pn/kUMTVGETeNPqhJCbeo2wBhmKCQVPHPHSDzg1yET+DQy/KBz+ye9v6lKOC
XW+zYiajJHUeN22CSoFaSAqvtJUqzPUcTK6DJOnY47yM0QnJavoJRiYTi2Fc9XLeRz8SWtFPBZ5N
AdSGNEEMxty7w3k+zen9VtS+PXVU4stowE+2m06h6hJx6ySJ/bN3kw13u5rhKk7oQ5B6xLfEV2K0
NrRoXx4UP0nVUO0/rtSF5Aaw0BCIq+S7jUtleSM5r2Iy+RtrU9EjwWfh1Ph0sGXJp2zc384P9+eJ
H/U5tMFIR4FHbAZZ7RyVuEmQcOrK1zZsLXHuqL8uOpe0UEOL2vhhjix/FvH/zUcSd1lVIaeGtyW0
xPsqSVShSU0xU/bTExbcebnTYh++IWJQJYZmQpcmd84v0tYemo59MWGJicHh+J7b2SjZv4xD7yTh
URXv7p+U4vfJOfaEMn8M+xbbPxgTzWLbQG+fRK/W0fga/1arw5lIV1G1tIx5DstSYOzH9CZ2sRTj
HHZXSmkktBzhUabv5078trFOWy18l4qhM2FS5Y/fgVhTlQE9rC5x/P7/8Bmhs8O7vQ9HB9YZMen8
HVSq34KB1zmM6hXhRf/qWEglPj81TK5/dwaI/I05ZocJhcRG7ACNikwrgMWijxO7pu085aDFd5Jn
tlNa+fFoc7ANfaBY94YeNuoKw142e/dyxsxtQS0Ku4YBQBVy1SQovm7qRctdYfCLNUIG2FD1PjLd
YD/1+d/EObGQtUpDX49+JjsfFwJNoplK5PNp5srEdBD+xFuexVRRsha/li0N3WpeJUH5OJPlNp0I
WSbUV/UUXZe2iedt2rVYQAoZ7rX4ByCge2mszutRMJv1QFLvbeMmdgwz6nbPQuHVmF0H4SqVdckv
OTHCg3qfUHkb0SgbeMLXVV30RF3hG9rOZd1qsxlttL+fbByNUCp5hXqiNJS36jZBVOtB2EvwbFe1
MQPO5FpbgLKZ3g4dzgRpawmJXUys/dG35e/1hRwtnNCBTV5GBFhnmoT8XAYbsRSPLjOdP2JqL0Ij
a43w4NGLKB23IrZi9IolHRNYHtqy4dumpQSpyXmPr81OOMuAXURdrkivGk8Qto8wfUN+TWvP0XY5
ibHLycoBEy5p0kpAuzPR8ORSZ0mivP5ZMFggBTX+Hp4pw6qju1IK//mAjo+qyuCjdHLUydR3Zmsm
IDbzK/tgV4EaCW/M/qO2kauzdSH988cgL860PaPrNdP37ceIrHtMlC6VDnEfSPxJlpMKxeIa7+D2
Inxv4I2yVr9u7+3UuEPAkLBN3uFPXT78kgEworoYI5A2Rn5f7hIhBG093bnK9lm69N+DTwKrVN9m
msO0g0Isi/nWC2BGhK6TQZbn+ly4DnN5cRnaRzaWSqkjtUmC713rsuWVO8rpNWYhUT8cEZGO/osJ
f3Yojou+I6OSOx5ONQNqlxcGHJjm+ysSZgETANfGOXc5oE6dmjVVmYKf/9LW+lDB031eJs25lZJH
d5pgLiiR53GLrKMMasP/i1Y5KHi6BjxdaW2ABxE3aLISjXkakXP4NmDeispFrFvkahrzkjBhVCfd
8AsKF3d9NUNaXwOxDYarOwexwTfUCn9y8P4+MX8g4o5WbUhhD8dY0Z3zgQ/RH+/CJUZX/6+Z/le1
TNLrtYgEwXupVWE8x6Ec7XhwK0YDveWxKSFLta9oLwcpFlZJawTJCFc4HikaemOLU9wzOkP1Y7Vf
FWNnsjm/D40v7TQtgCH+OihF73X4OgDoN/rBiCvaCPlvDSXAJipwAPN3nLbUFSfnLPZgbLSz6jxm
0cCvFCUKLfiIt/4lxbm9p5tuuXnslfhis0wmAofbK6Yg/kJh2k1V8n/jopfw26fTcowYF0X2f8K8
24Fa1EZnY8+yR68jQhhBONCBDoP6vWjVn/BwN4AB2Ewt+bC1QFqokHptFERLBwcv4ed/7vwyALmL
ttNCeDNwVEjrRgUSrIWhu+6FvnBfCufln8lf6w8NQtxNVBHtdzBauXyWmY6QWjYKUYUaoxOgfqIU
MYqZk0Z7c7NcFRlVNMTFLIh8LwNC3igEc3YPEh37YAp1jEaB7uCJ5vT9JQmyXhICnYBdOI/efBSW
Gb8Z2dMq1m7PyEIx/XFDeDzCRKG8J7Exe8xBmsTsBlL/XXxVTnhBf0iqgQWJgV37VcouSJgpHdE/
QJIYVR20H0rWd2dEKplG8YBKrK9keFo26q9Omi5GFoVpO259EC111aJeVBgRAWVJAHus6A/lyKZ+
ywjyC/ICgh/JWq10//V3bNVCOySi0MjJAY3pkGXR65iYOYGBfivQGLSOc/HMxI5+un9928ptOhJ7
bFf0YsnEKV2MUfDDte0Nf4bKd427rfw4megbRAfgzFuTqcuSi4Dv2lF7Hy8yFvDxpX8OUO8qW9qt
A5C7HsSsQT27iUuRrD/OGseZNOepLogvK80LzGj5AIVxABg+Xf9Fg5J0t5DMEUpzPhUn4PUtWz4K
fOm764mgXqX8lEvjXAP4WkWev/Q62tA8Y35/B5nDBlwRHC8pU8jCMdTbcWUWMrLrZHLqyjARCCFd
mp/HLP9h29LtacT9m+EvvXqkrFKr+4yCJsXom4BgYw3zPoHa1rvhTyF9VZCbaM8zTzd3y3/+bFof
I2IwAFkO/4yIQhR0apjt7YGsGb5Jo2Rf8Q1VhEjdPfLPOUfhSzzZO9eApINosr/gCe8E3Q9VMG32
0rLcwcyrKizQ6Lqa2QZ1VImzlzc0RoSugy+VRS28mqbFOMcnhlJOWjRydj8SlQ+rRK0lzDGU//8E
joSt8PJKvFj0irbFarwx3DVMDTvPszVYkf7oYiiniGi94o8UmvVYakBC6TP3V+5jw1Pna07vImbJ
1K6erSGAgvPxEisPceLTtQhZisZ6lS/9hdMJ1XpdgMhqFfIoQ3kUQ+shgVfyiAs+afwIPy7Aal8m
7YFEZE/BwNhgR7BaY2qHCvNszX71xX4QZqgX0dDSiVsI+AxYcVgSyeAjmUUgrkXyfUivR2Y/Zo08
QZZ28mNtOjNNk5YVj20o9/NlkDSud9PsNoflwHwucDf2umOGdzzEdh+ABTRE4JcE2W1ooaZiueSK
2NAMjtgdbijlKCoEnFOXpil9Tc50lFuEJXT0X1Qbk7y3hH5w19rpVHHhp5FJuCwud2N5rl6O4wlT
PaD7yA4KcJXZK3gs14IL/GSoawB+DUtO0ecT0TxD1Y9zG2u8py8FViyAFw0WVHqcmU3gdVGpDNJ4
bkSuH1lM+8HnA9dX35w2b4NG4MybMNU3ghJEFKt0+HUfYjRlNllJrYYsoyxu9d4jSTLTPztgyMT2
1VSwjtTGpsZJhxr5FPjIidFKmy+mghCfA2NpUU23AajCdT3i/PBVk15JVvmYnSgZTJpdk5wUkYce
WFG9abWA7caTeoWCqOJX+lnafeP5Jla+9DzNLtirNtRqve4Asngu2jeQ871Tfe+lU968NTCapWOW
EUQMrsN/CyC0OIvMS9R4Emd4ENuR7hacwTe8y5UmXeua2KS1YHo0iEGHqjxUmxf/e0Btb5kAd+Me
DzIg+0X87/OVgsY20DlVqI9fjtMrG4Tu2yBEblCHp/fLtUUPzihO/Qu7XCZ2Dz2SHA4VqkgyOvkU
YGSwPRRAOXEwtzRF1H4hT6u8i+xUMk3J+fKuvEv2NI4dk8E6dSyVmGjrUHFxe8Yzb4dcWuNPfliC
880hKlWpikMwr8WE2aF1NCra0Gr+lCbOlYhmA5Rp22lbypGIgQCEpx6HmaV5AWZ5T0iTczfuHzU+
/0nta1hBLA9mD9TJlnx7JJ/rCmNAnmCypDCZkH6QAZ+myKEZKiLpf5EtYshotQhr2c13CnIAS8iv
TQruv/bjVzI6zTocJTZrE+3Z1N9Tk4D3K4s/QgG5XvGPcSFNxw6mLwuqy9x30+bzbq+8/RclZiVr
v/vRGNSmzUxhwIuMeqRK0xhtFrjTr1KG1jUyc4JL4IGZYLbxs+ykbkg2uzgUpl5USotsvE4S0E/P
QCIoqBYv1jNDg2R9+HrFKZfJG8WhU+jgIAJz46cKbBFBnSYNT/vNrRwCIPjzrvHJOOX4gWrhUGto
LTIzXenaawN+xxtdzCI/02X1bKv5Y2RutJOw4zktJIU/tM+xQb9Su6LJJ5QBKfkoHBisGnUlDg/V
XpRp8WIIEG4f0ZiQCSEEAeyA05HrNCmPNat5WFclnvqGHHoOOQZRDIKDMw5dfEpEyz/0kdq8XooX
PM7ZbacdpOlhLz7//x4n67f4X/d0KrlHWNYzD3UbxVIW0cnyDF3ATPJGtRxjDZoxhYsuwV2kZIaP
Yu5dQ8KkFlxs+Pv33grr489lJMV4m9yd726XFtUyrQKy4jaYNy+h94Pj1ZzKf56MNl/IetpkCS/v
kmhAh0kYRXxIwyOmsR1CfrmbLu/PkuYC9zqi2MFuDWKIeg/NH/W/7tmuC4Wt5YhT1BaNym4YgQd4
dDz7tt5EToIjo6ZH+yuehGJTrrVcxjfzm60ouGFFwZKOXHrsezJY5OYx4EA3J9/pC2TGM++Vh3Uo
kwTvmdwWeWqrBBPM9kRyfDfGke99TqaU0QjZXgqJye7do/O9fPtKgqpkC/I+S9kZvXDMnfj6G5BH
fynIQyLnn7SWKAq0jE/gnla8qz6e91L3rZg3ZkKBx0BjB42GPFY6pzIfIJjULCJLDco/hMJY01st
z9VS0LpDBKbUUkXBNqZqBgTTOYbey7i2tf+p5hCzQply8h0oxcl+R/BFJ3LPi5egFjn3dyf5KljJ
KZMMK2+EoVdke8EIiQPes1AoCOHiSGrnhV3rCY/qmfj3WZ24NBPopQ4dBo0ayhM6xmllY+xbcEiX
hpM/zDcWmpF0Q4nFDOJnszDGO1IC3mSeqTixll2wXRCw+s/Ducg80h9lJgoICaXKHl2Xj2b0B5aB
Wa3H9b4jowetWdsP3R9KVsxnK26Y4MBR8dudMolOpMkmGoxJkuQIDMRtFTFJrOMZiGuPrR523lH+
5lKhwNWWfTUOy4L3BRfil/1pUYSrjnZ82xFP8foof4pDJ13hoMaTrj6Eh5LZXml+mi7bLHYECP1Q
o1jjdNjiwLVi1U2qM1bXK9iTobyeGXD6QAJu5eXJ+mv/gz3uO+V+YGF377f0cmOhe1Il+PJjl0Mt
+4CxXg+0hshVbCOqVcIB5WutL50BnyhIODbnwvLJR+eueXrELbd2tb0gWFCd/KXQ651wWBHTKbNk
hMVXhdT1VRKwJcPHNUGpQ1WQxbwTIe5DC0aoHfU+gPmbbt4E/uGetTO2pdr+qYWYJW+ufGsgRLxM
oJviO5AyF6FH/qWaUJwE3X/5KBGNnfrlwbYYChX9KYDhWvNgYiGX3MLPgI0Rcb5Pmw5FzHjf/TPx
S/NBrkJZAJ8tSrQZAMrntG/j/0wPVdpFF2KFoc4B9KIYkmDKVYav/1GtTIILvQMPhEC9HUNj2WAX
/K2iFIbjAu8mJob5yL2jWC9P9BwQjXcVQwkIM4fx21X4YuKd1d4yPqjGbsV0vykhvs9a6gsRQkpP
/A7fFB9VQm/cBYYtm3zBhdh5tRczw4lLWtWaLMZVINVXZCxMqWkL+fXtU9OXUfpOb//u0uvJRu/6
UdYF3TQSzqSS0ranvEZMd66BCl4KmQSOdmV+kTFNNpyrKtllUA+xJcbqw7bHl8rLnrPEiQni6jst
Wc9ScmCm3ksNEGwJRMCwhpKYQbNEoQrAMmlCWjCkZ4FV5Imj1BeK6FqVf7n0BWn7vxHNZ2kZ4z+4
NT1VpJ+GqBkL7cyDVDX+Sg8FCq4Nt6u6ylDVui9h1YUcvzR3oKo8QTmZDCxEBbkwki6Qx81ARk8B
ap07pKtilx0n6GCUrv+OOPhqIzL1603ZpJm8ECtPoI1TiWfCC/FK5mlxFTMXBSWhcfl58jwRGG7B
za8ZV3jrSsCKDwSA5rUbRxqjE1xMf4+v/FrOhZ0Rqq/wYTc7cl+a2JCl6hnVaFQpOUIGHZxR/0yO
9mEee2zU97JLxKwOoZGZ+whBi+vGPs3UoFY+j9okt9wSdB+KPWuaJVnZg/8wKN88+u8OJ9qDLmtA
qnaYdy3azMAjtezIUK7dgsLX3/jB9dJGPv5k19kjmdpkoxKxZGCskI+JXRfkbOoh6L8+I/z+Zq26
rs84LtuU8ue07Rwj1Naj9ApJUAtb/D7IwbpSQZRfGS2Tmzh1I5NmdlH2s5nVtIAQ5t5803+A3cNw
Aqw8mMLE4cwaaCLG3A4jqgP6RV8jx5E8z69G7L0Yjw+xUYzdbVr3Q3KSt+lqDE5VGBJGcherw5zB
JPjgjR2yZ12VNe4ZakuxGW93GiqpKl7cFIjw1DjLueu00oTkjqPIGGDi9vut0HEt6jhSVSukjtnw
fNmk1AupWCNNTVFzZ45awnfCrsIPRhCyCQmQUynMhG+zQssC8fUeCQkHBGGL4b4LkTp4PBk0hnK+
+Jl9HmpnIR5nyifWTXK4n1Hz/CRHl2LqQvvIxz1I/0g+hv9pdzT43GTCRz4Ecz7xHI35QHr13Kxo
qAHHElECb0Y3vUlcYm/hyUu6re8sbEs9XytHzstxmdCo5YU85xdKWY6a6FeAUR9GcboXeS96e5V2
OhTwvfQY+Q8xMRNBd/ao9ldlDa26gGLTpnlc1YBt2ZcXKMit/A7/GTxUaiOH1rPNOnx2OwhDRjDN
x7412Lnl9u2poo/hGeuQwWOYGMp6qLTuyf/m0cd2uzgkAEJba/y915ZsSuNCi7m8iM+TX0NbrUOr
wrM9itQnmCLchu27yEb8QyDZT2xpya5iMB+T2wMX9ZQZ84V5hrdqfbYn1l20rg80Kdl09S/CnwPg
rpny5NLhBuuhs4aCgPhij8ERJ0hsCS64m+WuT/az5qUdM9XOPPcKpKgCVE057nDPhwfkLay5XSIM
P7E9jChDz7htVAov6fq7OEloeh1+pMd4AZdxV467npzY8jb2rU+d5iaIY3EbXKb79U90ZTEzdoNu
Wdn8Vm8qA1kyGjpTKBauu4q3C5NxUjfLKV46rZxFvW6Uo53TXYqcEkKL1m1sHssbuGp/aZdD8Vsn
yUfl7vp5S79i+vXCYYUs9crQboP1sbdv3qjga7VbcL9btEXLZIwZtE9G99J0YQwbpc+APAb3PjcD
HWAZoA++i4kXIrrsr5LWdk1QWGJDYX2bilxyqAeP7KhwJPC2N7MclegZYwY7XDAhDwR2x3ZxjkFz
u+INUYBb620TY6wYdvHDQKvUpqgUOgXgH9KFwR3Su1cOaaw34org6zY5khyBU/r5E3nTxKp1AHdU
LkoAyjcjPAQopQncMvHngLWnF2GDdh8v2GcA5E8CCEu+r3pYD0oEKN7AWIsewua9m/IPSajObYip
7qENRG48YrBgO0fRWDQtr0eh2aR3JF6EE8LA6SxixwX7o1YwNqKYzEqVz3ill6EtxiqOYIGLhprO
1Va6RE42BaMFps6oPY9RHPyHkjA+useaQSssn2sHPup/ZsTRcIrxtrulcbGlsABmFa6/LHX5Aj6t
X3RknF6GHS4byrhwNz5ThvRXHyrF5X6wqtvq6/v9uRKzFjy6xTxOndZghB4dqk7/6W0Nfh4PuyPv
88MkeZTI4/4rTzbSfkZvyS84NJg0JgB5sagSpa8AtKsTcwI7v1gpGf6Xh/m/rJnwsRFvGaYCIR7G
I/LhB7+R3tgXzEED6tMwoedWL6rRe4XfRhGIMNBWLjRqKeHeVlqgsrz1AsefCXjtqFVEOcRp1OcP
p2kZMxA4RrirldUVU+ZKzRoZdCB3LCopLbOmEJaekxoMLlA4LeopRIwZWtlBg1KJdjjFykljElrP
W8mbIWRHpOQ5TxskfvkCYHDkiYvR82qdsqhlVfih4aA7BVW7WcWYB8gWldyyCXR69Ba+khXtded6
JOFaHOWVaPvmeODF0NbgUidTEakzvYscVBBoTXAgAZbLKGWrrqe0bV/iL6PwII63M438iRTucXOF
oW5RWSkrCudPON+/7r7eO1inVJ8J2zRE4QPw79aXUd7pzqDzoRQFFwKimGLbe/XnbCSFjHdyOng1
I4sMLniW/IPKbeC8wrwuG8Ew7FpSAvLu5ie36PGcpycAFKcf/fJxtBLFw8koL+wf6HlFlM3Jup5v
vf7g2DpLNfQG+2yHrw3x69jH9qyIvl/NoeBlAdKKG5HCGUO//RW/Fa+TGUCtDp2LCEjf9fjwpdR7
tByRLfBJ78ZtubkEHSYRu/yFQMg7N4ALyK0O2adIkq7RkyzSruMne2iotWz4dKRhnYszOZksU85z
AvCTj60Q3euG3bZSGHRSqbyimvnDRf1dWNCsCU85eLR74E+wlc9Hh5OH7hg1wfIzTOjsQ69ggTFs
05vClH1eJ3CcWS5aONt+UWACJTldmLIv1Z8lkXiH0Z5oJhrYDRrh35kgIDAnAi4Ef3ud5QdRGosL
9n2rVpvGDi0S3/M6sSS72GcFH/X2p3N0wwGcYYT/XZrr+TETmYovGMHLQBOGFpeXGeJqVrYHaItq
fJ4HuA0LNdRfLSHfMF8NTYPI9ks/a2IyB3JskGQKdUAlmSsBX4ShaTTSo11R2WrTO+9GBiedW6nC
z4kSLxewrxTI5FlkoPFJPKdDsw9iy5dGp/Pd3aoELeXxWTa68wJC2KGgV03vYHB/qPuYj0VfcW5U
cDuammxxoQjXBsveqMUN741PIt1nWhINenT2X34+DMxA2O7IzR0wTwYE1k9rsRWNFrKFCLF/PiBY
l4n9AIUwAZoxw6+L0XOBPbK6JfGz0bI3UjBNbuzxUMEFto+A5fCt2G1wFtKUCvY6kcwu2ia3pbZj
688lv1JATdT1RtcJaE8lvQhqTOEDZxzGcihaQ2m3KGWZzhnGDgFNB8jeBWHFKYSk1OCCWlZynndD
IqreOeypJp51JiPqxpAHNnPy4RVo4sVXkWZoK4BCWiExK8LN8ds5nhxMi9Ql4D+R0asKbth6yXR6
g8wVg1YDlBJMgFvZ7c3Mpd2VAdk56Ae/3f75ysApv+wo9nZ5LQK9eIuZLV2h2ztZ61S2tT6MzXBr
PsuhP42gQ3vgTerKaA+LewEixEemYLbHeJRN4wIzWLAubfNq2PSWWUnh7rWVrtJsnZeHW58lvfkj
AtUG29HWnqvkND97AIb040rXJQVqbKInCLLZTC9maG9D0xG4pn3j8V8AutgQHgH7dv6QcHcPnA9h
eKb2gVEDLRK6DJSBkhJyfNwepToYUFD2jvv4IIJo2/iCF4S9DjW3Busg9V4ETv/6IEieUqIB/Ael
zm6/PL13HbFPB6ZJI2bDOZP6DydFVmGdQaU0qzU6a2JBxvHQ/UCRJMPkAupZMR0ML7HROfb2AlPY
Zy1yz+tg5wqkUH+HncwFIkRgNlrWjgqE2D+Ar1AzjYzg1gFLlQMICJVIsCVeM84Xb6/9OrxlP6UO
dZ/PXVdeXgl1l0GMlCqiQ5mZwxhqDQ5f0l3L8xLa+7KCsMdK3t6iKIE7EevnxeiPGRjzCf/yonWf
lB5bvYthxCITu1pLVMKtpgJV0wkm71dpZiPTjbwb0phHl+d/i0fA0DKQiCsj7nVoFL5tVTgv1aSI
snzZw+9ruGypAFOUrvAZRMcNi1V5o65wuCFIFOXtATWvRdx51SyXBSXgMToqJrO021KkV1VBWzJz
EhaJBhlIzf/NVm5qxv6yEMBlmZLLJYyUpUwoYqCvlZRgw4L1nckTksAEHjtwM+I5f+BSdv4syj3u
QBvCz+WPOnh4l4oHsnpdDGLwby9/jtwC6g38xHhF5sNHCH1B469eIOnlDPNuveEhp7C9hLAW4Dk5
0P8JJ0IVpNUNq/F54ypPWzE2aHW+z4Sb56fRvz5GBn/MTfpk+6/c1z7JurXeuIM5gJJC1CMN9Qf+
6IaVHAdJ8Ob8t6wLwQjudQ5mzn5yUjBHfur3DYJT3zugjx6I+cMxdsRqfnlrrJVAokeTYYW3GHtS
jyrhzoh/RI5A+/h7fZYV71RQYpGVx7L3yKAuHk2sigP+k0KjfVEQwXtxay1zZ+1MdTgkcR+R6aEn
CRrWm18EMs+jqeKjr+6Jhm/mUuryW+ki5PzuZiNcwPJV+Ty6G5xHXTQiBH/PUK/pCBfmwuw8FMXL
z3aIjFgldZJqd0WNb+WdjdpexvmaS72xoiomhDikCNvpOvTC8RQAitOTMc71JiWr81M+6MHRQDyq
k8fgl6V3qlD5qOZD31jamPyO3lihkjGBbD9SvlCXuAVTnhITLLFitKKUBESwB3uF0ooMpmn6ftW6
0nY7yd7mhSP6r5aUE9CWPX588M+GawYCX/+DGwPrTtaQ+RkjGtqZFvdyHVZwgzlGxYO93zrpmzPR
QhmOV9Fo4vus0oNasXHTMsBkgeC5LG0WTJlIwHQ+4s4Pb3lFWyTCu1cnnJiLkYtWtd5eis/PUXyA
D0MpVFtMILaZwkODsDAEybjdvXYpov9WwqGAVzHGbLLTsbqgjbpCkKvS1qvQY0v1+13f+G0j9wvK
heBKER+BJ5HqTxVizESBuQe4GryBM1uNk9BLtv2gKglxxenRImgnltLcMe3a+p3t/R2pARH4hUJm
y+nBnVlzIqM164HF24I/lFzVuDao8pcJ2mEbXQVxIknmARsMf7fnsFjo9+vGnaX9KVB5J8Z9CFjL
Y5frXeOlEcroIdyo4V67ALofbUwP7RhHmfbM+3IvXpNQzpD8okcBYbCu5N6U4IEVw5cHLewEEiLH
mSS/c8JyDW2ApOepsf19LTuG4OTlNGAIWahj0mYPAc3q8UTMX4vQ/GD/DUThLz2CAVWDSdKdPxJ3
5lVeyNGXvy9nBXuY0RcapeBA/31TljOEVfj1S6RkymyJwb72gM9rckDBb3fpl+jZ7wprvGzoXhIj
t5WyqL3ddMg7094U98/68jlqve3DUWyVA6Gu+E4pjvamLlubYwcVUpFrZwky+eXQB73hscRPZ4p2
xvR2QeCC+zl3XV4w20HtakT/Fu23EYNLsYGU6Qrnsxr2JmjLglUOopibbJDTV6oRayOx92EV5B7d
+tkNTX33B/jLIeS4U3NNrR6wYkkdnGqWOwkzoYLkTuj5Kyfd2n7GqZq4gERRQ6UM9dj0KQdjPt84
lJ1HtFReBZHsCSuy3PpBFtHNa7cfgf4qqgFUNqXs4NTzJLLeFW62AMCC0g9Cwq2a5woTOziRURgc
Zov3fuv4L6KakXS5XGGArgFprPhLtzM+yQRuGAsR6e+c79WeXLtF9Ih0HpcjaLpfmq0B6VR0Lsx1
BhwmC4eW43TjTtYBlXreU7eECIYdV8OCpFFE54PMaiaYDKNdojSeYFF9oAjBRF6VKAsERSOMEpqo
DRrD1fHf9VW17znNQwwBq0m+8gLIVT89EJ8pFL0uGX/nxpRVpadHxjUVvyuYxrSnIM/N1xUFx22w
mDi8Ui1E+HTdusQSnvsoYDRB4lVWIB2wBUJAp0rIFMwVUSai0K3pv9+9gFkC5YfXd950r7kLAkwi
v1T+ubfgL41Er1fBlw0QyNO/MGRkaBLE8DARp/yyBzm1/56MQnvZzAqF67YSdH0isdJA5i/BI0Zz
kqRWzUJ3y1S2Z+xlQL6nlJUdAN6ZrUMrW9dTiOCspWqjBDfpkVog+OUo884onRem/IEMK02CDVAJ
kWUmd6DJg2+GYwbLlUA2FdXArdlTDmPLGbik/BMq5fc67TQ03nUVq80+WOFfW2KUmqt0xsnR/M7z
ziY7KcCD/1xwQtSF9hftOS4Hvo7E2z6+mizflBkHnYsnxRw4G6MqmDUotDDii+ai2g6Rdyy7eshI
hINCN7ys8trKwYXL9ERGR7erKm8lE+LU3XWnjOrw6MpXzt1jR239+M7KZJ2vSk7C+M3/8U1suEMD
gy5vTBctGqHl1Uq3vSn+43tdcILIzxu2ockCdcF7hHukV3+w6+bVF8R4OgH44Y4LQIXOD6SSLHy4
26D2dO/ZqDw0CASN1z9qZ/nosxnJCv37cQZVmE/2woVXsL4NIH5STY4hz4Q9GkFcj//l7/WpE6jA
M7HChoZvquOe7rGxeSt3NjpPM6FLH3iFnJl41yuvtEHB6KumAZConnIdfWlRJoqjVFiNPYX0gX8O
+jzPjK6g+RfMSUOMWB/0ZpeJ8k7b3HwenWZQQz3lEa6eKaN4LOOQhaJ/pgFMFpme/vE2bW41GXME
A+BDMKvBILrgWPCd/WzDKxy6fh5iLwaLTXdeQ73PlDVfriHCtQc0CxupjwetPsMw2yP0b1PyQsiT
NPeaz14TtR1eaIY+JOhTC67SzgVT/45w+UaY3HrBg/vK7zA4tdQve3jf+khCmkttA00T+5n1MzqE
PM2d7lmNw4LbPLRwWf3UjW6qSzQSTkhgTd4jDZMftxW8yuX1iVqiJOeBrmpvMpQcnemTthamKkoc
Zbpzd5AXwzyBGH97hF6S2afBku6MkmljB4pyLHif1sCj1JBd19NklsypOwLwjK7c6N2tt5RHJMS0
8tMutOyZU1XjC/oKYLDGnYUmpLDaWdlUz2RyI7nRELMZurZDkb2gAKK4fHsuK8zmj3iadyZOub00
ccnMWOxS6UIxdOhDYz8gLMyl5aXgZTqu2OPsx1CNiG4oYgxYG/Zd1o/i5gqZ2ToBU+DiT45keo+t
ojuyqAqC6yAhEpD5wd6RQ1Xl5N0pGqgCRutBetnwaO+FjmhgOjligVjna2rLjHZxmC+d5rPI8F7t
Z2gkvZp/PbJRN0Gc8O5/G4lz2RnIkTprhENn6cmMGtCTcwuonGd6iH87feWDYvTXV1sZMBQ8cSTX
mUEku79KVAsGqEvP/uF3qIZp8BDxFPr8Il6NCpXvMe+D31u95gIJpGEaeq8QVSeDPc1K9GseR1uB
LIqkJkaMqe4XBDj2yAD0dyENpPjjlqX0u+8ZRbpZaaHOpW7hE4lkyW6EI8pmdwtMPFWeHLTdj2j8
ZbVfAHL7tRCjXItMjjvD5Tl0MFWLfYJZMGGP7RKrb1K5OA9KzQSP7Un0ffPRSHz9RGPQj/KcQDpr
xOZxEdQrhB7nUT3kGaqZRxBbJj7XO8zaAlGlWd8+XroZz9AtrUjaAxSv6VoiWcskdIxEUWwSPVMV
aKrRvvVYV4MpP3HVq35WU3v7KkUSloZTznHzC5RPldUdyw9TbYFge/V3/x49wGymiA/AlEHn3ry3
k+JWoUS3y6hPckq7JyD7oSO0LgQd2mKLi3ab/eyaGdUAuFH22jmfcfAWeBJUf1ILaPGh5iq7DHNH
FF9Ioor3GIejuadpeAI9T1KQfmPkuJYwa4Xl+o0FO7G6lAV1LpRv71OZc1K8lE/X/EmsrZAz70g6
EO2pOViXVoXiw+OQ5T1Ougq4ZIsDdw23v2Db0+81eYfx9zjRjGM+0NYnp4lfZ363VZp/Lf/lZWAM
Xg+3i0brnXDLG4ZuVlaz1kdWsuAVfnREJZWm8hVUMlzisA3MqXiwIAFDnq6ibEnfEkWojBSIoy9/
lkqeczrc0vAMIBC/JlIL67obe0b3ZEl5yoiC4ObTNQJhotU2z0OFePzDv3RQyXGIM6QEK7dGKRA9
xrPmxyvMSOCgPEmtDtw6C/g6aD1kJjFGNCYwpbzZV8yyfluc7FOhSkiAtmfIpPeN3dVMf/sz1W1M
/kNiwy7ufxvwY5B7p8uukdoQ0nTiyIvsbenUDK3NTdAr7l/8tm7wxFbwCDh8z1SzHse2XN8GfY3n
ENpoL4vAMdBWo5JHUXXM2Z2R7xXg4XmUC5pgOUCryVsIc20Ha4P9A+AuydXFCSbwmSHv2cJmtocl
gIyHX21y7BjA+UBobQntjiQ5w8RNav9EHP0W5/aIdI9YcgLPy8P2S9nBQq86vDQrZhxAoEECfACs
38sGCvC0ZcLCDteOfo7KP41vIWMp5+tBPjWVOyEsUD/Il/Hcq1oRUyF9WdllvtQKWk6ATAtPp39g
Vht25NvVhbHOWdbTi3nfPdbS7AUAae8tChDLDUafJtzU7urt6M1PiEP0bwtUvZNWUyzy+z99ZAuS
IIGpwIWgCGOlZzbT90/EErh42ycfILLHpkzFc0RURXJAw6b7qVXN1Ys8Q26NYa5yjjvShqpLbwzK
ydGRFQDH3IwK8PFc3644Pk5/YdFq2YRRqEPPxWJ8uhHHo6VlDkpUvqImQ6zjnBrMQ/pnm+2sH3vV
69D49WTV7vFT1HcLLvzznqRBfCIlqbCnqbCW8Sh1Y7qwPckzcZxZEz9FOXjfM7XEILnIRDe8BUUx
oFgFYsFHHw7RHjt/S/BMXMV0tGN3tBj+UIoEzBgfYWhFPYMgs06Z1IsMiQN5FttZVPy+DvIF7Qh0
fjzp5py8hgJabHyDaFefqz8CXCfhsTkfPo67zNOHSoQ1LS68dS4qFnqghf0DjVzcIpIMJcVmfz3i
GgNK5HbegEPm/kYrcAP60mAHbfJirBmcB+5DvVsXZN//zsYiIV5pFjQBlpDnibhv3pUHWE3c+B8+
UC2HUbshjL+j1G1/h1Dj3I/TmheLbgMca/EDn070bcXw3190X+SgxOyrXdfVa5K00G3qeN2d+/T5
pCYHeiCNXUunKEjMSKnVBeC3SVVRz8q/nO3yqThSM1JocMhCrcAmOPhjlLnpctqqgJh3q9HWkqyP
5jCw6k0dGGoAj/ODJ5m2jsx3/UZ36hx82MhZv0yoCJG9IMU05tCbKlFhMaSTRl2jDKV08hR8Ivpv
s6A0DnxmSn+8gD+v5bm85yfxr224608plgvT7/xYWAwpjIBv3DTqlF737bpSp1umnUWiMpex3XeM
DL4oQeABUwryhlVY6Ir+G2r1Vbq8iCXaYVhYT6MXDW1o6dsHJwJINUISqHcRzWxP4t1c3Lj+R2SV
Z5hKoHXEhmSbg9lqNTuoU2aCr2yrfCEruVZ/w4TcEy0PMzjytCmkJmJXhcNo5b6z3OfaYFC43OOw
erRt28545EHqX7Y+/JK430sIjd/i5d51PWG3h+9KZxrF/VPqFwL6x7UILURq/OqpRPbAzqttS29+
aCc1mxGqthPlZWxZaR5aZFB4dr5F7GK7fcnxLZ7/QzGUeVY6vb2C7j6/h0fcHedfV9a/W6kQIQeC
i0JskGAdXt0HeLZDq5OjZwIGmWFoifu3qsfo6YX+pN3ygK3R76dDLk1mppsdPpYNvOQLThS4qofP
10KOy/hkHD5IdARSxHBoyVIkXVR8n4Hnh65V9v19gQbsJ+3/jJ9+isJanbssUoqYZdaxIpnLYH1l
noUDbRLLY3f6h2f9xc8o2I7XSyCtdeKDlMQffIcC6UsY2DZZuR/T/eSUxB6HsJQAbfWMsvc8VA/T
vje8AbHRrRoXKxLWnPVCzBZAcAUBdPUOzyyzeDLLWE6WLfNxu5bQDrt3/kPcgD6/x3l483Sqq6La
SNiBxADijD1W5lhP/Q+NwPKdNOykERk4yVTLOLUZpnDpRu4tvApi05VKJ5uP5MyQd2Tizd91xry0
/PO0K8mAyfsl9xLb+7bJsHeAeVTbqR0wu3rjGCm8rGK1AyB/hr7icIPROXxXWnj/F66e0Y8dewc3
iIhcl/P5l6S10RtcMTb1q/LaDlfOyLWQ4hJbFeNcJ4cu96buQUaemeF1M0Z+JxB3epYfv/LuJxki
VziAToSqUcMUlooGDrDoYPVfQ8rTauUVQJWrZVOjvVqQEvwN6DU7Asl2RpC26UoFmavL1rlW48eR
T0GRvRCzr5kDkWoA3IVWDr6E/K6RUhorGCINThBOV9d+IvsDWac7Bg6yc6ErWeIc157fHINNauMs
+gO5PhERnNmdeUwweXmXbEXSd+Kn5a+xIah4znce0Mft/6zCIIMKLfXXHFQzDqlMYRjAgJJlB8yA
qR2IvRi7Ha31m/XKJZgZyUggSIZ+dqvukyzOt0U1vUUG0mSt8P/XZWbirPDBxac+Qw9Lw8umCfkt
+bNOMufNE99nMwSUW0+AXNzBi7gsctNNpGEoH1F54703nOTIDFz7WwOrDuE1bENRrbXAMNWvnt88
sVfLLjdMwHv/QgpykG/Mzlp8vFNykHnqg8RDZm7Vk5LiT4/BOm1Q+mV9gaab09q6K+mYSGXFIE4L
A27QVLx7fCwN7EP22rXy7paQUDUpB0A1X6p++dEerOLoIli19qeCrO7yRjS/mruTfg06ZIUPci9g
/Wn9EP9hB4wZ01lmZ3v5ueYuahvHejunyklF7o7wC5jOzcgX+Ja2JIMH+VaXuT0/Ib47F7p+ZUqb
10qOkE0A8WSk9klTRUlJuzFM61iLLAtVa1U9v+v4lYAln2Nbt1YJn8qNBfurRKrkYGMNh1eoqFmt
ni+hq+gTLIwCuK1tgqwD5tfy/eNoPQ31lkjlb0/JEggEOrwUcGd/n3yM0SSUhziciYboNyE0kNBd
/YciUsOOANcbAiwE7nEKmzCLe2e2k7YgoMzZX0XU4DjFGihI9WRz0S0qfhc8O1aGIsewKGscEveF
KJdj6jQqGE8zwCV10n8SpEEeNzbS7j9Bve+oOWGNONXH7KPfADU3UfZK47QDEwjaf5ig14i3zHX6
nlbm6o3IysEfe9g4oZ7Z71pqFsddMEoOBkP368H92pVnjxTAEo9nedAdPLAhTULfIQC7D7qAmFn2
BhpsTPGAyhNYNZPru6i798Fpkg0H0cNlS5c3EsEwcArDIruiHKbZ2F2NwEGUl0XJq52glckhT4Mn
ue60tqMyhYmhq+zfecua3ICUcJQs5EiMyEMt7XowX7idUzE9PhyOl5oYtRPoZHX56cV6dq05qdPw
1Zf6ze3X29AS5LZ3qFzzKFcbLtY0+ZqISErs/5XkBqDZ9OAm4GhIgAGCVb2Vzxpx3smz/e8Oo2WT
V4CzBcgKhwd7u2E9So7VoLY4CuwMipVkNlCec+gLwX2NYHQj0bwqnaFtP/OMz4cKwbmw8gf86mn2
aZ7ktRM+suEmmePqgbTwAKH2pYH5pyvE2moBSOIYACPcvH6+KhxJcSql9wgCcbNpAClvK07aHfyR
6YJAie36Abe7SWxicECJckjgK/iLuDsoHVCEACueFioBamvU2Cd/JSV5E/5iysArNBAHf3uzFFd9
4++1s2zOXpqfIGmDSpk6W6vG3fBymUCj972/KxFWWumZz58zndx45jsOrJ14Ov9Fh6BK0+SbnxJo
1kJLL7Xb+by/xE4lEZvxG8xzhzetxePbk4MINb9dyO2RDwp90DKeVK6W1G4regO0X6qNgAG/92wj
Vz8Kiq6JY/zU4X/0XrH9xP+pG6j4fQpfBdbbhIgIgcUs4ykmb8fCHvRagjkqXtgeEQsS582QXR9A
CHtOP8PQT//xO5NFsbZmdE3ZXfTaiHSwJWn8Aha3/s4HZVhtvL2rBgqPl2GHtdL/rG/noOUZPCdF
ZOZLdd0RkaX8dLPReQHEuq4GJaIYqTXXI87sREHBnDHjlvxxEwn7IYah+jvM+nba4nChznumO0BU
Zns6X260cssX1vUtCb8QiMwBUIWf4e+J4mcycy0GEdy1JKkz9tzef2LedrRt+rcwF+gw07MroB6k
a4vfLN+EWdwU75stnRy2ajzZuEw1CN+K09hJOObtK3Qlp4BXmaFP5wnCapH/iuGPuoGsZclVp7l5
iHJ6zJ7c4l0rsUXg749NX6sXlkWg8v1YlNFxQ5rJPHsqI9tuEW6k6YGPFoN5QF8HRSKZznfWwzjX
vFrBRNlkOEfuzFG3cyNiRnMp6UZVgOO1YYXr7dd57fng8UYLSStU60dpm5NKyFPqPxL3tPyfHpM0
yXf1WdXN9jZCdPoffo0mIkEUQuU3EohqyXoR0liozeyL8nPWK3j5eggFaVn3IHaecrLLs3t1iv1U
639TwXsD27rJk1gL85sfQmpbBVimO7aykwsdRh/ioWE8dMP6J1nw21g/CGQKaDwXQNcDv3EYL8g2
xACkz8CUA2F/NLsa6N9HqM1pmEwovJ/unQ0cElE1FDw/kegT9VfaJ0GnWI3JFF7pj9blcGWzvA6s
swkzTljK6IvxgBBNQsyr1HQQNg+ZCj2DXr5tNiKLT5XlyDjhSufSmxeaKzv9TwYUbCAVobjUqtg9
2XtF/nPFljt/I1XTliwnlkgeuEoAqOIv+AUDc2GmQndx4Y4VJ1+AsKNy7YrL1PhCJv0hx0S6m+RX
P7OhVZxXwNORPJnMWtlFY6QIOeIyi34/Wf5pRozizatWSS8J8LIzOfVuvCm14r5LT6Fc4kdCtbCt
3fJC4Vujm9zR5A2DA0eXaVTbBatRt+JdKbWYeWFopp6cxpO2vid7lGP7jdImGjDC02h4UqrmRtEF
ev2+zOwIAMEPzZVNcG5QD6SKb/nduT3hMyXGmSwN3f2Wpw9v2ibgF7sGfvyp2l0vwho4yNRjPRcp
gzgjFt8L1Yo/RKMwKVyU0Ph1H9GlKayWKKoAH47hakts+f7ND5hKY88Ah81GrOR9Fi6/AmAzfPLs
rE98D8W+tjGxAkfj3TWSY2cknvBHXSefjHj3P5gwzCrPI7ofx5dfdwI/5HnzrgEooIRETG0aibWE
a4ZUmj0mH6Zl/M7kFhbukgjVLbSnxPgE/PG2JEsKDF/15XSMw6t1sIh/xIQgZzn5+JUo6shUxgIz
DLty5IfiAplKKW8nJWk+YrUfEPaluHLop36hnV15rsH5/zAI7kTWx6Y7tw2JXcZlSUzP+43PqasU
unTvhhmjBd4QbUUWfRfNzq7R0BZN1qOcTVCHtqT5EsvFv7TG4fI/WFr7VICCw+BIxtTA95LDF9b5
3X0T3Gf+IfJul0woMTDncT+ceBW2r2+Slgogxwk7AYkdyPX2sY4FeOeFDKUkGjYt1TKq4bUA3QAE
V1A9QZU52o6M92GMBaezaGF/tdAA6bUvRAB2Fls4UoWtmfd4Bb+jGP3TQ6Mwuti7MYdHTPfxmNB3
pxyJwgnigM2lkFHbfED2zYEQSEkJvnYpmYMgrl2XNBAc7HpFyNIQveSJkEtFJ7qhqR+N5+0r6Bk0
1wFaArrdVH8OIkd9lCeIrJ1K+T3DRVOmzqKlWngUdIiPrG8LHu4a965GyoNdj875W1rEpMwP1+uv
URGXdlz8JAFudSOBO0J22HMi/yIEXTSEr30aypyIMi8LqO+dRqjuU+AuviVjxyHFt5xIt5Fw0Clw
tjkJI6CHLETYnAvZMGpmo7TJ75ZMYWE4g3C45/433Pg5rscKzuJWnYvLyMC2Y1LJHz0x0JV4mx4O
HNy3XSXGUuiENj6ZPcmzUIPSGAdUCip57D+l7vqpbNfHEWZuYKO86i8nKe5HD0KgOF7QjrH0sVno
TdaNTvC8/KEmyKO3mWT3tSGQDfbYpXAPF27qznK5DyDj50rRB1qAXQ0+ScToRsTMYQ6qNmYJ3Dr0
5DoyWaiHo2I03MkzEuJ7WmUr+MV/UaFaEpoIjnDt89eEt4h82Hlfb6+TwkEN3Na+x6uf/qlbXW5g
arDX9vTbetJdW+M431spSpYrxetuqa4+vYvZzV/d+8pWMNGHtRY0AMpj7tFDCx7wRhVjJT8iSVGG
yOj1tx7v9T+taq0Uu+jGhBl/jy4CBCEtS0L/WJndEU1evAjGOFQyqnZNH8Wj4GQ3SNW1Gf9/knqP
lIA75X47vT9PMSYD4hJaTkG4NdZL/3qRevZLO2ch2KyPJD7D/cQ4ju1GJE/VTs+teYO4Axe40Ua2
UP9PWTKKmqxaCaoe1b1YA1HaxkW3LSzA0ln7LTvL/KP+QKaL2bOaoeFHoDyj6+SaigmBbSBOYei9
7+Bbgu9HeTuCfjM/JC1CSclWX2XLDCka1kw+eOhtHNaCVzLdhjFTSkxUiFmIU7tfvOej/iJPG+0d
O/Fw75kj1Y/s9C4D0aXPkZZk/dwzvkn+rIibztXxR3qojnRx/lBZXMglcX0ZHbw4mhCxkLOTptx+
eNcL7otwjioL4tjAamsSdITFjPZfB7d7k2Yuw0jhXTRSwe8OS7ca3BPOEpvlEaUTMqk7A1EoEhpz
rES/M002wTZTIRYciNYZHJb2svVIYA9sccImtxZlOnHqiPvBCTGwEokYz54PEMHjMef00nPnqVRq
DbC1kwaqWAZx0kIUpiCc5oSudREVvxPYsg1qc+LCYprnZPRBGn/CIPgwvVuEoQIdqJc3tTBNFkpC
h25Fiq+b9HFjr5m4HlAU3+lJg5DTlFG+WtPm8j3QSa5ZDBktjnk0d84XBuwiZ0cStmmu+R183yAI
lBGZof2krjKZBUgPDS8SKV2ByYgl9259Tz5+zZzPVuAUYPPpWdtrnVnZiQXZNY7Qe+gBOCcYCRuz
JHAnebGRKElp65st59WPPqUFFCgy2LxjjUgAv8ttizWNMeZZxDCB/Wb6iHSSg+Gi0gPfaQzISFaK
V9WiPZChxIlst3VhLl8QAeRMVfmITn5T4/l7z+rYxIDLGpcxWMQYwHa+mm6JWXVzTCF/zl99PaXj
DK5buoBG+pjK2FEGIr72Sn95O+qBJl4btH76gLKzAccyXp5i8Le83ek0TV0FW9ad7k5La9Lpta6O
SeFQUswRXwP90/0X1HUZtt2OJglfP75tsswNXQYnrA+YuY0ZJOS/5pYegBdxAhJi7PGpFPagD0uI
P6Kwnk95/JGLUprlDbb/nwNRDeKQCh70wDP61p/mhgv2+uxyllnAjlRv9petHAipsJZcfy8PKkm0
jRsxPypQ502/fGLcqBLwDD2ocd7RSNNqbHYyD1qGqsD7hOvi1kowbFWN6xIeDsnNmt85fQCkfbQ1
ND9pO63wmmKMVmJp7YE1Yl3m+evZvAWQqt8ttj4OxcBdMykkpPlfIgWDBMKt7pM0tHBRuTZ8WAeN
m/+jnQBsngm1V98Eo8UBkxpLHMRSTqSZHCTUSVthnd3Jz16NI0HOHnFvrPBbeZzHD3NwvqjP7zGw
Y4uRMLgDNwt3dUDXobw934xxOJVLu4ydnPmWHNDvU2CQCW0Uxurrm8rndazYjlRlJcSk7Z9qmFWB
crkmjVOaqgGh8RRIVbINwagxhr6IoexhgwinAAf+g3fW5VoeHkZ4WR3yzjORLsWILrYf9mReMLFA
WOCNZUEY+TcVe/8EpKdBt7JdNqqSPJ2Fh3IUr6IPb/ksN9JWu+jbhFXTJbWAwEmRyg4KBLnZl/l6
dLvbfdzefU2Fi67bCn+r289nak+bA7eEyPo31YzBUiHrMM2zrJLFn64LtDOySPT5fmtm53ftikaV
jd8V5dyV7HHhCRaDT9EHB7eLiFJz+YtpqlsVd0micDY9ej4h663jt0L4ElPqy66i+5lyLduo5jof
OLt1fP9jqnX67zBF1t9XumA+o5X7QDV/jqVMg8eXgP6dCIcGwS7g4Ws6n5wk3XKk3uCDG3aSaHCP
t/JoAJKz0G6yo1wRnR/RI/XN/sFVihElolmE9AUoaBxdCShBTHFVSSBkTAWwb6ibB6Jsyq9prgDD
wE5l8XYquuMS6Q6tfnC7qDXea4gUSp9GNbfpxhs8MSsiSSbgA2wumi48mWofryT/m9TzxNCe5TX7
oGeeSUEpBEilntYKVtuPeT1tuGSvSZlEeGagbYZxqjolJsgXpbKFs6O/uMm/dz2IJSFdlR6yJH46
+GCYlZPF4YEepcKS+HOiXCpZFsn94FsdmFMjkYE2mlbTap5b3Ri/LYtwhyGRga8LV3EXHtbo4RRP
uurZhfzTrQjuBSfPyu21SZMldcL5+VIQBFcfj5H1yw4kMgSs2SLdQWRYcs7W07bn016R1O+eys2q
yIRHfYWCEwR/T5d2fLaqPdkeFgky2plEKTNJkYcwg6AppiPNNUAgtKq/iAoButCnXP1l1Ou7cKdn
Vgvyv50nNu+MjwJrGW/35FiBBNLLPXBUHvDxd2OCtmoeVC2WMM+PISYk0CbUlzR1+qJLfRR6j6Yv
lt3cNYWHVc8P/RnF05htGOl8ds313o3s9YAmLKERWFtawoChuHR7BFLm4MoZBS86Ju6jO+nN9wQx
AnkjSG6eslV+rhhAJmyK8VbZKWPTV9wQm2fuQ5Orsxv+jvxhdSoUhPBJnP69AN+bZYD2QxxhZybQ
fSzIDiZpYlQLC1o80lIw5YogxoOsZ11Iql6HB/rUszWT4o8Yhz1RhvXT489g38Nz05q1WNZjXnaS
CESzEr/upALKsjLpkg7QQCE7QYqEP1SWkUILGNd7AB8JK7+JZaa9mip5R3Ot4immzdlJjYHKb+E0
6fFSWT4zegZUP0krAGnlPWfmoFofCJy4pAmE7FUop1cKk+7+NP2I75gJ4p7Av2iyaPttPa7B2ltM
j0llU+A+7TmkSc8jG5YMB4SCY6phVDrW9JIPgkkYc1paHhv488cusk03gDb9+xD3xq4dBdBlnNyX
RSHANF5V7O1NcyCAKSB8LULGGCaE0bcwFqtjU6hHgPhEm2rY3DcRqE7l+DpMx+MMVrhTxiBA2Jsr
+eOIntZNBQbKWItJ3rICxwlexakZBYURFMNNREtXadGf1Axzr6TuM89sj1klrTXDNKdvRJWxDHnL
A+GafS+Fuz2Mbl/+vC0LXV+63VQpB1fIrPX0Prl4mqyTKN4UtY1l8yd3Aaa4u3BhrB5aCIwHLYQ1
pAqWP3SkWyO8jaIAqKhDQtJtNhanbzVsCYfx4gSI/u+lLRjBq7LfSu79ZQniIeE7yLhMbcXeK2fA
kOuVCmQ+THBlI6VbHTIKC/sXpgDD8+8nZdDU7FWhDTAXzAqroDOKU+xrOZcy0LWq/i5LuD24SqKB
qx7epBTWPxH7JUSMyWS+3VlXTiMpOwMsrprHV//0t6/KPNUBdvUOcKWx16kqt6+OZ/cl+zpYnUm6
vm2yd3zMt71NHEoi5CfgFwuEIZXxxWCvy7TEUrVaYCZR3BZYuVdKmWoKPIi9pA1aBZcVpSLMGOXL
PYiT3p0gisgpzqNutXyFWQQSL6IIlc+sL/hO+AkyemCc7p1Az3CRiIOxykj7zewJ2w4HysiWChJi
sWitAzljMax/Dq+g32St0uegL+cUAxirZbxgUTzK5No007caaFpgXT08WfwaIsH7LhLmfM8KOigw
sEbGWHu4spw8eXCznLDWTcceVGDUfXpCcE74tYsQmwU4dHphA3JAEg56aHiYVzEfVCwGHbKULhuc
1dit5Urh47X0NZIClmgebetB4rIIEiwvsMIOSBSaul+juPS8uY289drL9bfThoJ6SrkvKIi61jTh
sdOntSkLfaXKWeQ1En5oAdXhR2nbl4fVAc18BxNuqOWeeX1fmfE2D8Bs3Q31bQ3zRoREjepvSDEy
tw5O7v/ZZhvP5IVkMFzuAuCneOXv/xI1xNGg1J52LjRELb2NpfF+2vvzEeyN8TLP5f/OkX1Ig0KO
3eTXh6CnMfnqgx/mvfQ2aLbuVPxIkU5OYByW8s1BR23fn5+NKY0pL3s0kogLjPrVmI8bKLSP7dXk
alx2280s0tPx+zCN+Eks9d+o2RZKBaNZYkF0elHwb2hwnH3qbnl1vRqgwRV3za4szMnxWJGYSaRl
XXXTboGYGfHMud9sKrO0gh9sQMOHLxFoaY9JKG0BqiBi+7hGExTcmVxCQ7G0DHZeZ/OCcGIZa6Rr
KEGRuIPOc3C0LYHfLw4w+TwwKbBJfHdcTuxmzRG5sNeVQ6cThVHi17tMX+9Lrk0X+GceyGFaAwjq
lZYs1PwT7jqsMpQ+lcaziCeVE9vxf6tbzroo6CIo5i2SVwq7kXeoFxUl6/5Wen3ChhRxw5LRv5WE
0HnbXlQ1wTOF1APB0+Pxe6FNKax4IBplXYjxjUFIjCycvgnI+KAeFRrdL/SiYjAWEUOc90FwLZFC
saemVCaPUTQ1rKiZIfz7yBTOtHKnYsKXUtS1NgXZjKlnuHjQbbMZ5Z77+36wyHP7eweWe4FR3kx4
BNaVaSzubHLBwFV/KFyIy5XcHnKEftK68Oq9+6eXA4+sWG6HIUHobxa07c9rJqIpnHqarliPJwaO
b6Oaxp1qiaX09t7DhJYTo0P4EIh2p6mlIuqWz7Em2QPTju6Nue12uGp/f7QXRmzV1wZGVtwEYB1H
8zrO43dLbzdaa5r8stfXv2bZ/biOFDyX5f9g2ZBuzEhe5rGxhNNsBDlodgT4BNj1wuD6GA3GlTMi
WS6u2SQgfrBunKq+NGn14DFKH3RNTo/llnNUeaxwmvAL/Y09taxB26c2qKJGXicfcNXvWvbWaPdn
DX+764HqBdSOdvUGrSIB4vbOUwCENkxgIi8QDywQJhA2XNbzGzIH7uNp8CYCPktbPDeZhtKCd1wS
xLztladWCV6HhN9KLjht0YurhHGZWb0FA/xdw0+sSQl4jChDqr3/Kksp7L+gqf7mDzAOVoyBLHHr
FjfHr5Et+N48kPkZ0HH9Ifzif5VmXBBbKZySI7jd5HLB/Pl+VSCCY4kX/39eakILAqfAl0CEEruT
ne+wAa/bA6Z8KfMsw8OVlJG43oOTuQYek5LmH62zzPRG1BY/fSxSBXjC4SRP4GQ+mIA7ip9g0LaO
lnRx7OS1syTblm/JkB4QvVaE9ubtDCykQpIixnW5O1qdnxO8KkSsTyFfdXhoPxK2ZQoA/Vg557O8
/o1cE47nieTp6/z4InbeZVJV4GNa6Dd7eosaZMEKZQMQsIGfbzQfS0MnF7hvwr5T1rpAV73EJYR4
r/QDqjZmnoYmoAKLqncyTIUmHnGeB6J6yXmtyfaH0RJ53hAfy0Dx748DK8JKej4gakCqU7EtozY6
xHH5oftdDNXRZhGWpoGgVHF8hnk4digw5QPY8KyNDUYJfWa3d4VI7FtSTlZDcGhpv9w4MIpxyeKO
IAhkXs9OcwPu+ndHzCiadk/Iw1xtnMlUapXsCeSaWW91h5NwYKhywSeyejjcxUuJUIP30eWA0LTR
db6qWM3SHdajwKRHG/L/IGxR1TItMtOUxqa+oSYV5ZL0mdV4uKhnZQL7/TaZRXvZEKkF9wp+V27b
8wh/p+PKo3l1mphq8RO/gMVZZp+giBWy4fOFYulK5zXvbfbncxJZ4kSEMR0x/knbGA9LQJGyWU9W
tDtCpY4wZtudcUeNno6gsKf8LbV9932gHxTBxoFV9NijcAZ58VgigeJO0VQfGKn1nwdDX21tkb8O
TDSfQnaDiJscj8exHFmdIuaqq5qtggHX0vC77AuFDEMFpIF9sUUl/GpYe/TJ3K4azS9GqYwAVOlE
vWMWWboHFcISKofkJPlUR4mnnKGzBDgBCM9EHm/FxY7or+w/tIy6cVdR/Ytlr2AivIo/ozNqIZTT
WJwFAiJWFBC8HQVSbgWq9WFGZA500gXSTwu30cT/JL5k5MdsaxWJA+75E7Yvx9KJBq3602ho6oIc
RFqIvgiIaoUcXOcm6FgrFFGBUmOErw1IztcVFtOhIwsUFH6I/9jtYHzZ2W2Ot4gSuFSwW+rmOX9v
CALcEFnZXgOTQnVIdwJ4HQb/MfHNdolT1yyYgn0ZGwHWC0bOukDpw2fL9PTYUWYLL/Frd2QDRWSj
Mvj8dhvmVVye6apoW7hX7V6GbZd2eNSiQLJ+4s8RP3D9PsKCpKxF/tTglI1gnLes5Cl3187c+cY9
M7M0SFY42zDG4MufL/iIT8Rl24S/CsTGkBb2nxv//RKRy7zGafBBrg5wIfB8sXCCelpi1pWv7sui
wVAnAeU70rhjAEM3gG9TGuEj4T1vyF/QMow+E3K/ppXn+eb/SaePAWq8kGdhha3qCVuX+s5V2aZD
YdmfxSIew6PSIg2h42NHyIPJad1oyOaUVYM8V21LHIVq2kWyrVdqzmHVeBDmQOHNFzW4diuRvZeo
pdKVNjs7EIlCWdXiZiAYFkd3lRgm+0RUgjzJ3K1qzVFK4tweDi88RxdVgNqqQMncPjRsxZqdT00u
7mCzlQNMHn6lS5zKfcZbetzKjfnqRlQA8H8aYlsMLpLvB+nxcSF85AEZU789cXVVw0yYgfGQ9enD
015SqZD0j+2Nc81HyVeoycOwHWuNiBeGPQQ/D+4TGGZLzfn0ExnbTlcEg587d38fjQy7bBPyYpa8
wyberLeJ6bnvFI+Qgtwd8PykvFTpIKUeFJGWweG3NGjZ9ZhEbeqYyKR5IINz49Qrjt8mAB/904vo
CeHCTBKsJF4BO3Ey1gn4OXfXaIwrSvpimsCrYCnEFFBrXsLS45vFym0ge9FS602F3GID8EmesDob
Bs/3Bag/58VX0J+e+eoO9NbCKpRU1vBea41KaL0iirusPmRDgthNu0+QD17Ku511KVdvsjaYE2UI
3M2TP7AGUA4HHRaOs6K8ad/3blt+HW0v9AdntNUj6FueIJF72TNDc16q3UbM6gha4i3BViCi9im4
bDoQqCDH67vy0/9zyUP5tgJ9ARQVFlrJS7VUSrNH0l+VeynPxbrT3opo5/HsfGvL7B5jo5N6yia4
btAreLENG8VR6V0ZRJ56T0JBaiU264YOhKZUmvgy3BiRNiLmuD2pQYWciSrx496p5B4Ym25/B5VE
HKME5ojMpVzUkLquztamCDbmDfmyWF8pfMCq9jj5lNBlnLTTq4wQnPL730HIAosP7XMzVmdxZhQD
3ErUBst+2I59OM3uvkD6lduP1q5MqmB7HYJQCFLkNvXGibp3iPwaNOTvJRiYqIcz5WWQ0oo0oNRj
WujAT6p4ZpQtUaJaGqpznbQSeIUDbD8j4AMW55sF0g/qBys+9hQXLe2E5zYvioCh61gloHn3IbeD
rEVxbxFVDbpJhUKHv5HLM/mnphG7lepi7LBHgrtCnf415jIiwNVPkJibsV5kYhrMW4UL4qe0X/Lf
7k9q1DYnHU1FRJ5chq9tE0GHhw6zsArX3iVoDOUWgyhu72MwudKh4AKtUbAvWgXyaadmb1M41mD7
HP0oC+zgUKMnNHRLWXl3w6bZnm9H5IpVbEfRq2JyavzsiqWhHcl1Jk85L+PoQBJEHNaZJBeO0Bwv
Nt+wqd0uAmK37arzLglfVei9bhST/TBugEBmkBEwAvCF60iaIXOF7oCAnToM3lD1wTWXDW5VaD88
mMV/QMTspyXpIT2ozg2+1Ab6/7Q1njEarLXONnTpNnW9YQvbm5DSNLlMuWBN0I8TZwD/QgFmQ6IZ
r1iUF/hGxOx+iaSC+qGwmfBX8gBeLZ+RP/4y5tKC3ED5s/W+Grs7FL+jSyO31P6SVVSnPs7A/4rk
kq2nhaFWjnXVX6H9HuBE/G2apr1SvjYluVLDiY2swoQtFcLFytp2QKgAk5eh0V031URGzS+WlFSS
nBfyRsXvnV1KZ3EOZ62XaKR92DXctJ/KhlVmORPKWl7ft1L0ULQOx+Dp/h640O9U1J7uxQKVHhkj
RKssmUlq8EFXRXGf6pHVhy1+FTOeOyrdZkwHZPOY9zG+4xqy3cm2zQwga71mi4mAsW5Y3j1ZY66e
GIpiZL3yf+UDk51/AJaW8vwwodl3+ec9EZCbjh8bnDe9idl6sqXkP2fxhxLlc6nRiD/gnHmBEe2D
x+L2cIok/oRO1Q03AZx/uNBsRjinzpzKbP/2xClUvrMYcx+Cz+yzBJ9LbDEVX6HnQxI/fCI8GXb1
VmeYCKqTqTQ5oDpehjBdzdYUAa5wB2fIqld1Cl8GIGt2BmA0UknbIi+9OqAvS0sPqPZ07iSBL9cp
vOJue5lcolw74HNJh8Q2Ifm8D7sPlk8svpyftWGG6KGcWP7dar7ldd+BzFtKrr1obrd4PsJEbxEu
7mEdt5Kx+nHpNXyKlAtWWWHL0EFkcmbfKLdDQABxFvLdc9y+BS5ryNap33gA8Q8xMUrx8KLu+jgS
fCq1wvU1u54+u9JqU6hrS/5RYZnLFtvGtTRPLh0InoBBB70VgDmyf8A1G+ZNpS7sUHwoL5m5JA8f
icwnZI2k4w/gU3JVHGBCYKQOx26BLYImzefU4bDeCNTRTQL1v8V457CFV3zz9ygcG5RBAvPXrali
wVJovWEEtYxkDrs9oz9J/T8r9KtF7DE8BeqVxzsQA/SQCP3Pu1uik4Xb4hNS2eE8Lt9yuTf9pBUh
FNQvHjM42KMhC2GbLEwwLrbC9EgCQrOZ+xdUeu1VAc4IcNDB0yZT7i9FZ16vkZi+pFGV/+xlTiLT
YqSO13nzFn1m9qyDnwzOrnLAUki8vSkssvpn3y7ZZVJWAJonGEFWIWYw5at34/fPVHS5mm/ALMqg
z32Ds4c+fdJ6STThhMcPSNSVPvIresZyb7gxOZIKYc6/NOGYbgy6hW3X/SWsXopvbrwVwZHp4wAE
73bufXy6mT8VbAUJidtpitQ49KjLRlEZ8yxwM21DCmQlZ3t2GELW06iNVsS4+B5Wopa/MC7+cTU9
oEZkafnC9qFL4TkDr6olkpNLlsHEYAQTJ2HSEphCMSa+vSmJtMrnyz3atai430sDdkPA8kxK9R4i
ljvldbKj0srg/KQwH7f4OQMPqTqlXPvnPGJZqNmSdY8s7k2tRMY0ShYoeR4vVL/silSFrJhN2LA7
2xk2buTquIUk21LB1v4DkQGIfQ76bMzrHLYN5MnGOQt7B2ync3XFYFq+mK+8qNtp7Kq9yewm8oTi
aOGZjt38QFisZH/3mLCFHbvWy+oRHxfY9njEhNapYpvezwFAB25xWzG9IwJMRiDB6H/f8GXiIvIW
FrRujwWc6221OEQNEX45/kSRIFrPRHX+WOdZYGX4A+f6chzyXIWlsbRKKbHn1zXxnxazu67IzlPv
YALQ9fLHv8YgfMoBE7dLOvsMQ8686KDWqs8lz1FCX4jHV8r1i8IrGOAoiJgCkKJPccPsYGJEkUno
uv06rterZd+Y/yGZkwx+IAoqJtQ/xGg01yeWQa1blWg3pIGO6xO6VoG8ebgKSB3+wy28/K2dZh2a
MlHocKDTApgVtqdBEYNcNSkWaAlvIb/sTcR2V8VfSLNMvF6Y935jNuOhUYhyq4nRbED90owcfNkP
YbrL0xVD+n4ERP4uweBEJv3pAueCwCY/1h2CvPcQjtVs7J/AAkbqTg3D0PG8EkEenfWheT9YYOxy
SREGbo13AFzDOyc+R8ExeudVMhb2aPqmOdzOewzhAd2DAVvlmNjY7mrcP1Mlg2sGmrGBPA+3RorE
G+db/YSOxDCYOCQlzzUfymjf3CG4e00YyHbz7JNgkGwyg6Q4GEq64cHyqJ5e5b/PgiHJ5+4afVCj
TmtMB85sljQnxGQEtJ6H5a36ng9rPlsPxPNhSFlsX2pLX4u2XODSK1imx+wCcpfee3vvo6b9W+23
51X0JCoJ1cZJgymNjxVAumni8L3DTNErnkVfMmanETZSNliIyBtEldegmbYvBAD0rCkKfPsOepyJ
+TVOLAGFjbZRiEZYGLrypWCpVFwG5rp01KMIcKkshT1wvfLpiz9BAf9BGkaoQ5RVxd7yd4sgAab5
vsWBczG5W0fd+PouRFJO3zv0sCm/YNh+CMxUqQPONKwmR13CPjvJlHYRDraXtVqnLY6X299pBFl0
27uPlzYR/ejLZC8nOUp3zXAVj0eHLpPHraNH4bWg7fpAUUTiNCJb68y6MbqjkDRvmsI+6QwpL4nt
46cdL1A+ORc8pe6UtLrnOeQ8Kzkumpl1KGdNnHfcU03EghNn5oMDnq7nxI1mgxjL1+/nzBuscKLA
xaxz3HW0w6cFeHXvsudeMHbYqPrsNzu82hr1pV8RBDXF2O/Rr7iGDN/DCL9bVyG906xpmhX8PImt
TTntHGK14OBclxx8ShxjcPQR2V4w9/zhrwSvD+bBnGqqXc8CoP6jK/D6xaEX2LT22VuYSab8JDeY
qE/qvTtZzSK0hnEfpZq6SKsbfb+tPOu/S/S4OHQfD4aFdexh3/HkH35uoZ/EmuyQbUOEVZaGb9yq
D5S4XwKTZJ7LDYj4er1NV8SdKjv7rndh4OJs8Jo9j8pTBNfuFddtOqDelNf4D6escpFCu0bEshe8
wRCi3lO9rlwuQia4/Df14gySDEOWjkO5f575ePmhSkNI6Xd7XVWDvRPClvQ8LftwpXkwsLtLraD5
IPHRn8xurHlz83oHGHBMJjw4pqIh92twtBHMw7lr8LOT75c3vFIPystgdU7GuQPNJIZbg+sJIprD
IZJ9R7BHTOBxF27y9AfSh47eIjEdQuKPQrcRqvC9/kCuYy0XqrKaoT1wJWwgaUT384KTXsvkeqqz
nyizTcEjypLjGxJBo09BIvaKn43JCtJ3vkgVk40V7WLZcYiwmuGJbHkzBRdIhTy9oaOgsugzqI6R
1tN3TdxIq/ctD23Id4MKGvhwdzph5xRNcs5IQtftQKy8L+3fiOK/nwJ5xnoOiGi1KhmyuCU8VvBk
2zJbfCZfRKEAfQGx0iuSPvm+QPs9tzfgAv97RFpRn4jgmexL3LoZyzBxzzt4SwpdQdHB/7uunnEF
PY9MJn3QFsa88vaFTzJzmtZ6D24ZCcnd9hcm9Pem2xmtl9N6zBYMqoXg2wjdJBFIbE8Y4kXDbdfX
hRxJ8gSvovy+mB3X9cA3dv4uukXXQ3F9+bc8Gfg7TypWnEcBlCbR1dgJi/hzrNCdlqE2aWfyyY7M
VBRDBDa6Nr/+kYKsj1rvbFDBS63ECkp9FRx37nxFqoM4POysofBqtISxPMpWZbGBO5XI4/77e7D/
wz1kZpF2iYqCKkXewuGI6lPRohGH5N5ZC6YQ3xy3Ck3OVLqNfn1SURHwNRRRIo0nPuUrXArIwizf
22m2xDaa42Uv/lPlKktz2ZHwDngSQp25ydju+E5raX59Mm0tGNpothFwngdqv6u8B9S3tfFfZdnV
pUyxLIN5LyS+pwkXdYrxOY5EAdCQc2hcT97liPnkCMptWQI2l7F1rtD/5RhQbVzNdbsYU7v7tJKa
vf+av7gx+DkDIOl6AVij8RxIph3Blt5flz5CVDv4dSOLuZp37q7nmUiiFC4suAMMRcGdoNIaWA63
wMqcyS5jcHhGmWD3vsIUmy3aQITk0smnhcb5I5TsbM0s27+2GVNOSbUFy6uzipF7CfroirzdKroh
hRMy29v6SsDXFvVQ0YHoOrDcHqGQ/xJGLu6FxDDD/1aJDJ8OWWwJLOTTlyRDTib0bx3MnxXESRRx
4udzXA0jTl8RaK9LEb5gKFzxaFYKHAPGrHHhzQ/yMueulUYsYpV+nKjbw4vLbcGWC3LYxjX7WAlz
Z8bFCb6jkmY405HdsKQrnJxtu6N/ulClbR1RWlgexbwtvDnIXgkCwwXDHyBRgLKRuLnigAKGJnEn
tQWyLWcdWoDL54ZiBzh2IevuwvLQo1D8v7niLOsm3NgLBHKrkrFnNHTuoTyoiNUYTcphEiYHVc/s
xg9n1G0yimz+tulVY80EEMV4TtuVenWbQWTRpyeRJalwWRlw8AI/bg+NeF5ehPvxQ0gUJBhx43jh
hrQUKKz/bX6nhcKvDuVFBE+OvCc2KRkC4AFc4gxfqChmRjZTP5uuAw8hYSguwMbG72Dd9NjDpnUk
CP2KCUkkG6s0dVP7lK0PjbSjTgK9Clu/ovSNn9B8peZfnYuY6agEq9NjTEMmm4iYv2VfM7fFEx55
V6kQIkc8GoK+qoGoOizfZy1J4MBQo/DCkZk3vl9+mTtuimp157zl3esU6MptZnCIgSJCQfhHSuKe
0j2EZos96vsNlmk7UL7TolF6e/AqpYBH/HIwt9lvDf8UGdE0t0/SJ9F37/0vbPYx50oh9e2B0cpn
fEyOstczTmoxAWCPZP9pgQikxSnsmsLb53MIlSvekXS2WJP02TEOaYMwQ6/Ls7dvAyxp2tKTx4Vu
5fQS/CSiq2nbIpIyjZe7BwdUUvuKcTPUlx8nSpYhJMzYez7oTsoBFOn2gDOcu6Tpj6DMrROlyjsk
YcstkwfjQh3H1EFub+YAxwIlHPfsH9O4gMHkSV2JI/IAsWjNcjudjDfA9HUtzy/MCyn3peuVKuI0
K1rtTXpPj/OWWU4uID0vJbPFjzA3fyGFNDCqI/tp9nIsQ6xCP37HMr04A5P6klnGDjsW3wtxAPFn
wI/v0Eotbngm8r4WYBc2NnjEgMyFiMOXLFGFYJuzYGRUa6Y9xEKKiHJVsNtDZ25NGOgm3dulGEe0
yYRU6V6UVwTi65aUj3p6lcBNX5u8k+kqSOJsCjyYDo4j0EFP9iluKOOuQGsIB6VSzHIB4iFAf/Ei
io9CmHZL7SyDcNLmSQPXNKJeuf/M1Vu5dLQATNtRXBOD1lj8VDXGTy54JcjwDZOvr006uP9HDXh9
HqGEZqE+Y7b+Xn//k3BmKc+miB2NsCT5+gD0rpk2BD0jak6F9r2TK7o6IHeL/D77Rd0yZVl8b4DI
w93dM0ZnVU//ZDtxbBKXBfvFG1CvJDmgDNociZ5WFiDRC4htE12/dHDGY0M4z8t/lBG7BlaP8Ptp
2BqD7uFxu8TkiAzITx7F8rsSkhluegSKhLDHyGsq1GxKIl4k7IzNShDTcVDh2YMvmbuvgk80Pi88
QO83mi8+oIiB41mSIJ82IcI1XLPORICEcLf4X0CNYbFDP1H0NQsajhQwXHSc1YvcOiMAkciS0QQY
tN7g1gV1Dgp+GWe13U6mRv8/JrL9Zly6zhFS7iX1CLaUXOaEAR5m4FlrVJmX86TMiRY2qV5DAh3z
kUABkxTnlCjNI/p3xUAH2sISbhRlj87KHKd/Cg2Zf5Lj7CVvGrF5YiSuOXpKkleQuCNWbDjl2zBd
ovHah7N86ffQFveAZBCmhrWY46IwaZoj2iWpDn+cm8+WgsgLR+BNLx+zb65ES6Cwu5f2EgCFGASA
tEWX8NKt1vZZk4Quk+VdTn1KzdcO/ytsul+rKkGeY+hhQzrZGzf2pNh7Bj/Gc98VpSRRRwdteuXm
oTtvR4uBIvieMgqxfvxvZjcpSNcbz6DYQpKwq4nqhrjpRrKJyLC9PuGoJI+o+0nAUeSpQIAcHbE1
Xiou/zoaQk5Dlb7vyyxzWCV2/5CEFzOM14HZIbYUtTRL8IUdxcHRyjbOm8lu9BVA/nQGL3cnM81x
ccZDp4fmflKj/KbKhIBJAZLDIohpvoEhL1dxFNIpIYQPuLclH388ioATWsqyvxZK34tHnF9r16dZ
fBNayh6zcND2MUIVrVSxv+rtEABaSoa5E4lYWJ812ZoBZPU4ZCo9vY/2JXlSilkL+AaX10KaUVgS
Id4e4Y7C7FI4aGbenS1cj+fOl7H99I8oHf7gPRO9c6bIN6vbEJC/hJJitCw/yGu0WPucgJINXRFX
rOv7zTp+H185kFN8smNT7cpeuiuhCYj1HB2SxvrxkmRiRTSGe1VPG0aeEiKvwXWF8tCI+tCeF1JO
ogWUQ183XyCSaaEuEQ1V1xLdMbC70Tdlj+lM3K+mJZMdo9pAWdvzX8WULwWB8MWcnXTQNtqCJW7H
c/YMpfbYi+UQq6rFBWWUxL18pxhEPXBal8+ZdvCVCEvNvItJNVwNtjELfTq9Nz0IauFBsXXoyUlM
vOwDSIK3s0hkzpblzzmVRf+sOkza2k36OqcEnIUha2kmN7uTAME3FZc4u2gGInfLrJlwIXniRPuM
kho97qBbCdsfyhU4qZoK/qVUgc1dfgLwCdRqyw2ZcfzW4jzt7/wPYAyLMJ97ImkyV6lif2HiAnGc
2+H6Da/BssCTy1xA5VXnhNhtZlAwv/Dw4LNL4B0pqz5ZUwjzdErpBf5/bH15ChRMvXk6dXuHS55T
7VAmbcJt576wRRg3Go0QcTG4V//XMRqJ76YjSkvRTI0WgxpcwMtTJIDXxU/ZOpyTikmrzpHXmCN1
P9BVIU+unpxg1LcOE6vdCdaEa+T0oTQNF7uzVL9EnexrgiHVJEIi/6ldxQ/q+TGwx16oVn/2kfat
XhLzEv/r9H3RndCIjZ7SBR4WvU8NBrGXGwzRmeVmpngsNJWQrG0jrMsIz43k3ya1RWo69WAFHaqd
AqBY9tRktg1pGZRxjlN+mFouPzc3QIMfwXi0jc85/a/mt5OzuSwRhX9JSc2dbgK+mdFb0+YaqBjt
osIjHvIaZylylmjkQ14IM5EvGiot4lfk5KqPNIH4V2GpmxbPv0VmDQ4YWvs+JvAkUijz0iH5xBxz
VTj+8yZaW78PeY7ezInmXKa19WizqGKqJZL4mIxNjDvCM5qcVCIoTK33XsZv3IcYtj0+rn0mTjJE
OiJOrDMYR8YONaXiKyOG2SVTYXmnOIVXZd746Ik8TPQCmGx3Ab46Ckprn84TG5e3JIddSEX3EMCg
kQMhpjTIVxn/pRd/mQRWIM/P5VyZznT7fctRJLMVTtJogZyUxGsmOqsIsc64ogWgc0lezY6+Y8YX
IcIplY2vJK1r1coVeEMoVi1GrAw0LT3E/oLpFxWWQEl+2PiXwZ/Ta/VL+tMsrGg8eGoTbD/TASCm
OWOmfahOdmqxeERf+CRzk2NfEtlSFiH11nWnza1BRpQL3sKf9xxejQfLb85JKsdSugawYYCZxesa
/MBZoiYBHRBBWXa7lSyRsN70NMR+YuLVeTq+22zlYet+wZaAIrAHArDFJN3OVLcoGPmr+qBEkOxb
UZHrnOxszinusqEp6KfZbRDsqir13wC6KH5b7PBcby0vEnqZNWiimLk48kdRWkcB+xwy5wQD6jbJ
t7iLPzVEbZwlgIqvQbOrgfP04s8gulJknmH29rORvZRPmdQI81pBL0IUTbnhvICRSqjFat6LA5xN
4P6MqSfe3OZxHgtmp7qbtGka/8FUbC6sEKaMIVAZtbEn7TbuebM9yUftzplaQOxiAASkUrTCjoYE
NccZgF//MjeXaeo9Eady5GnXToX6/d5F+E8L2hbX7FW8ltdt3k73pxTe+B1zn2QbumwzQ1V/HlPX
Bd3PaUuv04VmDxhLv2Umy4ZoE+bQfU2bz1xFtD2EIxqNiDREQbIK3JekRgMzkkvxxFkNv+ElgTod
Yg3+blht11bWceS8/t2L9O83t0yu7sB++Z5tBwQcxKn5U9YTcQJboJ23EEfigCJUtlkqdQrkcDij
dmDGqxeNDAs+RyWb609cE2oFKF15aKlDAwwOvTQCnBWJY94WtWPQgT5PXew7qhTTYzB3nYN/EohV
7gfQiDf9V5NI5UiCOWra/o1x8gHuPCuZ8kdzn6BBviYmqRJfKGk2bvRjrIH5GlKOkBSlxhoLda/E
nEVHVLWHC4WzudmGI+nmya2sx+5AFIJs7UXI9cmM0/TQvjglHo5E6+M8TUApYOvCsPJQCPh72b3m
VmufV24PutnXJgwTNkwY+VP2STTVPJuib1mp8EbWofhfpg98tvjKrUEoBB8bSAIPmcQtXzyUEg7O
ixF69Zl+mxgG+++3DeioVSg9PZHpIH5xXChp2e6YNqODhMoEeo2dIibxIOazN1xxwk2iAkZ0zaya
SpInAU7WBQaEdeJAAJFOJoTtD/+vq5IXr9QwEMnOgrErQ1FJ7W8d4JOQXThC1uIpx599wfB0JVcn
bOsYPpNvKAR0yyUQifzSgYnmSb6Pzh75kSx6l16h/M2tTkBx4wVsbG+PXj9DE4CGKgluEjAqKz/Y
Sk9/1mGvl8glXq72UoXPclQl9tFPGR66RKr//cSRoAisxvT9/DHpMI+ZIA5lmODxWjphK0D/YYGb
9pIPcbWYs8RUV7ZHCy7IfXiNemEBZZz4YzITI3iXsA44tGdLFPV1jvYOInuPGsKdMGJjGhpy5b7q
1tLCCuv8/MqvFlbF4/dMLfMgTx9VWmZIUOULn/DjSqt3ox2VxeEdsPfJsXzJizqBawzk8Ji3d5Ds
YEgiDhwaj4XeVCKwJ4Wxc79GVO6lnCeOsnHRsqo74oc7WtGxzxZabgIRM60U9onkX4LN+LbfnJ7Z
0JuB1be0WuudLllgUZsAkd+cLENy8ho38rXf1F7xaBLsUMYQBh48w7vwVNQd/dZtBn5Fi5vaEX8c
efoqMdOKhnfyD8MWq+hPNUj19F+F/u1Z1cOoR9u6mcpq+oW5VTot9Z2Eerf6ryoWwtLQzHrWY3tI
ILwmEj3/zX/tVeM9ly0C4+4XzX2n2O6vNcKcrHEl7RpfISxNJQBxryHDVu28lrpdfVJqtsXpH/DL
V5JaeN8QtKHZI1dM62EX/ay4dqVxy+WOPWRGlh7OfUDf5N4wReha6ufR2sifWpgyLtQgKmcQ/Vye
iKaks6D9Q7dKTkM9qmt4DNNNgUKnQ4/fieOPGloT563GQhjdok1qHAZ2iUXhE1pt6yz0cWsBpyDQ
G7myP7x33qmQfyWraO7A5VhOvsTZhnnRYZf8OGRIkpMN0ER0M7/7SdnFEDQJj9ljiyNZobzvAF0U
VXGsZfWdPDO42hQo+buwSM10bPmnv4GGatLNMqkVlOtcstS7/rZ9YM18F9XuCDE1fXB6snkU75Rs
YrqLKCYE8R50lNiJGd+h/p7FOdT2pu329O6qjWCQAV7A2cWHh5cQ/Ct1YyGw5GofiqWaLUKB7hDw
osKMBAvFeQG+Xr79HDlsQRXPMU/fFumijUlE+c2JkhldB9L5Vv+mHc0r4yQPZn/TQ8r//EioQZzW
ChBe2YphlYS2KPRzyvUnYGxQr1vehcwhjokZVaHshzgamJTwTjEzHZY7Ov1fI4Xci3WSZf2KQwaM
ry5zrz4RGbrsHUhnSKyLiU2y0/7f27816C0pFyHnyP+T81t04MndhyPcu2sKwo4h64Afu/+JrUeZ
AlbcGG5dojvMbRKdmslkrjLC4xys1HMcUJ1T908LdpDyiJX4jdPghgp1xvsqERoKVEOCW8DIe2oP
0BC054Jpf/P8fcWvQgFNDo/8s8HxrHzaRpcY7s5df7rpweduWig/ROSp1LXgqvNGRk95xwPMhyCZ
HM+z2Y8K6Sxjt12fIW8/EuGsK9JDZKya25XyCSZTjAEAM+xFnVjaqK/zPpz4qcI9rdQfd1BjQAbh
lrW7eVPL1MLq9OyrIe9ZbK3W9lAA/EGTQYLzjig+VMwl2WOh32v7n2AIx41X+CNvz/lCl0aySzCs
aGCRB3aTkaw6Cc1cxvJQDu2rqpKE0dO5LcbZmVmyhGIKKLrkHryf99yB5KSMqGLPJSzZhDOafs8C
O9WX1sSb8kg5IhRjLLZEkobuSxsRG+SW75+ZEtKtRJzvrytK1nuriNBXMP1qJUaqSr5Sfi0GaKyq
UD+b0qIfk5r50V4SWuDgKs8zaB1qrTxflgpV3iTGOo+FOK/pQ273yWY3ArbpnqWZKuyELHz0j+mu
TcYf89xapwmkXvrzKztrwWboczRbKkiXRiiTu4WJlbmv3JAkLtPURFVxjjjNOFHvjImYOy4sqc3G
cnoXQF65e+qAOiddxUnUjTSG8qLkl6FaHgXVJKyh/V8wxKBVDSBzNYpAtaTKPx2KOoJTGFfZ1QbY
P9I45dM6KiKr8nOEyyHrg+X72CvAIepDVMFNDN8VCaZcd5Z1VHwuKoFTXRxa0T7J3sRZtf0jdh7h
CYFtXfEP378qybcvPaYhLAOgTlfla2zVRuGaDxc3z6ya9Gxr9oufsPXUJvZHB3gXU9B+ok9CPrxg
gQNQOvDNJxIPQNqGDfqzycob3nMSC83bj2SzW1J0UtfUmwhCF/PT5AkVdjLuEdCrZnGjiiZyiVUG
XWvQajv6mxM1SzRkFU8tnTvHxzZXrfxL7yOLOQe2tPsdAxLrQDKUoGmfe8WGhOyich2tfx8h+hW1
yT3/KfIxmKusUGNGvGj/MYzoJfPblrjgqlvyU668iPNIJxMSs4tZSIqyUUWkE72zt+bd9slZGYvJ
0gwasqj3xaC+q6RPgiunZtBN3rJqgcic+wkckDJjHtgEu8GKlTVfFkvZ8e+fsP8bmoSEoYNnWMWx
XugBgIkqLuTbZK3kR45pOrgnSNDjrWV7bQ+8OicjStLWrq5XGgcFLfEjog4fb0HPJUhIrtLp4pFf
tAGg9D0q2tuS7t5Zeehy8XaUbxL76jsjYAgI/Z871mVRaJOofvAUMeId2JWRkfNwof8xaOYn0X8Z
XsuvmztiZ+8EFC2Zm4Lpg5+wwj5SHStfoe3x0wXnvApj7T3LhNNzSJuF+oZarhnWc2S7lqL2GsbY
wSJVLUYqcTIj3YOEP0DQAzXSb/tdROBjX7n9qt6h5NVE6u1yqQ3hDpV1/EeKGU9v8VOrQP2ygfyH
N6IdnX9nGtie5T2T89DeR859e6Zucbc/DatmFc7kVOQPZe4AqG+DC+ZuQvN/xqS0Qawjrh+gBgVC
u/yC9C1xFPGqM69BlxYM9Ttx6GdfHgAjUfyFJQ8sI2K3kB4sgT+MHeXkC8qvCwczrdJvNJc+4fti
e9EHeQ0AUVW8sYXJo1oVlniBJQ95mgE/VE+dIiKBYfEPeFhMod/2XPOfnS0RBvLoQRM5x/G2VUoL
aHYiDpu6jfHHFGakKZupolLrz2babE5lI52UjNjxOCjHlwMLBbNQOwTRLJm9m5PO9NxdP0kFkffK
4pJN45CYt+L1iObsHFA+TNE4P/+BYFfhbsA+8fLF5/iOfFv7JV2QOT98y5wcYKBE4t4QshQFk+z8
oXrYHrrkmBSFfjQ+ZyYvzXjcrZItNJlA+EO9v8gmgx3KeNORE0scEK9AmqyxCbmDZ8UHoVRGP2ca
yDh34Cra/vnIO0p95gvyuQTTNRhiHStGfoX2y8b4eduU+qmaVA/SpBNVaovYrsbP9N3RdO1Eca7o
StEnC36fOCalJP5qX3v9mCCy9os6YHgZsYp0BKahZACiHrzrzHclIw5a1gP4zzofg3FFk6gJOBpk
IOgOzACAu3WRdb5p776oGZgNRoWgFfeGYuQtJbCk4nrqX+3JhPK0CrB2fdznggrWjcA6GUtejCyU
hXswMaGpDRoe4jGHE/I25ayfvtZFZm1aMPvjInnWyZBg9KehwVeicGfnYgaDPWh0AWXChF/lqn9M
E4uljvp7PQyo8IRDmi2plNzRI+TrnzD8xVu+klQmyjDkC6EMpVgIIea6iHtHqfnqT4KCH+ho1i+a
4DTNBuNJGGo5CrYzvzhr0vfaj/R5dV3vbNSJH3nUhmNM5TAAWFc+fIGVVsPRHE89cCAj2cRfrTHY
D68MF0ZE27y1pSBVdoiUzMzXjp88IQpQtlpOIpxXDPz8SGaBXQVTJJJCGCDOzAhjhgQ1zvbBLVI3
cpGJuYO8hG3mgHZhtstIbP92q2qGBZNz/ssOock3jrvw+UTd+NttQSEULhNcMUHRwVeHv7LW7WGs
gVAEHqZ1V+bQHfeLW9SWaasrGaElNdNMpPDG+KCdpx85zg67e4J3+o0C74PoDx+xBISkUVIANBql
gkROTUsMaLrUW9jYFArXSJt1hrwLku+hoEYkkXl9VK0lVNyIMef6zHExNjs2iVlK2/hnaaE5yod9
K2QKOfqX5ExX32kPJcjTfeXNWQ6uFiyjI7Jr7UJWdpGR1i/PSl10ye1A2ju8ZCUg4atqYEK+wsfZ
typlxKeHDiJj0PLyaytpSPHq/nJxVm9Ah6LdPKlZ4SCTa42r2tOF4UXVBHjDxDzyGV9tMaBry/de
R5AiGwHmoAQfQ/mW9s70uZQsrkXXiSozLEyIactZqJN1fP3TIFoJMliTJ1JYqZFbqWh5RjaE87Ck
qNRUoFEUKGPNoS45dyX80ZGe4zcVZKgkY69U66da4mUh3DNxWV2ydknyeKE1Xn3xsZbPgiXYm5z6
0aWUM/PkCPJgLj8Nb8lGSq2tR7MQSv1liTAC7dzatPJbsYyEKqsPHp1qUzg9FpDHRxCTZUcg1uiy
lTMDkecue2YJAhD5IPCBuYJfOWjTQeXVHPPzRXjeT90wSscd8KhYGgdsHXJ8AqmTB6jthi4V3Tce
g21xtaH3zUKNzDHY6eAeOXmGkzhfJHGUpyYjlcaL45PzmMcg7jz4OumGZSb2RB06/Kc3TPrWoRR9
PuAhYdLpRr5sSBP4GU7Gwbt+t1nlfPFtGf6aTZrH5hCybJmIBxSsfHdyHQaRwPIXpV/VFKk96LVl
GpoHgv6XYk0xJSiZfg5pAlcmZvPX2E5ijOL2yKt4Ai/mtyCFokClJLhpqotn42DXMtVSiYW3O+aN
j+iNjsKblZRKMARwiZEYv3BCdMLilOF0h//uM+XD4OfJ205wne1DhvqHoCch5ZU2WWhiFstuGuWp
wvclqqdSl3K4IaZp6V9LlHgtNwi+kHtUbdJOhJOsmPVtzs654ctESOzpzXo0CcTztGNZ4UtImnNl
GidBv5+BrbfiwDXTacMHM+GfrWrm81HTk88ihMJyvRL4yCi9SjIseMP61F3D7RRXmdgVsrW3p8iY
DXAXnbcAJsCh2Zqa0pHDfR/yjQO3jhlKtvoAuU5ikkXW2fYYXA8CGi8OomVgC3rURI3YHbqPjKaV
MKBFIsjFAt8eZYLrdSnXO3a3RwMmjOaGJOhoqqUI3bBnLaLQj4d5wor6tY2iiq/ZPd6L6W7lYtJ5
cfqk21wcPWX+VDpo7ckjcueD+7LF1z49wsTYLOSy91irqCHu5Mhd9ExfFrFvER4Stzqfe4PaaoDc
Jn/0LQYUbK2i5fDt6UA7te5QPkbxVExmj3GVwjpZ/vjWahqHCzQaFVEOmjJpyZBEi/oxvXIAcfSl
sUZgWSWjYJHSB8aHorHLVzvXGr/yZen8D/bH9LlRUZ6Z4E2DfWcSzjaIOJObEptFBVpokLv+dmvr
gEI0v2uVuYZ6jVNRs2BJMRo0WTI3neL6co/eCV61ks7dPLlM8yp5L556fyIvTX0yPpAWsgqha8Ew
D7x2M8Gv5ojceT0/OFAWGMOaq6wNQdAHUzAYwbiq0n63mRTDEa3YRBN6S8KEj6lRNDtMEOEJPjoQ
xAOBWrRrASOrgwOJ60BKxZIe+EFWh4oN5ftt5G1sfF8QcJyT8vPirI9wtj4MUo2ar5XKe9lMjfM1
GH+ypUojOS8mbt405voreBSHxaDD6+Xrx8CsRBImJGBn6YBuHF5T8G+eKsjT44vpTwlrDcQI8x3B
O9e5MNxUoAlkj3AYrbJ1GxnYhYNBfs2m6do7EnMQz6b543xaOV2khfUjh7qbTUlzcNI8PWrsJpt0
628V1BUjoRdivB3XXQKo1kTJJLeozACx0pM1NGu0oy4Pes3ZPeFHQkVfY433BqrT7waNA0sziss1
nPgPqu/aooAZw48QLd8WnD9frMyEQdBytmVAai84IonIb92SaNSztUFb5+7uGBMjcFTUGXdyOiLY
QTNPFSKtoRA8KUVUqByM4OABHZCnvquZwM+uM+oY8bxITz1uEmB8QnoWRop+PIZdtnwowq2d9Dnw
5TtMudn21yzN+kPWSrXsfN46PKR19IwNOL1n8EVvt+4sgYM/6rc9CLdBZwpwghgX1u5mq0R/TTRV
qMrynfcXEEqGOtloBU/uGiT67bNI6bgznUbS2LjGaRVnwTXhY7bSYfGTOJ7+mbe2nRW/0EOPaGQJ
IYHp9L7Onc7je6U4pP1EaKVaihSPxFAHaFGIPuz+8E9JXyelFVI1Oew+XY1NJvsZFs6aepg4DRgB
qufhxXlke5m2NdMplfBvgTFCTn4wlq19Aw+313f4/xc0TVQpxQn1T2V778scFinEjSNhCDcAvq/8
4Ly7jdkV2ZRdmgLnr7XUhlFCRejVD1fCbZXtQO0kuxHkHCmxE7d8GOdE4OBbuV7BnT6pqgbffTM6
6T2icoBPaGiPgDPKbiRBRnSEMeSZ7/gmyRB6V9657fAd3MbRIIuolgZsjuR8PvJ3HF0Ya7zNDQKO
iN1mDV0t6mg88h9W464xywGREVzJvScyKhW9Jq7fx26vALHn2/jTd4V9ZNIyjgc+TX+PJJ7KCNrX
wsLory7ZvTX480rNVZnydjfJWYFWMDzIGZ3ShYeskxKtvy9YKc8w+cS42d5pKVHryWDzl83R6zqv
5j/Ef7gUonQfYyW3uwXIRM1GJBqI+1bogxcPJISHR9cSiVkscxakglneGRaCKk4Ik+EDUiN7MwEO
vSWqA7zZCxYvdar/Ag8m/i4f7uYEttFlqvImn8GHmCZMbR8jMquUYY9NaxAPeKOUW/3sKUDgvnrA
IqEgqtwRbefxxeq2S3LJEm18T+ejdAUKt+px6pZ4qg+7o+S2XGDxQGVCXg2vvEJaQgjTJu/1/LGi
S5/6FFFLmEqjjK8q/o38+p/LnFvN2REGucPWJ/3vb385/W5l7BE8j6//kucXEA8+7So32CeFNMfY
j1shVuAjUWDfoXu+mr45in1KbpGVgeRlWhWU5E5ieEaEOV50PatJByuJz+K1sCDTU38fR8xNY6AS
IwJnyAyLZNOKVXaAqJ+ncI/0QNua9jM73HMW0c7EtSBwCnk9Wjdlwivm3V0UT+a1xsn/Wcj0gu0i
9OFcOHL6ysElFNwQwr8mvedMEtUQugYgmPN1hvZi/yoMlqMZ8vo+oMs6wOPRSlaNnFV7yzEWuBN0
PCcrAaNQU1I0gW6MK8xif5gPQ7yDiUfrS/AOc/5Jtg6u5g/lDuYcUyz77trASWRSMo1ZbzDMrKDT
1A8f6Rrm+y8D+gjVmbl2nYReDjV9TumWIXYf2jLf4YrMG5TjKP6AOzvaDXJ3G5OLdaiqidhn1XnI
2UIrE2FAGjmaBjTHmqzqQ4YzrIzgSvG9rhz96bANHRfg6ynvB6jBY/1EusyNJYLWtBkaecR+mPY4
q4vDOYMVpzBc79rk6KAL49Ovqo7jOPmNfz7XFzh36nRhVpu6Nx+kvLgpAHdkIz/lqv3LPp0L0Wlt
eDtqymij+TzilKWCQom/Fy7P7B8Yh5//OOyiGdu+YxaDT5ILfaDUwALhjUHcdoWP01EvVSGSdltd
dYrBQzhX903PUIT+Ws+crzfH6BfWiEW2f0xB58W7ifSAv2HtdviVSqKANI8vASXpeHxryiZ0tVoM
nLytlBY6kbphjo/gg8BX9+YzxTKmC29718FxNbV7LS8HH7b8978MsZm0AYK2rc8F9Uv4/izgDP1T
ZENQxjha2JndAuQThEnXt0NqlV8Qv+f6Cs0Lhf/O/PsDiSutQVpu2vEMgPiBshk8dne/XFhn5Y86
rM7NjWipuNzQtjNYDXvKiNzw+MeKeojwaucGz4Usre4rt1FwPo3PHnss7IOSDzmKJIs/gcOT9u+u
uqmgEGWdCfma4bCb6x2yw8+rfhZiL1q/t6SyQA4AgRf+Qp6E2i6K2ytczvsvRS5DO7tkNrzi1qyl
cFEHSgflA4UKoWSFCHJbdAhFSKdllib2g8CcWsVFscO2dHBSMVV6c6gp4cASPKnqzrZmvFmSS5Yo
lfZZbPYoLGhpWQENbftKPX+WxorXszI1kpkjpgvm16cMUfjxDVl25sCGKqff2l/st0FbvE/MJh2R
QV5rWso85Kwch4Ifnrov+sbSeSOv5RYdz16x+FjeKXCH1lQAspRnKMvtE+pQR8sbuFvjodMDXdJ9
WQxslrCMJTwf4W8wnZPrEqXMCXAZ8QGC1hq25ZtrjN7aGSp/MD4VgFNfBpTrSq0vVsNMhqXMdBhc
VcgnhLjBFgK1/c2JzW22gVXMGv7Dvq6BhEUzeYZ6dcnFD3MZkXgk/HNPvG4IOP8lfu0kwyofjz//
clZCf3pHMW14vvk1aAVZ9fqK44VQt5HpJykkizobA8w+0LvfcaUHlobzoYVvSD6gNf76Tfs5dFFn
XXqstwxkX3furDKgbDO58UPOcAXrMMn4yqi41QtHRC/jxgf6FTm1nm3QQR7pxLARqoUrI2EcK/Jx
fB+V11VdYlJPIycW817ZMyAWEAwW7Uj3LD3Th+Ux2S7k/3MvxW96ba3PKJ/K/pjzCNRbLMW6o3lI
FvK2UK12xOjj7ULPWifZAo8Xy//HTQwf9hLHnjuZ7pEvdgLt9pzGjEK10lAzwUMiZcYSMOGq2v/A
R6MrNjFXKwoAbBOeoShXVme8Vy6WNogai8sNsm63NbRPuVEMD4EICP6RuHwS+ldzPhTr1+el33Qr
0TjtjZzKvCfeUWqgIFd7NJueP5gWN8b82n6bZPvAfi0ujmKoUJ/2ZygvfME5k9p2gLiXpU8lRuK0
ziF6jvksjt5FQcKo4HMLww1qYuNK801OTlM7r+HMkPvVj8J7AG5egnlROZaEefRDzdq5pHL345RQ
u6UA30xrX8r/+0a2/oi2oz70wCpn3G1M2yRBnK6UG8mBjlKCqYgnGconUK6am0fSMSadZ097VSx1
ThnZOwTBV/7jOr1u0l2F4cLKItagFbDVsKoQP8ugfXM2vd6LCWW7QdXOyu+q66i+Xlumjg5iTosg
sbcdFxhjVJKzB0nwVjzszPRCfJKlbCiPRU1RJfvyS54HOEgaNAdDuHmQxhBRxXMPSTUJO6MJwQdP
qUJxgI6QdORmg9nuvyyDVeYWDzs2NnlShgi9vjSCw4lVjPylua37AlhvHprDBRiAQRC5MFSNNNlT
zqAYVdsqOyZbkVUyO38w7vJ3xzzDWdDIugleX7gPgIsPJZMyvs781AZJ9t1PmiZhxONEY8w9beL/
pyELAC2FLqwRIflEZP0lnr6iiJ/h60wO4aKsacWhUaq6ABRjqEI71hroserrimeAY85ZORKGzWXd
6SvguFSLiUVC4IGnPj2I7SXBWXgP13OwH3k47VogGNU=
`protect end_protected
