XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� B�P|��;�2�u�\���g� -��O���T��}�����[ww٧C8)H
�^�h�g�< ��0"p[,��o"C�>�K��H�1�^H�c�~��|��m	MA!���KM�7��݂��x{�ld#�e?�:&nгl��-�"�$ם�,�?},ŷ�𥔋��������(����G-[ZՒ�s����DƄo��VL��8�4��vO���$�Z2{�P�Qbm�驙�3�z�H�J�`��e�({�o�;���tE�KX�]�^\����F��� �ך�nb'K�� ��]ųӪ0�~�
0|�)~����ը�'��+�������b-@�vj�d��>f4���R���a^��+��s�вF��Zlh�r�3ɀQ!y���^�dp`>j%��B�Ǖ�~!ο�9���T�mp\�^R���bjỉ.�^D�U��ؗ5�~B>��6�J�a^B?=�*k�dD����ɜ��|����q"�a�@tu��r��m��'���C�y
m(]�I�����= ���4/����?��k���B%�)���P��iyagfʘ�mR[Ӷ���$RB�F�8P�$�U����-�\Q���P����&5���R�Lf�0��3�p��������(�t�'\����?̙��C\��8�ҚN�(�պ�G�y�j"֎���5JO�Ab��z���2;� ��Ǯ�ö�b&�Mګ���c�l���DS�:c�M�ΤaV����v�'`@VtFfo��Y�v�%V2XlxVHYEB     400     1e0�~2�j������I����7�nC?5�҉��P�n1�ĺD�@����sIz����gR׷Uo�\�3G�7��d���,�*nO��$�־N�cyh�,Z*��݊=ּ���)Q�	�s�ϣ&�f@�X����4ċ�A�˃�>l1�|�3ڭ�zX�1BE�v��:�i�����<���"�tT�����0�Q{;��h�(����	NB�a����H%��c�.��>�`�{`�D�7&%��|޽��ď����E��S
�;$e��i�mԂ�c�h2�ŷ�lt�UZe���!���ܛ���V�	���X0YD��)Q~w:������zl�";��M.���E&���!ԓ��&~�yi��R�V�U%�>���g���Sa�Ԅ�</[�M00�gW�\ �Z�Fd�c��&��sQ�.�6��w�����"37�{un�9%�g)z��&JV~��H�;6��^��"���i�oXlxVHYEB     213      b0GJ(v������o�x
�[po.�W��tCV��E��s���ы�x�"!:��wS��}ŨI%��M`c���.��m��~�5h�Y��7AʈlA�6���RmJ\���C��d'�y�Y��r�<29$�,.�ۈ��=m�DpO�����t�׬��r�(^��9�-����S