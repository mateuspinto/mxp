`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
T20EIAVzZTnsYrxZKRJVsXcDYM5xMpzqoIVk+qhXZf2PUwSLC3WhGtyeadyAmrRAtrjzzbuCi/8x
mcbLLttgkefXxIm6h06oMNP8nF9n6SykgGPzkdCbsOZkYysroRwnf93q7nFBGWBljtMDj0g8aheG
TCJTOKRWDxy7joC0JFrjfpJL+BwVQxY7bSmVmxOVz3vLLmwnDFJV8MWT/6VpwyhQBYeeXi/lW5bL
KPpifdP2DCTv0l71b8pYAz8xJHAC3s8eaosZ6ojzeyFb0L8cozwxnpQn5fM90QLSpHJ+N9DmE6G2
P8tYDvrwJ3PjnDGm+yHktPCW/sWz+9w3jr40xk878K2V7Iq6PIIeAs4ZpOiJCNcuGzXOLZK1bPC2
LwaksJbI6puplpdJGrkXrJMmMh8SojnWc8WJe2IM6iZRjmbT1mk3118+rV7LK8pLC7cPIQ5fHfqx
/CG2WvU2YJY9G6FI8ya0Bj7+GPQ8OVWda+M0dMTNzGKceGNPx3ITMk4cnS/KP776dpaRsh3+Rhoo
ZYN/KjgJhshvvymegi2zfWgfSf6nIk4LcPB+OPSvcXx+M7T7uK9oZuj6t+g88dRcJRAUgZLUNxLs
KfJl3LqvBZjbGBeI1ccZTtpUmNGdPy+9Hpi/aq7E6VzTxk8sNG9D0I8VwjSNBvEwDWN3/EXMIB3m
aWN4HoFGX6riQHmt5wqjoGcGyZ/fGJ3XwEEhu1whQvInxWIEZwNedXxtHo2LaBB0xoztiLnUEBSE
7bi4YLhHAtY4XwVm9ogCH/Kdr88EYnRuFzHPas1ouuzvcsb1VJP1S4Vez8iQBQZ3qnKWjz+kgBbj
tVUgKHzvmI4FUUUW4j2dFm8zFC3UZrWYn/UEdsBMZlqUEYyiCgzjeh1vEubYcNUUeL8iqnnd1aKD
Gv31rkTirx0HAY20R+bpZrOzzxYRAEgwCSgVsGLlN++6fs9P2E0qAfkPg4StW8CVrZolXaXkzgq6
AXYM2ORwef6izXrUD0lEkFlnez0iHJtU1U+93hcbkn93VYUr9bph8vT3IsEwLAYca2papkGGhVSz
7eHVyG4mu+nnAfwTLSu8phALniDXmwZ/aqj8cTg8KmW7JpmYhCY5LAcK4dWIHDpRJXdZnkbt+Yzf
pdumuZE6dasK2RblgBckaLgw6I7o+MzpaVvvDElx6darpE92wit9IBCn5HT/Zm9t+xevj9x1H5uh
zxCl2nE+OpcPjrS8+0w47f9yp66D1akKEnNxREBtzVqxunNyC9d0gDoXeMT/XcLGwgQTYwp1BZ3e
Y9515bC5BcKSjON6HjmakgxHc+/cmlFOQSbkzS906ZssQV6ZhmchaY4Tax60MmoPceqq0w4qb4Z2
L8zIMdocbvoHJUzm97AkIMP3Ncx3qvMJ/goRPwIy0HwTb1qjs/uw9Rxf9paHMIJxy5LMbt2qhr4C
sLezBx+1P8Znn7RsRur0Nq744qVAUbWDNsw4F4Vz3OrPdLGI1gjr48hatDjDjlTA9mvLQuz05SyJ
/MQVwMi3j08ChGif1l3Dh/vno0hB5Bg/Hxuy4p2i/a8GLzkZd2mkbu5FaJltqGUN6Ek7FZk0jRjG
3E8oJg08JJT6U3Diyo/g0jmqMsAAg7GvnXbUaEFX0ANhVsFXxutHUTUVpnb+NhlSUn/xjmQPQXtg
ra0gqdO7D6hGxLVJR7ljSDLJj6Yb8QrAz5KfuzTusMksCljXSpieLEHWt9TeFJridrAXDOOY88k+
7XosH1JxtwBT+FCiruYRUhHsRjTm8UAmj5llSUB0D589MvmUIoMB5nc7i8RjJJF7Y5kHdpm/NRj6
WmcspgHgqcmsyvKnNBlQDVHiQeM5rqVDElEyXVqCf0dct95ZSFC5EtM6ZV1k6IKRB597H/BQ82XU
2zK9EJwmcDoI0Ealp5kQ/GJf9Zw19iomRPp81mTvDsbqtrdAFfOTM+3Hbr8fwuKSTpD9cr/XFBsv
AfP52unOr1yY+1tJRpF1BjAFLSTO1nnsMpnimexZywvjZYPN7bsVslOq2gv8TmLIvUcAlvLnRFJi
Ve8YG9p4L5IE1Dg4lZRuR1wkpp/jBoZPXYoiYC4XouewJZ2Iz5yegsWgxI0xRK8Xfq8xriTmIkCX
4JqxNSqePo1WtaHvVYUXu+Cs+kLkkjjbzdhBrZpnYflw3n5xoHjhvce39MqN6R/VIDHtCYHFfpL0
Fg/iBowl4w0HT9CSe6Ty2THXjk5ybADuv7XdjTX70SJqvdrjplDK8FTPDs1BrA78ivvTbMdW4TwF
tMfBAAqfO6XXEKwg8TwtjhUskd2mBQBLIQL6nqoZf17QgUvzx0NS7dl0aS7JhcjNQZ581XGh7Hy8
lTEWjrAiWHRSUP7DNg5J0ILkXSegBXYO2E7kU3wP/isPc6qlAh0UnSc/0msBAh5Rv9QFp4VtpS4U
tdu4AXo72D4iI/ThxS/Nk9dS4iSXQ1RmM3KJ/9udZKQQlqErqBwNQqD0PeffW2B6LZx6F8vGxXP7
j9c534ngNWaUDdEMD8CJ+fVXEEVQKQZK6fsvr0enZOMK5mv5PzBnjKEzRA1AF3bZE+Oct/6a1ujj
ME0QZHODcwE7VqCkvRzeNbUNOxLsX1xZg2tDmz2hNLGsoOKLIM+eh5z/CuOsvbUI33mFRuCrV4Fh
/Y8TWeaIfxOuvAt02k4tDIpuSwSAA02OA8J+JJ7z6NjinHAysiBfKTbMaMVpNqfoanUCGqRjSfb0
DlU0SuxIZxbvCa/cHEjldhh/QFSudWu5aKn/wqFGKAiMLKz6kOpCZcAE5MyF44GSNTd9a6a4moAP
NPrS52BRzs603K7Trnm4d9gxWIU6KrIWKwRU0LMCpSWLFyZxS09P+USkAcRMf6Jx6RwJ6ONdaCN3
3Ws9x5kzlbvnuPeF5uGGXVTIpU7bXp/EnMsUCHGbPckKHbKJN7eJAn6hkVw6vX0K96G4Y3Bj87g6
1dNCXE+FDDr4JpHH532FD6tGrbBu5pECtHBKU7nf/WsQ6gmG63ccYCBVm4teX8HWde7PXhy/w7GR
0UViUCTX13loAF7uy7DdK9egEjjXruteMR3/mL6qv/aNR+009hQ24Z0FKj6fTvo1RgdnILnI9dtK
echkLO3dCFDZh6MWe9nOFr5/jWYF8SzyaQmV2gNdzm3u9366bujkRpcYJsGj4LaRkf9A3C59t4Ci
bAXTws/7yY1kkMC4dsD+SJkdtMUI4KCafb1WI0V0JnqXiCO7iEYqWuI4Yto+O3tG3cs6x2Ie1BEK
6l/jdXud8PX7bwTc/fCQow/XssZFgYBxShTq50uc6BIBgUbKUxAEO7wqR9njioBxAE7VxDlz/2zr
eeSBf9SFvZWWpUeY12indTB9j3ueflZknGYrK5nyJ4skWd6v/RpAznm4Km9QH8LrnUtvTDIK2dcB
NiwYhc1fNg5Esosboa4MMJwYIQOIJJbUuRIxx1scoFWVNbBv/vNyCeVmOGHWV7bLj7bWNR4+acix
x8SDl9K4HNJGUP3xoaN0X/MoeElTHM4XQ0tkpIQieKKzeF1LwKeB8WprbzYIZqsP7qWKiHBwToR2
YoyO3J9011q4sQaGLzWDOBriucQT2zueCUFT+IdcJukefLiYwD9QozgJdXgDn1vX/2wDE28yGEiq
MJfkadzNDyRrEYHy8hjv6hcq4gwNWYY6JqrSzJy4sCKKI195MUxCp6jWd+m25Ux5/9cblxH0eBIc
7vDcbGX0fFD31QWOSEl9TTcQIaQ91rtKXr0lz19J7h1lF45axH5F3MhmoWGlQJ5WsB4yWveHLfbG
THM9DjYX4odaFPgHn9oY67UgsGtuy/e8CxnN8u34nyBVB3xUcsPWkR0oVLf1xpmI57lxWNZMuKa4
LuMw+bZB72h1yhjhaMq806yfxASOGdpzSl0Igpc0wVqlvGP1K8gTkER0WCNLOLaX5dsXqwoTUs9V
jyf/DdkotTDD7wsa9oDQqQXjqVIXxYTbBvmG2PdsxnPb0AqzBJBOIMVqX99IhrDg9tBwdoLUpfOH
WoFrBAFiSsr3KVvA8q0byiB79xF0solZDbSRkVqWrqN3fx/U4X0GGxidxhuL8nGgHoSy0f5YArLw
gFe427i9419h59L0JOY6djPoBpl2A+n81j4SrON81dxrW8yJqgi+LN7xUkOIm+MuZBbjj8NGe55d
3ONRAh3WoHIKBmVR4i/6jQ74CiSrYXkVClBWXn3Y3m1WqnNcdifvSc81T+nHLNKonXSz1f/XQrFK
dfF8sNMtLxe/wnQhHu3vOfipINB6Woyr1kxsQDkPbTcOgyuVrHVKn96svl2oat5ScBlVd5axKiWq
LK8z6Yhn+3zoqUaAybeWDhnXCeALSNLUZISdI4n34SIsuIC7VO5QRUB0eaeBEGs4X/XKMNItrymK
BqzQrH+AenqomeVK4zMhFUaXCUJrQqZU2Wj/i1IBQGWsP6bBQgcWFoIRvmDG+X84Z6andaEjD/yJ
gVuhEb3VAPIcCCS0AfT1gxP/Zgamh8Z3KF7UwE60sS8DOOVD1RiP9vjI618rsuvkbqeCRSHQ73jO
KxWbF7EuVw5jBjI4qrg9tPT3qkV36W5pCYI5ZVWaJvpXsadwtTNUNx95xzixYK5axU0NTobWExOX
3RPCa0Efk5AK0XEKIHOsCqEnqeTqAQP1Nt1nZGjKx0WstPefAw3LMCt/CAx94Xejrj81OJ71hKRi
Zn8e4SN0AFx5kiMrv8Z5kDh4lqfhZIoTO80mW2ujKVURWTnU3dEoKpMEV/m9LYGNddQJm8kd/PJW
KTPqB72xErxakAR9HeEaYaZCNvdq593VrTNQH7fgNUxuC9NBBaw5GrRDcCw0hTNDrZkNU4TPD1cn
GP6NbS6Fiq2lRnxKyiK+Wh1ziY8K/SsoCoCHssOlyTH+7d15RKQuzWCEHcis75r0yamLrrphLn49
5Y/DMEhK/xKkxokrq4oe0LoYBnJ0PRLukKgT9wCVwnA41cVt6IF4FSeQSVoElMlWgrot7finRCsr
e5mP2mOAlT4fVeg06GyMMM8ALNXUGhNH09kujgNIACrWjMO/wXtAC47npCd79FXgKaJmGGTLqyS2
lZemPLWyaUuZI6qTjJC51aqCkQIBJ/ibZBJzYcrjnl1JvNehSpmeD7DkrfQVyegYL10ABFfw/lOS
TNddz7ns/8V8J44RdxxNDV19qS7RsY89+nbLVpvTh0MnId+6o7jKjxF/cj9wrFIVRwgcCMcy6iZj
4wU4a1OLVfHl6kDT7Z5Vy+B5NinblL6tlZFjeDIf/kAvNZsXUdjVCTirAsMZPCKrHnsxo2ID7MsE
wOVsKodcb6XINjyhGXLtH2uIV/W9K2q3Bgby+obBVJHYYHf/WUn6sZkwQm6NOi84gpGN2Z4tsxqe
AXGnBVRhiRAODddGL/qftVu1eJmM3aUGkY1XJDS4GkNcB6cbhf66QLhTwArDoYiBJcSbAN/SGKwY
YU1ahoSbclckODPS85Qr8QSQEIVwStUngq5LSTl1AI4I97YlZ7EhJ725JCJrkpcckgPyikUZOaoY
iFKmZC1+92iQiQCRjsuVyLBYYchqtcJcXQGLTOVtTdPLWjKcstKYgGtoyE+i0w1phH36pf21Pw++
axCFvqpJD99Z38A6KVnYRpV+Ccug4ZMJXIxZV3545iTr8GAdHjVrtSpU7wK2WPsyrNWb8ogLDiqb
TZtj5OdRWW43FgeT3RVEdg8/dhDQTNgNuqh5g0PU6rwuur1N5MEZjAppRYNHllL+SA1tS7Evavjg
algDbD0BncyEGhMnWUWnhu0heDUqIpkgmjffC5yz1VHIFksaSPA9034ApVnbCuBDG6/+5mfYrhET
/BxqTTlHf/IkpRn1Q6CKL4J3Itx7nwRzVyXYv0Z6A2+lJ47dRSwpgXoOJYgbcfHDMClEBUd1guXY
+Wu03DcSuchU5oNzTu6NfDnmmvcyLR0WN7zPF/aP3Iveark54gUTAynCUHO5a8o2KVUFPO8yFUYy
KXEJyRN952vrpPeBR7YnCtZdRrlZiI/AIbFeznbgzoPnfvzEqpU0k6Hltf7iM3PCv8BhZkbG39/r
Uj36cULA8gIaqWUzHVdM3G0IO5urPmi6/txa9fVn43JG79gVkrSXdASWLfiuM4ERYiEUgL/LuZY+
TjMKIDHAjqo3zUvMfWetbg/iE3qtX0Pr8INPIprBEoZw8UjQ17u+wh/6sFmd+HbDDUocZzYnAqKM
SPNvtre5yE/Z8NWFyfaOuQ3JZcjluBvq4g2RhHHghq6+mDoTi5q9UaDPEjQXAQvWSCW/Xpy6qc8t
vXw0isDJGuwK9WJTzT7mYpxHbgf/vH32E8ANgR5nRGZtACqKzJJSvdusWt3HthItJbKjRTP9pAgM
3EPWIH0nhzKbNI7l+OZ5WVAERv4VAP4aWsLEFmsdQhRZ9CyunjJkxbgR1vOTBgZNn/x/vH0Pa7An
tLKUgUfcrQmabcRVOyqQ+yW5H1S3UPdhy/hgCAAzrARheuEPeKM8Pcuh8pvYSZvTbOHHpHqZEDNq
WbVmfrzgue3qN7vvXXe3V4PER0ZL+T6ZyVp4W/soc1NjPmXyGqKfutzVJ/MexZ5jiweOJt/w7gRy
NNCeyIsaMublCYu5S7Tof86xQ58u2x2Zfg2DbBQaC205IvlBDFMF9xItKIHHmTgm5vmxohM9NqDp
yRO2l62OpE/UCWRdpaOfOXMPisOdzHcOrfA2xVeHQPTtA9Y5/4GS3b+8eYlJDh5Y8VyllKNIj638
meXPwz26EP1mJ0LqXPs/YTJ8O5BreI9j8nwTFg9GXy66OjcfxNvL1zQlXXRA72Ssi2tyBwqixTLs
d1g4VqgBk6Uy6VIogQqWRDH8BltZPLYeZkZaWFC8+xCRu4Rj29ys4eK7l210MyrzvLdy8/bgxzHS
GJoVQNYvxX78d5ohxFqprQD52oaEWUTcGwCDDR7r/QCrEFvVBCdBQjo9m9XAIDsN9FpT14lvkd5h
6xLuErhDw0r5iT6Jjb4m5ZAPtjOi+VN+c9/siLwO3crhO4pV87UyeJE2zIh7V/hUSpca7Qaef4pn
mLvG1m/CdOfa8F+qA514D0uAyCjYcXFDBqhpabZVsSWHsgJ4jnq81vZC9x385J4GCAHa2BoBsA38
H65FHhm/J8wIoon0BE8M44bCid7iq9XZUXBgaYi0le6XehonI8ZcMMFfghSwGeP0sELgrFD3hndA
1Ty0UuAPm7zDbrhU1uwcqnKiiJe6p9mNGSIY5l1fOKVqzRItWB2yQuYWzfv0BAsfQVz1M9bSTOoX
TeuvJ3hOqqikzVEwDE81/r1ze7jt+sh67WohsWzYUL5Tv+Y2nCyzI5EVuiw9iouzPZrsBO3f1p97
WolI+boBy9P2rNkk24t/akYSG8uoSp5XRmcA/N9fAufKFBoLtT3eEX6FswW1dLZyG1SsxcHYO4Y0
qYXxp5QaQfNN4y3tH7CPUm++PeYHa5ifafKkU43gaYdGDBXA9RD//Vh/yjdt6YnuIztlKeMyAN/n
FWdBqMQXdsGpPhZur/Fyb3ArKa3/qByzcVC3kriR7Hq/ZrBQZQ5Ai2QuizHh+lkXInbewRFkahip
W8vlobmd1x6TEHSCdt1s13+SOpzcVWslGe26MzWotVvxjCKg8jbMQOI66ehM0L4LuR66AYo6w8mO
xTE+8vKsZqfOqXgYkwWuKV6EcR06uKpCKR8Gp6aMTe7q0TZUqKghDD8rmRvwKgpf98y9RdIKb2TA
GH5BNPREV0dhrm0AHD8CqkyQfjKARtISjz64UiekT6SHzHcDfnkSxTVO3ro0WXZUnWkvfJq5sRtz
foTg/VxjB08DB2sleIIP6GahXp0Jqfs26fqY4EC2kZvFn/u9nD068aDayYLmWh6LW0hPCrGuQ+J+
jlY0QZ2GxvLyFxyhE1jtxaprQevmp9vAMPmkCPqWwl/DU4DICD/1m74kpCPnk9BEOk6ccgIaIlwn
9xIPEqKmRMo8DZG8Ma9gquz5bYvB3TOEikiYvf0nCzYDzkKwWRfvmLPhBugCrG0h8CbROU8MHnME
DUhj0qPX1JpYIbmyuLfurlCzh4ZsqC4wZu4DG6HxV2NwgUf6oWuPfocIPs2iJYKNbtG8IfuKICY8
bPTZyR1+ylDQfQ3EizGsfZQ51oXQg5hBFSQxCV/AatCEd3WW8nhND4aE6e6D+P5A3TwRDeO3lBTa
tYFpqxblIK8TB9axaJANZa4HktjpOsSLFZxJAxXMVZZG69jHfULOrfMAK23EGaOhd/dYwfsalD+s
H7RQ6F90uN2I40WzxVQb6yNIm1LiANY2MEwGIQ5oi6/G1HifAxu953K0uvsZH2ydbo/PsPU9gGe5
KnZhtemXzhJ4jZta/5ZpQzkBhr+EGCFUGwzeKSrM2oAKOJm8azftnOqch9N7EMr6VLZM8v+nAxFA
Q222Dji3fjyH4JdbFl4d2C4YQIrPUxQJgu69ETqpQ86D2uqQ4sP1n4i2sIsUxSfgzvyse4AwzboZ
eh2lH4T2FtgKtjM1aGH4lpBwQtUGbhIg/xu3Ow/PJAiTbZiefNdfZ34Vh/LQ+M8Rs47wjJ4UD6qZ
BM74n1vqBze5agr0F1zZqeZjdMlArIjltZ4pIZY9N79p5Krc829t2DKxGB95x1KbwlGKcFCM/Ifu
Laamv6pRws/SqBlOkFKQZw6uvCJkTHfFE6TsOFoW93ll1hHXQgxU4wC97PvZVIUpcT3/rkUdNc4E
3segzl0muoP5VRyrq6lKAcbBMEaQIq0HdOyKARJA19IbVuo40aKz29aAxfq6yG/Cqk/VcITRenYb
mYk5h45dpGBEOLh/akeY21xI3n9Ifiop24woUZIT4HryVSQLCftwk9J3C1/81UhdqnvwhbWVh6jc
gl4hHKuqXohvoH0Xq4dC4fcF7DW7lAdoNZrSHvB27UPwOhRWvwSouad3jvITU4h2fN7jaKCdwoG6
qV1C3VqgeWy/qlXwmUPY0VGVnk8aMZXVwjlRPfhttu5jmV+HxDldAMZthpT5tjwJOaf6Q033H5Mb
WU9t0UixRt/5OcpovoJ4bZzaReXufC7WbdxC5l1+d6xSaMDnsij1rvDiqsY4MyLaA2c6HDzHj+it
O5uEu7gofSmg4fF1Waf7R525iER6UJ2ZyGoaoGW+7/Hna9OhfjJyPec5Q+S5yZJbZEKa1tVbzQjG
fq0eNzHAs4F4gp+1IjBocH7OF2sK4n7MTa9izu4+ckKMgNU1QmZ9TALYBz7cm0tGXUpWXUezF8/B
ovAmMsI/REW4ySvE7g0ix6KL8oJct3J4mQOe/BdPcYOf8BvGOgCMpHihDEsJViC/GpfHuoa5QsmH
tO5vzO72i69FbH+eyQMgWQ1piAXQx9PD7MUSBzTyHFCeDaI8fP4M2NffQKkWAyz9OfWuV+Bejnk2
nhR+uOg/OQNTWe/Jrl8O5jXn9pwqAzJMtUe0kPGmC0NejvZf0UBTwQLX9RMEc4FxxRcEi9R5w0jb
bryVEvrMeRnbVqCeHHA8ZGMImErL7Bn0yDwcZXthUF6wbyrOIJZ3fJOo4nANI/J5apMN+5P3FXTh
v7EyMS7cEiSp49kzoEe3x8nWsG7uFd1Cb+ed55BmOY+tuuv7P/fC4L48thwOgA2k35rDPP6l1m32
8xfiR6hZxaDU9fzA5FmBbyh0kXmXkfCXaFFy4F0cRCCeqcV3hTXot3Bdv63hSMPR2X7/BbN+6Rog
4KLrItbPkQBZK9s0uY9wahbKUnsVy1KTMnbfuiFgycAeoRuMtHLQmASCUTfTAkZC9BapD3y98d3r
loO5VKN2sb/ez/u4W2/C+tslFoCvA164q6KSgIJSOBu0QYFiU7cQ7eG8DT9uQtnaQ0cuYg7owDJS
iD6ALtqJh+iYWNNiIO6Y1i0uKAwxUxnPlQm4A71KkFgrQGrPQEPD+tsKKz4x/NdcRBwEDknQeZR8
RoH3Dlkv0sM6hfwJYFd+itrHydwzmhQMn0cIQYvZflMJL2ZGoTZ5qcloYCPaN2CMFgXy7j2vP8jp
6ALSWscpbqHZu5vOsI29nIRjz2EqlrW3a0JYY92j/kIvoezwfCKpiGunsEzaAn1lnwJTbal5U4uj
tTrswoxphOw+xZUIYOdab0FjvuHXjdnygNlStE1QZYYj6QiUcX5V7M3pAg3RGpIsSkAY7IqyHncN
tb9/qhahulV3LKEn/lydeTI8piTjthwfzcXk/hVhDRoVhCkG17XL/LOXwcmL1J/j8nis+OjQT9+D
j6lvcDZNm/C8PVotbqdmIm7FGyIn7Jbsi0ixOMSll/LWNVqju3QIJrO+dAKEV08tt5FjUPCXhP46
FAWCDxkzn4YmzAK1+elE8BcwZy1ZZJzS12+MiSmEtT9XqSLHRCPkUgTV83Ut/a2sRXASvfeVBQ6F
2ihdrF7C6jVQBANT4hg5TLJgU3sUAf8mfZjI0qDqAorndNrv6GO61Ji54EAmMbXR/HmdIq8VD2bk
jdp6msCln/83UyV+nqbtLpccU9i8jKTOiJCu5AVg+H4WmjM0kabVmIO4O5SOiHdaj5pJGcLj4aFU
PaKeJl34S4xIiWf5/xWOFTkurQoaeNRIGCNgihBi7IquMNM0kFNtWH9gBF54ae4qtfHjLL6eVuz7
xQ2I0lFQ+2pNpaWNhJRcNqi4ZmObS08WoPtdd0zEMvFi/CNgNhNl9qLWfwDgOPFpeawm81qSIVRq
Z0lPDIh+qXy2jnGiUVbByRAMbd8kVMiU1oNuIwadl2hGcMXvnORMbHpBJo7Z1N5+wTZJUejdAzCM
dzol7gyiG6KKbS288ugxY5/rCQij4CJMMD0DT1IEjN4oP5A6tIBMCvT4zPr37FY1IuRndS9niwhe
r2bbFovPQ5MOgFyCEYcp6qLvG+9qvvBHPYKn8OIWjH6A2WC6he8GYJivOaLPYqdvEjTIFjCnQROa
wBbICQEPNqRDgkFgHfz8GeVp2uP6LVaLNKVTY6PL4glje1nZNnHHLlZaZ7AyRwbW3IPRuBpho7GW
ngFu3XhEo3j+mewop0Z4ecwF7/KavItpBzAB4DQYoDqrSEXW7Ra7mzWV5GW6y8IJzu0/XyerSwL8
YKuC7AuuFbJuunvKdRYqxNhFGq7b7T3cYbm6FJSrqeAci9JkWVmh0yFCoSAJFHwg0v711FPVyBrf
EjbuqRhSa91py7gagZygZUxwg1Jez5H9Ivhzamf8O2zVnKD9hd3h2he/xpIe6lRYOF+5SS8LY+yn
yIPKFTCEksbWZtkkQ8DueanXygLra0Qvs+/au5ZAv3ku8r58vxgIZDpZQlqviLMZeaOEcMo0PZMb
qUKSRkWj9p9okqSZD6biBPmK7ybbKG2Rn6fL6UMWrSW33aZeOsgHssGANuIIEGY2JExRwQDBxB+d
Hq0jtMt+epgtaYAzJVNj+h3dXLw2moJLdlp9WtSZIwnyL7z5JZh6lhavP5DSTbEbZzDYhIz8WUfb
GPx7YT5gObHjAkN26NKZipVNSsrVZgeddMs6XPcR821X6cTb5QddVdHYVU26cplIb6rQv69bh+3m
bIDi89MNsOs+2DFMBpFWZvzO33pFoTmpW/eWQf4Knw13fYKBuvaeRPcuwrfK20ikC1Ucnx0gJmDs
CKT9a7abhY6Nw7vOJsr8E1ZCAW5SrFDcdsNNzBQm2uPWuxwmpuoHxJUDFU09D6kll+1GPVu1R5gY
O67B59/J0PU9hmyqT3FgPjDSWzz1MYyxKKwwBUE/YK3XrfzSskNJ0WmoJKaNGW8U++naWdaV4XyZ
JSrwUqprYU37MqgV1kkkSmxDDn/T2OGoAAJ+WFu9vYqFe0yd8NqqvLMz86XqkpNKLO3TKsxV2QFO
aSEHDs12aZvY1aoRDA/675431HYtA1rlpOvbckX99HS4aR2U+4tBr6PuBQgLPWyYV9OIA9TsfZgb
V38S86wN6t9wDlLmni3QwQTZDsWCVNFqRFIV4F9CsBAqGFuEW5ZuDVrXR338LfVtJMMKxhfyqDzo
CM5TL7vMWNQM2ueKJJjU6OLSepM+FGXB2Sp5L1WiLbKpDMWAH5W/UUpIq70Y96LwUeVMqsCpA4Dv
/tqPXKk2bF2cx+LbUlxXbar+tZa4hKg4Mo/vHl+ZVJOplZfJ2Ci0Rcb78L1sGLuT3rZI7feImVOC
82i48W6OXcp1+QeFRHQ5o4SWv2AO4Yb/3K/Tmt0o+xndBGKNkOxnTbiIURw1Wc2iz15B2ddmRZD0
NwRxvwLVPI9h/LEFiky+Dn22pf0tIX/VQ9kcrScA81poVo4UXQrOXpElvrGj8Jy6/iimQvPxNFnd
mddjdNgnHb83ixNhdp9AuVUXYBVmOIhsiVo4QAiP5Honss4EC9hoxGgt9vK/ig47/Fk+ElbAvC6K
B+QwxCpyPIgw3AtXy7SGIMz0WMzpVfk8z8083pIGUr3in/GjBXVkODf4FT5kIUtnTVrOCmScmwPV
GdCdaBTcf0goW/zf2mzDuYT9xU0QI0tbYZiYR2bI2+vIjC0+UhyBqMThJXrOjcY6G/GGLMbNgJYZ
pGd4PNDBf6DR1xlsJNXuQIbKwyKok+5tYhDYDEJIxjG3ralD33WamJ/Sj3+c69oDO5liOoux9qFu
oWj++TLK/nwq3YoZG7rvIOPaa4A9Yrz4RgGVlgov9K5oUxUqYA30K7pySwwJ71ICTAyu7uWRgGJK
a2/g1ozTL6PP8WHAy0T02151XzV065itWRgMUep9KVDSpGXQj3NJYkqsWfu7xaeUXXCFTqCxHPpm
+Fj/tR8nD3pBTXt8NyhoWU86lvVpw/0oIDoSrt6UXXmBv6+Qxp/hg9L+p11iHLm7lc2ovcvDNE6e
R9YUQqXk3JxLBsasZxEpZ6tk931j286dNJ9czSnkaKaF6J7qObzCXL2oiwtBnt+obhjdmb4Erqbt
5osBHXIjnv0kjbqQg3Uxh9dMMbzJpnJmcaJ05OPVGgxgxolNhrtYLtt4Dl5gRDTLiWoUO1837rSV
h8th7TsfACGJ4WUFb52SIwAr98Yv+YeeXRwwbB35qYEi1zdjRtOdJCzgT2SCR/Mja6huG+JtgTJd
LzeX6BPOxlRS7oIfIowV9pL+g8gNIEP237zrAXLQ2oVy9GVu8vbi5hyvF4jhGx0a7FSVOj6PBHuh
TBtt+qQ/eML46L7/HWrjOgmh5AwQzfRrblzxQIUYRce4ndnKH2SzHJJdY/Ma+2K/gmHwNbV+PE9w
2r6G0A1Emrmkfrb3fEChQyrL+BlX0OzdrcZTw1i7RNEwGwvzY4rYAA2cbViF9CRsV7spTu6SJXrz
u2KZxRo8TrMF9tlLDIn9OfBYwgcfMWBytg==
`protect end_protected
