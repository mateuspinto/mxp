��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����I�[RJhO8�>3(�̍e�]��;JQ
2b������)`�\s��0_�^+�����c5�A"^�<�a�'�o4\���S�N�tKm;�zK�K�4.�>(�i*5��nW�%Q��L�xH�.��̧��+#�s�&8�`�r��P������?M�U�|�\=��{&(҂~����A�B�,�h�R�Ę����d�])�-	!|�ȷ*h��E�� g���b1��L�X�b4(�I�����t��F�&Vx��z�)�EI%yYW����]��[�^�+5�j-��N���O�ם�zh���6 �'�Դ¶\`V>▱�ۄ;Ii+�_��:pƐ+i���.&���C�]g���*+쮠��I����@�xD�� @����w��3��k�"�)wX��ǜGS�,A_�z��g=��!�\�
�;�1mw8�R�t�r��6~�`4jvy��3�^��\r�*jc�JV~��?��6�5:�{w&�$�8�-\�������Hf|�8e�eRGT���13N�f|�5���d�Ew;���KoL�m�bWZ|�x�P�����-w�p��[T ����*�|�ܒQ�AR�(Sx�\�k���K����`
�r�1r�$��qH]Q��Z���Ba��J�6�p[�-�n�r�N�֙����tg�˷s;�6KRg��q�U�k�K-{E�F��o��ޛ	X$$��9�~�	��O$2c�O0�����mQD�==;��ȧ������>`���r@����R��wҴ�����)o66]�;H�6�!y"��r�%���%4VJ$���$ơ�a�qDЗ@q*���ݻ�`)4��DA�~Q���3��H�W�*����h����Fs�^9sIH�W�CB��7-!��#�����Y��Ѩ�LU��I07D`�j��yc��*}cK)_U�����}l���]Gw�^����ů(��c��k0�C���# �r��E���'0T�[��]�~DdÚ}G�H�:% ΖvB�:ۢ��ݣ'��}�k�9n�<&���%�š��5�|�z�+�ph�;y��������T� �E���=O���$LY���1ٮV��s�Cyݟ��y��$+���R&� XL���? ��.Z�Y;<)]C�Ni#���n{a_�D�(oZ�m1qzY����b��߬��J�f ��Et<5����k�%~E�O�K��Ҩ�q���[�����}'T�U���X��Kj�&�����7 � _[�Wj����Δ�t��60E%����$�<�JDn�y�V��z�Ĵ��w���t��`�w���69�?�v���dGj��0����t�X���v�Z�
�lA_�:{vy�	���r�z�-՛��F˅�9�
����v>�MZ���1l��2p��u2��f
�f�'Y��\zD��q�|Z&�X߻�(��o��;�g#�<��M�Z�b��h�?��|H�_�W����djڡ���Qw����u�g��MB�fj����ky�g�,��ń �q�]��c;h��Q�����v��䧦4&�k�U�Y���ѫ��GE�*]w>H,Ƿ�"V��+�(��q��5A�p��["�	�4l&Dn�T�c�m��G* !���(U���S���.�_��Y��kR�SH]5l�-C��s�%�
�J�����[�������2|K�Ӛ������V����)h�'I�O�'b�}'F�f�1�Q�|<x�қ�7���;Ř��Ơ�&�]�x�>�k���T��m	<ރN��8e����5�x�8k�^��Z��N,���i�w�^�4��&�!�Kk�>��#?[���1��u:���Ȳ["���Tp�D���UR��B��t�Ρ(��B�i�r/��(aD���]q��	��.H�q�]�p�.�)FGL���B8�.�����Oc������`�z	:�p�xEn�ŵ��=>h�?D�<���L4�K���>��珵F��&�):�率��"�N���ڜ���T��њM��T���.�L�c\������r�Y�:\�����U"�f�)U�R�b��%��J��y�`��W�Hت�5'%�*j"�����헐���Y�i[��U|�J-=-�Z>4������n�a�lYE"Z �D�H^�V�wm���c�o�	�
��MoGh�>$���	�嵅xђ�	`�.�z�ID���90?&F4ZA�.�
�d#%�uxk���r���+�#���$F�W���_H9uS�?j��[��R-%�|��}<�C�a�H�����tF�b���Ç xV��	b��aB�{H^�By�`����ps�`�S����$���^��Q��MY�I���������T�:�%�RC��5���#�}b8���K��_�jۈm%��1E�e��t��O!@�`��H�g ۊf�#C	���B�`,�O�gμ�����5J�۹h��9����<���g�9lN[0��@�h��t�:ڵ��	��S�@A)���d���K��4 2��]k��A?X��~	l�)#��Dh�Fz�rD���M�gKF4��ą�&�*D���tcfn��'�~{ '-ʪG@e��Q�f՞�iQQ�DWH��e�S�����(�q�8��YJ�z"�B���f��Nu�wỈ��^���ͣYM}7a@��n�MCx�l2�}[�r��\���s�����{P��4�� �@w�`܇������Ýn+�#<6����8w��_��������N� @rd7�y{�
�ތu�Eu�)�N����9�%T,������+��⛸Q8�L���Zיv+_E�N��h����Vt@&��_8_�	�E�
�M�����4�D��6y��`��|�"�y������aX&W����f��*�} ;/�-B��+Y��1	}' �
��R���i��L�UM����cw�44z�z���j�v�Գ��� 9��3����m�t�0-zk��à�kE�ഃ}E�8mۋ�𤂓�]Xk���@�E������f��� ��<��\�N�Ҵ��l� qz���S��VZ��c��ey3�G?y��$�l>NN5e���E�,�`�s�DG3�E>�(��	��'�*��/��y�����P�.?zI�RR���0Y�$��\} ?i��\�߹D�;iP:/�\�M7��(�]����i�ƶ�s1*�i´Ydfl��V�E� �! �uMt�`]����{�����C�_ݟ�NS��T�:mp�<�V�y���60���%Rlm��Mr(k��C�P7�	���v����s-���P��x��N쮍�UU��R�:�YAY����^6
�/�Հ��ԉ5� �u�*�T�3��)��xo���y�2�#����v�8��h�5}\�̱�M�fbM���&�՜1�ً{66sJ#�'6���ˑnՂGH`�����L�G{�@p:���;���NNg�Dk����=�Ǔybyԩ#Uf�[�~�-n������U_(��A^x?��/[��ܖ57:�6ie�oҐ0�p0�BZ�Z�DFV{�e����S����I
�\-������@Q�$�찔�4z������s�DV