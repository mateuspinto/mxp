`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
jIoo68qIfBylNjLC4pBX2boertQOUrbjyZRb4ae3WM61gLXRoOktYZ90kGEx+z5hoQ/+1HQmRx8i
cE2LBNiFK3uaICsuK/PwRMcxaJeCY4yVXVj+QfMPFJvawq53z5kAszwlyaJuiynI7h8Beqp9VlEy
pzX2iCwFY7OzIBU/q19ZC25aqU8MgIZwocbgf3WufHvjbhM/DLntOf2yTYu1W9bnpNWFBlIuTuOB
IWrQzeRM3O9vVvsj/Pj0Bz2NpBiIUwMcu+nejZu4yMWGezucGMfNYfGliSL859S4tz+tVmAPiBZE
PN2pGzFfIIuQp6PgKkxy2gLVhfiPYVXC+1vW7A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="QFype/U8SRXIWa4zsF0ksYYNBA6amGw2Hq4Ow5H881E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
Q+ZcTG0IqR7B9prz1cYiu7rDvbyYPpmHgDGaNnEeusmI39l7ylKhhK1gHfJ7N+PxijmG8KGfF5Px
Wh2l8XLSqQAqw1W1JAFTPfbHJTFWXgefYtQfYciMjh/TWNhA+Ps7kNM5Ff2FD4M2ilscfnuUnoSr
xywlcj/WUddtOTZa8xZAcQ08lg9oCS85xNNOV/3LB6X5ydJY+GqtSw6V0+ph7K8X6M3Z2fJCk/k2
6gM5Nz0ySiN0We9R2DQP+B9EjSRmBLzCpIHgvvcp0PmqbSGtv+4JlVkA/+lQwcjM8dutwP93ON2b
9bzzr0xL2WZ/QN1mbo8gkWOQEx6p653/wLDFg7JQLV8mlQI6aWCodQEP7Ydp7Yy1ZjLyIWLpmiKd
yAj8ZvZmWpvCyagnMkoaFqCd1kLzV1266QmBu34c+eN6OU2L5cRYqCOolK4MXBkgeBUWC2bf5H3K
+YKvEFOyIHaZBeO3P23jpOSd5pYbAzjBWda/BX0RnCAvgzes1Ib42BUa2W7RqbhQv3TmEYfjwH2h
pUvbfs0SskKuNQMIcHWU1LuRfAmW1a2aKn93QcLB8H6DppxxGHUj1EdRcHs6DFXxRV0EJKk/2DWz
JhR1MkGOI+RCoqOQ/XwTyLYY0yENXyyp/6LzVLkPPdLyrCDC9+7u0IATMoD6Qbq3uv4zU0Rbh6W6
8KDUINXYqoGcwZz+r/zvdNXoFQ96fJEoRWr28cDNq5xpA1Ldeg+gFvquKOhJGOgzo+5NGoYAtNad
U0tzL0+Ng9n3LtVTpyEqK0wcJ7MgCtgiUnCxoPRq6ivszj72Ite4eDSuoknSWr1zfwbE1aTRNuDc
ETXOXAZJwiIwZ6s4AoayWj2d2XvChby+HXHYzzDiiLjmrxTzF3M9xhzICCCI/nU1kamkoUiucjrr
ThBP5jwtw0Tg3Z8Ciq0yFyoE1T7x/ikLwDjUV4etpxopxysUs/zHuNOeRheI916CnunqwQizLKzN
P5nDSdYknX9qFgdGJJWZ6cToqOpbcST1S7fZxPSBEdF92mdoBSKLiDMtB7A3iXXM1r8I/ES4I/H+
i6DNQb1W+wvGuHfu5r6WWgaMM7/M2A6BBVA0lpzYfcJ6qrpQxAWqy30R9TcaYI6e10yMv3FV3e20
wHCv3HRsnRLIDv1gLaLMogAOMv/WiZL9DfYKGJZNXdzJ/nDdZIq/xkOBzfgVBB2pDysCDA6GjNMN
fTj19CFFoZ3u+RfGYzSh2YTzr5UmdRZmtR8WCLb4rYp3XmTVGul36J/HTkQmgFRsXTYbQJqFIR1C
g9JFx6ZdlbJoaGA6b2KMLdSPaA62h/K9S1/2ElzcOJQ5sbeazsvbDRhSDJJiCsXe0+taS2UWKsSR
opTiz14fUrdY+mnO68lmi52jJdj/qblFSLrfjJyz82HwPZBKHxVEwnEzMoizl1pUO5xzga+E/2x7
GbSbkSW8bMUHZTcWVjc7uh+z4OXb9zCFKKiSJQN8qJRcY9+KcQMUj/VD9WRI7v9lMx9uCZd5Eonz
pA+EAhy2/mveX21c228IW5TzAa+xT9FLneDJsseScIT4kI3+2YpBsLxq1ttaKp28BwTU1ESGulZv
+KyPOLAnvAZzqkZ6WoIHCnWxjg+YEFC9zLCbk9UFau6Tw2zoX2P6RJ3liO3srR0kdcpMIgwB7EO6
zw2BSA+8em158ALTwvn8j22zvNBEqMICRptNMozBb/S3H4E2tOtUN8wp+CS9sy91QlAiA4SnDfHy
9qkOtmUi7R1D9sel8qwXJJpZy+i2XsliC9K458FHAEgTcxKNxDn1GATpcBfSt9fHL03jxM8NUzNL
78f2HQiefBwYsH3dtiY2NaXblAxegpoUVzhto4CwonbOqpFhPRwa+QE3Cr4f36Chqz6xihl8M9oo
7nStjuNg5WLZrZ1fAAc9a4OhV3z4JEffHosSzDIHp7s00uCUnuaMZWSRwKin1kNwfW+hTabi1Arf
Y7NrIUPEU5ULpxtdDwzNdEt6DOoME3GuA/p9AskoARrlk1bNzpNEcd9SavP+4ktv+DUHNAmlBBN8
4VRtnV41/9ygvc0xFIqV+DlzDHVYgqLN32oTXxUB5HYZxkL7l/z2AK+UGm0U
`protect end_protected
