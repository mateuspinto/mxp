`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
xO71WvHfQz1Xj75GOsvgs5QUcJWfOg7RaQQT4fUrh6pQgm0CDA3Nlcpmzq9dFvttAhMS2KgIj6Rc
oTZQiKgwEYtX89ZgokBqoJod5Er1s8ndvaWt7uw5qYZhrYarEG+E7UWz9fuoOqrIVZDNxhpzxyCX
5iGdWfAVejUIVF1uKuy+ey/gXPtDuizXSP+xu6ZcVvbFAMFKVeoQPPofL1XJ/NHmZ3DXOpvvwNHP
GA2yyCbgcFByDmMo6R9nAeYlQSYiiBzaytjp9l2ckSvqUIqDDE1RPdIxiQYTzfCs3Y7SYiZ6/13N
K20LrHsfYBOnlhVuxb0YRjrTfMG9R4pILnyxmSVqcuSKGtzmVlV1nsUBqEv7QcuzuzOdjRcEqdfG
F0pSnWkZllTGZGdRUBMTNs4h+eZKciQeQMiMHDZHHQy8sXt108wX6acoycKJntkmOWrD9Kabeyj4
Ce7gbcOjFwvNb4niRHTwQpMGshLp1Z1eDT/F6bjqWb49sPvCPqeh9Lv21iXYzjSkEkfEwbbOSTwq
oOmj2X0Hqr5G3u4xCEuxrWuhyW/nZOLjv9HefR4FNqK8ZCsakeBFF/kuLQlQ/6S/dEuhlbeOETR5
pjsFrYo+0NQFNF8qctKr27FiJLzaIF9I/Lu1Nha8FNrpCCkfDHbSpEpsFIIPkvXaDpSmPQEuwl+C
vTRHPhXHIZDpmz9f4tWf6gMwWOkNKLdZsjFhm81G1hFDjYz+yVsCHy4yFXqPgBCbCuZ8eeMnifE1
/obKud1n9877AD1DAFslxgLQD+x6wopzN7u8Hao7HG8I0Mp4BUlpYOsJSjk9oNwOrzvS90QDz9ir
nWGWBy/5e8FX7xWydnmYxvtVfPjGezN3JgT9GaFpu2CY8QVgL5whkRSpsRs3LW/K5Yd7UG1XPEBT
PDCcsjLJ9k2as9eMtEKxP6VCZWSxzIJwKyzz2pzwaK1bAww/X15cMIY5gt6yI3bXEhgPfPRQnbPg
pPARuZ5tTQe2cc/KifK7k/n4BQMOHUeTZLmi3qaDnhjVBOXQtid8/BsT1zv6TQpDs2jYeH+HubAM
iWOf0TQW0lYBfYF1vZbbPHKCemN5Lhe6XIegv+GXdNv+q4A/cNu90lSNhIy6L2e8vUSNED67wrVQ
KFXUwiavC/U998bYG2dWiGNFPdiPhcHFrEP35xKRjQ9cokDYjUJohwIK0qhbOq0YwGwM0P1QxmlE
W5VjdUx21QLHIHutUIZFWIl2cS10Gz2N/qVofcwEn6WZ9VZGsvTktcEOSmaCES67eHj0fvpJlQ0m
LnSP2wnBNy2PL0WtOpznnfMHfKYLgzseK/0Vw2BHBjM5ftwa3wpBtJ5hL2wWkLWQJ8+37F6Ai6U7
oDwi2AQ/YGGcNV9xs+rmNkLSN58fYiP1RBKXHu7NeBgS68kb2+bvs50Q8r1n3mQvmo/shEMVe9fZ
p5kENyKf2p08tLfuQMJmScVwhZqAdnsjT3OFU0ZDv5POmZuk+Na5egg2JAP7AXe9o4uYFHDlxsie
QYzpVALo/CUjVXA+ba593qrCf2820j8bB/GwDD0MhX3WBiu2BO5OwLB6L/NFDlAqKAB4i5cyFVUW
HOgaKs8dAxY/hIem+pX6VeLhKSxy45RsSWcmLNRDbqyH/tqUWBnTkq0Ii9/tDDCaLdxNkVwpJR9N
y39Jvwkmy+8hUeTeBQa/Gkq6eLT9pvGadxXq7ijcY28UyXFSLECJtN9dE5rFAD7C4dRyHalt6QsK
DGdIAeZ9HuTrdf+jB0R+8rixhVMf4vOvwZCL283Wn5V4d6fbgkeVBTr9KU+SdOjS507V/1sTdGb2
SRThMXtcKYOCO96lV5KvFGSQdIlL0K4TGUVgZ69Mjwbx8Hi+PWRw/0Y8IZ1Jy8eGkcEdTkxEveV+
4BDxggZ3bT1zMkTo6SRhqK0kz2CTI0iEcW+tCpRdTz3XAJ2yezwJbRgdpd3TvvkDoFu7Y6iNfObh
SS5zY3/1f0XYLr+XIyvPF9/RotYJ5AG7i3FQ8x9cKcnztgzQktdoaVNvHDYZuwv75LqQgrt271F+
vQjGuabbz0VvwxOvcjbWU6YMQ6weGmxwv6GTzdKbKOBCbsVrgIqvIM4bTKKPDRTlgZ6fe+1IHNaL
qRQXO+lidTlBnebV/JxgNVL/rjk6f4lpdGp7L0157kEgwf3xc4V8QLd2smv2A14sbyIxHwdD+UgW
CwXCP4HewMZMphmRF3Oy8FsU0DPHZKBNZZ91cQp7eoq02o1HCVpANx+A+3JZZTN5sI/cE7iWFzpr
ctTJtquPHTGy4k+ZhBjQ8H7qFE34zIyXG75YoLBOA8g4waXfEGeHHV948wmd30YhK4S6bAngEFkh
zV9EAC72UNRR9SRjigbGqcJ0ylwl9NOcMyHsfxZUqPE6I5d0p4CwjMY5BcuPgQmOY2P+n7bSQ9m8
c3sJNDkastFqbmBOJ39trx0B+TXZ2tltoBBOQdTXHLsM/yoo7vO4SfqDx5eUxWGE73elWkZuPUEL
c4ED9AA0R2lY7lwC69y4HCZ4s7lqmgQy/GvRvNNhmXiO4aqDwauIn1DMFyqYuLiDfSwYF4DVZ7Zr
p9+3di662J+LChbppGV4BOWmc7i84FCLCaq3q4vnoGtE3xvYKFLY+1qppEwSHC1lt9uOifNP623k
bOB6Vob+bjITRqqabJtJdtZNAJ1fmiPuyS88ZpnkXSjvKPCoyMFojAc5VrcI+grNVKfQkD6WQIs4
fsYQIM0dMAQgp7J1qnQ5D7kQ+DxokQvAVlLHeGB6p3B/k8+CCN2gLB9Fb9xeRN+DJkUpJmD4S3im
KN4Ui3JAfKuISJHUMbYnfs/vfmOa0QVJW77IpcmjhorwoPOIQBMRu/9fOL69WufZZ+EhDJTw4qV2
RoAIkyNrlMKAuoycuJ2dkxjlB1PvqcaQFln4pVYUmEJnH7znWVNzJTDoWKcUfsb/zG9/wgYEFoR/
YfQYEqblqaqKaEC3PE2FY7CMRs1UgkKfVx3M02c3Cl64Q7VBWcYjuFS+q8ioZPRlJtGupdB6ATU/
CiAeSsf34ZiXmBIyq8R6JxvOai9cEViieBZxYiwJiHDJFoKRsxhzryiZaC70xoq66FYsUyIUBOjR
TX+CI4H+tLd8Ko3/ns8IVuNemX/aWmL8IeCFCaMfN2KaX1mHe5Jq3bl9lhPEM3HUSljIqYSPVnIM
0p585mk8ZHeKA3/gXuKeNmy2NsptO713wO+xZp4DPxHGbSN9he94PJY5eXBuKhJYa4KkiztdfZU0
T8L5qQgianNehQ0rnG394Xp+deFNYB8Xq5GcYIfVWJwyl1kbKLi16Mem3dv6yoWpuRGKV3N11DdM
Pxx45SnajkuEnNMr9yZI7JIG5axTJ7NOibtfjwEv/0x64urc10iHcAiRby01Vm2w7u05rIvwoxfG
zx3T3xAEMs+9Mj0ROlxXzKYl4c9IU7WpADvT4SsFfD/A2yoJtt5GqsyiYCDaBF5BjTeYRNLiK1X+
GjoqxdKzZ4YmDxYKEJTJU182pIR2nSiIhhuoKsVfqFxmuCf2t3hd2E+auX1m4GsRTOKuqaxo+ttb
t5sz8Gm8r92JQRfekLYX8ltIVpvmOoV9l1PpgHavrLqksbBH9SLhWUR00OZgThIPZzLj+htOIb89
3RNtWfssGQ5PaWotmsPy3YYEaNQs5qvJpjj/a4JlRxf7yp5jnKixs4bUcYz7wDBzp4ZVwsbtrbyI
W0F9xZwIHA/cjsByfjqkveXlKwp05cggIUZFkutagSuT89beCUZuHG91Mol4zHDv7xLX3Jonq1C0
TA7CfjnCUkZxW/in7qjVPR+A1aKOMwR28l8pgKKoY8JnAGb1WRKHRoKgKG87afLvGkJG/3tJCZOS
96QDczLwDQMXmGbeO+7OF5h5FOpHIXeAw4jKz/t04JX0IcANO1Fpo1KiFnByP3YnBmXmZB4UwbCA
eVwg4+rZp1Cd40m6oHdBF+u9MuOQCdBaRtVsX+RhSzbR/XFh8/zo7SC5LHy6haUyaIOaVNpa9fzR
kcS2h4IDeQ6++eC7rRZCh6xKAy6IpI3JvrFF0nwsHFiD7SQIIU+gPpS0CCjsXNNetxkxAoKRsAQH
hNOKYbLNQVy0glXevOYVaPQAFmSh0LjPeeGw3wkH/VrLC+dNivGhxQtOT2rCl6+mkutaOnsmNEfR
k/Pa2fzNMucxRnGJ3+3d51rgUgqjkwNeMz8BJlmLJd+pZT6xFqK0F3X9dbdmCuM5oslCj3zXA4GY
wnHc+Cav5MCusk2Xxp4BQ7hJHIXnKzVsPudhJHLHJ72EFPx9kWKJfgjnQm1iS7cMiTHcWtegdjjp
r0N55mlk+jyG/oaAxNsDpf7lIqUVrZywYBuukUV19Gj+iKZoAyr6z8UxmDykizyCUIGRZWt8Flbq
+oGmezpMzYmVmwBLLhk2JlFwgX86V1wcluqTqJKTrEUcarLKGURm0fi+YY4ftfloHwq9mjUyNUU5
RduLPFv7/2ygZOVhfLyRw5WbAmpHcFSZINu0ppH3CyWk92AUsDt7dhChLzkbQshiWhA7v8zo7rNm
0Jf7uSNtEQKvHdCAS8uw+02bZJ2Wm1AljoTGDVwz1ul5xS3Bz9ExZCOzZUoEisSqV7GsW4qU5uP+
e9GY43Z6n8VCs2h+iyh4547EKDudkD9a8LwM
`protect end_protected
