XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#`ʣ��l��7���k�R5� �$��%�@�,M���賃�1"K�V���%Jv�v�[��-U��};�'#�EP���\����h��~\S�ġ�NFɽ�l�+�B�Qq�F�7[��?B�4C@,1�-���a�U���E�E+��z�^�(��m�RR�Q$v��X8�XdU��8�y�h7�8a�;�Z�L�M҆j�8V��9�Hq��֧��>v�-jh��ֶW M�t��J��(G��d�����S�~'Y�:|s]��j��/�P�1�)��J�^P�C��gàd}�4��u|�
�x�k�B����L����������1��c�c\��l��a�h�
*�|��V0�%��5�ڤ������t�	�K���`~O�Q r[�2�� ������Q�1���-/^�B,C�2&*��7�dM�	U��):�|��is�l'W�,�䥑#-��f�6\�æX]��	>g6�N'K�����詜Ȳa�Sd�E��[��W���*ƕ��X�v����y%�b䃧&B�q�s�
�4utDL���m ��޷j���>�`�y; �VK�� �9.f�L��MF�ե%�0c[�9��V{�q2�z��!MO⪴S��uҷ;�>��n[" �������z�D��^
�;����&�26�6���K�X(�vrG��s��M���K�Pk�3��,sI�&���/~�6H���%%j�D"�M��K9�O��= ^ݒ3|�1T�izXlxVHYEB     400     230��&i(e��[��(��<�TU�˝G�H]6��f��,z��u6��)~s����q��9M�������^����έ��\�ĩy3_J9ϱ�OϪF��=wƿ�C��}��)'Hpm����!������z2�%u@�;�@[Uf%��,�Q`^Tǯ�)���k$\!��]�%C��G�0N�$@�z jy0����$%X�V�U�̱�]� �an}'�@��l�ƪBc��/�H�_-�k#��u�x�iŕA�L�����Dd��v.T�B�h]�,����z��ˏ�����4e�}��� 'a��?5��梊Cs��®�a}�Z�k�lǆ�7�N�A���5
-�i�-����g�Y?�����/���X�	s6K+��U��q����i��.l�ODظiw���()�Ds���Ҕj�p�J��L]�|Ǌ"�ٿԍȢ0QׁbG����0���>���?ܡ�ӥ��n^�����r.�K�:,��w_�Uҥ���9�ª)'8�\+[�3��*���.6/�	/Y���� u蘀�����BXlxVHYEB     400     1f0�v�F7!ci��`f@cm�NW��Jڳ�r�ϯU��k`��<.�°!^�8u��Lg�Kѧ�Z6ܝ&?9|Y�hA���/�j��/���Uc�w�mǓ� �&�Kj��|u��ץ�OM�Qo�l�)80y�Fh�I��ͼ���zU��گ��{TUb]4�c�p>�9*%,7�*�f$M|�,�
'��$�&kf� ���j��a���}�_���Gֺ��}������Ca�+.@�ө�S�Y�|B<�1���2(��t��0�MGPT��ѿ~z	N_�L�g��[L�,�À,�$ Y)����5���c��Y���F�RY�-�c:�=�Ȓ�^o3 I��Q��D_���d�f㪕Nx�<�N|i��^�j�`��-�����|�+�s���=�J��H�{1��~g�Bu��Ȼ\�FZ�X��B�l�w؉:�-����%hܬ��nn*�v��y �v����v�	��A���I��m��k;�����A�XlxVHYEB     400     1b0״n�0��:�z�u������"^�a��b
v:�v��D� x`)��<��e��m�58)���FPG�㿆��p=h&�%[;$D��W��.djo;1p�SG��'d	�s�a��Q��m����t_%:����Ll��{P�wm zg���K
�a^�Q�-��A@'��5{�y���Dm׽�&N���������,��oq�±�@�ċh�h��&Ō6�&��cǭLWz�s_�8	��w)��4���ݓ�I�8�gޔ����{v���.K����Fd��l��x��%y��W�ν�>� -u��N����C��4X@a�I��T�]�,0��OM�x���!,�?.��8^9`nfV��r��+՟P?��o9�����g�A�T���Ρ1�6$��?��WGWT���ڈ\�����X֝ ��XlxVHYEB     186      b0�c�Z�xަ�~��SQ���6u��+i�͇	�8uf�v��ف��
�X�I�"��0J�G�����
�U�)��r�}���i/�a�\*�[�`�)Խ���\���
W+��C2��A�?cz�c���U���bT$m�Y���v/�T���NX,�ʳ�ѡ��r^Z���!#%