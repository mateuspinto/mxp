��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���\ޓPR&� ��0��.m��D�1���X*]k�<&Y6�G�xz�ǻGp����-!��2�?nb���M�]V��x�5���S�I'�:�VW?��ϥ�1Ӗ����
����Ll�&J�4V���^ȩf�oԷ�����Z\ݸ�iYn��O���B������=�6�>4$EW��;5�A��"c_����X��䃛aEz��"N�+
oox�
�ۏ�Ԩ�7$���l�����Vz���+Q�~����::x�T̏�0ڼ�=��㢳�BpJ����ݴ~�b���X�!@
p�"g9z␥F�mdo
�J=���QH�	e*ۘq6S��t@����R��A��iͫ��{!uE��Е�� ���#Z*A�[Q���5�@�\���4�}��BG�p�H�c�4n��j��dQ&���Z�UF��m�:z�}	!7������]%Ob�P�-��1��z�� 1�s_��wu�`�K����kT���cG�EKF5�KCI�������=�M����F����V7,�}6� .@�_R�)_Xu'd�po<���qS� �#rHt���m���}s���ANP4�~���`fC)|�S;�J�-A���`J����,�"�嶵~�ɑ�9��|Pa�W�I�$����ǋ��7��z���H��'!-쟕�&�!d 揽pT��V}+�� \�FA��� J�`�D�Ǝ���Q�?]��OQ��y�������63��s��J'|^`�t"�6~�Լ�'ͽ�NKH�q��1sn�~zQ���7��Ƀ�&5��E��s�Y��l9FO�$�/�R��$-�z��Y����������7�b����!�/���|����PD�$��g;���2�W+��������y49��߀)����U�t�Xٵ������w#MN��k*��4�r:��O��]`�TU�e�2�`d�O?l�_:��H��d�9ܠ{���
�)j�|����o$B��撵�	��zBI���`�T����q��I������q���F�
uJ%�z6�F��w���YRo��̇Zd�5$T���c���m�`��/MFf���'�!wj� �k��.~W���P�y�_}�wg�[@r\b���QL���U�ԕg��ĲЪ���5�0�	Y@�y����É�S���T�������ԕ� }�8��A��2�F�� 縱\SK<v��ũD�}I��>�P�r��}�ypv��X��T��"RG�%Ct�Be�,'"_��KwS6.#���YE�O4��`�*&M��Z9�T�����q����{EA-#��h�cn啌��
�$S��D�#���J��1�8�It�#��@�2=Ͼ�]�9����:��\�x�A����|�@aEw!P��s��Z�{C�<m�'M�	K�e�tF5���dwS��b����_��5Xo��YO����}�&I�8���b�Y(G�p(������XI�l˲����{+퓼�J�7����~�DgJ�:�z+ǎ�S��Yb��=o�t��j}׻�'k�'E1�$������+Z�L�w0�$��xI?���N�?�Q ���Li��U���G	n>Q�nGjJ�E!����D`�� ��{|5��g������s�����Պ�%׻ӛ�n_JL7�	�/û�yǒٷX���"Mc��;�(����jH�U�{cb��Y��ŀW[�2	��@l���9������a��z9y#_L���Y������۠^��,�ӈaE�AO�c��F��" �\���E3y�^��.��K��bu���@�I�'�s�V�M'�{c*�B�kȥ��k�D7I��Y�6��Q�n�wB�V�E̖K�����:�#�]='v��튌�tb=��~el�� G�
۬�E�Mq�a�5���S�9��sŦTzE�,q�4�7�(o�~�Nh6���_Ô��$�d��ơp���	�:>.=�LA8W����j�Xk.�5�faX,RS���k,�eD��ݰz��<ܳ�f<�*��f|�5��I�)wmnpjĮY3;��ОO����4i����r�����U���O�?�Ωd�Jqo��*1ȿ�����˖�|�Դ;���Ni�n������5�#��qu��j�����)���&q�[�&J�F�`����W$�x���=='K�*��K�6��w�Wj���z��`fi�$u�L�N
"�5�����b�����0��ۮr�އ�|U\�3ȩS'�	�9ߡ��T��҅%��QX�8�,~e������ۇ��:��CѠcނS����)��U�G��&��zʡM(P���}Ӹ�^�m����Ag�����d�x�jP+�ߟ����H@IB`���T
"���ܢ�X�Ϭ����
��S�3Z�q��d@���o0-�|��P>3#�퍯���8��&)��ApQ�a������ƪsBĊ��
M+	����iz�$kc;�D���0���Um�?lŴ��O脖��a���-��O�~�����%���Kwm �Z�h<����GUV��2Gʂ9��Z���ek�@p�	��;O"%w�2|d�D2��Xu�!1mdC�׆܂�5������ �c��5�#�M�����T�W�~0E�1��E�I�N����:�+Xѱ�ߎ8�҇�#����I{*jN�ZY�_�����ό�����ޮK��x�M�n�g4N��Q�rr�	}I����l�	Ո�=��O<�������ez"l�8�DO�Bo��`�?����Xa�F�x�
>�M(��{��^�	��2"Z԰��y+g)��A��%v�����5s��[1��p��T��m_R�?'�:��i���1m,�\�7#o�7��5�ڒO��)�=2�"p"n��/] ��$'��'��|�M�	�����x��q���^_V���&G��U����IG&!���P�Z����M���Q[)}��#�^
&mF26+Y�ۏ����n� �R����^>�0�u�Ŋ��?�-*�~���B�l�tVՌ,\���Oh��W"e)��I\2$/u�>�݄U�,��%tJ�1w�Y��gs�Z������ºub'����`����5C�3ڸ��&.b{|

G(�ZqzX�:S��Qg�[_�}�
�9'+���zE����n���,�ݕ��z��_�`N�m�/rh#ν#J�ƅt��c��U��v&��%�<��������ȱ�&M,l�[�g�r4,��?r1Qy�4�n��<�;�M�?�����E0�z�Q�k�g#����L7"Uz�0��;��3;���0w�[�a��J���^��{06c�DZD�~�nIʭT-OH.d
����'uH�"��PȦ )imA��,q����4[�n�!ݩFm�����Ч3�KȦt�$�8�w?d : �Q�9�_��SO��(��I��>�Ș�]�)Sٚ|��]�٤��$Vn��=/oj�Q�g�R�����A�![���-D�\��B·y|�'�RU3nnnϨ�i����?ym/�Pj�v[�0�1L���u�I��_�
����+�,�^w�׳�TJ����(bO�jԄ�������FR��Պ�ݖ��sժw�� (�\����Mg��9>6�퓓M2�5I�
�-��'X7z&�)���A�"�T`d���_ԛt�*��}�����b�/�=8b���x�Y��bE��9���e�/1Uo�gb[s�w��a�sS�� ���Q$��NeY�񰟗���b67��D%��^V|��]�	x�m��n�뗶Z�HZcA$�Sw�ё��氡T�YO7��'Ɩ��ܱ����1o��5�~B�.�԰�w���8O��s�I����o���Ю
�w�v����rw����(/uJ�:���� X)8���e�}�&?A#�Zj�O���1�dR�M�C3.Z�����n���E�p=�m�=߻ґ�����g�Z��{�k&�w��}�P]��ÇĈ����n�ϗ��UQ���������;�C���H�D�]�+]l���P~���܊`�}��Ʀ���j�7�c�$i|ב�}<1�����A�Ȧ�D�?�����c���B_U��s+9���7��Ʋ)�KV{&֦��+�1$R�l$��� �b
��J/�X��UB�\kc����h�)0�9��&C ơ����J3�
K��P�j�2�3���c��_���r�J���[A�V;5����">��();I��\�3s�7�	�fb4Ԓ}��+Q�;A;��a#����H�<'�T�{!��&w_�I��)e��FX9�Y4NΏ\?�m�h�ҭ��P�.3�\C�m�Bye�u����i�BoW�դ68J.�+�B� ����5�ں+n�a�;_A4�7#���S2�vއ��|�rIg����|�� ��{P����q�i^R��%�pͻu�6��v�D׀t`
;E����j3)�����V��#�s��:&�+_ؿr��g�Ȅ~M�N�
7�KBC��^�	�j� V���>X�����::�{߱�C�DsC�� ���m@�1��In����bȻ�����k�[�ʏ=��1�PT��L�H��$fYoY �R�$��H�n5�&�A��g�~ܫ�o��|�;Xa�������6�#!�6�4}$:�õ�[�!�g�W�-��MK.��PU��yڴ�� �1_�J>!��Ǭ�{��sï�������"���1v�C)�8��)��U��!)=2fG]��rY(�̣h6hR���h��P�8��CGڿ�O���h����5P�����xR�!*�ӤT)��e�
�l*��g�7��!�QnqYY���_=W��Zsu���BގZ�bE�A ��R(y�5*�G
���1�.9�pdy���G��# #P�=##���e���qFÀ^,v�8�)�s?�l6�m誠{>�C��II���#%�G�o� !�f�4���:��	fl[l��+6�|����*������rO ��_�E@Z�e�xɋ��*v�#��I8�I��{D)%�22�%�D���Ʋ���q-703����p���N��Q&7��G�[�!�}��򁓩��0�g'���K��u�9k �; ��nL���3-*�{~c1��o�\���z"��e���k�ݹ��r"L}�6��g�b!���5��}Y���r�ro���VS��S���.�$J�y*69D�ys_���<�Z��7�5"t]R�b�b�!�c�{�a�m�&���T���@5@������6I����$'�U�~57U��梧z�'r��`A���Y��p885PQq�J%#����ֈ��k*hK�����VA��%PY�� �|yMdD�q��[�*��3���7�y�����k�v`�nm�;J]�:���,� ��;vt��ʦ.��&B$>e���|��(+)I�
��Vixڅ�Ǉ���-җҩ�O�un���٤�-�J�yj�h/<Zd�Y}�U��:�D�]2T�ۮ�r.<3�,��̸7>]\�:��s�J���tv=�����њ�&��i5-�O����G�7�=��d�u�?�/ +-P��l��L/a���ss�J 6K.DS����o���;�OZ݄���wA�q�r��''���43�&z�.j���	eg??�݌�c��>�6�F�B�����J��Y0�l\%�^�
X+��h��_�=8�q5���uB��~���03'���v�O����с�+��& Ы���HA��۠u8��E��ǔ�&����O�v?rE��/6t����2#��Zc����O?}����6���v:CBB��R�^�4������i���K!���~Oҧ_��oĎ�y�
.�!,(�T!A<G�/���6,E_�������p��\F��p���ճ��ٹ�9�%��.V� ]�<�����g/���hgt�w�1DR�L������	"��K�����.g��=���er`��c�y�hX:D���s5�V�]���)cd�y
�N��$D�ց�r���׺���Jь�1��[߽~�x����N8j^��oM�$���8b|`���.�8Y���,I�Qe�TqL�<*喅b�/&(��z,(��rc�}b��c*��Jk0��,�k1zM@�C\��L T����̬�`�0��I@C�Q0������g�g��^�>���v��8����