��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���]X�FwC^�_\6i4�4�ss��Q*iWģ��E�����~ �'����Y���wS���_�[�w�n�W�3iqx�vn��*J�;��g�$l�=l�+��r7}�Ȅ�Z�����w�|��F�
����p�Vz�P��Ϧ�RN�h��t��^�;�d�+�>.N�@�Ѡ��	����N ���8ըy�������v�Q[�Q���s�2O��LO���)4��N�-�r4�#{b}O:U���h�qp�*�M�G�J���ٶI	��q���@���b�����Zc,<jv����@�#8�N�28T�v�����*+z���&��B:��bM5Y��Xԫ9�Kh�/��,���t��]K&p,�4*�.�C��c�\�#@Ƹj�\�2Y��嫳,�-�%b���:�rl�t��Ä�L�*W2�>��sR�E�W���VȲ��U�"� P�C��(�	�ql�F��*��/w��7Zb@v:��YD�^pe�Fn�ut�kx!���R��I�t�?���d'"�(�;e4��j'~�T��k����W.�r������0��m�AA�M���b7�Fl���NQ�v�F���_�=膴���o5�������c���l��߯ ��fv��� o]%R�z[٪O�C"ױoz\-~�dУ��ڤW_io��O�>I�S`��SY���F�t�g#�ɿ�MP�j�N+��ۅV��p�M��8eĄ��
��>��]|�$��c"����kY�g��QW�+h���ڤT@�S���gr��}n�F8���yXB�S��",��RZ��Z=�zf[Jȯ�b��p�0.rN�����Xl���\�8���^ֲ���彍7�����AI��z�Cf��f\{9k��л��O-����>Ⱶ�� ��T�l{�Q�61#v�¡W � �e�V�hV�1��d��@��R����&ۺ�j6�h�M���ͧ&�ҷ`(��r�Z��
�p�,��V٫E������C'�~ �����e�n֒pk��l	p1�������S=< ��Ŗ��M���Q+F���x=_�!����!r�h���f��K��e��������Ԓ8c����^�:E��V�i߫{'0�3�(.���	4��Af�]�D�)|˭��s��(��[���W�QMq&��?)�]x61W�b�#j��y�52u1�GJs�VW��TU�;e�s���� ��6	]��U���wIeׯJ�.w�� M�4 F����R��d\<�����(�kSz<ϙ[|�|�I��@�O>]|�VV��}2]|���n�%�b��=����[�m�[��Sp���egn�PAEl��m�����ԓ��|0��И���|R�قa�+|�fb4�_�5d�۞�@�s���9t�È����Bi�<u6���Q�&����@�
��m��;%��F�IBb���W��'L�Y��D��v���s?�q�+���STe�������:�+�y�'> w���8c���f��5�Y�y�L��XIڔA皌�ʪ\ ܐ�j�4g��>a>����m�������
~Y�]qKx(��|�Ҝ9���WC��h�uH�]e�3pb����c�q=V5�j�l���d�g�2 �@�L�)H�B�WI��.��6l���Ŀ�7d>w��a��<���weO����dь/�7�GU�]�r�z�������0^|D�:�F��X�ڮ+p
��?^�V�|[]Ezj�ܯ�,��Uf<UM.��<cH������J#��Ln.�r\�l�°v��O=)�9?�
��V��3�;��X(��A�q���_����0������Q��V4[�&|�"�ް�ƷY�v]V�3���)AdB⻒���^�(��L�Üs)Ӏ$ߦ-L~s1t�(x4��Í5R���@~7y���"�N��#���D�Z~
d�j��V�T^R���&�r���k����D?��ۆ,�c�.Z�@�B��cg�,)?"���l��fixƧw�B�s����W�_��q��.pq�NI"�U W�e�B`w�;$�2�<�նH���5���I5<�e����sS����Ej@��>�*t���|Q;�y�>�K��tE�4�ymy�ͻ2��9șCt�E|)��&���P[o��>?&�����6��E��bs!@��
ۡ
4��A7��@� LH�&��D�t��tj*r:	ifґ�$���ߪDq��,�d����#C��v�EǴ�G3Yk��=I���s���jl�@�k�Z�+��e�_��>�U+HM�X�̠B�#\1��[�&;I��Ĳ�
I�ּ�R���7�B\
@ng*��ؐ�>�f��u��Z��E!,�O�h�]�Y1����a�?pXNJ�ۏ���z-'��.+/�Ґr	��5]��������!����k�|^������%� P�@��9[)��5���^��\��t�
Ep�����ר(ō�1h��R ڭ��ao2V�Z�_��Ⱥ�v%.�h���=�%ߗYn"sO�қ�8D-!���j۾���3�]S��+��~ �/^���p���>��Dء����A*���MXS�O�?��7Ý�8m+�*)|����_\;Vb�1���'���˵�L껪v�ks�fp�d�U
�'?�����꘰Q��3_����r��T�g����똝N�f�z�tE�$���u��^N��ՙ%��̺�����cf<jXsii:�Zƾ����MZ~C��(,o;�Q���_]GP������Z�H/4F<�n��r�wrs-C,�M^�l>�Vo`�e2X�ѹ�(,��^pC�'��-�nuƹ�0K����a��sĽ�Y��!��lap������r�7!�̒�X�Z�@F C3Q�Nܘ?�I��ߘ�/�����'u%�Z���+�K�"�3t=C۷�JB��S�g��-�
? `�_����E\У��i�t|���M��9K��t����EPB]�}@?7[T �D�s