XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}C�?��
�Sj�s�PWb@òo/]�$@@-��1�\�6����1Y��/ZE�惥]�*cm����d�գðW^�A=7��Sz|�4΂��U,�N��[������~6E6��x���+��T��4�6�8c�ԝ�������:��k��A�'Z<ӛy��ٳЌ̞�ʥ�]�G}�+� �,E$��vt�U�sjY蹧?�����+��D��}��W�����\?�2�v��Ī�9�m���7�E� ѿgɚ�<�/8���WJ�$�u��GY[5�mZnA+���1Wqc��(���Z��u��QP@�y�1���:[ nƓ=�m�'�����a�^d��NE����3��j?A��i��)���2��JUE�w���vc�l�; kP~�B٩E����)|"Ű�u�
�d���#�#��j�X��(ň�vo*%r�?��m�:�X�j �pc]��Ӄ��dי�'�|��p(�VS�����5d8�%��V�()�7-�+��d���
@��Y�f\�N-�x�-�+�h%(t�Z|ꓵ��-�1��g�9�N�_�/�����mL6�[^����s� ���ٷ�|'��H��z�џ>��B�����q���g�U��,�W����_�����?Y���$�c��/�=ǘ�����������)��:EI�pJ���L�/%���~����Wg�(��8Ӄ��n��l̿�%���F���)���B��&=���.�-���$b�Rɓ���*Z�ș 톦ݮ�g�c�XlxVHYEB     400     190��y�t���8ܗ�.d��h���W��WVX�׋)�����]2�SK�>�薡�`x6��ai]���3U��m^�ƻ�B}��]ga+��}�Z�KZ/t}t�� 
!Q��~nlt�ђ�/���l�/
R��2�������Y�Pv���\{�$+�C�g8j�H�WU? ���縫Z����!)H(8��
�!�n޾�{'+��9J���ր�:Q�Ç�����)(mS���c8̾��7pe#W��J��x��3�Y�-��3�m wF3�T2d]�
AUsQ��h�pP��0�9�M��u��E��EI�����U��\:4��G���CF7�u�J�TfN���+cࢡ�C��]�O��b�Kd�$��k^a�?�b�k�A@U��E�"N���_i�w[XlxVHYEB     400     170�2f
�w##Z�S�09m��zΥ�T1�a��[�I#8c̎x�I�v/HQ���c����N���O��P��>%�'��(mx�=c����c84�bYk(�,�\v�5ҫr���lXAm�`���I܅s�|���𮶙�ˊ��f5�!R'��f�N�.��ă�����, �>�t��}G�@���a�Qצ�~��هH{n�$,Йc#u� }�k5����#�Fx}�iֈd=��FQ��|�u(��&
-��`;�	��7�ȦF�ߢ
�䁸A��;ә@��>*��;�/���%!=Fz�K��}P�)w)���C��-�h	��=*����IuǱ)��0�+fK�O��@~�;XlxVHYEB     400     180�=��r��<&��S n̨���~����������k��.X�BR��w���lu�/6*:�k͆8KU�T����S9lJ�&͹��\9��#��tU���~M�s�T@���ӊ�Q/Y�<P"Vᢧʼo5J|A���QLP-�M[�Qlড়(�z�H�(�n�a�p+���ض��hg"��ur��d�ɜI�! {���x�K��u���gl�# ���P�fX��mR����݃ۆ��Q���������؞�-fΠBX�P��p���,����,q� ��`��:!#p��'|��!�N���C�'J��=_Kpw)r��AJ�҄:1�}@���L��M�xh���i��x2iY��?�A��С��Oͪ�XlxVHYEB     400     150��'w�-�����-��r�������.RҼ�{�^*�f70��Z������8��	����{2�������	 ���I�d���͙E-�tg���Q=���U�.吚�(n��1�b	��M���p����Ҍ�Ja�;�'���ܐ���K�%w����L&��x� �c��+8�1~|��W�!������}��~���0;�������xC^�/;���t�i��A�KO�n�7q�h:��)�jF\c{�a]��n�껺I0c�JB��c�v�{c�+B�7������N���н����FSN�� �"�ς9��L�I����j�0�XlxVHYEB     400     170��d���8<�bԥ�-��{{G��`I5��Hv��8�H�=�X��/�}Ʉ�B|��ƽb�ƾ$S/�n��̒)VE����<U:�̨��<�i�����p��N����ks��_ eI�Ӥ�5�p��B��"ڢ�����$�vKyQ�l>���ݙ�wt���nND��B!�C��X�WiҗH:�f�؂�&��恘_rAڿ��o�C��<�SIO�w+���=q�ԛ6��v�	��G�e�-��T?�\6���
ɰ�ON��㍡�R
�����p��h�� �Ĺ\���J���V�t���hlϾx��JE�9�+���ᣨ�~';g�$-H���SJ-��E~ցҏ����=��	�gXlxVHYEB     400     1b0B�8r��G��rw�Cԙ����T�e{��ϸ!���ŧsq8�m�\��;)����^���i��T7'�w|-0#�ί��֌>�OUojHqNۙ9y�G�v���q��k�0Y�P>��tԲv�Tš�I�G�3hN�ÀT�3�'�g��Ӟ��Q�z�V(��c����aO4#���q֛�ِS�#��4_��s^Ф�r���Y�|�q�����ft�m7��l/Vf&�d-Ҥ�jǌ�m{��2�h���J~��Om��K��:��h3�~X�t
�
O`
 �!�%V�������
�����V8�t2V3��V��sqQ�@�˺T<�T�XB�a"V�9��S�K����eb��E�~ʕyO�>�,�2�f��G�}��Pn|�G����C���q�Bu���k�p�&��`��XlxVHYEB      e0      a0M�S^��Y�22�<�X+��հ#!ׄ���w�&9��~�	������m��Ʃ�]U�O�R!�dnslc'��>A7v�����~�t=�U�*^S&fȍv��`�b_�GW�,_h�[lZ��u̏C� ��E��b�"I�,EtT�_M��u�i��
�ZJ���