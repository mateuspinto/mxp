XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a	�Tz�V*�~L7 �����S����ǅ��1Q3B��c��	����Y�9�wV�+��w�# 5	����	!���i>%_ޯ�Y��H����%m�U�l���T}�saf�[|�̕j�쌿���I�O�C"f���♻C!��>U�_�� WQ���4l�)�a�	b��t���s3�-ڪ�9�:�4|"<E1�6f��"w:6�!)h��Hx��Sп�}��cT�0'�4n&,.��Kwþ�����X/d���&�.W9�ݡ�Q�0�޲/�ɰ�i`\�j%���x�W�k��\�ښV���fTm��}��W�M�!=3��8���K	���o�w�M��|ݙ��N�.�����Z��|����ي���y��qP�'߄���5w`8�[ҕ|ڷ� ���s�^����x��߱�A�-s�&l0m�s��į@�T�%K�����e�?��{1;~�,=�������r�e~E-��w�.��ENe�^� C��@�����X�,� �]�]���#����}"t����7�z�DS���>{���gW����s�>���ܱ5�NڪF_p?����x����؞�4�`�%�>�MWP��%Y�<�xF��:�c��@V�������5�:p�|Y�[��"�dɗ��vՏ��-�[,�B�G!f�K}R�םJr�U~����,��"���3�f���J����<�>r,���A
�>|F���$�N?W<fA������0v9`p2XlxVHYEB     400     1e05b'�k�ʪ���^5��t�n����=X������6��]Q�j,��,�v[C�(��|�n�hC�U�,�H�~��&Q���q��!- 8���Z�}|&L���m��S�_�Q]�+ɨ����7��0���N��	�R�����buUy�,��lb��:����)'��,�U�B���?�X��)�Rg�G�9y����:�����v{V5�y<��[F[�s ������O�y��2�����N�r������B�?�����hD�O!�Y���v����!��pO҇�P,�DpB�'�ؔi~�B![�JƝ��a�@E�����T� D`�V� +�4��[DHZVCBiAcz�I�^�G�����8 �t��{8�i�]�aA縭��vK�&����c�!9��U�E�?�d�U�H��1�cr�cu�οX��g��H����Ji���B;un:�F�(l�&���,�V�A]g@��7�7*���)�XlxVHYEB     400     1a0�M�XH�e&_"�~���T<=d�L���9ϻ��4�f��œ�0z����9y�,�-�_��W
��#�W�3�Zb���Z
�ϓ�EvW?Q8[a��4�����)�%^V�(૔�Z���v-����K�w�C}:�U^}9��t�dW��ʅ�t"�«�.�@�Lm�zS,ў����o�Й�]�9ɣ1����y�ۓM���,��� 1�#�cZ�޲�z_��c�EՄ�כ��"������ѓ��=Z\��ͬ��}�m�=�hq��� ;��,-Wk���?�a���y&Z�#5.U� *ాi��O�7B����Dp �'��9q�,Gw?��晵�i� �AP���t�|m�a���ژD�����k������uY�3�"�b�J4i[��F�6p��G�XlxVHYEB     400     130KB;I/�-�Z��#�.ߩW��,ș;>}ȁ�B_��� ��<9Y�x#��X�l66&���\�6�e�`k.0���k1�ITS��O��@��iNg�h��Ǚ����/-�Hh�9a���#%'t� �f�ҥ��8�v�tZKTe �����W�>��a3�Ļ5|?&��\��ٯ"}��C��3�u� b���-�￺�k��[��+��^�T�r��RbEMu)7��.��q�+qD�:��6@��P�j�@m�(w��8�X\Rv�\-V��@��P�I��@sV�<�ث1R%�WQ�{XlxVHYEB     400     150n@w���@���灰Sk��y4��;�Lk�;G��ށ#�[��({sB���Z*�x��h{b�l��*:� ������.T�F���	lf���(<~:X�I�\,1Ԗ�$pn�@,B��q�c|B��p�jT�M#G#����UI67�������	:8^!��ļ2^�~���V��`B�>襕q�����#!:�\�F�ԋO�Қ�A��	�K��^��f��c/�P��,R��,��ɭ�h�c�=�1�
e�v�h��gc���)���P��F�{_$T-�5�~b;xP�yR��ͷI�)���o�d�1)��9���u0���29k#�t�$*��'XlxVHYEB     400     1a0΃�OV��@̷�|6)�/9�gܧS'sk6!t�U%J]$�idsM~/_��,@p���ٕh�ፏtU��Ȃ�Η���Z��i'w۰}���j�?hI�s��*��{�J���T�����U#Ne ����_��!����9���V=��R���!7��L�-d;�׸5�źd�a���"
ѕ��[����G������	��p�fs� ��v�ɂ���>p�����+�YR��-���� �g����0l�h�]�$I"u��˩��޻\B�13g�Y��m��3��6������Ϡ�¢��k�b�����Ƕ��;�I��[bc�"r�� �!���cb����7hD�5KD�:4�d&��q�޼[�j4��@�����D��y��d�����cCh�!�l	6�XlxVHYEB     400     180|��G�_P4�گKV�<!��0R�
}l��XT����y�=���`�=FTT�1t�j�=ҍB�=q�~����N�����n�N��RTE�
��Q	��l��GB(a}K�������l}x�(�B#�W9/tO��`��g@��&̕��Rq�V?F1s�ʮ�h�|� �U�<Vt�	0��#۳��/���䊯k28��n��:t�K>��Ԙ1Bj��kU�.��\�8����ͺ���<��b;G��������۽n���Y}�@��j~��Ԓ*�bdI̯�p,�z���un�"W���y>�`G�F�c	�&r����6��";f��׀����j��Bu�vp*hD� �@lr��-�J���~�8�<t�(w��=XlxVHYEB     3a0     170L"_���Ě] �� :>���w�L����Oٍt��fhBI��_�`_�,?݌�2�<{4��z+��r#d�c�8�z��,��V~����dx�X )+EL��ښd!]B�Q��*��·�-�o�n����#G�/�����>��#�)���@Wnd.��'�Kf���k��^lW��fÏ�Gl���/��f��#�h�'w	s�Y�%`[��؄L5$Tv�& }3�{?�%R����,}N�_����].�BC� ��Վ���>f:�x<��R��=�z�@#��vӥ�t����e����@Q�t�m�`v���:(���H�|��`�V-jx�a���Q�a�~���r!��q�QF���ΦG����