`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
0USWSUGxovGsyBJteYpEoZULTXO8M/lkrR88gj5kiv9KC/+dcuPtgbWnOJ9KJj/5yKBPDyWYIVbJ
5D9Z5PBYxQh/aXUUDQurUeMWpsvkMQAeH76yM5lLyZyi4JQCDNFakFpePXvtzw5+g0oHccB2lSPq
UoA+fAQ9cufYXTZjW3M+2/xt8lfLQyRC5GaFcfN67bUDGd2/FpPBvWmZHxjUnyTUp0HhYqTRn8aS
Y9TFfMh2Y/Rvb1jh3Dg5ah9+axL4M0HVzI7T5NHvXzPgKbT5Hsxxavh44tmUzOEJi0j4CXG3BgZL
IlhEZTtWxACzyIGT0kz/cVYafCr7F/0ZdIQAK97GVoZRz30mymjnfSbys6IyAPemFeishjozthoU
ItbUb7C5rafxcB2waTLV47N/ZzVZHl60Q7S+Pqkl2eJC0oDxM6D+PbWzM8dv2HOyLJtPddkKwLDG
MIhdmkw9Rd0SxzKCuCSbweeUscx76HuKCnmcJlrU/r4LYynnUXE5Fw79pBNOJ9l3qKVBa1Sd1oDQ
TRj9ebUMiz3jGDpMXsJWXgcJYPcuObsOiTVD6VRvLe5cMo6q/Hz43BKUe2JwuAv+KTSxlpR+U8dX
DW+aT2l4BBorZYgHn53MQsQ2/7aTqcxSf/nuCGcXdW3hm6FQzZQYZns3w0ZF9Af2L8/OB/o0eapE
3ODUTz3Ct5Xoqq3Ng++LjbIMwPGk8xH8M7bM+xTQgT6deL3srcAseuCjKWCmqy3J9N4XNxLJpsM1
k6AlOrhrajoWT4Fc1MnLO3NXcikiP0pb8j2RWE6iqz7c7qN++gIvmgCP4zIjGtOfrYWO7YBVwyiY
XP3dMTgYtKAdo2h3+sqo/rxU49dzL6i+E93NYlO65nQlgXPnVjT0gdeiTrTavUp0UVFC+AE5GlY0
XuUIM6B/UvD9YvvQUt49sN2MfFSjaGGCOS5bg3NCykBWpk74yHfjM0MfWFQnQW9W6LKinb7Gy0Ol
73CUlQzSNyL1XsdWlT9vunaMNUpwzLdozkLGcKynOaENrlOZ0rWmBLGhx+K30Io25GwigMWv+FnL
nmyiMCbsQs5G3tqAkVx8LzMna0XMePs7Ui/DiL1L08HRLHWvRcJZPIz0aEVTcsO3X/C+A7qBscLS
hJuX3mRnnfvzcuTVkRaWHMbuAygyi4SWKTvLt0gKzpA7B6OmR6cEBOnksdg/ERYS8N5BFYWCk0pv
PqDV3NhK7PNQVzR2p8uHRHmALbgItqmnvIk92ceKqKi2r7wc1jsOdi4VEWwVBfhvH9jL29xIBlmz
CedWs8JhFYJM6Ejx11iii2biU8y3KnwoexrgeNuYV9XrBwCnRz2yPjtiEh6LfolxBclIEhtAHly0
tNX5ruaKm+RWfp4E5po698VTQkUe73altDOvL95UkWtH2IuTArmYCMFFt9tT5osZc8eP8VrxLHOQ
cCiN9SIaz/7+SbbrsOmL3hQi6DzdLsCUdNIO4rZz9pKCBiVoiseXidKLi3NUyaG78WLJukNrv/Cj
eAhTH1gQ9f2O65bKnqWWecxRfPAzLr1c5c4G2F++KWWAbiMfbaU0qkGJtfvXy9RrFUT5tn2x3QTR
895RC9mWuX/b4lAdf2kBmaRpahtnurdstl1K6yDdEwZiYhxd4Ke7qiAtnxyJ1b78f6tgR2wLcg4v
VGrs3WlbltZqD92UC69jzhI8K8+IIz9sEshPt4tE4oK7X10uEyJ9CuHSnM6x9C9AMVIvbihucPqb
aP4zgwEJMfdKR0OulYJTLfHNwxJgk+Dv8WgpimftLySeNH0GIRRYcQ7pFsEBZ+cyWtOwvaTVFGWf
loWsuUAp4Omi8dth8GxB7DOpoNc2+WFLZQBud/PgcRqKNtQ+oyUB0nLRe2nS3q4fGoi5wDJlk1qL
8YXSbBXSFmGCAgt17Jzt5lijtr1xuiVCLM/mZlUMl+kDJqc9iSQzomlKgK8svVPPlA/nM0XiwwGa
/CB2xCpGypItDuMHj2I2JQtnOhynmyUfPGdVFpHiNdAVvsRrLNCSOU94A8h3mhnfJ95j2fFoYxAU
GlMNcIvLsAJtSfbj/d1d457g9nw6t41zUpgyZh/boj1L5Rn8Tv0fZe4MvmGOSBRiWspt5MiYnONE
ASMsY5V/9chLAoAw/lxqjGIl30TyKkg03TpRGke97db1W9lgbvywQgRc5HZo2ESVbD7w9grLweOa
MPS1QK6tqi8C8TxUUDVgq/uR1Qc2lKQ+3rt2482FUFhhgxjEYWfkGwbiQul9VFpH8XgBymuhJ8cj
2kdL7yPKswhww/G8dPf6X+7YIUjcdg8xcFckz4DR4T/BUewyAZ+vTc5TrHpeJcnlh6O5jcCT5E+S
WsV1A6RoF1ZIpl9OYPr5oUK4D8XTLnVJkKliLmKtUL0NfOGSUNG0x8JCK/f9Dq0u+9ycGsexhVON
qy8khUA/APtLQJDwnYUV/tYSH+t1Qy4c0oJ8IbEkoFvH1X6OtMIJiPjc/sS3uUsC4FWzuUfPKT+Z
FsXJDnI5bWbdtxJgJKKayt7WYTQ3JQx4qTRf+BYeRpOuPYa7m0SNO5rkZyD1uHBbB8TAqXWIn+00
3+7+Aq082P/GImDudyiBSqn4eDrrdRa+RO/ynjI8hKIbvAV6UzailXW40p7sZB62V9GhjMWzS1ov
6eFNeOa60areSNAeFPUZfC/VSHi1R9FVBt5JYLFW6Dyuev7sH1M0H7uYu461bZiLtLXzAonL7bXM
p19NArA1lkwTD0IT8qi/H/M7MByPqaz2cLrE+vheCvlWEITBtWUo8sOjVI+kXBz79PeoNxCFBwM1
kpytPMPS6B4M+azWWgDOmS/KhdJDuJQkv9kJe2XAFUe1+ntwCRevIvHP98xQi3//Eg1xJAbaWjzD
5jojiqlq+reqccWnd+SlsuBFcdRKlzCSUpbAqFXH8ZrHo47gWzZpgVbuBx5erju1N7At/huIEkjD
d9+L7IKgcL9w9iFpx/GCwmIqHHG1ZjXBh+M09Q/Zzi+g8w1pWEGtD6rpGX/uMZf+0K3d2oLp5YNN
/6rved0lERPKNFtXXmSZIgaY5rASsTAHu6dYE8BI5ID3GmH/8/afiIqSFdU6aeQDSc1zQOq0Wb6V
2DqCCiZ/bKulY7wn39Vm5z1DZqtO489WeGnFaqc0EAuReRX4GIOKac8AQaLVWRPi8GxRzapDeUbe
rk0vTDq5sSqhmza0s/BR9icabtumN8L4Yz5PLFyOOzLTmoJQjN5nU+1tTCLFLfDAU06tDv9TI/Bb
Lkl62kjCPsHSxFPVUQYKsfNlSyZ6Zeln8T7dTaD/1EXhclW8PoqzswdzlPiby/xwy/4DTa+7Q055
v/KJqKQreuTYDkkKWLLzOd6/lPf2rpl1a8zf7mPvuHUUiqd42DJjBB4Qh/kpgLaoZuhvQQeLNrZN
5WVSrvnd8x6avWyRXsKP9dxgq3Cy0FsCdwDG+tSUOCORniDZN2dfRjfq18oU2cnGLsUznhzKka+4
lQ0+1MS5V6NfoSW1qnD3Av4IbllXh8rECS2pWW2rvt4TSRZxYgCqpzVhCCrQhMfmKuABv8r99fod
iJ5C/2FrpCe/o/JyTd09oEA6iBNL/9gWkhy7UDAzcMYbEt2DH/I5D0FxzTGTC2Oskfjv3KTd4PHS
gwY5YYbEUWqJKugPhykjPS0xUFZXUN/NLIgu+aazmXaPyDf4fhS0TZUePJvcIgHcUdGiDmPY7zNz
ih9pevKiiy9/MACqHhR+4kFJ8Ior2Evv16xXA+zGQd9AtUPS0lry51zfkGNu9c1NQUsJsazTQbIv
ditTp29HKHljFZYO68OqTLq2ruxeswgsN9Tlg2YnVq6zFpvxYn0JyxTiu4LP2pVzfnZ0pVGUZoBg
d+HGafYHE4hLQfwczfCZ48j1Kb8ZXfrZSaCX9vF5R8HgWkUhTrrY0tLBcMhp09KUmtMdtFPtHydc
yWIkMa9GoQ5bzumwpFIhpeyPNzfsoniu52gs+9dX0cU//HYbyshXBaAL6fpiXBj7k1Yxi+jEneZx
HD8LEl3V22IHC1i+kIdAoaFpLZACYF9yzsLk308KJoUVPxH86fV5iet36cOqHDEFcjCZgJsEgPJt
Fb0Ydp2L1fQJuTiPncNyFk9FRwingOPRmjzmvip+yu7UglpLZgDVLSHLLOvq2lPPrE34aid+4NlS
meuNU3nz0JZEXsNXCVd8K4iGCRvLvP2vPVPK26tOCIkAwvvRAT9Kh7ChqkGx1E/bjjSwOp10T+0Y
2Udpn5CZlzDQsguNYiQ9VICD0kkjTLQf1KlRHqxrnm/XKYjNMeYi8HKrsksVmPnrn3htraVtzYq5
wckAGpk+uOv3np3h2crAEJWJfRKGQkLN+DQq8wsBePA1YjQ2oxjWh0xm0CJJ+M1olylsIhh+oluK
E3QwSZAaALDAopFHhfCeMMmbyaYv1LhaYgIktcPgSWAiClP9CfZdM0MCVz5km6kMuAB+hwPXtUFz
WtdDNdxvrzYZnhgQUjZZajR9LA8UGefIs2ECTo9kZ6mvIeMP8T5YczNPBbJhw+AeAp1jqMkXwkNi
VQC8fKVQD/ufVck1tr282WlYtXnTCQVEoRP32pKruW9+a6odn0ocK/HlmgPRB4Z1RC5IlwIQ0VhX
pqLG/2HnGA5C51O+USuL3kcUNqLVxTWBEt/EvwJZadzK8EuDvm53baezBi5jS7LesK69l+LsGv4C
LQpIH4381v9mrGiIREcN0REw5QSKxaQWYsQXw4TihmFvnNKff10zlrxtrQtALFPNvRYYS9IH4Bbz
TVV0AkiCiv/UOMat8NXkDQQGk6P52xvl13Iox5kzjHbdzm6U7XUXtGbs3VhmmOFZ8aPNdbTX8nWD
ZWDtajPS19uBO5qy2KOjzHzROHlZkYAv5UxXYdW8nrPcdG1PQgrM4iz+vC14p4f5rS4KBMR4/1g4
V+28Hrw4dFGFYrCVFpttARbPAf6ol7bNxkP3pvPbyv7VmwxUmTkNqRFGTcDPnCX8A7pJ+qEx9M8d
gbbNlsJ27Z3q7089V/zmtE/Joc4QF+GNEIdr2FIVBHxrva+W/Fomlk965+IF8wjW76V4x4qKskPd
AKNqAnIITzKf/u3PGRUoCIh5hrMqNYdnJtFbKuOQ0554OFOGpxCe3iGBdn/qX3hgoynJDu+8nHaR
3D43DDBmn5PhK7xBN1uGkxSk9vFS2qMKerlB0CsqBmF/2FIPpAnTyu0+1RGRnbEng0FNfZArg5/h
jBmXjcR8o5q5aiB8uGU7IfMd1oxrw/LZngcuVZOzzMcvfY5ouiIYcFRQDpIk8grdLtvpYBbUy1Qx
u1q//0GdTtVrdFDvcUR/kZtvmOMIHXjmUlWeAtq3TEqd9xx8hBDc+v5MqtuF/vMqlhUZDU4Uo9FF
ySuHVXah/20jkyxKW86p5af+iJTccz1M/NtSU3+TsKb3BlL3/luPMGdUJFV80X5YKt7EeJSHlqCi
qVmEmWFNFkaWSQjG9OOMqjZc/fyBA8kGxezklrfBBJUbNjsbCLTzPzBnxtZgJMO5EdkKY4wK33uC
9RC864qXtPVLwEPswpaI+NNn+wBQHoUNT0uGV76/ec4m6b04QbuuBkcCXBle9VsjkSsm4my4Hf1z
ssaO15sPQHM4CNgPiSESgbV+y0BDxFV8zF9gFRP9zpymqD2pN9EskD/lf4qERZRWSnCUs840iMAs
WSGFyGSBzEx9+tTv1TIJR7/2f7c3N29KXjHw9ezO0CyDLlQjqt79C1EFmTHN2gKk/khQn0y3dbGO
w+QwcQGbEDMVFrToxHe5fGyIigr6x08JYWeNv2DNsMeAAkA2tcIPM3c9qg5s+xLrrwJSFR4djyXn
rYmUh2JGzH9OkipeQJjvOF62Gpy/Dj1jXIK39wWAHG+RMinuAo+bKumr9tXJGNWNhoB1zo8nnrB6
d6yCnzPfF5O2h41du1UfO2Yx1eXI074x1m4spUvpUPvdDMv/Qz/VCthoeCaoNpOC9KtBYx8GCj6d
6ubBubjuORVUcfnBuvORvGGka7RAYJzCOvmo6g1zQK9O5/aR4SB0AR9HLDHRD36LbFyfqW3rKWjp
+MeQNM9SaGFJZUzjYflkBVRb/CzQhsrETpegPuVD9jc7V3X8t6q9fQLcm1PYblsNwf2QZhMsAdCf
v+n3dS2QQ9Dkp91jXU2jVwWQHUfF9D+VPYTbclzSET1FGp4qe59X5B06pcITI7o+OXHZoXAtidlK
/q0wHKMJVrQnRNkdzEVYQcgMWUs53MWjx6jZe3/UFA9LDasqcEnEhGtQk0ZkIxQiWzcyZXL6+8Cf
XMhEEton0EmilpN4/MURQYARWBTPe67f/pI91j3Sr1zYTnM+3hqWysZxKRwy19m6fhGQBpnqMLh+
/GdVmY2ndL5N8sUfFYszHPbhfm+6HLkciwQP3XWjSJWPsFdC6/0Z1iAhVFR/bsLtYGLO1rs9roOt
OJ0ddHSbs2xQWaroiuF+yQMgeccE2pHErh1sxSKqn9lJIDuAU7gTtnHF3LWgIgD7GRhs++UjReti
Ru9S/0101PrEM7dQCc0jXYCcP/wbszhL7ZGLCcLIV8ukQCoQGds0EsKzgn7l/asUhW+fg7AmcI/b
1eIPjErKBEc+fHh6YTj5FHOP0vYwRWZtuDqBim3iCEq1yg1H8onhRPHq+xhetHPx5ED0DbwGj3cx
PIOU9qGrskrhcR1Ju/HkLYARJ1Qm0MSPCpe4rhHQFPISnENIhw4zPzPAYrwZ2DQl/iEFNav+myK8
KSAUn++QpHejs2zVmy3eY+hLzb1AR0QNTt3ARn+5QWzlG6jyqKwMopGgXo0k0RD4IJyM2VhLS5vx
ZXcll20mEdDTf66MFuFi4qq11pI2z8MMLer6bblIVSj/nNY6dKMNXUUUt0lb9LCgdXkPRvJtjvQ9
iLYaOXPdWIW8+Mng0linr6HXKGLQH3W9hgJaSw7x9LupBGQWq2KQ5KmVj79i5MSJMcXpfkiA+KkS
UXjJsBgbbD1QluDnwiRIURYLL6u0jGUc/rdpWdHiXC8uWFeUB6WAT2IkhKe+VfqJFbsU1QV9siup
KT1xRr95SnOvu5prE+NtAyEkAC911jjesZXB/xtB3YL52W9CpVeSkOnEf65eUjcDSeAd+5r9PLSZ
KGCGLkv8nHBFWOLmOOJV2n0dwB7Di/zBCIH4QvAjMF31A0ySvoLIrRfy3flOzg+W0y6c8a3BIo2i
EASRkHmwiYaCIiS2wtteXZFsWHvep3wIPX1HTpfBadnqTOQOCeP3zR+zHHp9VsfsXt9idUOaext1
xkvpSwJHl27i/IdkMDh9yKQ3cUGLurjmVcHpIi8XdKT2OINOiC5D0U66ItDkzbKAWhixMDCJs/Xd
OcTT7lprw5ZkL6HFHA7I6aw6JCVspUVkh8nO5SjbgHDa10rwM2b0p9P4shVs3O45/fnO0tXJXN+C
zAlj51L5ERDFlwGEhmXQbpGrnaMps+iEOQ8X0amgIaN5+or9K53Dw9A0BQAnvg9NL1OnFODj0v1o
4acv7k45sX0QM6Jie/KMQUtJSnv7uDJLXysmBgVwKJvQGX+rbn5xMrYKrZ8tnT6cdPRkervod1U+
7f2OqBNeutR7Qbw12BPD5Zaw6Mm08joR0u3AXXRb5IwJ40t6UweGDA9TApnRc2ymxhhDXs05Y/3n
Aq70x2TvyK43chDio//38TEIYiriWJdUN5hAG2W27jEdBH5XN5QTlmA6ochgLxRQzFZz6ORcTBV+
FWzjdhbzYxsONXuesmvHVcLig2drduFfUOgL16FO5wwJuBV7XsYRnXJeC+qS9ZnkajgJGaJxWj0z
UlZa/SjE/bRTmvFxEuNylRbMw8/XpuRToMngoQQ8s66IK3zJpzx3QZ8rNOe8tYKHFSj9DC8iEJXy
Klp09P+z1Phki1Jrga9XvaoFxrn/+9GPSCc28bQP8PZIEPz6v3BOWnx3Fa4nSTgrIXoG+A8ZWiKL
i5zW1B/qUiamaIrz8rY5Hf2hRIZLw3N11QJooOulfokh6m1uQkC49FD9RyGVBn8BXxvl+DzPIR4I
94PKsDDBWOZYL9rgN5Ca36eS+eEM73g4tLfhiSlNroeRnKmFIxC7qb5VRVw+2YwazOJJKDc3kgci
Wygxq/ah2U3d4migYxEi/ndcfXEVknX9tF88oqz0FcPP/y7RzX6Y5+nTYz1r1q2MI5zeJYNzx78Y
arZIRKfb/EzN1I3A4x1mFB3Y8LqIC7cMJzGcpR5ie5eTGOteA2ppP+aLtAbU69GXoZ3+C+zILcgM
a/X/FLlmIwr8tH05JfsbCV40nfrs9C4gZvA1rW2a0Lwb4i9u5TkIhCdJzqc56GdW4SVA1ZawUS1N
No8oyElC/0RGyaS9B80G2fhCd9h4++Gp9YE6+StjTZZg/hYJ9ZC38unKBI7OctmjWUr9w4S5n4Cx
p48E9qynnmF6g6wJ7VTizCOimXzTEAT2fNToeoDdqZZo7raiDXFdKaGFahXARDyxNYxAU7T+X2xp
vVV1IBlQ1T4qRLmmnsA/KA==
`protect end_protected
