`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rnt+eICI11hLErHUxbUgrMs+hbWtpD/NgPopFxIfX9RuFjsPFjGLZBe4TbAYaytKrQj4ZRLXw8zy
F0mbeotM4HqNyMMGljRgfcZCnwZv1rO9Q/bgwCvK/F6y38+8PzxX1ZS4hPT8eI++mtwzfS9RMefp
JBZmJI9+sPLSP/W0iZJMYBZR9AjNVMWtHHwzydEW4ekpnWIeYG2fXo2p0OyRL+o4EzIIMU2FW0n+
c2StEKgLE3WxIPpOELYhmkjFPy75k4A+gEsSgYWwUouQ2KwQal6j3nq376eJAioxOa/MHZ2H8dJm
oSI8ZOoEO9gOKZESITz8uqkulRpFN2Pbt84XhQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="X8pQRTlgSCDDetM/R1pvctl6Xyz0OdaUFRtDknsxg8Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18384)
`protect data_block
k+BzAlYHzs60a5jYBFf8oSkpcUtjJFqSG9yY9mRA4KafYW4Z6JBIFFx3DvPlWk8/1NtiZgscgxhv
Fw9v7Vx0BhHAQLKBjR7+wEYbndU7RHY+7raoJf9m5tJclCwP1RvI7fUtSwYTsmnBfsh9+l2P+Siu
TcwOovve8ZdLq8zFenV+6KedEIoRTvmZh2cWxpOA7PR1r0aWkIYVjQq1D4BHiq0H0REaKDlgpx4e
g9DovtIdqt85PaY4M4a7ABeCRLo+/zHdKSGG+1uHH84AJ3OBe7HTx6bazFj8DTwrojzOMNOLxsyR
6u88yQYgzhJH0ZhT4dWIUI3qVCpTvbALxs1RHyRMpUxN+OWHa9PLolQYwY8FyFU3l2o7lUsMnBUf
SdYMm+MLBkVkcdiE59duTCNDBGGSO0BJ8L0bIk5HSy87ZUMjE4UWyUw0i9DqChRrMvN4vH23iYAy
4B7syHpPGZiR6jZ0u7D63xdxrRXyjeDXsF4HuTGVeNcK1jMAzAE6P5nJzQ23jpbwxrNiti0f6Nb5
q0DVN2ONfKqFYU5Qyi/JEHN3gY4tXE//cq6mCye++NjwkHpYM1R47K4Q7KbUkARSyvO2kJx+QnCd
5qhk87j5PLJl5yd70g9OjHxeamkQ3jXVFwj+6VQo//T4wEikcv7fbI+ztPe4sdJRF2LI5/noAW/g
B0Z+Esej2JXRN4WnE8PhVrmtt8eeB1+pi6KB0nvSM/7pPdHs+tj3shgezn4egLhXENtYZooUya25
M0GZsvP1EXBgrxUdR3VUZkgFyAAPC7xjNUbU7x9qz0vvqvKR9hO8rjuMIqaRfVn5/OLXst7mYnlJ
prX0zp3270VPNZb1vrR2X0JN0jyu1teJzL14GhPD5PO+DPXVsXzXq8kCnIfuEiO0cJhXNcqx2iHk
LM69zxtMnJEJl94ggVQCGWbjtex/ccDuEZM4W0ln0ZcgGG5PiapGUqXujrONzQ3IWRiLqQSka0NX
jflvoIJko05o3kkpoOQ5yu7wW6WBw+GL0oUGkQQKao1lWE6lxoSY++U1jcHcEdAOdlgd+k1nmivf
fGnzpr1x0p6GiaYbEv020p6U8udrAYXhXcGV9jsnKvm+HfMvawAm+uis9u0l7or7Xb99L2ckHYlQ
veEuoicSHOTOPoMnae7Q195CCVi1iLnQkD4i7cap/Is/HObNpHl21lm8+oWv+3SftTI4YKfrRCi4
Jjm4UUFgiP4c0AbBj1uKTZkr7C64IJ0DrskY7SH7VI7wS8gl4v9XlKe2hUkl+sgb1Y2QSUGR5K2g
gn7tcLCyI7ClqXWKd4APwcEOl/IbI8ofJ8mQZrUWQIUu3PCf3q9qLOdGCiUY2dXxpsIF0TgwsDvC
LvDpbu85g+Tsz0Gxsqo0lbS7YEHaBvzahlqPvbr6UGtTnL56fQOrlRckhi3H4lvduloq3XouNTY3
7sEUlloKj5mDxy6kW2q+nJu570Wa/1OgL4DotkEduhAcmc9Sd+eDEDDiSQ4F3lHjNNg66YUUxtDw
/0A62aStrIImg8eddZITNdSXOmAtEa+zYGkhEIejjFWdvgPsAPsCjfcfQj4MXF1f42fcGhUjPqb+
N6OeCA6giQRSyAorH1xNoqHvVS4/INExVWPU/+g/hWT1yUIdVY9SuygrcmnpC/d0bHDVZoeaK0ka
wp7JxYJGCdOEjzw7aWgFR8Pn+KIDicZncM0R8vWMs/ifAZEHcbSEwPgzOS1ce7NmZzuFHJPRuHIZ
krWyowlcGSYTq2/uWyVFycQ+i8bxb1i2ZfTO+IkMr5ccnZ4oxL/b6C/XiYWWhvxzvFMHJO7Utfmy
a/UotGNou+VEL8JsDamTQNCraJLBa41olI6BeZeUnjdkssBMyyG5ddYsoMpWooVGGLpc2lx3KiNX
YvHyZBR3cMYETRWwXsTI4tpJdH8v/Ye4HbgOZNWZUQaVnf2pMDLlDFOKZVJB5kDA5hVAayEtIpBb
8Ngw+NFToBVR6uudeNMQJNj3crA6tzJeDGIynDEAGFoLtxdp0/ih3rU5bNUfF4nehvfIDCp1KhVL
9H/qOT24FDVQAVRqtBw41IOFJx/XdSUwnMbxCLQwzFRsWrIaFN70b5MxwuNXcKbNNxTvMUu8dVfM
rGktGeD0//SrAfU73YhX0YgxSO87p2qG+Au/REyKlvoMICJVdreRTez7ZHA65KL+RxY2wB9sUCTG
TmXAERobiVXcrKNrLnohkJm2IsAANU/LlYbg7FXW53fuZnWju48Fk50/52IKb/iAlDfKU3j4FuOh
9imhs1DpydAAqxQvcF14GD6dq/PuJ/o4e8l+0ULe4JOh0BpCWtxryY/lJSyTDzFc4vOHzHuTLC3l
X+VTHR1RDfF1QnOHhNm1qsKaOHG0cwgJRuZ9sTXzrY5CcrFjK1Sfjs0ge3eKKahR8yGfKCR756sg
uZv+rmf3xnJ7AogE50TReKrBE6K8ZhKKTwxxuemzwpgNDgxVyiuj+5qnWsInaTDEMoaO6HwKLTSs
PBzCiyIt7HTf0rPL9xwUPUMUkgkyiTdj5F8PpiB4nmNA8gYQjCxWyKnOKl+jvLYzEAJ53aJcmrIX
N/R76xHH4H2IKG9aX9p092R7LYG7A5TE3E/f3JW9rqfQyBvhGIALhKR2VmpWNLDwZugfR9arbes0
0f88Zmrzv3U/6IuxOhah/k4XSacA9jtBwOj5J0BRzDTWdSZpeGoWeRLQ7xpc3yVFL5DvIGB5XLa8
5akxz/kySe7XB1k38643xdLO9ZXTpR/r71qOPoLLyzKva4UNfv7Hiw8oSKQ6Jk+7oktgJaA6b0wt
el7RrwwnMRI4snKKryEF5Sff0/ZOBQH8Sy1n5w0dtPPVjxjC0ue4peVKC64XV5ehC2RG55Ylt+SR
UbW7VNte0Gpssl6ZNUS+hOFvxLdthN5qzaz6bK07oQnpc+BYTLInsA72m4MD2OTLTb6KMDmSPZj5
h6V6M6CpX4SbfPmwDFIX+wfXFwQ9cPQARv4RFLXPWfyGMXVMFfvMjiL2YevfSqlr4AjRwNmTIVXR
OjvS84MeXcR6S257Nygw56TMG9+KZvS82daW2Q20PltJKw3WunLGfHEqApFV3X3p2uthZczhhLgo
wU9WyJ6j/Gt2kbhbqOMm+Ipa9STP40iYuU17ITXt8T8J5OO4cumpvQpvqE3pUIwyUzdOvDBD3cRJ
wWzMQmjwxArAY0bjPG7p/sDzobrlcoSTkPiSFTV6gGXFBbUPsmbh486fuci9HyMdE93JOH37y9xI
xbXdIkwqlGCruzC5vEr8/ETDk3Ppod913D3TMZIM/lrnyzmSj18Tx/8X8XqeoqNnU7w2g62BQOuE
5pG36ANqn6eemBc6lsnybE8Q58dNytElZJz/v59nxATSPfEsQS+/fexzpMBzgyAjsdABpAxsiJaS
obN1o1AncStXdGegjrhgPe4+tOHbYddSut9O5HwCl0AmdcN5p8OIBJCVJMxJYOyfhaInDN5xntHN
Uyq7P/JXbALDE6jYR+m8O8kTlwkHOxVkt/WVc0SblwnZptOdR/b0LXqHMzMw1PNg0OgK04yCwffJ
WkllObE5hJa5u7GJTe9xKgsIpgiwbK4Sm5WQ2JJG8d27Z6HjdIC4H8RPIlVs/rnwPkURqudNANnr
MOxH0aa6HgLFKAQZcxstI4FudM4bHFUFVXi3ULV2w+nqMrqB9AcAgBdZBNQRmFN9kHGTFwNIT4cF
nMM/aXVzWYp4jSp/A5vdseBgMkWxx6MMcXFUmpHKV87OkaubUb7K5WetWBuSCpKioLhY49XgSWIz
P8KGhLQYNRi+yrvVVb5f75i0CHavYLJyV/aVUohVLv15GM5uHk1tM04YBnYDyGMaupeej0CqTQNN
0/uaZ1t7WJ10GyWZSZFVWoRpO+b1aPh4LGz64QUBubHo2iE+9d+y8mrAOov8LZTv0/Gk+NO3uCuz
4aDV0rh+VwecOjUElVR0dATy4extMEoEPRPCMO0HOuY3VGpr4PnvB/zX+2iP4jnm54dv5XNhOHsd
ULgGDzFyPa3/+b8mGdZ0MANk/va56Q+czqNQ7t6K6e1032SxWBtsdUf5a+SmPLhTqZb3dycpvNS5
Pvw11CDpHPMikYZd+oTfW2rfpj/VEu1FmreNttry+icCRlqUX6g/WCo0uTG4w7ioQJ0BqKXrztBn
8pjoExRGkHzuS/Irclc/88HdKrInyc2Y7tmsiGWz4EJp18LDc9uIven0a+/aZVVC1vHftSc2fzhr
3vpiYEO9VZN+yn1NHncHW3fkW6KHa8AdZ5AH0cxo3IZCPM7GI/5afcK3g97X8SS4DOROOyCkB848
p9Nta+2ndPLzpuCGN/19GEbx2EdYMjT5xolxiAn7kjr8z9gbNelLQB7jHCKgOusorUPLJlFbDd0s
8+z/UduG1wCAOGmz8CDqFzOcE03PcSH3GOcFYqx/RIgzl/0i8RIehMdbzR0ou4sZk0u4LwB0Bm2q
TaQwhtBMW9Vo7T9vcmWg7KLZVZMJ1efKdclx/HYo6R3b5gm5rAcVoDcVS3TBHFMJOsNbuPiUHnn2
tjdHBcsWZzXDWswTXiikCZCdOQavHQmIQh1R/cczMYZ63pnSrCmTUvu4lyIvm9ISwFHClNfB2UlN
ig5R2Tfvt+h+koezbMbTBohw7yuwit9zFOypDhiFb+dBUVptXHOwi28+k1IBvU3rjerExywZ/qxm
PUGeshCGZyqW1WCYIutuQxmr0y9eKVz76G+21/UHQLg+j5YvZ+tL7BRDTfUTBC2HH9FQiuHRL8Z6
B1Rm8CcRpPsOQ3qVyUVCJlN9UPhkdA5Z3W4/cPCKJX3hjgqUl/iA104FMDBG0Igz5juKhjjaJh2s
ve6UAbcf7Ee3VgdS7K40AJgIt9NlV00Pk16M6du7jW4UAEa1SX7i9l+Fy0wEQSvqxqj52BEHhESV
h716m/2ooSzSjcIWgLrsKBg7PBk9T93ohKUjML0sZxXSohVyKkPaSp8X8O1g/x949r10FgQfTLQn
DHRAtvkDtRkBVH77jL6TGD7jXaTSjBlbRvQosGaAnpX+97PSf5Zu7y8xUCmq1qutzO69ThjHY/BQ
XqJ0gXo/j4BQNJCNYuRI3am4B8ys0n9fNwPXSJdpdVeD5eFo8cccxUUFzWyMnz3W1WYMw3N3T27Q
WcVAe5Gm5JDFPqCmsSa/1ebo5bnRfS6iFnxsTBlZd/GHCWUWgysRuDUdhSPoI6UqZr7YeGCxT6oH
x7tocMApNA+ooBv5WCLCNsfkh15nmHtFVp2fdmN1Og+/Ik+wH3yzZTwl657A1Z4P7Lc+9fISXJf7
wV7Am96UWbwy84fp9beK4DqgfkFCQSI+wgvQHks+7pfqIbaCZPGXAYDs7sSTzE/EoIo94LLx9k7Y
djHrYU+hsrfEWlulPJI6O/YxDmJSOsSunlaZfc0YvmdH3sr7PDWGAwFYFeEVYjVR9D1k3Z0JOYsX
hMopgbeTuVas3aj/LRvUKNmvMR95RmOXI/+VwhXZqKrpGNYh+VkmujrXRGsOr0WUnWlBwnJvrv6i
+6S4MhggpipZq55DQIn5kwE533KBaHQhk8Ak88Y9OZTHLuHWDKuBEv7LQVXIQ4IHsE2paSEvYBlo
agzyRebUqroakXovp1eToIqchXr5aq5dKZwEdtpXzL60FprkHDedcvVmRdgbVEJB+yw5A3dhOFaO
NJLD5KRDuxkojY9BWJE9+gRojl/kdyUpjuNbsMTDvwg9efJpZSZaX2YrRSD221M/cw4lnaKA4yZl
sPF9VybSl5j9PFLrlYTK5aslJZn3eIvLCzSZFpAxegP5U148+tprdjdsSXvHvmhPCpFcDV1Y4B2h
zDuvmWOa5SQ5sh6lqtceiT2aEOeLR+vWzeFfbnb/y8ks9uTrqe9drIBFBFMISt/U3W+oSSAuEiAJ
3VLnH55PpkeubaF4UWv8qUKFB21ZDo+ln8fjofeUFpTorb+ny6BnqkbTkWibH35LxOd9Kg/QahB0
RgTn1Uj1l3GvDbcfK0bYHntS/LAHYST4XJgEs/achA/WmLo01w3zSO3JNYL3PzY/2D668z3y8Y14
68F9n0NxBwcdgDdPCEgc4gOI7GH205puaGCL2x5V2DvuYDf3E6tzOxwxzGLkfzV1AI2+Cl4aOuxy
555XXTlzSDGMz7/cL4Vo2bSbuCiQvr1GWnRhp6vdvhS9pQ0E0omFUVECneJvS+QHG8xfPvBxS+yY
h2h4i1B31cYCMvGINR30FhIoJI6k6xhb5/Jq4t2oa09PoAl4UPUnsaUmcCwl6r65Crp6aBvYwse/
ZpC7h55OXepjabGOxqMY+BIU9RQbdaE24NadAbmAYOQqWxTcLoFOOPDxyYKjjAOrtvcBADI7STLa
Yz0//9aL7q+8dCRGjKRGtVprEjSjEKw4lW0sCBN0fkpZvtsH/0CM0bsxZCacPGIKu5EdAftxv4v+
MjEDy69nEs0o5MU3FlJtJFNS4M37knj5TMYlVPAE6apE0DsufdJy4dpAv05JYvtG9rsSrnX2zacz
Nb3pt+sBPLVgv7lhaRV8BM0iiE9nix9Fw2mK6ShFS0b2J5OAX1TQzaPzykkKFhTinOM/DetR/dxl
dweCijardYPXCfOljSzSKpbeNCSR/nQ2QlxpPyhirKwkI1GZ9Xn17S64ue00ywzm0s6i97RcFADc
HC8BlChmUIn9UHsLskLgt7tGo9sIr3E5E3kqxAXIV4eh/srbc7faqJ3as0ijEs+C9+JSXOKvnEiA
9E6y6QmlxEOWlMENtjyLGGB45fa3QKLp5lpBuzlPW96WAmWtHozCGAkfCWQsSltpuYLvhFQqvGRt
g6LG9mZX+65RUoe4uEObDl2RnPNWgcVbEThotP/SDMT/YN4kAHOf0fiyjp/O7pmHIz38SjXJf1UV
jcy1+fi1R/DZ3VaoLBfPr59s8pJ/L//0z/NQruOcmkEO42UltaO5ugnNX6TiDQy/32G4h7wFAXkf
5V8SBgme+Dm02G53FDvPBqpIG/gPOfXLN2d+XjNSD5q94psbmnLQjVGMp/+tt0SMMX/deIjwNSv3
WJ9dOdERtqS8B+1xdbY0TceI7Brb1W6aSs8Xo9s4JjCq5AJPDgwiQqcUXibNHlEWD3DgBrB6HhWc
URIjitcy6SX2/2EGQIMxLSvNd6PrRksSNucCc1ArJaCVxf8SbKWqrR8PiN6Heg2wYoVVp3rvidvS
xJ6iyVYZsBZyCMUM6/YvSGeIgPiM42PB+3eZb/r7abXUXIS3MDc3u1+sF3FHbUEocYmgTM6XzZOG
Ltd2a2oiHkJLkChIMuvoduO1m6U9yUEoICT9boechazinBeBH4iAkG69l6wYOLb3Zarr1V8SCwfe
EaQo074vQqMUtHbHE0ti6TJaMIY7YLQ2smMlE42zevbnz1b7nZDLUSeqyF6/im9wA9YIkSTXb9/4
f8wsr6llH/Q+9CVz4msk5hZJfQors1cJO9CeJ41RsdXHEu4OrXMUrONf5ju7w8Rz33YwthnF/OZR
nXd+6q6ToTpO6K+MbmVy4EIuBg7DtNAUfHKKwqFp5HQhjEZK/PPiM0rXFuSxNEjxD2UO8nrnYw7p
GFJf9tkdU7Hkk+WRG045JlLayDSFpxMp6q/rYauEb494BlGnox9qLw9sGn1e6QpppqsuePVBdvVB
jc6hwgYTlohsGBO/4VlB7IqgGsXQm3pNqfNinve1Kut4L+rOUISPV3sBGh+eKLCp0dggk7E81S+U
rR4cqCLyZUcXRps7Z5E4uiIZcTPUb6tSf+c6iVSxp5HGr3ppk2C/k2SMcxgHXcyA5I7mKa5NuNW7
D8ZIqj27JCO2B9GGCyT0Przuv23NMCbU5irzVe2i43plPtZk2BC15irZaR3femoxaXgqWuD1L38A
h9bbmTvRJeSKSQJVx6nfbkM/aiDCs8NQE4gRK11UtZNBzryTQ2Re8mbruW3vkiVt12Z2GobFJVUR
MV3LYsub+eNNm8qlmkphwMR4jLmFvo5vCVsWy77CM0G/6AEpFku/p6XX902TRFxkh2D/jSlZquqE
Y0F3j9MeZyuQpU9gFXnJxaCu6q3ejv4TIg7YZBAfqZXSO952IL6d/CSolIXNk74Zaf4daQkX17pF
jFdNbkBU/yeo9DYcgW391UinqaiRkev1ksN7yMn65yscokWS2JZxFWEwoG2+b3EoNmsPN+PtLpIn
ErnhVGYsJdJpV3V4TBKawIV3Wmw+gN6BhXkN132gplu+4ooyZVZoGIws7Ak14VtcXXHqLLB66zwC
OGGdg8DMl5V5jkV5ZJpRegoBsUThYqS9XEwbFN4R2jeobyN3Zb9Q4YkG4QmnODQvC4khOCo572Xw
DloxsUoP1Z7A22q1LlAITDXdi8zvzI2FcwYnGJE7cMHSIItQaAYW0Bmj8gDG9TTXuHQbPxjVtI8D
j6ZLNeHA0tgUcTze2SLHJQU6tOtohCnmdqa6ifTEgH8A6TGF8GSIjgTDETkdmAe/JdpEBQNxUhMh
bjh0Nw5x0vrTV7D/ST91uVzO5e2sbaMtkO+Jg7VnFdUL/XxeLi56Aqm0YEuxbDpsLVMXx6dFIX/0
YDIkQ3KRLz2k1qv1qDp1C7Yh7Isezx+cL8pJgoNzG5AVkWMLFhmSpiAOhiOL7yL+IdcIbpWpq9tj
/8SIuIP0PRESZ4BYtt/Pfp/wSS0g03yR0aYPVrnfgtXQ8Vd6GeZNj5rFggS5hCBgOUSRwMxIfAmW
E4iMchuyEKHo44GcBDRiDldjF02+t6BAt57OdZFEP0v7x2oM3RxXaGZfSnE1+o1gbcM1gmp8hgPM
F4D+kpROFoiZvGXD0ZWntYAiBgg9OomQH/2Chu9HEu8y5iVPgtLdvqnujLFTmRyQKIbVEXBzETK4
fcX+Tskb7LMXbZCzPdBgNXKzFij+fdlQUaZp0ReLmB6giMN8xKWkr8xptKqDJzTHiWujmYv0g6kj
5ii4/m/qJvKKsBlaRwJO7fH7Wbp0oYMGjag0zGnNfGpgFNg7HvEIswUdl2TUdoPQCzPGZJZFpjmI
FKHnVRYB5IRmcZUvcH5kvHPZKKPAnnaAjLNRFfRzBiLEnb7QLDGTG8oYzZwfX2t6CdpDSrZRAIIp
Wkub4S/Hb6u1ko/Se0+lABwM3QuPk5rogsGnpogR5xHngO55Gv+U1uILHoZq0VFkHtq5pclyvuWB
Psw8/KLXinhtqScpOozclS2hDa0WyvAwgGlBxqSwdYUkLPa7jb2q/Tq4eUvcz7ADV4KPg/eIIfsF
zVdLLkBVlzKR83UvAkdR8IZHxdDa8SKyoeAqVfYltcb+YimLiPCfajbag2fi7Bz+U1GolkbEjyl6
TEzMvKxAzlu22C90INWn6LBH8F5m3Yyoab6vbNHl560QthAnUcThAKCSlzSKVthnvATyXYkuK6lm
H0miuZ5R6rad4b3WmMO76PQWv8BSj8gOzWmRHsxpknCRSyEKdG4mm4Zw09HNw63tluVTcQyCodWm
Eohu+ikxY0BSdD9j6jHAm6JsbBcia7uCIDkf7XkW73pwSA+m3cr0JBSzYX9tJimb6UmniPU16EJj
2WnRIV0//69lrsxVL2iAA5+4GBnDaK4sgQO4QTkCOoGC4Bl8Lxsdl0E6ocLG4Rqxdh0OOSTk47aJ
a9KNUSDTYVjVLr4tqqJL/t7OuzWtL+kcA5g464NSJD31YS7P7LxCNOCGWLuF3CXwYRwrhVA/um4r
J1G3vPXjDENJzocMZLuCXfRTiHPiaeWlNzZW9c2AMNtwjEDKWyOhFgTB5osK/CPRVBRDLqYXsK+1
wh59T0JOEou7z/rsUKHOqah1F3WOR38ctsqKNKde48EImTsXJ0ZGq4x4wAkehKFJ/CBNy03G84Hc
XHk+Dl9fy3ZHUsp9ZshKpfRIIeGMh82Ujym2GmD7xL2IzKlhWLgmekE1AIxFK7zdlluVauckLwO8
BzYFznI5dBbpHLVUsEoY6cpriNZmWbm+PQL+L2tHqNBoS5FehiClIAP/UT5Qr/tlbuznj3yFPEdM
9izf2qJle9Hfie1SNFxGt7Zpbg93INmsWPEaU2dqNpriRc+Y1aUgxjVKoqZRDHcAnIc+GzUxhppU
xjjlfYVjEYDumWBn84i6vPg9v5uYDsxpYipg4vo9Mvrwp/ts2Ma3zCRB82tVm0LdifwN6k7ZI03L
VfK4YZPTMu26QbVRILX96ZQeqri0L2QGBiWdlV8JhMlPoNK1svSnDDwD3cntdZoHZ4NSP4cfiLOl
Jk7CFFpSUrsGNx62MTX80BDFUrw9LH29fZb4tLfIugN2JHbr70YhwhnKMRuGgKy/eytTjwa/CUGj
tgSS0X5shZiJs8501b7OMxlTVeMYt91a3fvJuwsNqsSjLrFlXmk35PnvbM6pRqWeTOk4DjD6THiQ
ZPOJWjfSLhxXpeBJ8p5o9+EcgMZIswz02EStv1hCpN9dM5GXF9CAez29i2tIZ2f0er+bFua7/NSS
QM/fNZOQOfBaceUc3CkFwg6nmztfmHQ+JR+tF4m9DwBJp8t0Q5yOtMRmL0JdSAE7t//k6PvWZRpm
6lcKEBjds0wIhhqzdzTkHVmpAScao9tdH1bUZqJO/dMp+I6irYS64RehyPVgqPEYNaLV95eWWQ4M
Cp9izeiJrSg+J1EWOBQsLokTCbuEOgOzlNI2TOpgV3g43mLld4h04IpX+asqGbJ0gV+5oxl+rzRC
pTF85vkMT8HVrMAzTaFwpzTu2Q0y5z7gAAAimHjSxJg2Bdiipjn41Rz2ML5zrbJEmR0E4YNEgXdb
69SzDcuE0itrwA5sptt7WS0r+ORcNwFZTPG6j2GQBki7YQQESCkNXNvfsUSvaCTr1s03dzJRQ/rz
XtqsSRId2YDWC2MBF2Bj0JehL7bXDEba+84oBBC0fpfjKinl8hcWSTLf/fm3sYbipgjWSvRi4oyh
9e2a5TJ2MeWhnjl0ThI/XJEVwUH851Qzg5p1sFYAPKchCCEaeBKKoRsCYFiaHdJ6mpTpVWTHWBHu
yxUyD+1lpKVq4aX9VPDtapzLjDsunTGwqJ/pNMg23Dr7cIkidiZxBNPd0CzB7IybqINwOrftDmiM
YQ2PRodiYiwx0WV+oJbNhMha3m2WX/qstzYxPWM+n2yc3YJh2KLJuC4zMt9BlIHz8YC+uanrK/2x
lBExXXQWKXxj/L8o/RNTekgy2QiAQZod5L05z/h6aAVxjT4ElfgQHAdyl59F9qcRSQQFkz+MlCyH
tWUWUjc4/A92ZecRmgadcz2HaBRDjaLK37zjorMExYjElAMZrwErKbpAkhguh7HOMoJ1sWqFkCdW
pwH6I5Vnl4lPRZ0UZjovRkNSO+zqXBF5O0Adqc3azs86xorCXnedvhJHPzYu1jtboprg7vf5n6n7
RNGdyCY2cKTnCgw5TKzZuIs46cWX5A1fIGMMmbg967nVZ7kcP3Bp53jLtjTL47lmYJnV10qKUCys
gr6gNGFDvWDAsns4IauqmKeM5bgdhv/FB49N8hVoxwsfwsEkhVJTxbWCHLfIljjFo1ybiUqTzj/w
gjgiIZL7+GTBWrr51Sqpa6XDrtju+RZHboB/sJLYwWZH1vatDNz7qThzvNTsS5AfXDnL3qsvkVL4
D1omuPzm4A2UWEJ/l1lEhjmT0bf8vuXVg7t2xxGqFctvSl5Em/n8yQBZtUMJ3cN8h6XoojyAAv3L
4tTVbAV+lti1qcH3gyCeCvmcEFnyf1XMAC6y4UMKKWXl+mm5s1JQCRW3jFDkvkynSUtEDihvGlTF
AxOOiAR/bya70t0gOfHxM77e67auHvB/Oy3opzAc1ufsGQDGwBqdbw9i8D6iTWkJnNalsZwJCXUk
1FKhfOm8FanUG6oo0hARnlF/G7uZeOwclC+2MNwSyguuD0hfaQwuqKF58Maj+FFKCTMy9ykOwqhh
JvNeju6EDwmi01YZoNdboyOwQ4UebHUc2Nw/Y25K1qgPDY7c+TEOxU47XL0mpxR71yn7yFuzvq3V
v7+trqCTwBoMmkbQK8Xi7mxGHc4+6W08RJ/KLLnK13RC5dYIseAwrcG1NT28qNMbLGx4HMU82sb/
dmibYf80zIejons3e+zfyFLOwJi8RGwsP7Ygxc5ei/IkusWWE6hIfWbMmE15OUQhO8P0hulVia/M
QCrm/SEXt8Ufl/qfdR+7whgioZvjiw7PtMy1ZgyBnjVCWhy9sJh6ZasZ1OEUcQPZZSU3sq6uXY1e
cNq/2lwDhBpzj/TKSILSI9iEHC/7JvstAvGmD8QqS0NSknhFTWpZNa3SXYLBWqTmk/9E/ls4b1lW
8S4+cy0jveSVXk7YMSDmBhdNO1OPamIQLvpji88zPSycbjhuuC1vnVg8jZ0I5QTSbRxWvH++LKKo
B+k0QM727M8ih15Awrlpz6MYDwf5GO6CZaI8fCxe2+ZuqK8/kXedqmso9w4QB90O3Rr+XX+iuu5s
L9v5RKZry5mNjhJoDmRgjATb8bz1QdoczY9VzJQeEuOKWtWxNNTQF3BLHyXttK8K6/n2GIBsXEgg
99OJDbgqJa9tffo9AKqJbTHfo84DZOgHxJCkzmrT9X+epTVGCMSOb5Bnlg06hFWAPnTAcHf+52I+
ASW4xA8yk6/FO+6Rp0/0FoaNOL8GeO6U+oX26rLTfI1bWS9y7e0Uh08TofEiYlUPOhSN37+BFTaa
mX7bf1olPYs+wN46slb/mP/Y/JB8J898CVVXiXxoWkKTOxaYMGSzjaPYSLWllHPzmyb4QLPtUUzk
CLv+b8OxbnGT7WIzKcty4spJDguykBjnK7amBloppFMKKrA5Qp58oEeI5b057h+iGrypnlw716PI
MhM+scYQBlm8TTm0com2bF95pP/tXvIuvPIOUvb+OupT2I0CnNae8csTBofOflFiHSMASB37WJeF
Pc7P3/ZmntNmKfcuLpaO4owDyV+UH8y158mxQMmLBnM7r/2ZpgLURuA3n6nnVZFDPJgaEDWuHC3V
i9BYxtHMOMKCBfJgHOBmQvTk2WjNehMzKiraJGyBLWK5ZAs6y3OqJNtWOAdjRpbjklLx1r0gu6HG
hvvv3e2JjNaFnCReDiGZ4HZ7kWgObf4mbQ28tFvZBzWkdY0/82kZ+b3llDzjrjL50U5+e+vn0XPI
VSOZl3rh7W12hMfRI9hE4KreO5s4Y2x6hzV9/rtYYo4GscpJFeuUyKA2raAlFD3aRs0oTdpYYieT
e2TAGUN3XgsJiLceoFU+rkNl7USwTsu5sCaI9ptddGiiKmSWdM+X+8ge6K2ahFHLGlOyvfGif6IW
AEDFTmC0ellcHz3wimiD4rUC7vk8Z/psZsFrAPqLTR1zjlWxaC9YakVRI0RCnjYx6/DATSBXnj8G
udkkk1lDyufoGTMphsFJocyjJZl7r2zIJnidpRSLcNyTWDvMkMYtk1dBHnQqbpelogAnm+zU3YWQ
nQ0/BZHJdhHlyL2c6tjVB7B2OlgYXEgNv0Lcm9812uYTjq23y7BQog77Kh2OQvQS6gMxHY0QAHh0
daKSSaCKZbamPDsQWWdgaS30hHK4IFHjjZcLc+nRkwYKV7ZJMcSL01GIh3FoBuoRJGoEZ/+J50dh
QGvi+JPXX+SU0k6ox9kgfUuZrhenK2FBeEPs2J8bPl3pX0pC9TKhQjtiWUhOgGO320LQgoqHYP9g
annmQxHpgmT1TdReX6fjzU6U14bMJv28mfNGmPrzh4ZXS8Jv+6OUhSIcCBynHjnG9+8r2ld5ubGo
ig4i+MngtDUt86Eqv8dPRM5W8NhMu6eK0CJSKqg8qs00BrgBHN/hteCFXUYwsTLk4L7suBQGyzYx
rQnqjWfQ6rJxxao1qS9r1xr/L+aKy9PjMBK+3BND6iBtYAIxLw9tGw0jC2oOnFnh9LUgXGr+uvt0
8wFUiFFdW63RobSw7RpWN3KwZAjlhOTpWB9SK6zTVfJNZjeaYOfPjS7zxJHYUQtAf1OOTZe54USC
Nfa/0oBw/0sLkr+LjWhe8fsb6nLx8bjOoQ+Lskjg5cyCXIm+/FoFWo/OndST1wsGS0wGP7lzwfS6
W7YBoyhBl9JoRBFQBTf6ARVq+5QNpiWxELQT+9bZuAEEKreKMjc7t+tQShMiE9V8HFS+YrVFAaSZ
XzBvee4PT6T/bKdTUBIbOU34BJPgOC5wOWvrwhWo6hyL2UDCQloXqPMLhlJO8adiY3TbZkn9ByHp
71aQjgc6PWYYWgDeZHC6b46TvfhpHPa+RXJAZIRNFwLsG0e8Qs0dyt8Xy42y15XV6LHA86OgdbcN
KdQ+YYBONDVnPLrttcvjEkC5hFsvZ22Tm+6DEEUMLY2+YKGb3TmVANaBeDsh4Itb0ZNDRUTRXYD+
BsDQ4KSIubGsb7AHe8tPowg/2DHcdlnkro5CxMeYyi2K1phPzeO7Yiv1rE81ikjND3q4/rZHCdy/
7xz7lhpDxYzvSznFCfzAhP0OlmUjElyZ6Vp9/AQezZrxMSgMlXITx9hbnI1YVf4vyXfQPgasnTZG
yURWLz6zRMRscvuR+pbil7ks+sbaL3WKVV8xrebGjKdxPRE4P6WAj+7ab/zXE2U6EdGy0OpcQ1qU
YXuo0pAO0sAJNFtkVLe9RxDmKX7oaoA9B2CsiED+DFu5wdIe0QuyPf95jHihtays74tWzHfgQvfP
Jc3MHXgbZjfc8YPUt4t/asRYYB9Sk1P8MRt+kD2oOdquwBfQLNO08xn3dEdxShoEHowZN5lazQi1
E/Ig9mFO9F5K90xiVxtxQjZaVrl/uxgh3Na1vdHgAuygpVHxxSXjD1jkZo7ZrhRxyX1BDhQcECQt
ES6e9LIhIHYbcCxaaiqHoBccyb2oZipLZ7csd/AQEO95C539tPkQiwLCDZKB7wuJRfYHPulEL7p+
KpvE7Sfdd2IxzMhQtVEmcU786VLRIhkQ5aue/KmgDvItyMUgjWtz5zdTw025Mh39Z3pMmBrACzUh
d22uOELB6Zppzct5AvdsDCQuqZvXucWJsa1L7Q2vNOa4doCsK6/urM7Qax2gkDIZNjoDdDs+p8f+
k3vo/utOWJE+SyejI3HQjx7c9nPoQOh3Ba04mQnrPjLB0xi48jaDHwaURFanaXplhnFNfIGk3oHA
6ro4aw8ooJdpLvZiLeuRhnrc+ROTSdw74ymEqPcIXPJRYlBFihnlhMYILCYhO4B8MJSVCsUst5y8
TjqKUvbnRYq7ShPpZcbD5SQYPC+/O6yuvAyGTYpUibdtL3fin7u2HvERdtIBB47XVeiHHHJofZaZ
8m2PdOxzFm3TxXWfV2PrKcQqYhmVPlXZA9SwNGc/H5uQONM6/y+FWTW4PIcL4bhEqxhIPn9zYq4R
kctBJqC8+bS4PKdIxbl0tRxjT+OD1jLy8WZFoAVYMLIa9tA8NtNh3093P6jxwV/848I7K9e0b3Zv
i6b6aGb2gRRdOgJiTkctz9HW+8S7SRjckxqzuF+FLgcEnGKW5dnuGt+ZdnBHC0IRvhZ7w1Emt6Lq
skN8LOS4QfIBIchjq7pOvgIqScWqRcS++602ZLJhHutHmVjGvFCt3Jg0VNXzcpFgw+t8qiOqmif0
2b6vfFcIbHlhTnq7oL0wrlOO2PYKoWvpjz4ds+Z7AVMT5esCfzKqv34DI6xjby1yFRocCj51D0Ks
NzFHI5IVJ0HWkBdxAw6i8JwOJyunfGO77jm02xWF9Yk2us/aIeq+HVJAm6Ww/EJcrneauMfPqMBx
WRKY1M4xMhu5gVCGuZMlDTS/URHGYNV5SNQIOsDhkpnxtENu3lw294XU7nK0bg6snAZeo68a1uB2
AQwZeB0iHswrodjYQZj/H3ArKJk+uj4oV5RVbtE9wraY12f2Mq7MxiHksY0gQQbJc6uVS5vKlKgz
FcHc9GWEJsfYi/n5pV4iKTabqC9eSjq7xVjSY32Fcz6l88kUBE3q9fn/tXMQsZT9IJaQgbNbcak5
OGTtRDTIDQx+UnReeln109WUI8YhzJEqUmVzHL4n9vvlw8IRDXPkHoAhIKKFigDg0HdprtjcbVtC
YO5mrsrFyalsM40WMyPo/6ADvL06rfl5rl/5CneLxE4h8Vncsd70BB4JHyiZNIp2YPDNvK2iA3Q3
lYIxsRlwNwfHz4ALEjIIpFrkW7Ni92GjxhbUBdNjxSZpYK5H31Ec4J7Tyt+WSEXfEnJoXxqxs3wW
opSNJkmk/bZljQwv9RM77Ke7HYcMIBPqTc/dbyMgUneDmmpYiaYiRWkFL6uNCB+y4gtJFjb8zy70
f+ucOZCbM7yIRuLk8jlFNiB7R8gibAGWw1wU7q+LkQqY4Mjlx8nPsFnk0pcA2oUUQJ1QAc2Idd1I
XiI5kcGnt4AKRctECZbMDCh5RWdUUuTN8ZXAlPLxMMUu5yRVQ4aZrdw+bl6E8EbQGHyzLRjSnzb0
4jZBnqikpbG97uM26EE2NQ4ZilNNov2qXPImGOySXHSWm72qiu24CY2+vOPIJqRpxnf8n+jT3dMK
MIVkWT84RPoP8fWyo+j+Esgl9/+49PYkqFzSah7rmlleYxZDbFR2VDZe+h2HrHpI3SYv5xFYKK5B
VhDj/XaVIm0xLI+45gzhsk+SJw7+WAYmpbmM/YNePZqtuogGaAKmMvEUlMtTsWlcWKmiaWGySY/n
FJabCR8WsRhVFGDJ+Bj/3uwVCUrJgp4djCiyYroajSnn26YvhQNxMmkCEsGCrdhMRZntxTpA/kWG
iTdDqkbJfIE4bZrA0958wfNEBNYF1fkC3qTm8ZyKBvFFK5SauDySfGVg35o4l1C04HPAyQCTlaoC
gwYSDGRPS6elIfZtf4CkUOayRAGgnGjdowCqzY04BoOI+UL1rP2t6Z9YBPebZaHLe0lAKMmAoMPC
hUifTAqP4v+fRZG5rVrYLOFzonQh6zUsddBQPNfouc/TqhezINs037vrCv9sqURiwc7CR1KkSmQh
Bjrl2u85uGj0rl1qbxmapOTbXEy9h8ELPi5JXfEsySZHT0guBg2iLmYhHylSIwXoJFQkacRdPk+n
bm9JKGrO+Dg35qr2+qnyeXpxfgSch5TkF0Qm6wYQtYqBd9GrEFaLefYoQXYtv275l5o7gIPFee1a
1lpC8dvTWhsDj5zWC0hBDAuMI9ZlSVLlTR32twpbvw7p7Qxnt+yMq9VzjgVmEoLWnzt9CeJoeJsN
s01mzbOfR0y/71SZVWKfQM6RHILxyvv5COwS6UAiXEk21/RzekDDR9LFU0ISPS6jJAAWzqihdYdF
5GLRfJs81JGYcL4osarLFvywtkX9eYuZM3H9xdYZG7KJxvuZ6cRf9khCNQTJXnFVG6izyk1mvILb
ozF4cVgBGW8iOZXRBo7UEEwBBORHsQJTo/lz6bF8JqOvEhkBcQUdwD3hywZG4P8xAWkPemy4olOA
eq8NMLE8W4lB6VQIxog3EKue5Mno/haGRaLbW94GzvdGMD0Px+SyRX1nGYq1C4GUPdIhICGca3PJ
ccwglrA1K7w/I3IDXQAdqWxBMqpUI8dVVjBaio3clSRGuICOygikzEI79ZAFSkOtKY1OtRKJzgo1
sIUDlO2jCuh2CvC7YlMpdhklwtXwdd2AySA/iGjUaQhierelcOcj2UhhiOmxWQfkzpyafpEKLzWH
xDzplF2e/Pv9jb1kXzAEtrFPJL0An8/TBgQzwqu85fVBUBWRh67PERf6WLZmGEYEomvxuu9u3l5b
f5ImLeqZ6g3ku9LZPtEVe+GSTvmgraH7d8OLw2y5yHYSkDDtpSUdIsF8VXrkGHEtMNngHVUDTzmx
OfWHCRxs9/FbLBhD+kHFNsTuy0f0jHS8IrFci/9l5n4+5YEgmVxL6jY8fmt1Hw37JHe+WEzgrzHu
mtaS8UgHKVf6MdDFtFYFD56B7gHszSVoLIO2f8FAC/eaDmJ8rkUmKf9QbP3spLuRRoKNwgs3t99w
dWDHB0QpX8BOpAl1Dov+D5WgH2jAbUjzU0Tr8J1l/JAthASPxl/wkyGGB10IndN+hf2GrPmaHHCK
9KVd6W8Yi3cBulLFrIgaMoiO1bsipOt7a7WP4alDEPR9iKB1pjEb5kEBnlcRB5YU0ziwNtYSi5ep
Lq/C7dowx/MHtZ1WFlADLslB3t71zksU6Us4g1eCi0DiFW7iABXwBN33C1BO2QZiYchUpv+obcv0
8foYvhaeFW6v1bIVIpMTmhHtyMP85FqoCmvpR2YfCmO3SJdhzwD4Ld4da3xcJLLKdgj5K0alXodC
Q0X4kDoF+7DAJlaWJJodLqpKotltiUC0Hjhd9gpe49f6VZ7tOGo3H8+V1Jnkv9TOfxNNb+rGO6MP
K8IJ4bgOUhEH4edRzf1wiQ+jyKnECUVdpX9pC3eqIvQer0Et9K/qjvG3cuoZ1J47akT4lcPTeMj/
HoMqZsK7h9vx/SBsfA+2k064GIR4Jau8f6Tu1wRF7bJzKbV2a1l1jOYJIqJWGfCn9cNsF+usnBtt
X5q37fej50jo24STZaXbSDJlJhmkBtk9ababDhE4+Rzzb6iAawNBRxzuCH5DM+Z2R4y1rGOekKJ4
/rS+q7+npah+/T5mZfZqqIWvD1X+pNLJBC3fOKZ/IwjaqqlNBot/hLWObc/5JAY2/lm9Il2MtGL2
gZ7OMTeiSQzSFRdA6d7YdCaSbl017tDrCyql4OpcMF7kHNbo8TJbZDDdSerRjgVKqwestEY77qTI
P8yN766jVh2k+sE5ManTvGx6UX8/NmrXnG6l9dSB8apBUvEu6N/7a13jmdeStWOuJXYgMA6XQGuN
o94tg9JWyQEotIqbDe+u37Yx9Nev+13u0VD8hLo0drQhWB6fhJCath8gOM1c70zJtYPGveayOgSO
7vot+c3JHKPzAqSxrVIkybPHdvVWaRRKuIjO2JfCpaK205f2x9M6GddLPbjBGt2m4QGyw210OaEn
9LO7Oc60VWOVD2oPCYY18YUj2UogPgik67DW77Z9Odk09A0tAP3QqpBe5+eODBtiuAAwoA/zl0rO
HIEeirC6mkiQiqc7yPJwE74vtQdUr7nbTLlkVk8V7MAjiMX89XKsH8HtRABInEX+DncMUWMHO2je
B4JET7rDIXkfZak9VvS2+6VU5FLwQC04GBPpqvaDgKJCZC5SQWlgeOQOFMRHU3JqmheXKZO4Vdbq
t8rYPUVyPS9ofTdapI6eh+9yp1Nvrvsyw0zCHcfAIteRDuoQwFl66nYAB59b4SbjxfnFHDMZ66V0
thPqhVCwE804PVdfHEhgtb12xg6aJgOUhLp1MAcIGNXN95N6xEz/453iaLiFVecD3LVTaP0DF7rv
9H4V94WOfaJgL8/QgbKTmjFeyu72LvZ+NjIL368T6FlsELEp5wQT0MsTPKTcacsHccusbAya0T1x
U/bbcCqD4WTd6GnSk1jgEs3OaeWgZGm76NZUqkHWUWPf5mEoi+76AsPQauWZcNjzNv37HSdxHHw2
DYBIOJXNbFS3YytgzmijdRjzQFNwSfFjKQz3HOSEC65VP3z3Mjb9Z4yeNfkCixPds1wIKW6h9FYC
JXXARUWPWzviQAH5qgMokRmTQymu8dUiXyJHBVAGz+nFZ119QLlAo/MCcArFfyG+thVCpc+Uyzr7
GH7w3DKZWOiGwzdEf5WqwjiUZQHNva2XgU5+NPdcUZ75Ijx4FtvxD3y85uOcS3ZZ1XmgwXEu0CCI
Z6My/8UGXOifKk5LcQBnOZzceD8Bc+Wb2g/RvfWzLE/W/qlOsUiriJ3MYQGwB6VskHOJybCqMlqY
iZxXzY0hVLNnnesR3E1QkktOdI/Uij7IOmX6/3hahEyiWBCCzjB7/hAX47vK1jmQLQIdg7GEE90l
EnQuKehLs17Y6Xyp1wt6EuE0r4ciQwLsbxGnDlKW9diPhdP3Fu9+m1f+qeZO6bcUGmVZQQ7+geCi
u0f3PqbeLrsMipJgWv6nZMK68DOUtelTbW/a7G5nLWUFo10Sj0XvCVaZRnzpnO897Oy49a996+g3
McMaR4e0JJOsw1Un0M95+CdNQV3b6nnGe5qnGCPOkzjhzxpg+CNVOoXxIzgUIdBppl6R7j/UPqrD
4SZV3X1FLuItl9ni0WhPeLGZKfv3jBH6ydivPRl92ZpB4bqxpkoYzX+9COfGXPy7QADHWgCilkOF
D9o7ZgBjHW3926gUvaqKcpBKbg9mhkRwKl9YktkO2rHLmkcx0NpRm6dz3hq/9Nms9RUhdJO1iAwt
mgT0YIU3IskMb7/Y7LZ0BZFEXK4eIamnx7KLrrkArbSvUHUnfeDhrivHg2JW7qst13dg2ppvJyAf
UaW4bYkAQVptqLOa9bvnPdNrMAUVOMwtElyfzBuM+jGqGvV56RFBRrNPnvQHgdNtUu6qRgNrzN5a
8zWXvJR4ooCETelaDcwy4yWU3mUolV1cyH4mPiDOviTLCaQPlBLLHCUhxBa9wU+yiUs+4aevyq19
W/jVZ9FeVKuijMz0+MnFuKQMUTiYkwmKEU4JEPknFL5VOfdgSQp1J9dafcQQ/yj/Gto1cZgqqYSN
9e0B5Gx7Kwv+/sGPQZFJ3WczOOfVweyEsWJNvzrebqY8DD+IrNjFZohATcifICatTMTvFoThZtPf
0fNZjy+Da6ZD3wivvec98MVDnai5vgygbs/6yJQNl/6Fqy+ATzYGxGL3frvptuCoUOfceTifolTu
XnUnn1O0kMKi/wvL9Ziu/J/0wtq423KkuQRwe3p0ABef5jZKHxr+z6xW6Mxpdz4PmQKfst5+dhyY
MPVTSl06KszM9am3RvDAvGLqrAUR+gQpb0aSTu2GWNjEFa5virwCiBNRJNRNqkAnP4+y+zeVbPBR
phRrIOs70HlZl9emwsewM4pe1lxfxZTTTGNxfLQasWTndY9Jjt0vdtB1sh8R8AwzS0zn2g+uZX04
xB8kc+dFg9tPe1mpfZ6Mkb/GOVK7xykmhxlooRKXLSH1PAh/m44+oZegDa7PbDnm4dDXYknW+Mn8
prDn57tDuOzwEVYBYmq+Xt/EgLDwh9bDdEh3ZFVmXc8u80CBrtl8YNoBRzwh15GwZ/Zk92oucfoo
SvX9j+K9fW4jvTtNO95oCNr144W6n2B0aX3SveBjUCWEOcN0jdrHTbv1jiuq+2HcKpuCm6VzPunp
H57cg1Fr13094C7ChKu/HvpOk8eg2hMZJi+JMUVyxjJNwvLEKvzrqygepWPeoqiPp6evQpfud1q3
baNRoP0ql94RtSB5gjGG22yP4DYjSGbVIv+KuS+bQIp46phWrUzPOPaeF7ZEHZ9XBfoJuL8xD8SZ
mv2X3C28y5ZhfBIrobQeuP2NDot0RKscY7oAsANVivGCCVlLXBdk3uaYZUeOeDIwRHuctBxcAzzj
eCgwDOI1QRar4quVSGRbczkwZ1xll0aCpWJ+eYE9gkemAHZwuWpXznFKiX1MMr9ITvDktXnDDUal
DdNrdt7YbDstnljSd2geDdnkPByCYwVXEzlCnVgejfcLKJb4jCqj+xT/A1uq2L4Qh8I7jT7WGwRP
rSMg7qXKp9wBCLiEMfvfsJCuWxbea6gPcBTYDTZqfsUQbO+awRu0hL+rT9Q7NMcAsMap9r+acwX9
wXNsR5N51W5nIsHHsxpCnV450rfQq04IJoYnRKMFH6ZMOVGt5uJ/zOilgDkoNrk52SgRYxTwWwpJ
o6CMTOjcc1CMVm7+eL23ePnlZvCnht72vavq6jEMzxcAYULXeE+pVNnlEMOJpoJ8kgFbl0J+yxMc
Rep2tvB6Eh/bX+D7Nw2G1CirxNbklWs9VsamAJ0I8teP1lMvYXpXGoSYIjedD9t1CoYYlJUt9RRT
IftFnXozB6/lmaTUt2LKC952508BHOou0mE/TXDdF8/OKAtSW2eNCwzca1fctGMOA6iH2lxw+BwS
Oi8WWLL6Xd+LIv057hN2em5jacHqV6b0CY7KesDUprXkOpTfHB/sJ5V/c1BWgkZQb+vkSFDXFDLY
wwntq1J5uYJpmdUVwugXCP1MFfrjewdsv1DsKGKZAssO2eID76TRNjxq/oYn7OjKcI9fF0+kA7fv
VwxKaoOvj3I/d6nFzTo6pcl+vEEODFovs8G7Ie6G1iofP1xKBkPRh4RoDz1qJmHa+pU6pzvM+Ymr
INOWkSf2L2rM+xjzM6an/pGyKn8We5bACi8xxWx1ncaTnk9Fs/YGZbJKwZlfhO/+SOYz2a0WbwbN
c0MQ4z6qBWdfzWfjD11R+Id8NnEScHzCQ8O/VUj7NisIgzc/mKTi7oUgB8o4SA3gbNu3id/wv0RI
qqOf7G0KWIvRoZ5eXLd68b557pKg3rr3Ufc55b/FevR6h2j8jbS83EwDCB+Z08o+Nyu499smE0zY
hnOjHa7YFS4M1sX5dp4hk9Pnsll0YegrYUPijq15D7eDoqQIt09mp16nUzHeNhC6HW7p9kz7VbI8
guHF+920rHOwphn/KKrdNDYF6cxaqF9brcT8rH5T64XfohafSEZvCqzE/llyr+2+yB6GX4Tf7NEa
ep/yYXlq8SR8H0K8XqoUTfpVdaPSn4ES9Bs3d2bPHDhr0fQoCZ2PF/6bDNqhV3H+KmNMGx4sL0eE
IyMZQNEXaVMCjWaje22LsgGN42opa+axPf4ehXaZS9pD/y79bUttInn/s+ijL8qinKnnkDp3WAOb
BYuXPm00Y1hsWOuzlXawhAek3Iy5xGevlvhkMHx9Zw97bA66qXmrTXaSQ1BBZ694nPXVfGeI3eSp
cTeGZjYH/y3UNjizqjs8OMn2BDqiaBxp8MWf8ZwD7kXSFPk3DFzWBxxiRqFNQO8K9P7gvTtBhCbn
kHr13MFuopOXBLA56HUUDjyHXk3pFpkYd2vXCIrDJIMabtLIvPCyq0EEmKOKeLV+nVezAvgaJh67
8odYG06kftHyi7y3JGqF1QRwHNIMoM+OOc61eojJbMkTNcVtynPAkZg4Apt9bbGe+ORfKp9YfeJJ
Ha2pTkj6FiT8sD3kreY1RCWiKgyWsycyouiPDrgbUReztW7GbEIUqJ/sb/7ThqFt1B2bZd70OsY/
2+5gD1gYyWrMMxKRcIU+XJ+iptrFM7cJF7Ooz2LiVHjS3n3V5lyvznRrJihIkmGDmgJWHKxrej+P
tcjpc5hlwqVZrStrHU0YnxAO3QhQVjiPE5hoCMWBOriyXLVkaoxr10Q4X/JnKMnmPuvVHUF2iGV6
Ryu4RsPDXZEQldS/D/pynOgpvMQsJ7HRYBtKGtvwtplMu/I+HHCK40GlBowK85xlX6MKZ2J1idt9
FmOTlP3dHwr4GJ8mFOokL7m/WyGCqkm2hNGmJfIzeyZboSB8/ELeSVXvhQY1t7L8Ijo+zxbIj8Hc
hFPUJ4tr3mPM/E7JSRNFeynLZ6FvqroQMwLKwj474FzBwD8gw2726sCXJxaWe0VyuKVx6DEyFqU2
AIRcJ8D1XbOqmJdnZAFTjIJONxnvUBbxAt+B7tvts0ysmY0sDJiJ4752J92inEwHSZ2UW4IJp/lu
3Af/mD5WdO6Zs+KRjlgsqN/Pov/IIm4Wd+jXmpzhzzs/V+7j4/VqUFeQfzTlFidnyHbZ3QvgHbex
t7umjK1oNbUdUP9gSxc6Wv2s9TAhc5RNuM6OYs9UpoDPZy6gxgENwOOp7ppxMs7P6ug6OUjQQ535
DEHSy8rJH6ekK7n2J82VFtcyjNjfk+MVUBYWwfBsyrUuci2EZKmsLiJuH7cE/6ObstpiGKZJ/KdC
xvnxtYfFiHbL8VZctuc9sMCuZrcYWts+IG08NCIAxwcyCFa1wD+Cl/NrpjpMrFVcezp8wq43T9V6
BqgIgbh9NKe2MPQurkwmYZWTXBrAn7vS0Lpzaf9iXlr/Ywz63NurKFYZutppiQXVyxjaeTxcBPg7
LY4JD/ZJ7w5qleTe20KPEs+KnUMPWcKNy9PjvpTDJCpBVzP925QK+FBkI//k1xr6P3YfeHyGn8uS
qhGmKdbtgx9Kio98ENp7cMgUviZ9At5YS4WRrFFYFsQTVZ4X1ooBNunYdbCuW5ecuBpTStLs2Mlz
GfIHUtKu7LxAbV1Q497utbhADiTTj5viUuEaFM6BBiVZi40RaqkJEE55s8OIVwpMseL5Xx+2gXcE
NhAYWVORGmzG8gukHfFpm8rtlrmYJbOL36Atbe99ds9ZmymchcOjzuDPQZnors2/20Q0AGo72ORi
olF/oyinzGikM5iPEScWx4UP34GkjmEj8c+w5kYsJm4IXZY7yVBzLFDU0Wubug/DK3LQzrTpW/Nu
xQqvrVxjy0Uc//emPPdHQ74+C/hGHlv2frV7Gb/FxD4jHN9jXO3MLiSlu/AjGQfK1Q5QydbF10XI
tRVhZEgfv1E41UcWeHq5+T+wnsiDuFLhnWGN8uYY1skKieZTpg/rBo7bIBRJRH9hNzPCq3NMFFxA
zWyar7lAiK2w/GAsCL4MbLdXdJJ/pfAk6L4RaNrob/OcPDarrF+YQDR6N9p1LQkO7MZ1HwMdQBVh
F9aQUAJWbOnIlJ0MowrQHd5i4CkIwOdJ++ScMACd
`protect end_protected
