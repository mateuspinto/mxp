`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
Tl6hXWx3hOqkKCUnmLYWmeOGaS0rpH3xGYoPCjZcVjxolKLpmVMQLe70lsMV0ydxzGQ7SkjfqrqK
oUDwLpjO5gvz40hwbnw3M7aLOSJT5D2lAzuXWiU5Fqi2yBZN/MiwvxzQMC9EAKvPLQjHhQRZWMq/
uBLkwJ1QkPqcL1vO5Ry95uXmLIknnYbQaMaiewTf0sHntD6TB/pRMeR/GOpOPOvBoTKQL3d8tiLb
Sz+3ltICnUqQmnqcNKwpqTo+mwJ3//Y3ZFDk+ExAlQcUk/QTVvMSWc3Wt6f/n3yCmEQG/mQ75lWx
hBPK2r9QzZPSybbJoHfIIDeyckpe8jDZl0tcOarGAtxxwHWorEhZUkCxY4VvW8+GLC9ugyZW8zCs
XXCzDYEH2p5OzRSeXSyrNcHk6QYGuq0KVUcFKshXU6GeBOi8RUoA6nT4N/gWAZT4rGG/yeQm64RO
25urQcO5X2bmmeSd0ySW+dKc8mIjSPli2f7hXUtmZegKgMQJGSU53Nd5s2B3QqfTU8S/j8JBkKR0
DcHQ9qLutzM52bHZnfCNw2OpmE3fPz0yyaxcE/KqrwEHIu3d6ijd7dLjeW/GZck1EW3UuQuSR0oJ
Lz102wFC3j+3Z8j7RiTgYThBriSAaZgu2lwuNYPHetYNFFR6DprCBRUqq8hbsIky2VGj0Xczd4q7
UkmPlr/gfBAgLVo6X7xiWD0XQGTgRb4OJQMJFjRRIt5DVX/VjIy1khU4wlIMdYWOLS3sJrfkmjZp
uprrCweCPw6oQutI4n4jEmooWkDG8rpXQ79kmZ7aoJV7Maq9R889vNpR1DFKNP49JzkmysUw+TkH
NR/qYn5yY2EeBHx8W4BVYGWYCu6gX3i8p/TEPHGVcbI8Ixyl4xoNw0CbpT6zzP/BA0RfvydMBdHC
3RI3v5/OCOPNGcAw6mnYaoF1gMZOufF7wpEffaZQVqBSvKeTbGOy7sycBRd2IusmaPvDEXewdO0b
iQc3h6oOGlMqvQHmyy69s4sfynpdlBBOR+pDEiPMNxGgvBYM9cropB4H4uDK/gJSU9L0/SaXW7i1
hukJAh1xKs0WbwhJUEtJr4PYgrn5+FHv8FyYSUoZcmUSfKbIC0DYbvLi2ORTNyQEt+TEPsweGJ0K
NaWrGrfyUDd5XdhaAS/A0ESOLGmK+rMrUgPmFAqCg+9mddAjvi4vLP0J5C977gKoa1ILn6S8afoJ
c/dIK6XO76fN5f5RJNoH7T5Shp6Ga/mDuEnEtnK8NbGvPs96L6olDR+Q/K3oI6y9Lt4nRET9dqwY
fgvt97sDOkBnhTSo8dvpHOmI+CBV7zkL6UWjDxyWwsi6cVvxCTrtgUthrwTDBvEuCyO6oSk9SQF/
u4dN/3JZDUYaO8Bh1PvspCMBwFYj4Sc4VB3201Ulefhefc9d3+wut3ufMYQ02Y7spgEzpV3vcrPn
M3sdfD0tiutI1aa9wOCbc38zY0fOEGHvKCQlu23gFazUhI/Y05n+e83witleIUsPeyO2BbOSfdO0
YXneMWHErKyRE5Qlo4QJhG6JuI0bAKpywHT07XqhfCGn9/5qXFWpIkddGTv4yWyApEwkpszcjBMV
npna82YlaCY5GDZfqOxRPUSOG2LBeXtnEGo+BEdq7nt3FA/wI+ooTA34kUBM8l1qbCSjQ7YY8v+Z
teXCBHf0uup7mSvhjPzhxya8ByDXYcT0pnOL2J9E8kBVvjrvTXAHXDvxrmjJ/Xylc7OrFwyLUHJC
ld9XizP5txSbrkMyfpd83K8b6PC1CXMk5w0pdkjOPEFVBkDqvPhfQzDFMR7s8hIvIognWZydiCDH
AHtoYaosTdPuxFEcPIQYIBFLXvQv1jpA4T4MyUzt7tkgUhSLMjucdDJlHilRN1XfOXrp4XdOzRZv
gGfZA34FgMZcd8RTh9qBsIlJT0f+AqKGnuubYR0OF7RUFCHBwPtt3DXhqcDCvH7tmU+/0OemjBbB
9qOOL3asm9ktroQAx99lc8f9i1LlP5xmPuAqhNXbWnZzNr1jRQ2YxGev7DXhDU2GZMw4Kauw5tVm
Cu2Oi0QRbN0gEf5a0M+Qwha2VAQCuX60npSzB4qqNJhHdN9QPA8FUy8rfv24Ak/P9Rmfg0lsfRRW
MnunCY5z24oj/S4BS4aA7Gq7bOAZEZ4o8SmAeYqY/DgKZIXuOVnxa7jIztOwuQfODt9Gvu67bRYR
r2Rp9sJxno+Lipjf+pf0mS6bUQtQyE/X/DArl0iJOwgBZfPIkOhXmV1ho2Xa/UAMv76ikCO/yJog
D4Uar9CmA0BfgiaLi+iVaRNDxYgrv5JQTAyPPhMRej8nQ084fg2v0xTaGkxYvEJcFl/zd3gQpgKC
CExSQmsDJFFhOJcnU4lVZ2MVcx9OqiNm6Mx/0XjFHPwdDH/datF6UD0dz1i9oYM5ygpVQFU19f98
WNtHdmzE9KeZJnXgNoTqSyonoQ1f/4bXMpkpEVRFKFEq2WxXZNKvbeqt45eiMSFLUq12EX/ZLsF/
ls9jLndIxgZy1kxvMMXduYC9SlxRzNGVT+xXiMaTiDfGCZXtKj6lNcml6qH71jWZIZgV3LumntLo
EiAACo7GrRm0VlR6lh8jm0K4yCbibrgBo6NloM7V//CNjUqViHy/YNDd4D3KIzG22vNXiJdl2SdR
uqOsbV1XEAvfN0XidM2JhOZUIysJfydMVCmzB58m+bDsJcgcg6j0/uV4qsQ6hJ3EiuEzyjxBe4Oz
VZvyQt1AXXQh2SmMuJGohlq7sLPJuSTNyqM/MTnP+BpnVkGcO5JzsypRatjF83bZ2Homes0NBf74
gZzrzCY92bRqCotdGrdD50QosJRX7ErzjPsnV4GLs2ZreaObXSLA4NQHe/SQvb6cKoZkln06r3hi
X74t8nUuEBLFmOfFb6pWhriZkDcILHmvzPBNM+xzrr852yVrLFagOSOdidwODQpcMwKZZP1oNXJu
acfvlljZSFzda6sDHhZQXa/Wn7N0yh/eWGa2O2T/AXpPxwFM8moq4etU5nwgAzKhiLNwnp01oYJC
T4q32x0Jd/48C7trhtczeelH/VHNb4fLrq/iLmc5xd3onmvAgIX+Cgk+LZ2OWr5Y7ui6CoYo4iIR
beCwx5wY4r0oL687I9BxKsy2Famm28zLQRjEI+K9TNGgW9RDhPdPfWe0NUlFV7sxaCGfUq7jWXxE
PFBUPODecKdsnUjK8Z9u8FcLQdr3ixKnXnvrmdhTfOYvI1vil2zcGQS1bEvE4PNOj/SbYWmj6U69
4LCv4CIjqGj6dBCjDI347sllRXn37/Ir1TpdeXM9sHPGr99ttaGAIFJf/+K7KjMk3eg8JE9rCRKD
sWioFLOlX+JavomX95ZcClGV25exKe8hzupNBGwxoBGYKDMjdiSkQ/3raaNZiPe55FtgnnZMKoJQ
VvwGqVckcT9ehos9vvE9CQXuVMNBJomiEDOKNOVqOrit4JeGCSqpAN4lkg6T5Iw/+umy1fGrRQ6E
X+8SHlmgk+1UlQtru2AMEWBBwvPs4l0RAkGOwqBWgjiBk7Z9QZ3niaACOKPBOQ+7BLZ2zyWZlYNi
TtXirpNFo3N3fybZhXYNr5xyOTQ7fWW6VebafmwhjjkMygBNVHi7CyEIlV4c+D0JYyJYPqk/bg+t
PU85+YBOaj3wpq2SwfsgxsRM2cpMyocdIHmPPx4fwYwbWJ9FOLI0tjYAp9yOJlr/Qq4dS/iVowJ0
SUc/1P21r8Htg11MTWctzPC85z8t88tRyK8eJwYCupX4ErODo5Vl+e76G1Nqd4O/qWe2oiLC/xdI
tkBUGkJ2QqxhJSpCp6/LoabzfAj94K1ayXuQ5pmldaMWrIq5wso/CwGDfcsW7Ck07DvB1L76urax
h43Rx43INrM3mIhwlN9XiiabI19ckAHO8tSD/XKd//K8zuDTyKlXA0L/7hSt6/Gb36c65s6kK6Oa
xzccX2yqJqc4FyS2984RE/4q+KhmPC0PJLJJyAQwxmUo/F/mRi8x1t2G0r1yLmxnn1N/8dXI3Q9O
J3rP9hKrOpkYnUvb5G5d8KNt5W2AOWoIN/hinMJ3TAvHSwU+6J+Xnbcwub9ukekZo2+hFhJV17iQ
K6I7X0P4RymXky37k8A2EfCjSc4RPEj0thKaSf/jB0zZqzLqo5p5KoX0i6n9uGdW2hjzlaPkJIwb
XYm+zqs6+RhLkZUFn6+f2NNzRuNAzpI8qsIJkFTYJYd9NC87wn5PjYjHV/S8Gri50ka0kiLkk9vM
DoDhsx5q/0Sr4pniBKhKnyTT6VkVpNIe8NR9nJ+nh8Idwop1lUTfw+gNhLZmnLy70v4B+ZnLCE/8
AWC3pzd+dccLuTs7ozmWn1LWrXIwpCIPjxVEV37x5tVDw8H2EIyuPQrU3u205iNFY1EehvDrWjtZ
vZRGnTfSCBYf7h9zbo0kG07BhO3lkF1xJdEP84x9+pzifBwtmoFKTTXHxq85MVvVGtghi27IMSWx
W1P73zHPoK0hcRYzf2WiYuF3uPTjw1Sr1GV+ZuGA3LzUTuPHnHbZnwDeClmezARp9GNcwUVFpwsE
oz5F09kD7HJhA56ooNXBl1UG/rDw3rIROtF6mvpsqkMgQOLBPei8Ka0eQGuORmX/qx4FSqMKZmkk
GpyyG3gMMrRAvvu33A38yMBVSs2hDujzufZ6S6MOBo6N+x/CNgjTB/nEOGXHyssieM4GmTOKfbhI
RER5liJbzTIpYIPsMJlEuMZy5Op/pMR5cZqj/5knSFKYDM/ewn7wzFnDSgljMtm0vrKO7EhCIyoh
VGd8Qv1DUynRo0lD3sB4IrCAG2h1cxKQmkPzsipm7TEvSunNvQWk3Qzbz+v/k9pccOaqagh4zELj
pHn4LwwOjqgQrvDwe6LLrUm/ABkyDrcsyvKrxDomZnieOFGEW6fKQGxITxhIMTzp8LRPhMk+6+NX
s72DtCFstigIYMCXenzs4w0tjHT8/iB9aV1DdVuZQh9cxxZkyZlDPf4tbt/fGScVmp0cNSCWANYD
bR4KeS9ZlojUeUFYBK+isJWJMDPJjbijcMXCFZnnt98PAIt8+4qLhMz0cYob2MToHhtic9GeXEXe
avXRIinXybCoTVkrv8yNVpPmUhX6y9IcMDRYc+PAGfyh6rms9/Y2atxtVwnf2Dg8UPoiGz8BONMq
gbXPuIk0/u62A+tWsKXmMbcuIp81y+YixLsm2CpXYjSDL1Fpw8WLEgQoB/WC7XFyNn4t4NI3EbgZ
d0qhwFvBxmA9ImaabDh6bqaL4kJDGJzwGE/an0Idahu8KAt775mXl5X/RiUjXHUdmcymTbAj3+9o
dSPEuVSk5gInOLkOCnlarOHI5rp+NHG6FLmt/K9fH1EppE9UaKIv6pveFkD0fQ4Q1MQl99sQEi2x
nsd2rSGB9V2cLR75pFpeJZOPnC89Zc0BT32GXAKw478MPHy2hhDv5nLjzsTGwryvwyWUu9aDR7TD
u6j7912nExNGWpab0Ij0PY5eLhKzHjNe04YuiidIHFT7cLKuzJd4WUUD+KbXUaFpooN4PyHqGCWI
44IASiizmdCa1qSvux85WTrwCWhuh8635GdxhW+KwBFoyEGFaX4agSpUzktHWYO/or/qq4Vy9XLx
+XEcy9+ZnM3RJ3RHT600BkRSj+StxEj65xDgS3LPF9RbtbaaoVNQ/TtSsEZQUKHC7oYGZtvfbG6u
akleTbRdGco16G12DwmOId7vem2bunJfBA1SimMjX57qKKQe0k40/Y9g8puaZpeqtYT7qux+xgq0
hSRshmUjmoNf/0k/ciIh1WRR7Nlctz4QZEx1GlLElIUMTZvs95LxHNsIaOnqncuQ/uOuqgaJvWc5
eA1lCkPYWVz08Ts14D7r6QF3k3R9vRMFoDeA6qtJFPlJ4u3fWp0Lr+mL3eNuJ5iIC/kenZbFAeds
p3SZC38dgLm8j5XAn+CxyVkKx7/TJGvkAprKUIrEwxqiR5GOQ8iDyQ41SXgya42Uw68ynHKmqPE3
BEoXkrBzYx3+Bn2SOgGuqvXtYEe8lgMCF5uuTSLnt9M/62LazYs1bbBG82VaBsf8dV+mtViAN4Gl
MGEjA4JAr7DFLWavKcn+/OvsFwkswXLNHBU/GbBdFGDbQyreDIuNHe1uPQGPDcUzXE+/1Rf4tt2V
JTiBLz7K/XCdv4TM3XxyENJLIo0+gfTt77Mk/uk9td3By4iHnFx7FfrAFAnYvCjQ7Hpfb766tOw/
4esG0GAWO5hFoqX/4cV+cvD5YuOT+P758IBj18rbasMG1w4G8u0WDmuxNgn28r9J4mMMgfq3xrqJ
SUXNei1mzOsr5hCMbOAcoqp6L2iXTjVkL/QsYo/pf11pViIrDqzWMFDAvcllqLa2pg3Xb2MbC4PU
QpjUEI5I1k4ddaD6VJqHC10pl5D6vYNkAc7uUmp9ewkfP6Ho5D0+gnT4UvUxqoBhF19MjhSFfhUP
sOrm7Tcurwq+uD+tTdlR6YsYAfpnRUGk/Fv92/4fvX6tPAnb70Esv5QXkNGA0GWKS986I4YykGZw
lyQJxBjGXLZkmS/3BYAXYyMPzVhQU3IPhg1AV6v6kdFvW6thqGipoQtPM58KF1rJD/6UsfgWpWIu
L3CqCaxtS34FmFyyYj4qxiWpJQMT8n98SeuPBk2F4oahzl4xxVp0vkg8YSAla5E+v7Ja2tcbVZ4x
GMFoYH5BeCwimzXhDUiDtc1Z7d3LCJHnxaQrBuWAmXWPPsmGBC2ZccahRU2Wn14rzOc4HDaV7E4b
02zbeQxEZcRIL9TAJJ0nCyC/buhgZN/GHRLknahOdP4VLyLCThZKlSChB3bGENWIQPJXYb8rs6nb
DqbgNgHOU0dfAg8kyWkfZNvAqyhyeQNr0cPEJ4+TS9awiidl7VRxiVqkYumkCGuu/B+DAP25lXfJ
SFI4kPjR7ES2YTsDoqxbCK/7BmSXtkPhTqDosE9BGj4BVDruCJvoI9Ztic/gELCS0oU6E/8L211b
JGFv84PmEhhgEdYUAICymNr7jmD3ByBGiQFCWU75w1Esh+tUEsVfKz5sD8lE39UBXHJlOrovfqpc
rsiicwr9GhtDFYU8tBU9vHIOpR9qpW6T0Yn80823JN+gqa2pb0vRoTpnnQAQW7pvK/nKuDTl+wLJ
GtRJVF44JSSWu0jPnZ/Q5PVCEGdyZYAgMAh89r+uRlYURo/bCIEdtPGBI5gtIesUVBmFJ/2R3TYK
ggCTsT22s/Movf5DNFF0hqEaQdrlnwlBU4ds86sUxEooyoyA4EcnuGWH+hAgAefc6px88C+cy0pD
tIvk09pGzP6I/5CgYrcOXmJNGHT0zYJSWZURKzea1VSwroDLxV6ArTHlylz12oXRUo76mzq1eGkI
OSHtbliZgv/lZ1a0g0+2kw0DKqR8QIhesGwEA2ggKwMHmYMi0nBk6V9kQW43GoFO4x/IsOy+AMie
tth6Ske/VbAoI1ca6QueIDLeHn4MrXoGSa02cRaev9RavTgth8Ru+E0V+0sfoR5NWb/jXxr36kR4
JpptizelpEuTjXBsHqPYFxVbqkDQjbSlwlheoSeUZPXsI3iL4evEbw+00lflYRO8hVIciQw6jUiU
riv87G0MXuMCwaAZJmr44I0NuRbFyDppHHfq/EIAilwiTcd7EPRpO0s98AnANAIU8hzJNQgKnDMv
L1RbcFII/bodfwCY3zuF2raRB8UvPDY3FVQqdKlNQcIpIyoW1FdpsriCyWZ9A5tkj8K0BASr/pt0
Rat3aPIt/oPqN/0mx2wvGbGyZ/cjZ0p6Y9Wgw3AqlfeLEw8h7nAY+PPV9XdIacjTLfJszhAsNCAc
EuCCRsCuMQ26nkybgd34yWIIBsE3xbSlJEE9zmXpwtnZCb9eun1R0z5dDa4J8pLd8nB58m+FZkWL
LN70h+LnnOWwSoPoQ12nOGj9hILjefgUNu7AmB34M+LH0k6dDTX6XqDwyyongzGc/pz0NYGsRAhb
T1lNSShXWPqt1m1N/V2BDOzu8Ds4MBA/wkGTGqs+1n95sAhNezn3JTw5ewr50so0PssG0AYDn2dT
16J9bkrkIXngIiTJ3e7kUSlaS5UUr/ONA55vQy/3Sh4CAmX/qk/1lCq+AN2LNm3uyjyiXvWEVJCU
m/vwgAv2hj8A8QvogILm7gspfahxu3eqdQngkV8YrB0AQXWECynchvv6V0uihYSSFf4AC8X95cAa
3zyoq0XYe0MCYHxtyZG+bwqvGCV1OPEICvVpH3KpgBHQMhAMvOX9QPdF+MLGsf3yXkwC/CqbXQFB
Z7iUZhmWTMJxyBOUwjRkHS4VHNmfo+Gt5Ghq0p0eWrPlW2Tb5f4FtT9nDw0c60ZoEmGdQF+FIr4T
B5RUsiSnDNoMX1ggFVS54cc8Qenf3Y8cWJWQllSdnJ89CJNdLHZwc7vKcMQMU/ZzEXyspsmIaN2p
bWHXA34XdLU7CSEE08T6Toxpj3kNISW2SZaVrHaVfE5gZpfY5/5MG41Mr0V0ArWQCGxoItQ2yP37
uEzMgElaF13LuEtO3VIihw==
`protect end_protected
