`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
VRbrYcSt66IlAyRdCkmAm2Bkw5VWCWC0c5Ah20BG9idXcJO27jT05bJSUOzlC6C+D5PXa3T7HkNl
SiDVVRLCixSXkk6cNe+3kPaCLT/1AFkGh/0St8KAvgyXiPu66HYKVtP0yf2QPC4bqeBfqxG30htG
9k04ju9P5txJ2l1gJVGYH/ShGZEIxHRJo3SKF81otmdckRqforRgwoLTtCg/jbjp8g83TuUfTWPr
egc4BDr2hcWUsGqTyP/Cex+78OBXg6P2Yb3qeOF8pQQqFW+fxyn10Or3RzvVyySlinIYYqJufXzd
mW4iuTSsIJUmbi7pht17wbGqcvkXRWHA+nkJ1fuKRnqPBcAhPagMCEpuhVIfBXMkrSuwTm/3HOEr
KtIh0nNsN3benk4iuNy05aE2uaOOSY4kGy5MP+h9y0VvuPJQdAw3CHgvOQxfyqpCr2I40WH5K3kh
VY8K4JFV4nXtJOl8Zk8v4kIApKuiP4FmfnX8PQASTHgdpmpn8VIOLVb8B8/Yfj/BRh4DJyeX/6no
OcaiJGt+Kq02375oGZ5hzdpedCAc3bnCK94R0f6ux9jw35FvXpLnEEE4Gr9sJzUtoXX5n98ObiVC
MP9/vpQTmVHo264r8Xp5TD0ax/FfJqkMaxctTHZ5XGEgwMjuZUr6ePCrWCXfia1ZwqIQo5KEs3o/
JBf4NWxgm38/44b51BfVetBO6P1Dpbsxf+jMmz8afVlrLUP+bj8Hrcsj8/gicsatJ6jaHq6uL01G
XtyYYA8YibynatWaWrCYbBtM0qa3HvxNfeYE67HpthQllw1jbv6rJykbEWTBz/2rAdZ9AO8EXTeh
L3lCmUZj89luymTH6FEFNJUamjAsroi/WFcRqoA+trSqGzpKtNYe/WHxTvgadNvFTXYXKj9Cgk96
lSjPSwialtkHk2cAjclxDZOXRQBNI3KFHk3hQfVxjp/7sh8KT3q3Hkj0Au2e0AF7r/D94XzGv6zN
ObkSflACRmsnEVFx9bYQpe8WnD2g9+pkJndmOIioCsiUJr40DdBQYCqKS4syI7wpwLXVjY4bHMel
V12rY57YaJpdEUfYctUPymSuZMhtBzJ/pXViKzl2rWnVJkQb7Mq29L99KiZRAEjwec7jpvcp591J
tYQymnkye6YL9SPbLCwqSajT+EVSw7MwLvGP2/ubyISrjDvp1EThL2lzpiBZlxbd5Lh9HjQQHZ/o
lQ2nm/8JkyqXkqSrozeG7TbUNhJW7K9iPupsenG9C+S1seT39IvgDq6Gd39k5aoxoBloivOwQis5
hRECPYr7fSGz7hcEp9q0P/eTlyPhf3TUUky/gbO/weEzN42nNUaQbI07K7pleLQcsvJXpVmeqU8o
LLcwnuZGy6MMlVbZRhgYo1czR+ebLi7ikVfhVc4qep60+qbCMdydWX73EwnI9RavO6LboozLvXBD
MWxUfVfGYf1PE97CsJQqtfhnRhsCl6MlinMavM8e0Yak5GkSRihkm6ny0kN08X4eC+MxlENigqMQ
/AHjdU2M5jNM6EWbDXRUBl0C67ZwaO1VojXYkn0IkVnuE5HafFQQ4Q5RSJuFuEji9dSD+g3hnJGA
XWl+g9R85hRYgSb65XHp07ThPfbuIFZCDT7yzE8Z1Xj1+q9u+q4mR2hjuTliC5o27dXitiTwfg8C
sSwdpCIiyT+gEwmAM1rbwL7SnbeGZ5d1RurB18m6GhXIFXqEpDQGQO4yaZIud7PH7nopi9hr1542
swNnV1Zqtj76qxzeKu7FVVtzyhzR6hkrN0f6Pr0/L0n5okIIT2drH5wnJ0uGG74zFcAHhVYT67gz
P+4FAJpVMcD4XmouiR4GsfZea/gH9oLokvinmlO6Mfr82UEc1fmozi4mRUVDgeDzMmzXB5RL4oYj
RtHe+DZ7aZicPJMkHgAourkN9ZH5NfVDrZO8qqeExx3XCmTRtsYOhLfnVeC1bEfqenvOpjA0bOrH
44ZDHvkEadfcwqqO1J8uPpSQGhcpRJmWvnGHA2jRqczII/J2YnfjG9Q1hfV89hLHC5+qZNLOhDxR
bdbCF0t28dsqSdlVQiveKW1vinLAmj9NCQLWMEGh6SrpZdmSMpblfIWoUe8xees7CHoxkALkt6MM
o09qaVJjlJ5ZWVC7+a7MV8DbZbqDGYDQ/ugSw9LUUgziSMaT7VU00S0gxlQtNdAwDM5aq/AWt69b
cwLibqbu9AwjrUTUogmxs7yHZD/07GgJjRsC6e2IUU0tRXFS0JydGsJf6TTxssYMPhMCLQMiNjVg
rjHBpYFDZJoArT/rC7fZZnElTOqjik6wrtm2Oc6jPPPbcTUwFCKN32HraYPThWrZ0+DN+FgnFa4x
BwYKwQ1x+6+rfq/kD1iNcKPIm9d7lDpZo7OE9NSdO8knj6hg5q2MmfTCEtbW5NTzgDyh0iJvq7iG
esGesf8UCULkEuuqItYwEMHSG2HgB8THRy1Wtt+cHTkFGdERv94+/Omg59rcdo6pCKClut2Q8yyL
G/Y8FkuRwVmz+WJglgSMky2nk1Or8j40kLrcJsOfmDwKNEscXUMdGxQFPbYm70d7/wKIHX6W4+6P
5/8EBwaqa6Wcp/ziAD7+uQ32UP9t7GE90O+Ns1QK9k7ISGv5M0UWdNy8X25oqoUvexML5ZCdBq7D
2V7ZdZorhRd8iqkE71EIQpoXG6dkMhjBWlwwB2Ca/FrFvdNJB4SNsB3kivgzI6VhGcd5VbckwJ0e
qnOWN7r/ldpPMYvpQKmGkHgw70oaPjG5irwSD8d5pgsfQDPTCEURTBU+pIqTWlNloE1DbUi+NRt7
PzzCY3NAv9caccQvwv9Z70rg53RSnG4WuPaAC3vXTtixsRs+hbpKiS0crfkfiSfdTXTWkYhdtk7C
m366qApkThpGSFYvtVShKpY4BuUuKrv/pHHmSOynNwWdO9Ia+MRmwqlLyAmKrC2hXNpS8t5Q+fqJ
DlFb5l7gwtKM/IOW0NP0a7SZJqN28LOI4blJXb0XnmTWHco+Zc81aAgV9bBuo+wF6UO+tMHp//te
NiIgrkeF4H14uOdDiCdv0yLk1DwPepCuZphuEHOadxrzaxdP0OgoiLDvTJLzEJ7Ak42E6CzsWVYP
BE0NEQKLk7bZcCHcASYDlgC4XLc4LZQ8qq7mUhxqlKHEwMju7FVxLz2HNxqbbpMmvr/bS87jUX19
KoJrs7mqWoAC1bhlmwhVpRRNlaQS5o1vFD+b3AB4EQahFS+vvv0RdThTotGFlsmz8TTOL4ixFPb4
KlamO7mA0DI7kHR66NIezZurTQSjXOkooCUrpBUXgmxGh30shOzPmAFGPc8XmbQTtlhhzv8WlT14
nx5oWYYwGDyysKT1xd7PrLY1jzfCWJvBs/aYsCqOvQOTpJ8oLmun7FJ01ZtSzb1+VUMcfx6GLUG0
hyRUszjZ25j2vyaiQcbTD5fJYAVP2xFGzemSmwhGiWTynC9EQh9H2hsmpFIIvC+0twPpJWwVFrMe
XK0OI0qReeDkAJ/iw9mT1H7J5q16J64gbixM+hwmAGN9iWlEVOY4HUDJlbWuDkh29yHRE1D9dDM5
7XAnaBZJbkkZfGNDq8DFLFMbqghrsYGlUIwUBpbMYs3O+PBoQZIKWe+Hf6ovKu1A+hVMBwRMnB//
KgrRNHg7tY+tF169RAGGPYmSzD8pq63leVu6P8F6RaIWACuqfKy12H4gsolIprXW7UDzmKtp/iKW
aim96711QHUW9K8XIr9XILjcfQaiJocXqL79OJ7PQ8Uyf3JvDBKbE6DOtWSlox1gaQpNlSTqFRIb
8WwlBRcx5N0pX/znGHNYZUH6lJr9+AN/fhXfVXZGZHa982r99GAsxjL4SldbvObTijx1HDGxaEM3
hfTtsyHMCxWGfii1vD7edE4IjOTNoy0SJ1HMcnn5Aq/5/RAd4WGSiOtI00rpKOqSuBDGZsV7Bh3U
qrGx9NPNJW2jDU11fsaH4ADchGchQb7Zlhqd7TmSiapd/SZWpOW0qwsm2bbSar5a5bzHOBPXztwF
i6s2iPccWIetK6j42vQT9VwOmOQSBelzz9yq+2dD/CKK3cJ8eWnsdQHvQVvjEPdV0ecfe1c/Fdwc
HKK8gWpayqPMRPRNhdgOYNeKuWRJjq5+heJrLcqeYBszU+r4f+6nqD7KlWAhwcWvLQUmqzupHOHd
Y2Zr0XF3dnH1DalsuzjHoh+7mKB/SqoD+VTqZf4kiuo2qG+vk2ojwNgc33prETR3iiCdMLtFkyvF
U0vbzPC+CVuXk0i91U776LTt+tICxf7o4MgkmeQrlW1jISmWyb32b6qlY5Hx1Pp/3Vh88Cs/RBNo
DtomW2gRaFjMCarvM5jwOxIAksQP1+AZOhb/ZVvijoMxWJpkOTKuIBg6uoZ4usjRVF+2wbCMBp+Z
p0CPCUTNr9uuCeK5vMoqazZIsH203CUpO4GlbRcrSsml6GZX2uNk7qeM8vnEfUfa+whABzT3UdL5
789L+UCUvCZkdWTt8JwiQ739Al3+sKKJUIJzaFnMAFk9mMEGnieVpVCEZ19NZqHwtZjcFqdByWsE
HicZ/VIfKBb+egCmRzUcp4gMKzO30zZq/4T0wsy551L8lWmUG6Xu6MgZcwgoGqadDtiwXN1Z98+y
4/tQvJnDcoRXU6rqy+RZ/rHjDmjlXrRuQaoxRLoQM+UjHNBcc7YjY5Bj1JROosZiqKbnxzBXn0+L
IrBpAMBQf3qgmtvru+I20ZLgMDL2dt47zMUthVlf4xODVhG0xlbTVtjEyJ0oW5wyvDScTZ+ahGev
je7xlDSwqT4382S33dbjPFv8w0n585wwremJRVdkG6fk16+gbuxrpx13RwEMaK63spRRIXUyeyB+
fvl4lKEMZWSTYh7XzvYJmufhC2P/pFJvY5abSHcT+B4W8XTyzFILdDR7pGCS2PI8ly1/uRo2g9ym
/DC/KJSExk/0TM52wQrhL8T6StelpnNKhnLbHnqYzh/dJySlbVWpmEe2XkA0qLi9L/bPwJiA9O+2
CiLzH2pQmYLMgvmbgz4um1JlDQiHEFVUJeCUmdnQlA6TzIPpaCg6+ANgR+DYUPz5KxBfviTuP4xF
w2kerNt8nYUeSKlYXY/bbfrHm3amDPwKMChkuoKKh8kx4qd9OM1fh+uqwPjOS/HRBp+7Po2zqAdd
B9dSyC0y+xcNko7+7lnnqTB/9OrCEGt35MbwWSGIWNfQeFZPv0TBgkazo9tkmWRXtH/1h4yR/r/O
wQGUXqsFWdmz0VbeID5dh22IaFleo3qNSVKRyKPVf12ecqXXY4tLy3kNuhheuao/R8oeW/LqiFmY
7uLavKd7eBJWlpocDkOznLvm5jnZ5ELD+9yrVS988d9/VCcZujvJ09lsLe1WFpVg2F4uVFt6HqLm
n+ERRKp/ml008lgeijTmfKkxGHFxoh10WNUzFDE0mLwDShTcvk/8ek5ok5ArIWf0PoQ7M0Z6Q6kJ
avIbupcagPy4zJhkLmQlFyeUh/oH2a1wFvBcnlGJY+LdKRbRbELQCx+gIEe1vdSFT8NfXzb9gp82
YJrM53Gzcu+ia+qxZLeiL4XWtpupbQVV0ZF1T5isxwB/IvvsTneR2+qnoZAu0jDLBlz8GxqtZDyI
BzCVXeLBofKzm1I4BlczBy/HWF8mWmwSnLhhR65kaXjcIngbNAKiqqnXF69HYLTBiPOVCJnaXqOs
Zm8GbOfnXrX+X1QmZGjojEvKEmUd8EstPwCuypL5H1NY8gdJDUVTeDNOIdLHlu1C3E7MJVtOm8t/
G6q8+9kRIz6dp3imHu+a5YLYnNFSdnPdIWrZZj1TKffavE4sDjg6aee9d63fZzNZkvB9yk7Bjp9f
KUB1hGgq5CXw1wNx/GSwGwBd6aeD5iZ8dQeIM42OwFgg8jlEBgC63cYYW3gTAwKk4Ne1w1zQsKch
cijad9g1XxyXAixTRGyl3BK8cMr+mYsHdhBhDpuGyLCLGhzvIvGYdPYO85VTRh+4YkVQOOqHzKuC
goQqfimr9x+BYvIvmBvRo1A7KDGfcVm2V4SDpjyHBK8VdXDVL8Odf/IihTq0R8ZZVV20mLTbV6eb
VFscAMsJCtwdbTgaevEVagDYHBKmQ76pVypOSyhA0Sujd4FEy5k53/mrgLmoVKul7WiFkBdjanJy
FStLeTuY672Ge1G3HIT8JMIgcpH821ASxHiex9aXDi65TI2sND5ClOiCgl6UPkEjR3uQAUn0mcec
EZ/D1aARmwnbpya5/vwMicV/tOygUqLMPktdOloBFl4SmbQG069EJtkVjngSaZW5tFnjMz9mpYA+
re3hUSk8W9i3Dm3Wd0GkkS3/1kbSY5IJgLYpHoMJCR2gE4OLvSbqk4LKBVETSp9OgxfAoSZ1pcl6
M7ScCstY1Hud0H0YbLHmLUv/fghL8hAX4XyI3DAIdqLuV9pTlfJawgYE0XtPD7CsvAYOULfL1VRc
FFiyv4ck10rLiCybJjXi3KKZUicrJFTKw/fJLNPa6eVgBgGPrr2RPkAFX9eaFU5FNol+mEo5GW4A
Wrk5GqOZ0t0ukZjp/NISmzRU+U/6j5a930YLx9GXLEHmQd/OmgljQJ+kJZAHC7+cwrkwRlGSyx1l
MEIsywWiP2PBQ8rEfRnLccFby3br1J8cdYqBVlotfauACMMwdZrQW1mEQLVKyNkai29f/N4gPxf2
gyisZBuD/ul2vGwl1nW45/055CeSuLIduDoGTif9LW5/MnUuD3Vspvv10wcYKHZ+x1PVtMlQjAOi
7e32bSBED4K02WgJ71id/EU4cBviQ0jpau0IIH3CKoaWgdnpy/Ha9qVGRywm3T7NkAdU9M3fPDtG
gbvSPKhwUL8dEkKjtM3asWO/ZRiULg6uR2+v/zZZ1Hbk1WFHOQ0b0Xe9VU4nL6Ym4cZdWYh6+dfp
d1yJkZGkHNqXAxe8uJQ0awsdmQ2WhIiS6wsMmydY9Hjf/JrDyHMWPg4TW2MkaZQlmBWpdNIX45Kv
7HUmteXJAy9tu2lUcrCybsLezsTrRLJZ0R4uFz/worY7I2ou2q3yak2oScABQT+5Kmes7Pbfdhsn
UefC29DBXRj2+W6nujaddQEE5NkvTAqHp/WnVk+wERuKvnINjgwWayEWsajhtDLlzwa3KqRDBipj
hZwralZCzRjVfwtWAW3Vi5MUbDQeBmM4pv3uiwLjuFVA+jfLGepYP/qq9hJ8bV6uWGoeg51VsgGc
9TexnY9LDif8bCsud8zm9PikWASQEgy45tTxxvmOtAAQ8Ym8BbTCpXAXTdc4pdJAIBTdGtvk9ywT
1GekdR7Btd+JfHv2qC90ceT7i8UkA96EJCwz+O8uRI3Za736zkLntLBV1CrD8lbx5QGpaw4/txCA
Da8W1aWR88Sie4wEs+ztYYvanls1yD+dDt12lNV1tf4+e1iVvAY3rRasX11uPvxwKokPylVU14db
7nXcNfb0C2m744Ya9FwruLP1I2LuHDMdhEDUAn7F0SANDYa4221rQMRtOvwxUai81lyyeMIqn5sg
ANrYMCVc/ikZudW6TZZyl/fqX7H51Xiccmy8N5gPUWXS+woYCDtWwqrPof12m0/ViaaaDR5+WvNU
ev+IlMBi/e78dzj9j4dy0f9zkeDhqwieObHibhNuhNh7HUpFbMMl5Pl7Vv9NA9diTopZ1PSS6O6p
Sakt+2+9FF6txrdh5+Yk1XygEOSyzSzMN00+w2uC4bL6mlSACtZk3nopGkil51GoXzKYUJ59O1Vm
7OYOuYqV5B9Is1Px0aExptZceFs26jsaZjpPl05Y95D0rTaWE1ZPD//JA+Kzzb0eOcvMACT2NzPY
pXO2uweq1BhYr8yHsxsZZrRHt/gijGL1BxtLTxaGaZTk9//zFcVmgUM3x0gBrU5pcPCmkJYzxzxf
MU8FNjsxkp8GZ4uEB2jPDQ1FiBzOyWJl6zzGGyRfsFmBRcbskmgrPTbUXHTlm09LuQKAfOgZCzCD
rkW/UiIsM14/CzLbgCi1KV4hpzSKUWGSPFW/WbAq65ahSrJto2YVcK8NfyB6W0u0W5UOzChQlXOw
RbHOo5WrYNgXXZu1q7Ku2N+A4l/uwN2MIWVdTNKnnG75ivoxdm6ssvJwrmnI9jHwG0y2Jtw0iC7Z
XfR6OHPzU14PMEI6HohcmW+fVXt/2Ly6nw/hoYsu9SSuNQ0TIHqbt7Of5qjd4ZDJAy82maDx2DbH
AT7tPqo+u45e+NRYtCi8Wt3Prkj3Mx5sIsTlGHECXBjHAzJieCxn28ZPVLuCT+fcxi5lbwD7F96k
pGr7lvniZqs+JxhC/JubTmmtFFkNsKWD/4wOcBRioe5rLbOjVNMQ1pC8zSqEap4RbZTu17X7yS3t
wWVI1IBnza4X5Q0gErD+3RSXosQ91Fx2SfH3I8V3BMc1j9zvqRFmlaCZF2fxuNu4qgwhzkqRwj1q
Dcv1firQVEbOOdoXnO8aSPWvHOJUJANPRVzOflP0+UyGXFNU7ebkPTwMpsNbrd2sdMKaZLbQBrk1
/jsYfCAEDMyI7kqqZayzDOgq7nrPC5Q0MtlLzg9a9hQKBtLBnUq+uHNAh95lSmdoGr7gz1r2poQZ
97LeRGxaSeGbxXvk/AaFHXbC/6JGALRBhfEUKVKOeXwP2Jj6wkoZY000t/jbMUzSc4surtdK/YOw
uSGRKIkvORVqdLSpXyKJqmZhlQ54snLHuZ19cxut/3IofYC5YzArJtsxK0KKAe3n0oIJ9+q57ECZ
UVmTMzvLce2yQqn2y/p5fsnTJRgEES40FDMnOWdNZ1m+HOApA6/wWhD97nDfY2Cwb3EsHQCqdDHx
3NgChzDwQNI4hY4dcnssHNo9gJR88ny/Mkg6411MCOyIpFMzQ88AhMTdhRyI42O2ud3ZC6A66Cmo
nDFc50fOI4iiiFDfY1Oh1XXoKC8WbJcH/0t02NiLDYiccCfijbnkN4ZcOrruaJrSvHbeeU1WRR6W
axx8iEPdPU0BbddDnlGRawS6XoLOpUMdD7rHrvrLZ0OiP+aeOVcqS47XQ+rE1jjVspLlHyr5DvSH
y1rAsJKO9MUmJbS9e0SdFb4fAmChnJhlO5fQaIQEpg0fn7Nv4L+hPmM7jQwfkpdNsPjhfCLb5jU8
JYApu7tbAFG8WThJ0rDpuzFq06sxJUnxmV1Kz6Fr8jCovxftM0hkbidG2wsiRO7g5FV0cAHh4KT0
+9b6Cr8LXyGEGl3QBajV7eSa2BtPS9lTcaRwrJS5zDX240KFEXabJeJAurKL+dg3kPoeBJ1HwLkl
HAOqWwHeLRd2k2wxrgooSTX/0hVerbUer531Vh7W+ZaPAwCarKd556YhHZdKneRWSHBL+icidCGs
HbsU0ON8fZD5sdVzrArcFE3biDFzT+RMb1NIKIC7BVJLpbprZYR7BTIhk1U/QEtzd7ucYbci0rQb
YQDeQyVl5j9F5m1bnuWeDiAUqaoJAcpB2LNX8M7IgLh11f2k/nWShNuyp+PbRbvAjy/WMoy9hT8d
4RstfHMwB+xr9ZL0Dj5oLPK/zdBrPn+XvEaL2PiAXOjJsSw/a6h7Im8Gxip9yd60nBc5gor2pAvO
O/HvWzqRGPo92tR5I92fIX8BHsmIW/2CzX03chtAVdwmbpK3MHksGVslqZGp5YPwE6aPwop7NdK+
3ZJnY88inY/ojsR6u2C1KKAkqJUa7mGOxqBIIMZDIhjZTvtrSt0rrCY5nwBvL4V59mZmgsrZNHIU
OZODxDog5dpfvSsuL0w3kzeGW8cRlMUPCUG4eqfl4rdm8G8Ym4nr803lRA5rA/Ockgoau1aGuRn4
MN8sl8Jb4SQhpMVElMtQw9NgGkzOjeXzLFjP0lAeJwrFeP+3GAYKLsK42LVbdpyjV0jbay5Nipr/
BYEx/K9tdj2aDIMtQHRFEdfkO530FW6gzqb1sZduUZ3PejGmNC/rXRsL7F5jeIbPgjEkV9lTdkII
f7UIeiJvDNJISJ3FQriXAl4EenaWA8hSeM9vThdW9wSJSPpXaBXhBWHwuLI2sDI86gTyezekFm3n
fGMo0VRQ5mPc5/kvsa9gHgPJyq8AAuhmr0eTB0dOZ34hK6TBtMUHsBWjEla6X3VSbnLJt0yGCKne
ItTRBjpqkA45dwsLSw761JfL5JKTuLN+zm7pGDKPm4Iz/Z3HZL1vVOVVQKNnPFcXIp1kosDOtTXt
sdB4T8MJwk21w4azcu6j5PLK+5/ti4EB6lOhUw+4TGFLEI/zb2/P2qlMYAKow/+PQRdBKfyIsUW2
f4m4X//l87XL6BSrUhInWYA7tPW1txrT6DAW7vxugS/bYlTUyigLV8akseBOHuMMHhsgw7GPK1d0
1MxDTNWeLM1VVEa1Wmjn7h7CqlAoLB0JIevQZE19I8nhPhbNIxtQRxz/ynizeMNWuKj3S90d6Ph1
5hTsFJbNPOewmEjoSwEu/ofiYhL97VJdo4nRdVt3VgdPrXC/dTxmdmw7sckTip/BrNVUYIWl3ZLI
V78Z/NTNzgScLFAeg8kv9HIqYvYFuMSf45zKHXr7Gt2InkGSyVgbenflQ/TAHey2+alQG7XwrKkp
Th+WpiEGJxI1uni0ik1BdcYjRM9TWjA3B0pkfSg9wO9gPJCk0YrVatHS57A5q0aaBYuEzrK9IN5p
1Gj1u5mgMChyJ5rjJ9Dyf3A+3i+uX+mybEDZgaSNInUwxa9OyMq3+2P1CS/ZceHUOkPH3MeAP9wQ
PmrPigv9DEznNnYg+4R6x3SX2itfkFGw0GDC+jYSjNIPU7s1wJx2rjjUfONPa11gMVfAivk5MQYz
UVjlcrk3+iEoaYQpRGNU9tsEmHDIlJJo52AZGH9ASshUO4PmWnJ3Xp97QCNkO7NcCLHVFUlr+mzS
eYK8M0rM4e+iHK9OZ1w0Zp3Tk+gryIzK56JEeaM8q3luAdFdcyGALnxOzDdR/jDv9s7SowDvADl/
KgCir1/eeQ/0onAzSj7yuLwHjFS2XFdDA2JocuYGZ+TDN+FyxxqVgcsTBspzJKOhhbMalN6yCkDX
B41VQ8GXDqqAwwMABgiVtvu8KS+yUzuUihEAqxH8SoNGiCtsGwB4yDBKQV31A1EodaZw6ZWcOjuK
/ukalj9B6VI7QJhvSPOFmIONKCLCSPyo9LL3nlqikqXRH+sPywDGi1ByPqBNXit7hnUiIVlNcu47
NXCbhipb+xgYrfO4a6C/97NL54VKspEmrewYEsrKvjsb9uxOwyfdOLZFvMbgt9FNFhy80KStnUt6
7vLVY+WcJvLpn56wb6RJ8+SNCN27cpAxV+LzGlOJ2/iF2n1RqFlkzS/Xrsm7V/g6Wi2PkQH7BBVR
SRnD0+k3uQcSYvxuGO3qhRINVQ6OSZHUD8K+mXTqwACuluXv+HRbW0O416TmLqoR29mkTKCNnHV2
ngE7QOZJjk4khpuprf5KC7jNRP3ePch7vvWFtxrzCV46huz+KAxtb8cGiRg8Vqyd2PoWghUrc2kt
CVM8tqOoCOEtnp8911J4ZT4ra49ZWj2QXa8JIh1aSXdXf54RNbwehC3LSiAvtRRS5lulr83DGwqI
04VZLE7XNY4ThVNAEhUVO5IeHh96PZAWtiFgjBJgR0KYvCDCnFLdgnPhcr6Xz+sCo/eo3XmUp07N
1zNQHMbcxEIAKIFMlqiYmq8rW+WOSqtKoL/Neewz8sRNdsbhXOjEfu0LcGMRXXUMpyEmqONdWRFo
4zP5NJwwqKyUnO8ER79hWTgl2vR5/6CiuYPstDrK/9PdcdTgvCfZIjez6wau3VnDzlwj/B/GNJyr
3W+g+Dxh5vsejDmlDYMNECDSFF+W0fXhC00xw3r8RwBig7UB9V74SYhJJUulyflCuAm+QUZSEbgD
FeXLlWDWWtRlpR6DUWuTVHkoOtZVgFvKaegG5B4/IsRMYKwZ+Qu9jyrTq8V76fCU1E5XjRKZ1pvS
aK9D6BE2f+uVQveIGLSYijwYynSfOUjWzKHlSQn2tUFBEoz+xzz92Np9IBktNXToaDEP2AiHsXSk
BSZOKhsF3DIwK8N88V/qH9NqPtwuRaqJaAxmi+htElPoLlKesZ+b0V3i1wMOwKySnZnP/Y7/Xq2q
zK5lbt0Hb+DCrwQxoBPwYy8Vc12Dh96auGb+6mlGU8nQEBR99OqLsjcwNImqpqXHToNKq4kwJqWJ
PqR1TqczZnki5pG7IvPQfF7Ffnfmx8wGPDzdNEkCk0Oot1BHNI6KG/FEX3gJ8M3sdbTww+MiwBGs
a7TjyURDt5mBb+ssvK6Fr1gpFuBCBAdrF2K7+zVsT8yo533G4Bxe1pSOQdufz/C4UXtGQ6+X1u4k
uV6/owRAAYxnkML/kgrXbg7tlOSfktrDkOScs7+kzz+gH/mmx+OPlJjlcbcHwE+r1NDnpP0QHHPo
sDMXncMiVArwamw0UZmvd3RIHg76qkMkVvnmaQTwJJsiOMSIG3kBRWBxuzLJi9ROtwKl3b39b6wl
NAm0r7cE6MKFC93ZFOB1+xpgv+UqJqfkXwA7O5Kaxhbwzl9velmOxirwpHO2OTbUwkT1SVtqiYAv
ZBvZb49ETbKrgkOY7RDMAztl3yDVxzl08dojkuMsDRJDEtRUoQo5GAlSm1QazKc/TE2ovkPoGRU0
jr++gssnaOKWw7LGPZr1570sVuz2ZnUngoE2jQATDuIEIG+VnovHQq/JgXI9QIHYgk/q29X8Kjuu
CquuzcxG8Z2ISSmJU2MOZThTTSDf8FCaCd8llcaqklQSU3he+sfzch9b5RhAqMkSu5ssDWQ8qFDF
qzCa9RmvzvP1dgr2GfkZOgsf8221GqC9S5h++HnA8Vn+/3CT9/J/3g0yVfZqjN7F9vGnyc4kSneu
0THYmIaR+SF2Y2rOhWdgE20esH+B2LQTGz+D6QF3pcicRGwUsJjsCyXOtSwYD+ZFTIdLDVSGoR6d
xtUCtTPCBB2WwCr+bt23MR0JdHkYZSUMRlC1sOg34Ey10RA1mIU6s0GH4BIHedq6xT/HZc3Vwsnj
NFcdloFSNQv41HAhW7NaM2f7aKyUGw/SLba2A2Oi+7ka2jAUmhAgZj/+tOgzea+J5/62GQCZaXEw
wIjQ9lCHJ9rrtdZGjYx1JBmL/Uym+uEQFjVOz34E4QuSigNZNNnf+3J26kVAD/QtxWww9UYRfX3o
F1LvUYeBG0u/lz9yvjK4qY9HR/bYnLEhD7AZRmlQ0B6gHYGc6rssvTNIkMRYfnrKT8vfpmb6PHyB
Pcs3W1C4RswtRAN2hgRZO5F32FdwB6NIwNAmvuqEfK6Xhm8ZCq70ovp4EgxHyIqlkMW2EuK3TdRh
DOg+J8vHU3vRNdeJOf6pQWOzkHM5DEMjGvbVwvcQJP209yVKUQmHPuiWBY9asIQ8+o0lKB37C61h
H/XYgkWsrtoDEJIH0QowWtwYbfzG9viPVcp+fJWgZBbuOiFLydv3rlCh92GPgObyeIBs9fOWg3p/
Fc8QS+7XM9XHgvUkba+9Za9etzJCnnxuNUTn72VX1ztrYFe8s79X5nJF49jcz0yRflWjo/iRidXt
GpHKpFY1LE2WrdMPvc57zsoT9k7zYT7yfuFKcnDdDp7f3y1Bp17pveSc3bwEz4CDhyAgutH2OP26
8f5tid47+wO8HgFnoc2y8FwJsdlxVlr+mZA0M3A2FBh++fxsyvzpkOvgj/cW1w12vsZ/ZnZXYy/0
dXcaIGg/fgZrovzQ9KlpCb2PNUtvJyaNojaTam/yBTh2nDR4rbBI+24YojiRX7vzAvyfbTz/F23o
oe6HAHG/AS0YbpPMngN6JsWi+WQDGSTEQDmpeQlBcFAOq3LNEnGhqrFuL88nKkUynsCyEAMvkFjH
ozZfseHiG71SMkL6Hw0flbNrenjZL9L+gPL8FnkA1MDIZAj7NepCtS/g4cLJ12H3/FadaV66bRuV
oa0Klky6UIBX1XorAylFIa89bCkJInxTkHiiznHEt60qTuCW1kj+bRda2p+njoOqwKn+0hysCALD
aNdvUn0MVrwKdZjNukxRWcsPPPLtgaHVbvJtYJORz+XvZ0HRQwtaXaQ9t08DXlrWsAXCWLvwvZNW
KmYhOoMyNvInyldAf+i99B/8pyBWsRx/NtpM+GZxgjVBt0qi8lAyqzJJhGITxknz5/V0/AImY8zG
WgEGwktUfXcmlzGHkjXQDakyn3rYot0sIreEoxe2MxfRYvIzsBiY692mMkLljuDLz45OuFmfPj9w
HxNWK4h1QByRk/XbFX6S/5+7EcczfKBWT/XmpPuJ/uWit9oVfnePvdOAtAOsG6/+NP/JTIzX7zW2
m3pYkz+PxjZA+JuDsgq2JFyY+/br6md/bg4VdNeXRIbtZGtUKPZFcYo9TdVbbT0ql/YvKWts64Qd
al7RT7MvlFdyAf5lRcfgB65nO5oUYdlP35SSoUH61cZUAm42QnbOPomQyPWsYcdTp6herY5mnTEt
ud1+54CNbpxskaSZp0GvT7JMblnpAZtuJvqEx41AF4w7PxTEqXkd4GCqhQegp3wxxIR4Ri6pGl80
NoUx0O1XaQw2FQcHay8o5uXKTaQGGCHxym0DY5T6RlgMjnRT4wTrTsFVfUIystzAo532xEjZIM2P
laVhJVa+09Jfrdx+s0KAE88bPOCyixt3dnY+woYKEMZgQj59DqLxnW/SQj93iepO9SKr71DqZ1CK
+SJAUymdkFAXaXVI+bNVOj1y85G4WZEy1NEibaOebG3tkqBIctacv7UJFtyqTaATZakK+++Vic+C
yelkJqgJGwp2Rhkuh7BAv1ja3fhZauG0oWk6XjZjmYJWwRddKQN8JIOMW34SpP8gvCt6NvvG+2mj
/wCajiuBymPFRA2NXO/Z5BQQl3J5Jr6H5xEwlvCi/szAYhtl2XG2qyZ0eljyIZHIKYr2sh8gcLNJ
JYc7GJ9bVMZEps0QB94HFXZ3mKXcFnTT0dyKmTB/qSYr+/OAvKbNhtvtWbuWy6AZZn4mDTGauhbl
sssnTSV5k8VdyqPoA/r+m/MC0X19O83TQNKq9LW/ZSnjvs5pbn3M1KJijdPDj6jLgNtHesbKZbmO
0dciYkQ/XQme/Bvbw8DbqN2AB+2IptRQQj4doF886zDEc8EjbHEEwBsgt2oy9OrCiJTYgSLP24HS
cusU9Vh19/o5527XzI8g9UYVFnCbu+sTLTbhyW51nAn/DFM3+4uMsP7Z7KFHriDtXuJTBC2P7kDh
nhRd1XONJGH5iEOTZfcXZlfdtw0S2L1RdXbDbNdHsqRRNXYF/biz0w67maewga0E90yhr8Icj744
Kp2/wrv6WkGsY6LO+nL6mZgzFBx8qTltWpaXfMS5OfYHZwYukt6gYMv5IiCsMAYmMzFwv8yy29Zx
8yR0z0GTM0eDz4WFuSyUNwA+UE7A3iuEWrsDrEBFxZpT16WE7tHA49ssv/y8nSRbi3QDDBX8d5vH
Qq4eGGXKQtya+bXMHR5fmeSUhu0Sy7Vk0EDReC3zhgNwXW6oPxHcwysImuaW4Xz5cST5b/DQW4+N
qWIqjZSVthi+w3sJ3kKSNHu9YAs9IsC8qLRSpdf6D6wWHJy60Ir90AuCRsarwbOOYwlMNFY09G4B
k+c9BvxDOI9fMG2C9UYlGmSK8IeZ2rrvX8n63e90MgpxveMhOF7AqPnSW8diNUJi1ty4/Me0gd/r
UWLMxhx3roiY4Ih/dXX/ZcFTgm9m4/YoLwbgITxed2yj5VqlM+BiIrJ4I/INExpErMXWQpZdJWyQ
kwFkRwwYOvAkscubVJZCFXM6BBykzfV4/sJiIkHlvHwFOwkrb7QY3Dbu7ybVf07Ksl5Dc6TryRW9
K72z6jtZ+dF2sYaZvGdsiPtUbltyfpn8kLoQo+bmr2e8xaT7ceoCJLma43rbmJmsQuD/DlwMXM9K
tXuzM/Cu5L5TMbpjnquhXbVUxxeYmyzbY+YCF14TdliNHjFXeo0ZSkUAWNoRhsORsSK8S0ZHFBCL
9GIyAwzABcOOAT8OWwNHtb1GCpL/IhZxFxx5Y+Qh1/Wvr2M6hVbIrfiMZIytvxM2U7Q+plMfTCMk
V6fuc5TLwH1rjgy7LQXhuv9ijcP4MJpP08/MpIodAGRaaM8sdFLYm3XYjUVjvMxrwKH5IxIgyhbf
b62l48FfSBPRjEH6w08Va6G9sHCyGUJZLg4KcDGu5vKOVP8YKumyS+DNFoAI3XgYxV6+pF+kvuhh
QAn/MDv3xpzJHQVnYYvrUnYT6hvzR54a/mSoZvvVqCuDhSyT/yRwso/atVP4V+jCKdabG7tEdDQH
e6c8t9kyq6wc6IxYOZqbe+AJV6rcVElAUdOlPMwfzBwj5RKLDKWldO+ENf0yiHOD/sJwCU5W9Cag
x0Qtw61g0h0uIT5W4MtANwJVFZh5ItocSYoRVI1XcMEGovCJoGwM67qFGzyspkmwwm9b242b3yIx
nhJSm2FWH+G+38WJMN8XF92X0QNQ3FJqZqpEqrVtM5YxLYN6PP7Vp0mAAmwXtPrLJdLjUC2V79xh
pIWGEknpuSUvVtIoCdVydwnSEcO8JYru8dCVXthshGUlibti4xdj5FlBKwv5KASK1GqPlqfYLrwX
FI1xnAaZvtKOb9ph1ZdizV9hOyZkItb8uc6CNTmdrmV9v8JO5eOrKi0bIB0e0m+nkW0PmD20fTA8
Z5xyGHUZj1uoBBSil4klIbFb9Y0EyvkzXOiOFx4WTrDeIahKyqpIv4h1EDfF7Bo7BHKH8xTmXklA
U9A1+zH2g6ikXpnESxRE+p1HtygvxMtf26uc4+1RlAuvukoVy39D8TVr2f4Q2POoeTqG5E7ntMI2
cfEBq/HCtko5Lt2FqQaRNbhgPk/CtRnXm49TQyY4JCabsWwaLSMG3mrWlj2DhYww2RSVg4nxX6rx
zrTwNhTS/6pe4IqFP103+hoZhl0S+A7pj/oYSi2kWJouPzzKKV1u8CDMV/27J25ywSwXvT6FAEUE
UJbLuc0jyQmcpnM5kaMhSBiwYmX2qnkkia7oC8uv3DcPl4iSGiTPACmXJ5Pw7xukQOiJx5jegrGt
sDpUbHUDieNak2vcl5sxcdILYRzw7IQtKMoItHq5jJ/OlZdrf15c2l2PaRjsNV0UoXs7w63Dgp7c
A3tk+jDLg1Aq9Le5u/CrQtARP5nY/SpFyOyOsHQTC7mPDbLQEsjQooTinJ0Fw24HruCRAEjY6pIa
GWMsisJChEfyAs8XjbV+DFrBOsJpA8NUl07FxRafjzvz3NLNbhUt5A3irgwxp3GCdE5rn5WdYgpe
Tq4qMITWf3yEBXzb44w20v0ZOiLg1WmkIlquFzoJbuOFaMErHVwcviXWpgGweFDtn+FNn6z55lVE
QLYh/mSpIJsSqDUX1syFBhAIRknX3i3eIx921WYtE/hGK3WXZIQLkMIvDsmk1KxWRIT5oSw4O4pA
oJRP9yDV7kqBTbQA518nQF3aD40IdyD9YRiXVR2rY19G8a9H+8TYyh+e3ILHGiIzy2AZefyQIYIN
OblF1I8f+BGm5nyONKBk+2i75Oq9NwhsheUqfCI9E6R1PqO7GDJaSC89casf3u39yoy/X/bMwTvD
WvM+uYQRBuGXuvo6bWi49tizavriqOXf/JxgJA+iEyjIAmOgnio5NK7VJX5FfYIpWWEMTKT79QGu
IvVfKV5pbSxtwerh1F4lIpxK6nyDcqlDNjZgCJ1eoi0GqY8RdPhpdRDtdY4VLneWfm3y5tIFxYLG
WuUP+teBKLbkz7qjWGI204CKnYI2ECBl1AA4NDJj+n1VEMlML0AQrv7qC1/km4JhvR//so7TavpC
1B1TJK2XVUMqQd3ivo1SeXZtUi8p85+6KQhOIR8qjPzOow7wa+gipDFfcJdKOUqs0FerQ87Wreps
38zt6Kx05OVcsbZ8pX/hYhg19bivyQh42pSPsfSw7qpRdFpKbWz86RejkLdJ4eeguG+KjBDVW9C1
xOWBaX3OxR+0ZdDfLH8bFmGsdb6Tfz/rJm3Wsf3+jFUac2PPjrYqs9UOOu1UweX3bJJ3RTqV5vZV
PmM1zf3lIQhjTKDl+6tAa5zdOiwbABBaoYR9BTkyqbkSj0y4b2TfS2/96cYAQumkqDIWkKFxEHld
/a3rpcgeIx+bekEEKmqy4MxVW+YJqf0orYaeCsKpHfmlVPDv+M1aiGkkhjYLjjiXv7oU8rQLazap
XUHWqu84y92VKHAWYFGBarSrbUcxXe0mukeHlxqAmT3E2CLT+4opjQEsrflauUR47QqGd2HpyPpc
q/L7uDXoYD66ArANkTAJyNka5+E2jXPMs4A4WVh0abwju95enpiZI6olc9w4OugM8R3HU0D0/NP0
Bbe02BHqbe3tQS2FOKv22WKUvoqV8YlVKXELUFL6T5BFUGkWhADjzA8DvpaMlntz/ml7KC4hAorB
98IUZswtZJJEyM4RY5SXXSx8arhJf7ODKI/vy0+Mo/5lfzPCFnY4uWTC/tEtgJXcGdXkG+UKls0r
1Ik3WFtFVrKs4O+63WGKgIBvQtgJLQLALkO7ma2uhuB8N6YV7lCr2e1N4l1y0aAlibP/8WCtht2Q
sdZRV1Eu2/6XX5HUZ+TyX271cGcrnOYWF8h9L6hK5Sx+GJCdHXINtFlHAgDVVLLw/CZIRjUmh7P5
tCE/bzaRWWByxLAAdO5/oKM7dVPfDD6Nzt9Cm6eNJzdRYGE4aFB1BRavA+ePGT7RUnZ86wS189vh
CaIunyTcLzFY8ZVJcXDKFi4LI+DmX+kyhDFhkoxEHnBRCpO79qBAvQ9y+ePM8byo81wbj28KH2wU
nHFJRSsxAr8fHAXOQ3vrQL9GkAI1rrItxuN5OUVZa6MB40fQOECiOr9juKyrycoh/HbrgBoMBoe6
EWT+cWYinkamWss8Uavx4QeqmE+j9dV84GyxvEZKS24IZ+IBv/yjotcoti4Q0KMr3IMXYD4UCm8E
FZesVz/Vc/cUdVdn9BhkENFj5CHQA+cQaoqOicEmGFi0f40E1c6M3xZjSkWlLjh1XG/7Hb7i1XH8
12xnZbTTx7wquSlAmEq6LQH2+aE2HMrmw4OcrV4vAsJ+HNGZTmPggahkkqFtv1Y0qJEiJLJH0IMo
2VgZXLKUh1UHYa23zTMb3VlUrozOGuy6cE/tvxbS3aHIV0f+eB7RRQrPxYComkfEpO5ruu9cqO9Z
0ja1COOGQDv/6o4EfCps4wC4v1wDh/nqsoMnMNb4exj3X0bIEa1M8rHzzA98POx8QC+SkkTdhLYw
4ZcoqwfjD2ZulY1CwPiuHUwNz/aZJQ1OKgoBuZh1W/1GMLnVO4S1ouP53edxT1rQJU+zFYUeDbgy
VRipqVKAaX4J1fPmzrtBSJ/GnVPFEzswGrUiozkR7cwGc/tkNzMrToJe0JJdy7FvelgW3pZMIJKy
jNGd0UQ1EpEO2TEgPrQsqIt/ZcHaFxKlndkB6OE9VycWOGY/i/mpSXVewTZqFx3wea+54wKF4/4u
M4NDDc9voxyh/Bts3/Y92YxNsHp89uCZxpaVNbx6AIiLNwjcm+rEpVmJr6iTAtkDRyY01g95FKiI
7f+33c6zAi60G9531aIx6DmulY8Lfbvsm+0KbfV5O7uCnGSsoEFEcTFhzpXnZnkEMCGSaLZIF6G5
lMWENb54pgfIO3nho1w7lbsm200m7+f59+69UlHBsj4DXeDrTJd3rii1r3Y0+AIjsHh8O7o3f/sj
d1EiJ5tSOmrtK+b+MUSFnodtMcpHXJbwWBnrXIdcWU7mFlGXYHDboDEcMaEhXIMGpC1t6fnvvpuJ
amznCbNmg8+ZUVPkrhmbqB3HYNEbOUDwpP5EhpLIe+PMZxyvRSTaQpzHn/zSaGZU1a6v/SfgQEhO
SdpfU0T6szzBo9490XWfZco2j6+78fk9ezqNQTyoZ2kjiBYxLpmwpUHbTLyRuykqvAcaEyolcutF
KXDg/+QarwiSGtu4SQyRw9NnI/KknHpM5TD8i1KJHCVFNjPkYOXQ+JEeH1d5EV5GGrCDXR5+R/tr
TRa7kMT0aSQyI+3JeUASkE4niToHd3Bs2xWZACC/s/q10SU3yhZ/AEIiHzH+MGMoNE16dcmt18N0
4xYVjQFoQmjtkF7SL15j9A0717J9jFIHTEjkLKHztmiYLXjUgS3kQL8zVlQduQt+hOjyONc3Kcqc
Haz+2kVMhHHO5XOFvCouXlXfy3s661cS1A9wqsbhbG2+46TNl7dZHA1+SoU7rysSCneP0MirG+Q/
M8uClIACdZudwVHEvotu9RqVct1XOUOAYCl1m/WNG2ncZYDhz2XIRF087DkzFx2Y213OgS72UKu+
y5946ENeGlsSG+XAuatIuVV1iJygdFAcL0P/sNr5fo1tntxQWxKTTf9tlmzgvmk7iAuIxqkV6UTQ
abR++KVdz1/EQmOBirSE1y1mhbIErSkuEGFiATL9y1myAiQpTP9T+0S94R0OYV+LZFg2SZ+sBqQZ
b9aEIdMvHi3E7XTwBWINxxpyVwlKyZqxnxvhmAFZvxu0J7Bj3ph/O+ElsButbj8f8B89zP5fw0XU
1WI48arn4//7Z0usB9bZrgUW0wZhIls6ylUBWz2qo7FuDdvFQ8UJcYAjPDms165r3dK7teDI2UWp
Z/08dUDByPQ18hse81vApDsbKk0EAFZEUFB/w9DXc1yc8LQBxJyRIi2DODIpJ4zCrjeMb68dJFYd
1A5LRiSNy9Q2qpQ5a+5ocUic0vdYYl9TIw1lCKhXBdtTYQl4bQHWmvPIc0ZNZM4Vckz8wrRgqD2r
FQqYWUMYP9NEBq2OcQ8GCjlFKkcFisuxWZ7pVyDWXUAqMr5flkaid/AtPXA1V1qvMYambvDoz6Fp
g4A9I5aIvwBnqyj7WANAA1NfWw6RXy3sBmDwrhrZMwCm4wHZdCiqSx31xAHSwiYebLS62gOGhhhn
0q2DWrbnZIoJcl7PMI6X+LDWT7ywXThD814atKrULsS9rrDLhZrdbJ0sVp0oNMfAnyrhmfMW+VQY
SiERH2r/hnRO2l3N7dqVJxRhVd9RP2zXGR7mldzVhLA52MK9HI88j+rEOKXhiiyFvP4RNPAn/FEh
a+BsNwE7qPX8tY2R95wF3JnPO62DofQX6GOTZFC7spHHsWR/5NfsmOZ+121FtmoKoaVciwHsFG0m
jHsbr9/sxwzbMdnuv7UcE3MRx8RGfGDBmLD3RmPhaslkDxe1+tC/bVTVkpZzpPLQi8xsKMLNRBzB
DzB/WZUay5utJsNF+OApbZK+EJQfoBh29qZtDxe0hUWwo9FIZ4gLXEm4ZckCsUTKx713kgWw3Hhk
Acp33TEmulycLwqPz2OLCv7+ekz7cd+tYLgssNNOr3pTooSa4bADt8hpckcmDG8y0sHrcra7v2je
yeeGIGzcVFCZxtnn7yEhaWG/NNPf/xD/rdco/+SyovKOnGXq+2sWNyMhreyaja1rO8FER8JSC+GW
ann1iIJQk6VOFui5kdSWnRBl6o5jr6pJJ4QqvbXYAbqBxuKS9RVXazGxWBQhJ5YnriNf0KcWutI1
K34de8M+0gzgHlwPdJwtCNsBJB1ageP85OIq+9VWjVU3TocEkSMR3x7zAutTpBOjXwUXO9lLpio+
FT9rbSaIt/GRFOIus5UaQPtF8JvdrlCMdbwf02d8gL10FwLYmNdNfeuTSFjvUuf7KM6Ahzux9QmP
D1QFay4h3wx9N/25PK1fWXvQDCs3gALVL6kRBZO5AoR2WaQI9Rw5Jwc9vVU9qb/Jkh43E/aOpKdQ
3H6QuJ+NVuBIutkOQLJksndXWjs+JgJjVXgvjuuJftNjHoTeiah53D+amOMgpMX3wOvJG8aoDVbH
k+p78AUQ2rfDG/uAH+W/pOJZJjQy+X2JEPLyUztMcIXhronS9caXaultQAALyHyHAlRMzBMHO3jp
z/wjSUTI/KnO1OaDC4xSV1pbNbzU6FQcZxjv4+UAiHfqU//NJNQnlABW/48mYvflF1c1dSbvCC8J
f8z4qOAXiR4vv2H1TxSeEjf8VWaMsFv8ZOgN2MhN/iOtOhR+hvQrSNcY0vcl8wTNdPvVZ7y97pdL
LOQpC6c0gShtwJEPgmYSy9dgvF8vLhBrXsQXC703WQ4NPX7PF3xVx4i1/Y3PMhUrNagfEA/Y4aPG
11sw9nW9CrrLU7hJDDMM7hm4UzbdbkGg3QXfO0a0RyXMXJda6SevQ4GFqAFqNsLp+0g3Ndd7G3/V
8QFeQXrGuVYYwL2AgEcaKf5RfjfSOcCM6PN3lg+gg53kg70cpysiKzsulzJG1kT8hWztlxlG5Mwi
2g1v7dbA/AKco3eFbsr8CnarnxhkhhQTaRpczXDUbpUMIz7kcUfdsgksOXoUkW9/TJe9by0v7iz8
UD/XRtUacksWBX8aB8se+KuofLCOrlPaOsMiwFqefTdasjpnTx3TGfJ0HEqoMiu4sFvOj3YeEpe8
mQ0QYhuvnGb6aPdnW/rbS2JbRKcpWDOkMXNZSUJe8+nZCM2tG4Cjj/aPtLN1bj7KoaBkz7KrnU40
K2arZ8I6GTLnP03HBP75pVCCT5il8lql8Ai+6TAy9IfNV0ivHZMtVYmHVO6cRa5SiqGw8ZwPywUz
GeqjCt4kpxINPZsvMvOp+yXHMmMoSe1UpCJHQVcFYRlya2/NlVJWqUCsrGOOhwmJ5mMNJe0sdTgu
HTEHeelnhfWljOX57YscZC1jiGWLSxkBw8i+1CwKXljKk/drIZU2w8bEd9XoKKWqjansD4Z+gGfL
IE4vwQMo/dAvpx7rvX5xwEOkdFV1irLSvvRS7wePXuFCp79aTUXxqsoneGXXzY69Q9Z2XCbIjH2e
ajlfMbcrsA6zWliDb9ZFPklPR0LvYuprx09z3PPutfRRUa1sR093Vx4hMUpTKWufdXppgdCIJsgW
yIvKmPvAacfzH75dVM4la2phH2xxZzVT06Qglywr8K6/AKcG3YonWL0i4PLVqyvwQub5Zz0KOFDC
WgkelDNjO10IqaCY6wR52iokw13VYW6ELZi5ODevJV62Wx8ItExpNVOwoAsuT0WbBC3VqWZd2DAU
TnqmmoukFBFmjGgsRYEnhl5pEWy56nO7+7FujEt3TatUqpfjgWBaZJnUnEHjywuWtdO01DNahyU6
fDT6vzmrtvxu9gMk/FuqfpxQCzHJUVMJS06oR0/fYNZ0uxWKRaY2+evXhFL06sg1yY9pi+ZeHt7K
x6bEX9lsUP2rgLpYuYB1t6A77EED2IBH2BtM5Ac9LqIWlYEtbNE2WNb7udyLq/Q7M9YZDR7pMVbi
b4cL21gu5XXSrpM2C6VHyQejw3FC9SeXZu1J4u2zML6byWfrqEAJUM6BmCy5+fTCcavvsOy8r/Nm
+uTRenFL2HoXQQzV4qeXaeCpMNQ8KiJ/dWcLPH1w3/MSQRiGylqL6YrPSz13E22u/rMd9MHxHXoX
tBgN9Hx9K8/heeK79z7cIqRxeait/TMW7G/OfepY/IHrR70k/0VgUhl7S5Jyia0urEDgJwzt4fWS
OUCKaSsV3/89Xk9JOaKE+mT8WBWHUdtl0MgfQ5iPxSGogBqqI2I5U4tDBo61r8yFgygITRX0BrC2
v+u6dPgm1kl0cGV/57t7U5+ieVofrBHaWH/Rwrpot+WxSF4Eck77lMgdJt71wGl69+sNZ3DeiLty
sQs5uDkgbYMGGLiQlfBToNRcniAq/bvx4MsAEGHNJZ7eKaRGJsr/8Ta/LTnI3q3HTWTyS9OIqcKZ
Ir2ZYmwWKUSiZiBexXKXYbtdon5gcBG8ErH3Ovql4U0y9G9FyJa5LiR90KnJNiPR+au8eRVxA95U
04CLOhu1TcC7hHCxuQyRe2Mxl4z6UDkG657BDEGxhZosdOMvtxKrv2oAuUjKHg7ZE7w0eQeHHuLX
I+4LhRsS6pilvi/vetMx6qmmkXlHo494P58b4el2CW2jLM+Ejie3KfhS6ZPmBB6xFYMUJHjivVhu
2DAkP7s0YI0mxqX0mO83c+iXLGsbcPafvTW/go9GGx9SJ8uspMAb4TMLkMfyQ+c4klGE3Npztc5V
mlBwiDDMIXRdyqqOInGJCuAqhxCRvRW5tNQ+GwN1v+3rJbkOgz4kD7dYmv3+WauWNqk46nn57ukB
eyezmyraXaQ929uysOrsceRXKYqF6ujcthZXN9vW1WGJM5CoLbLlBM7pWOJsmEREjtuiCHnw+xdO
mi6jDdKV70w5Tuohl2XmiFdvmQRTw4Rw9zfbu9xnSSSEpl7unMnA0Bov4IfYs+4S0OLSsWsbL+2S
JrXsu5UotqCq+FaUtkLS+otBrXwjsz0GSA7WFdmtDe/NdGXJGF6xkMQ+OqQDqbV/9r8OXic5Ub7e
bm2uO3c0PszB7mMc8Mkaqi+5RrtTu2ve56koct5ZDUIa0gR8BAQ2H6aby1OI1RGnnLYMz/E1et+j
KI8pDkfpL7TPLnqddCvDR2VmfFDfwisnlQHC9t1q1tL7BLK+1KzMwaEVFRrdpOb+xXQuvtsqQowd
UYu52UByzJa0BwbbmkGZaNe/qC2Mo7AdaTE9dTle3+FWvXMnM45dA1Ve6pARluD9giLNXI1Ltmms
X6SwXCN8JWa5TwXUILFDbuksP8v5F/ObpMnBQ6LdUTk/wH96tafEF4NeNSGB+KCO37YhGj6bDISJ
giGukaPPbna6OiDApWqR5SUCh7KyOskzBEz1B1mOLMX60a0XM9Fn7bAxIhSXx3oOu7cIYE7cUmnM
60jPr5FbKxwQm9SaO7SftZN32m3osF0Lt6W1Yp4uGLXIwM3eJamugiIJ9OtOywzcgeMU2Cfv8tmH
0+WL403F7PYFLwn8VJCxx2G1xUfKUDk7gYs7ITZGLpoIcflDPUkyYAL0peT8WezfRaeVqRz8FozD
z+ZskFK9zLL2XaKDCYaCOoyybDNFGvYm5vP+GgJwbZJpALJ07hhbFz1WiTf6RdsRTUyaMNsOKY7G
WED4gWz5oHTlcPIVAN08aR4O3dQctSTHY5c8mI2DVjUtSaASDtKXLPXy8UauWiRdiDnWlrW6isWj
UguG9XzkxgelCX4dU6kdYDQBytaFcfucO40+FUk7Tpz3Mr5fXYEyE3RqfusgKkBz7W/ArEkd4yix
Tg8BIEdfg08LqEj2u6AaJpl5mOFqqhANaruxnJM3R2eWaHtgg9/axFy7+k7NEYNigv7J62Y8aHPt
I5VoWbmcStT8ZAfEnhY8DtBWGxmf0raVi8I75HrgPPDAh0+jUihK843FAD3ndI8pzPDHeOG8xIjL
nOY3Gmq+bndJHA7HuNgYvvRM46nkYLrIZExIIqbhHw5BofFZTrpyMv9iLBCn8XzF02PB4lkCwoRV
oI8oQsVYADp2dGfVs26Dutd5Ns8ZZ8mJybZfxGIzuHYWjyJ6zEYWg8ZzMVsGSqWmnUwZjmuxNHIW
AkIjRV3MlioWEq3fvjSceyfCHF8j+C21/Th/6q2Etfpbiislq3Qalu4j9JCMj3oiyj2s3vn40gDa
Zz64AAo+Oiw8h067xJ1ULiG4orqCQrg4U311r7ZLuxg5azAe1mQA33nk4E0a5zs/t2vYNpTCOYPJ
3o5wJoh6uS6hcBIUH03gKtGc1w4mJE/AD417OtcXCNUj4iFPSK0/H/CPO0kvp0cBL3LhiHoAihxW
rOoU4osoZtxvs6ym1xMkkkxIe/ebj9QTYToWl3HKMTlbZ7P2uIdtBv9fYxyLRoWfo6aPnO395yQY
otkTIHJZC/l2xijI9fFUPp6QRnpamzmkefm7apWpGgDOI/s4/9ByFLkiv6l5LPCWNa+5fRMntBGU
19Tq0cAYFp7Qk2n7jnrennFJyp98VfJmZ4IAtpr9Hz91/3b9PXnQcwnn6LNnG0QBzCNV/yscth0K
0B3kU8qcvu6OHf1vaAg72gbULfhoRX2sj+PYRDnK8tEHowxQsfGTeh8fpcgVQZiufsjG8DrDmiou
DfOndQa5R4mhSoe3GuF+A5uAo9ToYnyJb3koi93IElkha00M7OS6VotaYgXyHUrWmH7qhE7MmsGN
3uv1Q5nHZyzDZGsYX5aH0z5O5zH6t+c4R6APFoRoN76jaUOCR+LzlrG3nKq4UJe1aZWPTaoPjd4k
DAo4ivrcyo/nyvrqrGakmrtL8h1Qk5VPNsv6ioKg3iqpA7k4b2plAd85VOW6L9B3K2m284vgRnZn
TKUabfVZ+LhPPOfkxlnVM7cfUgXJgXVNkrQ+hf6lv2oL1VkGoJvWdOdxSNM9c4rqJbf0YBMd0ZkL
sES1li8nPwtKrqWfFVegxUKRG8HSm1Fe5FEAisVV/AeuR+ahJGEpUCJLJMS2cvxIJ0RT0U60NUj/
tUjYIfJeQ1TroJX849WH4dG981irAdSmOcOmDCFRWxmQyAxF4pCvNewGzmoBApl34XubXaVTX3uL
j5kOdgKXWdg80i+r5z4rldhl6UbVoUhgMYmey6Oiibp4fT41a1KlY0xdSm05vhSjGimuq7Q39Kig
ayD3JtWm8XngC8oRcQE7MBZOpCueZ3OedhQMvwfLYTWgq4U61A2woHQ5mIq4r73g9He0IHFx+OKG
H40BmR1T7cWoP5GxiHpbwUykFnCV65jSXqQk01C04N7cPshRNVeJ+RBq5nsHz9dvGzRM6DeI8Vjj
mBBE/ZPgFpJlhhpWt3oTRgA09ffAeuxpuOkJu3DKKDCiKL0bQxMvq+3xVlEiiSZQP6EAIg0AjUDQ
g5kw0+Ai6umay1QDo6csjWj6ewypFT7cR45VW/b9eLTlDJRVNwCC1zw69Svm0QMiLYpr+Ii4y6zt
foMxNn5n8r29OTe1FH0c37akwZS+xO8tL+amY0Vfi9gYtDIAMoCfrxOs0gbPSHJtXWXGTPxF8zYE
AT5QsBoNzM0U8j3aJfEeCw4GdsinzM53Scx50kORpmj3m/DpdvBdhb3rKBZ1c7Fr/dYz5kq+Mug7
ejBc1hXrg/QcEkE4IHEtutLWdo50M0CBWk8XKZPHIdAq/SZqW4MbB7gUVPAVeWteM3PiAMSKAE/s
8SPLIb/Q3TurB3Zrqlr5/wwQzkeZ1F/ayNhy9XSN1PZVSQaLPupFoivkrQAT1ilSCVAAMTvkHfoJ
S/pEpBWxSQAbNmgSm0+fcNIfdq5rGfL3XDXNovYDOjmsqDe427/CZsYeg5hePCG+GXUI+RzZwjzK
coV7S/GiV3Km6sd1iasWRXgj5LeRTSK1svbrS2SQr5t/+hgY+diH4dTeJwtvq2rh8i3HduANPsie
lL3fjl+a5YK7caWhcZD96SH1Z5y8AzxqTlWSw1+vZKyRSt1K4zqBqxdX1bxx0Hy6TwYig4usWJqp
5Gxg9wHFEAMPInH5F+mAeAdWGLz7nj7FtmttXWSR3IL8O9DHSPPDoYWvxbqoxbjEeFr7aGHot8GY
kJ5jFqxAdoWw+HrCVdi9wNxjvHxpePGObbKDD2xJeqhtH4WQ9ae6TBhXJrGcD6oPe6iqxePs4oBc
VfUFa0W2wAZ+6dEtN0vNIP+sJtiggJpsKLjzWRfNQZ4Q83JIYT3EzvlCZBoxWOe/ludjgm20nRO+
81DYNnl935s+QttWDGhu3iZHQT8AQWXnvZUvIjOZ9lENExjV5XGxWi43vPyb8YoTscD8VbSmJu92
XG+SjIw3Sv5oPou2rZxa2rsO8YjUrUe0vQXhNNKxLMILoJ7BD2H4iWdXemz3fjHjMA3+tebTq77w
0iWCMEv8K6oRwyD1aLimYnuckUtMOJcAmNuUfO0kZk2dWp5nB+sAH9leWGSWIbsS+P2VjLQgEJZs
pJSrS9pC2Lq1m6hCgbEKKKNXsN7qp2PKrjafhUOs3wN1RS04yHf7yyRe/5hFN9p19+uxLCgzLXoT
elPu19gW6VgJ5arL6nixEKMSP0qu+azEPqwLOD2WWsXA65JggGZNOT2s93rSJF3aQ4MBe+X3fUYz
7QEWHTUkompZdcby8xMVRxGh4Z8ezH34p8HUD3FRAbnn2k4A4YCsIGFYzN8uz9GVYHAZLLyAKWHe
ye2cH+eAkAR5+RFw2vX8qbvEMUIN3UUdykFH3q/I0LYyVTiamfDNulWZHLLRYwMGMLO0QsXf0K49
m3NopFL4fcpYXyndALjTC3bPZJdfsEqR/4SB6we9CbYR3byVftFFZ0kNpXjiqonxEz04hHzEfovO
+H0/UA7Rdho1Dx1cueGzfXAr9UP57Dq3mwKF1HrhtH5INfh1bk57+SJhuByO1YCrjY9gNdc+Elo2
WpJvJPncrIDjnqCuq4CvO/53Ju/BwX+jrD/uGNx5ipSTC032drxReGUZtYeokb35zAWAdYVozahR
aM+jqzfKSgb5YedcBcZdohWt9t7X7vTtDwqqeoeUS8He/E4oFhl7Xy88eScMu/ivtXUFElcHA03B
VUuLOYQ+V+KvpsX2UIKYC3V+Zo41H6YRgIjU8QZ64d5m0qlGxn2Ryc39LxnsRvrB5ChCQxrmvTDb
OAY/NeH5TV5towjbfDAM/1RATfjls/3JdfB7zVnFFZ56DJWdPs3wARLEzKYeXxerDCB/ZiQOQTX0
2RxZGP+aD8y6kKC+TZotpmddKjGePtSTQci3W7FGgKPSfgdgknh5LLYyZaBpTf6IDtHe3xtcVKyH
8wXWR2MY7x+02sO/NOLrMkAualJEXvdX1t3JsLNkO94jHj6wLmm1X5FtRbkR1x9WGqdGJ3HxnWfs
Wb56E5tWnwaA+DKC432160U5+zhkr1AtKWP45hcdOJ6lrph6gbNMwaZnrghrawhCeyeLlZkF5PVH
ZFP8cnitsH6yjjBpHTIPVRdaMoUaHLa2AOW4Xl/LARZsmzGf67yhVmQy9BrjgGRAzSWvnDvB2JzE
0nYl7SSkOHJ6q5TBogiA+fcfx+YfEfpaZWdamd5dHZJcqMGPuUOyPZn1DaOImQu7P6LzOGRB45vT
kiWo7bWNnljCQVruHw76YjOB3yflSNIKyfx+Fp6VCSUyxpvMfvMMv30oyPTl3nMmTXokGWgcBUDB
3AmP63d+k/ou/1hO41y5n9ixmYEhjJvx1KO8oPzooKvM425V71nwUJy0xPCldWQfDSa7caexUA3+
63WNXwintLTDoC5m0Ww6W91DCr6KnrMGqGC8lDwWMOtfNKCBN6WmTVdfw1PjQ/Tdv5MJ/bO5rtfU
3XqLOKjfW56X08hWuzNCwPUc9vbr7yqOXBAgbrCfFL5tZ5optCenlPeyBJYiB0jRM3EVh0n3cW3f
UOsGaBzcb3g/hpk0DuN1um5LvtL8H4k18AdbHF4wSakfHr6KyTuqxDMEIMYw67YNw2zqMhhLAddo
KRfNupjdGuWMPMtkQDH4C+UBk4IkgG9CzZ4IX6nz6qOTWECNiIh2sl5OJyqnJ86cYLS1Kj/zI16V
uA/lS4mZDiM2x6QESfqtKVPg7uI1orAHjbKxBcmwuNE81RNRfTkcqQQP+fey/ic8Zd65Qd7k4GqH
OnTBYVFhwNWmMgUjcfHP7aDaRLuG0dhD0MN9YZ9Kip3mJ3BixbR0y2sVsdZo27YSv3i9dqtZ1kss
bq6uxkWqeWLEbacH+XPb2fIxzosw+rrGahHiyLwDjAUUbmTwDALiALZI6UFzJpk1/dWus6agQY07
y7ResfG1UG8PQaaN4VLbvLB+atOpY1IKIWeEe6FWiFU/9zmTOhEgbxMGp4MZ7fNKZVRFSGFSq1mW
nljLts/W3WjAB4PDCLX1WC2BZSJG1AKPC7IRpi0KMnfWzW8MOwlpL46CiAIj2/WNGV72uaNBYmuJ
rs7ohRDggPUGQ/Mv6iyI37s8VQsDYqH8IXXUF+jgVAE7Q40Gh5iuL32zesBkE8S724q1xVwlsLJs
ceBaZ38pb9ptY/Xzdq95DUnLWgs3g1qocE6HcF2QOFslEjsrxfV2a6BYX+gPR3Hj595w9DugztdF
EVq2NlwxaMDpREakGnIaUsc9aP9CZOXg/ClQVY0LArQQvUyPQl74teMTNjU+tQrk21DqU8+HgHtQ
bVUfs3IbXH3ZRl33o76CRpaRsFzFzwgbBylEov2YZpYOUvglQaFdHyJu9aAnRAzlg6A4qxmGe/Gw
mOQH132CE+ST3xNPlRyzw+KAf3HsZk5BuK7F760qJnkDQYDaceKEW4xPhQ3jdT8wgQG3zIUs9Hpr
wnW8dCHehLDiBqsoiUzn0pcIre4/QTNdXNGPK81olyeLzwjcW94bIJHeQUARw/q+dg46sZeU7ilB
68FBT/Q4K5hpkMBLViPzafimdbTaU0x/gsRoQxts6stUMx3HiukNO4UHAcOV/gsK9k3py3y0By45
U9sKVo8vDyBWqAo91F4L8adKuIaSti2aO5ji9qlkfj1YIiemdT7MlcOy001tzVH8kAOGPalW1MMl
hoo8GwqaXUSwxKpLqqfjunz082D2gMonF0K9BA2TsxGAfumK7837/ChlFUnInaKmk9AxZaDeLHGO
zptSEmlE9+7BUjkUwdTKDgylsEiMrvMeHcBKfiRrHFFnDEknOfZzEJMOmUXsZ8i876aXy9VoA7/a
d/X8wmdeUcSJgV7tg2126HtwwzTklO7DOSiCNgYRPTZIwpsYgSWBsgWMBsHEeF4MvQhrVIWkZnm7
znaC/BHrbwSPnqLjaidrd7kbku2ClCp6VfRcgaZaTSYEenv3dQAC/TTNDcXgQulcsKOfHJ0/v9u3
PF0lNGFw9DQPQoTc8S529yM2AbmU2Qw07+0NUzekrf7v/ZoHke7zl9/i13kietAUnIY4Y4e/cs7o
0Utneov7HVDg+eDII2JHJd0c38YpgX1z8J+obIVV9Rk7tdm6yJisjqqXGdg4j0wCus3XS/iJrzWY
u/k2e+7mSbUSVz2UGVszFqwieM+hIwn41VfahnbxN1r6YUsDaC7brAL5qoUB1Oqyo4XFxz1/iTGz
e2XR46ElClUOUCaw+61NkCXzydE7dlzmFGgPxfPxz8Pns/vhtucAkghLwwOs3NLs4RLn3d1kd4F0
xavu/5bVebIXu2Nd5N/huU4fF2EPzCkyn1240LJLcw0+d9s7C7zIZXgZbAsv0Uvz0Jz4K8dg50qL
VnAagx8kQqlsupSYef/xgfIkJ0/epRuFo+thsH7pjzlcHCovuYr24izRKBp82cwxXIXmr2CmsEOI
6SoDyIVzqwC++gDG+XwGzD9Itwr/rL/R4xWcbZHtrFGwgal4+ULJDsQAL20VHj4D7TUXW1X8qiJ8
U/egn3QVIHYXXERE1kVwW7v8G2zr9FQNP5fhmxOWdtH5CJh62WsdZkyE+KfxlYPB7gEAG9LZZ2mb
LFNeYknDVHm4Zh267g9APR4r8JGBi5Myzigay4BeVRBjZPJXZkG4GAHSz2eSh/FRtV075D+dnFpF
3XyGE6ACE+EZ7AtO3NOOnGZOLngTUMZhAQg5wG2I742Ewc+Fw+mw648WWUlueUhpjzQk/2O9sGss
yim/6XYJOU3yAz3S9dbhruIzKiaYOTzv6wwM1fGW8BXiToXDtXkVEu2o83L9ubREOntxKhjNbT6m
qm4UQmvdyk6UfiWXq8aJAfxDaer+ZmA6OyeO4YMBe4fPqWfHAymJXae1sFFaowDRJ3kjpGpnfBrB
MHob75SxpIXuacyyJSz7NKaSfmCndK9RhqxQP3K5PdmwfKzQsNuxJknBGoNWhTA3pR15GPbyEeZ3
/DVQwwTAMxaEGFxslFiAuLWL1vfpkpTbySTn35Lnbv8eY2sS2u5JH7DE4NB6gQTO3uslD9dW9uBG
3jSbspsfk+/u0XjbjqYivtbKHoJ/PO52z5PdEebqFXrxEmvCNInLl9QwPm/XXBVu4x6SOHFVnMpC
NqxZ0aQ50Y91hTzKzKzLykx71MOdoJai92e3fgLE+XEsj4A6GYkSJChx+lMGix1lym1uIrk76RRx
DTGzkvVWc47zK/gJq3UWKPZ6hgB3FMDWqRsiktXYfvQ4SR9G/pW2KyL1DbdJ1lsRswyrYYwBEhMb
of5fzsrYOrzKBicWt7YAdPVFGIQz9zmZr350QUeXCU+GEsUHttiBK2imcuu43m0V0Rohq1rAsHok
BWVWspwRAWOHUNdXs7p7fM3QgXrlkk5HFW7gcqfPWWJEiBJmC5ZpynNxhw0W9ZRZhZuCTTItQmO1
rUH84lYmMpYuY0iX2Ri3KqnZSt/5h+BozV6KeWecbGaR381fqvU3NsXMKyU3t5IgR43+cTVJjhBf
d80a9BeRPbeNdivWuIR/SCiLQcteI0EoMrbghgpmDtrn7uwPjnBFcxB6H3cCccczAqL2yy/Fjczn
/0McS7a1OJsAUUTBI4bphwSgsBAfVH9jzJrsXiewHgxi6XPk3KWO5gvQmwT6qQCl5KPGaMHTHauz
MezYoJ2IEwNKf1IhynuiboLKwBq1lz5FiCWIRFsq+dNNvwnKTYlM/i6BoWXZbNajsP6giybJKeef
sXYkDvAzniF4tVgVe0l74vVsxbmLB4wjzcTPt0g0piQITZZj0QbA4/I+8A3qW84dJcb9a2hy3OoA
CLe3TezoifDs/JGgDKbGTOFgP8MpiODwaM1mup5yQo4j3gFrFQM+Ghwnb1ZUVylbnS01s4EYhUlB
XQObrRH1YDkNqNmit8REYCwSQMzgQcrSCGBhb1v7bTPrg9zyTIe7xU5G5Nx0K/cKfqGH+9V9khFE
q+oEtsrqQRl7rx2IhkVOqfa2+XI0iSJjcvpOKxf26fzyp/19S+WJX5lLQfy26pq3wfzKAyhgoUDS
2bL1RQIKCZvE8opesz67vPZMcg2qKTSd4gd/F029CKBXawJajnaYMTe1luWkuzirDJ3bqV0FGW9K
2ST+Cxg+PtMWlnLXeB7rEwTGIci9d8Ad5y2DCXNmnAQUOy+NjNQpjkNI+5LRSNMhAr/TeaoInyE3
k7HZL3Ri7Xd6c82TknDJf5Ubug9rv6oeiOsXFLWyRjWO7s9YJTdbERTXnXbbLxsSxJsFirerKZC4
YuejriK1lz/S4CZQvJjK+2V7R78+USF2xUvBr6KFzl/T1IwSMvgA9K4WBeH8cxQZZvoZTZwliRZc
grvAJNUvQqdSaJyttIZlNREWjaqUraDokFWn7EqY5BIyrRjTbCpHiHkXcwm79KiFNk+U1WtqfHp8
zAdkQRv0SlbJoqXdocPrJeLHCIE3HAunCVitHQNTiAhnFgcBmy7Z3Ay/1MH3DWcsOFfPmZfltfoQ
757ZXC0Z5kvpZTETucer6HoKb59E3nwPaIkQY/hecDz//J63uFuUKm8Vyxc1FupprOeFB7ag9KLO
nPVrEGkGg89I1+HXK7Rvd/sYHgAHOf4w1CjzqDp3sWWTU44i/tURpH0nsZYioTP4YRWnj+t1qNvf
1UxLRPfmgVY3gu5D31YC0aSO52q8ielhPZmstrHjJI3XsQysC22Za6hAMYcxNh9c+ZB0XHHVVryx
IPYk96xO5jzrH/v1AGW22EUciNNTetE5/FcJa2iFqYwiPHqdTs0B0RsXhewEvtXm7O5yEfq2y4AF
Imk8jk6bK4+RI4t8aJG9+tlnmw79pYr0FK7Tat0SHvByWaHfbjuf93RAsAEyGd5FW1/MQd7/cqKE
e6ckt+bAKa5ll/19/drAPS/yoiCBuTB+81KGdpn1fc24Jgo4UCT5wFFIVIvgnbPJsO5wGRo0o8oK
2swJv7EsKaZdQUib+LHNpKu6MiPPcT/ltTLQ8zmuCvSHgvnaPurbvpu23le0KC9mq7TSlyPfoJE7
VsU3xe9SzMuZCCH4dKKwuWhrqQyZWbSnwhTBg/19SezKVTvMmR2bCoBtyLq2SyRYqgNfm9jS4v8E
Ywf1XL32g3XO36DxSrJ6Ai3MM4KVxox7U21Cxy4iMMuFma4B0HxgtA36OJeii+UhQWUT5vJOg+NN
KkGF7eaWI7dEPVQYO8Vua/MJXIyDOR5wpVmOlraaKKsjpWOpuxRDrp9G6otvAqHbOiOWNk900vht
T4izdw8d1Rg9YE8sEWGsHaLA5GVmKrpfpSyAq4dY0otiME0VRiTOmErTyTjOOZgE4lPVIQc/u5Rr
A5kzawyDuCGigaO7gHUqzV4tHuZ6VC+XIJqy86AjzM02qHZD0TYfC0mxC9YtZLzVemo4fLIBEnic
mTCKRuw8p9lGKo+40dE6om+5Q3HJmEV2WhQB71IJNRefSqtlIG342X347cqf4HElNf4GGafaIeS9
mZMjc4KDWKZp1pBDZ1DINiaZVNTYBGoT0Phz5KxwVCVglj9l9NitNw/7r4Zyh58CZkhXch+J9c17
2zV82sJ2p3tUyBxVnMwc8eD1pa2LD+WMrfJoflUgoXMZXlTM0ENqXiWa9uDXaeXXaOwmoTd2naEM
dEfjywyQM/3Zz+skZiL9aanFX+S2vpk77O2oF69Wmz3+IlKcKNnUa8a8CKg6bmmEpUaKG9Y53M3q
Tj/L2xS/g+p34ty+fjEJIs6NLFccNee9Od8N6s7Y+g4tcfMcFtEq4tL6sqTywt071gar5+Ciaic4
CmwL0PNGydXzknbXOUPDYaxDMegCzLtjNFkHCepl2K5v/a9RyE4B+Q7YEPJ9r3oLYAppB3N4uu4c
m2dM6NJ+Yl/QfNlAS0Y2QATPC9yc21ZNMXlUp3aQBxF/5W2gSqX7XrmYjfb4hTi/jHeX4ymru/LQ
rDRqZ8Iz7LF2bQBQgxfvMqHfVVJ8D38jdS3Swjv9UkWyrbDjt76K0ri0pC4kZJ4OzEoKNaS3Zto1
ul8kIFenaJCP5eEktrK7pI9VhV6pAJarlYTHit5Qu21r4cCenny9R9FZiqYIB0ykk4XgMWLH9Pc7
EFSUELysAyT3h/pr3sOqFl0iz8KWBDM/by6GCso6YJqmEuX5MneCGIc5+mND4b/49T3jvPlv7Ymj
nPrzkajd++NYtTj7IMJBOnc8RcbZHrj4/JWX8xxTFp4PkbGHinX9eIuh8sFEw0wgPTagVs6yQklp
amHWZuFfifEzOBIhVSE4bMSmTcDTT2C/EdcQ+aD0qcD0JLrs6ZsgswjD289jmjrxfsItBaOULSru
PdLoeK522jK0Sa+q6pCLwXXwJXOcc7V9jjffIeCZCfeK/ENyLnGXGsTt2nvZeUTf3SBDrSF60Omf
QrVo3yPy7rS5+IZ5f/9OcH/IqPbf02MiQkm284hUQDxD2ijUt4uVZRBLGeUtuK/NrdDHMvZuPw32
spqAw+VG9qr/RHT1FR1POq5X7aQ6MtOQyWiqXFTiZhUz1tkU07Yg/Sptqvlhp1FSqA3vf8+0iGli
XrF5hQF2YDrhCERdCUEDr9k4XRWgum22+PSB4Un6d3SkLt5srZLj3AhNqHXm3DVqVlyKGIGVTfTU
JWIpQQp5h2h8tMTzjdSNxtsKODLPlN+uk8hKspazaL57B9FUDckvKE2AAtpVoqnan9rz0iZD9B9N
xCoe3ALXAnl33H9ekyNCspUqD3Gr7wmf30UsccP1Bzq/Vlu54/hyftxXfn52PZA5uDxDMKAkeAjL
wv4ayCmsILTT6LjcZGqhWuY5vu377iwupBdhgjT2o+vrMZJDxbQPA5pJFUsKy9GqmHixcsWDXIkY
bDjycRHGCL2CtYxq8nvIiQUCk5PfR9hplEHRwZ5gGMZKGMjodqAAcb/WQDWOYQB4VmIOXTdi/WjU
J0IufI9/cmJSQjKWKc82noboe6R0M1eopYW+0dPMFajiPhP9qMIng1f1L7ej20GfBIZmUIaJ62F0
IUQYd7kAvucdb7hXJ6SlaCUK0NaAH85IomgX+X6u1nUiCDhE9NXL+QDOPYQI5V7dhrSQUrfLZirz
2HSqsZ7uPLLPF+T0dObu2oYNWT8UkkD4kz45m6i/V66+OyBzIpYognQ9dLJZnu6K1IcwNKsStzbK
QOL6ODh5lWET1TH7qxVc59q1H1pmowtk1ucI9oZ5O1NOfGujPlqvkJ0KWfsd3R1KdJPgVtih6M19
nfDUMZ0vRF9C1sblLf7pstsozksGZy8TtaadcFtvHsEwpKT088IK7MesTAu2ZKANVJv9au/LtAIj
TeL7SVzc3A/29W+YKzpkFjWYDfN5kV2+9h6NUpVc2mQj8cBOYv6vScyqorTzbPAbv8G4TCBKrN0N
ewXn3lLEpaJZQf6w7d4c3ckBJO33hsT4r2MFY2oGZfl80tpzB6eJ1+fQTYRTNFYrUbPzdJjteWnu
OYB+UdvnawzS4MgdMh2stoUF0LII1F9bpkL4gYki/sX3GaUTdW/6/LQPNmh7aHnO253QjMGBSx8N
yQqME57EuyMd2Xd/FBy0IWBaCO9wQpDKVAB7m9LG3mSbwgjTA87kHSCtjeU+cFhq3VFCHdLBmqa6
vWA1NCnRg4BSiuXrPtzaYHOyYJbY+YrcupJz+MTTmgeY41w+/wpaOW93KW8nJ0M91sqyP+BCAo81
ipmn2DNYCU2VU6YyOx+LlzXYVn1va9Uq7+0henELLs7U6xUISiQgydqDR/sJoVfnEKSkDsxuXlg2
Me21ySFG+QgZ+qwdmWkYYeSTGE+hfOUYMFIw2oEx4rT05R2Ma5L89dQ2V3kDuYFFo0fdHXyVYKYK
uW+5yfs1HL7QNe09RQ3IcDf6PHOmYe0/jDg14ybZlXnI5w9xdmfzbBuVqgL7ga1eZH48cvhTs2bX
LZgxgkSG+6x/f+5loXFwWhmKBK/tS8i6KFd6BQw8BH7/Rw6xRHSdPfyA1YgHaYr+zvu/ShKNib3s
47x7MzjvCj4kyEXb+RzR0pzAZASTHyF2Y3W0RkEbyknzFwjAOij7wBsZDishviHANE3qEpYLaXjv
3ClDu+ZAQfqfjXzXGePkta144USaCJOAWH0iZijSXtsXQBFlx9u0sK8fRkMslSTW2jSJgwJPh9WB
Vi7c2rvHZjU4B3tdGaj3hWO0Kc+UiMJPQEOY9ss1ZBY84qo7Y7vKkkrXDJTlwV0FdmnHa+0fVS9b
Um1aMD9VAdCSc7KTsYNbH/YtZWYQq5KNAheLNWBcck1fafJeg1zr+ANitJQpoyVrBgOPEs8TOXXd
FWoScdwPQLDrKs+JbcKBKx3dKAbBR4nBWmY/516uQQv22ZjLLRUiAdDZ4E1UOJZT4RXv5BwF1ANN
5luec8jhD4y1VsczJ5jyppVv1gS1qdurcX4v3PBNap9y97lkBBT5kCOPEh/ijuSSV+s/24+IK0/G
PyL61OL3ot99vBeO8ubw6xPFO0pfJbbb2xU3tovgkcES/7aobg38yG/6Mr9XS2pqIYahuYbZVG1y
rOklf3O6vXEAERRToMGDpmQNR8deydybx0QTNfTzRunvmu5Cq1nAjbdoEwTY9bdNY9kZb4CShYI2
mCD67a/x9BydLKAGGklU7RprLfp9Re3lGvFD4NDi90FAPkBjR9C8cA7fFONwRtiRzvyghIxEiYzS
gCwWGkMP1r4hKtgrG6q5Zz9r+5Z51czOYkaqqkGq2iENU6U7N/aeOXgzfOWFSaRhMo34QL8JXWVy
Mp0X65mXHUy4GiwkNdd9aF0w8GDm5N0gX2dSB1pzXdS3IrNb8ZsyNB22PMbspiVrbGgNYik6wJ9W
6fIlMFeHtL+80G8igNJIIxaQ0Hn3+4ujXMHU7m3nUhKi0oBeJ15JKUQ0ylB10agZiBKxt52mZWx8
MRzKdHMZLhY31h8issoUV124WWxAVfhuAhb/ogLLVsF+a9hlJ3ITqbzgK8yrqc8v7+L69q2OsvEF
2v+3GyDUQUOckhnx3jnrPQc6xgEZcTibsCniBDBug5he92M7eae097kO3edeEbZ9jKQIdAj0NsuS
I5fqWLZF0y/aMBsNhDUXHSnl5S7Cs3RtzfHBntmJpyjIBwuzXj+YmO6EKnsshcqsDHRvNpbnaPK3
8HRW/5YNXaEhM+XdgXTNqxG1AUi7n9LxtYYnn5JVEiVu8ZvNW7b7wOzUAXesDc+EXXrDS+tAjBDc
9Bn9rGREWJH/m+cdbzV1G7gdxC1PSpJqrbJUiX5E6XTsB0J6nn9fosgKzDa/T8/fz0VzHDNiqiOy
l24iIlFUfM9oISSIKqNpYhsqNXKJn9Hh1eTJCP+VPjXzaoMPRMq3TuxoQ4gY9OymdNdwvzPqn7nz
B22ZkFUBs4gLiIjFiUKIoN2xcq+3jo4gQBJjkfFCBgtQ9VJwX1bbPwuL/YgLbIQrxYEB/TmBGoxA
xbh5txlQE1Mk3avlxstJQIXQpe6FeWXLRyEspqv1yyJG6VJWzKzopzNf/J5bAYoZBSZQ7sRSKax0
Ug38/s/Wb4hmygjyhYy8HnkN/h95fZWJ2JAEhGTwcvGZ1ob35tooKBDts5V3UTBWwXIXablJezXH
qtu5kWMqfbgX03rX4si7LO1sqP2uFMHsnuAVhSktNFjUDMW4kgNLilSb227iPPWFWEIg2QZEChXv
bVOw9X2Wggv0AePfXIEFKK1tmcWeMtSkpLEbkXIlCDDhMaAdcgYGZST6N/Z0YPpyqOhxLBFzWCfE
5yNduAjAkjaHO6uEmHhbKXIaMasp1WFz3mbJpd66DjHhekMJXyB2ge2tHsQ2vTYccSdNksHx7uOy
9Qa/BnerJFe4aMNt7VM/MACvNYg5lCWI73g3QhgyB5wZxCCu65pl25/jn7Aa+1K6bwxU8pHiXP2/
+Bgfna9bOZ77jYCIH1Hks/leCoocWSWBuaadgrXg3Scn2ov2lkFhHTsOO/QD0s5Ot4FkIHRrYE+2
LZ5/fE9/9ySPV2/Fp0YritRZ5/VB/fmed4lVygfsLco5087YOc2T+No1z7DNHgzHInG9QBNiOShD
UdfkLU9YFLChMLI58ytr9rdw+COVnjjKvtrC0glfDXTjdMbKF5xQKhNsnwvUVW9FQmMfAf01APFW
M+xRwRuw4y3yTKIxm+eEvxxwTqsQOYoEMO+WdL5SkF3Zr4jMmtlOY8YRwV7di0vS0susMwAIZDDx
dOAln9fq6R7tXWEWw1a7GyjLCd7J/Kp1bR7kUnun6U9F0+BWb6GDPHcghn2J+fDRTAqvLqZx5G1W
GPY0F1tM4dSz2N9b2UMpH8BUFvo+5xKrW5nrHkYO9brNVjlCv05a3Y3loK4Tfr4QBlTOw0CLJfeE
H8BsZcVdUN1Qo3VORX+vx6W2h+ezaC+u7iJ3K7lqwopyiINYLI8EdVpUytNHUeHT1BWIdqJGPcZw
VxvvfJSDMMnziyPvJ0kL0mqBPdYJCuAL2sICY5Qf6c935tcfUCVqv3mnXYL6dycpMeqVVF7xEGuZ
ezCH38tvpVtKS+iSr4NFzLu+5/9nsaViqWVyWG6FjEdpdTKqYsEPVha45ferbeqaYMSlT2dJsh4v
nEqQLhw1C62B2j1hxGNsG9raKEKXSbvX3rmHWEiNPuG9xpEIrSjAGyAClVdwL4kzksiyAAMJ4Hh5
UnGqe+ldHE2yfDMtbYjCy6wGJW6eWv9vY9ZHF8YEFh/JLRl2sy3o/gmLI91Eh+ca3+GO8MP3D4dp
ZyLxuEJjkfAb8Bhyn/yvosbFvU2wD9Gf7c+vBlY3xiJLr6o3klcSHKV+b3wyZ8ao2AuAWYqbvCNM
mEVN82ITKtNfnZ+rUDb62jhvDjvTtK5W8A7WXQWMd7MqlV59UL20tg0Zi9SYCyDHk/ikAqmaLI1B
ZVeE6blAhfRdnSCGFh59E446pZFo6BEtq6Rw7z1etrMrc9NVeBMiMqfb/XSo4WDQnmc/vq+6v8hR
eHFDdpfRs5PtEYjmqwceoJJC17Pm9KY2WHvx9OnYkVPTsonWHVPPz/x+3QfL1WjFOxtn9bSBzGHQ
S4cj0sJxB+ClhnIpiBpU8Z6pydwZnEeKTAYFuw/8Ja7hSIFmor/V/QMuC3eNILLGg/RoJYgNMZ9V
DFIPWAy67oKtkYrpUnopzORmkY23aL1+QaK6GEA3hBHkbTTSNR5ffZd54xkUsXPv2M7ZLmuzQjSh
kcvAOpPd2/Ofo6S91hPP9e3r4sBMOIxcpMnrFJgfK5FIjUKdnTGfglG6/02LjFyM/WnvjigAI6e+
g8sX5JVPdZ8gaHhHTtkTJNyTmX2fwZh/+cB7FrMGLNbp5v22uiET9HN6b5v5eo8BBMBPowR8TaSJ
45GAMI6Mcxs4cMID+0BOEZHe/HUg5h5fftVc4qqDdb96WeH+DAjnYl0vq3jwYT81tC6p9inLfwWC
A0Rb+gyVS2oSj4XaeL3WDT7x8FWKdhyX2MnmXKd8DovW19/9vc/YhdQ9Hf/QqLkiZ69exgrHpcky
jWe4i1JmL3GwUodSCwuc13RuXdGjhYhHKJVi0e0VJWAXMZUYH8cqIm2yocUs5N/N/HHz9jboMhUQ
Ws2x5oaynbC38trvKZr/KUkPz4ro1H3gltIRA8WhvsT43ZMa5bXbz8zuW2mrIOAo6cCqq6xmhPa6
nf0ai1bvGwEVc/8YPMlg3U8heoui0Q8vwpPclrziVo5aNDt78o7Q5+mwHaCW24fHonGRx9IH9zQn
IPW/rKue7tTA9jV1mfny4o61Gv0r77a+UjTD3rNa/HlTf5MdDmOEl3AIo13K3cFopHdISSrQM4/O
VKDlJPiCJYLmGgus5oJHsD0SzSi6B2BBcxNoRa7/9P2WXim7Ke+EpbZgNrXx8odVjXpdTIPNV+Ub
tuxhdauG10im761heP8a9eyQH6npjykUmh51xRmlZiDyWRcj2quOOwVD0Hcxmo0e+RE2kMXKzvS7
XHWQSYJtxKVv8gVONxJObJduEliTQoKbsvULXy1te+Q9WVg9PLObwX4fO7eaS1k4wHm2yZidF7hc
yeWPjjOPrB48JAxQEgli3XfdqIaeS/8NmQI+1NrmtSNBkQnhTw9RAmcbjMRN4IETMoPaTFwR6tGL
a9TD3keTliRYyDlhMeIceAKMTsNEWJl7h0fLdgCe68ZCdT7GQ36bde+KcVw2wPSOwcoWmoCLqkSP
L1TXt4yPyCdTJPWpUKf8Hf8ZRZ+TWgDhyeX0pCuz7eilEQzB6ZIj2UGrMurmi7fy0TnKEe07STYj
cAEsm76p11/vYqemYAhaYNRlYmYQ3602LKy3T74/eKuLnYORzQ/Dohrn5PQgu7T5atadSt8CerkE
WpFm3u05xNjet/sqrkxmZQ15jWKqd37Vaw0xJbQwX+TX1sMqgTv3rYMsQWqtzRSB0luZsIQhUqvy
Qzv6+0CpWJmHy8A3XsrXOE0H490xRAEmxxA3AqpGrC/Z5Dt/ZnQDBaqtOKAh0rLSElQ4tWUL54OS
zrPXBPy+f964yE/w7KfEALZOquDqNEKr4v5Itoca2ktmAcDFBk2zUtylulryHpGbqQpXVq82iuF1
kOmqYGECw942dltMEvOOg4AI2ILiRTKbyVq8QP/SQYupGVzJZjO/1QufdTybva/EGQ9iT8qUiVB2
o6XhJ0QppIJHUVIxlLqtRKUcrovBPCdgOB9o8E3ee5Les3ceDvuHdNOywBnEiHv6bgWSoZ1wageU
e5v6H+jop6irF5FqNhKaB2eVpfVH6oR4+Rl6Ut6blx+RDa6/dXsr3ct+h4mdi/RTWJYXvGP9lTg9
66ILYtCQ65TBOEnVAvg6LTFrw9swJsAYgHn0h+2m6IDzDwFo6y0xoCarlrnYUE2cGbK5VJ9wh0/v
sMKufRt9kftGnon+6UCOoDWXiNx6StoqbhLLkLIebNHKgBHM5iZdamM3ytZ/K6kOxbiE+/UD9eHS
ADwZZCkEGPY/hNZ+L37AuEsxtH0HGfYiRqELDx9z9g7ECY0vaL3Z3v++7sMp739ZwGNS9q1jP5q7
nhrADUDXR6Tv2eJeZL9EfZZAturWYN4/lT2M+pERTek7nsVHXPRAEHihJF3J+HXO0a95hUn8p/2r
pkfpKKomCaGpnz+8wUZFs7CHap9Ucmfr9B+pFxyIMZjz79h2Jq/mZq6Ab7AvqNXsherSbaB+ybfQ
Wa2wWN0QYZ3Og89quTkH/dEZLskCWcZNLFwLbk8AAbReLciHHpMYKhlT0tzbpbgDluHTAZp8pCHz
CTOj0gdJ9SbgdtIdEzd3ck/9jlV7Fy0Ei9Z5a05mFQpLiNTa4eGrPZ3f9pWOh4JTZ0nDgG5myR1r
WXHBFvyB5aY0oLWi1SBkLMWNG/X8Dw41Q7vWxAyXUZnXGEMrovkXbE/QHx4S2ymS70qyU2xa3rkm
Qs78PQinp+i7v+A67P0zjbQ90KSWlse3ZKgNTdANrvQnyY2zDy73sSRtw8iUpFvJQYB2MeejhFBt
imgp3GbhQEzogow0ysnrXmzSHJOt3ced62p4DHkNePkopeCzFw8LgNJMD2cetBLoLqGgNyrKqLxS
Jjmi/wvnNdRRbRNGra9EdB+t7W/AM+ymKvpcMPKRWYZ04TEdPVfmcnYDwRMt326DGFl3aPTrg4bD
lF312vkKDDodiozLqSxDGcfR/TCJjgn27wTeJeJZuORDxLWlNtNE4uVDwqfyuNgYvxTKrt9IcgY8
uMnx1cou1mUCgHRyrpdANEWZUYA+oTrSVXZJwv8cYmfqgBXbsu7YvezIjvTUG+bm9Ru1g3NXBN11
apBitEx6KKC1mgcOWnJR1In1HN9vUwjuUfXwY/TJE6j8WuMbPipgrvLXflAITBbeNIEw3bJKrFQi
x5o2WnfIVt9zV0V8iaA/0na0LhP6NHC8LJd7354Mjr6zziG79apbWcV3B15ScGEn/s4PZNqLW+Aj
EUeun6bO7m219XcuC3wx9bi9xKrF+ImXpmwtCjNODXe3hmk5RC13mOb7Kf47fO2Y67bsbdawFmsp
WQP1auS8NlE2FKd02OLOf+a5TWTC/NCMk3rLQnfpYihvCcI8ZSSUuHS+27ionhH0eMOIry5tGiPm
w8gsFe+EeWpY3lwEYuzwc/DceIzouESmQYT6j5o4xGpMEPQBFePazMKPDwcsA3eulhOxyYtqyC3G
KZkARXLTK7JL7/5z8QRT4j6AY+1c4d+KLh+V/8EdNT6OOdztcF5cQNVozYoISx0M8qrPlOp8BSM2
gDBCCIW2x4L83G9dUyLxlsENjAR7mhs/2kmt1nq6YuzA6cklYKAYHZynS+v0mx/7Oyyj7k3hTYkY
aG7KCIzpZg7vETMiEuSMfx6eOoE2lo5Id1FvIDklhCzDuEGLBgPVYR7cRcL406XGUvsK5H7uenhX
K3mn47Ubb7lfpZGBw+XhDdnkYLTi0k14XJCmgAEQFVeHpkNFj6PvpNGYF29H98k4lEmysbwYKSJC
p1ygb/RgI/hfbjNF0WG3d9n17MogoVGvcsXUg9LhJxFCG758bwvVAU7WvKR8M2rLTTmlL6KkAClI
wBOA3x3oiX0Xr2LOYskhp3FwzbmqvH1IiTugp9EgwOPipYd3FvXXXwKJwc3h7Nw499RF4kdC3i4l
tJMSaHAsm5CUCsonLMvsYqhgOJeLNPnVNwQlXlpmNYoFkx4e/W2+IjoGUrWZ4QPf9+oj69egX/JU
fl4IwSimg1mavE4FeLn27vjiURNulz/e2DJfXMO3wndi9kz3Q/fFxeT9PPbg4vv1dPYbmquGtobI
49H8lHeFo+NUJZ1yGgG85cpcvmP9qtP+p2P56GEPTHSTEJEnri801gOTkix+ugTusZAt44VvE8Dc
covYipu+UqENgYqlqAoRjn8QBTNCS8X1fODmz/oYHCHQO+Hv9GCWmhqhjmibUsOcReHKdcyfZTkE
Vt4Me546nxIo72QYbmYp1FUGyeX22R5O41L1FXI3W2nS/CT5MwARd5W0AqidDpbMDN6bZxYQD8NB
m30OCTLrpl82IC5teITMjdHKkSi1YgF7e5Q1grzUUDmFuYJyVKCe+ozSHZvxKoP52JKbGLO8tlTs
Qech0UpUkWyt2m+6OB28IOOGfqP6ltcdwoQxFyw+27pkhSsqgLLi2SF7JFRLs669d9/gepNDyTNH
EqCohDBDXlrmTWU7g+99tPWRhKKFhPk2unlIQHBq64FzA4dPbtCOgsD2CoCkYoytv0/3bYapNtZw
wPrwtCnD8+1Hi61d6TkHrf+BQyvMdS+bMK9RSvJ9I+QfcaM8/SEqa8Y5xfxoQSZu/IQY10nAChlR
JLan+rb6Rha2Grsp8Qf/G0mHG84/q2ZujFWKofhcgHkRGBS3nG+iVsFi18tII1e0f2DNUJPOGM3p
lSkmHOefSi5hTIE+5uCci3/Mi2MN+eBGfewCn0RkULhaoRZsPlpLIzwdpsMwJQHWSFox+Nhihs4Z
06DQFleqSl1OgJP/xZ/mbeoQzYfU8gVPJIzEwFhnkCUgJkAKto36aD1Lfjy3up/8FLvNs5c5E5Kb
xagpbGJumr71mZtU+WXiwyHDrqSJOuhl46U64YavtjiW4xQhmMbBd/0hOZQGVn6SFz/UACe99tgg
2uvl2BZS6oNXmI9IS2LlmELFNkTlPlsqV9kLhgXhqo2o0SMvj3Dem2KiQX0d1z0U91VBER/iysTW
GyBxexmxgN1HaGvjd+QkfxUmON9jpaABwDF1AEkL2Q/nhxpN1TO8RbSxohhemG9Dg/OK0BzQlcpL
27ypbdjfJCej4q526FdCjMoIUv17f0aR6wFYm2UauBo9zV5VWdO4hUZWNHiT9IXUTyJ/JxBWhkDq
r7he5BThh5K5el5m68wRH9OMmBTYK7r5Hg5rAfOEa58ycDZAA6b4cP0CiFFrzsfjpeHJ16F/hqsk
jPRuLw+C+hC8VGZX0dQTVqGZYONIoDcxLHfZ1INaC9AZlCTO91RB9tWYaS4riNB/i4e5qVKbU6qA
jJbdI/r2nHHp5BJHbhl18zYobV/efSay8BHF7NfWsV1k0OyxW0oCEjU45GAqiUydaT8q/Knp87m8
Dto30BtY8IfQIb51Q35RigWXol7WSlfJShAmjTUMO64LpHllXeTXb00k6pOOuqCGrKC9Lo8iWXrE
Oc5rlrnHIfNpVHEXD+6k2N3LH+ue2KHxYMw6gc0KTUoBxJnqMxpP8b8LDfDAjL0l31nVYBHe8+hq
+dqEpH5cQJsqNphAQNpl9S5v7LS2Ldt6IJmGusmw/xjKmLBlyjYwrg8maIZ82VUbjK+1gbOXldBn
gCz6zKh9zcPiV450xEC0I5Av5DJ7mHJtkWiN+Eu8Cb8jLGvc6iQh3o60MSfvEyw0EoLjHN1adRpl
k0znLJJyiVnQahAnNj3MwMwotqLf9u58eyBDtJGCpVEkMiYPnkJs1rvBkeN37hgzd8hCr/pEozu4
O9ZKC7i1gjolzzfjE8EPFrhVdyfRq0e2bynZ+qV1NCEoiiUT18kZ6YuPKf67drBrTgOJDQlwWxaO
FrZl/3GTFuRJqIjsy7f6uAOkO/hhXdsA8QLNKylMAvHaKsgqMNgkKsYV4HPMP7m++HhwA0GFTOg0
UxBgrq3m5GgeorcHkEd4V1EkeEZUBEfA7Oyhd8W5XWdGFuiGYQCHvb4Lqm/apoNKCfKmQQk16vZr
NoCHFdPtM6xvuf3dmPGclEfjb7pniM6+b/4FPsgM1VgTZfHfLci/TEKCskM3BiTcO+PrCxZjbhrY
Ph/gRow8CvxHaEn67717eWwl5vuAipgSW/5ciH0+7FS8q9n6j5XekuNT5CCV3vPGf+7Na8iUDprk
92775ffKbVkxpJvG62mjYa4wF01OUVwLEa+Gc+7hQ9pJSm4vqw72TnnFjIMhsTz0yD0NIKAq4sba
83uOiMdhj9ndsv2Mxu4BUJn3cNlJ7QeWxTkWw73c36BbO+3D5ebBcKHeUMOJqZxELKvA5X8055+W
y1u7OZ4oDKlYeDArxqSpH5kwIHpJ/qz2IYeddWYphXza3joe8wQ21Bqzk5TJdUl/aUMqEjBtrM14
N31JK6FEazRnnVJjn4BB+gcsriWXeZq4xIyl9SkwFdi8vlLKlJ0xr82GmAcF/IywpHCSO2C0c0kz
QkAi2s5UXC9kyWPv823zSY7m57lihL+xYeddP6uAElQZahjTqyxGdk494gx7nWPg3cCSQs269c7z
t8Nq/UB08nr0M9Z7i5yuJhq7NzHOPu/3J+2JxfQ88aFJcOaiMAAU1BtW5SoQ2CyrQRrKIwRShN6q
7EbtoGWHC/J6qE3hHLQhaTBm3QS1kx3xHJe9GdNVmnMTtJDEseY6IgxkcT64CnzfqABSmgJJpzZm
v/ocNlKfu8eJ32dLd1maGXazsgDYWpYoyB6BBmP6/tDcuItNKX/5C+Y9QZSpH/a/efxrCyI2PFI0
XcYdwhbAhHLXci+GDSxcv22+arkWA1ynkYbUt9Ytx6mfZcbJeNs98ZJdedEU0CvzJBM2r0TRYoID
1K9N2/gBvDvhy5WUHCXOVC614zPmLRcfNxbwqEYZzP58V9fzXN6X6UbfC/5yl8CF1KALU7iZnkpm
tCLkNHmcMO9B6tK0LJ0pEf6Ci3fGFsN01/Pq8/e33Dv1pzyVNaPT82JBJODWQDe3eWqQt64d6Wpg
+szTD8kne3D3T7q0U0KxKNWvyV0FvHTqk/CXya/136/x2YGDKVp7wh00zYcHQ41G6zAHhj+pbY+3
smi4N2HKtAYf6+tXTNlLuiMgvTQAZqZdHnQzPvZ2LIZUk1aEKF4Nh6xwnyiHyINFXsj9m97HVxPh
eYC1H8cj5Th9AHMlUIUOR9HuaqXDjQ66CuRdRniCaeZxTlFfJYe2Tx0+CxbsfCpPGEYwpsYi2IWE
iFaw0cczR4VAeSXCkB135daUU9DdpujtqqpbCu5OsehuXgW0PUiZqL1cTmY02LAgE9Ab0hUKNU6f
9sT+oHte2U4PqaZm7knaosWlBmaEcMYr6nIhYu0a6+olzXIvSh0ESCnIvQYwDrKeE8H3Q64QizMr
L9R7zqqTPr+D/Ox+n9qc2+QvMWdAeVW7g1GkRkQKVScLInHWrUed6P4cJ30yyU7a7d1irNyA8MJk
FUPVmp6+qcTjekBeM3CA23LY0fNKfZBMbIpni09hUZPESfMqt+3/6DCmZlQqWBW4+PWy16drHe6O
vNAchFJOEG9xQ3Z2QTb9YKIlRokDDwUm8q8XPiN7F3Z2xbpiA917mQn/HrB7Q1GgZLNcXoTnqhHF
ZkEdfw1LQGLJ5lgB7CZaGj+1BIvaVjJ1iEknLdNYuo5BIj/dPMRbL6IofbCi6vpmaVbGhWU2i83E
J1SG4EB0RMqKSvOPFJ/FGrbx+T6FcELEfDCr1kdg61CirwjTSZEfqoBbevMWz0r0e5FlS8KCGjG6
eWUueNp08DdgzPT5Kz+hbBAj7dum4H+XEcFlErOEllznXAV9PwRYWG5/KAoW6rmR8PKrVMSkfvpC
ZyGr7KiXMge5KCnFqvLlIYC5iBM9hc5oIT15tc3i6SXJ2zJegSqY+ow31Xbp6bzsAKncl7wkDW6v
6KXvxB80xtpbDWquK9nNMByBZsNr8tiJg6Bv/BD2h6G0h550MwgoXpxtX9lCaCxCfW0U601mreHj
y6bRRmYXNdNyICvwHecr2DHt+N7wg/Rai0oPyiSvmqiJtahSBIMLX9ouS7vUbjTLwCGCCh2/NOel
FvzE608FuwbGGoA2u4wg4gkraGfPKi/QvvjJyo3Msa7wZWZhT4kOdpzSe2h/QbYCb/KwD98dTqAv
V4giHjaydakXOigu9BNMjyZ+EZWlt4PTV+hnoGVGqwfV0WMXjLOnQg410Sv6X8CBz2NB7w8eA47I
OLr4MuwLiOK4IkzdRWaKlDRR8ww5PLN3p/fXSbhF1cD5Bmarm+K8hVNiRoWnNem9/JN70dSVfwwd
/FdWySW2WfCCKI4B1kRKL3Cw185xX8x5n1Md9Fcu5T+e9LvfT65EBrC2CmQBQffW3sG+fo2UVbeK
NliXleWhnwiOPr6WallnNDs7ome0pfGQIBIWlc0xW7bQ6dIOXgru8VOz63Cs9eRCs16ExMK2Ve7P
hFtBB/G91DkaAOUE+VfgMcK7mHpbCNyrnDgdKH8PbeNF3ysfMq5a/9pE0FFBxD1JaXkevCTra9gV
1TUhuihxUkRle6joObhI2NTtAT8mHQ0e+R9lX1fh77rpACxE5UeGXL9QHc1zqv5U9hf072b72dKn
gbZvNb9qTNhbxTSu6D63tUfF97DVphIudv8o5Q+My4wXl56cbUZoN5YTJNdoLrgCwh29do6HQi6Z
y+3QzimCA+gkgsQ9HOpQwpztbk1V2oxj+P4K1/0L8lCnWRK09kR/URCESd4jJhRdeYZg5Sn8ev+F
YrW/hIr45yjBo1f7r4jDYSq8LGSzJelW0heRLwA2qMJqh/QRt6KvR/nj3dNGaMvjFXuDc8iwABHZ
1eJTf/XATylhhcuFZWRvKdUkut2kTYeVRYPBLVlmBcNbwjF2nIs6wpjI+Xx1GxqbnVvJvGc8bA5Y
n6JLyhl5CvgqE2bXaIhNGrN55F6rv8v1T6vH8hkCFxuGr5eh0jTL7vru94wJH13r8yJObdqLokTC
WkBjOoELPws60Hvq7rohLZFO4g6NRSnB8hLgTX9GQlBhk53HOdQPy3qwXTAMT2e8dYcWyIkSnoRj
iuMJ4Xn4SwBcbDEdhrdYLyAhtm6QDsiLVeHwRvfZSAjFov2PYWpagsr8VoMdcDmXsKkhOgOAQyaZ
ODaGojwKy7XO1yyAwndRzjds51s7+Jm3lmgP/MqEK4fTtPA3ZnDlJfx93N7D8W0qCDEr9zoGzatD
qIru81dQBzVESLRP7cm0WW8V/QTQKzFiq6oh2JyI8GlQHLHpTQPzkgtt4LXlxUXVQhOxeWYzG3rj
dshN56YUSR2qjq6sJbwWwjNC9934EaMK1HhMTjKMu1ooNGGDe5q5C0PkVtkGwev0HJf7WrOHhUoJ
8dAldYK2/hOAH1wDH7ow2BIfWkAgU+EjJz7iewvPHcmHq8USIS5QVzPUh8mew7MwEDfaLbWwq3NH
VQaLr/K40FWiEwe2wZ09F6U69Yq887isGN161Wa5lVpX6rGdXst26Gg0F2XK8aPTx16aNfYZZTT0
y0xS1O/l9jehDDqUbe5SkDN9gCKb4oebBok/6iQ4wo+ErhAbleo/JnR9g4FpIvdEGGugCN0ZH7KK
fknaLOjiIINKpHDCrtE56XmsmJyLcJ5qdE+XedNVIStg65GuAYE8nd8/GM17sHzyYxqCexGe2iBa
gX6JfHyyi8wxZE3PeNDR53/SI55QMKKTejkszkOmzdGy3WiEQY9dqbJuZppjAlD33bGGE2j6E2ij
HxQO+L73qlbr8lYHPOLAkABjoV9YhSWGIv0q/fglQD276x0900YfS+zi7CEEj4eFQ1KjGyb1jA1a
auhW97xD2VVE9avAE72ZgrrRQC1qTsWGNkgIhz7Sj4B606R3VVMoYM+1BJLG4osW3StnG4ENOuXu
maJ1RUS8G6KE471rQU3Rv19rc7Lkw6w+UEvc5xvlMea3oyf99GrR4z2uY8ArW3rUPZPQ6rFzvxV+
WLpuUh1vULVu4Yv2k0GPvCzjV84IiiUMKb6axvBq1MuEnqwjeKaT6tYjvwhvvIMVA5057HT+sP/F
3L3fuBxAJKJ8ml3YsWpuLgeV2l6EPC+xZvFpwbLXkN54W2mcG2O2FnZAYfQZh2vTnkzeXbSLhmJH
IF3MG7bFUnP2RoxIm33FRaGeIkeX0LfIo+up8joaYDk7tm4zTkmu6vvqC3Gy9e0r5bJVPkmT7c6S
dYTCOKrMxTQJ2d2AOEWfJI/y10RUULEoluLOQs/+AJefSfS5olt4MH5UGTYcP53+qBJ+qQWkUWc0
HrGN2mQMIxCq4oSS+rt9X3A+MEkXlBnCgdo77SWWG24A+VZQlvMUolULVunlMMQjOmtWYe4QVdaJ
gLING7Ox5VlyR74Mxm6HVs+9qE3jxy/y9U9p9P0xlpHkXiIrs1mpfm8I9G6O4aLREEonhqzOEvY6
G8Sk9JXgMSyQFgHvq4XxmBM+VDp9ssjOtAoYfu+AqAQe1Q5DqfHnDUwqfAOWeO/VLYy2CWMlOrDN
NnsK5fiKeuUA2nMB00P3TCVap1nL6IBRaCZjyZUH0U3csuBq9FaUmEFweD7O0QqpSd2I9eKATDis
WYYWLr3UFA8gnaJiDjcwC5IoXonKQpz4ouGfueZRBMcl+g7XvhkfDVbxzTs1QcDDtfMmheIKLbo+
nHsLPVOrP5kdbuEU5UzOpu0Xu0n98p20jeO4cBeP+ss7BPpZcHxjrhwCcaSFOGC0yTuYANtPBaA7
bS5CB1vsbYaplBKIB66Rc02eh69a/MXdyf3qogBLquk3LYmvsmcxGcT6OW7Fv+pzH4Z6xPvxAC84
TkzgbzJ68/8WeJ09FndZq1vyu7BdYEQrYnK+MOdjPKhBOe/aOjAtIL1KB/f9I1lQum1zdrg8hpzh
/BKlxJ9O5pPw5ABjvPissF/ZRUcLk3K2in2n8pTPfl09BFoya5xZmeeyN54M5dHIaxz0dRF/YpAD
ndaKzPeaMhgN4F4/1pYubO47Y3Z+rArDH1OyJwwr7JsmU5+ftdqoDETnchlHKJtCNTsTTYFfoucL
4IA7miOu9jsn6w4jMlxhUJtUhAn+wM94DhYQ/xOtXjUA2OtVbabgYeHekMxzL8KyHZAk0aC+SRkf
Tcm31kfQm8YFCkgE6ZD6Tmrhqnnip+2UYYzuSxuhfHMxkstYMgsWt2its/0ggwFzVRzS/2Rh0PHc
6KeFMNFQOY73Rc/bQO3u9H05W484O0NmlZMgV4yiaVgDOuNV2nVavUAP2+/rAVsmmAYMSNursRjg
XFK7BWoWXGmEIo/59UaWx5dhCdT32W6PR5HPUl4Z7z8xAi7ELOJG7yp9fv0fuPbM/liEvxNOgwWV
582owR4hBCv651CzXOxBVIOCDttjEg1buSoRRYSxQCFe+nv1Ydm6ITpksP4X4P2fAAcj8CtmEMy9
mwVkmHd0NbyNfJVjxxt2/2Aq85aEoUZUS6Q1q2efKp6Sohq+Nv27W5/cyZfftXbJy9OTs4Lx590e
06sSOfy/d7vVh5qCDvxLrqUYqhxeQ5K6VrkBhJYDYwAy6Osfy7ho5RFNlNivqHAzsPy4Z0pmNIJk
EQEndmbsiBBEm49scb9uFBEXhqyg7SJPcF4AHcE+orD8x4PiSbKlasGe6uEh05SrM+x/tPhxwWBZ
HMTRo0l3jjOxMQRY4IYci4ad633e6okNGIw081parZAyIgSYoMMtcOe37z+fjl0mSEZlnVGVZb4r
8X0BvMTM2YFJenmkCfhhuSIA3wwQs+mzw9jKOZhhF9UoSBaw+7Rux7/PGHCj4O/EW3ROVCJx5YB2
L6WvMmjvRmTlw8xWuGaVQ6G97oXWtsQMg6mh50YktI6U1ixkl6kNmay0ShYpp9WTPgSr/RpoejhB
WHh1DGnnzmvzcVhBdchb+KCNthyMB6wJzoP9huXKUskZpDqKb76YH1iewnMDcVcEcfJ/0B/ANUdk
onZevU/Y6EHWE4Xy/Qad3F1Zo9dL1Q39sxitpP1OIvNpHA88V8GtvvvlxLGNMYGDQrkXxkibYYEk
V12eNO6DBo+u29y7ZSiNnR8JRM6V1neoHk6wiZFb8VUnTp+sA0B+N6l8hGs6hqAR0LvOCBs8BEo/
QFzVL9HH4zSWF8B583EFHv8dAAthCH8q5OMDF1QVq1zPaQMJkqaLeAHChJ/sjWzbdKgBjNhehoTI
CLtLxsbvq0goCNDq9f/idR0aKNO98qKDdB407pqJsMRdBwwIdMjppmnEhBY9bfqomYfQujyujM1a
W5PQIVxCwud677fVybg4vlS2KPVavZhZ63EuNZ2544m/j6hcqWB81OiybTgO7/aagY8PaZeIPHmd
IKMQKct8AVUDr7l8iirjky92tzci8gGJzIB+dT4azEbXBfTgtd+qp++tlp9o+d3RTzk3v/KKw4Wf
XF7JvnAfWb7+pXe9tYOE+xUwV5fZLHaAcMxgNBU2R2c8wMcWSLfkac2VrCTc4V+BqrtLlMATl8AX
ffoMg/YaSRXH/Yh7RYNASXsAZUogQruWGKPQ2xD45F7tUrisISevdgJyslMHfnFy2wDA0qWJ4yQT
kfOt0hMZkQ5Igus6mhlUYYQ9huN/VYnRW+2z+7CJja/N5XyqbjGm1PP5UrqIWpYJzpYW1p7WlMGc
bJPTvi6DxyxJCm3cSOyDB2uXyJpDzSKZ1Jaf7UaEVQJRYyItEXF1eam3ETZ4WfFQljdhA+zB7zIA
Onae9FDNGSb4LjklVNJ0LaFJJGDmg01sM9ThIRBH2twxF/9l+IwEkgPHnwjum21QcRvWmphfwLIv
UaViLtAXWXu4UAqkNbKzIxlCyompThpw2EhgmCe0r0UoGNX1g9Wj/j/2Q6e/S5MO/Zs5JFkGiiZ0
XcpA+yCRubWCGmSzS40yB3lSY7AEKXt4vo1/TPDyLYySVENyycNf/+C0UWm3RovHklrkgww+/C+w
sMjJdw3S1dhnFvws1Z+UwP8qbmbI8roVwIUgOWYOqEAduiv+r5vPXxIHb7CM/GnYLA6ODQnaqfmR
ZWoeeJgFKQBd0srTGe5uqkmfGwzPA0pcdNZnjyOL1fIfPs6pmD9vYf04hBInnI9KHE6q4qCbPP/2
rVeVQXuW2Vwl2SVntLTRXuXcepuDHObLHuCXvdhZhX5AGyQe2Sy050XjylHCiz0jZn4xAKW1xhti
znX3JqPasNbUBAJAmyqDQD5eQ6iA1DiScqxIKayTy+CI+MpkrAScDYPwflG4djbq0sEGZpdylsMV
DtdwGLhCHYOGwRL9WgdbtlYWsBHt8bFNenVGHjvd/h3nqNN6VeeviDJsybEl4m+Kvg8H9J4UpZHa
jS32N1W+fWFEJXPvgpcmO1Xdshg9XmGcpq587SWBPlkReKywBslX8cG1u6W2Hu8eQ6ZoiHVg+mLC
RWyQbFwAogmXJ4HZo343/Bd1HEOrMd18F762BnSiTNoA8Wlnxyv3wBQOllwqWOyt4PzsDS5TtOW7
Vdi3BCTRrnel46HUQgJ7Z9iVqxl/ywa4iNhrZvw8gvEj29/9nx7rfAvP7yJHVDqUr975Q19i8dkM
ZI5tszsxZ2v47SLQ91NpWRPTJCLMx8vMAT2ga8+iNuLlcA8cIwHfmAp6NaNsnTt6iW1JwQj/6o1E
u2SuKBitCENDMT7oXwWVsOrc1YHBQe31ScVfMWx+8FO5axZpw/d6bTP3LfrWvu7/krsrwGSbE+/6
CBIXDVkfDMaIg8klIAjd7Pn0u4UUgOEnbPDg/7s2p8lxgEYoXtXuPmojchMoTdNsZ8YWO+YVbbh/
tahQaW6BL2VyqRSRDtreNWmcYQfIrxAQ58hYh/wrXm3gCRFrlxhrbyPXrhWEz3N3Lh4NGhei6tzW
3kdBTWnMDE8QNIVM0x2j5QBY3vWsUP3vSxXAQZZw+qcMe0hfq5fkF9T/ZsEJqfZTbn0ytKNP2SJD
TvPzJohkrrjBP/vpAZ3KeQ2JWyj9ThT02gGNoVJSm3tCa5OsJXw58UGOZae5HnzLPS36J9UFUhTJ
27XTIZkO196PuX7CyHCA5HfbJdOHaCmldiQmMr0YS7honcHwngrNrml2PC57cWXZ3TLazkG7vq4b
HWC9J/kfZldvDBgkfub8XAkmrTEuFi8rAHy0sB6lLth+bn4y3Ydavf3J0o2wUa299Rurz4XgvXJY
BSlrpXe5PJKtQx+eolTrxSaDI/NreHxm22fmx0AnLhvaQuukFpVzFlk+AupYwmcUVF7M+OllC4MK
/ZhFDuG/p4h/FDUlhAQUS7fJnBuCH0Dpy2p2Y1J2o7SVqecIOsdCSzR245WYx6isx1bzK54xTq48
htR0IU4Y+d5YQmspO83uy4qg2ndYBuH4GE+6ZIsYLncnSst8+Vf7FQM2UdW9WaZ1XNRmoUi03DwS
t5079yeRPWmDrTuMxt254BrmgKdx+sukmI5PzTEV9sPw+K6M0EAgrMS51MWikAbpS3xKUYWDyt0l
bSOoPrhJOFsXLR3JIpB+5Ec7SFSqeh7zUmgJ+sSxpH41AzIn7SsxTlA3qjEU2kn4k2Onf+TqxjYn
kxVhQFYw7caGOvxfXEQHRIlpPgAJe8ZOuVAR+/jtQ299PWZpE8foBimFt6UYuLyDxn4G721Xqa7g
hzSiCcz6ZoHcN0qUMgv356UM24JCohM+Qiy2Vk/GX+uAlsmVrD0f99GUj3xkZjdeCYS5Mm1tZMSr
zY3Zld1UKyEl60IOPXCgG9xfWOHoQ8og6Lvy9LbGlFiX3VthwqA1mmVMG1WIoe93mJQiIrqzuCl3
k3daZ2O303Vxhr0tNwC7ihMAjzsdeWs0YZkSxoWAn4wIe7dMg0iUC50gNFLf8nnbbwLOiznmX9bB
OOkxAz9lfkh/r9PHk4usn0J7kWopkBIrSUBF+aahhb5y8GoKRC+O/58il8+3D8GrMcysMXfNydXo
kMKfafy+9X1T5Quss7qTJaFeX/8S3KpsDJ3H3bkSHa4PKngN1sMR/nRoNZN/jrBNi3Q2ezVKCs9R
65WPpoEUThSAQZKz7uFJubhb+lyEtSN9xNfHkP4YHoPMTEJzMF2xhfZHHGpP2uRue2vfVM+Zm1tA
/7T6QATwfkPHR6XrZGpyjzM8Oiu8YhmJy9Xam7K1cGIT8DMlMl+tFanJ0AQTVwyAwtOB1+isURNg
uXep+RMZvKs4wj49MhaNTPFifXvDQoLsRqwcm5BJ8GeqCb3KyWx13iuT3zcC/RESGGtWh5NHGiOT
Ud+OaPVCog8tTgTMAahnYk053QaH0CMZ9OzGNUQPCgcJXfMrsSFqSkolZoUneN7U5uU6iW8ru/4i
avSgQ/vTe5RCtMtOvvY4RHW3t1lYduHP7zsxhgLs2ADiFiLKsHsSB8VrTXwaLlB8Fhf9JeteDHR+
xwHNFpTVjfC61SB04dy5ZXVsmM8+dwoCYPoutZrkL2gn5pP9KpKmvpfMi16QlQmPVL4h8QMNdOd3
C0nrGf0fl7FWMaKFnstHy+tMmmMj/owbucL3gSIpHdTox8HDtLd75LliE3fIxIZKAE6kzy0qXKep
3zE9EPLw/emnnRQAx5Z6v9O/cSi1ZcKF+/1Gza7b7jJiso48/ASF5LecXpj2ZSe6oh9moX1gBS10
2f7LW+SImkW8PlaOyQ50kZN3/jCnt3AArFbxnWcbyCq9cfGWJ4E4ZCjd0l8JihsHx+UzqaB5WiAF
3Uo4LFfQSzXl+JW3Z1wRqFJydLc+R+6ekPKueQ1ENj2q+TtpSRPSR/gRJZZD1r9TWvT8Z/Suw6ze
PHzRpyxRmAE3wKPFkBZtP3XEE7gL7s3bkPuzi0bc1nYVg8deEp+CQmgM3YYNLWz9ahDiGE2Gbygr
aD5zOuPRkreSy4fCfM05FCiIEW+eqgNNWVJ+1za6d5WxcdudXy/vS/4ht0YlybqTu9RhrDsa/yS7
RaU+hqFKWIDHZTeF9SjqqddjCKRx9QvpWyI0WRrhrsm7Q/EQAdoKKnQFuQXsVdVaAwc75PHgzaWp
i57vHj1Nl9ouOYCqCZz5B+a23zVT/l5KJlupvQOkWc9P/i+FrOI/zFn4wcVAn6cMs8Mi5gI/Pkxc
OXAUchbsb0ru2YZcYeMOaHx9mcRT2nhRT1v1XSHc/taHkPmrIEu5T4vF8oE3oAy1YRUVh7y2aQN1
6x6EUEXY2ieNYeTT0Imn7mdrRsHHmmmzfUg33rTY0+hYTpTrn8Fg0TQUU2Qw7GtoWZW4G55dO5ab
EtYSWfZLs4mDXDKy2iHszPwssM2IZM1gjeY9IqFBGVP7hbKg8JxmjB8TDiMLxK4BihunnUGPm5ci
+WGpXUIf8Asux51387P26/ovuPNTTLQ1ZNQ9cRhT4SYUxgiYbJ9cjazbtC/VZFO2r16aeBl539ow
PQiZfETb1ZyCP3iz5p5elbTHeOEVAgQftJ9X6zH11H7nmCCMRgIUwwG78C4JbV61R6FYdmOioN8R
vG1a9O4LzFHznX2s4GAMHUv4v4JPj0JzqDHjyj5/hdc9SFcRbgc8JhvEx//oJowS9oEuAvYxdR5D
97cYe9FzbScYP3jIXi3cnH1OpaR7fBzmQsLDeLUtTPo6jXMUsQdI5D8zDvN6WFrVV3mUpeFyMabJ
6+H4v9yCTwfQs2/u3Linzx4seKJ2wceLoAgcIi7tBumFGqrg70KbbW5ui6G8a+HIZRJ4vToASwtI
a1dMILZtZfiKIqs2nSJ/zts3AUbrSz53vDlysEla+ChnKJUUGCxfvvtgsgJ8Q25cObRWFulvHOVs
2llb6yemwalk5ArXZ0JJ9urt4Z8lUpdgbZVV7nx7Kyg840Fz/MfSN5RqFHecVFJriS6HafOll9oz
/taKkzLdhL4bTuPCo3RFNCPZXbvKcJsqKESiiOFRk+ci+FrvjlHjPpY7PwuC/gvFVdJa0CmtQiTk
iS6rcdtwUS35vOKIccir6uF1WbFc4fKqyHsnKDvedHnaXBL0GWFyvsZ90Rp8bqf8Khfv9Ekv9w+C
rXGGSgtHGcETV/Kq0DD8epDyWO9M7C8R6423ymCL0vyO+vaImJJOg/vLIZaWKl4aTCggvJ7AN1g4
sZ2SyRSMsO09S/SbZH43IHbulXOJMWsRiraf3WB1s7jgA7pRLlHSFLj3+U9Y+02AFMeVez4k2+7g
CpPpFT6IHUZ3SOnVJXx3eS58NDV2kgVDUMZXuu0ZqpLKQWaLi60xTDbonL8eqc/J3meo6tQ1z0Dg
MCeR46dDvbdE6VZjY22E7Vc4AiE2SVQanhuT06EIz5Eg7kVz9y4EToKGv+RZWw/UEDlWAjSFoXRM
2E/uXgMQPXRcy81ypzVUydqzGkpF4Rsl4u8WPTc6/TyRCMlUSTZj0406nSXA2FIvij+/8CUf2NW3
+gCmDIyUNTVzPmKSK+14Tflit2Z3g8CoSUt/fVsj/jl8WtAXS+Jr3ypPB2yK5/YnZFM2NDkz6bky
CGSgAPsWBHnGFhlEoleN1Ptbl0oGZRuGLNGkVWD7ATrk9MxdMmT+cdCWkZdq2XOXQVMXgelxR8J6
sCkIkfcOZid2Lw0M5iSRi9OGzB4nylPlv5e+tr1NO4T62NJCWuexkS8Z15nacZuZs0YCoQxa5UJa
luIeD3MYsKnUJpC7w3899BojM2ldd/bBIddUPcVNyMltBKHOl9FiAnp9qQ4kq/HbLo6NEw0aQJQh
DSNXZbL0L9mk1PstJmCQfwfex/0pW2qFnc0pmSKBKwXu+DP/cBe3bJyDAq/p54Rgbhd4k3aYlGet
omZvbp0VPYEkhNF+DXifqrl+90FgCuugFFLcPpyy/DVWLvpikRONb/KDZFlHKr/wzDF+RS9a+QbE
Z/+tLTya1ON9VcL1Rjb5wnLKNIZ40eHTshv93SGvVJhEvXYSFZ7dTc/IcvuYQDkwQB2v64fS9o9u
VbbwRGaMy+3nquemSMEJWOZUToszgW/awRgeaN6Fq8wRGcn+rdC06DZbl8uJWRMhCvJOjYHpI1tg
QLIxJBhJs7UKsEWnKcsl9fXBjya1IABGpCHwz4oCRiyjPALTHcn+fEoBwp6PymJj8SzAphi+RAOY
Ozh8mT24mCVZWCMVYtDbpCGFILbeTg396QE358tMSvycxb/3UWOX6ymsi4QZhsh8dzgifNEyN930
G8DBJ7y/ia5sc4KdQR8wkVAFui0gfjCxMnl095cAyeh+09xPud91OwPBLxhNDZnN3pa8zTeCZpIB
aXS52nbH62uhUBqjDAkruvZxvBPSix7H4iy/+KKQw17g+VoC1Tfky5BW5XChl5V8dLXHcanA61wo
egyrXmMPOxlfRJZmJ2A6KpQ9YKM4EmPEL73xKJr1gABss5ewOulVkcN43Xzher+8gr/1Ei3fn+xt
29O1kYLHW79GdWptKNZNyxUGFEfyhTeJ38FRTrxO54WloSNcDKAtLoP7ZZDjP1BcFh6vEshFOrkt
zoxCcbXK1DlkJOXxUNRggpQf3U562MsIIWL8Vxdu4nR/1RpEZ+WdAlZKaM4q6rptNNQ4nXyZ0iMU
B5YXR4nR4uj3XBy5EgOIejbLfheD4DXbfZrTrPPkiSjFzsKuTohmhL5nx6ynA0vnzuaG5UUtqjpb
m1zuwn+Wpu4z9+4aIm+7HXWNw5t9bpwR+BpeGu5STFYSM1VJEXRZUW5pVSkOwAIGXc6vGlWXWoWv
Be1a85RUwNL7J/y6hq+Caw7orVzST4k+QhV26fS89mMBArBwzLtdXYaETAkRLBHflXw5YvUrM6Du
K9sicWMk8ktZnvblWEw+4tb71I3C4bgAlvuO//QkXx1t2jdu00yCvy2Wpnii9fvOD20bSgRbCRKh
JTSEMM1GKD+nJvb91gZ4GmggHvxUiow7/WHVR44ikQRR8PchHcCfvSUgoYIAColdTQ6ewADCkoDP
lX3M2Ws3noSOhmlOTzp79y8xFJcLg275iHFRX0Q8A75jCPgoxxu/iA1+kLHlsO12BkWkNyHJvX1y
VVnGxzS8lOAtcFNh0ZNiPtkKSdgQGcS8UJpYCWYqAIsAHJPPVaOjTFRLURgCZ0bYWfQy9FryoDFu
wdEHUM1HjafGaxGVM6Q6QGvXaSA0JEbSbZBT7RNWJEcDrMocyHwbLfIpnEEzpgXwt2NQse8RpYR7
mcSGgUltVTtwxhw0EqxJfmPZXF20LUi9lOujQlk1y+E9eNVif7N+Q+6x1Mr/rpRnvbFxPCpF9xSU
qQ6hXQJ2VlvhyGSaGlcxzaVd3Hfu5KKO1DgJNx5TjVW2XUgTJ1+0JYGedD4xOScOfWsGIHlumyI+
HpM7TgWFg2QAG4E5NctuUwGwOSmdxFylizb3oscbsF7e5mq4yHtoNbFX8Rgdw7XNEpfGFVcT2U6r
p3BJQod5AdLn3gdcIcsUND81rl9WXnK809/GnpqDQBZ1HTrDiLGu/9uDzb30A2xIOx5/Zf5AB9Me
XjoHUcaESy2jbzWgGDduDd4arCQ5fRA44jejbULM+v6AUAJ0tRyhCbe5tGkfdBtn42FXStmlv/ZT
Z/AgJ+kCbzLrWxOOXpBJmTvt4vZqBtlZu6NulVdhkJ6ZA2RqucOx0NIkoF76lYk/si/HJ5ldEAsm
Hcoajb0o0qPHS2E5T0md5Q2nb8IHwB5cgtmYTh3eaN1gIUHlnxtEeWFDkMAigGlUtI8JLcA6p4sL
XDA0wWbnymKdrWAAewnRVSVGp4dlxu7K7WBGZB32isjhS0FAwpVekwBGOXweuhmFcLbFIg2w7NX6
5Ebq+mQOlBJBCm3HyyB5XvUfik6J/XSgoi8UxQOa4kQCz6Q+dLm322736PHurPuOdKUksridoRxF
GnrgJPsM3+y+eLVdiRXpXPYelZPW6/MsPUFvcqohv4o2GfpWCjX8GscKk92eCgVlYqPw6eyCU7Qu
+Fyf4qh2d0LT4HFZ5katzqaKzUQieUYIlCu5b8kz28ICUVLKV1UQ9qpUtyIAsoxvF0r9ZzQSi6yZ
mJ0JrP+60cR9gSTc0reApWNqr1yQcH4Ck/MakEOCCxY7k5Vv/WuYQMX/KnNxk6A1Uf9KVSHVigFj
NHy66UEeqCr+pOYR1nQTR1U0jAbTeeF0jbn88fru/htiMlu5BmzQXcabae2Gbuu+MQW7CS0F9x2x
kP0oDNwzgyknGB+RN9+2A+qPwmjWYb5wRzv+DgDLWEcLVwa6Ef06btDmH/vbcEmE844zqGI1duzs
WXzCYSx6Tgbg7gVO36QyyASbb6iVqFUHw41hOqSv6IQNIqnKry1Niz8Q2xBgql6yjtydOz5RamNb
L/aPaQpxFGkcTnqmWJFAp3p9Ss5LstUz+LxK5rwqmxk93e8fIweZEwM5CbRA2wtEavkS7S1Bcra0
gr0Of/dALMbLCosLqKUq4i7yBpC0QCd8izV7Q4Ryw5GZtlCS+ilRVyPHOYr9Mq/CQpmjfP/2MhGG
dTGOSfIZYndn5eazlSAhGLYnfhbCWVj6H9OK3RmhHXT1I2I8NcCSJ6XsCsXai3Mg9oYq97cKc9yZ
yd+RRcwaBFUG9WF5iRx9/PpdOkzwFTWb8aCcKpVIlR3UMOXY5fbtBq3totTzk/Edmliq7rCXbzMx
gyoBeRpqWBY/8CO2V+InP5z+1ZChnqXDBL2UK8mcvYPqXwQM0I06Wm61Fa7ouEY0F3TwB7ri85s7
xlyQo99n3kwqc3AskvZTmLYnu63AyV8NdWhxdTBVy6kAWrT/2rVqeuyL4ZssY0E2n5CsLv72l/Uy
EP1DhyctnM//OtyTXszivbRwzCoS6TsP8mScrcyuU2sCtBp1V/QejnJcgewNCEQBFnXYpaQTHJ5m
SRLTJfUpkL+YIqwc+gZqqvkyrIXmsJQopIMkqjRhWtTLHII/dyNOC0Lr9FJHuFKzwAeXBm3/IMZ0
MfZbg2NYbKrESDBBUpdYT6XH5kCc/b0IXRA3HsAH4wd2QtoCmPuz91OeGA46U9wpZIKhx8U9SXUn
t/ux72y/fU91nhkZLUIjhCkQNQDBqyxI8YqHlClIm1kf6Bgnw15JLq1BykNIv6cAwnuxeHiDb/oT
Wo0aYJURTtFNQ71ICs3R0k5KYQ82Ve3wqYHT6CA9jrZk8/5XSS2ox+Mk0qf6AYAvFEVBbiTDE/+X
VSC0/hsS0nWYW73flhHk7MV/j5LMMc8/M+7EZh9uzNWkw4JhJ0gxHLjANHX0u7R9qrCIpfny4Mus
iC0ug0XBwVuSe4TSx7SQB3ay9XqsOjawcnsaKsrmJyvAy1qXNMi7YPt2yVsEGGf/u6HMdwQYcur2
ea1dYPeJhGsrdXMI/bb6HeKlml1f2bVs7JzG5U6+16vhPsqyPBt85clnXKrWQCNtX4ZAja8m5zW9
4e08mBF+gHreVTn5If6gwv3+Xl/WRLSryYWHsyi+42fYtHI2kXLfhZcgc87u0RhEWcN7ya9On5oL
mxI8A9fvisb+5HNbcD71noklfqqBIBKbdRNYWl6KndUMaN5/XI4FjJvUShCCaYMIJxG+0ZrTVHaz
9fXcKms7PER+lSmcRb/0S9fXKBRzyGwifjLYkW+pWMiCGjR7KlKlyXDWDaWMdA3+JrTloxPFWXQS
WlgFhOuRPt7DQw8EgJfZ0Cjigw3x7D59W1orvqlVOeK6xGTLdJViBrBjyWM1nvj+LyuYxTan5asO
7zAyhy4DBSI7r7gZVi/+nkULx8x6iitfrmi8KFvaV9C5qIPN2hQKAjM+gmclzES5g7rYXnLU9D/g
+jb9mjgY9gpf2inW8ykphUn8Slfu8CMJN2SZz1BKhBZ9lR5qd/bGaHN/flWEEfZ1W21SGOQZCxjR
iQlPR/U2G6Rc/zVPhYTIS9nSbMQiwQj6YupMIr+P1PwbDWEZMLnIz7lLdspKENRfgRiXsJI03fWL
Tx8adQKBJYH1mSNyhSyXCK8GnS0kYc3Whsy7x32QDEbqXgKpSpmTurGFc2gEYHAUOZqev4/by9oX
mODwRf5xVcnl9XJi6CGua4vvTgV3XpRV8jTe9B5bIdm9yzdXoQDjtqB9bg9em9fHhSSLNBnWFDFl
t83T1zhxt0KYOG+bxsI7orjx33D7eheY96KbiK5KxuzKq7BCzVAxxV2V2mQ8EWfQLDlln0HL3YZ/
y0BVb2sMgfTuha3pZ84pvmhXyPOoveU/zRnkzSn4Ie4K46RAlDhwueISJMfMYzSx96qmpgpCh3Op
LG2L1wyvy4yMg56abAdLEDUk5vb1R1Gi0M6CE6OjQEoZgzGOkWWnuIz/s++tqmilEnkRRGNyjD9q
37GyNVKY0nw0qpYcD+XM+3aminqUhTGgXWBhC3rJlIfOR7p91LI52m5TDdp5iwvWjKUv/EN14KEQ
uUAJpqOU2+1AyQpcnnLTUUcxn2RbrV8LFu2Ahic3GZ6BLEJxj/LdKdOp9VEcak3OOM7yJEe+iH+g
G1KXBplW4s0CN/IDT40bY1DfSd1pW8YBWG4Mwo8Rp6pmoO5E31LSEOoXksmxd4bPAL7iyR1+YlCf
S9dV5xUfXwAD83bBXnUeTX3G62dNb+yVxASCK4GbkJZVVXElXApIZSCmsweSbLiiDBkewVnuQh4k
7sOB2kYT0unjPtvd8i9zRUj6qXLxuQtydPb9EUi7m72UlEMmLhHJxghY4biVNyaEhjZK/o1c4Vbg
12G+KU1wMdFEzVUXel5ta+Km+aDnPbHomFicwMeUiaSNhUEFZnoQ7KGzpewT3Xc2draOK4jUUN9N
P7LqxcFah6i22A3jQnQBmqN3It/TuZ6Tg28AB0135owNgd5chiijTC5zOLZwdNH3bZI1HwRBN3MT
PdtdtVofkr/X42XgYbO1fmQUMUrqXV6k0P54bTvSaGXR2o/bTHAHX9YBebuXu6JXoAZh7jvpJ9Mi
NGxnOzen4fj6JaRRGRcdnAb6Z/djO5euSL5FeM/aOn58xUOQPiuZZUlE0p4CZES7lL+iAodbjjxd
gIhnvJRcS/EtiFB4UBoBI1W8gNLGMS7VrsmaoiNnAWUGlN0mamu2QzVtwaOzT4clMjwab8TiCe3w
6uXojpYMg3TENIKUlp5DA6LRmNP5ArtbIn8pLuJef081MeJ6qm7zwTKz8cHB8AAP12TbI1hwjbP5
HOrS52oXRn8eoa/vivfeUTaSK/V668cME4tUERbZgdfCCmt3zW2AzkjtTh4GCu2YbbS0F2R6CJq0
MNZOBA1lNsAu1J3oGc5tjjXOe8rtsoCtAz9LoE7Am626RbpK9xaiUIb0W2SZegsw1uEFkXnJ66Cj
I7MiemPfcDaWNyjA030Kz/IQQwNglRiK1+FlhTib4Dktu0IGXAqGQYdj8PasuPMCCtzRTmoXCFXL
NkGIg3aqoHmC93YiF5WYiiW7gMAAvfQ+lvnV4jQ7oobeVj4Wq2o+bqwhok4b+laTJ1ouiVxdiKnr
SdrGe5x9hNP+lSzCI2Mh7wuWT3//gHMxQ5pI7JmXrjHbUWOCkD5pjI1HGWjYnNnLE7FemIRU687S
HcB/LsheidMV0Ju/GuhDs1WkIvIUjw093iKYe9u9Re/2wv/5g8rvusER9oAxDZvabEkRVFPm/t1Y
lIRi7woDPNxVmkNdUkUBuJgyYKxWLlmb6K+TP7HU0hJMxyeiGqREn5dXZKsnyNWajlxnFtjlC9GD
e43fNbyu+FM/CThvHHUe0KWb16gi/tcAJcDR4cBGdY0ItSKUQ+pAVzodpjxaOSCsRfjpP8v/LzPt
RifrpJjh8Q5j7QfKlhs4kIP2MRp52fFxhVW2IKhJmDNo7PvqUOygGEOioCMgJqB1lEnRyogAvr/Y
Fl8CstsGQlWgZOMH4gaiVtIJzJViliEsxPXz4xJ5CaAvyfE7uO0G+rCBNkvUcoTYQe1BdG5PWDVu
0AvBG/OzCwS8t1JpSnjLXNpWxYPthkxESPOFDsLiCXC5PHiBSsoHHiIdjl7cITFsFmr42OdBWsSW
0in1VjACFVXp2H98AlIQ5MFp/g7MZfkg2h9mcLZHSri0ztMj+Uv8YtfjeeoNiNp9XK8m2XJ54Qw9
GrimQbADhQo2UnTewuAJwtoMR4/0Gtzd69Pj9rKJ6RFC3TsiPieEHLqvBnjziK4tcv0+t2Eq2haI
zEC1m9PllsqRIWAxstHt83sbYnO7U5ZMaEGj8OELinczPNHKBH1bcrBbrXlcKbiKg0/VkUbW9XjY
0FQ7/1MVuaP47+fGC6tvt4gM022i9fPP425TRsPkDKmyc/+W4VMtvKY1T7OutvKYuzTKZ0BrRxiX
jTFVdq1vAqGqdlOxaUBi59Oxic4KNftyNt8HuF8b28twCbZIVRJbUPrt9RjUlrZiqf3wLpMoEVbY
lpGj5c9YWCLx22gRg+ML2OGMRuQmVRmOlALceKHMp6ZRsl/jCCHkoZetxfOV5JorjSBLtBprH1AY
xd2p7xl1lsqRlpLvJtxWT668AL7tfEWzDVPmEYhmXSo8hACeofyPM/gwrsxcm1eK4OlQ60jD0wM5
AayhJkGJvURNDA/WwKZI9I+Ryu/ssZJaWgYtVOg+ZfKnjqsZha+qjF9ABHOahW58dbO7t5GGCHvT
lZ43HGWGZ1Wm8WWNOax9EVdNfdoIPRkctVjfWr/1qfdigcsoKcR8dlHhJIfSSYBZH69tirIq0nEo
zL53VOQvUuzx5p+PPIpuNhGGWqfSux+mfV3pLI4zCh/pOjSEpPldTv+YpHEDmTdbUkFZYqzgKD1m
NBuHyg0tR+dvs9R9bF2ih4qpJfzT9iDHrq/SKOBrRashA2B36bZqD/xAUmRzp4iQE4duykEy6Bio
oLLhZ+yo9GQDvY/upIylQNL6Dy1UZHsl9SneWip/xjIBrIZncyY/HxDdlA3tjiNm+UuiVJzopaH/
pqmiOftQXdaVul7F4tgZUdP18V43FdiN6bh8LiFWwRwtwnvcs/ApY+7hZf8eVw2MDnTvjBiIidN6
vrrYVawHiIaazFtpkOR3McXKsTkgxm8r708CYFnfCUBF1ogZiu1yxNCM//6PRnY4kPW2GpC3QRda
z8LM+M1FlJGpfLryW2c00b1QbX+Y4Fyfon2dyB+5P+QOJBXmwEM+nmjNs1J+kjCND5oPkkc8dNPj
E7WUgJfTuw6eAWRd+3YJOk79OP2m7ahj0pdUQOUzFKRNwXUIbQOoe9ct+IuDVfVJiUk5CSlruYPV
o4/cNObnptldyfRla9AX26oVlwxoSoI/1Iw/MyLbSaMQ1kjkbexaJ5JQyyFwjJ88oqe2V2o1yr+D
Qfw0akRXjQMtrC1ilmorlc8X1kFXUJo1oqe7AXSLHsEWaK51Aci4/0vEG19/uf2v5DjkIOl8Uvl4
I4s/3vrCokFxBMn2nPNVJRGXsdy1/sEC08a8LAOLGI4AwGKVAWZspweQcsy8Ossay1YPKrwxrvae
gJMZ5mzgOt4ge+DCa3JsbC1tPfG8JFDgelcIGSiTtZ1q+vtI5lItGjvZYv8luSAVMrog2dOukLUP
k1TyyZetqJ6PTq6/0/wLmxJr1+kuImF55Hh8lm1JRXYsv8WT+uYoc9FAXsdUhvCs/d5VvD0jQdXP
b/VL+MFobmTAUaj0+51KPmuaN6eC5JZjyZ/afAn/VG0cKZxqPLm+UFtCtbHzFm8FI043zYTqoZ1V
S4b8RuV84iwULA5GOb4lKbo4WupyxO+dT+aZsu3k0Tg3/zXnDh9BbVKaJXfKmiZZ9W4PuSVMTqak
n3+lgW/rv/uh/EolT8r3U7wEqFL0BsTqvhgs4hBKPMWvM6hXKn2lNR7kfs1qHCJkrVi8TqZIQ7Sg
YBSPLlWSkhq4alvHX4mayJZQmYC1Jm9ZmvevwX4e28e5RDm3DWW7rQ8JGxlkJ1KqYzPBj70d+D06
w6sNHZ/by+eV8xCiyLf5aevHor5F63ZJc8jqAZdM5B6gEASrzsQeHs/gHpw12cPcCQIlBJcmbpnq
apSgLmWccV9mpDi6qsQsR898kG2SKkxo6LRoQnPhZPbkOrMVR9ktyI4Tvg4bC0KFHaZiWON1LHqg
OMtyZP4x04FoSy1jdH+KZ0hFlmqgdc7nb21cU1wiRiGPrJ2r5bLYANVxgrhx9IRFSzzqt5hTrc/+
tsSQP8hY46PJ9P5RInONlX0HW88gtLhl09mRHpkgCGVfgmT8cYgwJeYYHDSEz8IcXklmvashoiTJ
ihDDONxmOJacg7dG/HLihR1MU1STY2vOHaOHOdik2REazof2Cb+W6izLvgZFLsIyjR7FuDXqdil4
//kIpnRAVbexUCAuWb/gK7E7InMW6A9MEEDy3Bingim+86VoI1cJNChgqKv/BYLyPtttbIgin+VC
FggKJFxsjBoPAvofzHRBiq/zFV27Hjdnhsod+owjCZVXD5hE3aAt8DKTJpb+zo/OkemNY7xe5Z4W
yNq8dzvlhw3WpU4LF3jcq3o7DQ4jnwDQoQ587LNPFAhBuxLREhYrTlKd+RoU3oiz2lJtcHDq8dBS
g9lSTwKPCQFQF86RCxmq3kq8ODX+4QlcG28TBeH3uD/qFtKcj2WCRl07f8iNscjRFDd8Dej6moNW
L83gMsikuy3pMCc/mVlpCG47NcnBX41RbKMb1pPQFY1rTFI5XSxijZXofnKCNc+4AWJhw+zLxUS1
p7qB1VqQsxpmqJS0WB1tt1o9o867hEBRt9VMAOCkTopuJcWk6tj32VTKRuHkh1KUyPwUw5sJh2rm
gzTdx8BZvhBOIzL2BLulYDsQZzPKsjQSGpWAzk7RjdWU0mprUKcRYs/D4k7f4tlyo+V03tLeMSpT
4LRI/NEuO5i8/1GmeiRiGGdApH1hX9uOd6vm3yPEjXku1xgbVejg0zeiJD0nDK+dpF1td/fnLzQm
VvSScCZNxcagCHEbZ1o20zy6L6TyqrqL2vB6NGaTLfwTTsKF7ZfYOaOJZLcK4IGQO59kg/Yc3IZN
M2jCDxhZpk4UqxyZEfZbMo0dKt0Vs3bhvnozmhPbnd5J4KIwnxHD7JBpZyyEV86eZ6m06uVf/stG
YuNSyOhTxfwvcUrkOXRuRP4AOPuee4+vdwbanSD3xbhYv4sAYNPpTQ4q7VNe6lIiZQ6WPIF+O6at
M1leCK93yn17KXa9eZ4K5GX/Q9+BKBJFxdv9xf1y0HC9CWPsgxVYrU2L1aACU5W6eJQv0IwQXH2R
WU+9n6buEN13txGOjBtnIUxPu7D39dDv3jwAmwV3dnUQdLd2MqyH/gX4uAiSpUS59YOk0DGT5jVb
b/KXYb5kG58ZzhvfF3a4NmI6qYEtFNQAHqAaJo+AQ5SqxbJAS1vHyiqEsJFjhT50Wmmps694GciT
lURivj6gMUQdz6jdyR3T2sH2je5mmoYGhULD9sdPgWZugxL3Iv+tm3dTqSAOin7v85g7cCHW7WYS
FMeVlq60hVoZT+umLIudsOV+d1Eu8myyRRM31T2kyD3Ox5jWGDx25ulxTk+dw/Ft5aOkdnN2uTmV
Dzd2S+Y/YaNsjzg3qLWA2fRg9xTYWcGwyN6I0fUj3pRfVcMxHcfdvjjN2oMPfjgM1SEkpoI0CHPM
VEF5LEyz7SZZfxvGP/Qr2YMkh5V+5a3T0+KMSIVTtul5BAWUHt1D7BFgrPL0lA27rOOJBm/5oX2T
IANTAopoh6BuamQ9Sk7wlXi1yE0a/8fjkw+4JMv78n2VGg/ILcISJ+qd3MzJPl1zKI0NpyC3tiMX
Z6+GIpUAszFhwK62nSOmZ8Pg4uL+P6MrS1BfW9W3YhTvVlljlziQXwogUgdAJSgWYYsH8qRrALNb
aFT861F6nAEC8kuYNkG0EwSZ4Dvff8nknGGdf0NM6TolPqGTrg8dOGH0E3sRir/qWKxoq67hjJQQ
Ni2522b4raqmvrgBAa0QoPWe5dL+F7JnvQU3P5KkRQUIYRssoxb1/h+g9Iq8ZJTitrgSNazlMobV
ZBpKN6blm9YjhThh8OJYDGXpEwuLHD+8LT5cqwdp9ZxVVWKjeWTHxpKUS7BDKKhbaehabv+Rk263
laJLWc18Q9t0QzNtBm9Vmxpk5M6EIifvR4lF5Ey3Ar6AZ9W1GazpYbpcBi4j0r7mjaX9JzhWJfED
0EqIafAgF6T1OdryCeH0rGRihc6b6CezEqKf0ylzJE7MHr8hdwpVC6qS7UVEw4FrMwzo+wwHBAlt
v0YdO6vl8IW5tpBTHitpROf8pP2JdRingPd7bmYLfS+vlFrSL7fFmgl6b96KdQcOjBrC8ZTrdE1J
j8O9nKHwSftCBpw/bmJUyrtJoxMxe0DKKfkwa7LxzEdYz95V8KzzGij1oZuNVdYD8ygnWAPGIsZg
SeKNMl9AYP5Zl7gArxttOFVQe47LwmLnuYz1inioWx5Jdyo2pVQ6/u+fx2Gw5Y+8lUPotI5eBuDs
xLEMPCM7EW51RA/6RlSkQf2xxZOwpqPhe4gqSt5PdzhE+T3lgo6niAicPFMCJMQ=
`protect end_protected
