XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��idj�c��)�VK�mL~�Օ�ܸ
�G��o��ҕ��W��dJ�H��U�Y�.Mk�Y5%��~�� m�U55Ǜ��y���E`�x:�������ߌ���G��R'Ü<�r�����Rx	��su�����y�X�����
�z�LM�����՘���3��-�z�UH��8���qxF{��z���w.��S*K���	�DlJ��U�RE��ǿi�g�AM4��5�\"�	��4�J��=ye�(
����J+��:6;E�ϽnI��T:.����沬�t��Rm�4�1�w��mTL���W8 �
���-�:�����5���(F�X��������Q�!�Gqjt~�@
��i��3��1�y�����/����"�IcW|5���Y<��)�xm.c�ܟ���Ҹ�l�z���q����s��G��U�������@����[��tՠ�#�I��ԟ�l���Q~�I��O1t����{�O_$� �����4���i��f������k�ZN/Cg���FlRЅ�aH2 �'7�\�bsޒ��%��\��	�Q��1��W��]�O�#�哇���q�8��D�=KD�H/�	�t�vAue5� �������׮+Q��8"%�Ҋ-*Oe�R����/¼F�����2��,�,��)�cb3a��|�y"�A��YGU���H����8���V=�LO��q���`��^�U)�۔T�C`1���p9<XlxVHYEB     389     180ƻ_����!�u x��v�d���))
[(���t}�'�A�[�_g��[��M'��������k����t̪�9�����V	'���Q4�|f�<0�l��բ�ǮI���[���=^x�߇M���uA��ZI��x�m���:�Ȱ� ,�-5�M�r0C���tj�j�� �|o���v~�Z����7�Ixh3�S>��� ?w�ܸ]:V��*ҵ�! C�C�f��Gv�q[�ĕ��#OknX'y��pU�}έ��Dt� ��3��#V���R����ШQ���pb+ |��߸�ĵ=&v55�q!n�(�l[�M$��f]ꡥp��1���y��!_� W�F���M���t�#$���4�w�k�\�qϑ����