��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����vp��:�h1ePŭ4!��%dD�1�v��3>�S'���6��Eccᶗ��@��S��mn�ϝ�B�p���}d��{��A\4��t�c��/�r7P�`/�ֱ��Կ���8�âHc���N�R��+�J���5���|4ӥ^�a��ung�M��ؠ�C�Zs�j������B���[3��Zښ�0r�0��'O<��>9f��$�Tt@"�f�I�$�	��Ƌ.z�^�N~�j���^�2e=�N�S0�[�=&2�a$�rS�3ai"'���lcGw0�@1BE��@J�G���a�.����z蔉���q�h*ȗ���ع�C�D�h8J�2�n�p���<�&`9ܯ��k*Mi��T��K��n�	�~���8͍��t�[�ɒ4_QNpN��E����-���e�H���yq�N����0�����Y��}~�xo!e���&�^�Y�ۿ�}mJwǽ1[p��7��h��G�l��Ŀ| ���s��[���}!�Yk#���F��ɚK�" ��Uʔ�����^�R�9Z�(��({͕��k�����'��T �%�kS� E��q���Y����џ%{��B�����]��1�v��m��,���,9F߯04�	�߹��9���2����U�A�v[Z����}\E�[����mg0��d�����;=y��D��q/F��c8�N��O����Y8�v�_R!��~.�~����3�O�a�yY��=f�k���&�5zPYd��5���-�����W���%K����k&�?�;��Dq��uD���ڞ,��2�A7�U����Qz�|�<@B�L��]��M��T��3�v]���Y?�3�?n-�#��?I;�lȞ�����8��"pop��a�,cS����A�m
�MmZ�uA�J\�MQ�F����6�ЁC�h�Y}'YP-I�^�Fչ'e|�1$a�/v=�iZ׾��3MH$#}P���
������w����Xq�hG]�&RcL��ex﹮���(Yih�/V�Ū��"N��cn_��$�&�[�h�41��XҺ��-���g��/��@5w5��|(D��T�
*H�Ȗ��T>�ֻ�h��;��������lH�����0�Ո�ѝMk�V�KDH��j�n�i�4��k��+�v���	h9�9L���P��#ZJM��S&8T@SfC�]_g�[� �b�AW�h'�Ѿ'��V�<?R�g�k��$ԛ$G˾��ªǉO���~Z2B��ء�S�"��eD!U�0��Tv�~[�"�T�[�S�{���,�Xw�RcĿ�m�7�~�ʃ�eG̢d{��f��
X���w���A��#ӐX��ܜ��Z18�)yɑ������uB]J���ȑeͽ��y24�/o�?�)�^K"w-�o��kaa�����6װd)ܻ�J�=mo��ʾj=��|R�C����1���/�=���Y`����!*')Ͼd�W	(/;<�������� ן�h�5�Z�f�@�{�A�;J��Qֶ���z/ˬX��U.{698/���׵�5�(��~'��</��HD���Ѭ�К��]z*[�8U��4*�9�e���=�
e��V�D T �Yu9���,8IP�H&����:�eI�C�jv�CW�l��%���=�>(�	��C�Ӓ�/��39y;D��m}������s�1צZ$-�0l�~eE�h䇹�o���!�O�������91�d�b�[|�/���2��8p��J1 c��Alr��y8q�Y�����Y�ے�P�#@�^'�8�q��Xj�ώ�:�1Ο��◭�������}9�"\t2�t��i~���.���c��� �����}/S�Ҩ���*>v8�K��Z��bJp��o� G�@/�\������ɧ�K�H�����q��a4{�h2�� ���-.%C�U��G��Y7^Y�X�n�"��Z��2����?d��8qT��T(���d��A�<��2�S7�5�ZA�{
9���X���	�Ι_��L\q�;�H|A�R3�.~�n/���"
]����~}�p0����� �/���h��h��R4�˻�����;J��}��4�L�S6��E]�	�$Gr���{�}������PP���j �W:�Q��'q�eZ��wmą�$�kIw���x(^	�2�>���T���;'e��^���wI(1e�~bw9U*_0�PT�.njs<mf�o�w5���W�^K��%v�������R:/��<L���NtV����Y;���K�8J�.�q�ŋZx�mv�=RȺ�BDS1�`㪉5��ۙ�� �}�s������"�Ym1�%����͚�v����eb�!g�s*Km��j���]Ȇ�zv�'f�3�{8��35��ҵVF���� ����!�<Kr�#�p�Y�w1��1��=,�N�JW��졀brP�b�*��)v=�Ξ8q|xM	>�l�1@����z��&g�/�4��ZǬӓ69��Z�:0�Z�IϪ��?x�xmV`�a�~a����Ø{;d��aG���:�	�[`�9(��%7	q�ܱ�pp��_D?�6$�(7 ���4�D��j.��Z�|�Nb�d�wԊūYGgSi7�sp���v'��>���!*��w�2��������5��zPz�l8���>�,�n�=����n��?���1e�G��c�L�L�T&�g��4t�)$�[^��0�O��Mը�o�h݁`Ǔ~�S~��"'T*�	�e!��K����K�4�c�Cv~��ID�ᔈ-�Ѭ�w �d��������<
x�il�vHU���2$׈?���^�㭅QY�d��y���7�PK���c~}Mv;ђp��K!��R���N��E{+�:�f��b4Q-�vip�c$�{��Tgf$��["K�R=�,��PD�T����j���� ._��C�\����r}u>?��+�I��Z�v��0U�[��QWơ��*b.�����.-,�\�S����2�z�t��ω�7(,��o��3����S�1���J��:�*�@��b-��(R'd9�ף8c�w��@���w��3:$�&�u
�m��x�6��O� a6��^y=����)�a��i�X�BDbú��"������pw	�P�Dq���\� ��!"�m�Ԑ?ja?��������~�R��U�ǝ{���O�/F�/��
sB|�~M���V�� ������W����֯�7�2$�]��:'�пd��-�2g���I��)�����\w�/�(�e�|�m�%�r)/����ׇ8�j�)x�q�O#�{iL�p���|���}j[��"4���9����V�ܷ��(�mn��k�?�t��̤P}-���V���m	�� @A��>��m������\я��A�xn o�֒`}LP���/μ<��8��iY�C"���2�0�*���?��hB�����e�bo/�y�/�iD�&ͧ�9��I Cd?�6Vo;�v�`�\��%ɡ-f���8E=1c�h���C��-�ZNU�x�G�`���i�&�%ڴ�)6L�XFM|�o��N�ˀ>W��˪���`��  L�x�y刌f�l�y��t��?�/~���.Q�"1�b����cV̖=�@�:VXY���DqE���۫H/#%�s3��e[n'�Q����}lx�8�=B��D�U�o=%w<�ھ~O��J�r݉?#��U9�#ni^�֝O��m$�fK>@�*�����~��-ّ��t�vT\�導jM��5�r��μ-x���vQ]�b��h1D��[:��c�߿�l⢶�/d)��}_K�q��E�k>����q���� ۾�����--bI�"!�}��z��.�7b�1O�[c: �E3�^q>�1˾5	~� ��/��:�k��s%�]S�9��uVu;�S�<QN����2�+�k66*���&��dE�P$��i%a�~�vJ�A��s7�E}�,l2V��̩RșH�$ܤ*i��m���p��tY�)��n��?���wܛ`ӊN���NH�zg�7�K�93;T�sz��~�l��&���H���V���|��RNs��s�E� "��?�߭�@SW��ԧ�������Y�\_f{K�r����A��c��Rl(@�V��K>!.^�xD��/+�S_�MX�Mƫš�Y��(+�bf�m�j\��
���B��C�@���#l["\����v�Ȱ6麥�`G��K�Po۾���ŭ�P�?��H9�bn���~4����
�ƅ�&�(���O��6���������Zۨ�s��jn��"� f�W�+>���iN���LU�E���醎2����k��A��"��
���irk�M�}����K�$��G�$Y�=�s��h��T4g����"`^@M�LI|�6�����P�3��M���r���i��w/<2:�'d��������X!Wx���xz~q�k��bUgZ�2����P!�S*-0�>8Q*x��ԢP.֤�����8��q��:�t��#
�:N����� SF	v�ñ ��z�X�����f���p��b�Q�e�i���₌�3�_ fg?�ہ\�V���H��h��D'�g�'�wL����6x>a�}mD��%��%�L6m�s�
��¨�SFl��5Nf(6p�9A,ҏ'���\���E"0�	�v^���g��������+�
'Gae���<�ӫ8e$gV`��T�k�{;����񋋚�O�9Sy��^p����_��[�FTx�W!��t��9��^��w���P��|;T�suU,�gAۦ���F�YX{:m<Z�)T���7H�'g6��k���-����_�r���]��3ȱ\2��E�8XD/�ǚ^�z���x.8��T���������"��D�܉�O����\4å#|D{)@+�ٔa3r�o�˘������1ge�*x��ۥ?m�R�������|�93©4����j"�P�)�K��.n�M�Ӑ��R1�ov�uA6
G�$�8O�,�5U�GkȎd4e��p#Q�Kb���-=BK�=��'=����"y��Χ8Hy�}@փ��\!=ts�!�F��Ai0� �����{'9`�-���nP|�Gŋ�_�R���Ӳ��<��B�M�<����Y^�t���M��j�5vlR=���~1�����_�qV�NX1�CM�6�e�oJH�ؽ���z���)�߃]<K����1)�­���{%ϣf&�����_�����v8A���Eg�N�ɦ���``0q\��K��[�gn��FVV����#��DeW520s4�HZ>����6��U�>�������@���<ͷV�O����� �b�axZ�}�� Z,�^�$��$�X�2ȷc����8CR �j]�o���s��5�є�����Y��'O5 Y�e�E-���_z��c/"p�^D�o�[/�h�eoT��dG�-B��n�C��R�)tȂ;et�3�s��^۰0�B:���6�R�)[�5��y[q��Q�r�IF��|���R~��J���Z�"��B�%�;��k��]���a�Lg�ud�8��ƫ �W�9Σej�%��X����]�`ֹ��]�,�r�!��;�w�WE&��@�a<I�#�hr���R�>Z��#Ⅼ��ڴZ�E(�le����<L��w>�NqCȑ7x��t�0�;����5}��1� �����H�)8I��W�K�9��7�qؚ�Cgf��pB���)6Ż��־-���9i#P1A*����$��wՆ%�R���\f��W��	v��z7�!L�a|��]�3�Vs�zmR8�tww��k>���"��0���������	�r^?�����^���ˍ�#���d��<��b�F�#�V�ΰ�����_�^�ϩآ���`�����c�{rF�5�Z�������/�?�,<V�?�>�V2K�o���|�̌�wvo���\��KǤ�|rV4g���K����S����x.�h�|�~���d<y��	�
U�7�4�9�k����{l.a9�x�W�O$�F�޻�1�z
O�b�2�|�mRooݭ��n�Ɉ�͗H�r��a::%�w�\���,�N�R��Q�eK;��[�.�^�ĄUPk�ϞY�1�V*jD_*׬9�;#��������k"%5�W'p��c:�l�ݽ�
b��.H�P�ܢZ� �\�8��Z�7�k�,h�B����4
�f]v��̢���=��m	�BZ��H&X1�7K��8�['6�]���X[��o	�;L5	��	qCǲ(�A����H6��������!� |A���懭4jr�R�O���0J
w�������MRP�Dĕ�U���%��K��^әy��t��1~V-Z@>���ug]��Ϻ�����{%u�kcْ�EH<�ڊVW]�-A�q��PN��V��?Ԭl����}�A�|��G2�W�>��r���Ͼqs��W��S12S%�$���<DK�3&�g	�c>J|�B��R��Ũ��.#e�3�*��љ�Pʐ�d�5g�eDD&�t]�/uk�[�+��L�z�=�pW�K)#Ü���*#y�K5�R���6�螰B�|�5���E8v�"R`��ߙC	����Ψl�(� �c�˷����OW��#��A-@��Ej.Y�q^�]��M���S��\]�4��l,�-}��n�è$�q�@��V}��il�Mϰ��0PE�-I=@�j�M��� �m��7ӭ��%���kщo2���uC�t$.�\�uMe�C>
�ջ��[��@GK���D)�	l����wQSGWQ*<6k�[)�4�s�����p0��O��/4�U�;ܒ��*�`�^�K���7�U�UX4v:�q����.�O�v@��Uw���9o���,	T��I�|�� ���d���0�[�aV��+�(w1E�M��fࡀ�
�y�Sf�)<���I�bE�3���{=�ƒ����'�˚j�������Ե]�tg��g��>��>V5�Np��t������V��
� >��o��4шp������|$�ʬL�:�GӖg%�] tu��j�T�I<��n�u�N�|��<��<	kFa�c%5�jq�����b6��y�~�}Uщ])���3ɍs��L��\!E�B�FD'�w���0_�?��Q� ��~zm�ǃƠ�{M�m� ��M���eR���+L���&O=>@�y��I�h^���ӓ� a
>m�͇�? �q�>Z�������Е�ş�jq.�Y��AC�����E��
v $c�&���W�k�Jᚯ)�PU�J�]��QK�;Q"�����bN��}��}����'
J��=��I�Nh7�Jd�قI	��$ʫ��;C/(��4mʟ��=�?����
�b�&��T�+�,�2dJ�=1�����5�9�i��!��q3��6��5�w��'�Yw! -a#r���7�^d~w�jzt){`+����/�gDWW�Ewtg����K֯�ʴ�\�^M6\��=�H�4;T _���T��柀�F�ы��q��0�?�n(?�NK��Lxl�����_Z��GVp��=p�'��d[Ѣ;���}�Gtm@�W@/�z�����>�u�2�ɮ���Uߘ����P��H5�Џ�~�bMф��Kuhi�	����d��oAں�����s��`�o�*�b��ش�w&F�HK�(�׌���+w����~���`R۴G�x4Ӡ+��\ad��SW
�I��x��`~@�^o�� < ��
��o���_(d tS0/�������n�G�@.��D�6��;$����F�p���q\\� g�1�yC�A����1�>��(��]��pCj�o��vf+Rͤ�kRZ��$l�c����\3�ET���)E���:��h��Hy)>�	$3h{u���_���*�S_AȽ챞-E)��)YM�N�h\�p���S��1Br��Y�UR�1���$U��d	�zd����!wgǽ����-Vl�U�.�� �L� ��s�8@���;y:�����+�+h�� z07��dTBTp���J9m��6z>Q:���ď��ՑF8��|`�D��V��
��Z���z��\Pu�ٙ��T��	q vt@E��Dk�ŷ�`v����N��k;��O��5�/Z|���w�/5|;��%��o-�$}��Fd�����K �9N�g��os�H� 3��t,��!�J3;�4��{� ��v��c�!��'�>�X���c�;�1��5�
/�wz_�|c�9�L"��F��+G�c3�ҿ�����O���8ArRС`:o���c���#�vm8\�[�"h�Vsifq�aך�E��3�.��=�$��Tqs;�L|��tP,g�YU�6��t+Kd��&)
�`&�j�����+��ME]�N����O��G�BM��ձ�#ӡ�D��t�T�V��<�󬊖C"��7O��菱��g��
���Yr�٘B�RK��|�F@�q%���s��>-�ܥV	(b"m�-3&�^8Zjb�������F����u�CW���O���6��&;Y����꯱� YM��\؜8;>�ĕ>A ��R΃@��0��p1�7�דn��f��f��X����h��(I�ӻU���� ��M�����Z|���j�����B��#���	��N���j�L�J�zfդǐ�J��X��%X,��l�鏨�Td���[�0D=���$g_��
軗�Lh��;��_�e
�A#���VH����]p���b(f#6^�[�"�橙��#�wh�:��WŽ=�^Ya{�ʸ~�����mA?/Ы��G��A�������`z8�\rYt���U���)A�-*%Hl\
QIp�M�ʅP�mP�%m���D4��<�Q,���r*�|u���A__hl�jK҈Lh}[��f��pJVXE*���F���}��ԁ��f{�z������ٷ��^�S�Nn3�,�� �����.�H~~�}���'m�P8��۝��>t�_,�|��wAE���bh���\NDY����E!����Gu�6�{��z�zH�ʯ����N����'؝~9�����-�h���0 �	�����K�Kl�˪A�M�?h���j�:�bM�빆Z5�D����bu������?�|���O����ѻ�B�-��0�M=��6lE���OE��lN���*̺^�v'�@�"U$�$6bxR�2W���x������U^vW���x�Η�2<���pW����Nw�t��jUc����3]D~���n�ѐ|�^���_����k��*u�ԃ<��ę¿ׁ;�ϞlJ��q��,��
>A�ʑ�ɂ7D�U؞̑���Q�É����k�=i>d`xu����w3�r�,�l��*Μ�FϹ��n��LF'��`�ٹ'!tO�?��33. (����Mz�҅A�E]�tXc�I����qlTU�Z	�������&�͡��ǰ�,d4��e�"Ǚ��iQG��v	}���h��$U�q���F'���ϩ��Gq����@0�]�)"�w6��Տ�k�X�g�1��!s�=������O�إ�d�@��;���x�c0s�hn뜍w���̨|��/�@�A'��d?��c��mMWy��`I՟
 �e���Xj�Ѕ��ؑ|�m��h}�]J�w�9�j=ڴ������N�U�>�m{�-��u�&@�Li��ޖ����b����_�5�}�P��9�3~22i����>V[1Z�͑�|,��q�#�B�]���N��w�Q���غ�`2����_��ݤ����(�#u��uzjV�R�-}�(�ؤ��j��_��Q]�+���~�єw��Qi�r;ҩ)�y�X�V82ۿU��7F�e$%k8����j�����ws"u����QY���H�gJ�l(1�]�$�>?��T	�u���OG�Q�Βp#��d'�~�_7�E�6Op\�^aR2Pܴ�	n����F�;��*�������UI���(Z�TVd&-��a��O��It2 ̍����×<�W'��.�JEY�3S�h	?M94%�:HQ�[�@s	��D��*�ӸA��tr���B��ݴ ��O��/2s��Q_󟨛]�3!{MP�.��4<C�S�L�SP;�UsQi��"<�yA�82K^��"v�Tvጅ��7迏$�LO*J�a�0����XZ��-�NfP��0����xߓ�(-�1�`�]�1�W��X���d?��gA���Y��[Y����RE>��?X�wȷ�R��=���` 
�o��"�c��w@2P�zC�\
|CG���E�*�d������U�� ��d+R�@۽��~4Mٯ�t?�����R�Z5�[6��y$5摁>���>%�/���xu�LT������[ԥ�}�NX��T���a�]�&���n�.��RݒĨ��4ա���� �,��U&*vka΄N�/�7���˘Eb�l R%�������:�|s�oͷy�T��m�����oB$�pY3>"��5���9��%$���y�*�azX.�8����+�U���%��'�P9���ܕ|Q�p�Kg��E�r�c�Q�Wԥ���OLU�y��In-%뙢��"��G�; )�=#� ���q)�x*�ܱL0��"�{� �64|
��lŁ�o�p��B�eP���E���jR_�@!r��=jB��}�u1M�A
}(�g�`%PgL'N0 x愾�L��MTUq2q�.���$�^�z���{��<�-�ˢ36���j����
�@�z��Z���y� z�;�Y� :*R���7�cr�ս7N
Cʱ��<�O��+@
�͕,;���j�?�5��G�!�SQc,�KM��_�X�DGy���M�5���E4 %$X����nC�CI� ���(qe�U�����U�ᙫn�V�d��P��C���'+�-A	��4�I�Wj|���r�P�	7le��8��{�Z�E�"<����!l
H�u��E���8DϚ�[�#+h:R�D�Lس����G����f����l�(�T���2�a�@{XC��̳����sg|�I3�-�3C=>̾U󇄫s�"-�8/�����i�rH.-(�a� TX�,FCuJ�*����y���W�8�]Ia��x�1hy�@r@|� ���cS��i2�����\�3���HV�_9Dg�; B�ke��{�z�"g�[U�y�P�^�j��R�'�07]�Ή�K����M����(AA�Mb��An~�|"�߅[-�H�+�p�$��,�W%<�#-�!%;Y�/1X����Z�fI���Fܘu��.�r0=�X[����Q���	��я0KΒ��>��!��J��V�1k��TN����9?��n O`k�b������8GK?K����6���X�z��ɾO�1�jf7Ӏ�3�'y��]1�ܖ1RS��P;����6�pV�,c%/�@�ØZ<�L��t)�AGv`h��֡�)|,i�j�V���`.E��W�g�z W:6�-�I`�٣�?|��!��3G!�驮�o������6�._��Q�:���-:�����Ц�3�Ƶ�}�Ե�����K���i�Dw��`�<SU���t ��"���mt^���''�]l�P�O|����UN�������}CHfX���j���!0��o)ee�k����̑�f�O%�s�e=�G靾 D����Zˤ����c!]��OZ+�f|�É���Ĝ����a��i<X�fR�/{Y������	8_^�Y�*u��._�Bғ8t'�-��f&��{�hQ^��g�����ɭ��q�@s9\��Qm0!���*c��R�^��<�#=�L^=�H{A[s ���b�X���H��hH�_s{=�ˉӸ����wB���CX�0Ky��!��w���/_Y5�^j|Ը�UP��Rdׂ=@����.z�Τ�)�~�Y��)����}��r���R=%itX�y�u#%ڼ$��bu�]�	i܌-�xŮ������JteL��N@3�J���B�/�L�@o��0IZ!�Y��W�δ] ��	�-&K ��%#x�[u)�:I���~��u�I��M<�fs6��$`����nAC���ܴZ馚,�������qf'��@_�y�������M	�-ѥ�|���A�6��':inEO����?�Nĺal̃�yb��\O�3*��@��CD��J�X�����C���l�~��e�	`����F����W){\�Z����!\�
=#�=��Rl��e��x�d	��;�'�i��䣞�AѮ�A$��/���O�ߚ���[P~s��3��RaV��T�e
�ϭ��k:^#���a>���Xq��#AH7<��QV �e�ԩ�jr�[WE�������Ը1to��=9��@3-`�T���樹KgI�|��|ʓ�e�[���|�Ƞ&��xߓ=�N8u^��ƴ����]���&P돀�Y�7��+D�����.��ٲX��C�"�7O{H �B������'X�]���aZB�T�s�����M�,�'*�*�
�k����a���_և�w�G���*����6� t~�� Fg�i��A&9�2�}��z�����p�U{Ml!�]l�����C�����o�1m'�olN����3>����-Р	���f�CѧY��jǐ��q]X�7r�W���۰���0a���W��P�� ���A�Y�ca>�1�E�y��@���� i��h|@Ot
��*��绋$�����dFڔ�2�\�ÿ!�$��AJ�ǝ,dcu���W5��2�
��j�:�E��"Y�)��C�g~�~��<3�X���u�2�-��WQtJ��q��`F��/��M�nϴ9x2d1���Ŕ*yk,�ql��:O����q��Z���2:
}������J�����>�d�ޒS��)?��Q��Ȭ`^3�M���淟��G~"��;ة�$��Vf���-F���{�$�����=w{E�%㸜��
�pã77%��ES+���&�R�;��RO(�TIt���Os�Х�D]�d*T��:"ؠ��Ҏ�,� �(�Ϡ1SZ��-;�4$��W��H&�2�_�=� 	;��ǅϟE��mǲ�RGCQwC����:�W?Z���4������dLz��9Cxj=\��"v�>䟍V��䵪����Ki���o���Ҁ&��o�s�rK%��x���^꘤�\U�J����Ⱦ�X�f�������g����u�.;8�Y��ݺ%$��vZ%��
Ѧ �%��*���®�X��dq��W�ϕ�(}bMvl���,��kBf��y�V+����ڕ�[�S��;�&�`�iR0'ς�W�B�a?�<�%���鳍M� �,�,pCx��ޞ�߈Ë��]2�ޢ�v��@0�9cb�-̀.Z��"�?A���b�}4cyQ�^��LWZ���Pnu��5�)�4��ꩁ����ב��ʯ�z4�^�\I�c=XcK���-}��N#w
ZhZX-�7��ɖ����C��p?LЕ$��ʮ�f����}�4����3D��:��"��j��7Fr�K0Y7w8M�)��u6�JjeoԿ���f#�_��/��a���+��J�E4J�>��X2I��iZ�?�^a�;ՅQ[�R/�CXoI+��4��	W�L���V޺��mqz��蘜��ؐ������m[��^4	fl�d"�qm]��U������͞S�S�#QhH���`5p�z�\��g#�1:&fQƍ�Kmj^r��2,����7x�IE.l�uK�����_>1S���.j.}�v/I�s�=�@�`�L�`Oy-'$*3����7�<�*L�d[H�k��s<$г���m���O1|r�HB����I+�Pa �B$K�e#FPnK�;�(W�+�3�� �x0�]?�
�vYx���{�"�U7th?t���Yp��d���;I��W�1K�צu��p&I;�N�ólP�ME_u
���G��=Ar�����R5^.� Q���?�<6�`3.7Q��ʎ�[������<�ǲ3�z����a�pG�WԝF=`Ɔ/M����f������hf��B~W��� zT�*JZ�d0��YW�e�5d��P�7��f�vϮ� ؘ>��$u�赳��Z�;�g��:Υ>�f90
S4�<�MC�O|{� �����ӵ��8�=���_�hHu�i⊪��H�(��z��:��+d+A�@�f%/�9�%D��x聾Ux����Xӑ��Lt�����U}��s/�����>�rG�c	��XjE�#��6g�VL�0�π��F����r���p�\�T�}tK����o���C����=5'��������L��h��4ܜ�"GH)(���-i��Ï�\b	��FT_��^����98�8�f r�/��	R�S���=�pVJeL��&��%�f�����y���3�{���,���-O������zڀJ�y��`8�J����7��8�^��=�B* �Y�\�>
zN�kT��M�S�fʁ�v�vy�E[L�g����]v��tj�7��2�]��E5s��I,��Ķ�Eŉ^�4�hTj4VD ��ر+�7 �V��2*`�yύ���<:��`t�"�5�J�8=�Ԁ�_G����8�� �4�����<8V�����mk`��đ4��h(�3
��[��d�P��|gi���{y�D�Q�jZ/a��'e~ ��܀������S���c�_�;��Ou6)(a9�W�?c�~o�q,8>	Ң��*[J�^ �C�݋nų6o���N7��d�H�h��r8��%����K��l�0��P��ct~pO��yJ�� �K9>nI�|��Z���<[�6ܛ�8�`���}-����%cv����PE���C�>x��]��{�񇑴hc�9�i%�t'�����b:ﮰt8���bY���UG����j\0آ�p�6z7c�gj8��i�С!�U�FJYL<�����[�Ӌ�����ɧȪ?B�E�*�);�(jS��t�.�^;rM:��aB�JCf��Kɛ��rgn8+V۰ˏ�ټfT8�:��r�t���|KH��U!=ȠO�R�P�ٌ��U���z�2�L��Q����yV�6x���9A��w���G8 n:�bw���3��H���W��$�z��z����2jDte&g�	"�k�H���٧���ڶ���A���͇J�ꪡ��������K�Z�s�M��ŧC���^����˒2A���P����2��)��A�D�}���-FMm���������
9U|!c�I��*�g��c�h!2��X�E�4F��:4x,M6�����I��6����{�$����>s���b7��\���pC�Wn�F#e�� �~]�ǩ
��0�>�ѫ>a/��"%D���
�mT��(����7�x�~2��փ�Z��v�@�W��vǅ���}��Q���MMjQ��L��M�2Ad�ׇw��*���O�E3���6��~�q+e1~VDf�/�`�<��'�� E�A� ����H���wR9�R�`F�`����q�B�aO�
��b����2eK����������9a��w��.W��F��T���`�:���8�?��ڀ�*�c����:��5A��#E=_�-���&��Z`�x�2�u�[���KL��_�A+��
*��Y�ۑQ@�N���x��:��W�<9�9)҈�U�.܊�o��> ����9��9�d�w���{Zǳ��S���������*�:�J����Af�
0Wk���F_JGx����l�ֽ�5�U��p=�h��ǿq>P3˩���ɰ�Hc�	�ւצ��Sϸ���(�mɴ1(�$�����&Fe��E�8��aJEOf�i�o������
b�1�����ʶ��1�ݽ6d����(?6��*,�+3� �A`,�`d�3B8���-i8#|�yHi��E/ܛ���=�i��k��� ��s9U�f��6"�ZPc/���g��)�t(�fӞ�u�4���5������;�#Z�g:m-*����E���)�ɗ��7����_��P���ih���1 g�~Nô�C�o�8�VɄB�KJl܉�Eűn�d�E�F�v�2b���?W�)���¤S�k7�<��p,�{P��[ϴ�KX��_$�n�|�re��2�U_#�����6H�U0}K��uL�
z��22t��J�NXYBjaE�/g�S9F�G����+i˰���.���Pb:י�����!fM��n�'���[qyp�k����ץ1�Bl���"A��57�O��yk�w��zE��%n��L�E���\%�wу���`H�Y7�s\��#����QH���!4����R[2�Ǻx�C '΂$��8'%\��3��\���hD~Yu���e�,~��U��Q�a[/4�բ�c"c�˵�(�4G�ԕrb�2*�
Brտ;,�W��B^��_\����sF�i6����~<{�T2���M��*@ݿl��CUD��ꎇi���e�ˤ���{pf�����k��E�@�QQ���\3����A�Щ�
�F*��	�9�K|m����sd�_��,�C����S"��y)40	�8�r�!y9.�Z����n$ͅ�IOp��x$��r�<��QXa�e��>��x���d���r[$:�_�$(fo�<�<�!QIPa���v'�&��&�h���xA��"�)��<�Dh|�Y�����������R.�	BFlq/ѻ4gya��o_ �N���]o},.�@ߨ�|y�ѡ��&�NT�£�`L�˝1��Y6�5j�đ�K+��X�A��0v��؊L�u�J�3�ԣS��u.:9��;�#�+�fב}����c���v�P�zx���Smh�u>�ss�q������\l*���9y��<��nBx��,4�w6���R��~<\� ��C�D�g!��]wDAW������%����kD���T��� ٸaీ4��l�7��翇n_���]Q(�7�V�f��7~�Sk*�G����MN�D��q���)�=�.����"�(X�9���@�%�?U�o���1�7�V����*J-�W�+ ����|�[uI�Q����c�uX$���{�����ٟ5`ܞ�G,jS��I��_�vu@�NR�E���.&�1�'�8z�l�%|���T��/9�:q�1����鲡�#�?��{@��7��e�<����ͤ����9�7�&�?i�}��J�`D�~F��1ܔ�zP<�����A�AFsxHb��{�"߆�����j�>6o2����3��.�gk��3g]̯	��Z{+e���xD6XAw�y:��P�!�V���������?�*�1qgկW�������)k���c!1<��r��OU��-�����s�S�������_��rVλY8~*�6��Lʗ%e�U;��2=�_e�lO~H��d�.HqПuF��4�?��0@�������}����v�^�#��D��z(Ŕ����9���Zz����t���X�8�b�\vMZ_�:"!�j�!�����Zs �t��������2b7�,�Il��!{TA�e���
����r�KJ�ֽ��3z����M=�F�"��q����g���U����0��g0��~��������݊��0e2�D�(5�/�)3$���K}jm�"�^K4腥7��1F|��Z�X-^��O>]K���t�3���?���*���u۫�G���/��ɝ�Vl��SHE9��F�$V���u�A�+�LS�� ��m��y`:��bb��*� ��d�<z�jx��GX�"ߝO-�3Ԯ�ĒT�ZF^X���1j&c�X!B���k['T��?�&���A�{C��=�_;,ϗ���~�qJm}_����ڐgTY���H#�� ��1P##	5
����N5�a��|�{�|�.PG��̍c�Rpi��\Ԝ��P:�m�Z0UJ'p����kF���Ĺ�$#Q�T�����qb��蟈^_m9?�e}�R�P\orkbd�Ʉ�ֱ?�G���[R�Ӑ��j�B ���S�HT�x�4����C�]��a�]j�ۃ�F�����jk��*fo ��aT��;�
H3m%�����p���3 ���Ă��Dc�]���D�2gݷ|���o|Q���Y�N�X��s+�aa��G��V=��QávS�e���k5���n�{���N�f��������@�Jl�Uʴ�U׶0��(����	�����_�=u��qi&���8|;�X���J��^y�_��1��))_�F$���#3TeY}(zǚ������" �<P"�Ŋ�J;�)��7*�d�.R(­�^ញ3�	(Ԑ0 �T��_H���������	�Δm���.Ni��.��4�=����8��;Rl��)4q�ǢAΝ�j�����ru�#r2�P�wڗ*��޾L�����;N���S��K)�(������������ZA����A&+�'A�׵��I��b)ck*'yP;�&A��o��!�D�r~���g��'�F-ѐ9�g@=�>7C�B���@6��*HA���9̓LC4�����s���7!��
�OK��I�����d|�/�&�H����(�F�oi>��z��Y.I6�d�����!y�{�˸KF�0�.O�l�y�u!�&�v���ݱ�{�'aT�Z����TK�<�;��~Qٸ��a�\7B�l�,�V۫~1���Ϻ��/���[�7�+}2�z"�Ħ���2v�]��S��e]�Dkų���KR4b��zM�R�Jc3ho0p�����[��.(��6�PR�2�`�T�����$Ò��� p���'Յ�����@�1��Uf��'�5�$|T��h�i��\k�y_{�:����m'�wk����}�k�}�vߗ�>ƫ����8t6�#��U������T�Hs���K�s�+o(G��m���P.�6���W��q���x�n�洪� �Jo��o;g�|�z�:)�J}o���u'蝉��qB�"1���n��|(��#�}	�O6NA	�7*L�<�鴚�<l��c����MK�iԐO����L(P\->���ꂈ�
N��cG
[�����e��킧)=�������2(ꎞ�������E�P�
�ӟU�?�/�SJ�5,87M����o����x+����(5�Y�
����U..�Ԝ&��hJAk���Ϳ+?'Az6�(ahF�Y2�@�P�~�J�W-�8l¦����	���je���i�(���	��Tl�ѡ�|�L"������ݮ�J���ͩ����5*���77��?sO��~2�g^a��=���K<LdZk�'a���J��H�^�V��6n����h2�]������kYz�
Ͽ�z�f�W��zf� ���A��S��4��ǤR�F9��<��EεU6��	�hc�r�H�׈���<�R�7�Dѯ�Of*4�@�>8��NP�g��ᗃ\ �cl�}X��a�|�;!՚-�v	���EB���	_�z3�jm�^����yz�cO�=}��9�D�8�ѐ�{�J˟!>޾���J��􃬖{�8�!]j�ŻO��Kݕ;�&Z
��:T'��uX�J�'έ)���] �Ʒ� ��c� �fT#�����1��.���jM~���b��A���퐄�yV�﨓�%�����S�e�::R��.E��3�4��x ���Zm�.<�L�[ k���z�s��(<#�mUh�O�|��z.�s�UC���P5>��'7WD�Ռ���Z|֢����P�N~'D,�QY�<B��rs�j�42���gK�Z�V��S\��%�U�G���M �n�\�Q玤?$C�7���s����3�tZL�ӿו�=i	��G��N%�f?�<G��"���F�o(��1b�D��ߡ~�z�P�08�Q>�Z�) &�JVb�����m�Ks��M@����I��W� �D����1P ��~R�ٴ��QU&��$l�khl�OӴQښ��f��he���u�>�t_ҡ��W���J-Z.p<�7@�C��#�c;�j�yi��#A�x?�+����y�T�%��*)+�G��9�u�hP��Y��B�)�TB�t�Џ�{�p���E�V�!g�s�1ږKd�C����_tJ�?�޼.�3I){�+�,ۄ�pʎ���lia�oN3U�3m�;C����aS�Q88d��~�D�3�҄T�D0�>����
SE�v�2���r[��s+�0\L��W��v6�PEj�j!W��n8�D��&v�g���������C��Ե��m���7�OoS�*��ͿDq��������E�,�*��CHN�7�N10��l�?f���=��z��0���M!��_�`k���*�o�3Q7a�&��<8��]�N7��]�*�KSL�΢z�]�}J62���D	��������L�qP�W����#䠬���v-�xyv�[R��*�D�m#q~���óx,E�~U�_ڕ��޺â 9/��u	Ť
�s����}��1ׄ#��oeG!mR�wS8`xK,0�D���l�9��}�0��Ckǹ�yN�k��3W;rCܶ�C֖�����eq�*ͻP��ws炴A�N��sѾ�{(�H�mn�CE<��(�$(!L�xO�1W��|��� ތ��̔���>�4��e0�w4]�&U�D5{��?j�L��;'8�㗹��L���s��B<IҸ$���c�5�^;����V#C5��Wz��hqA�]���λ���B��)����}b��n�B���D����d����T�`�~�;�|���Ȧ0Ћ����:Rٟe#��4ߔ#�BƝ�Е?m��wX�����&J�97�f�?���U��j���F��;	�B�͕0컧�Rpwʠ?��i~:)9�Tu�^�aֵG����q^D�.5	����lq�U�AJ�DSLY�c�\���Z����~��]D�,��Qm~H���IM꽘-���{��#�سI^6Oan��7 �<�R��h��Y	h)�"f.Q O߮N����MlDFaz��x��Zq�u��g�*����&7 ?y�ز�x3ѪR��"�V��P��CtW<7�r��کh�M�Hx�a�u��d/�ż� �� �_�b��r��&i�k��"wT#p1�X�Xi�/J����<1j���)L�I�ޟ\���q�ߑ���dgc~wV�wzx�i���s�C,��@�S��?�?n;~4׫ft�����;B�^uY���;�_�������HL�So���r\�D�Ć����RJk\��wSjg�	n$��s��w�\<&wA�(M��Qo�&�gGz�'�u�ٞd�hL��|4�����K���N�yjÿ�K7[c��eL�o��KQH�>�����ۘo��T ���(�Ga�@�N]�t���wd~.9˷�sWO�{i� ���T����M�E�p�+x�
���UI6O<k\:3fC�Yd}�jY�����3�C�,���g�=F��bjۧK\p������GI��.�?�\wE9�c�H!ܓ��v����u0��|m[=F��p��e�M���ޢr6��Z��$�gE?�[��D���>�}���#Fѩ�q&M��;Gu�ժY�q��'��u��K�NGp��
��Z��_G�F��e�����^I;DǼ�	t��:�K$�鲷��8%��2ȫރ�P��:^ͅ#�Y���Js�2��S�6`+<�3��E�ڭ15�y��4��4	��'~3lY��37{�% У��b\2�8>�9ɲ/��9�K.�;�9�C����b��~�j����z��=�\nL�=��ޱ7�G����'/=�~�]�P];)�G\K��'�D�;�W������Gp:z %����Ң	����s�-����(m6��r�۱a9�.�׫�2 ��2|8��AJD��,k,��uci�ri!{}��^D�(\�@�1��U='�RK�n¾�r[���'>�.ZM��6	�A�[����\q����B��v��=Nq��uf��	-�n�0�yV��:�� ��+$/A�?�x��=tppW&����3�>`��� �Ԃ��^��}
6Q��"W�F,�m�mi6�a���_y�#��.��n�=T��'�x]N�o���@B��I��9��:�yӳ�E=� ���l�$�)m�4)�Kz�H��5��<&G�������;j�$w h����Z��Z���װ��*����"ю����LE�(pa
�D;��su">ac�κv=�S��B-���=�
�����T7�b�I�U0M�uѹ^���,$���Ѵ>kV�hR�Jl�)��J�{ki��Md��!N��o�����w�+��+�:��a����cI� >ʸ_��H,��S�6x�ܱ��/����֑9}Kh6�6j�E�,Z9������S���3��O8$Ў��ő����ÕŊϥ�Ш4з�3�Й�Xv e�6��c�����80{������7i�n  �\���7�j1ؔ����՛�V��W�ӵ��ށZaN�
�<��Qߕ�םG�#"y�=.�r�= ��m�U� L|MB
"���{����9�P����������nnK�}�[䐱_;����͂:&mB'4���$�U����t���ՋLzOzRեCT���{�˱��`�U}\L!av��ąv!CM��v�EM�!��Y&��"KZ����r�1��M������U#��,W��&¿K�#�t�`�kּ����e7W����ع��2� ��aB�[8N�4����u�W����|g�d�%��m�tf�������ï�e����)�i�]-z�֨k�q�Zm `���6�u �$/��b�Q���6`��q�6{9_&���w��#��r�z�:r�[nοf?���6�e�/�(�T��KO��F�*o�p�\aw��%r�^vDKq�� 1*���� �����R0�]��L�Cf��+<L��~!��ב��)y��� �&��vc�|Sv���t��P������n#�ET�UQ�gc���²)�2A���u����B��E�l�]'��۴z� �K� u�H�I�3��gȗ��wK��5B�F������ �}k������^Z�4���M�4^=ט��$����sl>���Q�T�镨[ܝ�p�'�ؘ��m��S���Π�+l�VI{�0*%��~�����u��G�c��-^�4,�?�Y��ljCYj�~��aL�Cw���w-��>���56@�R{������=\8������ٚ��)���+��@A�=$�S�E6ŭ#;>NP�P㘬TD8�����m;����L�6�
}ٍa7�B�,�]���"N�FE�x�&z����f3�~Ǭm^e��SK���D�o6��,�����H��Uq8p1�}0*�m�����#�{M%Y���\�k~��˓dvnX�Okt�!Ѥ�!��R��g�z������v!���fI� �Ǒo
3g�F��uM��d�w3������|=��F;��������V���;�����yr���n�J�ݱ!�&)�m��!�� �R���/�� N� �f�+P�P,���v�ei����t!4��^�՗a��Flgnqe2�߲�DU���(�s��~!8{�4D'��~�tP�\Gl��auP[�3�|Ƚ*_U��:P��k������H�/��]�w�I�WH��ՙ�Q��mzx^oͅ�Y����28P�1�	�/0l��� ��"�n~���Ӵ�e�cM��^v��f����i�(������\_�P�[B�wŖE����_�%p*N{{E�.\dGq�=[?;�*1A�1Y�9n�����!����6 �,���Ci�N6S�t;���ৢKG�,]�0-��7������V��n���d�Ӌ};8WL1 ��5�*�Qv՘Y��s"�x��d�T��u|R�p i��Ez��d�F��b��Rz�}ŬSduGҖ5����Zh	�Y^�]	�%ųLZ��@��F�15�q��6 G�v|����ᅐ^u����^o/HF-�����o�v���-�O���qI���B�'Dh(_u�r���/����k�<�O�>Hy������ɜ���_�,EG��c�����	�@$��߇|uL�"@|�m���L�늭ѢϺv���Z�!�v�.딚�}$J�۲!��k�^�����)~��7tbA��<n��W=4>mUcse}�(��TQxH�	n�7o��Ǭb������j��Z��4e�`\q7�Z���Ә����`c�%2nn]jM���>�1�N@��U�4f����2Á��H6��`<�*�Ƭuͪ~3�(^�T ������C�,�Ƃ���ɮ�EyG�9���@Y ��s��=ؠwv����(��L�����޺F&X����)8�%pr|<v���gk-ޕNH�'\�v�M����a~�|�i�M8�j�E��U����A;�WtWU��ʵ��72wﱱ�UJߚr��FE�d��]t�8y/͎I����޳���5 Lmu�t���q��"^��r�[Ռ��U�M"B�Gǎ�9��8�}��#~J���ʴ|O��blu�����0��h�ַ0{~0�yD����^[h�}�1R���+2`'��kq��sI�.���n����ᐙ���z��_/��Eͱ���./��#*�Ҩ�0r[}�����O���]��Es
