`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
ayTnq/xx1lqhwjrV+/SgJmZys93zGJmGDQEUcauywuUX1PCMq7ftloUHsKNWB3ckjjS9oQwYR/5e
mH/agoUozKRIq+q6JJ2CoRMPSw/67nJbqtnUEbFMh/u6dKtvlt4ylrjtWu+OPqNb6ii6i/5yMAtO
0G7KAlLSfmRj0p3YpVGtA6pr5X6eoZdat1v8IfB8QFWFp5Aso74zJcriFl3thzo8k4yShpe4qPob
aw80x12j25MQbue+h+VJnRZ7blZsnYPLDaG/y01nXWyzTGMZ/zmdGxco9CkUpgEWVyvKByQ4OcP6
7CcHXZfmguPr+ba7hS/+e0ilTJy+oZQgFBriTA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="C//hDXnGTj/gTyW4pf5yIwRrRa7fQ5pOPaVXw9msxFU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
5U6seKi31XdGpB83lRNY4Qa5ExFsET9hOsGg+LG2qZ4tbwPCmGfe53xHk4YOourLxeixSaoYL/xU
gGonK9cHtGiH74NlhioqQFBIcOsrHHHo9bsNR/E/Kgzu7KvtyyPuPd8q07g1KOr9xPfl11hvCdQI
63lNCTmy/3+sePG+EcG73Y7aRMWStCkXo5P/mtodJ1UcmIj75eZoXWeWRGVcTcc1RqqYLWUJSyhc
HjGF37GN7mkCtzRU3eZIHESMuV2qWMYlPwr1qsdIeWbAceWBrnlvpUnmmqz/bbRwbDaFPWwgjXpF
NDISCMscS/msJdF8hPBGa9UyISgkH8J07kAjVgd24/FzsgMKEN/f8QXOyibDMsRnmkfu8Pt2OkhN
PneGjo43G5/fTBqSsgYWxqARy3iwcSjaa5uevK6RMd9Jtj2MxxsqQGc5rTye55RetQmr5EZ45Q2d
Typ5lBLuH04wZWyVePgu3kJio4vR4iQioJ6vtjwU+Enhu+ns2XwwvjcNgla1dCqzIduhO9u0ZIYG
n0HUffngjXbinzu+Hc6wQELvYY1x3o3j6IQbRfmOrtvevMf4pdadsKli9+Np4Omm3NUmxfrT9wIe
ODQDIjC2CBpfHQe6IWUaNZL5vbdU/ctYEAP1HmdNVQm8rDZurQqe59bvzOgOzNbDoktvgnXggEQr
BFNWtGLkLwzOS30cGneP5kw5CCwydjPCtN18v5pEEgoSmU8baJpXEwG/COZfQTYHy4E+ogkG2E1P
i1GWODZTg588iGlaLcYGlscZ0eAf6dlPBRRFAmK2gehYmQYxM2bfziVpwTyTZYoJWv59D8yoM/90
bGVCQ3B7sGzd0vJ+EbE3uEaoPuD0aHFOq7G1bXTasONetIc3mAsUHMHYRhiWXJHE3CSQPani2Md3
y9o3GadomLBUIqOuTujtpqRpgfCow8SmJ8oaqrUvhBDIyPrWGntdGYWcU5I772eH7gYRKNTvrOg/
ZXJegbr+NLqC8RkRme1eePTkcJ5rDok0iZC8b83atUwgB3vjYDI2VmsuNYNaOKZ2R3BaIKU6qY8g
nAIJ2ojsojXLbNSEgzWjp7xWLwFeGEs1U9yV0DzXukeX3q+F2wAi5p4pp/Vu8npe6sjdrHXm7/bY
7LQ9phP+Gv1tmbUuIO0wUP0weFNFy/THQbW2zvCc1qDcDY3TthrP5dPL8Ieb88KlUsUBB0heZLTL
096Mel+AaF9w+1ioQHYN8lFIAL5Wt1cBr0UdC0qFv/XdSHPF6vAR1Wir+vOW4K5P4gFxEDprCCiN
QOZPYtD1+yJMXhPokVxaCQabtrS5xA6Bzd29Z4SfKu3fB4zCBZsIccze0OB7WOEFRX8PCAoY9fgp
xdVpNAFcnj9k3VSv71CFlP/dlMVFCW+RKij5Nw/QcpZyKmbd5O7wOW6GbUGEcZhRmHwTMlVGLz9m
XbBgSZFQCaP4M4a8HWybNzGtP8tXo6rgzQolqjGpW7rSbxybySKbYvBYD9+RVEQVuiAyGpvyzG4E
U3lvSFjbo4Fyy+Ku1YvcDYoexnNZPSKuZtT+qiGiBwDOO7WiXCX0s+xFDEnYo0e3CTmswdVU5qIf
owEFdyjqvnBueeTbVYTfhOIysAWL+heI203bTz95CYoEUj1tn8w3RqYfWG5t9plPwlbKaFRtmACe
Lz2hCGQDeZa8K7S+boERkfIoCh524Fn6TjSy/FuXTIMcHZSHlfcEIaCpu5YwwKNWAvt3PR9Blzz8
cAdx3v2DXzJsViBnyz5mdOThsnyy6oZH4liqIMDp69c9lSixr77wLOOdBr0wQaBgcz+h/Fbolj6t
H/OeHY4WFUZ5WPrKcBpBP0bvHOE7esBAozSOElg9lviLXO+qZhbYM6IQrcDKLhXnYNm+gqdvBPvA
tPSLP5PQ484fQhF1BFqR2pYmk8kOXOPCxrVu8sa3NBBgXxxt810YI0GFhT3CRnT+aSIboYUB1g0N
x0KHs9H/eiatmf560XgkYSQej6CDVPzsADAnG/fj1c6Jmb46/7MId2ES3LJO/Lx8tOLiTlIIv0Cc
5cZBy6XLtrjPrWhGIJ9lfawwmw2LcH1d9/lK991AFWU/DixNuvat53OzQKQ3LcQAeJeV1BxbKLSo
7/eUTKoew2GTKEVqJcXso147egjawpmHqrfEIvFCI3OrT/XJngH4x5TTrk1sXFu/357Lq7oW7RC7
7SKBjgBtb6x6RTLPRYKMh04Wmc+Zw7Rkz0IRwdrbwhW2597yTnlETRoRjbq3TtCUMOOyPL+AB5Bt
Hwf7KGprHNWx7WK8nNE1JiNh0fOTmX0oNuN8EaB+clFHs8snFjjO0j0eq/IuL2TJUS6jTPD78pbX
vwUhqMrhFdvfsPvmNho0K+fHdvdEgFDR/Zw7b4rA7um+9JGUb2j5k992WxImTQn55ru+2mEXMafw
TxlhupOjgqvYoAsQhCrUPPN0Oh8tYuEVlnzDv7hut/tU1vcwc2hNGX21FD3x7UJY+FLXt9PXOYrl
bxIBdg44rb3t/RqgY2qwSm4C3ipRIQgh+e5oJMp1xhBJB5NILfcU14TNPgWJoi0Zcdtdkq+1nF5i
j9NgegBUXom2rUWYgY7U4aHspahtjsTp8XNjdxdl3t+4A3UItlVXKZg13YmjcKWGKot5JHu+6Jzz
jXzJo9nIZqk6KGFL0wgngevHlTrIGPeQRY1U62eBvqfTK5QgLfiwhb3pbN+FofYgdbNeqUL50h+z
/1/dqIllzzHJtkgbYN5Ks0DPimIrWty99BL7lilVRGZMVi4oqODI0JzmS2ipNOpz52us+hSvoOdl
oOrbfPSBr4xHXQg/kcSDrtEF3DEgePyGT0d0beoQyIxjUwO7kTXH9o1MW7ifbRNGQSTKz9DqQCxz
a0iZyLmMT+ThJ5qzqJtLHdazM2IEW+l9rMb6FmngyZcvRpljc9TUVmKTKCbAb4n54eFYhc6POIcT
prnnujExLAxPSEcSViKsZBur8PFxv4mPiLXJojketPFHyIRLfQCmirMTFEqYu6oc6nInL7FxkthV
SMaOkZp8ci/M777f0yqUim1S6tDm7Z2Uq4Ce8uk2L+pVv8yGnoxeVSLUOyPLSA//yy/YbBX9AGFB
fok+APl799HKxbCgCZk8mNUPfBoUHi/QIzphy/halRbLi79VsM3i6hltDwXXYKaOCV0nGi+ym/oU
naaET5AatdBcDPpD8bU0+wCHORoKm90sqsuKtVAr1BkqWX2IGcYnWA2MARXuGzf6ZCQ0q+u+hzFT
BUn7foVSWYBrquBqm07ZWMlqVU6QrgmU8z8tcRankfQLDBkrNM81BXmcVnYTjIJ6t8M71UAcVU6/
0qoWaIVMSGwrfvcIlYLwZI+tcFBdEbRZ6qwnniG9t9RkiFYd+RE24j1/p9Y3xBSRI14qFTOsdrTn
v4dvgcOuPY9eL6awdw1oYpbkowlT4uqez7TJeE2G9Tp2BchaLXpAQHD2zjjIbx6LOgcM7gver504
GgJ5lPOp0BQDZkSky0sSjh+x77K0V6UJdUIWxVb0vbmtGrbjv6NFdmGAG9V8EcW/FGgdhrCgwb8t
GAgYcOUVjg4CU2shId3S5mwJiN6yuw2NekyUCGT/YUq0ximP9I3QakrXNtAspIyV2gyDTKNxJMWb
chswYoyJXxwbQouoV4zCiumuGHvGhjsOKcNnXQpzBWB1EV+lRhKw23TE4VnJhedFx/Qq+jbnF1nI
b6dspFDsneBAdCVfGA915NEooUh0AN33pCCp5sewbeLgN9L5rBAFTepXhkw57stpOSUB0yQanect
Ao45mUklCosaysY0AnwoyqD6c8Gln72HLCKSIOXXPyZgV8lmjtQSwoptrUdqVT93+CO8IUYOfySq
0NIMRc3UuJBJJ3Wf6exMOZGYHy0UJZsBIFd51FTHjEZgsAwT8b/fZ46SqVukK0+G9SC1gwU2pWfb
G6796UpniGI5ZLg6TCt95D9PBWDrvs8oqNSawizqwNIwPgVk3dhQBame6kULIV9Gjj0vm2ZjcMZg
6418hbRmxKp7IcswNYXmElGp0r4TsIN99BhlVj0N8wb5JcCpnSeAU+QW4idtE5eC7rUPbxLbL6H3
V+yl5vgdB3BZpLhPCT8WSySvpwUsYadDM2HVzaXo08fqDX95weyMTme1lygLT6tEoEpqieyxrefo
BuIoNE8eMm7MLmDeYlT4ZwhmyHR0rxNQxI08FJzIFbggb2Usx13G9TcikpHFeBBwW7ijFOpnzqPL
UzyYNW/9LAnlPeyN6aTYdmAc+GxNTe9BbJRHTiXOyUS/AjHf6RpMDPVtDZVZPPd7cMZ4ZbAJJuxx
/PtfJLnTI7qUfrccjb24/5APQIIvBwtyCIz/ZjLe5yJXtVBRMPgBitsVI/nb5p5sozNYfPa6Rw2a
/qQc5yyFNKx5UHvbQ1FV9+OmFLCmzoDRnxp2qtL2VXu7EGIhBJ24xQWzJO2RuNdciERfMeXRnGFB
5Lwq04RcWmnVKgeOUWQKKWkLqHLoBvoYwxaPpPVC8NDCOs7XnIkrFaDRd6J0OCWvnXBfaeVMT9gI
gNafoQEbEXoKUpOCF8+8zhtbnyzAqinGp9JQAhBKsLGVN03bx72vmzu5Fgb3TOH2vjnRLvVn4CjB
1PQaRFGjlNdsi8XhlSNnpz+QZ61AaYzbqROooZQs4ya15GiBywtZeWyHZr09cNoPlgnN33SZpD1S
tH4PPBOejVKKWrty4L4coAIgbt7qNX9YQgxDpLNglxH7yYgFBfrlj7JUFI0DkeZ7eBbhMaB3UjKx
sZ+DN//P8SpHaFDQkoRKmbBU3RdjzM5umaX/7aqOCjl+t4l03qeGwGhshKk//NlAiOA55bwcASJg
tteCizf5bO2mrAf2YJYL+QXR1gkTw2E72206AmbMPvCjkg8gw7FMZ4h/7BqckV6qFyQIglDdlXnf
o/yzEZotmIwJjly9DUwd4stAP7rIa0xNaZL9vMR6G1m6l1P+zuFF+wHMoWiPiBnyqGjmoch5VMDt
OG1x5cUHwc9iNWd3eu63yIvcEprnXBU0XY+8TvnBbvZI+juiaErYx/PmHIG6GWQkqO/2RJlqFrRT
a9tm4c5Yw+Oq5NcBTPtOtSwAhE+8
`protect end_protected
