`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
UEZH7PgNAQ2/HJij5N9ueuc3sOZsVQGiA8iKl05fRr1UfXbCiUXfXeCfTeJbElcCnnbbxZhBxZ/V
kLqKu2KZ7KB8aW8GQULKrLI7T/b6O8rtcceYvbPbp1LzSxR4F07MmoFxtLpq6sSQBb6XggyP8ux5
bea8inuHl8yfmkeFyDHpnZUxXn/byjvhy7BC48IUenkhf2RvcC3bKRxBCmjIPH2f9WOO1FyqFkRa
aR9AQhuBd9UnKkee5Tkt2Bk9CT0GnnByF3zdTSNHiemMqkGTkjaGDCJErGt7mw6DkGhxAu7IaVrB
v4Bz0/ZZaYe9icuSi31IUuoOJ/o0QK50teaBKA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="V7kSU/F6hVg8FnUp4P72qHa/HxGAoJpN0IB/0hOVWLU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
f7q6sr2Bj9cg3K8Ka9sW/reL+SlBj8ckpP8wRJQ3Pp4ovpORAI4wwEHkkMP82V8GNqQPJ9EOvPeE
h2MTv3eDp3GjHzLKy4DU4lQ3onr0ZZcSIp9yLGcCjxP98I/Fcfj5scp9VzaHUhbu+zamP0TvNJUD
Sp7SZ2tGGC+mmSGLCaC1L1Ksz+NotHZl5HHiv/uAL8ddoH3E67eVUCTHJeKprEDit10sfQf+183c
d/ovPlFl6FMr+qbQiawQoLXlgU7bPx3nwiYeAjj524N071yr5XUTrMqX+Oekjh/Q0JjCUgE+6zbP
8/3LTNKkyEIQowuMiTY+r1FRDBWRS33+Nbon3chdf0WivwSI2gJlNgFxPHsTRpJ+ioB0sTvPpeYz
/RyLAUGdG7JvKAyOUVRFVdg4bHcSCmEiijiGUfCDHCqHkltZFz4I9Y4wtOwbF06Fw75LjzqvVk8L
igR3ZxaFl8TgvJou2YYzIY/DgcL7kRCcUOD4dVjfsR7UaCArr7faJQ0zvbkHL+hG/A9d4i8dHSlJ
1uvLMYY/b/fDa0W8LqOYda16ugaqYN1DNdXPAYm4wauLJtlivSCLb6ih7jlGYm1tDSYogvE51r28
LxaTBNfAIGLwCxzvAFuAoRoJaHAyEEbPHN6MwScQACSnNGGvF8SQSvXHkqvVFdVB/80i8MpACUdO
ClUAtiL0dYeF6SEBzi/x49633VfQX/lq72ZeH93MNVM8YPceWIgeIR32+AAC1p6VcjVDMmztQWvN
04KwRFyULVnVYrD7maHFSI4Fn8u/zIJL1HMB9VleUzihi4GhM6/yZIIMZGKKxU3GlVA7s2I0NTBd
o59VgmBP3aaDCi3sI0Op1UTOho4fkLtseJrFpfdX52n3puwr+16toyJfQ7+8vignXgPvlrTRgiIs
VtcsmOlkDlKaJmG5/wV35kpupvz13W9T8J8RvdyOm/xZAoMLww69p7hjTYY00lFdgvhh0+I3Sb84
Ng8LmaMib6se68mTGZHps69qEkfEvsBsCWvPQjvBUl+tjBKs0uZtO4YAzE6dbYn6IZlilXFiFsEd
WaGAaNsbaOt9bwjPcq980/eb0V/vckhJEyZOD28LndWwLJfOnmk52CIxUTy2qb45DiNT728KuVMB
LGsYg3S4alb1nk5UkMBKhVSnt/i6fR7cF+1+D0+Y8wJMjtTQvTJ2A7a5LOTIOV45PeSYdEpV4NlG
N6jYs92liUUYSnhMRRIdRHLVeoWxxGvn/xb9tRtXwcZHVZSvvvs4EOwfXwCLvkdTrIQHHJLWviAM
FPuAQM6xi6Jb2odpbrjj7Qeixtf0XrMSz/Qf/T6hh+6x5/ezz1w/nXDZXSyDUQW5AwhE9JC0164q
xA1H4WmXgr80Eu7KI28Mo3PMccsLFSTRFX2bELKaD/LnSK+sIyoccORKTeuVikW3S62Fc6gkZQRG
IFd5q2tKryplohp3XKod5NFQU6WwWLWqjvU6vUBOtruLRq3jYR3/+gcqGZOi5DXFeHEMrMRrxIJb
7XnNadUJZP3jazHCYB2wPI8MEPKUAYYPQ5hLluSFEAGqImjJhuPUs/cL2yrSUuxIVKe6yoOpDsIP
7g1Vc50GQahk8ZskF/KDD/nonf4ywCoV3cIWGGH3SqZkmqNGSCLq/r9DBPo+v0hrJMuWEigREXUl
3E/YuA7RknSzz3CAKZ9t5PTVjJ60N8modvD1CGDzb3YTwD9/JlDr3r8nqPIqo7NzsFybmGmLZgRo
PNyWOIaFp1hk0LkCz8SZBLZxRH2EOJTPAylD0TxckE++sDzGYxdszhe7YV4Ux2Ru0V20YRbfxvCs
VGZJVzc0dj+IBwYISO9KCHIQQ855JFjTRe4mz+4IRYW/8cI6Z7jQLFzxIHn4iLCq10OP7Q52QcWT
Ppn8Q7aKw5Mysa2PuaqVbr5E7Acwmkx1tLypQysqDl+6o4SUIn9Wznudhn75+aGcqicQ6hdlGJEN
qepbC1/nEV53SCn9QSLH5sYScnS8CIKi4mCl1NK1OQYZ92bNnqLx+xDmah81/Su7w52YeiPm0De+
Sx+w4al5RSquiV8Mu/UpWhgmSBXMmPpoywLUq5CjKS7cGUIekpFtEbFvoriYuFTOHDsgUKAnztRl
diGRirOxVBXkdk9OK8IjsQif5chxum8kx1hYzhs5baH8mLre1BhFkUTq2imo2BgONzr9TnNgzdai
J37XWckZfE14fxr2ayXFg/wx0guwCxDHtcJ8o+uMEv8OoWMXi4TcmgViz0DvSBEGGWOqCjK/vGZ5
/mNeZ1yHM1CnjFBrg9fFntDIr/3u9rcWxJ7dtd7M2GC1jFB1sqQ0hH1XLPmvfYdbgNa6wmv4vzjB
Ssfa6bpyZ5xZabas/T0vjoE5haOW00R86rowkadwH9oxSwzZHg/Y8NSrz83iQYoHD6jqdKhgcEqx
jVkd1HXgKSLbUP0L/JwtJNvnzKjoDXfvlf3A9RquVJehgnkn3j9vJqb2pZvJ4m36HuAtQqvL32yw
AGDIK3GVadXBzRFh5MkiGSrgBkG1UH7PI8awVbjIzRxPO4xHfmaD3EwvBbBWLvVNKR+tvkqI2a6v
RY28bxvVHAg2u5iIiUlC9S5Gmmps92UHQsug0rxROxWuUemHZ3D1PiBBdt4eCNaHS3VadNuFlyXl
nIWOIcFm5x+PLWvkP8pWDbpp1WPkXawNBFhkdKba38t/224HpwxZmvVTL522dirgYLt4zerkM+Vu
xsrEiS0Kgqdcq6eUpeSFBDmbZxbnTkOP/bVKUf/Z55PJakgrSx9WMnVpYGiLaxb9IWn57oOn2L+D
qT4HZgXYgDyb18QLUkJhThRHF6t87jZ1s8qjNcf5D9iyOSU2WyaHDsqJQfQwrS0iVB6wh7lZYXrG
iqqVh+OG8bTbHfPYZAqkPxzM1nB15JYkpNURqPpZoNx9iKYv1IGC4y0InxbfHfJmS+NMKL4DBWzm
X3qweUMZQSqc6xe6hq8ZMf1WLR2BCBI39pvz68tCxO49aabk/gaZXdSTduRlNlp8exdFfqdlgAGB
rBg571jsXv9xZV+wKsisP80S15UbQy6Fs2YTdcsYFd/SnUVVg0xZy9ySmOVK7CyoASzZkCzJv372
MASkWpi/B9+JE3L3kX+iwIIGJ4Sx+2o+EPhKc7BgVmtnf2SA5Xf/7GYkTmwJ3Q9oKksQNkL/urtI
h4Iexe36gqQbFjAXXmvk7mn+5HiA4h/5pB6CjQhQdbS03oumfRm/pSVIw1i8yXCbKKUfmoTNb1S/
4IppIlPJ42ezcyzleR1Jt4KvIAXee60YA0t9kxIMvRC8v17IXtz0ltks0TgAJ1VIXZmQgQqkU1i8
YmVPVfjFgdO+rqKgGrYstr1YwuMLKznHXusf4H4lF/6fenGQTvWgxM/zQltcsOyII4SRTHJhlkea
cTpSJUlTxDLLH2K8kilqxhdHGcwzlg8GU7v5/RqUR6eTTXclcdKYEZBo9Zh65IWmcc5jwxb5HL58
g0b9sO9b0A1ho3b0EwSRwb8EQWN+yQA8cUTQL6MDoV6c0eh4EECL7j0gdYELBI9TvIZdzUMkVPcV
/BXxKccixso3gQJwb6BnGLO9Zl7ULtpUfzjMJncxJlF0qNhsktaaaH4sS5QbNpxsvxBQ17wLKunj
ieKFwXuB1WMqVL2ugBwOJup5l46ccIfWZkiUafeU9Bc/TL0OrpHcGgj/Oma6f08/qD/4fNxM9UeC
7MLx5ZnP8SFYKzMuanCdr9SPFZQBTLn57l8wCBcT5krIU6plKSeH5hUy4tEJGITR+CvIKcRI24q9
2TZ+LZs93DG91oS8IWyq9ONvMOp01vSJk7KaHArVKNsJzomQKpcZbwIy6a8u0fX/h4QvTKBKvRW1
Mr2kq6H+hqaOBqoNoQi2pqm2LMYenpM4U5C9Ulmztrlj1lYD/46OR9phOh4Na/3N1HcPWN39V/qh
w7FLBTVrl1ASLtbhOs+F7hxcUis0uhNP0WRAAWIy67YR88nxdE5cUjjcXU0yL1iz8UnBZVnjsKLM
xoy40hC6EKajyqdTUuyG1oUiz8dC9Q6UN7F9bEmgf4sA+B2HMBAHT/YWomM6E+tjH6GJZ6Y2cZFH
9dq1NSEr+WvWXcEEs4auLOBXBrGQIyDnYeRzm2kqJF7t+V6dRBlahErULCLMukDpB5a7LhJPEcMt
p0+5CXkjFRAdfCp2kTDPS65esDbdOiv0jH4Yf5yxtEha9an10ZofBJAjlV3oJow2h0fihal6BCAp
EiMDuNpFLkBDtUn00v36yVyAsXPDpbVJKZbFsd5AQf7TKFyGBh7rZf4eI+wbfvPoDBge1XhCDk/O
NFWfXaugTdiM4MaMX5C4dLyawnrVYKmM2zN2kMjoqoecvtI64javtr89sBGDLwU7GeaBPPVS4VPP
w+ThHS5A6J7IVQh0wTvL9tICVQFB580uR6bHwvxFjlfaPow8O0xdr7Hw/jSK9AzX/GQau45HvlHq
8CwomEoeNV7guuFr46XG/6AJxLn+wd6LjPP3FNmEqSK+4Kwg5YScLrmlQ6Sk3xCpbZnjwF9cOoAt
6EoV03pFrLNb3+y3wJ+j4jRTW5dp4LFO3RKm+lpFJzu5OeL4+ilBx6qPSIRlX9+erJCXoov3IGzk
Ln9GtF7B116wXWkQkASXCTK0F8Ldi3mXc6+ctfc1jKGE8LDnK/ZqyuojyJMBP1zApZcUoQG/Gs80
b3YzgiAhuV+mEKjFWq6dI4plm7yJlKrg9sl4oETHJcdgQ4vQvIQveldgRgBf6onlpicn1/rUZkmD
j7SJv9YDNAIP85Kzmxem3QlvVnvFzggrDvFU7268uYTjvfIAf986qd8tuXIJnZQMVz7tIv0I5R9y
jv3k/bWBltBv7NzCPER6Iui1Ng+5RqTYHnqbxWYAEZTYN8lGqXbG+0sAlGmtKdvSaYpTTkEDaytg
X6/JraDjZ2YIs/GwVDhvRuFclnJ3tm/ACetW2nB0acP7XsROFmP0il2ZC5lS+SMIm5T//kcZXwgE
ZggOeByR2VGvNWZd5EaFh54WLAMjZK1Gjtz9PYxVIaNedKou/lQPaKzhTR+0sIPpQ6Q60LqtoltO
30ZsCbdqCWNOJB3D0aQZthuDQvSB9VWGvz+Ov2iYhLg/V5FcAgYJQ50ThuEdGvBkbIBRvxCC1XzX
gYcGZJso+E9RzNp+5g4ojhyt9wYnz2dnd00y31AOKi6U4j5QUamh3CAz1+DL8xbLdxaAW5VI/cJl
0bmAKKiJksnNMKAc2QZR+kSwwXt/S+yaDDfwEUJMpHfz+XlGBvNF3kUJZBuSdlmVnPS9i8U00lS6
D3GVYRWQSRCH9zAZX3PjMNCnbJLenkFx0COsqrKwbzF9vQsaVg+SXnB7cXeDOYTcYAy1SqJyl5ML
Waq0jprH4JJJJ6oNfVzPA9nSsuc0O5tAF3D/SQqAGxNnQri7Mds5ksKZIk4h5r3r1ZqavISDbkKr
PsyAbFsmtyWlZcVamzDbX39AuSUDy25JMnbhOkVttqVCaL7EnW34/XWpAj8nDDJ0WT9KeDp7AcUS
NthuzEOVlzsNMObQWXWG3FM/C6ggCTuDPnKdyP+F4NTcN+Aa+dAuGoCl/WdYcW4PknyJPEVK51js
k1zgi0AzA32x9HGu0roR7vNQl2jy8SqUIxxK8LMvPuO6i9fcwDSGb+sXnJPjaiXWW0hjcKFfULQv
25DaGToOSGP+W60iCIHDzDro6p/Kv5yWyMUhipcc0JgxmjF0/0t5Zz0zrYi6T27yCWx8CpcxWAJP
CfH76rejBe0tdapMbChD8qYt+QFeSTZLyWhONJhZM0/KglpVHQ/SB6yc1oHxcb6n4zvIDTL13/dF
+Jl8Skfpv7MD9L6qcKQhvaf5wW1BReGzdZfwEdUhdw05TiyWbczfD1THxFJIpB392zLFIJtlAXOF
2hjVIQML3COcQeowlxSTOEOQSBoTzZtmBNO3g2lTi9G5fzZpoHo7O8mo2W6PvK8f7G6Kd+YJSa9r
hAGzXH7ljZZqLwCAzSJKUmEMQ5AGeKQ/2VohfR/VJfMpL9vjWmK07YtHdvP2144eK7n7fwhFWktP
OFsJf1lCRNmzVh315gDK8mtbxSS65ahwFNSrdWZkLJ4ox5tuRkH8SRk3TcYEUd/fNeXYXxvk4pCQ
oG+HBDj9Vs9s3az9Si8TNPbWaH5UcYb+cnRF9uTJe0Nu0MzY3ZpuKfD2rwvjUNIbMFu0Hop41PYs
Q0krNo5bDGpCzkGP8KP9P1wbfFmmPj1Brrd5oSDv1uwXWhKhLVpbk1e5fNkDStUwS54E6rYXLJfv
vAtXBJE2zHa1WTLDS6vOU0fWm9VMF2OgNbPepgXe6dcvxBK5V5yuB2vS1JwoAXq9Q6QFFbeexNOT
bOa0D3l2H7ovINFCCJUYWe+bRXPDaqvULatiNFBnR+ZTfzBRce+JRsnQBlf4f+oBQq1xiWFZ6xoU
ZvB51ySw0Bs9MbsvrtqfNlfMos377stJsKtbYvH5+yUZj0thGAcTayPnOHjMEK56JT/aohtK0dbU
roffFTzRLJhqWvEkJ68wSu+2ztju2wPBE4cH0l5C2eKZQMbTZbHzYIm7RkrYXggTVx3GV4BCBqxl
Ew3h5C/2BvXwN7VhqCMlYPxifLtoaSKMlr2wJDnlfYl+jL7wnEvAHgHwdpoA487PqwH72CixbFp7
q/TTyifFDhlxoenICEiqf21rqi8TSIxGBuYSC7X25BMk9+E+OdAuTARrBQyxmKty20U6bl5dnSzU
KMtEVOnDHdoQH6wYJSRrwYvrc5s8sykLkSr6cIBzrzzC7wvZAYjiI9AYH2yNjGY9MD0ImSDNoQJS
dWVmNadWMwXroSA+OeVffp7nzVPy99T4g1jRxPSHMbdtmENe5zDNFw46SB36fhO2irO80is1n6G/
F2v0sbnXt1dLl7m+fWXi2VUrUstNuPF0vaYlTkMh2F92g8C2THvnTfMt4jhzpjEnnSbjlo0Um7dC
2bN95kQLwNJEpeyTv88aT6SeXZrg6osEUN86IZnvHcUmY8oiEQlAsMxq38wcQC4XINdY5YI6kH0b
p3FrHDsbcFz2atLAeQKPnWplCglv+WB5sVX3bTOuVV+sJyDtAEx3s+0qUncXSLV38xn+qsRv1Y2n
mWcDBpC2Kw5lgPlDOKQ+/RNQ/67MQOm/aO/3Ylas76StLOv2cSUtJBhoLOccZXLI1Dbf1H2XwefJ
ubTNdpjiXRetS1ATKyh360osMy1TmFzQFUyyeSTt/08AkdU2d9WcVo42+OlLNuYBcpTpyDORogAD
XW/WFWBXKI0QcedU/xek4yDw8p+PuFD14KeELPAj4STQ8sUp0qcvzVlmQDz66UCodBGPSkAE7NVq
Oj18QVoorY2471asEptf77JaNZkaFtUZ7i1egALzYCztHImSHxxdT+/mmogvOgZT0ONREyYvXfCt
DEHmjWaElEeg1ry14p+uAtihqg21jULqGYGvA5l0HLFhbZjkISOI9VLynBEAhHeyJ6fr1caONeBD
GLrzeGdmE7weJ0EeG0/KsAWGJzxudgDXWrcF0Ln4M3ADTho9CplTiEBXT0/+4wcxN13VETeeBFaM
2aajg06hf02soRe38mX1VrU1e3T98qSrs9MyFFA7H0TA9elvg5cuTIH3F7wAT/+9Xh878DVPse5K
HjWfMbIR5lEnURmIHFnOHrFfun/eDPLikCxRP7e1Pz200FsQnn8sNcUV+lRy4nfwRltAAipGgTaP
Y3202JUDlMcjzRh9MMNMGSwT8bcQZzkfo7osRx0GoWzmi+tbrVtRX8l0wCZEL9YtIYNtHdZ28Rwx
IuieouiQ2rctbHtcVRTI2k5Bu1RwXaGillmDLGKl5sk3/g/Jpu8dH1+HVmXYzTi0StLdnA65LH5W
vTv6VSsACmqVsf0qLAnQpzBsn86evXdNkxTbkOOrcTqY/Fh4Oz6ly+97+cN80CN3yYbdwBTCIXro
q0ArLK9Nds4qnbhYaSZNhFBMjccuyjT8RR3xVQh+xTmV28asGTegXskcrlzyYPhU8x1mLmgyRhgK
68LVrCvLryCjid+Ib4wY2RiA3616rPrT7qgmP4DrtmlbryKSPnyMnE75weHrNY+89pxPOkiFIs1r
pFORkdAV7AajDVmuC582drwrtQKg6YIJTPFH+sY+OVTBliuNPM4N9OtrhttKV/Nb30gqVPJgMZII
XrBulJehMDm//tnTApo4WMnIGkwjvz5Dn3YQyDci9udvTU/n/jUpdqApDQqLGzb6iwKgE2qZA/GA
ZbLPIbbatTowAIVscTNp7nzD/PP4SCUmY+6tf0kaHgGmFmDxHGmWrQKK47RGtDiURUIqX2Qx3P6Z
yMdIsjx+jgIeg2blO9awTfZlVvu8XvWSinwYVC8kNYBpguI+07Rbvsy5qL/iYVOMmRNk5j89mXfV
qTilDG7dCXdOnBlbnzSTB1TrEu3n9M8yzHYslsxeQlRO6sWaduraaqK28A1Me9N29P0Upim39BHq
wDnb8QCsdMI9bkM25ElpMA==
`protect end_protected
