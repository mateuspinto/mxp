`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
leC158MEBuQ5PdIhFCHWjBsvqgcC02ncNyDhuTmB/zUtonlMfX5tR0fB8MpBYQPKKhSY+OwGKLJG
VpS2olYFh046o9LN1yCrCT7YTJ3GXmhcyfiSEPINO7jssx+88WLscZDLDV1C9xcK295ic38qN7KR
mckzqp1FkCrrAEytyq72lGLCTcDCvb9xlWLDK24W4reSYVAVL98dhd9IhKwnEHPsFokzcYfYb24x
yc+lRtqRIjTBBLth5zcWqWfiB2mGYGQcpUiPJcivKFvQ7cI7xPl1HhQfEbtzcCAxbVB41TZlzojl
lVUtVCpsTUAQtWdNeHHZTsRrl+jrBRl3EgNzD+FuCkMGHg/89gqJm+VGeJTxdPVm9bDCKXRqbsfM
ytKiHOtmHIaAw3acZ1sZrqKXOPy7HHTkJAudYeO+d1AnqonyWHxYC6OXyAFLPD3epBxnZhOZn7lW
FXRV5rkvxP/hkneExte79lJxj86dNp5fK/MXhwfYSAwUa8bFrybu6wwfmYpcnl1CTQ9qSZ51WfYz
PjKHDsCr5//Xi8VnP8McggDAgSNlaNXqxaAu6SAgpGnrOXf1p+WplAI6vlHqIYbHkPDxjrqdit13
00ANHuu/v6DWFO/EQtJRgITVVCzyUbJ21UfPCn+8ys/aKXF0mICEJi33kqtfBAZaoB8nkFCQDVUu
rlukKmUABRZVclOTuQy+keUoYGPcDKOkDm5SFx9cqJDX1EVuxHsz5t8FF0kfam4z94Hz38CiBUzv
aZj9J+CRn2NzkG9bAbMFxqBBnF7c37u/z3vkGPXRdO6j9hZWL9g77lgMdbWnVuL7fpyU374bYcoN
EKiCCyysetucVx4wWhqVlqduUTV814trbvPHYG3AZ6LLyeNpX37HDgOnvabX8IEE7MISEugISs8O
91gnb5nqvtekTW/7BI3xfxTrytU5CyBEqWxr+VyLD3rsnH15tb+4VtQ0WiR7YidTP7BQ++FH0H+R
hBGWJ5vKct2Qxzp4K8t7thV4vG6iiMkW3jHlaTRXbPpBUDR8ULIzKw79P/odOMWy2Es5BnGmCkNJ
g5m4jJa4thIdqybgGcokxdpCyoCZPpi+RPIR01TJqQ5H1sIqQY2DhgFCgaTOgh4cyT0ZAbqcyU1f
dmpIaQQklhssDXSNzVDgmy2nwiWR72ATjzDcSy32JhqCTvq5jqqGQvZYwAt082v25axnOOSVvuuf
mNW32UVr06J5vUgdHgsvhCKL7O6ZlTxyD9mdY7qjwwE5Z9ZySshnAyvUaJJyMtPxgogoYrOyhVjO
wV51OFk13N0gI701FvGpX7fZmX7HNye6RDnUl/hFxpAl/wgL15jWTnVEbb3kI4+BOpGq6ddjfsH5
/jIJ8Q5QOnMyg/fHsgGJbNmVYxyf+Ix1pq1U1d9rCidfc9qwJWgLlA7RVBlf83Ru39Q2A9WfNmtP
ZZ6Sg4aRlbMTWkkEB3U1duzsFyP6kOUNwzIk5dxMRw292Mrg0H4WYLgM6LbD5TJ0hwq4/seaw1Sn
g/7y8y6aiWkvWPe+OWwzNLcQ5/t8jtiEil6QWa9oaFE351iQSRyk8L4RT2q0kEm3AErfbElYXpfz
u6ykKE7Nc+s7BJ26F9xTxe4OKN0znyk+oJiG1JF6WffSjC+ELjbAG14E9QdFpU4WU9Nzsuqq0Qxn
wyxzZMm18V67Whu9ClyH/jTmnUKR9g024F3bs73uHcr8ZXFBFK+OpskBtnrJTTvlbDS7ewncYS0A
OU8FCDyDGEpgC7rSdlKrjgfey3qICvj6UXvpbioktWvcuyCJUAZ5R404+zTm6uMDW21d6nmR3tfF
VlLfxPikGPqjUUnOgv6hWHjziqElABhscDQoxzzeN4I9/vxUVJ0U6N2a16K2qMUF2livUYVUJ4pF
Svg4IjYhADh4Wm+O5XP/TYwxWW6odzwlWggvRIsWDq3BkmhY5/xNujEOglQ7jW85PELTIbNMRkij
0elW51TJF7LyKzNgZsAs8gfN+NWoyCIrT9vBkTpNGXfu4a1gzcCWOo75Gp/7X2VYIE1qjLZ4q3wV
J4AgfHKQbYDdCIKs5ryXagFTT5P2C+w1dIWzXJxi5TvzwxZoMQlabpPS1eRYaTG/mWXrxVifCmtV
gyUL8mcRo2KEVmcZ4QeywaNSldPHQDlDYm0QNuvrRs+XvhAHcbIdw1+h1RjBlpW9mSkfYYBzzs1j
3rh3Lf+veiOJcvj3p7u9YnVCaQhcUw7x4eVgKdLYitf/srWcaITGK4MEL11JnOpNFMRzafDbMDMB
zDWH5QSlCgVRcwt6Ay0H1Je0UlHO0PWFzpXRiGJeMmIE1ZSHEsz3KvLSbkeUJF8Ir6NyUYgtNPFD
otdyJNDaEE+t1ux1tMZ0ckpXzAnaldZHZeN2aGJUyf4e+X25KWW9a0DBrgW/1ik4PHIHGcI8PKO0
bNx1yZAjyGMw13i3zFByzg9Ry2d7U45Hppjx7yfvvmzEl4GWVQDhzye//dZ8Ms/tRw21oqBoE2Ln
mkDEp5x61V8isMJ8cfFHh50+CDHZF5yOWp+kEbWvVeaBkkwtgDKL6o+nOFt1wkSyVPWXdeCw/alv
y84hHF1+svVgIdeG643Zie8bQr3G8wGrUV8Sj0gWmAg499lqbLpukzDy5e+P80cczS0X6HefjNIs
YhvRRpqC+CrN3EmN/wgtJ7d3zo2ejvYOVMfkpUJpVMDcvwk4tUlALNM+pv6UbkQFj9g/Sgh8ofjy
4RiKsKNnlCeWK8rPZeEOLJmNlDA226N/n88JppG3jnyU9jY2MDd/5fiRwnp5C6qO9Ahq3ISRh7V3
Wz/IlAAWziO3tTlT1g/85Ec6UY0Y41RVrsgSQ17C3QasmWcqc4LkmvffcUCXB75FyiBH3keXD80d
HriWYOmvxHMZHlcq3RTT9fHvEtDRJDvPNJhc79hQyg1Wvd8vWEh1HkRBKoxM8vxKyQbUnNklcpaz
0nPWgVo14BxUEGLjH3rGCxplIcKjVmwnXk7Fkh9cVNqD2Hm8KXzSOtYymrdQrHZXGuVXBlaBMSeh
mU302JSxc/275U2u5kz91g6YuKDIgu0EFh/tkSdIQvFg5xssbxjvCluOVZfC8S6b9GsCcz9dMKVC
5S3e0dan9V6dtm+NqNDwtiK2eYycw+UsReWSdTWzQaOhezq61i0ECZkAxmrSejfVYR6J0ntH+YAm
H78aIHDRVB733yPtDoMfImrdqCuVPgr9aiB1psWymiOrzQIvqKrQf6to29edwkU52RMVaukzOoU2
n0tja/X61ywnCgbm98PvQA393GPvK9OObQlZnPDcJiOI9Pgo59TvfaBEJDuBDMQy3Qp3tJ/G9eLR
Gd7vkt/5/WCptLwH4DbnG0PNueVOTI+dGxy7y2PTeVL1OcPQ/Z8rbmk2IPG/L3uFoQvNX/OmY3lp
nxzIhECGwmG+HqRVqhl91CRy8D+Q+IXb4M4wI3CWXXlCEQFUfc3Wvfj/8uQwwBlVucSWy07DD6by
QAUwQK0bm204SpKch+6qaN4a575Cfc9YcaEWAmq7U8Lr5HW1tR/H23MoytaU5OSfVK3tF315/heT
pivqfVNsCJAljtxUGRGCAI++NO0gM6WG29oUriPUkIlAsSbmWMdpCMTPqPpQIWB9JL0wPeIUw+ec
5s+qMsDuJCMt2Ai4ir/sZVVGGISKAgM+E+jhwkzGPtkzTniPww3zNTUuz2N5wVWkaf1FIxwLNY4U
0UwmtclEBgqbTiuVkiO6KcunWlBklxpJ+WlOAyZD0SfoE9h1e6DygCc/CctBSmauqH0spnPAIAcV
SFF94jijR2Gq9LL21pL7EevYjRogq7I0rPW9dxTicXwAYXdTfh/v1ShMY9OUod20tb6xS+9leoqY
m9fI5zD5yLJYvq4vzi6iiC5PSWpMY+21d+LuTsUyPmgeZBXrgNk95kR9nB9GMK0MpdfB6IsU6PCz
uwtCZWQPHblIgSm3d197NKYYKJ4Dg5n2JzatLOaGQxu3Wa3bBJjxoujOrWsaZr/yFnCNNnqSJyC+
iVlgFjwAUDSxmqTOr3Lpiy+9jmzkX6pHzyLc10d66R2Hq2TfkuMb+/ZNDcvu2CTbhb/EZo38TnSh
zL+AhwpXRX/YR/dbScIMXJbsZkmaobuKISPHjbjupBwLtge4ZnAkSn8NoBGu5NWBel9Qf1MA8aN6
YIJBPhn0eVhkOs2tPuP+ffwlYFqeeQ+BcEGqos+vXrPgmIgfBWSkRihbOrcOnJkgOW+QrIdbVWJ2
w1w/8sjYWwN/hvV0Yy4Bp+P6kzXGMKyTsVMpHDmQxExOb+tV58Pa4Uo5jg3/2b9V3H/WEKekQ8A5
N4W/Bum2dlrpabFbVA6kasXwZMjNYraGCoyhnZpTQsDOvZm3Aw2pL8HZzGq7T1JY0T+41cM+rD1N
5C20wEnsaFSvNvU083Boq5ncgzVZK6JO01d8h323zJObXLY50B3Tj1BhRClqYNC2wC6zTDoGBD13
ahu7bKU382Tz552ET+EsiohQcpRyJGUWiAyzRLfyuysKS86OfWcWn1Wup33EZwQ+zsyGDfvSm1N5
JvHUSGcxHTmneHpfgrayMD27HXnmTp7hbCUeTnrLgEsv7wok2vbgZzA/o22napQbozy8FW5+Rj8T
28N498hQj9O0qYWsKpOHu9kinGRBv9FJuIaIKQtoxY58KuHMwbXy4lfJpvd6hZ8F4mxi3Uyvub8H
TtyIXmXDh8Cu3XH0ddYO9iXcPVwCrN2T10RRjdrQI0x2os80UYJxzuJTokCC9u+SpavuQhULBJaF
8jci/sbSyHrBoef96++GUL1AukUwNZ87qeSsRrhkJnBEaLnORsX8atfNmRF4XQKgpE3JcSrmOaDg
6t2up6Jn/v3qrRK18nHvDj3zMV3k3DwH8gsh7GWVRPxpV91pKLite4Dl99f5HwutuP28d66Y7FgX
9qV9sEJkEjeYUJdovTkrW14ThJjuTUjAanTIfCCC/8C5N0K6C6liAnmpcdeK+FOqKH5Zs92PkUc0
6+nnZWbxKyIjdw7XYBiRkPQFP8vw0RID+lt0ReQiPcX6WdwIG7nFdYZQmfGc6QtoDto41JlNTNXS
B9xbhHEKDlGpnLXELpP8OVTReP+t0uMj/x0ucDLPYEtc0HcNGagI5j0jXdSIs3lN3YJXkx3SNQSO
MPPlo930JVbe9d2r97q9/KmceSXoe3yTy3ZPPH5z8aJvXwNnIuUor7UiTNJuEVYwrG4Gh5JXbP/8
k0aSBizImpjvzyluGJd8tM1h2jKxx4pmXUTiPihX7mWpooNCEILu2+ywzZCE1KCx4K5HNzLbIvNS
FF7XJ/csc2yCMDdPx1rsjPvf2fnrWoTyOYOmkQ8rCwYv/pEDL3t0qYkxVGbq3YxfaKN8xBYZSihW
6Ss03jpqRYgzDnsXclM60b3Bn/j025hSsXdd1s1EtBJMiv7A8STLWfoTVVJ/c8+qiO/TzUL+qeem
9nXz88iRGGzvrVMQYDQpkc5QeaefvsKBAc/Ue64qhLjG1TuLU55q2GNGV9Ov34puUfLQbun6ts/n
qEyyjZCl82ZbmsJ+KQ36NzyqQoYjphVfHw3gWNamitjPxIjfDE1E/ZoMh6TNvSyeeYbTH2WJvC/n
qMQI1N4kBdLIJ6G5SKk5TwL8V6WJQETa5q0NqYuVMc0uHIRR0RnD2zXgRqZimurLwM+d98h9ysRn
Swda0t7vJ2hId/oTxvLY0vaNESPTyhTOtY5IaeFQrrb7ySsLxb7fUvQ2mqfpJ281T773XuqlOEVh
TSEEH/aW/5XA1EvhB8zPcHoc01b3Z7EDBZDgHBjrooMl6AcGZJXdWNJIzvsxoktN7qF7vOFzEm40
sfHxw9D0IctcAHuzq6e4ydA6ywhta/Xmfr1u0bcnS0TMC7wsD5hYI/3H8mDK7LjWoYxgWxiJEuxX
NxwW+mNRGpKShno9eQmTt5QUp27Nk/UO7Q5pLfYqdyEwp6zYtfixBdk3KBJsUCEkSUSnaDlwMULA
uW2LlTSIljqoTnGLc/X4C1dLOSMNxkyfAGHrFfm/EhDXqBuLEVLMGs89PA0TK6OteTLUaj0LU55Q
y7i94E+HudBleaY12BjOlEsQbf7ykVkwLp+xzm/gqEBT7Lx22rrhhNbzHOznuOOlRoTVUeTOUWsi
vZBHw3yZmM1K7NiKiebE1kl9vBZg0JpCz/uNAgiHuHy4xhlEhdaBEQ8cxFUJeZXELRze0lWhYa4L
l2Vtspj03Bv1dhFOQ23DANVjb2xj6QCv64J63gZojc2NNjWQh6a0PPnyCI6wA2upeVzkWPMfRpk6
WryjMduUW/5UtY3pDFjk/Jm7uwXPujn/CYNeyGeC19zjYB3M25X9P2/vcJ0Zuo0NZn4LrSvlQtFC
wZct8GKBHe80W+ykkB0MG/kkuXMgtUda2h6PtM/1i3VB5l0FenAzT/jy5xk7PXYmksTPi+4ytCzS
htcjlTyECMXyZhnD2kWTIhxgkcPf/18cbBiN25Wy+INNOUZMjDLS1w9jqFkJNkBcVcH9y8I7XE6q
GSKzphQ7tlHcr8lm+RCXd8epd22gh2gwvLdiIteD568T4jAqxE0RKCxL86NV4sdJyo2YPQGxkDZQ
POOxKtLhB1maqU9fz0sju/HJB1T3+Hd6VCNy9DHuSNIwZZDT7H0fZIE43TMhN2yteUgYqThbAloq
ijQ2zL/9imyxSN1/+NUoZf3Q6GvXN8WDMBsZ5NcDw+VyKA9Xs0cJ6jxD79esRVaGghkxwD827To3
u04noEzJq/zZlO9wfledm0RlAKOU1p5OCQ4jv9ZUOK/4aGJMTMNofTnbTgn6UAzKw6pRu/reATAg
bHG6YPdIqEXzusYKPhaeWl+jJTvSxqAeS2xBQcVQI/0rbzrML4wGMhso7FZ1cGCKlhlcH2eYosXO
f4Aq74e/7UPHgGBdviGUStvQl+hjVWaMg5sPimqRqNcNmf2J8b8OKBQDxHPcKDkC5/FB39IgAMrH
nxkLYrrqiu3PNMtl/MorP3sOsyeCySiT6ty/DQGTAc3az+6t2tlKKBsVXn0X1LgQu0pPlR3g8Pio
YMTY9IkwXdBThPWSFyDY2+piJ2uQvKCvqqL0CUSMaamSEjhGAQNbFTl2HWUggjd3WnzlopE+Yze/
5cY7yKbxTfcJcAOLTjKYuss5r9DEIGxPZtkW7wV/0DKWP6bFGCQ4DTTfM5p8HuFcS84RkU5lsuG+
95Ok2O/+Rl0ejhDgxJSxtFTSsxOTPpK4bbgJE+RPiXYVkStAO9TP6t+NWlth560KUB4iXGKAq7Ub
Ressqvsv69/Cs3cjnlirFRMQ+6g4hihaUYRfhtahFR/0ir+3NbaKw0r9iw8/rNm73GgASg1/1S2h
JS3I9nwOKplgsQHfCWVWptq4m4zQUl0bKhqyc/i62Zta0E71O1F8f1j0bkdS6o6W3gjHe1KIq5ea
qIlp5dpbXaVXZ+Lqa2/wv5wE6wkIlvTmAb3WzWinLqpam89Zo6QZOZ8/k38qiN67F0MdTHtLmDBh
0ff3kyD2T/w8wGPiGWmiM4GNEwQq4yD5MRsDRbzX1sTaXgawESrtUrfhzd5YVkngUjSKO1BRi9ez
yE9RB8NzFsXzZdQ3cjZjDjbdcguvtQ9jZsp6I34a5yEzPc3/j10snRWqIG2sEzJbdszWMV/9Hmeg
FK/RQ+UT/7DDqBhyDAc1tnhlsD+orL2qzPbIYeHCDxWbSR2dDBIjqtygLkUvRujqNkdq7i49LCnk
hf3wYmmYlqavse9S/3OilYGIg8tcpZoI2E6Og9W+Vjq7gycYjlVbdB6rATkc7nP25qEaCcBZrI6E
R2KbUDjHCZ51YNyhvBluIgBVIqznFtl6F/GIZg+C1c+FogSWApfuDtscQQOJJjIFA/8dZQaj3lmM
aBBO8CeOusdAKgTlyB3ga8ej2VrEOrZi09m0nbfC4gJZ27mvBVUDmxOOW/UsB6Y9XsufW5XRkJRb
FmWIzoIV13Oc1NmytvyNxiiP4QS62y9vFmlvOrzQdSVt+ielOybQIIUjlbX1ghL5eZPQKRptr1ND
WdDD7Q0CRtXMZZ4e56JeHjnP0oR2vnNshRmPj9z+NbfJuYxOi9nZHxd5TyNHTPngE0TmZR1vWQ9X
2RlkNjcm0mafAd88q2tU4YkqgjiagRcuZcj9oAXoA+wnjLTWU3N3dsX0G0+pybHmhpL00djQpVvY
f5vGdvlLMNQ3rkMU3v5RhXCYcpAnknscvIyNKj1J5TXC5mJs5La33ra9IJDw3+ecNDsAsZd8KIH3
xXI+zmNb09QrzhiejoubEr83SBIKDbcyhlDtsmBpe3TlKAGl8X0s7vHamxSHQfepw9osXOmjDSd5
XaW0PToYzI6fHikKEjdbMef86dVpGsF348EeHEdJClo7g3st5A+Cfn39nZcd7jlnZBcdwxdOBFm1
FuhfYJ1PahXh8VXDmqfMDeaRQihWYUnWXZh0+iHk9sn+44YTdE2tt8B0qD2eOBh49wIATbvI7kfS
+YujuNYu+saAfId0p4m48U+KHc4segz9Vyl+FQuC/flkVx0agzKkd85jj+TQQOG4ODbcXw4SDPrt
r0P/eMmQdZt+vP8v+2R+J2qDCc8hGCfhWMr33AkI4iCaxkhxGo54Ct2GnjIdejYzpO7J5yfCuslY
HKQqH961mv7oMPAuV/Cq0aqLYt7IaUEnwIorjwOxcfZ73zreFJ3/M139jBpqx0P37oc+6wdejHO5
wbzdQHMQ8RRdqZzXyR3Crn6z89Is0sJlGCOTB9j5fsTuDL+OohcgSDnP0TJ+verSrLwfMiLXM7mJ
GNYL9hobnFRKDCwjMcxZKk7sX69IMYOQ5gGjSzahVes7LR3sjajzmTfMfhg1VSGZ8llpGCK55B/p
E+JNlsMRc19EVljuYLBans9t6WBJjfx5nc+7miL+Bjr9E663xbD+tuZrsO+KBpCfQim2p068KuZr
Rg+PlaIfb/dBwC7mwzXAAY19gEJmrELU/tymia4ZbsIq4Uj3eOe62KK2Vc7PmF032eeXfAn3N51M
QcWhBOiHAvIpi/wGThn0w0O+CNGsiT3jgOQE7KzE7rzY7HNImfSgCDx2CKvj/NXBkasNv4Ld9VAO
AVv/9GBtMijHtoc7tvNkA9jD69NK4uDmIQSINZwqWzr//Gdyw7bcaqOCs3dj/4dDxOIMKV+Vn+Fp
HqgRxQTxMoWmcS+mY4MDR4ZYsEd0SwhrszQxGmL4knBHwnCLySWaERihyUXXfyRdKa+q1BEYjtA5
izfnhMlKjvy5qo6TA8IFn4kfXHOhWPt5aptzD05qEDH9KOB6G8ZGRryu19eVlEuRoardx+o994kY
LiZIoD1Xtu25viylBQUA9IuRuvRKuo0jw0osMUruHLVpkDVZLWtRAwPI7uFNoHGd4X0pSbSzttyu
UMg4wnfHcLR6uNfg6JfMtpOfJeW67unhXW5F1TSzV49xEbU7WkNtaHRl/j/7DhuZ9mf9mAlsHQbg
Fk8GySnUrW7oLcOayRpPdP5z2Owh0Jo/+sTsix+iXAcrOBSeKPg491wEwJqhjhnXNjLw+d8k3/Ey
FNDxkcVOCCd6031CmZPhM/Uh8FMY9c2KmiqovgpTka+dLaS3FeU75li4+r+gWmdgWrcQgDDDPfgS
rlzpGsOSFqXyuXjr7V4hjaEHSTyXJdpWGk5NQySR6ozeSWiiap0g1g3pCRcwguSM2cIiqUEtqfmS
LNpPmmOPDc9qBClis10Xa070gdPTgfhp/5tOEu6BJnQfHyC25jPchyCzxxg3uW/owkDSsq70keuO
d90m2GQEraKSvV/kVw1d7Wz8xsM1+JFx4Ne/cquNCA1F0YkiogxyKDmIhPZOuqKMablQ8zZdvq4l
2mdNgP/sPLG5Xx1OoIx94zdo8BGdiSK883vFCP5KEzr6z1NEy5WX3iR9BOZNT8tOfsgNS27TqwaK
HZ3GV6ArSIrOwedGHeOyJiZ7O7e/iIj4sfB1fohR7BdIjrebdm7otBqqYrw1y1r+cd8pKMzTS6Pv
fwC5nCu9AR4i/dt3JE7DYRSCzaxbZgSz5nzCh4Sig3QPorJNXIlaW+eFGRKxJDGkH3jYcPnULqcf
/fKAKguGCznGx0Is0vvidRwjrPDc68RMhzKIGrjSzfHE/q036e+SQUQLWeLeVcKCwWUlfVzR126x
ew3n/knVY0EbWxeA84265mTd+SPOWw2YFEFxx7l1FzERTaZYGY3XkyHvKiaoGyL1tI4VgqJFhDI6
TR4rfJPpsD4Nh53OF30aDRkl9R59woNIIeKVuGzmxwrQoKflfrdBIkRmJOnRw1hsHj8YjJLaW48C
TDgcuo6m10spIdASeZsZbzdhWWjhC47U/fzcW8JCO8kxKFjBXZ8q/aCs81VsmHIa6WwC+f2UvYEb
qwsF7QMKVQ0HPQEMrtsZy8uU0YSW05Y2wQlShe6q6Sl2B3yXWFguMlouiVS+yzak7n59fIHYc9TF
7mp1Fcw0H+NhZLvvL4xMC4FuKLwexYk6A6iBvJIZKl5/3QgjN7H+TwkrE7Q2okdOvQHwea3ieT+n
JrR6/AM+1weSPWCcITmlciXRPhB9NIdkJnsyQ/aVZudAm74/bL2QJ1A0iMwiDtEvqQqo3LfSQss+
C7AyHQe+TIAKigo0poF/coGwYdOSvio3Kdxfsm+G9OORYD0/kdIY7Tb+ZNU9R08KmEg0lG/k+C3P
C3uZFEX3nRdOeobTTnIFUPUpKan1INlG24XZrf70TQqM1hLk4/3QKjiu6VCOSuEuadVbhS64GyIG
hYOc6Ilfkk+3Xjpe+/b8DoeQJ1PWuuZyoM1SnL1ZiOGvivJCRAKVqvphV6ynYqJfEfnTsYVkOnpl
k8f5aC80bKcUphwkpem0SOlUoJrpNsVYYCxG95Py2j3iyoxdPLdadcPgs2csYSyT6KU93xdM6+6Q
ZOmsxINBDx6GziuTTvkIQxD1Gjmmd9lWsYS7KbrhNXoKGRxumRXmoPsRTxMi0rOPDUYFJ3L/027t
a+aY29wjNzJY4JLUeksUeAFkCiPvudWhEIgH7lks7LMB3HRmK7J3mcSTJHlpAdLZqH7hbLez3NHV
GOEWTrf6CXyagi+qXtDEoh4WvwB+8OuEkQJvgcnk6MpCzTpyCS2IY5hqa6l2CP8RT7kJjPM9vu3b
ZYhRTIPln3pAbGov0j57XNZIdxUDSKM2DNYY46gh2eztaxe66ImNiEncNsBmOw3JXzBqAyYw4anS
/SuaGhGW5KyPpZy0azclnb7inegcir1jyUyYsSkuG6LM1zWn15fJiNjUWpkoYDU85dAzVMFSTaWR
isK5tJdRLrzECmWq2LSWx/tL2DKwz/wuLs3/WU70YqgZl/x9FjfJxwt37NyKEP8w4qm+GdYiEJeq
V/wdq4cZ1YgWwt2NCoYmG9RbTBcsLnlLUFSGCei+yFbzjJjwaRJKxGnxDSduLBKGA0hv6p+1TVYI
eSfke8Fm5wb+ECx+7f8PLNN37cCTZBm0LIut0rKtRd8UvFBDc85L34zSa4hYe2a/wz0Q/oDBMs7+
TXXWq16MahCILmvz7Rd90WkVbThlC+ExAyt+5Lyo6V2CxAz61sk7lcSJpF1G38+nvJSmhsIMJK6k
ta9M+w+3Z7iCcbeBKp6xKsSjcJTzqtZ5rMtKYosqT1H7WvuNg0Gh+CgaJfAzQPLjwkZXDI/mkbvV
23DLu7lBHilghnSS+O16zLhI/c5mFb3vH1s3hJyoootPyfXER6O7UOpjb4j1Ptw7/VjxeWg9qMgU
x1Vp3b233acz3hEGjwkufrFYRgyxonKk9EI508U4seCvIO+dTdGUwQSu4U6W/cCeG0jqXfPpufjv
fKw6/5BBV+gIarLp0yWzn24WQYPZ1wXhggf0Rwi5Y5UP7yVFX7cPoitjy0xA1ty0atVf1fG4oU9V
YbG492DI9joyFgaLGG3Yb/VXOkLSCfqwxG7zBVr4qY9ZRotuKMEAQBWgWWrgCnHOWUodGqlwDCwq
QxRcULRgF4v64lUSBm5D56nvHy1BC0yOeTJDVtzjmLo2hAsq5NcTEWF2yB7ZhCPmXAJCOnlzQj3T
CIH/vFgMbcSkQlBy3uZPCol1cX8pE21ON+LnWEl2a2BWmVPOVh7dNFrEyrvFrbxcoSCCaly6NeFQ
fSa3W7molz5CfG/gWUUrYJthbVPg/YZOEWzyyFYnEMISF5bBzAuDk+NDsQZgViBBMIl6am4ccJni
3vaTqKrRBMifQESRA4nLQ7mnDl11l2ujIVpjqr1MnY0sc6TFMVKzhj+vGj5sx5iPjuPtDnrA4nAs
EQtfsf5h8Zt3I20Agb3m72DjzcCCoJNUz7GcBXRxiQ43gnOu2o2gLFOrI9HTUYsbcmTLrwqwrakT
wQIXuRRSRd/cSj6tSvYb1FzFh/kFhZO6HtXwbdT160rLf+2vIYaZwmU8+lZRUgcivmHb8nGE87uO
rW4FpgOgIdmzJ5hCkb3iw6L/dlgAQEFTOwT96RrQAF7S8KQY+6IGQjtMV3BMc4TpjIOWIziYchEx
4JBK2mq5RzDV+4m6WTpmKHv7QOYW+ttg4DZPozh6xP4XJekldD8a+wwHOWH26nswqy6A6Rdlpi+K
lRr3lvFeMPtMv1Rfa0wB1LiEnF0RFi5iLnKfuslABqdKjv+SHkZ5Y2sMYt8UCHYcSaY0idWqbyVF
PS2+vijnjj1Cmv0/9YeOEYpFco+8kJYtm9pdBiLhjhjGkcT9HNZBOWAcftq8dMkoAz7uPPVRTBde
F5V3unfDLwNb74SVVlT+HQdEl4OZLRpnMrzj3zYUFur3yGqfhpFfNeB7Y1FlT8rW1JYGa3ieybQV
35FqHNUu6A/gilpLWPuF2ApNwix8PgvSjXGzN5Dr+I/RoF4HdGcLqLMJQYuzmZdzrz+TUnpdLzxz
b3KaN1QLHjx4T72E5IJ1a+O1hL54ah7/rB5HEWbOViF7ZCQV8XrAiaqi79DEDFQwu7nB6bTyTzCH
0uC+d5EQILVM/f99j5Iqo8jFbjh6TZvp1RavuCYBQIA6TUTwavx+OIR6p1tztF9X/BGpnDZX0HcO
LfQSaF6wsVVxpPPu6ilBKvnBgQtMG60xOAhGp5KxhOLY1G/1a6Q00Z4NNuMDjAfrUhmtd9gN8bUb
im2pA59uPIORPQr+qeOMfkQtnw5qOPWdOVkvDS/fKeBNxF0Wo2MjfSgio+zBJ27XLOqiVtUP2iur
aV/1CzCaLkWZgfXK1n9oxB7DQc1jFRf0u0QU0BAKnzl19jZMjBwkqjcFi2cf67+wCbA6ALUksSID
YTCrzn5lVozw6X4rIQsKWPivT2cfjnC+T47raejCp6IZPzIi/mj5aoMwOXOGosYX/mCq2Lau58vp
R7cZgkeA6GBm3dIR9h7vXWGcqAByNNXDsVhVKcmXXRFnZeQipK/c1qlF9deB9BnDA0atYV/kaWjb
dyFHKS5YThuAAtHuEJa8Yrtgq3cTkOiMV4HfrHj+AtjmPcjA6F2PBoWeHoi9nU6g1IwoTW1oIWuc
1l8coJMevRkZL61NQbH9/Wmm5rWW3NqCJCGGCx/+DbFUvhon56Su0ZpWZsOkJ2N9B+4M5fJzz5r+
hAhWLftghkvjTcqrpUoebWGeJtNnDrGoU2LaRK/DX3ClSzYcHODTuJ9xKmsqpCp3vc3IWfCmXxhK
2zbdnFszrj6qRlYOoPpbDqWK2jgklZHRWwL5HF8SYtsMuxegqjRUDK1P5QBhcoqneVyy9Vw7x8xx
wzVaOBrjRGEnvMAcbHpGwHx8I5Mbl0wIjgxOmKPHm6zSl2PJqZ/jqZGWym+z/ilQXGkOf5MhWe66
C6qoKP0+DOgiGFrtFnnu+ldj5LQjQJ1xhkpQ9txVYFLDiuCRonvOCwBMuSBtAS/GXg4caScAfta1
kTzNS8uQhzFasAHYNCxE/kR5vVCKYTbiJ2ceXwWkw+gH2L4vwC3R1DScCHm0YxEkU3DPVPLMF3Z7
b5risuPofFoVFof/9r1Q9wyZ8Vc3BI8B2U4oFza6h/epn/VxPfMGHAUN2Zujtpp+ifuAXkhrhX4f
Nbs/0qDnx2mX4qzni/8g7mz3yONziB91vj9ypzxczmxRZ/aMN7EAVB1WJuFI6BD2E3L3vQIKcswG
4Q+q3tN15D4X8tJUq9knOa0nnCQNWsonrxMEtnCdBYc5lgYkwafPM05d7LyqrxnUg9Lo1y9c/vq2
ohfe6U1+jyzQMpD7f1OImpyGXAjDK2xmP/8luDsWcA2rGIO3ZH/eMGUameTk6rQm0z0V+2Q0cJ6Z
OKFsE1VFBpCB5CR9A7bbGXW0dcnR92ET51r/w8AmTxcLdKs4ai+yUa9S9dsxYkk4epa8JddTq6Cm
4Yyn+tBAy9Q59wZK/Y5spfVsGwDNh/VcQ4frnUGIpvtig7erhtcF5yJnkyDRx2MI/HpNE4agSeei
KAKbRPJ2tE6XDsbq/7Pceipa5B+wwxD+GJe7FBGec7ghoVmW/AhPPGGQd+WMGfhA/5WkN03zQz3M
/u7tOiWIMuvg3pshLYWEWH6ReXWTOB47Jjec2UFbPsJqTBmVkTccQxKy/tVsbKILK5EaK9pt/aRk
+iEa4366n9P3YxViUfE6bd9GK6lYuec9lQ7DFlQeFpYV0rfK6T8f1/EU1SSSreFUEbIGBYZxwcez
lNGIh+24iEpCWV5FnSohVpgRjkUr3CVYt4QHCEyZrGRsnfTjgW/Hl6Mys+q65eZdK308h+I+jcju
gxxLQklPgU8dUwtf+ZeISc4G/H2zakJSQbqgAQ+/4VfiYY5pk7Cn/nJuiu6CQY5pyI75eiAPVhWq
uvarDORQQOUzCRd7wIaUlJUQ3p2q
`protect end_protected
