`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
hmaviAIq/PTyWLDcN4Ltm3LvG5tt871kkr3m/5w+fgld6T0h1lrkL8esxItVzGQM/czoeJgCIH5T
JqJhvIyP7KqPi2BRrs/DqcZEtCTkvpmxKZCFG+JOQ+WeWPNrs816Iry0/XvgjAjPnVjNYcghVfLu
WAMRxJgW8XJ0piQZodG3G+8zWAh8Ym0JAWMULP+PGyyldnzM19y0aGh5gRYfkZdnK4jfCJpxen9+
lpd3RE9D+/OHS1t7LBiQJqE1Z3ZP93MYOyau34FJ6Omtzy2Z4rv8cAUTZA08FP3VffzRnznBElgR
Xq/cpqZVdxxxqQLy6mRpXWFv96h51fJKff3BLfXANPN23mZh89Xdk1/Kki0B+aExoMGsOusO0K8m
1XgaOB17QHf32cixPtJU+tw6m5oxv1x1ZKHiSG6/31p4Alt5iCXWiLGFtVSSZKzCGp7TrGhoVkqt
9bMc5s3AgCED/UjmxsLW/4A+gUSh7VRqlWLIWiQPKRckEjeJ0dIBXWOP77awwQAfj9PTFL4l75CA
7AZLfezM3XsorRgUC2TFFR/IDd1K0K4c0YoYlurFFWu96tnVdsvNBEMqvE3shgfgEL5EsU2xuo9j
kJ6JmSNrjQDZccpamigDIvo/ZufuSw3dnpUz9CaZtBnKoidBg3BYQ1YNNg5E5IO3IDeCAH9Ccxtn
yL+URe2OGNTD1RtsSbJ7lasIKyrt2RpJaIovIUQGdsSCo349YNJpjO1kCekVtaPx+u57Cd+I+SGw
aEAd3+zsCno5iqIv8jfqsCi/ezhpqKDBCue1VMCv+UjrR910xwERdOnuGNcJWF1/5X38CLIEOkhJ
2EUqdwtfbRVbKeNckQs9HJ1dYBZB6xvZcwceQTxQYAhKAL/Fl7gHC+Vv56+9kzLzEUMoBT8OZX0N
w9H0AogbOAYEVHd3Tm+nUSGODMv6JVT9Iu59NdtEJ5xIQlYpL2TlwEkYPUpG9QMjnzygCzy4vcEe
/RgUHtXqGe/bwTyfRI7WU/CfR2xyL+fE/jX+zeAtJF53eVsrxyEZHaGNHRZi9+js056ZbPE8lBRN
UFwVamIh7OpGNtAjWRdyKs+hzCCyU1caPCmxXKv8iCfr/LA82OzZrAReqfYDk8SFMSZxJGz9CUa6
UnyT1NE8Hg1fiO5JMwzR0jG6TklfEHI+51uAAbgg6qThyKweodTxmEMubHxYvRLuKvo6UGrkdfeZ
1uYNyhsZquIYTEo3w5xsshCWAsSJ5qXfD0SZb5y8A+QCngDMoD6EGjFb5BLHitjR54H5yIRwkRyF
Xi8F26qIz9YEZMpajQTiCVZXrJa5MCUYSprSdNHm91WB0AoM4hOXHskRbTKkc0fZ7q+X6sz5s4CX
HYPzyaE4FIj0HkqTpHwjCSFiJRYu+ZXwNx+EVeDuOBQCL4RaG9mWjRZfJfBIx7kCNEsN68WlZUEy
CBNa03782YprfMQ4RYlMlwn9yYuWgm2rlYBKWGP53pBpB2+0DIIAwrctgTEAcMoLA1dufHhER0xU
4JrwWD8R0x4NAt6BUllD6QoX8hvZb7/5C+swDxuWi+EOs9hOUMOtCvoQlsSsa/ninYtrqQLHAVN/
ohQEapskul6zwBxUqnNvkj4ffRUhqZITxQRwQxsnSBf8EF5RTmlvZgrYFMZramjl0+BpoGZSNBhU
2PmBv45AgqwyRk3mzrerwNyXhtSrXX0yIL284HHa3afdq8vIulrl9pyhFqDTW/R8AmqSvUv3IXkw
qeAZVPKtSjxWpKptMrrHnVPFYiAgt+65ao09GqbJ7q5GJvMS4FS+aq5vXx/PTMLZQ6R4xJ3fGCTh
nN1gT9nf2VbEWvXnS/tWS8H5jIO9/ylKZo7qsSTIvEbTQJxnSAGlhoCq9aEHcF8KAXIfc4z8AVBV
F+VDOYrPQxhsDb4MgDOllgvlRPMR3wFRF7S0/i4rtW2C6KPwNH1NbMakC0xGrx1auarCigKCeLS3
nWH6lpDfmx7XOv3ZK2T/NdoSOeln8i1HJmS3HZPuPvUtCjyxVQAdcmSdFCGbvxyc/EwEq3ebHUwr
ngx1WykrcT82T1WJlTa3CIa54IjKAecPZAsLNvfTP2bnAg3vCMH1iXTLhHAt
`protect end_protected
