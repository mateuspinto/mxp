`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14864)
`protect data_block
0USWSUGxovGsyBJteYpEoY6ezBqBpsJvN+td82NI+p54p5mH2LjJ1CaBFI2YBlLThWmCbwgm6TFf
IRJqOgQ09HX1dvqrGX1tzkohIlB6n2D5urdniM3MrApuzDacT27N0HXoU9wz4gZNRif+tGqUFr+k
ECQ4rFf4Cy4OaawNh3DZSjEQY57+FgwGyidT3cgGh//p5bjtM78ilDYa98ULj8FdUIau3tPo2irM
FWt92EwV7vmF78rKG8HQB3UN50D1J4NXH+j8mbJVzYYMw/hdyF3kgI91lAfgAWOe38kMkrxZyyMp
N5+g3O6JRRzZ6Uhrj35gT8ZRrXJNfWtbChKYjILlbfZ6I23lswUaMqC8AzB6fmsDDn+ipuZ2q/94
YUHnljj4uEk5jxU88N1dmQdXPTYNXUehj8WC4ajOiMY4QjYWZxVR0mVnztqID57LweEJmx39rNoN
ZWTl0A9vIAOgXn0fh8bvTkO2l0V+VPNfdvvud3BM2IiIpjV/Pi7SD/z7PsPM+xQyj2R6zxdTPZz/
27Z6ZbVOoHKtD3e/V8ZvEc9G+vyFkuX+PIWeaxdd16ewXIqLC6KRjq8ALj0kHSyZoKaHGtEsxPzY
7uSOOPceezSlrAKuMGB8xv4X4I+KIUUIzOFDfiQGkpi4QJI3WIWPLtfrTX/XacMhVC5RcglUihMb
PNmzIPZgAAE12UaYEGxqyQalcYFHTQWR5+fmBkpmVhTYFFDPQk15jkpWiXA4tXHJ9Ts96pBG0ce+
Gv75AQevBMXcUnstG0eP8z12uzx3z513ZkUl86pS3yi0kJgsTCCiNW9UY5sjIE9HpT/cbYwsYr/J
HeoUoRhmZue18iLZhQDs3vg71M+Vy7UlKnDbjZ6q8kDRbkfF69n7c/p7DSILjZgGhu8v+e+Ppi4v
lH2CctPrThxAeG05KFj4BnKoU0QjIPTYscLShdtesc0eOMs7qVOEYELgwvhmL1rXgAUTPTdF3xkl
R8C6mcNY9jPVFXTrHaL5wSANDejmCCXBKNk1o4g6S3Z2Lo+wa6oXpsVG0ulVBc6FJwjFCLT7L7Ag
BkKqJ4tJ9BPtymdp84a1Q6GTWoj8H97DSbAvWYi8q6j0w4pgong/xXvsdw9v2S7NWhpt6Mh6KWQ/
bsFqq33NkKm/t/x/lx6L2VFuOMe5/iN2X12sEySL5XP7LGAbv0bNnOzR7d7utIOgDsVF9agJ/6po
ckY2ztIik1Ryu//FMY0Vy8DiYCsuyZrlmcjzrMuFfePmZyTf8bKIE+os+yuGMmw+sTxQC/U09HuH
gOF2PHdc8rCz+u2InRpVpRvLn08mNKcBITossaKjmVgLiXZomt0uL/gXty5G/YNiFuOdhOkAdDbZ
a1HV/S2UcypZGsLG6hr0CPWzRbwXYyaADX9wSQEc/pGtR8PwUfvUK6d+ysOnjojc6YSTbudnO0+l
7xcmEV62fnZb5/JKfGrTp5bfX8XIpCppPFrzdFhxh0Bq2UqAe/PqLYNCuU+G0EZFwbbqXf0gGeRl
mcpwpZEpNeB4yV/MPt/5p503TA8qBSU9X/4C82LNxLmXtOD/W4EW8YEButuJXuDqlh07nXZxoTFj
DUbiXdcGcrwCm8sXPCypSFGcF55y2NwwvcXv5D6n53LKt/Gzkok/cRCajUSqcL6rnDO7G5yNQ0lw
pBwYEBMMj+8GElZAucNy3rSh6FxRje2nEj09cvUUf/EfnPHEg9qUWFpRcdUeKYXeMNh7NFDEXqDB
dwkPA2pFj7VUJssegZj7hwbCNcvL6Kh4QrgeVaSXkctoXsctwlVrJclFF4cmRxXz37bUkYovIJsf
GSPu8LvYxE5SwkEG+uE37vZP+Jda2drtKlsM1dZ1dBQQAKB+qCTjfQnutVkkPkGbWICJRZxgt3gq
wnJmJDNzbUgeYAZ/Juj7IOUgWPy8fajUkJOxOBBtnZ9qZkT8EwiaWQAmMHIGJmkBZL47pINmeO09
5pr+sYt9DreZGn8qP3vTgud85HytPEl9hKqmJYjfVIIwA0RYTZ+ZPyoYN7ODmXbswvx7htmAMS2S
FaC6Q5tq9XVLwkad7SKIFsXvbjXF2COXu5dJJtInw5Bk2CsQgalIFfH8j/5mceIV1hmq6Tivj8r+
SH4cGH0HO/Z+6YKwYufmRwbc0nYu5XO9RFmXv5F38nEknOJnEXhcKLtVdRpUxGACPUGuoBwFgiBG
7a/pJW2ysdxYXJcQWx2o/NfsUMwRaCQDueL1/7wC2gyMr3bD4fLL9ty6TE5sgYb4HauCCGn/dtmg
PM43001+e6RFxrz3O2z53ICNcfHWWvNArtbZmo8jTmmCCKgVu7Y0oaLvbpBA/epslOb5NwA3AK6d
AB1M0RTDx62l8/53Q3eeZSC7Yyntg4NQFdeVIfP5W7peCeQiQpb3xfqfDeBw3wtLSY5sMlAnsGZI
F6N0NwBMMtENFW01b0e8KPKvduGoYLCyj9xu84iFRXpsfgbHsbz7mAIQOJy+2xvgi0Ldjw9K6S+R
jmJeOOYGLiub6uHFEALu71l7pd+yZDerEeuq1kWQXCunC4YvZrFWj5ggoXNeO4dhCjL9ZDgT1q0A
rs22gYQkv6wb294xL2aBTHqujodR1Fman4xPxkUmup9AWX0hZpZrrygBbDskJviwkgCB6v4pRzZo
NkAENfZWN34dHbbbfIXozBptYxd8T5lTw1D2FCiZ2httJL99SbdWL9OLWZ3BSY6hTTRgj+O7LEMq
sr/yutXe6Ckk7dAeVmh9t6RnkkrIHYw1z+DhEEBKi1ELA4x1CoRzk8TwbUIB8WKepeJfIhSPy5On
l5mrMZx/Vx8nn4zor8zYRiCCuChGIvm04YJBbSv56tRsXjUVx6ssKtrtSV+xZdEFUMxxeM7Qg4l8
Dcv/z9Qz5j0uWHVj7OKBlvLEtIXd4CPBmONxML72Aw4DWQ76UEbAFlvjFQRSRskFc1ncsVtrwolC
Ub51+S5RuujRx4Bv5rc0QDjS35ZW9/M5ofgD9EW5CS1SltX83F9Dv/cnyWPk97Pyu41IdQqX4cev
cHoNjbpPtomrxW9oNhSIY2M5SKeRtT1aVm8YFJl1vRlrXYjNfPWiEFlwGfdWhIi6A4/5R7feIlVg
hoN3Ht8Bo7DZVe2ND+kr2UTY6i1Z/bnWefWKSMiWg20hle2gcwxP907F3RZfuXkvyUcnpTj8U5Yq
ij8xVcq/tPLrCKlkzNvTCt6JCKbVk/FoIN+5iJSrz/zuilo3eJ0JRt/sY2UwsnaCTQ4zcd6Bh7QX
YPoA2qq1BM/KethKrDb81ETfDD7KGl/oRMgdHlQpgOAzuMTcKCJHICynlIUhKxfGBR6tLCArW+F8
Y//dXcl9uaOm3GsqyVMATHhcCP2nZE/uZo8JM3tftHFOPoeWJ8xUuXJGYJeVfV5Pas7eRi6NimWS
F39I7SsrTDjtL2qWIHgj148UbBlLiq6jNsaPSXQLwEiDWUCz4FaW178S0TudGxxo8++eUtvSWbzK
2w/VKdL8aKdS5WS48TdnYY1VlcOtQzyMoQ4gf+/Ang50ObfFWtldWNNOWNdUWFz7u/0its3lBSza
4VpiOiqnxi35CIbMJGjHAXU6hsVOit7L/W7RQ5NID/ieFYMuC4qWyqZbfWk1AqrX6lMqiVSkkut+
ehioGTe2Nj//zlImaWOwjD4X4EAVMYb4qFmZxSrXPjCdQ0cq/eDfnO6JyoW2f7jC/ifWus93KsOD
MQxf3G8LDT/D6otG7XlTRjy9X5O2eN+EMIcZOdpldDG2R2Tsfo7gzbFcXFa+DcRPUjWEeuDTTeDq
I8w0xx9nVnq17b/ScT4yHSJvA/MnTXXI5kX2jZ2l0QmWaGPHrPJ3BjCcSWuXVFRXayVIqXpi/B4H
DgwwxU73CNlh7+HXHmoVfpeUYCVOjMLoiyUWWeBThGkuh3xxmILiOzB87NzOStzphwOWVJu/1GPx
BH1XRXPPEaKIyQvVFyOI6KdgyuKT5wB0+63fAu0lfCEiL3CZVzyerI0BTBqf2FbpfhQqCPCE6H1q
Oprh5uarmiwZUg8CDx5SP4UqO0d1QQ0ZoU67AGN1AiKZjRmiHDaaKZwZYypeZPqSBZKzZkZbimdc
TKilbz0TrNxXzRwIP+2A+qhYFnx6m/H0ga7FZ2sHABgsqLgD5eods3gGA8l3gx5dL+EX2KlHNksw
2n+iUZtVOahI6CJ5wyQrHwArKj/zCkJBtR/hdlX9jW/NsniGNs0LfxFyPpZvxhvgwTpq0aow8o4G
6+1kqyN6Uds7v2HRgYZaFadPnc2AxYsJnEAr9GPQCfSjmQgWrW8Zu1n97u3cxZN+P24VDhhQ/WOy
LeMJ5xZ+9hFfyxnxlS9/umWwvOXcaachGONVBFZ1lzw5JQmp4YkepFcUrNs15vR6FJFuH4mb6IoG
JSoZKZIW9+Zc9jOyVBOz9TDJzhpQwg3XiXV6D4bG0F4IKMGNttE/uI16iBPhczBp9Q00a78Au6mW
VmXkow96OC++LokmD5Ke1ssUUVhgX99fSf5NLctKn7nSX4/g0fpqGkXC9mz5tAveAvC7d1SqYllp
Yto/ZqBvMFmaMLTs6snaDYBUdbeLMmWenAUjSir6ZBsXYC4m0Yhn1UlAzDYaRB+GhvabBFbDgo4+
xQ9aa11HMc1MfJz8EIwvklMcL6DF7zZoMSnsujD669g6nDvlK36SOYrdEmMMK1cOFqslACxr5fWI
flysR3QDAuFCspKSzp+3D5b8sCEHrfywqYAP5ySiNK6tdJE8e/Z1e0CzzbAPyHlMv7VEEmtdy5Km
nmoX2g3trNaTCgfsRoBGREKgQFuphsYbJol+wIYfDzQ/fH5TP5uYnKmQ6eeT3t7Agikjjkq7khFU
3A1rcHM5F+ZKS24wrFliSd+7wZKQefEGM4xLmlp7d5QuKDZOhE3ROm72P2XmHE8HEtdFOW559jlu
53TkIBCarx00PTk/+TgMuEhZhkAaxykovC+ubi10Qclzqo+IuxlwX6rMIrgYwOsd0yebhYsAB2Qe
vUsKrNsvG4ItCcK7P+GdCPQLe/vYcqSXsXqaJtO/h3PW9fXbDlcZd6+YQ0hgadr45ejQDwsxPh0z
4CEJDNUNxsnvK+RqW0okGaxB490Pucp4SMSBog/rpuWPdifZv0Hw8j2NmaEWGZqpLFLS2gjHAE74
27Kn5lOMjWp2WqbIi35drPjl/jnFH7rs526GUIm7qkIxWDYICsbRqzCEX+1Rrqh2IAz3JCMCXnTI
Csj9reJxyDAApfkIyjHtXqgvhrMkBcXXVClUWUwh/Sa+4OLzHIeQVtFlQeE0f5+UVYL4B1wtDyg1
P6XPKPH8NZ0JJFDAa9OztXru0JjzfayPw5D8bnPmrd8kUIYlmT0murmJGdGOBIJRSyZckHvKyjkQ
xzjfpl54FL4FA1Kr32m75vmA/mkjV/2p5cRWbbXlErb96TOMzqJHWYqIlK+bDuY3edvOTk/jU8eh
3uirgP+NBifJ2o8BfU0oc4leuAUGMcydlRmNtYS170306HncsJaN8VjBKzzA94DH+cI2SyTLCYlm
Y1HAnYNI4qakamlznewDMyJ83v2ZkoOteHFNJcpqxko0MkRY7a48KjffRtoTxJQilk4oIAt1/9QP
QI9gDYpMFDt+ZhIwHMNhital64DEItQQxH5LVDhQMb3P5p82XS66o78OWB2ZUzy5YmuevsIwBV2h
44rv4Ak7cNcLHwVRWZ/V8/qU+crYgTms23Z36yJuJMO7qQiHXihwQ+5idM65hyleSH1VdEcetbcV
r3wnRbDoGPw6p/u3nX6/JuHxE7vK59UGpkycf8MtqnJk14Rmm8FWTUCn40A/lPdP0v3gvKmsWewM
m++5YEAuG81n7o/4MECkBHh1+96nL9QDe5MnBa/YxEexRNa6Vyq+tVGIKlmIbnWatamm3xxojvLD
RwaCjhZHGHTa/EhelgVy8WSToOpUH2nX5bN+RwJ6alP+JY4x369I+2W4vTGvKgWcnoPsgnvQVJRD
7P4PY6ATU68Tbs6tfA98UtsB7vYLJmdR3iBFuUOvmoUVtx3Bf7zV/tuMhFHDRKBHDketX0K31fX5
/fAj1v677KiSjcSw9GlgI8NCbJKI0LILD1kASi1iX8Q+PloIj6quFUbLDTD95lWwmERc9S9rbioL
WaY6znYGI/O2blldPejnYY7CD2+uNMLO/aTNN4B8yXhanE1Mk9kSvI44BlQ+BMZjcFDmkRJG/JB4
3Rnxbcz8uVNAwDyRhbFuVFJiouCa4Nm0xti0/w0JxpaduDLRlUyxb64w8AQmAnOUwg22mTvkBvaS
ge7F7phWg+H3ZChGT62Lvuh0HUpDE7GiXgjqvWaBf5bwt6S/aeoUI7W4LYalfKh+9hjwd6VkC1eE
Tq09ijeRSydzuj8+TlwOzNtzDHosqddnpYNklGSkaclSVu84QUgLMcpIXLBe7h1HDGekezNlr3S9
xZ6Y4TjkT4rJyxhCfwBnqjPaC/pC4wL1K17Y4JT5U9aQh23aJ0tK00yy6NQieVeOCuScNtAytBDE
IHRtWgy9H63mM/JuaAS6jLbMPJ0JgMYcj+EmYaOq4+ojAK6rSnE6nCXuwC3kmxRd+4yYbDSPvPbp
aDndfdwD/nScjmZDjHmrnZ5PvjyVqn5JgznesNzLeC1N6TwSXjGKh885Bms/sXgVy3Fb/wyqNffQ
ccMhjsa9K0fG6mOQeyfC5wZe7TbPWmpDAjYCSB7i5jmExnJDmzs7EIifUJ59RH8h6Ub+RsJXIlKY
eDsWHUPCqPSZnQC864/ejmsRjIqa56moJP19NcvXMlpNQRrjZmez+66/OWclONN38h7/0c9K0Mem
liM1KLic4b8Drboxz9HrNi5ACwumCQ0rG0k5memwOXSUTL7AIkpcfWLA1fYIql8k1QoO8JA8xhZA
EmAMrFjCaGBXbavhLjRUIjYjwqiFVSkajImTLKZH4v8foK1tDVD+HelrnPa2A9925KpAQ0Yu16Pv
JaxAtqf4+0M5+adYTR0ZMEzlKX/byBK8krlMsYWXNhxrLq4y9gwGNiU6kboc79wePXwhsW+3hmht
oaD6z19Gd68VQ7EtC6ktImTOAb0v6G29+NrbI60i7C/YlNEHwCBkIla3yVbsEAyx63s6nZ3CgxOv
86h81o8/n45zhneTphqv5yzWub7rPean6gDOA1qdL4PG48oAUs3JPgf84+Wm6Ew6jwa8JTtuA6gD
TELIhvLmdVM0mWTsZqseQaK07/K9PvlMh//5qlLt9D4/wFS1IvKAJyoajKxnsKj/DYKcxWzZLqkN
Gsu0rQInS6U1l8MxZWAFoZX7tVIDSwC/3Jhxi8pODGT8MuZrwMhwiXrQ1LmqSamSBBEdnqA0aeeM
Ypva4RX1MX9Xz5dYvkbL3hG0JlBBeCqOmkPwQJL85esxuADGlh1Z4y+IpuvQ/U/liZzRkP39RuKw
vpEjuNF+b89VO91ECFXKzviUrV56gjM+uWePXOzm+fi0OExG8cM9PVQDtiINid2UHowibXQHe+r3
xwvcp6ybElZH4gLeQqTJSQCDfj1IgsZQWE5ZX1b09p8ObA9nTkNL9+fAiWIj55QMPpOAfJQr+MIE
ypGXI9HKWbZwDfqDLffpmhcn/zX6k6nHbCOpWzTm8J7ZrkbphH32SOQhiNBpEOxaCOScNAmVQZcf
czvPtBXDZj7YPuo8/IiAY/AWJkh2Nc8Njg8SSBsqYq51VuiuhlVdqjA4K5X7A2pGXSmHNROof43b
a9GNfeklaaBTCIcvoKONkkrCvfj3juS4/2HHpsIpruEGZg2f7GFk8f5wtTjbqvztD1bJk42B0Yxd
t9UN3v3URq2o/0h9T9ZnCfi6biRzrhcyp2Sj2p2z+k5nKiHo1zwDG9toL6ThcXbtTclYdwXYdf7u
RVRMBftNbvXUGwp+QXVtEBFBXYhU6diK7fCNxGGtUGKVEkNEzf2P2Qwr76Y8MpAhQ9XmREQvRbb6
y/axScfwMmGgQ4eVuXr5uRJbEQ/yLsBmaFPjIUSzlPdo36/YKPdjPpHI7NerCnvbwyyhE2q5u8G1
IvFH3IrNMVCObSdBK/AcEz+wqthZi+39wCCl9ebdruzd1hteNuGSs58vJ5UlDoLP8TxtCbV49lL5
RXFSdMSSybWNv634/jH4P3olNJSEHI2732A71uuHQobQbSmOBQRCLWXcAt8d57GLQmpXQiEuosBh
w8Yr3bIsOd9vO/OpZ/WlYykYTRZsNsLy8tl2qFodBmy0NGLo244/O8mLSP+su65NeTBVsDfP4Jsy
QXp6pAfKkxJ3fpvd5/FCn4Bgp7Iqj4uF25zUhW9U1SLhloxaBlbioNu7alZoRpQQQCww9wZcBvqv
LnqsWsISe5CAjqr3weuyAYp2+glvfwMOl71o12DjYwAhd5E2KFFk/4txuqVUzxaW1HKEjJBYG3AG
FYRATI9lnl8fRKECanVDjmkAVzWm28ns6OD9rpP2fZKgdQADJCfUbK1ja4QG9VFr2dGjmK38auq8
1pLW78dAISUGosoUf+1tRBBKGAhub1o5oTTxOGnHep0dyAd2EglEYOXdzfKAhhqiGVuxb5XcZIyG
y8pn235+ufcxqI3s+El6Kdz1Uatr8TzrYBx4sy7BqqkWfj37Pre6x2iT1u8gdGhD8LvfIV+LV3o9
He55zQAe/ygDjgmAWdrttz/szrWEhi9PtsxAg1leIa4BSVUtM7Iyc01i/fJsJbydY7Fe3qtVHvou
h6SVbzeGeITjkpM4PQNJNENo8Ux6lXpUl9Ah2g+fib33yqIw0o0y1F140xdnK0gtZPHNK9oGkJ9u
67Qpx8Fg+7+EE+WAKPLQHFDowMRosKWhswseQQvECFr6K59eT/0NejWZSzNlqPkO2UBUL+WdAssi
nNdTecaMxAMFgKOJt++9F2Ree2432r/RIK3miNhDT88IUHReH/enAIOR74b2l9XDolfP3bakIiuA
xhfAzy85mCzfC6ExZafD0U6xwQVWTrip2Sxcdjkflrzlru3WFMk6TxPlTI+Uh2P0HD/bOJS+ZfQW
ns+jFdnkjFs09WNu81qR1khMXuYlqbSE6tfLNIzaAHdLDhz/zG/OZ+lYjT2lgt57rs1F6B7fHfuI
5ATyHghWWMRDosxKMl4ZDcQbcZLLawa0D/7cjqwbHhngHPvP/k3rrp6pFttzhYVCLOujxJTGUUpp
0S15+06z+OJ0WXPxAItgFfYil1LgFDttaCoUVVV5JiArUfQ7OaAvxNWBCP2cdli3brxRecakYuYZ
oVUoXM/A6RpJxQDfjj8I9a2HB0ZOzxF2YftkGzsq4reWqHlhKrLtgCCIquQYWSKsU2onmkSF/1gD
/0dg0nXYYEzADxI2gS+7TWOZb+4UOfWpaTgZRsgm/Y3LJ+gT54fwJo7Me7FHt72Xgh0xcIAQDDx/
S/B7i62g7d2kWhDO7G/qGPKPaW6bpxMC7O4bhiQk0gVVs6zREAo+WQEA6jtaHKk/Y/2lBTGcDF8v
AzXEH37Q92ScjOptUHifsV4Psw2LpSaNsCO5AIwJd3QopihyoWrj41yNNdEEMy3qvnjH0+li5JL8
sRY9+Hrn062XRBfI4CYjDEqT+OF9r5EpmCYxjpmKQCl7h4r1YlrzKcKCcNUeuz0ELvsf35/Ipj1d
3Kt7mL13JUy785FMi5mpv2zC4oU0wfTUgy1gRsyAo/2RUg8/81IxnME3ytk+Fmpzb/dsZM1510cZ
UPSX+03psnNyl+IpzunhXwJu8Tevy7VKf3vBBF5DUaR2/+GxtlLEeNTz3toQ/yLFF396JPjLBITe
hNozqFCKNllDK9det6I3vEElyxtLnynSV9ybjgu/tPrG/8nUvs4M4e1jcUfss5QN0C5HrUNvgj6N
MMkCxiyJWPWKbrej8+ODRetXmUuMffW9/sQnBs8sD1vJCc3pjl9Cv9jH6s4DbYty4dmFEoTzqj8b
iQyxZcHtqeiWQgV/WmUBEmUx4nms9pshqPahc7aopPA47aw0EDNz5NZmBjc1aOd7eU7AWGXfBBZO
38ibCJ3yiXT30PKFbT8dd5+Q5Up82dkBZHjsFYSHofsLLScs0ND6VYCxrerdlQBBMB1H+diCnfpl
jFXVJEBMPXS62uZJ90b/f3+rwNdEGDHyeGcjdKn4SKwjNhUO9IZQB6kVkE0YgqSyJNTfwVVyAczL
24SqXG+UOh12A9XBM+CoVCGMS4cuyMrukSfpMipK0KcIIxsYcEAgyZ9CFWtjhu88Tunb95yQl7Hn
0Tybdu78bsvmK7ZB4Iy+BBrOIu54YvvfplNASoUaUZRFsSr5JUEftJMPJ5jmYXS7IQ/P5TOqMllX
C5eKJBqyFy0SI2W/k0lX4btu+6GI+M6urZcFHSi7WVXInGDf6kZN8yy4osDEMGiBAhK3ZCTUcyPA
LJxciFsTpByPg58bgsp2szfriZrClEFKxmio4Zz1KMKKhzTSc8WJ6qvxnc5vp3HREbS4cGYJT6/g
RrZLRpPJoa8rMBc1OxeZ5DTcz49cjG/1Zmjmy50wKskMe1Eq71jz1P9AmDSDO7LibWGGptUAnZxK
HqG0z9f92Fk5H1xePuQdwGSxV1by7IoRwXpWCXzWlMqZnqVL2ej49gG9C9QLA6qWUPezSpIDteAk
DlSrHmgdVXmw38qwWB6S2YQChBVPgTcjiBJ+OL7S+SSOKoE91Gj2ayucTOJHDUHDZ8dOjIS1kEZs
6HSrFNRSWMeA5xZ7Hy4DjCP5frzRbewlgetnPnTy4hXpU59W/0wPxgklsrHu7PQPFlmpnT3YUOLf
C34AkbJdzJfe3+DkEbQz51UtmdIJ09KNyUr2N91/2pYwvqmjPx7wxht2qoKrKh5jLPoe1NV8H51x
mrQahI13GjEtA5OKtRVsYwFdW0SC3QQZvDkENfi5iCK61da8gyOM4NUAu5mI6YYGnoC6zDm0EZYc
kPAh7QwjaN+R4lWtEciBg+9CaEeVLbNwPQ69TM47vQ0z/NqwmMtLX0Xafpe+A93PLS2Cu6SRxVVG
xOete6wp4g0hpZGs8463mCI2eAnscu65sLEGhqTZDpx0T8hZ7GbuJuqYrDMwX3+cO0tMwPNmiqxH
vG3dc4xzAirGBlu00FnW5ITUKIJ13+QtQ6eDNJtzzH1reLraUhex1LxNGXpNzzknZ8Qm4prqOMep
akxpKGvv1Qcsa3ooRvk1OdM2sM73w/GaCH+5ahNU3KulkCQBqHda8MZ+sVsF+PdesVz0uWirCvnN
84E6qcWeHDe/E1w6HC9+yVaCFa7n3bbZkNMb2shrx5UOv5K/V3yulmQ052ZFaVLb3ZTc/On5zEx2
5AB/diNJ7EfEl/mcaPp3TYzhf9fEQG5/uW7qS4mW2SEeKfM0h0Jum0MgxPqczK1RYLX1KmCpIHV8
K3enwRqpB8dMMaWTofvxxbCd5L2PuC+JmEzuNuRukFcr5QlIaBipGd5ES+VkfpXLOLb52WMCIrAL
qjdEAVn8rnX6WWMsNC94tOUjtbxeSHfa+qwLWzHe6U/J6VTDHs6Vuf1MrWwDv0DJWQlwCP92xTIX
G+aJORX8KJGV/8JTMBDhWTrmeEEjMwIKlH2bS5/Wi6c/EqFBOnYEM0V2ljOqsFHO9n4QZgSKPsNg
3rys9Q8+7FhnI8Qq/DvDQAqIeRnebIAJENbEGKn4DmpphLQy5mwww5wmcwddYCsVRKPFawsvhuia
RrWf/1H6S23QgxGEL8ODZcfZMw5OE9Suy6Sj0+hZr7naFX+JTqtAqJz0l6rP0kpTYPstruGIAwM0
HFOGOnciL+8oIVtSbQpct2A7SAI017hkgQNbWx1xW1JadG1gtmfEzQGb8+gmEI+hvKciOdW7HZJ4
C1kS5MKVyCnr3YafXvd0zRZwKQWzSQc6xYPABJ6iUqEYs5XXPFQ+eEkLh/0tai9WLUQNJ5ZdJ1//
3max8kTuTU5sF2Y9CAsaL0KGQtF3Nu+sfnE7yOeaDRt/KSHC0iyGzaLzJhUn5a1U9qwh2N+xTj45
ph9ztYf0jc+gerDGYPHkUEN2a33j5y3mxVEjHZLqsxXtCY+JB/pcNsGocyvzsZqHKfZxYKJIKgq1
I8a+PkZOf/eWecnRUpLr1Fd1TaASeBGoBEqfLYX33+Z9ku922Oj9mxon948nypVr+X74jTYrt62A
JiDi1WK4dcJ5oSGhUEyJBAJNmItjaCKJh30opS5C1H7gHC8ruze9PQlJ7mVGwKOlNprZc0iLA3AT
K40Hdgnm2yHY8rr386Gq/XXqr2MonWojqv8sOKRvPClTfxQPAa8CipGJE8KCZiBEtS/CjUFYRsgR
/HsG8UWzg+RZLiUBJbzXw4Q1eXrK4xQBVHSFXmpfuEza8gcFTUoDrqszVEuMyfdpiE4pZCRQ97tH
QkS/m14KMbco5iJ55NBYNe8Vzn7MNaQFTE4x4ILvCgcAzdHmHY6ZvXYn1Ltwq5kkRBNUb0ACxQ5V
V7PYOdDST7zazmh1hFwf9HsBo5tmyj2YoZYrquWZy68p1tZQts6tuzecfd0yC89yeXc9VQr51mxf
583eA9vtsq+s+YaCd5yGU1ha6kT10ZkyIsuAJdLY6bvOx+47QyFiOdsWdaGdWPBvwALycrXUb1uu
T82v5QtgRMbKSMB2F4EHYZ3u9aG7Qh0EOCRecE5p/5F9dkJ2fKHlN8KaDf5Wf/PClqyld1W6TLMu
hgitGux3LxFnPCrtFwDgIlFdEEoPHQdXXvXK62Yk9Ch+WH21G1xJVYneaHaVb64zNddlcR/OYVH+
Z8luo5DaaaXMe83pQIoIfBiSu01x3FP6TxuL1pcQDSYh7Xq+sD+OgNM2ZeiYyjATKnJBJzCp8t5C
2vq4IvI+T3mohghOG4vUVUOH8zv6RXXryPgvLwU1zosCucGKSOfZk9hsdsu/tD6Lmqm+P7B1LX67
zhtXZsz1H5+5v+imt7rkzpvCbasjAt2ao2RXqaY4r8jOIvOxCQhREPP/p0fGXafrsffYwQFT/EoR
644n7/OM5gUTRmSZj+eX9ywIVxfO03XbNlfuIv7yqbOQawLw+D+HeG9gG+HiqRTQj3dgW4ae2nF5
FXYby4f78sYv0+s5OOpJDJTXgZj/sPqaIB//TocMELtQgI5Fwtuf7o1ZxVSQ7cjPWhHWwA1vDV7v
FzIzUB8yxjhTeAiJRti9giF2lSqvHovro+gcIzhEzmB6SjA/EwWUKeC5yLkZpfQXVkOTZyqnFqy7
iOJrlylkrgD9rXHHvuetpCVAJnZhu+OD2OUCzhy3czo+8daIOrrhMVeLpT9elOaWRCs0bwMTZ7HZ
5E3pp65PEdATWAAtvOsdKrp8SgmorqfO15wurLeAKvBSZr37q2Ui9oQ90rQ7qv0IwSMdBPbHcY1E
ag1WMqV49Byyq4H4fTU20cfLv8BwLuKdOA0PR2HpVjQuisRWcnFDta1dMm2M0WFPv2U5JeTiz3CX
q+fX5rU+c6V0zHoNtf3Vh1q4UWNNUX/lqOy4CJWUkXKjFkGT928qX4AO4fyosK8p9duLyTjAfYyG
ET5PZwGNpzj+fxjzN9ns8M/VFlKsEaIzAok1pZLyQJEKAicjUZVS3G4TXLKe3MCdEs0ZWF4AInTs
nW+aiQxnzrA+Q/DAX16fJ324m2zbpftsS5H0zZX3S891KD3AF+mrWWnNGwqogYdJc6005GIm2hKh
Lb6lT3Yh2ULaeKkMZE3hTGWg39OhZp1SWDwvpXg/76f8sc20N4UvwdgFnACUXuFfTNmM4ktpSnPq
WTNuRay41hidRTSqxr3+rv8NGVsqerRFMRm3+L/sMd59YoI+S5ttpC6Spe5bSb40Apk0wEAny44I
cJ7g7vsdoOtMR5u51XYxtK5VI/pMbDQtBGAsR4TvIIwgDZbF0YZUryW3Oz+lcB6iJApWueyax7Tv
srGtHhVJDckuBY1HiJLJRFI0RT9l24EYiCL4830uSpEAPnDN6eMGYMmCg0WDN699egASIfNDffr1
v7htWJZgjhPcA5Ug1N1r74/ZseyP126/sUYYduPfVLblr0ud+0Re9XxQSec+JjkZ5u3pXaE7yulk
5tYpCOuGG4OpYCEFd9w4U3wvVTEGWLByKwZwvD6L0/6B/M/5wRpqRNlw7c+aWX5oKW7upS2GzkD8
TSE0soFlKvdsSBsYEsvWEa1mFYZbfDIUa62l0Yh1fyQTZE2shifl7v5OeTxC2UaYO2j+0D93ixw4
nYyDrfsTz/lrWfzC6kkm/HX8Urn0aERuiBtIskbdqgb8ArQOb5CGnLEsYc6XKfHAZmhD4cS++JAN
OXGRO+DYF3O/ugxDMGDkIecQNNk8tOkLPqG1p+o8S3vaJtToctVanZHiuRVQE+pYhAHqexdVYLmg
jFIuDNMAoi8uOeyqsdebx1BGvjLxJscPetWHQAj1h5w9DVQ7hfXAw305xzcZSgLAOJcB80mcDeHF
iLrQrZ2ZopMd+KZBIZW30cr06NXQ1pkphrqRxWSQOuW1s37OtMmo05WcG9HpwwyxvR8KbB9u2R+2
E4GTdVDmK48n6RtOx0uPPfcenKALHfDmN/wltoCQJtxxWuwRDaYrHJ8XctBReZzVxca8+A9KaWSi
xQ9eVlwMCNFleYrHsrJgjwaJ199Xjikd74FNB96tof6Al05z0Hc9GuHE0hcqwJVjzfrXV/Q4EUHD
85P6hVWNQ8+ke2eTrlK6m12U4F7R2iJ9WeXyhJmvsIkuXP87tJRsQVyOVMxWwq9feo3WteeYwKVo
9KyG0IEQaPNyhSnEPTaj20NSxxIIYbLLYNenUl1K/qdbB9dYRRFa2nSCRmEvYAb90eOocK7a2vMC
NapwJzY4b3XsdtClj31ZqfI8jeIGrY+Sm/OVhOcuF5kl8ez9BHEA7033ejzqZqIkQvBXupmev/1o
4N5/Jivue0ExpOtvqLC/RLeRWsdG5RIRSL/GqBIZY/Q6VWUHflyp2naiHgkjBnX4ZrJLODinLwcF
N7J6fQ7mRjJ2XDXvlGqF3F5nCemvthOkQwZhDV7hRsuxBS5zfJFB9Nvrb1LTBljDUNPDme0ldriU
ETuyVuRWdrpeYZlTvWxhLFVxJe/IPJOmKmmX7CQnv1hW3qdBHvN7rhQfTlv1IlwuPEDW33o/Jvmv
thR3miG4MCpHm1IRsUvdMoBQ042qMaf+iRY/ft/95XWhKsWfsabbEcuOydLs+pjC0lui+S7Dmh3y
H0s0Brr67hfGnQQiMmEOhHbyRDucyjUgjeOYhi4VxG+i5gO/9BTgocgbKRWxWwb9wWi/sWSqVhh+
6fzwxwYCU6eBmQ6jZSoSWpcEIfW0jSLaurQSDoPgG5x5mLA+EIVXKMMuAdDfLujxhXqaC49d9vZU
lW3tKQveJZcHeyrBGwT00wpfa3JF3cvlIrPMyVONjblFgFtxlsek5Oz2k/QHKE3HJTtIJoOh9q8b
zDE65ooLWyy/GJ0P/MYnlTbz6aGEs0xYS1WoEtlJqScoiOkZ3UGw+TB6GQ8HzjfxrAmwgoQU/msZ
tu8rXCe/vpmVoiXCGZCj57sOYhhjHJFOKenTMXHIpjUTNVwvswDvG5qLOGnC7NyWPRlrikgPd7zX
9DFNzz5AEvoNju8O/Qz2WPlp3mG0qM+lmkYu9qXGE+HuK8yKn9AjHPsOTWloypXPH6JQvm1Jw9wg
jKm3nipXjPNBOl0hKeQpwfU7GfKPZylyDEeNxRAMYkN207LrjXcJe/7aMYGv1NQ9XBicZaJLDSDN
xqO2p5KJfvKxgqtPihvzFXTsHRpy1w1j0P3+gexc3lJclreMd+dKrMs2wQij7HDgvzlTt6Fj59eq
55KYKzo0Y3LLCebRQqW+DyReqFhb0PBt0fK8qZeeS19O7mMtjmmX/8SAYpHcIVrGMUF9NoU1ubrj
PI2WCHoZZwVPNKlAO7cdd2HryzTFS4/JcnMOigVuMzGCiutdh8kjLVHgjfmI+M9vMw+TxWQQWOmy
oIi2D9MYBwj4FsSwLc2fhkaHXTBgfbFdAZTNqo/+1W1stINMWAqIISgeFa8hvfNOxTBt3Qw91L9b
63V1vRrXM6H+4sWg/8PRe5YLYXh4Qxaa43lJ++eDzlbeGcb2hEy22A5yCfqkEMqI294Ui2vhD+zi
d25XTqcDP7jYKJ1xgo7JQeIFVscHYF+C4r5IWnJRjf2kjyiW81++SK2ywBFDe357mctqI7LuXFZy
+4OVEYfB+yQ9siCRe/MfaKTcwSKVqagkLERWGq6AmcAYmostju5pYFs1ACn47jBOs1TtrzGlYeXd
HSY0JqHU9SH2GYv+4Z943rjRlBPI6/27dB63pHvOT/i0ToUqyx5X3qGuqDHLRGXvw+5/ijEVTcNh
YZ2Z/PmqhgyxZOoojxFcqouiWLxFCeqzc2VOiNG8WbTY9jVjv5bnh11DTxYn3p5Y+7yZHqYB/avL
cFCs3o0A5ijfHTcABu3X05K2Et4tlQ4Ubn2UcHgXWYBTToLg+8TNZ1eRmqs3BAoxlYGAGIMLsvse
Bzw3pNpy9Rz3asV8E6MBBvcLCdM4exETm56+2Ex8nscttdnJVY9grNwNwp1s4A5FMRgzg0ddvyWM
kK8IJnrv5C47abKa5tcEuyQ+OgK5i+2Ow68lUKdL/lRNaef0F9fpZNSj7e+UJORWYQEMmmmXOFKr
f6MuliNSasL37K8Zw+j9HLC+dCb2cpVcArw65Xjwsr8jgczU4VOWZBc70DUNhlmiPXbsfsH0b45f
lDC26FNqm2TY/g51qGkFh9QW8+oYNXITG2nxM5smBSgX5BPzVkinSmEQHTNP+zffghfc33rpST1H
qWY7rMCWu4GgJRcSwagiM6/lF5b5pbfHi7nVNeSqstnp4XbnQGO4OoMMtn146gk+fTG2QWorm8sB
GUrFaciqxkW85oXVpHNAS7GTqzYLvGrmf8EBPddyX2eV6B40QlwGKyqis6aRDXAvdSeKeCeJq4Oq
fjMONiwMvkl4dbKdZH7pH9RVdoX51kaF+0Cds0w2/8lx08v897EZwf12cNzXOnEKhAtCEoq8Xjbk
qQ9ceNKlkVExolFqqi3NHWm20eFURnSOUm51u0z5lsADJsAVCbfz3Nijaht1ShVPCBbVB5FAShjv
/5T2DNLVRsdAd8SDEMu0k+v/+1FSD5TjiNwZ2z5hY6WeOblMnzCA0UiYvhcOGFA6PO0E0PDzZgOJ
IWYbMImvHD6gkargFmQwXGAScqDNIOiKw+ud2RXgf/afJUfnKDXAJH8Y9W31KiAthYCJFIFiED0D
hYYnPVZ1o54ptN7deInKpv42YyMBZM1jhEOawjPb4Ep3fPIb6Oicdx2xQAtyOifFrBjx10VYpAWQ
fEEzk9acajYObuC78LUV143bREIEr6Iz8KmHMxEFkr/v3ilJ26PNyWwld3r6x+PWN2/Tq77LVa/v
wUUlxn8EfnURbRQwexmLs/p5p+TdsA5esxwLAczjNmY6fmDnr/apDbll8gEylN/tsCGbEWd76ohB
zKnDMXX9yJT5tPe5b4NaeZQ4JpPxaWYez1e7mtKKHMACU08BnfbJC4F11f0gq8bINEEB6fAUYXz/
uV1BBCLsywnyJAjNSmCzFamWWewhc41uNJjIqtmwyAw6ofbuzwh/IgsN9I+aDZidSFgQTCyrvc/k
pBjogf3Ysux+pz8TLCXDMqCJMQBYISAW+v/4gPswg9dISOQhu6llHY4M/NV1YFZw19NpQHbieKOX
Jb9FXZeyjVY849J9OKEGw4vgNbkIm6NUKCkVkB+Qk2/cAmw+s8aiSxOa0W/lKmcsWkUnB5AqFpqW
Uma26rg+FaveDVF9zgVHCJkyS3Iu63ddMTYz/ENwrAgLwVUhG3HjAeS5AtAzEVugt0STptc6nrtq
GwunpmGYjKXDLD+yHH2fOCiOrjp09cVVFKfTAZJ5KKQrz3NTgVFke3slF6z1jvCevVHTmoIib0KN
Km3ksGH1251G1EzzNvegOmFzGtcA5EIuwd8DmE5YowylIlJHVCM1Ln4j5YZEBRKz6g6U84rVgf4c
06ZEtEVv17dMUECQe6pENuZ/DRz+wqqdW3nnjSS1oorHbsEc4D06+svBpUvF7yQwqnR8ppw/pnSK
uwT977tHtR6y01/dW7h8pxxbmMcMKYOJtlNrl6slHCR8PX3FYKUP+EzCrt4PMcMMAZ5P/2PMAdFu
nh5fOzwBDygAbnmM1aNq1PmxdvS580CnDWC83yEWQfG/u0qtWFgxI2QE24IOKACGmbzRdADLfmKX
/8cunDqqXjy8QmsYdJokbiEqsCiu+oUVN5I5Icgvmd4LUTTl78DBay9J9mLjGdSTxC8wbf7JVf1A
/iAThjQllF5/Umb7fkOl9043ZE3LAtfwNI2WXnUWgEU9/37GBIVbNTSUiFLhNIuGhlKhfJHt8Svg
W1tKlZoU1JL+oM5FPRpvxEw5E5j/oIxP0juOE90rnvH4sSAZZRx7EDQm5CoGcTAbukb8dZ068kXc
9dP1P3Enf7VI6XLozBNwjzaumrR6UPKtCM8F3oE6RuMyVyZJRBcNe90nK0xyUZY7HYOn441/w/LY
/JOrBAehLmRP1pag0IwmCepqhmmSU7pWKh9usZ8+qgBwLHhEWj+4ge532SzFus/3NvOgZtJlIraA
7MtHnoCTvVMoEl9xP7lFKItta6dDnEg458o+gffBmO34XPjM7EHpaqfxOoZlZpBupN6OUj+r+M5w
SsrbCJmE5Fi6m6nur2sNQ680BOsHDovWWisBplB4tVKK2u0EqcyZuAQCvCFxrSEm7hoh6ZSrXlxE
/rZ/xHbE9c+G48DM28CafvAi/EbA3P5U2Rq0aILunFb6ZG6Wx2uK1T3Yn47zZbyFMzFuPe0Rvaiw
T7gpa7A5U8Wi8GD+MgoFW2mJvOmf5WGYXVxDTtQGd06EXJuOpLRdn1AMm/taq1r6j9rplGar8eye
IWqZVMzs6Z6jHqq3yE1zWMs/sIwDrQOajd9ZJVGmmLZQgMtLg3WqPdbvY5PI7vwHWFWEswKVNdZH
7ohSFEUOKHzVoGJh6cue2vSbvmjjKU7wvBCs6J7V/10hfRDfMXetEYsOGFCj8w03vsM4Qmbp88yg
BNtQuxH3rBTCYmz4bt6oleqbFrBkr+F1cgHuPgq9n3wbS8xp4Zjsf1p9tf+HoXvjqK3NpMJywqKq
/xjaxfBQgTkQO+f6T66VvBTjSmewiynwGSLp5okodrU4J88cXaF+hEztO/VlUxyydnD9RnNbUHny
2pa1NH1NyAgoEAlavtDRavzZUhhEpWyedEc5mWkHoKjHcKtC2MBL3kgJHbxPkK3bdEBIL3eeFqJs
VaECLaSpQeljrzS70pzSfihHEQqmVxT3X+NvJNcuRWCiNYMsYbLR5YkKC8EyCPjUjxdzFMEbNrpA
K9NnnVNy/rH2MGPGZgEtFocoDL7zJe7rhk34P6gA1HFAqflpASpjRSki6Rw2vdJznf75EuDkHymx
hA3PyDadKGxx3UOEzFgUwQ6aaWgdJGxHqblPPMQaTUxYKTgVeAIpqMhPqaOyrPAa1/G9wIbghZuC
DPUCeMeFUpx9UVkDM6Y11OSi/xRPjU00AclsaIl1JBI6/IufyeomHISSz/KgYasNK8xcS9++vQCL
H6Qz7MyymBMIuI5+jQhvCaYgE5LK6DRfAbycpD2I75Y2pi7tne0lVZwD2UwEGLTZ66ZzyUiCYpw8
zpfKL1ZPuzCtbW/5qx9CW0khd0rRBeEtW4MCViu2BUuqa7mrXmufiTuDXM2I62XSWZQXuCyqZLFT
ZC6l+ydems3Ntk4pfAPZXQlOMBcn2N76EeVPLaELKjhOeRXetLeXNKEqhIM=
`protect end_protected
