��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���#�Oҿz��Vl;D�F"����*%F�����N����xL�(��Ժgb[�0*U/�<��"!�@��A�:���Ŏ��_���1����z�p��s� �>s�jK):�լ������C�W\�}��|@>�1�;z��ڪ�8�����S;Z')Q�BDȱ����$�[�Z��eU�C��䚒{量�C[�tfY������x���U�.��ꇟ+)���YA���.���9U@ԩ2`9才����r4��ʌ�n�%u~� �����f�ߥ���9�倠7��H����z�痰���4�kqzF���U�ꠇ���jU45��`�cr����\�V	�-P�p�j�9�H@��Zwk0m����.|P�v��<�TN��h�tM-�ǖ�I���u	U��-�tbGݖ��g
h��M�zL7&S��ʘ_�M|7��I�h3"2[����A��D��[~�0��P��
����n�r��V��ߤ�}��(��=�qO�k;ܺ�waړ�x��5'�W�C���˖8/B[�8��M�Q������F�p0&�/χNz�$g�@F�I@5�U>�o��*��/�\���%iޱ����W�ȹ�����7vr���v�p��%ȡ�����
�F��1+�����$!b8S嶎���0�3���.��v�s{V�zR�aο�d)�1�&AC
��p/\]�)#48���ir4�z�!���2#R�����v�A9����6���l��`�����QtfLO�;I�����|���JC��3�ޒb��C��u?Z���t��D���W���9��g}cs�N������!��Y9�?	02ʌ�z���-�q��vğ�Ǆ�蔩>�-&��}��=���˚^ݻ�&{����K�����	��Ĳ�,u"�b��r�����rјwV+�µdG��U/����xﳕ�������B���W7��\�{����s������.�%v0z���qF�0�܀R8��P����c�カ�	b�!6�_r5��N��Xr4�K]�HC/����"�\Ya���eT� ɠ}��'뫮
K��1O����`��m����Q�m�uEj��{S��>d��\���ۈuw�f��/ڢվ��P[?�����5>[o:/
��%�f$MH���s�g)Nc�fS�`w[�b�y���0���K�V��o`�@8F���Aު#��<i��K�!bbƨ)�����ɸ�@��L��`�
Q�E�v+�-=�uA��דbr+
n�{�Dy���\Ãe�+������D��;e�nX0��;Teի�E��	��iPkI�(����;��ӯ1��4�JD����U��ǡ�NѼ;� �`��G+ ��Q���0�Y�S�w%�n��
�ι��U�*a���Hn���N��t(�=�˅GPs��6঄K�b9��Ʃ�g��*�h�{��2 ���Yz��a��Jޚ���?��k'��W�N����,�Z�ãn$$L�U��ۙd��^)�0�HO��&�D�0� �W�Ä��K�LYE���A�<�C��y6 ��;i����