`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
R7IQXoUsWbZFZANcwqR0E6E5zbli038zPJRKphKXuQpoM4R9e1oPESq48u/uTRggIsnpj3NEJ3Fe
ZLcIBNcIveeRaOWjBRfsrRzo0dHHXqCDxK00JWvn4jT4eoPjyNKtBxP/XfM+BTr97Y0OURll0AdE
S8u0iBVq2w3xzCnRj+fQPHIf5J89RcbmyPWS5VB72trDdWn0fkfIeemnnVmuyDQLpQY6riMhA6A4
XyjYhSRfBmtv72r1tV5YC+Tf93lHmodR72ni1pZWwQDax9nbKSjVzD1I49JrOpvbZ+5pXpJABI3p
Wd4/OJwqsfGIquNyrYhuwQasfZNxUx3OdRAbs05+H/P4A1ou4/irxCroriwQCeP3auQOmUUISXZL
4wI5soPlm+3RnqDdA3OBPHFk2l1/nUwc1DmZYgQNnQT2vZll6S//zkVsUxp8lKWxnAmbMR9HMe/7
35pzPV7OX3a5/8P7xgVeH3GJeWZnmiU7FoFgDvoMTo+Lmo8stRX5nVjNc9fNlmDPWHofeDwb0st1
bE1d0VFcY7dnEHOJ+ca2BDxczbAeJPrwzECWs73M5XBtAiMH+c1hS1+w8cJ3t2g+2DbXyB/X3wm2
AgYvPb3nPqPalZVoN1ls7ktyR9N/z5ldMGoHEHv1G0ffhCEm5cgcxg5MM2CPBy6nOG6Ccttu7qil
o855NsXPGfBb3hDCNEtthko3koyUlzsGj0LdNee/YejNtj+rPK9sC7NsX7w+8BphP8kNQ36AinJU
wXBb5jAVhKvESq6ryvuVlhSeVYKlEEnf/fXkzbBUMu8x+h2in6br5b5bRkmvzSB//Pzg06BLZSY8
NfhwQTvkP93Q3KG05vSHlPc5YGCLK4B1p6zjjT0sKXE8cZQnb4Fki724+1oUpF4yRjGy5CbdJ3wb
H45OpNvy5PrcGSUBnnYiijKHruZzyO96Dw0ytHEnJ+vhVstmU/GaORaYI3qgWPYjPBLSYxY6HTA4
1vau/TAvdz60JwZJFMt92FrIDyjteEDXiK5vjHSOFMQxr65kUe2ZwGjzSXoAjXqzoZOg1h4twcBc
TFu0IgjC2OF8IItB70JHHXgs1mpQQBv8Qx0UbjPJYMQjlVysG3v+TTniXVA8XCfQPWSOwcm5osh6
WqcSS+nmSdJ7OOGXuF5RzhDp3oYh4ft2OY/9nn6wDu9oLjLtTPcGL2frLDWVNcwNaucTp9BlQHqT
Q846UxjoQ+H65TH4mYZKJ+e0pQxw2dt6NVbPfupFv2xPBSNd9+CSsuuzMmFep5HNtlizOSIlduUB
qfusWikp0GU7xQkI7ux18ZfqUXHWvfxwS3EyKvxr7aW2xn8lof17cLrEBiuV8TiqMLbzUzNDk4dH
yh7/xRDVgqrtV7kSPzDf1sKhmN6AuNtrFGVLQnMuKpXy/1r4g+62a0xHXa2dTqxKBvnr3iZauGUW
ShMET96+O+VXVwRvsbV3ElDNH+M0RdVO7aEf20mQXFiN6H084cMSrHGHPHEpcy0zW3Dfs1kJfFZv
+kiXUK3NgbW4HQBjoLbWwIRKCQP5N/l9/r7yASpiok0u9Kc62JuBzubgsfdgdm4yazoZzwiFtXYK
28tmYe7yYVbFAc5QOWY/rwXADusZk2oL/VbJxFYYfgypcUyb06D6tdu5CNSwYGGedltMA5p8ohmD
W0gKL7k71Y46lS91CO1EVDcdEzNxOffzH4/f/hFQc/QYsE+jwNCCSzImdVN+9EuSNCd2wLned6nm
sk/rQdvmwkadX29+pUS8u14k8dLSzICDh25YkkE6mFtAtcgQuLtSpgNJoJXYz5WhmNcYWgWl36Ac
0lKMvhO4yKztsmlfEDvk5camfjI3S6AMlmAM8gHv0fTBte3nEoA6sBMjSFck/h/nBz7uyE+wAY54
R+f6EVZXL2vdRGZu4Sj+CAvN41DHJ8Ye9OiDvhp32IlsDwRxCWkX6iee+Co9Eq3RGsiveHLvG+bI
VCAkmtlWbQ4VHLs0gGcNCY3RfLEXiRe+NCKa2JbyxCceX38+BESJUH5ALvxZ+z62auCVGtoXPl+4
b/Ln1xY5FJKIT8iWq0CCtbvQwzBb2E0H43/OR2zw6KEF56Kf8gNbGfxniUOoUmPpkMCBnm78sQ4u
LWzMjPZoPKlAGj4vu5y39tV9bB3mO1+DwqiQdD4ZVwKXD6b1o7l7kkSH3wVf5ZjE886cSBo4Aaza
YDejFmACHeuvrRFzkphcDNqCiz6UOZh1CPc+Gdprt310fp9Zeaf6MivCsULj+Q1JGKUVe/+TAtc2
5AaY23u9912PpLif7mQ/3NiGUjApeMVU33xOnE1eyTGur/ZBwbcNmI47EQ//ubJOtl407/rzTZnP
KiZrqfXmhledck8gaM4OIchT6MkElKeG3Spq16h6DRi3Q7HysiOqJwGTlft9MIPXhrzoTi+gNjZ0
lgK6eu9rrB67Jc1hGoCttCzd1JnLjcacEs9K+nWTA9p/Zafi1dRrVxHLNe3svnmB6OnYFLDMeWXx
EwLzhYYxPyyaitVQYQvYiKHUx0lvyPxW0fPUDuQ7evVSgSBVqpWU009wDapT/3sqZksWK4yy875F
h8fvis3PzPgpZJWCYZGzsTkkijnKs6TWlsoRuDmZ8YJOD38BdtcEMsWay1tAX/+UclbktxJor5ai
z3ECjt2AkPZZPMeGxKNU2xrmsuofuCjeJU6xJrdR0bdPtn77ucbPfHSZxbVK0EueFQppswQeQTsN
lUvCKExNrypj55SwWqK29ARm2KiQNAiIhemSXvbI/8rx4zDeyZVwTbicSovd7/FzpTwNbrS13GbJ
EHDSGU6WndZ5KiKGJ72t1H0BnyBkqz55+KO6+fjedx19o/tbcWdTaXL4KelIEOwGPGuuNambNndW
oRVYhh3ZrZQ5C0Yd3bJNU983eZSJ0J/lu2uSgWv2GJL/PMMX7mWqfd2ZRq5JWepBrvfjC5WinZ3l
ihohP/phBxxTMS8C4V7CmrZe/ELtcR5SZbs1FJPN/F1+fur5Jn/9qRWxRc4oMjuIaBp/H/CtjTpt
YK6MdEV+riE0wULyS0xIbKOetn6Yq8HyWexqMeSCJey6DG+AECyIUhm47iaRoGILMZxFWivxACdj
C0bCgujyH4Ju8bMKSIFLX4Mu/cDpSRlIieRZgVLV3ZLgYvYNrI4hqnNqmYyJau/+KGR32w3QNYbT
6JeDZyfyl9swxfjLHOOp+8ofwtOirGbkG601GlXj6EOwKkovOd1FKHEfEvSMYEB73IlVzpgrTvpt
OAqCG2hHbp9HSGpMda3Q7ZGtwF0H7A2awS04t69F8C3w3SrVN6s6R2YqfsXeIz/PGLaEKXqJ1cuo
Zs3Xu3tjN/SuBonu0CWjQZJKK1uwyODUyg1GVKtttplzBZjRg28xf2jX7sUFemobzYeXEEtFAiOZ
nQZla4WXhLhs3qwG6r8zCi1MBSfbT8WSm/Rrfbs7v+d434kg8oBADnmR8K1Pbqh+fo0UihUif912
1VCg1NCMYYObixz0+6Juhl0iY7yCdFnuJn0Fbx+cZ5/YhyrO+Aao//4ICZLXTmDLuF+jL1rJzMBD
jQt3DBZRbbkZ2w5YA8614yKttYprZKfyCm0wesfwX6+Fe6Bkr0HoigUV1FOwKnkKja/ms8tfS184
a8mLXRztdYg7QQmBTGjBOXaTi9XCsMDlMSGktb+k6LCn7Wtrsdz2l+iL8UIBowU+N+CxRhBiJn7i
VigSLwvbEF3I4lUnIZYE69R8Zfx28LAJ7g2E7/tfslBHjhjjepKZqeOtIAYy4UBZJo8MHkrsOEEv
YwcYWATYy+7VB/6tZz/aA1Jb+dTSStXsjzPkQjxEghmTi6DibEVPmBSk3D0wMwLJk6/tH5DKVelL
nnjea4cvCFHZ3O+IZ7BPPaUWjAdAUJgqs25aWv0DQoPNDtijyY7aB9wh8Ybi0RA2x3eHoqjSKClz
qJ4M9sYUgAI4OFrXiIIU3hLnxmq+xI9G3TT5W1yuQtJ9y6M7TjaNjzgSfvZYeBFHPn+NP7N4+VA5
1eYP+d45abg653PnAZ1aGfFpI/yjnN83QbDYDA22TvoqOBctQ9p7Hn4SJL5rJ5M5waih1RD4oA/k
u73oUKYJ1D3RRGe+ymP/ff5jFxHqjs4uOYeW2LH3VZHCezs9CQDMH9aefggfxYWyoS+zm+SLsRDz
ppxMHXzqOD2Ts34swCqjKZnYYJJ1r8cY2h43wUxHWYYp8U+nXqwHACbSS9k/KwoA0VXX7rp4LES9
nw/dC8G7PzJOqRQ3GWOEF9Ut8bmLGe4qASFQsmhLH2dWz5x0ETg1TSXz9Hmd62My3CxUEZIP+n1Z
cdA/hi4fXM1t/Ns9i17sRLSlXelgwx0i56RaeORW4w3GYHYwOpVm7VcUdd/VVsivS2D1WW/NYXK0
s43apFu9spM6wk5xJUC/r+0+wSQrofNpQFp3znIh+1WARUS65/Amzba2LjUl3nqgMqEOA41nYvh+
3thoTkUYMciKeTrhKfJzEJvHffJLXHxFurLqbsW6V0ReajvxIIsdUFUjp9AvvR46zdSsfo//iGI2
/U13klZsj0fJTnQKxo3qQmEMz1XG5MFzPT0lSsFos6AXd/eREDfi2ccHc4740YZ3MRre8X6gGhZM
bORAZnRk/8QiOsuR54bJjoogUrGfO2FmchV0uNx7YVPlX3n0AhVEvDCYd6DKhYvvCZ74YOvCMJ4w
tcCgWZv4GougVTTmIsu3zpXLxyJHVfmFxSWhB8swUUPcyiqTpJaw+utkvevt3zp0nhSakdxIUiu1
Y95TVAQicLsLq2I9H5YpTS9laZr9WWqATSTJEQm0FSHg2JISyrGkafTalYH5A3Nk+ipvN+W7xQ5r
EsKjurMiU17xjjAW3d/3waW3JvGTU9/J80DZarlJGShpDuusub+jfZJv4cSLbR0jthrrU5zed/+V
sjI984aSe6nb+R3OdreyxU+vuTMAVBeHgZYV9E9pZlU4SKoLqWjZ5cjJV9TeCCv0bW3OBcbTb+k1
lWF6HZ/GLzuX5l25oRkWN/0X/XPtzQs3qzfk5OFX8apz24it4YNYllZ6swIbdccONF2qdtJ0pkSM
ukl4q6Gu75vbwm2bBlzP/jkc6/63fE4TgDhz/IA+hdruLVpMX5knPbamJT4HEqbzQHh5pcmbBIo1
tXyRKkTwKn/LsZ3t4uh1kc3mbaBAas7uH9sT5cVNA7GyYjDFEyjEwpr6U20qcNQJEq0AfCaKWnVd
Lcl4h/X1q2yV3zna+cuDAojx9E6TQBrPa3C3h9Q2ev4XLKY/rnAL3bq+na8IF5qqfMraaEafOikM
WhRJ/K8vXxkFEp3XQa3UCVU9+R53BjFbqcjUpx3WRHjYty0ZAhjZbhtyvrMlqFfrJOA8mIn1fQOd
UqxZl2imTouHi5Kvyw6yRdNpX1r3CUwUIiCAi99NYsiBYGpmkcCaAQ3E2gVTzO3KnwDIoU6dKnBR
OhK7dbVT9RmFplfpeCS6+sQtzus9z86q85MKqip3G3XSB08bw2b7xGsLQQKQttVw5lnd5rE8GB7i
zSyOUbpfe7aTA8tm0yB4gxmSIWrH6M7sK/79qGhze0RpAUJaQKVuZDouP4yCiK6mi40FrOdcrvgw
E/GXCwo/TtDfvNR4FAfP1qebDjI50kyCw+G/We7kLy4gvTDfEbmJUHGW8Gvmln0r7YS1qvpGcdlp
CLHRT6IjO1IH4kk0M6P/jw8fILDNsD5vv6hcdfH5sgDPVMyOivPPbleOtCVmbWq7SeGCmtCkJ6I2
Lp1bijX3PtxfrRShyD/ZFQqkLpqsrCzlFiDrJCUcif/Q2frA+l9ThuZ3gPMpO/VQ2wZrGZliwDHX
D0TAZyUBSWY83R8b9oCHfd89bJFLSoig+oJ9wVpr8RdoJRMCMd5dAaHGxh1CbvJTAhDDeoPWrQkr
h70mHHBzhxo0ILYI1XmZnVdlC8mVh9vzH7VgZH4dG92ZScjFb8SLPLDt0OdrjJ8x0l+DC5r4xzkO
6ZhjCpSOjROpOyAC5DXfgvY73MJyaVbecUKN/IjwKRDGx1WMST6LMsOKi/Pir8KVcuaKiIWhbpq3
iTQwQNXaNIGqSUJh9xATVCNQuqLrQYYeAPSAQHC5h3br+G40WEtsAIyJjuNdSXwxXp3p1V0hswag
McQ0XxmMkAJ6WKjlVKZ4IYsrgVLKnCaqFUKu+Cd1avoIQudSvn+i0EFXBb9U61xuwUn94zDQ+2DO
DdkI5qYs89u8NJkhJKqh98gi7w/hzPK76gEWA2S6QW/hTrlQOi1qvc/MLYR1nLRuQbL4P4n0N2nS
yNJyVkZuWnr14h4jnOXK3iR1rcWEMIyiG1b1uHxs3aNsS30A+SkqgP11YPJaTmCNxaxFWRD86jm7
sbnP3QVmiRz5ycF3O3hY/GGbAdsdG/bC7wWXb8yXQHUz3Lg2BIxWhFuoYeCyiIa/teOMr8zAOUax
rpf7hgWXkqjgLMQEKHMJbEKqp+PS1Gpfsutnq6zUa/WEF2islHv/TCkIOqOn/knnLwaXcw/uKbi/
YenL3FHqust6eIDjHzBzZRsaEhqL6DZ2TgnVpauUxHqh6zwrnOXv5+T/QmWSN3m5M2zv+HZbIj12
0zrDJWclhwa7XMrhe70VsnvFLYiMTKL+3nLnilC/GJr64HGzdI3C2/h2JKH3U664pfF0hwEa4SCS
RIv5W7eJHFfY698NEZGyz+pdWu8dtozwAFLxaUxrHlVmGrJE21yneHHHEXg8eEPZtX/iazohSTFC
ejSMciT38WG+Kx30O+Ux4SLnJ/1t/Orgj6Nr8fTW+r34mcliCrnP8hZw8lIQd7CROhlR//N05rXq
jbAdSx7O1iFN6UOpmRoVk+E90pkiH1aQeJwiMEbQ8kr/sAXR+xqRe4ZOCnhPeOn+rQm1sMmQYBX+
vGYlmBHphLZUwwOL6p1nq/xzpe3x9KJ3uslnTZ0/+iwRvd6p4XZcZ2k4VKOuZztkEorauDqUhq88
0kDemOl3Uabte5hj556d9VdjWvqj1Ug0TCNRI/CUSQXa+m1Wk2jbwSiUy79qraks47j9JhDvjxc7
gKYZLQGFAKtlfzU7ORw1h7lBWuJFskLpZggzTRf7hMmIvMoOFlSRlh0ZvSp7KgePeVBuWFvHWoMC
wD/xp3+8Zj+ZJ8YOi92vLJDHYs3wXyR5gi39CUQT3HxLK7ADam3xCSSTyRBTkAdXRYswumVocov1
SYThgUtdRm/oCW3FdjuleHST0JnHVFIACOL7A09vPIe55CK4koBVP9rYByxfKX4oaLf7GkaqLThC
nUXLgtCUmgV+dYT8XP/Mt6ei/wTCUcRGIJ2PHgvtaCvZHJto+6Jg1oplDAD3/FqW1XcB7O1YGZS3
4Xmntz/F83LIucdypcoiYy0MaHE9x3kd0DwC/8OF3F5f7t5bWb/oDtJgdYGI6ofIsIVfS8qCrT6p
Ad6Xi651L6fx1/QBbCeEwrLtsa33dHY+5vHQsVuHIfROlW5o29GvmFHnXSDpwjFOY46R1gAWpUb7
LddPw2ZYHonBG0V2kHC0WTjyGOESqt0ofEcJcmQnpES0b3mvvuAKUJBY323DcvJZMcQJts+c/y+l
l52toVF3nJUJRQfI7VCdHMGO2CIQliK4abgU4gK1wb2nl1Ydf1ruqXxTNhL68OipUsES1Im0nV9a
jrBXe8XSor3HYFwYWeLXEM5D7v0Wpi06j2phbFNSMLWaX13r0ZHMHjC4j0HC8y1NdrOPGpwaxoj+
Gj7y4Fl/nVp9Zp9RLkm5PjIhmvCrfg7Eohu7KKzduq1wQcXRb6CqA2Z6MjEkuBbkiFsQQnpviAcb
7h5iQdsU4nt29gtkXg35iX90MetQcOW8ivzXX43dIlidPe7wnOFqz4iQsrkRMRp2LOErFZKpIdqg
izhLy1Ww+Uic58T4AmrrdNP6p2SVNDDm9AiXHbWxUMdrznUdqyud9BFQiKz1tcTI2NzwJy/ZR9mf
7Wt0F7QfCFoGWZwcaYbx15fvOzXYBZY3MK8mh2g8y3EXe2DDzkWSh8ZEE8SLH1Q+Dl2DmDlQsz9V
9xlXJLPAHviTRDa7Ul6xrtUbw3gTI/EJeqFqwGJQG0SQ7Z1Btvy0gfdnOzNzl3Bt/sTPZ+V69vEG
KIDK/kl9V9i+icPsQxo4hWIkFxvR5c2hwfojrsCdiAk2UovwRNcRRF44ln8OqouKX/IrSS69fnu2
rglZV/rKe5NtCrg9ZLHSHJw4Zi7w9P5L6Z0vD5CFfGZLh5uJi0a4dE7rfZKNimZ/sB+2O0IQRPHi
BNE88iUxSqbBsvwmOIINtl8AzwpKbNboSvJHMNhBpYiEkTrODvOSRhFBBvdP0IfYon+0DdVcDcVe
xRMKdMLi4vqr2u6KGrs1UF04lSQkwzEgHxg3IFb9goUvyeIKEDyKbJiLmnQpaVPQQoi6LxVMTlFV
hvTCbH+ZXtyvY4oerp3ipdF15QqHdpRn07Wx0zok7X0HgvQxENf162akIMLDp0yNP8D4WhjnM/CI
vo2zgMWIGA3wLak0Ge0NVyEQ5Z0GgmVn80gLr1tW2YoS4IcYkUBjua2cylQDV96uoay24pZ4IvEi
3UgOFgtpQLJsHqW/mi2K6B1cIpiual9y/yDyGFuMjKo2JHi57LfgiGQ4br2vJRQ3xWTTN9EEvjfB
veRPRoSV1MiaoWsuwGRXjGJQ/BxDtrcL4dANxD+ZgiQtbpY8fjmPv3WE8uo6HWHFzdYiMbQtNd1g
nwHj43x1KbJAp6q9tjAAVUKQ0smFqTCuiDZGsBrI6Y9WxITEg4VTDjRWOG3MOXNlAVQhCC4nfpcg
WHDOw7Q5l7eGmioamdbQ+zc0FulfWSRlVr50O6AGm4l4uvlmlNB9d7M25/VrMMYP+7d08/s+hHsr
LqwFjrxer0nsjp5l8Yn/VCxHxy6dI3X2iFWTIIazwWr60EcjJZLGwcZXld7LCO2pVjC07pQXO//m
4mx/KE4dgVODGY+LCrKD2g/Ee/skbjKsURSRVxRIPB2/JUnO8SzBPbps0+2+J6kG38TyayeEOobE
g83M4UClntlWJ8ijWbNsj4xke1D8v6vmfQacWmSLh3r8jqrPFaTBg1jlwshbEjny9QHhRyS6W9mn
OmZg3D4CXCUHdb/+Tk/bTgSwyQZ74PnFKczXbWyoVgV1aPdzPM6YQgFvdf9jhQl2xjoH6zM3ovSB
G7aPf0j33wjcu2Nt17nNDzxXpA6K87f9tGqi29/rxMkrdauKJOtxSjub8s/CtYX4Zxbcrx5t1U0f
PawTE7onLmBsaIDJFDnC7RGyROsCntZ7Xd7q3z6P7ubnZg7A0+sKOOZYO88SuuwJzHv67eFiyBlb
YcOuhfaQDMK8pfmTZZjPgDu/4ec7AIzXin7/2uhFWIME4TZMibu2z5av3pkSdMI0/ewC0gwhIy5g
v6dTppyUQctohCansuHWocG1/xVtRf6QWNQ+/Sfp+CwylAZOvqpPBSVI7iezEvmN/pfaf2fAKvrX
Zqi/9yXyPipbipX+Gv792kcq8XKAyH5vQ2Z2BVIVnNcyswhGDUTrRJg+Pk3f/oVFpkU7YI3GaZEo
MUj1618qYBoMbnLGGa3R1gfOqGyCYQmVDvjlcHrig0NYv9igJsU5aqBGCii+i3mb/GRXG6InD9cr
XAUmRv9GipORIjjGoAxw3fsfvtFSDvfYQqTFqLncWpsJLaE3+BJ98PsY9TmugdLStdQ+TlyxLZR6
CwBtUz3m1fRxRpheuJdfp9Ft/Zp+P5lPxUQy13DhVrG1hhV9o3RrfMwIYnxQzADDaKINn0x3r3xo
SuJNW5e95ZbxQUrN620/AsjgHFtkx1ym84dVhokNeuB7qt/kJBhnMH8zt7yK1QpPuqk/FDRKxm+f
lPFce7Ibhtb3EhkbdrUs+5ysJP+kT3mQrlkiTw5NohMPm/m+HzZS5crZcAvPHjIBEZCLOQYLzTo0
P70bHLRcEAYdTTAHYPzG/yxLsXKe7jc/MhTN4QpQ6KiqD+6aqxIAcH7ftAyfQbWrmhe8NJbpi6hC
JrcaLUZ5n6la3FdCPLMJBYnngkbWfU7oKRT8P2utQSZ1yNXPk3uaGjtypTCSamKc6VPu1mrU2mMx
3FZlkWR1INJ99hOuBa7D1tjTbTmfglW6y/onkb/eWT3biPsypoE8EWu+LjM7Dl75n2OH6i269vmZ
XtrpWuwZuAdocSpLrMrXWpP/6FN1ZpRq2uLNAiQZimLuIDd+GrSPqPW60Q95yNml6KhoZlLMGstD
QvyQHGkjXVbo5tz48QU2Nd/61Mpozm30Wh/JhZMrO40gMbJaFVCcOT0kvCjpEY33220ZkU7KrkdD
U8fePNSMEzAKVVYB+QRwmFv4D783Z0I5MwUovq8QRMr8tDVQaDcWurxNqnLOgzLsGDQzVtJPDYLc
+F+N0m4WQA/YFprDcr8ABTmgf7dqJqpDrfibXOPkQ202oViExFTKzy/OWXULIk4ARtM72Q8e6bIq
N7StzWD50C/Pdi3TVw3RVUEp3HNyqOXjaMFJMlI3Dmq9xCnjMN2e9KGpeQsRIfse9BVq0yEWA+2z
gJljnI56/F65Foj3ztapqZsZOwDEjkn4I2Fefs3oVaBFo0z4675QecJpZSepAvkoRDwnW5wz4QCx
nPbLuKL9igPYt037LX68lNzCleJJ1QJxn+w7dm2kQDAlK6lex/GaW5yAvncC0R3LeHq3MjVRkFsO
eoC4rgPybo/FHKYxJAKP1ugP3KNf4HHtB1YtKqo4X6J4aTMjhnxQSVQGlG0ADWYT7/NHNH+SPZ4S
WRd2DMEXvNBJcmtL7Wd6BNrLvcK/yxjEYQKdp7LZj5TRFaXasy0rY0dMuRr5nDtxdbmNWlS14x+n
n0ytWcJPhfZglbSigxJGypRP36Z7m+0F/X3Okd9n3ob5JO43EwtxRA+AlaWJ+jTiZgiaNWVpMf1n
BdBA40F98SdnLUEo1iICzIe8ajKugg+sIE+aPzUDHSPYwKhMp6kXXfFULu4Pbh9NNMrYZG9msEkn
cwum4fge7Mn1SzrWQgaCLS6dk/omTtHOzjh5Mzp84uVaUIpJ3J0m3E5Rfqa8tLjG780okqAk4oY5
A/5J+jsudHTa02f+nRxfDvQAjhXnCtb2W7zWYpo0bsHwwv/hdFud/+dkhFkcNQKxcxZ6chDQ/bpu
N98qcDTOZfJvjDLQLtr1mb2DirJ9Fx66+dmd+5E2w3rPjLGPeFuEItT3OkUQaea1PyXkgvzHGQXb
cINtTh2NdU5vKQAwCSF7VeUKkdkcP012p4VWDbLzFzh5+P0X4Vc6ATbV6yN1jy7OPU27gE0KFgrs
tYGnP0xM5cvmjbGfyxMbDAieKJfSy7hAB6z3KhViinn9XKaRdzy5gAbDv1E8LTb3Hwrz7fv/iius
UJ/GE8HUKIoPnilws1IIELenOSHCLzmDeAtxZ/QNWomM6P6DENDhE1FgvgBJt06cs2t7BckeMSIF
ftqy4EriwM9KhESj19fEd474HEQeWDTX2AJXXG+WFyYxn+kQomGSeuKfhewLcTcT2vX7ns1Ifkz1
feaIOGZfLNKBEyJZOno2/hx+V60UitSi0cdCG+u9HZQ8izZ8uDizPYAFSnNo/qcSVgHrGrDkszdj
UppAGiUKQ1XLrG7vT5K9ttLXrwVvtFX9zrAXrAqrMrz6zMd3pbrFgxa7l9l7Hexm4hQ28MIySraM
X7E4YR6dv+hWyu4ZkwXi3dLBfHZb34mtl2x2de1U3rmK3fZw73jkvOy69u1E2NHyIwEX2CDP/GUn
KoK7s1FBt2WS5LZw8GQQWp5OIrEIlI8db23DNWmaNCnC7sR46Ei4oWVVGxTB/STSGZDYcRAp0qLr
TDtAwjqKXZS2hmcAx0Be1kLwAi2eued8t3rh/STudu1ww0VeBS6cFdNWRC5SbPluyPVgiPUIxDZF
xKWLkUWQ7IePTTQQ46Kq7zt0yhroNvueRDeVQHwZLK3bqjeKg1J1BTWK5bMDcrtmO3g9O64Q7a4o
5xu7yZL4kUhHjWNG/S4gHCb3Qvvndh+KB3mAUpiW72ObttHzDb9gMgfH0Eo376nuJxpQx4/GqSSo
g3TzrGXiJD4dX3iUg2A3d4hhUTK2RmhQiMfrTlZbFhhEA7+BfeRG5gbvzfENB/wAvmunDGwFrVlD
wW8Lc+Q0b1wG5T1PylduLsH/grVtRoFiAiC1UwE7f+1rKTXnczaZzYYgM08pqK7EYLIJ+/P8YA3f
tbcAowMAu1Ay2+1z/ADdvDomVfhSTFD/zaVcvNIKsv94N4krLw8qK+Xp+xu5hLH+0RHLU9p4ecHy
UJ8zt36OkxUOer8EX0oklGNd+J2fUyXDoXm4IDXWA+LYiv8np86QTdJzate3l6vqRqqR2heoZUR9
srepC+M4nyAUeICoMVwAL7ELWRYBCmYOs99n/u81T35rxKJCKgaKz8cmPgZIlIORQsDZxOQEqK5a
Casu5WhqIdyfIz7wjYcsk9zYN0LS0w8hIPST6d0FjIvu2FCw87CyWM15xO2UDp4wcZx6UtFuIgVg
dFGcSvsVgzDPZ/QPkTinstiDDrczEJnnZuYH8x4FZVXYMMa6urh+HQ8RaTj8f5rI5eGOE9R9zLPw
edZMDCejYhXDME4k9GdhKTAzLaZ5ogVqzDArT+ypjePS/BqrsMU3psIkIkME+esp5ocQUvPdFfPZ
6BcKaRVPjywkp7qTIqR2AvRgI5EgO3nWaWAxwN5fyutUDyG3bKp1skoFjndu/tgt672c1/6olOQF
qRMWzpgcARDsA0bpM6ioCMbHo2j8RWu/LBfnRvsY3wUcIYqU3eQA3Yg6c0oAOYHYNP3ie5H1eCJF
qCx0lh9kEagLU0hm8Ko1mcRhX/we3LveiEQbtdg1TJCqQDFI6VnbKcMh1YecZza4Ct8ISSkeT9Mv
dIBqM6NRqsC8oFllV/BckFc4QXMtwCDTiOST4JmaaD3AWGRbgcdWcd3uG1YWWoGOc/mbZ15OmknM
DZEL5EwtpytODxxWif0Z9lFujMDyuKWPQF+DCSJsdeSELhwJ1rjAk69PpGSkkvbdEjcFsViusEZh
dIMGgENO4J+Cu1ZJxUTI9UUnD9RWOtm7gs+fLfgufrET9pBwajv8DF60wBG/Ioddxmon9Tj6eqVu
bmMLqKJdj3HjG48YMqkRc45AC7ZWzK9QlRKhIN3oRNu9TgS84l55+G+w2SiMGdMaRNmt8HSv6jFW
iijvoG6ADKRsw9yhEeTuhdxcmCiAgzxmUF/6uLJDSX1mZpYhBK4qkIlnek8cT/2Deocuz2NaBoly
XMbdTu/630m1CIg7ZzCSVpI2LY1KfEER/PWGrjgqZMXwIKL75jWFhV9Q7DTcwlBV4e766u3UQQ46
VGyUKtw+eD/45l6kD+jO7x8yDCw8cadD6bKxXn2m0IzB6PwLu+htZtkarnwcOM3PYxEFEZyL8p9D
0wfXQhNcdXLrg4dbjkMTUcJ8iIEW/uu9nvvTHm7r+niMF8+Ki7VtyK8jHLnoE4WkCOynM6ofQPUF
EoybjaKOcOdH/njEwj8G33f0qMQ9s19Oi7HKoAAQZZ2Kcbf7pjRZr+D2loyFbhm77kbOmI5n9Bd+
gfg+OS8WmCMAQKfjvw/Zb64cLF5wrAg+3cJkPirNiwXTM3tmBhjgLVyyZAUjWPvS1z58m4qrpOOm
UHqg5C361jby4SemHpbrZOfq9gSKAuE2zxP6EM7tyZtrQ1xGBGkqwHAL1h/f0UJk6ujjX4NkuAc5
Zg1Q/PS97sDZqEkAoaoqGTLZuYmYovD2nS3oKscGHyCHelEpQzx+yTIKCnFOOhQ3TY0cwwEQM3ON
fgMH+JfcA+nGbgrIHmEaCOz5fQ01MkywU81pWsXwg4krFqpLqxbSbUGsQ7SQtIWcDzRisgWZ0w8P
nMG1oDbK98oWI2efTLclefEvRCCqrZaxasjAc32vRInKO8fI3VJNpH2F1RNQZtFufyksS6an3ipG
fPGPpq7aQLP+SRHhAhjnqBB1WvPUUaRZ7ky8AH/c9AXcjSd44STCgevZAjrFXi4nRPPTPaPVK8fk
JCNYBTGuKgPSiJvUKUTIFTFcs0vW6nGE0V2aThemleUMG0OApuXNmmmGBtlgBE5Kle5d7T8cq82B
ovePLFs32u7hotVt+MOmlhCr0lhzQFPX21pbOESkMWXYbERjNSn9o4yq0DPwajDjR3O6HMtWbBza
EY70ZpYwivgQpiwydBu+axrE6jvEbFvu5aoYyL199NjiIR2m6xmiOvhSiPc3aQBIghIzccPI4hkW
slteBUBI/6RltAkhrHdw2kJocHn1sqaFxIwvbrB4ZJPF/zKFppTmE0LEn/g/n9rTlAYmuwhlR/LN
hO+7Bs8JTAGzawck9Vb9qOOdYovJ2wtKmZRX9cPjNgj4NwSlea+bU/l+/ZaC0KjY4Bc6oC92Dhvm
mT17WGDCnj6DdymxHp+JaNhjKsDj1wTRz5PqzeFT84SdWbON7B3E+JCi8WubpQ6yMy7O0kyel2aG
ystbqeUwvP2mHKw24/VJZ8OlPWrWL3UXIuLt57QWhb/jxYeGnwKSnu0ZEgy/o1qu7KJ1s76SJDXp
JUbQC58sbjjA04iRKi9qnQp0tMWxU5D/mFLeCj9KLSsl723ic6HWF8BMsxQBuf26t81Q2y4ZJjr8
azWoTuXcgql4LASesV8BM/hWZ9ZshIkttBB8um7LrMqzfhtCYnYMhA4eFGyDpxEoQ8L72nlHlvHJ
aDI4r836oMAU23x9k2SHbkHCFCM19ZXpM8CgPXAU1ChT4XGCo+1dAqn0LtRKEPy48rzB1CXr8v7p
wAus8zNoxrpUxtOw5NvVcphm03iuvQluSP2L6fJJoUlHOD/78z4rkEknzeS5RNSj1SCJVG6ZdaaR
fkOvUsZaez5DB0ngLKHEbCyRD+e+1aycFZPuVvcsNXseiY5ARke/RTJRJoc2XGTwTdWULQn8P2sB
1HY4cjMMegNRudKz5FtYodftycoG4kh/WOxccnHRksS4HkKsEp781cLlwmbyzG2ORBdKFOJ0iSF0
ZQDvAnYBbw1o11CZAkjs+CKcpdMPF/ZgloY9fHWPdBN0b1VnM194pSyjEVJZ3qPMQGQQ47J4W2OD
pgxw8lkVfgw7xhtXXifrJeRnW7uHzqRbAOgD1dTl12TNzut6k+F6OmDfBI8UdPnUKYD84jT9btu3
CWZv2JH+SmlgIXV0KpBzTvwftl9DlXYhrNlltZTfRqOL8427KUhg9EOweRsON77LmKWJl60VjPW8
2Jmcjvzah/SWz/1jdKVnRloK9zzbpTZn9lZYSJlG+ZAsIb3X9yTxiVmv3CI48BnS/y1kI+H6w2J5
EUO2jivJwUi0WX4QRTpukJ1JpMREiQSQ1yERyn25LRM7G4MP8WJgowOZy8H6dhyqcuMBdaraiMK6
9D7qFL0PQMJqL/S8zp3u4Xwgy2QdYvrQFes1tKuU3u8FGRR+QwWeRWqy9zUY0Hik5zT2Vmdqckh8
otpQSkqTR1iojuWORJm5Li52m5BqPC1iXNKyh5fAHEuKsP2q2RogeC0PtQH9lIzsK1m2ls/CG8T7
i3qDe4jieWw+Ush9gDAH9tYAIwi86p3Cd4oMJE/pmYq0AE/+XcB34XxUcWzbRRVfHxJ9MHDjQTRM
UTN2GFrn8e5ft08GNVNzMroRWwe4gsmlT0yUE4u3A80kdDRDsqStceiBep4x2piY/mqVWR34+ZaB
/GDnLhm6Ae6iG0+OqrNnYoC7AriwvfPjE10qlkCOfRSw2sSIN2XcW+LxHZSr4S/hnnxuttlh/BIn
+iVq2zSCshmbWP25/w3mhqXMabubIZhZSvoYSQ12pCcdISEcDEcdZwQCgwZ3FUCXnbA28amDLET8
ENl02L8LcgtE2SzFQ19bcLIVf0EoyCGYnMo8sXV621dB8FvNwuqAQtFv0bWvHf7ANjdG2hq97sLs
f7Wo8XRd44lW15aT7PuixRmZQHFN+V6FyPy2TLnEBVF7PEdyD6msqyWM4m/Jco/xzp3+G/JsMCkB
5VdGJ+3W4Ts9c01so21LcgW04rwWsgxQhhyKVkylHo/wnUVQAJmm+Z49q+6t/vfJ+9ge0vpzF2G7
OdJUbMIZz+IoIabxyEYdOWBCgViI83WFViZVHC7A6Hpwyd17S8FlvKX/jKxwHzfTTRXa2f6Plh4X
f8turbiX7WJwBH23tUTkGuol27TveuhvYPvX/q9R/8Z4+324IhR/YBHhgsjaDcv5pju1uG+eBlf6
8Yp9/01ZWLKpVDF+0kjmDBR7G25EUEXWC0/8BAKvcJc4H0yorB24T8ltzMuUVRCUNzLmJ3fmpPZM
MAeZVeSnuJ8KXM2pi821Cq33Ps2+ZviPZILvvr7ODL7fTFi24GXji6AeZPo8ZBTx1XjgOQ85W67F
QksDjYrq3/fWBe8rS59ZVugcLnMJjERKP066aRhvk4RVfH3e51eYvzOaF5r8MvVlp5vL+/BPKOsY
z8cfTZhHvxUUDKV0pXrrGcc4FgdywXIA4kRQ9KCtZKkTd/Qg878R3y9/vJX387D1Ryybu445k+HS
1Tpu+QS5oLY/L21dCfb/shf87ty0bc7PqncmFaem2ye7vnsgUXg64oHvuwRfgVEJrYifl2/n6Zdj
wkBCaEbUqFco/JmjQbDxbdS7KG1J8jfgqQm+eXthkRzVivOijld19TPc7Out4YA/+uNsZw3aoIJ5
jKJ/39F8qMrxUJpXtruLa6hrD6+E3KF6M/FQZmKzoY9ash5tAZXcib4YppZOy2o/FjaKodxtWclk
QvVNgoa4ujDZktry5cfhNI3WB12tf6ctQ3RT2MTkyK9gEnj5eWWgp3hNnNksHy2V98J9BBF0PMrJ
uGNNCeielcU/SFcKr48YFQYorx9PZtGXNMBWLNEHgjnpsqTt1AImncaZY8jYodUg5bKbIEw9qi9T
4FeeA0FrI7I3NT8vzXiCiMVZD/Aizg0zEqyxsKJKY7yt+k+ZJaPoHFOhY+w0pS6jyuQY/OSo53Aq
FGx4J3UAJvy+MPr3a/j6jgi+d5XU27QyXlTjUcRCWPysIZlKswX3BFbBtLRLFdNLRjS6WjWUPNhM
i44Nmbm66n9rWmskv/R9W8wVz+GpM1wrkj0zibqd5PrF09DwBADSm339sC1a+TGCMz3kJAnldOlV
CPp71/oPZjtMCowPQs6yVw8QEOignx8Ieip+524/fSodbMVArEk7kGxfp0ayxAJxmFCKC3wmL061
vdPDP1yPL5MLGkLYZ4rgMrN8uoSDj63d6RHxWMPguB7CEvDQzDVG9YeTfxJT0QwQsExXCcOsqUkX
8zbJbfAAxemWPl9xAtcjl8eKe+U+QaYofB+CdcfDx3ifDM4QCAfAPCOgYiDZFDYjwm9+mdqU7w7P
zrShgMpePb5w5aFYacltirFG+dvITuctqq7MYXqqrLhymUycldbiFh9JCNhROXmWykJYEzOIZ/JG
zLJZDGJQAm6uP0hLOeZjBvMHjzl2EP1L9Qu3O64a/QsqwohwEn5l3Z9+hquhHZ2UWKXeMQqfgJM1
hv/ABwLjKvBTb/Saew/fuQhHpx1lmc37qROmPZnv9J4eN6Aq2Ri1de4/ge+ucHMkXPFUQ+rfi8xR
SNZCWE9sbejY3apWXQZVeGW0378JV33aOFLnrrtJTUQVvTw3Q7Q8rvy8DdAtKK/YxMJJhEcITHe7
2OUcgvBsP1WukHERr688zK4d9EPM5pxq+TMWjYIfGT2LeX7j7D5VF4qvMc9kgt4iRy4YCELQjae0
jBM2d94H2x5tKTcr2pCxxVm3iuK2Oi4zBbAe8quV1JIYGn4VeSp2NLOm82vn8w0xdjPqJ/xKHZ+s
blS8uch3ILrZAlTB8fTZ+6Vif3mP/GXuO0Je13sxZ2Zr11tuACNESPoCv1ByFm+5d8XS4SF5UouV
7548levNZnV110aXaQbDRS4tKKUYA3mdzUxcphxidb8PDVfVELewzk+j7KrP8YHppr+tLUVWSi4+
GRGOFvBwC3VTLDd7rxb2ecDpcUqc9zBZy7WQapWMRPgwXZKfFFUU5r9470kKG15NU05FcFwTr8bv
5jsQCqKqPj+AI73hXlf97Y+okiPKGS5XFYY6N6uUBsWmj9sQ1QchKQvWDqk7T7vaLpM9xA6WNiqh
kOP6PTfPkTJOYVHzD5oURCQkgWXb3kzddvSUTDN7yR7CuU0q+pMfFmR9Nf+ijhBAMXT/0OdOF1Jk
gylqMB14LdB9Ak6c2cvyrWj97iWlnyYAoaJpzwk20Cg/bVxGS5uUHJGXh7dJ34HF3FJLNzDNhrR7
phKc/W7dlyQBBEAWBXy/vIC/iQLuR7XT3IuGbshTx+QEdjDnavaXMAZ7m6BbXeaRlHc7XZrne1aU
9aEqzSRCknQucHDBReHO5ljiYB54xrYD0+aRXFTVmTz8t4UPKuZ4XU/uN2FVTTvuNr16AZJNiHpL
g/9pA6Y08pePpcXhu475XwoBfeECANoZh1bCveYSuVysNLwiGAO3eGKRtxKGGE6TkL4zhxv3I16S
eQmhF45ZWwuDPx11lQp6ejRNPWEqIJwv/VpaAYQi9Gb0wMFBHsIwGeM/29QmzTGQhr+fYlTEv+I1
V7gBO2e+iglUla0+6CoRZRyzLSs09NsevAfAKlQzQoNg6Cw29hFvlDs4yyhlfrPtEfoFXUIjlf4D
jnLLNtqEd4wm/6eTIetH2FRdpqHeCWn7z7yk+At78mwSB+74FpngxVidPnRvrFp9/TzGTyQceNCI
WsfFEwrIuz64EofjYBXozSpmuXA89l4kXyJ3dT8mm3+8dAmksGrV+kikTehyd8pyJZw7BI4S0Ceo
AmIe3Kq/8An9PwJy/4V1q74uRZBaUYzKjnPPfcnJh6wEOYOTMqH+9DLdcIeGhElKYZC2jJrvHG8w
FJAUScrvaFWBl3a9BMz31ffmB7O/xfTJT3tZ2c4BzGSjXFEDwQUbonccc58TBeTRAlWNVFQDOYcA
k/6Fj3ltfYkeHEKDdnuA1KGhk4EihAVUQ8Nd0KvW82TCAS2WUekbrxYuwoFkj0HavilVxmWHQclE
ctM9B2Hpdza/58kxAvfk6yaJPjfKNa4v827davlg3DrpFsuj3jrtnOCwfu84lyJbU4fEN1EVB3el
KJQKVvTYIkRSCVQ+wMHpy/qL3fu/Ziy5c5GFmMwYh/02O7Qo3/VkYq6KhTsfJRxF0JO62TwA0XSz
hKVKUHj09XmR/me6Ce1eg/csdIOgNVRlCjCQgM/XlXxbB4RlFb8WaetJyUTs0U/gz2emNx2lmToH
bLd18p7Xf3N9GfXxz1QBr4qgObv9vZng8lttB+pF9hKIzgZM3h2W4FzbzND+0lyGfEr5Z9jBcEhq
75dq+Isp6xJl0EjyyWtdIBeYKPBMUmXFOrGmx3qlbDt89Ha2z4AjhNxsBh0k1W33AFR1PjVpyINh
fRbEFb75xHAyZgiN0IJ1+FuHqTa0Xy71WqKP0jxFVcXs8Opw0pJb9R1GFyNfVGAGfm/nGO3xSkfd
WcQpKg8hZ19Cji1cwsk7AXDPg0FqIJcu9FA9cgCzHkW1KmeuniVF2w3bRUibYYyl/xpDqihE8UfF
KIpkd7b3RcX9cN3eSRFxzj0kFXPKXFO+xEDXBefTCHLbpIvjPk4TtVdz7rYnlwyoPbXd9NvEkk2/
Vioy501f89WvCxSHApOHjiLENcJt0M+CGBhSXmNKEm/oubEnDa6S/vZ+zVdxFbsfHuXjrUpLGP+T
SGD+htluuOv6li/kfqCnv/JOsIJG8D4CG6KI5kd4KCJuCrC9zYhfU9ZU60TZKLVOYHv2FjOH9rds
nOQHUgOxZKnKyRt39ekyBxppzTPluSRODN39bzwJwlStKz0LAONAoJQqlGsf1WbV4ErQwVP7NxW+
kkTq/2QPS2PDRWZ8oaQXtehXFIoRYHnrDy9xxjfFJj1uj2qm+AKsQq6vVZDN43jBY26vxLc1/mmu
/qSTJrH9HNteQmVuM0wK+JLXDO0Hp8jnVfmStngtJbflShKHk4N+C9L/KH65MjtliAU2SAZSebGK
p9gCG+FIC7Y5x0gWjX5IH/5b9s2Ik3m7Ew0E2AyA2oKGOoUnBRPCzNrFdKieAimX5o/HIZmh3dFO
vbpcgKmawg38mRtz9QWy2M6uV6WnV35s31EAgKLYzrQBzlN68Gyj6gRo5e4UULZ/c2zbYRfwSK4z
J72sS7XpdJyKRw3RMt3zVwvTnJ0vrOrKzws+Dkf0wGvjn8fsgNIzmOy5Gc4Fy3ioem3pdE0hARqA
XFsd06NFZ2FBfKcCZjbKWREYSgj0IJCAclgS8BA3ytOI/tdaWbsd3tz2EAAqiTtKy7ozh7P/qrgO
ovjV+0EJK8wJc18fMlHLF1mj2tYh/n00HIQTZJRUFfvPl1Frv+e8EqorCaMuL6w0yBkd687+VMW8
Pg51abPLFivaBI865TQZrtz5tAJHV8hgrDsMBsszRaKDNbA+voWARfMTs1GyFcMBy43m15QJ1BKu
5l7LLnZwDNRrVPp6qk+bp1pck+jS55zXzJiZvqXPOy4tMhewIDSJDX6RDonJx+wjYT4uHEYnGbf3
aCJW+23fD3ALkxThAz1rHf06PIIWgTHTU/pkr16ITZt1M/5SUeBfftK4mZLpsXCHE/JQMBnaLQKF
EOZXcVbhYZJLL/ua8+3KYBXcFphaiNFPF1HCbGbLbXnaV5Sdv7r5j1qDIyy5ScE2xsdpq9jXTsOy
jM5IojL3aJKk8ijwQzUGdZCknCs/ZPTUcUndxVKDxuWpqvVhJMRDQg7DaCRmNJua5WnVzhCXbSYi
fOjnIr0n1S5wxy6r3Y3Qd0ASUkbFsdCOeYoYSZHBVZ6KKPC28+nefYlYyGc2EPTLUbxwiICYQ4R7
Wl/yTOGRCdXdANEYIEjGaBTdBsGJ7TDGNrUp4ENORdsdFuvgxdHXCOLG+dRrT2yZd9WdKbUvcI4N
WzYa57ZrHLo4a8hnKyrYER/bvBVzCcOseaPyJ7Pf5rY48x/H2BxmCJ7he/T4AA06iQ3cCnXXLWO4
WMZFr9H6S0G9imkpfQSZWSGHFwEF3luwqHt51rUPet1mXh8Vcfmcir4YAPVpZGEN4ex+JXuFDfIs
ms8m2jZ3HrgvlohVxRbNir2WRbuVYH1vrOBi9CXmpC/tWIpMPEQe34NeZfDuFAIvbeICXElDtSs+
ynVqGMK6mr7JzRCIc5uL1FOfsFlgJapg3NFWwyol5RfmNitHg1cNrj+f/Oy51B0pUc+uS97JmDu3
VAVusTf5m8lfl9Q99TsKr03yONwIxSmc7R/SxnuCe2EEpBNPDjBCheHlYsqI1f90dN7ASsIqEWnb
HTQLm1OkbGMAPKsiS7JrLyhh2zkaJ/uhXOcb6OSvtMSNRDUSptsLQGxA1yf7MY1vsJ10yDMj5Ssf
otIzvTwiW5jBXtrCc2eQtMQt7xQD0BkRHDQJqzD7nhYLZ3CY3wva6kF3avUWpNIRmtSdCzPZ3ADr
hC58qLvWVLgadI46gHCee82gukm91xB7A+7N06B73nsaV2Lyp78rtXNhPnIkQW9apk0hRexhiLhu
/y61WghE7Kg6Rlh/kYCUQxK9p/PNUsRAmorpQiwa5CQEaBlhG9YSDrPKOX2BIIy50qviGMfQV7xX
WBB3npCtQePxQ+1SdFdGtJ41Uo70yhcSgH67ZSsbtPifV+NzQ3CDKmgrTgSrjbUCq3m+3jqYLoJr
0DrJiRYYEgsF8ZcMc3I9WujzwCIgzOG52u8xgwsW25HqP9IgK64Wb2xbpCKJppuJ66AhajnGNYnK
wGf3mo4XgRCd+TkD/faxE0+ulGF09KOb2s7t8ugrAmru/8WwmTeUiEgjEFDr5s3RqFPzlKF0DXII
uBZJ1ixm/rSoL9vjAZt3JcaG+7AcJyXnRwheIMqyIaT4+MVbYl9Cf+o6SieykiyXm/OLuG5x/rdm
PuJVBDfILmj/BhabmvORAJuy2pm/016JFdHiHYFSSZX+7/ItimnIMION5aj++yw/qwAhexy4xrhN
FaS6LXnebayspQPOWsu3Lv5m9Co3f0M5xR5uLC8l+4YflGu2n6K1D3R+jeni7A012u7f/omh7Sj+
P5FCXjJ7XFI4WwsXX13uUw0YM2Pw6+fmo8m49RmyGY6bYHDzKAnQ5mmXWPtSZ4rzzOPCaZcmpfjx
s5ziDD1atFmmsCv0R9dYwfmtzLpqUMbhgoAFgS0hsrOGVzKjTf3TKmfHjSUhjWN71xPWOzhV2PX1
Io1z6uJwdDSC28OKysVB3wOWZPwS9vKCBdqYMiYy8RQ9rQBg9zEvKMa6PzWuscL5ZKZVsO/VK1fI
4GwjqLOdlTMbZA+MFcWLbCAypr8pmfGVn3kPj0nnknMuXcP9NKvEoiEL4jozeC4ujxJWb7L1OamW
UNFFInNvOluwNbGSzydPBxqVtusZCtu56kiSx3vLFvjvzqc0kPv1jp3U4i62mXI9uI35Gfq3iZUo
rCfoJG8RhZVPtRxCozY4tPsmPxxt6XmaamVqzpi5hNMdQxdOAYprdWI4YJI44zGsh1QSJXjsUMpJ
NVnC1n1Q/k8LHAWJ2dhJuuvrgQ9f/ajkkxd+hirN/veztr2zg61s1sbLsL7IKQYDBGyuId9IOQnx
Kf7LtpLBfxA1kS0I0gsQfdHn3HMUPU/wJ9nm8YrFEB3Dze1o+Tb5XECYILdDxNzgdw07GiR6jPFG
2oESs/iY6WLySzvdhaWkeEQxmKjV49Onkkj+0/qaqBAuLyAcjZE8dBcbPVcpWk1uXwhjxeNJG4tx
M4Tj3k4VQt/A0RdJXt9ZwByvu8Zrm3Lqoj138/GHb6OduEKzxrcAbSuQi//n7yHsE817ltz2J0Sx
0+Am7xXv4s3CSJcxPK6GIQ4kdvLRHzRV9gmBUffMDzpVpR90kgqYhZy6pcHoeRVHjvVQnSM+qTGE
NWWOwCPxAjerBVyc4JooAK4aG3kKk3GS7HmshHMtiempMKd6uGV3d6BYCweSglcwU0/+Y5C0Xz7B
2Rq3+6rpugGDm3g8NeNRsnGZVjlgHlK69x2noE+XJBzEmLWld4jGNkVB11UYlsUddbujwGzrLtvw
K5zQyC2aS2KzgOZQIlKhP5IJaaHwzuLO2llbkuESWeJdzEroUhULZwCKnpVxwI9ArI8CMbHU8kAO
ACizdkHyy/2AitltBZYDjBzTG5MaGpFo7LGzq46eyAJvkF+sizX1hrsqW9quGXHBrbUV0EWz6/Mb
nG4JSlgBhe6X9j+x+6Ni6wfqNDrau/VeqCTliK0iI/4ksfjVfwkZKdHKOfGVHriSxJQWhD20isM0
QbE434T21MNOTwZaRD5eAr/cKrksJ4lgCshK//HRKmyny3hxYiwSVJEW98+WNGWDn9+N8tbgiHEx
B9Gv9q7vtHoKo4M2h/8RZicFdmryTtHW7Es9pMX5+Qm4VyuLd9UqrlEqtFclfLJdwOxNKjafwEqo
/ByepN2Vs85wFv4HLn5HrD+xXKjTgWfJBwzwk5TJSvEiTXFuN7IgDG7AU26kWorYOOxJOU7MVpKt
SpeHZQ0ps91wzhXSYhp6vUK5EolBgt+8+by988BHXMb0D+2v/SwPiSvpHgyyeu+jjd9Mc79zLEzE
2PM30gQrTpiseGbpXDvnsmKgn05uOornEKdz86TjSaXPU9epTGzY6HBEDImFqElIpyIVQ53Oz1nl
C6ir0lIZmUN++K62NQrZF3KexMk1N064j+xrLWhJXTyEIwVh/sjazu6gLyBFgO6NKJLawwIaDMON
5fMsxsAYZlfgf+Yca2ClBcDrbEl/bFrx0vFAAZfJiNWkefs/DxoJXNcpcGsW2bkLdKRjmyEsepQ8
mRY0uJ5L3Yqeo1jJBZ3lMkGyW/QU46FxGwsaGNGlAQRO7QkcWSWmqFplQtkqJ9amv3r3DAYcgSX0
gYc53vTufHaZHe5rk92eSAdZ8G4kjSWCxVQUJay/epOC1rBg87CNAwcmdJnGJAWXZuRKP6hkYYDW
Nje/0sTccaX60wgw7WgTF5VfrafW6WA6fx975i2KnYKRxFzS8GB9kHaP/uFevu1q98JO7bkZ6Bx5
z0syR7TdmDUQ1KTpmxkvHhI7BcvJLen5lDdTGagIF4HDkRWYgvQ6H7ZsISPvZC+TfkH110kk1i0U
dD2fXb0X3QqUk0rg+i1B5GvzPWUt+J6RIkJjrn1pnkGYw4EH+F2GTNHK4aetlHqhl8u/WPFlIbsy
nRs5Lac8puclQUiv6R3t3qiMApr9hVHshahO/gOGhDp5J2FqvXY+GQNfJlzLLE6VKXo3sjJJH0Cr
8Lz1Wmrv8Ah1BuecmbtiT2hWCRLAAtAO58hsRPEk5s8OGgU5Saa7f9Md6q/w3NJtxAg57L0PEL6S
XJ3ygzf5hOxk++ZcijL0npoFpkb2js8m9IuSTduGrTlH/H7NkinhxSV0kzTiz3C8iDLfxn4BubZp
95ZejtBMf+hsRVA3Hbe8IInolTMTTFzrYpiMtMfgiQ+Ssav0YmvRa6LpsO8+sSuhKMSo2+18LvrJ
zzkBJz1ikgQDEAPUhsDY2KTZXAFnYs+G9/dkqEUSs/62N2stnrYeMW0Z58YQ5v8nIVRvgWzN7AuX
wiKPYJW0Ihhn1/H6v0YdU+41hYOlrx9U95AhK4vu1JnfgvF1pCSSTIiK/fPH4Z4C7ODKwkoJxdSK
PC8zZ2AeaMSzvRj/lhQpmIMNlv+leQqwLXQlFJRIw4XMrgwy64///qkJTwLzojtewRbMI1aR1W+8
VQWtAkDFia3gZAnaA8UM+hFacSD79IbFiQ+BODvrEsTUnO82WOamNjQaobjx64LjaNzKk1snhxHX
yV3Vm02ivQgswjO8thgEzL5/jPpNXVMB/W4pB4S8sRRfYpDyMc6vPAPOFNwNECk5DDChTMhwTpXc
Lqsd6O6exzexz9dk4OOCFNG0MUBbUkW6bUCmDqKHRm8WKZPmbv/zxdso84+3Vk78BfnnVXR76Jjo
mvNAELZU8645IK7EGb+AYPezIBbVdEeexxJ8FckSsPAj5k84SCGTz04RV23Tv5Q5f6kJolceQnvR
amWhIFgz8t1LGGOlC6S2EKHewG18CRC2bXHu2gl0VnhfSVkT6KyT0LYZrdIfs5NyaVw2KxUFM8w4
sEQdVQGhyApyZDz6tsLA6j5j2sHiaajy8s/zrcIG2ZzJ3udB3v38j5Hp9Q8UVMkOEMYnIDPuLqp2
Pnhn2MkIOvd+41y6d2tyOxFfA1alahAGkWXBWyXKHdt9vRhhjAz2JDvsFWnRrM10aHSPQ9oBFBku
wt1p6lDzRmBtDbDOlU76nP3Ch6B7N1S7nZOKBgjtWm4t8pPWN6hFFHgTxC6y3Ch4fFTz4z4lrCgN
lF+OzR6OV9hvt7MY44j3mfRMgLpkfKEhwI7Z7PqEGuAYn6atgpZscdgxx88vmjf7t6IoeqtLdIZu
iLsfj10vcUdEqagO3a9g7hXmqHOIDX13C494qHLj+0ESlqwHZwq91fQADwznKU+fQ0ZifbWNqwnA
cnkhReKze0Z/A+n59/ZyEqJm2CiWWq3/JVyYXznuSGhE7/WbAGOMgDJOuPDd1K2j6rTQOBcdLeib
BJz+7QjIxbV7Zg2cJ+DyP9LSFAEQTEHoooSqNgCRlazxYFA/wNnLd3jEBLqxkSDzdfR9uDZBj81S
7RfSzg2mk48s+5IT25RDPeXJT8ohhPdN/VoK0TddwnClPEv7ZMrZjj/qiFWScLfCYXT423mKU9Y4
LdkfzJ92//9+tLn2EKnyUxI4clpHLJ3Nq/WkrybOGK7Fgc7yiFQOYw0M4DOHJm5cdD6Fip/9818M
mV+POvwnAIdeWJhOgjY5MYhOXIaPDZA34nYIZ6YvXzilxZYfILIy7SnXy/jbHVI3GdvoD2PtbWLj
6FMN0m2+XBwuJlNqkDZKFHTZbO/1TC/+1TFH3iHFtu3vXoHiC/5mhpJguQjGcEGLrzNSQaRD+KPA
UiaP/FCMJJWpVuqdigR0AHxLOnc/5HYNXE5Ig15aYBKcprVwZdeRKX1YuI394IExLU6tll3sH1V5
RL1aKdR+bO56/IqDPwRSaILRg+rb8YSIw1C4MlPYsXXYfDbiyjDx0tnKCKTxM+X0FukecDNhIT2p
MQ4gcR7OJ0L6xCrp75A5AzBonYESNMz1vrpFA78yLhcJH3uhGvhbrQ0Cfi/odFdHuNGirMQ1z5Tw
PeQeR1GtaFJ8zEBrBV3iVgRiUOhVXJW8ggRwiusSWOi/5ASgtjU5Z3f9zlsC0r3OW3JXCIefgMGy
CCZRCxwn4DK2GqoOuAqoqm9Lm7jbJKJUXI9kBJWj5HlJai0eTk/ChZoerxUfzmJZHqC9yjGZk2Vs
pSdM7gN+FKp+srm1gZLaRg49B4XycnZBq6zC+b7t9ViTBp4uRyz6LbkO6c27zMX+8n4xuvRoC/Et
2GvFS09y3ujaKrlGgGtyAg9lU2whWckYPII3AsRuihk7fgF7AO1hPSFoz6mLr+59+KvauYlvQp6Y
oIyyA6aCpLpLzTwAdfMuwd+1lXbGRHiEJa3qK1spJXYM0DNKf1TvBf9GYtktadTzHioIlDADFS0e
M6LO5GnF/NQR9DTl/2OvLw0GFYvuYkB9AWHs0pYzoWwHQGNV52qG4XHe5f0bP4p/4UmmhSmzQSdK
RI47UGYv99NEA6nAz5kWMZn0RZaAgRBVa4BcQSU4/YJhiTocKbxW54NL1POO0g8+FgADrGHYaa2J
EQH9sYPTPV65PtT9S+Tl/E3r7xQRmFwC4+dALalvILAr7vtDrpitFl3nyJ0UbM1g5y/fLH1Ff9dG
NfaksblE7Q8oDCgTpFECT0HUUM9y+IuMleuo18NUj53Uscib+dgi2m6TEA2gzCyqyTGtFm44ce9A
tHvcXU8knjf6P1U4awDX8KALzIK7ezmxBv0fOLCwF8CLAwjzg2eVWvj1QDGdIChpWbcgezdL4X/k
toGEhHpEa7nrAUVDQjW3Qnf1SQ37frVhar0Z8vMp4sbL2Oemrea57BjfqRx/V9kGrTHrzbAEd3xi
wZEZlFZvmOt2f751ni693Gb0jOP9VBqrZiKUcm8OLtPBCvbOPRmlD6MxpKsfzYULPFy/SvvHhpXH
Pa9rt5SirJU2xSnmLdEZv0z+5frM9nI4ALQZTBYCAOuOHHXhw0HV8xoD+kZ/aI0xooA8h+cngygu
9EUttjJAGsD++x/Tsj/D4PcGNgcXLhYlUxpp3C1wB1N4lHq2Mxrb1YbfIYVSYWY5A/N+DA/StJgb
KiJymvcssxanQZIlJCNlextu9IVoRDjn2rasmwMffPO8esgL0Jd7HTHpp2fW8zk2ztOiGDa40znF
6ywpVZ/pq/ACZxBGHgUNYXlCSZFQSabtZNDkdWNODibTYG6o8c67n7XyKQSZT3/63DZUeMonaty7
eEitSEomVXbgXeciFrfW+l6c8yp564B8v6ruSHlJu/kDo4y3XPi11FI7v6VkIdGXR4rRvaZ4B6d/
pXLfrlEOh/aXy+zUGPI4rCv6R+DKS92MR3KdWVQkeaKR+9ifCBCbOQndBbRJhq4p4QSC1ChW+6tl
by/A1NSH+eVZy2c5Jq7B4TM4O0TnLChz7/mb7WDrt4M80agOqKBxNYmPcHdnuSHLgBGaoyIdVlcN
30rPSw3pHZXmjpRccCxISBOZxNWYgOhPm8NDHHw7gvjpXkJzRgAbSePvAlVtpxAJrHLPChCR/VCx
F7c52qOGgNGVFTrJhijVKVnkwGq1TgOtvgUb6jDnaHFr2QxFRxEBQZFWV2zLsetlDt8D1vypCohb
w7kgqhd04C5x1slK1PT9Kn5cm2SlUnAh38LDSnp8SSDXGR/WvK0wHeMdU+n4xBJM4iwYgdTJ4y7V
49+KuFkNPT/uJvbBq/UNe6tY+BvOhBAonMSgShJm+uNXrG4Pt4LPdLfFwajuad13jbi7w+p42tFn
MWf7SZFGG0IMrIfg8Y+qJHqw+Whw9vwViPVysgy0TNQmmARocwVA3cpq8gG87ni7j4xWLEP0rN8k
t+Kb4Jj7/355LX/x09AmFhWgl2GroXuZWp2gT1MyTgQVjHq89WXpSq73DTWpsdRMEQFFgXiqWXt/
MAL26EXr+vFk0V8TMDc2U+5z4h32ZG0bGR95NID0fv1SzENEqhnNpypY1UeF4yre1YsHZz5/4cN3
Ilf52lEHZ6hXlOS2nSMWhhgb+3hUQF9uQfOUUfH5StKpOLQQexANsJEvqL1L9roZyM5rX5nfywKU
0OjnYdImwoJQOIr9tn57+aIhGbvEfLbUIwWBoyUVK1x7o+GX/+7/9SE+Cw4pLIRUBN/2rtuPYZ32
SXbrqa7DgvZR5wJgTByIrUK/mhbpMr1rE9aX2x9nfNXXwINKtxfxuCeeOFgLuckHEN4HqHdafzxF
cL14dH1AjatJ9ChbXoV538q8ti4f/+4GYeiK3io4JsybbOhl5sJKPsNi0RktN36wbl5j3aDtIScX
vFWcINmZyDZxQ1oClkvdKvlbMExhtYQDp3QAnJjgy7MDCnby8OiF4OWmcIan1g3V7dMnJhUfkneI
M96BAvhLnql6GMMRXJE5KvGwwzWX4LqwQldbs4PuhGDUUEG0J+MB8OzzXLMuNWhPIeqpd88ri41D
ate/4FIXYhMf74eJ8OWdMxYwMUJdnzf1ppjtKj8ULCqfNjh5Fu98Org1Jv8h4yyJ0LgUj176LEmW
9dXPUvVoXQTVIfckc2H4cHdci8AUWGIjfpjN1/n7HHSpwbSFWi2vkDQl8I4YjLsMQr+cz2DzltX6
g4A2oa1qupWSK6rRHgdQUG5aZPaouHF3gr6XtJxS+hgRRHToeY83s98SkuL2N2R5YtPOBKsKo6wN
/vUhtCrWxyuoQ6Ss02ASyBJGOKa3gjh6AxaEpPbVGoHaPI8snywoE1YYhb8e/q1dLLTNydABD//i
OtC2J5Q8ytlVPeMVjGvV7SjJrobuNBiGBlg5cupnGGUV73f8o5OcHQVf5N0rZmpQsd8o3dkLq5Yj
7AD7CmShgnOXdA1DgmTLCQC3CPf01dqwUG9mJd1jChnRBMznoKOuUyYnKVY9aBhoV9xljIIs8cW1
i9qPcIVO7OBv1opJMRSbbULkoAa5nm8klfd7pkKembjC6Z5i9zQ/owv7sWkxrcnqq16t+SKVw57S
cuLjzWRDSjqJIcJ1udKQMzpjNkWdyerK6WmxvtjPL4+Q1qmQqlrvkjg3FY4C7OS2tje8QeyPmfWO
L/snZHTIAynQ29fQWL9F+0EuAjdTxR1g1vU6CCasR0OmpRuQVGYJhYbk2ygNm1LNg3w+YtjDsm7T
AgDlOjJ02WGbLFFs512alG8aY6hgMC0FLxPnVPkZuJYrmND+WZFZUQGlqJ5uGE3JDvWIWazYe0Q2
c7R2JXDVWkYy82PTuvQE2XkeagdUtnxkEELusf4orX+s/lZeuyZ6R0X6NHBajV65YUHj987MT48W
Jn/0EhgleUFoj8WqjQKtffaXCq9X1DdsBJy4CcTW+967ZQhLmVq5BEyutFW2Cp5Y391UCK/1/xfg
Jm6D1dPR9y0NA2AUXDdO1OEfma3rBlf+Np+to0/9df8wNTHAKR8vJinLzPjsQE7nyx2Ui02cjctz
vZ2Oms0Q1mUjhufSaCBubiTKXFU3+n5oLipJrhquMFVkirsi36/ucx0w115TyLqQtv/d8TKNqrIa
KNpTx4pveIaYtXmt/IUJIubm9reqcg6/op63t0UrFxgVtB+DvaPrhMg5je0nakRKuKc3IES/agAL
SqPjWJ7tf2c5QJfQtlyto7eERu6NCsoCR+tfraFI0YD1N4lo6/UZxsV8bsG0jqd3tSQuhhxuyxd3
RfQdfSQum4AlaC8wjiPNJ+mDCEs5uYyUBBgDSHxacuEge1CdGHcYQnxqaLr4dDwYm6znE7kpn8Ob
Vk9ifBKWMiC+tUs+qsIao5D5dGxovMMpqxetnS9e5vuYIqkNJzHAJ7w4Zgu0K51R49VkykA3zP+m
Q340AY+W9c6VE+4EAOCEhzJ5nJ0Ut46aJX1ZVX+a1NZYhZs8/eVaAcLNf55Xo6R1g5xMErJzgbOW
uPvlrSLt1DNTrKv+/mb6AzeHVMq6Rsu5hH+B0gkjRkm1zDJ9jd/c4hpsMCoBbwHoC4BTjVKd9zro
rrR/mir676eXB027j4VPm32oXV+ABl8BhT83OxKMLdA0DbNAa9IpdGLJ3X7u5s28wy3lshu4qeg+
ZAqTzPFKEMSAIivRTbToTqV569u3/sLjnF/XZM8SIpcoo/rnqWPVCxYPhWaUS3xZqV6hYImk7Q1h
G8eKap42Ue55+GFhq5N6mKLs/1CzdRu70fQ+D3qpZtEqpSmaTBWIxjg1KB2A1ERfZjBw0jlNAi+p
deIMAKf+EuAgHewSd5MGK49o9T+Iq/Pg4k6kmt57cm4lWuIIuUTkvnEcX3M1m2OnM5ZaFxSiuqZc
Lw5LzaHl5NpShXuAEUAKsL5keBlrDwPi4+ZNX8z/9wxOhFf4DbWH5uU7Pu9WD9PZ2hvWugYIG/mp
NWt21SldFBrlN/WMvRyEJy1e4c6Lf73u8cmD92lVhSom9dV3c3hCaAPgQIMFtTodD+hstsWRCxTb
/kAfV2GrCejce+ajrkKlDZJnMJV+7i6LZ7rvYts3UgW/d0efn+lj5Fg6rWhxqwQ/11Nwx0ZtiQVV
ztkHEZZnx6zMaiRebwz7WAv3jNJXWRSUjeQh1X9VsAzwSphDRFSVytLRFVFWYAdE4OwITZS5mIra
gX58LdgYGWCNynApzTbw9jTYVSXhuoYE2EZ1iE7ewB72xEpNDj1qCH/I4W9TC22L26QgxAvPZWIu
0na/pCrfkeeZ3h53Qj8uJaLLKw+Vqx9TLAh4XnIirJlC7j5NVxUiCWB8A5+09yb2Ed2kPUQdt9WL
TluWvddvia66zvBtCXTb+JVe7CKzUeLMuPIUpssWGdJvo5qBb/gwivjTowLfsBh22jYdMZlPypAB
+pTbXkSWOk5jCmAvX2YzV+zejAj+bEDl89o1OesG9Vc/PoaFmWuLGujW+L8+4S3KC8Tbs9CJYcHW
ILtElfN1/kaTOVvgHeo7tIYEfUDu80ubhss2Wtcmn309uSev53MY45VYj10GRJuG6g2sxUMCBJuu
wuXMBB1kqG2Q4vE3S2txnRfk9ltCp/iDVZv5XVUeZhQ/MPMowopMmdXlxg9ukNIinkarSiFzqa9t
+IMUA0eVux+4ZCA/0N4HyKc3i7A9nfmEpGoP6LNA/K+q+P+e5uAGyKjhp1iCzOcw0+79SZLcw0Jb
3SG30nERXIA2vzmcoYX6Q5WNG7+MIPhpvzXNGaBq+plGyEZfrsucmTz6xOq35/+jLgfo15kRuYBd
sOO1u93dE1AHexwYfczYXoLAVFwYXHCWDRi7pUSP5FjahrM7V/0hDpffazbzilLSvSCGMdwbtSLV
ORxY0RG2KjESzCTXXKLSPXJNSDWJ86l5fg4g04YZi/IoFaCeds63JxRL0O6LXGaqR6goOKjw9GkT
D6wAyXCp8/EerOCrioffYiQptuZM+PttrQxw9z3PhfarNm5OxPN+xflJedT/sQHO8vSADIOom+LW
NAIxq9M+OXzYbnj4Qnw+rPLb1ShmL01mz23KY+NvnFNTb/E5LWIYuGHa/O0AWechK2ZmoPPINBNP
S5jCnb49Vp2KUYCOQUAVK/r+r/4i+l42BSbO1l56l39b2uCpn6csINApvC5NTe7gwwVZKnLN2bpQ
HmiWXyyA/oemCaEOTVuK35fpG2oo75ai4hJAyCPIghl3NlrG9Mv+Zaf7Ej1ElTjaHCxA+fudr0/r
YvcKpnyWdFh9pwXzkjV1bfQ3PihT8L4yhye0pIzfvVWseAKt7exi9PJjc+GRFr+ZPHPJh5l8ypMM
XpMRnhpGfx+wDMilIW08bpUotyyYHyHxNLr/C9o9VUIadbkL/E+pJugZdcGuFBT7gH2grz2OZBKr
TPiueIWBatWI6ZHZQFPW1UDeUR1LUNKPtezt3Ycy6xuWyn3rbC1mxaQb9wSK6/MTZVdkzialFZXE
feabJfju+GwD8xybaMqjzBRqWpm+1inmRmcXZxTk7Ky5f1+iL5WNHUcGSC4IIX4v7vXlaSs/mZwj
CkSaNjslpnqCs0XUuk/ueHk3dyFppcYuiLHNYpHnQc2/b3KFBhz9w8FpAKdvwGgOGIAolTtIDDou
teKqQtkXHW5rmnd7hdC4J+xzPmunBbregdpHb59QWeFLwBwiesfoutsJZD9WzWb1YwqhLootzPVQ
nJV6ZEws2qfDfl+h91VWK130c29wcaBEwrAEw7nacUcVStDJj9OKkvxkW3SYMiIM5aCQ5rVRhtYI
lcb9aG5RzcHUS8gigARmK0RAGo9A3gFKQNbNFC1NV0jsViP0CY5e2fccocc+EsK//gTQBhOfR6uF
HoEGwhQONYUhzLLlcz11JDg5g4vHYd1VhHb9jBtpbp27Fil24hd86o1NBIsCRLZV1tFmHVCpPeLm
wyG0xaeqv57cpTgNoRLGkyJ6fegj5Q94DLC5UhjPTgWUNlVjz41uskDlV4wX2vLUfWZj+tYlsDug
nydzatYqzfIn2mDN76mS9a3gFHiZNmR7y7ig1T1DfdVE1pgGUL1p67v2kQ43cB1Karkhq7pKxyB1
OKQhPzr+Ze3jx5NW0I4noheSvVOdRaQDe+5UDAhEefQ7lO38TJjiQmOv5tdWbdHjvly7xO5D1rC+
Q6RJA3Jrye4o2DKnBwS+T0RJw4CBuejpqACg+zCVo0KoQ5QlOSaRSK5Gpei2aKWj3chhlj/Mq6ZK
ZxFoB/L9ax2apu6XVEe4y632b4CqR6v4C3CgMqbU8DBMPc3/DJcFtCkP4McMZhMa06Q+cejsURs2
Nr/e2QFkBgCh9mZyMR6mSX5WZVEJFR9+1vF5/hoWBhcuo37d/aMyCVjEnP8ViWXoWBxcJysTNmgg
ZHf7E28qmJz84BFDIM/bfzOr5a0j6Acu/GPxeFk5BmugIoyCIYNW6n0YnSffE+wae5CudGIYlnQV
XakNXrWImbAlSmRJSKssivnU2z8nMPzBmVW1JKShqScznp1+AHBikjKprdGMSwq5mBZq/upoXphV
7+kF5dpT+1BWEmW3SEx5r1fwX6tbJ5ZIPetfapJ6EdxTmawxdQYUmrzr0cgZNAYf/XXcKz7kLfgu
y8l81h5xjCWX085lHIeT/psCaN5at3aHgyRGocWmVtW6RNF6sLkqGr3x541Bfj9teTgw+pgEbdNa
fKtHDpwV5rD2wRnvNIJ4jTQ2J6PahR5kCwImK/jQOacXIHAYFXt4AZHCuLTnPhV4f/fW37iHEgZW
TzBli0mqBB7CCeofmRHMwvnRhW1/QJ39WuIlfLHpmeBeq/Q/QXFOENyKx+iFyCqoBnPMd1adV/w9
mDONWzkg/Ph39cHaanyG7rRtKE7dpKfqg4JW6JSgChQ6QBXdjFPd6OMrk4amyxf5dL9udKGx+drb
KoK+1LiYg3ZxI3IUWWhOyzcJrSp54hiDFu1xcJkAqA8TwrPLrVkY+flFpFZQdzLiSBvqyJM0uS2n
7v2MbmWHuRaLsdLk9oKmEpOj/gEEEiT8aDOJlJsXa5ecev+bIc0bZVmcS9D+vaQSTpbtvHK66AG/
84la9q+O5hLTLXa/ogpRw1U9ZZT2VKvUhC6iBKxFU0AhEAFI/QTiPh/dn5hMTVXM4KvDyV8K9AcU
5MT2B5/UPtuWqDi/mdp4RpuKqldpAbuu5uRBAMRwVN6Kc6LHRFa6ceGl/laXz7F3WFMvEiHFl+P4
PwL023HUzrxh3KHjG/UbLb8YyULIjWYSLfCqLSFnRm1HmqBNruHszkND3SdEY/9Rer3xTXSwKJDc
Wu1mLN6D8fe0Zp5dh4REj8IQx1h2CWgL2JAjd3418eW3jIowHbN3rT/ph3ng/XuEM/oz5iz3Agi5
cBrB2Ia4BXmqrxKMEo6pISGnH9pkfJQXRSM4J/uBINUwbvn1Y2z2Qah1aK6W6Uy0u9zegatvdnie
JfwQgZCWSzrs1f/r1ZY3BIiWphThmCbfy7qpTuJax9ut8ieZq0KTBrjtAtUMkqPjqVQya/Z9VqIl
geBiEWxrlq2Tb/T3rIyG73I0LM0Xyt26AmU2J9amt1ds7kPEISoKo99hamYiRD8Qwpatyq0/kNFU
R29RNA1BOtTS2PlO1ODonm/HTXcHR4ReK69W60kHK/g4FOpdAGoXXt+/+5qrcMDCoI7XGpIu9Ked
R2n1ZrCfUE2y1L1+TJNsvTJBKRcgtzFOmGwZLcvLzwPOAcaUVxVyuoPO/QCnJtpJTccimxAk5r+A
0jkL6spNc/NW9TH2IAJS14RbE3bpwTMBvBF2oUVsJjnfEqv8gcj0QhSZxFoIWoR7ZmpwhUAwhoSW
OfhfNqhP/60XhBe3Rf2pE7SpB1HQ3nxIB/Kyk6ENk0tdQWF5YtCzIhf2kY7Xqi5fDlrCJkgrFpgJ
SCM7mbiFpwWDX6XSIQEtmXujmxgCxuUjBnCC7/Y4N4ZABv8FVeLqiTElZdiu/xkn44qF3V/urHM7
Ft/UndISaZqzWPQGV8Og3yqr2BHiutEAZ6EuK+yb9Ptf22Y35CHGOWY7KwnB04xjv90vlXT5Shv0
TGKO0FitzxoQD+LOurvGRp6iesBSu4VV7T2FURzVW+hFGQOOjkn6L0cVny73qTLdaRa0p8cQwXs9
OLVfkE36Fc1FIlgxJInDBWQiNcza4n7UsggYxKVRjX+jilZcXE2mcLUIphxEObzMMcPCT5g2I51d
fdVkgm7l79IoHciGDTCD2bmbzd2OXvkMgAb3iRGkUu6XE004oWLq3GTV4JLTdfT+sU3IZgQSAB71
RX8+jF6TUGqW8Fxh+vYTbW2+McgoR53w7zk7FDDdFmlSHT9+OwFaBgoXK04g+Optvzhka5dCj6tY
s31iG1IqlRv4kBdtj9bUitUTQmyeJLMFHk7tjtQUzntvd8My5gdb8G76CdmWosXEASx68KkW4B2G
BWukAd92ilHR9hbzWFstF8hzgNueBbtZNWg9kn8XV3KCwsfqNtu6OHY4oIb3AXECN/+GxHoXgVd7
l/YbCXj2d3eQXT1jQrse6swC+IMH+DX4yfr8xz5VwOyI3yj4D2PSiTPmDuEIjoGi6D2jD/zp7cUu
VgcsUIYiOybBNclkiceDCWHOIGqXojJ/NqcM+j89f+KTSfW8PKvPAZ1NG7+qu5kYS0Zlo1ZYISJb
scz/Ynn2bEwyt7OU66LI+arwaQ63msm+Yr8MSv2nmu37IQaILbXpscPCFlKvRSaX8RhIcrIUi1QS
hv+MB4SDC+LQ6mDFxB5MeoCxqbhFp4+0ZV6fjbgY6ZeYbio1vUq2q5t48lgdv2tE0jhHq7IZ69q8
3jK5lWqc2cAtdG4DLsZsQ3OJQGm1ycyo3bfFNeWRNLAnZncQRZfS2/2Ck1GmIb5U4IuyYhse6eCz
6TDoPUhl1JjTGSyD4YyQmWpRhzMfjdgcqNENZCVmzNARcX21gqvjNZ/+KJSyGpW/q3LPOWpC3ZAu
kwQwe70y1nIwU9N6LXADHcLVsadTOnWqLYIWVYhGbe6o4TmD98j4CDXBvpt/S3vVvz/Whpls44+u
GTKwO+EcITM+v1VEiL7XxmKygAPT48b4mKM/mNodmhbzASMxHNburoGv9cJS+FFD6S4Cmsc49Q3W
0chONaKV/yxnllxycxAs7ZtxVDIKJVAcIE6rN46gCG3bn4Brt/vS9oaZY2nFKe8rznaS67Yoach/
k/4AsZH9dyOYioMqcz7MbChIZBYN2flFBkafMD8flYNEqNbFrTDm7c9NEyZSpLmcB5ashrFkNmUH
8YFmRN7O+Uv2UdoN1kkNUPxQyHNoosYI2e5D76KeL3nxuAh4WPNM8bCEAsygFjOoRgU+Njz7H85u
F3BTvqBykm0zGUQ24XX0JnvH/3u7B0SFBpn8a5Ujyb5+NM136vFd6u2CRIooYAYo5O8QYZIh7Cc+
AstgS2DORpahVWPjLtT/3ST2OnNYBpg5vvSAtz7UN2VzFQ1JvaAQcZcQmTt0gqXv5zu3lx7yHvS8
ybZ+5LEavShleMDgJya99fJcnCst74qlb1ZDQ+hwPSOGiOUvtUW/3U09r6ZBqLo2lHzmsZ2quHqy
neNe/kRzy3AQ2sk+Hyau/qYWrlzWfq7TlsVFUzlQrHdsux0grXX/+V3nEfDtjmacLZaDqV78IKoi
JV1EQw3KXb5TOm1lEH+UY41K2gzsjU1MK4D0gz36EFX/NrqOAt78SNGn0NL7QWzPWoClY9MpGwEX
n3NflxjxfeQJu/2bPRlV9iuBpVDndbcUBGez/1bQ4G1dfRUwQR+ORdlJWKcqX0+dEE4DbkDMQwAx
KlO4MaVn8dO58E3NtfVlOv7a0jAyLNgP9DcBUr04LWq+P6zqkTJ8vnx/h5AtXcKRHj59cDcKOMvw
zC67VqCB5zEfse9Gozo7IlNStR9Aa81y9t75z+A2RJrbb3mN0cXbj5clSAWk+HaiIJ32XsOAac95
a3GGGYKUkQ7hlnJCPJ41kj030q+yqxJR4qvwC/9wJ86y1aNWA+AWIvYcQZVi9nCX8b/RFhPQrQtC
W0GbRI8b5ahid7+HIuiGjmYNqgE+rVgkTUmIzpHF4efh6NcA8/jG5kcqIhzKi2FPyb4xjNtUyncr
M2vwvGZcrtz0OhsDIBvT31oQ5POWrldM+weAqtA53p7Dbyh7Pp9OWxhymoqeDjTm26rIGaN262Ds
LVaiwhmAzzkrHo1Zi60Fie43WiFkIPTn5v0r5X7h7F62tPeU8eCu7Kij0wK+7Wjm2v+gB1J1iWxj
8CbQJDKax5flyaW0BCCCROEKBMCLsnthcCAImU1t+0AYwXzjOW/qi8gYCpoCempVEBYlFZJll/V+
gUNogxXdu/sg8ZEjVXs7Mhj5vVDtjpHSpOMrTrjAPo2KdMld8JiSSD4i/rD6n5/FN8ux1mAQjnk7
0enbJWtixjJ6FZSWC2hbnTozDPJmuzzmXvwltq9R4r8OZ1/ZqDifyVjiqzmJyBQ3FFG0vPoViUNq
YwN/u0X5z1ZfBP12/fA2DfvUrtiTjfCFGcln8xV4GGMb2VRIcyh1IX0QT6q58ug7x126esSfKNOF
j5xtzBKc7AVJkm8vJ1VUxD26uD0M30vJCpSOWWRbjuCcKtvc+5KEp+3MEDI7rQXrfJ+kCwT9yJAo
CsNsYq/QKp/BkN/0/dZs+Nu3KJ8KwNe5yq8xj1K1UUV8BqcXHg37wCgIQNDGeEppXdxau4sryPck
Ye56p8CCoF52OAVnK1Ol7npoGK4YqffU4H6nhMRYxsu4uipaSZOry65kgzokZv8jLYbXwnsbgPSj
FeA1TriY2CUCGluWcoAZw6zNIIijM0TAvs58C1cdEDBBQrHPT5+liLEZKSBsK9f2edPd2V0Dcoxf
LHXmkD1VM5NP3D/iqyR/YqASpL805cfzHhrvG7WHWch6pGnL5bh0nC4LLVFbPK+Qs2g14mR1WqC/
XwWUVrrZrFMTn9ApsL/G+dj9xrZcfUNqJzWznkAJ/OBGhdjiAh47sJzC2VzMvx3Sf/6KkU+w2Bru
OigMrPpWGI0BcN8E3nS/0Nj17x4uppc7fZSMTnM9SmuQayn51OzLFyekn5rcoawqgU2K3nNHlZeG
diVUqCpUgA9hZKvKRWOA2mWtT9dosPogujDqlR9BPZtnxUTPmNeP7HCls/lSo4//slo3lD9onPoL
Tn9SEy8zv3XZ3jgMOI/EtHQNnkvnzgBiXuazDgOUEhKEnhg0Vib5YkWNJ4rm3+RGccOQdRUODZ5M
Q9Gu2FoIfIocwX/BAvQt8a82axOesvB+dY3yqqrBAQIPJI9+dFuRJj2rfrkcgV89rdwaF44KnBUr
FIUseAZvowho7FyYYi6R46UU0YB3VSX7jg5pG92ex+3+qHq1K6sitKC0PJTZ/K3vmqe2v0RTKOuZ
9Ubtdx0J03eSJb759kqNevp72rujXvr+8FhQVlj+Wgj6iC7rfAVXO9F+burFVs5evndMDDF/HhrT
RNWozi4/pCfrhPX5imb7f0GRopxN+ZnoRvexIc1GNuhU4jLaEmkZ29AD5UyUO/ETD9Dftl3O103I
pBvMGjEBKcNxnaYVOtR5Qxnj7IXWWh/u5bSXgTQId9Sa7mcE0jBPT2apg7ZQyZZ44n4CBJQZqTOw
ly+VN4a5Mda8rtVLzHlqr7onz/R8q/+Xbr675lf5NSXpXil5P48fBUK2jnDVK/m/tEEP0wA6cUXy
9C3bfxvAyNXDlGH+t1+A/oFPo5eXWGm+RxezVhaoKG4l8kYswBSgVzSIEe4SdVdLzqCXkRPIvtLr
y/MRoaKGKgeIvDkhva+08GYVOHORjNaWBL7GX7S1ww282/Te2WqR4WFWjmALNE64E/dMKpm/tiAt
yHDD+6lJVfhky20pZ5Py+LhcGx8vFyAkMDTvuUaU3t9RJ4aMQVW3KzAGD6aZy7O351up2NpDpm07
VuC2nsZxExPwoS0h/QWFD8hZXZ9mJ95OOcbKkiv8D8ezHgzuCndlucNxlB9CSYORTqzFJ6dGPp0f
ZriB56muJPNnIP+s+PeUogfI1lNzFP9lrdy6FJCa1CeGufie6g6I4iC2mpN+qTuHIu32sFD/y2qs
HewoDbojOKZltyyip24DisBP3yoSrAmhnPxpaDgtxosP310DugByErR3VaKurg7tn1oEpT7M5kX5
wEExWARxuVRIBEecxuzEse6KuFZZKs6shooGrc8tKLsrjgFJnlGnEghTm75uoKfZhi5NmDibGQmy
R9OfblwPfnAzxlgnDNS2uP500ALz1SR2xnHbGNw2r7tiZ4AaBd126ULHpKbL1VVeZvv3fFRkL3f4
G8luZwVwfY7v+GpQjciIciDgRRnWUUd2WiTRIdpRpS3a0SUz4eSGFxV/xM7b/u71FVafAcqQeeNK
oUgQkToLKdtWr9HYwtIqINHMnHSKWEMmyc27EZ0ml5EmymAYyOqiN0M97Z3oRH5I9Ql1ZFTiFmKQ
XH4A29rfTMr1fVSJgSqtncqqxbCMNVdrH588mXp2qiz2mQ2MsPLxFbXFUAdbpc32U/VBhNwkPnMa
1iHR+lsLPLX+ZQFj4TLl3sMpMR1aDmJddDRD1j4lkNdWyerg9DfNPY4Yz0F1md0WW+jLHtOaNTFk
rslQA/GcDmWhOudg+y9Iy7e7YLMFAnldeq3wK6dM6vrway/rdIg1NAXWlK1Wsawot2l58LLmveO7
ti0V1RXhRk4fBfpE4yninf6CDb7RmTooWEf+pYmVNc/r1WLvzR1FP5aFfaBmXoOsX9KgspPh6rCN
e6nc4J5DEuFppspIe3GQU1aNTz0o0LZsX2ioTF7G1VBVGylJUlU+c2nxZ2+qz+K3leZpU5PcUuSq
KrX1npFiWRGATkOpJx+9fJxWMpJoL4Kxos/yx3yorpKRnJ1Sa2MYSuOUQYvEv32rWGTxvxJ1jE9H
1qs4XKCuSuzQEuRVNEz66BTfJ1nw+Xeqgx/bm5JRANVAwhZvXu7Au882khXPybOqiEWVficz8oRL
+4IAh2KGA4nb8P/FejGzUoHFEXkOkTf2u/i4CEXPsMAkVc5iVIS0wrAwb/1XnJHdX89KNki8kmYl
jd62RQqq4Ue2LBXLMMX2gEgWtho4mShX1rbaIhj0VpNTKrYbkSSjDq0YBYUs5BZHhMdg18Tadf13
lzMVv4GS9sC+rhuc7zklFhDdjDZxH15JdY3RYLm4+z4XI48IM9SPPFzycrVFFcJgp9cSE4Qc/Bua
KLaeXA8zd5t3QLbwLdm7QtvMbiPwwI7CLAUzPrFVJBzO7044H7xwXZpL7iqNNyPyKXlYOaOwj+oq
TfoIsOyZrsE2rHUT+lHzNon0LmIDwL/ySKQOMBwWHlHNeXz0a1Wj5v4mxuefUYyOr2sM5GMre/rp
p0Ulvo+S/V9UgYUCv8dfdgM5foCxQvHclUej+Y6T4jNRV4zR1zqhLEOu0kHU6MJ5qzYZoA+frLHR
WJAQoLV356D2iqTebPBNrLcI2Huq8KrugGnh8DdB0i8xWBhHxKarhJgYe07Xgp5v/N3F4pVdaDMa
mfAT+qEeIFyUWe6qZuVuOhjM8Y4N5rZ+veQ5lwhmg3HNgqBAcxvKKZumHvm8YQYBJJDT/gGCVAy/
n2KSpXkWHgV93Sy3j23PpWH8oJiGGsMtH54Fq1FPZTEAh1nTZnuktljdzdorqmN/EKRxpWNroSnk
2MwI2SVvJ9YUGs+suwY95+ywrT1QU7w88ReLt564bJ7pksuxde0aOUJwp59oyNVx8K2SB7CXHwuU
a73Gt5yxCqusSmAc1COWIWUUMjErOl7GKno0MkPYF/CaR/NNu3LKI0HStYEK1Zi1em18KgBiCfYD
/50NjTFCC/ILlOqYIacc1xX4nDS/EZ+kw1uiQoNGtr0sbTb4yQCszhKcWHdHdKzKOUeT18rkkpFf
iH/gcsf8P60KGc44lmZiSPE6FoE6eTij0kahusv6acD2OPOxiZTq8zW5qU/lQMPxtTaNrsA3A0nS
V+20rXxIQsNroWj2wC8E6pEx+VNeC1qN/LljXF7fzo0YbAf2l0fhHQvve3TzSF8Sf/Lrh5uRudVB
4RJMXUTyHBFq+86lbW3ha76BtlY+PhLMarbPeNBcEzQziib3NSFQ1tUFPcBZJYfx//Iu8H1kszdZ
33OGqsDQDfyrfWbBZXoMMONlu8d6vDsUWy0v4mPbPeZg0dS4y49BKc5VH3r7rqMsod9rt/jGSomi
tvEfrLa9EQQN0zNplx1d9KNKTEeCLhgRAU4HpyV29AJ1qK0HfseRFGKYh2NiXNiuaYUJuHGaOsEb
QucyYeNrNK+e68uIViKApviNcFWchH+5OlcvNL/NRp0/BBBqoWD/xlbizM2Sou259NIG+szd76AL
lZZvl6rift8JmfhjsWy8+RBstnnrMJoEuKm6Attg0oLE84yUqvAoY98TQM+qy1Xnj1IYMgNC/A84
R4KnPEoXuMsTR/LVHUDNubpDun9GGo6HP3LFdG2ravpBibgKtYKNpPTGqpm3ePNFKsUQ0FrtPPP9
mhQM9565q1dvMmKwavJVzEU4SfAMmxgFMPiK0WRX2msalsjaDUHma1dAIOw81wi2rAX5ToPzq3mS
kYCg/qKizR56wiBqT+LAOfEkRAz+mDpvzfpmjdpMaRuuhMtCFSt69qV8FlI1LsaZcnK35JpL4awP
pzM4P1tdw7d1hk/cRdrdNULxkoCxM0A4CEf69EbI24FniBWiqADKRsS3heCGrOUZL5l14vHSyMqO
57PsDmQaixcUJ2I8xVKYPbfPBdeDjAp4IeFYDHqXVPkBDDHVMHuJbbX0bCm3A/HQsJqN3r0aK/I5
4scT77+Jy3yj6PnAt59WnBoiW2N1N/r3kmlLubMid/7NfDiUzdjg54ty8XKA7kVObZXmOQMuJxvT
SGxME8IqNpGkPne2mVWDuudV9HwAbuTEL9CvezTh7I3mJ5H3lJbI/3MeQaW+4NQowyXNTT5XT+VF
Q05k9sduxdY3E+X34fXszstr/1ki5DoWvGvVpXhG5pLuDekJKzAghfr9UGgqMJ3+om0Vns/cwINJ
jQWAqQhr/S2AOg0ha0Ns5JIdc9i9wY4bBitLY78Z/3+2vpUwxmbam2o6ppeqYwuH1LkEJQkvfVv6
B45PYyAAq9ulsLTnghc7hXRlGltnpMS6Lq+QtF7ioqQoSjb6fPXHfiAJB60rQY09q0Nh7rBuV8si
WG6QMNnwFNodo9bYiFNrpYbGtg6o++lQAFtsx2Djt8xuYTkW8KGzC+AA/9zuu7By1vOX7839fcvw
IDqR0SkT4GO5gwZ57BxCUNRjPYEpirT8Sk5uetMl/RdRO5vsMT7QZ96s2cP1UN5Os5g6+DOcZLAp
ScbZylCiB7HOD3utJ7iGPpwu3p7Km1wpQD3Bji8LVKUIdreckH9UVvf+B9ixon59RBDvwr4U7G9i
yxhZ79T/tvU2l+1LgFy2kAUbdXhN7R/2ER29qRItn5Tdoe23OBoMRspYPsRHkmx2VXtH+NnN4k00
hYPOQ/8QfbkYuykiyYsdzcKM0ABYMqAJtLM8BQ9HRE3IBj0A0exsgKy0/w+flo46+YiaUckK5WEs
FcOe9UNDyWpGPdRCeQl9IxwpNzM2hjnuaOzaO+GZ8rpBrxJYJWivzv12/P49dGInog3jAD8X2jpK
q/gdGa0Gfxu52kIScZqP29QWyezuVHEQXrsJR+YCYqqmqw9dSCYku5FZifIEKVwEaDuVo/f8pGOw
TVTAKNQMDTGyR/QwAxTAUrJOnPJ4sIA7PCSqwzwVl+uyTI61ufGICezgzLnNMCfgKsfXHO2XUc5i
7lTSUDvHg23J2Ou7Anivy35KgbO3YbTneQ9Y3jUi5M2rbBt4mDWBlqoMgJpsZSN8UrwgeIMOTVqg
jEtGOfOYsJsCCKrk+lkN0sHqFT6BNDp787POL88+phAlnuxVAYRvyewMnKt4bBg/3EEPL8R1jql6
jT94OSfHbL624bQaT0bgWdGfQ5lYfDkgNkiBWcHX1aAP8z28ATrL127jJ/V4sqhqxqTke0zN+Ijc
N8cUR/9hvRF8oVvvWJ9bf7Dr1m6qnfCt0XuVg6gCTi/pjOpiW5FZLapGcfS0YMCh7F1e73xPBldo
gkUAp/QeGmtgm9vtvpqZEjwPof/Nk31mMjDZ81yy87FvfzjtioJZQfFV0tyTaXoCu0UtA7TiFzqL
aE8WQZCVjW8bE24M6Zb48vjgh8GDQFNwtP1GTzjPTJOjtaddfQQlJ+fvDYeGZXgAWvEoU0aquIN0
nkFoQbv1JKQFP5k35IIW2FVdLyBw4HEKrMnv1SvGmhnCz17OoBLVqn1CrPkJ6IYA66uWmvBrD3HT
P9U84sOKQGuKloEG5gZJveg6BzdDe4q+42R1MQFxDGvKFPB5KER6rZ+XdFSMA5hE0k/pCr6eS4WL
9egi8O4KV8nE1Da+mThZHhVw5JRjP18RaIWjy7s2ZpHhTOCbLmcoDbZ50D3lHveO4+VTGLOVX+K7
HxNNn5kAcl7tGgWoJf8xNJtlm/JenY8JpvvM8TWA4DWO0oLg/N8Aw+wkDGUzhjaHnNaOelVehAfO
J12jvcY5J33V1CVkZhtb5CPCqu1+tJgx3gP89i00KwqwgL96TN/N6yGessJWHFFyioKBWhZZ+HTW
Jztt0axhTkeARqArl6MWRzNdoDfrRY6YcNjFMcNzQTlfe18PuiZ81c3U5RvCmcfDSsoVJGiNNpTm
36lNQhVAV5RpyP0pN48b4EgB0cf93PJpmETg7YTezwMEoX8/oDHKFZgJaipzBKQF5vlliciDTowO
o8yY3UgzsfREIxx1fUDpz2HxqSewuaUisn8CQ8P50Ek6aiaanwdVjhEgT2UVkbeMcAHHdyEB37iX
CFTfaLX1HFu+0iMyTfC2Kinq8Jl7Noy1cTGfF0nV00LF/pRvaK67mMefrkiF3e0z0lG7iQzG3l//
ePXxx9pWuwhB9qI1qQqt/mWpp1Gs01vvhPkZgifQtiV3p3a1F9NCCOKd2cLOr3E/tktbF3Pa7nqv
SZoofxuq8p2SU7pVqLROi+BisnKEPAkcqGKoiEacBTCKBN/K5kr9sAvE2O5QsngBtzO0PveSQL1w
7+w0P+ppccE0ZQG79AZfTTDscZpKDmj8YZj0CutTWib19wpwGRnAdY6BsGnOPMRGgZ/lNd41Epz/
hR9NaPx3cgGZd1VebzLpZMN+mYDmk9fmfNy6Y7aTpAtPVKWFHnvCUsDQ/QRfjWGqrEzoUvSCqREy
kI8MnKSuA9CvQs6Lzzd4Z6/UbaxDdSBClH4rtJ4Ohznv7w9cRdnPTiW1gAyUfAaPGUlBFZQmvyN3
iyEeXog12CuA5Ugds7RPoXxr+J9Usk97LCZt/7BjZXTccA3rNHentC5KgK2NxmspVojrbjg1N2yY
TciETEbThXia+DpI2IGGmNZ3havkFHEfWMlOx0kn4kf099eihd5xTDvvKzCk93RRb/FTLOVU/UxH
4jN9cZhakPA3+Wn2hvhdZFn0MR0StEUrMoeJpspitliamPegTnQyCKCf5LP3FwbIpfna4oTt06KU
ACaM7nAd9b1RPzrcEjGw3AOIKl8r4A1gjgOtouhIrIU/fQEb2CW5papjqaIe+/B0d27v+9VP6cY/
wdIKY24evCMc5T9xYCSgwqS5ttt8xN2+ImfX8vNXcwdE+iMDGq9/EBvzGyoIF6MKJXWnN7grAFdh
MbKkBDVN7Wp4pFe9OUgc3Tj9VufXedsUCQiS3sIqnJIfZpipUpC4veaA7G4oVdCGw/KoLRclMzKF
tp7/fpdGD9/2gdtMVNo0VfJZ+Wy34BVwO5feukfOjCQ+BkBvasEldhaTlKMM+uhhXlN7Jjyq7TQG
aBAw4XFks4sFpSBXuOuB4Jl63w4HdaFqT56T1nIinBmmzSNoSUL2+EZHapmYkTxG0Z17Cj0owqL3
1LH7equJ8lwFvov18asYtu5wT7s8Ti6cmRBeo0kqrNo2/8E9nBEVZvuKpoKDaivDGNPkV+bNjUeD
4Nu4BxZSo6YC12cplY31MhpdJMjTWLauc+gAu5lpq0hF7TndeXHDio0ESZVM8Z7rrUOwFuisVxp0
UEo5cVgFH85aCFSNb4INFXnEZEuIF2KrPf5mGessZC87wej75L2x81EpjXKKwEkR1dUHlp/9JzCa
xIg92h6z8Mv/mUAyn4jt/NKuaj/fX/+ocuwz/yEozGzkXzB19f7ErVFOigvhH7CQQzylLF4YCg3f
k3TtOaQ7COzkfnhx9KD9FKldZJUlJW3kB97feogbW7OIuTJYceKs6qs89b9/QP8pPJb/PYKF9piZ
kpp1xOZIswtkTSwxoEWi9rAThvK/7dDx0IDhIxNdUfFO6s4fA+T5XI/Lz3cJidBW6dIwcSQwkxFj
djGMdSkPMGQxD53IXG9jOaxpikwNTanbDPbVlHY49CYAl4QybjLmkBv02TtZJxcLkZ4SnQxG8iet
ZTl8b/I7fOsmbArDkAywvsbKDoOVIrOpQgEv4WuuRDiNJR4xR2U29N/zT+VyjssHPl5/KSRQ0JiY
wKamP+xfZp7ioimdvtAHMPYn5pfhTujXOwBLJnYKzkRhQ2a89IdvMct2LxHMK85/fLjZy9ZlB0co
LHCAcjwI7jXIAFr0xz5z23pyE/H6K56BQ+IsNxcWlcwtWe6az85y/kI2Il6NS1H7VPbjMNaOe4GN
FfW3ibNVOoIM8xGVk9QK/eV/H7hkVgJwoBLrnMbaVxVHoUuKZfIuNO/3C8f/GKEUozIgBkN0pHYo
/QZiFHggmdF6Q2UcoHBSIp+IC+3M218EnnjT7Pqp2Tt67MVI1cPz+xaFiUMU529gvFLTgvCQ4lwg
WoPo3zohZi44lJxq9fozSCd10JEkp7Yt3RmVZGgKvwImGH2Yg0iq6CxoGiuz8PH2TqNrK55U2ddZ
+TIxEyYzzgiGd6zbPWZ6SjBmKO15JwpOX0GujxyMVYUJQ+rIyanl81VRAEWOFBnTJvahTfEFSSC7
eQRZQIA65g/gPhJOXzt+CC6YKgj9mY3y7wU9ZQGFP8U3BjubZM2VdFXGlGe0wHaHafjKjmupLNG/
N7VEbEoQFa1dcaftYsgX4+F/m3DY8BQG1zqINon7mFNJjEGa5PfyXsWdPc7ZfXKGUikgaDtkcOeR
dCaKWX1rkYsnMMBcx6TYUVEhN7U2JDscY44XbAi/BJlkIlnzySXrCy/L+ZHwhfhQ1CfV8mOfwJrT
4EQcWP00NMjaOR3GyhWkRpJBII26jWlWA0hJHXGxOJ5XXcEtxQQT/lDRwRa0e1ESFsrSEH3VAnrU
Yac3lYWxNOsIiG3F4b3S2OvbjSXeGbCoHuK4amurS+vCPY9qbFWJb62fHNnZMLUFt/OLngEg6sfO
e4cyYDKFgI8xFyjTMfep12SX8CqHpqnJnIf/S+24uvQXpToMpSpsNmEzMBSjB/tuPdfXVoMSW5++
dFn2LAiLkfqo4grbWlnMiTygfrFgl5W3ngEZaqSglqi1zKQWDeO9INMHrKnXbbMNr1uW8+cRRrnF
EDpZeaee1o+vr5FcMQdK61TmRzL2IJ1s1GlAqULjOzCdmQFYB0ZeDN7uZpAWBXhdtZoX2d/S644m
+qwt7wU2Rxt+pgiw1Pu/YPb99wJTGinh3tEJ8R6qNrGVCGq45/79Qx3FMkX0wRYm1gdLMyDqZMmq
piocPQz32uEUFsNUlOfgJwOiV2CJln8cp9APfJFOx5WjcN2gzmgcVfhu5NYM0/V9+6wlMFf96IgG
5pf3rj/lDYI47+SyIF0TCZC2/GhDUHpvzL/vCDhXfLfksawoyK0POQWUzq1nKOrpLIc2yM7xzu0F
vZOJsNlfNu70jX6PfthO72EWof9vK+fStp8rIHjBpAe6ySqxCV0qj8SEbhcKZyLXU0nyvr4OY5jn
QKG4868gMcZSQRBWD68eVbawUAhV2x+FLYUNc1hhQIlf2XF22JucXParzsmPU+3OjprEPxZyAg9W
0A3bE43RkXoAe/mRwitCbdeyuEnlLKSsNtWTQcFAKf82YiC2SJVo1Z36MDLvo3RBhTcwAvOov7WY
1M17Dg86QYcBSTDAL+rGnD5d6J67hmfTxEe/Ed79s9ml4t7ocVsASDbibwXNrktrN5+GkoWzaJpj
lTH4ier9359z96O5L/DEis9xBa+sblZEiKM/BVHXnAEm6cTFh8fDBCIJh+L1A9N9KHsTpsbRPTrK
y5M0Kyx847Ol4QHaecm3YwK96JZhb6sHlFJYocRo9ibLJs9bYkdFrdYIcP/00GhM/1NmYJk7H8Aj
MmfEMpBPW+tIzwFlkZx9KeI7On/YXlkLmDe97XuRwJbSro6wi9NR3BhOBdkrWlxAXo/jxseqjYhp
yWjPb5LMFCOqhQBf63pQgWMnthfE+IjwX7xRjlxWY4RLrA7httGxCvf1AAo3XKtZjwWQIt2SwcU4
36zg5t2Pj6d293OC6hWdACfUzRpoBycZUJyPA8lcuCRzt7g5LleSJcBzah4QUZy9tXULbaIl18Xt
8ZfUjEyQDOg2Ro6H5rs77MmXQ5pFc1ayPatzqI1M0iomoROIkJ2y7q0CS36v6ZHx5Iexx1d47diM
ZUNt+Ow1LGwgDfbqr2OifX4QJxF54daZaneVm0WibUeFwjAczpYtHfl3oQdKsQwvyjKYAkpiVKe5
kVHGxD6a6j8dGhjxa4l5hVhxWstEooAVGk96pVtM5haFRZ7oVhw1BcaHq7VKlVga/eNkUxr72hzC
Dltmek/alCkCizcAZTp/gELpdRicxTfExWL78K5ZBWOfAGcljMc7H35vlqOx9bFotP6t4DHd+tAc
jUERmIfe/Pzu4oGFxp1woyXkpoN/u2jpjDQ8RKkUXx7IiHaVAsXo6UByAiEUxxakVupkRnLGvUXG
mmBz+7I8muoP58LmitHg7y/6smTAIoX9aHjm5/HtNcAGbFM6+eq4NZ2EI2ZcRlB5Tz3kPyxad3qu
eIxvQWmaHpZ5Vx3Duq+APeHcoTF5aKpFGLbV7V03uchEhUmbefAXOHPqAwGGcbBRnqhu0RD5sS7C
QeWMCScjN79jXYMZtJV0/dHyztH1xJ+9t2k0I1l8+T4P406sjUGydeXL/IGbPx+9lP8aSBbu6orO
4cKW92EahFDgrfcYwaR9UP2jW0DnENC2kJc/+48Bdn+Rh/Ph7KRfwn11xyzQLI2Tneeb9hXTxmkg
vTJRYbWL0vCpe58bKpCNLOxKC0mEAV6TIYcY9k47yMPLfsFguZefIBATc39oexOHUYFvTw1wM7zh
ivsLFNtRxNWlmwCDiZEpI3IL6mI1EcxGIU5JA3ApKuTGai6mLuFHw5ZHqf8qLRDFXq5NPjynWx/e
P46BIESFwPZ/ET//Olya+FjcyC7zXM48lcnPSiBH9MBRMgwynPH66Qyg9EF5NkTLRe5YrAoVnbo9
R70jMDZBJqFsD5B/dmzwv+oxAt6gAKVRdXRTzuj3to+EWqMh/r420kc/fD66zwR07CEwKSNnO/Fj
aat9flCNzS2hyuk6VjSrGnGZTeMfrdGNzM/oveZMESE9MqF+1Y7XMzCBvttHPF45vzg64Duh/21H
4A2uu7MLXRm9EMejyV/q/TqJVB8gyGI869fqCvUZxM/DasdMuf5fzJjnx5OHdk8Yh6dR5Akyrfqh
RZaGpgVNfvomuf7wlZwG7tI+wFMVLYF38yfJkGeYi8WaaTdfVVSHM5hHmjEATmMWqZwFq+PAhxQ7
OvXzUb+E7mfbErNcLlGLU2DBoiFzNAE0KIwuvHZ8fX0MTf3Imv/ZhRmLgW8308Bx/klsjVNdPet/
BhMalIfHotRJUjFYHEeiqTFwqmsJHBQzUrsUEp8Yfq6CTQlgQpEXjI+9JTv1F5XRYQG3zet7U9Bt
+CXgUfFImpmXSDjZOJYSe7y8jTcxhxYWxqHZrEnXUhNjzwNjUxzOW0vOTHu6H6UtkMs7UIJswbMw
dSKsUmdMZPmd7evBClITVJPdVU+zmP2olKkiPz1czoKe+WxirDR9AhXMGxtbHl/lnK6gEqxDkQpI
0VOrxg4sk2Fxjo5HPTuUFhxovVuK1AHkOOguqkUcnYVMPENbqA57khwpphaZcmVR/zSk1aEk0NPq
Ov11kuu2E4S90yNkf0OoEJFw/h85/iqnagrEzfes7CSL3D0oc3zvuGsRf3l1CT9EVR0B8zgMmBq6
FzrtNd1uFNE52jJJaSTvfxsXeOz1xMnzBy8XnWj325/BKEwAuEYrohdP61V4sHDAk/OFP4ib0A/U
iL/Z2Isv20YKXXQr9Gx+JxTSZiJEu4wC8hSWdo653YUMcXkieAR5swnAf/tNlLewYtxRECZHrv/6
mymsyb5diYYjcnJ+hNTZkNUuyzi5WY0cFYLrjAqJpkHyy3VtKugR5Ecu00oJKhVqPj4ZFm7zliD9
RCkly+MSVGNefQMNB13qsMYp4NjlHBYzt/w+w7Z/uNDIYdGeawani5kFwWrRbxqEOWMq+bKxwfGq
uSeRB9OTsIJgzDbsIYbHrxioLaF0JV+1zmdM+AAZ1NXcnMo93pH2FvBv6M3SHnPxzEi+Ss2vcFE6
rpnaZLrWr7qIyAOLkiPNMXZVtMdxSTa6wMyYhsxcRywDA6lhN3ZRWOIVA6CeyPY31KSK0Mt+paEl
FiylgprCamTBQdcCRzYwxaA6SI1uHDZA6xRc4GjNbtti13yFa2HQ5xTae6J+15ubGb35rJaoQPsF
WhofKnWA8UpZf9tShzFAK8kqI0tiAWuBmmQ+i6HTecIXT69WsTlGUGJa7kFWOpYlpPAZMxLpQUbX
raEm8kMilVfEde0k90h92AxCc+Hj3GhjLsUjr7+5RNv7kd2PSOSLhK2TkqnlbUnr11bs5fcOL3nP
s7sA/rX+FalYRcYrlwBYnElKQtOd1yic/lshDVzYbPHZb2ebx1sQqnOJV5VAUoyEHti59PLZCmAq
wigkhvKE6k6vpxGED6vz19ZrC3/0tRBBn5bCLiM6W2+VegpGZaXsSILJmwtZH63IaNId/rJBdriI
572UIVFSzY3ao6IBqbpZOo2WyiUBFJCZpH2O57ImS/8QI1QaXOVslw7QSTzaksQoTHmHC9vaaHBP
DgOouGV15MK6qzrqxn54RJ3ejnKKEk7QG7myxIECKwzs9l+9W10SeqtJMUb1s6jKBe8lQfZ93LsK
mDoECYmuemvL/EnLC+aH2uliSO3DmVlPU0oDhxLzNUkZoHs1rz2A5MnWQbStByLyAwhSJWTnHg+b
1nVrd5iWK+HyqfC0tSqkNj9gQjR+MYKV4F678+acwUTgT+noZ35MxOdPFRgJqVtl6I7AYZA6V/uX
na0DkZGtE2rWwisHx+and4pamUEYcQHVYYbmDFXosRd6CM0GSK+pk1tJsCPga35t9cS+ej66eElu
yARdnKEE0zRz/ZRiVBv4Ktm0IWmPHd+RrwKB+fvl1jSOvnRbMlXGUPMffi5E2EGVNLaWrc0dRewV
KA0nxZCZobDFVku+utFzorMskhVvdEWXzEXd4KgY9fNgFkM5HeE/X4WYe//FIXH7rSy6ky67Vhe2
EVCZFtHKWIb3DpqvSA6/v4kFBwWiLugpvRLpjqTwYj8YhzjQw1AYqaG685SBdATMrWUWcOFM9Q2o
XjkNfjCWzK3BmXOkfBnp0d78k/aCyvN4n6Uy1hMsjzBedsREe3V9BWFdD06DX8U8Cm112tcSqSGn
pFmnBrXdQB2SZLiXGmH4gXJwL2yl5nPXaxxcU83ZLCW7brM40jwf/+BgIANE6b2vzBig2OaPOeUP
dejAn+KvUF3K5McAq2+kKTBoUwlMdXyG+9jxVOzz7XmJ8GOcUkEj0qXUCx3jNBFRdS9bkiifhCqd
3/KnUBTQKVi27ebOzPHJWbq4sBBAbjq4TY0gCqFSZ3I3GZ+2uMYDj1VzLya/DpYrtTg7wFdK53fE
oqT6vS63lV3Lh7DD57ESoCVCMSqUHhIIaFMh7Kv8ovNEGK78+cVDDXO04/WPIVuxLsl+BAa7Gyr/
LnR5CBzug51IXvWzyfP/R6TD/0+1c6wQIOymPkYpRPMLu9fKDjXyvGdpC2bRyAsEabz+mmIHnLuE
EA2V//lMizg//h3nFGrnZ5oHRckB5COzbBsI5oCKPlrKw9slrkGRSz44zX6rsZndkWkkxc7v5q1b
8cjAmDUaB79VNThhCRJ7h/QgNgy2l/oab8ZXU+sh60qyDcAMqNfZwXGZXgKNMst8Veen8B7eDOOx
M3cxPGb7Z2BDfGHEVaWCpJVeuvFgQEudARVj7xID/BsmOKg/fpAsSxTivJADBox3+Y0d9OryVzpo
0P3jjmUkFiDl+nVpvRDV3TWepKVQQhnHMT6TlmGS5ek9ikilD7WYFETrpu2RUwR7Ug2Qz9tQCMV5
8ooKk00ZsV1QaAWDHgHL+HcWK8wvgSvDvgXq1jme3HjOrkc4SqFiSprBDTFG4oTxMLu+O54xHUxi
26N7TJvY/u2stbQ0Gg3K1pFgP7b+8IbkWQhikHE7Kf353/X6lOKAZ/ptW+j+3UJPKrFr8qSIu7IN
B/p3+Z5z6jX+e0bOZgpAZYcxpRROwNVS5Z4fnJHtHRdisr5/kEqw6reLOe+N5k4KU4idrF6thNyb
rX/XOg/01jXafISwDIIuxcxDmXRnpzbPprNsUGq7Qv23j+FDD13nkp+52IQ10GHMhTqqUEly42K+
nKgQ+CFl+A8hNpjilO9spyDKZ26fWgLcNB20DkQsHpcdq5tuafzZKqcsqYJTGopGCTKbF3g7O/+4
OWkwO1Qn1RbMaBOccZN7CxALXS0PIIzXFNMwhU6cgPZzbAwX9p/shv5dQ/OA6xRzzGI7md9dHseJ
aOndQxKJBfvpcYqbcHGnY2PA3+xVfFOukVSsiTs2LvsILqm5UdnEXv1lxXhZZ8feGuOB7dS7wjwC
B9gb6PrgQ0nfO4nsQNNhlTW1cI+Bg8DYOQ6P/tQGUF6+xaaBK93LV22nVU0tlf06NbUn6SDSQznC
2YeUSgTaQYNcvvvl/YGFppD+j5h0uXhEZtkVSkfSCOZUtnC38fl2ey5gf5MMtwqLxSEcbwwtdqC7
BMnFMYSlWH8OyrrhA6TrDmlglBvwhRO20kK+MGDnIPJ1GluYj6gykljVbuBHi21GXkRFroVaz3Of
0zsZ7m8QgSq3UKwnOFOQkuxXfoOsrmLvlRJ/dGbR/+DOHcDLTR5D3owuyT5X16fWBsB18RXfb12b
1AMdHbOrgvdQQweEkPp1zPmzima4qiu5t7klnJAc1GapcB4J/XqYzUjecPjUAR618iGJJqLwPzVW
zDY+m/ieT3MSRyomhMeF6yQkY8/+W8K5iHSWc75pbe7omzGhWWHGS7ZG8SscsPyzKWJisaGMUK0e
VXEZrjR3dmkYKgMFvlAuVOxb/hryXUYAuZ5aoVcjaUFczyvsA2pwOQnV/Aj2sb99nEHOjtAy9BGy
HjY9qfWopyaYj2tprnidOFFiNR8lu9bcprC4iWGzpPGZtReYaFIBDOE/QXPzUAF7pV7TyIotQPGX
l0wJZNqJSkYVtyxJdZHWTTdzA9ElRyPSLtdNJYrmgU9aEkqyJTtanSg6eWxjxlDvEEuPQHko+zCK
yDCe066QH+iIqxyuzF7dkFbuC+saGHpvPXOEcJ4tfr/h2bF19MxHocyHWm1fp9mHgSMbZRRtH8gD
b08OFyTU15GodOEEnfiCGrCTV5uh+bBiKWSAVJ00Q9PjVXvvfP9co4L6fIowYv2WtRQsqy34UaBW
tADHuXLXjlqIBZkob+pKmf1Symmw8Ywab7PRld/hNKAdpdxbzPei/XwCE6VYbDRTrbO1dOarbTa5
WrFPiDQ8nW8JfW/aw/2GNHWe9DL8OSHyuSQQ/v3jz2DAB5qUYtSmPYYIvmbBcz+vJRQ/l3hV1f9X
BHMYxhOWo0BWrZ43BRNGk0zeCIvvMzJtg+Wv8R+FE0QIKLDftzccz4eFXUm/48d1gSLWISnrI25/
rmgV+HYJ6JGHeK65uew1rv4R99Az+YxCOhx4ZA4HRkfbvvWstBHp4mgZwtqecgIUayZhvTPJezOT
nXm3DEMhDcOvCDayJsOWXAx9RR8sMtDy3CTqTDfon/BojjDN/1iQb0A8SEXD0v1SK9I/psvNiEgY
MDuYq9RCSnLp4c0t9YpAvOM9pMUJDhyrklRs3D29DUwyB3ImKKxmfPL7GerfyLIb3+CXDetMyiFJ
KNpGGU+/ObBs6aswxIZziNkT7oMLrM+kfBoKMiCulgGdpBsn3xScr+4NBbol7xlmQkW4/MmKyYDe
Nlk1JxXKmS+Dc/g51Zz9eBGGC7p67IefGpP85BlewjJuiWT4a/k9+tITo4GEjTYet60hsw/qJTgz
d/b/UO9e/dU/Cd733fMK9Y6+hRc5FrUgysUKVWPQBWahxgUTm6tnVu+kWK0QyfptrAzb2AL3ykmv
ozwaD/6nynOocHgECCb1pBznqkMkf4hZxNnugQ1s/oSQNKzewaVM1BmEPQs/TkUftYFPzO1yZTNj
Jy6t1Is0BnhGc+8Fasyd7A7X1z9u4gjDhlYIp/YRxKSry0+0NtcOB7EfeoewhZJxKxSBTCT4p6Am
HHwVFUvLRTs9eafKOJ/qAZxYuNJD+zcRaXxCoWQqV5WASE2qdFL/RIIpw3lqpNk9IlgbAbzm++SQ
q++qtOduf9Q8tAu2NSU7iFmatVouXMJx10Wx96mNZNWhISEvVErDtAe6uvM9U+JdZyEuECRM20d3
RTGWOoF83oMfIEeNrq+lGD6agv1twlSAkewrxOXGFBXjjUXlVNV56bnOP0WQnJSO9m/suxensD7Y
ytAuS6FWMmfuZZJkVha8Jo7mYVN14S4qzz4bu5MN5aQY2mUDcdP8nJilK9n+Ddj9ipwcwPG+HyrK
wBbtLY47FrM5vHOVTFQgpLUZXyfERaEY2DDm0pIKTBFJaR8H6IoGACnw5l5Rb2xViauvu4BBFVxg
+Ypgc0V7NiKdfJutzolE7D8oODVne/LiH9+KNT24taTQ39RxOoN8xnDCNzl7GPykG7JEBw6xnLtF
t5bs6vEzOJ75Bn5nLAJzzgqRcuZ225GXDQsfNT5TJuAJkz8Vn4u8yR3FxVaPcSIW572PoHjHRqsO
PBZh5q8pYkCbHRxlZ1HFpNY/5ZMvvTUggZHrHYklpYxajZxm21ArQu5spCeZMBbPzeIlL8b0WF4K
Pe43eZD4jNqfWhl468hEbT6t+MHd5gSLmC0I1IgZNdtsexI85g5AFGXGtnAoIt6H5EqOdXZOpOHL
aMbefUtEfMaZKtvdzou7UsejL0BxMyR88+3Rz6QqI0yN5SXVmqDdFHNlkyxpyjAXh9DHy3qhd5Hs
w89zkWoVZzEwTntGJM8g6+lsLT4WlXgdnyp0O4OgVm5PVY1jBKgHq8rOxkwm5O3ezTNsdT2P5VsN
HXuX7OcqgFnptAyEBgasPraPrYdBevu3anLec1745310l6CoTP88RIVDRFEfDSIAA7Egzmg9Gw/O
uR3E01fOzODNhfD4TTSg21xTDeIwZVscIVaPcmuDVych76SfVJDAPojnJeztKnY9c1Y44VVo764d
B0ABhbnQCqBcM8G2xy5dv6vJhrFbYe7SXqh5+DEQJjKCeaImrjVqg73idkBZ+3XUOk9J3PLdvkeo
qTONGFm13pwjMCZN1cIGZIIZVunu6ahstmYdhAzA/ICQJpFmYQONiv3Fa34xgDdZYvWOY5rjw0Xg
G7p5rSibw1dA+d8bcFIlaO04boajfe9AJNSmbCBig3dGoHloIR+Kx8CqzVH8wrrS5k2z5V6KmDRY
3saoYGaFTmv6rlD6SaH9HNj7if9YwJVJGxVklnM6t4geTJ83GjxgD6/RbRW3qIjbAmjxEUtPvnAe
tclYashQ7jLqh2lR66CD7AIt1SYncWYVu8GXGB0OyaT/5TsdBsJVL9Q+tAYEIRHIMV7xSk+xMK5n
JX95zEkzBzk5Dm65GE4U+T2ak80HmXfAXl145QxoGYhwaQCShbJFaY1vnafPjYWqR/R4ioV0I62c
xLBcWQeP/03t8rIZkY8/BIuk2TtQyeiKJApsgGWAiMEOY9Asnw1/U0vC7b8Y8m6dhcCDuPsYxBNv
JOaoTo2TsJtm7EGo4huXF1ASLpDPtOwK8rGQqhfhU8009zjNKPx2rNdJiOUDzmQsy6uQWoDlPfB4
mEEzmJ3yNxJAUWTK7NkzbshFDyzA5vw9q46qB0L1oHWtwmMcCmZ2H7HzvD1EYi1MB5f49zDSnInm
S8zJvIlh8po5AA/5MlrKwr6SlIMmFyAtQrNlEGtTC/5hRXP9wjA6I+A0ByfvfRtWDTpTMUaK/SRB
y0limbaqaJUn2XZHhQlPlJa1klD836TwH014Rs/77LAOo9jj0XH7wfjq7EkT9A1Y0XOYvWT07vPI
7C43HTNg2+cpJ0MhvGcIdc56JKUOBQKCbJFRtQwFrbRr1YbG5+GCLvwPMfT1f3WYaaBOa0vTHd+E
lgBQX1W0MegLXugi3TNDzfP3VWE/Z7FDAD7bgHuMnplMiWZZ1093TiX7cmWI2aouktZN/Kj7qKTh
zO+7J0UJ1BVUXLRbNDTg70AggpWmEqIaaHxgOwzdT+/446aGg3koeeGK5KR6GbUd074jtwqLLapE
M+NDY1AHD+vFWIq7uNdr7iu6r1igLA/bdLOmyAwfhFPHtpAXfbtCxaog1HG6WIHLjVocdrkkOJqL
IzWlyvHghMjBc2igVSER51+Dk0gvsAGMpkJxdLSVH+xGztU2CboGmGU/Eif8bAlFnYyDD91ZIxuB
suo0T3i4saELCaA7N6CphP8II+bWANkUVn00HmSY1VrMv1KyUHXYqGPoJPNE64X0HchP1wSCVHlL
W1++N05ygw3OgFOQnB6SpEB4pWLR20pq2m0YQKNtLiI61me1mTg3wh1PFk0Vl6p3+qSZS4W0th2l
Nvaf51mlvtw0o/Lpp4VM51MwoQ+oIDtbAf9b+IGfNKhi0qi0oAqRBTYfBpMcpYA248bw2Kam+dzV
422Ok9H/P1oqENTMVKDdp7U74bMFwqSiHD4/WjM+gtKvFUj0XplsdrXq31+lkHSOxArXffl2tPR6
KTfe+HNosE9Q82sSRnixei/l8g9IJpGlO74HHhVq2cv3PzUjV1UcNTJeyZn1O2BzKlfjnB6f1MRf
JiPw+LiJB0VrkbbFEWIR6whj/TeXXAVDFRuxpKT/XyuHdKdO4U5jDK2jPiDqt4/dzxURj65ZamXA
B0W+VQQLEVRPhdQhhG5HooMBpF+fcHY/0M/b0Gi4SojIlcqHvYOUJ3Jo13WiUZM1/YEK8P46tNF/
0Ygo2bqWBIXYJ+V1EYZslSlc0hPm/5rvpopRhgB2oadvELcPK6rtd5lYrEO4OBtrmK8ZLNYTxXYg
5zueqRi/QFiLsdS0H7rIh0vXKpHzs4TsCwxxvbDhdZxaZZhoiV/QID6V7rPDViQJFdYIPRbk272s
Wl4zQ4Dn+ZK4ZAqoZZxNgZPDqr4JUdiS6vtVfidZxilUVHKRaBUc+vnggYCaC0CX4BxAqExoPOAL
PqvRFm54Wwep4HrPkOlkCgtiBUsI5kHTcD/HXYcOeAaMfIwJw8C9+UBC1Lf029KRkOIzZ9Vbqt+d
om4qoInLkOjAc66e+v3dNDcd2AwTLisvdgjqWVJ60l7gho1K9Ou9krI6d0WrFhdLrrfEWWJvNy0U
t8qhwQOfQm9Xm/OzBZ4c4qgzPiJrLIUvhU4ctDvNHm1+5IHq1HFwwKnE0dxZ9nf0T81KhPnA7sLD
nn1sxLzYk6K3zfz56BfRvnl1HqRxG7LdD+GZ6zEjn8MJZAOGq5kNTntL533+z5JbuyYbJW81HhhE
Hx6zbNbTCzIKkaw0f9DMlF40MQyKk0+nn7lxqjamQTSfPWP3xYUhqM4rANr7E0WcjcZr07hy6u59
P3DDDmrtolJXb8lInAhh91LsN1M4IJG9kGuiF01osodSMHx9ytCsp3efzIptsop/jROtgYNfGXVW
sOtrbj4uuJ24eBC2OMWirw9nWN0wcl9QyxsZcSQb0T2larjnR7FDQXrFA/vMUrff/u6AqjZcwZJs
vFe57RNbGjH6TxB3CxLn74lnBtdjKbysT4Kkian7T5zKcI/cL0aICrhGPksvXVBydUxf2/AWiLcB
OlH8/inK1BIZf0V/zoSu5vQBadtacQW3hAK0Cs9Nb9O+lnSzy+m5gxivpHhQStJ3RFcyD1l7zzi1
PKuz2eQ4YKjzERQh4U+4QE1pJZOYSUbL/W1maZMRqVi7orTJomLI7OwrG2j9CLlbzfqE/rtRBme1
vCV8UUFHYg84LbI9NqnDflkiIN29qFYj/IbvS2X3OCgKQNuJMo7TQ98T4JxpmvYQEkDQFXs1QwmG
fjq1IKNepWSe4Hxffyh0usMrT5eN1o72N7ZKeS8oxEQgawuUFXCnypE4+qK4Necd4XYqKoATeO5G
YrXeHKMgHv8PHRi2WrxmyubLYjwXG6P/Og/zbNrqLqKGKTfPlk9sfmy4nLaQ97DSIAZdk3ywC4Lw
/ONEjw9W4IOA8kZ5DZYtED6K4yIu5S4IiUIZGczhS5OSbQ0vcuPC9fFReYxu/n8Mk1xuyUtg8d0x
Ip4k/zmJNrtmRD/SogTyHTGk0DaV2lfprsIbsRzJlYtprgvLzvozYolxXbwLXmWia3zjR2r7Aia7
Wp5cIx8UxW8w6rxVOHxOBTbbGYWFTbF9t16SM3MyBhs4QiOsusvm3ksZAhqjMaWIw+mDs4YBVP3K
rByO9dIHfYfHqZk0UpTAk0OL2tNqE+6ymQ/PrORMfpjI6kvkLCy48Vd1y0o7f7FDCMBspbz8NRi+
or9E8BapsbG1chlGd+rrnr6az9beDd1SXrz3Ru87BBL5KFzB6VIHZrOTL0R3I1JDUNlAleEkj5gc
QZE4UtI7SwDHTkHrx0hHqEwGtkNVPT7OlYwTYSOLNl8GGw6iFx4x5JNC2tsM7V1f1o8Ifm8Dxlxq
AtVUra2FzHSTgGUm1rW75Pl3n/Fwv1xzH8zP5chw2ADoUrM26Noz36syHPxs9ySOVPAabOsOKILT
mUO6C+8kfktbaMKn5LDud/VasM3FvOHfB9wiTgJRZECO5m/P1V3AuBUcfo4cPHBA0HaWeruytcI7
h5hpYlVRNKggVH3nAjiEz6tj8is542bEQdTn6awkF6lh6JsNuQ/WK+AjPoLs/L3zRiUARfEtNmiP
/1SmFK6vES6TyJtYutQr5CG6Vaz19HRDan7ZRkMNDpVqK701wc4N5XXQLG1oJKIi8Hxo6QVeJ7QA
ZcDfrbN4jridoba/oupNkeMXF4T7Ik9T4ocLcPZaPrQCeDdTLc4R/9jZ3WTXoKcaI3aV/GAxofTo
1tvGGGo1pUhKcaOw/zlUarmI1q8pw0M1H9sSvuVEzKtVejz5AxK/NlmFJWboAppiMPVNblNpCaie
MJbTc4iv6LaeERfyNx6dAHlFMiodzHMmxcqncN/nqLjfQKchRNMrkfgbEzMzSIxMKfOXfJ2MdSWt
7cQF7xkcXGI6zm0KAsaJzXbSuABj1tadW2FalnwlLMXSgAIe0rQ8V0AuCyv0GM6h2+CgwQMcaf9T
Q//5m6dXH8angpFjceB+gQqyRqU1BJhqiJeRiXlB87MQHG20cswnfEzEV9u0MBHhtZQnjS/BdBHP
r93NBzUHTr3FfEE37jPxc9p+chj7Ipz1JsP/6nivW5dqfXv4CJnFYbsqxgMWC/mBj29v2YcUVcWQ
2vmRs3GhXSdrUwPQt81qAa3XIZdwEfVVb736enMQv0pY09aJVE/fr9/p1Ufj4TfuqEoGmIyKfEri
tKuHSnUrvjgwn4yuvQh0EkN6IH+pa95mwK3xXwXxYd9fTZYe3Mdcy6Tg/pZ1tloSiOow+9UsnAwD
RectaQNdSQGq0pPTTWD5POdRFZxci9auG4E2jP4uEJzXJz/JGPfmi1hVEj2n5k51PS18wioIQtui
KeQeafyBKzyHkF5u42Nzov+pi+Kxikos3oqsvDSbf6+JGYk6F1ORfGjEpLSbLquP9Rz5CcTpmY5D
+bfdQQQdcekslY75ddswR7LsI23cMNq1OzL2FJTJb4+S0/gGoVayeJg4v180/lBK4tJYt1kwHNd6
7Oop2LbgtEKBEtU+ZUn4RRefUetCstGUHnTuflDaeoECMHhkye2BKO6Xut9au8/q4im7uznZlmYT
YyL2uGmASmg/zpr6pmwFje+UdR0ERRgWBWJ7FqNe0qlPZ/3KLAiZCFObVB8u8Stvo0tnEZnhCBE3
b4lYH65CztAIZkgtrGMH9xua+WvKJDGbr2CVokylXJiP5rlgZNk26hApDW+FVrrUn18LD0ucmcpy
sAM700BcldVQJ8i/nNRciAJiwg+KL9DlyHX8+eNVQIQRlfWcJ/tStBEM+IdC+Cf9I8gv5X63mmoH
7U5cOfjYi1vF1N7a8PjBTuWNkbQI8fBIjWAesaYShxIokPfw7QyNyUV7frN/MzpXq2BLf3XhIe6U
ssOSDMcLh2yLPMBcwBnrzOps8XCd7dvfPU6+rhJ5WqiDazXttFPl6NNu27NnzA/e20C6KtPZgIKp
AxoB+1Mw07nPgkBYFaPEppM+CMP9tr1WMDZZBeeciuBfXI3/2z5hTZ4pkD73kMogaMeuQXds6HdR
5AxFG+/o+3aCu/SZx0o1Xzy1aRf1KhaTsMpmSshQI5H6b6T9HyqxJqbt1mS+ARKedrPcCn2I/nFu
/oA2ch2/Sm2fv5NV+Ycb19HCg6QYhHdMnUVhFp+DJBdThO1lvzasIhdQ+OxOiUAyHQcg69krw6RJ
Rk/aK88mfXqmH7aBxCwgvBICvjlOyRTcAwztBqI4vhbwLFy1TtbhKPC8mEqTT1LV1r+PStjwfQuC
zfQWfyee6c6PU92IGbSaFbiYYeppkPp5pjVjhnSs436w9lz9TD6XrpaR8WJldLIb5YgLtE8vq4py
Brf9PLyIdx822TrY6aMJQ3nvfXknzy3WuLCX9UVgMJKK9Az0/yFSvId31YpAaWjWNp8NE+Y/2/fK
1bSjWpGw1F69Ono8HtGJLK54Uu4fmbaAhJJ8uAJ8GqLPqcScXPldIkPUum/QZ7TRnAmtaTtxiOr/
LrB2ZIU4F8SBBCU16iotOCspj9HLZMv1dcxHrT6YrYtGzosw6b5vuJlF9FJhbyvgEwbt6ZON7Ima
W4b57hK4ThscjS4qCmFKdeZ8/O4pQrNo3Eivcw8tUHZh7EZh36wYtiwAkK/fm6mRQCPoF95jwTe1
RWVVmhqnXEmEG9Gjj/wxly525r/zPiF9Zzf8yAv12wOaHno6bGb6uo5gVB4u7ZMzPzxbD1uirBKF
5PpdoMQ072wNyq2if/rS4a0kjSV0WDW4P1dUfd5FGvggMBDaYxijXu6H6r6SMpM9Wsu+xKBl2PYA
cN8v1Vsod6yWau98Oz7z/pR18B0+twhslk8QjVhi8U26YGKm/RCnAY1SnkuFI2hy+QA5qDhgbQ+a
WWEHxKWMc55sOFSRhPLlp3SOkumz73J20X42jaxfMeqgvO1vzQwNbgD4mLq/mh49wIuOHvXnvfC2
SqWYxHkgN2geejOmEa/tQZiN+tJ8sgsfepsDSMxkWiGhJXa820SiKlHA/9I9KU0g9nM2MmawgpBX
scblfhBHcJFTiZAUF25ditk5cBbb9GNBigPUdrVdMf+678f0JOQOn+3+reOGDVi28Uc3tzZTe0n8
60QvCL19cMu/S9fyPyqKSN1o6f7U1ksxUzicItP9de8GQX4V8YYr3+71msoxAoZStDP3WuELtz77
3YmGmaebnXpdBuXfFN1ruLxMVlsQe0B+dodasQOP5fCs5zCJ3JcKJ4H3/GlfdTAbEzEZjNl51kE5
jB/NbLkZrB5ACWBgVfyTKYDrocOxchVrekipf9ipvvsq7oGaa7YpbjbcB95lK4a9Zr+en60VneR+
pBS+Ubu3fgSQ5fEmVQCOiD7qVy69xcQRR300/5PICTgu/uOzRpVtVKuC/NDa3/PlYgW2dF2Jjodk
H7FL4JBamsQt4ear5Q0AdO0IgbSFU1XvAU5Luwu8hGnkb9ot5ZnbG2/ilmIR715dr2DNplRs13s9
gZqNAH1aMVe5SW/IwSTAJ0uKI6WZJtxemo7T4Dc3TlJ9Dkt01/2rYUJjokBgO3voMd6gyrqJhEZj
TpGK8TTYV9o8wdcGcN2ha4mI0URaLAL6bvEn/z3Ymi7Yvy2IVaMNoaQtJY9GuTpC5zbGTOQ8OGjv
Tpg4QphTY4MQ6xjS47IUIAKTrDJfM9VAOxlWNgCH0H3zl8lxTX/U8eKWngyek/so2UfB4HyngwXz
xMoxrfshLkeecTzS5rAf2LWIfyxHhsD/kafOPOfYk8d7ULZRCzqv83d7BcQJjH0OjkNv/4zH7Zj8
pG/791s30ie1O8s0Upb00pVALAYuhpAQGxIEs+LFN6wzgQgU1LK7rA2InUTH/2vBYf3ZDbksbk/+
D7xJv8fhUhzEi9fygzfB/HFcD3PdOo6SNSXQCitV+aYqAm+ojJjSbLwfw+pj6h92+ulKiczKdQ4I
0sS0tjJgBJomIxlU7FTszsHrnnMfG9T1b56c+33c6sQ0dqpTslsvGD2hE/G9zppMtzOHBNkVJ2rX
tumima3ThDd+CgLm6BCPrfo/xB79PTxqjiRJZJeZhWpoDIApsEbkXd4l9Z70CkkkjEGVhkxfxnUy
BmjN5+Z2sjBmdx272PycUEeRqkeJZGzvrVmhgwU939LlvB+zhvNyMO9I8TMciaaOixug/1aHE3Qc
JDHucoLg9vh7WAs1dL2uUzSTZTqxrB5W+4E4U7t2giaOrL2KkWtW9xRKAK9KNvIU6vFOTu9CCYAY
yW5uiORaR1LI/BUPruKCeSwHUAA2ovxKX08uGNdaMCVQkvU3S3p3MPGhwRefUy6PdnPYr2wFIDDl
YqTeGIBlJ9r0FaP1yJ//IZrWM/vTU0CkeLKcMmiJ1rg7p3xz/TSvmr4orng5tWKoyfwvakIsgvHC
ox7NoyFu4KmHExsE69ixw4IeIYF9XGE+XxXFqHDPSh7sspPVhjb5a9qJkOcARAFSLdRWZkyJixTH
XLC+76we7Br8uogk1J3+pE7n3SMUVauwI1XyjSipTPjt2tbwys/24ff2U3Cgmv1bKoahpLEajmtr
1y9ZFO8MSfjwX3TYDbZM055i3b47l6xm/2i1Wwkx68Nl7eRgNjxCALtVeVVRf9ljbpkKNQ4V+QFZ
5U4MLq8lo92vJ049SDwTM5aUAPCsTXpj7o4gS+QndLtD+SYwhxmf0noWDiEK4aKDOi/7WalWjBIA
Jnqqb3euXaa4gaNzN7gtLWg0Jr/egPfNLtWF+/TdEc+fth0cpWEl8VfFHGe0APoh2Yov6077O2w9
E77ayzAuyHCUImguD/alMIH/ErVtNr93KPDU5aU/+uBUwtNC0HpzpkmnVOQSUpOB1XAH6MQcs8TX
UJPVCaKgW39qSzL3vYtcSmhy9g1UqqA3DWInkpqzP93Jo/RjlNSE56dqPydut9uCdvjpleVjWHso
+lgqOCWOk6uq2Ads3P/zYQ1CxZU4k15cJfHm25LHv7j8PjKnC6moOvt1C7aUT84Q2YaZMy2jPxM4
NIbYLP2eltBiu8B+tctTk8R0TKTayOgqyC1fpXYt0xwOnnAyay8pzTCzsBC0WGXGBlkhPKdz/dxr
phoXXarQJ7XegyQ4RlZ1gs+vQp/2iUt4fJEaA8k/Q3aygUetwUmS7dYEU+tS25pcV5FLvdDynwal
UqDNXuBbSnBXjQPuKitR1cdujX0dpKQilaj1jXCxSSPyg4fOGMPUcfSFKAYPBTWWQn5m/pHAr+59
DsPreynB1YqgzvDzDN4kvxHDZ8oaR/EoWRbMENuLu9QbRSy2dSmC4+A7ow5evORWkfspkYoWSEGC
8Vitx8EI5DzTvxPjHnrzMmB1Spj3TDkXHRBw0tWD7Q9wwaTzmYegfV+KFLVlqPSCzp0Du9XUeMbe
q7ZrGW7FiKtgX8CspOQSPtRt6X58bbLBx9EHX1LDxvOT7N4zYP6x4nivVuonEyC78uH1TZp1uu6k
v182KQwmpkIRLcskKgSnxFW25Ey8ZC7Kzdx3N9o5EkbzNL9hI8f+j5tzKJSsHAbA8g6oYHbWfaYI
R3dwRXl4uf5G07slgIVWgIzVbCvaMD+Hc1FRZoQER51GucP7N0FXNuPty5zKE2n4E1qRZU+H25Kt
eI3Xy9iinqrF2P6LFRFYfq1sH4+fDMLJtq4jlSBS/VR9Z3KLSMRjP7o6QPYHuaqZa1kZ04WAryGB
fgW57yYXz+187Tft4IQPi0qTcmB9FBU9HLiEL2iLI0c5NfjTlMgblrtQN3fyMUirikPfD87HdwmW
4D1hT+fYVnfzydI0PvrI6Jx2082Ru3Eonyf4NZ3Qos9lBfZflWK27HCTPkegE20zt+XPzCLThXpW
WauuuAzp6zoW5jc5QMEL10z2s2cyIbDmKVzcRMtnV9U+A+sRWjBumGEuFink8I5qQcmS0EdzSU9v
yTJmE+T0iQx4bBKlEEB0srFrFYPnOqO49M7EDvLfPpZD+cxl7B0hG0j0u7BTgijNsP9erAIUaV/0
2gn9IiWfkuh1ej3ZXCMr+y/OrEFKwiG90m3PLEaqFNPlJSae68WDgAnLXtdAPSaaKkMVaUIq3nar
xUH7T85Sx9k5zg2M9pr+1htuVUR4bJLtjo64cOMsz9jCunTBHLK+W+LKD4STkFCQYwyh2BFIIwaf
PHY8G7nebWS6jeNNU9PHrvIdlMJCNtI/RvgGf/CIhyoHXCa4VfrsobVEktQBqhhln5Q7oLZhbtdd
5ktrCE2sinKqnqGZj5dXScufuvR+sknwDX8T76Vs0HDFTI4IcBWyh9zRkFHqGiCUq16Qn7rfs5v4
sMaarEVIUzjLfgXt1l7KRQ8XLq5ak766q+RkCNzOXd0Pdb/jLQihQ/t4g/Utg9mGcj158jurmA3w
QU3MEjLjJb5TJYk/Ft5Fy6+rShlxNtke0XdSBQX6+STpOXpmPFxAAaTHBGnty62dWtVvaEu1/8nF
iXbCuJIECzMyRlA3vWOwJj5ro2Tuyw64eZDH59QVDsXbO/6fs62M38L4iFlHeXKNvVFNqJrQpczr
5q05VkDYwq56fZxlUnKBpKDxtjj1LHN8sjCJuvgSNMmJVKf/LnfGbzdxjpZtNQ7E7ZskOyiozUGG
dWnurD1W3luc34PH/ITNSdktjgtEgbZtip5f77Lk2TDTLv4K6ijg4TIQY6BHwlNI8P7MIDYxEYn5
cm+RweV7gLbWZhakWiUtdtNDWV2EQUs9gexI782S8XXcGPD4fwOodDq5LqbJDZWZPDmQ1xrTRubQ
8HVYPq6hpUqESiXyDOaO9KonlUoQBbYmT8E0DSiVaE8yqf/eOyKzxgobsMQBX1iMBK8sKW9x/Y3a
yNYGQ39TyvAWJLgwwv8qO1fB2WdY7oDGJSJXC2tQcu220oXB1bjpJ9TQnkiQ/fcJ6HAYaLNWPt+Z
+dyw01vvzkox9hqrOzEUjibCua0Wspxg4oCVGJ0fXQEJIQsuwTYv4GLfPN6P64D6h9louAnoJ/yT
AHjTrIVZ5W18G3GCyOUY/WzkNkIbn2uFXJSJjm7hNnxXcRjSdNTcUPyVOD9pSk+JqMA8CUEekAwP
xPOGyO45hpcigsWSNX5DZBgcBKS6nqg6kQtaZ/bSKzMpkOSgNEW3bryeyBRfs0k5VU4K56A+yu+O
LvZHHh+5F8MTYl9ciDl5VrBw7E5Hsb3fBaXw8g0QD8BNijzv2i2UAjjYigjJb+TX4BxtBLJ68Ms8
EyAZnZe4aIBZgoTYg4BzWQPjnnru154b9r+ylUtUr8R63XXUgY6CQeW7+QpTZEYn0wV5zhOJ+BVz
9C1Cl2pto4nGD7jk1jRl3zK3CPjfMwyJCoXYm+ghNlTOdgg76iTnf/t0e76jZnqTTapotoFexnsQ
M13JnJdOEaC6xrDWzznj4GXKBYG79BQ+ezPIFw2IX3PkcIJK+T7IjMj/y4MjRnQn9cqmczI375Pp
fNzsA9iDp7CFgQVvHPehh4PFkrX/gdL1eSR1FqrMZQU1/3SoAgutfQr0KaKXbhCZB+MeuNxEye0V
pP6+Yxw0gV8VWUHSDLRxcd2Sa5OMEho5D0b7LxfdR4811PW4/qHWF0i7EZ7i5UUelwtV/ohRsrxA
muhTvGqOKQbr0htAMO3Tu+0rdRrKrOA5phg2/IQrOsR/ONQeJ0senWBvDTr4RO2U0J30hcp23kPh
hFxAGb0WSG7bXb9Ih7SNwHS9VphA7CymBhMS4taCXgWzJydQ1Rq9GHQC65Dvi48PAbfGDoVo45Rt
UWYOk7UHUP2DOf7o9l8svFygDPjRKcq8zKr5vaQrKB1bRbxdcYgs5woM9JspBv/I2C3pjG4XzOjw
QSO/hgPQM0zUnNwbs9StAN9iCu8qDmimJ2SNT6qjVV//D7G5fzAidxOOMzQy+IKWSiUOMtIu6/1l
xqR71phgwJ0GDP3vbX1BTMP3pFkR8wwJs6vMFDlpnmikcofkoCosxCCF8oMuWnKu11OWAnRHeoMg
u9BlUym5mN/Agc59i5xSc8YuY6mSjNQLa31TG+FfntLFL4SHy5Bd3furyDxOQqR/yHFTXnKzRqop
8Oo1BE34EXq0ECBsr2JAq6avrxw67Q7j6PcT/LEBFK98/OHInn5Y2WwqbqsmVMtH4Kk6zlzOXZPo
qWyTf8tKtcRNGuWlU1OWvizCPtQUrD+6IUBylGqAPrpcgBNmA25wCU3VjK23nqofIDEzdHty3yl9
o1+Weu6UkPbPBRJyohLz2TzgtjmvXGIaM084gBsLLyFmgh+fPJJMGBifWG1OqucvV5fKjHUzsF3D
0QtGqBUv9+1ltOqL9gp35xSUScGhHHVm4gZ9hgRJYvstnAm7UmCBZFmIbMgQY36IUNBREOfviIkW
b1C/Hzg52DWmhQmnKdYX5qEw9YsICfAAL+Ng+AFJihm+UndmCqAo/bX/0Sss8UfAVJlffzht2eiW
qzqQOMOhkJXGi6NVdQRb7H9isnZ51jUp1q5CO1PN6DsI6ocS4GJkN8eKJu1Pj0TZ5x5JFBXEp9us
Cr7PGGYGChSnN885mef14Zs6arS6KH28dSN4hkplDvC8iSh8nkuOtG1YDRKh6aO4F6nkRDiR03Wp
alrBCnqTRDPc8B4XWU7ubZry52OaHplkGNrB2Ev1PqRtlNnfYnk02u5MEVJL7CeF4lLRbsU7w5Ij
RE2tFX3yqBSz8k5HJg6B2g67Pt0l8RgY85MPjDw/Vev/xPWYzAc201LUbi8rzN9MCtlVLIMQwCxi
PGrW6FvS/aZvNa0PauBDaID2puX/1cPzVsYijDqf1yzsKYybPMz+2KoxQNjViTW9jVOXEMAkiiNg
zcm1nArCUKsY4uKvMUgcypHqr+77dR9kue6bPGXE/06oJ5NQSVqqQk+leEHdk+AJRdIhXNFxCzkk
RuCuYkd8+ZvwpfoJTjzmmdUng005IOwJPScMRvfezqcuVLIGMsmXNF+c/cWEgJjdV0C9i9MlwAq8
fFz1XBN+320Rlcn6tqRryWpNh+bEj0txRFbaZUK6zgINguQvNKmX7JkRY+MBnsQQqkw8Okf6xEP4
6w1E9SqPAuxpZOQa3NkpbcfA5UP7r8SNlMXxlgVA2mDx+4gv9d1lYa8efGAuytyJsY9H51ciKTb+
IWyFdzJApMEYvJw6QWLA84jvzYHHdCCB+jCjNreqA2kRyvXG8eg3c07saOV8xTGwFlZpWlEPfmpN
bwPGxEjUL/CnBPzP6SWS3RczyO3wR1BYgiewNCqREd1w28eRCK4gTSWPyWt36sotiMJqfpVdJinB
ocdENslB0UQf7SylpbbFkxoSlR3h+SE4xZxy9dbiwgju4EmD768dAxBxSmKqA7uVfGQxyR3ofopw
EsQTAr8i8JB/xULAappbYgnDBNnZ6pu0C4i5hrm7QqJmBxQHYQpayXB66tvD3vmIq4noTz782jIK
k4rDzWZl/rr1F3jT5x8Nmb6L3JaTENcKVTSciF0nQ5IR7W/+9GaOulaphz26FuXMs5c7ZhCY7QFI
z4+tbvLCXZSerSD2DxDruyuTL8tGmWpa1wMqjnUtpFFZC1nehuzRiWuBWxtLmMi71iNH9Id2C5eI
nftkBSJpADK0jRLOqdX/nOT/5XC6g+8AaBSN2VWpiYKmh8gPXdnQGVBg5ytD/JTRtrhHWMLwkPwL
TeZPJFBVUq1mOnxiaCfmRha/xdB250OtH6/smtwWH2Wrrtd4c/JYmNxHtnGf5byjzCwVrNX6b33f
eym75QvnEHi8pKBXo2EGc6CIKNszNp2V6CdeSHDgIydhbWWHom/Yw0v6gfHMieWnMlYnEpxGmZLl
JAdMuiSvEj+mBzLsndpc20/PJAW1QmAWdkls4qQGMbA9NxYfR324vDUw517awNJ5pEAU5Gupwt9X
6JycPAmOK5RA7fEd278SJXD+0IXe8yEkCk+rHxoMNRcUi39Bs11aRg08GLtHVbqi/93QZcxLfGe+
PSQ039Yiqyv/1Jbrn7pwz7Li+bgoQr35MLdg/tFljZkPx+YcUAv/nvoQAkz0j2MO/NXJPfmdM8aa
6VSs7TVeBIZvBm6FUIXT7BeAzfxRjGita1teobvxK2M9uREzFXrkySmFh68rREEu9fmvpbQluLOE
zKAax/qFNvptTuzdV5EkUCJdsn4V0SIlTT7yeAdarSRgzwm2wjuxzmaSP0Mmg0uenthu6XHeu2Zc
S+oWv07Wn/jscNmFJQdA0ujuhidUFsl+Wdw1vIkThX7+N9XCNWmkVUvS9HXDOYlnL2saZv1M2WFW
3/+jnPcZKOoev46wSBN8K3b8lGOf3xSn3bSU/h6GW0A4Pe/GKnXsr6Ztm4AFucWfwJt8B3zv3NjE
xuQjrAhQplJxCn9FkNUQvHZMCuTuhDIj1AO65wW23ylm+Q/Q8tMHoFXDvsbraW7k7N3tTJkIlTX+
4UH0/Qs44Ie6Xjoq8u41QpCtk3kk9yz6yuYHhhDntu/6AzZHgoFdRo8c5JMQTkRLosLCcndJ68U9
9pHsuC0zS1p7rmTkM9LBGCWI8ssmcdozFx/qFMmUODVIaxJEHsu+vdeE4NEMqonaqL34uAtdoUK1
u33PXDTsTYnHFEjv9PIsNHXNC6gJqqLcDABWZp7WKfwTOkVfK7k+nd058DttXLuUFTgTOp2PH5PN
KMvBb0Y+YvnQ4S5zapZXBAzeAV24dguyc+SgXuWaiK1sz1lQEmXyltztqY61DNuggDUEASFcP7tK
nQJLAzCnGhG+TpsXSoR3Qv7HkdOJ2dkwFs2vrEw5PsthOCcjz4U/C3K+UbNgPbjq8vO5iPEVobPS
yHlxyh6QS7wx6A2ASaJNfzeQ6FuNvLryfnUWGFRnlGdIdkL8GmKp+Refuc/jW34wgaPUqC5ZvAY/
UJWH1EKp7B16CJ/RcvvAcIxIe5STgCOKTjTq2gaeUtBCYg7p9wniWhQlW5bE1HfGStrRSIq1hA0d
L1qVEYYoY4bpVhhVXDMRWtllxOyYOaJVIelcpch3Wv5B9qdd3oARoP7j7ATPUsEY34PdDbhfIRIs
F4iC7xUe1Myg/ia4kYbqv5U26dPVN3rX9RLk//0UBdSanv3EbrGSfXSIbETOAOvRvZL0sw9ugMng
Zbu4KxgIQ2NXE3lZFYD/f1HVeOD1aVUrX1CFGgfF2bPaVVBxy8emTK+rj/1i0X/AJ2TmjI8zzwHQ
XlBxwwVuUVVM3h98kxQzrR/dQPsK0yLXl5ymvm7yDdK3m9VvTMaH1321wuXjSw6/1EfqB/c4TkL7
tns1bICOOZznh4zeIBThKdKkuo8SRxjN5JTRKsdRcVPQehWs6DdloSHWgAbTmTnqBjD7rBfWBz3k
eeinM/NrVLSr/TPGbb1HTUIthpDFVcCv4nM72yiChwL2vqrrhmt7JDpjvmWdITsnA4KnUoR9+Ig+
aYc261u93uc6HDXJs9By17UKYRjaggost4eXQnfOcL/Mt3E+9A6f9Ldy3iiKqHLD93C0P8KqHtTG
pXtDkSNK2cHhhKmhQrbr8sbn+FokzEEqq3SmWJO0MXYvmF+42mWoiRmon+KWB3BicoFEtM/4fi09
1ufE9v3u8vmt+gXKhhDL9lSClE1jDCaVbF/F1gMnCQQjAWP2CSiTLzCbJB6Y/hSqusI4TLJpZNCP
o2mLb9zhuVsGiQwCXSRsEpkCyuo+xBiQq6gSSgjKHW65VA4jagmaWzfbF2Nmr+VLB5FATZ6hqzTg
AFHyYSBbGo0VQURogn594rv08VlocFnOODJht5vZBGevJoY8YoCtfR1l3Xm5qBcYt/87nJeU+wlP
ciu21GhLImRaq+gZZrL6SElrYzDE/Hhw6ICmse0S3QxnEJO1Z9e9Lv/jT59xtH4GIhnIKb8WETXI
Ym3swrkkh1Np0idIaZmEhUfrmdTrB4Mp0tBXxduxKy2n5IGlsZEU78svMPzepjgcu8fCKOTLauYA
p3uL5YYrjoOnXcZ7gRLA+PLpOUacytYx59Si5qD0fQwAsc1H2ex/q5ocdQEJ5Oqn1aBvpobsRQim
eIw06Xi8VXRYK+BRK5m/B3ShEXM0P8zDRe260DoO2uDhLkh+x2t8JGyDotK5eb1yfWBW40TVyJek
jPn0cw7Q9dOa9xx6+qpOYvNkvdprZViZgvxeOLYvtqv++dpvgZXOs5gaWCL8aE53MvyLHaETvQ3b
8kmnsPSiRnYSjAx8jkfBmLBu/jrL0wpJMAJE32TZAYn67QDHo11s/tv8LWsDjPS2rmW0tsmnSfIR
CKqmM69tkk8QBdybV5HlbT/DOvVMHW6BBbTwsPp40hvYMq2/oIK+4iuaMgOzZiGsX6iGPjPIV6uA
jGJVzfVr+SGN9HXTIC0odPP3EZVIl8dwiBqnu5SdWjhpiEOnnKNjuKGq2jHc4RYTreJYV9hjzpU8
kEXRy7gdmV/rSqT4pmsjFLz+U20Oy4yxDTR+mOwAHZCDZk5/PQQOiOZ3H6hr/eOdV1af66NH9+19
J7XNPA9IY+7cfzc6u0VabdW2lmJ/JBnvODbPqVn+ic2NrhvgbIFUxn027p+J8sWWZJm/6wHX3uKh
+1pryoQ+bXeQX0gVcWW3nIYWTt4F0oaZLvM3mUxsFEY9D8L/iY6s+gVKsG2Yg2VRoS/JXyTwPyra
xLYEegX6or7mAjB0BEjsMkBIMGZoWt+ZiZIBc1B63NNoEv5UJkYJDWsGXBbhEQ3/93t7v3k0dTWa
b8UIL0eKvGfyMTgUNzVHrnxl/SuVqpz+PWFhEmpG02InlQDNpvVXTUQ+st6so9PwVLePlm7nohyI
m5AEr+RIJk7aD8lQzIjI1RR4TkGCyXlIF7a0R7g9JtUxdFI7XxQFeRoTEuBHUs/sFl5IV2P5o8UH
jLhUnZ2YiCWHvL//KOABlnidELiFMFhGgzfKZbBJGyE9W2Jxb7sViCsJsk6rpxl4mVTsbWyMUSCH
lUV7hNno7mRk3r6WOoLsz20qxJEplZFPysJ2qBrGSI9dOJagu0C0foeyt6KXZVBbhZAjILTb2yK8
9CsuJ74NMpxpWqhVKa88F5yhKPCL+Hgf9GlqHNptvfHRPuT8aTXzCQj1C9S0yQXLzPAjLgrX7pH0
j0uDylra3Y9SxCTgzlriXAEw3HLldkqrqXOlC2ph+Ig5zuifBu2C32qMk+8wN3P1CNRUTcKxkxdj
9YsB8GixNPuWlIpVX6whWPxSOks0GAla7DaTU9QW/kBIVx/wNu0PRA7pYzK09D43xBh1rAxc6e3R
z+XrhfvnF+0p3i94J8OODLaKMDebExKxyEQI++0SkVugTHqxpfenJeJmvw9ukHs+LkLrJrLXwTph
cr/enwlTBNq4X0JFlYWCRi8yKA0YiusSSoE8smOuxMNNMg6Qt0Ngn/JMdfNRo/ACr9X86Sb2G8UH
SDHzTJI9RdSNKMGOqqSPO/awz/nyKO44ONI5X5r1WbfHvR3ZiY8WzTxEaANgQmfH1WpqPp5yvg0u
7mv37sc56XPdzuP+z/RpfRS1yMgaWah1HCf6nDZW61swidJTAlYOFrkY5n+mgUCgf8KCKJWYcQ3I
zd1Dl8PWffXkK10tL/kpg/zbOApqTr1sFdGy0FzJggeUeKLNXA==
`protect end_protected
