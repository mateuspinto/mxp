`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
0USWSUGxovGsyBJteYpEoUUrsfTewzRI1cIPEgOtz6mh+Dsaq4or48CHyq/JeLeCLEYgZuy0Y0ek
+AoVJzSDytI34FwRcarhDByvVu9XjHAoR7gh6Yp70zxQf3NimZbWp+n6t7H39IurXzTLrPMynKmZ
r8CyzYQYn5rIbUVpXIK0quNjPMFJ/MFoMGg09XtRC6sPuVldD2cSMs2++rJkRYAPv61BlvacpZ8a
i1Dfj26gM+0T1CNUz7JUuROa3Vli/jwClVHSlbYhPrj8IFG6s7izlhcqtEmcbDQijjeVUi6KUIAA
twoQcMdJnFIgilS3PHM2JPOLfhks0ZcQyPBRFuX9S11u4p+I/PfVgxp55HwjANb2CH6k4n8VAZ+m
6ZjUra/X/KrN3UddpR9R327/sXP/rdTlHmTEN6CeMJysW9By42yYxyEYvOQlgbsFSCniT64lM0mh
P9lLmwj/VG2jf7t65GPQaBFCCySBDI11LC13FfKhwZI49bXMlQvPReCyi43HoL472T+dQlqgdxZI
a9dSrvkb/J6WPUoDoZrVft4YXH7tNieVxHYbkJkKwmzMR+6aapKL8LR8ufslnswN01E9veiEy6l/
rpI1rIPU/+3h+lMkzyzidw1rPhtHF6Nf941vukLvG4/KBlqy5G4oM55xiNRIuW3Z2NIJteJUtXHl
wS2++yVqW9AwxbmuLy84cTGIY71oorKYznEcfq9M7ISHVvSGxjC1GTnKUbF2n5pJFFueT5zt3L31
OfIaGeO8S+7IRrLarFkZpv422h9y8h+hsrqJUmnjzgBiUGAO9W6cEMja30fVzKe/XkJmR1zYPAnW
nGYUnrRb9Dsk608lYgxm4IsyjQSwIE9rUgOyuORSRA4sJbf0PMvqnGzFiBnx5fFJI7n16+nNc2uD
nsZX0JRR6pM+BDdf1NNw9PblgNiUzMya4qdFzhxUODHDpTR5HGIBj3KZE3T/M/vY1z4kNvL9eC+j
nOP6WKHAlr+NGfZ5JP8uXNllikYmnJ9viegh0jLNkAU5H4q25eTriOgeTkJVhioJbS5IVgrFFHFA
exdZYoT21YWS+1GwLSLhtn7Yvv0zf6L7muFxzKZfQjZ6IbqavD+i22CKlycbqlRaWKFfiqNm/czp
vlMwZJ1Ton/EDZ87UFpaMVnb1A1+FvaGSWgRA0IGkAKz5LOQ1y8df9Om3fDVz7buXlnE3g4KfcZH
ZyXaQ5Lh7MEYXGLqounD/EL4hK63VK7i/s+D3lTSxJFadKvJZKpmOWb5EC43FY0zy0niNsf5dYbN
Hhj86ZIIhjaTmBauxckP7WEz1glSxRRq4hv0B/4e7reLH/BzkxRS0NuP+5T3zDrTcrfxlrDBxe1y
VXuqy2B8xkWiQaWqtDWm/ra4E+E0xtmqOcCDNwK5t8irkW4hodMghJHZ7xJP//ffEFzgQQC8pTrO
Spd9ujlc1dFCV/CzXuHe3U13/RVO1eu6YyuzeHzYP5uVDdg/X1GSNeQltTZUN35mthkHzvwJCnAP
OUu/L042iJ72qCSuAVDDaBUpWfYK9iPs/WOF4H+h6ZFomPXN7jtlLTl+7pbrmxYqEQ8MJgP2h88h
F/4gJIk+lvEnA1kDJgdnBd0Or4f0+ah1jpklmQsa9k3N99WTx8UsCyHqj0vF29Dl8WAeDIV+M7mW
bzHri81bh8R1NtmESbpGQEAItJGXsW/dSCQNu8DEX/XjcduQLqFgnkuiAQ095mVCbcHfkAd//HOZ
ZX89nSqb/OZ0rog8yQq/QTATRnO67wUpOwpOAU5OpWcwj166+l1Sp77zw/SVmu0SWsHpGYDRit3n
t+9A3Ft3CFdAyHfsH4P8nuwE/x6de57tB2IXV+T2oS9yPObnJOSfYU3GKsorcza3ADVYMcQUiN1a
sdpBp+HUEegKsB7im0YYv2G4yDQsXQ3Yc2AhMEKHmCjpQiyQ+EPgZgksP9V6J+Ei1BdkWEZ3u7N3
jqoXZBP+DasDSg+I+6Ttoxs5tDvVzv4pB669VewNA77c9QbJSH6Q7FceRbsEl9H/m1bdcJPMO54v
E4oZ8qelLvyTFLRrmdN0MgBIkV56rzjZ4jQpCl+CDENMyICUQDEWDO61ubnt+jqno5q81scJ0o/i
shLKU7ot4GD0k2k79NzEfcko+bN/AsIgTsPxhBKqdXLHXteF6qBqA6kNTfR6gHSqPmym3eB+PolP
Q2XCcxHsb2XeJQivFpFyz0Vm5xUhiHWbICiR2Rj7WmgQ5tno/pq2gvPwfY8B7ujsuXTW4eGfK9qk
aXSDGvvmutWKBY55RYYr/VldYLdkivQiWssVYda3bMcLLo7JQ4sMwqo2RaqNZh5AsZB+feRcz6fR
k/fcA3HoJrP0zSWkUB1tWjIov4qouzaRMEUc/W3hLn74JdanpAPDmTvh8JDEL2Ntgvjpr+f3aPtj
oLCPhKGWoBpC7agYJAbA4SQOq5u3d//fbP3brm+JgY4MsKjigC2AaezwMySc4gTOpITZUdjIqhyx
5oeHDmBAmu+f9d7DY9uN56jK+kAMVBfAJY5IsWxOJ/3knDRFX3RRB3jao0FYrB7hVb56UXmf7h1A
atsXqLqxCrxG2Q0pHgH/eBqBXqRMk1LBmCRgoyqQAPV0Gyi8GhVpycb8Vvvt0L83oonk0PZWRMwX
9lWzJypJ81/gR7jb/MZyDOSDRMsaPlDbdxsU37vretvjGStksD2l/NX+3QoczW3oSezumzloBVZB
cBXIEfFm0D20EE0Ar5qhNt7LXUsfX1pWfDc0pGsHHbjbxiSJ5X14cKH40m0SSiRFosFk5+DqNgm0
/gDU/A4fEwagHKeWmxETf+rIXZjaD3ltXcutjyq7Zo9oGHTpdlulNKsvDUkVgXo+SwkKaYs6Sqsi
8OPF+Id5Xb26VhwuBnRPT26UdpVMhJKnUZT6Xyx+No17wx1vBpzQphOPminyjf+oYhozCvkKDexg
cMILuXqowPYxZtaG/1vkVzNv7Ju2WsFOM7RaoI+WXxHMCXCQ3oBpU9uXym59G1ZrJM5XtO52T3uj
NdqU4LfnjWH6gmQuLeadpgJJiQ+ac1E/pdXEDa0chMq7tht54kL8TpiOhb19BWTm3BOxaiDXlTcN
sTlYV7ZEeFY97Rdqe42z8P9KUVaTOjnVeXCiA/iTaMQgdGP+VIhSVJXrtOxNFFQ6zALfyOW8yKu9
yTOIzoSDgAuoYIqlZrwjs0QklI+EsPONZwreuSUjReP7lQllJnT3EYlxkT8OH39i3RDdXHo/p7rI
wjNktEksRd9E/0Hy3QBHaxGS4Z6pBHuhmeKLkUPSLRnfaVs1QZnfuHr/X99ozpCmEViyEpGTcW1/
Q1mGZq5FvvHEpnWa+GO+0qEF3TzHV+lCJcz0KWXnBupss9q0+R1hiFbSRYpczC6oCZSyP83ptVPu
zWcc0llGcT1B/q+qozwkDxBw8pMl8GyhjF54ExkRxR2WfcCUnTyFrGGIWUvOOBAHJPbWTVyMBnqo
56262c4/VqLujYWk+MIOvQ7qkHB2HzgDzgfDv4qGKI0VlrXrovHAmSHdsA6fknp+5vjPKf+X4CG9
GO6hOr+VSKVu6NKV5vre+hBOauVzIgNLZztxOshHar3fqu+Zs/HDxgW6X/fzv/gHv3RoOgTY9nfr
jqArwxl2YOqzeC8jAykP7NqTj0Ekx8na6O1TpEkrmOF+EWMKxCYehTcG6jhE2NzKUojzcoIyaTjA
XaxVzpVY/mMpQQJi4t2loqp4vcWEprnr7dpYNR5vt8K45X/kXz+bCt+BncfvdNv9iIuqyhX5kisp
qYlVsgs4YtLx6Lnuo9GDFe7FrzVHjEguC3zpJ/bEx3ihTXz2FjlGbvtd8LVsCqAdmMX3QNFNN3kO
WA7Vsx6nr0ZDUQPEO5EOqccm6+WhfoaafosUeFRkLC9QuE0TQ5GANereT5kFL6dzFBJ4HybJODl9
rGN4lUdd5iChUnI4fTyTxgXJAjFGuGtuRquwPnbPzJ/rmtKN6PAzcrX6cky/h3K46cG5Az2IEXmJ
9Kqq0Gg+PudwmrjgCnPFcBlK7BhyNUHc28xVAPmYiRPSyleMcxDC4hyIOI5wfH6RWCej3YxUNYGV
yqYLuOC8bpdPJrULg3o05k9cEwA8zZomVDHdvClOaem3ZM6dFG3d6BYND4maX20cIdvYx0sRMRnw
2Z+EGrY2D0mGnjsu/fjuARkMuUPavViAkxGgcaQUQe86Um+YMl6/+XWx3z8XoXZ2Q4FDQRhf/2I/
j03Z21keixbSc+/1vOFNtPtHp51wD9HRGESjEVFMXfE4MUZRnQbz916B3lmyPelFb2vnXoU8Rc5e
Vyb2Gf4xnMNKTKuQkzJbnOaaSg7Xh6bdl67ItZHBUmEbWgxedPUtZOeswdUrRrKLNBOOukgdMkE2
bmQ6MpQlWjraIUpGevqDOWdSABGlFmZMjJQHaJX/h4zGCy6JJVaPZyEgpsqFE5PwAA2mrkVR78SU
1UdrRYkUkZBhQbOsoIOtYcCCOm5OG/Xp5z80JlMAP6WnKlvTnJQ7XwQAaahs7O1vAFaE8P+q5lLs
dCxIml6Y254gPmmIAqYB0DzomfouB5b0pGmlo2CVBPSxeU4yzMVSqJp5comeit57IVQ5dBgdjmgZ
SJMOKCl+pcEtMvAns4LfduEDqVGEB50T6w/0S6EBU9bcvpHYbxI6tiyWYmqqD1sXggrL4XiL900H
EFUUuTlZQFnl4hwB+inebdrV4z54Z5pJnGvU+8QHtN3q7yTk7kpl2wO6+5CNLeZCZ0OUrfICJpgp
1sdSrLq7CPUp8YrwklZZ5Xq7c6Jna+o2DeMsG3dmiF6SuS/0tvAoKPir32aAzTbr1Q6p3YmPcA7K
SWErLghAkYqxny/u9rCnp3lXTwrQdZPkNA4kGJEFroO/gP9bwxmEXAeRLgSEz6aiM3RtSGgeCDvm
RX7FKRl58DU+VSDx2TkbZKRbXtJMSdSJx7F5SQhjDTUSCfnOHlFL1ajOB549IxiLskzyX/zxUn4+
/VhkqFHYeqCWbRud3ElOtK5mge+CsYdheKSC4YQTANvPtW0esWzfRi56B10nw6A6nR48Y5qR0nrm
hPi84IDF6O1hLAZ2wkjhoou1jgBGm1K0y+PZ0zBbe/HxJhxEPGw+JqHx1XRRF4JaOxrJI/qQwbAe
dqg4zOv+17tgYAo1TOvi7UcPuEE40vM30jo5vMHVQago0vzed0oHFkQcNV528Cxk+Du3wIrrw3bZ
PIAaDkBsn6unuRddNIJdIxw6SHDXBsxXcRfB16GqKYJGCQf6xvzHLBQlogtu7BapjgbXqzmsTja/
iANezDqLbfXUb0BvO2uDs9EQCPSpl5EVblJHZQrHEbQhtkXb88zI6S/YeLOUkaqDcO8ymaZ+yy6B
D+uv88Q87yCw7ZOOGw5EaUKDx3TumXx58GMy9fgVrsEKsvwa/kCHwjNmD9if5Ci0KcvZAdW/3uP+
hQb4+FHtm6TufFhIWLqVwo2czyCIZbW1PiWOIh1/3LAXrUjQLbFLyXbBKZLjDPH0A4KvcvBfq025
IcV/ww6R5pNZyAtqPcjWbURfpE8JiSgudgUmILc5ejRpCGnGQsEO7rxuTpRF3pFr/npgoukIJtkQ
dlAHX4bteBXXO6TaB48E6B+rgo14TKPcOQdLa/1Q5xLl1fae7UVaueY0zvBGosdlOF1RnSrhVeZB
3JkW+isk85rLPqhbEZvbpQf491DaGjoySgYXxdVcKSjl/VKm3ZDd4QqkEvHHNqLuOC7tHiz4myYa
ECl9rilM2IBxrbKIVZIBGDyxB7xVRpg0OotBynq3rOE5AUf1SUCNFCfstz8b/SdVU4/7gP9Mqk8o
uUbVRbCfu6nqyEuogwrt616UQZ0qQ0K5YFX3vs0KPr+IOlq/xHxS8JPNuOSL28AXbikdcZAv1Gok
L87sYnofGwj1hhG7zwtRnmichnkyobds4gbXE7y1aQonEkF3eOioyLaUVn8Y794GWnTjg72wJ9nk
i91uuwvy+/15VjCKRXNq01eaumIpw4mk+8IbtdRYxKFQL8KLjfoQ7z6IVdXqjiCq6iAOsLH+qBtZ
SCxOyqCcp4a+ZFGhy4MjMLvGmqIoUKddeIqeqPpAVw6RIF6hp1bxBGpnwqW+RDDNjaqxHtD6a29s
lfVxTSh3svucXOgKRccfPlbjTKMtpcQtaY3SdjO7lAceeAAGN/FG8UCD9Nqi1IxTQLPZ44uvQAWe
Dy5fiPir2F6rMzMnSimpkrOOXPuoU0UodLQkrEFGFNP8IveBtf6P5iDY7LrfwQFrWekRpPymV1KW
Yn3DNg8B0D8KbeToI+XtFxMwPqvWEEamMvNQAAPklrj9m+5dv30araokHDtBEc4fFgCaEVk0+p5C
2nfKvz9sTBVmruvu0Vf0Bzz8swkGf36an8pVyxn2YCWDmliMsx6TQ4on5xzSU2ESGaCnEAt1DfW5
l38yWtXBlb23yVntG8Vrbeb7LGLDRIRMiyZ55NXCXpkBlIkmi6zGLT9odOEKm5FGL2OokAabnCol
+2IOXefrT0H+HDg/by1vEL2sl7g8dPoW8Zu8SJlzKKCwftSD2OfD/54WuIahKRL6feMLYu77UYcE
f3wHdFJdrZ2rE0AE500t7c/EOQh0Opfo3m2/jXjzkOqXsPLvA8p8+SYzzTjzIR3hNopzFCWAe+W6
tf5CAacfDfBaZ+tTNaKvHgkzG4Usnzn4spL7DNQslKUyrtiS/NhiO6CQgldbYqOQXTOilnoRDWvB
ioXbXB+FVY4aoh60abXJyFZPNMD7TPSCTECR5truCsRbN3RANZQfZepe/+4aTvvdJqdao9u8fpL+
JYiIKgoovIBfLdBeA/8TZhvvNw5P30pU8BSZ7dDlLdXes7KE8paCLBnucWcjOft/3+2brFSxZJJ0
LNoYdduQP+A8N9N1tSh8YUcXfidktZttqf1+IBiM1BPhWx/Y0rmU6lPetOGxQsrFTFiM3mGCRU3z
ibC0Bx+Yk9GwckSLKgLayrNfaJSoCuBAUI/ytsFtMYxXs6e5kRD0NH26o0Yw4mF+Ij8wFaZGormC
2jPmuiSPHmQ7+POyL66aKssXGgkzyI7mhzzIIVpUyvCM2nvEHY6/X3yLjLs1Nvk8vTGh11Lj33+t
Xosa+pin5gQpBwQpk1sq6dDzzb5YgQ5Dl6fEqrSA4AlfxUXrQW7buwhKk9vrtpb/F1O6WhRyIjnw
n9vwzJH3Pq/dUtHCcL4LWNLuDjOfRTLAp2xtOd+LNgHm56YMB3/+CVMO9SLB9EtNbjPJDSCJyM/I
OQI6TK0lMLbGXjKV7PfWDZT9Lnq/oI/JO36Z+BAkXk/Md9YaGcb7rpdDu4zD108HYxK1C3JPQOoy
/Fh2zWyH8Uw8nuylUmqUQEmegrM/C8WhnTXjaBophcWY+ZTSS16LALFXm0b79lNcx86m02D8MVF8
+1Wj0xoa1y+janRbRVGomJU7v5S6SvaP0xwCfn9KLmZPJ/lv2+4/Erbyv2+wHOhAtijSIu+lKgMc
dUHhPSQq1kljBAylyUIpjts0QmtcdO6lrw/XznQ++eldZ5A2lrKF3qeeWdGNpHbQ61JbTQA+pQ+4
MTIKuMZeSlNPbs0haJC+Sc/WxD0ubBEsZw3R7bMjYkI9saEfk5/KLnOqBkctS0jXgnWptTA+BnfA
fmX+p2LmSoaK/c0jTvcALJn0nd0m5lqVEb6qptPz+/T9E+LtmrLn248Qe8ROvc+RrwvNa4raKBfG
Tph2v3mBNqG86wW2brDgle5VdLbKT038Uz62DHIVn/k1j9hdDIaW/kvrqX9kO/ltfTki6NSAFWt7
sXV/Ql/CblVRWXVRa12r39JYrnSs5onHQv4Uto3rbUrKT7daUGMjuaQb2QhfRdMzNMKVXb4KdBZs
SAEIvH7v5TNbp1pOCG2W4ystcrL5kBF18sH67LVvm7H4eNsyZGfXtfHvoURH19PLb/SeSWny59S6
W8WqhTrGxVxxD49YdboJCFUV2dHTfn8qGqhBZdUXDzHCGbFcZThGD6SxiKAe+5FHwTePAPbJmIJm
ky3KT0dXEoXaQta4QiGUhcmtZwc88p8oknHBHhrRYEAv4aObTCrTC++Ux8ypT0CJ9JtLTUrFeTR1
eZz4NbsFjODGFDPZO4z9toEsm3B07ljdONxlAxRuOh7k3vbiwaMW4gy4B166d5sdmDw/LJ9+ms3t
zGcH+jM6KZrew14B28Avd2JoKXRa7rdurKxHdmWfwkrUC0JRjt0v9nP3Z6UtHhdQ0JZwqlthv+nV
P6lwImrH8xx3u5h2kmV7J6oodTiC5zla/yOrVh4ZmA+ZzbXvgM7J+gzWykWdM9NCqj2b0HqhVt5+
ClF4SaOgVioICIoUxmVnR/eHIP1ITfPmXqh5iC1Gocw3gtzsa9ePGWUePb5c9e8X1bdGUcT98Y4H
RQt9InZeJiwPOSuPEzqY1IMGQfJpkzaFEtoWNiAsrzBdvAwY5An2X0TF70bevdUyGwEubXfkPRuG
vqNv67ZJ77mcxiiRBrmk2OsiMKLOQn4t9hdho8Hb08YWwfKDxP5aZySB3W6dNtDR6/RqGRs5JjP1
Cq6BtiRYiQR/D3w0t0/T3mvVKHJgs/h6r0TwbkAdZ6JV1N4qNDNbhRIQS6qm3JjWzeQ0sRXSnnYj
AAFUnlpRHBO+9MpDJYHWRMCLz7IsMJHgsKpYILPgWOrR6SMopsGZ04qNo6F2HGScde9Z7xsjUsqS
ta8Jcl7Wv4zZFCASbJj/1J1HhzLReC10rMjosKvPYiXeLPIn1pmPiQM1ESdnt8sKCYK6u/ST2+1e
eCPJVj0zxwTI2wZ0KZAp6R7XL85bEGTAdAA4zxEdLM9NaAFbwVwg0MrimUtplmJvzlQR7ENWhjEU
sFsHxzwRryXwZPNUzq/6K1ouS6xVfi2JrNL7yzgqp3B8i1uhuwR9zAGIcd6BNBHueuLAj//rCuh2
3CGC6hlKmoVsVmQTUy9GqNdgemC4mA5K0BS0+4wk8r6c1avOsshB0gWFiBBE2uTRVMYKVwzdBTmU
YisZdKWNxDowMhqB6ig0NVZZ8hjHbDABp5NLqkVRZ2UuJZD6dhDdfmY7jgiS1bPKW95JdwF/FTP4
8dwKwBPt64KQ5MZBzBa93X9Xvqcd1XcTV3TMPtrxuebAXEgxRhqrdvcOWI1pZE1UQfpyf9zsQJEE
msKPjCayU430hpyRlzN0c4msAnbQjLTmJtp7nTQpsOcp2SyHctAD/jEtpOXmegMNJwqeE0juktPi
3cXwh/UruZZhV9Rv/6lZhjM/NW+XIU9jQKcU1w8ui+5wv4YIJMxeyK6N4XDBTDhmK1vl0w+Xhew6
2CWEE7Gu3KNCXQrCT6ePsP6oAr1ILznOn+uP0OZ02lKtX18OxlC9pVCdUMPIr6+azFwLgiEEETh5
rcMxAP8M2PYvW90ZzFtcZF6USTSwx4c2qQOJV/TtRmfOv25aE4l7XD7NrUNfSS0S6HTiSxCNXp/z
DBS8bzTcNlO6+GVqad2gOHMUtsnPtYu8V9uEUbsJvQ/Lv1q7TJ0n/suftxyI9H0YM1ChpqBiJF8m
WJhe2ujOIeLuJWI9ehqLMK609DSTUQwbxjVTWNQvHwD13qe2pSfEEas1LfLi+SOmTuAgSQBGfN2H
dSPk1ZAm47pPWG1KTt+xKsqHEo+TW9AtrwSYUA4BCBnT8leWKymdTYFCc7GODbh8TyBwlZItcaw2
tJHcIZTslW0vHpn8WVtJSO1QNK5PMhkN1rKs/DGlo4ohwRr613jA6AlzukGED2kdXRgKdu7dduqB
zuL1FaCdR+ROJ6K6yYT14vxswqHs72XPnNdBdmRTdIXzPx2eMLU4OpkqxjCK8uOwa/gsTj3DzvXg
1gT1Wthr+x46rrrZ2J7SM8NTXMrlV5mlYh96Jn895mfI5WgX6Jl3kZFY9mzL7SpUCHE7M1wlArqE
vCSFtDOrPAhCcPIvxv6iJY93DBOH4wSRRhw6XBYcwiqRkfjxla81kddyTPpcOPqgWQjXtPzx9qga
YZQCd8pnhfJWQwBDiL5/OPbbRlehkhry8SN0QCCogTJydkEyWFjWrgswTmebl3maF3alqZQf30/O
7PfDgT6KUcNpe/UQAIXei9b5ZKgX6tgy/Au8LQQ7Q23uX8TgQ2gD/Qz1C5Khfd0Ju2elU8SLfULL
V0FcxLuix9fNi1z2LUjdw3i3cIca6B2TZ7k8Xj3N1O6AHvZx+7s6ALxFaqsHkNC14rYBOai1OjeE
Redm0za0RkKXdsUAJgz4WuHkHt3xjnE9E0+abayJo68THbpPzQc5CZrrmKy2Ygl/rON0sa8noWc8
qdK6R20ZbNcpTpg4ghZK9g26r1sjLtykGzFs8eyOJmwPNz5SUGXFZA3UtiY2uiDr0D6TDaTAHIr6
dsYrYcUkg6oMVrsyOIO3cOXY3reTLU7Olne1RaYKs/eQ2whdok1GwkyAPu+DtyaqbeKkKbUeB72U
oqVxdnUgHR3/zqwc9dYyKiLfMeDq1lcXPrDnm4UiqfdnOlwf23IvzqiVZsyRTuBIFA+tnYQ+OqN/
VVx5yxZECRgSboQawIh/pVgZJ6joAeOUm3TCoJze61P9soRPegGI6vrhoLm7vnaPc1iz1aq9PlYe
snlkgp4i+JGzPfYwIVhjdU6T7WG7udBKJBv+XB+qQaDG6aaPf1FJNxkEgQyS5K13rCUZMgy+fWJa
mmxhXPz3C1rsVOgPHRQMW3m97UPviGzIT2izSFARNk9V3ASslmKqwfyyOOgQebO2GVVar5AxqRG5
dTdYu+3ydb4+BeTog6Eh9KNjVU7dOpB1m79DmL0JbNUpiR1NmojZwom5TRkLqwtN2jXc9YwE/Eoq
m7jcW2kxtKPCfRmNuTafZRd2URfmR2JgiQ8h5JwgF3dy2V9uBEstk57oFbvhMFBcdv61UfwRLHPv
JSKfKWJ60NyRmL8HT6Q7TAzrkF9tDjKeyUdfcgfkS0UOPCCZI5D8UoU7Qia3u0oZn67aChhpn/EF
msDzSrCh68DUT0bE5qK41qDCxXX3r0/OGZrRRCGiscDLrZqD0V59JXc2DKHpNtuFJsa0tbzUVlOi
wrW3wkqL/DD+6DZbm3r19kKwEsNEFsF3RZkxP46n/gqxotlaekJDnKQuU2+WUA7E5+BsdBJnGPA1
aLP8qUj1IWVtYaKd8rI5jjtpIpV0XHWmxRM9Nq2aZ2CYc5LiPXDdGE7ENoL2a54f2G2NzJWHSfwC
7GOa4calf/ta3Q+KhCnCHJhBkEisJvmjXRkq3gntLYpJKdpnzsGp3RwmvZoewxCoOrpwl0nhnhjp
Cll/mYxxWBNc00e5RK5ZFwcpOMNRfnQ7MbuvpusQM+b0qLRqcEwQ7smbVK8mva1MJJetlUrk8tt5
ZqbKLsF6A6ULrSpV56t8WdH4ypb8SdrzyzFI/VTqxADHu/Kw5l1Kl7THYAaSkOoPtgGZRb82aEup
owN9aIHoPWqeXgZkqgcnfkJ2WmgjwkcTDzL8oekxihACGv7l7QDrXqebfC62cCzBna8CxjwLPa7p
8J57p4zFYOOAo7y5xB5aZNytpb3aa7lxO4ga17MY4Vc8Ee3DIpWddReF1h2f0ecwR0QQ7HJ4KUgy
070/XzLob3tN0xbK/+Dd3bDopTulSZY33J1uiL8qV5tCLmlsBVCsCgVsw1yi1P8/JSdHsxj55P48
AGRSjAccz93PJGsUGVqCoP21e3GgW/T5kDd6fWd53EzZclmGd/7YXh3xSErf8wFj3qewBTr1oWo0
+PRGGye4OZts7GubRzOfnSPBlWW2OYQEJbgRyANAqUguEeOdZf5mHiGqSOFfAxG9Qy+kOmptnFyt
0JCWnj3oNxwudlHwHFi7JbBakOBmEngmdSokA6lgkP+wPj6i6gXDF+7bJi8A68PPbRH6hhIXAR1j
oio1J89doaHuCpfWhBuLAhLcQF5euSzHZD5+yfM8gj6xhmUAMjia2SJzhW+4JUNIHCIvP3jjhiGk
Cf1KORxuRWDmKqCZbp8/Uc7+rpgx+w53dP6JnUAIjWLSGvn2uyF+n6Jx7/KJ21ZvC46PpQXGjmYU
zOzrmMPPE/QBJuwX9PbD+Qb48ogE9Ts0Bw56zjCRwvv8jy8QQqIO2cl05OLJ4ueKde00xfMItCwW
8EbfVuWAVWRuhqJM3OhjH+Tw0sv6VIvVRQtCGpnMGKqt9SS4lZxyPxs1g7jVxt6XnoOZPRwfL3Oa
IPv5GPvK1QW9UuafrYYeE9K3fn1DaqIZMwk0HhGqfjW7ccaOyYhNVbdR9yaEo1cDQ0StwzOaerY7
Arpcl/99cUOaCUj/U+a6mR5x/brSeEUKc4TDBN03afoLMrsNNTX1wCU3xZezFGU4WUlOl6eberYa
ulVd2HZaPgq77icM/5qozwgUcf7KdIR9LojTaxOr6m0JF77mxslY0zXyQAYvcRat7mdKIMDM0O+2
sS1e+chhEYPLZglRdCceriTh2nOORprjdH0arCPrFpSRm4GoiDPV9vO+8K1XEbcdibHqMJYRxu0p
OBoTQxjIQTNU+pYp3yHjNQc564APojItJ16UhmfGZ2SF4HGyyp6Bk9+b0w4sAab0qFeONHfzSPDp
zjBaG0pMv8lqLzRyhqAHpVdCXxn5owL6LQOpjPQcIDAjj9F4CK+HfOj6DonAXt0Cvhy7otKCHPWr
QLydWKI4g/6/OekcISqc+2UNccZKl+wbUGDJkOp96ZvljIS5gZOMs+AA/vPYqC6JRY3sKJaXH4Ye
+akUwh5CqilOwVdmExVmWALXw3FpvosGsvamDBzYQDS+0wG38swpKekXJLhPc6sAgoV5l0mZRYg1
lRX6C4hLo/hEBNoSFYZeTzmTg1qjotS/NH6ALZgJQNjTwATxmbwWlYanhD9lfxeMgZODwT/MmJ/n
xR3fLC6Zqt9xXcz55U6xPUPU90QWVec0vW05QdELV1gJmcfb5K6lzs2GoiX3PI6QZL47gs7dBlEz
i7c8XVUGbZLbScgmdA/SUHPfbl463xK/Kf9sla+U33lNBD6FjGGPPanHs2TAhSP+N15K/1J0MmKo
l+BJ8C8mikIiZRbyv36PsN2lMrBJYqQrlryaoMl4VBUmM+LgdljcA1MBXtDi5fpFx57GDSZt5HQM
gbcgztfk/+XQFVQCdBe/Il3QqHbWHEuyzeM7exRSu0ruKSSM7rnbuu5n46iUHPyaeHfQ1Dqt7lqH
afKAmEJxbyGloOEbM/T+R4KgUBIRtFr6uPAZ5NIC4NJwcHW3+M3XKw/wOgplrqf+6wUEIcBQgWgL
hC1JaolkGTqZMtq3TLBXvD9eDVQ1uVAv7w==
`protect end_protected
