XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�ho�x9�� ���#2,~d*���t��\c���ᏫB�k�݊�Ή�'�އIYQ`��\��xX`�#Q�@�z�5j�?Ūn��$s؄�e`�N�
8�	��c%	��uk~w��g2����N��B߂6I١dV

�&�qY�s�R?�h[n3���SU#(�A�t�?�Hc�@`̽��Nu�k�&�e�m�eE�]���ou��/��&��O2��˼���B�����@��ۖԯ0وwɎ��{��kP��$���Y��p�w���%�
�wcb�hǦ,�����}T2�D����;q����̟���K� �<���H��{Ƞ�����	�wn6����\:�R���a��l�����a*���j�؋6$��2ȇuz��18��InG\o�w�9���=�I�x�r��(����ۻ�����1�[~Jq#z�������@�߻j�O-��x �Y;$�zI:�/!T��=�~ ma�0a1DOhtgK�S&`�)uA�(@��6���6��md�l5�, !p�+b��yNmoO$�4G^d��ՙ����gf'H-�;"��K��kR�Xd�m0+l�	�I�W_�W���-g��ѻ�F~�c�d)u�E�IVeG�xO\�I�Q��"B]k��	L|���7�-��Uк�cӽ�����k7l1��ВY�3����\�2��wE`����&?B�������dn3Rk��=&�>�v����J�nz4��2����D�p���/XlxVHYEB     400     1b0̵L�E�dkA�w�5t�U�Q�_�	�s���/~#<Z(Ϫ��+��R��ZVo�}��I��mm:ph��R#Q~G``���A�t�&8z�fmZ��0T���D��� )���ԨT��Г�Fp��\� ����/�%�5i�Iե#P�P|N]a����<��j&�M�� �&�т�c�o�y���a�/�5�us��F��H�x�Ѵ�nCcN��N���~ƞH�Þ�1��CNb��j�r�q��Έ��ᒝ}u%�O��Jd������v��G�-]43S!��.&��ѩ�e%%P����"".����^��Q�vՙ������o��ʾ��Um�H�J}P ے�64&}����*Q[�f���c������ҟ�	Yv%�i.��Y)	��˯���A���y�N%O�k�7����rP��6���x�=XlxVHYEB     400     170c�o���g+�t�ūp����{=�+Vg�ZL}��_j J�/w���ѭ3l���.��qqd P���q�_~�~�^(�N:l�V��EV�^���aO%F��;*���0?��]�m(HA+Ztox��꩷-w�馞���>%��B������`���A�u�|���&��9m�>o��q���o�O��J��%]��Mp�/�~৾�T�e!uOSO��󹲺��ߪ��Y��]/\���.�3����܊��a�S����� �D��G$�����DQ�܌J�b�\�ܪ��2���~��p�;m�6�)�I,��,��G���b���Vɋ����!����λH�y�x+q^BXlxVHYEB     17b      f0���ؚ�JD�d{���ۋ]A�ٙ{�}Í�����������2���T��ox�'���E�����Q	��=�]��'=P�ȦS~L�n�����AC�:�pJ2afQ��&E��/y$OU�q��"�g���m��.�>�H;�:�=_(�p���\�
�fG�'Yl\*���dir�^|��d�"�����d������5F\*s�q	�50��$`LۉC/Ҝʒao�պx��X