`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7216)
`protect data_block
0USWSUGxovGsyBJteYpEobrh82QgPo/7UxyqmAdCBDCXQ+/vaeINhHXnCCt+8gFawS87S22qnj5L
IZ7rbkXK2b13WuY3/1oJT1pU6A4YNVvvERKxzlf+cspYPYfUgLmWI4GMJhOvYGhk39uc0b68u+kc
pJww20kblDoplYeDxg/o7/wm8b4tmmZm3pAI7n2aViW8NEZygUQojTAmvQiVMihjKTWip0qROdNC
+i7qNAjBIfmA7AbzwqwF33ReNetJJt4lqLNCkjF2jltwD9bImz62DB90YOt9lhNiXoekuk5TLQ2d
uC1s49GTuz76gQe1a7R8qwW+M1mAxSGbeciQ7//qGEWYR4his0qrU2GnNYsD4ycYmURBQjZ/BP4l
qx0niKS6fuziHzT7ryGsBU7H6+geU58GxH6bQLYkExU5Ny1zFU7nVrNKeACenTq8k+aif02XGQse
2bTOLic/EPvWY4kitivMEs1Tc4jb7zrMBucOGEVLUIAklo8s1PCZq8hxyS3azGHeTBZ8M0oORvib
Aq2Sk/Gayu5SSd5uBsHMv3d/hyqh6ZWLnv83tX0VhbzWabrWnNXpKUBwNWCuQFT6Bc9r36OXxiGl
HTA2j19jKWbYDgyOxjEsE1zwoyIoFyV1DSKcl5KdUvVNGwI1EcnvG/SZx1l6G2CuCw9pF0Lan99a
V+cNzSernogrzRPBW1m/Fj+73iilsSXgx73+w+o4f55Vn8vBdldCeSwfYRdW3xbbzVRpZgFh7wBq
euA7evXiaVz6bZwjp7BI+siRIibwpoqRjXAbgPTGxVWBdCKuumPHCQrGUejl8osWC8QgvwU0aBYu
OGFbjWFubL2YL5yk29Zy86BKm4nSpO9utOW5jUMBL/BqMG/HJe9muakA81JhKWEI2JdbpXoGngur
Vvic/khxkNl4Q5aX1eqqEcOi9/PopPqtAQuqFK1NucrB/rzxZm7WA9zEgdNerRthxyK3uKUu50aW
zbE5rckbKswM0pvf0QvXHia8K9vguPXtXitJNs4hGQyALwq2zYUrhIsAEjuwuaqe7hZoqQG/9TDR
se4UfzKAgCakX1gZS6m0zS+rtlSoJXxNUpEnhwmkpaGGBbkywW15uNAqRaCBs3wuTSlkBiZS97sI
6UxFfuP2cwGmWKueniJ0zi05d27jJBQ1uy5k32eIUucIVUwuRvIj/KnLZIJuVjQ7v4fu86xr0l/7
1vdh8fF4qQYOzLrNmGaA7xTywSIlRfRgNGemlEpXV2AAcNkuQGg+PlbaMfGqa0ujwFn+ut2Hb6ou
7ysyhThmr+CrprSIQHShzNGq8d7WVeLfvhlkz9S+KCcni50aaAa9nkJoasvCS1Pfu3v17Z+UVIvl
PPXYN/uHGQY2BA3VHVz7lnP2r3TpaPifImD2vcWdz7iICGDPLcE/Mg33VJ9cl2dkkEKc0tBisLt+
ysHIqC+hHLaJDy+Pisp1wtnL3HpPuMq62j5uLkEQF39A9aHftNPBtUwWthUejA4DyqwdNFsxFxPw
zebH9cr1PzcYv7WPnGbbg47YU+lA+V3DzgJxKVlnfYVAYZB+Z0+IXmQ5jlriVduFvRhjSMFpTxI5
sGVoFp7Q1i42I+6WzH+LJ/n/GBMM5HIsmXNJK+JGAjnWKXmRLt9iRinIguMLsKnnjqelDeh+ZWNz
RveCTVXv2Cyom410s8wZxH1alFvfZBQOSdi1ef+tr1NLna1D70vJiiHERWjYvKyxvNYNZddjjMJ0
6Qi+n3O47DoGmOoTMNM4WmURQc0RIgMbWQnm0GSBBltabJjHEfJOWRCzRAnvZ4+S8J8Ykz95v/hE
5h7xvUx86FhRy9ZXCA6IiVDYg4VNoP/Ehrsp4xI/FS/f2F1UfcXbSXNtAZnwu85uLYsBvUIdJopW
9BYF2FImVJ1LkAsThHNOqLq0lSiay1U53uGkm+3pdSylUgGdUM+PkmR63u2P0m2+V76186oPqE44
5hIXjjbmPEWJn5aNTo6F81BIQxSaV5FAPlAHDHpjJGIr7O0mJiWMYUXV520A5XHtjqa7p+xuQCAL
bKq8Fmuvy4UH3nqJqqSV5psWpoEr3CwO1cRWbfn2+viURt6HOQjYelva652knDqEqgiqqn0AMFlr
QeT8WxB7rYWySTAv8fMcAJxR+mjWK5Qpxm+pH8SBTvEQGzYKhHXqKA1wxXDNHTDSQXAFi+df8YbT
izNI9sBoIt4/6uMamIJExhXrLI9B/hp/0hR0bob736Jl61pQ05YPkEoJqDLDamzM0qRmPIDd4tS8
er+jpi+hXRA+rBcZ97nX5gxmZzteZ6hUiTwQpnMy+tCeARxEwfhkAGX+aETW+kRwAYCPFWwj7cyj
rwC/g1aeYeey5j+c/ihMF8ftUvYlpo9HwCOOTH9myA3TM8qCFa5y3O+VRVBTEzxZFEp0T3iGbd2l
mNjsasLlt8f8Z+2wQcpJ/d6sl2Ugjdl0F/v9GFdqrytlC06eoEwv9Gfuj1JioWPtZ8HmR3cuzsFL
5bXnTlxdiw0GwRlgqUM7UjwCN7ZwVAAF2u9QnhJE3qexrhSdge8h1GRnTwNdR3FgrSKSHBcMYRSc
2LM++BhkcZNBKsE9HB18pheRrgAoQUHwRw6PdU093zpG8tsyVoy0r4p0RrlDqzkRVMegSrU54ivk
c7994OLOd7kaHPcfEwa/SPDA9/f0P2ynMAs9XmKP2jp3rAtFEqCMm/qcNnYG02CCStjv3KIcZCWb
r4mT6GCZbI2J9GvhMTq/2fHELt0rEEhwrcnTBmvWwbwP8aA+1KcF8dFsNriSN9vuauYKmMtDPFEB
2aDOgJqhkeNA0VhQhYT6FHaSAkyKRdgdsP7eSEdyhQtEajSnpuBu5njQG/rd/dwYsr3f8FvVBLXk
+UaPgod4ReT9OOLBW0okZTZ0u7Mn80uXOhgxYJvJdLO+zighX5NKqUu7w5AaPFqss+M0pfB7/HOs
YaC2kiVGHtIU8BYvU0so4XKSS7l61gsyKdFVG4b2yzO6icZ0J3aUjOMcz0ZfQXZ6FyXadvdPSASo
wKPooLtQceIYyKEa6svMi29xJh8cxdkyCJfyUAhRc44+CabE5TWMThLkp70a3JsHg7o3MPdUIoKl
ZzTxYda5SxLbSNYfVc4assnODNgOuaqecF2QxqNC+2dDSTEiUomvZFPf8nH2ZTQrK5IcDsC1due2
Bfc234f6DJpP2bV7TlGgaepaFdX4oiLwYANEhhM47oCxe7LmV+ix2CScFJIk6JoEqS0C7boM4Nq3
BNgf19tc5FgyHbdsalQDn2tRsdKHpqIrsLAar6k/q4FRFQbScRudrQnLB5IiilclXxqFIcUFcrGN
7i6K/hVD7ablS3dIDwtJhAZDp2Fzcq66htaw2fMTblmF2GgvQOmU8S7kUUULOTQU5xKNvGlipBZ9
ZwlK3iPQstLy6QmW7TD0P8JrMD0UhLAIEFbvoEvT106xrD2gnROWdWh82ZGPMrcGPe0Inx0BTTbd
LR78SnIji97P0jMufPievyMd1O0aI1zO4mIhDD9qG3E08CQpbXSDt6/WjTkxBsgg9Fx/1CzqGScR
9nNQnoQCyY7+5XOD7gDqx0TW0sb0Cm+t9Utw7X7Hycz5dyrg3eDp3aKHoSJ/coU+K1so1YrNPklx
BK66vQxpFp/n7qkbaXxEpa3nXo7Gk7LOAkkq8yyA/FdCbaDlfTztm7ossFvjsPhl1+vOUI0R9E21
aIO9o8fP+Ce/mrpqqvlnN6VI/87WLILQJB/OYz3jZ1Xra3hrEzdhPBKWmRsaw3Sf4n/gc+AapvuI
v9Tg6PWRR1Wzt36xuWhuW7q0j4cLh6bfM3OZwuq+tfSf4fIQ4Yv3Ni/PsjbPGQp4eDGg0jZydkff
KFyxXcggm8mKYY39jLpYoK3UYfkrnlhA/pxw2t0nptRQX6OhZNEBYWEWo7hIaN6UCUyl8YnIbJCP
txp8+bmgPApJELUUlzz+oFY7vPkB81gZqX4hP3x163rX8Bpkj8LkwDgmtDdF+rPlmGqjiiQhdLFg
lMPmqEiNqZCUe3gZIND8bmpCMztjSCQ+bsshWVB3/oSrUreZrIhSA9OtC2m0YiZR3tlY1JEkLdI8
qGzDw201eOt5G+wRmbmxZC99Mix+CikdHmuaTvnPc3hnuNxOZGrXFTPflDoO1wX3Be7peVDU8v4O
n+GdP6xTsiub+EyKvpZWeBdSmombCjnQVw3y1qRlZUFwy0O3Wlhyud7M3DjW0z+FnJSSsg/rG8qH
XkM8KWpP3+PxFg8k0/GI4VhCu56XV/d64pHsdg+GVmGKTivocg8bIilxz+6nCvZO2hOmK/i3xqaH
/7G4kz9TaWDoXTxzjZNRT5TfsMe3jT13RXkcTmE5XU84q30VvSPYubtrL66ATPNC1oEAUkkaH18K
S9wc17poW0pMMox1jTIRBNuQdCYrLNP+obd9xh1W5xoAqtUOCJjdDkepk06sRupExaNn+kAaX5yI
3EGIaPEsWWbwlF0pTshI92o4mHXARR8deZXw3g1Br5iRBz0zNDEvvordsiyt5Axm5ja6bKU7sAqq
02i2SPAtrNIas1VPXyoL+fEx9jO3bxkthXz1xJ6GC3KvIjnBTDlDBcRzpRHqOY5ectlZYfHrZHN9
eNjeYNpafJK8Z/EBtP8P3DJwcwajy+A2PybLgI6vInUcyeqHvDCjYMSGUMdbT48ZtrB92bgXle/Y
YqVZnnNsL1Ya6yrt1HoS+hmeS/iRrxoCF3K48+tlAP3DvySgkpPjvVvDyLI66lmOuo36Qw6IwIQo
8e0qSB74xOXD8hORt3VlgMrQDNa7BxaDPPcAzTzfbTzAJitVEc7WxVZ0ZvXU8AXoxgHfStBstbem
y8k1hVsXf0M3J653RcmqFayurzQtCBGi4P2PBuyRy428LWoQSTJXr6kslWeMf1DqaZoouh18cBll
UZ1kE2B5GTEUWScVX19BovSVK44sCL8MS+lzYLhSlPHacPYxCLVJBhuIVYFErI1epHf4NT5YYlUT
6OqYvHPHGaD3KbuSuJ63jYSxS3FTfR3IW6F8HcmdM39X2JLclP5m0d5LuW4cqw+5rQINmWwODAW4
jwMNlnfB4U++afjgucsu+8BGbplIHiwhXNj+wVHzTSfW0xgomxjZ8j16KpHPXNmse+oh1R4b1wM0
z59NQne16KUK5y+Cm/bBTQ9TAK/Glne1butHJUh8S1X+f9XRtpB4i+gB397SqY64nWHRUYpF3dRK
1TP+Nd3wzTJBqrO+oS2vNTIimaI7myYGG5EkCsEjJTGOyx1KkDOXgX+WYAbgI2XIpXzshKei1WLp
BcUWAsp8WNuIH738j1SUoC2fpOVT25WGqrPeBvljCvXeI2joehCkkCeWNE5FX8hzdzlw6hlDT/Dr
812QdskNHBL6tmMvwX+sKU9cFQuFNMH4meLq8T3C4m6ytrlvUW8XD/pD7Zgo4lid/zrNhCFvx9p5
/Tb+qs80IhiFCTMpkvWPwe/7uYwcOdi5bBfIha6bPdZFO4WL/Nw2CerpdpuvqC91yBp7qhkS1Xd1
ijg4z2JEBX/kzYY3pFhZmu57WOkeKQr6fHKyBe+D55aVSbtrEGQ9WPbBpSKH/C//RcMLPoePIhk/
w2ijAiOtbXlYEd9u9gfUBZqlbKQLBCWOFC/tQ3jzx+XKBltEJy6zf5asSJzGh74IPotM76wQpwg5
Ypz/QF7XZXjzGgUfsLZSYGlix0yjExUSvpCslUimz+aL8UDlS68T9RoYucOWD1de0VR+0h6pOy/d
XUBR5yhQewPDkXnri7yGOk1qtg7evfYKzeVhisqj9IZDgo3CJQ6ZnWB0vMIQj7vkh03SB3o2+oZT
j+RPo3fDf6IUxliAfjGr0uemimwsbwBZ/tApYEsmov4TDfKTejzaQb7v6tlyS0EZHnCTvziVgely
cYvJdsLW/ak6p6GNTh4d9/hNgWqDtWhHDImQhfNxohHzYs6bZtt04i2JZ2xtVKUUMlGdUVY85uGU
e7YbFV+4x3miBtr2/c8TMZeZLLGZN8nQGMLP+u6v65Db+VwbUpHerzdZ01fZPyGn6yBJgIh+vFtW
bW7+o1aXKbnUxxRYwFRjmdZ27sv10moRlbMmQQs9GC2FE+SSBEnX0RrjXl7G0ppJ3gKNde1nl23i
X/75S8pXDyrYSqN8yQgOl9McYKf32RXMRXHvk7xPYN8bAuepC0Koc4geNLAAShnhZEcHAxkdx2Ou
Si+9BoAixVTOlp1pGI1YnkuDCBzmvf/ypmVhQb4qUg3GnH58ZQBYbPPXA7SZxJqHKk9xAMyEg/W8
+O1Kx8/fVBisLxHNH3ndRpcRxt7T5dsulPZVXTdeGHYV4Sv0OBIJ68ayWYATkSc1SK72A+68ePA4
oo/MM3imJv9G5FezKwk8c8AXdz47zkRbpCFnrt2bXgxITNXK2C5dA9qTHYDaO/OmaCFWZEUzBLFc
cP3mre6muIlFXTZWHQ1Ro8xhUy4EUbvokPyKFAnWeSLilLNCsZ+Hk+1euh5cCOxbFaq1I8GSw7p5
rCfAP3215OSABg4obrY7+8P9JJBnE0NfJAhvSRD0yTthgfJ6d+OHBL7ww+zXjJOAg1dZEeSTxScs
kAhYjHPEY348W9QnGwQdYBr+WEce5s+LyDejhwOJvial9Hdknglg8r7i1raHcafxuBKvMc09iE+r
644NphVjyRggLyXmLRXCj4nwtLaMBbBkSGxA/JGTIWOjK18vNhcwNNuBrd9ZtUUnlR4RMzFvEOWJ
gIACru2ah1Rb04l1FHbykwIwnIJM0K/ArmxsTgd6fD/yS80Ji/MEGX3gVXAjcHxpcLWj/8s2U32f
GKjox+Z8aklyHv12caJeY2wx6BUZDWQrDwDJxCEOvxDuDlHahYh9c9ys/Kp5okpIYtZPMV4HXFW+
5zIBuNFtmA/389FWHrCNdUmq5dupUKdl558oi/kaavWS4OcZD7TKjCougHo6FY0wxuTa/eLhuU8F
Zkz7NpxumDBsOWMJPvFqJpPgdqPa2qX3Vcwh8q6sRS7npmUDWibYqUApJN2IEZeFb9Llb8YAYOJZ
9y/AJa31wyjs50NTCi7b3FuwvRu2QUwspclGHnD+r97mW71SOym4bIsfOgWZTy0LgIlS+YnAWkzI
FLiQ9ZD6s0VngcvDiL7SHMnjdeHztc5/dhOpeuBYaiW27qtujTKnPOp6+NeJAmNTh3m3Yu6c+9UQ
Ca8htH49Zht9YKIUKDKMunin20gd1C46wjjM5EE5WHWVXtgE8MyBb6E8H4TGEI5zvdcqu54SoUPg
rYyDo1tCXMghAc7BHELSit/PLqx+HRz8ZFAUBv8YuUt7LFnGc7Cl00hxv1s0//c82su4lWnl3yfc
Z+B66oE/h4LN4VI8SaTh7UTp/Iu/0BnIIokZyZ2WJzSYWHAPQozRax+HCvTuhNR9jKtThuJLSMlb
RBoTx0ig0Hb/zbmTSBX3jhPtmKd50W0/2JFDQWTo1xD6xh1rR9vUhfqtLqMcZjHn7rWEArvhv0zk
MEdzngqMg1sjCl16q5J0uEPibyVu0FRi+2ezhcBWLrxotn/77lRWNkRe4SXV/IIlCa6M1n4oMzDq
2Yorg5vuwc+GPbU96/heR8BI3f7wmTNiisnidcnQyLemivh3X9uZyVmS4Fg1mAd5fEq+mQbsWK03
z1ulWsYqJbZsb+1H47dzfwmHspZBoQvWkgVpFdWvGPHZJeXZ53v95+8fr4TGzFQpajG4GozyClZc
Nb/KQXYIS8Z7L6MmxPyqh+6RPJV4uXsAxPvTKqMiMsFNPPhTCO+W8+QKP2s1rXUTeMcYVoUfKnMq
kr2bj8X54FzdAVqbUzWCJNLxUSbZFdIytUp1L/jPlT5PLZ/exK1iHijQfljK5UzRTPxWlN8nxhcA
jCn8KGUS5DuebnCp95VVm6sJd47ZiMbU/soxA3slfOQDGlsXu4aBDpWKGAD2Du84vOPqaQ/p6yVT
QlN9iq7bPPtm0mRA9UUq46wQwyWKuqZUFsjpvjB+fFgPoWmzeXWRkHJM9qeKcvpr4gYMwJM8Xfem
87AKnBcN6x2MchucBTbw0gmRRHvihfNsM7KtVIEx2VYFcjDOIqQcH7rxaZkLShnblIpIg8O2XLdO
oO4MEYF2uz5x7NkBolepYMNN+rueu7gRQlBsQDqirrJmnszEEJfqzgQf8QlZZsMi0bMoS7yhwPgk
gCWQ31+MD51go9X74Tn988pyGFIbSF2ILOfFpeZfZU2TSWsE0TjDYPvB+BUIqFTDpolAQXnmRKfd
YvUdjD/lgWtHH79kcUa4LXYCgnbsdWxRulKExoYPVjyny9+wZ/uF6HbNqbd/z42G4M7P1MIBuJUj
14J6cbeiIddJpGZY9p1wIlbpTtMPUxmbQ4TZwU029+VtD8062YpdVe0LT7dRCR7pKt/+Ri98cV9C
Ivwoc9oMdZMTRfDsAUxgqbWUsExnw6/g5LSJdSHa/ePiijXnNHaT+zWjDX8IUrPEUPD2l23Tdwsm
4eSqi3iWwUte3zHrUasISiBGWSrJUiZwRMKNZ7ebvDUaSA09p7zCl8mxFkvJw+22kEK6a3OCjUGv
J2BCXGlphUcrOogtal5wSH5rWqX4HcwJy/sj/957FDwAYSsH51HZHHKsmSsaXA4MPgylhBQKfEBE
KoDX3zSxH0GDNXXv5yZdnymzaUyFbZk7cGlMn01vcjCSLDZ4RaBxtKXSC+7TDQpcck4jh02gvYcH
YSGrqEQwIYIdHZX/LhsX4KOowk5/Dh3sZNKn4dUersSK+hhdxmIzmYH3o2Z7/83olaM1VwNFh7FR
Me6KzBi3uJBRe1Km9dB2S/DuL5yM5QzgR8i+AHkoAEthZOkFDSlGbRjkYad9lnJT2SwJZq2O6eYT
mGubhAGB9XUJTZqi4mOJ0LywCFqmC/2f6P8beMWrEjjd3YpfE7BudaS0freoX3bvpyWy3UXJWJ9P
cu0d/vGgDHdNRLKi0N/mUMPaMxJaDMuvCIcE/zB5mU/3xYjlOMSvkQKIJiJuysuHj1Hg9t4yOvK3
D3JYQelr5UO2Dso0+RzjtLBOQojD/Mw2ifoO112C/D+Dgw07IzOliMyNaccoiyQHcXLPqwXi/xUk
tZm43joFLXpMRW2tdUbzoB4jl9ImL/w77ERxNk3p/mBz+OLvQxbCFMyyd0kgfScAP0t+5olZkUk3
9t8vhKmxyusO6ZKC5AAChXTPMyxpLCswmGFVhVa+bdq8rwqn3Xvpf76oyxaPYX7jK1euZBssdZlH
ttoDHTukAgzWTKxo/7kV1TyD7xBmN5q+GVIhGPTmvn7edMxbU70AsrMtP8RdxYFMiKnQvbLtfnXh
4ndyR6K1HIkju9yEyOBfXcl+QpK85W8ELLUZkWPD8vvRaC+DlafUNbfXG6p7t60yN3U07LdQm/v+
FbUGahKFzpTiKZ2E2ZCVk6xHQZiPg6vrglRxPLnGTRnWPiHOj4kKG+BqYA3SSXDZQYNK38JlDohn
vxXKwBJHtZAUvai8iMRCUoIv4A7/SV39jQcMEoYLVTqmxB16ZDglJsY1XJO3F4cqcejrL9TFNpYR
K5MLGoy3k3i0ilkMUL63T7u9hqNKxUKwys5J/IOgZVF9XA==
`protect end_protected
