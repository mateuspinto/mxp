��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�������BjZ�K�nGD�${�5�`iFo(sJ��=�J�����H�p��"i��H�_[��eiٙ���R�H�Y	qJ���7��w�Z/6F��,�HC4�=fw�q�nWZ��1dK��]�:4?wD��gτ�N��:y��k���3��u�y���Z�6�TZ&� ���p*�XU��ķ���K�𪫧�t��X��l�y��"�/�g�,Kƣ�؝p�>�|�.5zs�(ٝ��3xdZ���ܽ�Irfl���l��l���&;��z,����@m�۬ŵ�6�r�����:X��+,78
d�Z����4^��������Z*��T�B�g� 2���.�b��5:�r�q{v��+s5����AP���A��-����M'R_��
�s����uo�#�Ϡ�����pɾ�.ӨN�9
�J�l�-�$Z�ϧ�4mK �RT+�_�*m�	��ك���|��>l�:v�����O9�E ��$ե�i��!or`�"�j��_�[�ui��M�v��W�(2�|-���C.<b(4=B?�yf�ᡷ�ڏ4�Z�\J$�NCs�� �9���5����1����Vo/k:�;����cƆ�3+��pA9���:x}�&�o_���_ڙ�$���6��.vʇ��qX�.f$�X�f�R�`���ھ�`����K���֤Z���.�,b�����lU�~o��׀א%�ZG�/��)�lk��VJn�Y�D�U�X�xY�k@	?/��8�U��LN�פ2�/��3�p3��2|r��Q���n�a�}�ʃY5�a<���EO�:��۳����Ȑ�(v��~WT%pg�G}
#��[}aDu����L|���F��Ǯ@��Q������-\�V��-z������x�$CK"^�vS���I�=Wf���Q�A\t.�Ed>rm��a�����{m��j���b�^��;����6���Q�״����ج��,����g���*�+d���� �(a���M���^Al���(����m�`=I�1�^���$*I�Mڅ�=8Qw$�)�v���g�eNzш��"C|جQ~<�y��_,�<ޅ���}4|7HEA�)�T&����Lw ���4F�T�>�5�����[	��H��ZQ��"g�MMjn���}CȐŰ���~[&�2�.c��ɘT�ɟn�%�@��c�VkA����я�Eˎ�m�u�����N�H%)�+wEc��8��^�c�*�a�D�ŝke��Wz�%$J���~<KGxA����e��G���A�c{�g�_�S�1!�y"�GegP\'�7B�/ ?ե���vM�ѵ�r.>�8��F+tb�:w�N��z�p�u�y(�1��ԋ�전���Kw�eA�<4�)�$�3�]n��$A����k�\���(HZ�%�s�aQY*Ś�-|N8��;֤JԬ�_�Y��9o���`��ȝ���

uh�ɇ����0����4d?��"��ׇ`�|f�lOVp�߳�I�_k`"-v{W��q�OG��Z8乓=��}����-��x�c$���H�����0G��@�Ύ�T��EB�Fa����
�������ސ_��0��-U�F���rt����Po��<~ID�i��� �^��T�q�8�+6��Bh�4��3�b��9_�ml��l���l��c
<7 �Z�f!W������{�>�n"�^�W�|�!��+��ٲܝP��u��[��\�C{ye45u�Q�w�����'^+|]^0.'�WH�!��I�� �]�BH�ՠ�([k?imђ�eӏc�%���\~��pD����ʋ��U!����ҕ9l�B�pc�1rG�'�s�X�����I�����xLY�������[NW�?�)����3K�H`ƈ�S+��Z�<���BǍ*p4=�ǘi�8�6����<��u�/-��ϡu�y_�'�����[X�^6I��8'QT��zd����A����\l��6�P��y�l�����aD l���A� P�L�6��V���	�^���n`JZ��Q�F���1'���J%8<��%�]�n�S�a�8�	�UAwo-|�5���#2(D����ol�n9�B��K�n˰ƽ��؞dj�!9��!�X���Ѳjz��f��"�Ql�������R�R����W$R��'��u��y�[ԍ��&>�Ӿ;C�jԌ� ���'SX]�K{z�st\Y;A�T�9b��x�(4� =��Y�oMk*5g�2�^3OY8�PjyX�ܦ�;,OEd:�{��ŵ�p{������o�+�yV��i4
�[������\�P\��9�O�gq���b�xv�!���߮��]��j�����OivzT��]8��Ke$WX��꘺�^��%O���$5��d2G���m���u��x�^�6���t�o��WV����l�F���q�A�]�Up$�p 5�v��>�uէ�e���gF�4���3G�K�㻋����7z?�ū*�bp��c����I%�D�a�7-���[v0R�3��NX?.��_<��@�'5���?�*�u�����eD=����~<����l�a!Fn�"3m|�?F��f`f�+��D�Z�ɮܑ�/�@����T�A���vH�1���M�%n�RfEV��/�	�9�)�uo�f� n������1���?�M��$K�<׼^s���1
]=��ց���K�[�i��0
HF&W����%:�\�9+s��KOH��{�e��j���x��ğ>d���M�ɷC�^����e�V�3���"S���֛�MM��,����R5}>�覓u2(dW��˓�a�/Φ�-�P�"��5�*̊:�_�2"�/m�<_1�qO��i��A<�L�p6@"�XE�;,.��=���ak�g�6`���m�}#��,���아N�������5�!�
�e�j՜஥X"��r���s�Y��0ߙ:�Xix ������|�~0���8�g[e�q�|��m��ӓ�7�PV��Ն��JՎ����G�!������y�9��;�����j$�$ŋj�4?Bn|�xжz�F�o5(!������G��~ϵxv��$�Ѿ�xG�T"V",:H\�K���%�D������'���e���%2إƸ����x��5 �O�.��]s�˟X�7�DZE&;���L�L���8�&��q�2�tn�>g�"�g���эBz�ִ�� V�I��b�K!��7��J�_�����Z�W�z����z�����s@�>�m^]��S2HZ��\�Gb@I!SE��ڰ��$2gߛ��V����ǒ� ������Ug����?e�F-��b�#��m�r�=je1����×�P����&�5f���LÈ53bGe���$EW|6䆊��Ē�~�/�F�|t[��5P*�&�S�2BhQ�C4̓JQ������8��	*k;���`�\T{��7e�ԭ�P�I'�8W�v���;"�L+4��Nu<�\���x��^�8S �^�om9,!)�S���x&�Q�z��Z�2��[g�F%P�* �6p����s8�n��'P�����p�󕊯L��ZN�x���?Z؍�0Kʙ��&|�1�ռ�<�����i�e���/���͉�o�9�u��G�Ӂlz�k�������G`�����R���J���5m|�0.v�Ή�Xu�A���5��㨐?�z�搪hN8����v x�k�$�6�U
��|�]��Ǐo�6ļ�B5B��  �3OH���麊n ���G�-i�01-�
eÒ��UX��c�˚+��@��EUp<�9��ut&����B9��6nXdw���D�[5 �	�]�H�O��d��NR�E�$��Q�ꍘ\��[�~Ջ8���S�a�~��?2�k8bϼj��V[	��[.�"�Q�.��f�s�0�] Q��]��Da� ���rj���O�tM4H�J@����tK�
��\��r�ά*\��p���v�*����i�!k��w�J�wV������X�*¥O�ET�l$n��f�tC�������vh�b�lSI$Ԥ�	���.��L� ��S(�ԩ2ژ��&#�u��	�����ڦ�������iB,����v��i�C�`|���%�4����Ԙ����!��.a��k��E���{���{ĝ�5��&�MWKʓ�G������m��V�P�ï(�d�f)�s�y.��(��\n	��	�>$��Z:�;��唼6�e"����^�1T�R�,�hH�k1�e�nJ	�N!������'a)A<�#��|��B�d��z�SF��<kf�z|E���.�sY����g�(.t=�ڨ�ҍe�c��Y3y��scQd�=:�0�,[:�]q8HF��Ȟ!M &����؋��o��G��^��L�u�s{�� ��yAU�+����D,g�}�fW��9���z�n��xe8~�^"�yGNj�h=GE��u%<J!I�
d�!#����ؽ:(�`�S�.�����e�hX�G�S���A]��W�IK�}�"o������)Ln��s��M�,�k�Oi��I�z��o�R7�T�-����ѼF]�}z��ߙ�^)��)`�T ?�F�7�$dCS��pU^X��f�@k���0�%T�S<M�Z\��hT��B�C��+V��NK\�O;��k���C����I��)�:ttg�l?F��L�]��h�i�O�2 �og]��PUb��^.�)�x��?}N3�O�	q2��i��/,���@�U� �]K�ĀC��+�E��)�qL���ك���$ ��0Eva�
���/P$RDvhT�	��M�u�'��Z{EX!�L>�t�U�;�'U�xd��ݧd������²'�,���T&�vU�	���Ǟe�D�=�&���d2ݝb�ϸ��*4[N�d������L�LF�"P�M��~�i��@x��0�{aɂ��A߈�*s�hNAPC�xr\SXQ��ia�꫒	sC-h���pӥ�ɞ��)Id&�{��=n�߾\��G͎�.h�ު˖��u�����X���)�ѷ'θ���-�N� ��l��۳�m��a��>s�����+A�xkٺނH�ר����Q���4�\���[�����Ĕg������B3$\Q}j���]sz�ty=U����^�~���y ��Z��ؔ������9���+��^�t��'5�C/��4��eF�YXr�qK��`t�־Ⲱ����䢈	������z� �c�0����Y�J�bt̗!�I�=��R_10����
BOtЛc�ط��f �b���(�T@�vW����/��*�М����e���bR-F{�S�y~���1āoH�
�%	��t&�{~�$0���Վ_�Sc*o�D���U���/6nɗ%l������D-�Gz��!4���ߨ�W)[r�y���zU�Щ��0ŉ7iKGE��Y�$e�@���WR^H��Y�@襻�a0�jPҝ�V(@��1�;��6��z=��Pmmc�E�몠 E�r"���4>��q�m�TGn��f�J ��*&�s�>`Ѝh�� )�t�ڨV�����$���f��^���y�r�o�m��!h����P1.Uy��<yk��\O�\:���ڝGqʡt�:a`��0 �H���b-�l�܃���CgE��%-��Q��|��r[�nHgo)w�.�{���!��*�k�K��k�y���q�9��Q[8h���/��C�/k�,SlMϲЙa��S�O�wF��б�;vfycD �F�HL��Rx�^UnL�RѶ~�7�H0C�D�?�����K�/%��Kk�,���\_���U�ܝ�j3������[���o@��5�.�����d�(�flAV��˽t�ȟ�����@5~UZ�$�#O���}q~5n����̀X��07�y�\Y�\�v��������|��W�C��cn�u��-B�|,�+v��aqvV��s�~������Y6��OW��R��W�K�2���deo٘!eм��J 媖G�>��t����d�8"�+���K���b���ikBl�L�Hס�m�_@ޤ��X ��%E�Vv�cL��T6�����I��a�{1qx����*d����:���/�$��m�b-dp�@IP���a�@�0�S�GŴ��;u����:��KŽA1)�����6��=L�dk|��/��c�8V��@$��1��FY�Љ��dAE�*O���r�6r���Qk����ܶb�j0����\���������3؈'P������?��}��,H���VY����/��u��@��&� z�+�r�~��i]����u��,��z	Lp�t��� �H���uR,|�ky�D�Ё�]�i}_�C�ف��'5�m�
v�S���Q�T��j��2.�} ��=����R:�O1�w羄橩Q�5�L��sSg�Il�7��C�J�M�5��L�S�y�+��Z_�>�do+��\T�Y���h����6��>)��!����B`$�)�Y�؞���9'��ڽ�������*CP��[�Z�D'�OD��ד~���4ϼL��6T^��[�=O�v��"�.fC���>1O�!n)\��W��s��A�=�@������1�"+J�U e�C.6~�HEM4-O�[�g�a��sʀ�d���7v��7��]a$Zn뉭�p�T�kûp�Z�Ğ����Ӿ��JejYJ���'��^��eb(2Ds��|9&����k]q�%h:[�@�{nz��35�=8�R�1,�SН,���
�
J�&�����ԉe����c�V�7߅U����@�6)����!���ڱ�뤉���Gn��	\�l��M�jZ����7��'�5	��\k���ٲ��s���i�>�$�u�u��|̞avp,\�rN�>�4��+����"ݗ#ڠz�(��'�_kl��)��JrQZ>��ʵ���^��u�5%B�L��]%��f��|w�/�Bh�T.I���c#����/�!��E�x��-x��o�r�MːfHoޗn�r��[��9_1�I��-�?������U�m�{?���҉����Fڏ�
���_�ּ���V<�{�!��c��Ϋ����u����H��=j�8�|*i�����E�h=�����Mm�Y���=\p��]�_����v!O�SҪ��{�*�b���e�J9Ľk��+�S*n�䁧�&%ްJ����߱��-�>������:^6ٗl51S�F�����[?�r��7���%z#�0x?�y�S�U�B5s2$?�4z��*�@�,�_�H�|�����6���g�j]k�@]p����mx��/�<�`7{������љ�| �/V����YaaH�����H�𞇂?F% J�ؘ�9�JT#e8�֕8��s�����V��"���R2T�]�Zm������H�G���������m�i?T�׹��C�۟,R1M�O���RJ��� ��U6%�;�MCR��D3ګ�������<7��R�IL�AhG�w6���/��"�����\����/HUW�N@����@��o;2аh5a�̀
,,�BY-��i��nΒF�=�.�t�0�7�Dk�Hܩ���*���F��@M�US��Vg�q�VNq���H���=#ļ�`�����ֿ�k,�4���ʕ�Yb��g��ж�$а��ß�b@�;V9���<�r�P7��� }m�v C3���b���%��ˠ}�~���R�9�Q;��w�� Q�e�D��%�f���R)��u����2V�%U�����>	kŗd��;�(�����h</�"��r��~�#�M_9��>�a�SG{��%�;8����G�y�������H��6�Dfnd�NE3�L�岽�T��̈`�|ZFճ�	K���k��^���[4e���|��A����Od��e�K2`nv�U��7��O�����wFy*~���ϙ���������:���Z���J�1�F�`����G�=�p��Ȅ3�<e#�&R�{�X�/Q_&��,�����U�N K�\�N���n%�*���v�&
c�ᘊHR�M{)����h]g#�[՝x37V �0:�bFw=�p�*�*��SÈ�\�C�א�>��>�v߄X���t�nBk]IѴ�T�;�!��r$M�d��@��b�X��:��]��&�^WM�ѣ��L0����%��]��%�=��fYϕ�ϝ�c5�^D�)��Z�+}�8��6yA{ 4(���(L����v�sD�vTy:�)��9E�P�ߔ$q��bmI;8pa_��37�F�`�ئ���\�;ҟX�b�]���*W	&�F� Ҿ`	�����S?���f���l@�w��YԨ�)��3���[�j7�i}4��Ǝ��2{=ư�$�@ w"�v�+)E?����ӥGi�7���r��p�Ff��o�)�Z��iU�PfTQ�����/qr� �����9��k��2*Ņ�gD(�q�:�RҾ�C`�ؘg��j��f.,/�j-�S: ml�Ζ?���|DW۵Xe7�k�]	�=��$��<�D�V�)��[7�������%��ް.���td�Y7�b�?1�������tTe����w��5R\�vg�~��Zx}��s.��Iĝ]>�$�>��E7�	3PI�m�2��
�>߉kf� \
{ -n��F�e�[[���2����UT./>��f|��q=jV�����&��
iM���u����\�W�RŚ��'��<mΜ�a�p�2�R�xn��T����!��<��*C}	�0,jIx�ƏuW]R���4�_Vb����!o�*9���e�<�Mѝ��؝KXmL��2�%U�4�A��H1���߷RQ6����Y��=�`��E��yǈrs�c1���pݶ���T���w��MIz�,y�]~�<�T��	����m��w�5���=i�p�Nǈ��M�a#��B�E'��3#��FWZq��2!]��?��q���\Do��U�!��3H�i�_&i2��� 5L��z�5�?�57˙;F���J�qO����$<`��?^U�u_q��47J����^Wk)*7�����ի���!aA��F�{�#I^x��_�]�k�򺮜ωt�=�)�h���'�c879�5d�_�*%�fU~��G�GRP:�VL�C��3�����5:v\H� ?vkl��v��Z)�#;QL!Sg_�\�6��c�6+�hǂY���Yg�Ѿ�7�m*k�E�\2|*��gռ*���Y�K,�JdI�5�@xhL����eד]�'9�J @�S"� �U1sތ��p[Y����%�ɗ�F�74}�a
t���v� �Q_ʸorfhJ��H��l�
������q��R,��	U��J�j�X*�o'�钗��b��u#��q;G|n��y��{I�������(f-c��B���Q!���\/�����\pfaB(����r��/�G��X�t,_��b�O[E'�R.�ᰑ9� �MGZz"A�K�ti�f����$����`��;'%���wj��q{M�g�����*����ݶG�+[|:�%WN����7�@#Jiq��!��\�Ի�G�̜�����Q�o��=S��ǂ�+�^�/�g�xǜ�`z���`�WuoU�t�`B�͝.�pˈZ�}i�B:��O����#ӟ=h��4���,w�����G�OVv�AZ�Ho!A��u��>u1ׂ{jMHR����� ���n�i=s��&h������!tt͗J�*���
��w�e^��[}�l�I�[�U(*�vO#1EF�ў�A��F��n�xX�|I>swb	
�CZ�L1�@�"1X��	�	�;i����j��H_�j��{����7��f���>�>�EX�S0��Q:�L��I��0:Qo�c��,f�;���>����":)�#��F?�ƴ��X��z3#��j�زu1�$��YGM�n��Y˯�35ܩ-�cE�B���C�Xy�l�R��4�k��ǹh���SY��BF)6P�������(��`��@kÇ�Ss�5)&�?&����7$S��Z���Aa@�X�{�l�(xNa��U��[�%v�(�+�}0�:,Ț��,|ǀ��:�08���vl7����5�^��h�h-S�P��F������L1�o�f���ȭ��9��7�<�����X��x�7Og�$^���\�C��m�z�'{�XE| ��~.�ʭ���Y�w��&yJ��\q.*Q�a���T́�6��f[.m���ָ�&��O�?�w�,��Y�r��ex.��9�Y�<u��*H=B.�(	�����w�sBC�}�f2�d����qROa�W*s�1�����6-'�F��VC�E^=��ע�_�! ��i>p���{��|~ʭX[)�`u�j�vs�{pu1&n[a$�x�&�֍ ������C��<"�ژm����{E)�Ɛ��K�53ߨq{���ԥ%��{@�l"RU��qu;_ǒ���az��Yv3�-�O���1����0�f�U���[�b,�=D�	��h�7��t_E�@u�3=�T�V��|g���^��ݦ�&ɚ3����7��O��}k2�>�Ԏ#D|y#�NSj���L�N~1fW���O�P>ە��B�+*��	O�gD��>�ͩ�����������6�3��(5[.P��e�4�:R������
<>��4��a�ܢ6�Q�-ػ3<���Q���ҒjLhs��2�HY_6���K;c�f5ԖT�u�g���J]�i�TW�(��d���;�I�t������[�b��P,�]v�$�o%��J����.&�*��#�W#��&��7R~��,��G.G�sR��`ai?�P�\�>��l���8�V+b���9��[�Pz��a�D��XZ����҅��s��tH���e��W��N�&���U��|�>C���O���&�?�=�}J�+�/4�����6`jx����^?���a��G�ALV�j6T��0F�:{��\��V�owa�PB;
+�G�1�2�S�ܛl���F1p[&��Z(G̕�����D��SK�5���n�r��(����;�Ժ����J�W��o�H�BК��D�Mb1#����C�9�d��e�P=�S�ҸJ5L�s�P0���w�o�$<���HO;qѤ�� ��D���Fή��o${n������$Y"�d��'�+�Y�19�R&O(1�$o_y�ϊ�.�:�x^%���egS"�5V�"g(�Qg���2�(K}\ح���CT9w��:^�����F	�ٯ��	���Q'�c��A�� ��TP�,p��R��*u�=O/Њl;��#H��5.P��Jv�y2ߓEQ9�S)��t��݅�=��&�9�z�{�*�|>�PURĎ#����D�� ��I'O�"x�A��4�f���ύ5��sP�Z���r��T?�U�KH��g���O��_>���Q��]r(�P���Af1�<���<)�4�d�f����Y����ݖ�ޙ��ԫUX����ĭ���:Z�'8՜����6���z1�[z]t�,w�Z��b�qg����,�}�T����4�q�Ï�t�`i�5��"pV�"�aPP��}���"vx���E��n��KT����?p�����L�_/H������q4\�W���w���7%�gy�3��]���^ص��W:��(���7�ޫ%%T̄Y�G/�EB+�St���CO��+��~�N�i���h�H��	�&�f�E�f���{t�	�R��`���?�hUÂN�̼�8s�-/)�*lj@v���c��a\v�.���n��h�12�L|>�HLfZ7l��N=
f���/�^Z�D�:G}��;�p�K�RP��zS�m5N�`�l�ۓÈ6�^#"���~z�o�a_W��֎~df��w�$�
����8/MЇ�`Zĩ䳳n:i&Ěd2+
��ل�5�b�.x�֐3�H�q=���r2��-���d|��<5K:�A�2�����u�'����޸Y�u�_4w��I���ʻle@�����[�6gaur��o���]!-$	��줣��#^wke6|�:XHA��������AB�ǿ��.qB��gg����r���HTk8Tx,�,:l�^�JZ��ѩ=�����چ���C��Fm��S��BXv��8�l�!TQ{����A%"D�h,��P,Sr�e�F��{�c����2E<�|r��qeO�zn���1��K��s&Q5��q��	����B�?X�U�L-"O�����}���	3�ȥ%�f����s�l\����(��'��6�L%4�P�ȋ��^��^ĵL��P����0�M�׫�|w�d�3�i�9KA�i��e�R��`#��N�7��]���E�,ű�"Ў��$��N�SR_=��6&@��ȝ�s2�u�;�}�F�I_B'�[uz�
`ic�	�/�t^ �+�e����`VL�hl�)r��Ɩ����	�f4�Un��G__0����	�O�M�<m�V������O��� �*4��n%
����s��L;�S����=��/+��=w٪�4[z��lf��J j=�xc�L�\;��C:��TdcKX8�<�A�Pj��Zoq�2"w�cXu�I*S���N�(�%{�t�a�+@�J���J\j��C�棬�1's�S?���𪍅�y����}�E�Ssy��y�M2�ٲ:߱�'YŜ��
��c+U�������1�"������T�����!�Z��֯9��iLS���mq�)N|`�c`ю��9�WԌ������\(���!"�E�t̍yW^x�[�B+Jѷ�*���K�k����f	����8.��&�oβe��,D��A�?{�P?C�Nw-���ԇ�#�f/C�_@��j�w!�髊z�sv~�kn^H���/2гm�6�)�8���c:7�=	�W:�2�i�B�5л�5C�.����c�5�<�y�q���D����;��lkܵ�0o��_�d�/D�d��P$�a�)�y�:i�W"t4Ζ����8Z�_߇�=�R�m���[A'��&b� C�[\ސ�R���_�n�z�QE���0B�TbݶN��$����f��jb&c�V�ji'5�>dV+�a仄 �q�f�b�����|F�U���x�7E㞴&�Jhn��*5`1����+Bl�0F6�-+��Y�e.�y���h����WN�ʯ�lS$��j�g��v�I�Y����Xwf�S-�����d�Я���{����(G#���8�z͓2��;���X�7�#��1���Kܞ��SՖ@몫v��AĽ����5r�	��2�Y�J���W�x�,�� ��G�C�]��U�@>�G����VRWN�p�\20�0U�=��b�q��xI����Eӵ�9�҈+�����|�N>��l�E�kgBMA��00����Y����J+o�?���P����,��N���	�"�A��S8d.�VG6�C�0DK8�n+��$�e.�������i��~�~�l_*������"�D�4��x�+u��u
�?��@�Z%�B�GMld���_A䘿�ѵmؚQ��qR\��٥ૅ��G}�^����	��|M��eI?�.����C8�,�O���_F�����涀=K�S�RT'�t��[/v
J�Z�WJ4�7��b;M �����,�Y�`F�@�����lnm���c��&������Yu� ���jPʽ�`J�I8Հ|'{�����O�z�~���rj����!u�gʂEa+Vb�Q+73q�K�����sf~����ܳH�^��e�V�q`�zA�mT���j%�ח�h�m�r����;�y�����6?�r�cH��e����a�n ��'��(doý�Y�3W�LJ&�0�gY{˔���r�������R�r��ƥ�M�W�DΓ�ЂSH��x>��77T�C�&>���m��D汅��PyB;MCF��6T�/~��ｎ��)���Vjĕ�LB�I�Q�)��(���L�'����jn��WR���pq����j,�7�:�z�E����V�x�({���w� ��n�X_N(�̙w&�F�d����fA��:��{ч��y�
v-�! L�߮+I0���R���m&��0��[�f�RA���o1�� ����屙�N���P��p m��E �=��Q�*�/" {���K�=�	�lշq�W���!�Up���E2�Gff�@-�z���9�ʁ��Hd�鍝;��΅*uz�"�hU��<8o��
X�.ɵ��F���j�Ĕ�d�1��̲���'�r� �;a5��H��>����3���x�s�#���uD
u����t�ٹ�\8�����q5�W�V�T*����I2 ��NUL�U���B> �XA�o��ݖ$�E?z��4_:�t���E&��4�[V^&�1���gB'@Um���lqNy~�5��<W�Ni��+X]+<�u�/�۪���x}����Z�����p.�Y����^z�;�����v���">�5J���c�QD"/{ӓj:�[h	�S����d䒢*�	A�����;�q鳆�!1�Ӳ�I�	�o�	�����b{�V����n�U��h�2����[��ܳ���fxk�+Ԝ�(�rG՞k�>��ܖڽ�`Gϧ�VޛQ2�oٯd<�JUB��'4�L�~�(E�u��UEƳ~���T.�_޻g�|��
.j��%JT�;��H�-�X�
`�"��+݈*+wd�ށp��\��*��5�#(e ��ഓ���2B�ԏ�iH��|��c��,��(�&�ݪֳ�u���Wk޳e�6Z�aq=���~u��CvWR���}��{ڒ�fg��� t���\NB ���^�"��O��C��,��f$0��^���u�WQ�h��  �%�!��n�H���*疀`�!&���R�E�Q2s~d�*C?�J��y
4ȕO!�G�X��R>��'Q己?�B����A�t�����tZ�C3�:ӔI���Y�nhu�Z�/t[<����h=��a�����:x�rbZb��	�"��bL03W����q]9�����sc)��_�lxu;�!1x�����-�Oh$qu-�ǎ���q���J�M�}��`�[t����2����Ys����|yU��*4 ��'�#�+�����s|J���g�͗Ҹ���B֡�����P��e!��j��l��T;Ƿ8�Êy�>�2�`}
�s(%8���#n��ub��"��kw,���v\r�w]�Ն!)�g��Eᷫ���LZsP4,����K���!*�\� 3��8�%Q�i�O����Oڻ
垒�z���q�D&����#?n�d�9#WD��?�^r�@)[��e��8?g���d��pb[�CS�-9�W��g����B4H��l�mS�ը����23�U���RU@��P��8PԾ�����מ�C��Ӹ� ��i�C���em��BbA�sL�Ҟ�Mð8&�7$��P{�/��������O"��2�i1&�N� ��}��q^i��Ġ��B�J~.Q8g� ����=7�W�0{X�AA���]d�[�ra�(s��7^]O�%P�>�'8Ծ���%�d��Ƣ���홉��4gI�|�p�L������_,��q	cq-���]��O~<Y]��dG�H1�k"�ͭ��t�Pe����
B6=*�	%�پ�L��1�W�'���	8���!���_��l���5��������5K�D��HW��C�s�I&�hKc�gK>�$�+��A^��u��	���Ù�@y���Cgl3��)Y��צ�NYUB&�*�RAi5-��}�gm�H�7n��7p���F�~+BzMUl?�����!���S_y�8k�wsI��E��5�v�:������ھ���5�m)��8Q�26�5�/�A�������b>��Zj��{���f�tj��|�u�O�^앑�Z��h�;��c(�$�MSK���&V�������-<ץ�-[��m@v��!r�ǫK�(C��,��6��$}�c�$	$�I�r �1���Ξ�����*/\�P"m�L�MAH���;�RIH���s�vt@d�Jo����Fk��*qq���8W^�����-���\GH�Չ�o)�9-��)��l�g_Ԯ��h��+'��ٜGp��A,m��2�j�/�V.���ȹ ����)�`l��þ��X�X�,�9��j[�ńI�J�`ឝ�?�P6+�x�@6�([1��,qouF��!l��?��	S|l�	+u�0G�9�s+������B %%�&�x������RC�X4~�!�C��A�9��(w��=�3��T������u	Ç�K��K�H@���R)i��:��]��'�X�/�n�)��1A\�Be��:�[�[S*Dy,�ɿ���un;h �+���i�K";o���57���"�s����z�s^θ<����~b�oc4�`��.w_���l�Bz�l��<����u
H�������XD{���2U�ύ�#�}(FX�n�e-�>���f*v���ގӳ��^��HW8��.ڻ���F|�)�L�M�N��$#�v����=�b������2�� ����D�`*�6:�:%���~���� �G�z�. ���O�/Z��c�����!6�m�C��O}B�����,r�r��	�^9��]�wZ��pm��"��i_�%Ũ��l��f	�{o�g�ߺ�E�d�6]mp�u�['F�Lrpj�Us��\�@���g�ݡ*�C��P�-��.k�*����!O�(���`�
�J�����ߝLS���r�	�M�,E����(Ce�K��M�l/���Pro��T�7�����b����	��e�p����~����:�W0�������z��"�#��"��dN=�o�[���!_]�YW*zu*���aq���R_{w���Q���8:��ʎ�s*��x�΃%�=��E�%��ɏz��E��� Z�_S#���yh�7.R-�]<��u�~h�9xY[����j>��qD���ēJפ��bp����?�����"]��m�3�����S� I�<����C?�2A;��96^S��:!ݳϲ��ᓽ:P���k˜!Nn�2�X�����ȥ���:���륵���GVά;�F���L
M��h��a�}�E��Ro5ݴ�0�0���'�W 9�G'�PR$�?)�)���<#��	+�7&ilR��j7Ҵ�'G�u'j?#�S�(�6Q#���E��
�1S�~��}^�y�?x �s�J\�/�!�!\��gLGܿ#L$~�<\�U�JDt��v	���� t��trD�UBD��9��<s���+����A�H����v�����f����(;Z�=?��XǕ����x���j�;�^���=O͘��d&�SlC֊�⊦��HQ/\�D�nN�' �]xh�\7cuSps��u�{f�z-���LZ[��z�(Y���|5�>}r��~�h��w
S�Ψص�R//(��Ev�El(�ϑ����^<�JrZ�6 �tj늳f\�2Q����K���b�B�/!�\�Z��oY0������� �8��r��I%r��	H�@�
ד��-�~佮8���4��*��?*� ��U2N����,����^��S��7ׯ[��)\��n�g0�g�s���ǫ��g�����\��k5�}���BF9%���/r�;��q���=�֝�^�Ljۂ��9�$�nS��#�1+.ctIp���T����� Ś����;ª"�h˷nǂ��L�w�}.����:˸���}�=*_d����q�cӰ��DJfBw��g��YS]K�_���4T�'�A�iIOd,�s�tG@�{=X�|��cM��eEujY�c�E�k���2�]���?�7�����m]��S�>7j����g"�ZWz�r�X)�v��2k�.��N�-|�0�6��~��?���N���^?�$�fN�w��l~���-YG��!"b��,$)o��j؎M!�b(o]о>�O��\�j�L��*X���lQq�e�\l͔��#��F/b���@L��B!7aҌ_�����u�_��Qb�q�e�x��t��댘_=��Ō�8���3dָ"VޞY4g�d���"�phH�y��!�hz�A_��.|1VPh'&4"��~��Y�L�g��<Ar�KEɡ:bf����+*���d�ųO�ش���gY�� ��ܳ஄�6�F��e��l�Z���F��(�L�.�.k�Z͐�� |K��
 ������~���.����'���vO��=�{��u)[�7�6ύ��+�>
��Cŧ\�@	"lĀМ�[�
P�ǖ�5�)�2*CKG�[h>� L��v|�Wt�=W7d��\x��@��l�H�d_c����,�ӽh�瑷�Tހ�R��Ɏ�N��Ԉ��R�]�z����&�n=�i��}\��DƣE�r �8m�!~��� ,,
���[x�%�b�L����K>y�)�8��Bۊz�
�3q�`g[�am����ji�������=�6������N��0;�ݬ�<�����4>@��_��_�ZfP�	�(�}�#,�Zp����M�\�3�x��a*���b7NeU��!�hΖ��u�!4S�L�ym�,�ڼ�~9�py�1�q�݃�,����94�I�>��Ο�� ����(w��K�%�?�b���fWy Dڄf������:����ա�,[�H�+�D~���;���V������\ل�N��f�!�7�Tk}����JX�m
�_̛��ȹ��$߆�m( u ��5#���kA� h�G���j�e��������)�n,��>���3ޜ��ޡ��䢖�����%Ø�F@�P����+�������ӂ���)��f$��R�ä`�`����4�B|�'�5{G�Za���KG����B�ܩ�:򢪛ҳ�-���b��Ϸw�1*��W�Y���<�����	/Q�?*g�9h�����T��Š��%�i{�����5.Q����K�^�Kŉڴ	�z�J����qU�I��ቃ�6|ve��K~�/�������׭�L��G~������v��O�	��I�����q5���{;0i7�z��o<�~�?m�N0
vm�&�WL��4���[���p`�G�&��+�f:_L�\��C�&�32����Z+|��ve����(��m�U�Ҭ���iP&X�wk�Tz�NS�A|����=�fGl�i�5�x�M����� ���w��%4���=KUT��q} �ć������������F�Q,�33-m�M¯���T$!��u�hngy�"%�qBo˞��nH.q�K�¾�4��:3�_�(9;����D�|J����L���U����v�h��`�y���խl��L=�������@�pCw/���:L������w�9���f�˲IG�
���ʆ4O����Wd���r9}h%آ����)?v�&�@N�rflI.Fѩ0e}Q#7_Ҧ }��&D��N�i���@�p���<#�7U�ѻzp�RJ}��� ?'^p>�L��!�`X�N�h��QC�o�s֚�Ë�� ��s�=~���u�MS���n
z�B�����9�ك����9�>}J�TO�D�;���n�Ej0X�N�����N-�7��̘[V��M'M�dq4̰2x������<:g�t���%��&z�'y1Qw2ۉ	���ZH���3mXVq!����i����.��Ģ�{k1����
����v��F���l0Z�'���k�"�p��{���r,��Bp�y�!?v��b�3�B̂@��c�\8r��0ݼb�*B�w:�˟�G'\NS�r��Djr��ԑV$��kc��l�bf�_>�����D�n�cƳ�PG|��v��ǭʉj��E���ױ2�mD"�:���V��.�![:4�������u�t�I�`<�B�\�u;�ͫV>����l,���4ʀ\?U"�a�F��5�_�����rG�'UY����=[Ǳ)>� ����=t�ޕ�^�1�-�U2	Z��p�!O$8IfO�(�����
�fe��x��F��B��ʷ�`�rr�=�(d�rT �rt��T����j�}<X�4�a8� ����7���T0G���G�dղR�Y����qي�����Z�n`���;��ʞ��]��U,�/��}�_ƑV	��8~Gw��]���5�g�uǬ�sE~���$��_�ޒ1�9�jp�l��N�58�O���t�������Je�0_#=�Q㙍�\)�X���7�	��	cD/i��k} N�'������8N�։��Ԇ�&*#K
Ð%Գ���f�l�c��!e���k� 8y$�0Q��w?4C����A��MP9����1�bS8T�CƔ�4ˁ��V�!���y���O"�e
�A��RZ��OܥU�h�-Օ?=�u��<��&�Ü�̳G��
T^4D4M�Dv��O�{��:���|�� "%�����/!#⊀�j1�1ƴ���oFW��L���oԚ�w3@rxjw�Z���Q�픰V8T7R_r��6�Cj�چ�J&��ee]��(�h���/�r8��X2LXx��}��e���F{h�Y�J�5�����XH�e������_�i�%(�6��_a��FG6;�'<����Lfy��)�z-�&#���j+ݣ��EM�p�6�g�z�9��j��<"z����|�l`��������i��e���H/�:Ahc��F�=M��B�{�鯐GJ��`�3!��9�Zcéwph�S������J�@�s6t棾��F�\_;�q}f�ܚP��AҠ�.��烔1v&E����`������+oe��yJ�f^�n]�mio����!I�Qv}c�R�p��잫��B�"sУY3�2/�hy�ALx'/�`����Sٷ��́��̽�*7y��ՈYs� ,��I%J�;�~O�/�ʳ����ׄ�i#� u��\����@���t6=�����Vi[�a9��\�X���� KKBα��HxDLy'U�x�C=F"	�4w��a�َę~
r�'wJ�K�1@���X���j+�*��m�%p�Dޗ���I�r�X�X�î {�������G�V���<�$����Y��=Ұ$mt��R	D�}��ɺS��ƾx�hg3�XP�DaLiY"xȏ��,��K�=��S]��i������l�_?Ճʳiw��������P�Q�^���j����)����  _:�fݺ��ᖽm��4�����G0e*��\��z�z��5Yg�#��R����%A��;z���?B&�X���͘`�|��Z�We�3ur��D<�-�Ui�+�z���E�T��p�x��C��:�����g[l�_.�ҝ�=��B/���ճ�Β��UH`���=�1���O=N>W��x��s�WO��DHwr���W��+����`���ٖqSF&��E�-*w�o��3�ƄG4��x�Rt�F�,�y��-�᝛��p���'>��r�lB.�&!O(P:�=������$��_�dXu�bԅ%���웲�V� Y�"Vj���s.�N��_'����������6I�V�T=ԂԤJ�`2ۖo!�m
���Q�?�`xo�4�6X�O�i����M��� �]b؈��T�Eo����%·A��B�r6�D��P�B ��𖔃:��5]7;I�=͓JL�2�k̵�٧�=�7J���K`��o;�s�
�Z���)I���e[�Yq �.����Z<+���pj�hs�w��)5��2��/lS޴Fꪆ竼�u>�d+�Hx�Ʉ�k�|n{�w$̧:s�)W�a`��b�L0G�m������4��
��)��5��r2T -���J= B}�����1���q���S��y@��f}��9hx��,Ңbj�n��=��~wu�ќ����p�i��c�i)ԏ���^`����U8"�>���N���cW��D���%��&�4�3��� ��)"���U�1�T�T�jV�H�Rt!˞:���M�?�rX�(i*�-dR��W ��t�_�{H��R*��h���>$M4�`�0v�P,ʛ�|[]�/���
_(*HgzƂ8�L�˵��jLr�ۃ,�B��m�-�
bw�vc[�p��o�^X����ȚtWS�o�u'�$}���� ,D͢������I���T�7�j���Y���e�'����Gc%��~d9���<f��N�tÔFhY����5Esߧ�2m~X%�=#Xف�������y�u�n~h��F3Y�n�wZ�Ic��k���C�����S����N��q�/�����x��5BM�?mO��yýD�?�jM◕��2���v��L�-�%�����c���c�z��$!/QmX�b��`H^�@,�o#v���JܦO���%��::����M�(�^�L6�b{Zkx۟��<w4��'*̛ˆ)�
u6�q<�o���m�(t|߮妑��<�;�K H)h\ =h�:���hCk�Mw��ONG�&v�
�)>�0@_�_���龾@@7,��Eb-&�{)ʧX����:ʺvK�9�,�y*^�d��ԿtX�J��aP9#8�\���K7:���Ι?Y�>1��j೾]�lh�s��N�q���So�v�?��cg
Q+V����?/����7�pK��M���|E�sL-��㞑��cDR7	~�-�W;�n�\
���O]Ǉq�4��w�ˊ7<�كX�R���V�D(�^����e�N��*ep�F��}��ӓI����)*���3�ҏ���|9g+p~Y�_�Ȼ-��J�mz���0B຺̋����4*� eI±A�"�!��?��͵�xQx_��{׺ԫ��F#�������s߈����6���pB#�
V���o�L{��� 9�����o���PJ�V75��(�Y��ŕ񰰰7��(Ė�z���x�
e}`�S�������?��q�M�j�MY�{ZJ8����>��BT�F>>c�x%|��f�
�s*#>�L���	�1)�1��@�#�[j�0e��u����.eq	ؼK�6{�2H��KL��|�]�D�W\Lļ���R�yËǜ��o~]=&��Cf;I?������h�a
{��\Yy!+�(u�}���o�I���y��l�7Bm�6��,�NR�I��S�P�c2��
����QD4�r����6����pr����a�J��a��<�m��c����?���ʷC	�<�o�5����t�z�"�;����K�H���s����hK�ƅᡞ�pیT��O��� 4z��^���I�0���C���g0|��5�H'�͙�o� ڈ(��D>߳T`2�V�L�u�1Eɟ01�4����|Ț�p,��B���Ah{��#�Fq!��`8�������hf���0���^f��Fvĕ�1�bo�J�H�
��#��f(�,��:����� ����u�R4�2��M��ߘ���;u�Ԩ7j%QACqaW#͘��=I���W{��rYϚ��l��Q,��*�2��DT�vߪ�85�����:]�L�(Ƶڴ%3��B�b��c�Q����vdzH��00�P�L���2"����$<RߤM�6$  i�If��F�>�#!�A�"$1`SI��P
�:�絗�z��}�����q!ĩ����
C�/LŴB���Xj�?�d���d�D6��Ƚ]�1���F3�b�s���R8i.�rv!�[���>J/ɚ�,��t��Z�#=-؎�A��hF�N���>H����R�F|,v_��j!S��'�
��65�÷���q5Rk�2���Jbj2dT�Y��l=��� ��o?Z�w�ܰ�!U3�H�0i�q�����	'�
�T�y���Ǎ�e��>>H.�:��X2�T��I�tE���'c��K� nDˢa i�y-��2���{^2��Х���]�5W����eebD�SX+�4۪�g�F9b����{�LJ������x�AU�OrD�?%��NEP����\v�S�L0&{�39�*G� m�M���?�,NT.B���H{;c�Y+��L]6#�88Oo?���_���*�u��ˈ;Q��6ڢ:l���B���Ѯ�xl�v���!et)(����+cPn�|�?~�C8W¡�ދ�w������C E�7^�1Z��p_o%�֚�l�C�̧�O ��ʰC��M�F0��<��2�ߍk�`Z
�2�����{��]Յ?��Yq�!q�
KK� (��\V��%%g\�_Ť�[W���� �<]�4-��(c�j {S��L��H�I������QR�H`��-����)�CܧP�^�R�E�ٗ)��*�:���Zr\h�s�����wޣ�c;�_�4�����{���X� �1��	�:�7<Z��C�%*�N�r�v������k��>��-�
���<l�?��R=�e���J��@Rݞ�*�����ݭѮ�v�����4x>�2$�9��:ϹY�3�F���oݚ����E�Y������S��y�wD���#�|vam�=�	9�H�r�E�U  �����K\oHw����X��������}�\ũ���oR�}�Z)%�>%5`�D��^N�㧰��D�*���od#��XwOIR�P�X8��g-
\�v�[�Wـq�{�������l�m�����C�\�4]��@�PQ�5��t���.�$</:t��'�,82ht%��?e=�����w��C+ǘ�V��,uX-N�� X��р��Rn��mJ��X�w�Tt(i�HN���F�煾NWr��S�����%�W���K/�� }n�.���,�=Ө+۶�,u�q%x���PpL�*A߃̓���:J�;�+Td�L(��WA�u|c�b��2g�������F����wp�t��:l��z*Sb퓔�R�a�$�%==���bF��7Vջ���(�p��=�)0L�139����\70�e���n6��w����*j���N�o�%;�x��6��u2�@�S��ZL|/W.�i�*s�,j
�d�`t��Q �]KN��z��7��sd@�9��96%n��6�c��'*���KV��e�=����ry�aŜY�����|�H��^r|���H!LQoAGr������0`*��ֽ������͌���|�F���Չ ����7��W�J�F]l�o@�P��4'~�o~���[8�s�4�|���'��+�;� 
_�˯Sq��`i(����^xA<����V���M���;hzc�	>[l����MVK�����X�NC4q��H�A*{s��ɬ
l@���Ͱ�:R��e�-�@-�-Z����)�1��{�D�,A6�μhR�?�W9_��wפ#�^�ytX���h���	J!��|��H����\Fu�h7o�H��=��!b��Q0���Ӕ��^�����#�)�r���מ����m¦IDC�46�Y�[V.�쳊�ફ��� ���'Q~��*gZm����Y�ƥ]������H�Níέ|�	8�бKkSo�"��,J9�C�����\4���c�'	v�!u���W��'�؝j���9?h�0*���aA}8�$ޟ�Šr��I���ќU�M��r"��+$���NR�2L�C�7��MS��(� �;���=�����o*vq4r;�Hh�͈�L0��JDr3ԩ5�y4���m�K�9�kښ_��5��d��L� ��:v-~yfG���Y�@�U0HT�$6=*+*H�T)���Oۏ���K�8C��V�<�=]��Z�T�e���i١"�O?پ�<+r@}8f#�)�uO�S�<f��aD����ז+{R#Ǉ�؍k�ˠ���.�h��m7���H^\r��k�+��2���&��H���d�2�ɸx0U�X�͘�S(Iƻ>�������ym.��<r���j�
4.˞��P�:�����NE�v���D{����4n?�Q��������dR�v�6�Β��]	]��	ֿ ��C<��)��D������f۬� E�z����?b[	�P��g�����%m�����g0�ݡx�� �B��X� �9�w�_��Fݩ�yVR٫�S�h����?&��,���P��/���E 9��<� @\(�pa���ԝύ8@յ�,)Ys����q�"Fx�0Qފ�]�ב�����򜴯:��=���#����T3��b#���W��~z�q��!I�+P�u�|�����gt?�>#�@j�!_%ˁ�., c�rL-�ދ���4���dۘ�'lΰf��˦��	�X�K�m���ѥXv��̪k�*9�5��@�$j����-ݺP�u aȀ;�r{���K,8�1�g��*�m�D.�&w�^1-wa�Sxc*��o��r����릘��͙�%oeW���A$�R�洜��=^અ���{���Z��*��K�%o��{�I��ia����s�j#�p8)�	�c��#X����*�`^����Ee�c���@7<�`�_����!HA軌�#Ǥi�,���=Y�1M�E_�2����<��fa�jI2�}9�*XF�9�����Ck|�=�<qd�Z0��a�"�!q/a��W>n&9���-5���h��~:<4n��I6��;D���sF삫?�l���N�r�8��#�moz���$=UݣP�}R��z�Wۂ�5Cң�@�>�y�/�X�%��U�"������5�t�Q{Ń{�����X��/o����A���U�1�C:]���s��_3��o�� �C��*�,���^��'��-ʵ��X��F����,�Lu �<X���)"�tw�/6�)�PH��g��":\	�]Ķ�B+���|I��3�������C77R�1�w�,�7����%�z���FjM-"�K�={�.���:��d3p&A��4�MC�X@���G��`5��j(7ԧ���p]�����S
�N��O�Y�AOAUGj�(��	 ?}9�>�,����8V,�he�ļ�-�zs-ʷ�@'vt�vj�`?�U���Z쀃rc�F�M��g��F� ��BT�m�XgyG�a��wՂ���*�[<���y7TT�͠w^:@^e�P�3�$��_�Q��mp���MT�A�d�<��O�	���SGy��(�S�*��)(φ��]Ug��Yb���?;r{_f+fкy`��q���?�U���!�?���
�ͽM�g�_� m!���,�˾��l"R��&+�A��q|Q_O.�a�R����	�7
���]�K�A��� l�=r/�r�h5Gq2�~#j6��D�r�s3ƀ��$�o"�UX�۾c��m5z���T��=2�����u��(\�i/:|;P��<��cSB��<�-�2E�K��2�|���+M�Ľ�O�4�?kP��S�\��6WR)!JN2��#O�}��ҵV�̍���'F`��@&
:ꚬjX�Z�Ĩ��(O�"�]�Ui��{>�G�)�M��9����ɌѾ)%�"FG��e��S�;��0��nXd�
�[Z���(��@�gD�I6DM�;NqN#
������.���u'X��`k�";����:;L	t�P��D@�v���%8˙%���G6�V�T
$u{B��R�a��1Fs��o~G�^*1X�X���D��*�C~t�_޸��G~d�s�؀S>J���Q��k	�pv�Т%|�p��D�c���؜���죤I�]��_����㕤��9���'��� ���^p���4,Y�����h'�H�,_��c����{P3��0dI�9?��|~�fc�n��n�>������h"�Dq�[�O��.X����EDj��v��+-�&�.��ܾ٬�/�n/�*�'�s�̡"���cea���[g�u疋���\)�z�k$)��L��_U_�2	5׋���qcJ�pmUW�wC�q�J0Vv]��<�s��J�{b�y:�/�uK�ɖ̣�K�>��9\���]k���
��|��ƬQ��)s]B�����P#�lٌ����Ac�O8�wɌ#^�ڏ��,�G涛󝉍{��0�5�ۄ�[t"�:�i3N�;��ս��g����k|5��g�n|y���n+� ������U�8>bFj�2�&8Z�.����O�Y�itaJ�c��,��׻-�{��a.����¢}�em���ܤ�� �r�qLr}�*�lHC�3���/����t��k�)^���������oD�6��a&l?Z�<?8kkj��^�6���u!A#��B��P4��b�����'�*�IZ���)m�4-�&�)
3���sZ�C���6� ��9!�n�''�Ho��i����	/�?��
����:/Vi>���3~>��*�n�J1Q���
>�gR�mk�ǫ��?��۳s2��8˵�S�t��;f@z�j�6��43A��os�(VWuz�� ��R���w�bO:s� ,��� ���I_��wYd{,�.6���1�����EЯx������n+\����w��.#U��v�"ӛ4X����{�]6��6l`s{��	'+�D��z2�w�p���1����G��Z(����Eva��%t�Μ��.^���9�>��*��Q����������[�i4)i�ty|�{>9�����8Y��@��ѭS��CP��e��� ����%�\�t+ojf��[�B���ོ�3� ��ч��Π%����#�w�}�<�G��.�-<|�l��G�ꦏ�󥡝"�yUE80�GK�yc��9�o�����}�ɧ1S�����A�nڷʃr���C3'�cm9���l�ڷ��좀`rQ�<��c��i�>G�Thod@Űf��0'�I��3�;�����j��*of�Êp���2xLnO�Z3�}�T�B���tb����U�u��
�;P�������Wp��h%��4ljID�E�̖�D�7�Ï5���s�] ��B� ���k��Ǌ���8L7�k�_�x.[*�Lk�4�����<��sx.ڟ`�'"�\Čh�"�`�rD;���Ï[�z�-�Q���N���V��T¸��rs��ˋ����D�5�l�*m�,��� �U"�+v������W+����CH� �40$gw�4CY�YP�7yhaN�u:u�l���/̎�8Y@�8kJ4�q��Qp�ɡm?�C��>ͮ�e��@���i����ٌ��/&fT5�HWJ�E�O�Ze���@���ę���3p5�
$�hM]!����=>����.��mXw�
e���셌��-��F���/�E�0H���:��ݱ��)�ϔY,�ۯ/���5����B"��ʃR����R9&f[�z�ae�$�w	�$�C��i���E���hHp����z���>v�G�ʽDo~ ��c��)O��p�1�b��2�X��0��q���@E�~��w���Ud���0P�Y;�̨�f�@J�oR���[�8w��u�z0��di�<Oy���,��9�� �X��#����A���kl-5���/�:���5_ȴ�k�%��˹���[���/)w]�������/�x#��[��Tm�o����݅�_�%sM%7f)jb��L�d(���/��� 5�)�ja���.�*|�(�����tq���F�4��Va9�˦�D��� h���,3FZE+�lFV��:���H��
�<N����.��L?�u�cD�s_��+�be�@)��2���m,}��q[�t1����%2tl��񂨚��{Ԥ~A�����Z�J0�c���Ťi�4m*������[�x��1qm�q�]�p�H�h�y������<��r��Bx79�ݘ�X����e'�?�ӹ��5�z�H�.�1��~�p�=x����v��c�!MH��V�3�|�\M8t���U����}mnd���v�]��-�ݰZP�赯>�HHJf�E4G���^*ʍ)�f��i?ϛD���$Y��$;��&��݉��w���6޴#1�>��w�1��8�d9d�X��G��\0���:G'a><����=��K��o��}��J�1�p�g]j�l*���C���C��ʝ���݉���*;�qm$!�2�P%!n�=��C�i��#()&���������2$����C;���Ĕ�ݾ͆��'�$"!p	<��=j'�G�I�G�+u���w
�@�BX!O�Yx}��sZ��-p$O��">�뮯z?���.����F�L���U
��Q�	�ϸ�r�c�}|2a׃>F*��)ߜ޶k���g
r�=��F�(P��R����R`{�{R�YgofuL^�E3W��.�{F�~j��=�`eҩ�P��~�ϋ�߸A����S]L�$�ʴח���e��eP���2��h��'�]���z�`M֋�zߴV/&hFM�,*�������L��~��Q�	9�K���(���kq��zD�fN���O_��d�/S�b�Ժ�٠ 9[��-��߯�!�25ܱ���9�;C��@d˔~u�\d��EF�!"�d�T���L�<�ǚ����dȃ���@Cb�q��^Ɏ�2���}H�n��q���1��q�P��Ng������=3����IǗ�ˠ�f�	7Ґ����X=m���.?<���I%�n�i��tڑ<���?�\����<�y2K� �Ӫ9�2���/���a\zH��4B�{"������������̤�j�#.�Չ���ٻɡn��I�W�B}mb=Է�KIه;\ƕ�T4.�ݚ���.�U���E9�(`(�j8Ϛ��G_�&hc:x=Ɏ�8g~(���6�����У���Dxz�A��l���T��� �2�:m/���S�����:�='-hz�t�f�R#p��m�U�	kW��N�舳�)	C���R��� ��X�)��� �8�їl�َ��K�D�9���Xk�;������S��)}�ú�����7`����кL���ؠM�m�������GK��wH�M��?}1!Y��N�U���(7����EaD��dPq�H�.�w��?���Տ�.��)�S�孍�g(-j��@���XE�	ŕ��^�O{`��^�~���t{���uWxL?�*QHA��Ν�Aj3a�uy�y*�2l���7�\�9@c-�zQg�P���[��+k$�*���X��@C���,�p]6��z���5�t��V�k�<A��v�I֪��
��5|��/">rX1 /��Z�ԫY�ë��N�1�Y��s�R0�@п�.3Ki���'b�����)�x�Ҋ��Wз�)��(���X�5N��J��?����y�����d@��h���v��
����$�p	Y�,�;��Hi���BG��pO�Zl���j�4����T���c��Y��V=T(s��u>ۗʎc��}��C�eI;������ 'Z;v�
��]'�nV?�p�fr�ӝ�	�n��z^�mS<���kU�wS��m�����8ƻ��5ԉ�#���Q�B:+6�����K}��-��`���< ���\�C-|1ŋ�T�O��Ud�� �Ϥ&�B7$n�	d���p^9�Z}͑iP�?ҹ�� �VM���:y�����n��X3��Y�>�m"��b�DS����V+��gΠ���T��e(/@c�@&;�J羑�j��>+\F�ٙ�/�3�^��3h�y4�E�5��:n�2�h��t��J~�/�e,6N�]Y	�=�t+u���j�*G��/��3�|�#�K�]��y�-���ܱ���
-ئ�"��Qs��m6|�=�����?>I�ԾFN�#�V��Pu&������E�odD�6��mקw�n'~�o�����{�����44� :��L�vz����xy���Ss�{��%.�qo�����Ŧ�jG��6��S�^��[#K�8/!�4�1V�fw���|�@�T�����h%���e�6� �o�����6
W�oBj�M�h��ڶs,HRQ�"��n������ؽ����z�B/0�-���U�k[E�˭T��* �w%ӧU�]���3���R��Q�7{�%7��N����lM
�űT��A�� o�ѠzI��܉p���S�n ��*�N�F��z9 �O˙�V�j���G����J�{X�G?ʙ6�}+��6�}����8�lr\�e�8'���J ��P��*�_W����B���D�����ʰ{�np��~A��,<�䝂ۓ<vS�r!Чp��$F��*��Хf�X�[9���#� �z��5��B�B�b摾��O�(�D����ţ,��C��wy �e������b�{\[YrJ��Ra�@�f��q�,�D�1��2@�Ņ�l�U�b r�f��ޜ�)�m���@Z�v�P(3>D�
()aX�DAӚ]��+3N����>��:���T�.�\�9�|"!C��L�P�_����"oI��89�Flvg���X����LiW-������N�c�Ƨl�f&V�;Wi'�Кs㰰�5�
�2�e����y%; �uX��E<% (�5�6�8v���:�2�:�Ʋ;��Ș:4c��q��l��}��#:ğ~�?b���`@�**��f��I(w��&�\�rnC�Vb�U���dEKZW|�滯J�ɵ�������0�t?zi��z��y*`�խ�cLP!rA�̢>�{54X9!�ʑї����QH1��M9@����P��z�[w�]�{�cs�K4�r���b�;��E��G���g&"��*��Wo��m�Y}#)�RHi�W̥x][���i��VN����X��,���q�}0d�]�Y��TE���~�������>�/9�n:}���t21u��R��=�bAY#�	�����O���9-I�i����������Z�&���>�
<�#��^��7> �8�	?_�O��Yz�3 shkO�{-�<�Y��GN &��U� S���_�+#��ŻʽKhR0^3n�{OZl�*Y�Y���h�c���nh(F�Zx,XJےD��*�&��qA(��_���	��Ya��j�oH��yc
�ށ��l(��^���*�0�,��@�]ݛ���1��!��8RBifX�09����́���h�#'�&�����oG�
�X���d9X)�"J��1����>��	��7JR�<
-��A��@E��Ͽǹ�IZ?�k�Z�@�Tk��z�:&|�Lڐ~G~��'t�Ç���i6�t )�]x��L)�M����n�6�.d?���eA��=��וv�@,�E�(FC��Xd{�*�I}.�/(v-?��yϑ�nb[r�m��m��J\*J��h�.���(��R������F]`L"'0�2Zx�FԚg�6W�?��Cm�Z�7	Mq�l"f� Kb{S �#f���`mR�r|?f�0>얲IG�Y�Z��*"
�g�ٝ�IX���y~���Wqd�-TeG��o�^�������8�r�B<����MÕ8�g�7kj�;�����K��etO���)|� 㣲��i0��%E6L��.�zZ\�x1qA2<�A�RɔtŰt��elJF�����3��g�Z����,�]�8���"O�7g����,ƕ�ͬ����{K��@9�h���������k���	=hz�d�MN��y�����	����F����K��a�r���>u��D�,��r�x��W��B؝>Y�w���6+�}�����:p�RW\Ҙ��9׬�.?=Z@4����{�����}�.�ll}:������Z���Xu.-����b!d��������AK��(�o5q�ba/@�������^?c%AL~J�
���J�5�a���/�BF���"l�)*`3��U�R�s��X���;�|q��srn��k��Ej�L��6����$1Փ��(K�"!%���_�AK �HNTB���y�Z��-�i���V1"�U�yl�J;�J��mC�E��*�U������k��.��\oX�I�ְ��U��)G�\��Z�k���#]���gƪ���0��(�]_�Y3{d����In猤S��Ë﫯���Pm�� *S��g+�F��� KpP�B��l���bhqf<��iJ��s<�UT�Rt����Tl(F`a%ޚ��Ӛy� �C��`S_L?*����m��G	�oFL���&,>��
����Z��V�A�r;��K9����z׺��m�q�iyg� DLW�,�B�+�r��F��j�I����m eZ�'.��vGF�{@�Wr�X�%ʟ�I�h��չ*C�i������Yv��A�ls>+]E��"�Bf�ψ5���N;�cQ�K��잤�m�$?S}�f/�\<B�I&������J�ÿ !%-�R�_�����ڈ�o%���m#�	��>�ی.�Vu(��Te�_��Јl�4��-zy�Y�D��5*�=�G���@���QFd1`�)Z���o�]B��6�rP�w�=i�$W���`�bR��9�����企}Y��E�x�������f�G�+����O�H�,2ޒ���v���a>��N�{&ݏ9W�̾xҰ�,�����fv���٢��b�Te_ ;{$��2^8og�uY}5h�6�=;�A�3
��D�%\d�W��T���9�[�*�L��M��{=گ�%J������<�I�ME.��P(�A!��w1n� Ai1,���=}�D�hV�{^ �~h�t�����u;�����OL�P[�����aCmYyb�?��S!��OI7���횟@�>TO�҄�^w�mR��[?�Oh
��F�ev����S?8�{���u��?�$PX0d��)@́�ʓ�Y��&2��0�Y��Ӊ�3�L��XɆ٩�n䓴�:.�����H��0E��M���3���P�+r����S}�� �y������;�.��q�'�D��[�{��ȃq,� :0�̗f�������t���(�5z(`��F�kx����Q�P/+{�.��4}$����})iꋸ���(G�&�@�s�{C<9�8��o}Sm�f�W���m�/�<�qY"S����}?%q5��{�A�)�:�T�2V�G������q&���9D�˰�/h��U�/b�����AE%h���:��9�iq���(^6w�JP��|=�Wr��e��r)Ad�ľ��4
B/�u�O�mw��_ީ3���S�;�F�ʊ7��!�.��FB`���j��H1}>�����5��m��l�Y���C̈́�p�h4V#���'q�Z����M�1cM˷\p�钆�yy���1#k�f|�ks�����>,��� �iك���+F�geDY�����q�6)����n/�Gz��`���>��	�%�NlI�C!�VŜ}"��A��w)"yA�:��Fg
�N�?��0�d����?"��j24�_�({"���S��'-Z�¾~ �դɑ��'�1,�w��^�G�ݜw�R���P?��ĔQ��L�2��������D�xV���E,?WA���	�Y:��d���~��j�<��z7����Q�տ���1s�S�‑�����")�ˇ4��',]��)J�O���Ɗ(�b����M��3ꭥ�X�o��E[�e��@�'|��J8E5~��x䍶HS�Y��KKZ[�;>�+}��<����I�.�q�%q��|���'�m
s�o����󣮯���D���I��1@n���k�m��|)b{Lp֐�bm��w����l��r�����#.\ԯ��ТSV>���]v
�ǘC�ɞ�2���U�Cx��'P�T��ʬ�ٯ��G�L]�����0r�����¨.�Hx�����^�؞��A���E���/	uë������@���bЯ��cXc	P�dφn���<�$�֬y#���j�e/��J˭Z�	�����5"�]��G��~M+�h}��^}���E����.�>�,c/^�0�)���	3�О���x������f�(=���^��P��CN�0��n4��O�j��D�S����[����3B��b^z~ �I4A"2�3��N�_��Iy�E&���ϟ�[���РE���׵J6Zl�C��k�i��Op,�?��4�VQ��ْ/��.�<GǮ��/vc֤5yq��]a¢�4�U�e�[n=��������m�r��~J�S�5t�W� ��)ћ {��A��dpQ�v�2���0���|sR�{O\�!�����D(@�L���,�����U�kȕ��E�$ )?����ZnI��
���lq�0��rS+��� ��&�5Z�l��a }L�\0��9�9���e\�@q�>3u���W!�h��嫬HG��|*U�,�����nJ�ӹ|/���H �|q�����ՠ����IbW&"�0���c�Z��\��Jʬ�SX������g-<���J�/���t0�?:w� �gN��9mlu�S���ÆXWܒd�5�Q�MXb b5�_�%>�;����\z�&\vx��5��x7�?����} 7�]@ ������BE����c�Ц�����Q��&c�L��H���Г�x�� �bh�HkRMע�V�H&߷:
�=�!q�T^�]÷
�u� ��<rގ���x�+���.��v��g�1"*]�&9Hɤ�S��J�d����QĠ���!����<ʬ��ĝ�5u�2�_�*g�sX1�u��x����%��zzNdK����=�lxE咳+\�W�<+�t ��=���ʫ!|�,�C�9�~ml��0�?�l���10�:V�M��2�F6_H��A{�4w�Q71Ar�����z,�AUo�t/�F��6��	�$B=��GV�7ߕ���^����#QoS��Ё�f�"�6`�~��3��Ou�h�	�ݚV[�j���-��*����0U	��H���pl6�E�X���c聜֣YI�0I=vս��G ���w��̊,�F@~Y|`$d�~��h�B�e��M�d�ڣuS�G��Hrqr�`�Ѳi�i�qf%�s[����c,3�U�M8�\�l}����;${;���uܦ+���Yp�L�[%��m"P�R4��戰�y�M�1�*N0��#�G(�Z�$�i������C�f����vU���#�J�eOS��p=Q�3�~%t �y��P����>wzK$$V/9U��><�e�L��_�`
�}�&�����,$92,�3��_�ɯl&�Dbx�]k��Q���Gsy����ec�d<���Ln��'v��RN���̈��1,B��,t&J~��s�0r'VQ�Gj���N2�Mn�m\l�?�zJ�`\�����L��"����믯=H��c�`�	��c�Y?<��H�w�LU�*�m9�2\�j��]���C!w�F��=z,���wO�]7H��h�f�a�g�E��Z/�[�\����)�8�Z�;@��2�!zG��-�k]�S�����^���r�%��V��Ws#a���!�!�_Lj�i&il+��AngGn�#��'5 ,I��뵐��+�ݽtN;:H�Ń8��b�ǫ}���'�slX�`
����I���_k��V�  ����`��0��Ǭ	<Fm�m�0_��E�y _M�����؀+(����a���S�T;��$j�bYF�Mi˝��;�5W&v���#�&'��
E�Ы7��'$*��+jE)� *	09�(�w�@e�f���{��帋�+�!�����sZ_�m�G��S׸*xl�P�i�,��6U���Ū�=L�2H>ax0�I�w�U�z�^+��Bي�AJ�-�X�JUJ&�2ۧ��Jd]B���Ă����8Gm^>�(�U�����&��`M����?�Kn�@ڱJw��.�4HS���|�
4�����u{�y@�1��_�=�;���9;w�,�-�͕�Q�\D9�h>�.f4����k;!3�*,�c�Ԃr�pa=�R�P��Q>xL�ít��M3��(��b�`��|e/~������f@?��7�D=����.��M�����GI�/���s��2|@}��zk�+�b�I�}���=O���:��K<��c����:j�ݛ�w���ł t���^0���ķ��rq�ފ��f������˙B�[�L��E�v�.e���W2�FF`M-c:�&��H�z
%����2��&t��o���L�<��n��`�23|�{���г�}�}�������5�"���\�M�Ѡ��݊܊���_Yf�ҿ�����%�Ͱ��Yޞ�
`�2&+�pU|W֍Z-T�A*��k��lc�0���R�dT26���!w8�(h�~Բ\	mB�Tɱx#�>V����u�7	��|��w����y��}���H��̣(����7J�� I&�V�3�,�AE��=n
�N�L��z>M�=��zV�,������v[}<�Q�s4�Bdj�����h�1��4I`61�q��QC0^
��X�4g�*0+I�u�z�$��~��y��K.�e8j��^G�r�dUM�g�f��N7TY�'�~r�dz	A�yd1�a���,��iq4���/P�!��\����ת��	o��]�W��� ��	��o��r�gs� ��Q�?+Zom#��o#8�)��P_�Ϟת�4�M���ļ�3<���v�u��kF3{Gj>�#wbiG�O��ڞ"#���쇅v�OW��S��ig�W��$�N�E�%�m #�.$XZ
)w�����\�t���u2�b�TwCʐ5��D�Y+zɣ����F�3BX�w��X�*�8��t����2�w>N��O�6����ɭ��"��%�;Ca$گd����>� 0�6v:�R"-��r��HT�t��iL_B!�ڮ�d�Z�������{��;�2�=����h���: /���m��	k\��Ew�����.�1©������X��V��?�枇� uu��Y-}�]�u*)ۿ~�x���!k���ރ�K�:Nq�e5�fݎ���m�r(�4ܜx�R>S�LW�%��U����c�����`���Q��ynrs��۔��0��9H���u�?`����jZTrݵP]|�uGR�a/|/BEPK!dPY��#�gu$���àP�fvI�N��K9展�|9B�����
����_�Ud �~E�����RƬ��U��e���9�8�o����_��T�=�z�g��()�/�B�l����2`�	�jfBԬ;�$���H�Q"�~w�?&������+dXQ%�vy,=��^'cMTS(.?�ŗxk�'�a����3:�ª�r2;�!�;���2~��DV�X�����1O�@J���!�Á�f]�:�>;5i�J����娦@.&�͔��N�NQdE��o���ɨ��u_��m_q(�B��jم�f\�;Z8&,6,�32��L;,Ԣ��@��,JN]��q��{��s/s�O4�#��?`�K�"^6�H,ݬ��,h5����41=�K�|���<�z�<�����/�s��!� ��'����=vÒ���πh�R���d�th�n:���@+P�Gϖ�=����Q�7�{Q3w�D�쌦[QW�)���^\�R�͈ Z�B*���ŉ7�^V}�	G�l��ả��a��k�� a�y��ñ*,�Y���A*H&|2���4��~���e>V���� 1�����ƨ]�n�n;{c+OD�#Zh�;��0;�9w���	�j��[���^Ż�m�(��͖=)u-��gSX�k��W��2r�Q������ 2_�p�8�@���=ixo�I��;�L�}u\kko���IW�-?���?FZ��ƶ�9E�M�;	���������M��#�;��QZ�*�)�b��-�2>�gA}a�_��p\ȅ�h\����OZ���� ��Y �qZM;S�C�L�ݡ:���3�R����`�R߼�.���'�	
��,Q���H^�{7��B�ލ3Ц�֢��+�~&�h����J����műfB�S�|)�����`]\3�{nYV�o�Of�=k1���p�����ux���>e֏��!����Z�I/�2�'Ʒ��֙�ɷ又�P�_n�Y�F}�0f��rM��+��l�%QW�]��i�6�VS4	R=����&�
��~�˅�6G����[u(z1Y8O���u<��Ȭ��B#SN[g�箻_�Cn�%�4�Q'T,3��4�Z�mF�[�~Y'�7|������U�Ca�VՃ��;��.���`���=�(pc�IWi��M4@|��d ���L��9��d}���$�.���|b��鷟:<��Ů9�*�g��vٺ HN�~��!�1�œ_�c<vC�I)�H��oT�ń��v�խ�|�Ec���|�;�aI��Ö˶g�� c��&ӺN���a�~��Z�3����>�P�����AF� 4�oH�H�r��P�7�_�	��tߏ�{�`)�4H��� H�q1���
y:����br�>����Gf���i�)LA�ɭQ�:S�KJr�d5X����|��=T\h��sk=�%��[4���
�Ǟ���q�l�t�'Ő��k�r0�1��Z�b[(�N����-qk�!���Yc%2�%c�eHgP���1�=����9Z쩻[�iHv_�7�<;��v�D)���y�����9n�G^��M4wW�sϥ5i�
�	��A�Nކz�"��n�Sr��Y��������RaZ#��Ψk1H��P][i�?m��Tꙧ8{<���(���T�� dyn�S�ԗBr��?�:$�W��J�����B%Fi�g�p�A�'HN��͟�ܺj3na(/5�j�����X�W�L?+	�j��	�caS�_�?����<�1�g牡j�Y��F�+�Kr�+��ӏί��F��Υ�c���nm#K�|�A�o�CN��559��r�<�흺�S��K��h�<̩���i��;��1�0|<I-�&:|��*� 1	[��^͜�xʿ޵�� \�fHv���GB$�Z�\�� ]�>�
�ex֖�w��Am��ڰC���%�5��'9ws���H��ٹ����_��W�,5vw�'گ{}W���Rt�bS����[z4ۦ�P��1j�d	���t�=,.j�.� ��ƅތ[�1N�})$��t�Q��@9�!SGWJD,�JM�a����i�U/����΀������j�?����8V�6����>m��+<�E��S���N�ƫ���������O��zx�=r�ʄ�}#��E�Q��&7v
��2���"�W���%�;�8�'ܧ_�>��mӬ:���,����g����դcgZ��q��a���UG������dx"J�|�X��Lp��&�1]UXtaTd��<.���$n��L.��?a��(e���Gƫw/͠ZS��B5�,ẻO͊4;��k��:�J�R�n�6��̜J[�d	)<͊��/4`�!4�]���5M||>�����r=�����$r�zE_(Ĵp���E�5 F���Iƻ��sc<��\�"��,��ĝ`��Z���#�u|�b�������@�`v1W$ 9��I�0#�9��'TmN+y'!3�w�G�i3�K��9a�m����s�nA��)ֺ��r��p�'��x�f�kN����i��:�  �����o��i6�b��k����o�#��c&*ت��%���v��|���	���O�0�LjC���d�`�|<Q�.�6"F�j!��r9�$\��_
��K�-Z�=��4>ι�`U��u�V�é���?��6���|�� Q>� =I�%�NĄ��J������i������ e��,��� ��X���I����9hR�ƴx�02q3��)��̓�gYH���
�=@�3_ ���xv�<��$fK�{�6��i�.���`c���7S�G-�WU��F+Ψ���{v4!;2��PH���?)$�I��c�7�'#�2Xs4G��KfI��� !r}eo���5O5 ��]7�!)(��B�Տ7!�l]cw����|X�� ���(*�IG� X�N~[�1(����$�C�̊�b�]ZC�xO�$2H_��mto�P�]k,�$4�.3�����"��סsf�E+*��}���j 8�L���/�x���*/X�J��~�q�x'�*���Xs�� ���%z�C�!�̅����R^wa_m�f��0�5T�e���>F�����io�%�%B6��Ρ�;)�:�`�6R�0���T��r��I��6û�c�R��d�l�]+?"��Sَ�G��S�d|�!	�c��[K9N�`�ĭ��<"̩��� &�<�V=AT[���n�*����x���p� /ٜ��p��L13��OkN7�:��)�+������v��Mɬ�o[Ps��*� � .�AG�A�(s)5w��A�v�o��
Q��Z{�%Դ��a�������	k�8�ǩ�(�~��ZM�d��Z8�Sc��9�;Q�E�K���^Ub$:̀�������7�m.n>n��鞟)�l�t�Q~B"��F+��o:\�d��ɤR7�%�y��,�w�<]h��*/1-���+�Y�+�FMffߢ��\��v��`Q�L�"�h=�V2�p�~U�8̋�em��N��'F˱�,|g#oAD�<\3Q����Q^�'��mcc����<�o�Y�>LS[�Ncկl�)�#��2ID@��ݪK��4���N$���gU8X}�_ȏ�n\1�� �A,���I3�-��Kb굆�gKg49�lw>��PZ=��a�9�n���(���*'�!,�)�7L�Σy~k2*�9�Y]`���"Q�z#N��QGB�%xV!�id�p���G�a�� P'Da��.�2�8j���t������9y|�'�^G1O���;��˸�����dmc�9eK�X��P'�!��h���9��(M�Y�"��W珲NԦ�@�3B��d�a�=s��Eh��
N��E9�t����& l벢lސb��S2� >��ү���$��I=
��(���CȁQ�*H�n�����X94<!��f��X�XÞC�\�s�Y���I+e0������Ȭ��s@�3�51��D��s�-�̻]
ߕ��fׯ�!�;��6�'��9۹[��8ɏ:�D#��X����G��5�֢�y��������9�0���=�慘[x-�`�˅��t(���?l����|�m��:L����1V!�[��+	�'c)q�kcY;�/P���I���n���L�b���|3z�_��B��u���!�x}�B:�Â��*�������q��G����9�>�n���z�HWR��0�oLU[^�L���c
������t�l	�?J4i@�ya�8r5���e|eA�f>���.���#����xu��M�oj_Ț�U�DN��naϩ�aB�I�ie8�\��G
W#~(�c� D�>I�ZIks�4�
{�*O�6��lV����6�F���f��������?^�'B��� Pna�.�����ؒ�ތ�q3�1{��2G|2۴��R�q5G}8޵,���&-��+�;~ �[Գ��{���k�����O,���u�<
q�%�K>`=i8D�h*�B�S�%�:�AA;��c�i�9���b9�3V, E�ؼ��=k��o�2�CW2��5Y�J�q]�Ok9e�>F������yLWr�;�^^�c���G%xH}2"
���\�XT����_ bs4�gm?x�fՠ�M��N����X����0����d�:�ƶo+��F蔡ц��VR��,mG�'5�����êeD�㶮wO^(�r�����`��O��I|g���/����a{E�Y)�q��-K��1�(`���	����S�!�{T��]>\}��w�g�*���߲�%O�9*��R]�~*��=�ț0~y�)!آY�4U_�g4x�Ĩ[I�,g�3Q��?�����r�a�`6|�]�d�JcH�5E�cV�����;׍h���w|����S����y�+m�W���ŤS{��NM4#n���?gυ��C����LJ>G:%��!�x�N\�: A��%{�����"�J���ځ{�C�&�a_;�Bb�9�J�+\ސz'�_Kc�h3j*���N�:w�N���٠�����wr/�����]H/�b��^�h�%�_3�Z�G)m�V��>z�r:��s&A�wm�ZiZ^�	��?��]���甆R����#��q���u�cp����-r�Lf��~Р��#i(gܤ`0�4��Bg��o̜�x5ְ��r|(���ގ�{#�"�9�ʹ/�5�O�t�:[������	3Y6�73�ԓ���za&c��gG���e����Wk#	B��C�lN㯿)� o�
+�o,�^�-��>�0�����6� 7��?�
���
y�g����Y��U��u�*��E��4���sx�v�,&�����>�=��>�I{B�#�����P�B	K����ss*����8�*��2f/kϰ�v����w���[��_h��t�h�Ɂ���j�@��کh���xE��{�G�>�J���3Ҁ�;�a��<�(�H�X�jY��5�JԴ�� y�"4�װ4gGH�%��Q��8qk:�0Pv+�;�XD�n�� ���?��v�>fu���W��#��R�E�6 �B��
�j�΍n:�ə��2u�	4@ӂM��p:�M����m��� ᲊ�2�ԼP��&E����3񞧡��r,���H��j0<��K�{�����.
��ځ�����nlw�}p�>~܍���)1��Ğ0��\��?�؉�I�����P�SX5�4��ŇD��P5YL{�3:T�S��� ղR�T���/v����j�i��D{F���kJX��O��O�T Y v�9Hɔ*�8kӺ;�ǚv����n�T<Y�A5l�+�70��j�L�"@;n��������`�lN�è_��u1-zMi>�Ѳ��Ͱ#��O\�@�3v����t�Cfh���!��'�h�h�+0��MQ7���o'^�������et��`�Sھ����&���WdI`w�r	bYEq�����2�1u���:�Uk�s_�C��L*�"���_/d�C�N���l]�����c
�[[82�}`�őm+͈f�g�j��+ED*L2s��rD&��K�:����D���ޗIkb�	: 3%	��A%e��<�]s�rV���A�YH9U
����G��]�ɗ�C� j˩7t��ĵp��I���,C�[�u���l�iS��w'6��_~̝��&�ŭ��\�a!��-S;]��7Q���v�C�n���V1ϻ���ƣzGR�je��R�����Q-U�Q ?�*��A�< &�~lz��}g����|wg��,�i�Mc�����b��	9���M�p���ӌW��G��n�(��RZ7�L�웛|EԄ��=6�s��\�on������w����l�?�.<��GҷA]�X��:�r�j>��/֌\�)�pW��ϋ��d�`��K�s9�v��4u���d2�ᬸo|)@-���s�޻X�ж^�h7��k���H�in�4g��anJS�=1/5u����VR��3[�Z5a W����i�9ܠs)\ą��<B"�*��� ��`L�1G�彉1 Qu�WY'q%SƗnG���k@s��g=V&���!��}� t1�5��P���icB
e���o�R���Aޅ���%$8�ͧ��.�.��	"�+)wk�*�6���8l�;�8�E�_ڱOr���W���ŀk��:j�'�fl1t�)�k�˛�{;��,�Kj/���C�4O�:y,{!5��_�j}��);*��̴|AT��qd�H����t�5��\�"w���4��)0Ycκ�`7�#�����fg�&�R����8���3Z�wH��֙\J�g}�����
��0������l��w�!���E
wrj��jyA6��-��Zt�l' W3��J�3�3���E<�{�i_�&$�H�`�>:Y��V�����|���@u;��[���%�kw^���Wv�uA?�[t�ډ:X�
��">�(���d9\Ot7�&j<��{�V��������=o0�|J�f(i'<K ��]�#yC��;�b}��2����P��7w���
�U���1�ˬ�
�OX�7��
�[i-z������63��T[/.�N_7�sEyS��u�U���|.S���n�'�n��
����+#x�s]b���YkՕc;	3�]R`�S��rC!�.����_NC��@B)���Ǵ.)9U��X���xp���9�(rmj�~X�)�b�����F�l��y��͐�fqK0�%|�fz\�Z�K��q4y���qvJ˩B�Mh�8����RT�з郭�_�|��Z�R�9�o�õ�A��m�՚8x����_�,�\7pv�D�/S�����)]!���0��I<�
�"�r��P���z�Aa�d^����J��|�^�XJ� AUj��EZ6s4�{ <xZ7�7�}����F8�����A\�]�~���WK��t�s� ��6�B7+��~�YYΌP�gg�B�I;�� ��e�!�s��@[�1�hA���Uۨ���<�p�v��k�j�0�=Ɂ�P p�� ���3����U�tRͬHB�}۵z���|!wIM��ѐ�/��{���મ�=[7��`)ܾ��"��Q��D¦�}ltx�t��������D���l�z]kz���H%kp94�����0(���!+�oH*�E�����
u�َ3<<��h�Q
�)!�yOPNk9���ɂ4:��W��������v���<X�E���RW[* QeY�62W���ȁ���j7���$�3�H��fTdByW�2�w2�]P��C�p#/��T���;'Q���Q6��1�w��Z��`���X����Lp�t�`�w:3��
��N,� ��	h�k@����>|\
��6J̈́�r]'�����2D����u\-�2(���sB������g��R9�_v��i�;4�}Iu�dȾ	+K��*Q�I�T������ȚP5V4bP=��f91l �e)��/Ipٻ��	���q$��!�{Eס_�����U�hSD�Beڏ���CyC3������V��l��/¯��ׄ���nQ��s!8o�@U�+�9Z�:��ő���ѝ"�-�A�'=���[V'C�E�̫%X�W�";�l:��q�)���n�.�z�ؓ���Q>�z�(��#V(�q��T���p�>��
�}�I/�^�ϝ��~�VJ"ꫠ����|�"K0��ف��ЭcS�,s|��4���H�-�¹@>�)k��{�$F_�J��L�DX���j���D��F�ANnd�6�l�گ�E��������U��5F	�-��RI]3�"�L&�"]H˶Æ���˼;��=�äu���L�wr��I-��������iv�3��k��Yq���%�l���#,g�B�o��m��4���q��*
�)�l�)p�q�oKi��<�9���2=�{t�ĕ��HZg�i�i�����V�$��qD�
E�ۥzSJ`����GD�PI��b�� �fGtJ�
_�f��ِ�ڞ��R}6���v=`�u�>� 7-���	F�o���|R�~K�S����Waۢ ����MP�H�h����m�Rn��çq�d�Ff�xh%U�mR�2���.�役�dΊ��� �Yx)�T��a3%��|g�$� j�.��:KV �9��{�����5K'��הo��Bw�������&�$j�d{�1Z��Wf�dT�}lO��&Վ}�'�ijKTŸ�[�;���!.nU�̀2 �Ti���x�����Z43/�ˀ��#�p&||MF�+�k�8�E�6����ȡ�^R��X!���=(&�������+���W���]ʛ�b� ��Q��D�������R�����z�y�z!�g2�T_��ۢY
&��P4��&�J澙K��P���4�:��BS��d׆��t����x�����L�i,��_�	v��F��^�44��SJ�'!.Z��5o�Yv6U�5��P��J����Z�w��<H�qP�=���^]�� �0y�C�����ͮrx��TP�yr N�Iƥ�Qx#�7!imr:S�'}��O(��	��荖��kLC�����m�ϼul��HB�=!&�>rW����QJF�;�C>�]{�� I��RYd�5�JB������3�q�E�V�8)Ч�Ҫ���L��G�UM٤��c��=�>�M��rmiY�e��/a�f)������F
�k�/ŵ��:{�[pl���2�Y*:��$^�D�VbbǧnW?_��/���3�x��ϒ$�f�MQ�W(�ۀ� ߖ�j�TŢ�W4*��/�r���w\�M�3��L;^��)����=��4t���8W��¥"Ȳ�M�6�Z�����>�%��I�:V~�&�#!�j�X[+�T��T������%B]�P}�ey��(�s�طх����矢��؃����>����˪{��ٝ
dM��>�b�����b�q Fl��3|�iV{�l�l��ͼ����<��2ԍ^�*uҡ�8�@C�LCw���庝Ĩ�2��IT��ٽo+��*3�&���8��1�i���S\H}�K��Kd2t>el��3ф��ɔ���Ay*�x;?���v����9!/]94m��;Y�df��{��}*�;(�=���E��σ�{�Vu=���L.�����`���9�n���EW>���}�����;��˦и�L���Ͳ���-�7$"�8H2\��_�����`P�ʏ����0�H�+N�f���T%�Y�o�+�]F���5��+|RD�b`сZי�����cv U��|cU�c�ág$h��wEPǷ��ԓ��`;��T�/{/�^�9���z��^��޾�e�T4_��7��L.Bc�Z���'+����X��69m��H�z�i�~�1阵�������K�m���=ֽ� /fVK1+ҞW��tNZ�~8�;A��7�v�S�d���ݝd*�2��'/�r:*0D��P속�M$��3٥��>�y�놌+G��9W��Ir-����hj�1�����X�'�`��v��r�s;�
)$�Uzf4�'<�3v�Q:�[hÑ`�m��Z7�@�Uo�{��|T`1Ht� م����>8�c��$ީ���
�
��_��H9��h�C�v{8j[��90�ną8x���V��7�Sf���`��5q9K�j� �dk��̍�R!C	}�� ��F�݀u5H����[���fqCkЫb�avFlgG/�7�3q^>�r��X�k���b��OIw\����|+����0�du�=�hD0kQ���z��y���;��� ��%�DY
0���z��̒��}�'��=�|<���b@��#h�矛O4��S0?���)��OAg�~����M#�����m�eK��E;��H';��{0�rL0�"
O��M�vAm�1$\&˵c�
�+����J���A����j >���$JP���M�
���P��6'�T�k�o��qv\��W�`�a�ٳ��q:�p��,�K��9$�g��S��B#�9�TT�ָ�fB﷕\:�4x�W07U��ț	�*yI�GC=���Ǩ������e�&n<��*	�U����b� ��w�qSy$f���	�v�`�%ˉc���h �G�p���Iu3
'��_�-{F��Sp7��uP*�M�Lw�ӢSu��_ʦ7ϺZ�P�˖�WF�`�T�a��=e���:����*I ���I�v܀��'G��zk���wW?��l4]���E2P��j�f�kwiO(�f��0ԏ]�{T������aG0D�y項��PUח�=]Pq����!8I�j�u���:�d�:���NOa�c��e��VH8��o4.I�q���@L�(�͘J�Ṡ���"e�q%ڹjFߨzΐ\��:h�H=�����RC3�5ˠߜ��ܡ��cq�1er�2��Yõ�ڦ��x��N�-?R{��h.'�h)��F3e��d[����z�̀Y��9>� �F2!��6��|�4�Lt��/?m&U*�dY�{y*����@��V�}|�Q�l���#s��\KVG��ak9�h�3���%�_q=�������P��\ˢ�gR/����as��~!�� ^��z~R��v���NT�a�@d�v�A�as�{�	���!ыe2͔5{�=�P�z䧦���7��#҆u�����Ggu�\��r�"F��I��S����M������.���O��Ǽ� ���:�w��*�ɐCă��v�>D&(�V��@L.͖��3+���R��Y)!�uf��vv{�T����:12A~����O��H��Wi�6Ѯ5^LCCd7�������5�6��)��v~\&8���$a���$���A[��cspj"s��ص��+>a~3�.�0�IP��{}�f��Y7�G1Z|�Fz�SsFCD��G��MN�4 �b���s�(���ï_U�S�%�3,ߗ0.₮\e��uK�yVʀ!O(�����|ǹc���a�p|�ꐼ�oL�VJ�?ú���BL�M@����o&�L7��&�@�1�;;״Ü� �1�a�S)��d;�����x�v��l@��Dv�g�{��v�o�>��