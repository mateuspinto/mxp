XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F���濾��XV��];�J��6��(Ra��p�q�`8SnH���8a�����($Ce���_�Ch�<\�������J��-�:���#����� .��*M3��4Q"��:���]n�%4��d��z/�ԮN}:J��g��A��s�f�泴�Vl�+���l�"D�r�P��m�������%[=tGȪ7Q-7�/�+]������D�B�]�Z�\I���|RP��>� �����+[�����f�(6�������nw���ܮ*ѐ�gT�s�s�����-�z��T��VT� ��+��Z����3Q�a��h�s[j�Ѳ�$	� �xX3�+ �����E>_3Qh{5�>~*?��	�D:*5��+�c�uCTW�O�d�g�6##�L#<���8$7�Ɠ�s��NZ.�ͺ'�"��H3q�2p�;��b\��>n�Ӽ}���n��5�j����f����~4�0����]��Lh��K*B��F�X0��mH�:�@N�;���ƒ�?J����2l�ߓuVҦ�K[fs��^M�&G<�UM�����	�w�Ѡ{l�9s򂂰�H�	��E?6����"���!eѡ�D�ńY��Fs��#WI?�5�/�xkYp�sG~Ϳ�ˑ�N��PY��R��횅*S���v!:P�V�kI׸���~Fۘ��{O�V|�P=n���O>Њ���ṅ7�ڎC)P@,�A�w�EvbH����>�O��fء������Ʊ�'qXlxVHYEB     400     1c0[��6���!~��N0���v�l#˶��)�b~Aܖ�=C�!d1��11�8$�����0Ϥe\nD�n����1iN��.ϰ���1�8��3Hy�WZ�|��P��nAŕ
Wh"����_��X������C{� ��L�f`g���>�2:�̿�x/@	]��:I��vyK�LE'_ƀ?&E��ڧ$��o�{�K5^�n����Ҫ^=�c����7q���,�=��р3�
�s�\RF
�ed�^�5��^��R�����%<��+広���UG�GS�ޔ3�nLհ��Ǡ��i�]��?d6.0�p�Қ��fXk6��8�u�
|@�R��y%��5����G�S��W�s���G���Ɯ����k:���f]����5���f�������ڝ�j����G#���l&.�Ơ�e�,�,�̖�dXlxVHYEB     212      d0�Qr�����m��H�)vV�>����A���}���	��#,߂�/'6EF_�﹓��
����3h��S��f��ǉk�GE���O�Z����"]��s*(�S��0��h�#8���d9�H�5��.#�3��VN)�F���Y�}����#U�_��IBX+�$�S��?ۨ�W(k�K<ȋ��}S{FA�#��fE���o8R���<�iir�