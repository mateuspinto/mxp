��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����ǎf�@�}͚�|ET��xW�(����2u�y_�5�ɘʪܼ*�\w��c3&�c�zP���^��G!N7�1p�H��AK����s@To}��]�#U��Σ�$�w�*��F�c�Wf��/�5��Ca��b1��[��b����Ad�|R#�O9B��̓�5�+l�f��b�to��q��x�V$8�����={�P���ڷ&�i�K?pI���w&_��TL����;�O�w�pQ��.� �Z��� V��jK��9��N綷+��[a�C��S�2�?�܋�0�=���΁v�S��+���mz�/A"�v ��-K#P8�}O�]	�H�f	�?ʞP���up|����?��ıN*N��/s��$��w�"NY�N)�.�W?uJ)���Οyշ���%� �	�����ZK�
q�y�dC���=���8��>k���g�
�*|���!}��T�%��Dx���P9:�]#�j�	�9/�ǝƼ#¨���}��Z&0����ۤ]orG2%�"�R+��qU�q�(���/�7a,���i�2����+H	�4ɹ.�E<�ɉ��m��P.�`����z�b�L �O�"}u6�^xe�S!����.
#�jkXՀbYC����$�eH���jz%va|������k����S�聇�tNĵ������؋�A�v@��@��1^"�}�xf
	��3`1B�]����"]��&�����ki����ΤuvU��`>�C�KO�$�� �ӂ>��
�nG�E0�.�t�؜K�h,�	?B�Ix���ƴ�7i�M�Qe�Ekˠ� ��H��!�X~&��LFm��%�~��7I��pv��u���񸙟r!�HCJ��8t���om�J=T
�l����]���pq|��UE``h��.�w9���b�{s��t?����ϱoX���O"����G�����_By�I(�}�����:B5�5wR_w�uua��NÖ�w��w�1�u*���O(ɞ�8�,~8�q�I9�M�5v1� �#�-\:���yҟ�8���D�t�`D)��"�
�2FM�>.73[��L�	��*�}p-V�-�������h��ن��/5�?�#=�vFZ���fv��������f��m�и�9���VE'Ì�O_�9��S���2uȒ��࿷M����+-�-K����^��D��Cn�=�&�@�~�f�Y�@F#R �l �H?~���T�
��xՔm�A1搎��>[��4r��LT^��μ�~ 9a��q&RK.xg�ڟ���Z��Z塿�~�T�g��L��bM��+����}�rPC���7�䗀_vL��T�������e�D.f=q�bZ9�<q���x����<8���s#�@7�M�L�a���b�R�����M�[7$.ʉ�js�e�`)Z��թ=�v���N��/�Y!�}�4$�� CI��jj�S&OD-6�������%`����+Ddc?#�y�|{1��� �q���7���V_�����?I!
�L�aGP
�� e�W��zw��.��à�)��ԟ��T>�[�M���2?f���z�Dħ����o΢@��e�|셀f�y�"c�"l��.�\�~C��Rrq'TG	V8��^؛j�ER�9T�z�7�d�o��z�,ope�>��:E��f�2f͉�-q�X���8��_��OQ�1� /.��̧y4Ο�~@I�3=�q,�kЮe��MY���B�q�P�_I�|cs�;!"136�g�0��LlҐ�D�ִ�ݝ�q"UN�$�n�&�^��dg����u��0�8|3�t��|���d�����V��&.nj�)��s���!K���O�e��B}֤5ё��z��)J�>�K/�*��ѭ��_��kT0M@�(1�
Q�Q�T�S���l�I'/(EӘ�$��	=�N��f��)E��Lr�^��%^�@�@	'��G��6�#Z2��Y�3�q�}�; �%t�-ߏQ��Ί���ӁE<�b���TҺ+����\�>��8(��"��'��ez��^�m��D��<��k��
�3���PΙ!��6;��j����
�+�,�!G��by�N"�	�
#1e�M�b��Dȵc��t XTG��+e��[�vy�%K��q�dj{�HC��6ixG._����hd���#c���y����	����5�>h��L���{��ŝ�ݝ�W��`�h��(�L�����jFx�`DSv��\V����s��3����U��׹	�w� �d@w#l��	
�?/��d��QɈ��SS����E�J��0xz?��i�>%�'֌V���~�\BZ�D&]a��l�w��9���S�j9̡嗯�T�h7�����o���vω4� �/{��}��>S�$�wS�щF�wւ�Aݙ���@��C0��(Y�[>�{$/W�Ĩ.닾Y���l��6�eƧY���0({���̌0#kvl��fyc�:�F$>=<s]��yO>I�����៸��;^����� ����%�df>S�y@�ܒ�ڗ)����J�����:?]tTq6��;/�]'�C���y����<���׾jdbċ?+��1�(�2hw���$����9�k �-���	u$���4!X�vGJݖ�C��oI���	˅odے��fn ;D�,#��]��4�UK�*SF�����
V�Z�='t�v�PGŁI1Uwex�1�q��ov6u��
g�� `&X4:�,��|����Ҡ�ԉ\�����ۥQi�=�8��MfX�;?��?�d }ѓ���.���y��.�)7Z(�ܰJd���D�84@l�VČ�d�;�TƦ �{/ܦJֶ�Tl~'Ƽ:�T� 炙���8�Ě���K,���-�_k�
MSXF���1�w����g��k�qt¬b?�"���
!�����G��:�N����e1ghD���5�����t�ƧE���I�=��W����J a���@�?�Db7h�AQ��ҎU�4�8�������L�IDq���K�P�a\Q�}�`�H��~j��D���%��W���R�j$]��b�<�m�4>�)�k�-�ۨ�k�E_��'3�����/Q*�^y�j���Z��
�S�~��˯m�u�f��#���Y��	僪-�;vc���Tdj�{Ru�]W���	C���z=�̥;w�LFgP�S�kG3��<;��F
���˨Կͻo�g&���!�Z���JS�8�ܰ@�P�+?(��	>.��J9|��}3�ݟ���M��9�|�}�JcR�����	繊�U}b��!�+BP\54J�{��~�9�5����v�-t�Q�Iװ���w�z��T�#��,R�i�����%e�� ���1��Y[�\�ـ�N+1��5����li��g���_��X{ǂ�spU�<]�ܘ�k�Aq�sK��=���I���O�L�h��0���0s�;>�%m�6a`~9�D��R�G�	�mD������@P��-93C����1]r8<L.L��^x>�r:��zP���TK�C?��CiW�^�v���EtDtAF� ������p'獌�/R����{�}a��w���WI����O�g��ϝP1�O__�a�/��;�ws~��x�e�����G�xQ��:+q��	���0Խ��˂�9�Do��Z5��I1�Ad0��Nk6��Y��*��io�� ����3���ћL��ۂ��f��0�(׷�5f�޺���w)�Y��`�V�Ȱ\̍+g`��3���ѹ������w�����gdu����wwX+�˚�7�
�Zd2Z�[\�Q��Lّ4�ɽ��BX*�*Y8���=T�H���,(lė���7���#��ye{j?q� 6ES$�U��a7�!}�c�����Vt�����u찋|�G|A3���'�`��O�W�:WD!��]��V�iu�'P�Œ|ηS�a���
������Ai:��P�������|r��P�̐�˙����22C��j��5�/l���M�Ǐ�>��fVl��	�ރ47N�z	w��j�&�rħ�ױNTo��j� ���Z7]���v�'��p�����>���E�N��Q�xd���*�*BR'� ۏ�G���� ԋQ?��Z��x'gYyz��J�2F o�d�ۘ6a�`p��B�T�����/*��%s��"F�8��7wa�4%2/��<�����qJ|���
��c�[5G�p>���.���B�ty�h�'�v���E��;ho�K�}Q��U���`%��4��r��U��[��L%��(��z!-P�9�qJ{'M@/����I� �gh��L٫eP�IeW���.����J��7jEg�Ӝ�D�(�x��?�1���fPC�~�J���.�V����H\l��������Ts?�������M}j����<%�u�~7�A~�H����}�*�'i+�xh���l,s��A���TN��%��ĉ�6�4n�-��ʲ�FR6�I�w'�?s*�ةm�K�<�:]Q6�_��d���!�u�%A�?T�vNR٤�${�!����
Q�n��f�I��hj"���}����W�
Ձ�Ob8�&��Q؏r�g�B���@�a��yց���'�vV�'7����PظC�H�J�;Q�<��id��(��4�ܷ����}*t�XXUp��/���� VjI{��=�J!��2d�Ќշ�ƕ�B^c���R��e�,�/9����6j��1�Y��*�T ��n怃�]���7r>�8�؃?E�.6䰵�3} yLMy@�%ɷ^|�!$'�������He���2�����_�޻��~PZ,��<3x}���+�Mga���j:�O��J�kW_t�N�`%=(�2��h��+�_�6/��@d����4�0�Xj�H�Rs� v��۾��Ιi݁��.�u+/ڢ�5��]�)�����J���ܬ�/,,��Х��:�Ȝy�.
DJ7Y1��0:ҷ?F����_�)��N������x'��e��zp�%h���q�&g��?_�|4��z	B�����@ԁW%E�����6���f�ד�-O�_W ��J8�69b��lpG$�	�C
i/z��z�
~Vc�nb�/��Y9���;�䇨���I~�<�gP����Btx��܀&t��� D<=ː�~o�#Jla�J��O �#��"@nG@%�#b�k�u]1GvQ�c�	�`�-���!ς���r��F+�ߝs�������d���J��*,�vPk&-:n�mg�����e���P�
g���t^�Hu�~�P���c��7]Vf��y�b�]�lQҐ����z�\�[�u��YqN&����1D{%,���k`����T���6��K�Z��T@*��5�_�'�D���3Xu{�K��>�8W,�-C������6�q�����ꢐNE.�i��b"���_�-���\��3�.��B����ĘLԪ��&ڄ�U)�Ȫ�$N���Ɵ�T���l�O&7msxyE���si����\npR���F�,�sNO$˖�,b8;��}C�Y�(��}{F2,�B|<�̉믽�3��Ѱ�%U�) )`�C�Tj0�6F�ąxU'�u��s,����U�n�Cq��	&�Őo�f&B�����ߠ7BT��x�[(S~й�T'�H͔��s����wɶOE�~���ٯl��2�F���H�%L��*0�gȞ���W	\K��WG�Εh&V,Ɍ�ڹ�.��L��0��2] �js��)3�σ�6~�,�W=�ǟ`�X+��r\=�ϻ�j��4ڵ�G����7�:�m�pT����7�B��@�O�oC����2��S��\[�np{��ߚ��%��|VZ�j������*��R48���P�G";Xv�#�����I����5�����)�cӟ s�����}�QYO�t���@b���X������ھ7��ndI{�S&.y��"�:id��YD��]� ���� ����Z������ab�y!/����aqR~� 5j�9��Љl�����;�i��vN�M�&{�B��6���tv�ߴ��g� ʇ��Χo
�-z
�-_��|q��%@��]�R� NF7$�BX-bزI�x�Z�Љ�I��$S���<o$Lobx�o���(�мv.�-g���b�<t-:ȶP�كl~\�<�����4Aki8�������/w���;`�U�,��׃%_��&=y�N���t�	�_ޮ�K�J���?Fu���iJ����rL������͊V�g��2 ���z��8,y���Gq,�zs}��.uD)��L������Y.w�=��ג�9ā���.iaRtA��)	�G��H{�� i�d�ɬ��nO�R�h���֭;�� �F�&_-���Ը�ȳ{Y�$�%H;���Y�C���|��wS�14��Ė���{Lk�c�
�dؼ�:.�5�=1��Ѩ��up8�$=��Ń|OY���o-�X|�Nda��(20��n�$�*9��\a��k���Դk����{��Rd�kQ��Q	O7�5Etˣwo2���'tp*ժ�vV!���Uy8����he�*��V����[xA
>�>4�LD�!�Tc�d�x�Ȱ�;�,/⦀ƅ�D7Y�)E������ߞ�Q��M5��r��AP>S����$L�S�yJ�|���h��e�P���?�'�6�>F���ڿu���}��hG��CK�Uߏ9iG��Y�|^�鳈��	SP��;Η��'�(�qRx�q3W��$g���U.�9�b��c���=�S�ty���&>(_��x�v���HK���W�
9�FI�h��U��@J�?���fΦn�����i�B��Y�3���m�6���ξ�scܰI,�K|r�t�E(��rj2L�)�U��o�Q�r�lli�b~S^�U����_�S��7�0(�����e�H����u�Sh	�G���jiϤ�)��_nڿ���W:I�3p�m Nĝ��������cvN�S|}%4��1 G8[g�A5k�R��9�W�6P^iΌ+�oU�P�c�{*1�_0 %�'d��/D����P��q����⭈/�h@K�8^ޮ��n��r|<�Cl3m��c6�1���������3�+/���� ���
�4����81S��MF��¦��?#�)�?]A2,�sG��C 8��	fb����e���ǎ���]�˔rw&GZ+���D�$"i��
�Կ�N�3�o��1�QQbnb8��¼�J�l 4ɟ$���G�V9��������[��V4�I��e��a�EL���+!�i*Y]�=fC�@U�)�n�<k��f��r<�&�A�9�&��90�m9fo�qaJ��S��5�U�F��̽`�|o�:y:��M��R��Ĳ]z�L�8�Qw ���׭��]�!X��+䁁G�.���� ��ن�RδI(�O�5���7KR�}�!���Ɔ�&�����u<a����d�ME�/`W�_�;(� "Poc������<��B�p�.8]��~��M��]ݩB�?�0����sKiM�5�ַ
��8���	�:!� 0AVO~sLoP���eP�*�/߹�N2��,�0����: ����v`�U6��p�ZO����+�聾ؙ�a�ߥ�_Q�M*\����Jt�C3��[���3��
�{�bЬy|*�� XC�%(*gU��;�]��>�@�C�n#tl=�+��T]�KUu�p^Ѓ��ݧ�k�L��=�-92B	Z/�ppn�zY�^C�\I��9�S��~ױ��z��������J��]�����"L��ʒ����D�v�*�~��S�/�{��o>�K��l��A6��վ��'L��le�v+�r{HY�;A�fLk,N�a=C1����${��=JS��o+������8���Ҕ�a�S�/��Oej�'��N�R��'q��9��pJeo��d� ad���L��A]ih���F�-�n��yxJ�%Օú��Χ�Q-�޺g����TtS���_R��A�����������R�N�����]H�����Y�.Ճ=uB��0aڮ�t��dkb���kw��)�:}�V����l~���a`��!�.�Xse6Q䲐=��M�������.�}Ʈ����'<�v#�
��3�.�ο7?i���	��;���학��)$iv�t<�ǘ{��
�@�-X�  �6��Q��f��^�d���z�-!���
���*y)���yvZK�c�$s�jj���x���3��5���.�#�O�A	��`f��\g�����I�	w���� _��R|������jy��xLT�A�wv��u�@��(�y�J���u��G�|��������ha�I�	� ��Tb ��(*ihZ<;���ky�D��2�ք�[�.�"CO��MMX�]�>���޿��o��lC~B|�g��g᮹�vq���c�-�Q�7�P!�\I�)��u$i���n'��8��@�X|����������i=�Ҧ�YJ)8[絬5KN��#�����˟f]�z��¶ߖ���b	��%��h!��8�K�m���^+��n����q�sk���Xӧ���_���l�K��X8�ak��J�
�^T�_{`�*���Y�lLq]=xl���/���&u�A'�ۚ�`z�C�e���^�ۗ��Ǌ�[���.�c�Pa�C�5)ijN[=����-��.�v��I������u])�t�ٜ��w#�큪"\^��B�9����h�>���uMP'�5}e�W�t�<Τ<��;5/�T��8�T��s�=�W�i=�7v�C�3G�:++���?�$ ���:S2F�=|���N�v$.��6�2��0�����b=�%��Jz�8.,��<���N�Rk��jM���ZPb�mY%��7M�Z'<��������d�o"��5�	��{G6슋>Q�@h�%@ӽ�;/.���g��٬��0i�GxPk��u'���u{��9�6�if*M�o����[(0�yj��X֩)�;�.bC<�-@+ն��Ȳɴ�$����k��R����Vw`����A��e�	T��
��#���S�Yn.��0��܏�����$��t�����L!�Y+K���p
�)� ���r����MELԴ��<�^ *1���)n�x6��z�l�/�q*���W{=�݄��ԙ͑mk�����Ή�YT����7+
�+bS�����A E��~�C�d���R�v�o�#�}мR�}wytn��n��e��s6��]�ࡖ�]xɆ=U� ���n&�@M̑Dsl�t?*#���c�A�O�%�\II�z��Q���V4x�c�K�<Y���F�9��8Oo�k�kL#��]��������z��3c4jU����YS{�ŋ|f��_"ѫgj����/:�Ā粘5��!��	M���k�	q���.�W�����`}¦�l��W��Ol�j��u�ıK��Ӓ���[�}?+�lk��8��2[�~ɮ�'{3�(��`�2V���P"R��-�6~���l�M�T1�����2�~f���#�L�)�5E��������)�}IR��=E��\�N�x�������ӈ��$�Mv��!���n����3���}�q8���Z�m�˪2m�RP���_��U�7j0Z����P�@�7����=� Ƿ�i+�Hi�ͤZ���L� 5�F�m0�c�i*vu?�Y�V��"x�&g,5�H^� �,:���_N�'d�h�4����,HgkM+�����/Hf8D�����A���r���1(��H����]]̽OV�'���q5��>�!��L��_�+�:��%F�r�2��k�`Y�^���ˇ��~��X�[��nX�(���SL�e�����׺�N1��>��)X9]S��[�cs9 ���_)�v�����g���vC�09g�T�,� |Y�~)^�P�8��s������XrD��� ���-�"�ԣ�W�g/;����3�8Nԭ�ߡT������ԙK{p�"�L��ٙ1V�g�z #���Ps?%�=G�0|B��������fX�Љ�o�K�k�± i��m{'Bl),�)�����F�C���(�b�?��a���=P'0�!�D#��x��A$Rw��[�6'�k��x�e�Z�h����G��qh` �}���EZ^lH񚵄���V&�Z���X���z[#�����.��6�t|�.B�:��'��0�SF�ы���?�)��R"T�-77�;�D^�'���mCU�@���;�)��������c�="8d0TW��_������ͺ�q܄0��2۾�rK�!��aӋ�D�;���g�>{PAh9��CyM�G������5ϔ�ܸD���!��&y4�{��6�`"�H��+����8�=�
#XG[������H�B�B�ߐ;zҪ���v�#��:�����7p�,}��h r���̛� +�ژ�����V�D��7���w��6����8i����O?W:Yb�*}A6C�L!��o3�Z����n���ҩH4�Gv`_�,q(v[��"��$���l`�i7M�DY&_��P����g��RC�#v�o�m��\b�� �l]�jW6��y,?brܐ�N'��UJn�A��)!)�6�kw�W�/�$J�i|�x�9��Q��l��dR��:J��0�?��i��ޕ�2o����T����ۥ/Z�)GmiZ�P��K����u�w��'�7z����tu�-W�@�$W��-������m�;�ɟP��ɟ.�J�1!�;�8�k��5�WP;YC��"s��"�R������n���(����ƭ��T�*[����9�Y�+z��!�|�ե��tО�[����5S���ifM���
%��=׌~�T܉V<��Zr�52L|���al'�`�H���M���sVh��_���x�&�S�&��&�~�L ��L�x�k��޴�+�-�r�s��5�� �/���I^M5!'�=-�t�V�TL�>-w���i/�M�n�^���jK����E�qf��fL-�?в�=c+#��B��K�G�� �ԋp�b@�veP�*)ku�2Y�ު�^�e�#���C�Uv��?�g�L����'��*��1���^t#�;f\��������T(.^�(���XS�3���	WRA�)����26�dE�[a��R4��]?��&ٟ�!s�?�U����*^