XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����9��rp $�:��cu�����t�Y�c�,��?J���{��i���KQ�bW�l����궶<��m7�}-�wG_d�����]m8ű���:Z�
 ���#<Ǌ����!�.���	o>s����Q����#����Iz��":r �f�ljd3�ya2�Q=�;׈���⇡r��#�O��_ӊx��d��9| aa�C߻����K�8*�	ld��q�;�<��W.ryq[,M|zǴ,̦�x��`��y <�v	Ƒ�<^b�c9u��ކ��6v94�j�#O�8rK�&?:)�6�����f����̫u ('�}°0tt.�mPI�������\u�>@c�I7|L�sD�Y�������sb{�sz_���"S-YoƲE��91���=�bE\���?�>,|��*�Vb�����UI,:�D*�^�7EO�2i�o*es��"�&�Đ=�Ң媐9�j��L�3�;���
zF�ε��Im9Ϩ���{G���E0��l���Mʾ^��,{�p�7wÕL��v�G���( 3��p<[6uJ���ZE+�r���7����^\5�K��KM�F���qN��q��zf�t*���2kFj���������qa��Cv�*���� ���˪�e�����xM�1�g"`'���+����Sn�
κ��ǙҏL�7�<YuƸx�dJ&���E��px��ڻk�O� �1�Tv��4����&����JW�h���?�)4�lR�HA��NU�U��^��.TP�uXlxVHYEB     400     190��`��Q"ԣ���/Z�J � b4�����4�V3�d��?|���eH��/G�,h>��/���z�O���9K�n�J����k49��2#>�v$�%)�KVē��HK��¶rnM�W�ƂZ���k��	�>tn�c�������ߦY_�I��-��s�F�|��T��0����i0p�CVp��>Z��/�A�.bD�1Gg6�}䌖�W�6ǧ����%�(7��{]�YZK���,��5ҷW�gw���!�t)2�o���q�"R ��ҨC��u2���Θ�H�n(w�0��R��`�oʥ3����,M��.es�w����|�m�$i���T��~����nY����b��}��$��t�ٗ��EBVݼ93X}�D1I7�F���XlxVHYEB     400     140��Z=ܷi�9�@>2����?<��w-����Z"d��7����SUȤ�ֆ����O8W��	n�QTRiJ�D�N��^b�'��D�O����K�Ŵ.OJOEp�UB��,�
u:���}n����D�GR��$V����T;'����6u������h�`og���k^�	
E;�W�[ �|��X�ͧ��>����}!=��}��X%��V�C�q���>%_
+�������U#X���Qq���q�e�H�'2X,��t(^Zl����h���\1��\�ԩ�V���{��P���J�J�*��E����XlxVHYEB     400     130O�>����س�an�s����q\�
tu��,KvvZ��2tX)i˺d��,���u��rVh[�,�gk����� ]O������g& �5
I�+l���l��� �;�\�
�x�Q��D1�(�J_ٻ��~�=��1:؃�˙��x�K��T�e'��X����M�7a��Z���⣙	�\n��RmǨ���Mbҧx:^$߼S�8�*��nG,��yQ�;W���^i7Z��P·�5ԵY��h>U��1$$Zg��z�W�ht����Ut1Oѻ@���t�3|�(����;�]y=����H�P���XlxVHYEB     231     110�g�i��]ѭ��X�{�R�㽡R���i��ul�sb���8��A�.�]���ޙ�����ڒx�#R�D�g��W+D��dj����[���Sv��'�F�X�Q�U�d��s���l ���]����h�1hnK��/|��P��,���Q~�A�q`���<4����k�i��Y&j):$�qz��ʾ�,u@qFuJdO8��lZMǗ��u�����$ٗ��{�Z����q��$��f���uDg�/&2�w��	x�0:�"G��rʽ