XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���*?�F����s,?��h��/~�BZӡ�!�d��,A-�Q������Yp�� D�1�Ɲ����n#�8�<#�quch>F�e�#e	(ɩ%bgm֥Ǯc���������@{^{��%��r��c7d0��fu�]�jŌ(��`��zO,FtO�_�J��|����q2Q�3����z����D���ϖ=V�P�9�紂�3ܨF����>x;4W:f��8p�7V2�@�(�,��|G�Oib0+e�sѹ=��3��`�0�-��:9�m֐�,� W�!(���gx4��ƇL[����I+�Z�X$��T�
Q��@�QI�*�m�F����V�!��܎	�]i���� ��Uຎ[P���<�B�e�V�f��RN��ԡ@��F�ч�R�]za�m[�EdIgY�1p�GH��Cp,58А7�:���%$KFy
e�{��-/��Gvo�5]�/�JR9�.�^�v������-��DeDcΪ�e+���b�ya#�����qv�|zQF��=� ltyd$�=���s����w��et�ڦ��:"��� ��i�ujV�.rn�6����;�%i�#�7�y�� xE���I�,,x^�.�i=[�S�O��aV���)��h́�aoں��A�s�ʚ���.\��@�-.l�_��"�1���	�2��s	=%>aV����,prn��2��r��	�����C���p�{0���M�e@���������k�4hs*�A۷3�3���P������0n�TrXlxVHYEB     400     1b0��kG@ĤQŴ%�3����Q4�WK������S��� �n�5ວ���E�t](U �KZ�[�4g��r�.��d��TX��0�	9���2KK�<�뮽��ZKɼ��j,d=�zS�!��uC�g5n��	?�ǩ������y5uGR&l%�t��Tȝ��Xj��;�RQL[�2
��Z�A��	"RQ:\Z��������7�Ϊ�M殦
�V�Ӻ]�����1U��%�bM�������&��@��t�R��d�W^�%��^Y����������=� &`�{�CCR� ��_�v�+oىi�Z�hL�a����hi�Eoi;���F�P=��'�g}���U��|vL�^0�L� w<��W+��V&��m�Z��j�<h���8!{�Vq\!K��K[i;�[�H�[F�|S��o�xU�r���}VݍXlxVHYEB     400     130��uso�����J�Ӣt�>m`f�>����i�2(S�zl$,�w90a�I�G�;��Ʋiw�J3Y��n��/�Ɵ�	=�ۏ�������v2����R�ӣ�=��f�\�9��Z�K`���cQ}��YZ�L�J���*��1�f�?T$�3"����f�i}���?�	��5�S�(0(q{��yJI���c�����W���2<[2�����^^(U���xh����,�}�4(���F~�!���F+�e3b�b����"!�4~t��l+�/��9��I�w>i*ED���d�W�+�XlxVHYEB     400     120q#� ����I�ҽ�X�j�Ù�l�CPb{��gg��s|�n}�[�@�0*��|�d;��YV6Ɖ'����/�F�
�~��7#O`=R���ڨmX�����5$8�G��� t�������h@�'�z�֔$��p�V=V���+�[~����a"M������=���/2��������f�w�m�M���-"%!PEA����C��k,�(��cV�X�69o�m���'"��ϖ�8�h���%���"Sk2Lh������ҧ��<�jYh=�AW^�XlxVHYEB     400     170�E��eo��Ξ�����O6�d�Gb���J�]N��@��?���`�5�%b��^���0�gWrg�U�y`g��aOS"R�����!�f��s�b�f���ZGK�ݸ#�Ȓu����8&�zR��� ����F`��NG~�,�@r�Nk���z�Rt�u��*�"�T��H��*���E���ΌD<[O��-N��*���~�#ou)�e\��iy��5�v<u��p?�,�D�/��Fͮ"�7e�^N��w�>�&������ު�5$�r��Nz�i*à�6C��RH��e����z������_/���NC��/O/Aoc����KJ0��|�|x�̕n�`���>�XlxVHYEB     400     1c0(�[힢�����6f�rku���u�Q��^b����x�d�r�Ћ�
���E�{�]xkR����ZD�<ZY�Y�HO�-b��:ZTĶ�ec���y��a-,_���h��[v	l�p7����_C���`��h����8K�w̌\�끼�}��dRe�
�%-2�<N&o0ɖyzk�f����7{��x2�7�P𗭂ū�oK��̗qX�4���Kw��@~keD�*�U�	�7��t��� �G�E��G�d]a����
�}���e��J�H�j�TO^^=$��Ud~D�^������/���eƘ�{ .���Z�01�S��!�<��q�������I��tq����ɐa��]h��V�He�3�-���:��Z=��~5���*gjy��ҝ��!̛��v~Ia��pX$-����p6�}L�0%=��y�旒ɟr�XlxVHYEB     400     170�922�g��5<�D+�j�͌�;)�^�+��,��X�e�0�d�9G��ʐ�.��2�Ո�9Kf�;$̾w���%��Sqڹ	��.�/��NO�/~=�Bb�UU���ΞV����a���̵#x�k���b�C9�Jk��?`����D�ǘ��r^4E���w�2�LO�H
�҅3IL��$gB_"^I�/��D��"uʥ��f�jYE��iG���z��OR����Q�"d�Qm�N�e����2��UI����¹��(���V~�h>�+9!��R ���EQ��L�@4���ѹ�Ք�:l��$��Ԓm��'Ǯ�B�_��	ɮZ�Cf��Jg۩�]�n�iȹmJBJ�XlxVHYEB      5a      50��V�����c� �s����
�@K�Ш^�i�c���~҂hs՝�u�%�x�t!6��yDɬ��
���|K$p�