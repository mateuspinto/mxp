��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���g�"u��L�k��	R�&N�Gc�݈�
f��U���i�<����Q�j�eb�ttt���y�lo�?V�-U�W��(h+����z���=h�*i�g�CS�bXpc�M�Y�x�Q-��{|�u�� &����5��wHmaU!�%SP>��YA��tZ�wQ���>-�Z^*?���*�;��^/ÅA�`��98��ܪ�Y�K#���/�y��y-o>��A�~��j�d��ΦT-�"(=�U�?{���)'���kP�5rI�6�,�y6�H���`�='ٜN�&j�B���a}jQ!K��|8>�Z�]���0p/�ąiB*���^5&RHG��mj\�o3|��k�'��,��4�[d�2z��+j�M���=-
�m���D�	���������J.��'P�i�-���=�z﷊�i��!4�A1��k�-�AU �I��`1�y}�+H`0.3 A!dH���b	R�����GI���?W$n�3ͥF���� ^��=^Y�_��m��a�ɤ�73h�[>8�������h/��wFJ#���W؅ݯ6rbRR	��CߐK*�-1=T#����v��3g�yC��������B��<G��9G&A��\;��mE�ʖ>~�y�PFZ�i�f�~
�iL�52���+�,>~�^iX�j���G�%s�b,�˟���Lk��=z�g�/�Tv�,z�l���ߎ������v�;,>?GtF�v� �9o�S�����d��n0nv�G;�{O~XH�6�&oh��1�i 0��|#f���#��	�E��_�l_�'4�]��a�C����E��T[�x\�h��f�֠Z:1�] e�8�.�zV�!�&3[�����H��i ������vp&�L�󷞫�Z��I{���1v�K�+�x���wTos�K�{��D������$p���[�O�������������ut�<Vs�N��9�6�D0�e n����*L�d;�����6��kBaT�o�3�L����Χ�Xx<>��{6`j�y9s=�`�v�|Ck�[���t�����O�|�4��:����O/]��I� 'ʁ��s�4���s�Ŕ�!!�9j=�ѥ0=�j+ ��P����:�OHb�}�l��ִ���4�A��l�	�+|�P��;5��6�.��P�K��V����CD��"DqW��rF��MN%Q��W�t�N��k�LC������f׎����5�{����^d��6��v`�"�wt��g�e�Ƹ<]}BCr����>��ɿo[�o��D�0q��/��7��b����Z����xm�ivmv"E��<V7�?��ۓ�D����'�>Q�`|˳9� � l�Cw��u� ��.	T���/T�,I��Q��(a�<ȩ�.�@P=p�Y���:(u�����BlA�T�_f#�^�0مRV�ԛ��6Kw9*VTle�c�7�*�h��7�����?���"�Ϩ�ˏJ�����P��a㈳���E���9��ά_r�`7�����o�cxHBqmr�����g��E���n8�!5�;�T��[WS���^c��m�3�>���Z ����oN��n���T];�����4s�(�BEQ!��aN0R	^c�Ŕ�d3e�d��yӔ�+8���ŒH�,9D�Į��?��E�}����|�B�.F͌zr����[��$������<���s����a���(��gg���_tW���v�8S8ޅh����D�o��	uJ���C����kf=_�������)WU;tp*J��t2�?�� �-�A�~ِ�R�q��ΖΉfq[�Es�z0Fu�F9�/a�h-�����Z��߳�h�?�`�i�l�������v6���"���Gw��D��Q��س��d�;%I#6B���E���2d�7��V�N�J�Z�	[4�B�m��L��-��a@mo�H������vn��2��#5lT��1��_g�?�'*��S<2xs�l�[󻒽���G:�B���7��g�Bx<���j��AܰMy��L,Г"�/�b6P��y����+�?����t�sZ��|��G<��\ֿ����g֣���E=zE-d�*�_�'�k-�ߐ,�EX���d*���B!��.������5����8��x=����i�o#�(ţ���Q>�ꊣ�R�Q;/�*�X�,����ς/�_����*�ts�0F9����a�a�� �K20�ɠ82�.����i��yw0a8�&��(�K��AC�P^RK@I�̔���V8N�}!J�	�	�YҢ�c�"�ĲQ/K�H�0]�i���|D���	�;o�'���@�i��û�`Mq��3
����"@���j��ZP�.���绮0@3?ؤ��)�P�vˎB�lL��l�<Z�� f�Pط�l�������ʏх�Cx[��2��£8�k��)��PDX�-�C�"�*G<,�9v���N��ߡNy��3bu�� ���cVd���y*��IFtϒx�}�:o���_�EH�OC��tl��uA�
A�L�D���6p3r�I�Y� �<�^�����a;yz�Rw	����A���1���(��+���n/!*����*�T+m,���)I��3�߈2��
xm^��rU�j�]#:��Gx4�"�O���ZEo�r�9�,��qI���t���x��||#ƃ� KF�+��J����p�0�Al���|°t $�:�0y#���xe�����*��5�>�+Ŕ`��z�R?ʋ0����o�=8�G�*S��zټ?�eh�H�c��"2:fU��sp��l�A�k�ݩ�5prEP�EVg�6���
���;'�7���qg��Z�.��P�EZ]��������qG���饳�#�fU���v��K�%���@$��ڬ2{-A��{1�A��X_�X1)��2vAl	�I�+�R['��{��9�_�W����쁘�v�1�,x=�o��`PxHI���_�ѱ�M��^����x\�&f;=�|<U��:b�b9���'�t�m��ظ�w�R��Tӏ#ĄN�RB���$�v1S��R���~z3��Q��wj��Lnj�����W�.c��*M����ca]sG"`����	��ea��U�Uf�	K�}I�g�����G��S=�z��ӓ(`��s#��lr�R����}#���Y���E��ѥ�>���+�;�r��U v�~�Mщ��@���	±��_�[����	�[5��� �L�˝/����)K�]�l)K �"�#��U�C7����:_�(dN̝���W|�EUD]���2v(!L�4n�G#�d�\3dj�xRq(}�x�� ��rz�������EX��J��3&��>��\5� �XQf}*���m4�w2ڧ�i���W�oڊ��VO��?��T�ë	<?��YZ{<9����		4��R�73ն{�R�$|�KC�An$&Q�Y0K+RzLz�ܠ�Ww����@S�D6��=���_3	��j��x4x�孢
�y��O�K;���j�D��"�����n�_nvRr N�R
ȇj'��1�pa�Їi8���ݑIvv��<�q�򵉸�� ��l��Db�a��)]�l�_䎽�M/����z�Y��k��.8��$��W�i��V\C	j5�(b���̝��ն �u�v̀��pG���1m78��!���ʵy�u�tB��7oK��2"?-?n+����`�T�r3=�OoB+��:l�MO�w�b?DSۿo�fc�p3�Qn9�-ڂNK�t�mO@M+ߦȒ���\�F�ű��4K8QC����^Z��8�Ul�*���gE��y͌���B�vAm[����2C̚���(ݛFZ�o=�GS�C.�M�і�����1��Be�����<���]$��~o�I��;x�6̑�z��Z�/����mKe�$x��-jn)��Q�J\$����rz\׹�hw;�yUG�)��Ƚp�:�m���j�w(Y����bi�J��r�z�ʈ�Z�j����	Ҝ���	;��y��+Ӡ���=T*M<���|64ړ����GW �2^ ~'/%
�w��P��������B��gWczu����Ԝ�n13ۮ��A#?��E�4���PV�<��c���(�6�zq�\�]�y�C[����K�ro�@��p�Yo�ϲN<���&���̈�>	Z��q]=OH�&��Tm_���P�'tW�?Z-K��>�{&��*�\��B.�.h�^8'�&%w�c�ǨrI	C<1�[^ oLDN	6�wl� ~�۳�j����*��<��hyY����C�/:	4E:�)a��(:[��:����Y�����jO��&�֨��2� �ږL�X�4k+)#v�B\䍊�A&k���7����A�Df.�Տ�� �Eo(8�=R��P&ڹ޿�"wi�k�"41�H�S�轱j���9�_%D����� �ʪ9{&X�����ĺ�*,:��FiU�-D�l2�c���q7��W�[�>���!�{��߲�4�F3��=dh.�v��� ��rL�k��o�I����i�[@����e���S�R�!+٦�
$O���u�ϑ�=T��~'����{S�jsFQ�3pvp�\��7���W��@�p�ɇ�E3�%�"�k��LFU�N����RR¾{Ȓ��|��:���-Ơ|���jT��hPJqh�Ȍ6��������?����v�r��
�j��%~h�����nɚQ7���#���V�A����rfL�����-�>��O"�ٗ��쁢�v/�sK��Y���٩�Q�> 3�w:"����8����J������T#3�-w8�Y<80�흺�pBA�K"g���t�k ٫�M!�B�Eg���uܱ��1�_M����9(�9بH����Ϧz�o�\�K t
yn�Y؈#��a����ɢ�*Maz�7�\�%K�u.Q�2 	ay�Ψq�`�U�	���[�L�,*� �t��O>��	�*�`��n��+�N�l���]���.\K����;��ľ��@��/��k�~`R��$C��f��V���6�0C�Yg�,
p��A���11���S{x��"��n]i���OCX+�d�����l���&����\���N���+G
ؽo�Ls�Ԇ���ʈ|��4r��1�ۇ�x�ԓg�٧{�����i��k��k�����b0��A4�b��N5��x�25 ��f���g&�%�|��O��f�+U��h�Y�*^��q�v-�.av�'g:{>x�[�^�����0
F��M7�tb��_��0B�ZH���qgCџ�\%`�_�;����{F>���I �	����J��
x�(��`M������я�ޞz��1�|Â?5��ߩ��>1u�Z�iq��zW[IH�w4Qq��/�~����Wr�i�1k�CT���O�ma�]I�M���~,�=��a���gO��Xq�r�r�S�6c6N�:�>�-�,=z�0i�)D�Xs�vʆR�kk"��E���ҁ�v�*o��"U�����վ�A��a��Z�P��5!�w�Z��Ej�M���ZEW_��H�e*�lKl*\�\$�ggeKJ��_��%�dl�'SP*��Y�|X9����w�J*�8�J湧��8zJ~;*�WZ^�YǱ�!B��?�PU��ӹI+�U��,5�0v�ӌ����b�0���\��ѻ���A�Wżf;!�2.:/|���z[�p��&b�?Բ`
� ]��P����~9�	��Ѯ-��ir|�rS��avcg0z�l#9���xx�zаA��J�1�_����enH�� �U\�a'�JkL鼷���+�nT�S[�R
�����t^,����?���^M��}+l�6r�M�8��.�Ӂ��$�#\���a���ɗRn�zM�v�������$�m�Ot����*/Ӂ�z�#�,@=˖O0[E�o�:k��ط�4���zZ�Y�>pZ!����0�
X�E��1�,^�<P�D�<(���r�vr/��G�pz�1*S���Z���[vR7���i�PmN+!��G2dcAk�Ӌy�TC�M����!8`�q'��אk���ȿa��z,!d��E�5U��/������k��H:e�Ґ��8����_�<��i<�oZ�o+�����[�8�'kx�o��>,N�UJr)��B����̐n�gg�������s�SG�@_�.@S�h�-���⹰f��x�bv�p���k4��n�IJ����/�,�i{淖���u�ѩk�b3�����<��$�,%s�ݙ�Ma�͉�8t!��\�'5	t�q�=Ś�	ΓFN�ܵ��M[K��""����:����ɗ��vI9�̛�+ٜ0@�KӪ�H�`�S=H�'J�"J�8�[�V�&9Uj�r�9XX!6{�Lc���҅^���<Z��'ݤ�����d���ƞ��nd���/���l�ӑ�u������	����\p�?�8�����%�V�F���v�-�v$ʻ�����@����I;4a�"�v�&��+b6�c��M�)���,��#�.��7c�/�D55������v�l���S_x���e�P��y�~19��_���%U�U�g;��$��=)�F��EDzɍ�����(��JwT���}ӑ)4��ə��z=�p�`fZ�h̿�j@{^ڄ�b�[(�mOU�=#0�`�1$'�>4h1yRK��9�� B�Cᢳ|��F�81��pL�rAhc�tN�'�qcGC�T���=�(���br�2��*~?/������CÔ
c��qd�pˌi�X��:��� {��7/�B�\�oEEe�J(��D��Q��S��	�%�W�4x��ι��9mRթ�&:�X]�OW�G!�{��'�G��6�߼�{n�%�G$�X.W���ߍ�_��_�8��X���!��e"��ђX�U�5��ṳ���v^j�$��ma.n![]�n�;���]y�s���X/貌��-Ɏ%�)����`s<�:�;D;��)ݎq��K&�p�D���P�i/�Dz�]�/��!~���{�=�/�3T��f�x1z���h9���Y��r>l�Gc?����=;h��V[��=��r�Y����Wh?/.�$�a`nP���_?:�(|dF��{'�q�ո!�2���;�*��TǑǩ9�W���F.�q����x�?%J@�/m��xT8�q�ϣ�3�r�m��82v1E�h!��G�s轫�L=�^E�e��{����2�J@�����ذб|����@�,0Z���^� ؼ��<�Rz�rԋ�]Ȓ(�6Ԁ[\>Y�I�aoX7�	��]x���1԰����l���"��H�r�cz%#�s"���]rv:K�?F;><Y��.���D(_���}9�c79��`�!���,��}Rn`��·l��]�B�ʬlױ�Jq{�$e*��5�r�Ck���`K�9۩�!���5��'�ԧ �l]�j��a)�i��	�Y������`��)4���x�������U9�nf�� n��icjMX�f\�����#�,t����Z��[.'��o:5G�Cm���պk\!p��^g�%�o�܆|����qP��v��׋o�ı�2_�\d4�cI
 cw�`'C�p�C��]�>s=I���������Y3���a����� �~�����Zt+�r2��u,÷A�Z䱘v�A��p���H}�[��4o����M�?q��گ�]YF/����إ��\Y�L�D����;�_�1А��YqPs������6A�᛺�̉S�T͹Sm@�<�e����+R�\(����G�f�rB���m����m$�Wk~�B,��	o�.�`�d����F��2"J����Oha����N�#��y�ֳ��/����U�}�9��D����#��g�D�|E��O��}j�����0��$��\\�m����	WY<�1�s��x��y��*�r���ϭ�oK+��t�''��Ȏnl�b�0���%@XC�ɴ�)�4x�A��h"��?�3«a���c�T�i/U�$��T��o��Ai,�n��l��d�"W�?&~����)�`���&�*���c)�#�.��Fqh��9���D#�~����tʢ��KK�s���|��7	�F��sk��kc�7+��نT��i��Qg�;��7bS͏9�6��Ӛ�\�G��+T�i↜q<Xw�r��r�B��4q5��w=��ܻ7\?7�FD��Q����qS����G7wμ�btg˞Lo3��������kh2f�^�vuOФ����d�M��Y� �G�4ͥ�.a�O�}X�R�iB�C���:u���atá����r�?k3���a�6h^h��(k��M��s��mO���=��ƐK"o��#4ܶ��/���ȵd�.)-ŋ]�i�}e�5�Z����i/�l����o+����ݦ��s��PP��jsD����n8E��#bK,�m�]Q����=���Yr�諃�j�p�ȥF��NKkG�#���,oǃa6j�;�'��;۲���Q9��$ۥ�P[��D�S�{d�.�!�F�����vjS�fp�r>D�%LC#�I����`T�9:��^s��|����	��@,�#X<�s\�ӯI�1��P;���?�hW��X�e)׉����fO�Dy�
���v��8G;QXg?.xs�J$�rdY�
3`�'$˖gT&q`�9�7
�:4�ÓKnN)�o+���|� -N&�r�Mx�����>���6x5U�Tfັ�:	Z�Y��e�-�r����x�kY�S�����	�7.�E~�[_�1$D���/C�l2�˽ʃ��8���'j8W� ��@G��r�o���z;�\��PE~$��)�f��[X]���|�Z�+ ��J���Y�n��_2�T<�f?(�hF�O ^ >h��aҎ1'�*�������[o�u���I��4[��L M����቗�TL-8�+�w1�����M4B]�R�yI���W��i�y��%�� 9$��/�sMG��{4�o�x��s �v���r�ń��o������n��4/P��6v�*�r�Ӫ�u�4��1��\����i���ד�#���A�'��]?�Nl���5����=���9�բ�QZ����D^����p-������fgm*�c`�íV��]|�8�1�C����ң�"WH�,��i�B֗;�2�~�1�:���E8�fj�b�����*:�ޗ��T��|�� �o7�-� \��:w��J�^M�u��o��]��:��W,.ݎX'f3m��<.��Ch���$�)��a<�2����AW:\�L���c��/�[�O�XlGD�K,�/=��
�����$Nb�^�l�pM:�����V)0u��
 'rnq���yRUqj�M�~(olr��692�E��[Q M�#�V7�u�_����&M��Nז��yռlW���RZ^�4�����+F�]J�n��W�?o��������yK��M�)��s��lUM�=��*�0�k�.@h�H#�=��g���l��d��z\�g,ҳ  ��@�>�J�$i)U��_c�ހ"EH�|��e��t;r_֙��cV�˸�Nݺ�g/��]���ʉ=��˵�=/4��.�v[����s$�X�Դ��Ð+�mw�x?\n��+����;�"����w+���A��1-���;��g�X��Q��A�]�//ņ4��~6��:�"xZC�I=��	�e<��w G���9cY�\�z��+�k2�r�ڭi�ѳ�/V����ZݠϤ���J�h��?)��-�:�C0�ufOJ'�٤�1�+M�gw M8�"�h0�.I��_�@�Jl+\�쨠=`ْ���`U���C�.oΫ�������q>Q4eX�zJ���q�(�"��a-*����:�8Q�������A}�k�x���I�^daȯJtҳ���YjLL�=�;�P������Ӽ¥��3nKѶ"���?�`"���k��aE���%~�8�gS�ִ�v�ѠH�܌�@%�� 0��"s��,�_��U����-L�<빞��J6옩�e1��&�A���۫*��Y�wM���y���jXx�	y�,a����tra2�[|�׏�GT��w�61$
�Z_J�,�WO�7:��'�,��b0��`�^�}�J1j���'h9��s���lP�q���^�jS��K�@�]��?<��Y���?�y�o�����c0>z�r�!�ݷj��s���!� !Ռ���ρƫP�o�Q;��VmC��V0�f!4uq�no���p�#�㒻* v D�j�3�C��4L{�[�o�G��|��߸\*
�2k���K{�������N�Db�ח����h3�ű��b�@_0����C��>�P ���;��#�f��hk�@��s�lD�[Y]!u"����]c,�0��8/�jC��U�*R��H������~:����l�2��٦�'����0Vqx�b���D�۱���6�K]ă��b���3�Ov6�4��p-%{�%���kbZ�d Ǭ-Ѹt!�B�17'���6�M')��e�<F�E�9�4�f���n�Ɓ��ll�[:^�u_f�S���Q m8����	�3����u�5�sR�e��x��QR�:L�\>�s���v��2t�n�8^�R��]���z�UnW����%��8�_]�����F%���">�+�0�R�(�it<h��d�Gt��e�ZNT�� ����+��TQTX){ōk����~���):����e�M>h��\˲� |́@דk
j�a��G�@ٸQ�85�;�M���yYw=+��Ҩ�?2Q-&*�ĸS=.��E/^���,A��o0��Q��	��;_x�#�0�}�̊���i�f7|)�#<7��ȼ-iU������|����ȹn��-M���̹B�*���}tN:(�����䨓�?tS�2T˶edǅ����U��ﲏ��M]��#��%da��xb�Hh�me����\�6�?�iy��\�ԫEE �����4�̰o7�ڎˉ��f5���Ģ58n:nW��5�� KqA�n�kXG�k��� �X1M�1��,�����k�.��.^��'����O��tnmv&�Z�Gash����	j���괇�����k8u�����
K�u�7���Sbs��H0���0�M?<U �oed���f�rxr �m�<���q?q��p�cgH-��(5�'�J�D��j����&E��m��j�*4I
Ts[����H�C��,=����ݠ
�c���O*��CՉ&����8+H2��b%I�
N��O �~A1��x��!��έ�m��;�$����"��3�ӟ0R���\Pj6��0��f$AB[��*���;��㍜i�Wt��W���<!�f�:���M�.E�p�J��Sߛ]�G ����� ��r�o�ȡ�U,,f����*���s	pcK�-epfȾ��!"5�n|-y������5�i�k!ƥb�I�,�9��� <���aί��+���\�i%��Ξ*6�Ź4���0��'��Jy+��Tč����i�Ѥ^>ˏ���
Y�E���-��j���Q���s���` ���'�Hq'�F{t�^]-���c�I�Ȅ8�����ɯ��5ȀZ�K�Q��1�q���:����E�����ܐ9�{�c�F�F���C]���ˤ�:8�y6����X@C�_056�jE�/*�.�1���
�iv����,�kOY`ީ�ug�VM���"�)KZ� �ib:���|��ߓ�ڃ��=hV�[F��y���u|b(u���R�D�h���`ᗂh�G���>S	W��C)F���ˇ�H#D~
���#��� ���(�$3"��;03Hy�Tl&u�h��Ou�2���\���}O��y��Q��ZW��s�T�얫klh��Wk��UNe�'��*z�kR��H(�*�P0/�%��tJߥQk��,ѱ�)�w�.��w�d �D��Ub�е����`E_\%$!��~ހ�OZ&��q>���v�?i5����V;$zv�-�V
�u[ћ/���	O[�cw��R�ā�V�t3�<�ef2�x�\������!�V�;�[�����@J\�)+�D���G�̶\����Ok�`i�U5Vz>�W�t>��$,m(��*��2������J���X/�Ճ;��C�   �U$�n�ںS[\i��ڣ�!`As+W������qK3*�'��e�G����v����Y�����i�B ��PF<�ly���I	TG�G��k#�XS�c����p�jo�6�~�#�v�1n�;�paX����ʒ�UQ��>���pb/A���9���T�e#fO��&�(��è�@�aMF� �B���:����s��C�L7�"E�K�|w0~��~_+=OgQ��V�U����b�E1�m��s�&J�'�;$�W�������ƻC���v�}q+��.@#t�����T>�x/��S��ڗh�c^M����8I��Uuo- PP5���)��\�w��6�R��]ʳ�k����x���r�="�,��I1�@گtո9�����"&M[s�_�/�@�kT�'/�[�<1��އZ�/��Y:t��>�&F��tL ����E��W��{�j�<X�)C��wyH��l�2<�u��s�;;<���e1ga��O�%��n�c�=��i��:d�z�K:��!�u�����&u�j��4F/$���c����Kϓ�O��!y�mPڧ�$���6�Z3���:V�a��nʲq��-�BBΝk��bAt�C,�
Ν��i�{��,���1q�f�4,D�P�*�f��R�+���M�G�u�V\
�I:�5�qa{���3q�e8*��or��.A�F�4�4Ԝ�7��8 �����7Ҝer)��)�� MI�E���~)�;P9��p?��td�|��6�����D��G�n`�>O�]��Z����i����)cyB�d��{�ն� �}���v���Z�Й�R��Ohԡ�o̮y0v��1k���z	QqFA�d=�����wn��Xl���1��zїiP5�k��A)x���dOf��3�)i�p�09<���&��N���J����E�hdײ�t۞���E��q����`Rt]�W=�3���^i���i��Z<&*$�U��аA��}u�'�X|��W�Ԫ{�g��k5�8�]w���v���F�=�*����
*�կzqeit�"߽� t]����͖���ȳ�(��Zz�Zgڕ��(�B�����yS�ɲ��*O$P~��l�-����$�nھ^�0�љ�;gR���C`�(�d�C-6���&�j-�˧�t8�i�� �iv�픋`.K<b�y���|ξ�H��8-�.jIe���0ϐx��r�ox?�ꈛ�'gNaL�+�;�����.��r��~9����E�oۡ^��3hea�ߵ���mel��s�P4[��̂�5�����*��e�~"�֖-�Wﺺ|��<q/��3�,,/��S��[�t�lz����Z�ʾd�7 �y�B"=���L��H�'���	��_�����o%3��P�ďms.+�;�}Sv{^��R)f��Á�M����{������b{��ۅ���7���\��:ɝɑj�ց��<�;+&�ĳ^�̬y9,���t���E�F��A^	i���*K��u��F��'��L��++�z	�A�?��p~��M$�p,X&�r�ٟ��IL/-|Y�c���ZG����1L�P��ӼM۪�$�A*a���@t>� ��nd�� �cv 9~Z��G�^�����m�e�e$� �eZ���O)܋����H�����OW��u�sO���̸G�ێ@W|q1��՝�|(�2�i�C�=P��:�Їq�:8j���G�[���+�	7ı$���FM�P��Ҳ��"�	���,�:��]��N��2��h�)�O���=�L����x��M�up��i���2=��O�:�Ѵ���H��n�=�_̏6ĀT�.��������"�MIf�q�4����j�Tnp��>�T��Rsh��q�
p0%�D��	�Y,0D��\'������:D��B�7@3	����)՞�����=v�:���i܃�T�z�T��r1b�g*5��ŗ��رz�X�\��Z�<"�r����K��x�W�,$5�I����	8ǐYQ)����88�(�-ġ���w4�A�ͳg7���eiN��gN����:(r\#�B�g!L�k_=���`��W]/��^B�z���j=�JU� "@7��r���7c�*TR�l)�[
�|��.�t'����bd�d����I!�Rc{�L�Q���j��X���?&��,�ǋrT	� ,�
(��H��Z�n���2�"��]
򻟮u+�њl��(C<�����U+���X1�X}�~�� �����f������xO��C�rQ(H�{�4�ǎ�D�]��{��]���o��@���Y��z�e-�Q����F�3 �=��b%�O�$�e��ǵ�C~�a��h�tT�CO��ڷ�@�-(�jf5���R��q;�c�PM�ԅ���e���`�ï:�:�������ƌ'AΫֱ���귱��S\oW�l�`��֐d�h!��m�*��4i�ض�3W|�Q��Gf�s2|�>�)n0�T��c�k��M��6�@^V����a�2��4��M|Z
��E"x]�j�$�o�|M�Լ��2�KQ��"N�)��^u*�)��Ÿ�?m1�[K߆��1�&�	����Q������'XV��t���L���w+e��$g6���g�s��+�D��2�bV�;[֡��pq�4O�����0L���-3���U��1v�{��H��we�n��XԔFP([Mf%D���b�,��D���jz����XiuR��	X��Vi{�v����9M�(.��Ge����ٝ��lM��"�x�o��TW[A��zCT�g����B{�p����X��0��L���TH�n�Ņ�.�k����-+k#H�^B&V��h>�����Bu�/-lbF�}nS����rq���S�\6?I�!&Kk��Lzد�JQ����|oɗO�]SM���8�L�Н�Xˇ�\#�O�И���<@2�~S�㕀��Z�L��UQ@8�p��9�"����
HD�G�C�2GU�]͠�� 5�J}�{�Q1�^2k���ԈP�� �a6�#���|�΁����Vc(
,ŐD���P�ǜ=�,�L�&�u�	�Y'���|�-F��ɕ�QnEt05�z'�ed�޽���qq~�D�o����+("٠�p�`��|\<G�������g���yq� �p"h%�� ����G�ѸLH	[����z^ƀ���~I/��יP�8�H{v�Ι�^$���r'�U���\�� Ex��5)� /7�nj����l��:���׹�B5�#�qA���У��}簌#��X[R�����w���e8ͤ��Ҵ5��R{DB�A.�i�35Q������R�eߠBs�p�x�2!��3o�i@+�&�7���s9�Ҩ��P��ۏX1��V�Eg���lqR�M��
ȁ�`�72���C�{�\j�+���vf���m�r.�T��������Ĳ��}�<.���
L_{�-���|	�W�6�z1����w.���Dw�Ys^��+:޿ҹ}�؇�����ǣp������L �)c�e������ް��s���r�C�d��)���.I���3�GrBKJ|��"ԾYx��V~�P	f��N߇�1po%Ne�����H^"u����H� 2������U�ei~�7�x�ڍ�Sz,*u�5��.S7�G^������#P�Mw��0wwr�LЎ�RPf��LZ�����j�ۛ*�1�Nk8�fP�� 
$����~̤?�`t���"-Ϯ�4N����J�=�݀  �"Z�a���Y�T�mؙ/k+ �U~�������t�i�g���zz3�5���r�A�*�6��Oo�K��e�q��sQU��K���[\	.rT��x���=dփr�*o�s
��%*X�$&�m���!��h��2��+�3���!���:7����:�Tb���!4�͢CƠ��\q`�P��:fF����+_g��� i��a.�<�O� g@���!�60Kz ��px}D��@w����\�J�T����Z�t%C$��7�wߡ`��0��~�"e1憗��,@�M����cm;�[��f򿉧b=co�}�mDJ��(���I���>�$W�-MΒ��*潼?�#Գ2ה���I�D�T���9� h�u��`\tt�e�H���0�}	Y/��?�l�ƹI5�������,n=v�3Zw@�o�4�aLVڲ��'oNߠb��Z���Z[ffұ�X^=xi�cd� 3���	 �����Z��zr
�oh�.�H��!s15�5�Z��'(�V��A���H��ۏ���_`�?���iZ=|ïi.�� #3G(	/��!���ň�-�ڹW�'� ��J�*�0�>��G����F>�t܁�,)���tWn�X��ԃ��~��5���n�5�g2 堨J�ᇳ!;\�DF�Z�H�ܐ�ޅ�ԆL�9ӫ�5ɬ�n�������(F�P�*g��gƱ�b2y��3X91b����zz|7�S'��
ݜ��Cb�Fq�W��2�0��u�猨�{�T�x4�b�r��ey�d֩t晝����Ӻ�_��F7LMi�H����TK
dk:�E����/��$]O�h��!��*�:��sG1պ��+T�~3o`~�3���Mi�Y��/��fzxl	�u)mcL���#��5���o5�5��,�CW=c*:0���x��WDL&/:-�����^VC�����t}nOt��B.�Y̎#-������<���$X��,"G�n ��RSc�y�V{�7^���\.�{�.��IOn���t�Ei������Wڻ�H��:N�+�P֕V�啣�UFu�O+q�H���A�w�����"���l�Q#�xD��f�R�k�%& bΤ�Ig�30J��RDD�4�Tx�bi�
�ըy�XTO�ph5������ȕ��S��\�r����l�zG���,�UP���/���d]{�R�#��n���Ep�~�c�P�{��G�j]1��FfԪ+t�I�=P`���}4�&�NI�����0.�Ƹy�~�8ٌ����âȤ�����׆�@��x֑�+\[k��F��<nձWrx�p��m��Kc��wt�@��_τ�����P�bO^����XI#g??O)����T5Q����
aS�kp�2y���7x�� |�u�T��j�Оl' �n9o�1�KR�+�v��]���?�i@�(��X�o�q8Bz#�k`Ls��Y4�Y�.���Җ��<��q��uگa��8�PKNu!{���' *[���B��#`��ұ�,n.�F�N%_�R�'o��JO�O]>SQS��q�˾��'p2�����j��8{s�vB}��V+i�X�����ڊ?��ɰJB�:<c����GI��	�%��:����e���dV��c.j�w˚�se�4d��9��mX��Քz��>Qy�x��x��S|qd��)�u�/�^�~�bA0�������I�վh/��U`[�@005��`p��*�q(a?���P���v�$Dj�ښ����JTV0��]d�R��4���f^���%�f(ǐ��*�����h�� �뢝�hllŒp��`ȞG<���;+�/)>�_ur����_Q~0��}��'4��4|���
�d:!&M(E��҈%�����1OY���-�wh�*aK(1RV�z�Z�4�qP]|���R�F���<����4��#o�v�E���Ch+0.��@�X���(@�L-Y����YWPU�Lz�j�b9��K��� '�qix^�Wi�c��S�1J鳢N,�CO�����d |
hԏF�l"T��oH�Yfh�Fk�\@� 3���g.�sؚ�,�WZ�0g��
�}���d�ӟ �iצ�)_e2�}7���s��׎7��
��&n�1����=Qc�x���HB���Y��4����#׺ۏ�⬸r�F��=��{�[I�|@rbg��������/�X��@HH"۸���_I鱚��^�ޗkY��e�����[k{тi�s+
�;��2��G��$R�T����	m���<�S�ZSן��h�}m\]���q���[p�u�\��)!)ZF�H�逆x��T��r���������_��|�Zŕw%����k����Áã"�2tB���8(��������j	�:h���b�t\�vi�����e�����i��4�����b�l�d�	�*��d	 2q���~���fv���E�^A�;����j�X�K�K�{�	?�]�%1��_Ʃ��`�c�d�c��$���ʲ
ˮ����J�޲����N`Iʨ��-��o����2�s��DO�SX	��Px*�����Q����-;�ŮH� A.�f5>�����EZ3�F��������$wd�t���Xti!��R�����	V��I����6�L��?��G+z���DBEޒ��[:]�ɡn�P9�)�̮|��^��ukّ���o�/v�LQC��ud���[� �P��oE�1�z�Y�py݂wx����3�%U�n��2}�߂+�Z���H��������Я�w��������}�������ƭ-�M���S�'�̰?,�B��p�5�6,g
�wT4,�R?��9�-8���3<�Cy����Y�jA�ä+��d�/�`��� x��7iֶpZ͔gBd2���B��L1�;��v�W4m���-pv\[(�û-�M~t��d�m�[�-b�YY�.����׳!�To�d�4�%�]�q��2�ڼ�U�����~��V;�lW���'�K������a�^9�t��.ö����ͽ�#�����n�֝������C_T�J ^�6Z!v�,�X���߻���6ˆ4��䲅.����ɷBו;�&���ɱ��
�jS+���B�)��sa��1OBD�	��G�Ԇ�,�N�!�y��|�u2S����;�@x����o[�T�x�l�p������{���xz��wC����ߗMD�[�:8�+�_,��Ō�ѿ=+�A�y��MZ`�W�Q�+/{―�Mʆh�������C�v44-�*�=��GQ).��df��B�D�r�)�DE��_*C��d�{�=qD�p��ϖc�r9��L� U�kuQ�T�im��R
\!C�EF�I��c�S�~�c;d�L	� jP9���������U�t�� �j���ϴ*/��������q��;ɴ��n�'$�c^���	�G+˭�إ������WI�v˕�QXS�B>���K�?�CiQ�-�QOZ��q�y٠i��J&�����WAmK�5h@�j�W�0w,W�r����m���s�;?��$4�!����I�Pt�;��o��b�L�<��FqM�O�>��\c�Vg��kp�����f��Q3=��0�3�}�u��tm�II��9��(���mN��"��]ڰ�#�����l\���t����}x�MP�b�̈́dV��1��-����7~�X3��~)q�*�����{�m{}����$�u䈵�z���D��Z�'j�GzԡN>-��O��|��I���c|����B�f4�H&S�}z�m�D��qg�=:N�ޑ�,P��Fu`W<��sƮt�H�_��b��\�f�8�	�@�B!�&�r�w���PR���w�>.���k+í����+�$:ad9ᎅNO�ۭ��u�k4����Z������֍Ȉ��s@i�������Z��f�B��������^�<s��T�E�iDj�==�]p�O��k��~� �>Y�0��v]sE�Y���q�Uk��9�o���A��Q�]6�!t�%�jO���8}�ɢ?�$�[N����:ܽɾ�[�|\��>l�F�Ý�F�r��丣�	��itcN�J"r!�~��t�=]/#����Vxl�@ 1JG�
�)w���<8߲#�HcQ@'<5ǚ���� p|���>g�,�Z��Kd�D�Sr��~���`V��J�u\HQ�`�P�������Q������2��5�	����II�q}���v����1��S�	5�2J[������:ɺ�u��fJpYb�%����&�O=������������q{��L���7����\��(��z��}1N����P<�L��C�
\���S��(&�������kܰ� 

�����i(�g�ox�8|x->��_ ���,	�eׂ����'���GrBd��+��T/�.kt�>����M_DU'���KH���moj��R����Va�N�]�l[/p%K�Nqj^�JP~s˘�!���Ct,p�1�¶^R,��)o�H9y9�d,ѱ���@��/u͕BB~�tp���[�o�!�h/���A��$�7��:�Xg���=��x6[���� �2� 72�{.��6��w%�۟X�W�����:��$71mk:���lU�/�q����nD�}�"��2��%�yfQ)�65��Wl�
�y�j��<�:PWx��֟�l=�R��c[��|mc�- �B�^�/�U� h�ɵ����d�cu+���6%	�J���ԙ�����=��%�UhT[s6z9���H�N�oʪ��N'@E�g5�tB��bHj��o�'"�Ώ�����\�~�"��9V�-�s6�G�iFo��[����"#
#Y�@.Q@R��Z�\ m�("]�c�MS0�/�%���{n�>���z� ��9�(��؀N�M�	[�;��;4�v�uI�6��[�V����"�'���χ'fd?@� �YGH- >g?|k ^�w���U.�Y�yM@7l���,kL�d�I�����_t&�E��s6�Wa�b^�V^����S����-%v@q������J������g����1~���u��	�s^.��0������M���DNWZg���^k�t��"�5�g3�vH�>\�@d��y �΃��x#{額��)�/Q\^��	u4ū�����7�f�ރ66�$H��TDĦ�pJ���PC�}Z>H�￴fYc��$�U���G]�r0�I�P/���b��o�?h�k��)qU�rY���" ��3���j�iD�T�H/j�N$��oK�Ȗ��I8p��|���K�D��n�}5��P
R��Yv%�q�//9�y��{��&G�Z;��X�� �oz�[Sn��Z	1�l��K)�%Ϊ�����P9��I�}�	T[B��9�������TH<S��%����@�>�ݓ��$��yيÂF��㴽s*��NK�ˑ!��a���Q�A������Ƈ�<�U�{�ˋk�xu�p�7��=����gw�g����J�72# a?�-���s����#� ��b�5�bU\!j���ů�{�ŷ�_�@gA>��x�F>��W;�\��= �uY?��>@	b��V+G����M4�P$d�5P3�����$H���!�{.BM5��?��?��J�M��g�������ۢ�PQt�G�qi&�w��<�V��ZT��Y�e���PtJ��*?�o*��8�Qf#m��k"���R%���`�(�]-l�Ԝ�HL���������riM�[i('�޲�>���l�H�6�W]��j���`y��� k�VS_u��ZY�TZ�.(��Y��J=���n�)Q�\"8m��u��p)��?�aS�Ƙ;����-;�V'�1&��6�.�'K#���OfY�:�0'ťW�X�iE���.+��~]��FI�n\���I�J�|V5n����Ddb��?�n��0"��8fnd�>^���d�I[8��zL(zv������C9�����.(�0_�������."Z�50a�BV.h���t>(���3�X��Ƹ������<���[X{=,ɵ���M��{�� Q�(��<�2м"�_ǳ)o�o?c��|����E^�
��5��������r���y�P"�	�Y
Y��5�I���W�� np�]��L���K�v���	��vI7ۮV\�+�g���N;��c�$F�/Dހ�Տ��(�[$���i�!ll�5��$"8JJm|1iY�M�6�M��GD���˕.r�Fv�;����nݲ��Zd��$X�7���g>4e���8�>�ʫ����\h����J0��=�T��҉q2Tc�� ;loԃwd�9�	Lڜb�ւr��o�Â�T��=~�l�h�P���N�
�.
G3�ŮF�J�o]1���	�ǂd��P����"����*?�$� ���bXg�W<�MI�\�ԭp�5�[Lͫg�MV֪D$a9AcbGZQL�}�Av��c�j��X� ��M0�y6�(�z ��G�a�aigD������g� t��N�5�씻:��>�Jl�т���NP�K1.<ʘw�{��x�e?���ưy�T�������_W����c0N�q~�g�r,��Q�ǵ��;�h�#-{�K˺]�v��r���x�ޅPkg-'���V��uc��V����Z�?�x���e�(���ww���	\�������H���3�/1B'�*{�QyP���;�i͜�����ȁ��x�4�L$O=9��f�R�t�����4��9�yE2�"nr�i���F��C�i���a�[z��ʺ�V@�q���n����o$I��{��T�f�'a��}�kt�Cv@��9J�D���N�����+o�IS8�;F�E6��K�(Lg�i�!� D���d�mS�ӆ����֦�L7zg@�l�O�m�5���u��;�����*����.,CyJ%=iE�#�qߎ�4��Z��Y��>����پwL�m�S\Kc�Q����rSY'�
ն7mc�B�k�lwu���$��\�#-�WJ`��^������*��8�?km�ь[������%-������ˉү�2Lp(2T��ݙ���)&��j1�p�����ZbeH��| �����NO鬔�J 9��b�%�Z�ț��Ph{-�V�m8S��"�R�d%5/"��SJV�W�d��������
[�	��X�Ɗ�4�.���yl_24X�C�1��qR��S&2��������>��A:h��L٦���1�I��W�7n�E0��5n@mCB�2NM������)�g����Ґ�I�f=�?��G��P"�	������&�Z"�cNi��.3��oo���<���*���}����_�'Z�3o��'�*T�k�^���>L�<e̔q.�N=�<cॳ0U�ФS���i:�?��]9��M&�nߑ@���j!O(G��������x[m�^
45�$��n*�~HL_h�x��p7�5VG!����0�-��
ՙ�f^��iyJ�I����2�3Ej���Jyĝ&J�;C�-�EI�#�$z׎��L�����T$0���c�c⚵EК��	/��7�����23���?���$V�C�u��$�8s�;@��E�4�񩇺t]s)�ͻ �QgZr��G(��Py�!���1v�x�gGG>�=FbSG�������B[z'�NXP��7��Y�9�$�É�'l�_���l��-wippH�|WR훻LW��?Å�Z�_%�C��c��;c����r.�Z��}�P_�7||!������Et����[�×�m���s��$@ea���'�d�W =��\f4l�_�l��"s�;���)x�� ������<1�{S��5�]v#eU �yB��V%���%�-X:"� ����$�a11i��9�E�Q���g�O����$2nf��1����9(���f��>��d���vӋ�䈀�l�Xэ��rn�	y�����^��� �����j�&��n5�)�]X�X�FgD�C�nK?U�^���A3jS�ύ�)��,\���%lwk��N6���a��مq�M�{��ۓ�ɼ���T�v@��~j�Y�Vޖ�$�2DU*ɮ�<J��倾���(�F^��3/����-��:o��V4�s�/���d��%Z��G=|��n��V�Dbr�/��i�,��X�HuQ�Bo�b��-��,�>U�����b��[���hs�^�M��:w`��]1�BT��ȁc�x�`�����lW��iRAd�='�/�?!Pڵ7_l�M�B��
�8�ٛ��<~��g����=ǯ�Qlΐ ��4��WP�%k��:l��ZV@'���H�������L�Y*��"iEXٜx�~�����fr�k�P�a�-�*̝��vTOy��pO(al4�G��b�� �Q��(Qi(�����C���*�*���:*���9�
���D�u�g;��_���6�]~�z$oXw�;5ez�M>�&%1Lx�Pؤ<��5 �JNeoPP���٬����[��&���Q/=�]�J�%Ŭ��|�����7����	�D�WC17�S%����+�o@�y�[{#{V��G}���>W�LiXY;���gW2ޛ"��a����/�.z6>�LS�m�s<]H,�T�
���>T���Oa�a\&��F=8�<���;I��2��T�Gk{�
�z�;@�.Cm���ˀ7�sW���:S|�X�kz��p1V��&�����o�"/��t���xzIs�6��P����	D7���Z�v�6��ű�EG��d��k&#jk!G��Y�@���*���C���~N�"�t�CmuxhdG�ɡ)(k��(6��8�_� �ςغPil������k�;��	Ɗ��l�V3(��	��Iռ~gde�Ђa$NF.Z����Z�v�
�!�a�e{����+��Ζ�݅�~�5�7��C2i��+��`�^���2G�ڢ鸊�ҳ!9�	��M�7��]�~��6@�(5�u�c&�D(go��H��δ��[{6�j��`'}�v���ƪO�z���7�Hh��+Ф�cv���U��.?�;w�e�d���/t�8o\g=�(��Q�w�i�To�i�a�$�z��3������gŵN�����Z��h~N-"�h �C�� wh� ` ��E�O�~�RS�u��վ�`�fD�(pW�bZuf"rބ�A�Y<1#��/|�t�}W������x���"���jl�j3������!+���T�v��f��G�p���_
����p/�z�I�� ;SJv[o^1%YP;����̒H���S!\u�x�I��qK�a��RX����.d8���,�6���hEM �'|�����)�'QIa�4�	7�0�2
�~���J�7���Ԡ��	�~'��L�\D�y
{����d3�Z�M��T��M����v n\e�Qk�����VWW>{i����g�d�.�2
�� bPʄ$��JBGX߭�c�Q6�s@��cj��E�Q/���X���V�M�y$U=C�V!��i�DE��u�E���7"jtc�����j�还f/
>z�9��~�����97���Jq��Rb
'Yz�(�������[��{=t����X�.v$#_�U�8zI�1�ES%��|�/���B��6�Y�ću��@|�*--�z>�������D��ŋ?��Ϗ�&-�mF��%F����dC����z��nA�Qt(��_#h(<�}�Kœ~���(��qѪ�k�i�a��ʅ��K�Wu�{������U��`gsr=5'��_�4��zY�`�urcF;�kO����E^��¿T���pN寈��i���=~��M��
k�W�:�s!��~�����PX�DNr�osau��~�Ҿ��U�]���\�O����J�橛Lc/7���޽�Qt���,/]��E�WA�vH�R��Nέ}�NPǥ���z�e��xX'$�Sk�1N�avI8��L�DI�"�ȑ�_!LC���IyhYJ���+�ٚ$ܚ���p����]3�y�@@�gJ��h4d��;_v�2�}�wq��d1��| ��bB� >^��f���-����/����x�"މee�D��K������0I�^�f��RQi��X	��ɢ~��d��f��-�����2��5��\?-�[o;���B��K��M����ҫ��e��x��nC�12� ���������W���$�GC���քX��O�ΒA�Mހ~iӰY�S���Y*���s�F���:3�w:�� �c�_c���%���MG�ܯ�7�`!ˌ�a��� �|����F�٫��ZŔQ��hNZ���E\�δ_Em+p6P�MKV�A��/o�CR$�c�;�2�t�L�ɂ_Je;_�@16���N�J�[|���Ĉ{�mee��T��'�7�E�����98�NU�J�r�ҀsOl`!�]U� T��:�-�W;�Me��� �9�O���=�]N�B����E�uY��y<�Mo�������k=�Cv��ދ �[eE cM����+�I���+�=���f\H"Q��_�o�l0�jk�zvq}�51B��X��6�4׳����\n��
2v����$�旿8Ux�R�a6X����ݲ�������܊�^γ��IT�Q��M/hJk�^��oS$��]{O3�|A��޴o��=��K�'�!A5��G3�����MP��S/����q㮐�g��Q]�ȣ%�!@��-��[��G�:���$B'R��t�4dzcacpB��,:�A��[a�n�?��(�=U{W��6�J�l�f�"S!J�h!�RX?pP&�ۏ�"*��<��`�|�I��Ò!T!}gjj�Dx?b���\&*���iLG�c6a��nd�؇>a�����p����'����uJ�L��9�x����8V��ZX#}�+U2]cr��ߔ� 3Q�eE���NMuR�g�-�j����.e��j��n��!�6�˫ir����:�i��k�:AW�V"�;K#nH(dqNc�r*Mb���|v8��:Z�x��l
��m٤'T���KF�dkV&��V��~��~p��:��3��}{
!��{����<Y��ex�ǟ�\��)5�w\lC
~l��������PF�>vR/q�= Ӝ��tW��7��!�'�(9i�����4����Q+�qǖ͠:��ry��"ٌj|�9"4�)�(ݪ�9��n�w�8�,�U?}7,Nh�4��,��рz�6y����A�х��h���o͏�L�{�<1�wL�)}[�p0�׊�E0n�x%�]4���=��k���r��&���W��d��=B���x��B���C�,	��
v�|	��/7#l��b&��d��|�5	@��'E����.�W��<��d��>M �FԼbzUr��=`�K"E��/PYm�������3����i��C�ƥk�?���`T�!b81�Uˁ+�=�F²�m0WC�u��)Y9-ǝ�y%cj?��n�[X(	��}���:>��F��\�~G���H��/����Xg��Y��Q~���s��?��m�^���>�Gk�T=�������� ɟ�� @���3+΄T� �2�kj֪��/!K�<*C�|�>q�gg������N���XkwDҰ�j�z�����\8��l���j�1kw���u�jp�j�F;��wKJc<	;���:�>��Y��ljh�(�� TW���X�<��U�"?V����8)l0}*�9����Ցo}��c�9L�SR�¯���č���V�,��o�\VBBiz9�f�J��/غŃTtJ4��aַ�GQ`�d׉;}�����o��Z$O��~Yl�Y;�(��ԧs�zv�%�y�F@�~�Y�{ۃ e]��r���b��x3������0v�o�v���>U��$��CQ�Q�4���:��G#r��SP}�r�T ����O�g��y�r%	@�}�79T�@��ޅ��w�5{�'�x��Ot��l�τ��n0j�ҔӨ�g`�/�u͜a{Zz
)�ǜ�¥�ٺ�
��b�O���vk���g��MV��w��;��Cx���x-�;�wܧ�+>`�R�qL>7>�"��唘�S-6r5s�� �d �xm�t�y�rTy���"�g]�3�U�������c�*Qo�S8�w}�:e$� ��U
�R��Q�E�>+w���^`A5DnQ��B+��C0t4ͳ��@I�V
�G�V�x��J97��4ױSA�<)�i2d�a�'�������P-P)����^tP�����B�7��nC��(����`������P�UCg�K^����fqQ���j>-�����'1x��m�TN���.�\@gY�0ĩd����?����6�R"���ѝ��?G�T���:3$�'�!�S0PW}��!s�{��BR������lN
2R����WX��l��l��CO���!sBp"�-$s��!��*
�q���xc����4��C8����I�R��0f�虅����wg����.�h�͹CG�0kG������P�,i�V�{¾n�E���=���j��gHM[ >"H����Q��$���pǪHK�����ƫ�{*_�P��TΈߘ%�w������Q}����V-�A	;?b��>�����L��������^[b�s��C�LR	C����5�j�i�Ff>��_�@�1��#N��p�Y��D������dQ�Q��XWuMH�y�T@��~_7I�9�1��O�$��!�"dF���Hn!����}�;k���r=K_d:�\�/۞;˂��?d�U��8C�'7�~���_K�&lm~]����tUv�8\TNX]���&q{��;�J�*B H�)K�]�c&a��R�#]��ٺ�uD�{?Y]���Ly�6��f�=��I��K��׉{To�,j.״+���"vZ/jJs���h�AE��V$��v�V������u��v̄���Q�B����H���i(�#Y8*���0�-�p4�S$��&M�]���ף�,<h�K^�����E�`Lj�E���,��G�mH\����tf]�ݰh$�ZT!�S�q�&A�]��a$wtn����xB?9Cd��������D�M� �T<��(���E ��`i��n$x���[��$,r��޿�-c�C���X�'ܿ��)��Yˑ̱Ѝ���%�����S.M�b$�X�R=!����a�E�����i%;�h����(�j#��$� Z�V�<؁r�/B�vQ �c���p�	:��~�T�q��L�Lq���^4�4c��/O؜ېH,����W�D-.�����-+�P7'g�,^�:�������pb��JS�zD�iz���S�L�b`s��v�n�#
�c!2֢��P��(��%�9��k?@�3Is�p�ΫMظ׿a~}���_`5�_D����g؈<$�ЗI�M��e��c��P�O�l�5�X^qv,SʸY�m;�c�C���c��ہ�!a�R��{1���Ŧ�e���q�T]�����K�X������K�_�x�g�c�fS�`9(j���8��!2���6��+�]w��; ���'t,�d���(t���`\����A����^S(roÜ�Uևۄ�$����Vk�fQB��>
�^�9�1���}0]ᜮ	��S&��O�&�Uۦ��eh�g�qDrg�s�W=�A�͛�ް�t�|{z�/-c��u=�H�+e@s�)nC)M��0����U*����X��\)�j��gL�{[��h�͆@j�Lz#q듸	�g��<��фv�t��UrD/ӷLyr���G�vEʣ��?Sg����������;�2�W�2��~�v�������{�����w��W6	��I��~L�8�aQ<��	P��E[�+�sY�T�@:����?�6��#��?�"�.����-��.n��3H�,��4k�������o������ո�FdY?V'��T�,�b��S��� h��-}u-���}�񑷢 i��ō��V��'[|c����Wt1�W��-�$ (p^�~�o�=���ݬ��
J�����tEg�M&L�K{��$39�ױT�0k! �|V��Z�U��#�|��kz�'��5/�2No	�y,��N]�Q>O�hd��WC�=%91�#���uЋw��"�xx���0y�\6��լ�_�JZғ�j%�*�zI�� \\��w����NN6�y"�	?=|zb����9���7z�\�?t(`6�T�%��?�L��RPvk���(��*��PT|��>�k��D��HFV��S��18�RbmH�nd����O��M㞀|�rX^��:�@ٹ��!.I�B�5�8��t*"K�lO#�s�Bm�~4k$F�Rڨ�૰k������,�>�m= �s8 ��q��_�Kp��Uk�d�^l��\�c�쿉�Y&xSN��d��g&���#a s����d�(r�Eg�P��g8��n�o���FݔcƉ�{��l9ܗ��rjw4��?� �ݣ
\�'a-�_/v+�lv����L/}8��Vn���o�4��`8#��*�η��W7� 	�v�-�L:�f#��B�5�VO��oO-wH��tE��)�B�aλ�+k7���+T�Z��f|��� �����GG�^X(�/~��mf��#���e�����	���mVR4c��|��R>Yk*�%�F-�����(V[l�T�ҕ�ʐ�K�+gl	u��[��E�13II�J��hVXT��޶����}]w�4�4��R-�y	��+�/�|�Qa�}��6c\vh��gdD1��-����@�^7݈�`@��a恙ȹ_ڌ;�+G�;�`��NP������C���1���L.T���W`�y���j!�I��_ia~��6S��_��&ԣ�\`��z�Ro(Qx�ɐ4������O���d�g�)�MT�>@n��bXb]�!���T��eh}zGR�!{O�k�Y���:g�*%�(J���o~�'ȓ��r.��	��a �����$�� ��=$B�jy�`��<�a�T?��	Z�T�d��N#nsl	�ԧ=X'A�~�G��q��<PKIY^8a0ifM/w	<^�����j%O�л�ď�<n��{E���hl�� x���^	�X}Y�����Z8�X����m�CC����j:�G�����&�6�a���e�{������D�h�����JnY��r��%����H��IF@�=Ƥ=Yw�Y��=������eY��CJ6\��&078[�V�Te��w�|^�&�c��Z{�eJQ��-_�4u�e��&`�~?D�h�Jzk����E��t�ё���m�r��e���F�1qD���P��\�׍���}&�Ϲx�7h��ݕr�Ϫ.�آ!6�͆�����Y����n�ģ=�ND��LZu���8�	I�M\q�E�/��dͦ7W^P]/������ ܘD�uM�o�r�r�8|����\7�ͨ�����7��v>f��lR�>�B54zܜ�i� 
�j5�Y�T����~�Y���wݶ�f;.��E�L:��6�� ;����y�.R��h1��Ϛ�(wY����^��u9�� �^�����&���r�|� 	޾�A��{�`3+0-�L�����KC�c����E����T�V�,	��b��Z�l�ʧ��zT��I�ٽ�3 ��7���7M��{]�/�S�ڂc�.(�$�1kc�����l�W4��G�WefJ� �/�h�.Y��ZI��t��I����K�j~�{�5|l���UT-�D̴r�]&zԎ.iw	�C�fD����1�|7d��٦]��5�^������gr
������_�ӣ��3�XN��!8�G�� R���iPBt��0!�5��8���G� �lEܝ#c�&�u��6��D�t�˖���'VAd�Ӂ��kʧ{�Ju��n{L#�s�osr��@p�L�&]�.M,wr��\Z=2�X�t#�g�I��a+Oo��;敭*+f��}��a��Rذ�s4&}�f PƢ2Fk�DX/�#$�+�ş�^o�z����cp��~�4(vf���z1��*�+�2 ��h=�r����'I�nJ"��m�4t�HϤ<�12h6�ɹY�Ml��ߩm0�g-�۔�����C�;��!�$�	,�m��Q�̴��6kM�ᦦ `fሸ*r�*��I����xB����,է�X=���N�!����X^l��3t�� �i�x�t@3�3DRV89$���dM��ދ�ךZkU�Q��SmS��j�3�W��U��1b ���aXTQɆ\��\��Ѿ,7�R�.��/���"*�"ִ�����9�_8D���pvOWk���4OEb,�l�wR����&'�uC�c�|�sg�>^�dF\�mݡ��<� �|ONp��h�t�����E�� ���'Q���kB�yu�-���U }ٰ�Tj���
��>�^3j���\j��^�d7/�&ܘA��Ȗn��;�h��V�[�\�Rj��VI���l��E���#���ra��$�D;7��iĦC��w���N£-o���r'�G�<��' ;ï[���WVĖS2��
��uTƷ	Y'���y�����5�|�n��%��g4��Y�TU{���W�,e_���n�"B>�nf��*Z@R� Ya<��6��8���k#��2(�g�&���b��xb�!�0��8�̦ 8[&dVQ�Z�!���N|Q��}��K� �C�K
R���m�&^ap�"	$Z����E�=a�F�Px��&@��jn)�;g����$A&�K*������#��ؐY��3�"��O����=�z�1���A�e9Y�AoF"e.9��`P���?3^g;�3#Aì[C� gc��G�n7$�=�?M\�_�f��:�P\�B��60���B���8m�G�Q��ZrO���:�}�ډ}�>N��c��@ �]&��eۨQWY��T�2 ���`���&��1����g6ڻ2�v-7_��^t���X�+I4)b�p9�V3��R�{n[�T
��*7�Q!Av^J����~�hFǤ�z�@� H�wx�/S�G���d�_h�����%-|�ʉG-��q����2�m�*#
��-d(]  �
[�jH���W�B/P�L�mpY���K�A����V�����⃀�w^�.������MZ��o��m*g��������+=�]8�����+���P)(��=@�����aE}:ԏꝖ�r��<�i�t(��z���e�<�"@��W`��)
����{��<������XB�;%��tla�o�n��*�ׇ�C�O�,+A�+Y�*(�tE&𮕰����L/�~��~]��}�H\���dη4���@�!�`*�ڭ���L˫j�2���PR$d������jt3>���./;)�.u�ARk{ҼbD)K�V����)>��t�Z9Ǘ|��xڐsׁ>����0r))�xQ�<��H�12��!��4�N"�i�	��>�<�J ��Lq�üXT�H�$.)vz�;�Iw�6��5�tى$���U�Ӭ�P��̓%&z��g.刅ܠ��C?�u��M��(��wt�eZ����\d�y��.T[zF�l�V�"���!m���-E�Ϛ�F����M"�(��	�z��o�K�z�e�k/�V�����7�$�(l~A��zM�=� T�x+O��� ne����e�\��K�
Y��P�:G�Z�L�$q`�	R�X0W�)�i�"��V<w�{��0��À[CIy��
t���.7�C�HS���0�����ha�/�ǽ�eO.a���[~�J96���ް�2�g�8���1S�?1�7��'$���) ��P\�ʬ�Ԕ����\ݺ��p���8Q]�b�z֮�3#�@�i2U�EU(hA�V��3�I�Xt!��S\}p�(����V&�����?�n]�@�yc�SIS����s����i��K��Q����/��.��Se�{ȑ���>�0��Ef��g����,�)NX��͑W��r���Y�`E���#Ooh�U������/�,n�Ľ+"ي3��*m"+�b��k�m�ECeD@Kh�8��=�[�q)@�<�]�2���+�|��˪	��%���l�,4M
^��W�z"�NM�|8gN!�tR0}�S�ԁ��s�:�kY_���6�Hu�br�z�[�Ζ���q3�Aab����͞��DUD��ײf��,)}����nA"���
Ҡ�Z��M��Y;Y>3����H>� 0D����nLv�j[�,)Ky��0��zV�H�JT��2�/�N�&�n��w��3�U%�z~��k�d���ﺅ��9���mvh�z% fr0�y�m��
 ��s��z8����f����g��xE�v�tp��f��l��ݕ���0 )m�?S�6z��e��A��NӶR�hԪ�Q�{Ĵ&l�<�<��p.�W�K�oF���Y:��|z�����b PEA�p^u��D�QľZV��k�
��
����"�`#��:�[�c�*�����,	~�:&��$-� ��g�8u�֐znu�\��K����#6�o��P�ȝQ|��(��6Է�Uc�^	
vve"H�UX�%�_�B�1�./�t.�]���{�e��9~3{��a�Y�ʇm�/0�X�'�Cm;���@���a��>H��U\��j>~�]���=Å8���[Zm�6�O�<���ٶŎ֣ꓻ+`&��qEG33b���������M+.$d�<o磹�
be�8�
�"qβE�b��h僸�v).}�f���BmC!Z`�ث�*�;q��,���P�>�gL����}g��{��C,���wI׺c���!���A�YZ��e��~ICRb>��j�~�a�ᄹ�3]�����նѸ�~�"�q�G�@�Ἳ9bk�#��E��� ܌��� ��;��8 �tz\*;f��v)7�4��n�
�C]��Y�'��љESw	�p�H6Q�b���=J���Q�ut���XJא��{m�h��m�Ŗ�D�UE�o}r�s��g��(Gu�OI�#�{l���S�O�8��)F8 �΋������E%r��f��I��Ѱ��n<�~k,嶧�L*!�w('~A[[O�fw�Dٖ����|�,�w�CI�lh� F_;�`j[��V�=:�,�o�y�g���;�J�߂d |׾�A�I���\de��yC.HAK.�\s���ϕ'����#B�ʒK��l�3�:�Xa�;[f^�)���gQϳ�W!<��/�����FqWX0����M��^�k׀���-�Ʊ������J��.kY�<�����a4��ކLr��g��]!�4	����`=��������d�9gz���G�{�>ӓ;T<�ӈ3�9(�~�@�:�1���@j����9tt���e�� �v���T2��
GH���X��
o�P%�g�|R-:P*��gwm^w�[Fa�/!M\%�]�����	�A�V�ш�F�p
�^|D�mK�&g�ޕ�������׿��H߻�$�9��� 0zʠ�KX�#u�,Uo���["^��a	zR*M�zc�1�9��L{}�t�ːa�V��q��qT+���J���ީ� �g�[��g��!R� ^��,�ɸ�QA.�yMz��X��ϣ�3��È��ox�A�\������T�!�3��uU"������&|�����_������>+�X��-�yZ͂k�_��o<�R�V+�W쩹X*��J����RrgL�>��ݭ�RG���Q�G�s�2y�,�P���ʻ���lt��������ۮ���(�VT�ĊL�}�*HC;W�ʧ~N¡Z���F`h(x�
+e�t������XT�v&��&a��S�<���L0��g����A$_,t��2m�w�k���uCF����%��Fᵠ1����f�I(��ץ݆w^�u�bfd/\���-ߙǝ����K��0!R�����o�yrA��y���Y�����T�����HLۉ�s������E�oI�wvj{Hj�Gť!�<�G�G�=TTy&We�ܦa�a��d}[��t(	����:?��A�� �?x�ym[��.3�Ei�51��	w�J�J�
H�LPm�|�	����v�'��"&��n��X����9���ǰ�V0b��QO���2�X�А,�fp��j���V�ߦ�uU���ݞ-f��(<l�x.�%h�>���b ��ߙP��|]����VA��0 ���\X,e�e��}n�΍�/h��\�Q�Oa�����Fc}ݟ-��p���0!8�y4M�����Mm�^ૉ�>���oED]X,`�]9A>`7�#:z�+��&D8�{W����a��ǈ#٢��n�4�pL��ֈkn@�6g�m���=�˩_����8���c9�>��l�z�=�M=O�|EU�*�u�YAx瞣�V��� ��8�E����m_1Ϯze�U|3q!��j�>ڈ����O�Vu,Qވ
C��Z���+�$�������,��d�$�' -vo�i��H��*���u�j�̜-�������H���Ή閕sn��{'{�B�z9���V�.�[�v�SE$��V�s��A�r����¯J��Y�w�e5��	��rߨ�����̲�k��~�� ߲D���ҽ09�KS�y,��g��IxŽߙ��兼3h�4��w�]7�aMc�����}a�l@)Y�ږ3g��17��nt��<���V�]�n�E|�V4C>Cf=s�U�>��a��iS ։°�JU����c�{�nBisѸ��H��q�XJ�UF��sO��e��̱�M���ދ��*���rZK��~��i=��
�ŵA�X(]r�ͼe��C�[\��֒W���B|����봶j��Hhvz���c6��z]S�2�T�zZt��X`�Z�D<��]|a�MȺ�Z�e�܅Ja�B�G K�l��mn�Y�W�]/ݩ�t��Ԋ[�x6�hj�J�5
����Zf��撒�^I	�,���6��B�ijq	�NУ�]�kx*
���ŧ��)ug��T@|�u- ���OWov���*en����X�;��U��X���lK����Ҟ���ڬ3c�3�a���I��r�QuX�z�H���o��)��ٲ�c�Оb��	l�/��'w+��Ǧ�*�����,�g޽Fn�1k�:KB's�d�>c�n��z@?����0�a2+]K�Y��x7vH*U��P]	�]q'<)��*L-TP@������J2�~�-��)'v���A���1z�Og5>� �=��G� �< ����yw��Z�/���V4����=��?��t�o���!�!Oi����n��hG ��|�ܯVe3�PG�o��D���1Cl���2k� �ZY[�;l�3���q�n�w�y�I6S|,�8�)��c}��?Qn����u�1���� 5gh�B���DMY���Z�D�u�g7�J��P"�k;�p���~�w�$����B���}1�\�f�
ȊS�Ot�Bռ,�<��V�P�G�!��3#'6	�]B��5h/QS�]ai~�9��
��w���0�^�D/�o��R+}T�������|����5�FX"�"�5�6���լ�SGOXN��+'�(Kc��!~�	�@q��zR��Z�;LQAq!_��[���;�=�^���Х�^-x��Na�����8�	�-��{:�;�3�>@"��mϼݢy�Lc�����n;�5&��l���J�6�1��u�L�#gg�B�0�ٲ���o���Gd[a�g
����v�3${��6ëo?�d����P6	G�>�k+�O��l�9������_��,"�X�=��xm���Ats.!T�b���vQnl)_���y*��0�s#���5���������߶:�	���^u�2G ��� �y��i;�뵵��<'Dj���xtq���2��%���@�I�8ל� /��@mY�P/m��lZo^�~2F��i%������|�������H� cO�ǞV`l`��=࠹�X��7��ܲ�@����
"~6���ouՈ�Oc�D�u����Gw+J�$�p��	�t�v	1#*bZ��py$��J�FuI�̒U���~�҅CͶ^u(�Q_S��*��z�T��8�����~?��v�|��w�2����{��5�"L¡C�.�=�3�|� (rE�k[�2�2E�Y��ΫdZR���YqZ� ;�~�oШv�c����"�����r	"P�}�
��y����/^"A�Ynr{*��+��k+I��8��(/ ��X}�Ⱥ��mvK#E �UI�]�Yj��5���#�� ���p&89�ǨS`�� ?q��Z�H�9+}C��L�)��3�G=��X#o����9�	��S���{�D!h��4�K��g��a6���^I�[|��������V�.�!����L}?}�65
#6�(R�@����p}ߙ$�p�ˍ�
N�^zg��K��4zɾ�wk�Oe˼� �ju��9VX1���p�H����v�����E������'&�o�߄�k�T�M�$@l��SN����r���̆����&��yXo����TK��6&�2F�F��YR���#�f�B�J��������'�=��9c��G��3�\S�ARq�1?�!>�tg��}�
үδ�2e՟EF�	x�h�l���(�Ŭ�x��l*�ߤ.W#<�F�<0�:���ݪ�����������⁂`�[�Y����-!�L%В �_d����׆�!vc5��M���n���Z,n@����v����H�n�ϑ�L��˰.�اfV��39>������FUPk�Xz�}�ϡHA-��wH�Zf��,A����H�E����%F��ĥI쁒�JG�]@P�BD���\���Y�߾w�� n]��3���^D_��ȖO��F�+�B�vIw��5��/s,�p��X�:��{`����E� �mc��5�s�P"V�>�f|�U(���OE�3Fq։^F��Ǖ�m[����XO�!*�d��D��T��m���Ч<|�F�o`�C�>A'C�*�1�Õ��>A�zT�T�f7�{��%�D���c�Fd\�O$��ّ4F۳��ۄ����i��eN�H1cp9�v��(����5F�1~��<���o=��������8������G;��=6Y��q@�6ZJ��ہ�{T��X�#Sv"�X�&u:I�ѿ���Y	�S6;|PT0�ٯR�t�~]��5�IzX<!�'�AL�K1��n�w���bG9��i��(A��E@D�=��`Τ�2��u�Sv��峝��x��*���Gf�Ҩ�.ӉsI�"�[)}L��`d��m��'��m���&�������<�����Q�^O�Y >�������������%�M��v��rɉ��u��������S,�\U�D�K�C.�#�f��f�V�2���g���w�/�#�ՄF�YbL�N�Ꮴy�"d�Z��V;�\ՙ̼�R(6�2�xq���z8�4 j`9ce_T�Rԍ���ֽ���d�q���w�_~���vWA�Oµn�O9<pl��B|��6�0�iJ�(�i˽����sk�A�էO~̓o`�J�N��H�es���ULr��mY�\�Ԅ1šQ� ��W�qrK�,��0���W%���*�ג�ټ���>,��ݚ���OȦ/
��*�XN�P9�M^K�t��i�������Pܗ'����:���V���q����tN���!��c[V� |�/iѿ�1�<h�� ����-B��Z�rC���|k����g����hu-�n_u/��RQ�����RV�iF��QB`g��EN�P�:�9�%0�Z��)N�.��񆢭j�����g�����sg�wp�e����a*�ޓ&M��?�[�{��̤�ZϹ�������sHg�$�P����2�c��"�e�o�?!��`A%/�\q�^M�w�����K���Cj[c�:�ֹ7�.���ו�-Јɜ\�*�����˗���c��U���r�P���C9Q�ȑ퓦[r#��U*�#��Tիz��|y:׎�0TcÔ�v�<�`<B��IF�Ů?}�V����6W�6h~���-�����ߧ� W��tЯZ-,�;!���$�h�!����8̦�9�N��~�N�fA�쥜�*�+�M��tɏ ���A[�&U��.�+fg�d��X��$m�(���F ����%����"�E���&���j(�����1�;S�������g�,�V2	i��5؁�{{�ף�}P̓�G����Ø(ളc6�����	��X+�X��T��2AZa��H+�,��S#��K"��=��B׊��"�$�x�Ia�/9
V�$ȑ����9�Z*@ [��g�p��ֲV�U�V��J�Zu'���j$��U*���W�.&�ߜw2��V��c47��E��.W�睮t� � nN!R;$Ү `C�.��Y8�me���`P!	�Pmwl	D�"j�(<{��I	�� ͺv�=���Y�hOn�t�辸���y!�i[®��Ho����{�~Ͳ��f=hAbBtIi��X�ݒfaٍ#,��F-wnF�,��m ��H�:�=nt����6�V��G��h�p\
3��JiZS}����B����A\ :�pq��; e��Y��v�FTtnVL1k����=���2>O����f�E5F���ȃ�F��&wN �v���2T�]�s���[<�����D�A�V��m��F�@�>Ӊ�^;Jb������%�@��Gc�B����u�^x�7���[���ȶL�8������\���M�U�lb)����¬��H(�V`Oz4�8壷]���;z�����z�gXrQ\��T��W	WLu�R�vP]�̚_�
h�ml��Ֆ׌�D2/�1'����~y���U�j�;�������w�z��"6�Q��ַ�t͈��M§�h�&�n�C
b��	��y&c@����vX�7���"Ǹ�>�c[<| M�kN�YH�A����=����񚉮Ó�h���k�D�l��т �$N�5b���kI,>Rhҩ�!��ːHw�r]��gT�b >ſ�M���)[{��v��Ymκ%ʩ_��L��qi�{�ÞRc��ٹvl��T������R+�Cz]����L�N��UL�h�]H!��$#��p��8�����P>P}i@�]���a�7����)x[��O4>�}�~�N��8Snzc��9�-?���i��S�����;4�R�Z F����!e��kv�t��oČw��@"�2!,"�k�byZ@�j[�2��T��L�x8owrQ��M���<���1qP�=���
��j�C5Y3��wǣ��~������f\&9�b��}UC�Ѷ>`�;O��ţ�=�E�ħ�9�����!�*���`㯐�_ʏ���C�6��P������������)z8�Z�z�o�X�@Hi��i��₎2\)?���(7��b�oP��SZ!�24��
�����[��NQ__�.���F������x�I��y�n7h�S�IӠ�D�;���|D�O��O;��o-$����a�5'�T��Ĩ���+&S��TS�eK������ħ�I�4^:���Kw�]\������=���C�Qۅ�@T����X�Մg�xl��֛ e��zl���F��a���E��#&A#u?X�5�u�2�ў���������!�����[3|v�희�A�3$E��~U����P!����IL�z�����Fs�)����;OɊ����f,��f0���馴���?MSL*�8J�&7���ۋ&<Gխ�r,jt��k����~ZF�x���b�rP�m�/|�6jU{���r�u�4F�'p�{� Ee�&$�z3�[&pD1iLڍd�լ�d$���R`4h�x�
�{��XS�-�1�:��eS��W�a�]�ڭ��ޤo3:���auo��j\������?�D��3'�p|ף��*�W����x#B<0ԟ�v��QD��_$�f� O�c��W��o�\���7�i�(z��N��ʛ�p!�g^TTW�-�k���@WP�0�{�؝)��I�eK-	py���b7�q��$5Pk����O�Np�س�ZL���hػ�v@�͍��os���X�+Z�Ņ�G���,�w��b��z-0:�6���Hd��m��#.0CF
˖���TM�$��An\�H e�3����c,/t%Aձ����z�ah���f{���#�CAJT�n�w�Bh-�b.�Y8�JFy�7Q+_J]�LZ�a_\��tF�H~z,��?0@a�l��1��N8�2Q_f^qh�{��S-Xҏy���P�sC�K�C�lo����U)��-r�9L=M�\�:�m	��>.�o��Ϳq>��@�q�e���w.Lr@)'[Xh����/�X�5ݸ!1��Q�4�pֻ̨��wGk��V��!F_���jӡg�VH��f����_5�W��F�2�!b�c�}���_,��<��U7����Ɠ��������Pu�N�����H�aKtkC,��8no��vn�E���q7�;�[J�}|����ip�X�`���� �;�^���I>�����/X�t d�x����Y��$�ä�N�q A��W���8��U��_�3M��������7�o�F��ϻ�f�b@K�$�Ts:Ϋ�TK~��ו��0���x6����u}޲��D8����� ���������1XN!�@R,�9�m�	�z@]:�Y��M�`�lg��z��n+=�JE�~�^�ʘ�MEi����5����/��D���K�?Ln���w��p jW#��'(X��wrͲ����a r!q�;�j&T������ᐧ|S�b�E��U�ǽ60�tғp��t6�Z��H1b��!�Q-EVO��RuG��#�<"�������W@wu?,�Г~WY���z2��U�yUH�ohX�Coҭ%��i�b�)��1{շ���j+�������d�9�8�a-o&��������c��԰�J�(]�r�=��W�"���\��,c�?H���S���H2�1.��1�lK�e�3�)��B�������k�f�#�ħ�W�ݨ��,A�C}�w�_�t{�+�����x$��q8������K�؂m��؜�O��ҟ�b���y�+��u!���H�jS�� d���Ê΀c ���k�n�
�x�60�^%0~m\-����$XmT��=$DLap�l�]D�(��*>����Z�0˴!��e���Km?o���(�En�5Ēv"��F�g��&�p7o�/`] B�ص��kqw�,�Z5�!|�z{%�gx.�u[)B��Y	5�2C80gǀ&	�����C��Eزq�a�LQ����p%��h�谚K���9B����x"qՉ�a4TWĬ\2/
�]��%���Kq��r�S�j��@�#_�ú0����].e�G�r���{<��HUU��+���A���I���>K�� f�#9+��u�vy�ړ���&y�d��s��b!S�N��:	l�Z3��D�Nj�^�nڶ�f�8QF,10�l�o��0�i�d��Jl���s����)~'��bI�0;��|��~ɎUTV�JIl�h3�$�q�)�VL.��Hqwv��tO�3J�,h���ʬ�f���F9�- ��흂��y�K1���G�KӒ���u���"':�o�F��Hȫ��ҟ$�9�4�ʓX�N�x?��]��/Z>�,�t�f�O���:IK����3`W���9G�bݑ����>�u�l^~��УB
��?�e�*�#'[�����Jf<}'���h��B�:}|�SPț�U/���Լi\Ӂ�{/İ疐���� ����M��#	4J��n@%�TPػ���W�w��$I�����ho��B�J��Q9]�*��	�<M|
��*���S�8%8��0$ Ui"�Xm+3�J�D����������
E��(��w��Ǯk�j���ZQ�<�>ί]F���H��VN�"rKNq��0XpscZ��5�|Rԃ�5��ġ�㐥�,����#�.��t�oeO���@�;�
D����� �>9�O�wUћ�^U���F�������3"|�=�;�q�R9FYM�� 1��O�'��|����Z�P��L	��"����r�A�|�!���j�Ԣ@"`KPL�ϧMr�`�1d����zi6����|�/&���jm�	�#&����f��NF49 aH�����h)�v{�R�+��H{ˮVk��7xvR���a^k�G��m�b\�%%��1��Q�$�n�16_�U�d�P�����߰��њ�9���g�S�i�)R	�����Ps<�d�$���	oN��}Z��M����6>�s�#�e�I&M��z7�.+� Ɋ�FxJ� �kҙ�tvut����mF���ՅmL�;}	pvޫ��;3/9r$��$\���2���t�"m�e�8�Ī��V���7�9�!����tXo����s�AY��҄G��Gv����*d�~w��+c�����a����s��A��Vd|A�IP�P~p����Q �#���-�����.��q�O��(��G�f�h�#E]Ty�0gގ4��<r�2��m���9d�A"[�	�/�Fռ���1Z���%͉C�o����#(|=��z��3���^¨�{�g�_8�pI�N����ؔR��eS�9~��X�%�%i��fp뒪�di�|�k[�j]�%��G�����O2jm.��>|d�Ƅ�Ȧ�k�T�&uЭ����\�2���H{�%:l;$���ޢ���jA���/Z��W�l�}5#{9�^�&�l�J�(:H���߅#& N���
a�[�`/��;�b�j�������.P���)H��B6�����Ҡ��iw �A��RI\H疅(�]�!�I�?�ľ�� ��H�
{Q�q������A!#=&Y����~���U��uu�X�Z�ӏ�~��c9�f�U��1��\�.}�<�l�LOצ���u�֏Ȗ^i/H h�=�6J�_�hː)m~9U&q,kWl6T] �8�׸.��2��7s\�d���l����S�<@�qߙ����B����߼�S��$X��!h�ڒ�m$�������)��`댬k�Sv�;���'ů�w$�~(���T����# !Yƀ�����D] �]�z��t��Mv��_��4�~��M�I�6	<�^�r|��ZxJ�*�q�����S�+����";#��o>쓨��A�Mk8L�5B���!,<^)���t:�~�)I��3$�l�	Z���GJ�[����#G9��i8�2>�����ySDzQ������~˯�7���0m��d��~�G�^�ѳ|����,�������i�DjQ+�ܥ�Yn�];�U�����s,l2����;�jc��J�h�}nF<i�Q�D
�$q߻�d���R��C���;�}Z��jn`��<�R�H���8bd�t�!Fz��L�y�o�&W��Ϗ��r�}���қݒ�t�~���+`�����Uj5�|�	�VdPN#��ώ�e�ĝ/�:B�1�)�xb6<��ԪK�v��F�I	����ѡ��ئi��RQ���F�`A������<K�7L2���]hnk��nLi0;u�ք�H�����B�2���K���+W)f���?^�U�������0���s�䁠)�#��)V|#��f�5���n����o:��}� ��m{l��@� �ї�7�1P`��f������S-E�T2\�׉��]?� ���,�2��Zf�<��Q��S[��>M���p� R�����(�1(�	��&Y�9��9����QC���VjQ0B+"_��#�Q����|��~R�P�xj�
{�$k^��.��8�.�ܲ��zF|�0��hȤ5]���5�3�0H���z�P��
i;�Ц��6.�^���5wOHQ��[,|ms������qI`B4��"[	!�#o�o$c���l������
1}P�lc���%����u�wg3�o���9��ɺ��H,NޑPj�Cm��zXyb;��E������\Xv�����Pu�N��2	oV�C��w�3S����D�2��h3��|�(#�\K�J�O�t�c�`J�e̩+fR�a�a*!hۄ-*M�2�����i[�u��C��=���_�k�_tqx�W��ǐ�w�m��%^"���f ��i�@r��Ze�+��%w�P֨�Ȍ�>`K��R_�p}!���ۤ���'���@�w���ᆙz��#YL�al}�K�%V�X��K�N����r��0��V��g�O�٠
x��9��d��r�CFL�~P���!�k�� x� 	��j�5��8���Mש�cm\�|C9B����|ᥚ'Y��k_����9�3�Ts�4?O�ܣ�I�������ʑl)s���g�k �h�f���"F6���)'0�A*ZHh�}^�,�u£.14�pj.���#g,W�rka��Pq��(��F.�昑w���(錀jBChSYk:�Oy�'/�g�w@'�7E�+����kM�����ޙ)��z%(T�`0����r26�Fx޲U�^�k�C'����ԵQ���8�{17N[���5au�>�z�Y��Z|ꌢ��0��?�x|G�	�{��
Z�"ie������zy|����G5ǞjI\�enq�}��f�T�(�y��ɹ�/�H��_��NNk����V�h��5�kS�Fg,#E7��O9��"�}]��{I/��x��jP�T��� �bT�L��	�Ԇ���'�F`�y�D,g��e8��hk+8��/�i}C�!⾙'0@l�s'�T��"��_�~z��U��V�H�:�C������$js�h�f᝚�`Z| @k������R�f@�-\S��f�sK��H���i��  ����B���U��3l���i`"Y+;@u��L��֬�$�)���]x���W�y��q|�WZ�M=PI���N�:����
�a�c��*�Y#!٘�p'`*���M��WdH�4�,�aEG�/X)�(��7��i��0F!e�$��'(�5�X��ml��3��A{r�N����� ��T�H:H�拵#���f{�V��z�2q2YD!J?�-bB̈?��u�۽��M6�KR�ɒ�$��I��H���!���pmFO���ts*g�1��M��Zxzy��S9��7A��.D��|�e̓vX65Y����<:{�ig���Ƀ ��0�Y(�>Y��@[�����\��0����4&�E��Lۏ��e'�������z��� l�*�ED��:�[�+���L�$Q�|��,���#iQZv���	Ag�{MR�Չ鶉FNkSe�/�����ͧ���*�₮�B2:�(@3G�'����m�%�5F�u�����������8��Z��F�� pZ"|� X��&�����_��ma�1zN��0�qGn��bHTp88�,��B��j���j��2}��x�Sh��L�)�����@v�e���; 6��t�AXP8S���$�vN�dR�����KGB8l�̊$��֫�������j(�.S#wT���g��OS�w��r)�c@�I�UX6-�	p���N@8�d&�V
T��#V�P�j���\hea��s@Y�c�&�=g6~4��"�],I��]��"G�wnq� �3k5������0�S ��FF1خ7�\����?rԳ�E��"o�=�Ɨ(���G�3�t+Ϡ}�U �{�#f���뼯�]����_f�W��z�-���D<��������
�$&7��θ�;���r�#�	���/	5+�<�u��4��_�Y���~O�_��oLq�1�Z��ɣA0)�<.�m|�@��� [3�3}���F�����`B7�P�?������ɬ���K��I߹Y��ʞ���ӝ��4XNg�����&CC}� G�;d0τy��,
��1�D{H��>Q}�ќ��+��bv��݄Np`�$�2�E��w��M�~�^����}�s�³6��xd}�T�]?��8�7�u:���w=�#�L�5
.΀@���[�x"��{r[-0���Ң=ÿG�B3/��O���_��<N��7k�"x�2s��Y�:q�b�d��)|Zez�b\����m\��qZ���8vg��~`�� |���OlA�^4X��1�����nȁv��3zo<:�,1���d�Wd��������f�#����t��xeuK��Ct�,9,�m.jA���~�� fd�������C����m�u�!f��-T�1�\������Z�{˨±6��D���.�]ش�*�tr
��_^����yp>V �q��Id� \��Ͳ�l��"�i	���ٱ^�'�ڙ�琭�J|Ӧ���똪�&^�^˘\�8��+i?��#N���b�Y�T�eK����	��7>b%���L�p삷�c�m������Կ�Xc��v���Jt6�e��`�`-��.�R�Ƭ�b#��;p�7��1��F���Pi�#i*�.MF#�If�Y��c�
p�wʔ�ˀ;����
�T���~�E���������Wh�BFw���_�q��,���O�H6"���`On<:����=��������iE�of�6�\.;9�a�,`'��=r����/�Kz��;W��%DOU��W�;O,���E���.��ÚNq~�dhoq7Q��l	mI:J@��#@-3�����?�5��^$�箸8M�0ej�)c��Pn��^81� �F�ILuo���(�+[J�?$8�!����
��7����a$��ԋm�Hf����)A��a�@eص�K�ir�����e������H�	ua8 ���XX�۶,�E������2����7�U��[�4��z�����
y��A���0=l���WJîl�ݣ�",2H��]~� �	���o*-H�*������z�(����k*e|�K��|�G�(+@�נ����8��Yh�5��ԛ���Lآ�Ҏ8=9�^��en�	�C�4��>����0/��Rp��ޑ�N�=4�O�݃ⷅ�`Wo��Doˮ�3�J����UT ~� zao˪���|�c��_�������d�I#�&.JUH�6�:/~#$I�<X�����%�Fē/��mK���bS<��@V�<���x����� ����|A$*w�>^6y�|e�SCV�&�f���L��0��$�>b�-H��?_�+�n�7�\/��y,�6m%�Qm�S8+�S���2��<~�u�������U؍Y���ާ��<"*�3�D��s�Ⱦ��yI��bƄ�,��_�r$��^2����6���1������z԰B�#R�^�Q���I�]�"��rٓ�]\H�<�hH�Nb��&�k��y�^t�T>����;�aJt�w���fK3&;�G���c�\"r+���d�x��GNLE�v�pV��W���Ł50�м��DJ̩��jU}�	N�K��W�͛]o��b����z�A��&�������4�@��Hx،���,��"�W�k�l�T{`���O�dz����O�����;<��c���	th��q�3��"8��i,����yf�� �ƈx2v����7�kl�P�3s���?����c81G�ܥ��Мj�Hy��G���Y����(���s ����