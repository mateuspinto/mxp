��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���mQ� ^$�k��Z�.d�/�1�<�3h)�W3
�v��O���q��ï��7�Z��N�bq
W�g4��n=�|��<�E���fw?���u"�X4^�?R8��(�$�Q�k3��@S#�^��%��E#��kw$O<��	C�gPH���)�r�OQS�M�a"��VPUG���b�>FМ��0�Z���ĺ9�����]l�<Z\�N���pv�|̳��kŉǂ����}W/E�(\GDR���~��gt,'�hV�������:�-]&���}���ߝ��
��ݔ|Ϥ��71���u}Y��������"~�+�g���T��f��¼X���U3U�U�w+�#t��<'��0�D+t���q�|@���a�<���Q�����I@r�;xM���v�j�>U�-�1���Y�O���h˞�m�5u���J��G|�X+����M�w]%�.�����+�Jz�Ͼ+�]-:��f6���͐���O� FyhM8���֜�e�¾_:TC�j��a0��ht�~5V�ԘR'[��7��+�tC�!�r �0�l��w�%.U*�u�G���3.a���@��2�V��"�)%I��~WP���hm�2���K��m�X]~�M���O���%��<G�&��p�;HQ�`�ɏ�V��Kc�D�|+�����/nxQ���p�+$O%o���)��5�]:��Ʃ��MB���2���3��Eܦ��A���ϲ�ߓ�XK$Ɵ�ʈ����p;��~z|}��
�v�֌պ�V�����<��s8�� �q�o�WQ��vV���]Dٯ���h���Rs��7�Quk>(C<�F�Uɐ=�θ����:�R�J�d��\w-��l������M��\�5)΋\T��7G{*@�TQ��\���Ւ���Y5☇A�q�]�˧�Ŗ?g��=鲎D���a9:���t��W`��bP��;D�j'����έ��<S�C�x�+$�I����ſI��`��X��I+��>YҠ&hU��ĹMl��6}�6鳈F3;��)H�gޝh�����^e�`C���끛���=���B��D&&Ü�d�G��US�c z �ABi#���a�J+Mz���YMi� Q�[A�7)8�L@�=
BPkA)}:�-b�@y�.��h���{�Ք�����<b���v;�혙����` KR5�����8�1�O�r��!�]�h"_N���-��^�IHJ��v1�k�	WWp�e��k6�a���a�XD�%`D���}�,����L���و+9�c�{P`n�<4������Ͷ�ꀥrN;��20e_a0�� D��h:g��WRΛ�(2Ea#�_�d�=R?z�|�"�c�}����-[ND�'��A�Ā���,�E������q�&�Ò�Ds$܌e�]nW3p���0屬vK�!RG��癖�5������D�/�`"=2�s�T{�#"cȆI��>v����z�zǵ��x��T�X�n]%Qg<&�C����d��&8���8ad�(y�h�vs��]	��^!������R�_��؆�¼d}6���ֺ�'!�\w8�w=8�����~�;��8�=��D�4k����p�l�h5��0B2�E���Ğz}�\�Z���'�O�?�����IA�=���`€���u�|ՠ1x�`r����Y��2�>r����WU8/%J���wfr?�X��[�>;�IM�v?MW�s�g�p5n���4<��S���c��ˊ!��B������{Ýh��;���Ҏ��댈F��s~.9�}��x�*>}'k4
��Y"��L��r6�a�2����+�do������9��q���~ݴv:+H	����Ŝ�;�uS?�c����ݤ���ѥ#���W��-����z�_]��ZWF��o
�[9��Pu-������|;� 8�>�5Ma�q3(;�I��x��h��wͽˀ�Ԑ�I��