��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���=�^���{3�%���\h�:�0x�஑�Z��:ԊZ[�J������a���!�v���0��Ȥ�O����h��B^�Zsχ�����֫d�odvw��%k��W{�{y���P�J�������ڋϼ7A��a#~*P�7���!�e��m�"�ɞ�4�d�U|�+\u�s]��},�F�M���i��P$�ˬ!�2Y��o;�\�������{%�_���u�j�~�sŰ�\�Tjl�[b�o���f D���G\5[������u�g�2u��.�h�G<�EÛ�����N3��>v�6�7�ޱ��g��f����­eb��؋�d�c���|SD����8@]�[�V�h�
����yL!5�NK"���|}v�߆/��i�br%u�1y�w����1��\@DY�X_J��-��S�?ݘ����-s���rZ�����U/j���4��W�_h�)k�,�9}��_���ؽx�n�G>����IG�q+��;7�̲�$�����bO<W�B��x7��� ��j��������3�]�flXW�VZ�w�Tn���I(�1�B�X�tb��-ri�l�نk¤�����������j W,E"�"��.e�o����3�ꈉ��`��~I�D�Ѥ���<R�K��F3Sj��<��ľ���ء[s��*�t��e&��N���i�^����e�4�j5��.B*t�Ku�c��"#'&�ӑ����W���2��d�띻B`��(�Ii�@��������w� �	��&��AR=�Bwq��/�Bgqf�6|ן�����װע؃D���碌
:��ghmײ+Ijr��U�5����&���P��T��,?���2�;2����Ŕѩ[e3]h��p��}�]��9͚*�?DiƲ����i�q4҉����W�d�K��}k��D����x�R�-�H�fh��5lH���w9Yj`Bj&S��1�ء:t-�ᖷ&�潗,��o���W���JR[�G�r��^�ӭZ)S��F����7�y���x�
�~59�Ԧ9�ɟ���]�L���M����S�{�e����7Tΐ�2����;7�C �n����Bb��vH<��V�(~�hU�F����7��ʊ��a`���b1%\��>V��p�vs��|�0��^	����pS��*�dP��t�����£W����9�PG�H�ג �$tc���=�kn	%u5 �3��Xs�a4���ߒ�1��G�!�p�w o?v�q���:��B�/I�vW�A��^j�qh��:��^x��Ҧ6<���`��J�!)$~�o���\F�C����0��7�#a�����_����3(�Z�f��^u4>!Y:e�O5�$К����HŔ�I�fbިE��#�V!�f��"�������f���&�}���ܱ#�?�z��T��,���C�!K��k���sy���"���_��|0��=0����+jj���q���X��Z�%|C��V���Sw���+�s	c�65�-�uu��t����K�C���I��jڎ�O������XM���t����>��Ok����\;ru�~&�4��|� ��Ǵ)�0ﺮ+���]v>[d�/^}���4���B��[�̟� �@F%Rd'i�[��6 H<Y���Gͣ��$%�X@I�3�g�A`7oA�e�5cY���nA��ѕ��%�Ot�'W[$��9����rWR�^�����Q�?�3�`��;�7~�R�a���MLS��Mc��6��%a��℆��4G�'rۦ�y�Ϟ��L��N����;O{�1z�ɍ"���˚�$��	`�L�HbL�ѺU�)��H������S-���Q����f&��:�m�-˰P��em �"G����4vt��!��x�BOY���v.M�y����ӗZg�ByT"IjU�1R�V
p�2!dK��c�����v�W�b�Ҕ=��%�}%_���?����gV�uWg�T���U���Hy��j�q��sn�v�'G�^0�Au�F@c���0i!�nK��q'<m��04z�
5�Ⱥ��[�E:Z;��5���Sa����``���C��#D�S���}� ���Rr���r��t�q�o�$�=f2I��� �ܜ��/_	6,���2|*���V���+��5>
߈�5�g[}0w�Pql$ml:O�rky���b2�7�t' �R�����o���31Kif�J-���]��[�V���,���������@��P��i"�7�I����hYv{���nk&�:<�#{}��C���բIFGu��C�ȃ�6�w&Sa��������+�DVuk�eXs�p����28����Ƒ�����Ɗ@_�=�������[�9�T��n,�D�fN���i� �nJ�3Ǝp������*~G�o��a���I���rf�i��JO�D	*!��#����2p�lD	ل�B[8�b�Љ\K������ZMp ��N�=SU`�*���V�����k9LM`���?�i��M?E�S ��٠�Ȭ���3���[<v2He"�7���4����x
��|�V���6���p��W�o� �
k��M(���d�+*�;w��DW}/]��'��'���c���#�?��f"jW��	������d|�-vǃw�]����I�M<��d�܂
����o��	�+f�J��e�>�"W��;&b�2-�n���C5�U���\��h��<��E�<	���`�Y*����[y��#�$_/e[7/x��e��C׏��<���@�^Mк�Cv��q�����Fe�MI&y���>6Ie�<�����<]����cD�#(0��yw�?��Z��҃�P�4����c�D���������)9GK*��z����������J*Q���&Y����o|���B����t��R|L�ф%=޾��l��b�_#����>B2*����G��?��i���<�����l���eԿ�=a�9���_Z�B˛��Q�G�E����d��[0�U��1�i~��D%5/RNo�؅��X5�M�����U�Z�/�vZ�����tʆ��b�\&/J��>��4�L���q�,�W��@t�gD	��c�� ��3OeA�I&�~������X�?@�1�4Pl;!2<i�ᦳB��ܒ
}��-A�2�HI�]@�ۏ�ܓ|Siɯ�i������/����n�)�E�ɹ�V �����a�|�Z�;��)�-C`o�O6�f��][�0@ab�����3j5QB�Tg�_��@f0�uU�h�=���1��8�s�!���Y.`�e@8����?+ғ-e����ݘ?��$�/�,��F�G�����y�ҟ��!�|��B�ޟ�Z�ӱc(	g�FZ�-]JYSgW �~+~"R
�-rmB�'2����Ri!��R�v0����i�ð���n��5�2MKĥ�p���30?w"��O��RDb�d�0���)O���X"�p^��9F�컫W�}v�����<t�-�Wh�2�Xj����]+I��C?��������O���������(�LJg���g/ IS}�^��Q>g`+A��/Pg�Fr���m���:�7a�oN��N��I�p����;��_�W��F���ȇ��L����|�k@��E�3�hܞG�|�2#Y 7�^+'���*k�aN�]m��s��)��g�<������?=���l@e�Iü%P
��p�]�Z���|�r�=�`*Oj��b�r8�Zw�`�	���{%�K�������b����1q�K�U!bR0	g���'%��ơ:�%��r��Gz	� ��C׶l��U�4�����Kt}�ŀǑ�/�MI/��
�]�u���y`�ᢉ�אƐС�b/��m��g�\��@�	���̂���t����|�U~�P���@�6���I�#��G�3��~��f�5L�LJb���%���Ө��ڸB��_Q��K#�Q)���b�x��l�:���U*��}�Vɤ�T-Oue�Ϊ�E�݃h���c�c�x+q�ѦI�~_��i*����(�a⌡�
TiDG���ڜJ2�v�/6z�����S�@�NԽoy���AE}��C�H ��>_7�)�/����$���l������ի�(Fy~����Y��'��S�B9�s�	u��m��D���I�'�w7}#�b���FcA��5E�A�]?Kܠ�l�Uڊƒ�Q��jnn�n }���w��=��ƫ�4�[��=l�I�.�$]Jx���$pIx�3u�$k����Qa�X��{L�q��l`W�/�7�|�e��ZG̰��fbѐnKOZ]P3�x� �	F�^�G��ѳ�F�3�[���ڿU��P����6��c!�JH{�H��6�<�Vd\���d��3����mo�&?QeGX����7S��B�s0����ߒ���bW����~�È���V�8$�;EiN_�80lө���iГ�Ț�g���#M>,w�y����{ ���L�dE�/*��'�2Gn�53���8&f+��xki�� ��w��%�H����Q ���V�YFuN�׳f!^�	�# �$�7���M��,&51"����dl�Kd?�z;n�ʉ�D���0/�{UZ/i��{yJ��W3;�q �@����،�p�8<I��d�O8(�Bl�o���H�|���7䔒�<���Q���C��|�y��ĝ�W����c�F�V[�� o��w��k~]��v;�PI�9�O*��Js���*"��:���_h��+�I{^0aQ$@��]�ޝt�����A��}y�mc�� ��O&5�{^��3���.�|CM��!�ae0z1�k5#��$io���:7nt_{���|���,2��ߵ�Ƈ � ���� Ε��&P��?�\�>�h�qّ��e��"1��jYG&�� �G߼���,�����$ʰ�z�:��J�v`� a��ԙ�R7��sү��u�P�P(l��)����=Y�A�qp�ޘ*]��K"��u��Qf�`=rJ(�sc+'��;�[�!�w�h�M
t�Rᦄ}���1<�?-�M�:��n�I0��6'��o�A|8f� )񟇱-���*�J;��R����*���:��=.� ĳ=��ō��}����(ó�]D���:ww��#��@T���ð����u���a%#�6J�l�&��B�,�ٿe���O�����AG֎Vc&���׶揪y7g�F���6�!Y�>0�"ڼ��d��؂~�4��X���#���M����,!e��֢>��k�Ԏ�-���ƬW����76C]���[�_�ն�+ �j�|u�"�\~���_��k{z�X?�2_R��_�-��1��ߌ(�L���4X������ճ��ѭ�1�龁�g����B��A8�p�6�y�f��\��:����S�Zg� �/�wC��a�%�Y|�ݕ�|�vV����½��G93j�\���w��rP��Y!��p���s��zY\�'g��ς߹ڬ޽����Wķ�`�V�t�s��{w�����,m�ݽ�
��D��;=�2�Ʀ��/4���Yq���s7bg
Ԉ�Z��)K�d��Uعej���N��L����iS�Hڲ�4��dI����x��l�٭$A؊j{�n��SKͯ4F)�~��I�[ҟ����/�������I�CB��l0���0y|����
/����n���3'Ɠ�����|��J��H�{~�OĄF�Ϳ�A��_��'�O���U#��.C�y�VL��KPt�T;B�9	����aTI���������Aw�e�����q6��7,G@\�W�&��e���5[H�C��\&���i2�/<oaE����j�m�VP�B�tJ���1u�C;ܲf�G 0�1�:������1RlEx)�� �<���*�@�Ϝ9C���r�{��*��+��f�"���\.�1����Q��-,� DI
�&�$�4��E�Y��y���pGy�@�O(�}(ॲ����Мb[M���u���=nY�����w굡�*)�>��C�M=`
��]��5-��)�j"��G+foO�A�Yy��>L��f .1��5�o�?rh��V�� :��W���p�l2;|���`�pJ���������J��M���U��',��q ir6GO9o��Ĥ*�kB�^ ��]���0]q����,j� �ҵ�!.�^c���MO�8S_NH�z5�p�Cvl#���>��9������D-:B�
;)õxs����O��S��CS�!	ܵb��S��՞�P��	��	����cOA@�βe������W��fFd�e�8�D�Y]��x�=#b��%���2���#��aM���a�X�(�o�����t�l���J�ڝ"�1?�V#ȕ7�����L��A!5��.ߍ̭sjlC�D�K�}�˂<%әj="hMy�p��Lβ!��CVG1�٪���FR#
�/k�>�n �gp�+;.�v?T̰�P\��dɒʳ���E�iy�m��J(b�eg�x�+1��:+ۧ<��6�1fU�=/I��Z��^�Y�`+-"	�,�7�����L'p�O�|M��l����0P��(3��dg�Ph!�}�D�n1}0�4ZV�+JRYP��4�Y��e��)�6f	��v�y3�dp�N���V)��q��j�ϭ1ﮮ ��b��ΎEc��,�s=ӛzE&:Al=Ky�$vUϡ�}Wڽ���`aO�{������H��E�C)�+�MM�{�/Y%��l������l�bE�vz���a� �P�k�.+>*�Vj�-�8�xx�K�m����]� 9�}�F���¦x���0��~հD:2� ��U�PJ��+	��rLr��J�4�u=8\�
�d�ƉOCFk��p��p2��������P�'���g�q�>]��l��#�{��@]�$fn���s<討8)qvuP��W��7A?�f���\�a�3�Z0��땙Cň�M��J����5v�a*��t�=�t�5��*��n���)��-"�ž2X��c��hK�"�+(:���g���b`���gk/.Sz��yZ���X��UT�߈�]�O��]D������żK2xYiF��Mxs[�=-k�n�25�*��A�����U>�@��h�iQ4Ue8� ���??yԤ��|�`]+�F�^Z4n4����c�҅�+}8�<�[�:��D����)!0TyJ�"*� Z���G^���I��"�Nn[~��O�~��=n��tj
�@�C���s����<��zN3)n�H�Xɐ��r�"}ZOd�Za��(�c�ǯe"����zu����!a)��e=�RFuS�O=�G#���ʕ`��P���ځ,1�E0���d#�',)l�2�=\�o��Kf~�h�&w�
%OX�]��xgb��>e��m��3HpJ�R	�Bn�$�*ۗ��%_�Cis�\�ubX��oT��ed�mZ$#�`��e1�I�$R�c�p�(�+����QYV@�GG���5^�n$)R-�vE��/���p/���]��{y�noN�g D�s/���Yk�͏��R�R	}'�;��+�pCQ�Ge��~$�7W����&���܏	�O��-%�`L��M8�i'�Vw�+�,R�M5	O��$HT��}���u�ne�L���N��G�n������q�=��XI�x��\�T���f�2D��?>�R���3R*T1��ϩ�s�H��ڊ�uo���%�" � ��d����^�U%sJ�@U˓��CY���T(�'$�0#S:0+�/}6�>���I{b>��Ԥ��>��)�$$�7hA'3�SgF% ��gG�j��w��w�3�
�8�8����AC	ݔ
�6�y�c�gC�h'2K��]�KP�a�1��o�0]�@�Lp�	��qC�����)��
pg׀u<[T�Z�����ش�r0���KSu��<A�i.z���-5d�@��x_~a׽�ڠz0};��PRF��k.Q���{�*~?LǴ�TWJx� r� C�S���*Dg��yi�,s�J���%��щw#�hN�_�N�K���)�}��{�چ������h��<N��x��Hud�,���;1E��s�����i�8�^�Wu\k��t�
\.�{_���O��I��U -/�Ó՗ej}:�`X�!�$�kK���e�A�s|�P�{�gH���Ge�q[��m�-t��7u��m�V��en�P�W[�������a#S�0��`� �-|v½��+��]���k~�-�����ۛ�w�rZ-B(9ɝx"߆�n���;��y�c7_�"/	}�q�Y��LۅNp���8ƤXT���VNȾ�?8��M�	_A�c�fi�-�?��4��ɂH)	,@�xIAԶZ�GdI �j1_�Q\��"4ъ�eFh��h�Q�_#�e�� � �Q΅.�U��d=����t����>�vG8�^qSr���<���B
���ɕ�)��W�F&AF�>u�V�z������D�Q�Dr��B�y����y$P����Al����-��xW~��ۧt �#�c.kJA�7deт�R,c�A,�)�Ɨ'�x�@��8�n駃r�#��z-�����A�N��R���q�]����W��N����
GF��Q+�O�v��Wd���R��Hף�e�1�#���b9�`�W�5ݡ�+[%V�[-+��èe��:���պb��>�&j�e6���_��m���ƻYDؒ��0�M�����T�|�O1c6[0X�����U��D{���X<	��6�X�bn(=��L1��I��i�n]�-��G5�FU�a�-(�]����k�T�z��ъDދ�*�r8W�	�ԣ9I�AdDM����xm�H$!0c3%)�7�s�6B�D����~E��y����yl���V{<�	�5i7���	���Aw]4No��4sv��|�V��9��?��'i�o�"�aC*0�c9Q�޶쥬0��1#�&��{M`[i�t���,*�������ԲVe�m��� �Ip`�t�#��H7g�M�ny��R�ٽ�[V���Z��%o�(q-|`�뙫daZ\��n��Ӭ3�9��9��B�kA]{Vl�5���HFd��YG��꫅/�wj��^����/��L+n�ӦmP^NT���l��y���nU6S��HąÈ�+_����$��hOs���5�In:m2���]۲2��z,�.�=��t=�9��a��1����g�Prĸ6+�.Ҽ�����R��{�&!޴2�`�XK��!��j����#W�ȕ�}�����f��+ibj"����;�(�E���!���,K��ѳd%@���N��aVη���b���!�c�ZTW냱���G[�Ďc�����������XS� �d��9�U#l��� ^�kXx$���	���c�R�Qg����A�Q�2D�Gb��ٰe�<��>s�x��S3�q>\d�Kà\3��6�eM����l�3��ڎ5`g�{zbP���Y�'��(����=r�|��Zg�/��kn�o�H�M5YH����x�e�T`�$н�Ru���m�BlR���ڴ s�tt��(��/q����I��1B�A��jv��k��3�_��C�}'~Er�l��-�Su�Huy]B͵�*�Yh8 ��f�~���R�n}�Y�������G$��]�XK餀��� �5�l��Pt8�o���2��t������<�7�%V��k�Q����1BW�b7Rt]~ە��_�7�`���f���́��%�>�/5��}"��G*�ؘ�0\���)��ؑ�31&�Z�_���}�$�݂�$/}� '��QiS�.˻��k��=����LGG�>ꭧOP�<Ruo�N�L2��N�<��i�uHNMҬ|~ZQ��`T՞ى�]��0������V��M���C�ET�V±���Y0.�_�@�3�R���-�ނ�w�m����^�ݻ<15=݅���e�A��)�d�n�ċRP��ͤV0���u�H�-�6��C^9�	�<$d��z��[�=��\��׻���]��rz�q]<�^��e��BAr��,O�9��$]�"O&�j>9h�;�@z��ү:� AϿ��op�a������?�
J^���T F��)cNx�
�vJv�N D�bn�Ԍ`w]��7��ǥg��O�ԝ����ۨ��˜J �%�)�ظ-�w�N�
�a*��'x^�.�D��K:}���]EC>U�#=}��u����&)��P��emx�$_��,�u��]������m�]�
P�����:��n��Ξ�Ż/��*��{n�sO܀<�fFK��Wh���Lm�nȶ��F,�\ee�K]�x��r��,�Ʌ�N����HH� ���rm���Ej܊W� �� �˞�\�tv�yl]��;~��c�r�P%Պ���}��~-�D�lb�o�2 M��v�@%=����d�Ow�i����(�b8$�*W�Q�+�!��(漚���Z/��!��J�[E����8����\,�g�������/]�(�����~�վ�4~�-f9��L
�{�L-�-��1�}*,��D���Ռ�H^��N���Z!|-"
�1��� �Y��>et.l����րh9�e���'�1Vy9$$���:�L������ �H�F�����4�1���m��eZWq������1e��Ll��h�I:���w������� ��5+�0��J ���u��d��f�Y��Jta7��ؒ?���`X
��=��^l��]�td�[W�],��<[V�P�?���iPi��71M�Mb!X/e@S�B�����nL�������2�����Yr�)v�꥗M��?�#h�O�u����!�*���o��������7���/n�O/=)�p{�?��;]��:}�F�Z�ٍ�"qQ�T@L�������E�4��s:?�k�+ހ&��t�io�'%�^��r�v�ܥ7�Ry|��X��˥��r�8qw�����+�Pvȝ�"���v��Y:�%�%S�c-�:�7��u�xl.�&3��;(�l�B�I�SHU����o�a�r:!d�w�޵��`� ���'��� -�͋����)���Z�6�v��ż��JZD�2��oU��ƵZ�w6ػ�
G�
�A/��6���<�m�4��q�DO�&��	y��k~!�b��`��l�[T����r�'��|��t��Z�|R�Ck�uX�U\##Ћ ��%�>���⭩r�ԅ?��>gd�ԍU��t_���Mѝ��Е(�|a��S�V��Lt\"��Z �"�>�N�t�8��ո������a��܈������~�#�a����`������Ӹd��}�)�iu�!���eYBx�E�y齫�e^}���w����i�+�V*����4�(QUq95�Mŉ�gj(�;h��n�"2 ��ZpRj�4"F.yt(q��o ;zӶ� Ü�\&H����l��ݢ�2���~�*Rft��
�U󦴠WDt�J�:�� }A՗�+n �O�-?��%4���J�q��b]h����m��g�Y�(֧��3�roK}�Uf���G�{0�2�I+E��(��Im�y_,�v��զ���%8
���5��?pL�V�n�r���x9\�����I�rPo��Y����������s2 0h��p)N=�n����8��L��;-b�m_�M�+cAǟMPD��Q���0n��W��Ou�_���;V��|����Xs�+3���lN��������0�bT�;�KRϱ���}����G`�lH��'���=�'F5� 0S���*{�����u�~���[���(�w��r��� ��f>Ff](�C��X?ڸc�]kQM�*$!C	��Y�p�bZ��d���Z_E:le���qv,��݇��X��GV9�h��{�/��D� \�Ġ�����i^�{�b�)�_H�����8�UNزX�
�a?
y+�=�`ǈ���4P$�����,4����W�ߍa](�	�wL�Vi2bʼ@Q~D/�:i�?�pb��	�%�7ܞ��b�?���#r��,$�	�K6W�*��%��)�	�	�"|PK:�z<�V�DP����X���M9���K���2��)�S^b�U}H� ��5Ў�]����1Ḽ�t4�M����t\�W{��O�����fw"� 0��5��UZ>��h�����G��!q���#��C��v����tt��&ej0��k�`6>�~9-4T����1($�"|�S
��go�j�D��ht	�nY�~�JJ���M�zi~���?B�ѭ����k�#*�͋ɥ��/C[�7�_Kr���!%dz��v�dur��܊=@���n�ӂ�;(<ٙ���+z�P��Lqu�וh�%芣w��Ç0;�y�0+�1֯��_&�nJ<�e?3���8�F�lne�i�m����5�t$�Zd�9%�\�iO�\���Ԓ���=��NxN&y�.�.�
ZM'BՒ�B�Y�B{RW��k0yp#�w_Ė�Y{m���m�Ԍ��(�Ll@t���D���jłL1`�|�<j'��-w�yg|5���絭L/ ]����o�����,�̛��լtP?;��Ԗ���H�_�<|TlӸ~���š�滇W�m�v��E����NU�s)��c�Js�3s��"��ƨ|bp��dmo�{����x��@F�M�&��?�Q{ө�B0�9k(���:يs/tee�@|�y����;ִ9� �0���1}�y�Z�ȦEE��;bU'�X�\���sU<N����=g�z���Z���g��=���Y��j��w��_.�����e�ҽ�3<��5ͼ?��Q�9�(�RG{��Fw����݌>:��K%��/:Kq۟tO&Ϝ�w�l,��/^�ɋ�æV	��M=��7�!�WݯȼL����>�e��~2%J��˟����V��o��m%��Yۨ���$ܪ�J��^,��
�x�Ks�[���K�C��p�Q�ڕ��׻�9祿�gT}f��oL�7��"�ͧn�7���v�-e����=靷"�1���]�LW����se�9Փ�R����	s��[UV!�f� ���{�.��S��z��`D+���5}���+���JBqY�
��&��h$ÊA^��G=�'��(�4zY��v�F����Q@�?x��/H@S3��QF��:�p�� n�%ǻ�����rj�o�Êڃ�AIy��A��I[��A���'���Ft�s�H ����tr$b�4F9̏�+���-�{�M~8�a��똷5��Q���gb�L���N���n�;�b+��>Do#���+���r����Z���=���b��qPy�[�Z1�������։x��������^��!0�o���B����>MF�����?e�Q�%�Rm�I�i�ͺ:��4�^�uL[7԰��1�v�� � ��U�z����k�5	�G�E�u�3�ܕ�6�p<�
�tLs/0lN}�W��	��׈���*�����ߜ	C��)��M_����@���Q��Lr܇�m�7}�X�~^S�g X���m�w����C��ݨn�z��=��&2�K���n��y�܌)@�������2OL�F���	�_�D(?�ߥ;�-�G�A?��g�$4]�?��Byy��"n����D��KϞ4^z/Eo���T�+�8�U,�y�Ŋ�j
�%�b%㈛A���s%���|��䗠k�?�9*y����ǉb��0��9B�I��h����r�"�v-<�����(�`��w,�������"����1Ę��;��52]��y�{}��R_�s�	O�Q��
}���h�����5\3e����_J�.}ܼ��'\��gG�$��r��Br��b����nY��B�����o14�A�cK���r���]Z����I�c�6�Y���L�.}��0���4�-���A����.��9�u�ش�H�-D���� ���D�1�`vȋ,0�s��r�S�W�c!�C�1�������0,�*�Ǟ ��d*\o?�?qxu��DD���� �i�O|�a�5�&���Z�_ ��قNs��~,����Y�IL5{F��{��G� ���Mk��3�3D���S@��.�U
��ⓑ����.f|��ў�p͑iӖ��b۷��"
P��5�]j�+
qi�.�$�����/3���K�q���E����k���W�'��$�oT�Ny۠���ts4|կ�H���k5Wɪ1T40Oj�(-|�@s�T�CDV����UF���b��ED��61��C(���Dx�E�.�z�ۿLb~�uۨJ���^�"���uo+Jr�����
�$X}��3#:L>���]�E����4}�;6u�~؏�>��`qgug'�t�F�;��.�P����'�]�ɩ�r�}fƞ���x�Z텹��or����\�M��w�&!��ym��+�n�\���CV�{ի+�7��*�V�	R�(����M�N���af:�🣡T�Sf�|�V��)1��H�U���6��r| e���IW�ҬGnp�nS��[s5p�)��~��'s��Uh�(�*hR�2�^��Z[k��ʁÙ��h>���[��B׺I�~�cV-_ѡ�M���ѱ?Z��/G8na�����ݨ�O7�ì ٥����A�o4
Y[�Y�l�����V�����`*���h>��Ҫ0����"�d�%���❟�T5��CT��#�����bG����e���i%j0�B� �(v��u<c��}vQ��^�K&�������Ö\��sԢ_
˓�X.p���3��,1r�L�n}8e��B�Q�~�Z4�������t}���pӁ1����,۬���5��Ъ#%+�Y'
� �4CL�1�[��DQQ�vRi	/RD;�����^^i���ķ��7?kj��O�9(�&��ى��b�QԸZ��	�f/u�Z��2���u�ؕ�l^e�-�����˰���E:u E��%���2�ʑ j/�5����X5|�o��i�����K.f\̼!ϗ��Dլt�o����`�#������5��wb�}�\Ζ8�x�?VL��
��5��~���a/.A������x�����W�(�3(�DD#&{9r4t��gǗ���V����S��>���9JՃ4:Ns ��۶Y�[c4`3������Ao٪�+8㙩@�Z˧���(�\��s@ý�%�q��Cu��@��������ҡ��wNKI1�Ik(��GI�3��C��&)�܇1��)�~�&Qh���fZuZtB�[n�L9� ���矝�����n�I+o31�M��n���R�Ŧ3��Ov1�1�{�Nj^���^�W�_�^oG��Ыs,G��J-���i��NH���%��YL�s㐩���H�`��3��P��Y+cYd�vPMd2f�@������<Vm�4������΢3�,�h{D��,]ML���xӏ;�� -c�q2�rI�I�]��4�X��Sl�O(�N�=]��؏�7�x(���	���E{�����g��������3�ƌh|�J��
�i|*~�G0+w�d_
;](��퉯����t9�is���!
��e�2\Um����+��v~�t��l��W�"l#��5�G���Ca?Ӈ�q�p)�H�Zo�^�H:4$zM��C첲�x�Zg��	d���:-�*�Q ��c���A����]U��%Ev�˪����k��RI��$aJ2F�L6W����L*���Z\g�-���{j@�}6,�'8��_�V�i�f��v�m�
G3��i^����H9�i2������@�=� � ߧ.�K9�r�;DU��]~���-l�2��`z���oڄ��n"��`��ң�\ē0�7G�5���d�� `ۨwޤc�y��ӒH7+W9����:P���dj��^uN���BA�. �G�׈�ŷn���;�*a�b�!{�}[�5�WM�q�6` ��]ܭJ��)>#��m��`@�q���`�4�N�$�A��D�����8-ZQqYW&)R[��.���"��Ӌ�@�!����0�ȋ��&Aҵz����.�Q�ˠGtW��?��4�'����M�e�B|�Z���_%��M�z1�4��#y�p-Q�m�lb��ӡ��5ʭ1�$r�|��Z��G�����3������xT}�#�!)�)�Y�
�ڦ�S0n!GW��t.C8*�[W��n�Z� ABGza��jU+��TV׹?:3�,�D4����ڝ�F�%�'��0��lҁ������zyHޡgø���`R�#��X�Oh�,b>�$i17���)Y��3��j�{����bZV���*��^�%��K�M��V� d����3A㠔b
2�O�k��M��#�ז�-��5Dz�R���L�&��"��0�r���5؇^�0�p�wʑ��,	��`,{�2���ޓ�Q�TE��ڌ(�]�����ڳ:\���^�2�h�H���F_i	��n:����u%h(��ԋ6���Fb�n��>��z��n�[�[e�uz1�[�n��K̿�Ј�<��4ri���٘Br�᱇d��W�?9��4\�������q3ȝ�J}YC��cݶE��h�f�=�+������GT�[\�7y"0*����x+S�t!;��l@����Y���~m��,'Pְ7?�;�9�т�q�#�νsb�*_(�t�b�B��6ԇ��R� E�,��S$9r�ZYZYI�`10�	}�{�J�[�_�O�+"�.�I��r:1Ş�.l#�`{S$s:�Љ���)�g�zܴ��x'��^��$Ή(`V��u���R{n?�)�ֺ޺r:�_gr�p�T;��?�T�	�@Cn�6 ���5�4��
A��s��Q��O��@[�����c��a��g|�	�6�FӖ ;�1��|)��ce�Ԛ�툹N&��T�ꪑBM׌e�ד�x�T�W�O��ӛ)c��a���|�Y���1݁.U�t���H��<�z|�W��M�����i�2�_�;�!x�ޥ��'�a���}�B�ԟ���U3^��HW<ru�S�Y-E�Z�K��
t����Y�}Ok�z5��R�U;#�=�֒#_.S�x~9�x0j}�������4d�����H=����k缀^Og���A���-F�_�T/N���UZɯ���Av0��c"�#�N��?������A�°\��ܣ\�=o�Q�ԌfU]^�Y`^�X�wH���P5O�G˧�3)����ٙ�#�r�S}<���<��%y;���Y�v�~ad�"3�X-]Ćs�8�;z�����39�"=z�V��&I�`��i��Jj��~�{	���_�FRKl�]*����e���W�O�.^�3�ַK�BK��@EȈ��Fc(p���Z+u�Z[eV����*�x�;x}�͗�r9GN���;|f��#4�J~���e>;3�Y=ݱ�?�ن�RZ�G�(Yw4ގ�A@���_�U����|6����9���fN��<��D��Q},��7��t�OY���A�VA.k7pi�(j1V��Wp�K���u_���$[�%�*��B��W��p[�%N���� 4� �B~�E��7)"�E�|��8\�B�g9�zg̊�u���x1ʗ��XЂ�{��`c>�	��7���RiM+p��_(�����M��V�b�iq	��r͑�obr�:+���f�%&.�B;v~�H,u�eY���BF!��=��V
���t�k�(�\�X+ї���s��:'�Ş�ϣy�db[����(����O�> �M�"'>w��m3�%�w/�E��DĞC�i�4�� Ͽ]/��t�[����_(3N�3���O3�d�$,�	�������܎m���8�ދLDt_�_Yy%9�uM�4H��]�h���!����0A����2(e�bNN�[>b��A/24cvDS�͛W5Ys� u��V���Hrt���6B��8E7�'41�MI�P��7�"¨:���{_��{9�l7	v�U�1�~�m�8.���<�Y{�m|Dی^uB �h�n�-!�}�� �X�O��p���Oµ�qb�P�ձ�	f�5Z�|og�m��G׼�i�q�"��eހ�*��	E����M�!��6s\ R�VYê�t�9@WH{H�M>���１�}�`�c�9��WY�IV�ƺ�7V�7#�`b��pW��>W�t7�@Z����CW�k��%�řC�IB�?i�s.��g�'0tk�pѨ=�����u4s��w��6ΊV�Vɤ+4��5���A��jAS��(	����!���ӿ+�*��[I�H=���ٴ���42��c��do'˦�����S��	�+\��i�%���1f��%~�?t��z�Z�<��{��%��g	h��L�q���[�u$��a��T�0]�F���Po{~��TX<*k����ˋO�y^��{:K��ӆ�L�Z�ʹpO��^��a���9�q��<�μ��H4�⿕��Hoo0f���۳0�.I������'�=�h*a�N8\}��W�����Q��T�t���B��J��c��[썪ES�NS�b⋋?v�l�!��W�-���A��鱜�jE���)1�K��	���䵵T����@h	.�T>L�M̦O��Y]|�r� �z	+���dbt@���yCQ�P�9�kp^;$��|���,���!�!l�:����Chݰ�"c�{��F<��4s�R�C�]_�T5�e���| �щ�4z��8�)&Lx��Ȉf�}��CS�Ux�R���(�JlT$����u3i�ʟQ<~�Zg�;W���]͛\�h�S�hDs8 ��Y��>�� L(�QI�����|3�����p7Db]>��5�;z���I��y�jk��5�z����\	G����_�a����	����G� �дS����|�\1::L�L�/��a���e��%sOސs��D\3�,U��b{�zc׼��(lx?��=�#5/���ϡ�U����Ƙņ0���T�������m���+XCg^����%z��f���~���Cƃ��}7B:�.���g]AGv����Hu�M�:�"��ʽ��P��)H�����F�� 6֟�W�B-;ȣy[�*�\�L\����4�PL�p�N����0�jJͨ�{-��PEW��"��|fP����	�[��.�Z�s�nü(�1�2��s�9�](T���[wd�lU�����,���� \l�F1�(�8{[1ͫ7y���C�}��}�J�L���^�p������8��D/����U]k��L�e*����`�񪧤|iZ��y,�q�G�l�{6y�0����WX���d�y�D��9�M�(*��(���l7��5�?��L�"�s�3�DJ6R�B���JG�t%�A3X�r3qGU�O��z`�gHT>��|7 ^O{ǏtK��]�"��9x�EUHڏʲ�Xu����4�L�2�u娆����dw����u�O��q���FL/Q�E$g����V���!<Y���/qE T��tW����v�}��P�mH�/�o�#�t<I���6����,���aj�zٝ�-	R��*�����\�v8j*��p%��Н�S���W�F=�A�+���G)��\��rk��Z�vZ2s��i���w9�m#z�z�h�6�;��`��C{�|��D�P+O4����1~�x�y�
����j9�'vkvĻ�+�>�����)���u��^��&�P&�=R8f�4������r��T�jʂj$9����4��U�k���Ϟ֍�{�����c�E�[Ie��~�� ژE���W!��F�mU¶)8�Yba��H��=�,{l�]�B�^��V'چ���A�CF"�M��+x����]z�0=��}=��T�D�}�>�A�Ї�f��`'��'K�f�cѸI��`5H����� ��r ���:S�s���!��v�=�����c"G"�:�Ji� ƛ�e�g��*�C���Tsk�Ě�:�)'�4LM��r� ��d������o9te-��IR���Dc��vl��r&⨱�Aޛz���ú�&lA����#l��}o�I���{�j�m^�V�b�.�ޗGe[pKlVQ��d]i�:�3m�E_r�`XPS���w�0;�w������c]�8Gc�k�[Ҥ�^p���s���ӯᦂ�F\육~
K�`�Mm[4�6{O>���6$@0\)���d�Ɉl�#<�}��a ���[:��#Å
*�I��$�a%��Y �,k6����R���ؕ��k��t8�Y~oy��k�1�W(#�sI9��D������?:�E}�k����#������k����$�C��D�+�p�c��^NQ��=��a�Z���N>�Җ�������/^��~��eB���X�݆	qI������e3���H�.�����Դc2�:���}ZUT̳� �hc��˖�y���y�;z�j -�\�M.|�w����6���,���r"�O�;2B�[����Ѽ>y���N0s)����Ѩ�O^�5�<_�m?,����H.�.��`��^Š���E -Ȏ�7�5H�U`?��?��o�y�&��_yZ�x��g?ϖ��j��q�EE���/pxlk�?��X��o�ǆ�dҏe����F�����B��'wJ��+� �ӟ0O�aҲ��u���,��D�A#\U%^��By������6�[��ZJ�=�#i�x�Wq���ȓ��������w��nC����BF� ,�w��/�F��'t��ع�J��ӫ�e��a��^OK{"1��mY���D`��Hþ2��z�˨�P���b��;,tvS;��^�`mU�s���O!�a[i��i�a�˽�,CD@1u�@W�)�Ӗ��/T��M�w�w��(W��.f�t+�K�D �ML�1U6I�����߻�%\
��jտ{,t���!��lMy[ړ`0{�e��W_�(��v�G^�ǎ��*�3���߿�k���3(�����4������sQ��Μq��ڍ�d��s�����;�I�vd�
Z��<�Ƚ�w�4�B��Y����$U��
�W����O���v�"}E�ĳ$�gj�?�D���*<��s�L�o�'�
���wM�%sE���s��#4�'���8�%C���̟�xM���H.}��S�du�ʏ*	S��W[�q��)@�V��=A��5Z�8���0�#.�
i�N�reD䫁�;�%m3A�7������g�v�їbMY���A����4���D��sR���<ݷ3��K��p����r�?���>�����������&�I���"4�j��u�/��)�!}��J�T���6L�qa��.V��i��I�eNt�Ģ�. U���3�^Qw\d�嗏�{	�j" Y��I��E�������yV�61e-P�2Y\�Y�%�ч���v�"q�S�����r0���Oh�^v�u�.������[�$��&ǖc�	&��*���I����D�5�p�]��V4�eٖ
�L7J����+ǽ���WE�����t�f� h�{�k�o
�HKU��V/����-X3��U����l�@ғ� `�~a' ��<��90z�͚ ����@?� mK��5#X���-�>qO Rk��-D� �i뽿Ɔk ��Qv�2L���V���cA���"se�oI�D��7�.��O9
`i�$]!#�fag���0�5�s����P�|�e4��c�����%�0��

�^y6Lh��l����z$���{�,�Ջ���[��5-f&H~AE�kVV_�6l:Ǩ�]\)jj�d)F@�z ɸY-
�xw���ۤ�]�y�&#�$]�*?�mR�5��Ö"�t1d����!�6|
8�8����ց�������&��s�W3/)�}G��LN�dڋ�{�#i�,�4���5y���T�U�$��M���ED�nT0�誣��O�lf���T���X��ڎ��uZ�TSD&ח�ef��6?��o �R����&����<W�*��ɿ��mAoOqD�y�|�B�׵�HM.~��X�T"G�8�j/�c.��Y�J%�����a��>�1��QR9�]���_��t9���U����z��8�΅:��H��4�f3�i=�5��]�� �~�`��#	�)��Sُ��F/�3#��U��K�>�@����������$��}�}34���L� ƫ���T��=������a���8G�j|-ά�q�x��s�/���i쩧Ujb� �"L�r��P<=GԲ�����؛/�|�]�r�nj���@�WA(mnc_cu�P�Q�z*N/��?|b�4@1�xC����:1B�G�~�у-/���L��t�H.V�c�(@Z$����W����*���8s���?9C�������%����)}r��\���Pz_N=��7OL�x^�ΛgÞL�� ��y,㟀ˁ�."@2���@s�������~�*�?�:�iC��s�5[d�"��~��i�KY�yʪǪd���#ѾN�lٳɏ ��Z:���.U�d�Mg��}
���*7*��O��ge��a��Nm&	�L@	��(��=K�eZ|GD��2�?�6gKt����y���A��o��?$N��C�DrFr���:o#�3�˨r����R�l�~��rDN�+Gat�����f�ċ�[��mՈ�ͩ����*�|l�4M2�������>7r�a�[ц�Z#᭄�Qq,C.�ˠ���Q�RH��y7#�y%��o%{��j|���bb�G�>���A3`���j$icJ2�i���������(_�<��m�U\�)��G���Fl#�k�����I� ��\H,��r��u�	s�����,�������, �����T|\��\D��}j�{̼=}�Gh}����!A���V���\Gդ6I\Y�i.�����(r�ԓ�g���B��ޑ��ҭ3s;L�Z�����)$" Z��64��}�4�)roo�D��t��S�-jt�՜���ȱ�Z�2r�0��U�Bs����2�Ay��P��<�=[��8i0n�n�bJ(���m��ڞw�4 8��Qf)���6?�#��^�, ��S��-��kJ0&OEXHC��[��}�(��܀��JqG��o�n��$O�͑���ID�!�0}i�G��!�0D2}S���j���Bt�M������K�4�ŏ������.�Q20])��A��Կ_bR
�}Br R!�jT�%�P�m5�� u|�/���@�K���,3�w�6��hd�@ܾe���Z��O�,�4R�L�[8�nb�< ��H�,iaq�񑮌p����6�y8��<���I�54��Z�֖h!�HO���ч� �I�� �]�uAm��x�I0Y��+f�9����'��}d�A�V�q.vY:��
P=FFǩt�Pin�*�:�o�?�'Xa
���t|r�ˆ�YD�܊����i����N�>�c���oκ��v�(R���F
�����J�g6�e<�U�LѰm5��-"E]ÉY�\�wuw�殀�^Kn�����%�޺[�3;:�|�{ �WL�F�|]_p�I���D�R?�P;Mb�����]�M�I�#}~V�d9,S�h���PU�cuއ
#�,BM����W�mm���{������d���Mlo�g�@vQ(Ŧ��~j�^K߿�H�6����>���v	/r���%��e&0X�9��җn�_�T`a�:�t? e�%�~���I[xw�R�����^e�3`�$�
(��-�� D��?!2��O����������ak.V�-��U�-���3�F��G;�?���̐����?�[)��恇*����^�"B�����ݑtY��Ŀާ���2$5�3TTe-R���f"�Q���-�]��2\�%=g�[�����y⯰��trFF�Ѳ�So�O1����ao���Z������
T�p�T�F�a3h��_7#@��P�� E������k��t��IL�c����gu�hX�]N�UaeX?�rh1�h��g;Npܬ%�;�=Q��,�Đk1!'"��P����c9Ke�h��|�#���9(�Klxك��y���(/s�y�ǍW�Z��[c����P^L#J�Р\�Ӂ�G���Q����Z��DC���n�8^[fW�/�Oj �$|iyQv=����~�E�a4�+'����<eR��bbsxW��i(�9���Y�����[<��p�S�$�{�/���E�,T(�Xտ��p����o���7*�O�ʴ|�?Ow̻���7�T6��Y�%'u�sVifь�U�"���m!�.X0cA�O�9vudBj8���]sW G�N�1��B���0n�C-�i1�G*v㯄~�	��֙��-������-��qH�![԰M@�@|��_��Q8��5�x;ЁD{�0���bs �+B����Y���/0��-kp�!9�#C�Y2�(�Cx��+�&�Y�{)�M6�+��`Z2�3�r����>
�������"q.���\	^dSn�A�TS���?O�������؀z#��Qa�W�>-�8t���N�Af����YL���C�V���R{��`�Wδ��@��>��@�n��,Θ���
�+I��ɧ���bR��**{�A<��:����,����5'7�y���}k$��k��0���F�U�̵��|��,U�.{����U��[�VVzCJJ�#o��s�� ED��O�7��H�B��L�l6��z�7e������F���b"�8�h:IE�	q�#EX�('�7m�֦�����4Z�;�v~x샓�y쫁���ȣA�L�;�V?O7��G�IS��n��g原�?�-CDG��+T��W"��|���}��������N-�l�^aF�*l<�q��ǼV�/�Il׵��udH����\>
z#��vG��j���}"��X�
q�������Ab��4
���
��C���}[�3�F5��̩�!��?�#|��.�=|M�Rc��k|����
�����y����3eGeǊĳ��~� ^��%�vv+��ꦃ?D5����>i�g=͖̭��*i��T��%4��w
�-�b�V*�ϳJN�i=1��902���:sU�E��Ee$�?�U�����=|D�>�F��|�vq�=��:	3i�������x��fj�����AFt��.|]Q�Kj9�L^�@�ET�W"G��H*-ޟ�wKVR�/��YI��C<��n�V9|�zD�S�Q텙h�g�{���ʛy�*$�~�_ٻ�y!ϮW�
�IKh��q!jb=��v�`S�Tb ��ԁE ֏��L��U��_&;�M��P0�@�D���9��b)�'��Cd��S�@��� !��7����ƛp��s@~�Ѿ��w�`k+V�Ԟ�<̰Ĭ5-@jՖ��j١����/�	���{��|�r,b����`��Nr	e�����6Y���_G�s�/�OW2-n�h�:�
�$�}�2'��~��$<��g`$�i����Mq�JP���������5=�0E��5f-,
����x��
�� 4
a��;��,ޖU�ېo�窒-9ś�1[���E ��~��~��ɶŊoR)1���k�:�.�S7��<涞��I����$C�A����Ay2T�9W»[A.�D��,���HFcM�Z�y����t�;�u�����k4Y��J1@���m�X�V����� ���(��L;qA	�^��9��4�
�V��6�H��2�Ѳd�*�0˧L�>�^Pf	�ꫪ,0w�t#�*-�]�2qG`hՙ����~��#�.8<F�n|p��޼y�,��Q9"�g1
�l�d_����W�{@�̌jKV�j(ϫV�`A��'�㧨ҫ���J烟�j�q��^��HDh3m�1���+5Y��&AL���&(cE�H΁:��j��[&xu���3h�~7��{\��-��z��׼�6R�r>O�I����9� !��QULn��j��W��*�r���,����60���l��i<�Z�����M� ι�bt�R�i����C}z�,rG4��)[�U'7g�Bl���(Ҡ_��n�ذ��b�`|��H���K:���܂��� �����lZ5�eܷz�	!,@���98i�7{G�UE`�UV�ѱ1���]5�pe�������F��zٝ2�-���"V+k(��8�6���OW� �eLK����rߙⱮׄ��A� 2���������3��)��O�#��S㔪�o�ֿ� �����S��L�*��E�������HEb���B:���/�ш0&�E�^��l��:���o���;�S	���]	���K�j�R>�M?!��9&���`��r4�`Y�5�i.�Jl�|���iA۔��M`R�]�ȧ��q�Be�*s�Pu�-�h�,)�@9��/$��r�#T_kn�8�;����䇰�����4p�kw�Q$P����w��p�I��DB�q�'�sO2n�ApJ���+F�}/�MJ����H��ލj��S��+�O2�(Bm({=�i�v/?�b�$����x[9R;:�OO# ���W�ـc[�d6ik���%1Os��nLky$�H�`Hґ	�DlK�@�Ek�۴9 3>��Ǚ��j5��.��/WU�Z�pq�1U�-�{��2�����9��"g1�fZ�R,�v�I9-��S���&%��^4@�sf��qҿѶQ�%�g3�����-�Qt�d�p� �]��8��$�n/����$ÑԪ�Q	��^�v?j�D�q9�4��$��K���R�JX ��=�V�<�͟4��g7��TR1�z6b�eU��߂��#��;��0���֮�LS�|hL�#}�E�l}�)%Ue��C���5��Vm
�q3w�p^]����� �ǋ?��a�0�Y�i�E+����"9�0�S�SFrs4�+'p	���(�Z���W/ㇻgH��y]P�����mxl�YN�2���{��*��ɼ���M�]���Ѱa���
b$��g"#�������1lRB$��4f�U��2����O�T�1sb*V���R���Wf��j��B��ViR�X�h���0�0���ч�2C�7���N	�G�=vJ(:.ڛm�|�/��n��Y����7)�y��`h���uyR���O��E��e)�,��gpٕ�l��!�B�B./?r��@	d[�e�rV�n^��H�৒�@�����&��X/R��3�(s�:w�fH�ۮ�]���4�x�\��4k0�*ղR6��O�L�� ,��,	+�젖���m��r�n_�>ڄ3��XK(��tF��=/���["#Z����෗c8.�`t�А�`f�Mܲ@%�s[��ca�ױ�xNɱ��l��	鉤ɀ����1�v��_N�:�70/�TT�70Mz$3�<� />�4�/ly���c��3 u5�ϯAm?
��3~�����@	b#��O$FSP��Š�&}��i�<�_̢�=F'�!N�$@CV��\ԍ��ٻ�� ��^�^��W�%)�]���fm	�&�8���w0˚��
�"���R;�5��˞�P.����aw���L�������Jq�^V�W�����NK�7�o���ڵY!�VX?�/������:/S��.z�(O���� d�$�Io�����G��u1&�I3C�X�)Ė���#o�s���L�ou�I�/TyX|X�>��U ���e�\Er=��E��}�nB6xA�a�@�~����C �X��5F�����<�����%Y>��P"�Fr\$d�q�r�+l��8�|28��d(G����1�P�(Jp�]���Y��Y�O=ԩO�6���(;��5�������C�F�N�s!�����XӒgٔS7T�PN��:�����|�X�e;N���`;zAV���I?�/tڤ�f�P
z���0�������u�j�a���#�V/��H�N)~gf`��U�:s���v��6���x��C��c)�����HJ�"�O2G��!}A��oE��4��dN8U�m���qฤ�q8K�]����Č%��O�%�ֱ�^@����*�&4�B�,I�6ۥ��%��u�1����駮U����8^w�b���e�wh�"����p'ho|�0R��W��K�}D$*��~�+
�tQ�O���N�`5�(Ԃ_%�{~a:e~�UeFv'l��}bW�%,�1"�<�vfr|������)�lK�Qq\1}�'���?Q q��+U"A#V��)ު�pYM����U;	�F�#^��RI�zҠY�"���+�fs�ܴ�� �rl���+x+[��r���'m${���̲tR���n�h!@s��f�/����b���ћ��"7�á�#��{5�!�:�D��>�9�y:o.r�W���:.�Gl��#��`�x�'=4����c�� ᅬ.è�7�/��ZA��V��+>�p	G�7�?�O��94+�t@����@S�I���,j
��|��͟X�70��WA%���=�y,ث��_1�oB
�.��O]KG������D�$B�	e!��} �ˡ��2S��Ok��q��2��L�y�������aAzGr�A����]7��%נa��� ���C�������%�r)�Qr��g�7�J��k7�)w�FB}n��Y�e��]�Γ����1YM��/oh���'q�
�$�%�m�+4��L����Z��u��-F2>w'�%���֣���nx"��i)��к?�i���,}��5
�)����{�1��A]�kOl��(y��@	@9���E�';���	����@�eI��<C \�ʰ�߮�i�,v������k��ڮ�,1��o�J���f������4«����Z`��7�\!>Q�z�U�ү�K�f�nW��� Q�y�dK��~_A�W�Ԟx��F��Ԝ�j��τ[���1d�x>G�؜�3]��l�߻�K���o�mR�	���N4Ā�uAh:�E^�z 7O�����S��OBZ��m�	�7�����׮��7e��
̾�l2D�BK�%����e� �\�딺*R�T��p��Z/`��d�2p���Yb�S�9�Q<��`��˂O�2��q��PM���@�3�,R�
��ɹ1˷�|�����"A?�J�4@��ݣ��#,�8�3'V۴Ӗ���ڳ�5�O��L5����m��A�� Өh������T�#��_-��aõW!��M��oJ�g"vɛ���P\�ؾ
�dp������9mqd���b�sNi��B2�tX*���ݜ>y\[���8��IC�Z�@#:bAN�6��d_Zt��4�P⚬�8	�j%@�S��{��^�,:�-yi���Gj�f���[�5c��!��8X��ૌaP.�s�=B�OO�h�ɚ��R�'����-�����Q�{)m<����7	<ǟ�w3FYѢ�]��&�2|�
��0(�:6�~/-���Z���3��,~��\'Nt�m��@��iW���Q�E�=�KR�y�����Զ�)-�|�zUU�?��y��n���Kn����3��M���@��ɝ���>�&O�q�/�ݟ�PGme�{r��P����`����;+<u? _�;y�f�Eƶ~�6�K$�ʭ�A�'l&���踕b]�Uz#�$F�<�ؿ�ʃv��K���r�YpX fg=�~|�
ۼ�+/|�xX=t�񟴔o�����>�v�zB��P#�P����U(���̻-�X�B[3���+��[�qQr���7��}>�uc*EL���F�)�17þ:d����pZy�I52���}^�# 9NMI�|?'���������E�_�K����7���ߍ�xӌ��D��s�\���W!+��	$��@�X�g�ܧ���Yq���o������)�L�+���b'�Yw����GwnىXMJ����94"��P��)�������%��J�v�����D�uE�Ϩ�/���ʯ�v��=%�oU;_4%NJl��|*��8��׳X��v�ɼ8t��#%�Rq������a@'t�X�/�R
Ttdt}�'愠΃*ZX��3���`�VQHBY_���-¹��c������_���<jO�9"m�r�W�	� �?�B�㎚�)���72�AL>1A�d�F�O�X�.��d��+�F�{�U�r)��{_��d���;���Ў)#j=�ds4Q$x���;���r�LT���*�d���G��\\��$!�i�9z�CL�@�&w�A�Z��!�]Xji���Sŕ�eI��_�蹫2_��aMv������? �q�X�t�~s�!�\e�8��gm��]�T��ƽMb�x�W�}5Ⱥ"=t�I�%����&V�A��@��i��x-�op��ݑ֑���@�VTT���z?������|jN{�վq�b❦���b��3�>���:3/�Z��� �P�=[{��Z��{��}*h˭\�|�}X��I_08u�rĈ=_��o%nv��U��Z.�mj�����!�^[v03�p��ɨn�;�����;3��4'3��z�~u߲��7G�Uw�/��fS��k������~gك����f U���ʎ��1������zW��M�[�;�B�ÓE)�;C�PV�2����u�l+q\��`0A��}��'��n׼
�T���-�&��֫-�c�%��>W�p
#�]����
�<�_��c��N&�#�Q��j?�T<���/v�40����U���c	����bG��b��A�ձ
юy�]�RƜ�kRZ��2Pa5��x�������1���Q9�g�^�k�y!(���s�M��~sVuc~���\)���H�#��б� F'�����S� ��_t��6�����K� [�7����E��"K�X潂R�u�y��D1��YxEcSX�8�6C���{>�`&�4�i�~Pz6��ι/�i9b�����˄{�-H�����@K4����c����vc�_{�I@Z�������SI\d��rӂ�6[bE�>aDڅ���F���|�� !�����fx[t�G��,��K�6�����+ �پ�����Zs���u@y�V�N���gg���}�K��b��7�x�0'!��]� ��^�h�ʌ�p>���w6k�P���$R&M�å����k��q�Q��h�H��h�tU��3LuN�3ٵ�3�v�N�'�Y~��O9=N����[�%�~�r�V�3c��鹅##=ߴA@�׈�	e�F��꿕Tx�KS����7�y�į�dn�s����/�¾��jקL�\c�w�8 t	��ag��I�9�@)��������I۲�S{+f��$�"����z��PTU�<����C:CZ�Nl��u�����0k���J�n=ar@'�>���ZtN���+vaTA���F���_n`+�JY� iǸ����a\<v<i}�x�1��������4���=�C���� l�����S�^O�C����%5��ㇵ��/T��'Y���D� ��)�\�1�-�n�Dg=-�ׁD���CA�Ev����j=EaнW�an�5Ď*ш�~�Y4�����~a�'/�"%���N/��tt��s(�Pp�ӂ�GJ3�ַ!�Ņd� �L��ﮋ&G��d��}��p�gAF{�,XU�g�'5��!���"�����m�U0wW�7�]��$yӶ���N U��y4��GMn('��lB�6M�szF��=��2���X���S'�
9n(MzΪ+C@��2߹��;��GdM��6���� �J7@?Qw�J�s}�BY.�a'�/qpq4I�����Qt��+I����cS�<�Q߯9��e����Pܱ�� "�tQ|�.ʳ�����i��m=��� X����`G��t3bj>�
@�K��{T��`���� �ݶ���[H��Ύ�?�%^���&�C��F��z4�R�IJ�ss���W"r
��A�[^��x�\� G$t�[$9��o��䎅�y�`��Di�ǽl�
���7�c����j�1X��7��FF�����$ٳl���2&��=����W[vw�x�&�1w��|X��m`P����\�������2�*t8�=�:j�3{����N�(�I�ɡ�$�`�CAixe���ّ�9��?�(������P5�ք}��N��RHƓ�ׁ�p�I!��X����Q6����O�oSf�zi����h���7�[�(��u��-s�Z��m�}𖸈� �:�IK'컈s�����^:U��������f<�ؔ�Tv�d�@Ah��J�y�*5���\a�'���+	V��o�&0f]�-���ԛh7R�l�~gG���R�/��*Hd�a}X��֌0�in��M��\�!+�y�}� ���� �X�b�+�3���}����7,R<~�m8��K��U`A�B���2���^i�I�*����4��5o�Jbf�&޶����+�,���|6��2�1{���A B:0Y+�/n	��l�{�5�x���)�	E(H�.�U�~��v���95K�4�ˆ�Y!����U^�T���i�vD�{ɢ�w�!5FA%������:���a��'y�I�V�i���i*�A/�7�3ɣ�;�&�ih	�j*���H�k��heZ fO�Bg�L�|��T��ܻ�#�]�59�jEV���g�=�<���g �?�YWU��43!�f����_�Ug����T����j51�"���I�`9�Z: �k<�9mҚR���2���*�w��<[-�v�1l�o���|Y����╜I���Y�2I��#�x�c*�U�s�'I|������@���2�FHb#O_v��B�VwRв��+��
d�U�敷$j&0�	�v&�O1\52T�F~�fv��o�N^!CxsN��{���a,��=�@����	~@]ߘ���ȑ7�@���6.�G˝�7݃c�R�:�¯���tEҾ���*�,B3��5+�x3
���x��O<;�(�"�q����|�Έwt$�������H%Q�:m�Mx��Zr�f(�L���8�]��L\�=]�� �D��O�hi����OQ���u"f�{P{�cU���`J�B�Nr�.������H����ﳍ�'�n�c"�L�dP��A��d�?���������W�N����5�@Zuu��.���s"���i���]��"��!�� ׯ��v:Ƶ)��4���<��E;�_�Ԫ=�!?���<G0Q ����ʖe�?T����q��_6�4�Gq�
���A6�0v#��S���ǭb��jĐ|}�.��bS���aL�rχ:�%C5���F<����Uc����ѐ��3r��&��Yw�/�0�i
[϶�akh�}���֌㣾Nk�5CB�O
�m�ͤ^5�S����gN�T �m�;	�]�H~6ϝ����EZ�M惍�6s
<q�[�b謥o���Q��W�g�j)��"l�.z�p�~��+��kcs.�u5t���h�|��2��mD�a�aΨ�J��3S�Ǭ� ���/�6�W3�;�3��%���y����	E�YL���+���\tRZ�
���$�ϯ�S�7�Ym%�??����A�JW�ꈨ�GD�q�k�5Q$d1��������F�=����5�>RD�fO�*�6��*���8�8cB��)Prb^�r�����w�T���?�泬SH�Y�eo�{��P�N�SI(���;��CH�cR�� �o?L����n��p+�~#7�	�~a���
���aa�-�s����jg��3�Eb=y�T�S��<eR�+�sr��\oO�f+l��h��{w���S��)oPɥi�_7K3��GO�KgZ�2����V�qk�o�A��&KhZx��ވ6:�U��6�;X��n&� ��k�='$0���f����7t�2R�A���~n���w}��Z;�!��w��!�_U��&�W)�g����GÁ����k\�G�/���:�-������15��D%�	h��I(��(��Ԡ��zO����r����тZ�z8Y��7W�F?��Y��bD��Y5�s��s�[�D6xH�y�j6�����
@��mSt"��5���i*���4�JE���S�ꃁ��b7:�
���mr��Wg뛇�s���yo�ya�~t��w�Q֤J��
������˸�2@�(;~��ң�|��_V�8b�	�rI���N����m��)#�}|���9�����ȂF��o'V]j���ڔ2!n����o���v�&�U�&�W���_Dg,�i6����X}���>��Ob
�p&��1z��X�>�"�|�����A��ʍ�� ��>d�� ��]v��"��]Gtz��x��ș��g7�VE�[���V�4ACP���7�m.���v��0�˽�����;I�+1��+�!��H�g����?�-�6�_�:f���󂾐@-�o��ڗ*�4.�"��
BY�
d̦�����LG�ذE	ԧ]$�����8`����|��!!W���k��3����%�Rr:��τp�`$�y|��e��O�<d{p�4Q�
�AZi9�mR�0�����s)-���{,㜨�y�d�b@�>�����u�@k��ƛ9��X���cy�ֲ�j"l�h"��{�M׶�6��	H��Q��ԗV]�U���)yX�Mk'�q�{t��M�Z�8J��`�����b������/�����o_;���QI�Ha	va#��x�����*�i��ۚF����$�"ʱJ��Y���������6�;�^�͔�W������Q}#B�V�6�ƨa�+�DE�5��.,:�K���8u�M�2�Ǔ0��j��ϷMe�>e��.n�y=j�Úa��,�n�\Q 
��拹Rke�7 eE<b�z6uϹ+�6j�>��!$��>B3j�V#uS!�C��v��c����O���s/��{���e�=DicK��ÿ����WT� ��`�[Ɇ�KB0;�̢42*'�td�t����yxBQ�DD�$���njAs�`�P�g�-�j�:���1}����T��u���7��1���~��z�j'>�RQ^������7���t��?Ks�z�E��m/@G��!e��!ቾ�^�	h��y �Dfj��ɧ���H�P�!$��S��
��29��T�&�l�D,
$Y\C�2s��-�x��ϵ_n����.7k˜��q�pB�����dU��I��1�t��럘�~�ϒ���.��e]h� ��E>~�?���k�Ϭ|��P����J�!�����aY���:��>�	.�\[Z0�F�ɭ V�Q�� �6K5�T���H9����Ew��nI�d�BA!�OD����w�T��MGm{�a%�n��RC��hmM�5�ǅ��d�댨��yXVV���g���	�I�c�1�����l��l��f�̍]I6eI2��ymӜܶz7$�Ϯ���p�US�g�p�D�f��ڄz䣄K�5��+��A�E��Vv-�����S~WqZhC��	�_k��,��hK]rR7�c��1�f����s�P��q����3$Bɢݓ%��pWB�ݼqCM1Ͻ�����d�]h��證Ç��զ��^d�a��7���3躂�B��ia����먻ЬRva�zK���y�� �JoP8��E	����ǈ|Tc*�	t~�������Ȥ��O�)�nd�{��������KN�&����+H�ζg�[�׆�\��g��(����LD��˩1�อ���)9���%�;�AA��)����HK6�(�K^���+�("�����k9l���{�Vg���|���uĸ엚M~30w\��Ǔ�	\ϓ�^�N˶��}F�TZ7���C4x�
/����e���k�Ս��~�[�7�1C�;�//c���'�_'��{�#��Ac���K�bi�xz&��A5Q}�.C,V޴�yjIK#bknc񛴽뫜*t�}��П>�-5�ɻ�z��D��Ե�!�CS�u���s,(."�`)*(�;�s)=2傜Q����4�����>����G�Ӡ��,�s��o�����D�y�
_<��t�������=ι�n��Y9���{�A��U�$W擻C����߰�g�s�~���W���v���;5Y)'ɕ�~eO�HM��\�Ȓ3N���o9V�>���W��9��s�����'4�䮢}��v� 8�hHB[�cô�x>�����NA�;�0��IȦ=�J�����o)eA J�F!�(R�T??�5���"��u�Q�R��c�\��yr_�U���JAK��(�ҷI�����B�ˁ��e7��P��:�L��]͢*���0Ԓ?�.i�A	�Y��k��q��f�cZ�y��7 ��tV �Y'_:@6�&t"�,X	��>�Z�Q�)���L���9Y�I5	IA�㏗�L���� o�7�+�ȑ������	70�~�:��U��� .l�h��úT@�G7Q ���1zBA������HX�8�(�@_�=	�1�ɪ)�,�RQж)�����$ �FO@��������`>��/�(aYV��1fZxm�E�#ɹ-�pzh�0?�zL���K �n�-��[�d�N���7��`��% :��hqH����!��ގ�B��Z�-Τ�[Q�;c�|� ��u|�Sy�؇?OJסZ�����9�!�4����9���RkI�v���:�G��Ȫ�9<%�������ru��j�ƫ4!H3����	�>d�U�Pԩ�6�&S��y����`#�F�9���.4�֢N��]'^�l�A���Ŕ\�8|�_'�:˦\Va�z�xR��+�h��`o;"8�s�\+IO~�>��F��.�OL�������4���r{8�K���Jc��������զ�8y��6zO��9߭��lr� 2�z"K=_"���GEy����V
%��kfGv��Y�܂���7|;��:еr6��TJo6;�p��`H�i)���-]�o��<W����Q4ۚ��;�&y� Qy&����ry�����'1�3������.��2�Sh��k�;(�_�9ʀ�OoaSΥ�:Cr�R��9�;J��ڢy�tz�]�d+dv�o �o�FV�����+�h��؆�@���M.��z6q����-�
*�5����r{��|��mIkg�f�Ǉy�wį�*��Q�mEא5�Th�3GI��N�p���ӓ<�Ԣl��^�k�8r�ހ{��!���9�h`_盢�ƶ��z�D�A{��B���ǰuS�8�hj�25Ѽ�康*�7Gki]_BJ����$�UK)�P��������B�W3���uu}ՁC������ 7�q9y1�?�>_l��e/ۂ�`\p�p��^۵Z��~������"y[�˾��I{h�Ł�NG�-}h��%kS"`�-�b�C|8���9\(��h����	�m���3��SK�{������l����e)���1��n-�P�-Zl�h�v���N	)sAh&�A	Yan�X�lGu�Φ(���/��?�~B�.a���{��F��8�M�=�9hp5:��D�p��g���T�����F�8\�����87�邡�j4�C�5qLq�~>�aWEψL϶No7�X���m�fi��ƍ��a`֪�~|�y<G'���$_E�f����x.�{*DNb�#(9�4����
iq��*o`���{��=8
&�x�梍ǹ$zW�*KJh���0#������\�ՕR|�u�v(�Ώ���\�:)+�ڋ�k�㼎Rf�$�<�?)�a��i���)wfh�,uuK��o���=��M���T���N�����& ���& i��;�b��L��=^Ku��nf������2��m{N8J��R��S=�6��=�v>L���)E p��W�U,8�����U�l���n�Sf��YL�z�_��mҳ�
_8���Ķ���|��(5d#�_�V����W��P�[K�Լ�zŎ{�'U�Pdy��Т�6Q=Kk۔�W[�Y���y=w;<֌����y�����������m1{h9T�Qֺ�\���L�<�B�2&�O��4GY�޵�c���'�˯b`�_�헬ƺ(��-ۖ��
����%�Cxb͚�:w�]c��J+�(qd�ή�|��i�+�i�v�zU��F����8H�M�+<��e���>��I���-ư� Ы1,m�g������j?�¿����7����w���pB��O��,��2y?��+$Vސ�R���|\]x�V�_�z�@њr�� �J��}@�5&s����>PEσv@z��`<n�b�p��"W��*��z�H�n�s�1�Hr'�x������h����O�a
�%�Acf]`��h4&w;�������zX�<R㏇F�~ߤk���Q�Џ�} T8�"ɗ��/���HE�G�o1�(��I�\���Zb6��<�*E �#�i5:���Q��th+�Kр}��v��Xu{�~�}�,£��]:WcJ�>�{�sq�>�s��_7��T�Q�;�u3��O�E�VjM������,�fy�G`3��[�n,������ך��3bP`�# n8�h������A 4r�[bg@��?� pF�st�c��g��-͝�s�x
��#T��۾�vD$b1n1�L,�Z^��#r흩�jL��6�4���t�!|K���62tB0~�L����̖'W�i�Q�M�SɌVE,\��@���D�9O.���=��5ߛ��+�L��'���|֋�E�?�s���GBzӋ�u���!7Hk��j�x	�)���/	#'���}%B4P��y(_*HS\�oh��}{S�݈iWl��V뽢!���<A4���q���6��jxy*���2qjq��IY����9}5nJ��1~��EB��x�����u����:�{aμ�n�E�v
T��̐;>Ҡ�gN�O,
	V���1��vv(�u���Bk���%n~�z�s��v��2j������y%�z�� �������!.����P;��,�⋏�D���.��oaNn���H\�5��y��By3̚]qv#���f����a�b축N�q���$P?s�gM��6�yj"��m&lie"�����4]� �^�t ݫ�Z*��,�Cg_��(������Q�΂���,�1�-�����V��k��(���8�'��e���@�.~B��Ʈ ^��K�`jewB�y,��1�������C����
�j(h�k�>�i���}���څ}��x��WEppl��&�ž����i���'!<�q��@���������/,�x��l,���6frޢ�:]��u/�^�!v��ʎ�,�s����U�@E�TL�߅n��za˘�l~���ګn��"z7#��r¬�DbI�$r�&��%���|W�AZ��-��4��'M�^�5���[�c�^�QFF�)���4���~g_��T��vP�M�,�{�.�Rr��O{a��z����5۩��� �����AhUq2s�W�*de&��.�:�n�>0��Ao��FⲲ�Q(y5��J7 ����~�b�y�����V%���UK1�>�>:4���{������ ���a�[��	|��{; w{�S 6/��ه��a#�^�$i�����_{ �-��e��D�+�*�
$�m��h_EBh���
����5�'�_�؆M�����QҬ�e�2�����R'�_�s�tNLwz�=�N�O����j���}0-���8��Jf������9���)��"��í���?~��jQc�(��e�]�P�Cz̸`asY���H����}�n��;]j���
|�Jm"�t���8_=�7�m�Z�X	٥y���e�[m_1\�{w0)?ZF_*W�l�hJY��*���e�Ƶ�:�������CZ6R��E)B��G��/i��8�/m�ef4d�!O���������g���F�^�{�"�8�"�Z�W���;x�枆$�\�W:��h=�8z6���6�m��=h��|/7ǉ���~����%�ް7����9�[�H�Wd��v���a��9|��}%ɏ��B#�m�G[�d�1O'��|���l�b���c����Y�υ��
�������;���k���X`�N+�`�H��\JE���v�f�k�7+|��+��
=��=�?|	U�,�8���`���3R���z9�V p
灩��M�V�������<���R|�ߤ��G<_b
nt��M��@��R�];s�������d=-x�'i} tKy\@G���T�6T�⦉��7�5�-jj�%�WkjƐ���Z)���	*H~�X)�R�;�����{n���]V�HE�[}����"w=yݲd��Dg�OYώ%%t��	�\��.|�H7́o������9��z&d�X�n�������,����/9j��(�ı��/,E�;�̋' f������O��O��E8��=� �&۽L_��S����Bm$����������� ��r�8�n�K5ԩ��-='�#`O_��&�`���]y�&����fgwg1������g���	���@	Yh���O���}
�G&%�řⷾ��m���;��!�Wٯ���
j������$�t��u\�y7D\T�#բ�$�d�խ��rQd���TFѮ���G�F�+�����m���Ʈ[�~$���(�P>V���5}(#^5:<-J������h�ۺ��}��`����v���%H�e���A�3!P�U�Hx�x}�q��[��'$��oZg }��J'M�«��/;���\�>*�����#�� ��{Y��hv	ϼ���"]�5�
h6�v�̼
�=>?1��f��2����ڦ(��f*I��f�I��+���"@�_��`���c#1�����&,(����t\l��f���Xn����rm�M9�:�#��6]e�֊�LY�m�Ro�ق��^�Ŗs��m���!4��me	o�$��8���[���Ua���{�yc:��o�,K��k�»��-�2_�=ܐ�����nR�[ ^��C���C�:1�ǵGl ����(a�5f$��9�73��h�6��$a&�'��D�¨x"�H0���4*������G�4��fƱH��>j���^�t .A�!��v!�u���e�&�+�/^��k�����J��G.���@��7:��	_TAD� ��H����9�x��j�|�;�i�G[��z��b#m���^cW��'s�S+�e[��#�DK��}��Ɇ�|����Jh`M	��TV���5ys�D�� K|%�ɳ �tj������[� �l��u��h�F���`V�鴅�������%pC[ ��|�y�>^�_���E7�g���߃Y�K������*�h��f۰����s�`0�C�l��&,#~֌��Y��A�>�ӥq��
��9���^tc��T@N�㰒��O��KsV�
�����F�l� o���N���[]v&��y�C7۷p�����-�0��ʆDi��0x�j��~���@�g��-g���aS��YT�|M�# FI�J�#�0� H�����&y�`P[�ʪ�Փ�L��I8ن`G�c8��r��n� m<������c�~��WR���9�rα_��HYU8���H`����yD��P���|�օ��bY����(�<,!_,	ߊF>����h	�faIe+ R�B+\N�k��X��X=�.H/m*�O<�C���0v�ib�$yۭ�ci,��W�/~r�t;>�u���҈(�����ЫU����߉,�4��p\h���S��td��$�@ki�]����I���������X��H���J��\�R���𥑮c��6�G|�ݫ|�+����u��w"g��|awF-!�w8����^�.׻�杲������Yr��d�\���:���+4V%�=ӵ����_�BexD�2a��*�O]!ZJ��g�g�xk�`V�@)���Rѹ*'΂�/f��!��V)�bD��!F�|�r0�c�lx�?��T�;�(4?ydg�)�������J�I���X&:)��_�lەx��F_8�q���h���Qݽ��bi� ��h��(��-hl�*%�9�����F���]T�PbU�b&E� Ճ46tb��S�YH��@����8u��8B�N�-D"=-����(��a:un�`і���K3�W+�[f��l$�K��/�C�z4���D���e�z
�L�03�`��<�?)SY�e4�Pa͚G�1�2������u�4���L��W�Π'�`�=2��3I���s�&ǥxK������ϺJ�Ib�`��x�<e��ś����{hmI~�=��6�ZU�(������N�C����Q�=J^�	� �X��*�e�E����M� � �L��^�ߐ���Q��}3қ�~�t9;2Ke0/�����`�(5�����<X�AU=�M��VB��ІUfGw�z9q�ׂ� �,�4��R���s1{�nFh�W�߄;��l�	�����}h^�(��$�G@�m@'��)���ʌ;g4s��P��4���� ���v%o��C��"(�uD�-D�CJ��XB�rw�m��bN6"��ɔ�u��<����2Y��}�hP&C��%|�-`b鐚�ƫ���;����:�B��i�cR:8����|K~E	��B�w�B�٦�Ć��LW���"��@I:C�1�<h"�����S�v���HY�3�v�n�]�{�����l�)���RG�U{��P:9��ÑE��-'F!���#�����n��h/�����P6gQ�/�������H[�����D�fҾ\����0��yo�ZYyt�D�#iKr'��Q_Z���s�2���6��h��*xā8t{�a�C��2�[G���W��{=���X���x�YfOw-��m KXh��O�'�6d�ln�;��j��Vj[�M97������(=B\Ӓt��i�������F�s$n3�Թ�F��`;��j���B��2�
f���|��l{j.�m=�Zڣ�npD	��}^�V���e����_���ޖ�h�����7:� $�J�B��
Z|j���}��{�h6��x5����w�YLŕ~' q�9�Z��dC����)�$����B$����֍�C`��\�1�s��]���G}�C{����D�F���d-@�j�X忱���m��q�i0-d�n����1�-�z��5\�q�V�zsY���3jO��;*��4~��R��#21�G^1=���)��h���O��
���.��gƝJѓF���<��|BA��!��=�Ñ2�7�)}��O!>���+>�{պ`���7[��Q��]F� K5(y��/��Ӷ��T�1���r����bBC���Y&��ŷ"P�6ݛ}#H�_�v�a���g��;Y2�
1Jƹ��0�_x�������\���T��c݂�:��:�G�#����͜��ހ���.Н3�V�EL�ɢ�qt��,Z�ب�升v(8�%R�7�4Pƀ�Pt&F�{��'���Őm8�\������ڹ�s�"�٨
��ߑ���\�7.�c�!�%���h�v�:ܹٽ�����`�JNm��h�
�/�i@�uy���prm_F��k�C�5؞���'b>��Cf31"������#�s�O-�F6���1��\_�����en���\j8�[��=���i��hޙ9��X���:�0���qL�']�>�m��E��X�0w�n�.͡���t4+��\�S��| g>��I��Ƀ����)z ��=�����5��]�_DS�s:��ݬ�z �]��ŭ���CW~�u:�cŔ�8P��d�
S�_�n`"��ln�X���;�k�z4��쳣w�i>+�'�AP�t�_� J�Ɣ�S<��6�(F<O�*`����S*K!��m�|r=y̪a5�t��M�UC���$pmmŻz^l5���He<���;��W4
��1A�M1�����@�� �6�Z�G�����sc<N��6� ��N���ܶs��$Q*n���~����\�봶�z�\&/*cse���zxy>�����5^D3����q���J{,1�c�9�}V���RpO��Q}<����q� ����Y��g[�^c��)�!��D��\�0�q���+b�Y�<y\��/2�������d�����IOnݗ)���k?���u���>)+}|��V����H������[v��$��R����Un�� ��&��%
1�W�I�F�[W��`��_��F\���oJ�i�h�x_������ ��N�K�/���]U:e���de�@R|���F,�+��w� �{�'�����nſ�nk޷��rW����@�.����k���RV8�����G�L�ΐ�R��r�\H�o��f�H��ci���������@,�e��
���Hw�-7n�P��Gg�^w�s�~�'��fa�U����6��R��Y��i�$��{��4��s�^�M���|.ߝ<�_HF��$�K�z����C䐘�M9կ���Bw�_�XF*`-�����0Ls���1D#����U��׺4j��m��ҬKup���Z��| �bEo�#��1��2X�B�+��
3�]�?$���\�W�ly��z��c��u�oM��-Дiβ�D"����u�͹~�*ׅ' ��1Y/�J�M66y�Ɂ�A5Kdd����^�t@�]Jߤ�&�sd�kj��;����=�^�%ȣ2��'��j��q���r=�X�tz��ʖ�?%E
�P�L���VrZ�_&zme����dj%��k�O���n���( y��2�u��N��v�[�;Ą�����\������GY�!��z��U��p������/���u^��1���*þ5�hW�f"Ö�=��#��y��~�s�Ҭ}u�Ɩ��a�]�)R+��ng|d�_qH�T� (lց9��0�;�Z����s���>B	�
b��Y��WK��OR�\2#��;���X������c�	^6�ۛh��W3}HG���hV&Ѥ�ޭ_j~�"�:j�鏝�GG}��"�h��>8}u/O��A�v�D�|��H�� �ҕ�{+/�s�v� ���Ո�g��u�O���;Om������jբqe�scJ�z���e��sz�������i�os�Ƽp!��rR�h���u���&��*ߺ(���{���5l&���*�DX�%�䐶f�b�s-tgŘPK��>���v1I�x7'	\zv��߮��!�p�FU���M�km���V��Ędo'��PӍ��,(sD+9�\��U^(�N�)�#�y��PE�݂V�T@�H*�˃v "cg ��W3{� 
X��Y��U��(PYh9�E3X�l���7z�n�կAUY�7�PÌ���~pA{�t���+K�����?>�Tb0H�j����Q ��З��l	N�Bn�Җ�)��L��fǶ�-hPJ�X���F1��q�FE�!�l���}y��
��M۳s����tav+�J���t���6z�C)�-��[y;f��y,��|O]L��2F~�y:qh�6�7���,�o
K}��~H�%3����{�}�guw1+��!�|�ֺ�;��7��p�T1���q�~�(�k2$$f_�{�*����Ɯs:�"`��Տ~.d�4� �RLyO�y޽������G�-Ug�Ot��p���i|���x� &�����Mn��J�F$�r�����硖��*��1V�f�-7t��x^���kq�#��N.~�xo�N��J����/�j����(:��a��c3s5���v>FY��eƎ&t�1��b��f۴�M�P�뻍���0�U-������l?{��Ɨ����N2G��k���O�^ɿ�����JӽJHwO�Ԋؗ2I�>Yqj�� ��a�W������$h�H�	T0Fj������G��1���=(��;�NӴG�*�^R���'�Uu�߆0Gx�-zT�T:(�8��(�fh���}bO�nR��9DR�ho.��ڈǫ�ѩ�;=�|�����_��r�?ewJ3�C<�ߝxM�L�<@�l�p�9�7�Z�_����� +gD0���3����o�:��5��Rf��q���u]� ��/��b��z5��/Y���.l��FW�pIA抅ˡ��Z U�?�2Y�k���$�D$�܈&�b���Ej���a��&2H�~�Zx�K>�x�d5�(����K���̵8F�ᛦ ��z�md��7����,|SK�Z�/�9�/�������nFݠW~hA*�E�"~�
A�kG�����pHZ��5[�,�@#�ܖ�B��1Q2����&��-R�8�&�w�Կe���"ˑk��QF����Y5�wLͥ�|u_.'�̌��i0�4�b	@��ΐ��̜��HCr���N)��q�Ί�9�㷊���۟x�ufe'0}Q)9��m�|�7�D����*���2TƘ��T��|.�}5-H�YX�d����<O0�\"Lg�KدP�W�YHU��������]�h.�'�Z�u;��Wd/�~d��o�x�Z� �_��	��f�)����(�?mlMΤ����n��5V7*/�շ��ȍd� b�)���Z9��k���S��U��"�Ar=�r����g�U�0�)oY����Y�:'I=�V67�]�Z
���"�r�ܫ���e�-��Z++���R��zz(�ɠ2��E�q��w���B-4���Bf������*Gs��KDZ�"�rMfo�n)�}�o��<;��V��9�]02U�$��k�������Y��"��㜠dh��A����_���W�����t�@�Jf��K�l�r㜇�$��-f����%=����]��n2;Ϛ<�x����U�C��Y�42�w�+(n��O�G5&_�|��4���e�Uuـ�v���|)��Q2z�_���Abw�Xhꋓ�I$	|k�[�|q��o6�oz �;O�� �^�����~�7� W��.��hC8����*I��s�v��£����5q4��i��_�|ez����֞_M���-%������8.V�Ԋ+�߇��88��Av{wjk*�ϴsѡ�-�޷E���o�-s���Ϧ�� W�����΀�\����]��m(^�${��SR�TѴR)��V�4���P�,@B���Ce���B�G�a��\gq�^�!.y_|#�'�jd�x�Y-b2���(`?w�$�h��<U�t��D��E���߉ʇ����<���h?�o�6=�n2Y0�=��Z��5��Ç���9��4�o]n�*v8��UQ=q�%�uy sM�zL����֌�3U�9 ��u����Z|���<�-K����@�T[R��gM�1���|4��W��wb��XVsuP�n�t�2nc��uҦ���X���Ra��d����#� �8�r$��_|v�%�����8}�,���)K�V:�'"�+����o� �s����ة/�bL�v!'!d,���R~B2���Z�����3Z9�9�6����;h���["2�60����i��6��mR�����HV(�Ԛ��F��q��\b��`>�f]�k��1���U��D�_���S-CG��D v���5�c��ן�U:���P�ԃ �B�↲*$��^��M�fs~!L� +����Ⱦ�s磃���	ׯ�o��~�|;ꌙw������������BJ"|���Pr�N�&?�	��s��������[fAN�߉��ǅ ��~e��.������>2�~2𵞇S�HQ�
�ߑ�P�>>�7��0�4>���l�x�xya���HWQX�o�1
\���!�^��'�E'?��4�g�芏��
�L�7���dB����N�u�9܋�h\�gk�}�u/w$�[b	�����q,'%��^P�5�ȢOP�<a��F%��[
hj���"���ox�l���+�E���6ak~��t~�h��M�����i�I�gm�:1��eչFs�O{g�ë2 9�[���4�y�|���5�w���q��6��\��{�	O���K��LL�(��qJ�ɥ��~v:�驽!���J�L˼�se2����b�����,�|� �P�f��M9g{�ň8k��򡚪��u��q� �