XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$�}�5�֍. ٞL�H��H��P��(6"[�j۩���T� ��0OK�,�h\E�mh�"a�g�i��6:6:4�����+ى�6fP��W�f�-<�C6�����l��%������m1�_��	쇅��[T#@ʃ����!F���@�-v7���ѿ,8pZ��i�H@��C��N�̾H��ⷓ,�Ȇ�h}2~�<l>�� �X,B������E�h�)�u�$`9�y1ŀ�J��  �VIW��1�5PHP����'ή:A�����2O�wL���W'�)��o���.���l����5Ĵ)����8�}Y�����y"�����i���J+p|27�~I��Yz��S��Y������V�-�b��$4�dU��P_�&�a؛w�3�$N������<�����a�R��ac�w&'�ݍ�
F>��#��F35;(5���i#
d��'�*٪"���a�X�,��ׅ<�j�5q�8	����-��N��#��yG��4��*�i��̔�D���5�� 6�E�%��fZX�"͎���d�=u99{ gI�1�h���f�և�[�oW�����Kt7�Ç�6�^�O��Ӕ��K��pt�{�ۈ
�Ve�ޮZ��i��S�Ҳ��\|��] ��p�q3��|����Ʀ\&�(,x�E.���{5��ݵ�?��	3���#g�S�˽�J$ͣ�`�g�Ko3�R@+ѹY}��f\N	��X�.9\s�+��x�]��*XlxVHYEB     400     190��Z����Y&�*J�>��i���O��J���0�CС'�1FH��ܰ�e�n�,�Â�<�fM �/���QV��:��� �����o�Yľe������&�__�+LL���x�゚�ɤbu��)*%M-2,�� -�	.��q)b+1-�M��sqL���;�c����
Bw�%�����<��<Wu��� �#t~vFu�~%Z��74Iy��/g&�.��Z:�`����Hњ�Z��NҼܼ��]�}��E|�e~Y�r2+���8-�F�|\w|8URedn[�s����.��U0JD�tF�&s��	�)�#M)�}��0<+�z��.:?�tL�l�uHw]��l�苭��Dғ�*҆,��k��3V��?�!eZ����V�q��A�᳍XlxVHYEB     400     180F�2˝ߥ8m�*tͭO5qb�V�m��a!%M.>�{��"<�_�]ޣ��zy!��`)��1�̵���R���jt���������h}��He)��W92�3�~�*Fz̿z�h�J���D�xT;�n�
W�7G蕅x_�9�X H�$$��D�*����Ȯ|4"2T���"� `�e�Ԃ����H>���ЂF#��ebe��D�I�۱зn�/�ej�=�:�,���ѐvg�$��bm/$�w'R	��p����S����H����f}@.*��*BK�ǀH:�ؐ����%���js�b,�z�&������L�(��H�n��2�����:��33�0 -q`�-����I?�A����g#t�	r�x�H,:�G�0XlxVHYEB     400      b0R="+���#��[�c��\3x�o���k4��<QN����I�
���x\��R=錠�'�Q�T���������yǉAG�h��L�W}
��r:�	Q� �����4�D���H��NSܐ�Z�~,���k��l;�V�)y2gW��5�bwF��9�{J?-����;m`a������9���n�XlxVHYEB     400     170s�I��� ��~ P(���p@�b�C�q8��+b�q)�s{FF/��)����� 0����v��[d@2��8��آ`d�i	}F��X���:�`�_BN`7=�z�PܞZ�b*  ~���i��._F���<?�6�am�� ׈�:��Ø��I�{�Q�˿��(��6a�$׆ܪ��ҴZ&i8@�7K˄�R�1>�}Gov$��͋�2��&��������J�P��|PA4��W��]�ٰ!=�_py-��[]����*��]�x�'�uQV>��T�R��=��l�s��&/B� �i[`�4��ѩ��/�j�-�h��Ĵ�u�/���Ό�$�WV�#���ԇ�v1f!Rn��pl��]33XlxVHYEB     400      90+�,籧Z��:^tēA��W[d�:`��ö?�Wq[��4�.ɱ)qJ+����YS�m�;ͨЇLôi/G*�$`��	=�9 /�81<�U��沷��_�c�������Z�{�|��be���	a�P˒�{E��D�hXlxVHYEB     400      90�Lr�OP�]7�jʌ&|�����z�1�L�߅.�L�#�-��#$�w�l��C'靀���`Bv�b��;�uh�-�����Ȭ��Z8�FA�'�����Gd�+�Pb��&3|+�����&Ԏ�
�Ȝ�5e�˿tCC��vXlxVHYEB     400      90�P��
��헝�7�m�Fh�|�;����H�Xܣ1��Jʱ��� A��iI-` �0�g�\�8�w�!ҫ��R^�c���	�r��ꨐ,u���7�(l��ʰ��MHD
�(և��A츁
�l7~�������XlxVHYEB     11d      50мy|�mar� �f���[օ׸�0��BϨ�������%_y�z0��Z��!٤��8\ͦ�o^�q�Jx ݈,