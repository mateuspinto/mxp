`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
3CzOE/1m/gqj3r93kk3YOIAwqx3lF34HTdcmMP6l3a6evl6hYSR+nMSZBE32EVci2Gxh5DXg6Egk
R3RfNO/MB/rpBTNhQjbDWdcxpTM+LWBhK9OJ9Dfh7WetqeeQHi4NQYYR5aNkYXlmKpszBWapguJK
Yvvbvf3XmX/y0HMzFteQAPFF3nxnjMxImEQ0zYivs3d8h6pHMwuwbZejwVZcBAXL/eAR0QmzkJj3
cvejgdOsHhDn5j2BKI6aVkObQ78wy+BuUbB2iZCl0E3KeADXlmJT6CIUd61YWiwjvWjBdwIZlglg
eSH4Wrkqc88kYJPJNIg51S2OkCSjyyjrjC20GFyNb/vjNls7KE87VqUpcSzWoZ8YCXkQnQuro4RW
DIxXkx4By3IgmiY2Tr2G98bd2fPsJwqe6l8UXE/au57lygaOWbug1VJYkVkomBCO5gXvkpjvHHY6
eQEQ4AIF5gtuhfs+4yReHE2VCf20RA+UKQ6p8f3q3/YXF84htC5Flc59SQkt7mOe49/2pzfUr8Zf
GPnjFMdG69f6L7zT3+8Z/7MgqVvn3P18eXqjDJc4pWsXMosJ6HLMJwDfC9HCe6GYAWYGat09l9NA
LDx5Emlh8K9TYX0loUxE+LihxGMtMHZNwH/RVb0Bob0o1rA109/l6qqM+aJCCultjPjHL5xF294s
Axf8TuLqqylrH1cRZUO8+89XFEjOHjpu6UcfdlWzEsmAZvI9cHbtAenmj3+eFNe8arX+cONwHoWK
MgX/MTJ9J0OySziHqDdHASVEQeyT60+1co8oajQnSpZcWu557nFD7FivF2Cq8Vf1sMfKzK/7CcY9
u1ggq6z+6CWu88DheDJf/oPXVxjNVyfRIyFciXi+prTzsssv7yPgJzkTqmwdXe/FztuZy2zi2mDd
OQ1o9BEIAFB0HlrOcW3rmhzsTiwt/6R7PxDrykAxoc5bzw5BkGHgnuyJtU4SKKLr6bolhrS+E63L
ZrwPcJnADQv9R9wverATcZMo6gBHEj252wABI2lNnTp6ZVcfHK1a+4b4ikOw9ZCMy7KrVR4iwqIM
tIVvZLrLCiQpCvIJVA0GjLVtMHlTr6Pqk+NwkJ6UCNvOrhqvo4miSF/YGjwKmsF5ix4SnfjTJJds
8txFmo9EMdN1904VOQYm296cuTadKKreKwr4UNFNt0mM20BZOabqcXRSdL4rZbCP5dk6MrIyT1ZW
SgDBqXl9sSzn6aTAqN4JwX75Lu4LO2n+aZ9lQj0NIM2d1JahOoMidTpEAIDqdsV+aQN/uWgNIIus
Ui4KiMFJpkki3l/vi9l1fJcVw6zqiocVwj9Ilp3Iv0pJ3hINYuyJY46HoeitBuXQZEST2YBR2hH/
UfvzM/ymOIYES1KFhTHjReJrpPGd27njsuwPce6WuForM/67unHIncLsGZG1lvtzuZYmTQwfMdcU
qQBh6Zmsm9iQmSDwSNuIdhJh1Aea5WbYDeiWM0eJc8EJNBkNyAToEITD4kGNAP8BtVY1a4qffkGK
9amWhlKaAC4PlzOLcLlbxYI/n/IlJoKzLUHX14WOCJDkNgngh/w0ak4TqzfzgDWb8IHsaJN2R4bj
SB+n1TqT/sIXT96Kk4YQ1o97ZNJHrXV2BtL3/PJJIGdAhxUBovRgstgo1NDv8gcEGKuZ+zHLrIe5
UMECKE0EpNbfNGoJiqSK6UnsbvcV1bIF50bpIPKtXBHkw+FVYBtXAxhQwNrO91wNVZgIkvn9NzOH
ml7hv8K6r0Z4wYj+F1IIRsK+j8mRPat8TVmjhbprvbd0SxBF1Xb/9z58S4qOb7/k8fbRBeKu0/+t
rdCr3Dntak26S3bjeBXqKtC00Ow2zswfoUqUXVo0Pa4YybsXcvIeLOsvPX41hNjNLyewOxaM2+W9
7YB8W3mj9yyaJulaheYWDPBSKB4Gq0fCeIvCNp8OVauwUtYKpTnustPD5ImajhJrc88s5s6rg9f7
DyYm7eMI9IfG3fk1kI4D0LutQ16Xm3sZLC3S1bi3lnjchxtRoMpHRavjQMnLkWun7S+I6GTu0LYy
gmbV9+aqa3QCFqdXkWll4DSr3hXN026HjFGHtYxXPGn+JygY6WmHiaibRUSLBBdaFh/HRaLX2uw9
vVD8mXUN70i3dlJkxwo5yDvqI7ULFNn9TzjmnFdrqpVLucKlyptuxowSQEI6kIqa8OF5wtZcRwM+
FqZ/OJqVrK9wkLTA9EHhxpkQdIMjO+fxdH1Bhbr/gfYgcshtniqP8SybREBs4675mj8lT9kMSEU/
IDEpkMBqqeHIbrB2t13bFIr/fXvxxM1tb8/5Jp6Pu2guQJjBStqFnERBaamhYb1dY8c9tHs87c4v
VsmbawfZKVmVqh3HDV6thE8KPq/WR4jHgRZhb5fmr0PlZB0Ro1b0YQAPaKATVZ+U0sKHGszyP7j2
YkLMX2eHEete/N1bwAu/t2CTtOEB3AA8+YWiYoF4OIjaoJXF0amHPR8A0ei6M1JntUHPD0YItYxx
vAhXiHAMjFkgMshSf+avx2Zck/z6t+nv0Wc7yC6jJOp592kbpsmCF6kGIobVcTrw7HgF9Vj8pvA1
0tZaT8tljbcTsHz8WO5d0JJmxRxNYruANMxWgzZCxQPSpr3Vu9GJ+1F1ylEkxfXCdccgT98yTHn0
iIh94XcIPM5DkjmswpQoHAdRu0/0GNdRjIjQRIUFUqCdVkfBOJoSyoTPh+I7nYpmPIXQWFxvG1zY
DjmvvPlm/WJGOdZ3zYeuTeXNYGPN9BZYVS0JcuZgf6jKY2lZyftELw8eLRGJ716fSpBgOHsPVSji
lWzTXqAPyM2s4Ufv267kYHXpOZkWVNuM2eR9rQla8qTPTAwk6zTZnTbDJa8ayNJvy39oDqldCNPs
r9XDQa+sEoK5TuyUSVovl2OSfb3m0TsvaZnTRJ3JZW/gklaNyEMjCkpGGvw+NXv5YhshJ8frsx9S
ju7sWECXUNJkPFx6TYTael+2F9RYkoxM8JjGnqHseVzY0mfz+L3CwOSTF+mxHjxZFb3yuw/oKaiE
eEZLNYpTkFL6pzGGTeJzCSm3wWJrcY4fk5yQ2mGPAQCWLRYPOQpjsD7y4aA2bvfRlH52BIYoiIe5
cCO/RIeIuNkZZjyoUH5eyupPwwFj/8NkzmpkkGyE5pMh8GxhhB+thF0W7t+hIkhnHMQnhNcUkLvz
pf59oA3vuzQic6Xb8EKlJCogYvr+md9smRpbiZ+YVmWjadmw/4qGKSpH3DsCcQlhFofo1IMuPXLh
W6CWQO6iNVin8jv0nLb3MZkC6OZzgCZasOYAtwV1lbd8Hbpqx5ZoplQN+VQ5WVuCxghhbgkdrSIM
n6v0ungW0XhVqecxCtvneerhxYHn1R42fhZUzKwJ2gpcTcTdkqSYzPfjZAFaFQKuePTHfPRkWrUV
PvTUZqXmJPe4HwEJ/YUEW4ZvDmoeE3BRy7ebFSnjxhUnS1gxceimmR1h8gQ6mN3FY5ctsPbPm1ur
VyztC6JJ7A8QE6tOXlDF+O0Mm8CQaK4CRBYWB8Q/6JrN6exa5NWxnzGcO+TkGL9mWqmVq6SwCb8i
HrZNjKbMYvuZhtsxQttOFWQuufjWZMyRyWfdyC52+Z2jpb5QHDjxj54w8flbV+O2iE9ImD5EFEoU
44Oa8mcE0xg3fNQ+StREeeHfzVXU1cWAJiPNB5Vj8frLWGBS0WgqpG+QYnzpz+yGwRSGcWoayYpA
dXmi6YJ5Dl0UeMI1nm6XU4jZJ+/VvHQY0pH2uqA4efgykYiMiEJKiM9CX9RyB65k3wW6hcOboX8y
L+KqcchwdgnhM7GeT/oSZHV3wnfNZvab0BUBSeVTNnIWQ4nYaeiQk4kAwhxZo+VU8OGDKu73aaAq
aCmY7Xo7CgGBCVPWFTyXXw4YDXlQUrxwbMkV1X1v4ONfpsRmyIYsxYZfcsZN75cblczJVjo5+g4/
3sQFz2KoMPO01eyNYEo1OtSTMmBDIdzjxxXOm7T4Ci6dsnsegHzzUajrWJWpC77AhSU4+Q8No8Ci
0i2MWPmZTvKKVx023xI+3HAv2wjltKM8JhXz4Dapr3goITy7DwOgwbtFNnwhnEu9aWGM2fGh//qv
EPqD23ElYsKuOWX2FhjbCFnfVnT1FsgX/fXvoYrbfwHoh24QZhjw2fNQlJkm2mceuOJK7Ac495bA
nVruM/DZ4B3qEJEFSnpbKGeV40JsNqaJuQs0V0RSQKSvv521Dz/DHh+ZnJB7MXDL7MsJvZF2jfCG
M9M66olkQweQoku0blOCjiEE4tyeFj5L1igmksSdV9tvLe/nFdey0SxzKgLKBglAvooWCb1Uywtl
Oj8HKNS4zbYc7hv/TpKnm0q+WSPjPp0UReByKPhynTcyRbGa59a2HkD932qb9Kuko32ScslvLBGF
y3yebtPvAQU0hhaUwqj7wFbDNhgCQGUp7a98IjiPbEvom+cwkwsjga2I1Thn9xxTW0HAXdpKWmxs
mjeaPWGZwBnK81eewYKgdk8tXTrsnDRMR7MRaAj7L0gCTWTY22MteX4ZMjfc2EJvmU4RsDBKR8su
upjzNcSLlIMiAvOw2xWqqwy+KBH/UrfWy9A2vMnJJhxyFRvZOoTk36DlqV7Qm3pkbc4jGyMtL3PV
RgSBN2F/sMeqjiMshQSnkYnCVp3U88Driu6ENa+ExhFGjW5TzVmIg76TdvgtpCG9bSMKbQtHqnOr
n0Nb1dzRQtsew5ax5KvmDN7sAg2BxjwHZgyUL2dhZLIABnKvJ+vKFoHTb9k8BCzVYyGph1vUSMfv
sTgZcDX4Upz38pA16loAKvpCA7fzyWSSY4Orj+7du/rhPUbGnzx5HJUIIoDt/FAS+/oayXTFLnnc
PEbhby3cwWC6JUESCuBhlasJu5KR3kr5LO4MA7pjXK4j3+aoTdCyalU4SbMYuuHx5MZCSt44SBjn
PMAHz6BuZFm3d37ZdcCvijqf9es+thQdd3kZLDXNql12iQNZD40GZ9eTi3okzaF3YLO82JStsv/A
y0eQ5oNC2QfM0YgW9o3OkLO64AMczXcHYnrOAlQsNT1y3Qcf3vOyYFGOgpKaMWQ0RbxmmwkScAUz
q45XYuPDWtQ5D3HV+izQLI6QJHPjBdmMsoM5otMgne7HNLEELuoA8NaGrcYz5Diz4c9iPp7HD9eZ
rqULeDN8DUswc1Jn0rFWg0sj9Ed6raiAZtsEQOarrH/mTuwbjjTV9MiaeBjn8Micr65cfnITxuf9
p5aDHspd2VopNCoN9Xc7er1B2Gfcl5dakexBrvnB768eFeISNC8fNzfXDVTZNd9eGo7m6NFd0FQf
ZOKxOF3tqn4TCsvXewfzqXHAcghK7Mx4VmDTcY87UTsFHLyVyXlz74KPZn+f8lnzAtbj86MQB13t
tsOayguGGGhHr+jvmWfcBqdrvjDWyFPN0k0EffbccqEvTN/heira6LscDvmiKAK2edcJ0gFHZLxl
fFNR8oepsWYPUxW9i5wU1AdXhEKUa731EqiGtNvxxcls5AD5vldt4dHkMRZkvm+/Fdouel6fJ3Ad
tE/ZTu4pU73bCysrK8Vcg0Vprme0a/PToefcWqif1RM1aqkWliUXGdiLF2j8RPqee0TGDM1rVDnR
pU1zRVlMH/+LejWMwXtQTvIFP/P9kxb4l4V2CW8V55xi9K8rh3kvD1Gaqv903tanbA4SwUNn7KXP
kXvbCKm/PEX13s8PTRmd/Fa37dl0P/R7o70B5b9BLXGY4OObynoLf2YWWk/QOR2l0XL/3p4zOaLp
WlyodwINbsHKyMX/Z7L3MwN7CUIZLoHPIhsV5bpwIRV8A40s7z8seGXaQorBaUyhtv0WLdk5iS68
AqBD7NIIdI12Pf6hVKB51LEDfDuIdMOZJ6p+paqeQezvyW/mU68QISxq+QysBi5nm4IrPkBfybu1
nRgka58fj4EI6zd6yM4+MSKq6D10DW2ZAC0PexJhV/qhu3qxwlLQTVzky2DRIHYNZqJa+PB3s0sO
HZtzf1buxgqcYFJFx71AHCq84FDtMOUgDk6/A4Q7K1L+W86lnphhhJb4q4X7oYWItJe/c+yMX6Vy
EE0oudvCpa/hxGYmomXqqq0ZBPm6NHRwvT4AgDp2B+UxeVA2pkSkUyc914Qs0kN7gTrS5RvD/Kll
3TJ7FDPt1kbjNq6beHkioCz8dVbbCEjyHpg/2RLCmdB/A9+Ebi7ktEq+S6soq1lWWMRUHypRfrGv
HClT+adHAXMbuSaIdU1E8qq6n/m9StV+daGDti/D7h0kMht5QhwlzIq6yDurZlywLU9iSTBiO+Xj
mvts12faR2V/41kHVOLA3NnhtMQds0UKSRIyOoztxDYo0UQvigAPCA9/0H0iZY+FcxmmoHtMsLxm
BozOgT9ZbyE28x+KZdYDYMK9Ehn7iy2H8On48X0LcBj7wsDn0eiKbKE41Yc1COA9qenpRxMj11cy
g63ck78kDP+W6dikQBlgnB7ft2hlIsKw/hHaOvHRXGW/Xp0AlhHPyTaiNLT5VJW8q5MKrZ2/wqMd
AjE12vlGEP4XuBicYUy2DHeFC0lHP3ljpTCzc3XHGVM/qXM1fDyeKBvOji5r8Y1IY/Gk+Mg34K/p
IiHh4EE7nD9AHJ661/5QH7yWO19Y1zxtZ56RLyvRtngn9JRko5I+MI4GT+yDJIZofQ9XyNPYZNk1
z6jWXnDmOlO3PMjRM2FhVMrcVMhmR1sxqx2jFSQHu8Go+grbuxAzZkeQdwxj1BXDmT4dybAw4pn8
dM0mZNEnQqK2W0gkblOaUghJggBXCL4fvKWVPJliePulQQg9vR2yj4MldYkWpQnlRe5+xNzdYbLv
H+CFEUZTVtCmvV8cgn1zIcjnSdPHqON0Yr8sVPB7f5C+Hxvw7kfDKlsQSN41/Vgye+3FAjdEwC3B
UYpifLc3WdLk1TxoBzpOadgV1zogN+81e11VkEKp8MG7K8+RBUwXdUnz8k1Jv7Yvaq87oLW7yJxl
UHQlKvPuBlhEJQCQm7uZPFfBfElD3bGMdayfRxKlPvakvkLJ8hXETeaCatqvI0d2geILJgN1sI+v
KNdJra4xnLiDLx0sQPuJxgLtKCdUEwM6qx725vzRS1kLhDoMRDZj7n9LCuSf1z1MSPsY/sk0D/Mb
NGxaOndebqlk/EwFyDomoxdgbvRPEdbJeasaWFBkt4pFJ5+pP9PTVHtHjmQkeMszkF27Jqdzy+9U
ZHc9MOg6PDj8KCA9AHQvvWDqYXJoJeVQY9S6jjKUJtdq12XEfLywTQrQdJiJWfWt2n/HotAYGeg0
E9bXa4W6OpwX4wU616VA+dXV27JxKzk4M9Yds7YctFb1dGbBt9VFuEzHuz5LYWlHocdrfHe/YpMR
r1PdnSIF1nO6xOV7W0taCGsZfU199PO2K5jwh58z8EcxZtp+UGdnPFTc8zZjGvz9Z6vWzSTaZvyi
FBO4bZyDwbDHw5JV5m2ZZRnjhjCr+r1c8paJmw4tFgAcznEeo+zVatq3eqAcMCpOy/yYUfGWV7Mw
nYr2J0rQgDUThIjJ/PNznXEFXw4zoOo6H9lKrG7s/IKc34nG9wdu9J3UZZKQbM12ai5J7uLqDhtQ
znKLPpSgtBWALRZsggqPf/b+zbnj/diSEqXuox3F1dL232UmGWEDkkU6vqH1pqGjKKToAWU/bNSn
KT2xrrx/za2yZ5P1Om6sl6C40ug5Sx62YUINrBMFgUTM2kk2gfDH//YXR5r7silW2qxip+Qt4SQM
QAp7GlQfXfirEHrB0Zy93CzDG44iyJDXCDR9emWlK3oEMqBSn1RCCiPgjRAjMbSPBT8E5ZURlCnd
YhHVNVZs20jEG7eSD3l37naK/IAR7v6XH8ZAmuAlm2bf63ph1zareV0eNhfAVXBTazwhARiyXe5m
G6BYBoVvNiKlrY4BDxNuJNlT+T0PhMJKfQlqw9UwK+HG6IAWjuc8J/Ild1aX+ekI8gqkrnTEziMm
3tuLT7ukLaMq7P5rcbj4jm79MTC5Vj0pb2h6kShFdFWp1Nasro/qKE9w1DOjBFEmK31LGRdKR7sJ
wWgIjMAquwdCyQxxfi1kYwmYkdBJmcpCrR9boAvd+mLx0Gbw9qDBBOYu2jBjpqDjfWh/4SpDFvfz
wqroe8vjFp8g7PTB8O3TuKa6qCbeurii0oWj7mQhW/ROzK7Q/tySsEgtkgm9F2K46OkFE22rqmfk
BodI+YbRJgu1A1Rz5VEgk/aFuV91s5gBSj5LHuMeDe59NErRgX/cSvAK4ffmVMP5V/Q7ybtc5toE
Xp3+e3nhoEgh+oj+8Ja0vNNZJ9u2Nyhg88Hg+2sWjyAVWdQTT4dPclVjewlWAqVu15d5y8pQ4eu+
ES+FTc3ixTDsAGsQMNBSn1y25VSwknmVrMyX1y7s5ou/80ytQnkO/5euUY5pAP7w9U0vmizkeQ8G
ZGjLp8yqm42vrXOPTkm/2JVVBlQbPprvjEXdhdIsG53HiOK88ByB96JhoeRRBPG4q4QQ0Y7sMEf7
3leCML81aLYN8hnLAv+erMpIhh0Ys490yrXEMIhMDN5bunqfeZwvhaa1l/1py5MqmIMXw0nJWp9e
iYgUMFobnqAph13XMcqDJQrPCSc/42FQUS2DC3bYDvMTi9BTlnJUA+/Y08nY/ZlKQ8ZeRKhe568n
Q09wCzr//36ka+j0m2FwVMVHGlgW8QdZ2RkiJH3yT39TSZbd9KyzfJ0b4so4jrp8hF/dUE9XrOBR
hqWvUd1xe3h7oHgSjwH+QnVPx9ubVqIcIrbuXp1AoKPZCP5b6pdOCyFJXmCzCErrlO2NRKR/TnK7
cvrSEAHI4gkUySruIFGHzIOrkE7/Ea1j9ce+BDVhzLrnv/tzyl4aGA8tArLuJ25FotH7jaCzqqLI
nR1EWCNdwDxCCziDvktyBm3LD0CsPveXfAeb4ery6+UU6QPFUNEUgMGuTrwtA/Wput94bQkx+Z4K
BjTaOuXAp6Znc541/iBQ3uLT7V0XxIxQ1zQGslnsYi8SUyoJXWAl8IzewI7fghwHUVavVRE8+WgA
YWwRGqgoaUAXTvYkauMvqCVEc0KdIUyKE0DaoHhHdQcTA+ytNcPffWo0yP+MOLZS8ShVnc85bRWG
dz9j5J5ZJ/5LPbboEG5OflPcaw/t2PLc8YN46ZH0KV9MNohdxGyq2pQW4X5nyNrf6+S6vvIm1KxZ
kNDz2jaTUOwltSc8iTiKyfflQzLEXD0VgiyCdREP9tsP2aXN/5FHUCbVUTqDvFuaB40VM5202SNu
VWo/VXfSKu/WCbKtgODPmPjjDlA1FiIG7x4YLAndnVj8aOO5eG+BDy5TrliKIVdgs369SjpnI53H
zzpUubB1hdXFGkNMgA2B8we3qfmBiuQR4Hi5LKYpCrJJy9HxFRkRiJKDVPdswMnE7iH5twVds6Lg
+B86aWJPfue5GdV2omK8qHT0houqSYRnLlgmgHM4mJxkZ9ojBEisPZKnVvI8cR7H5HAkc31X6ayH
WFdzdaMKO2HEP2pkqcXyTYk3GJWMMI6nxXQRwxn2m4fYgPfrVPrjPYpFMwwDxSG1JBFeYjBNHafy
RErOkJRx5RML27Wlk/O0HiCQbtSz+7CO5c1FZrCUpC984TlV6NVzLRh0zOpIFJ4Hb06KTXBH/zvq
fqxqqn4xTkUuovoRh0qQRMwIcgYAfet1gkR+MZAlZZtVVA85QB2SELNPDhFO7lOdTqAJCpOp/1no
zcCnY6MaAqFom0eOL8ymy6a2e8CdTexd7F2s0YBOvIXRHal5P+b+De2QAWf/rhxdEnEii5y5Bb6o
iobCmE/mTcOueRxksRVCvAPdxlvPzQXiFJl8f60yVurYVZIx4B6BxVWCbSjno+AP/gyGc32yomTR
UadOF9Jjvzt35NERvUd/ounSSrlSMltnqoEmEt4z+hUk2iT3/5RWxGDSqJRfUY47JERj/ndGKT4f
2/MvJXk=
`protect end_protected
