`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50912)
`protect data_block
D/65d2M4XSKZY0fYfX1QWtVYpbOeJLQOFIgCnCliWwkAIoWaviPi9uogyErmwAznMR6fBcaEn/HI
K1UdO2wXOuCFiYC/V3HpdIFamEPR4AhH3uIQs/c8b8lmIuW8Zfh1smSgfo19QmQdr+YkQeOcdLfO
pjDnQVQK5n6KKyIE8H6tniYZOqDB33XqEf47lUZpn6F1QSV+mOrN30HKGePcWhAB7/TGnphSH99P
4C/K3EW7Nc+lGxg95YnF7wdQ2NvFqsQXjCjsmZ40X77zi/wlQ7sf5tRgKrqdJETDPjrWID76u9QW
E20PDw/9Keg18sJdXZwCWtFoPysO2z1Jykkozt0uMMI43AyfoGhTnEmYiAsno+gcXf+xYRSGQeiV
4FXMswS80gmfYb+eL2xQHziGyuEvGgn3CnFfFihAsDllNsMeRpdXnrNhVidJqm1CRwL/fDhRvbVr
P/UbvAzh1wJexXj3GbOtFpXdGKan4IzLTB3+DST8/JfX/8had2VlC8jYkDW26EDYG6jpGYO3XOAR
HSkBo2hp8sWe//ouC0Qw1wQ7mR70AHfphq9x8aRPlrHk/3vqo1S0fY7I1iEoc7ZGLIvAMsDNGMz0
q9jgYVjfUZtqObJwMscRp3yKRnKGy5t2J//M7y0slVbwpjVZfwaFQn8MjDSFP89kEH7blRKo8yzf
rrox714Bk/VPSlsEN/BZFCrphaQ0GhJHdQj1MPphK9BgcI8m7JpDPK2PXuShUD5AC79+1WhoELbb
xB1oXO45+6/81tZ881GQjgfMW97/tsWLH17EYky9fPXtf6DhPaP0tnvMobdC6o9SKuLMUjVi/Uu6
khnpu+GfkfAyP6//Wk84re2B7QbJB007ElPqOWOwFVpdGTCkLL052kQCaRCp161ndzglEP6v6Utg
B+giU9SsF4cLHCGYf4d5HIAgWY6MK7OQU5P65rQChTLTj5UFaa/nyD/Uqc9GNFJzP4svFl1WRhce
40Ng/NsLTPdLXu2LT4DfqApBUK195CsdegwAHEf5u+HrvMNFRBg75Z6Lam3SJ9ePVi02lwkp0zsW
8fUxMuHmOYm5Z1oAhZ4Xvv09ETDW/HoqluMWwDbwOAaDkRxX4dizD+KeB03iuz0c/W8MKPajBue1
EHh+YQKhw8sdTJiVQgjNLKLJv3OeoeKAX6K8FzZAeUwCO2RoXu3GFdObqMDCFge2p35yCq/6ntB3
h3vFwoe07gUe45/w1vBFKw+BRzsv+RKeUhr0KJgbLwDSkkfwJC0NhvPf5j+ii0qy/2Cg8t3GEPas
otUMMVVQo4Z/YB1MuB6dR256oG47pSpD9QT6fWrru8SDl/2CtBJGpboqEBZEHR+Aa+8klStlJrGa
+GAgQVzeTk5RVTL3ojVxKdTT5THpmWo3VrmW+SdQ79bCXPrS8zlkuAQJkf+dDmqHy/+s/MOoEEcx
Deif6AZfhxCOwiRY+EVr8MFtio/ShY1Yej/Ivz5fi5NbWpQxKNhszE0KsL0Da7PjUXv38zua0Dwt
TCqwbJI8Y0fwRG5afx93zcRYdFTQC9UmWtDfyRPhZ0PGEjN6IPBWPJhi0R7FZ2r/tis3/4xzov5U
c570Qcjzoc5H/PVYmyrsIZkK0fa9xuGRvLYa0/B839c0/XPhxPPwobdbDB9ey2+ZpzoSX1UlHdT6
hNizrpHV0hZjoCvKi372XAZme+dKAUcv8fVDOUlNE6LaaTHcTNpvF/6slCJNYKsuvTB2NFzn1dmM
SQqhkEYRIikps3w0x8Irj+En7gaS3RTh7ygoRbiGrgo3X0MNnW4G9qmUxXOMH0nkuzFA2Uw/aqLz
xOIHTEWiSWcFwMxYWgycMp413hdn4TSBAhuJ2D6lpWBZqyHnS183uu/vto5B9pRW8kM/NBwDDF/G
A8QWHksnwxcG04Zz/mSMIXjqvovFebQ+lwulTXknNNGE2nsi0yheKDMWgj3O71phuX87QqyLYH42
HSUAfelJveRSFMnSpdlqrDIIS5qV+KqDNQU/+5ty1BL9hN3TAKaFTU1tOhQSA9H4kmpyinA41Yuj
NL7vCLWJFfuAfHaj+b7m1uN4ZMqRvfdZpJU7Umq9Q3GZ4knwUVDOYK/pCVCluVcEboZDIRxwvZmu
Wx4nbZhtH3OkaNsVZlFopd6ibjDvH/zENTMKq4NDcZeBc3cbuwzHTeBZ3pWKxvCuiq2tHJ1zDWD7
A4es2WU1lAJ/aALF84gtRnpF168+R3wTG1C1KqHJtj94TK95J6Rag0tMqocqb3atOfZW8g0i8v8y
Doe/gDUXYqHrceOqVaeONkkGlEmc+B4N7AUEBe8EoKKGPgnMF+QmmoLVPyTRSqu7L5OIKxfJEwOz
zmDb1adUA26ecVZ47OK7lynLmwc1o3blQVkXCkjowTC1v12s3nYqwi0R6EXRb19JDEhUHeoVwXPP
fZMdFleyJJXp/A5Ka4Tkia90W4cAsECIzl8vlgR+4JNk/dsrat2JAaTIPYXAF7I8yTCncYNxFj4S
bDlSxFY+tDENZSPELroKHj08gPRonMHAXS+M/OjWICLVZ8rMnN/IwDHpy1OdpgrkD77S9U16xuUp
u5ZZXisDpWlT3YMVP8MsmhEVA28zxMuzTYqPCX6u5IFX3CQRsZhcu09THuKmCQnqAvL5+6mk/JxC
Ffg7x0Sjy1lbvgU5AkxbrRlBEOw7wVIJOZmnYtJxlND6ijGFyoXcaCiWltuGu6k7bULGBYbHAVPI
C2lKl4s8XxbY8eGpR9IHviBSm20CXpidsMvwk98MnBF0sgJbavEka5SPWOhxkgxXxlwUUX34ehDT
d4+nqafpghMM+yvHnp90fO49aU9F0oIlePZ2l0+KwWg03h9Ab/rEgWrfQvgwIiFB/9EB/jJ4s/Xv
iLnD2FtgRxv1R6UCG7Z3KNcFPmk7xzr9FxhRy/29m3aPamGAZlRK+tWJtPIjKDDZX5e0PQ6bgyu7
EJ2dxpp9lAxWa3qqXu+KpvlsqVT/6YO/GLbHsoos4Fn6zVcnQSuqXVfndbzGSjGIMX5RmlMUpkp/
mtkDEFZilfQ++24vZ80Ci+WduqfmvpMditlTp6jKuJhd8ksu0rWiUVbx5m6F7g2hrg8bYy9eGgL3
JzqL2obZqpnWtKpD5T5TkNCrS4sZPDj9ANhDUnRl9+LFGmm+0c+wvlNabOFAm6PhV5aWdX5sjoih
Fi1IfxiJ0m17x5E0xNloCub/F2VgoicPFpR3SDTm+yJinAs1ifV5DCuElATxq1LviAQrtaSydAlt
r1ymejn+ijMmDaeLOzkcIAOCcxWDo5dXVe9GC32k0VEXn+D4cMUEHp1wsSfLzOXkdxSe/343Yb5z
2mLFTkoRmhtNO/sPvPCbFGWHQ+42TqAwGca3G6VoaiEwCJ9pPdVkMGwHn8vws30LlDsJVTPd4BPZ
dD4NxZVZb+tkx6kZ7QTXOkoc6jgCVpfS1h6fvsqq90eN86rxF149QkfxeEOkZ48hLTahF+tkkQJJ
kDS4PFVJDCVskpB9b/JCRkW22ghcZoGMRHONgI8KESsRpCYRsCFsr0xpxAM8QMX7NlT1IgEN9k5p
0+5XLw5Hlt1+WU7IWlgc8lp4pEGhOKeXDR8/kAiuXtpCo0AFxdhtMJdtfkbaAf5w6956UaSjOa9f
H8OGgsDDVWdrjEJjMUIjwPut3Hy7WhYAvX0tRPT++3422HrlpT/Jz3Uquy+9Cz2pqKnTvlo3rVsc
50Sh+JHGFDDDJGFSOguLJmVeZEo8k17Mm8x6W4H9oPRrpqYeAGaI/tHVH9FFocN+UMTKcYJtVnZ9
y1xbd5VVQxRWJ06f/fVO99pWB4trxSbbPXnQ/hNm6TGzeCsbarQriiWT54mrQ0Mrspkey37v/AFP
/s5zAR+SlpudTNEEAVFyCBPQsZfTuedd0k9GWsd4/IWUwQEogxexEv49S6vYvaXlqFA9KW3tNq4O
+SAzLx54iZTDit82n1N7makAqyRZsyXwldKzDAYqlZW/GNQAOefwufmEPceSbTAPjDYtucTits4K
kvJRr/ZjUnVlegc98fhNMx7naYBOrrY+JLL0gT1sfoXTkZtNvMS7k3nu6bH7nNN0ohGGg7/t2/Xo
dDhqedmbsqYKFcMssb4v5uywHYo7zONyN7XlwV7ZQ+C0gtuU6g3jZYkeNd3aEgLUOO6HIh/mRhNK
Me0QjvW/bqwmAtodEp2dWfzmkj1jj/F6CddxmCqCzFiNkztGC5NbSgUyviz1jtMv8kSVMAnq9/KU
/z4UN3zgW1V62oFUVxyp3I8fvsvLeH60Of2w4yxH/H2+fLEBkXoR49nWy1BqSMMHSuerAX6CWwHY
CvPJRkUjJ7wbuP5k+23XQ6YvdhggQSGbQg5conVec/+rmLGQKhqgpI7/RcLw2zY5h+ECz8sxvN0y
4PwUdSq5UZjokVqr97uJnlrZSEVXe5CDuOtk9FneBf0R+fF7f2cfuSY+rZWNm4+ihbbxwGj9iiGW
6RM320gFesdkZ/OMQgazzusj/rcJt5AM8QJx9X7ghkTNk2ph8LXQEpIXnorqw4pstA+aYD1zE6Ca
XGhnQNbtiNtbX8a+rYz1z+Q2Ju0CF9ILbvPYAEFM0ue+2YijdAD+aU7DmL3jPanP0BMTH0aauXYd
1Sggo+RUsa7rU2MwCjH5KqhD4jwqKHp182WSKyOTUZQhtVKdOoBKKz2el4QHcnYejIPtJoYhk+32
oJ90QAIU+gS6T6t+iNOpz0L4V56H05eVdgIrbl1Mc4Z9b5+8DoUI3kDAkSNwrcPnxWKBcrbp5T4K
ACYZAcrN3bsP5Asbl83GUdD4D+zYXDIiM1UGSTieoWbzouuosPluWqJclXUL5YtSVS6R/g8T4sZ5
3MmdxkDELmzodYiyREfyi2LI78gsNI9YGXlSiJU18QP9Q5ICJJ0PxzXAzAMAsieJl2K02jnHuH73
J5uCfPnVmWO7HBXXzcCWwKB3Uu7ToO4wtvpDrGhW0uRksj/XXXKenFDSgninTV2+fmR2RrSrxeP7
1/K7LWKAYxJXfNTeultnMaVdq+HKerPqxEAna3Wdp6FooNq8MWyvGkeHV+i31EZ6XuJcF2PB+FBT
uW8t62jT64OFp6Hvlg+N46LhQt3YUbGzaCafzY9iXgxAMLU7W2mSsUTyYwpOa3h5B3fX5atSGQln
0EDQHu2v4WfLPV6iv8LqOBtMbdw0LlpYUCZEJVhTZWmuhc0z1xydEd990snjX3P8uchsmN/PdFdU
3QAhbbX3fRDq9XUvTHhMhNLZX0uuZsAnLmkZAH8lJXAEANN3gUH6gTGu9KsbWEjnPr3srvKT6vOH
lLGuS7vKcghBan8DLf/P0Sgv1X1yo3/8s08gIKiGv4/+S9rGHtu1bOXPdE/c00GfjgU0tphn7FQ3
UUY+707OwPVKDqwzMhy7lv3o2naf6JiGYwdhzhuApCXSU5E1KCWOZtcH0rC7qJcIXbivRfjOa16h
lJ9Dh6+ULoxfCR8m/qIaaBJ+uZUqq+RhmXmvz9vZg4Cnd+b05fLJzi+lPWtL1HoLHf96ILMfYdQ6
EwmzzrhXrAfRIzVzaQHxwGlhE2DkK4ei1NPjvY51ipCrxXAerUHHSjYBgW6AIYWw0mVENPRoxHAu
hyvBcVw1g3iqVTVc55LQtBHybV+qFKfXqsgb8AVJLBA63tRPRz1lLNmOQW5Vg1oocRB4YR5QbyFm
f3wc4XzGZ5yR7sGoqtdyo2jvaxkeZJBD1XBbW7ud8coJoWVTSK7ampPacZ0hq8tbyZYY+8NI8XHm
8xlekIEJ4SHtwG3dulVndlRkF+isqcGO+cWLswL6x3nqXu+V4gtspV2XWAd5OsN/Yv58FMYjTfYT
U2O3i3Oe3G6Dpdct4PdRR+nREwK5asQgNzfEw8LYBE+e929g4RqlVz6hQdore7KPSPMOXrWdCUUF
JqO98hA2x4IMNI4jj6oGYJNsXdAVSfV6eZ79+MEBK1zNZVnKklC87FAGhdi5n3f38VwmrQO3Tx1d
gVpKpj4Z+B21fouWy8BZCjdz2DyfqwsQVMKVxsAzu6SRgBbPmuk/4RkxOa7PPaGhhB5qeE0LwScB
Ad0ABQSKQ8xuggzMld2MAsTFlIJpFcCU/9Wl5wEtCLe4L4ObA/kdBkluWHtmC5lGU28Prym0qEFF
HzEkRb1qTPU5ioKa1dMtH+drXuazucZrCSvBsBhHt9ajXddFThzsnDMkuk6slqfk/f3OmXj+6WmW
jIVGDOZIVwaJFxTFEDEOt2QHmAsWeRKR1pnzu/nOuRmLyiyRcgRq6W2oEQvCG5kUTawIFCyn1eWA
7t9VuOymDCSyIua59AR38bVdcsgFhsE2dYkUh9+SplsiVkKLX6pJ/yPh/bC8330+emaMpm9p6I6b
Er+H2Anj/labvtboaArKNllV3AYcf/AMilEKiRmS4f7CiK6nopRBkVqNNEOExIZSkENmZkQNCzYF
I4wFEAWlbdesCFp6FKrNQlb1kx3/UaJ38WCVrwmyZHGRJjQpSZNgxa1IW70AfaMq1dxCTCwr+dAq
UdekVx+2P+zSkdyMERUKNlnD7rJkKkTlRS3Nt9o28xwo6BXfZ99lf4ccnS1w4Rd1+cy+B3pTo4Ch
wAPVY3ZzsBcYQcpFeL3h92kaUQUuPGHHKFuwhIXi0XebO8xIl8L2rfODyjT9Y9d2x2uMp5/mYSZl
WAQxz+ScCj+rk/JEJCoBIsC4y2dhGl5ZHVvyJdFzheOlTu/Qvycqp2Y6v80uEqBG9G2rWwKsuPgd
GmS9JtqW8cxwezPQD34ACWvX42dNqlyhjoX36s8vLYDp50gQ+f2LnudkJIvJVlw8uHhigQBLltAv
KEdHYOtvQFi9WS20T8LdaxQT9bYSm9nILCcEM9Mr2EfBJWlXeDTsY360bsBMvH71FuQiOPpKkicj
Hgm6J7e7qihqM2TroQBaOxk7/eFtunn3JsJ/sKAtMoARIw1ShL3rkHyZjDO9YQ94bhjPE7NwvFgE
59wxL0wC6ZLbZRfc9vbSbfQ3qianOEPXcttzCMWbwSD40m0whYq7Cuu2Qu+URwFZZ/W5jZeAsjFV
n1IKkAQQMI73eKxvPHXfumhITTeAFVCFLnS13LoePa8IALqhVuFZ2NqHwf0uST3ycLMKN5qe2muG
apbPzOtGy2k9qpIVcZO5dFAcvSMffvcQkwp99b2pbou0Upe07u3OTzDoPgokW15k7VAzJLbCybxk
5a5QMnU7cv6jAEwo/9pNkaUzEB1XQzLkRszRTiS3k+UOVJJIQKxexuUs7+EHeneDuSpTGqYf8+if
hjlKw2yJ8gKk05Fq1I9didvdteNF8vKdFPHr000qT/kYNkxUifYvpc/Iews7z8aj9PNevdj/JkVx
GAEyutPT4CyWBcyuslrOeBxucsng4Srtud6x8xtKhhYqqu6hk1GtueIyI1AkrL+3A3aDfVVZvKE9
2Ek9CgoTV/8TWucqrmg6XE4AhL5rI3RMrUo2cR6yua3z8iXhCXuEVXbpVRLgOa+YB3/IbUdXDJsq
fVWPaQhbPAZYyCP19Z+ovILIweeb4sbcsZXR126im4bdkU3xNmbgTsTIlZ/psiLQnp6OY5oKM66R
r5Wmt0j4uRSesPn3trTeICdwqOBlbp2ohI3gydH/Kg4c7/Dd1a83wxvRZTxC0bE7DVpNLEqfS7mV
AEYU9y1RhLYC1bhVebuHmQ3jUVWwGen9HMp17cm5fU4YrF9DlNbH8m0CIlm0/aqdbpVIm5sIHN+K
L58RRm7AZAhXHrcnqYLFpYwnsUoQRm+wv99YRH7qllwCZs0DOCf5c0BpFk7o1oRobMtmvkItQZ0g
ImtoyVmu5DWdfKt0NX4Qf38iKAv4b5PAXH87bpK+lzmzVVvxV+Qg8a5Tij11ZxyLyKg5REuWp9kQ
+wOYjW9Jr/umZdgP0CFFU/VKKhGmO4viQReudPIXhsftWccReHTZ04dcLsaaYNE9b07fCap941q7
7CDvBcJpc+lzmTEEGPBZCmd9wRa6oMIux7xOE7+Z0J7JxyC0tmdYywKggPt7La3IVF7EeTzIBq0l
u1UaNFIHcBQWxeRHSc0vZwd1Ji2hgIDlCeVmHPm4Xv8V26o2stTtQ4dpauVBi/6kZupbt3RkpMSP
3c6mW91zfqpRG0LoV+jOW31Qn6RUq5vw43Ug6JduWBVXffzIBpP4D55BoWJIw5W4bEVYPUcE0203
24jw75cQWiRLOXkIE135oQr6Sw6EU274gZdyT+TkkrHtOt5SN6PodeNou1EhFqNXYatKRI0r2U+q
TP4qPYbmO0aje6Fp6hAeODyQlXmslageuWWJ66AIq+ASSSTftg/8sMpttobf3zS3QsKRI+8ZrR3C
YhOMkIyhmv8blqAyOnNo/8pQetTDe7nv3pUJKeTfkJ/xVFHwmJX3r8NLyFQUISglEZmGsXmx4xNu
R2gcMXNvxAv1Im2s9DEe1RYQIYeNfa0lDNKhk+nobfTyaHCisEdSIb5cQNikSjqMarCGJQwGGVcF
O+VgL0xcDltIVlBY5ODhiIL8m2cfiHBw7c19pHa27dXly1JtJy+BTDDkxVM5yR5tC9XWP4RPkOTk
D/7QFsdXyt7wzB+QdeFYA1GSav27OZYPtiDgCXTBP0t1WE6PBqzc9lyAzqG2q0/9SQmNs75mqMpQ
yLZbGSKaSe3nWXHMlR31ns+oExY2QEqMlCCzX08mDwbFESjZjf6OqSatK5PnWNMNwSS8doyp32Lt
bZ8E5XChYUa1xLF+xThvXgKcsgMrPCa2RqyKG464zts5XW0zwMVwln/tRqsGeb2Yixh6nCXfTrAF
OMsQ9ovEKBr6m0kSsMd2NeyB5GCOA0wE+ScgC2sFfO7gb9vPhuenLfWIxP1qbGS7Ym1cRhivCNxK
mcl4klx9nVUdSR4zG1CV9tWxa1YSkAAkScBMfDo46tsWbIs+1M8x2pmY7NLXsrVLHuKVC973Lruv
3qgpocmKjZNxB8q/toJJcsiwNxipAwdX0+8Y+ZqWFajgTchXDgaLLTH7QuQ+rl0fcWMNzVXNYkdS
zin/Dsu0n09mP5GFcAy9zyHI8NC5IpYukbzsiO7VwKxBjaHk2Lz5kQRGXKiuHLOD26rmwmVCNw9Y
70LcF/fw/ZzdWdz24C1QpRp2osZdNR1lssfQzEHn3esFZtxE3kIUKpMJCZq6kujyuEaE3IaqGx32
aPhFp1SkZC8aImLzKT+38H+KVYDYZjkd7uOTx77ODk4AHWIX277QoO9gR4AViXXBUc0Im4F7l2nr
zVZPq9tM6qZQ89fzbq2484Y0+XVi3n4RwlnWgyujSmJ8N6Zqk2AkKqoO0VwCDfKC8OGrG7FGXb8G
HkpKNaUfkWTGoWvp8F9y6s9PzoTRNhJnqYt3kLToYzvCqfwNJ2VM3NC3oAfEVNESPLKPSGCL1ujl
TIyJKBBbJbUUWovYimyQdr6i8Z4nBBSQb7QJbrFzz2e3L2s5Z2JMkMDX1bj7lnV5hztRivkb4jtc
fN0HpvK9mNb336doM+UWLCUuWc1VMiGKWwJf0ZMDm9qL8emFw3JyN5t5caQOhVgA/HvCHHcBT4aX
Rn+xN3u4hSydtxL5LsADqQf6fOwzZfx+OGHK/zjn8lnGJdWoQF1vSHtVru51Gl15DboC4CqqH2kK
0gvAsKKmnt0rudieQZQ78vmeXxfUc9yNmXA+brv16zHt+Bx3pIK7YG5P6+qQcgwzWwaKcr5+lmoB
9z9qLsmQNHIUludPV7SBA6BMqsF57RM8jl5Mj+vKHvRDpdh/as7BLmjigSzW4XLNrgJTJPF2G1ep
Z9oekuhgzvBSgrus3zm7185iHVGLFSld2MXooq6H3CfiUxcIbLXVgotPTUYcbXD8RHdfr2yDEt3Z
ezmnwpFk/9xGfl9ssfgjyDqbGrkpoHVQtweoPKGBny3xTLysP/joNMeMHQ8WKtdSGjWCxVPOEilG
O+oxT/GK2j0ox1yOCvYg23/Qbj/XQiM6ug8epgK78sMPX5a0bbV6Xb60yP0MavmCYXsH50lFrytS
HuSzkihmkxA5mz6ARgl71aRrJeb6wfrWhz+hdugU8L2pumV+qHRhIFZ78k8hCa7wTm9znqYyrvei
dP/dshjhgMAcRSqSbMOsuqvYYb61A3uphGZY8bmTEGyXPykBfY4rtiWyecI4n7zoXNknoCsCUq14
3gEgXvIUZXzd1NWgrhU02XJmeh0j4IXMZ05K/eCX8z9muDfdPQjvCkMuPHPY0nOs3b0GG4C2luYG
jBNitzaTeGVffYC1fWdj+fxe7lUYZP7iWVMMk3vBrHLoGbFenO9dyz6kwDtip0qSAUiIPCuLkCsE
HFAe+u+Y4winerWJV+W0y4qNPo3NHMMdlJV35kzoZGgiWF09tjSJ119JvkcwGQ5vJfjAvOE/b7cs
8xeLyUuSar0o1+uBqHQarvSeEY/u30qouoyGQsFgS9fj7ZsYTGmyLznyLbuZachCIgaR4XqTn9AD
PnxQK8ijWoKTRSxO/mY24FQDUau9MTb+KtKq0sSSppv+BnwjXQ0PkYghkr2l4S4wLAV3AucMSj+/
MFvnieB6ScWbZYxIClpf75dAW+LLjFMEh219Znxc9gxFzKzmiMg4S6t7iMOIUVVYH1lA3vKa+wZf
Wpt8H0bV2VtdHqJshpZKEiHNq7JRUOV0DadJhxY5N+lFofNLqLDbVeL4zYdb5Hs7+kulyamJgkvJ
iroR57BlvMqA325wQHKARwLX7BY0i6xZspzCB7ndWT9EG9fXPBIvDAJYN60cBfvG8bNORCqcjd4b
soNIPRQdr7LJgdL6vn2eLzNXkKto7UXHYVzBnFM92osN7gmJjO14JJlqBML2K7Itkoa9q+z8iOFN
ItqC1CEBLmIa8ALjtC1e2AogIFfmjYsC7gYfJk+rLqSVcPbGrQ0aTCuzw6BXHh3sNOUs9fCJHTBJ
30zPoPiiiKohFifadESUOIbe8UESJbxS6AiTvDgI6Xs11OQEPGircSzGBO+dBoUIRmDtC7dJOOF0
pSw1EVdtpRG8Nl8TyBzPHmZtab7bzoz4WmJeqqTLeWcILw8hf0yuSesc8Ssqjq3Pqk7IbGa0ZJ5E
ntWA0mCZzXyYW5KfuHBozLbNJyO591JfR5JhxGEFMP6CBSheeh/TqNd26Yqywv/4gnYEXtkyWuom
M1Z7gphOH7XP+9Nkz7+uLpCfsujGBtUORo1XdCAaL13gvf18fXwNfjh85IlXGoR12KABdoimDTMW
EOaC1uJ5DQjJZ2D6l+ndul4pLoCH+FWD1bADCca85mQ+wLj9tkSqZ+NzMjEAwmjsr0Lo8vN9UJCt
OL0xu6gpyuv0N41EqDZNpDXZ1uenz99wOOmx52LSneTiOzfTElscSKG/i6U7ofe7NwJzcbiUS1bE
J2ASuutZspvc01XOFEJhmhaqY1Vq4UBq4OPwb+gqUWK5v9EE9mg/9imZaw3yYM7mJPRE1cfUEFyf
50pZQ4kbrjkEp7ycz2tGl8xyBK9Wlx7pjde2vXfTaKFTdISqeiFqyGDq8qLVNVheysUxRdphEzmf
fSy6cXU1mhpJKP20UrLVfQRuq02OOJAf4zTSnR6lbiAgfmZTSDip2So7QQTJoWDepTzXcJftW4/T
zlKyUQOTVoZLRQne73nZ2z7ES24Wbw2i6jKCJOEZ6rQ1uwpO75BvYfteAP3B6RUdbPVGQEKj9qIK
PPXvcOH2rVUBHSQqg/V4pu2vejJYsOJi+BZh6+MBKO3jBCNCnfoiSy2fSkEbXOEGXgq6d2rsrrfd
jWWf1u/2nLG0hyNImtZXL2kHjb/kzgRZA/mojJAze3C02M8UdB8Vn7fPhnNuy/mlkv0RP6gQqF2e
NLvxFGkq9gH4zCmo1BDPQ5f9rB1Dr5OpSFBbdmCuVZPwrz0g1aWorP2gHSlavuEn3sC1Fg+FJs8r
2H5SCDoI/4o4Xna28ez7tq5CBwYf+mHmEDo/gi3bIHz0yFWvBEBgz9xg3OWEWwpRJcgXVqlZZvuT
iDW+AS/NEkodLRwg53ZUJrrIlZEFie4Dj3/0JPX8UDaWkYHC4CHF171WLDpsEW5YlEDOQdgKJjYf
g7RzAwT33S+CKkbreehTXWlQShUK08GvgZE5YN5cyi0xZUy0SZSXFX1gJnwJ4Dy40o6asJ9IvX82
/h/DKNWJCwOVk5f7y/gVFr3g06loIMbq7sHX4MotJy2BwEZXlJpojiHOAYK2EOejjV9ZUT3wGAE7
Ske28stDPyL3LJxF8iVx14/5mbw6YHhTGYb0JR1XDTLCTp6B3jfjMq1wEkFtAYgT8ef+Pqr5rrSl
IKHrrmjcekkyv5zP7r1xCgZLH8tyquUzH5GOFpbIxojWnFtSIA8+r8ezDpFZ9ontCkx3zKMis/4n
Qi2f63CjfH6EbcR6ZYdCgKGIKSvLs+9kc6YJWTp3WMnGZNYlDWvewXgfVQDmShugjjmNFE2fZpzE
OpM57LUQATlS+k40ljqS3bVsFNJKRvMZRJeJNcC71MLPkQtKONN2dBUJeTev2HUIdsCWlwsleZQo
Y7uQ7HO4i6ljSDsZAjhoxb+FNo2Wg8M5LX0s1XpkwWMqfuobZR17YcBe7Sj9L2mDKw63FEFEjYc8
2n8OwMIrtxurZ2gWhZym+c3n1OxsHQEmzGQW5kyNlDqiLo9Ct33EUMUQ1xFqVFNg6Eb71FnTVEmZ
u6SxZKRzhMNzYVRVRoO3oKi0BvdLdp2vo4+Mr0eUsclukgnlxhgHOXizRUdNvBHKuOgKeyhv+KEQ
GO1eu6PHZphVqMuQZND3+J5Os4Z4a19VxmpNm6IjL8nMUMdQj5UXKZr9dKROt6G1HNgzay19UxAK
5MfEdknlmOZRoWr25J5QwfX+grAJHnxb3Uz0/N39nP7iU/3kvLT0UQplqTilw3xOIRKLuw7k9fuZ
1TaYZPU1E26GgggPcJG2ZMoHHPP5Lm/4SewGkrPuukIAicBTxIs6g7uc277TEPw2O5XEqOaXc8+x
xNUujSgwPs4wthamuXKb6xxu2BsS9vs6KkUofuEQWxykI5wrZ821Klq5SjM8FIbMCOKPLkVCnW00
qwyJq03QEZ6h6z/aRyFRgPiKvjOeb/KC0nyZJHylpCAgN1rSyOKn0jl4a5nvyQIf5oLxUC3mJWDh
WfW/rsMCRwfxtNHjS4TUh9P/pxDUVDvs3V1bvYNl8ZzGjzdMz5WBzcEAK649dcN72A04g/aDIln9
FjGsLh8hn9vt8wCB0+tXVFTOuJB2yrvPXrDla3UH5PKpAbcJLx7HL4tyMnYEKdGo19DpO4akq7B9
/Mq41e7FMA7GzcPrBqr6jyWIM8eQh29+ofRoqH5RrZjFiuwMDnqACXdZWGIXnErk6qGZqOx0bIFl
8FPcoY9Vvu/ueg24g/kB3aet+mTOvQ0j+84XntDpH20k15jGm460CRHbi6FeJl0FcmK7yXUjqDRw
svAZPqvjGXlfJ1r9J9EmO5g86Bj2YyCKNFZFi0pGuWuYT3A15cBqaJOR4anfZOVA+iTjViOhmGVk
snNFud+PlJ7PlH/Rl1L8btF8W6ay6mpT9COD+imq9LMo0dd9RvDliq4loGkkRtdLeZMua8pVXpLi
CK4jVZs1QjsiCFd4GYE5y4QDFVGtVIhbPgxd+tHjA/c0E8+/R5FugSV9wVTLOBxwQxHHsGVQO8XC
PnjSYJojVE2PC9Cb/2yg9HuRfgfrNbki9W33YcgbLoTySnBUnnIrJmSs93wFRfg/EQpc/RC+0T7p
os3u7rnH4hE151LavspoGJygvMY8huqwgyKPEO8i+5hoggzV6X6bZA73ul82lxB+ZI/0dHJy51EY
Ft3IubQe4LnkhLznM09aNSGeTe7k8LlG4J/DIXMOeXvcb2Wh124JApWtPsNES0N0wsDpG5qS3MpX
cUpRjAWkBQ7Z3l7jxTCvY009CZKHT8PYnFZ7pSdVRFbThncoxyVY6d+pHXl80bYqfh8UrErjBqWD
aapsHMpfTQ2MeQ62wpQZ4WXY/LnZbx8ZONHqZKDGuLolOFMvK6p2hGyRFP6w8l7RwExWFFMtEtVy
QxAiczsrrRUz/aSd2KM5/LLjJRVKFPadTUNA6/Wc80zToUWSj6i+0h/VS3OdRuxo4GM2MTcLhepn
e5s/UZVzXUja5+JPLxNLFQjMPp9RaNeYyMZzrLniU1WDyicGgTqwGZs/TCQRSf6mRzzMhAyiTNVB
3M+rVcaXH7lwAOCNr+agR+kz/dNO0G0nvy8SaOaf3mAXt/iEIqqE5EZVFs0vp9LKjW0xGs/xm+en
VrnV4+ME6vfDsTFKrSsFIyvsmOnfeXP8/iNUMNoCgIDYo0mxUvxBnIdRfBondqN3inXHFnb4JQui
enkZ6pTc3Ozu3XzGAN+c4HX9aa3Z4FM9z0DcMXzEQVvVlKOEoyblbN5FVPtAuC3zr7j6qQ0DJMoU
wATlgK3mT5kdNs8c+zvbQmI09km2GAZ1sAzzmC3axDMY/lbpuu/Np80ZO8eqaZG2UYSIpHyBqXjG
fb/7G4Q5YhZncKlPAJBe+Lz4qvNqOt7vE88HH+JxHf+ZzftnI6RbV5L1qQYikjIXZZLkBm5P9RIO
PeDT4vfAHDocMc4iuzr92CfA6q1IiCQJJEj7Z4lGxGSaRinoXAvhxM5JXDxRGlG1rvHbiknbE1GC
Y69Tqc1+1WAJskwYw/BdzrvxXc5nZStrWFa0HkSml5bc7uppMrA2OgOF8PQjkRSX5aXBevAQWD0+
pMVvt7EklPN8y2pUd6IoGlg3YOxnD8cUV5NC6fIP2MXIPO+Ve8KU5S5RW0pxHuwaOBZ35vjFlTRH
FrZXZ0CSmtmxH9oPdtlmXwnh/flGUjGcMGo3jtaKfGTuEY4nnoWlua6NEaINvdWzyWKzmJRLcZSe
Qk0nZD2hhskmpk2AWRyreHtfMy8QSkbxYnmDXmEyZVVQrcN5wQ4nmHnwy7fV32w/rn+sRy+ctH1q
KGTzubbtC6KZRuN8a6Kw7ypaJoI0WMz5Z5kF7ufntQxxE5TseeGZlDId6YeHIb+LorA6w6NTLSkJ
MwXm3pzgEMQpxMxPWEUCZ5eRRuG1a2yjNgggE63RI1I8seVQGFZ5IsIpNAP4Z/aGEpMQM9gShow2
FjjzGKvOk2YAVxgcoqPyK3cdfgFfohuFRUmbo0uZxQaQaWzUXlnIsF+Uj0hLB1c8CpnMs3R4NQ2S
cdr8MV2PceEOa8VgCm9jSUJoK484lcU2Y1NqR2NngarSg+7MSgs6jZt/WP4uyVs2ypF4/R87Ykrg
L4ww9Qq3bNE6+Q7tvbVzajwr7ZpPIoyY2tgoiBFUtkv8Xs5nI8f+gU3YRT6fx6oBltfQWSEmW3K/
WapJJzIOSz6IfM8dSuhZD5jOlilttuqtXxH53GjeneOHdzm666Xgr6dmHXdO0R2zSd9dyTAWJBax
t3KYYEu5+J1bxDxOY2GX+oFLfQMc0St6WMO0dGeIvp616m9DoijPLjYQE25fJq7UhrdqI0p9OTBC
s5elp8k4TygBCPgM7dZa+L6nSBbNgHnIlQGQSir0HwfwGCASNFqcZM6DySOAERNY2ga5596dl+rt
BaZFdTSqLpLovpx5kjtQayGEwCp2EgIU4t9u4FzlU/ew0FIJ3hSBJgm3g9C/P9juJO6uuo5NfHcL
NDny2ZW4ISfMSsOvyWFS/WdKRyE5N4UMqaghcohnG9k5sb8QB48baq5T+yqFrYW0Z6BzCF2zT6JQ
LU/0ewZ948JTmEcLmkRzPOg4sdmgGNwMKuAs9sXfUgunFpdVOO7sOs8tbu1Hil1oSld+xEJB/cyW
qEsuAySrutcIByhCbK4SLvBQhn+DQYzSRQlxjYdJuWBKUwcnBbd6oXA4o47a3e9Y6CAgTZpasTlu
XBxztFRYEzjMO5OnOwsgI1m/PB5Pk6TxnSvB/vCQaI64cI8XPAfKbVBRwLG8KMyve5vVvcP4q3P/
5oyVeNriuca3xBFWOsSx+AL1mqWrWPw7Wl5NPlZGh+vyt/XVaV9M+f2LJVOt6kfTfS4LrQnSM449
iKyXBV0OGLeSNizcSdUnlWEqJHOp7DC1fZ6rgMNjhEw6caBfhGyr0mMC5u6i49ACyOm4YXvlZp74
emE1vixGoVJZaG2W6QdJ92Cq2cytx/PwCW1xIw0FNhEh0+F4c7GWugkPEL7vCYbfWUcIqJZrTNee
/feDwbBpaF+/ezXVcHiNM15mfSuvMeM7U0l9C8S7Q8GKYv4ASI0t0Y71AvZlaieF8X2MZwsosar/
Aesf7W61i1zkbyJtHpy8joa2RPBGf/y0/1l6rSoo0dCxr4vaNbLlI1K1t7e6dSt94lb7JKQkDqwp
DtFUqADApjTEYkqPxLAzz2g1YxETryLiuvk+RVLGtYDNqVPvMEII63MMTON+DtUVmQmCHJrvDezp
LGE9zBQwi8JZcw9ry2ffQ47SzqVGgr3KC7kTwlsELUhv4yiBCmjKhA7yQLddatHHgiKNCXIAPRyv
FQPyNpTFpq9Wau2lWGTZlN+Tk910PTGrwNLb0EHoL1gNd2UKUtSWjl+QSty89wkrbgJiE1Ng2vA9
Z/YmSiYHXFfKOfRAG/IvBPKDKCfmugi3sNRqch5Q5D3ZnQUh6DXIrn67y4BCj3D6zGVBF6+rL/hL
ugtNCdUkXORhfZZ2Y2JHFoGHKKR7jL+Fm7dH4NZLbKOX3CiM87Q2A0eIjdRn2Y8Tn18XxKEbHsaF
0ZeqJbuNV5G0uGeYO/CRRiTs2tI68Wa0vxAad2QR0xsLczS10D9hQ8+FV0AaQEJM1qRv0g50WKlK
DwTotPNWAtEW2gRx5KtEqk47IhtORqwa5KPtR6mtUf6MkGDkDpqWaddOd4wPKaOyQWluYLAAPD95
zzSpnXMxjjnLylX9mspjKY42QSsizEicxIEGhXZrIZ7fGhzGSnArLuNS1YkFPiSDJcU0A/Be12P6
3o3X8pTe1S/SKfnXCV2q8CTz0tq5WdwiT3SmarWakyv9iUowboUo0pL5Xmn1foD5pAhNYKQ8z7rl
AOj+5w69EyeJ/lE8q+2itnfg7Or5oiF7OvoA71I3sgZ0X48GEQCxLYyjvaUfQQBF9zj74H3jA8fH
MZ1xAfEMt4g+ZJV816GjAxSGy5kzTgnv5l5cxfgQ7M0WfgugUVeukhQnXUntuExbYYXrNK8SdTRc
yVDfGfrxycOg8FGsqKB+ZqfQPSr0tteoDBDZF3kxVZ8LiVRIDRQ6BGgybAl7pVCWe9r/gq0NLsM8
dn52A/MB1kyA9BUBdosPp4YVR40MQP2avfwM8GtVXfZibrizd3WR1HK9c98ilp+gkNuM9JVLc4o+
S8Gl1vPACRqwfuUfk1cAXzPQ3rrPhvhHwwYe32C1/E3SAbt9w07ZrsMjV+skoLpe2fda6aJCYkZG
BdOMS4f5egt+Bqhg971iC+xA38opE34Qlh8QZb+j9V1ZWhw+NE5yPXfKN0aTT+TB5/694H5CgK9U
CDaal/p1JEXYHGwo9euLC3Xe6fR5GigLeGRiIR+iLe4iQJBYX5a+OwUY6RKXCVIpGrjGwZ10PY76
O4x11TapE21o/Eor+5lpFGFCs44Hgnxax5CNGGUG0GcWnyO3VsGsmyJ5Z+SR94LHzNHMHfw23RGl
fbvRAUDcjqOr/zag2WB8VqzOpn6OzQci0hIf21dYZHN5rarw63Tqum7pCWCY4SLOfrnrjCMy18lp
N4Qyu5vHwNoPm2WFY9769ifW5NyR7FKcN001qxpFwx1qT0oVTwYTdPcE6ypXvcCJg/opdIT1H58f
ND3tV4Q0LTenQy4GJjWqjPgNpTghsUWScAvFnCaq6Jvva69+q4ISwCyO2SiH79CB9qtTzxjyagEp
K69A0ChqPTqMguFVa6tsoU4+wKERg4lUaAwiCBCBLVBlLoS8Vl2VdanhfiEQ/KCybJ31mj8ELB60
U4lJR8haiNoqaQgwpsJKp49/yBRdHJHI4W2BkJsamXFcszyUMOiHe68HcRtheBRjHa1sfQeSPPaj
FqG6OZxkEJd0vmZqCxDVS/koSEqTGKwyYW+t4VKrrSgzwRtql6xz4ebK9oSEFnA3vACPXoWJ6Bcg
VelZvQveVrU9ZbkgVOVk6dQfGNZ/jQZrmq9frCHvGASdjjhTeC2aXtS/BbPmMjm9qdupDSCgqIfo
+jLRXGLzN6zx+L0sCHqseg4M1dHTgAlN3bVVy5IWde8d62AjI9RkhD7s+LdkuyRSzk/MabSG1jXC
v9J8Qi9XbprjXKHJhEfFfNeWZsegEspC+I1vRaS5R/neBJAG8o4Ew75GbLknMVV6iP8kxCwBlxjW
cuZgQit6sl1lJn28fHKFjY5vnTIlZZlj1/QO3M1Xk2dccx9ruWH7jlfDSss5BB1+F9F3OPm+cSIP
u3N7xixs11+21SefEqJNEExTHnYUSF17plsrIlI4aN1Bv4MQgQjUmlHLqCSJqoX5aVwJljQNBihO
aSk8+vqQ1J1Vy/cK8V6DGTU5E/paISFBATx6k2dCbBbKc1gLEXsvjg+bI9Bf4EE61Fj6MI66bC9e
suVkcuybkLYCHMCTH0ebnH0XFEd4wu2U/GxlzKIKjCKUavtmH3vYtnUOnR89dCrROGDHxX1YAIsU
8EhQL5VRWMg65mtMASjG6/DJbRug/fan1qgPk0gpGGvhzYFyxtP7B7EKJ091RbEzZ3wc56J7Hj5f
Y60IAkWXIsQ9JY1wlXFikhMJKCrD8yHTNEss30MOOfSHER86ctLP65VHFtIDCq+6RbkEQJHV7Boa
nVYbm7swp9mSq+aO/DWvGXpCbahOA7+nsKKe6lTfG8ZGF8nJxMPBryq5QfVUcOV1mvYpnSMHsZ9z
qf+SzY7TaM3+WrfKarDd6XxzAiT75d3xy1i8ougIaRTOAWJCAn6I054BgSSxh2yz8nv95k6Swzij
M0OynPtV6Z3cPVFAUg5xEyUEB5Sk54z+jnBhdVx7jOIr7NSGYdBkjV2BVyYUNOMrCWgdyavqoM/M
PiejT5uO8uEBSrcF/ZzAOk3Tl20YDZE1X5B7+TKKyn9SNPvzAPx/BChmHRhuDAhpclFWGGNBz3pa
CiyLJxwTpUMKjzQCsQtpfbsiBju+5mtjSjzH0xX3+tgc9mTl7YtKOQB3xlKJezP9Sx0zZTYsqfdU
s0HXNxkOkRezIWijqJ9Hhze63KPWGrHBqu/0kArWOyOJcK7iisqUh+S4RYz8/ugUi0tCsJA6fllp
9MdN8NCoueACb2iRtvkb3+o1wgYSroR+Ie7Fry5LwMV0yD3ai4KHexz4e/1A8bfx/qzSduGNWMiD
i6cWjKu3Vc20iyru9e4aOd09Boi98hd+yOqcKmfZl/w/LhlyE4nHyDA31cgonnOse+2KMrRKbv06
HzR4K0ebqQ/ZKZi7hw7AA3z5bbiKstqFgYpcEI3pkUxpARrYkRy3U+rvxAGwV68xiaVkbv62zqWh
S0+5aCicLO16a54qDaGRmxJuir8f1clCnYB7JiS9+N64GuhyPxYQ2vQXTOPxHJcpzspBo7s0e2Dk
SMWPDHVbcRKL+WBmnlPa+3AKVqQRqd9bEqibXVSudWUDarlwsaJShm3cunsehGP6RgQO34Rg9DrG
fw6m5Xk+IPB+L1rodo4IscUdZFG5k0GX/11ihB+gw90h4Nj/V0sErIJrJ2PbapwmfProp+GvJ2wR
Rhjv5QHujdZ3JIF4AlS013kq9aWReywhlS3Ix2cp3w0Dsntp9m9qil/jrS0qofqOA8NMF6NqIxJT
IoOORK+tuslkF510R7efzhBnhJdcPmO1va5kJtw5ym7fUtCzgbrv7t6r3MkgsWEgJpo9dfG3yU/2
il4pSVCHgWXob5hqxdq8HSGispNtmeTSbA6lU7D07DqJ81UweRXJkYAyaZjGqkvhggyAVkjMe5Ld
8xXE2DeWIkCN8O0/9f40Bc4rzQXiEvjjqGx3l0ZJKx6y1ivny5KE/v/QTe8fEzrxnrdMoJ1Tf+LY
9pa8HLoYY/EX6ColaJAFekrBmzHtFvkYcD8HTXK5793B9E25JKTz0WtNwJxffC2PmQasT7b7D9+I
R9iBzgFAD2I3d5OmzzHcsgZUzXd0uibn/7LZwr95S1prBMlNreqid32bEZUr6x/urHoKQ9z2Evpg
pXHzaHw4LiuRE3X+6P/8c2J7p//vcWs+8XR/8IxKyPKZiXF+KP6MrW4Tdax1MXx//EW09tneTt7r
d9qh2FyXY7t9E4Glt6PqPb+nyYq1bUBTNKzjwZbiu4AdLOu/BsDdDYfX/WOtGQZJ8gV2kuZmwJNA
BO0GLgK3LXAyERO3mIxrl7HZ4fU7X2RwbJIbZILk7V+/7bk8vmVQTGu8UXlZ2ZS3xp97wdd/WEZQ
5Zeb5B7F+h6+pORL/IR/sx0hxDZWj0XmMfgw4iVG3NZIvADn1HJMpNIZ7spkIIQpxpPXSBJnExOW
dAe2kDASAwxa1uXfc7gmwfIg7Y+FqwI3YXJpY32lDGK1Evtw7Dgi/XDSJHM/qGKiNNE0TqY0zRhJ
RjdBZ4E8LenKE0LTr63l8bk/VUuQw8zGdMaIZePFQxo2NeIsipJjnBpqVs0TIjdnOg0r7w0TrFLY
sN2Gt3teZMe+jZPCYvOmS6RB4y8kQGcQd/rCxQ217b2j15/8biF/Dk/v6+V+ETP1EW7YeIWojodu
RZ+AqYx2tIZ5Gs2XdRnVcAafmdInykrUhSFTodAE96uhzYV8N7lT9NXerk+TWzUkthNmEwsZ0EtI
YGHOGbO1CVQCbvvewvFZp8gg+59TwBe34PJLRgjNZdRVT7e8r5qgXiBY+8H8HosbOjUhfYQ3QfYR
7uH6uX3HpblA0Ikn9hGxGTkEuRBXlhF8uQjjdsRZoHIVrbZQuGPHTrShtH6GRcOv24QfcKpwhBvp
RIZqurnRaCCDW0QXaSQdQVDEcdYhkjrXySKr0TeQCgmUDKPhwXAf79lIirA5hqsvhLbVKir4JmMX
M4zMkTt5j9bj6dd7SHcX60Exo5EDW9MFsNahbzZu81Qhk1bDI2D/TnqkALVfcBzyzOqQQe3gEZNr
hlcgXKIigKigbrJnMvAQswntYoID8l+S2gtmFgV8LTg+RrvyPvc8n89u6nY8hTe4tVaMhpSTdbC9
rcsqwMRaVmvJZjW7kRe/cpPe9V2Y6UIbIvsasc37XFSyiMiVl+7eX9IIOapMzXWKgB8FMbo40fn8
f6wNNyb7p35HIiSuykvs/ZzUw3NEc8cs+4JwmUfzEVIL//gAHyq42a4aDPGqRD0YXqNOQuWiEFRJ
C2Oc1swundxsfCLogssIoLf6Qfj7CH7rYSe91MdUWhj4TiREpuwofL9O1IrGpZCtDjtyTL+1iRjp
LBrxjErPk4tBgtjfL+GswmdP8Pz2qjSRT2VlJQjgUoh25WJbtzW29NIHy/kutPFQ//2pSAmjGyiY
CnR1sxmRRMOlVjolvqd+GEQIur38/CVYYCSy9tNyQ5lRVIrjxriG8ntXN/jnS/3PLGp+Du+/1ibk
lK+n4+zsswuA3q8s0gU7quu1SgA8/liEtNpbfuAWzA8IKLE/PJV7F8Zie+4GWngLKzK2/z6x2Nas
RlZ3Qhh9dRaU78l9dBLcfgBrOHekNptWnNKhLGupB8pvj8dwEY/ZAwyiUWHp60c/yHv+XSR41tIi
rt/rBgs4rynLevjGFJ660rYBz09ImiONlXNkVzkJ5QnqvRFFueBUh6dPfFGdxPz0wzH4woNZQfPW
mO4U1K1VtJBkml9fNipk4GtkLuy8S7ndSKKTEUOT6kuknXi87rMa8zD7bmJDimsAXcZUc8n4E517
PoHvEmV03PNVNrGxRcuPbCbkQTUiFmuDqNVajtYypGRmIV58LyShCklA4Q1IcuV3glpGDha6aaPZ
782weDyKNBRbJl01d6Zz4SNfoVBnIaltNrziu95eO1xmrNii6gNbQ6CFvIOZ4NkIjFnOlehney7E
7utud35zYyELCzaCjOytoB7yEoWBo3ocRGlgqGouqNYuzhDoZ8mtejcHJ00f01NeVtxIQcZrqsHz
XTb+hTlHNmNcbkTGRFYreAAML1kp6X3aBNF+B1qGnNwNWkK6kgcbE4/NuaaKLqkNaCUKUdaiW/QD
Uvd75PXPi9LKBnCnZ+MaV5Lh5g/ki5JA467cfE3UAaIwVQgsoCEQAzxbb5Oz8VIzQrLR+y3jKzIH
p0ewce/3mKPZmDYhnqMpOu3+VvWwgNotASiZCTjaDQZ7tyONNQXm/rxEMZP5NIhftSdddtVR8kxt
cTRuBDucRwOw/vTXU3b7hdgarMTsaOHD87obaA5LtDU73UnUAj14SmVnol0NM1GCQyG7XgJFQp0C
/0CWBMO1EY2X40uR3PJwSWiaEpCPhGh9VbjZxqK5pPeNGiv8yKEeA//8C6h+XFnVxOi4S6o9oTz9
CPKEq8awICMvuRLZJJhjSy+3ev0r7040eAqCIhDP15ic23rogHf3TOmO+FSiLymaKC8nii7g6wgs
c7ihE26uZL01wdRwucJVcjmWX0A06DPFFVuFGOuKjhWSV83tMKeRAxlJIVUXJV2mGAKfTbEdTA/V
72DoIS3f5jCADoq8udbJSbyFKQS2k22hBYnSAsMGb9Ek707yMlg1VO5siAH/Nx6VmjERUs3QMGiA
Yiwszxe3j+Zq9D7NFCTrnMVedfEFFmnsSxNdW1DskBDKrK4AYJkEl4lUOHpARsONdJ2/EUILOq05
eaiis/TiYAXJX0q56KPGCLTD1Zl74wUra5ZQIS6w//gC5lp6ExS/e6PbKfrTwW0wrKnBHp68sUba
Vl4K+Wew7shshMx3czrGzYYDfdeTfMftZAyGuGNlxZyOFZmSDWdwOI8okTY4ZV2sP0C8pRl4z6RF
KcrJH5wA7EdL1qnsPYf51OOOdlxxjbEJ9zOXXeMGHyGGVXaAYh+UH+0moKMAWS8IT2m8L5Ah4RT+
2dYidN5v9ApLlOrtzRewa8MiFnqCupkDTxaInrpEbpoQx+bGfyOzQ5dvSZPHqCATGV2SJuzrAIn+
A7vmW9s9kD0XyzmahZGvuKZ1QSG7kO+3G5pU20pEgRBIEESAElB6QiQdzgWW7P2FHgIom6Q3me8L
ND2pV3f0VxumicAAMmpLILrXITPXrsz6NW8WbqdzT18Q/ImToyXyEFNGvWW4GDRO8NMmE530hQcx
qiAgV3oUKmW8zebnFS3GDC1pWd3rleetPg3QVPl+PnX2A0mRQbrKLLm0merYMYqoHk9CxgEglGJS
9y+cnebHeTj5g7i8NV20VZM/Id3I4eZcnitCIl+T80J1Qrldv+JjTdFiwiDMTXec75DpS9ZlkbuX
Oq9CpII4MeI9dDilcvGb8jwJCqRLEdCQ7QquWgmF2KQRhEC+zo0kUtSMNz6+D6FRS5gJzUUyJC85
1B+ynTLPbz+N+U2wXkGiLz27CzugW6mU9bGiH5Rglxj9TH0MholJExVBdE6F2HY83akUKHYGC7x2
j4HVcuYKmD/WMhlSvcw74BVoKhJTxS9jcfELoouhhOScg84Mpl6r9SqRH/Q9A78dbx996LsTyL8c
f6qnc+mbMt9MinJUMulaBhKXx2RIUs61s/eUWLuRtrnlr86XOBLrpKMUJ5QvDdMoL3hhWBGomfI6
iPhJwDG72pcy8AkKTpawHAI8YM0YAtiSoI5XUWIlqv8itRbUYlU3rnhWgu7amw0FZSxX8WKh4yZb
807JI+to1D7F7wo2dSkxVEWKwxBG/g8ZygMn34pte7g/+c9jqEKy0c/Q4kB0qO5WeEKvPyHqkvmS
66u76n+gSfEMu4IR3LEpBTzsiWO4TBT5wfYQz53fjtbIoc5eQ5uAfoPIYFHh9Ao5uT+Jw6WSYXWT
SnGzaFiSnEi1Nepd2C4mcP+8h4C7HgjDCve4r3zzz6GMgc3ijd57OQpyZdM+xpqntPe/04OFPXJj
Clsu/wbwC7aPaS+V+iRGD1ba8lFeoZWN15Ay4UP3oJkwdLdVzY9P8LaqBBFKvi949NKSUQRlTz4W
l4qYo9TUydsx1rQhNuMr4d7/2ruH8MMrgK3eMwX18j8o7O0hWRs+ZAmHmI9rKtpuIeDPzCKCeV5o
rxl8Ue2JL0wbQwv103bkSwk6+Eokw/Zel37KdOBgcPwdlN5lwCTy5yLqPONo8eL/UrTP8wt6SsQx
TVlq6jLZ1O3i12KMTZqGjjuLZo30Ej32Yh27w+hGUyGDYUb3J5+NBtm/Uj+11m6Mk8lF0oObG24F
m7FhjMov3cMr/EdLfH49ROCGcgze5T2bS57DG7xrtq5/rh3I9lX+1e4iD3OciO7mChiasRvT+ba3
yGIQbMsJzo4+ioB5s3XlUNDHXGA+MW1LON0KZnjxCIKnNMUHwZL33JDsEXDrhXrKR7bzPUyPuuov
xRbo6GxeegtxJkgoT2G/aPMH5jdFHIHD9jFxJbSFJ72alnruMCy5NDZR37GEIirXovYB3o+HPG1p
8F3K8sQKhhmZ+nt9YBvw5xSOJVPBrHTA+ysXlSFYcFKbeqWALejx+9UqpX8orVWkBoEYIpARUgGe
AGeys34iugUMDse/igxblHPV3gXYtFz7hzvWyE/a7HEfUODcbDq23+tSpdRxIn6TJ5A1ycgIG9Ih
MTCnPnpQbtA1flv5M4VWSmfz5EzsziEbIVuJNFVLoU39g2PEtRfOYEne7xhAwVYTZXJ6CWJoA9wX
9PpXyEW3mHgnKIrtpJh/lDnKkk9aMjvg7XjjfumuhVJAechK5ttuFy03pDKnSBstOdPcgTSraGBQ
5pKlSofkgRGzJybkN7HNKpl091HgHmI5ScXzo+6qvSi4HysHnrUvK1TYkVHhZBEt9MFD76aQIQfk
FNKl/2Lh+GQrpHyYmzwLkrnav82+sQkO7NfRFFWmvUAQVYWxoI+xNgF8eIP38MjBFWWmPIsITbjj
EZJpnKiGv1QynGwnJ0tdEHvtgn0tGGroUuVOl0U1jTeNlpX/FOZCKkMaP0ikHqpX8OZy91sEcwYd
1hk64ai0fZ8B+AQOSFI0+nhrN5wJfvbS7znSaxfEqBFFY87X6kEE2yJ8f48j5NDPmg8GsHX3XnlQ
hEhefxeK6MZfUrIFKtRqyHQFARKCo3Cqp9KvBMwiVDtfcOaIr6OPcfITCBY8p5MQm0EdREamt07J
Nsz0iMxnbiWGOmv0QlRBYbhXdz3EOPZdm16hBfaRGczf8MCFLtEn4oXxbj/Alt59sqey3SwLuy1W
sQQ123yvL0/uENc6Xo5KHQldWvQa8S3OIE0keiRyCbvH8ypJqXa+1whtYXf0s+3nDhwGYUSikWi7
2l4iHVyUAv+AULsLF+zwg2aQM4B6OYH1MManYIQa4+2XsuJRUyExJ6akgLCZ+bIQ1LM3Rj5OV3OP
nTeBUdKdsgmy/3XgFTTVtL0BW84rorbfZHFRFiIRwMxrxVtLNXJyG59HRToC0zwiIo3O3rKJdhUd
OYh8sx8swzb7cBnwFaTVA+uhP+N/dN2SZaQM4w8Cektg2BCUcvUl1T3K02NY9hqrfryJ/QmVXOiv
Yt0W+1eP8Y6xP3AG9enVkt0RZ72a9aWsB8URyxE3jpIpO2pkQn2rGWwIEe6p0LSx7L8Z520I4Ftj
Urz38Hj3Gl3qRSSdiZR3fK/ww+DQgF+E8+1i7c9XMPiVImEhmXN63/CD1mQ98XFz9gxXa0+F/iMb
R7JWL8YpgpMszCBfwolMdSD/ycR4ZBQZ05/PZUJgXl0jjxK/5c57YeSRcu+qo1oDS3FsvWttDTRx
vi1Ptfhz/W2utrxPYlFxpLomphz69qdwp8V5DUaw9FEnspZWYjNswHldwa/5G0pmb3tfoVBH5tBr
BcdlSVjpi313dTf7s+2zX3E9TtZJAbijd3JE9uLYhCiKAg8GT1UyleQw/iSCusxowUNGoRVqUX6Y
cLVuZqdETngLBMggJwwqA/rshTjUmnHA3QRG21LIteFCvhfzMg4kuYtzofS9feGYck9CKD5nTy0j
OFVlDcv0taMI75to1Pc9k6GR6HSRuSuiF3PQwFUS0bH3RdtrTbzA7GrSaoB22NrV7Oodw/Y/0wdz
3nebYKbSryta38DolUHWKNs8AROfrrIjOZCfTE1KO+WTpaurqhhlOibyFpnxvRCQ0bv2erqQo58L
EAfHmXyjBysPBbItMMM0tqI6Mw3ccsyyGpcZRcaoGW7K/P4iNAhbDvgmVLBIf/m3kKm7KOkrbyy3
m5hiIBJiuDNrWt20Nq18cXt8KNwELrvJprqkK4lQDqDRbi9pcbd5apL7k+r2spXzvyCFsJh0PL+V
fcUONaHEpvu63A/qXYY0hjjb4CZHHqYpV6KEnuW/zpvvOfTSatD/sXAH7wafI5EQCVxtymo+p8lm
uB4KE6+yBGbkFjWltP2x3VG7s4OhaZXN2sDz6ZtZbISr6k2PnMaLryVNlXxXimCo909hMLy0Um2A
XUbB90emGwKxTXJzPIrgreomV4A9FoMmVL0jWALdIMXCZmVJf4S6Ub5c54ZsBw7/nYPHLyDze25e
Rr9I+uyLiIbMpt20iO8v+7mvujx2v18g7m9+oB8Vm9IS5XziTtob+mKmLRC3gwBN/VW8jp4lMVD8
Y9J+rCBLj9WF8IfF6H4cPKTv7/TVXrchHEQ/ev1EuATpSLxeVwz9zI5o0wAcEYZP408cRYtvleIM
lc4x63oj+RRHyyLFPfZaG1nqfp/kXIgCIiO23O5JQ0c73TuYoaaJI5yjWhBgqYJhTqqqI+nuBi+v
OunsHCxiEMHjCuqzrJbSNSmIsCAOgrtfVOoSz2Ae+4nS2IzZL+8SsLxBmQdweyRstLWrSCtKePs5
otto6Q5wu6ydx5uqe5dIXokGqylmdahszv6NSd2d3hAiBc0jiAwFl7ZdTILlBHQufqZMiXg1tbLA
sUsF2sorEuGyqrMSJy+JZSth/0gnsjV7U4JxxV+tXa7HzYs7u+LN6cEmv1T6qvYqtvfhY2KFev5n
60z7AHH74WIHtnKq1RQ43ovYWyJc0E5hhYOl0KPUhYuqGCN+TbDwSQ3S03082znuV69saMPcALGi
Q11pwIZJcXgCjtFxQWetT7pdggACkjgd5CsHMikD6ypJVa0KSoD9svj5rRFRuRMmP2UPooWRMbfc
NV6aMlKoOZtgZdpQMVPfkg9iV5lFPfM+xyBDDmGLx2tcuFL1vGC4cgkMzVRiicuD3B0iT6gwHpix
wMrPkKLjUWhB2Oioumqhce5rcDp4i01cyN8OLggkl9wYbYyqvN7joN3PcAS/YmeYcnaKZNAtrE/Z
bcNYHd+ZN7tFKVcr6/51fHA6uSjHL0SOumZgqLcB6taQoAsbCInXmeP0wgPxSG0nGLcXEpPic4NW
w50083jfebSB5tjCukbmcRVNm/Q6OQwbPEwP9LpwGPY6egT+LH+ZwodYVe2FunFyIRx05CW9BwgL
z4MucXhHWyIjsRmCWnxhTIu4zg7bz4Qw/nEBmPxZbc9zMOT3jvf9Mv8nCGymFUa2w8XPIdz5Q98X
xSGRLM9LkKWfUV0Z1x92rA3s6jX9mCBKd4/uSRUBzZMUf4mx92YTnhptZaBg020aKx6d5cJVGY0B
fDx3r6v3im+d4ocEkyoW+83CCFUEjbytAjNTMBjRK0eubbECOdmwvsHJS/AtsndCpexhIT4wI+j8
SKLovw8kTTkCQayH2Rv+w8lQd96bq8U+aAPInLb2MjgmN2dQZc2e5TI/ScPM1NK9YmOXk5O7VK1n
OqupjkCqiYsWOeeInXoDN6N9p/u0zNwWKjuugWeC4lZfOh35cg45acdfAO4L2ffPpNdbueSpvDBq
mLyYj+bFvmp2Jhkvrx4NhxYwMyMZAGZKVlQ2+qgYCGqsc8lP36/AQykZlgKlrguDzou5oDI12Tw3
7IcmN1N4synnX1eVLfsDrU19RxN7ObAuFfwfChLl0H/yYjgUn+H2RSRU7FuAv//5+JQIv5V7BBqJ
jFFp/CR7Q3Zt8LWCUa8y1GIJUEaQ91MNF+AUMQ/K2/S2jwOJoJ166yV0IfqyAA9opDjan9JWfOrp
IZFK4fPVlRgFJlCurgTlGKFgphYnX8BM21SgJQDN2+TeJUPBofmVpD/mOw0PPPGa5fglVel47y9a
vKQZL8AJ34aLV9UadDU9JUl6ZRLAuh9EZJzaw38uz6h9yP9UwI9EfMiYz1HfdkkarjogLhccWTS/
yeCnFzwZ2/8h2//I+vvvBfeKKqKqsAob8D16eZv7ckbtNAHvnvDW1iafZ1QptWkjj4kOQKXQ7zrP
9vXGBkSjlB9QGrvJs5355owV8onOZ7yUhloOMDQT51HE/71NsXsvhPFZnHNzyOnJRTTTVKWmjq3U
AzS4tG8ND7DWMFqmrpxr0pkQZrgjT33TpVB3B0Q3rahItOyMkYbJGFhfV3s6mm38BEeY+0XfEqLW
ANlDU/LuuFKETbNQQrsBWq+PzVx8k3rIyKV00vu72iFWCmeDTWk8o1X5C/xu31SxA81QqZSmJNhn
ip6dElZYcgRLVx3BP7CFUZG8zY4jFnXG/dofNtcHFEPlu7N8xOk4isYVLZYb07IiKT/hBQ8S6edE
t5fkSVnWG8KfUF41Y5swfGVB2p83C/dieUk5KxOlp/KP5/eGMllmTF55ePfBRpSck/s+DAdVhtUF
eoCTJbnX8dPif/bYhEzf+YZOs5B6eYgaWHtsz/kr3RJExGNvCZaqXHg+3YKA04x+zwOHeSfecD14
vQ+es2jmZ7+zNvM/GFWNWO2GptArZv/67vGLTvsKi3PZgfw8XLfxkgg8kuvUgFlJs/jQ9HfNtUGu
5M5WgGBjmkpwV5QZwv+unxNpxoagF/cqllmM9vOKEoxuCWua4Asv89jDEnbG1m5GAfZ/1TbZwrON
G6fDp0FB5c+p4fxoCo77VlcotXgj1THbRl8ZS5kfauuAaD/B4ApWm6NRLsagzibES1LkvmMlGR9v
jOYGvJqlCQ4tldVDEICx3Y4tiKvP/JoW9f1FhTxL68cP7NRCqPm+1nV+isHpDevkNlJ3t2HnF1hb
VuG2TotNjo16D1gvjekHBwDLulPB260gGg4eIRyMzxhY+7mt6z9XJ6z3Wrf/sme3Ake52rUbsImP
y3Ut0yqODiKi4+MWqC2l+vBca2cRXCv/3K1nBA058Cl8i7IWHW985shtV8UoJvTuUTStIPBEAtf1
YBjAscOeTYqdjLp9AEsX578B7ldcN++9tLzbDZm0zC5Ommh68SIunvPRghjRjqNDjTBI6lCgA+GG
hFbiJLwyhLo7WNtTCtaPRepn+AdROwkMrkxnZeazxF9iqDUdF3+OCmZBt+e4yxIF9rG/+gsQ+S4Q
nEyFC9Jr3/1l8tqrG8kolR1Bnc3ala8jnSXeUuZNJX/5OH1ISvjwXP8XpSE2phBeQRTFrj15u5ZW
AAWSiy8Q8hQGL35jLREFwemPvH4I8tyQDrCsRn5i4ANzLEH2sf9N4Wk+f3c6VpBnzhTYDC8vEIFc
pZ4QjT/GnbNseFm+AQtvRJjhr236t+zWicUWQ9C5j/cFoYfx/9DDGc9L1tSpKhVbt5u+FdbRTGNI
LqHt/lIL88whWc7x6KqjT8dZkqbB1OMke4CChyOMpixcmOQgANGOrKF4GFf+XIhnN+VHKlf35L0r
VBfLXxdpJBh/paXoBfdE6E6kTml++cbe8JLq0XWijCEwB519bTFJ2qyC4G4FsbiSziSx21cwsPaL
PJHPOZCS9y09SbEfStki/9akSStClALpzQiNNKFILNDHf8+R/aws+IkarQY30mp90w86pQC0dA74
9P9FwTKOAB0hguhOVI+RfACCdi6P2GQinKI/Zc9MjNhHM8a2uC5QvOgXmI5bc3BLIGUm4CAhrC+Y
OA6iLgtYC9DOAkkZaT+p+5q0L8IqDjE3dLvmAFdJ8e3n62A3MLGF5tZJCVuTpawp0HEeuWd3tClE
+iMc8lybSyocoQxLge1KkfBmiTWjPyv4Ez6EkWzmHPib1Nx6Z75rr+fMJV3tOAwSTc05of9zV5Id
riK3yYTyYohVkBstw7IU7MOPGxjtOroiWQJrVYEZnnERkrT2c2xdUtBGEolI5b3fsSlNwS5pUL+n
aIb2mEQhkYrF196y2jnbKG7WW8y6cLKR8HWZ7pOKnuZMbKG/b6K1bbTdVJ2paah3BhfzAMHGMF1h
JVubqb1S/5J4066xgMEOwAzfb9DW0QrJJadk1f7Pt+acJ8kCACkVWDnQcbgOA4Cur1xh332reryA
f7DZGE451gQsDAkBI4Jzm0beEUe6abOW2df+cvZGaRiMepqAioMRsz0xlJ1fNWKpA8j/F7wUDRo0
IxmTfNVYvgh9OOPiF+i0RD+tX6gXuVu3T9a2i8GRF4elPJwodQgHZM5MbsCa1kggRvj3Dfqd6eO1
K2oVlECxjVZImpBXtB/QCFXgwysj6kCubQVIzejiQaUB7WbqpM3De4QPv8lSu3dp1D6kNPraVZTr
8D10HTlvCmWrTCjk1vSIVkWrHxtds5tI5xysLAI3GO3S6fYONIzU8Jp2lk+2AtZKqcAKwxP6XZK3
t7CVXs24YrmaIn/Ihuuiy4R9BNNBFEle8hCC1lXQSdz8UG0IS1f1SBImmqHTq05zCQPpr6kdJUMY
jrH3QcxYHpAo3ToLc+Gkr5Pg4CRkZS1uC6FAyAhygrG/LhLxeHOly/FGs5SpFnTaxjHaCZx8U+6D
2wza8Iv7owS0UqQgu67lUKTjVD6QLbyXKLQAFfcYPWAtAE5Qij37/ggPk2jS6lNTGO3yJKlZznCZ
gx3P4qisl5lN1IpnF/Bw4/3QHPN4TjJfM4om9d55mdKgW3UBrUFFitPvRPpJN/5+pTXI/dD9Qi55
igyhjsZ7GJVTwkLC02OaSv7M0lLi3QkVl4+Dx0Bz5p1YAJ1pgtVqAPvZoFzn0pHIG7nvKn+k8zWb
nkSQw7MFvm6WRTYlq92O40LXDxgZhGNV3YJUhbZEaf2MfK/ZLddImAEvIZOgx/AYDj4XS8qaU4ho
NHX+Qi6iAx/FHKVFDNduO0By+C6+luY8aDsihT9Pde9V+KWPd1B4fG7IHWdPN2QdXbW2EtfZE6fw
5uuJorkHq5wAFnyNKjxqhY4ireE17jm5p95QWpNUm8m3PWZsNWA8vgGhtp9spRa5su4222aGfb5k
yNNFc7jz+p1vg26rYHPeOMrzq1u9+TDxG3qUm8t3kop3a4OdcxWXA/nY0m+Mtw7AhGSTDrgXusv+
yOD/zdYQ2z7jABp+G7d8fvOKwhgHGwPV6SXUWs7Lgx6XLx/3a4fF7Arz9dXgoF1tyEsyIQO1fuyZ
J4Mk+P5AAGfjBvPXg7BevHensB87ATiWkKdFqzinKvrUold0aSzlffyWcrRKrMSaItU1uLt9MvFu
pH3XSQ9esahc65zdv/97G5M13pWhAR+ieQS2YTjOb8LJ+P1oCVBAKtCBs0W2VchyZidokW5/tg7U
TOt6nUEtswLh8/Ohfs0+T2MQVNJOodaknnq9BuAmrAZFWDYJW8Xw1rOQ/OJseUkhzSWRJUxEYL+H
b7H0QQB+XSo7Z3doLytE86Af0dHibddwTiJTdR8x2NJ+Z5pGW+/PmHrJxnijGiiNmAh5thlGWWH4
8k4/8igoluyVD937j+YipfSWdS3zVzL00T1ZHWiWg2BG8DZOHLTMwSwFoUajf0DO/Hew/U1AuEdN
D3wK9Jr6GP8PhSdsnHje1LKO8+dZQBwVi5AHsA+K72k3aRf+ClRYspOTBdk078SlPrLP7gBA59sV
3UhmBUzCetKBRRC44p1bQhUEoeeDgXV5IlisgTFVmoDhq28bKhJukw1X5NKufAK8BAeMtJHrTmf6
BYceRXjLKz+wRgLGxC2gwqjvhTcgxuRT+EzO90IwMynUI1ivQivG3pKc5Tn3gUS8j6IHUcnfu0mt
gIW+Ui11qxgxrhaqGkIxo8WooKiBqGfXK6fEjpi0y/OsMrUm7Hj545dkFvpS/foZ9rngjcVNBpCf
c7sMYvly7MZz90S4K1uE0zY6TCjTtEhmtNKCTCViGRCQT2onEGDK7+IaAgKRzyfQtCrMQqXq5Blw
XD7YLl1zxMCd8DRK6fVYTmm+YkqOno7hpe8NfrJSj21DsdbKo69IqTBoUbQRFpqXlCRtEXgeRgTT
VcLjXlHIKwmjaxV65XMpCtel8Fp4tdOZ9NhnrRnob2aQ1lyec/xhwtdkYAD986OBLamuech5ACXy
V1ukC0avG6fAfq5maOBf2tGewqWTuhMfynPtBdYdmKa/db6OgbouGR4j/gkT6YBGjDTweqJCAUrK
WlqZBT7DYc34r4dkslSK4G1LiWw5VwwXSpk5H09Kkkt3n2aLXjj0a/QwShW/m7efd5cn/7HRFAHv
HHHbwgeV9gFb6Odfw3ANKsyi/ebDv15ZFLLEvBguAQz6d2x+MPUuDNRpupTc82mr4lB1+Neh2Y6e
7nPw5uDar+Ot2h0mT+qo5NNErG1yCLfsyaaCpdfO0DPThykonrqRVfEIi8PeX/ZAQ/PbpgSgdb05
k9Xi6CnQSkumhIZA8u/+DuLyWxnI02MZdTM9VDBrJQ+1vUpeM0C6yBmzdOFobIwD5QaNgkyzeJoT
UvBaO7vAmE4xWzXXUrMZYWeODaiT/TtaiqR1twx11rNaBlhBAOORgtnhLcmP0xxiv1w+xi0PGV7I
W4NuMUXYMlgjYbIP2E1GMX8k1P6goT6exj4g3KHcFbBOFDzBp8MMetZtG7bJBLJu5+uwhiiJbhKy
s5ZoUDTEI/+qlV7EHp88CgaJEMNj1onNpqtavp6wfx9hywG/yWyqRRaJoIe5c+1O9r0OUDV1B3h4
w9PWvRK29EHkESo5PbbLPA2nzh6v27Q/zl3lF4NHQA5Dymkh5bW8T3x4BvoU1nmh3Yb+uWfoAqnD
lDfFIOp5eXTnRX7mU4aZIAhCDRcGWre2P6vCIzNovpgDnR599NtLcRtiVdKmnJw2ioPC8rpH+Tuz
eb8A9pQkX4gvHzYb1wDo/gXzBF53eqv14MN4AAK8AJdsNtr0042mPRpmsACGzZH9SPsYGZEADxnD
vSOMOI+OH4mcT3aeaVkhGzeWyU6HBoEgb2CkW7+Ule0S/vT6sEWm1Nx4ehNtyDJSUgwywnHCuBh8
92FwVFCpqFGp5plwj96OFKzf/k9wBw2ZjD/JvEXnpPhfwB5OjR6YcoaF/1mHb0bNFK7qTjl45eZk
mwMyKmR5b812d7mKATg/0e58jtj/sElQ8JQzFiUqWUF3i78LdCCYNOnKrnKlN0mrMJNkY7FHqQ6g
yCj18I65ZS/cEqtYLW0HDsppvEVQ1UGMrSL4HexD/pu6MGcvbszj0xQlSPrzDcvlqyjEq0qoLEKT
Wqf6R11DxxgN4ihLSK0y138rmxEvbjLV/ThCwq8gFp/RGpoYDxKi7TPlisbPoPqLY97N7r/Sjjf3
rQ/JCErXP5ZlEn0axmiV8iA1FfAFBxoC6+z2Hn/xn6EkFT1YvtaJmlBKcVFweQ6tkoLI7G7cU83J
7WkJuTet/dpiIy5r5RsDPWIF3Vev9NfUseEyl7uuV+Lt037TtB5K3jJ62LVIJzlWrgIi0lEdzZkt
Ea4Z+LSGKRnk8GHHGCd1NqWeKkwqmQM3+SL7XvqUJw9ehRkiDpvAywTAvDuUmpO+NAlOGVieheKl
KaXESrhafcxadC25nW3ZaJv8565xXe6hlWOmO128LOYuIx6xAJ5cgJuDQZRNIHJIGBWnDA/sadTu
nzBGKAKpNEkAjD7SKss+mXOl49+/3JmamOvxF0DPiESpyxw5SWPQw75IoYbDuRWk/aFvyzX1dqdQ
jBntm7XmB4+/IEqAunSJT+wxbF4Fe5b1PTRxjHMT89LvgTtT3N6JF/WALy7xZ7WeW5oVeH46DUS/
E+IMaLEO1iQACG7r/orVsi1FOwX3mKVomg9Lj99c6igRXfKykohhilGLdIuBz1aTdxinVBGZyR0e
vbVDpnAy4zLEK5GAIGqtxuTEnMCpzUD3A4s3z0ED2xTZkLmJr9b0pznugphQFNp+7VKA05c/8Pr8
G4Zj7uMrnNt78WOM60JwCwBolQTTPs+V1DcZvss0IbQ2k0zkI53DR7E3un5Bg7saLpfhJU5h/Cq3
jJ57o8PLP12N9nE8waYhz3OQaWNhgggdttl9WgjTHEED1IXPTt/dte17Zjv8KXFhN6aAml1QZxKs
gYYrWyxv8dOYXoG48dNILcotvkOR7NXtfmOV/9Wc4igK/qmQ/r98gMLW+MsSnnER8Ai2g6bOgE+F
PL25HjfEgISc9ku+iTx5wNBzE804lCIMWX4iAigjNGMaRSxAV7cBcfn5Ludam8l8qqwJ8a75GcnF
I9N+Gc6lo8St2PVsWbRl9e6j8aJO7vvDlSOMw5qv1JNN1BHhbh1wWLTd2CshjkGzZjxHA+OtKmj4
JFzhW10YJUil5CU/c3GbOexCNmMkOm+T+Gyf6CNg+KsXqB4gSigmjI0tOwrykuY1XxUycQ4wSpD2
oPajatFBOJmRZXt7eTWWT03SNt4VN7QkOLWWwZqn8o0qLPupjQCF5uvR6+rGjC/q/0++vwyx8W5I
uVNb/jhafAkfpJdx8/n9qSAASCUxoiZPgIavdg7QjxDZPGTgVd40Hjs/4QypH+K2yaho4h2Ripdi
Xgs00eYM3QI3beu81RfGIvmxFgdN3NM+B2YZVxcO9K+6dJfo8qiqlSgdh5wOOQXrg4DLnhn/fkJq
v0iK4AShqpYNCGGplS+3T/C07akz0pnaN9WVkZMyl1vADHnotxKdGaq8dVQ5tupfCj9M1EOqhmY+
N2fs8r3CXOT26RIqKrxrQ3obGmUxd2XyQwjOtPMNot8ZKpAUpwxnka1RPUMF9Q2e4HwqLpyoAv+q
f5ip2DGMH5Y3rmWNLwafpuQNLpNmsF9EHzUYghAXEEmcqZaPtbCDlYGJ+cMUtFRwBykytevYYYYu
nceiRsUQ/eJh4bNluGU8wmC/KSJv1qLv90Zrh7VmanlOqTANiseZQEOtsN5fMb1KAWkOxBjRxhBU
DBjr+Hse5JgtS+rL8zWKdUhh1qLk8FYUiAHZQFd5KOylzm3IyOUQo0cu87IVowtJR86CUn4Dwh0C
nElnptnNkxDQNJdGZ9qZj/HdKv41FhdRUWxu8/AWGR+WoYPoMQPMDv/H30NKBtJ5ca2GZT8xhyW/
Vv7WNgG7qGcfDMKwyP5VN5/9wT/8UR2d5XijALsUE1dKwmf/TD6kHLuOSA820sdE1VkWixL6gGHJ
0G88LxbUha7auz3a/3YdjN8dj3Mxkibt5zOpaZYwl7RQenP71X/MSvTKeGramgVIYs2k3YXNGWEP
CvOKv9UGUnIzxQFskP+9IxP+mmsO0cirJuGR1jf5jLfJTcwS9AZzeaas6Zr5erprMQB8lapWx37S
olR3zS6036Wvd4yNiL2uclkkG14B9IqXHxRpiKgWIcW78O6hlzWHm1RyvTh1zNZ6BqoHDy6b2/xz
qTzlkoytGxMKXrqegQ00kRV2K3ZriUQMtxBmBFjBfxgDfIp6y7gyu3YRkpQpag6HwxgIFooRJd5q
o4qsxtAGSl8NIFluUcgikAoQy2o/51Q0JHZtyXXzFEH9l0LXL4R58DQpjdxBn8umEEGqPSsMnKGg
j9IUnpBYzEkpplfBUEKP4zdG2dTxbX05S6Bv9kpd0iueIjercYpN6tVAeHbnqJTH5eXCSXMvPfFO
LYDmD6+a1d+eR0RYNL8YxzK4bv5ioWE4wLgit9fMtLlg/MVtn8EwazDUv7VumfxCllk+d7kCtuvN
+UmfVpwrl70HzP4s/iJxzQMAM7O7VQsixJyicHlc0vcbTultFE6ZtSEtCRc70+x4xX8XW20TDLlx
xzMWqXIgyVADnk+kfL9PRJ7DkI13TtvFibCNF2XLwAt+rxO20Y1M/U6Sq47dspQCx9OIr/eXLwR/
z3kp6glLSCcH7cyVXEfpDtn0XqZMneCqo2svQZY+1B4F1slic7C+O65NeUQhrKMnVu0DqrErHgEL
w25MqFaGBvErKhHMXPg+h+i4QLaQAoaUlJw7pQXIosbl0l78gwUx6FMXVkJBhvkuV3XYCc7X9Fwb
mNUd88gR91r584NXPEjlEry12XfkC3PP7FsBiScyjsNgHL+21A26Txf24U/TlvBTNb6+wqYBu7xR
amnfh0nUoMbszulDWSzsjiG3Pv9+v/YgZLgu4fZ/ALMXRB9W0VRDmwlysG/y0cL+Gi0ntLtTe+aR
sirEWOHi97w49OEQWzp0fJcwTbEv8ptBJOwzKPJS4CrHYqgMms+VIM+/55p4BqDjZX7waCV6kP0c
BMyW2Xz5L/8rvagb26EO0+te/9RQ4qxdcOlVN5g+71PQuKB7scaH26tymWHPLR19Ns8n9t0Qrht8
sQEyZy1sW6HZUpPdxF4gOtRG5r48Q9nE4Y5KB+RwUFoz1+daPFAI2UyUDijE6JOhOVDKtdazE92i
sA5mityYv5Oc8U5ozTrilR85x802NHYayfsZN92s4vZujuqvfMj1wi2zT7JUsuJpW5ESQtuTENVr
LujEiJse2x6j9u7A9bvpJ7sPl6+McDtOD9VBcsoDS5Jc1lAxrknoVXTxezc6k1+2Mtt0SqD4f71P
CCP9Hy1j7m0psnIJc10AGAppfgh+Y9WAfewo9tHEjwoB2ebuepMfD1uTikcTg65XGf/U79VRY9EQ
//cCUXx2DWPiRbMScxTRV+S6g8mnkehzuxVeXIm/GmG0F4teVK4AKzBDvLlNzDlx0uMMkC3L8pXS
nYIGAru+WdtcjdCz0r/x+0OcHc5Pz3EgXi7IhAYeRaLMFWG8ZLRjZ2CYowLop3W273IKtj9KteQQ
wO5/eJiuemErAIGtSjeRJXWRbEbo4H18EYr9x29O0zcXFfaxBtFmjFhXVKq38v0rh9ymliYumxwm
JaZRZtO3PNdqVV+C4hypvFJ0edp7vYSJmftx6r3SycFyg1NXdUtBc8U3oymyOsbKCJptiAXDSQYU
KQb1RdgVY9Ba9zZx7VXWroW/ZS0u3q7TzJ/YMiJysgYN9WCwHGV668O80QT8vr8SRZkD6xKRT1Cn
WPKzB0dvZAQvSkRh/oDF6tHAMlBnrHUTbQM1pWUP84vmHzP+9LWv621xBMsdH6ufPIRzwTmPGyr0
RJCG6RscYkpEquNCLvRkITJi0EGHS7kS2PDuVQ/NzvMjcpC/es9R5vxC+tAjwY3eqw1u/WXD7giB
N+jvNHYZO5SD8HceViHStdFBIaoN+dbzcvoqJLk+YSWp2xS23R8S2H4eaml74vf/GvDKj2GJDApP
qtCRSN24poQ5WCJRN8DZkg4COj66b3tToYBMO2b8BRft7Glglgr2PLuiqWTqIVjL+mR/+zqUwcx9
JFwjYDFlrdfcLsQF/eP/j/M/+f6MGH6mf4hbi3g/6auR0WGYYtbnJuOTF6wHeEDDTwOgXoNPkie1
jcfF01qnroP+j/lDyYeC02Fhf78RyOFmFm6dX8dQlpcpDHih59KP3GW5rlc1zaSoZ0VTmMzFrZC8
R7VP9d21A/18B25sytQkpeukkSIimkmGyD+95y5Q1bSgojzqdjX8IteW9RaCyy5qlbKRsSzS6g/5
iGveiRVpiBlVW7fwJxJN/MTzQ2Dko4aLgzLPVTwb4PfVKnfnKNocp+CCaLS74bf6z22Mod2yS87O
aeYXjAbsTHiDyJSiYx9EUMSAFoCx78SAFkdu315uhAhyTLhHCU/XCnCJz6zgrViKKhmSUrJDK6+b
ak8uXCKeLEohmfW8Whh8UJPTLtxr43jAceICdlJDkYFZoFBl986dk1lpFdBhHNxYVlbjBp8fi3JE
sLrOhdOebA7Ck7ZpHF9/87B8mcTtHfRi13cdT52H76/wVo/gHBPgZuMBAQnSXl1DiSgJfVt6TCEu
Ct3tETHvpVF0lTRWBWjwE1Ok3DD4UFGQxrbOdPiE4SyXkkZKHBPJi97Qew2hXad7D0oX2p6NU8rb
yWzgWT0ygSTmmfl3bDviyLrjKZqAPQEyHjyaSw7oBSKRPV473ke5HNHxpclnXgrN56H8ALQ/4RrS
XSeGev1wQ/+76p2zmARHOrQo48sXBkGx+8hRt2BNAuFjFYSjPDpT/9+eMy9y8Q6qPewLWN1GsqPt
eJTnCSX1gEGQHp49ZMvfYYhJVY1js7dkHex0sjUcqJXpD894iJxIztMz74REjEXFyhpNaMpbg2dg
dJssRQAT/0Hh8Aj70fvxZ+QuYGDASu9T+gza8zxMlsQ23pV7YY0uslLgrC9qKmIaL4/9CQIJ0ASI
P6uWlUG50TFK/Dbfj59jZlbEmQA85cXA0NMhB9viR4rDV9czIyiB9Ad405hAs8H9oxSiycjc5nm1
knKFu50HPSCWJNRIef70m+857LRJIczR8lYuT3sY4I26HO1M3TU2uM73mZrSSR9NWyW5JbfxwB0r
MlR+qI4BIWjKVniYev/Q1JhKizWJXeh/6v5m2wIgbOqw+N/lAfoc+6xIBbpx92tXbxG92w3zQaks
gQbJd80hrmCwvUK40U3sdAgd4UQtU2qIRxGjWtriIrmoxpPgSai5rFlVVRMdCnl//5lRw+Y9NAGQ
PtfOgIisIr/WremC/HfYxDLvxOuxMj7o+QnzvJ5KaxNNZwDV6Ni+CE83N1FVBogUr73X+B31T3fq
7IIJZxq8JnMVe/RFXVB6/JF01AqDK+uTZzawQK6yiKOBJsiUpKfBPpKzTGI3wzIjJ8zM3bGsB7NR
67MUKP2mRsFRFaA70gqYwkR0fmJQvJYq9mkXi5ASaAwNwgQpv3lxepiBRSGXX31OtwF+JUlwWddL
q7sQ9mSvD6xCyLYj1yaPQgS1gvUMXZpKnGhsKkxq2IJrnFOvTW2IHpU3eqxRWv+v7g3OdVzHho0b
0+Jtw9GIAx1rji3kHbHxxZmqgtR4hTcNhDDVTO+hW/1ARjYeziMswIcLHcVF2Cy75LNoVcRYpe0x
A2aaH8JdcS7/2TLQidETm/q8VvI+7Vb3CcGQraaSY5Peol1afSbR0U3NQsfL9w92Vnw6q7JSEOdH
icBfsSXp2zPlEQrq8TajkUNni9DxVy3x2KTvT2pIXf/p6qN9KAl8bUATf5le8J1PJzqa28wA+YvP
wLrpCFxqYzzIfTtMbulpT11uEdmwsCeI5j9YABc6EA+T2qXE5stbSAFS4S63R64ySHyP+uFtLF/j
JgbprvYRjcIPlmQsEFDGYc9/mklEo/2hWk4nZEGqqvsJufX7UfgydKv7Qp2jcqQPbs4nIoiewPv5
gS6clkOkw4pv4a4clYN9SM/jpMiXEUq0XnqROfAPiibaR6COXOhjxge8I/cLqit8tmKbJk6hzw19
POJIiNyQOjy2ew2UlkcifvTV1a7hUdT9SOvyui51MzqxhB+UZqGiOXWes1qqlXd6vVivXfSOfYSQ
0OC9OLw57OrpXIgFdxBVLOarrgEEXBpR6CE3MSFN0aaB5n2zyCRKyf1PWxH2Y2g5EVeJyS7vVcqV
aChpnZ1urcpBhgiLnX9KHc6A4VLviL/ULG7CMt+JvkzIJv9z4xy1R5vbza3dLpGgQyK2fpWv6FVO
cOtrO3KRBgX+om/tOpqfLpIJY5z4MfOX5AERtLDiOhKNJgA2oUq7h/f4jfF7mGaudGhVMwQGLkqN
6SxqJIsEM3PIEH4Cm5a9oBT1b1vPTAjcU/belXsheNK7kt2Waih9lsCNGj+3o2V8uoSrTgBWraj0
bb7+Yh+n48f90rPDXlcI2ZBfsujzQ7svEnMXupcKTOg4OWn/nQ9lZEXPpdgVlXBhimZvfnqhbGwb
mJQw1ZWsaTF8ScbD0/CFzouMx6x3PhWZao6kH7q5Eskn8X2VwxbuKGUy7crazi4UVku3E0mPQgOI
E7q7QBmjxJNAoVHjcX/SyzqciiTZo2e0VMW3SX76m5W9SA1GMUwWrwpmdzh2mqqHHxKtv5nH0ZSx
6unybQbuv40/pSVyjsv5bhAUl46rfMn0a5X5YySgzsTQn965ofOEFsucXMnP9qE2J53ebH0ORkf/
sxDlPmIfggGzTIb6eV0A0CcgNyPcoDaYCJoADSa/dP9P5hBC3WZNWe8sD0DESRfgVFusSLGcX3DY
gU1xPyrJIRB8jHWaoRvWgb/vTfljMyANSGI9mAPQDYmJelsbXlXG05Go1+VXo2RuYVHlpZcFoPLz
xI5PEn/rLgVKjNsKBhYcpPmrTEbviTmfU0urUrfuqsaM8Ne2cSLr8gzYyLVp7uOBgnKoqteeHjQh
RhIRg5xWjmLj8D913USJGNsvW/ELvQUuTUHxuqRz9+iOIUSDg4XkpNTBPEaHrSMeHMM1DnS1KS1u
FXZnYvai21upg4veY1RP99HLnDLl1FhJuxKxO7t+BfrMsfu7I/ZMZ/geTqYfoUvUQ+EfjBo6DU2V
n7l9ilTGjaByNAnylTGhh8qXwP92EINhAUKLp1Lg8Jj706Y2GU9SjZu7OtqdyspLEjMkJQ7N4vsL
NAGcerCAFRZx0+ayiuCC578pkTZHRsCJsOJmlrhrG8qFImDRyxsGAL65IENc18WLhbVjMEc+V5mZ
uUKxbZwLAezKqP+QXdIEQ26vVQElQHt8q58K3kXjy3t7oSH2ijQUWW2F501zALwh+IxuQlWQbGzd
zCSMejp0WLOWkugrOr1EMTia3ddi++6sRttgp871Oq02sC/kuZxWUUvBHr+9IwcH/PitSuuYNAfu
3BO6wDaBpEJ8KHySTc9ZGBG9KxuAUBib1TpcELZm4m4TM0dGtL+wdsrXObN2ZFw8FrgJdVr5va7I
wwDjq3NAExsVve4qpQDz397GMcn7iHhDDZZziyPFC1Bllm70jA8r4Z4W+dtEYh0c15KopSnFKRiR
sum0gE/QwWfa6fdtwSNzswB0E7sKDykGDCF4jOeHv56iAryuE0v1MdUmgdLOnt1PBTD2vJTeE1mi
EmvMg4y/NCaxG2NOuBp7c59jFEse5yNN5ZWBLs0RGNZHKuKXHOu1Zu37Ll06Tzr9TwWCSKrNZ73K
idQCJzw881IN+5d98GGPYDepV9dMLzuENcP+I4hwnXbcXEEZs3iDqc6Qq0AHMkTiO/bw7hjMY9r6
0LEKrVODdh/LgXW/7H5NJM7HsqbFLlCQFxvbd86pguXytf30BrIn0ctFKKJKzvAeSA6AiRHwZgkf
qAsDES6BzeHaDPvPRYwXK1anMDvOnJrrpmcFcssDUsxntoJr2IkOBTJODPr8UwQ+iflLpu6fpKbZ
tuDyfWFxsrN3WTjyErVmogilJk5bQBakeLYKK8G9ktCdfYCZkfQoewj8i84obxppCs3J03z7PNkM
yvwZQ9CbiLOX6KUqO0TXPvfAjqbwGZAMC9bjUljTVsn3jcuLzqnZ4SlnfCYRekQ+v2Hs2T2cADqZ
mMwMDkK/h1C6zBsOMaQlRVzlrb0T3Ydvk+knNmHnawfQZzh7ikMmrsp3x0Q5NjHIGnjkZyuYKUIU
S4uYzP6wAF53xkiNEB9bzEVCS4sG1qnw751LubDgOsZSZtqEXoidTyDe/aSLSk7aALVQ/o6CNUm6
aOylv4zHHw16B2gGqsRlE+EaTrGUZxqDc2X6PmM2JDeSYCGf6auojcq2CPPR+6VAXSmXgnp4K8ml
3LPLBYiR162S0imB5yXCcPT6hQk9wm2GDcLe+gzTo4Nq58ZBuJUVa3gIGcy5WfN9ux9W0KyhlWKG
g35IyVsE6VE+djNNNj9BePDdJ5dEbmZ12D9iPuDFFiHAB2YDmHwUgKbg17g1RY7D36C0YTIQBB+6
/CiWSlZoaAdTzNOT9oBSE78SSfKqZpFpuHHy+fGizVzc13gKZDZdylu5MtgIRz+5yvLqjzmipArU
dKcFSHfX6OgfptyD9dq/4eDuyQscshk2zVL/AaHkxm6GC47qJABy0ulZu1IG857xhnqJltUujdDn
UNLRvN9kjsRWIKgmwRdKALK8QN22fhB8WBodzmbdDi+VGBHqfOOAe3+GHv0Jv7eiS7QU3cs5+lGs
lZt8LkK9ybUNsWPZ+2hTsiSLugRPTfs+PoRYeE8z5p+AbmK221/c9QWKZ54fVyDnWFVQWBTACDvC
GThgHWyA5xruYstS8bRJc7D+m6/BiZTOJe8VOko1xY0Vc5XMETIxkzrGbqgp8FAXMq4Do0xB05Iu
l7y3becCfBiPhUeDKo2K/HO1LVzulZqRko6A3Ged1j5Ak5147R0TtkiDUg3i2RDYklXFly4b/EFc
IIATk0bNGQhCRrOsBSZqIFNSquz42S+YjgXIjKEiIMt577k+Q/toCAXCXbRzydlysDAQxdwXJobE
yKg9OZQIw5QdL1Cl2uneXoCUP4kRmDx4D4Uo+Mf9rjuffxTGw1qk589UBZiHWTwLSILAjBLuXKyT
EbJBG+hmpIEzcvlXr906lhzDTtAPcCgXzV/cOh0g0UPTXgmIfrlpDxKn3qKRAA0EOItR5q4x3opD
rUijJP8avXM+r3cGNK2GSSkzWOdlL2U3jrj1trMM9jlnZRLRxdTSr32WhEz2h4+gCh4v9RHgS0RE
5szShJLda/gHILVP55M0jkC5+t/kPe8Y0YmdO3T4G5B+S8NJUY1n9WQTAg5gq4EEAci/shzzIqEg
M5HgGBFhpbFV4D3Ov+0RlrIx0p8N1Y89JaYZQ/HuL5KgXmCuRVQqd4BRMKpHiGi9ElW0aPvoJzV5
ES9z21H3tt+8pnftBfoc3W2YeYx1G4gkSpO9lEic/ozftLvudndqqU3ooxbi2iKEdXaBbyROp5IW
lcFSNnRAY7MFtgyUQxDIs5/cFYnqhGkHDotJws4zTMkGQn2oXOjJyDTHTxmYHINi66Xh29C4AFA2
ZbysYs9t1a9w4Ee52eg62m98ndrEhlIfC0BGxJ045iIm9d95vdjAeY28JDd4Zpakju3fvjf82bg9
wZ4Gpz3Z31S4F2TBHTqw+SrPK6EkBdeh1Zbpvkxq+BAVenOrMbizqqVpXKC1kw+tLU8q0bn1XS+u
Yuq9QCEIVMilDyhG54zhoi2JvIT5ZMmDtGAScXTzgRp90e71+nYRvug5AO3pMMUhucb2YPTvwMJV
+YKbdW43uLgyTCf4FKpeC1WSfohnzlJXrCPMwBvIth6Lo4E3Li3mlVk96ndSX4eHCBWRw2ANJOqS
fmS2Z9LzSzSWQQs/+YRyF8gSyaD9T7QLrsusrKGEuk9PxeZBqgJoXecAzVum3B+8wOyB7HwIU1XA
PmzTTuq/oJc3SX+XKCA1wMa/qD67rAd6iIkGCxu7kWgsayikOHsVxF3f2MSC3i3TjEqHr2LumCLk
HppnTh3EJ9j1/0Zifion1zhNRVS9fRBJhrbo5RqOofZxO+CWHO2AyrfWLXmoJEg1qqOwHVvbdSDE
nM3G0zpVE6JImMoTYOIPih6F3qLPEpElI/LPn7wL9UfyckvG78p1qMFJBR7b6VKjD+qDolnvEo4A
uCSoI9Hpp0yVBlW5BHSNmBwyvu46SwbriDw6ss2KYwXEZidzVJURRgslrQB9dPzycqiA1lgP61zf
x6y2QtA2+kdSts74jEXwPJFoBUNFrbr4EazbUxkGc/TRPX8jgyzDuOHKEdjm/36niZqapxy6yLxp
zTQ324pQyIQKGIXA23qa7Uoni+gecdbpDFSj3IEUjKJBGBBOepRBrZjjUukJASP7kbazlgA4O1J4
KZI77vLtRBFuWe5Bsh/3W6UOt0pgVzmWCAAbNVLIWEQze0jiKxOGySKX8RK+TnznP20fqd/9A5DN
4ORgB5cwyi71ViDYcOT3tzkJ7Zazn5k2fb7Mz6/Wo9Tg8UOBhhIwvHem6wKtYr2TCnSCapW24zpL
jZNvF/gFt0ZXu7T0XwuyvH1oacIM5IQsZUvKi4apaaZwLcdEHHkvsesAl7i4UHfQ9Wj8BzSsJCS+
GY3MqHMsEqCtwo6wsHOfRjBAr4EKWeKN8hDRGX8nPzL5Q4oFM3SHnFszBwjt7b5Afp6xOugwVXuJ
FuaYRF7VGl0u51JvkOjIPDzGuI0LyYnhnq6GZQduGU3JstkzIEmyaQx7GglwhRQJpa8RtLYlWO62
26IO3/XLfzGnhLO5szygB6Gv3mBNZTdI34k/j/Rdj74H2/36E1h2lc+7TEQHz03iub9jqOf6q5aj
ABrttT9bXfTMwPQ6tKQEyC9P4Kuh1a83WTs9AUrb1X6s+3xO0JIRn3qQOcDy60xjyd+C93fH2YRC
xNOB7znI6v07ue306V5ThlGmGJycSR7Q3NHFOuExTi0vURweeM/MPhDDSL9FT3nit+n46liaJ8uN
B+jbjH0IE1F8vDHEv1dLEmST9mnjlIJExVDb6mG6L68bnLXoWXI/vhfDQwV4b0EMcxzOV9F2MMB7
s2zupF5dd5a0QbBvDGfVhntUrqDlWdloL9XREA5kNuDlgyVfBlGI8dDMfxDBlX6mLLpcpis18cww
jqh/a1ry4mTrYajObtn+QzmP/DGKbrh+OQfXnpRUmL0khWCaX2ZKs0sdMjPid/nvrga9Nq09jaLp
+ceKJTEk6K21y3imMOSW5BaCZKMtTcWKIhWAK5+8LdUeox7NwbWSWf3hXLjXx0V7fTrTIhfenYdN
pz6vkDIfU7V56rW2lC1jkWl7TCWM/OuBMkMZa1ruPVk+YwiMosfJ7S4sDe99yqVqV/JMVtgFQlM6
vk8PKbvU1dcweKFm3p57adVdPhqQ2Y01iDVk5+5CGHCYqrs7X6qGy/QFjT43svi3qfEB5r+Q6Lfj
yMLn6RREmsrf7leZh7pwPIn7+/Ovcr1aN+N9TEo64VRiZfzp50ybTxvPcD41zx2tSmNutwiSF8Xr
a0rBEzyF/gjKTNJALfDGDcXzvO7fRG2+MDZKE8xkufPMpeMpzMwgVC3ZMAhtJRxKHfubcMf6W+En
MVvFRbNP1rb7NoVzlJ7B4LakIHfAOS1RznJ2pks/EfcvP9w0t3j80GzS/7MrSN0UMq8n2U5QMpqD
9c6grSbAQt3/M9k/yAKlXushjS0skNQbxe4V2GE6ph1SmlGhYfKKqdaXQAclYFl+oTIFiy9XcRtF
ewgWTuIVuiUCYVtW+DNCCfC+SgLI5T9oeuGirDdg/5MXRFYa0wrNCvjOTD5oRoZrMHa1Qd0wJOZD
EzlF1ZqBiBUQOGFawLUrJ5CoPHyWu+tIBTRQ0HGf5XIw6Yz8wn5UjS1Dvu7j20zJzq6QKSXsZcRP
WCEwnM2ATh4sOJT8s4rQjHxgNIrf7bKYQwuBPStXf9RXMVTW7wR9qqpW2pfxlx94rl+ob+EUbgm0
PFPYoeeulgLoIqmfnjOl7PCEIba3PDSoMR2AYiimhVgj4Wy881HqhDZyGE4QSqxw/nIJb2ySEwGR
AWhDQLsVcqWNTOkHuCHggpUxVjUPzhTRt5TTMRAd4ailU3aKnHjgliRQAh6P1h6+4XPZnrhqCqpM
1SqZ3AV7YlrNBr3USIev1KtZXRNNWAn5Grga2/hXBtiFSD7fYMOlv5taUeEyZ6TxYyPVkmMglXfM
WwVkXLnj+Vu0R6YLkMsXYuxlB+sA253zx9jnCupy19BmKLne6AdRw4p8rX3SbGcWxzMVK0nzWw9E
drTf54IgIOTrPuup4CB693BuQmVrKGirEHDTEchYJQVNvLBDHoGbBT4hkH4UGLM7r+kDy9tHYqn1
qO5QtzzbHMpyJC/nxdEF+NM5jS3Zf8n4jBX3n9OBTEyw9dGEza4toEBHLSBJTxZlqqvEHc+vac8Q
RGeZzm3Idr+AI2zFSdac927gEvQPMIK+sxD7ywj5D8vMACNx9a3Whd3RX2M8aTkgLJGFy9FZoSge
SjpGVtTpDkkgLdEsquRD1/GhlOSfvvX6iGcfQBvLHLn8pt3xE5EhqjRI62ALWxgpAlYpo0N+/EN7
eBhZ6oxfhQ02JDGFckiFeiLOgGSPeMxuZzmyls1XzJovcGW3bIsdGpDXAMQ2f/Wx6X9A+2eEFOan
jUxCCXRNTAzlHCEFbNxwXUI9xucH0vkj1njqYVoullIVmEsS5YQSdld63MHYgyBGCf0g8eUwKoRO
b8nd55odMLCsxCCcl1AUGSMgDhtoSM/owa41zqB1/5vlaPyxF9bzlA94Nw+rFP0GlKyxPkqkwQig
4GuiCfvnh6wcBYBHa8zHDKarddMCXSXiWwS1HTfoZ2nYFXGbPuFUucebjCPAxeH0eaYkFD/PxcTJ
Fu05G+KVwf1syZ4cF4UTM8DVpwrwCZplflLvpnk1XAHWNMWCm/+F5kR1VheNRg8n45jS5Ml3c32a
IwykEkpe4jCOnKqw9KNQf3LqdLyJQMP00Vh9RoOu8v4DVKazaInEhkgi2A08amYkZS+wSnrERIAe
cxX/GZrFMzunPVWN2E5DSP6mNdmH/HRnFoFZUxM51XPAsilkfwVylq4WnxIfXytnvT4K1B0AC54N
ojFxVEokOC53LXP1TXVvH4KITcnIZxHJn9PyBriLF4NpnN5okm4+IXF/+KJCv/ApsaWoxXW95skg
yY1XCR05hQwl2VSmwil54gVWvP8ChJm18kAHOB6AtFpoja2XGBhm5aI7wxlUjr3kWVTlrBFeD8Na
qC5/phyz0yqC0fhafYq9VpOQYSpeeCsyHJU8D3KvKSmqWrKz4oUv/t3ZiKKkbg85QGhlIgqKqGni
HSUODGdg4+nbVLx/mnECXiNGkwgdDo3nlT/gx1ppjwcVA7NGNf1EKXOknsvg48mzUbx1UCWRClHa
fSXA4ltMmS7I1XcHXXO4dmaA0APNbcgjWon0cSoRFXZAS84fblodDGbsd/srgeBKTFiZMqS4DQkr
ncBoAtFsETkfk+8TuO80GWIGd4zSwOjGHM4bs9Z+2nNNS16JiKWZIXcaAJWv+I6PyzGI0QMcEU1g
ajNFR4M3u4i7cuw0WrA8Kdvr5AY+i88kLdG/rffwTcp7IxM08CmYLC7pLH05n2ueQj8j9bAU5emR
0cBmQqYAt964LhwlH0TFmqx+zyLc1fIR0VFkjvBQGFrpIaEh8d/TKSFxN+IVE/yjhuInH9/wv390
/E6EreUjDZCIGPCiKTDPWYyYbss1HzEzLWure0PsHi19sbGG8o4TSOHJEQhLPaoPr9kYOfraIuXl
mvWJp39XK7DouGcu7FY6xGxXT7cUbWEAp76z8MdsT+ln4C5TqRijExqsFkBPSdGx2FbzVul+qnOl
zHU9wKAYAx+Yz3tWwGx9R7gs1iBhsZVQx5McJxt2QTqTw4Bm+19Ymvu/ojJpD7YiPI+bN/QylOyJ
N4QcAm6sRL9kwKIwH1uUIDEOG4oXgfUdWD87kvBqAtv5Vc88jiIeb7fYqKICPwceihKPTN8IOTpF
gT8oWhYWgo+cO66ny6Es3Z3tIzD9Vq4Mrl6QaIoAWHZXE8+Kblm+YK9jUcljaM0hVysaqBPEkOMO
VjYo7BFvLwO1jGMnPfourgEwuJAZPDTu2RWEq1gw1Ud9JqNHJ5krW7ej3sh8aamIpz8wWz0Lj8DN
RYhizKFNRX60KtbTcwa+90S9Qh6hY9GnzgL9jC7I6LPlVMKhJU3+ISyhRndZMH3+FKKhmFP7djdW
2iHHMMOJ13NWctwaUmX4v+Qx6m4/318Lxc7M07GswOTUAhdGDssg+qMwHywDVKsRhyQ5kA87lBJQ
Jt+n8VZV9Pp4fNneakmY/MNLb7BAQ2WXACikZTefaDKEviwq5JBQMHZHQcb80lsMtEHeaeg/W7nQ
Ds2YxoAch1cf0VCWjnbsc0LyDoAfMwBq0cykGcSWQwughJygU9UQT2/Z8lDKSTwiXjT5LC7bFVne
p55He+pvxXxeXytSduVhOnquOL1hb0tz0Xi8u3l4Pe8VPTV5QwHctpdYoEN93PNymP0GzWhsvwv9
ewJ4kYcNfqSolSk1PxpUhSMvTUliCrG54uXSEKZczgUTNXXawsAbGhsV1f13Gq1b10AG6+celY/9
9fnAHGTfQJs/oho85IdoSvAKVWUG/1AagJnpbSTMNA9fD5h8GTqhmYqiXkGf+RroH8yT5Q3lrgS+
ngMBKUTVpEgP1/f+00aOxTSxW9oc/IzB6el7x+fqbKxeAhQI5nn7Yrc/R+BSE2AwOQJVwwjJW7UL
AlDhEdXpm2ZqzqoZT4pN0ESq5o3JC7fGMPPGOXuYRZkIHt2o/IfqfKyPZiRCLxC458tnsvwBAyzC
VUBgRalA2LpWWjVZObVsHUUfhG0EwXxNK7vjMtkF02zt6YH7TF8TeXWXWxJ5YpQn4ZukThW2UUyF
R841sKkY01zctBkLSd4qZG2hLTUSw6We73LggjVcf58G4mSMKmj4M2/w0kwg2xGeGyK7utCfgJ2U
9pMJGOEWx5dOHXHW3FkmJP4WSMNL5o/y1KDUa9Vq3Ffb3bOxPc/d7ghPBHy7kHSn1JuqioKStKia
hkvRJqMzzKdAf+ApYa0MXaVIH5ItVg9olpLxH2SviuWT0B0EcdwW8Lqo5F3ITsOiWdWF/SSANd8R
YufSQu+X2h09/gQsddmnnTB8/lm2BJHrlG3gXVKrIdhldpgtl5B+Wi1JbKIhhx8M2J0siqC40/kc
0qcV1Im2r1uyIGRyeEaXZMpKzKRfE/KzoDnYdA8srOp+1Lzj9SWq3OnFBqggF3Ezy2QFLowIGi0J
Hvk0UxQID/jcQyedDF2Ae8fzn7wKhkBI5x08LamcgcLSjwWNmkD7Rcnll2x7WxtD/YvmA46ztOdA
NZyfwVp8boTiaTCKqFd2LEr7JrbTyyp9kIljtMwrcCMe3E6vTxMnnSYImhDZid9H2+0gXF4SRxXe
cvVKZlVgnDT9qWXcc5GpeUfE0ZPG2s0kipl8N616whxfzj/oNvwKu6aDxa5pFHSePOTpsS2n7mZ5
37SIW+8JaAHn3aVlvu/cGPwXWsaNYaKnB205CGwUv1SAgKW3ZJg8ZqNBQXBA7kq0siRP/P/ZPvEW
jDFon7jiF4Lhn6tu+fk3rrYqdj2jgXzaamItiRoofywzC51MUkuoeOIMChJi2dXlVtPmpyBq8GsT
cR6yU6G243XCGig3GNqlfO6I8H9fcrFbTvERzlvxbl3sA/mG8O4kSlyRYoeGzACqLRRNOAyDjI31
9Stpt6wfokqQ5XInkFqiuCcHoItJqsto1nF6UuLtkbhWAhseMsgBDn4psZmlceVf+NoovnocWPik
JSVR6t4YrffsJv7w9XBMo474IW1Gu3LLfPR1z8K7OSo3EWu1FBZuewsJw/c5hDOs00wSsRSjBgTT
/x7Nzk0oBe4MrTvjnQEEWy2MWUM9x2NRHgN8quzP8TGhz/RJXbn3vx49HX5lNAwzkIyDWHVHhvSz
HmEXuYEIElloJzR1afXeieC4OSmvuYdHvX48Wvy3TqU6WkXfFG/hRozwPq6+0zp0IJ5DUghJrODj
iPCmit3aYfR+Uu5wMIjCBgebD2ZPLmp6h5oW0bKBbe+XA5081S/6Yq3ZVuYNcbP3G5hAAZL2kVal
ngZv2G/tYuMiHmG9IkBWJrmueKW+XxDd7QSAzOeDrbSA222jf8Hh9YN+SCqCxmTdiYeYe5Dr8COl
FrK7KktT9YAlNSeJ12RrY7JbOzyQd9CH/4dqw+poRWip1hQY9xyvuov3zpSNiI+fnbHV3egEVLI3
jdwtR+BeszxsYeyBrY8dQwxrucWGDQ8SUxoyGiIxIH+qqsWhvH/0AW8Ge5OXBorm+2qkzq41MwM8
ddN0nzq7fMRi/bTVCsU8MRLGNB3JXguaJcUYiBCIfRJlXdBSYNC4iQIhg0GwtBpNM/NSEpm6xyMO
hf3J46o4PQrdSw+ZYo0xUJswdvxObZZG8Ufstw2Piy4UDpM4K56KQUtaADGLtauI4X91AQMBcjO2
ehtIS9uxZaYkCv3i52AXKm53Mj1NzT0ZbrQGRr+0j5tTacSjfzPM5vYPLSINtUGz9vvcUvrX2LGf
Y+rx0qHtgiyhN8J0WqWODSsvCePH+U2oU0/I0y3A674Ct255xX3nqvvsIdr9DcPuojhTHPQVj4ph
tBUegbloFL3yTrRED+67copTZoe+Tw5L0yUDaL7zyIMvgs8qv92dB+GHq/vS+SK4S8e4NNhY8ZUf
5UiiLIa1kIe1gyqiScY0MvgaElJIK7fU5uyD1IzIuVjEmAEDJn+8TDOWDmCyPncZL7MlJ0RtBqke
V4rGwyDjrvVjfRatlUfNkQQRMxa2RPAlfPq7uEhR4oOb1zLRJvMCTgSZ10rLx+FkyfZyvRYc9tHQ
vWwceTLrhdQOu2E1QpvwQLNmKmU4mShM8vpISSBaRqQb3kaRe4gPBe5gwDz2PfVFWnW88V7UrzaM
3yDAgXS0DQ7PVtw9UWL3SwMizS3HAwac5r2Jh0KI0Xy01DJrl0Ar5RG1N6e3lF5LUtf45TwgJLBA
W37+GpqIU0DPUHDxRVp8I0RmGYu7K8F+XIuDiy0n2djwDAWVM1unyGReUB+9X5vPNMyhS0nmS7QW
OBjqDbo66lWh5uEWMBJK9AqjIeI+bmNq0P4ysW9vY+fjO/enGoiigKLTJ1WWa8NL4+lE5Au4qSsR
9suZAN0RLaQzv29y/i9nl894H7auPx2msBNlpMLwNBsWfqpFVsJNd56IScJs214f10W8b63ZqjbY
ZSnawiDPPOFRAfsoPLSc7Xz/FZe2ICd04BEg4YzdtQUDpO0JjMLlmsPHwtd0unOzFi/CmJpZCnNr
GgVGjhTx5eiFz+SmnGaL83pFrfKG7HpmtKCQPctN0mrZKeoSbrsvxFe6C7IQJQ7DO7yIO5/ltA93
xCK17DbSHFe6482/pkpDTcG3abRcVi7gW4KHmOo9rGOy3pWR5Jfyyggy1r5sO4uLZ+9zedEFikwA
hQkC8UgjnBdpb23r4kiDmb54am4SpPDpZYhPdm5ACCtOxkj0is+e51SuKaiaFlB2RhDe5CPuC6TZ
znYTcJnlRm85i22YDW4AlK+Z/MFaPztHd8h4GwFPr1/E86gNtDFrcl7dwFhLc6fLoDpRAQakR81N
jyRyZk4VvLnpk/BawTT89DveZxHP2V2A+Lv7Nm0hpsPl4yLnunzjegVJ1jqofgqfNhr2aDhRE97b
6802eE9yvATfyI5eZb/8KLYeEnnLa60fBD94MRXoBKI3f84CX/fjospeMNfFyxOuL6ckPk+t3Qes
3i9sfo2e6jQ1Pw2XC4Bxp10PDo7qq1Z3yqhTRPehBbhCnC2j/27bDKctfkwsfsyN8EP/YYf3SKL+
pnBtY6rqXQPN5C32Xi2RFY+h59FcyWV4HZOpYENtEKIgEdyzSGFAX7VOSoQTe8qjDdpOtwZKJvcy
DZv/TwPYY4mppR7YFQWyS3ZTdLkkOpDz2PlaUxN7SMrYf91btn+FmFsb6DVvcJdbKLf2xN93s3Gj
p78gPAsgzzbyHtejRpTIwpBAUv3wzl5riqBoCtfpF7IX2yYu8mieSzJh9bKag+7mHJU/i+yRhN48
si1uEgiNz3ZoMRIQfuPHEU04KOxS4OBeGnbeb3e6/+RRu0avXF3LAGzcdqV0GYKjGxuR+aM6D+Df
eOlIlwQmuwJQYTJCH5wBJud689fzlYP+/KiUyZqS7KlnUGhdte9jMc2UXD9cMtsUiP0uEIT1Qthj
wFZ8IGNrmNfULMpmZV5HbYRANScrgH4ByaIq5bBMaA9sqT+nsY9HqT+ZbJpsCmR3sk9OYa/EbBlQ
Rl416JCqYXHFXtrw8+G1FEJkDThyS5zvaxsG8sDMU6V57p7LKsvVuzPZfjJXaKzfLQw+JbvLpX5X
lqkhQzpsjPI5smvghqXMeCCWXQxHJMURgoZ8E8xJGwxThIyiNOzHo/M6qZ+DjOTSDN5ZdmL+MSHA
bob8ms/uoq7PRRMR6tC7oCOuB+ZwKcI0ajnGT+G6RjzFUkTznytn374kQnJ8h5jbUupuVWunyDQd
Yat/M4Etbr2XaLU3aZhlM5psZ2FNraUgpdaPhDRe3aF3hyWbYo9JV7UDJU51XmoD6Y/XU44NtakO
TNDQ1qk4GKuqjAYnpQy7LNqDM+qFetTfiO3jtap5QMGKprJqpYeWfvyY9yPLnMFOK0TL71SIjddL
Sx1CVuvhJCJpR+9znMbhe3imZoMHWTggAFF6UA255mTpUPIGD/bAFFqaRDBvfGr/lz8dVwUeBZyg
ndYE0M6PCvB0CclGhb5+uJ5yezlWgXnjE5SXPpNCJaKHSltr56l2HEsuztGk6HwbF1NqqKV8XhDX
Jt/vrjhxOkb2S0qo9jaJng4l/xVIShe4AJyWv+aWp77OzCGFIpMqKvKi+ZHjECPoiMXSmoI31Moy
drOTBTbhD4ulPyjL5WQzY9iUlVpYE5ecIwXldQlSIbrGV6/p5KtIw7Z5apylV/kURQr00UmHO87C
RdW/KSJsGWoOocd5d4Ut73BUh6A7Ix1E+DOnWi1DHqED1AdA2BSBBzS5ZTfTr7Vjz8r0aP1Dx5P8
IYEKLu9fyNTLmPdYiL6X6I1aDuGIuvc+PRMRLeyhjMm9hWV0pAUcFQeAYsxbZ1UcLeV5fTHsGJeX
zagkRpDtuGQPiPYYiHh1ErdIp6fz7URCIJizWI97Fe/nkqTZf/qcPBOVDDTiTJhhs2e9o42Mq/Sv
uJcW5NUL74COAw+UnCLzliB1/jwUagtyIefATahcszzH1ok9IftFGB6yXNzqUaS7uYqyKQ2InKVZ
+3CXfT7sFYMt0PSWi00s0SGCgievwbg4nqpPcdkXoQAQb3k1J4q8gDMhH3+fxYEl2B9ooQ2b3iKw
XVbO45RDrNTt/cQnCWTCU0osUBl3wKOEMVMeuazAt4V6k2dGSVGnMhb9h/T/sF1zXDifKB4l81kT
B34Pnl3wSes2sQ0SeSBqRNFCT2BU4NxaPn1SCw/N6ds1LM4Wbh7s4tilzZxJAgZcgYBogAQi4qtd
lzFeq42yDpCwxL0ZOjGUY1d3DRaAW9FM9Rdx15Ut8Rj+MLVW2DrrJUrd4jM/D4eZUePC82TBLIzG
aHyH5bg3vwZaJDQxCgIvFx4if6yj1T1qZVP3h3HLarZvhge5GxEgeEKaxmM7d76FcY5hblrl1qtn
IGE7+IB+KoI7SNucO28ECzQUpPpJgQ/6wLQJBExKIO6OFIjkRAWeguLCwTbZkH5xKvzaca+eumsm
Rz5moIc3ha7FuDh4qO6egGr8D/av9/3RU6tJ/HCP0Kz39OYoW5GVUcVlMyjvoSbAx4+LeVOz2dJd
48VK3DWUMNrSIx0SaGZi3H46QhKT4EaJlEzXkTVkBd9HSn+81mYPiSZDA5qsunjiFOHkW1p+JJdq
yaVBWeoGjA984HKuEOU9cdmSbvavlaQm/mGGUh+B1/opE7CFbp3HLuUqxXE3tNJJXtgDGRzuCL9n
PMynv01RW5dYL/o9SRzkQrEi2fxzqGSDZaDHWrzj1Sn0plXXPpTAGbpU+LxHNkgxmJKU2AcNA4/L
sOFrWwFUMgII7K8XGzoVSDEjN1MwuA84t7FycJJKPbSuAGA2Ih03r5rR50OiG3Ye2lar7kmOxPAZ
w5lgNlCvxeAxHeN5YYQbg78zwyiavEHgRWBHoJieUCMd+yaPu8UlnKnCclLK//04GcVTZ+aAtynV
54IiDdV4pUuBXwslFdiLgCxEZsNqfl9rgkBw8oyNe5oGmWTWDwlYBnmwPl524HaFGEG9ZFByOirW
QGQ8DzNmNHwglucoa9X482tAOe5m1t1Atg1To4Gbn9ATbDNcy/R3nP7qLp9+DRcHy91Kp7iRYa7n
xA9UsPmuKdR5GyMLhe9pJIYtCDeC2qXfxQhnLQOYOfPJ+jvbZyLN0/mzc0u0SfBSlP4MW1Fl095e
y4BI7G4LiOj+hayjiMUUC+Y4h8cORh5mVs1FMd5wsKZsSc8PVBzrNBQo5xxVQOTfJjW6JVHan34t
c4AsQCFICIab836ZLADujFLkm+7j1y4yqoN5lNAxUh1TNK3tlT3ltcQ1khVZ5guQXQUc4VvcJNaJ
z+mfpyAsrdruJOp0fUNJ1OXMrwXvjzoWqJ36DxXHthHIKyu5g3EZRna0b+JxTAEWSosa1sW84yCF
9ZtgYs2hP3oNPUkc71uwC9ohlnW20rJCfjlYDRIun0SBqsjpq+XQs0InCAcajkhNZhwgPfp3pMhP
5djWz4mlojOUa2RG80mURQIKo8BoojNbSJJQpCmRMvOYKFSYvp7Bb3txaoeMyID6B4VR+N9BDzDK
o6H1xxW93J1pqXPGfJ5uK3bt6PrA6a8ZyQQaUaLq6eW6YCsUL75prSpSWgo3i1EXhDfJ2lG2994A
tUhiiMmApKo4lOlUQgqes8RCQ1XgEGA7jCiKwEDv5zT/Q5C/JA3OzrPJ+1Keh4895MFGQwjbdXES
EhpKdr6TnQ9KBSIfAiLVUrB7VMyeQvW9835wtRHcRUcDX5OAw1h+SwsQebri3emF9tH1ylHymRrt
M8OW4B4aE23i+CuJmbUMhXeDuZO5LOj3wKRZyPdRZxzEJGUzRjA/4L4yLBCogDgvJuSRGeOnt/UX
ICHqclUN29KoZ3lpChMOXfowSCKAN+abkHAq/Q99+3vvTXSVPQTJWHP2mXHh/4YDsXoionj1x+q7
2y4ukFkXqW2oaSSZ/dd32MtYKpc4qGiqeRi0v2ByI1yN4kzC4wOlBjOBL1oPHoeGmxa0IApVLCnh
EJ791RPC5Ggh66b79JbZEsJXUhijaK9cSvtdIVkEilym+iAM+EgT8KT+qqeLAiv+aZWt9yeQaUsR
nv78Y3wd3SN7Yih/eNAubG8M47h0aXAt+Qjsco2qhpv7STs7T8y2tItnPL6XI1a0UAJWeDQx1GN7
6wLqtq+U7GKcE4XaDch5ByzC//hkXUBLXsH0yKLWR51F1avIQN5forW5/gynx/bnycEVil2czo6I
Rof/WynzdiJX7cORfsvzaWhhBRPSSkKe2nprSYo3u0OeP2vMaWGdd5J4OTuX91YbX7zz4gQozHWo
4njEIwHqyWYeKjs802n+lm7OzT0nJMcGGXCMeXw1L3YdHK3zQSe9exZskoek6u8JoTLVeYVE4xnf
wgliQi+SNwfiZW//97hnfFhjPK8kiTZVALypVJxmxIpK9QpTsPqrKDbU61ac8tmEPUghfBA+V+qO
C83hT9q6OGV16LkYo1GLBWSh0wP5agLwtYx/IMaXCeWhC4uGE0vap80/6wdnE3WrF/9vCOju5U8j
HLfGyshYT4NqAuNUgGXBs5nOiI1fmBeDvzTsoQ1hw0VwGxQQM6VCwbNAcfkusmTFeoULKOc6y4hV
b4MAiJeS7NsYveshVo0NsPjQJAED+E6aKArgENW0l5APlPatnA3hSJU2FKK8CQ8dbHj+9n0OVw/7
o/9aVWnGl6ON0e9QUQdZ/uxwB+XHyrfwsXcM/lg2xujbzCvMez4sCRIonidANOZsTuyKo8hSjB2P
mL7VZ/GqeA0T9WU92Rj3TtdCIp4FJd2594uuPzouZRrrJXtIeKCjJkoJDp8tyhkGZevTnIZ9jr3Q
bPUfW5rEJXZtCxiyUYPb8HJOLlOJk4SQ2lPX6pZAK0JJx3lgFAco8KMvb99uSZeBJTixf95waXgu
RB5l+69WydiKj+FblJ/NinGPfar3NFmqfXZ6GdewC+aWs1Aow6OqfHES5bbxWK2NBRI+qByDKW+J
vqNPf+PtP9rgkptRb68d6qUKPqrMAerfQuk0fTKBigdYl7m03wCkZJBXj4JMbUqlTeKMm5D9Yw81
TdlJLvd6HgG39MxZZhD9uXioRIwgK+CTZKhurP9ACPYcVJeGZl4AtZOwEhc7MK8nLztQmIRRvxHq
s9GHuNK+CdSAkBbL2n2rsaYGxvYGIzQ33/Y4RCOOLl+Xv3F5bzzq8N7Xl1AEofxqfklcHdsZWwaQ
pxOtwX6AuNHf0hBkac//wGNb8SJjDLWw+hiLyCdJ8uz+NLYLOPOk8UIxvnuHL1gTqV63h2IL/2YA
NvKlZN+VSYcc9tovNbqSNK+ZzMv1Lf3u9mfMm0bVLMeMHvHTLpLWJT6UxRJjln/JXc9VBhIT0YKK
2ekKSg7Him3QyXikxQugIQRDjK6IZjliVXpl//QAlH5JFsMd0NiCLZ/ITIdQcZYi4M9jqWoNHs+l
hdeHCbxlRg/pRICPkJnder5DNvF8Qa6d9sIsJY6pl8TQdCXcNYeJeE5G/cDGLhCGQVhN28lORphi
UuFHKbPiD9ZoRmLGzD+HsUtyo67qHfJ8MqIZ5uQeT2wiUZVvYZt/oZ5s41fILuPEsq2d52R6mJ/y
p9hIKRsAIef9JaNeuUTW0slTflFvbMnTuD3PLkJWKsM+aauDaZsNzrFwkN5p76PGu1z6DhqsIHyj
H4f1CPQgn9MPkpvIpCyKq5btqjFX1jhfmgGxvMBWImgATcyWzSqvN3roGbLsrfmBAPgL4loTFOmz
rI4ek1c7NwCDr5QyScu9BUGoqpBiKIIA/thhEs/lpPzO8JQySnKa9YwGVgAYRLUMYZ3G+8CMa828
/9z8SLhgaxDrOR2+ggsZyJ+oqgZU57fz7rwRQgxi/KJyAdNtMmecD/1VyxWRCjycy8ViDuNsIHaa
nivj6whnL/vv+/QY2+SIeXIbMhknEGAhwoWCHDn0JKbg/DMNl6N0ifCBfBZEsLMYC/vwjo5gCXyP
mZHA2MbTuQsE97nK5MlBF7fQA2nEkwVg8ca/4TyZTDSBp3NYx6weOADBOQhHZexzgt6dmqBd5BLG
Lcvm0WdhYjTUv5OlbMdiwBGg4cNXVv1sE2kHfO7umb3NOFoeQ9tIfLmMSMjYmeEhFWTwed18b9FH
70tTZJTh+C7PvUOvA4FVGPKMeH86dZBIOP78ztQdfqTYqv7UlD2YDJ429GBtA196FjQ3bI+y9gMb
4h3HR1m7UHE0I5ukf3usff7RjdbWkToaJBT8z3BBUnRqlbNJmsRv4Um/YjWqUozVXZbHSLA8TCIB
66t6LK4J6nZ9QsUqGoQYAgeE4hwQhhiaKA10dqAPXkXMvWo5lnG2OfN31CRbAFo7mdjrQOfcfuS6
+1IH07VuUN0EJHlKFdSq56FQLsPZ7Ve+A3E8WdgxQJsZjr00QDIrtyhb8xdKVIsyEQfbNYO5GU5Z
wfxhUGB6eXQBo4oA7xWwEq/CqEt15suApkcnvJHfzyL3eMn9QLswabcBDS2cF6kx67x1LSFg7iU5
acsWjrPqZBUSUsm4JuUbCjErWZzOEtWyLwpwEDZ2zjyTHE8L+kGQPIq1N9nArHBuP0YIOo+gC+zO
IjOYA/ZreeJS+jSlXA3LVQCLTxbfOD1H1SzfHlymfAETBjtyij/wEUG5M6MBbpfH8jsBbrvNPqnU
8S9/ebjbziULFFL/wtkaW0absq5OkSjjx3Gqf2dmUZY0QV+7x6CBm9N71p2GdCVeu5umI+/kD1+h
kIcCq08piBNQyDyQfQnd/n3PQa2NunyHEbSPFAgl9ZtL2yaifRbBAc+Z/7n8nnFF59ANttbWTjt/
hWfmysUIDEP+MM9h0O0Um1OgbTI9g3v5M80oFe87CKETgaMUwQLKw5besRUbcyDWkjeQDA4yoWwe
7FOXM2Ol/XKi4j+noXNKDhU0bO+UUvd+yntM9ol+3o2hrRIOjgQvpqGf/qE7SCPJ39Y4SDh3RaRv
QnwyytEdYe0jqzoJAMIozzPY1nRfQB7AlZDjpxezkrnJBbTzhuFiBw/oGDbv/1o784+VWx5fMzO0
80HitqetGS23369kk4kB6dq1vE8bIb9MRAKcGUxKu9LgRez/zsX8lAUyvBB/MDNVka1nZz1c3NCx
uQZlBIi3tQUdfMORwdT4SrQicMSpsaFRD6YHBJ2TyB/5wTe1Dy0XUOkiCDWMVMO/HmLsAeTHfabx
OPwC+hfp9kP5UDNT8CUuvxRebBjJmJvBfqP+R7HFl1deOeZ3qV73MkrRgMU1buEi7k7ie0FlnNBw
eGbuWfh7QaKQOr1rOhKwrOmljzRlat5MFsyE9vjtlq/gmWlHoY/Cd/OnX4Gsj4iSZimze5DLsD/+
dKXxUYp1jCH+WM9oiOVZypsH8wIBIIRZIrsGtkj9nndgrPFrU9Eqz0KDchGKLiZJFknchUz3hPWc
2le9VFZwVlAuYNKYrSavmDLAdD702vuPv0eEV0USq+fdcvH3L3sVfeGcxNYTKu93uNLkRTlh2Akv
GEY3Ps1QK2jTKuKH269mK9u8s6cij4Unh1uNXV3citzbp7lFjn0ucIyhiG5CFu5LtwE5KgYl8ak5
VteL8v894NriKimrfhjyIEcjIEsZCRhOf2yeEuogEU0rEklgzN6/OzE68fE1m9z7umLstKojgR1T
VadXkMIZaZJuC0NZXY4675OjvOLpgv/gQeXO3MQn3hsqi13xJndUdKP6tWtesLODjIeuVCHw0SXo
1uYYqBWyh1+rETRypjWE6FErubAHhMhobhsXaeNMR6bUmQ23/xlM3HR8FH3LNzJZKDhI4kDV/VKq
cJmbP5yb5SV9mEqDLwLWudBxHsa3xPynHo+tiYS7anWK9mzxajXXnxjIFvnGqyUl4UwQ14wj9ODU
dHmQJ1objl/BWa9a0DMzSUq9unjgV1YyUKm2/CWtSmc8K5E7t3qwuBmqSIe3mzaG4TVqSZK2+Qwl
Te7x0SzwzUYntv3u5YTulkibWYxgkL/tQ9FeNNsojluxZCqKS0dWq8Y3ZrMVo39WHKTjJND6f42X
O6ORU5uSE//n5wGdHYBexxDDShwZAV/DEO7ZyoNKdo+e2l/cGnAgDN6U9dFfm08YJ62s04SRxIoA
rNSYNB86wSCAW7JDYnUx17sq7ML8dCncc2lMyW1GysLzM2BJqUtGprGGvVdJoSkJgIsugl3IXu45
8M/R2IvqG6sfaluyosdWdNf7E0dG6WPSwdn7J3o6+Y+Qw94xFbdE9+Tq8EZg8qB2gjDJlrVWrB1f
+meWAiiWpLMIdkE8M/y3ceFwqi+mZXDlaJXIWPmcSk6AS096KouC3tl9EmrDc0wK5ep8ZZEGpJ2o
pP8f4d/QEFYbnw87NMpZx8d9Gw68Y9m+iWolIrBbraGCQdhwK1jVJTkGQWd4D9EJRa8b0YFZOmew
hlfmKDhGp8/5ZmiUY2vFXfwx978dwvwg5GBHoxPteO66iiMTArKhLIVqPYBSL93zgQKZux3Pz/Zy
bZ5fSMD1VN1R7Kz1I4tca0HkC3rD3Q3BD1vcNQUGiAcHYMWlyfWHtOhdsLQMcP8m8BVjLpimwi29
LW+Hc1zlu0Qc1Je/DO0iA4K40D6YkDV+QFNa/1o4MHHXLj5ItDf5Ao9P5o6k4Ene/ndAUe4DxHJq
tTYLCCxGkP2EOIWTEtJ0sNi/YtMCo8D2CV+ngXz8oNON1vyIPUG9/aXbJtMN3UUdDG7e8PtQJ6Sr
1dxxlg8Gt6CHzo31MimV7K9dYw0ArGccljr4vZRYMwfr20eeYlaOraJ0gf/YEC24ZYugKjxR7/el
kmlKrsCzhu31vwa/ZNvfNXxevhmKgLp6BNEVD0GpUhOT6P3gnAwDW8XCTzhDt/LIPUNbYxB7ocvy
H4B0bMf6Jb8zIeJWHsy3pB45pjKgePYE9IOrHZjJ/1rokvA4Jb37xWLXkqgi1FrsUf7bKwwEyDRJ
tDh+iTVVEcdYB0XmtOG3qqMrQOSpHudFEnjPzwkyhmsCLfIw3EUTGwum7KswgaMcFpkRDJ5RhKO0
rYgwFH73xWc1zg0Ycyq7nuVTmUMtQoGF/nmjkJq9stvP4G3E/Au0GXTv+D/DpoN4VnbsftAB0rB7
cmAj3WlNp5vTP/TNpw6tA+7qNvk27DBut2xY4lbxb+HgHyhqZEnxqyrxGVTgZakvej5inZa/ebRZ
6HEECR5Ih+2yVZcZPySswKW/ROYLUrrMqkgZ1tf03ZkQZ6AA1Od/Ns5dTKhl7E/55WuBf2/bXUQp
2xpCovF9Mnw2baarUSMWn/aNG5yXxkIDAZyvBhmSAYol6a2jgGKLyCH439Cf67HdFxWLKDMfoMr8
P7r3hTjYG/QAIaiOTAeLDR1gv+GRjzoX1RoE5EC6qr60Unkqa7J1JaJCa1VrfLa/gTgiSdOdnF0d
P/my4QR3t6fFByie1zeJom0JENQRiN9GqQhCTG4vBg6VimojRxvt4v+oRGs8Hb5VbKmzlPN58yZs
lgK6iLW1ePlHSwJhdjPB6D7GahxukTIM1sQVMkyVWSxHcz5P7WmOKqXdol2Jto2trnGhE7us/M1g
bxuhlF1YmvfjCKrHBIGHr2t2uY42OM6fKevQuf5FZbwqpuU21gb4To6/3LZqj3vHu5uC9H4PNRp8
+D+f1ZL9WP3x2n37UR93U2iXO3HCGXBNu7UpSxWwk7P3ToUyBKN4ZGZ8RJnF6UtR06PDMHVV/U4Q
byt3JW7EYTOP0ugzui+v/L1NSkFvhsD0IkRErbtwAYrd/PY6hUIAJswqBOmP9igAf/HYnoOeQwP0
mAzTq1y7TcnlYWfshRQxRsjdsAof2QUMHaozozuk6VhnDTAAXmFaJWtDSOpr1Zta1TPRV4NmjEeY
aWZjnFwM/RmqeBExvJrUsunAhvC7YqMP4cMPBUCioBxqGJbtC4Lf1Ql9FDoW2eehRgwZkZ7KLjnr
3lEVFdRDjERTmyze+wInHNSICDJHHZnJEPRFjkUqG/Ecc+oC9BpXDYD2LokrYWqeuIhuo4LEOSOO
UQvVjtSdg16C6GYSWIaBsFdlTz/P6GF1ntciIkgN6sa+2i6iSoNwCxUpzMzEG7h4h8+Fkv1Vv9xM
KBdMMk7dpjozN3fvRMiav4Hp/87tUOcAD+y2yRXUBhcMKNBfr48JRVUzYnxWAQ3BFs71lOJZV1r+
nMgqtNU3AfiAnlTAaSit0AeNs9RJmYa3H64ByHhDuhtqdKjRenGZ99Pa70h2IFE0j3xd/DtVUhLU
NyLsZST9ZDkkVZwEq3mBWRrexBwD8tOTFJXEtsSKtwY6G1FzoJxew1eGVoZZDquyZ9wYeddPoTjR
reLnTHvo5ehKLRC1Y+kl10WgCxrm8JlcGJfOycNsuF8AXwUzoruOH51lb8uznBGnpHnPTvGckq7Q
outTkdOpiBi1N/4p96gfD/m/3jBMlJS45OTL20aLX+Yp0jMxxxI0EOiRwA+WVFG45qRbG6lNw0m7
Aq6D3JgA3xeZCCqQffPBOXJBXLkFhtzLhBXwx03ivoXVCEikSPxt24Zu+/3Dj+qFr6YZqkiSrzpn
V7oA4hLuJL/EY3q9SymqEuHuREf0DZkcBXMIm+Nrp/BszGns5gnKVomNWjElNABuvgSFeaFZIF1x
b8Xi8TlOgUoO1cTPyVJEzGk+WeWpFJzPbGaeCE2l/VzmpAQFTxoweRhcCrtLikV0I/14IijeA7vM
05juXAxzXpmmz38yy7w28iLYaMQA06GLwOjrwgAoeFFBsfdZj9U5D5R1q4pC6Aa9uOv5jW4tl8H3
NOZ3vASMwoa6NCzxvHS9Hr5ezYgXGPykfb1DhFQq57Qan7dZSzw33wK54FwDXLCGk81iwfKNcqMg
GUhxb1m6W6PLc4vJOofOu54/i51lW9ISRu6Qnft6/c7NvxVer1XW8LYgtJ+g/vMTIbt1gkrJzTEA
sTh34yTkJK/jr59/6DZN4I6UsmOgJHGbUXZzB+oNoL7B1RaQoICV52cukGAfGO6oTLgKXXGaS/+1
8N0YWtDDUgJfQjHuet3CHlYo8LE3MtX7SElyUqXoOF8niE4lkD5Kj42wKKf7q22gO+j9oxHr8VOe
xOV55NaMWFdUilFgCqDkoxNEesmJfT2d8iF8p58+ul/LSTsD81P34GlX7bmlUXRe+A47bEjXoKSL
hZo4TlRyLFonX8TyfXKHFrNoog616+rrdHiyitLJ0B2ltsFIV/VHKW2UxAWlN5WWd8/UmJ9MB9/F
y6hs+69bfDsswpbuOcASdfQ/9Rm32oHsG/s18yKuQ9nPv2+OWFaMwv0q06+5gKmNZ0bx2jqrIcGX
o+bPJP5vzfYXEgsAyVbBWr6DZwyA/xBWZciOlFI/PwSB0SJEyOy1sscQDxk0tswHtu8hFeoSELEt
TqjHb1cBA27Q6gvWV8dpqVCcJTBju6y9eteg+8PdsSZ69YVeZeQ/xkGkRulWniquBOECv6m0KQLq
k1hJ3YY2ozeZtSiQ2XI8aRDcvnXt29K5T+3B56oOD/tiFCvCGFIlCCO7oq8uT44hSlkW628Uaxmi
Uj2/90fFlDxNMyRuhBnZubk+GQ02EkNwqqjFBSUxXhkKwcB4IJbDwO6iNKWCySbLsBAL5JEiqUR2
ZWW+/z0gxVm1Key95phWnMUTcip5GKbh3yI2rhcKcjaAVsULS543TsLhZOhImO/Ka285nffkGaMI
FjnAJRN4a4zfxLpXP8oYNlvPK3DrGMzk5buTFBtH1rjAupKgoWH+2T3RGPY1vRIdckz5dJPT6EIR
l265m+7Y69ZNx79a7Vbd+R4/GFmjQjK5Os4XS3kqUzalNzZ7iDB5WMzU1doUeiRDSSnD+G1ayQ5U
AEja805mJ99tQ6rfaJ9QW8E6WbYc5PNtU0dc7CkpcrlbzQd+tl0JcPeV2X5PG6e+9inmhNmpZWQI
95wS7TE+GpdwLw/9maUTRgfWyewmN9DqdUJFOTnjYF+cvPMdIaCDQrpdX/OPgtSXxf57lWhLFYbO
31Kp9EPE0vADnxGdSotfM502izPb0SoRn/2YJbRcxY3+m7SldIuSgergcBHNr6ZIDzyF09JJK7dD
OXtANTl7bbuBWAKef7cWfeW/Ino4oOxQRaAzEwE0p2OE5TC0ZT7SWVpzckJAZXujg8op7HO4GFGP
8t8l+H2x1Vo8SIuRze+fE8cpFqhDY7ZiJFDgtlE4bkhW4ZpFrCxc4SPlN7aDpv4Hb3E1YaPbfuR0
MtniiQsU/5OWsl1hbi2Vn2ZmrqO+p7LEp0u8FkjdOM5demys1wu97JfFRelyZIiny0CnS4gwmRpS
hM28RzHJ/QgMqNaPLKq1FVnTmGpaYa3deBqPBfjaewVzEW85fgmHXjdMclwTlX4Sy4iQWboV/JM6
5AJX2c9aDmm9GPBfFn1SMR7pzvQi4pbzU7k4VZaNuRfGcW7cZSJy7K/3V35XJdTJF0dR9memAs53
igLZt8TxG6mhbCKwkM6bqg4GuffTTfV37ITo5nokgs0K2ABKEZza/23YoBJqCjG9RxzZM3xPji92
dAEcPhmqxhSY+dFEKJhRfzmqPSIJg0ib/zray+GJh51GKhASIBUMI8OWpf4E+EsrUc+P0BrdEked
ASWyR5SXcV8x/GjrZ8qoWmM5oX75tfk7FJmnVqrjh2gpneRMdgk2yJJlzGxXKNTbTSsFAAUyrvjn
dbikZmnthdAZlu8MDzhJ5ua3vqi94hJsmonEukoPWkoke+G0GBjSdpeCqwKPUxOpO9KsGYMunyEX
vVvTLi0NusAkJF2A0tP1WEw+GtYAKbkgDDpV0nGDMzeh83FNwmVBqtoDN7GHIJexqiwJkf8WINA3
6rIx+d80GBKIKH/HSZn5uUbT9OF3fWb2Q2B7ODZtmsVq6HCg2KsYp5bzSyL3f4LhrI+QCb68xoGU
884DsdMwwY39MZysWHaPyQYxXlKzo0/dGpbZy//HCQvIUR2dft6gpNt31bObhmxneuwCTxgcyevj
Gz53rCqheEKLNY8cFndpWF61xQTKNbEsMdBVeBloT54CQCXVx8JkfTfprHeuf57ErP9G5/9RkVyt
CKQxBVHZaOkYcV019hgXVn93cBjIotzoH3XWwn4pT6mwCUtPMyks8NLEAFe7Q2+Qux5nu1fdt0my
Zd8q7kbiwLwJKkBrFjiu3I5qS1PZkp0Bifv7aTmAW0Vyz8UP4Vl0tqcQhrVVhA46kyfVY40COPQg
+yZyOQondaZaTaK+1VuVqbsSSh0YWgyUZkpidpmB8PDJmkUgWOzRiEZnN9N/XHNdtW1qkws4hxA6
Aw68+ndmYlf/RILFdlRycdbIU0ozX1RC6+WMm6DjReLHS7fT1SJ9yoagjKL2lKeruMapon/3u+5d
Rf09e9I0fAP6ue1b9wZ+VBhs/NO+tjQafvcPeP8VPF8MjQ9yclgM2V8XPyP4wvC/VWvgdBue8Zvx
sHkGl99HB33fyh43ncv2+sYkKbeE248stMDoqUekb+ZIk7APjBRmam9SPviY4thp0sg66SfKVsFS
4EZIvDxavHCSr5hZYrSaqSauFu7rsA9/CyzM3wA9mLW8wBJQR0AKsws2j8FgqpmnR2f/cwgqUd7n
/1Bi13xEuK4rsplK0lcyAGqzHydhvw/FhKS9G9wPBqI6UlKOOqUcjf86ChHKx8V0oRriTSgcnvYp
FDXoMR6/aJNiDMcFs4xQcbrEcTF1VnhaVZwphNljTVCj+WIRplKj1qsVzPhqsa8AM3W/CvyJUSrC
hzhmc15WvcEk3SO0Bbv4S2og1XfWjIuJHUh2mMeT9PCYN/iU7Ab1yWJU4Y76ZeJddU2vhkOx7itK
P3D173hTWrX4e4eoq9TiFTqmXb8IU1RwNniLXoG93e/05hHUGhx/AK8/jtEXaGfBqnGsqvxexbx3
RxEj3loIxr6JjwaDAUz+v5mAsg4fDYgEa2Wo5/6mcllN6REB0IaLfdga8RXhuNgVQkPAKZ51GnJz
tL29pY6KRYcJvvipAR6SsARannBHqFBAE+hs0x7w0nkjPirTRupg3DqlGOfUSLiNyW8m2VJyIrb0
WJxBvkoHx4qVKfAK6vq2B3fB5EkyzBgY1RioE4HZLVL6IyzrrDnx04r1HKTXWBuwhZAYYQWjPOgJ
BuTRWslsw8nD0fAGBUkmaWmNvnFFAazmbNarCYCGN+LZm/Om+nlVepCB+kASg9kRSFhyVIW+YxVe
jwHbLK6cd2SYD2EUr7HndZIJf4T8lyh1MrlUMR+EieXlmi3FEzNr37uWF+LPl2wt8PFYJURqIPRB
bP4fwyS0Uaae/jUVqooxKgtQ9SnkVV1lGOm38S08g5A9g6m8PMcUzWlDV1XD16omnss0xmJwABea
WDjjFwH/qCCv4FJ9JNpnNmI3XLdR+NS38FVjiSHBNoRLmJVAtgnWLqhG+RWzLMmpCzUqDFXUVeTW
mz4YaDqAy0MDUTufjyZBGvw6ks5HXWYQFcKAn2chY/uC+zeXGvUh1RXDov1Pt50sqTCr1qTcrvzt
MyUCy0fmS/zMtGNSLE3E266fJ0yZD+TuA40P/fneutTpInxbRr7AIs4wt2BEaoynFMvhkUquW0jl
HydeZc5n0K4imCONF764/Zmt5emDbMrTw1ZE0nDvP6X+CZfPSMAqTGoIWKnuITgNzf45EZ+npijF
QKWvYHk42/aoQ+vCy7AYzCiQYterKiAjRtBIrXIijjxZBTUyQfMVbXnkeAwu82KTS7FJpElNJ9og
qPFq+Gqy+0iP+KPY+9vzAHLXXrB9Xq8xR4vDFCvd1Lgw1SAnAHpFwNpeTnkdCuc4U9vy7cSbyRkO
/XhXvD021OXZRw8a4xdg9ITYXHgC5GQ4UmsFhUTafxKm58RyF2bnB7z2JfXTKNN3+QjTIDpT8d0k
iOp0XQDTGS6ZygHKNAJiytTJukKp93zEtrqcVuNPCv/YC0gy+8r/hNndq9aRJ3a1w42z+zJ2J6Ij
64wSgRQmoajtngGgztZC871lzCzXfnXOEu9R+3fK0g9K4iY7L/H6bdXV5cUqUtN1pn480Ry4k/cX
EOdYlbCHatqWMj9cfKSMsiOv7X8w3m4CUUwu46nEwb4xm/GhGb8hjOFwMTOwrhSoJAHiyiuSccYy
61+GJ0T+diHD94vuzJXcrd+h3IdMP5fXCIw0UtOJrvcLQGnvXbg1+v3Qiaff61nxRjy1OPQAvfwU
16OITixrVwIk153eoC08nnEQirSu8F4Vt1dvGvNWnIK4xzcbsAm+JM7kJqkau7bYi2RfxiNgK3lV
PUGmCemHlmYa4C9UgkzaLo+bizTHgLaFe7jWlJyYSYWXY1UPno0q9FI1uPGstL6PcDrUJfBVdtdA
ITR4mFveH+yiMMFjw8CrNqiDEWL8GkEw/OYgsMPuhbdBcPX24HauRggmFwh0DrREcnrDWQE1RV2H
QlO24/Aui6I7vWAbauJCudo1nSawYopYDYk8+TtqIHgM8O2VerjGDUmxB/afrQ8nn1hm72xsLm7F
xSRjgR8+7b8vl6n/CdmwYNkX3LzLvjQZr+AetTEPGRiEOECdGLwUQMnZKapU6w5Le2DMpVdZoJZ8
a7E0I++y/DRvW9fUCJ4qdGpV63hLEmJqNzLvad3En4Fo0H0IfNNMIdxSyh5MmjRruhVjqZ6oBIFM
G5NQ8HhtI0bhDaC1Md9lBYXfU2+BhQ+mjKoAHRAzqCqzGC2wDzJmhpirkc2AMrI75Mycv6dT8utC
RaUp677bjUZT0IHatCdwSgYl9tjKjzc48muBmdrzKk9G2D2JZg/HK7YM9byZj+Yhx8VvTZ6oglY4
xvUCFisWeSZUN89vGP076RK9miQ9ITvdJ8KZtaNb828GMHPJSWG44LoX6lSna3B7sXWFLKbYPkKH
2YRboSBCyqPIHVbLLo1gqSFVPJNMr10tFL6TRC7hm+GTndvzno4zUVk3Z9mcjsslTKLCf4z8sCuo
vJlCP8yIOjydcZzoye11oCrWbEhcOLRcUf3cwZ/6qrTyDrZOk4UkK4yJlxgpOuX93krNh2w1d4oN
C3gLdgEQY++j4Mp/btu896yHig0Ni8UaJD2d0ux6Nj1M6k7x7AC/CoRVbiZ5BI3LdDYATW5uyikp
rlBfY1KYwSjS4Uljk4S4HqxxHtPV3YQJsQA0lJeDUxwPADtEnFlYt3PWbeKkPaVHyddiHzuEGGKF
kKxWrloEh2UBwRy+XJ2jY/D8ccnQtdrmC72Um/8Y4s4RPfjNGj5Hx1hFPbcLiCjuvostoYQohUp1
EBgiZeWgEEky85FhdBn4fK4QROQZcX+yhjUQj1AeDbGRbsXADErUaqc9O9dknNFGRCxG5mYfGErA
6PHoONOaHEZSmx1lsrWSrIMTboL1Rip0Zqa7Yp/XXNGd33FcjASW695q90LtnEsORh41BsUBFrQH
GA9w8kgP675/dg/3gqhp3MIG4JzzZZq7/Dam3LDyWjp4sFvmeSR1FbvGetHOTvPISeygkdFaNF27
Si9Sadnscw1fuqS4ACTkgR9k/ZTnUsQ/oJrSwpqFZkIukrLhijoAOjlPUmntlX6K6uNmXAm82w4g
gqfpEsAG++bxZbPVZtZ4xHDgWsJD44+TtqXb1seUPa2sVx2TY3vjmtDQv9Ir4BeKjBSdgclxshmu
VidqmiSWQ46A+YWOzfPLai3ViDIIB0DwtoK4WFdGjt4Z9DEdAsrh9bzkv18OcVu7B5LyG8VFMXaV
C3MzktlOOn+TaOVw5+1szEGuIV6PbtREs+RT1vFft7vbYS46N/BXl+9uAZFPtFxTXkmSRkD6tZrZ
V8GWe1iUdl5lzXR9K7od5RXe1IMcouj48GNuHgqMyedEqpX5Bdwc2gQadRMD5IPblAoMqFV0uxyr
7JfwcC7ygT47y7EUsh3DTyaLyV9MS4LdQCX+vDxrWr5bo7uo8udJnf/Th37Hp84PRn81nSl52s5t
ASzUbJnP8sGrF74LCB6gAoxY1OIznJkIQwyDDMbptrbScbf/5e/RXUgZh62vGnHwoKVer5NSxfTI
92wo7Hop0s37LFBy3rEXsKNDddUyrHDmK1uoExbwm2/BI/ZJvezfX2OLLaBmhbGSQ33UVS6K/+v7
bhg2Gdt1IYim+7o2uWygVQZls9/qcPZyQSzVm1hG+xrZz/gzHw9GUYtnCBDe+2xL9pf2xQn2TRoA
wUuueunIEgxY6cAI66A9RUJsFoVLWBGbg5SG+mwUoWTul91qqIS63t8j6OTPprssYUNF/ndnQ2EO
6co4L5BFD4BDrJU=
`protect end_protected
