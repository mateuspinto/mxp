`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
AiXZmXZ5SREFS5BjNpehMuveNNcmUTLER2tqN1XNTV2APMJaKY6MRzOJ+0QEXZQzDJl8ErEMIBOa
5/0ML//oOoZPg6EFf5ddxoNp/5Zt1LMFeLDzY+7DCnZH8VdQAHhbI/F5mgAmvNMCaqc0pKFcmNv4
iz33+XB37z+iuvF5J0CtJ+Ox1kVeASTUjzOD3iQhRJPHTW9i5L0qJJi+/8u0oAMkI8+9yF+y3KHE
yyU5+3BfKhIMz7Saj7RpSFpz6rtRHWPZNf8V4CuAdjW87ruOcd0rxkCotY/n1M1lj0bqKL7KTzgm
EKyeaF59pG/vOd1dnEFvqRAFCJzfEbC0V3R1AvPyxJPEoeiUcmbEetCCDfWzS3MF1BXVXu+0vKGw
cbI4jClq1GSrlbpTQE7IAnmttPKO1x4gsX7zELXrTaZW0fwCChH073AmeIHCuQvXKKZORJVtm93L
/uXQ9cTnzdu2D8uDf55HRiFRzHrS1ZQrGhrXmaHvaBoIorLUIJiXqfQWBc1+njw7aGpTq2O1JJ8X
QK1FdYbsbOz1Qbn5vfjOgXtlFnc5W7i7MpZND4/T0p28B4d+wbWYzYmbZgmqX63adCJK7gUVsMUN
xRVrmXRBS1lvZqjlFN5vfOc5nySoNiPFI2SHvLdPyCg86UBj2p6eWrpWKc1UFkKPbg8SxDGxhWYn
BuADjSC9O1UQ0SvMBlMLUQeMu8GdwWr56VtzNHWc+3vvtfEsPNOsD2fY47HICabiCu9FsFMwELfe
cy2skzDawacnGiSHugDgHFL/QVwMRS/Na7IcvO00Qw+hOZwabh0lZVZsS8gShRlLbyaYvXxrJ+Cq
MbrUqqZMo9iRPkGH0NKeCCoGyPBSIzH6QOjveB86bgQg13GQUocYWoTtaRnpg1bFSXBjOxYDJWZM
3Bda5Zh3lGhd8MGuLqcLmmrFZQ8zFhTf5QiMmRS0HGBQRdJvJ5I8J+4IUlVV0Jb7QAxMX6m917ty
GwcWYbRcYQgWg4Z17wnViiCaDr0+4XPUY38QtYcjhl8ZVBpLAwM9rJAhny4LbjPigbRnboB8FzKF
ifZANKPzLVkRofPn6vhLl4OAyCcsM9HovLWb5YT4fEHCTITzWj9VAe7qam7wqLL1MpYV4b9G/xSG
IaLMWGHa1LdSwpNis9Yl81U4WeFFXaNL5ZD+lVWdN58lWbXfpUVjkSU9GoKpNpqQHnRgtvufwGlY
kxCCEb1WD7kB/1GkIb84Ilw90kvJUYpzNCqPfvZjVom0Rvr8XSIIQhc0VYwhJfRDm4HXmCmtLuk1
ii7/Huspc8mcqrw0RmZNCZs4vbDAmrt/xZc7rTmxPVq89BPhI0A5t+mYCkRE9BkWqGqT2JvMFQsj
ODZxkA9mHD8Dtb0AkF8jjEOTYRdBvN3YR9RehrgNz4KXYspXrXwVt6cEHOXt9oO/RTznKtJCM3j0
Wt9qTtAc036Yai5SS+u5OGrvl4+UBI7ulkoZBn+Hr4NtB8i2+KH5XKvBA6JRf7wQAWt6ALIda8Mp
Rkn0nZvJZ+aQMEebqigdUfCtj+Tb3atc+Iumrf2873oazpQSgBzUm0RqpgGIZF39VaG6P6S67Q1C
+gebDFjMkz7uPgqAKgG7nJBFAxaXhKt6NqnuoBL6+jduGoA5BNAqT3qsw7PIVLJy8Dtf0+cnCxJo
45wivXhDQCuZgJBvqcpCQp7hCmr+lZPZgZcJhyi4P4CL/++vRiNG7eKXRwIFwOnWBBlVuDh+veQs
7+IAhxwRxWuqKcdj1o9vmpWhKgtxVZWaY4JIk/EgqDOzCn97RZlibIn/G6ClYBIGxaSG7TWDJ8H0
MdAnJ186kofopIKNdwamlhHZr/KktkxmbnmBDMsE678/FJIY944DcxSNNLT+kojOTCB6loaUu+np
tyKoxhsuEUdXNh4GuOLw6BWSDBwNQpmPqysguOZQ4zYV6fzQ3tHPJrD726NFMgzeYmn2mewt24ak
NpiiJ8ssnbcYeP7x1uYzW9T6S431XMPoy4uvUTNtATcZzltMOTEZz53FwkgWYTXiKIOnneZNDfH2
N2lDdbLqeyWW8OLeisdaRWLPzRTmCowG5248hKw6y4cOeCMacVappPRfqgtL+FcfhFwcLq/ECOVH
c8VV1rTYO8POc/gC/L16xfrUhp/gFJWelDLCfjnuoI48HZK64SZOKButbdoskn/+knXb8zIcnxPi
vzbMzXOooieBaEfG3ZZkXGu3xS3Sm59zmJn9SfFuZYBmtSrB5SRquceFEP545KYEywDM0Z4yEuXw
am3VJK2l/zchtxgzur87Hevu3Yb8ahkii6rDie77rQl9c6XNcb4DDT7v4297H7xAA9n+ZYkv9VSb
bDfUFflLPD8Qv5xuNer1xeLVWOhwD6LcjPDmQfSNE2NDEHoE4DL553Ep/uQVjNYMx7kJkgr8t5IW
nFNFuYOjhMEfk1RZZ+bS+zLW7Pb44R6GKTkOQeR/6dSrh90NAVXar0CJDs9yl9Gp8SfOWx/qoH88
sDEFllbB8lVUMP1M5Ro9ttu4cCsQvQi+j7occOVWWgXnJsWENW2mnKg3Bmqn708pMz1X/eVBYlX9
5gZugpVQCYPM08VU5xXP9pKL75RENkycSvy0CVYjdVUyj6ED23yoD3PHRgC0pH6/vxQtJtySFGXx
nO8pITC5pSFw/008cDfkzSi1mJKun3HGwhko3pHLIl0Hn+8NzepyOP7AMNTObEd90e12jqFnG0Xp
9+RmFwO4qAvc25DrgUJqhtY7N4byjzZmZ9YShT++FmhIoO6LDyJmBr63B/uMnEX2GK6gb8YEVoux
5yFbvKWzU1GAgK6ul93cJwGFaGtlq0cnRZYXmr+LaeVQ6OBiL3BQL2IpmEgpLmXH1/PKCnIxEyTa
ttd69Gcjw8LV4JPpSV6lrY46hhJ9TI8eW7W7CnZKkZN/vPuqNJWhG9Yd7QDfOwl5m7PAv4tyhS7L
qCHKo7tkoMIvdXWVbSj54cJOZeMuGXrvPoArSx30gJKKyOmaT4VhflU4r9260xY2/sVmkiChz1v2
vEwWeBbnp991GNdmGAQSfxxf/+Ir/2+apQn7gd6+CSM+ZBLRugH3eGc+IAhrSYsMqY+tfbx7ttOG
5XSVW7g7QLz/sTJ7bJPTR4fKnhmtSS0zrJpjjW7xPB9EM61+gxnQ9cxD403BB9OAVbmQ5RsuJrbo
cuW6RbanmtL0VHyqeJt9nrQF5BshaBN8d6maEcdhYWWFNwVypsxt55zO5tNJXEmZJmq3a2UkgHno
QHAUZt8tny0c/UdXVVQLJruIGCH71Gl2kVGI5Kw28SKtm5ZGN8OYCeYWai7VkOKJjD1Pt8ppdao7
AaYOTFeKGG5pLnKETI8+20IU14KwMFxxG0xd+j9j3Ht7wmeogtK7q68OJAapyaddhOaqRBvT3Hye
J1CzZ28dT+DIxjFu2pZgfbkGfP2f9EEKlHd9vUiAYGGa2kfD3NDlzJ78lpuTDaEFTFOQ+HY/N2HO
YfrO5Xc/eWAGKfGupI7GrOMY1ESkaJyAUROIeCooJmO0buFh2Unaa+EsAKl9Y/FcXwO8fVYca8wq
kPiBaA7kz+eM1SDh+jqSpngFNdnkmA3/eqr7xaCoE2kcHSZP8/jpg4gi8dghhVnG05q7MeeH27Xs
kFad9P2kHUpGLalkvWtILWFRwkSFMC4/GNi6we68PeLbtv2CPLedA96xj2YmilMPvkqYVsjAU3p5
ASFitXbVJNftZK1fHorMUkf17aLXzPww8I1yvhot6hOYckXT/id+vLQZ7zqeYR7vUycZ65as0h1v
ncL+zAA7k/IfpLX4a5V+4FGvlzAzmJqXMUNNlB+qxf13F5MMPnKwdkkQnaN7glXCLiT1srPBJbYK
gIsARoRT5nedMAIOdlAqQwV9/Gnks/apCn72+M0ntlnOIS0RwPZKF5Vl0s99nQAJ2ZI1yX7uCTIK
atKN9KNVrgfsUnDTq6hZ5tMACGuANdTvB+MTE4/vczBMK2lAeWnE7t/qsi60T5t4gXv1h94jte0y
UzDNqI88Vbd5IVvE4Rip2dIfmbptsRmr/5W8uZIg9JnTL2gX5V5SQOHcv8De/mTJt6TCTHYOSqlF
WtczE0TqZH9XkrUxlsaO58Jprhr/cE9r3AmPDcXOocHX1qo8mwqBP0eUXvp+aSni9hhJCuw++cSu
lVz1zcBvEmZ/4Xh1uQDULlIUUccn0nRd2ssqZh9CxQdKf/++Y2+k9kZ0ud7q4vArRKGEMCIwboJG
Sy6PuCPGAZ2ZzxpaNGyBEhvzmzmMsqayERQQdlHYGuFjPRrhOREZg1Yy1nJopHkxTJvh0Jkzfl9v
k5VXowJ1m8P6g0DocQH+1dezwocIJshrD2B/efHFiAUkNQxDJNs/VsZQ2vMoy2Qfv4XjyxaWXhPg
HVZrkYVVyQ2sPIhnndKRY19UJrdY/7IzeFa1b5DOFyldjJh09nLIJdQRMLO4Qu2OQii8/vHbMIOd
qTnfOPcuB2805X5QAe2+L9WF7XzWw4KRpab1egGxOdu39xNoDAwpj8bGlEQ+/hft7XyRviHQVtHo
8w0pb1Eilkko3Sdw4B+ei9mG+LnL+YhMcph8gBCE8x2WXeiPiulPk/2CvNfYnjNAcseWvEaPr2wV
7NzvJ1R5yTfjUJe40bQWqdhoAHTQjzK6PqziRwXhyCuySROLqqefu6moQgm57MJXFv35ZQb3mhP0
vBHeZTRkSh7aW0MWnGbW04wduW1dDyNuWz4ZYwwqDfdnx+tA9UGaLnxHnxW2g2Ju1KWnfoNc18yT
bNYOWZezQN3GIfAbfNBLEH11Ins57/0eP+NBQJqgRacGzJziHAZ9xbKXpcYxlbsKr7qLF4VjFwgZ
8hVZWeDo002qz2BUgbjChxUHpHEUUWnGJRzd1P5i8ZELdYXhb9sWNpvJLHgauHyhqWrRF1N43TWI
SpH2sDvocF+uiJrK3XulNf7i3b8XGJcQeP3LwdFmhBZHuHMeYceKEPIdxjuoTBNGvTHZ86SSdb1W
pWTGcpEENaLihUqHFBggC83cWKIQNr8oKZQrU0fOGjxLZXbRYqDm2qsBFp+IcB9u3/8OKgb+VlOz
RS7c//YRYtqlmtX0ryqE7xsJWCjQX6fc0q3e9DGZxR+IXmghRfTdJ23B+zSYUfiUntLx9XVHtuN/
mKRZnR4Rju32c1VpmXV4lyGtgVR/YtxjKXSrd/Iv/ccRdERynzQNuNeoQpbWeAZJdYbhqAliwtRv
XMrqsBN1wg1unO9JGWIQxGnIt4WFf7LjbAUSIUiG6J1F/B4ZmAqITP/5z0Seiqlddac9jVt7Syaf
rHT67ZB4Y7GrZ0vE5IJexmPBTf3hMDK/18irMhx+YnokLeN1vOfBOIlI4+ODxXnhdvRf3bW0ZGCH
mmSHBoWKWcc38MvpaKeqLrVOtIeniZiROguuovXyeHzrrbyxSL+FH3CjnJVsj1/voLwrfNSciaxy
qQeq3EFbEAb0GGsYlylsENOD1Ee/MUV2RGRe0/8jBSa3nuvB+rhSZ8V1stcDxjEIP2hHvBftItp1
J6NPI6mBR2YyhUGzR9WWDON6Nxe45yt4P25mB5Xw3a0wg1ASGcTN4gsRe2Ugk6xeaR8YWz3Hu3u+
pXE8LEUJ9rSUEDugi4KJuoib8f7KK4Twpmw1CoT5v/vZEDeHYpUId4yOnRaRNs8KzZvlhkrOrIcB
CQ5eIKwJFNHUh/5W1Na98s0scO+LucDO/6uVLJ15z2RGjsfe9zs+dodixZB1oNsV4sFvQlJhFlws
cjkIryuv6UMsJ5rDAP9UWN9BQcEoST3GCFUUwQq6ttdBfPDXCz4xunVAllXZeVVZXTkVK4We9E/k
9qfihlZJ8ddM+iwbAAVSnPq6lhMHy72kSS958w5igQas5ObBEoc1h3iPYfyoD7iPGV4fX8Tx9wCZ
etIXzrH4PdCIeTZ2jdEOtv550/yD/KZkQjc6XS6UL/OmTl8n3HoYway1mrjraFpPEet7jh7x81r/
IJxHi+yiAVPvt2ibKPqQOfXaStvQB10nXS/XlyOOxGtXEW+IsaCmubikAL0+uZP6v1tqNSUXdh0H
B1OMja25sqxTMhfZoxuMajgxh44WC7uS/SsV0XtiI+ynV+8iJGH2wY20HGLT6YvspGfjCY3IWnEj
COH3zF//yyO1DVzYMqU+QQZZykO9OHqoFYwAh+ZrNBjfxPp8wxEHRTOSNLZNJ8qC+rCIgGi3vbxq
jTQRJNUMsPlhk/CIflAWtI8Ts5dcf34+Pb84Xq6N4/Eq8GYh7L8kf01oEt9yDWNpjp9QdLCIQDFm
x1bBhvsq0BYdaWzAendfpXX8CxudIPlLfN3Gs5ixUUd3GlOYxa4elbyhcK91X3HnpvpBv5PEvsna
5eIkiixghSFcwjwE59kxnCawyDcDvwwnwjd4hUh93DtUrC3/QIWhQvV2pBbuogRSXFA0PPR9A4sy
HdwuIzFeo2ogyPkuareEiA5elFs9qDfeiYpDxJgTgl1yqLUOTGlL/W6zrp8MugW1ROB/7nJOvTfL
O1dcwsvFexvvFu4CPZQi6d7X+s7psxI/Dk7Y4pY5iTtmtrm3ke0fCC6ZoJMu6x/OWLB8CMZ4Twhj
/SVLMnzV6R9TAKy0WNAyxPfImn2yJCjXqyA5nk6RB0ogY8zhYac+X7j4QWvM3J2ZZ780Rzd1BFDU
8VX3/efoRexSmX67wunkR2GrpRb+kNFqp+dN9AMtMmcygHvui8bK1PwtvE4gN+sfBNtlO+DpL72C
Z3okdMypMokySe7UQWyJhWXqTTpb13gXLXRebsny6b1L+ulBymyH4bAMkPPS0huuKTQBi1uJ08ui
WfdUgpQfiXXCtphFF2MzSLAjB13+t2DVRb0mtjTGCg5sOMjpQboY6/9+YfP5+8FzQYuJWcC7WyBJ
nkFP9nMXb2kZrfzR8sM9Z/gVEWy+rueBh36mpTRwGRzDZIJ9RGMfQoEjbBgaAXzkfkrzCsbJcqtY
11Yifo0WiesWj5w2dKBXUW5O5HB52CBZOOm+so/JvswoiR/TlksDBjnfy/1AH4IY93Vk+DMntfle
ZLEHhrCM1cu16ShImKR6p25ujZpZ6z8pDiNlZawTBCIQAD9vDVFdfZLPCI8Ng0CBfSpG4yHPZy0W
3Z+Rc23yv7E/WlQyeMBL8fJcn5VHqNQZ6IdzUDFB9ABWmX8XVIcd9aJAQEPa/LAS6+a7hdPSa6v/
t5G5RSaV5fUKY85sVLDkZ3sxiujnsOm6NDYigGEKlckiPlhMrawtQs2gGAQ2nRbxC6eZfUs5N+y8
QIgkjlhfgAft98/nYW59bc2hWqZVasD2vAPhFEuZX4HBQLF4W9CutK6jExtswemPwT5ccodzSMcx
2q6NeTAseDcixEkJpSryJHogdkEaaFM1H9GEtVgYaN80j3SgvgEGc1Kxn+72nVafa1wJAayyZri8
XkFemCiwg5GXmiyLIRHWipT/Ru9pfEtY+hDiXgJ/PnkNw0eUiWxCJkfqtjXuTUDQBT/+jmOKE+8b
yxK/sdG6bLw6uUKAS+rIVdToax154q+tKIvuo3t9IVOhK2up0o6HAW8x/WCX8cu57JeWrPBObUQN
uWA1s3f0L+2BMKvZV5kPOugGCzU8qrd7/EM3tqWvhqAB2tXuQx34iX+/Nvk2DBYi16ifsuBe4FdE
vvuH7ASsW3FUnOHN/mPmuQqvGQJHitEhxyBy1FUe8y604m90wdrkKC1b2WT+38Gy8Ng4IpMy8gb8
wVpbf4VD/dS2MdtOvw5nOYrhGjlV5TsvMBJpYo4RKnT61Cj69xIs00fKQhARpS+WzqOmNwLKoowl
09O9qie8kRHPS92u8d1M7IYE317u6Ysmk1Dgy/6dmDXBssHgs5z2hRcyp3t1WI85B931fOz8JQCN
GGuEUxyD+LsdwelPjOlPVPLoRXhWkb3mbJnHjso0r8XGPG+hoebA6XJaofLjPAN8oocnUwu1St1H
y8hnpr2VYWsegYQqlu6I0vghY7YqoQyj4JgbTAn6c8vG4+gzgpZdGDqMw3IDbCD1rhiJO6KDa5il
YjRRzNkCHvnJTZh1/k3CFLB2BZykTmT4yMjySyuostiSPI84LeOITw8SN7UKVjgyYJj2C0AnWj+u
gYw0dGgVL8ChVY9Zfiby2equvdmiP4P+60zyZWQpUi5CEu/yrIRJvMgllrT1liO85wiDas3KjknT
rcP+UTP/OfLDw48/lTn80J1GyDa7MJJ38KLMTob2e+kOGTn6VBsbDzKWR1kbqEUFQw5anP+kXunw
v+0A3t/96UZwR+lva7BD2O3ykAgMouRJr3Z5EMa3IIrGXN562hl2NWbUfA8ecYPteBSFV7Q5l8Ts
B43wQNVRKCLdEv5dBAJpqGEujRcwhOGbmuEDRX3ow/v35FJGUO2q81RSCpzvNh9S9/q2Zhjal8jd
05axMXhyAcsFitK58xUj+75FgvTfrJD+yCPNzWdl2jUi2/pXhPVVz8C96LYwIz0hfp0z40oVVtKR
eaa5mgksxMRtbxfw7RiWoEWlYp1TCQgGg933FexZ9WCXNDbJI372S+iDrl3SwIC28y2D5K7Eybpd
VH+Q83Cex1455sVKVFBNMRh4OltUMDSvGRUEaJCkkE4S+0hAri7QPyC0X/HK4pL09v9YvjwXodgB
3U62mCnZK4UyPLOpkpfWtP35i2JnBY0IjIixVJcH23IoS+7DLA/sQmq4dzKsfEY4yA+LUSm/A/BO
nWLyiZGyOdHYc/245fL/S9mjk9I+6qnHxRXvbBTH0+3+Mx+Cizp4ZPdkB5EDhGiBockyjWkgjimo
6A4W756ZW8q0Yg7a6WM4gyLIZbHbI8zY+d1lulnZPZ9V5dLtMBgxaXPrhyLszwM6D4U+TvLDXZdB
AO6dduzu5p3CtPeyqefuIw8Tyll04wW+T9r7pT7dnUbegTFv4Nc7C30iJkrpQRvfJx6hax4P7GbG
akItTN3nZn9myPARTTaydaX6VyrtrrJ6Iw6SuJhmWFootwJxIVniPMHoUkhwf1ZX7mx3Yk1a0Y0i
PLn1likceFxHHZpI8t+DnLE9NZ3J5LF0q9FKivMB2RKDJhb/tSOonV/J1X19wPyZzZcW7VZDXOlq
LmnJ8bYXVUpUsOwUG2W4/fmpS41nzrE/7knXeDhmKgsYKc+Tv+VHFqCavOyuQyzxX6Sb1OqKzJBc
B9ZcUVIN94Sqclyn2BQa9aoctl8i1RYAYZIxRtxjxrBeju6CBzUWUTTMW2soCWW65YK7tClXgwJV
g6CYhcM8kecjTQ98BEfnXRQ0C68EwCIhfEAzFhzj2mgFvLPgC4HakjeZZ3cmgGF2XTa+mz1SUaCn
UUEfFq85CaIyj0Te6Zk46SfoOl3+EPqddt562jQJucbkkHI5j5rAh7SlBYdhaN8o6Dvs8jDW9ACG
cKvBQBhiNchBrCIJ2ki86TDxAjvDVOvojQUsNENBVGHSPuEuCO57Q7U78QXDA4NzX0oSx6a3Ktjj
3+hhDPb6xKcPHrkC8NuFNwGWBtEYCUNwcJ3i289FkTrBGIpWSVtgPDvUx0M8b/C7jAgdLKIcunZc
JYmwiTThJlWPjfW9KgbjDjQ6KehC408nz+8nj9lpN66rGPtGRdFums+XRWCttlonhSMa1q9tJxKk
y+PxApSl4Tbd53eF0k9V6vJ4HtIX+qkr7E1v3CE270vLgCuloTA4IDzbdrU7aVEpDsgQRigij7dK
RFi4mPnxWa4n7lcaX3E+usQQeR9ecdJGdkXu2VIlgKW3/id/vs7Wzya1KxzJ0eX9nlZJ7nY0Ekkp
p38B/VpHKMlM502th/yJLitUnjxoGIEc20/YnMvHhe+wDnW9iSjoz1B5LfyMQNBM36PcnOzWjr9+
96Ch+TEMq8Nfjyx9/c8R8x9XibyEywhMgWlIdgFONLWFUNIYs5iV8v/WRSOikr3fS9uqA1gyazhM
ptz3wcZ4DaXTWD8uhxG5cXx/kcHx4sNwWt845jE7DL1pFf/fitNamzFf7KsVNQiJgVmEmBSkQxn3
DhdNmAAvWkP4iWVpOhGcj0xl0bSd8qVusq8FLU24FtB8XkGHzxneFUfvEKUPw3eCBgQu7YUsQRoD
cxYVwxwmswe82N8gqCFOi3NS00BR7siSRUlmFG0vNuVPil2dmHYIg6TjQHQu1vQNPVvtEcQmY4gs
pc58ESopxCnyFCHjAJyu1Pej6huLPFohq+meJV27ofwrYodguvUZwgOAryPfMAHRgd/r4XNJ98Xo
PH5frtbNYrMjn3b4UjyA3p60i0CgquEAzTyzSOk1oqEMMFJB0USYDUC93BDI7TqwNDcvUCUlcvZZ
HTnCnUr3CFCGnqCqn9n6oV/fgR9SDWpCvnyBZQjLqVWJ4gZKc6EfvW7xcOnzuHHGSSrEx1CkOOTB
IGZiin6/wzZ0ibgGNyuNz6FgQWMiFQ/6kv9WRxbYuZaNirM5wZkPND9fGS4dKUmfkKBfLlAONwpI
gTBQu5hc4NrevMKhHeq57KtOSp50Q6C96Mz5CBT6ge/zGURHmSmuEdluIDvCbHcZCeU4VMa1c8du
cjNBHmtZrE8Yym7aVrH7XG/g6RlEzWgRubpj1Jm5J8jrVkeY2HvLob1pntNmf2XRfZRM09kJBc9+
GnkP1U5xAljq/bhH3k/IDwPKxMrDTJ9IWs2dhsVOvnvv1/8ySmBLl433LFx12WLL8Ub6tTJzIGqc
KzmAhW1HB62D/Bb5lAVvNlo39DZ7u6BlxuqYrVAs5KwgnFxnWaSZUcUm21ALdjbRdcN5YBWWxXxz
yqah7SbJ6Yr2lZjmw3VXXYXyAAWQXhTEn5cWhzzPP8Cgmo621tRuAvmr5iW5dsHmLv57yHfde3j2
NciAvC2e44QxmKBBf1F15FmK7253GS8J0ZFKhiDi3NmHkl0zxSGtt6q8cW7WIf7H2MP+v70QuJsX
64gDyDI0fgM67zFsCuhjxK/BniDBe0+/Ns51iYIUlakXa/80U1bwC7wb6ckkpuTyQNE48gm/C3GW
H9+baDUX50tDeiCCkM39dSsbXsfkCgqpsso8lhm7IGIT/q+Br3fClPU+FVDtjEnSbnsXM6UV25Zb
m6ma6EOxaddVZIOFtqAal1arpKtBMmFmQRfQA19Cfbdk7P+z7gbxfsZzUGK/b+G2Haauasbzosxs
rBp9pTgfZ9BrNgBMrA2WL2Vz3vjmmeXucszzObhcbjissI84MEbhWD7MuDgIKCvW2SDLd5Je3NS4
7DpW4gElw2gJMrULQiwC8zsBUKD1QvoGazavUizhbOM/l4+IQGzTxiiyQnuaULLLExqwCIQB2Bgx
bM9qgg6OAyBpjga4erqc72HMRBaCgOhN/JILkWZr/RlYymQAESAO4jZQI1LPsYGlh/MTMXXRmX/e
GOZW1WEPfKfTRjwiqT3Ctrp6mwetTfKCDwIua/ju4cEOl6+YzwzejU+twjy8urbRrUrtdBLara7G
2OVYsjvXxR4uSIZrJ6MLylE/LQgSZTLzbDx7v8lWmAaWxLxWzea3Wn/rtphd9nGnZN94QO8BEdS+
2827pcxvQgI2O/yMkiVf3PShWWZok4FMLe0CEP2cgp2L5GpsU7iki3vTZddSzh+bb03olO5v/yG5
e9Q1BX+buqhDEZF+6WNieQY7E20Hcoggj/OoaAVk9FiSfXuFj99QvWEaKsE27725UqP58YqCVORm
DqgzmLFax7h/Fm2H4HEBlm2ecCTI7beJByJYvZ3R7FAbqCohKL3FpM/KAk+DBbrfQWyNzfBV/aXc
byh1e1rHYaVdulqQ5XmVrmmSKh7km08sat0aVQYvA3cODvuI+wYPvVYrAK5pYIdAjFu1cddP8zVw
2Y7D+Fmr7zgnQo1AIUIN6I78LEpeTCcfihnhj0LtZtXwEmpiroBjjLK8Xg1+GV5aIF4Kz6YTG//n
xAZubyCpKScrTYhhLSyC2B3eKs7G1T46YU7G+DXaNqt7/R2ry6Uzq+H75crKT5EbJHie8ybx2mgV
AcvMxbe4GAVkHVEpQMuRGojzuo3oMKTicA+/lkaPJ7PCHPQtaKQcqeCGXetDyc20j5TecumLsT34
sOcJWw6B7ngcbIQHyLUqNqMl1RMRuIrs8R8JRLqBfDZpBtWJD5T7nsxV2U5eV0NAxQNmJfjKMnRG
9tKrg9dLn7sD823K8IxLXLiKMORvrXVHqyQlgZNyFOcchBtYadIr3pgzuOnp6BSHQAcnk2ziobf0
OPk7fO6rdFhVvQxwVQRFuAfcr3EmoHYHr2BWyLt3LEgRajF08Vgn50H1qFlcWn9+YEjOWM2oBBEa
LCzof9hLPOOqe3wfUbZOimecSbLHOCGSlY1fRCZ/Jrfc5m402y3sCSwkoeOScaLP6AGjJjRIcUek
dZBXWW8mX2I2sU/9SpNSF+rXU/7QmE6R3y6LT9eAXIBfJXKlPL9CdjgTIHpPhtRTrfv0AvwBFeg1
tP/uZ0Pv+0kGCTc7h+Yq6mPZciMP/ZWnG3Xvh8SPkhaMAk62JdBmfb7Z6n9kONXH7uM1KvEQp08D
pFnwJKuLxsrBIAbdLE85X2LxM/cb4alwd0HQ8Bu7J72IbNAI/lo2amzmC2V5VpfMdazic5cKI31v
mRgYN/NCu+gzxKy+8G0j9vFPkzM/LIHwuqxqMJbxd7xqX7usTMbOWkUkzIleYVcm9zF9bJ0UN1P0
FiNzMF9cOn88/XAYgDhATZoe86kfL7BwmWyWCn0O7N79wjxQEyCbK7xZLHeO80b2krcEoQn3RJlF
JPTf1pevVHyCFM8rUClxahHBSZZa9wx3jerwc4py+tM4zICaWqiGsihOfZpCSUKiB/yInlY1uo3q
F7xuzJ7cMtFz7d5CTk63BEYZ3Ovl3bNcBXAe9Iz5uAGm2Ef5ztU9QbdmjaG4uQICtNWdxvrCOdDG
Qvzv4cV7gbPJ1Hzpds+Kgsk2DP17jrvpFqx+OrcfVOL1fYo/bSKutB1IBNjoATGI7kM3V3oxKLB0
//mJwQ1WZu0Xq+tYzVQ8f8VkErQhO6wzPaPYTgOfYjXmXnVOoTB/xi0Imi/6ycwx+Nc5i09bWbe/
vQotPS2SnJOmCa7JNg/SaWxVhiseV4nIfFiUEw0fvRa+DVzjDiGePU8FBXcmI9mScUG1O/lD/00t
ZCgDIfmDZMh7OzP1epENhZqyvWbBeMu0Ujpp7FW/MbDzRBY3vh5YjXVD57zH/JioJ67hGxlktDvq
rnsCBjS/AvhWdijzv8jWHAjNqWPdOIcr85X3LQ0lOQe308sJFi3PAXEmwVOs6DTpakqgddJEfd1c
c8ls91DPZpGGzMq/hnRsBebVCsbunM7Hp0+WO5qBRaWAFXItJInT11YNwLb1tzwt6/UlfdQp8g7l
0OAvZquvDOOz78vNIlFgSuN5c7+4lYAR9hg228QHyL0v9lrdDnmtHSkccWWqhOBf+z9t1MOGUsdJ
bDSvf5tan2Sv1XXhA6pPs2W23HxvzbZr2xm3l/Dxxj6cY/NebiPmaTZ+uBHMyhrKMebqeATFZloR
QLlQlBlQUMePOwCHZyjZ005LXiqhAUZ7DRHywVvtyeKy2SKjwiKdbwc+pNt8Pl81KnWygfvzxkn/
2N0OuTDJPAg0y+Y3nV9X4IVd5rDBlqkQ/x0aGtwCoJICDQNqiLo6ZrWPBiChyAs5Y043VfXrYL9/
mVILs84MEn0UI8lf0kTjR0pxxVyTi/bwW1FT8WD8bKOzO/gBmtIe2n1egoEyDhX9V9K3b/6NA8Dj
PCfyqeNHkmjrwfpJKnhuSzUTF8wItB0a4Szl90XqBznbycNv7ocIPfEpPke4O1s5mVlo3Unhe1Y6
STBUNVYqm7T12Tsc93/BP5DmtiFJKDmxCAsEoIqoyhqCg+RibvuuAaC2Lio4qkIAoa1K4fX5U3tk
YW8ZISUG1SvoG7fYCK+v4Q2mwAi6dCxeZlRrpgrOmPTiyt++M/LCAbyCx+qbpDqbm6w+0wOdNEHw
kucD05yAKPbchdv1nzWXi8VVTSJcQG8QikxdzPRG8DaJaP5y/nu0bj5yl7jbm28N/3QpunMgzlcY
MKPKPdMo8b8HpfwFvP5+F7IVswKuB0Etr4OrXk64VukaQRP2yD2YkZqsvnDMhgUUnW2cRdIMNF1K
HDl1w6IafC3oGqjSjVaBwFrxgk5PjAQaGrH5yo2KySHzelhmlAwRUSx0EMBtZVR5CzIy1hffbSeh
FRg5yfHfvawCL7ias8z9qLBP3/aG1GWhXwtMykSYMrWNvZQqdAQLjuzYng6HNYRbUdcdQFoGcdP4
bsqHeM+F6bnGECRULlamvbucGiwD4oN7ALR7NMULOBAB5M6hTsruQXB4fuPaKWxiN4haUzFj6PRX
Ic2JWC668puLwcOPAq1OFDUXlC/HcBVK5TiOzsefwDDVOn2mHKQExipoPUdx14il+MLaCK9LbvFu
k36h1tMUghHDxpRVDPw8BWxQ9G5WDgR3Kw2lD2XEmoDZuvX2S0OblZrNQEPcdix8rgDrAxgzNrkh
R2obYLQygV82oVPCdj3fWvd83KKTFKDK+qkqyy3bXUdsnpXDaAzdS37NHwLtaFQzFZE08WplNLDH
/Jm73cWMSO5MPetZoGjgkGKz1mKzsgkRmDdvmW4wImWBjT9aELrAXzMuXhq/0MkZA0EtBJgo4vzy
Df6RQ9eooAV89UnaDTWmdwHbED3C6YF3yJizkZlDzVIJrcX7hDQTcWxuApkXGNvtPS63sRf7Hdzh
ZQHtJVTCtGaxK5QtVLEo1Az01Bw52dpALppmZiD+qtbKHBo8GPomJfmsn+hGs5Os+RGBDlRlob0G
KESHPXfq/N1ez4gNu54EvOeNZ7Zqo3+OVacsxPkeJcEy6t4bDrnfm0XxVhbyft5ucJu/EbJNeGdt
cNK7VAJph5A94iO8uKxNX1z4gxcOUm7jcTK8Zm7XitmOoohQls2nyC3tdkv8TgVmKtQYf71BtfWw
AmODWf/mGUmCzqIsD83qvYRobstTz/6+2kB7gAerFSPey/IhuAhuuhbP1TSGEOPJBYoU/mWrQKH1
CyKpx74k9nO5zCQjHuVBTLiLxD6RjBrsnnenP4PTJ7ED/fVcGQTVmqCwvCT17rV2GLKpZ+lhFjPZ
JMlGgQWLL7pzJd26fW5T3vdGEG/3ldV6RrxuunaotAg9XcNibzKFM6YUENInS81GeN1KuhcIvmLp
BRRzkwJBvQe0nsZ5APTrgLpuZOx8Wo91KEKk3vnqHSx1JABBW5OPYVYmsP7cgPTNf9e+wf/QQz5P
V47O/Mg9elk2WnwdGKJnnNu00F8CigF/jFKYlsSVj9aEEyR10CUQcxovKDcpTGALPhU7SrZ3cON9
ucLlcdrQNJxrQPPoNES2xhUygKE9Q3gNN5Z9G6gh4tzT/6r9udxpT4Pdom2KrqSDZMPXSrZR7RJv
u1FqIePwZOO/7WB0odIacMtbDuJfcGaKGiWZI+Si2vMsjmYzCdWj+QhGnKLsMWyjRaGK/1Z6fFo5
2YD+ASHBjKyTksblZfweUFP+OJNpfFsZNGbm2p1nBdLGZYyxe4wOgpH2fbN06ZFMwmeE6LtTH805
fu7VGpD+1e0Y0V0MCF7rtx637Tw0I65DNGBKRs2LWyUwR8/SfHULvmsnh9nAeNawghllCLc1Aj1G
xnc560THVsIZ5yQzI4YXigpBQRKrV1seSsAA2ZkkG7SLgm8UMHrRYi7SYyc2zPbRMgzuyAiMglgI
DCNOWZyVFQyE8Tm3YGFohcZOfHBwifmQgYYouMX3RPwucN0cfgQfGZgv3FElf90HgWoAiAwW4HFA
yGD+OqWOXk/ZLWzLxvAqgm2CxnTBslnJL2r0GpqXWlsJMUZBPtCzJQTJLtncVvS+TEpuCEzjKDBW
kAoDG9eXkviNv6GR3gcA3t2V+taT9opVDY5tXtit3lwMTwOqaoRi1ApPddtTdSdgCmk9s9Dg1KdL
EiNH9+4NXWcgPKfcc1CVZtIvVbR2sHV8zvWxbMPI4+/SIidN0agEDCMJqjtn4to7Emghoy7+YhOE
e0ocUDR11Ezwz2J6ifgKhyamgm4Hlrc9WLrzTQuCputRG2Asg1Ae741roqVCMz0bPO5HUGGmh1IR
PiK6735rj1/Vw0WtTJiGqcLPYbFB8duU2FKIyor+GdybT0oE94PUHAGq9GHP+IhfPFO9+o5JwtGR
CG9sYhvMiC7Sijds+Yx7JrBCvEB08Ws18wyCq2cB/NUA2/PTkeGx7K2nU8tbWdEvqWx7VmocUKby
y3bjsljmkSIwePxXT5HwsVRyhCmbjW2/qdoVJwLo5jkGPM37aZgf1++QLgustLwxJihvIKw7o/1Z
CiR/bRIybLKrrPLu/EJvk5oqFt/E/W01P4NN7lNZx6jMKKx4702Hb0yPGpIBVNN3yF+VO8ThaREh
rgFE8lka0zUSHglgvk0sGaFyiKnUp2bg+cxEAPvOUNWezx45WNR8KtOV9lIddJne8GZxojatQwm9
qbwHIv/TMBS5B424Lel6G6RG3BZH82HmE5siUIY9ItdsLzm0eBJknuW94NyM30SP1AyR4f3VjVnl
gws0BU2MigeHZeS/WjhMF1p2fJhIrZPCkEYQEHP6kNGRNsWeC8k9dSNfpM0OX/aDko9IPX+/1fqO
PKsfd55PT6NagwUtRQCmqEj0bVz73KnTwVfdgi8tK9vW4XkRDYpdyEtD2wVVE+jgEkoZw395wEgZ
SoCbAl6lt9vaZ2RL2O6dREGNeNuGLqAXqVheqexRixswxaRNZa4+PuQbBSJBgTdkT9uyYqRgBlwy
gknk4Zh7mRoyi07CTq36c7ky5kQg6dECXiBcN0fNEoswnGDEEXPk+y1g8vkKbZDUwXpyim9ClpUB
NHT8Zf9/+NG4VsQ7LrD2ITeuKGtpyRRUy1rIX1Tvv6iB7whM90n1/Vl0HKFoHYf+TsYp15aSQGHn
+55RCAFCCOEwy94AtEJ5WSRDU915Ta0d0iqU7806Cm/nr+eVxZWxL7iBG0aJkKDz7vxVRnH27G2s
0Za7b6zgDM2QgQt3SDPKWifEqYNuuvUmCTnzDa3zTn8nolydTGsqNmNASeI1rIUQHjpkb30f5m0/
raDkqHLqkV9CvZGDav01tsDH3FK40ne8t0XVro0w8ZmkHx88onRTxwCIHPmgdbl1IBRSaM/OYYJJ
VxbSrLmkH6l1Je70cUGQZYjWBX2+EcpSKBd2YOljQm9R5RCj3xKpgKE8dJQu1YL2yJ2VPtSOQeen
gixjS3vLSdipva4C+Rc01YBCsUPnmSbU8PDWC7PjKXdWlvI0M7mXAjOpDPR7rBacvcFLqOYMq470
VpAsyEHDUvpeqd3wAEajgDxG8nHihoDuyJmKVRRYJPuWAxb+ssC1WW/dq4yPfu4ubfd5hDCenTXN
Ss7HR8B5YSWJsrNXZuSFzC/6kaSSNO9LOknuTJg+jZG4zvPFmvWexwAmHyD8r44keq8JOjnvp7zR
14zStQoWgqgkda8bNOwGfS/yjQ61HAaz81qxUgICo51hLT5Y3E/q4ZQ7hXQaBvvWauhxo+Wmjtmo
ROy4GKClxYflkXPM2fLEDUj7JY20f8v8K4yCISmDud1nts485aY+v+UdEsc4aZ47XTX6+wwGwWfA
prhfL6KL6/RZJJdeO+dNvAp1M28z7aTCFhMpTROSvgtevuBoc5uXMkdS6i2zW5s7GtZQUgF/H941
jHPiG8qPJI3kza2DmJAjDs1aA9hRtdtmRzEa5V+fszdLcbl6FPFTpOOD2Z0UMc/7DLpQoVoL6NDz
vl+7o/UVf+FoVySpHY2KDTnszRusicxXQ64JHOfZi2yRE8L8XIyXjJTnNWcEvUbKP/e/bPGQ3yl7
e1TewHujaKmsW2UHW18oixBOGuK3jJkzEYSJiwl5jpLLvPnwR9tR9kFu9ePMXoO7Y7f3riEfyb94
hyGzHEO1JbxGFRrvLHh68gmsfwjHrXNz+z++sU88jlifPXr6ySzMXNGeWbXqAYmJpqYrO0CJRVxl
XmuSl+GdF4Ko+9xcvr76Zm9Rdg90PLfq/JZ4btcbiEnUb59mJXfKaRRUnv1ftO7CsFY71WuZI4Wq
d7vfpEKoPkaOaE5+mA+hFlUqPpgk7Vggzy25PP4bkKQLYJa2jjKfbQZARxReqhsUb97bJBvNz5pd
NxXbxj+NpWoVGw310LmzgmUXix5jSQVnxb0x31Y0esVvHhqLU6PbtAZ/OLP7UyrwhITO1OISz726
DCuWZg96K8r0GN6Oz1mQMnY7DYzcQJG6ttNeHcgLzEqB+GdttxHKB24fNdO36u1YhC7CKFJ0dVvq
CKG8/Leo7W2WThKKYnom85Z4GvIL9U+MJUjdriuxOHAlEjXX+pN/47h6clkPVbXBg6Eh0eS+AEQN
tYGAVnqqLsXFEa05CrZgRaOUZHMEdH3bv9zUY1+mE3ELvcq3EPVTFjWALE4G8XMZbxQZtYL/GuTS
B4oMPbKDTqmNnZ9kUcjjpqeYo+eB50tJdZKF/NQOsuudjQnz82fOSKoDrb707Z40RU+JUMfJbuta
tC6gczzAZm8hqu5sQROP/204Dv95QXly3C0WUCHq3+9pxzUL01VSWTo5wSZSx9r/MEOACqO+w5W9
RoK9ZmDB0u6WSetZkDVVa/M0LNQuXElvEOSiYSVMASlpuW8ru3sk3EuMbRVYa0bdfgYhMjGBUJ+b
2iVnSZ5V1AIWQAAMe93df65A6L2BZfj3gEtug0zYHKg+a9b+rY9TNgZfCHcYDu5wTGgfknIxVQ8h
7bvk4tAx59HcD9f8bdnWlxI1q1lplpgAtPyS/qQyOVCs3AnHCekFrVqxcNWCjNBp1oExIvvwUxYE
BV2vC6Vtb9Wfm+mNOSuQcjtg76AzbifNzPT6aq33wdVlWG1RHunQXJb9I6hn4x5/JnjAN1vHtZub
wvoSKYyUh/IY8NfYCiNCqiI1oDehkplsy4iSwK3YHQPgrt8C1+2QAm9OeT1593sq1/b9blruyQoa
CCWNkwBxRY1Iip9DbMu/H/8ZYFfkKccBZdNEQGmqCnDaf1Q7bg5tVIbVa1icc8cn7ixWzZDbJp0A
3ooMDytee12vVpl0dL8BnMQU+/cAtuu/+7s/gfv7DGLfM2fn5pARvgWO2i0fEynDAMDM5DMk7KF0
O4aGKDAV2iTvYxI+BO7qkfnTWLYovSv/Xw7dAAvRaACg/XHg9m6VdR6Ow5F+PSH+mWqchmVzBOFm
rL00NQMw54zLbI7+ZCPRPobN+bk2UGFFWSxCDj7Ghu1npteCU+bTPO31Tu5RW0gkicu91no8PDLb
e5YnTTQ++/T6BOwTRdrn0uVU5dl4NQoU9NAS9PrfhTH7zsK/ew5rQZz/ni+5lVmytyKzfbEpJUP1
M6IgD6T0XU+HZu4Wk6SMRMgNR2C8vGhSO6sVB8VAzmQLQckKDMnC4fXQZJnOgz9F+jZ9Qc8Amw14
zaWoj9x8ith1BuV3TOoo2nK20ZmnzR5iQjq65YaBzza2k8EKPK6fuCZvTFdCTbTGk0cw2yyIuOm5
tvpMmaP+EbudrFiexRrXUIe7L6rXnyaKTws0W8smc85CZjFtN7uMyMn+gVzbQbchrKgzQvfKJKlk
4/AkNw+W2C+gfpW+vyDxv37k9do9/frhUt8S9Ey8JdQQdZ+O4tk3u+3F4Vv6EXb8nv3Y7yGBsyuA
f7PL/kLISAVXEIBv7Euf7wVvQ4JYSqklVIOmSogOh77Fa5tV8Mwv6nq1VjoT+tvFEi/Qo4RqGGbg
d6xNMghTneqG0YiPM/XZ8ZT3NpOMS8+EAyFUEysufw8EEkxD8cBQg/UBdJ1hkqkLo/W0sIpapuqr
SM9eHhMtkSYn4c0vj11fHhyeJToR2qhY3YHZfCq99w4OStIduWZSp+6sDkHmNByVLhSYnZ+q2hWB
tLbXekcmjVOyICPoUpuhCLVSO5UQ63Tql1VHTm+jLSS77i74BJZvr9zTSELXgFCz4eIP8fnYsQAI
kLpUcRyXjVPCOe2mAu9CmPsvbyqk8n1cpVGTfstBnUkJIjC9vkl1JFe/ecEgOpHY1/AA32p8lQg0
sz/TteP/4Lowsz7lsJXwi9dnT5oNcb0ZpkASh1P97iMlwDXuxLMWZZ4xjPPC+qGrmq2fHjI5B6BA
yOQscJX60PwXTU6fCKi8AEC/W11KT2JjpfEZ57niES7HKufz9P0IicuiHA4rde/KURr/U5o9tzRC
HpVw0RMlKqTuj9DXJ1EM0A9vPQDmcdc2OSCHkcQuEzmOFj4tjcz5Dat1sdZ2qxXtXGtEIw5H8EFL
Ct9/nZqDsedOMAzh7CgV7pXORe/XkUKUGniTr8IocMoSRSmDfwPEdmuTyZj9xMzyyWPIGHAfhZQd
Cdlg6CY+f4tvdYhJp9EU5BRly7BhSUSjDFljbz6Z7YweDy6iWQmNj93diMHQibUSVpmbwNhxqiZd
we0YLDXk5GViQGFIeSkUFjp7QSFXiDui8auhtEosKG6WYOe5XK5BY9AUQOUOKQNauenO9aOFMqsY
B13052n+jL8xLZeAxXGmCCnFRzeoFPC/jwIUL8xbdP4GJ3xPqDPx5xtPHM6d9VPaReT4BI2kn1KS
+Hn0kHsJo8FoWH+f2/fDoHvZccJ23cCHzmRb965wjdcRWzZfdrpNknGxHR0PqXmkwYRJGZqlmpAt
lsyOVNrEdx923VjNFxkwtQHDWMfroLq6L3F7rGg0ysaFMdi06cmhCWU95A6fXicuLJLEbd5aVWuw
2Rb0x+utNshuNtOUSs07AK/Vxa8OtYPNhrNfdhdGsryRC9FznjYxdjkgUscakWujfC3cgBITqsE6
q1+CJE4e9q0Z60FUiaBKYAXlSDS69ed57HjOgOdNpcupjoRN/jod9blLMZXazPXquOtrK5WpoaYw
s2doE1B2nWW4nU+zt5IBCI/mVPItGGvz2tAPq8Hr02x7tsvdHnBhI+VkVRGV0p/faJm9yIINpX8z
ppH6K2jC/RyIXZxkRKgN4FA76RmmLCi46TwHB608atzeAgivXgDH6A53+04iV/8KatvLOn6bm2Tm
XcT2BCayaWkctKlAM0Y+CJLiPF4nQzy8Ig7Vq/ookQW6El2OHY43YSshRTtqEfSv70zlfZNdpns2
p9SfwSvFMs3ybRGof7O3d00VSJ3LmQzrdZPD5Is4O3Qd3V2eJyrPRBiXRLm4zTi0iRGYBbx5jlqD
DQd5dbOSqrRFZh81Eh/5NDnc7SMIFWscTjXXqzH3GLE09PgbaYZ8uUKR3LIsm/inxLMuH4zQvJkV
dnmPIltsQaT+p94G7p37HVeojjcTLRT40mbr0qZ7wYgVKvsg9seBVkyH6Zbxhh49L1WEIn0Bc5MN
c63nKpMbV39u1I76g5vaJSzZy2/jLOc4+4/kVlqSTK6a/6QYv1q3CQMXOrOF1mg3fU4F3zYcp60L
YVQm6igIZpLYWylQuAjXpcvoVLy2kQChUd/JpFhMzbIRk9Jg8uOC3Vlhud4L1tczyvNm69kQKYDH
rVEjexZMiCeQIvLvd7F6hDbnxWVak06Ab14djWewZy7gC33mTBopnhDLU73dV5MxDeqRJULcU0XK
okfsYRxE8zJM9JPZoJSqSJY1QHj7xdIwZ/ieu8M4wRfyBFY1donUqnLXCDONz2DQbhKAH5hdwc+U
a0JZF24BDj6VDZxDVVqpqcdKXIulD1Wn9R8OpqxTt3Y5hXdiyfotllIxH06DIEKwkEJTT/9ncu/m
hgF3vfYPlD4PkGLpAif62a7w3QjOWegfEDIRVVfRZkKcrIQoiW3MhDSLyt/zZrNYlH4XNwXd1MzC
/h0lVCvARj0lY7gIuHDzsJUqukeNDMI1BFhhM82QKijIkLmClpOYCct86kjTV5NmzOGqDHMdP4E+
0HQD27FRjebxQq6em041eP7UAtcL7uMtvjsmJwjECPiXMTX2CMYbLNxWQA2qmdxCxh1ddow1zGB0
VC7UiFyXFYn99ksUaF+vm8otbPh+FDSag8DZmWLflgwggbgIEg0x9UxGyqR0oOA9JysjSUMiN+i5
D5cL/PJ2QwJUF1rpC4FdPOr0qmrL5OCz5auKnc7T4GDnJrFNbgS1wE3KeMusQwy7C9G6TqJDKKH1
c+4CBWw5SH1geLtuG+QCh/csFOvJfqrLC0j8TG335wwnh9auwzJytKVBzifl4qJ5l2Rd/xaaxy9X
GowK/Kx1iJP0YLvoRhBuL8LWKagl7lKtwkbhxyHtvEZwOxcTaXdplzp4OF+4UOk3K95fQSLBNfM8
4cL2S1ivZ41wZsZhsq/gmp0pQs0XieraHBaQsA2hCVYJCr2hthgzR2oSvp12aOTqMaTyMgv/JE7M
xx9lPs8kEOfMDQ+Uk11BAK6dpRDjNNcIOOkPLRZk1xHADhYeQtPe6EjsHzZURYTkHnCXQVcoyhYD
lyMzXqOooP3EDf2XMs4+FK+9gzd3vB1cb6nwXGrwkYwu6vnuoJHOTb7O/HLLKyAPeIt5n8xOpT6j
V+Od3++8sW8W7nbhscug4gs6r3MwOv0kISQcMNIjq5VpeF4aPBUQjh/ZSaAG3LzhJ8ZFKIQFlyjv
HfY6z2OND7X+G+7fMLIDdQrWa+FZXsmjBJm5g8pfPhBiSl9Ystu0tgubbyVqzd+cGXvKp8iF7IVJ
/wXLjdnwE/tFjpBvaNjZA5ZLXb9WuOzQeWf3rp+PnzHZfgCSEDbNQrKfC99AtG8r/JW+oXDHE1iT
LpqkFu+p0xBo17vKGZsbrs+Yk4uA95npROEyIpQB006NXopd3HM0A6+89+z+yqTUdwIg3Xbq5JyI
p7Ml2ZXRPNpxIzsLFJQ7Z9vvlgiYgG511mZ4JBsI99P2z8a2VJKh0tSem3/rHAtMP4BY446+++cx
LTAcbeyvw/Bo6mtrza0oyJEPu0csV6kw81jWQ15mpx3LUBa4Qz1vZ7tQilSoMV6FVkxHg2c1RUxn
SEK4xAb/JV/I3Pj38j+rMekRMSorKGNYc8haz4Idyq6XFhDINrYhI2sTAta4WrsiiwS9uO+mmim8
AIIBBKq6FoMUn66x8SAVxq7juhPR2VEdjrwGnHc7e+/+4Ve6Pq5Td8lvKnzSe3Op5cj6M5/ZxgmB
judEyYEuMNNUFIYXBWCnRdwX3QPj83Ww4i7AygpH3erKSKp0clIiJEHl6HsrMKqoWL+QjH2meKMc
4bRZATrCZCKjvS0N1lQYqT5xwOwHQ/vZ2XBY2KEK2P/AZzzsImCFrJJdoEOjIicbdOJAaGT+M0J0
h8f0JjpuMXE5dN4xoBYBEEEwnOY2gEySPWR21Ed8VwfnYWLFsdeK0o5JCIVHFSp8za/oGD8Ay63O
Pow7HB3A6ZPeFz+/MCRgRyZzOMrDuI1WQGSoUoDpLTwmKQonzMJPApzzUIV+0IBNvgY3CCtmOp8a
c03z5l6Ir9sDTXf/TsyyQ3+04IZJEsCm2SQZLUdoEXa7xzNUo1zFBU90BZOYyeAV1o5OYN35LdHJ
EQkRRGGPy5JrWSWmqfGqzZftakZShsoaF1ROT5qClHACbDtEvSU1fNJ3eBhbCESYbs2HSkX1lqT/
7b6rmcHAgJM4H7lWc89NaguQpvt35g/m37b/5kX5qu37qFTrGBIA5mvM1KpAn/VgKtekzekjHpVx
hAy1GvcjgIXOBsu+rZe005eoJ45JNAnAwN6Rzx4K1OtPlEVBbP1RJ5TxfPe1ZjKF1Di+aSVyHYyR
2PdNC+yeJ1uk2T99eytso5QU7bIPJPaScYreV13ftMhFFkT453mFW0t7ZjHVVjYW8co7b92fmLbm
ZbVg9A18A4c6xJOmo7vRAozfvAmKeF9HCfpOhn6U7e9coabZMWCQdFKkPbtkSLDyIJrZm6P7OdXU
HvKwNDXKJIb0efIB6meaBbu8JeKOVBEAW9LRbFTNMk4YFB8JMgniLrkhg3l6WgA/NQZ+44+M24Ij
VvFO7avNjMNYpiQC8IUOxIBph2xquSZX3+8z7iScYQ+udMfurU57C3mL2vDSA/+Qd8VYoaeF8aD/
bAInsJTKIXprOxf69W6NQM2GAOWv5p5UowDCNkOunGWhjBMQGUmrv2WC9+D4uejGBS9Y9uCP1ls9
saSWOTf56PwX61GzRioK9bKNXaCvCCswImD4/rLhiDtUt5fyn642YUp1j7HY9N6++MWhWiP9Ga5T
OzjcvKzpMvKeokEaIFtidmmaivvHDb4bC81lhqKPcru+/oq5WXyIvsiZ4ZXZDp0DYXuvfRJEBjFz
aDMCbkr9fxTHECmDzhWpegOSBOZZTIsZ+nmo9BTRkekB/tL6AiLTyvXnWjQPKd96zEMQ6h2XTRi0
VRFigjSVdAVJY1ZPBgpRvbwNM77khRi/U5yl1Hp89wtUwsxQBC+owmaa/IQ/PyhE1vC16lilj593
VhokVE6aSNK2t3YVuqWbGFTg2lUn+GVpW+erfvoquxb9qL8Junx5Sk2Hpg0U8FCKj9nX4J9E/5Tm
5HbA7eUhqEaWIKkdeCN9unmM+lYQ9f8+3BfS9XNlZIT+3l7PBNgZw2wYu6K07niXkivE4lonUMh9
8cd4dEE4zD3ae5G96g+KWIjscr2E7QWHEtbkOiIH4AhZYnZ57rZqGAZ+RlG9AUZd7oxz0d2XKQHl
4hupI+Kahrqj6oN7rP27scapCGJfAhjl2awQgn44bxISdsbjf6UZyKFV20WTXjMFuAuC91Nbk6tk
yTjeBTtCoqd9PB31atn7xpndeCh+OpAz4VbQNm7MFg+5ZNPVGUcCKNVghX+UMsPkh6j+Lr8KMRre
t4Tu1Yi4U3rNbPBiN9YxcvSp5kPJgTkCuokwQMLKcppXxvUEOQdT5myMfnbnNR9NNbD2qr6u6zPa
fqszpH0AayFIB0zNvI1Iro2xfFr2uhy6xFSQVUIY86dH7IZmoKBRzKXrfgzTWUETcH0QL8RBJoaP
+qyn4yiKylUId7lH6c/Sw3vpSJFn0+L9X/M1HrMMdODJmzgClBQn2Df10y0tiA5NXrqfTHD+gcyG
dqhSjVnUcVWsObekVueB4O6fjmf9W1C7iTu0oUM+SvdQTwciVr48GLE1ZDc04ixKoeCEoThel0q0
dIlidxvhAfI9MHWYPOREVJEEWtVaBz50+cW8hl5YTYw2NpK0VKe2UFOqH+qtOkwUYUDGgCva27Pg
FZID0c7rvt+28btw9EpPQaSuDqHSy8QtHnTMR2LbtG0uT9WH8zsd77Dgc3LG7FE3kEMPXFTiEkJp
9WFx/k+SZmJH+OFipLXgUuQjqLl/L/y3xEJaIHpGeUgKZ7SR2/1ftwq/8PZJ8dSq6rf+tYtI2JPF
zFjZ0ybCveTx7Ramwq8tF3wFBsNZybE+wk7bvVYRs52iSDWkwPAKmsiGeyg0pJ30nuqm7dVcLj5C
7gu+3BdDP/4b+Mf//JICyMxQM7mh4MHaSc+oTsGjXsGwXMEyq2QDHWaE85N0lTXkGyybWEqVypnV
VtZLsH0ZoIUCUOjs9hBRDSS04WLWol1X8ytGzVUon+m2oWfYoy/4YwcMv8+MLkkuBq4PWvj3WLM0
mTekmJH7L423aHTsWWRZ4S6yqP79awqN/V/7U/hpzq5FvLyCPBznsTUs6/J3C+t9DgO7F6fDFEKY
XVEMgL1PjKPjF3z9Pdn18M/myC6TzIuR+ZRVt7691r/HWpEQMHloTHyilsL9h915qn55Y0wRcMzv
XShqLfMvuarwwptRn26MkbK97SHxvPDXCH9fih9gG1Mvnbn87YhI/JCvodAfuHvRjGKS2uEZv5zt
bbyXgy+dkinauMcaUJtISJLRlMqvB3KtoU0Ach/mUo0YXdCl66h1e/CqCcWjHu12UOGqtpc6zZsM
E30MM6I1ogAuVJXchcwxQAvMddO/FTiInH9eoScVbzt8HIy6eXRI2MZBd6sGXV2unWBdbLmptp6K
vt4TQrrJ6chpvSaOGD98PaPZENRZgt3rE9xo3lt12DEF0R1TrMEmS1+i59cPZ/B9haP7PEjHms5E
s2G+wdZE0iq9OcGzzAPN+Fns4n9ocI3WwmIzfCXWgALtqhPdIcwH3sdTingEkbGIykGegbI/0iXE
EeGvsRDSTWBA/tes77J07SoRLtuU0ULFlRrmrMoTJj60vNsyz5JBoAcxLvENDdO1AwMr2aZRG5js
8dy/vGJ6fUPoy9tafA7hr9wYjDtIeYc357FSQVWuSQDex84WJkI+jFbW4vw3peaCG58gaHiGUwlE
NSvXOr+MwSnYQQqEgKx3KB9HknNemWOltfBiPsiufZp6gcCnhkYxF+Nf7cD9QjKgn4xzwambps4y
39j48idSnHhiGWtrzULeQv1/1nGWQFrrOoQWife1qidCyfxZuIbX7ZmB3gzLM4ipNXbsQE0ubL8A
8rwKbHYT/I6pl6fAL445U+ak/gslrPr6dL9SqeA/Nw+zNeqIHU0pWLlhloxqh2rH5TZr/yvo8uji
0fDxZy22qb0e0SQmGOXa76hgmFxJ6DSWDv4GL57/jU3eHYGthgjgYTlTeTf+GdSK/CDjYwBfpvyV
/FtA2J8dNsH0lKo9NmVfAPg8y++67Y/adB/WZ30OiCbtbyX7fUxdUYS0lRdqTqTyb9gdg2mMppx6
oiipdSdgWdXaiQ6MVVYUNfCbH6jMBj0OeW91JB3wVXCzEg2ad1IQbq4m6IQP6s5L1T4DeLFI/NMl
0/BA4nFsK0NsYYMQQ59NQ/pqlSPH8EWy0ZmeewUXcWhEIsO0jwPVnGSguQyConfMMlKkpdl9JnJY
vccelumVp/7L8xpaxWYKuqScEH1qTGi+bgntbsfSOSE4mUo716OfNvIRyUXoGICgffmXQiU6YE7D
7L4r/+TRuJTdS/axNcacTWWpoXC/LcdogzI0iyZbYO0nGqHTvs1aarnSlafmDvDTruKCIFkUXhXO
sYcQP9Y7QU8cKOD3JE5MimQ8bFv0uMvo2NwTi4guUVDwYQGRVFWTccUOadpDS5aMSxuHkE6bIkSu
Ix76uOaQniC4adohfOZuf1fdmQaAXTDjqw2+S/P7ZTPJCX9IDs67CZgmMX3BkPZ0/ejmAl/cMMY9
qzevjMzKDbyjDKDA+Bni1iFDPTljrBTXt9wJKUOcSF0H+Cyaap4zDZrQzipBGmJ9j0UTm4UHxQCD
tJkUFJhqPr88JF3zbRHmVBmMOoKMALK9SzD2eFVuX+DdlJ7N4aauwzEIR4/tENiFlj3BBG5Ws21j
TMIlH0G+PjIMFeW1jPIsJRHDwHUt2q2c0N/2bBNKeFW66J7sDaos7GMloCmQ9yUyr9ziCiBGTfRJ
jUekFysveSLH7URAFJwruNE8vjSRo1YkuSjI05HaB6/CQ2HVzolyKJBTj2FLIXxueJjUtLfGnPu7
PPWnraZBJdx5p2mHK1sQSk1MiPx0tP01/Ak7b6oQmOZml2nPpqPKfmTSa2QqHIzXDFXqH6E2ePHN
oZV0Wi/wH+iGCiIGwMVUC48gi7fpg/rWVX2QjAzL1tFaYOrEratwl3uAU1ORv1yWJQDXPPxQo4wc
jNcaYDZFYQRGdSwHnstgE95ZWm7cm8n2otELAsl7Vs3bujnrLC7t0Mz4taQWXUZMkc5OWdiT9dKj
RLk5MZK40t+Kn8FI6AkXOAtUAobCgzMXj+9YffKW9xhzuWxYg33ilMicY5GqumO6/l/MVV7NsJav
4LTqPaqOYeaxrvZllL2OFMqtuoRRVsXeAPx+MvTCu1qTCXdTdlkdi7QyufDdEUJfTxgiJcKPlbAX
QkWWh6gMEkzh8B6s+I/wB0M2BmJJuw6Xxp9tiZxwOjg3PcbXtZvRDTYGDlhdLCGBcjtgbbL4ZtWP
qSRZCdQ0En1uwktbyB/kXbfvjctHl4iA0SYzMx/NVGuxIXSymYBjYUd1HUhdV8wuDHPh22NvgWFu
VCMsbu9V4AE/ebepl3GdHQjRMlbcDWe7ebUI+MLVHJh+EAKRifjr3QAhn7r9qJtSse/f0W2EN7Lc
mrBSS9uOaocRDq8ANnyhxBvz3dEd9fSS3LoIOr8wl3UJ/f4ruZ71Lhcus7OB5KiRsl/D5BulFETE
jI1dh5ieTNXinVm2aPR2l9PZIi6oUi8xKgpRmTTJKO7Y5Ej9dKCLCzoZBXNBVILnHBI27LnknVjE
BZGpZwWqKAqsapp2jYEyZQTxv5dxkS1bhNduWTIe0uXS99euY1ywV8YjEM0PhSCDpr6dJycW87Tt
qcQeQ0GPjmrBWeCzk3/OsSkKjf7x/oZGpX3vy1Srna1IEY4FgPntYNR54JD2gYJRMXD05GHFYTBE
BLGVNUzznJKwQj/SMI8NCfcvzczm0XJVZU0GAU0+bJ98eK6zKr8FkLnR5m1GrRt1BbngWpBuK7zP
SG8yqCn3yqlXZQXf6PMsM5gBkr32tdWp5gRzh0NknZBNyG1rz4Y0lVOwq7yhuGL9xDhsR9BVckQS
iIymbBxpS6edcLQ7e8eAPVI9tkvwBKGL14MKrVT5qF88TEH79uVUiLxJRfxUK+kMk6gADtX5SHT8
yROMlpSxhE439SDJAbRVcu4642u5UXbKVXTovxjgMuNZD+nwfzDKt6nWeVlx5VqIKKF60ETrTg6r
1K+wKrh5QEhvDPeYxwknXethnVq20Jcuyw6C9TMvbGO77PUSEwVoKscRt4iuuFB2VRwBBBRwLVg1
OxiVyK7BuZsfIjn6x2RPYjdkJD/o2//ObZ5XzD5oeRXQFXBIxeeCspdxsW2jnF2UHCX8O6bWA59I
hffklLZGUYGPp6z8AWH7/MsxtKkShFTpHjlrF1ZeChkiJ9D6Fe9dEeeioh+z1sczXHRHjotKJmvv
nEIbxFYbBNSOXQsy8Hb2lWj962Qa5pbGi9Oh8eiSiWYPTdc5J3qfvHfTUIobdfFUOFKQCGRpjHka
QgZnnWpgdd6pGznSuLVg5XP9olBxlL0QIZsjAzMOrfMULd88XsMkOpQSvAF30ddx89zsWbE4EVEG
ubyj2EHkY8FgX8K0IrxUfcgV5Vjyyh3dowfm6Y1GeQL6eqG+omsXkGwVVhRzsl5bPnRby90Rn39E
B/FoydxxJj8rcUSLqp3D6krKnH84UodIchDylvgzcEzQa8vXaSmd8cE6XXMHdCbF8wt91a+qB+Xr
naY8RpNxaXPZsyXXkgioLMRiuuu7vSG8ebjuGbtgS9Sy3+6kBLN8pS3rTLcDHrDHX7hZtihtTbvT
sEHqvxdnlz6wm6f/6QKT2hSwRRrjONbGt3Fa0EYrwusEfnWyMu6d6MezxCNaEsiN0tLp4A7WtKql
gJDSAOgqBdIRbbFfOOGJa3VWoRtkAKLIZ8ZDf2sqQGNtNcHbiWTC4EzmrXGF8LPe337tvZpN2/2C
sXt8T0RXnR8RAgF0OBilCrjrAg/dv3C6shnRTavRuKQwGgMX1PATzKO2xBtGN6CQoWLYGeJg8AIC
F0B1qNGLXkeGy+S5OAUHLHgNVKV0DdvyCZph8UTa8ax9FCfZcsInilIO2pM1y1UGJFRVv2/4QVW+
c8IfYf8qbtmRzxXoCHO8VImBUHdOzqdUrs8m66idnu6oSRtFmYKjWBRcSIM13YpD1gEM+xWTs5/5
lt/DCy2l8xyjZ41YxU7VzQwxe3v6tYZPIe1bJXjX4Ja8svNbTXA8NA8BYplboIIploKd02LGaKbg
EcVk5kyYHGF/hHWPyqOUZl9yWb+rf29w8S6syncJmdPSAiVpzsY6TiGCdG3EmIBYllkwwiz1L2Th
J4c2ID0OPFE1VOggWtiDjGpNR7zyRPk2INXIoxn2D/oSRo45WqNJ9W9fqhj88YVrBZHc9G3dXAND
ZQ7wG6S6QQKBaRFOHiamJYbF0JdqSYcwJUpEWAATzeJHfll57E9dVUnU5BFA8uOgYAKIww3ZGnRf
jwBOz/A3v6M79pHekXUzV3y2p4Uhio8+3pNVyyyskjV0BlPZz4rWkgmZWzvpJs6//GYvOqWRvfSK
k6hWg83WDnosBQotecaVIVPVLj8rrL9YURzHB+9A7hJbLNZhBk2jaPuCjZJPDHAXtnbmo0hC+X1D
J5Knd2ytFBUtgRG4W1rWlsZIAK6QdUz5agAKzxjsuU6YvH/t/r9fmMDBKnZWuO6gV6droC5P8lwh
lwgvmYc60ImL3Y4zhuion94aeZqXigOI812v6vGzQk1WHCBiLuqLETltXSZmX0ZW6jX3PYmrtDan
AUqhlXa+Efbkv4XTpjMQKOhBS0Q8wRr9knO89zUIgMTG+NsMDN7DNZhoJflVkAG9n0yG0akxPvlb
2giCI727CgygY071efFKKv9qUGIrY4FcUMtXM+NOsKiuDxtSFmemo+jbI0fC1wdHHl/2vfuD6zlU
RADE46xvZWJVPWOdO9APW+1bdKGokcDvpMCxNP2KQ63PZTv6ImbLlMwS8pvTzNmSt8YhCtxCp6jT
WJDFaqAK1xHD1faFlkBmIOIBKKNJ0c4rKrfrsjHDWJzmvFUlDQY4zoPfQcZP/ZU2PkReJSktjQI8
yp2/LTlvSoNNYjriTYqo25z6j1eH3tXCr9m5FZXpD/31VOH23OP2BWgkjc38mg5+sPem1D7hz4FL
5uIvqOGIYsSqViMAsUtj/bZ8H6VLsNPTf1p4lqSAVTqapaIV5C8rT23sRaDAr/4kvdZxoTPBaMyQ
YCAlXPLdmZbL5CBCeWV6cdDGiQChDiZwk0zX32VhwCdhcTxxmgJfLmBCspXSJUHk9XjeD4K76qfa
BjzG209W37yeDBjqg4enEdjKPzy3Fmz29Hgv/MBIWmNj/lVqws3id+tctjVfm0N/NLPfWd7RjwW0
KH9qmOWYrR4ZRDcnsRi/6MMos6ofc7h6btsVZJY+P8/p9PrAXdxjTlybNwr/gSD2w6m0sEAVkt9j
z8vHdMQaDzcfRTPwE6B9c8wapbPtGa7l3GaFyhmSf3M+NRApp8SD7u2SKpM8ihgikop3dF/mklR6
c8rNUATuuvjkA2ysUwyImLBcNB1NoAu2EidpfVaUrDng1mUokY78JyuhMSXAq4/KIcu4Cbq5ZJp3
5iVOYJ1DXgMYYKLg2YwF7JhJRxP/boraFME26tltxKUCboscCMA0cttd/NYyMW5sbtnzeqUdvpZ2
xV7rHQpW7VvSaS7az8tZsnQXJs6j+K1GgX128ZQA517PZpfh0uWS/1l2KEcpLKxceOWmzIDqC74V
ij4ci7+0g6Mt2ZX5Hg4YYIEbXZGXH2/wjbAzXpeb534YkwdXsV2+R2nFK4T/X4QiubeNuhPQiZcM
iWV6FcwHJxo8Vgxy3uQjhs1Ifqxmf8VvVeDDx5lV5ew8y0CMb14ewyWj7o4Ph9Oe6smceFiiCqVZ
wg6BymPh6JJp8il6UjDFkDqSjqg1ZlWNZYHRtvc1vE9Vq5BvFtrRxzeb664uitwYECqVYVFxJF4v
Izolkan7gC9TjNodxOK+wWBpWHTL8N1xkHn9LNbYfH1dg3xzoeeFb82l/7DQvQIkpZLHGKIWKAo2
luTHXJCNm+5AqyjmwJB1uor46c+sUYlzskKIAQYWwVuk1HXFztAkmwlFdbwh0J9DCUuaiXaiqaY/
K/OZMv2GfmnXAUfOVPKcA/OnxuJyqvsoHG+BtwfcBLQcLZTEw00IiskGtcfVM+iMJ7OONHyo+adq
ZPJiNulh2IFU94ZRuIm0N0vfzLh2r9SjgArVdZ8r05ZzMU2heWoswjqtnWft3+eCyLiOU4RMcmCC
3iDFS5YdNlcZD8Dy6cfMuBbosOPP3wI4Z3r2ubjOmiDiTxDUQeTkaSlgh6x3nwgnE3CaEG9SY4YW
yhjAPsJ2+X58WIyGejbsfQl14G79c8hSABoV+eDWT3XxGfJRtwRVT4OkCzxulXNs76UyBhpmWJu4
8NbNbFfLPxyA5CPc6NMMbuZhxVYMkM9kjEzOE9qXbKi1WrozBhlu8M4Eu7tI0/T+pCYG5U706auq
/CnBLz0wyQTrqw0TizuvUdWKmTpu1vyRcqRx8pfXzACE5FjeOaAgtbKFvUpeeuNlAN/ic15RYhKX
o6wBXXUwJbdxvQFVcQN3aDXWEbtVtkyhn4lKexYhe39X3V07ZTNSyVJnDKKywSx9UFf/JwQQybp6
b5BzDm2y0vAcXnxXk7jeyLEDoulXcJ7pEjFCeaqOZ2DuBJJEdt0ehTrHm37lKXFmUYneXiA4/wgT
DIKu+fBUrVd1oqVfQ06kw87OSsG8hLnKJKQCcu7B5o+yp/FpKi9YgyGc9iqjO5Xx9CsnUFDkxlnw
paeLm2i2sZbSN2vofZdBcwHvMftZqM4X4J9J1pfGHfTZbXJXk5WkrfcE5F/Xtf8cgCHsP/3eVWJa
FqNkK705dYUZ4kUk2FBU6khwniiTwKG6Y6BWWxNysN9sMo2keaaJJwPIJlnArkx0eqKjeNS4MuHL
BrqWMo3lYRJ3f1MIHboSt5WUvplOrtSTai3SJkVcuINVu+Y+hjrtMR1Y+Ww5bElfW9RkboOSt2me
GuYAsIgYZJ0cL4UfF80zvk9hG8SDDD9UmGLGAgphXMrzs6ZF9I74Cb6rl6nbU1GrgFVzfkYVM8Ft
EU601GDVzu1Uby8kJJUV2Vgpjb1bT6+/EcfF1dnBLTCMsr3ekKiV5iIQYK8NiJPSafzO2ZzS1nuR
tUZgrBtcxXd5nSnG3Sue1c62oe1ZodA8Kvi3Q1UqEwxLTv1wPOu+LEch63dtLQb2NHpbNmPj+tkl
5iwZsAxl3XZhSkAghcovlBclv5Tzpz6+4bcY/Mw09rnLWDfjXsmMQUSV6RB5r4ZpkXUIK9FNBHAR
V3Hb2U5TnBmcDmMBTF1Ag8DGNp4NXWCY9jxh47QO8pqBkMEEVgIi0knUBXEzwKWBJDjHWAZjk7vg
lriT2TaVyYy9yXTjorTnj1Fx1kJvWRiLNwrxYyYW4daaYYj3gVse5RlD68v+gtk2FB1Cu+V70EVv
84cFCX+t8DrwpgUv5eJG+nF6svMDvNEezYYF1uL4kr1l62qbdACcfpVvJfCoRSh16+ZcKTttg9Wg
8Eo/wP9Ku7Kkpgd0mWx5oKjBIaqfP5jp8JdNA1kIMeEp4NeVFrofzFYLHZnLiQ380m5PXPp3k54W
34VPZPGm3T1V0ECkfLgGMVwGxk9rTXQEZ8zaCDb0yXrVEyVbqb5NAoEximeltdeZuS05TXyPHgkN
OMcZqtgLFqvm2bBmL5sOQbj96UQ0BcmxfpVFtS9UTWkRSUOWtIChv8+bTjzck0rvDgjRv35u/uCM
eEnnusH3PLsPJHRO9DlQGKAZUB9Lzjmh3KMJuD4uBjCzsz16urwTmhct2NBN2xVA+xmCQVhS6xZz
HOKOTG7Ub/m6+1GdELKYXbP0HpaUuhCIGdEP+un+8ftsgztXExpq/5TjmFUg24GZMQhUdEIvd+mP
brAZysel3lfAocGpLGyaxS4+WaUenbG17v1cnksCNv8fDYrwm8C8zfUJDvldntzZeYXV25++2bUL
BcSCM3MbeBqNOFqc6BSr561FI4jrxbJu1raiqaCS+6xa8HKo8pCGjQ+LHJjg7t+h0038vDrf0QF2
zr8Wft1V0kNJ8HwT5WO7sx/sTtmb5rgsOayv1p7/t/DlEFMhnch9bEk3Y8+XhgMTUwZcWxCaJPRU
ONS5PBKfANBkq3GRymU6b0ULMAKZjDe6ifo6HCgKtr7KZ6OijKme91Ir6Eeg7hm5xs8BjEamIRDS
xJRxZ0X7dzUnfLsRvatE820G0+YcVHbii6hP3yZAu70IGNfd/owDTUSIIWbU7NjUxobKZ4LJNN3H
rol20dleUKCLzUuapUBV+k+ygMHzo1PmjmJJkaRuujkarOubN+5zaR2Ri62ii6+QP/5iI6JVcmxi
Zafy70RwoG+fhW+YCuS6MNuEk3ptfo+1kA7UVmghlyk+C7LbWpbwJs1wls0mjPXHpSQRS/RPhY0D
Rvozh8JbLziaV69/F9CE9ZN9vXvyAHTTrXCPK7i4V0x7taV6JaXnSWhdorBSJOomZ+ehojFeyTtS
TBnmrg7ddHqZC6HLzp935MSqele4nTuBVmQPktlrMLqWzjUVeeBXY5XWacLfp144hVRUgL0P5lo8
FCld4kKrI4bzQ2MqDDT3rvy4Q+rO9+V2Ar+n8Ra+hbNjrfGh6WG+c303n5nR0Rp0441CTqzUL15i
yKcoTu30T1Hir6ZiS7pkeeKxvIpWum3Bl4+198vCxjg17Hpr7fv9+xWjCwJFEzHSrphmShB5e3t4
K2D2n8bD4444E89KhmIb6hrnUMzmWZKHkq7VaCcCTYtxXwLEzO5C+hE6D4zovJ+tNVVainzkYcLv
nVyv28jg1yOC0UmN5Va3ZzNsn80RFEKiujeSx1Sgq1x0iWKH/kY/tf3+BsEelREohToClQeA+cUY
YC9Fo/rUJFzwNIgJqpVQo8IOFE7R9ngMa6Gko+qhYE4cyuTdZk0YW/rPAvHZrvH71F0EYf4rh/1P
7qdKWC5PI7E6R2VeF6lhPDJV5XmTsjv4MCSsV/lNhv8xOQRVx+QUliiXIDukH5JyAe2zf2zLLVw9
NEis/7J8IXcMVBrPLGSrJ+jJ93L1IbQsx5Gr/j9MxsTntmqwk+yxqf6c43GXq3fTYGjnoS6dZdUB
Y8Fj9+kmryuiUPiCiY3TQaaZIhu7lO5/Fl0sV7c5RG79QWE4S+59gShK6b1MsNSnhkXOBv170H2H
E/vt5R532Bi/bhfl9KelQQIwktkJhPZ437ka3MaZJ6j0De5wG/WGKvcOfe+qJipNY4ZPvQCL+T96
rocJ3nQNa7/EBnHqBj2gqjEGjhsSEzGweZJNoJbKeW5vpEyknoM5lkFVTflFzBjQau426pTwCN1z
qIKtnhZ04Ty7uMGX1CEIpp7w319FP7uRyfZulZC/5BUtEnBlPLGMPF8aewL/YLKvtLnoKNodc7L/
6cVL9gkezgHgJGTZPxX6WDDnd579lE+OESBWsgxtr/HOPT5k+k+yGrvyrET3d9Nr/XDIm+gXDkRI
LkkNTjdrIWr1KRwP6tNAy1iI5W5cmrOQ1fIJFBWnZNbXdNkhJQu06KiXPgG6rlyCpPsLf3qeqQ5Q
bqI//ATpStuWp3C7qvfAWm6c3DtpgsX1i+FtbxYt3n4ZVmZvUd8P9HznuxTT0lVND7j//b4v4Cv/
XqmZTPx6V6By6lfVard5ygKB9BXd6ezcWmR1e1IwDGdvtYGjtvPltsfVVlrwxKE4VqPn5ME3eup1
wxXPxD93TgaFrtCTj23LGYSLStV8JyJTHdGy4D9i5jKDHb9Evq51T52dD3ySva/seo1io6CFbWJb
t+9Euynlx7HAEo1QJV8I8njAKYiS8xIicblKRc5jGc1IkVzWzjSquwzB/UZ2HE7zujj0LRj++IFb
TnL3zi1538gKdklGwzRuotkYmp4J4DhW0mcWo7EEseXRjXHRK/wBsqSbMh0Z5HYhBOd+mZbIHOFN
kovhIXA5HcQ/8hgfvQ8Nv+Xaw456gqw3cuaV5YqZxkQyPnrX7zUg1WbOZWVnBeXWxFuJJb+InYfi
S2jVhon5H3K+72D28+92dTWIBUxYDq16x6wsqn/u4ZnCjO35cs4ZkBEn1tigU4FiwLMQkhkDEkql
XtBjcCjUaMYUle78LHHnf5Qb8qiTy3PqeZIutowhTQlQoHRgLKuh+ejAt8rKlHnCOJSZl6s5Y9wS
Yr69LUJmqMcHw6ycJaW9JSXbOa+1V1ErZRBUFNlIVFQ0LzSTLkpFPHwPdoWCTFAHvVvwBiBGRf7Y
3+v3p4uwV8OtwnJUEcTDmxdUwa5vEPmI9n1SXhfLjRanpBWqJtdptivrsdUopEQ5tENI2YfpSPgk
kwG7tz+1KZQSzY15tZVOaciSZ5I8xE0sLCgTa4yJASAiqltXbeoFI9GbvdXSgt9GyXG+ViMqC1XK
DrR+7qGUsDVADC9Z7EjgR5B39gBk43P0zhaqnUGR4Yrdp1gO1BTsoypQlUBInFU7N/dqxoLmaM1Z
7Iy5awDkxS4kVbQJPO668Vo3ieoDeYmySk/Lr0sR6tQe3jW6sa9i9Zbo2imjI9/pUVzE770kg+2G
u1J7znG/tmlGpfTBezDWeIdw60l60jmUPO8zKjfVJp1CWquAI7Da2vkdtVvR20C1aTmbtO5RTNfb
T/FmWpLlMTmaknPeVYeTiSDFhSGx5TzMNwtGmtu0x7j8LliUC3vtsl5Hjm+MNaDaZqV+yA6bL1oj
bVbpBQpnv7bIEdpiConHr6MZVdlVioVWLQ89MRqx6k8chsiZuKf08ud2aI1lhKIsCyePBgrx8bTF
J9LEhgbNnhpAQFWTwg3SM5h5nL59MZBX4IxHucsAacCxCyOXp+acmGUYUY7g+UeITlFMEIiKSWKb
RKcZcFl0EFDi3+kTr6YXADrQ7lXHbU4CN7g8R69wGMu4gLZgKVnnxXip3QYf/lebY/yC48qD7nEp
sQP/Vxnc/IAh5e+/6xW0ZjRzNHfYCc7TSAxa4Sf8fi3eg0NoTHxP7RnBCByoxob9oB6Hc4F6cf27
DkYB1j1hHhRO/Q1VKtk8uPBgB0GaUGDSt1IqgLnx6Kw9RnLVlmeXrbiamZ6eEFaRLvx1YrQFg7rI
fRgdFi0v38ti+XZYYAvuXSjalx90Iq57QLx7F0sADDtcjw3+rOY8QCnTu2LCEHY10FPx+1fvS0Kk
Z047YiFOQLEXP+fs0lzcYQFR17lb2lXFkitoxncq2RBV2zG/kJYpH9kR6pxb5tUnxL6WpdcRh05t
WZBj1+TLkQ6KCdsnqs/wGdfrjK/pCEW+oNiWTyKKu9TLxVIJRAsDL8hfLfv2tQaoC5dvd6AaDIYp
VV9H6wDop68hpfkTyO4XTnMu4djL9Rs78Fm235LL6zvVGCr04lSK+pLTuFrDFg/H3JqLCy061sGD
BqJEcA4uoF27v4hwnoEHc+PjtkQ1pU6MXN8dyhwO23SnVmM2RStn0HGbmk8RBaghbSpriZ5vlTwY
RHjO+H/AKNadaaNx8OlyUdM9dVacPnyIiTQvApL3nKX0pHM4KDXSm+662nZgn0vcoKK4oKZCS3sr
UXVLfQH54qT3F/DJaHfIP/3TUMBzTtCeLnTHVgZRLm34nj+I+SmhWx2MvPnjOge6fDyliUpRfjc+
Uf4ZwbYW47/EIJyxEsGx0mtTEgDgeBAh2tTYjjSsE5NNCoxbGjNaXCBPO37VO/Kjfh++Seinjv2F
9Zxc5mZ0oR7ULTlZB+LAeN5l6oqUvb5Ej40xWJ3deNdpq++wv0cCfQYhqOLCYDdLT5e8QQE9JBI/
7Gb4dezYTog59VX1P/9SlpBHdkU+tr/24ekMIO7QmXQgHz0VN4Qbif7FH4omxTC5c1+vCE/J2BVG
g16mouDJ91RzkIf6/XKL4FVlqFWNr8bGeEQskGGNnNjkvI7VeTQX5+Ky4CMBz7fpgTIb0Z7K6dY0
xxchUeN3RvKbnhtd3KTUivMN/K7mALksGOzR3kklODN7NCG61RiE/Zicp7FHqxs412LfguW0KaOi
1El0LD7G4aCir0njbxiAyvKLU8/SNXVt2Bsm6AOKiyHdUH7O0kSSp6zWbkuZ+Wp+seZKnITauHYf
SCWOZW2E7yepnJCgYndYAfY/0q8PBKBS7tIWh6YTy/ZmcdRKq8gUuCH94tOVDOHoiVXMg7GXVzuv
in5RRKPU9Ue8BekNJsLwzcL14TpRLnQQzipf9R+3l9Mlk7xZpMunl4x4BfjrAcLKM0O7bP5y7FSe
vFHzi1xKTDzI4cpLgtk/FM2zSqJ/reCa01oShnVNjrYWIcQrQ7LDc4S4b6FLTHEttAGGlFtMDz31
edncE3AdMyjNR1H3YVESo85y/col6nEm4YDJfKYveXi1RGlIWk9nCeGa+oA4/HzvVvctt2f28qVB
qj+8fBEMLf+FBtPCzNmzw6d139LqihgMlalM121MCjXfNb9fUTKW+xu3Ss22sxLyQ4oi/Ygnq0zN
SBj2F73k8FC4I/gZ6wufu8+Rt5Oi+CmcclnLDDpkBS8dvfnZyaXUtQRolJBDrd6NkrYZlT2NgqhM
uStDKsRogPndRvmspFjnDFNTSE/cub0dvxJs0VqLKQ3LuhZLDIQ2G/UDo0MLKw6hDJOe04luTbwn
qUasI16NX/MKVVkITN/gikB0KYAExYhZjW/GDpDYiI5lXKZzf3bWJJH5A7vBvskqYmcWJAZuBGuv
K2lXnj0oSUscc/scjCULZ/wv3Kn7kOaOj5q/EvtF433874Hy9gW4SS/NP81dmjcKlxNLqiQbWmWu
C35CdSOF8sKsBe8QOqAP5MgVw+5Ny4x7Tf0vlSVClp88rM9SWSZ3lyn1A+CG/0wQ14NJWl0X9kTA
neM0DnFVgmsNCInOTD64ogdSkZz2ZVfR5CsA3x6+KNi6bp7skpCYL6PBtAwi0wE/x6P51xIyrqMH
leV20fT6ETLcuGb9++1Sq+sgCu+Ghd0/ezFXSPxcdujQoHWCPXaqNtCKfVbCI0lXRsAHyYDFKaf1
XTpd/a+Cmp2KCgZv8X0/1aJ4XIMl/TDVMyrTZbDWajeUBW98SgVvTDVFfZoHNLmm883sX6XTSPB6
k1/tfow68CLtQjgSAmifqXt0A0NVOVb3ojCbISF3irJzEV+iiufLWWEnOf9mWMwuvODn7Rybzoxb
HFf8FVkQguyVnyYOtcbaXj+HeIgucXKMiLdgBMI8YNaj+cTJ6kcbi83Sg4fUItajdfd/t7xkUXmu
vDgNaA6GcCpW6Xd0Ugq168cyti2BmG0UmWV27C0s/amd88bO6VmO+7uk19yegwGPWy3PctW1PlER
tnKCIzm0WgNDbNzyz6jhkEWSuUcu8NYtFW9VMFbE4OQFk0TMosN/YD/W8ZE3tVuID2s5Iz+gnAZt
gGgOUaXh0gmsBpQySsdDqaoXYlEVQCAfujGCmiZH9WNrcOoE9ZJFpSGboAeYZPi9AYaoPag1uloP
griGnl6xNjzMQny68IUusOwrlLZ2EWzVmIioai47STDm2OrnBO+nnAPaza+Q/KTA9b8yY1I9fRmd
B+8RPwLEHmAGw+tyb3oqq3ROsfQIz1R07T3wd2TUZtXZ/TjQM2yUM8T+RNqiAZSekLVW26x4OFCQ
FxGBlfYu7vmDHVbIiRP9yvS8wEOzYrY9iZg9oxD2R1XW/cVLAEPekNVNgjNEO5q+FCJYFtij4NZI
Sn+zhS6JmU/itYQf76DLrydqtQfKo2VupLZ3lzx+MIw26p56akMbnGyFkEnjc7qxxOGD24g6XsaK
7lDhmyvkBU/p0huA9e6FloejsNz6PlQ3CIHf+zMY0Xk5c4eH8eQnSy7kgF4YwbtWUJ+D6dCAH8IL
EXi/vi8qgBt7ePyksPHyP4s3Ao01cH6gsSWOmWLXNI0ElK6jtLgqtkFP3T1cqzfbUuMyRtedzgxg
eP89bNhfX+bRNhr1XPqUh7TsdkFgyMbaeCkyFiChy0C3aCotr0yCLpNpbuputzw5B+BC1t8n5l7g
G81alcwlZD9O4sVmQkyomb+NzKWw5KRfjz4QFUNoM5YI3xHdclWa/HXS7TAd5/rS0UQB3912dyws
uEtbyzkEWHzBwGYlBkPn7uqXjW49vrLUpiBffcESrWolZP3IwRGBavgZ1vdxhj4hh7cmuZqd4EUk
9KQZKb4lSEC23AQ900+3suxvL/E1YkmbEuqK+tDBLoYdPGXog9LnCMTJP5UVPgNEdvg55EXTBDLm
PYT8oJ9MPdj93LhGnr/YcYVDfqvRBAxVqySkgtKmKcwwyN06MIzXtra35hMKPUG6dJH/dvqYnooW
SUSclA3nSBKTEdI0IzjG6/EtCNeEBZuhwCWRfB+dsiVKpzfjASO31iy0QPt/799Dn/Cx3eaJcemj
edat1LpNvrcdtHE6nCJ/mrin2qZEyx0o1AB2ETKM/V5ndAellpd9rdHPXfBsN3A0m6fZ2qM38xyT
gUhonKAvZuBIeEHLbNGQErHpJzHsCs3oyangk6Zl02ZqAzm4ITql4PpqzCSSVyMn/NgjfINIpqrf
c0LTAOaS4hWabwEJf20P3/WJJxcQ1COeejnw3235Dv3pDXemwNKg0hXHh8hI48ymY6XepcSk93Sj
WhYJeX8UEt+W9NGsFzO58nWfd0ed4kzM44T5DgJEGjQhAWfCj0QiHfXFp5RqP4gTQX+w4MyrjfR4
57pHdPb1zGGjJI+IQe9M+kMx9IkJE2zzuEo5JHWDRwTyzW4qY261QrU9hl8qBF4tOr9iRiehSfsS
z+Dvr/rEeirUQL12okRi2arLglEFiPNNYbJxiNkVjBrSVTdk/+X3Txorv6VtIsan1h9TFXn4cq/O
rGpa/aRZ7Z74RTux4rmyX4xRDLAKFTtmsL3weEJObZ+ZG8oty+ZBTf040vAzn5x7M/HO/+I20JFz
e5CS5OL70BIk6+Y0YMC9RYjfVcU/Op8xzkCVQGolGP0XnFIfRoEY0U8WHZfXScAyX8h8+lNYEvP9
dshGpExVE62oEuEQiDhDZ6vprqdveTK/53H5R48j37/WKJp2I7P4GrhlWGtdUImsRLUjDXUDvm66
K1tejGQrSWYsqpbkHIpwH1zvlvSXG5mvrJXI171mEc08kul3gQPeuS//p9JtUBGiQnM3Ej8S8fQp
8yiwhyl9sM0CkJECuXo/n5mliXwKJ8QwQAKN6+RKSx4efc631CVvM0u/0CTyaLb0MNUBIexd/Ec/
J7hraq+wqLBUjlboPa96M9S5pedRrUOpJyKbciCABV4AxCN1IYfDZioxQP2sLjpJxeTP/lHCuC3c
4KmgqwZnm8M22bkUY1igVgXt1VOUjGX462VutxJe/1LgdFJS46+za0to/aJm1o2bkqV/+inSM5j6
XknD1j/svB1l6OhMkSK8bImLGsekL9/KJXCHvPkxWRQSRm1EhV34TcDTg1g8cYyI3VmY1zk3Abs8
59yIBRkMQqFV5qa5qLtBaWyv3VE99gQh8XHx4gcYiAKf6I9sStOPqltzhwRmGzbszs3YNkao8yuQ
TPakDY1KbLQnvRTkIB6cIyNPfwQE4klrvhfRgOnAkon1GtofOkfSJGqIOjpAH2/aRV5chTD0z/rm
pxKgdnTIVMuWzG6EPkYK1ybCFMXZpeCOizNnGwalXpM5+Lu/y8akIL37dlrzhccLq/Q6nkf356FH
g2FMO4FT4KTfE6zWoAE6OlEV8o2jfggyhTwSMgjyUjCW2TDOZ7bm0bod+5XzCdJ+1x0N5XWb712d
lBQkmm5Zq5KH2fQe/ysPlkLLwdieRS0NfNBrdsOaeDRn0cWupPmmMizHfJfj9uQMigbMVYzBIpe4
pyoJE9HfgxDYIrFjvDaR9jRipKqPyhN7M/vhGvTE8GC5JpYzre5Fuu4s+fxDMSzurjGa/0vlwMl1
MSfZOILm/I7A7mmmIdZZPpOuRLubx8nrMn/+jOW5NiHMNHdlUE6HjazMU2XKWHfzjGdxtZOcZbs5
z86KYZ2G01pOvD64kQW1dqYX/OELqDOGfvOp252juMm2zbeSTpcdHHf99tGxlUJPBLAQmHKCtJQV
CUFAC4EP1cbtLaft7PtBHvtKxub/PUPJ1lz7ny1xBxPpgG0Y+785HiKAJhK7ObCVs63uie9KZpN8
1bbdVP1/mE5z1RqXX25uYFAS9HP3YE09TTZA9/b2t0np6BmdYmDJcpbLshMGAlVsIZQV91nDG2QB
QqI/vYwxQuELgTjvYJp+AowXy+VMsvz26nPoG2bvV4adKQf/q+cL0ULa36eTYvscRPxH2eeMeqik
WsS1I2dJ62xZyvsvkymCkhfV2H4oc/o0+RyIeEmHSW15DDDkl+gdYwW+CeBBY2DE34OYTF5RLqoH
cHw/MjZJnBYNxmu3hNexdv9Abj/TreWdnUjA1U+zacAmmHpxXoi3zYUrRUyUVF9CMBqgGoLc/dtb
/pvD6GuO/KX3vHR+qnDw6OGLQ+8HlctcsGPh6Mg/gplJoY5PqL6N9PHi/BLFDflh/KhwHGiAiPNk
O24ARnsGIfMyY2gOv+qlhROeZlvWriVIVYnx+hmB0nKu5tkKAjT0+veGKiDplDn7n92sIMfXztr/
J/oucpJD+4raO6ppiBck+i5d7hMhfr7sqJIT3bD7DmmDHnag0qtxOAokNrnJC8yUMJ0/yS5bxIQU
rwS3HhjqPjT4QCDrvMM5nmlVlESCcsPzYm0tejx6mc+oK6xVp1tWAfDaE2/D+FAUwBYXxLdWISxQ
6uceT8VlihJ/4WVEwaTNOzqCRBK345pFvrzs+CpPco2vXn9yIUovC6i4jKdNaiWlqspetOjT3w9J
f3PqOxvr3vJV7yKKHeD8gsxB0aIpdgtVIxL57uuMg0/6uHKPzoNu6dXU/XhAETPDbiw3y3gzgGBf
EHiUydjUrZcJOIinDXUBIQBy0PXEuoXNeU1sU0bVwUnftWmiR7G5vp9VVgl2iEupoCopO+DX9eBT
2uw9v1L37UWvyCa9RorIZ1nrkcyiaatyjnzrLWvbxQDts7EYDm2UlWB+VjsrdK7C0zxm1N2SQcC+
XOElcZ4VlGr+w1TJkAMDDXkz4gZz1TnSVstqYlT7L4gqxdZqKSmyDJb9oayhexUcwiNM5KdxssNm
nEkiKt4+9CF7wtDXLJuSwSzVCi6ua77mYLVdpWLb0ksdLvgmF/hmbkKoR06RETMoRV9eiL5z9JAL
ZQIfVZ2itzXV3mrLWj7Twd07oT3/BJLqMWoJFAYWa091Vw/MjDjvGCHrx27EtkSUPxZOtJG7EhU2
a6AK/v7/EcUK0OTOCfxGFQjHlaALDxvsZhk8tUR0dneM5L+Vb6WaGze254y8turyKMzm9KtKRACc
Yi1jmBrVQwoKUiDip5M2nEnYj8mpaWGx6WyXdnTaSz0rjMvEphFpspdTvvHW5vgF/WWDN9UWZpy8
/oa8EKLe9UukyqD4PwNeWsVbrsKGX3V5J++GeQMTjVatU0Vwz1GUoBYZWn8tnqnR4kuPs7pSQIUv
tP6uv+gyEX2gLjl2gHSNDbPkjGbsUwJLEJIeNzH9T+nMWd+efe8UH2AjcBYT44aVRz3Vsq5HJJua
emVQvyn88/e8hcSVy7LsWFTcw7k2ku0OyoJAyCTyuoPfatkVZiLFu2Y1E9R95eCOP9r2onCorEmH
S7EC74LS/EhewhWj7D/r3CWabOLjTfBbfMNX3QKHT/4rQjZICZeK46X5IKu8LZJD8Qy+Fj0T5tc8
81+w3JaxqzcdhVog8sjR/K9MNlzFTVwMsctMsLnJvrygTX1Lc+OC/IQNDuskYEHF9YG+ZFo+yuF3
H0qWIMB5lk5UdRswiWUXBXLsojr0X212KLWjZAtUaN0jgAsDPH1rBTvm8ZvhZoJlzhHxt1+i1vyp
PDx6jxJC+7mn0PpWbJOr4iAMUi0wvacIc6mKGGY9O8yxiirezsZGX8GJEK+IXcUcrfYq5Qev/Hhb
/93ZpWvY2eUweelCJSjWWubZgn1y6fNF4s53mClGrrWo9Na3+cNvAi8fEnuVeuOLAH8yDbVLObOn
BInGkbOUD+Ghcv3vN44ay48Q5LaDW35KuJJD8FcPk82rPoP+V2kUN6utaOB5CO6q7xfQXigh8HHx
hhYM17bU3IbKSSCBecutLqo1tzCBfrmTHcacV0vePQ/9/rdbX4Cm3iCErpw7IVvh0SdTgN5tjLfd
hG7jpr1treas0tKtUmtyoL12jS3Hw9jYVWZjutnGc9y9UU2yrwFNy1318F9u+XsLBrPoXnYw2u0G
xU2eKghdTRjDrfdXS4Vb/BTecrRfBjeij4vUKHeNwoq8j3YRBSwrSXv/gGVcs2cWA8wZubvbYgOc
1McBKBhkthLh+ReOZ0k60mj3umngp9XygOLQDXgr3l107coiXr3+mbP4A+pymMrCAex0GaHqnRx/
ycVZhoJ42I1EtoSxDuJYUwaG8q8e10GgkPIunc0f6tBAvrDkkFmHkkUOqk6BVnZC5QFHld19yvcg
S6PomFNiiz9+9WciuqCSGupueigqmZOZ1hRWz+UiijrTjRjJZniMA6jZOgA8gshAJCosBQy5jVXE
9bkvXUDKftXTrrHUYhuqGif++3UGIxOkHvPBOs7DE3Datg3vn1SV3VMLu5EtlBDTBVXe4iPvbEw0
XtR0c/Ei/HFC95kAyedLVHaMTob9QmaMNkVM9vLOsbiviX791OddoQ74b0q6bzaRKkIyU8zPZw8f
tn17RetaYAVWP9dfjr8y2rLGO+dsMEqC12pOAtraub4aMd0J/rBlPkNuImW3b3oR8psGQ152r9Fi
FyifS4tJ7xgc7OvT6+dEk60QtJIOddvKJTyDAdhu3nEUtUZ2L5tYgkWxG5An8lJ+B7Acf1/ApnfY
tFheqDYKALPHHv0KactkhDeYl5awLVp07bioqy2MRAMwIjNjoYozGraBe+WHYA7BIivhobRiWUey
yI7OBfvHtpxednZYT2Kc4+4VriXqvxwt6ot4tjx8ZoG8qLKvxVBp137GoqmpgFCz81PyIrOQe9di
Ellwd8VBEAYcCf/yKvWTa9Gj/rwP6TCfKhoOeWoo32wm/dj+tCwo+8oC6m9Bkpf9c3dOsJHZgtes
s11WTEPWmtwRs+n8WVLvaiSqN+WRGeB8yMQ+WShg9ZkLPtQRjIS6b/Q3FfNkIwnBJvUiSDvBJSlN
O4Ym0cnyHiRxlezExivzVdOGu67yRMhXz7fgssjgji8hs0G2vTthg0t2F/LOjXwhrdx7JMvXl+Fb
NijWGpesZgqTbMlU8IAAVMngQA4p+Zv/23IOC0dIVaOKJcU4DQ3ZYreqa5KIfZMES3MimIAu4Jqt
7mLYI7N02WtArUWd9clRf1r97dnCgladpg3W6j6UUbcHIUc3K1soi3PZPGwe2JhKoP9YE/aOGm8j
33yIdl8I7lwCEetMxZ+qBcM5piWI/JGRu9Bk22U+plt4GR300oY6Kz5KfadzZIdL5VU+k5PJmYgA
ZRGBqUIpYa5Cx7q5K7baK+kBquNlOGLMbKhyy/jWu+aCjNYPtvsKMPhya+zNvMtdSz5w6Nh4rmB1
sqekpcaDTbX7UqgGlbGTo+n74F5cbxn8aHnOszfFJZyjBHtikbwMpuBhNPhPJKMxMeiLnx45A/+K
3GTmJtjrhUEMlD+RL3biSq0+TpZcd/e0Rl8c4s8xFzcw/HsDSZkXkDKhJzBsmIBlI2eO4mMD8OGs
Cg/PktoQDjLknR0cOiu6u5O/mtbmOrBuCk3jEjFMKXDXJaYKo4Zg14B9j4wB3sEnPau06At08wD+
wmyqOvU1JuWalUweobO0/0OpR3LoqNZGJhGbDs5uCDy+Dzl2bOM74uUrcOVbIu+kOP5ZrT+7rt4J
F7euRTm1PkOARwObV01fP4Ct50BDEa9YKYx5i9SYrM4KG/0+rlnVs0qwJVCYYvx9rmDYD0ia9Bao
qlgCc6WVT0TWO3UzKYtjZCdNih25mG2oQJGnZkMd2aKQVRt7GfrDviLELJ2ppVVUG4UoQ0pFsth9
VE4LtmAQSD0hy2ai75MeI+SYpIpfofbA3PBkX2KZxenqKOel7XoqqY7nr9uyX+zrYbYX/CXKuSUc
PIz42InsnXMC4VHY3YGVGvoD0zpV16kkRt0c84bMKrdBMeb/sYz0VpK8PEAZrL1qqwVQh6TUFKsA
jnmAainafP9iGmQPK3BWDHV0HtAnMW85Z0DayxGoPhDDqANcNsOU+PquPSBfJsgdXCf+Gr/F9jOB
IUvy8lobQxj0LIMiZuGKpsUhKd9D/pBc6sC2uA+M+vnUq5mo7BwI5Eah8Pbb0Ug5bB5IAfJh4BRA
8hTuEts8EFsIvLn/7aFZISHWigVbem1EQxFQAXfIjcucjo3NcYR9HtutiHR3sTB9ULs3DRyjrFyt
Tevu6xYUuZqbSUlfOcser8ov8aF4ofVEjiT/49AHAP4mYuQ726pk0ali+2CBBKZjlPCZBXC9eeoc
+FwMV6QLxtW6EoIuN1VhJR43EoF/Xu/MVoLAKJDufXtbRUJJBRq/aNER1F1twNfUm3GAHVSybggc
q4ajv3ewrGg1e9amJrj/kRzYwH+mdpMOPVPx9zfnbSqnH1pZn9K5eZyTY1+ITgMQMx8Yf/AZboze
4+b/05jpitAWn/feBafMu8Yl9ASdlwKq6Z8DQkMj/9P4ryyB04tiTFPrnSOMF712uLrbCnSi8dCs
S1OzE2zafhsvV/Rm36X/29gd0Njfao4G/lrs33tPuGwMuZTbWkGlZio4vIJi6nBbZnLtTa0rEzy+
MgvM6U/XRwjl5Q8qXCZahymGS5F5qgzTFrKsnJd6gkf1uxViJc63x3kzUL+MPMZRNKL8g1sHH8Ea
JNP+rEj4qBhOZ72J2hhM64zDtp6oNeIUiJjheflwtwltMRdVz6TVSRMqigXpr/Sy5S/Cf8VBfUG6
jHZ9RBlOIiEeei1p1VzvtafUikdlEufa/en5b6P27onbzfQi1F+7XPvrJEOEAbiy+WzX+0Zakgje
rRuhdtC0iwQKhlKRQp/qP6eYCKFNbDuxSVbJVT2zt9u2+vTtqb1b/8LCJlOKlgMRkYrC6zAY4/2T
DgyAi+NRRhIkMDL05NqeWzYEQ1sGSn3Xu2QdrXsohBlCjg1UT6JAbjyneMexBdW79jg2y5F56iGm
IWuAfjrcnNeVwErvBlbTXcF4WJ96ma1641avv5wrdUspwF1dcsohM5ASMbWgnP0/FS1IFR+9YacT
7VoNBIyBtU+YD1ZPM0+j2P2LGaoUCkhfg87zi3xpBJYJCEHuBHrP64RNwd+WvyUjkUiIPj22EEN8
E6nbdxUfWWp7G939cAKfNf9XnK8ozigqh7/H1ca4rDcBrLlbr022B0ZHJ+bWXu+3iIcg5dR60H4L
DPSg5r9QIGThdRb6E58QZKKFmLOkU7Ep0EDTe7jE53kKXg+BnbnVy1m2heuqClLJbd451UFt7Ivu
y/p8rk+7nZV7WGFXFxKSRyANksb5KQuMNyZJLdI8opC63LReCTyqvKfgjDeB1RleGcGqz2eRF5i7
E5WiWjtDT4+pL5Zp3wZkOo5vNzQ74nP9HFz7ppOxSdOSHmR/RXbNktKRotSEKlYEO/qZaKG6lmvg
HmGbxy5WBv5S+AjaSPMjO6orxFKRDvth4A18SvN/IwcS6nCOw2CpIkToqIZfne2PJ62S6kexK2x3
JsRi8GfZz8ps7yFRgLv2+wd7z+SRpQzKifIbntRIlw8F1uOgnnGIzPs6xUwQLuueXw1ujPqu0k0f
kU7miH6Qk0zWS7KeDHn1AJIhtMY36AkWnRV+0LPS8I4QSbMUowlsfZ6meBANGLNpUrILFNHfpRZq
6y4SL/bai4ydoexZlb5tOUfJel6ui+peMUEVGSA5/e/LnJNdV4n5fPf6+7Rj1HfWTsrdGJN5jX7C
2F5G9lhXeM6zxMt1g/2uv5ngSryH3wZZ3u6RBdQag2ag4DbcQgXPak/pQ4iHfYokCvub4BeLfsUN
cZ/gwbaOn6d02UaKGu+C2d97xGhKVOfoIYErlH87rpRZBpYfG+UUKqwsnHqrgmfKxnqUROtMlQhh
0UkS5s44+yDIPcVIz8WSGC8wAUQ1WRgYMgYNcNym0N9wYG2fDGHFt3AipzC8arvT2l9nKstpvmDG
ka9BCPvhlik9WKW4RbSjicnVNrcfLJuV4hLRNdeUgQ9TPmGZdfXlhdFE6f0NQRjaPRUkddGbYelB
9AppIMdcRq2OKd6X6JIfhnYcoHhkOnfQHmIYCMgB/Z3o7bqL8yx90JiBiPODmAcmRZthwS8UKxbd
F+4R7O01sZX4EypqJMtsUIrhXyFAIPTuXmtYdbZmTSs5SWZy7aneZrs8uyFCiQ8TKMIERIYSKdo/
A5uRZ3CXd5JW9mi2G5R3yLW64MqaaBq0qQYJpDpF/uZozSS605KVR1h4ZniuROiuMnfgUdUEken5
5/GIDhz6bT673i+JGaEj7wz9mOE+WeY3boCZa3pvxIXYE8yhbX0+GPT/74esVWc99tGtDA99mpJ+
EvPxLxXOi4+UZuOFADx/qO/gkfg9uRlRs5czTutDCTjDYTTDM9oqtVsSxSfpqqE4/AwJSZtMPdQp
5av3tz8cUzr+JdPTMg//LwfNPNwt8QKr10kiqbf1mnbJn40WwCOW1hB4L5xtWjXj8Jw/GfVZr1Yn
tv6rZ3MXpuueUjmPq0zTtjWduYttzb7ArVQiRbGtoG++luHOlhApT2vhFjzoyhRQGDRdT0iYmoEh
kIT5vwA7IGcSakW7gTM7kJrX15H5o1hYYohkPFYA7EEIbU47p9m1MNKQzoAXxijQ/dVa/DuOcqeB
XF9qt/x4LfUoLOBIDzlDn6+chjsi2PBDtUt0kpmIDmUqh48n5sKNZCpvB0OpkcmFC6oQ/PrmZ/54
C9lyUtSIqVeMfSrrQuVbfSF7H0Igehp7znq7TDzeSY5peNGvz8wc7DksCsh5forPvWkMGW3/DL1/
oLp9xIaefzVVJfRLpzVHmaed7DiZ1wbEu+WzW4YSIaAiWyJlHBjWUIJL2auly7QBNblhFWyBZEq6
HwYHiKnfUWLMusqGQ1qXPfOcL9O3yi2XrKraJ3Q5vV+R3KB09KD49CwgFmHb3mPfjvmhYm1KyU9g
bKFNHUoDM6QRRu1hjudbncB+dvFVC0gUXANiZx2cOrfKYvQJ4SmeQ88zpJ4J9hn+sLJUf/CuZFWZ
RKqfTlziknb2Nv7F/qgokuL5idLaIhFuJWxqXRYiPrzUpejEoIDhbBaIlxXz0X+Szh2jD4vuGy9d
p3prQY7kz9YJWEZP++xqos4i32O+gzktAzau04vKan6W2wL22vAdv5kxV5Po3wpPjsBHARIOpgNE
ZBIhEa2fC9es7dHVSR1vHi/5rH8hxmwcmaA4MvNd9Dez56kc8+yGZLbUqFP8ALRf5rkmsPE+FFbz
msdm8UsR/KkPxeE9ywNXJQARz/mJvo3StgeVRuGX5of6pvWvjZXHcJn2K4W4bfTBmIMCnOeeQUQz
z8J7cUDbcmdP7grDr1MBjFW+DBAJGJIxmSfArf4gxTHpqxv1Kn8tnc/ROn0Og8fKJhI0l1ko/z4W
nzGIq1tyyZleZkshNuX/ww8V/F+fGAR4gaX8Zf0DUH/Zrts3RweazgKH73Lowjatt7L078yEYztH
OrjH4Ah4POaqp8irPviA/jK523cUarKg1R2sm9yWnGU26S6GoED4pIF5G0zTaGmkdG4PhO56vSaf
vdSB4kvmmUvsvsLSS94qi2qxpSJaYoZtp16uYFBMhl5ef2JUQl3j1RPRYrMiWZXcXEvUCu73mZz/
KZc4cfk9P/k2bIfimIROzNZQx6AHL2+/YI2EDfVfbPK8xlLt/bvGD1sIXP8HJ5hq81LS4ZMuKlkP
K07EQJUWiDg7e9xyYPOyk8vi8PM9G3XyIUMCf3+ZY06A1LOAKLZybERquesghos/9FeORClwuCkM
4riJfJ7tQS3N0mQ6VV6+Sarz6sql56so0KeAO3VlFiRIEn2MPUUrqrmLHcFgZGhw0EFL8Zr1C2FU
CYb8joXecUqasGijwbkqLb5tVJuAoQG/A7SXMxB8tV6Z8pOSdHNXPUWKWuTIhqBvIBzX/jajMY8W
OQ4fI473xYncH4sQVIei9u7CveJgd9N7M5+vmLPZvkxdOBezpEUZ74doEQkNkiJy0DArTEGYHaNl
yEoaLe6QjYweOsvDDlIWw4F3GdLP648w7r/sYBBRqQ6H4oSSPBejvc1pgH4/6JvogE/llflYCpqQ
NzwqGiHA5WMYCLJ3SL4L9FW+4ipFUUPw0IZZBwImIkdCV3uqbYfsyo5RGAEcLwdFcD28/bMfU8ia
HQ8kRQvFAcgJRKnHUgAurGgdzlflrecVnVZmqMkMC+z/6InLnFkii28mzuxKjqAieHL/cC70v0nY
fOTTkX8ev8Yo76uiFFaYg64wpV2fXOgGWb7Ki0AKAseg5K+LdQwXNXLURZB0XRq+P80a7dDmqJO+
Sq0cZv0U+yiWIbyH9fZ7c1Q6hEx1cQ55F+ssAE7QlNB7cJNvU+USS2iH2B5Bo9uPOyhtjKSrL9Iq
ZoQuSiZEOWQgvMt1XRt1PEUHLNrWCwIEsgMf1m9FK6hblVD5d/U4nX/EQ2E5ryTg0dHUY6RUbPUH
K4L+ecwT36AMFkhj7mqp5OACSToMglOr6IA7ZIbMufsl5WCjJ1iGmJbx0LfshPgY5rOcw5uTI5EC
ZdpfYs6g0c0YDMsqJV4ELvexk/zc73j8XQdRHBHjYqjp+vxFssZZ5Y+WJi2dmV9zThQ8zwtCL3h9
Dm9Peme83m+QPatOsxVyWoR0Pw02H6kMQzcTjhOkUPOWS+AW1mVxb0Be62wOMvSz1LW7lQibVkCC
pGPU9fOqSVhihAAK14RKCcHtdGAw1NW+Shc+23fCt0ddYbJDDp4iv4y369L/Lhbusg2GWubEhamI
7sYmbZf0T1tNL9Vpzrw1lqgv0dJb/txxlxIrycjfPzxsro6DYylg0XKl6rqPoX/Jfp/z7T6g4Z/G
pqvoCdE3bGyeV1gbJ7HfQXCzF2npJ46Uk7nmVtkLv+6pvhwp141wr6VIMA67MRbf4N096EAv+kCb
AYDDwbc08isrixjMlE3l34HVWLSAIbVwfmKocqu3Vr/Ma1oC2ASHWGuDgCOL5VUrpjj+B2p5n6tm
zrZeNFyTrKB9hcxNIT5w1zuQl96zB2+I0mUUL3N4sDe0f6o27TqLMIClF5d+ejsF0vq3BSU0HOLV
d8GKPx2eFlDMaHzWJyAy4oj7v2tchvSz2oQ2QIddZdN4PMY7VJzeR3PyJIoBDKTRKp8ob7NCelQz
y45U7vywmetHDhy5/QZdsjN7tzUy5Wea/PHQs4xT6hKs6oKPEvJOPu+mHiNyxKdWQv9+jeOL+x3I
DNTEfLlLi0TqdHokwoxjxNL20FZ3uL4cIQN4Qe8KRUJVC9nDxBWYrBK4wrJ4aHnDnlalzkhoQMzL
NLVyI55O343whJVpy1o3J28LZCOrTdVQv2jzrJJw61+iXxBd+5aMIbnl48oixZkOLg3Z4KhSCl3E
ekGFGktR7ePYcLN6gOuvV9XEb9DH/c7zrB4ScB3AhzAdPKjVX/bRuQxk25qZsJMmh1FOoKdP2p0Q
8dpxMpX+hM6TNVoVNh6v64bTvFqCmwoKiZfgG14MKloSC0zmyezqpqIQ6cHQRUvSfYJbN2pnbupA
o36EXcfJgVv7LjfMsD27ZuiG7gWyF9/9/ykpsML1g+IKD+j57FbQx4dz/cGRRQ4NJYIdQy6h29W9
fSvAl3F5kRCZwPc6at3O21xpzql8xq2Rhh/6kC39Ox6+yxs1UtI8QJHCuFD3LJYf12OBPUfk73Ah
6k4GEkYqy8Nu7mrQjK398n+s0qa9oFXQ++Gm909UJXNSRQUhOcm4eWVoeOkDQSQz88WMs4J8/Ap8
codsN2sgrjQdUlYpe4Du8XYWMSoK/cXV1yG3RdJZNQVbuC3XwVx/YXUskqVuuCQgv7/9Zm1IVzR7
+H+k62p8zi54DPeVTJ4igvshGY6ss5Cs9UQYrxciu6DaVBiIZBQiK4jKIyX31rP3mIohRPgtvnju
h4xudWxYpinY6U8xzi3WI6CCaNUT3MoEJpi2d5XTXEYtKW/sq0+jcScxWIfyRbudaLX/9Rfag2JQ
6EBGCvrHDEo/wwcA7uPn24d9XgrEEUHK/rF/JKvVZJBZEM9211g26y1vZSgN6cS43VMOyPjpULL9
fd3j85OrD6H9ylRT6qpxreN/5RwagRz/3Mp1n5NYlEHzxuyhasMyPoVfoj0+5J3KFvclJpnQSjYT
CRuq61kVU1CU1gMzVKhOlBLB+pm4jw1FEq4gt3ziyQxz4osKvT2Vsx5UI/uS4m7/6sNBXE1pSe9n
t9x1d4oRKbgGy/p4eHuJpDpyXHxh0V4rCopAX8LEI1v8Giov9b10fD8hEN8osmh1pazBELPErV5b
uAxMFu+CWPecvkZ3uim16CQDk4Jh3/ptkb00dq9d5ZfNRxEG+DSwnobGuhbHxV6yEQV9YzdmDgEA
puYa2iIOFJVoalFsR+zZbTKzXX6HaUcAIhvNHNIG+wLS5y3CX1sWcGxu8T6pn4SaLXlxkJ113C+I
KKo6b6XjX8rldhHtjb2ZzJ5Pzyl1dVokrbfuzbfdFeyI4p7Aye0nqO049QC+nJE5UiPl7SF4be2i
r0G26V0py7fRJthkWYuLo4J+d0uDy/DQdqaWawV5mhCsnfgJKqPMppOusniTroHpLAuB2qAK/XyQ
6QaMYBEonocb+WSL8Bbhpr9KqgXJ2GJq7PZZJK4Y/aoLdEUNTSr96VojbVC2L7kSOeSRCOpAHD+c
W5zOBL4Pr3WyEYfWdQ3xb2jOC/YxRI1JEs4a7k3yA1jYqHfqTH/umDedwZOdLGKIaj4xql56F4ne
6tOQN5uucipcf9S50QalckQUIK5RmcfXDJdieO14imR5RcFw3mTYOrBokrwCVpvPSc37eSqZ9ChX
wIRBa3SBK0SunU8QHv2GB8m9fFtkdhaK6Slef4NSdi+wWGKpVUyBXKYVAz3qs3xuabKQhdNNif5g
YVhZEQtS3NJ2qqeFQz5GdVxKLKV0N+LxY1YgVwGDNEkH6/WzL0vP66zJOkaEUm8GS+McdKbB4Q7D
9nkkpgF+uUi8wrG4cBNwt15XTrThzdaX8vd1kmkxoJkuqJFx3syIKK70088Y4mh3cmwTnZCFT/1y
qdJfoUwUJtEtx4T9PwLok+u9a1iakc9dfmKu0/3+WTQIO1HZk24g62aAw5NUCcUClRSQwNqs3v1Z
XT22Vu3e46OYgNiHP8L4Fjw5BhQR30x8Cs/SiXS7iYUzHq6EF6tckp4b35p30EzfekhhOKHCi9PD
U3ugMFT0YiS21E0jvPxits/+sPP6rqJ9VMGzzc9EPyf088VhYw2CWVNEs1utAOSOTH1LnHhXslsj
h0ruLXb3AmBfVnryMn7HC4SO8dIshbQ7JFHpAH/V24KlJtZC9k3gWV+0purk2txwt80BV+V3+EBb
jf38zpXdLOgPDRwcSefp8deV7sjmzIIOwuiNCSl9Dn51794DgXDkYltifJRoMDMj3VtLixofCtIN
AvluuHlZo40+cnWjaNCldJbtZ2Putm6+yGHoOnElt4/hWIVVeJJ7ffTXd6F6Wj/ZR5FkgYkZsIIy
/rktMROAEpedR/QZ5iqRTHswx+Df/B3YHgaGufeFOc/j967k58MO0TnrWQ1Os5GAARnZfwEBHYfJ
FqTi3r8q7vYdOibR3oQIhunng645srFQZ5WSC2uLa4XmH6ktUjxdSPDEjF2DytgkEv/35rJ9xn6O
QnK82JJwuxtVjaCw4o2ihXtPvr/sMt3YC9WjkSu752jH12Mwx0FQaAPWHWe2aV+YfkYIzni6hExP
2ARz5b9pHw9GdFo1qGd/mfKZYAhIpoQr19NrdAe7NEN/aE4+pXkiOyUT6THSjXlLWBFg7Pym5rHq
8Pcj8uf1PiPU4dDVSkKm/iPML3AeeVzcT+VqoA+buphalWPyNfj0aU7XhAGdvsfs2/OAf3sbVNVC
fAxKBFUft9+vsEPLQm/hISwYzg3NFxnoD6NYRXNp4Vm1ZgPLZDiMWpDvMbiEzj7HrLDOiTFYqUgH
Tbwkh1PlL0JvolHLOvUG3kD3QXpMwfrPA495TILXBU+V7t5CvobgN+nmK915dVlLl8NUq29yA3K6
IaTW10zAw5tAAdwtiSzxdUD2QIQIZBl4uFXAOc9nXOeL3wtidtdGAqDAmA0wLyN3dHkGNkGCaAkT
UPg+cJN9TfNMlWQV6ewqwsseVRSPy33CJVHBL8hnFUbsPmK3feYjW5fh5kRDxyxiTAt/kzavP2jf
5+0mMFXh6se3M46T7g4h7x7gixv7LC8nSSZZxTCB074womqWo7yBuz3gjmsknK0QFs3i4irV8gHa
lqe8S8jeO6I+mooPXtAtWOsvbPwaTNaTsuxcPTcG1I+TFls0jJCEotWQkcArc15hSZVJ+JYIJ+XT
Mt4iGPOvzjL/vcJx7nsxzVAcx0Zn8MZG3aUVGKChCd8rV1WMs7KXltQPh9ckZvmgLDuluVDwcTcw
ERj+MRugZiL7aGwye8IuAWhMWh8B9ySWPn7yC12EuqpMZz9bXpTt+6+x+n+c8N9ohTIoT0+dIhMj
ICrsYpwzmA+nwJ2o8C8aVOHKfooGTI7mDbnhvBW36b71I/mLJH4N6FnMBZ1eRdBXkHwEBCxgo9ZU
Ufp4dMsZntWPE1x/ZIWHWISi/QrhX4zp/MRoZjbkgnOhOmkM4xpT9jE02pBXcAdS/5+I1KC8uFf4
o3ktK5F3avrfqu9jr5T8SD0pPWQVVma0yfZ9FfNw+fWwF8l0AJNLYEO1QambUBY+R0yGrBjM3DeM
ZCzjf28qptnIgJNHibMXMURhtZEJXRrYqU6tAM1CYED5Ibwp8IevtpGYmfb1QjDMkOqVtIB55eNC
opQ5+2trlNH5xOKcU0RpgXdtHb6iQkjxBnTqSJjOXzmg8ktRbDrjtRo3J9f5VPlNQqn/Gf2dXAR6
jGECjl/7gNiau49AfSKlHbvm3WrNCqKdZ+V8sgFdY//NedjYiN2HhqHv/5C0pmjfLL+YMBpDJGo6
n6RkZ6nNmW8p14Y6g1lr2iRSusmnT7mTcm7RrE72JiNifviHd+4af1ZBUNd/0efOHE7T4hraZ/9m
CtnnC7o+4jgku7Ah815oVN24JVRcB4LMQiM1xgCdgLWUeRPAiMFZ3XsshgdQorbtLEEJeHdm7pbh
B2kp99raDRtqumZ8gXM5biJhdW5NjPsEkDTqYIZLKRe7DG+LtofvVklQPUOFyI/vTD1l2TvAbnTh
5ZKX4qPf1DDUt7LS6Aj9qM3mBJndVkDqHQkPp2q/6f5zj7OcFRFdcwCYNUF7CSmz7Eccv998ol7N
DdPNgHdOANex6vKpTXA+Mq4A2jIBknJgQ9qjMTsXPTyYIy7IVc0C5t7RAW543uN09ffvwvxpIhEy
soZg9kb2mDjTHgNUbXWmHsCKqrtco59yh4vjsL0d5Wsq4PKjlt6c8nUWX+9whhDTAr4nLpiP/4hR
AffECBhY/XmA13ctMKfgUgf0U3mPYWsMfEnBUYhPq9Uq+UfDgrgsREXgZn3aXmygawAXYIgZOz13
CJBWKb2+eb4OdeqY4RnA7QMu1r306ucqX2xfoNEODGkSEZGwcTdfIT3SBqK7h+ogy8Sbi3F4W3B+
GNJswIMJug8wFR9okxKkYxtVLBZStb9HrSfFqNTMddNZ02OIYfp3lO0r/3rtNtgSV3Pk82uFESyk
PbRbeZMxr1uYHNSefoUEFat1LdjG9S4ZMYdUQVRURg8gj0p2gs4dL+2HGA+/YvCrpS7dMUvV5BaX
nyzg2GWIpSu3fDuz3tGFQZVBrBbdaHl1dRoX+/glh/ZGy3CMyeeAl5VgGEh9HItIyrfurnNxsCk5
GQ3/MWA8Dm+QxfGFfJE/OsAlfJknKeHfqve8pC+3NcrLFv4zB00rCHOEH1mD2SvNYtDn9/n26CiO
sy8x6+E8bs+UoU2z1MdHkQxdEPo09XSTOGBCLrSe+U+EQaf3bp5U5LOrkeFO7/W/vy23PwHVBCu1
lkIG/LwEOGu/8CAqGSCezJATEUuqXZAi36ZXldsgqzQ/pTc4GvGSGWJfEAjfVh//dgzi+wnuFWt+
CjaUBBQQZ9sE2CJvL/omWAHNM2Rae9uW7CRexNv8rj+Wkxc+3+DHi/EUsI/U70KIKTA6EAjAHp/d
DorNItlQDEp2jF5RpPTcrNjW/VRAzY8e1mQiudyrU6klM/bLYTfH4YHmmBVvH+ld2rpL2sXqM2iW
In6XSqfczezQOHUc/+xucnoyqjWoK1YJDu0Oar+5ttL5k1i0n+vG9389OPZ80drtsBKoUQ1LY1MT
3XMXb5MdAP4ZvvX+sDh+cM0evUsYUW583Z4gJw1aMipOUJ58Lsn4PakJZrHhXlnb5pHg7JG90Koh
SshPFvJxbz6jt/Vrh1XVngbGY5Evp4J3PEeqRv+WkzEDDRQNsYKkyRu/eQCe/n24nzJvp1KDdCWP
nVyzVgrIE4n5I0vEyFD9xE2jVZh8safAL30TQd7YeW57jN2HmMCFf+rocsOxMQhIhHVLBjQ/pwUF
FFb9vvI5SRiqhHGLv7f0gzpsu+8x2lVrDoe8dXx2Wl+bRLOnkoCYqfOMwoRVz0b3Ygi+3M4GWaVv
/pp4WVhSfFeFSvTRrQBq95Xh4OzmNfqdST5Y3dFfob48D9jqM2MeHu0+bSW95ICHQwEgNgqi/4k0
JjsGb6Vy989bNsHH1FIlIdjFB/Svx4dLxhkjlzmLQ/ierD9iLL+StDn66inDFCBhNDymcMg8L1mb
zwcZJPrSYiF9SU5g/EC8gljqO6KCH59YIrERvyCZpDp0iF+QqvI82mc5h82ajCuCjwOHG3G9NP9w
LWeYUpEuIrH/eGg48d5pt4dk59+MrR7zSleN2UxOwwuSKBK2D9vz6Fz2ObWjJmiuOpwAONw/+lg1
n/k/mEyWFutnHzSU/JiVz6MTXic0SdtPOKEQktMop6UAHNAHETf7izX+xF4kNJlU49MTr5KNVGtf
prpNrquIplZeUiS5BV2/GToEHDOD3lEdIcsFLv3enYl9HEyeRTLt9tGZ8IIO/LSyGOTb0EsheI9l
QXkE86Va+z/rQHF60+adrwSmRhf1zQWLp5LrV7FSsC4T9usgkHvDMm4tAPxxPq7Wtd18ARINLwjF
QbvMchziP/O6TyAh2CHOu5Jk0625dku5X4xV0AdFRdOgdfbSobqz8+u2CPyO/5mNlBfD/g4ZlQFr
5U6qwhbYyQvcK5+yq3wtNMoj8EAHYBJH/nfwPzhMLq4hoo76x/5Lp3P+VYRC0ToVw6NEXqRY33Vl
py1HZVwV527QOmHLtskX5Bk6gGWVu0sqQdWP+xh11NRUZxPYslK5gQ7cRO4Jpl5w8W2nYw1JRz52
BJhzqehZsWdb2A0FHvDFFaESSw2naxstHgMUcZcOjhiMBtFX+lv/PxFgdMxXYnVOCWMB0fR8miHq
5blibNjAl2n6QQm/1BjCTj98CxMA0KQ65Ok5ZP2V3m4/XMaNIiSPK/aXDH93Wc1RpAV9eTzCm8+U
Hs2xyAe5VaxpQ2SkWXteYZyCiRaYZBcTugtYcd1X1inm8aIVcFgLwMrhmdvkmHKImVK416vmmvoy
7m+Ne16cpsWQZ8qPetdotss2bfb6XFe9oxCnLOqqLftwZJN5/vpWLtgwlO5sdFozgOnzvnBBiGqz
aLVu/WeU/dw3/2yK9QsSjv+wpIM8hxdVhi+kzwpEblmJAeQFieRLWR4AOPZKorgj3BYvfvkIqJpa
jdJ1tEn+B+FDFq0Asn1VbbwBtHs1W6F3mmANEl1Lx7NFJrVJ/Z3X3qBhBSf1rMzlhgAPZju590j0
o9HsfcxJTh5xp02F54Di8BTLZmMVyMAYT3kC9Vm9MXa/2RU7u6ruoyGOXcHf+COIoR8tAcB+YXpw
Mpq1MEWJ84JQcPKqdLcLGb4RS0mZSt2EwBtrdQ9G4Un5Rk5Rfm7mDH5MqSWMc4jsU+i36B8a6IiJ
7oDSATAiMznjhG56nKgL+Jv5NtfshJwqBe9rT1CJo1GujHttHwpUkDQQUyim5akBon4G+JcprMoq
N0IGmDHH9Hcqi5w0qb//+OtLJ/yxSXGcVPXCTiHy8hwM4m7gBbuxTewTseQWC0zrrAJXAY7eI5Wu
ODVA+udRJPNpsXXJ3QGLROcWC32YGCbcU1CfrhD+NdMOSmqoIYlht1d1W6CxDm8njCpKYnwEpEpG
lDP6uO4ox/FWMsyDgLbEreTVu1OgbwyQ6RzdVSz5UpaeQlsxODR5CyCe0x1oEezYliJ4apNYUqAw
0/ijohTvw7Z/+qEPzNBeaAoUqEbfL2BXtaIm6KQP/qUfggA6WKuJ1OOlzPBcEDwUXY+Ih8JWQWQI
mRHor8uLJ7EdjhD2ULOfxL2+lAh175lzcg48BkkSnRAg8kLvl7Qwb7h3XMonvzGA1CYnQRL8prEW
JoYQ4PvzKpZrLda2ffUUXPgIZ5cN7FD/3gLhmk8zXjf56+kCNaU0xdgCbcbBbDnY2lFDTiHVySqv
jgbTpbgzXGnhTe4DEE5MFUheEkwtukS++yv68R2F73y2ypwxPRMkoiQjcbN2eaRQAPfxJcc4l3CY
y7vdI/fnOBbZjnXtf7nlB0yRm/JtOp1M/pYsiQ0h0cEp7u/WwYEHNQa5UdhbqQx5mRWszp2QXLAf
Bmy146BqHzXD/PVdhRryyV1Ewp2XX29tKID84OL5fo1QDhZm6irl17/k3/4LxakVSl1Wpk1Y6SG+
hRAcBtknD8tC46vSH4dBa5xvQBlXOfar9IxLkODjytFapjq6APTwvmGOnXarPkY495vkcKke0HFL
QFQkohlOCq+wF3pt5SrMyhpDFKfGrEvTSG5cFPjgFikMg5Vp3YoCPZqAtIVAHcjqKlaVGc0uv6Cv
yXXURuzxd2jU25fLVml4bfHM4zLQ04d0krFKT/9XFnHbvYL95ws1H21dnw8x8worNyj0YiLerfK9
GjrXpNU+qKDzpNcCwwpm4fQMzKcMhENh2heVWpCS0eeCRxsQ97NRToODGt7LuOr7mflQr2PAALbc
EwsRjPvGv2ijMb1WyRorycggPP+yA5onRAtOMjKpv2FfZT7hUnrG+MYPwWStaz4TF+mryF7/HgZ/
ao3Kv38CEACWHOkoOo44sqjHjOeHocNT2AVvzuNoaSt6Y8Hh0oyu1afaz28UzGe8fO/J/QqycK2n
/tp2ibeKWJZYxFdyJK4H3IzCdEmJtlnGzWCTWCsPRYOsqQ8+QxtDkcZKf6HOrVu4t6va1Es90z8X
Hjpnwu5u6qxLTU6InWTuwB8HwM54WBWBw98DBYcTi+2rthPvLEudgcAYwd/y/InwOb0X9cp6BUmq
qVwyybldJe+bIMRov6BJD/5cphFLtErdH7WJYjaUv5cydo7A7CN5eXcZmdaY0rvZ6BHyv7Mvxatp
P576xYM9SAFtIXMVWp5JbkQa+qdRI9Ylkab6d+7/lD7TRRPCDqd7VzAJ/Pa561C7EDzvk5oIGGBe
U3sB/BGFtTBEP0k8w6j7KhRtMeylEnxY8/FoOBGM3HOl9dIxBnsnLTHMbp7XsR4EoFau8kryFNUm
fRVGCMPuHtKzW/X8mUkAROH/aPlZzHmK5WV4ZEt/IDed1DdSsnc5aBKObgNjHYE0J1GFVPpAZ3+y
Btp75VVldZzsFcM9Juh5PzmG+/1njUJVSWlNKwqi8hg3HqnYwwU1mJWAPMTI+1nFaecYJP1uDyRj
nOIhMlcb/scWOzeVR9pdIK3Wj8zxrMaTQDvIZu5nAeP8JU6Zk7E1ocdtQwBhl0nUVHnvcH1FRX3V
KnBHfZ2tHA2S9s+SgjFfEHXtG0D5Mte17RvP2ZAqidxlnJfIzZRqa7jZkG0Jutw28Om/7iKgQerw
U9Z1di6MF2EH+1CN5vkdOJByxQ5vFJPwdc1o3pYLR/zzg76NDuzdTPNo198O8optKMrt43X3cVVM
OE2QMFO0DmzIFmlfMnl1Rwk1f1soLpegyR6CZJPvvbHmxWNr0dxZWaoZ3E0/22uR4hHHUfg5rC5r
+HF9CfaZnosw1H0SqlNsN3SIKbgSlh1zpFLpHcyNAmbiPjGt/H42jReKHrc9BoJ2U6J/wPza4xp3
6Hlkf85gdnuUfdS+r129dZaHMbFMq3jwm2TmTkPhrAsch65axWgGWKfa42+ZPK2X5zX1BgrOmmAo
a5JCsc+OLBvL6GPnOC/6nUW7zP0nJL6kBPBXNi8JZ58EHHD9q4vfaKh3mC0/gRgGIYDxCRJSuBnw
bh5PrYkARN9CtRiVrpuug1hCCDhEZUkGsFJvlrv6U9GSdLLPrJeoOl9p0n4bdwpqfWHQVr3aC8OD
JsBBnmr6wRyNNwbX6OMr1tRw10SCA5DnLoyjHdsKoIGQKS3R0SEoYDGYasfZWs1Wi2FgABb9zijm
tj1eWiYYWIYTD+z8kh3aGauTpqtzXJCMXmxHtpw+TuYpgFr8cW58vi7gRVDUkOujjM9WQZXLs1gI
SzQuiKsxtosxgym6AMa/sfBi0giNOVcfITZ69g2o+HZ+dNBOe/NieMmMFAzkEaLOmBVHqZzx12/s
mdW2bBxtWD8C1UGpVtsYiBBQJS77pjTqD9irIlsVRwUHVSgiHfPqi/59GzfJFcKYcCp5Ltho8rE7
RMR77nW7rsof/6UOXtLOQtlt7+LW9+lBTXP9EfURIH7UDECxm9zo93c4G2Xg82Pi2+/Ot0Jn4UUe
XCuLIuS3yjretF5KlrfGti6h3vFvLPs5tIb5MjYji1vJC8t2jW7QqiecmqNHmnHJjKyEwtCLj/zx
mz5hwQXdzguRbmHL79wBwWXvhMuQMMdPAraFSCJ4vYQ5X0A+IRxGtsh4VN+X5SQFIIjxOAb2cxxP
ib19hiM9WiweBOQgiBHsSGV8ZD++15jcEJBMfaPM2V2nnW7mopELuFtfxIe1g19cvghoLSKaTYkt
NvE86UrcinzdyNf1wCj7ijQoPsexOXqctli463iSm3/fZdD5WbYDOQhZys0Nw9YCWiHDefxG7TBT
HaQZ8epo8DKjsNE0yD7q0s5lhXITYvd8iJACSXK6piUxJ0j5Tqu/WVIbKz/nVJT9GUxWrXlPHIIg
tmzaZ3VgoBZoARwN8FDH6BVMrDN7UWhflVXVHUmLGeX6fKVCNHtnvRLpEhms1D55Xb4VYcWMdQg4
HRN8E0aVqpRywQYmyptMvVcvVfkCTiqsws4/HI0M5VD+245G6l7aUpTX0+JDTZY4JanAo4fgyF+C
qJY8QyXQeb3tb+P0t2ps3fvHIE6hcbHf9QLYW0u5+Wze6JAuVf0z+Z9xKADkW8XEYgj1Ux07Bzvy
I4nGjTzKePE8GUeC2OO9q+AT+Jz+6xo3qqb0u4vwNqY34ZVBrQ7pgShtswxLA7XkaWVITYXvya4b
oxilGutg3yQmj19xlXbNbGDgRJi0o32DJnkoD51FYYQMjruOL6FH+69J9xP/BVbJxS41D8yN1NVy
yJhJ/OdXC41MR9OMYFuMpM5Mn6jQ0A3E4Fua5M7p5/os3fheRXCP7rLLJ/u7t3QE515qQQ0SA5R8
nRgMy0vIxSxNJ2pp2SALqmq1mce0+XtfzO+PCWcROg6bV7OWVN2Bob5H7CHXV8rWNjgoxf7QjPEe
Gb/xzOuSdDmdmmYU8g+/1MnW3Rs7V/vpLMqy8RZoWvChI11l6yhRYHwljCc4o2ffyG+ECem+cOEf
IqUoLpXCeah4/1EgB3KohDz8Ne6R4FRuC7ZBsolhQz4l0xtfyHzj1CxqgxPRWOtiDtx4saaykgSB
oFgrvlBmyr3zfYJoIcgU51GfXUZYav44HxmjOhSkme09N0Sj2YV/0bw3svKJX72Gsm/ZsczenMKl
blbB7xh5+n0/pXLhtAPzL4ZMd6yW5tOuDKKGKJfDzs6xDqtn4sloZHmt/Lxv8NAwzTngWlv6mOhY
OCJmzDdR/xJJhA6uxSf9wfbZBdgpLBl6ZNN0CXFF22VyDPH17rc7UMI3CCENrqA/lWr87t2Y0uLR
cXGIp/b+Ep6FI99XniMyHkWVz9BbeCqYdxH319IgtUqYpLbYAh+D2NW4Wby2TTvk9Om5RL2GD2jr
GPUZ8NEeURriF9OhGhqpERQ5mbuphxzC2XsI8dOs5s4DmPf8HFiUzZBy5j18Jk6CyT/n/zASMjQn
4ClF82UkuNXlUjQgQQrMw3/1FQlFoaIQjGXxE3NJocu1m+Wi7sGkybGRqC4IEj0R+Pw0F7dfLInu
5fWCM6ipbWv9Sta4yNztNTWSgYvwfYpWdqLPnP8OIccONAdIXm091Vy62qggyRVgFHylnKGZuqfn
xKKP+JmGrPSzd2PoqSTabgIqtAKvtMpbrZjx7CWD6YZ/pRFJC/I9gfV1jCa6RE0x9x6FwgoUnTG+
nrM795drZLsy4Za2ciKA+surg7HkHyoSDHm2Ox3yozQoZYtFcQx01f1DwshlKh5pOqA8EZH/VKmd
LqD25oAiB67LxKg/LZ0RytHrjXuiMgIzcCPrR7NcQkYgH1t47etNv8VMYzuoVELTD3u5Zg96z+16
rP+93DHPwcgzGZ7fbKQvtllGc4Bp7cwvTMhWhY3HKm8Xy5jE6T/Htqf/M8My5dcAziuDh54txHBk
ifhXjuJ65+/bkacjeVSt2HKrbiHGe+keD9qgp7kLx+4pV7nmn+PsEQ82JVF/XVt1jO5UBtsaZ+uB
SdNST+fNJFlncLn3mSpNlPgVQynvk5sGptINTucYCnXYVyMM2K/jJOOX9BBm/1FAyDbkMY6TMlza
qMHyXr5zE/w24KTbdk5pTdXuGcCy+8QRvPVfLaD84ezH5ykLto/MSJzrrG+xneGoXyNNOCUrQrW+
1O6uAINtPx24oVpf9+Mb3tZJtWIW1jMNXCIb3a8CMcqnQccNPyR8zvtNAvw2fTf2F6H7tP9cnADq
Dv+1Mut83PDIt+JOfuardkTEsC05Ph7zEGO5QvvvasBsZuGhiLqnbV0Yyvalhb5YJTCHqZw68Kkt
0xDKanjQUXG71gH7DMvbge/EJbci8jsIvxq9kE/+qCLR/14c8TPnXKJurBXuyhQPLQRTqsqP93uW
I5u0riUlAnZfEJWHqyxxx23U9zCUR2xsQJKuBDPWD+VVccvGQzaPwdxFXJsN6CjmeBgKTlAOZ/VN
OLzw4Ibwy8O5nZb1joDVuuVEaywMT8sA1Mor/9KUJVP4GV+Q3MKIctPwFtFcFoM7Qj0mHXVHJQ02
BzGtValDml8FCjopcN3wVHLvDj7ki6ZTgu81pHJvB7kn92E/ZDTQSIG0dPkiahyS1He+FbX7JJwk
TV8hqDk8CMAkiwv1CAfrt/7Bn4kbXBkmkoYW0AyPgEPYFHJZ3/Dpn6mZjPq/foLrZWXqPNqSR729
nxExx8bGJgOaK4DuzvyyV/fISliIETcCMFrfFWhfMSCkYJq3zYrNMN4AEylBjXKVkJSK6drWKfzG
W+P4rCA60D5adlqyfXfo4wjnPdE1mUIhCla9UcK0qojeULjxFNAt4xh4yyIBCeTFTp85R516OVaf
SwMaU9ewR++8wKpArzAv+vpzupouT12svA2s0hxYw4/JN5oop9/QFMLUIWc9R7y/cKxA0nIu/umh
4DJ5LzFfT4BTHtKc3FDmHeWeIoJ6AI1dKJpqpeudUcIXZ1nY7bL1UmI1nuwOS6s6i35Adg42LXbn
dUdu4JF9X+BRxKY/L5g3oVof+V55dqoZRWZCC72FJtR8QfESjH92HI0ShvJWsdEzCOtOfhA2lDA3
3C3xV791ziWlp1atRjeFH9RMtQQ4Nw8EPs60YRFikSLqqvepccmtBJ2R6ED5lPdSxhIcuAaJP1vU
pAJ87QGxoJUVICzAl3w84CG8A2ymyhi4fVZ3ANcLd+9OMH91rYkL8SpuQJyNddw3sB/3UrhQqQoO
AUPTVZwedauVomPyBrNN5e2KzvM2jxRjUKXaEUqpbvGJMsBWcXnWFnpRU6qR/61lb0pZ7L+JMaa2
ibeUIyfjltINexI6g4tS8gJ6R/gjXBsOJvlR3JNQkJ4xfx1deoBN57STjz8bCFjgyu6K4v0a8tEn
bPGTqyI1g5WWGfJxtjIIOZ6/nLvdWWrtYDrIrdlu0b+WH2/lxuG/aqpvu06Fs8+hR97cW0E6HuCn
WX+u73HboUrAmyiY4YSM8+lA89ChgAuhCHLaMR/wuNYB04c++YnrjrRIuTctlZm2Nfe90mRo1ua/
aIUH5P7EUfmwn/+d25PyZplMzC8P3kh1qcyOPf2uJ3/uhEFrhyfR8CZHg82gIlYzxlmnJLDg6TPU
s5Shnil1Bra84UkmsMYNR75gg8iFS7/H5u1Ub1NS6WbOSpGHj6n5xrAIka/vy4oSzBg8Abm6CuOK
IU2x6j9XJXlcZYfFaA35vh9gawjN8p59ITGYkjZQaDAcxbxRS2JNrHa8c3vXxUyHNDvKPNiHwDtG
jW+1MdxNRFLaEpksHXY8ImmRku/V/0MynaZwrghbbIH3GIaiTf8SwByL9AjWQKdWGGJlztb8Z3yi
kcocmYmEsQSKmQo4KOD8HsLucz5im0xRvNslTxDYt2YaUGjMxPZYhtssMlL0/MqQOkMwQSYK/m9B
qfdTQnwkb8qCFCUPnQnmeeT4Il5bIojaEY634J8+pZTxxexyRUMTuRXb9E0lOiC9UK+gIP68Pt3Y
rHRT257TqskViPFXYUaDY1UHUaboolWER3NkvBWjGjnlO8a4CUHBg9WI4X6yHctMQwWbFm4GkDaG
fBAgNmi6hvqs31TA7FLyQkbmrGcK5q7rmMOphb0V2XpnU8lu8XplBsrNE7nalL5AOYuJ8krzYfY/
rXWj6CT+POngfFLrkLMJnnx/7poVRbfOHablw9FfpYK3nY3za63T3xAt/nniP7oEKKjovu1cFqbR
pTLpzHg6xRA9hTCOdQTouBDjVrofdC81Namt2rsYhgOUUIlmZZQ27Fu0GH/29+6v7m4KNdnLrDPO
83JVzagUEKOHAuWaEE5AkO03DACi3BYvfZBBbgbUyEcDEIcYJzRuhoX93oxP6VJ+RzxTKnwx9b35
3kfXQpLBu+80pxbmkaHoNa3WCjExIY+zE+FUzb4eXhHXptybZBT7fnfbrBIT2jQkq9YUqFfTBj4r
K/If/LynqebMhr04o/SFQp846wDxlGK5bo+hDqwsF+ibFeXaagC0JLS4S+o4VTMheDR3hmKCv4P5
1XF34ax1i6D6eFInYEVFljHxl/fkxlDG3EH+m1DTrhMAtCm1/A+zISphKXcJ1c5QUXIDoxS84QYL
duqVDWC0zJ0oKDod8rbPjUPkzoWA76b4CIk2r8rVjB8u5HhWGa2/LeHr2HzNcRaHXI207lget+FH
0JXW5uwucPxbWlba6sZ6rFE6o1fgL2zfl/xQdDN7Bd8Zur90JSQfIUmeBzJQ936qNlnub6k8Jg0T
0j/eNAPHqInj21Pe4sjkk+lpd+Y5ixh2xFB5myM3vLWNr1BeQ5i+lvitvBBkgNFoyaORwNgbbU+s
wI7i5OEAuP6d7XfhITrsrUkapJBpP+0hGxu0yT4OdKB+4vomLOqRsrhCBhjMBOolaPjLIRgdxao+
jKRr7SmijxSAwKQqgY2tlDCGE2sXlsGc51A9kvGmI3CLHI6UxBH+Ikg49JWeLfe9IDeY7RvbZKV2
l63mEZbK6Bvwie0ZJFwgpvHvQmT5R1RF+CyTcGTMPlR08BCrg2DUdArZ6/8pxBn2MR2xj0H6kI0h
jD0hs5mdEl5A2jkwHFBzyBnoXWhtukgA7bLzsebM7fGGr04fLz26YliWZoDDb6VU6AaovU4WalzR
IfPQb6gg5ExyfMRKEI6LgpTqbQcUFMt0fTRJvxq3zVZUPrlfpi+AQfuKfTqLGkrm2De73xUZrO5E
0gLDTjCc+WQu/Jz1NVESNpf5yliRo9x7uLxehT2gak/WienHgPDBIA0jfsDPyAtghZOHIffUp3Fr
wr3obLGxyvRemrXqS/god4MQ5rQzsu2KJh6AF/w7Nintt3XIRIyibhnw7ZhMFt3/ORkUxTwx1l0w
oSqKVM16WnC/UpfAJM4E8uBytCBmgIksf1XZ3zMPtyKXX2lAZRzVGOeTdZslJcaY3aCjsh3HWTWN
ffE4q++05HSi4rvw/m6TOR91W9S+zv0c27pu5bs5AZr/AGvkyDZdTRsI872/R4CjoDQdvJ2qF6od
dTwEEIYTMc60fhAfg0ZqXSgDk5MGrlrq0QRHVhyMfz2xlNK9AohaH1/VkPDZz4jZK6zNZTydvYRD
hxOa8lTqDThFrEeVoM9LL4HJUoeZRrTuqY0j/xOlITq4EcCeqtuE+MI3mlDLVvBHcczPGWTUZEe+
+YFm5+599BNJHVoa6/05sImv1jXtI8yQhfZpGuBd/revmcGMJ/9lqCgpLWyZoubMOPKLiuk2MnGD
HSC4RxneuO7nxN7ECdmaET3x2QE6f5rarrAXQtfGoy+rryFjMdEj6mN1VqZByl/uJKXSBw1t/qQn
wokyw8qhNDNgV6VWGpxB3YpAcsCCCjY8Yn4HZp9Cfcz0cJnvziE2Wy1qtse7e2/wuNXX8kjXq7EL
jtorXb4LVNmGpi2PgZ4kqMaRwajAWKa4wAPgliLa7wdb6EeMGxWG5xKyoQUPxECvfn1JN/U5Yjh7
Q1iynkRWMOx9itjl+XdOB0huW17rWgM28NfFa5TblUV8jp5QMi3rhc1oSxp4co/0M/4R0CiAxEvj
SxQxyLUyiOZwI0qYlOuPYFmZcGE9zaZdztscTnMlQQ+Q8n0l4ta2+mf6Mj7MRR9p7oAZ1QcpiGRY
ARwmRIH6klmMqE6yUhTrQ6Czbqv2awbMmKnYq+Oe5IrdF97ZQqmInlVuRqRwlPwYcS3+645PbBU8
QgNEyltMixPBvTjLY05GLs51H+qD+sDd5dNDfnFcC7VdSeuSvRB4XBqnZXbKszfplOwfNB6s8wl7
0jcaOmxCrftcS96BsZVMmxkWVA2A08kdweU5TGr03TCagLPKpyBpI/qO+qcTjB+zjaQxUIkqw30Y
E4/V4/6ln8Pw7FEay5vN/Tb0lJsmD42ImaLik5L6yoSOk1OPk+NwOwJqVQwk7rKq8YcEmnPLiLGE
4gK7SZZRdyUVJI1QnS9LkIaX94icrbYfRbpZDgCrhti/R9Qaoqj6xgYCAhLAYjASspVMCdMqTJgl
INQONFdH9y0UFVsIf/QHDuKdfQDtn4TXPVPayOtx1zeHtWZgThonpdvksecncpMrpyHqmbXk7v3j
GzgnAnNzpSH1+P59ZLYnxnZqT7kPajw45kDo5mzBskf2ir8BlWWouL6F3zcuV2Rzf+t+Z5X8rzzy
ckBnWs+oH34YZndtyKnwPxJH1P46XNDaPW/kPvCNjagm6M9lIFEZGULyjqAF2lPR3bR1uGzVDtMq
4NSP2HmITijQ9w7F+HhTm1v/jo8+vgo8+ByzBNPtIn7RjeSnVMwhMFxdBuJACVMkwg5kIIpMZ4XE
IkbZPpFkjozxL/J/AmBHxHI2D9Rmo5T4e4SeNPls8DWcHoHjbquQghznRsIOSdGLVXsD2qTBk1iA
ydZoAcdbl8YhvdqUAE39Z+v/HWwi9jV3m/sItqe5Corx017qN5AHAcAD7De7TgrWaW3bNGfduOpX
joT5B6AF6jw1DWmQZlN2uwvrGeZWmLnHms1B+gFYN8buFHcgmdlDdgtfIuOE4TGRTcCZ8M7KvmQ6
ayvsxDOTzJLxn+82rCWC9N19pT+8kIB9X2NjqeoFeeTirj075IhPdIv6bV1Bx06qwBoKQg+YmnTo
3YKpEL2obogkY8NebQIy31zhb6Y4oak2wd6ekvi61ozqOFMdD7PcJsUkcuXy3xfsumMSJ4EN9IG9
7DkWcoy4BI9JzPw16V0Z1kLowCX+Z7cPEeuuR9yrNRFNhHOpsA6iCMQr5yuQYJ0N45BiSy64l67E
W1oHtvqayhFl71q/Ideqz8Fs2i1V0Cw3QmUtIiU6EC12T20JtVDMLUgfWeFQ+Iuxfhcwki1RmZZY
fm7wMwJ7+8Shysn5c9WS/A54XRk8n23xyX2CcAEq02L7V1xz11whWSbhyPamDl3O0pK1ckcWgsXH
z5szSflmX/sEuPdwJXCl05sE18x7rNcWnMxfmq4j/wI8HBDxEiZY4xX49l4JML8y5YuBNSARtU1U
SZcqVrnWEClYJ8xGhtitA9XyGMWs6wSyIJPRQSZAB2TFm7cVdetdL72AyNdSWhKWoxmXzYOFFy+l
x0F7eo2cuCFtK7inAwP8kDc++pY6D0h2Olw7z3A6Pf/IDP7L0tsbaMDaIGZ0nGp5hE4Fg9OfEIFV
spYx4wnjS4cbSDwN+xXDX2AwWBARmgCsGeF8Br5HWuzQae7bqGEjZ4HkEpM6bzXlvSnK5s5FUTL0
6kMPHIHesBkOpDM04sQcq3LHgoUYy8F7p/il1vLjuHEyikonzmgpOdWnfokQaUlNOorWwZsDcSgs
+d+L82P+MVsD6HK74XYbVYX4sFsC6REUyuGL5WW0jD5+irOV5zNKq1bzgQZGQZ166056rq8uUyzO
rclfI7vmSvwQB1CKpOGGaKP68rJ9hZaY0WmBN1wztmpbPg5c+0mhTnVc8eB6LQrpfPC8F79t2Qbc
vFqHRBi/scuZLmhs8m4lt68uda9oOWvc1UhMeIrFooQN7wv1gkv7DgoD4qNN+XH2ZH7a8T+nrYR4
bdlKaRaLxZLvqnR2iK5WuFBEVqqZ7S2KjyU7dWkpVSNRjpuLEwPF4zBPbqeldTYGwK0337JQbe+a
f0ik+QoxfooT1qPYohDDF6Z3qpO/mgJG6klrVOBjw2NcMxIAbY2pI2CJDebmkdW7FzO3GsZ0YPt7
M8+qC46jNaD6gyayVI/tqYqAW7Ic/3dqaMwqGInJmeVriBNXbXSeGHJDDORmEzcFIt6xao/rjc/E
W1RdxAoRUvb9L/EHNJZmPCcZ4um0iEl+sVb/j+lLboGFTsE1C7pjPXRQDTa1SUF9Y5xlnlxZFhRU
AJP3sH8PRQlf5aDohjoZkuJv6PzvxWtYPMPRtjyUa0vlNalPDATA92u9LmbXyWBXCiJ4ftbfOfsI
KZDYWEflsjtO0n5T83Vq0pmC8PUpXbBTRdIDUCGyI9LrrJPFcY9OsJ6NCv5rI7hkaYvIiqSTIQo6
RqVVvaLo2dKtxvF397YPlxMOiCqwPLwRl9H1mudREPeWYsY1KGL7n+cmP2O9v2tt9vLyVFEAgX4U
4OVmUN+KDxpdtDDHFQvmPLnflXE67Ulb7OahIn3r0k0Ofu7fy+N//7SNIsQNMf1R0Ak32hCvRNM4
CoNXmNcSdr5nfvv5mhBOo7hhkD2M0ARuu06hTE5vx0JdNzktisY2vb5F0bZHSj/3EPEq5dWyxboc
K4BhI46Meo1bkaqnQJiYvmmLNnj+TG69C1Y02GccIrZtFD6NaulWximBnCkbQtaXFCmFn0gWc1kA
vHgWjhyNYWKOhu101vPc5+GqfpHxak6qMdzFG3yBYnCut7jTIV2XgEp2Uaoy6qThBTfALKGXq406
m9hYMXkpXOY93eHl6B+63rnAb7wuKzgl49b9CS4MDB6jwQD4UIoGQWoGYmGz07cdkOJiSB2+nkKD
ZrLLQkF+HOgmen2UUv1M3U25lNQ+ZiXGoCvbhCw9HZh5AynUK7FvE+tsujlc/u2vvq6hA6Kizbwk
qmqjfZAfey0X6pLW72Age5iR5dAQ9GUjKpTVqveQZz0nyZam68NWZrMnLXfVocTZp/lccRLqMfoR
ushtaFIkX6lx6tEpVGaS03qgz4NG3ZsUf7nQOl0DlxglS3wwbd6T91+gF7KSyrMorEOc1WmKkb0T
nxUK6gFwbfoUvQbfsVKhjKMEJWCa4zkFeysf9FKnIVGqQXGJYtRj0io/CRaLKKt/bcgRPmbfYt5/
zVybl5qa6zNbTGNMhBlmtkg/3s5jgzzMeJpQVM4JCwFn47IkaxWhWseBD1Nu2BTypHAO3Zy2qioC
x5/+ccMSZ1MjiXb/KEqIMFRKQqseHYbsT8C8mp/vZG99TbPjs43NAj+QqjOwp7N8thSpSiwtgPWL
Jc2pc/+x7YI6gnxEIGh1l1CEhHZes+W9bj4AQuJ3Cg8mTnNymm8meB9KVBWxi8RDU6Tj45XstpgJ
3dFNGfOENgYcywr5XHNeZxNT5vrbeXmUvU2uQa5/xjcMscUHBjo3dM1xh8md5ZuAEoPdl4yeh8ak
aFUyNpAYzRM08oMvF1Kab5EKAfakKyB2FTXwiu9H7lU1GU6T7R30ZYQcFyRrM8JsFVOj/bum68j+
XGnL43z2MkYYg8Jf24asM0Juqy7+ztm25MoUjmADqhkV5dFO4xm8rqSKrECXISnZl8PulyHDe8mA
h+KrxndMQx6ashbiVsoBD2Kgf5IWsnvH5iIocR5BsFgEU7gMCW8qA9KaowNEc8Gx9ygYrWbJe1eP
fkRjSccGzQ3ULkOdsNU7elf29mAdLpKky2vnaO9X/McH6GX4cyFqYXF1ur4KAKlUGfE6BL7w7ADj
FFc6PERNmCH6OQzmQ7YBA2JxJiGSMYeqadoxuVUnhcZhryzyNobpj+HcIWpche+1YVZXHIXrUVyU
3HP9v4GkuX9rV8llIY+oXGEGnWvrYpivoIvTsApxGrA4XTMCrr7agUTBtflqmSRTb4KIEkVuV4rT
bgmzH5Op43IC98GZLJUWkZmmPRyS4ERm+DX1XutGIQDs2alSiz22AFX2XjDGw2mpk2OHa3DJV3wi
lrBWsHg2OKkBpIMXgp+VAZcboItEbEXITos41nRpjEoY9TZlq+f+nzm5BixIlv4iIcOyuiIMruzK
fRmrjfxaBPkBdMaj0B3ET5FOuxFXTElqaXbl3odHlhMl/h6RF/De9E8Dsyy7bCnyizVFLMVLCfAU
h6bYbKEmssrelQsM9097vVY94AFJHF58tZKWcujg0Ec0ulsx3mdvo6fH1R3QYbeLUUQ90i1NDPb8
aSuJLlGN5KXXSVvvUx+8/Zv88OutChOiplgKGk5VZHmcCKYBVXPwF46G+8HgCUVNibFhaOyjToAM
DVojSeSAO89hmec1T3M0X1NwOYXlHJ3EPdb+vBYxGcZNdoSqpbnvAYkqo/4+3+FwoPkAAHwbNGQK
bmGLFYd4COmxKOATBCNfhP5iu7tWCw8ZwOUqKkhP6sWy3xuWNVD6HbOp4foCcFhfFW+nibpDsHvj
02I4mEmQtWCxv0chObNniVoEZHER/sGbG3u3nFLbnw1mTiTvHlctzWwjJ06D5Oh5pZJk7Yyx12L6
7ezRNt71i7THoO6FjdRVB02F/QxR3e+unSrHUmdbe6K/nt0BUlG7K1bOFzzu0RgGh1XvVLGIsOje
KnVS5XpkE4EEyCQ//sG6SlrojYLL6Os5/9j+8LgBT/FD4Ec/smIRFwytdOGNRPErsexGGUhl/0QD
BaD16yO61wp/0c0adZsre1MQWUAIf0dPHnLaZHomtA6hlQHNsWAWseGyKNfD5DUakzjAM8vwtSLa
LqqEmtpbyLDobP92eDivFDuZ4ibzkGvtB49tdAI/6rCq0/gE4QpBaf1NItGZwJbFqkYywQZwU3OS
/3WkeGEjAkOD5dt4lqjKMjHs4wfbvVFCCDiNpQuupSL7e9ErFu5apldFeoeQP2e2w3qjpmbZVqzG
NdhD26mNl/A3GYiVia5nJi6+0sFI+SZLowfKuEKlwwojnuHrAqekX128a1ryR79+ATr9xJF8oqIS
U+3ssCiaJfGRPwdUB6P0EE0F7ajocXO9gW4v0rFPEJQT6khUOwLXeG/QvpVT99W65KxECIiQCWnx
UME8WtckbLjpFKpBO3WxEajappQ4lLn8gOgfW2fVDhHMVM8618lMjE/NzeRwxggiIXMCerTne56s
yLCYW/W9XROQ9lt0Dk/OHiBdnU6aDHGgMujB9bwYMcq7zttln/zLockHG+wgsg1RNlV2kZgOAmcr
2Ft/groJ6nGYQoU54vWBN9oF5mQvLz/LB2L/PqUqoelHQ7cEsr+quMWnBU/N0+gZzbRG/luTAzlA
pIR4BzjXpsCdXrq6RR/9YrPpPWse/ncXLZNMmwW5Ve64NsBN1jqqj85t/2oyF5DjJXgXpW/u4o9x
Fzp3FmscGdXOI+2uPRfSLjecBZAntJpJmubx+t9Pe2+zj3BwGUK99VL1wOi1nBMItxmFmlnRT/oc
cdMhFKOf2/oD9sfYyHsDXlAoDoKtsizuVwqgtIsN+NOl70GmUUiJb3kOcVcR/DnrFXVF/TSlfCHE
EnKOFCxYaZo4WnldC/d2UpG94pIy+a/shdQ3/ca6yxJZmjSr6npgSw5XANTGvkghiBwVBxdcjA/B
bAGbCm5fARdaIeYKI36W/eDm2jimV6b2289dkVH/ABn8dskfcx2dMIhSsNAfevQSoj9ZZafATblK
rEsRhdl3b9+EN/S2bOqfAMLqVECfYmw1HKWhk8yb5Yco9yzv6irpxudvSkeMKC4YBCCx6Sq4B0sW
R3hl7Kj4vEXzUJAji8o5kh7sQWHtuqynAe9FcPczhP/YIY+K3/QfWiNGp5nFMGCNUszuSzFEB9qc
hdHbN06dFrgDD/Ot4omTbNmygQbkts6wgGqpZbWHLt5mbP3sBc9bUl0GCZTPTRLJ3a0nrT3qcQuo
wRao/uQAmNBSfJiqeiTDSpOkjmLlF9H6H7V3PA8rDXnLwQ2ToU+QyNXRIlKJ4u9o3qVo9qBJ+NZd
1gNRgX76J11VpVeCs0lwnUEluX38xREq2b1cUl+CScn6MKAWWpKMGHYBlukK3BAsh6WoOBMcGyy9
jTsTvIwAFSGH5sstVowzrGA6o3z5ztNmyASrQw9RWiVUsqBXYkZTpcnq22kwPDvsxyFiTSlB/XXz
M62hWm9iZ1QOTbAd9oaZjwS7OTxhUd+4bxvLNKjknkqYLu1yVsX1BM/2iqmJiIIkhNI7TNROqEY3
hY7Nw2aZ+AdE4NHTtEgcv8/uSwhwnFEqBLU+9AiSVf89zhTDTeQKWbfKqCmlsoyFGNQLmG91ebIo
OmseMWziiA4Z5xSa9HRszl7r+6S6NpIj6fgERYGzPgsxzTbk7ixznhWiY0B89pNl3xNVTxV+DYRT
hlqTmiR5KbgdopBXR2qb1JtsIC3lZMzvM4d6FmQfZQ7Qwm1XnI7C/2a5tLubTk+ZCES6l3Sx+F2b
4jMDbEmcj9I1iRwCNYrvLGxRwmFPLWlzEdcTe87LLckmYoOFOwQIjYwYTPl2lbo9TONNupk9GG9H
WdQxhuEyivKatJHb2m3tbAGs09NehaN3D5kQaZiSOdaQWGTRVM8uLrb9aZ4DAC1d1lumMfh7+iy4
DUkQpk42lnITMBrlaN8he23XkYAeczAEmBqookOR0q97XaTpHj4TQi6O4fhOCr419bi38ymF4Tec
7+M7OT3HM0XmN5BtfsmXNvViIgOuB/RJ/PEZp32lTbrKBJOILo/YxVyO7FXnX98yhZxVMITTTL8i
/KZ1+G/u5FeZHu0Dfrmx4MnWfS29oxLLMpYnjva8O95y5DQlU8RwqQsmO9i3nyvaaFhhwLZpU6fF
aVQNSrH9u80SsrbYEKSoRvQsUwUdbttyu1lSNM3U+cbIzLbzgj4st+haPbt/Q17g8+KRA7MAHfiW
c/kmmUi8WaJKIQM+W2ZgrH+tLpWCqTMhLcS/tO+4S7aYBgMPL9wmLF0PQHOY89DkqnCbX0ewO7wX
vL3GbYKGPl+YNZbeYXmDkBSyZbItvui2K7xiNuE61AE8107/Vu1dkoAtLdy+veMWTz36prQBRHRH
5fqHQ/rgUWq3uuogOu+3R5U6q+Kob16PiFBwraK8bS4E8txOO/0Xi8upnP5oMrzIDOfmYF8rT04N
nv44BTR0seusGfmaVfuFo35vI6Y2yDTauyxiv3npGLMCNILPkO0xfOUrcziV0eEfZ8FQKumzqsA6
nU8BgJ8EWr+WUtEoa4rHJOrBiLGGOVDpITc0NWASjH/avKHmb3P7V2QvpslM1P3XrYQ2yUFaBEJ+
lDRptupSnnguvkbDe7AZ42hS4d5SClKUtACOMVJbqqADl+8ALU0oVWb0FVotjij3eF1kmAvGt6Qg
VBfWjDynrrdtLD4qziUMKXr8sVfz5nPjrJmh70mto/FkYrlaPEqaY+ONMV5nMvFlrbcA+d8NZL/N
Yh+XRyhgmQOeJwa0CDYRIRUTWrjcQX1/ZKsPkhxIGcOmJTzDx4JLOmy+PMHDTLdKjiuvC11luRD6
BNSFe7x0Ng9/FobYlbuHvqVTfYNzSLtiAWHHMDNCDPXywQ+jHWmqtwuyc7hwYTIB8cx8dLITzvUE
/WIVMNWZD4qX5irsp9qWmTzwJUTApCefnGOBku+dWLViIObsk0ayexCTh5k2sxDCQonSI5Mdt9qc
n3cIr27Qr/+YzxvfDIuywqfHxT/AOKGwpoS3Hr/BVoa3OD/+mf7NyPxeAEBEJrkKPsCpNVnkBZRr
XQHa0eB/h0dbvrJ4YITk3XxBNRnVwXkCyDKsmIFyg3w5BW2acyTFzBJ9Q3ZJpxMxbvUBqEPNVrlE
w21ldl8S32KAubSDb473gtLwvY5xLdM7xwixnIa4WobeL5XTgocqNdKzf+HOq3tA9bQ1rbUCXzTV
94WxrlNC1mFzqksQeRpql0L+Zd72FmIYKL+q8/Wmpi+PALG+lpQDB5YSfMzNwyYT1vWnIA/3Ymbm
ydx4Z9mfXXuucmOK5LCVZNy9zL+qfrPW6xZwhW9WwSukU8fMWa72b/lrRRFSYpIyAD7b515IeGED
ir9m21m+RnybVBrd8FLZFbsVqvrGkkdNwbdpRgkH0mcCVO1W9xmpo+pTcwSb5YkFMGgJG8a9knRk
KjHKrQZTpsCJ/wFLO46WVQsfQ5LoL/T2fxkINQjTXguizKhmuNjM3u4dSZ3eJWg3zQO9FPfRFueQ
iXAmvz56rtE+8wcmGx5XZXri7Cu4KSU4i/R1+XwiMYNbeF7n67hz61ibbTNBlwj83cNFnaEqWSAs
tHVvTZA89OUEDC3DL9m73naOLQ4m5xjWuRjgAyapu1GaUmwAw8rgIG80vs+BLBiF9e1rUxWjF2XZ
VrUVw/16DJPg1UUyWa/pNcGLQR0cg/TzwLs82pJucHzbOMfAyP3zFbBtiNBHQKF56AXkCAWRB/s6
uahZuf33WTeGl56qH/sELfEGUl97ATj0s9XtPJLvBMI0TLbEdYUuZbcMqg2OMr93UrBFSoECA4kO
VJWeRw1FafX7V6b0t7f1I0r5KTs94p4AZzXBsacGpIRy8OmjElmqA5BG71nKlAC84FaYwvlFXvw/
HMWGJFNrIEEhpV9d+/i9oP5xqIzPUoKAdizXFqSmMk19qGevstdVyZqKyh55seF4iOqfcjBDuu0e
F2ZeHUiOPIx1taNyeFJ96akf2OqzCh4zkGrYF4L8LIRpFtdEjPv8nGCW5WAdLY+8Na8IJUYgTUuj
f8/tzlL/Qk6cNKEqs+TonRLcIX7WttAiVzQ1wgTnVc92n//TgbOXYfWRrMO2qo7W7taHAfgaJHwI
5cf27TWB6nHj4zUC5KXiEhTGZ81NGOiYXBz5tKDRSWZSLJZ0obhk/5LbhwlmBB6P8Ze0gFWHuyeL
W1O6T0jBI6v4zJAOSgzHZ3pZMbhtf3CB8GQDQjwD/gVnAWFyCwdH4ScB6oM3/XIk+748zeQh87+Z
pMLnzCsyo/fWkyY6rkyl8dSdiQu1aTa0+NMM2Ow1UjGGnskQ+dQcC8JBQNwfZxwqAbD16mCqdy2O
BFQI7V8zpusO9LfEkfuIg2I+Ivt5UYPpmI0jo6kLRauIVJXp+WPEMj4hf90ytOh01HREIlhK8kd+
e0UIHM9vu1ppaZnirlvVVH6IdYoCRHusNlh2/eNEyLob/vlpZvQWb/eV39LDhS+7+RExR7CkJf1J
++7NN3SApJHw3zRYw2vZ6puycpDZjHHFYzlCiHPOZWbtHe4YP2hyRAb3cusqEne39j1TbpP1+FpN
ZcPxKiYwLc20Ds6oqq5/Gh/FZilztWZ0OyIAq321EMZCoyPeOr/gFQSgKw8NvEVu6mQmdW+fCl6Z
MnUsvJ0d+3AfVnoNc3eLqa7wC9aLrGzx16X/CVTQcYyLURvRYoCO2Xy8ELC3jGUtRYMT2FlxOAlm
JUNrgxSwG4b2cqG97ti5hNL85MdzUuGGUfh8ZAYufII1V64YkKaparirh562ZZZMsUvCNwaiIIyn
OzKqQLFpvbUWjY14i7nEL9tBE8ywIv+v5TZ1a3m2NtfVRgsp4ErQPsMtI6OKT1tWIBPSRa9oGKec
m1B/LZ5GKumM6IUUINmzWfq0uuDD9LSVGaHn3LY7njntO7sVYOhWC6vVdNC+T4ptZ/puSmk3PiuF
kqO7ib0sGy1h66wfholMzKoV72woGIGiBbtHYGT4qb7VnRmnEF+3mGoqPDuRuQ3dO7i1wIGu82bj
CA/sHqv6SOJuhe5tyk60NqTAcrteMjjf7zuzyVVoSw6eQScvd0cBk0DgojzVDx32kkBXVh2R+cnv
PTCrLmisoYcLWtrrVC2kKwJiZn1WfOGG5xwPWCYIaCFv3CXG87+S0q6sywj+Afdqkw9occBXwWmm
IzGfVhF36fy98wg1qolVz0nweLbYs3713dnJtuyHR6QcMtdKCcv01nv6dPs/CKAQdYtWucmc3pc1
e9OKezt5Jt5OkX2DFs8K4UlXyHXzsyctKjf1Qi3QMwzdwvAeNPoPkKmQ0WS3LOGVOEryOkulbPQ/
E0fVFqlGTuZigUqAjok0Wq67NgehxYhujq1HFZpjzTiq4CqND5oSmoAFzQxu8BwjILPFqxZwaen3
XuVuzTSv1/+0xQL3oowcz49Wy2sRwAjy97hRBRHHgGty7xmsEEtxm2UWJLtpgih/XQJBtqfIFzKU
42JBGkUog6BIfNY0NT+UDu7dnQR7wv+Ua2UV6xkEZqS30Q7QQ6qJ1+cHeT9h+4d62bl6W9UxB/KA
drc0N9gPs2aLdHhQVhMtnci1u5sVqcKDw4UKcZAAv9Dnu2irL4fKj9fBsmu9IbAyTpfWlwD/c3XX
V92DgVxkSnU6CmmgHVwsiLnITtT0JJeY9EmfQULvSgeWfc3PU6jq/qZLGD5NF987YTeds2etsf2u
eW3lS/yZFKGLmvRo8pd8s67JOsm8CxvVr2qap+XmFBgbvTmSTVuBMxjN6BSPKnSFaHadDBQXmAqH
sJWIte0W1HAB3HW/Pdj79XTV5ofSGCQ8Z1JJpcHIsAAwvoE5tFpq5LSlsfsl9cMu0ge0zpkiwjTb
UNEqoBYubBnH/rl84NPXJHcwZ3IsLDQJo7B2wRCZhETH+e0X6nX569acZcFM5wEFp52M6YETiV5g
0wNdHiL0YrPTMoS9Oeff1FUTnovGjAYGjA7J1BWx9caFGIaiV0bLGzWGzGRNDJuIA3/ckg514qdL
hgYjJ+/ELnlbPMlJkfDq7WxbP1n1CqBx1sDSq6jgURFlVCe5xefMf3m7fxjUNQCvwhLio/3URquf
rysEym/zjTZHugtU03A+nmMfoCjrY6OfPgeWrWOH0VOTjwRTNqqry9geB0SK3Iczz9IivYxDkmZd
JKz1WHKlEHgKnRHIZJ0V72xZ+EUDT3/BprmaSRg0mh1bKUvhaeCnLTv82Sxu5DKof6BicID4eJYF
VTd4l359gthZWA9JrRrlATi5l+75DuUWzE8drWaGJ6fQO6mCJpkwScp/rk5pczBysM2ZFtKudpLe
sMTufxg9JwSiykYuepuvSTqnqLzRGxjtAwYuCuBkbE9UTTiWorrRLd/s/Fpp+xOK0lmwrvnHeVlN
C8Mlq2xlzlm7ke0RcCfVOFMWb1Y5UYpem8zZMPLSA0vlJoe+aSO9LLLuJi99PfV0w1gA4FLAa2Em
1TKCkoB0Mvay9VX6lqMFJcTgZB0mC0tZkEqnr24V20GGYV9C6NaZO/aOY99BGBtdsek0X3qXcq7S
q+Vf5uo/jLSjpffVQ9Krg/sIjscRIK3aV7kl+9tNPgPURLGvxW5+1yf9nNpi8UMhfy+62AgPafhV
PRc0rQY3B9iHylQI7YUaNFJoRgIJtX0XT2En8YevgfyPtMd+qBFzE9XyvDBchq3aZLg4MMAwLO4d
No86nBz4huRvFpxW/fWfzj1gs5ZsIMLKI/IeA3iAIo7XiMR2d+c2FXVXgZalTJE774g+KS5G7SMb
4mbj5zi2mGeR+ysoSYnBzF0D1lryTMEswA1fOLcOmPYE+OFndo4qHTf6J1eC97SdPoHrMg7ET55a
nXRQ6xFniRBoAw1DrMT7wjpZxRxlPGR+zl2Q81xae3pzQHPIBzztR3sbktBUgzTqtgeMQXULhDq4
YNTGhuktXkL/XSWpZJDL8f6K7pxUE44fQwMGZWpMQVkBGHSaNt6ZL8aIFIeETQToWYqHJzPQ0IqU
yi3mIzjGrYNBuQHjzEmS0jPCxN+7qe9LTEzygVXsUSdU5TS3dn0s+h1RA3ZLrA1DBU+K9QwosQRC
jZg2uv42KKhpgPrQ9y8XnHXhwQ9ZvxJKb38rWD4YbwGcsCKwkRQxmOWHKx815Cyt7W/Ip3SL7q89
WFe7waPjJuxOVJ0379bRBOx8erhiv2A0K6fZT4LdkZMjkipAfQCavUuqtwHfXV9EzlEG3j2cxjAL
cF5YHcmORckafdfIJY4mL+LeSO1JkvF4bAmRweLOOdTQjlNpGZl03Da8vB/QLV4k+uLnHEJtTKp3
95TBL41a22U40w0FUhSwVoCevI6XzDZI4N2RmIzCwEgwjWhpvyHvQcMNR5Xuq0q7vTqfg7GbZmh1
m+vFDS61cu8AMCVq5xnbB5uR2QPaX947OTKxaGqxsCeAcUhOgDZ9MAIq3qyjRjH/UW3Z2i24U5X9
d9y5bc1KEr+1zygAaRRjC4rF7pbqUAJb4FlAVs2rW+sGtYS6OBzaIRyuSYrF81DB8/M16vK0yhIG
fxI9GwXFyHVlpJIvlX0+JOD/DyVx8lf0Ya65jjXqfqGchrF7D0phcexxsD1Ly6hLS3yIz7vwxdkY
1DlQ0tSeK2bcvcRQPMRzvJ2xxGGgiTrnuseHlUKGH2QQi/R4mZZOryv85ueyNTp+bP1lT6k4riG1
fBM7d2U5+a5BEiQkmQXqnOeN0thQklKhGbbawLDaETq1R2WULnKE+m6KfusvM2hLBOUQodxIo6Z9
GqNkuLDUwk22IjXhCyR5+T4hiB7rYOrhxIG7KHVNZXXCPU4s2ote6uJKiTOuKiej8cioEmF0JL5N
K4D9KWyGBqqSQ97leSosyApMrU+90oGMxnSljpcMKj+AUcN6pCdnctKey7uMBUQ9rgBBac6e+1EF
W49uxNaVeTT8l0K52Bu5Q1X8wCul4RBC/J4LLq/F9xszwG8JnwtvU0J19k+Jz57q0i/FTFU50aZl
6yfu/PetwbQTS4KuSehSyamUIsMeGJvereeFMY3LmDSynqMRBaegAJyK9UMJZnx7xwRqB5COpoF4
2D5nMs3lHDomdm8iOjpKbjDgZv1Qxa0HmDV7On0Vxdr5I3oRM2nThT/fhXCN108bHe/Rr3QakKN4
g9ZjyTCahTyBASwIEH/j53cQmp+07gOiM6O8Q7I/q1VJ7YPB3mnBKk/10eayAmRkJnljEQf8cdrV
s8hhOk0WTAB7gleRES/pSpwxI6cdXlwDfZWFbnv9h/OJ2JPW4/NRnToJ0/O+Gmyu2GC/6mRwws/N
YJZ+kitHSDxBy+zNJzMb9tuafUMyTMLbW/LJ0QUZxWBLh394aWW0dDWGUB7SG5IGs7O6bp2Bfvb6
VqGmlT0IhhaljIR1QYYKJ7E0bm6GMrJfwIEqkU+S760Q8nLhX7t6gqiBe7laXi6m0EGSbnfX9nbd
evlWMYcQzQgA7X57y6aWDz6QLxNntyFCyMggxQxY9cDFQfivunP26e9Oz7oeC05TrNogQD3c9MH6
su75Y1TkxE1kDDhBqRX2E6eUESV0kgrCoSaFQmrVKVZgsjhy5efAXbCCu8rHW66gCPxZ/0YpUQDi
qdq3GtHib6xD9XrgQL6VSkRbakCpXnsZ+L/Kk9T8XJHef0mtp+xHbGVvDEskWvtzGeYxsEzbujXL
yv0Xi0O3nIsfCK0mraozgwJ5X3J7im2dQ4JEXZCkx6jlGGVjuHTkInjsByCWpeDWEh2Jn66epufx
zyVlmx7b8Ju5Mpn+myTYs4zgcHPGj4heLaIpSBkzx2UpN3N105VtNkaUOI5f+nKs4HK2IJYOfSB7
d7GkD+rylpu2u5ot6BORX8mMIJgbzxr0pEjmI4EQH5Y5dQfjrxWNDhTGwkgx6M+/Gc1VqiKhDPfM
R5Aeyui+f0yMm0Xps63zO0xlVu9EdMBO5Gxfae+3qU2d2C5euxKu4CJJNWuCOWN/AGBuWYPscj81
0RSTl/I+iqWg73gU0D8fbJB3fCpkJvhxUN/TDgQP/g4gf/wOGN4bBNC9S4ORbMEJKrMzRzfrACkj
dyyQJTAZBMtllzUOjFNTbRakkWNCVqkaYWovxRG7QhA84CeS0uCgiPU1Uypfv+0BIvMcCFFU0siG
l2CfCGA68fQKAPtD5BaSEXfvuhvZJAFzC+T0Nan2nqrFZU0AIBQjGPvIS8O3qo0TazccmRaVzm/E
MQiQSRVJvIHX8+12GARqL4dEGrTEyHd/XQq9mmRQ1OLygg3FdNxJnUlzeiuGzo+IBFxiZBjNwdVw
Md/JKCQ4Ld5oBWIesRPhcSYk6Is/JxRHnBbktC10U2SNV8tmB+DoSKvLUzzhLLZahQMvuLrCJWPz
WJBcYgB1TOqK8y96vlJHBZnxSZkgE4HwwSzrQ05WvMyJJN9Uo0uqW08yYliexw1QZCqzPoG76EZh
87awNBPNOMylEtWshtq/ipJvQ3ppeLKzFM4QYscFWsj35DujVyNErKLzCxTe964Ni1usqNKE0O1P
sojts5VdYJxKPvG41k11wwRMF82hFrDKoYrfEeOcV0uiyyWA30EOM5hg2KgfD8B44NHepWvhTYAh
c8wsLcQlKfjaITFi0bO9sMhNXRUcP9H+ismQmWchXAbgdEhtUgjAAFXWqNZoz0RM1QuFHo/FB7c5
jG/YYRObZmvVesy4QXprHgNKtyABZoohPt9MOS2h9miXj0LxU4qIQb2/kBlCR/TkPf2R/Nrj6cD0
/bWtAMZMCVs17EEMbWardGpM3s95KqIrQZ3oMxjfm/rp6rQUDsuLvFbOSiyiPuzMI91B649iI2K6
Y9zBMR0aaIaReQZyL6V7gQzH3c/ucfugAHYvR637iSpmByuKSh+wL4o8wp2uX1YVaJYva93+l1BZ
f3pyGF2O/s2fsKFLS2hwsoF4ddzv2DHQktRPIOzUG4NybnSfkouZlmnSGQiDyOraND6lgnhb0e6g
ww31Oh1U5vn+9/Ayujz68vc7/5WygI3gHtCcH9vihOlNS4BfXCZZac2pE3wYjfAmX+LUorluZOdJ
YN0ywNJgl/9TnNZWv4PQSdewI+WlsFNO14VEcHIgmpF24o0yAffr8PbxEJvoluaTFJ3UehYhOC2d
ZkB23VSrPuVjTUUEN78iqpIsDo56akffEvcUu/f17M77O6Dos2qdTFprNEHT9Sq3NnaiND9Ap2Hy
jAX9ergSXoERa7EvCix8USxEwFwVXigqfivDI0yFauSN3+KHbOahdClCboOftGyIOKtT8jmZwo2p
B9sPP+/DFKsmey+EulpAEDdfqLQkEmUo35hnFE8HeUnEVrU46MFFtGhuQh2VpAJk0K3u9E7v38Iv
jzQsawKicSLjBo7Js5rKrH1SZZm7yv+GVlJpmWNkrRbubdsheYftQzNPfGRLlSnCPNvhcHPAWfYG
6yWvWdOmCnsRCBrEeQszddRJuvPtgJDoSCf0z/qa/BvBFv76rMT0TeKrvfGosyzvhipRzO8AyFyP
RhfwAK8Ek8DGaUfaVBq5sLIm0AO32IbOMiOpJNRwe6kajN4VB4ZZXC5KH4dBGIdZKhVR3rSqaBbF
TiyltSP87OaOKRT7n8uMN0UUtZ2x1hkTiArp4FGKvHeRon13a4CyFcgb9c5gt2UWAYe8sTC0Df5j
L3QZlltxXqeNkeN6Zlbq55FDJLfGLgi6pKyLQiMiLH4qW+Chm9Gxe1Fzn0HA8DZTCgV8go6+3w2f
Qs17FMqQkTiQM0oAsN4MHsGopI1rtCvhs/8mewOW/GHtmsxm9wp7Tg7ioNG7rxbfkC1YK2j+ZCrT
F5rNx8sePG80dXL7H2XT3iX1bbutNDTrewfjORWeB0b56SqulRySL59wytsHTGYlMU1fgXCLJa3F
JgRxtFXi3dBGVbYXy+P0U2bshtRQ8I24vpAMiTVGLbqtqXxRUz0Osmw5/XXeuyPpKs7T2v0X0xlD
oit4EnR1eK4vtqeIy6pMtzmUMZnDz0FqD8rttkf1us5Ia6a2p+/Ax2vTIbH/zTz0tDnAlL6nKdxg
ur3DE6vdpWOuC4TyOsJysB1N2MF8S9MuaTkPJpmFxCmeERqloLX3kqRHLHyciVPd2PutCtBIRkMA
57XUbpWl+yV40SF749K3q+2rTnv+dAHHSuXPdHh8tyY4Rys1ZiwpnGomZssEXMT7/FnuaJq6D4kS
ZIP5IFsXOh7e9FxnQ2pWVgp/CfbJVirLSoS2dQEA6QNyWs0W2PyNq8fOA4yDK46kjxQdrSa/S4ZG
6xXpOJMvS4yf71NZXbfgC0G8rGJuWC1TacONiDuGNmKnHhjZVohkOkNYFvkMniGNFyhlyn/I7WBg
5YPazpkRGWi3zWFVgolCfKKD5SeRXmtu7gHPB65V9Y62iTIWctGGw12+yBua8vUBSlZ0ZA7TjE6B
vHxpG/Z2D4SZ4hGVx5qcN2FwKBYRwprmUya7BoW1BmaQ1/9sHyoXe1idaa76rUWUK2piyWGhFdUW
RxX+QLpnZecV1mTk/6ugo4ZD76MIa1Xtz1FaCWuCLswQKCwc1yoz0aRRflZ0w5PncVhFERSSe7ol
jBKuhZoJ1efdvlfV/OQGpe5cg6j8tpVEJ47EgvXDpCYwJ3/1/CjoGTNxyjPk3X1fpfWOS2b0JNwZ
J+VUznThzrm9EcvbNlE5rRpFPzPdmw1jZ9J909yReaPnvviCgLkwT0uUyb6LJyfEjbH3grSNZpH8
c6cCAv57//qEMsBpeH+PB2fAi0bnYexaM44F+1Pzc5Obp6eDnw61MsqW44pFFIrc4TvIq0MOK/SH
5aKdmE9UBkQWYX3R/1GdL+D5QfTqwgPOqUhElkGQ/rM553OTi6sSZq9us497OgfL9VtapghshbBk
TaCIwqIq8EuelmwkrcwXSs+iR92fZgZ7UysHPkdOqKP2mNfovcip0uwc1q8e5oYSr11ZmtMmAnkF
BXFGS63WQR45NGiHfnonvy+fur4NCzAx/bjgNyXbzOiJ9xG3LTyoYMu+2U2xQY2jKQveOi0Y9DKf
NISRLWdLrsyS4m2PqTgGhsO5iz6GDx11mqUxZMVDCLre+FTT/cRW7uR43xkAm9vkGPZCrdR/YQr6
106zReUzCrWWXWyMlM7BhN+GOZA0GFPFPy/MM8mEg5N/sRsfEJ97R+4NpxKO4pV2iyR1H0EnXCum
R/8FgnnCZFTVDHk3P18fJr8QRzNdXktaZEpR8riZHB51imEr42xcbhibXXNpuNgZ/4Z7dODAfAXA
iz7j6wsL17Whz3+JrZ/6ILuAHyERQ+eyAa2FhePIDS5H6I2Np3fU0my0LXjtz0sdKi241a7OJnlh
bdnGoyO+8Qam/fli3fddzLHe5vO6OjJ1ycZQgD7VutUL6IMVArHB60lNVocjV1jYNcm9MvBn+1JO
OTR3rRNkcNeKqXLWpm0lzrHhccT5NZwAzMy3qnUiTA53gNH43820kFx1n0NMIkoVh4V7ei7TdInq
1SOxX3x7fy7J3Cp2ID8S5Ss0INX9Gcv/YxBKfJOl5Qa+26ieikwERvtZyMEs3wsJpB13URu0MItJ
jPxov9HCbKiF6MkkQML5qUIkylz+JgY/JquxiFY3LXiBIL4gAu244aNB5wPEqX23Jvx2pJGbZCPb
l540YDxYZh+y/h4B0FqL7Z57Q5/+y/oEyVIfXtQs34OdWIFAAb+y2RL0SA/LCHbKHu0Zf9yr6onJ
CjjpfOI1tV8c56BPKugmDqUYVE0LNN2lTGPw+/s4dmpi/CVndQpDCFqYDjgOhzuxMTFWRT0VHUtw
HZvYuB6ha67J7KwDL3xkwEG/UOfQpwNszBpU8sBPSz+zxKPokJFkMlJYcwGAhuzzWQMYOLUzAzuQ
l2817BNN/6uf4D8QjUMNBqZZu24BLDGKmpoeZ3mVK+ben292RLH2syEn+/D0Pqh/gVmmpvPHSdoL
rbYV4mXq+5LC/1a0RMgpijT6+TLuawD1O3l3PEL/2pVRxkq9WjKs2Bu8PYF8HYK4vHwYvMxP40vb
5n4RQPHfmruRR+wOnhS8eyEhcNJbvsPCsL/zypGiq2a0AxtptxHCZxjsdTsdXF7EKNDLwaUJGnlv
N+ZOMxJOqGJIsNQ2D20XLk1+jtAfIE+rqdiflI0RZwtx6ZnfOKY1ql5RevyQ8FkzEm2NvdVuSRQF
Tyb+E2ihHQzYyzKC6TZS0+VLAaaEtzmeN7tBNso2U9OiOB940OdnKxoqeVjtPZUwKT9QRX5CV1Mf
EK97vST0ZcRpjrMZ3lI6nqN85siQg4OuiQRGhQmG44qj5fXQUj4SrDCWox6nBnHWbzVpuhhurd7t
zq9AO0Kmm6HL2A81FdS9xh6NFT1Zs9tocTSyalqBgh6kqoMxSkEntFaCadSYoKIs/MIrVFUKleTc
QkL5pn4Wvf2rowSYQHWvDvLieXD2SKNvnFBiKBHJO5P/PNp+xXl5NJzyO0RA0YaslYlD2q82GvjY
gD3AoRAGbF55OWWsuz4yh4Bb8lhDrzXl+gf8PSp5LkSmZ0HznHgkW0YetJPpFZBByfTb71+2PRPY
ATCmv8p0LqKebCSWKfFaXXAeKaYVqAtbW6Av20rxAqCgVHU5EPgG0LXUOiZWSs6PeOrozjAeawAb
cyhpqylWveDb8otX/0oNLfvsu/Og+NZ0d21o9uK4tKQnY7Llvxr2gipAV/NWecEmbY9tyVuhAcXF
ovWVFqr7tx/74/yYRfhhGpd+7EKvBwpmR0rUu1aSQpqgTZKrjC7+XvJEMjTEOE8uSeP1FBHbqbvF
6MPZCxzCHQ5JBvREprNX4pm4oTakepRsk8pVsuuspP1jBZjANuZpgQfclYXDqCFCb06a+x4o37em
jmN65EaPe464pSCy6ettNv4yEha/GQQtId+XjDjlOzmSyE3xk5WcQOWCA61stNgJC60UAuY1LaUD
aEUxstzeWQVoZdeSL5vlOxzdqjKWACIjawC6PEjDsAktHU7mmmVmaEK9kD7km5VWLN1mdbc21x4K
P8FWXNstjqptgXNd3MHxjeixEHGWbXEsGaxrvr+id5w6AQ/C6qcas0iJ71LPMNTs2REHFs6dVkS6
teeS89SaBYi8ZnNYhSUiPk2iGvXnt+HqdSDFGJU7KX9CZfeegjPdmpaaOqUsIIYOiEORAIHGUwY9
G9RtwurBu17F4lsUihtZL1/+P6px/5oeeoholpL3t25Kfx2ofvmgdz163q/dsefgVGLgRHuxh9q5
FTYZvo5JLfgYfjXc2JFYD56GfvNbKSwrRkSexWXuEi/qiXaDE5Yr36tFMEANS34dddL/a6Fg4COL
EJp6R92fG/KtyFYin+6YJt1aQW6RBtO38GnLeneoPfOA9XnGUGJALLDjgMUpp6uIktEAfu1pE4jq
78xZzjBo10wqaSwBN2xBecAup/oSgbTnZMznKDTW3gtrsojdCs/ijlKrJOCgZpa8YXT0qUg7DvAK
JznV6soX/fVc3MFw8XuzUmtztnL2NQLZP9bkN7wGsyGk0KkfVOTK/QHOFv/0tSQww7vPVrobDeyj
NfCmI/7Pt0I03HyPRAbqnfDmWydmhbegBdkx7lCgn1vbBdgaPyCTjfN41JOpdZai+afKHObmhsW+
3swqSR70DZgGGqRBHtMu2AklcIN7pty6MA3jtntd0AeENJCqyT1BumzuCdtYnr4LByADK0jFACV1
x93jKDP6xXDeefxcLl73qKmFkIQpJpsHq8FWsbw9AB4RGXjl7cpt2JTX0VVUPvT6hZCeoJHLG9Dt
jK/ZvmmwDVPTW+NYe6veU9Gxhb9ieF0/a+FIS5Fb54TEnxNEUmikRLOh0RrtypBmjaH94Bwvo+k5
9/2Pe9yc2X3VHMwywEAPpUdbBJvk9MzCGxZWUsv7I0vHwa+hc6feTH2WFa2lyRr+JigimKSBTCJT
UIlhmUBaCiztDzKARGqeMSkcVpgWTIrlEpSGfCdx2Iw1n4aZGzzQ+/8hViYhExKN/d8g5wSMMiyF
DrzhN8ZY7C/YgY5/XqeY2FpOKoQkAHxwxLwkpGY3vWTIJR6BkyTQxsNqQt3hqb0BfiAwZx9pdyOr
44fquo1pdDdAFR8+Oio7dNZ1KYIcCf6JJHRZ4yQUCDrrSEm964aI3eYsBBdCzds4uO14LyB1D2Zv
gkIAEsPMGTIyXJdpnGlLAuS8TklImWZ7JSO1J12Kpde5pIE+YiUvEUUzsQH1lPvjH2z6sGQm3rd5
5jpEpIj1WJB6cnTtQAuYkPuzbJ9q9+0Ls4oMkz3q1wfXRy2ZPvoC+S7+W8XpqiUUa7EJxor7f1Oa
uOZ43BxzahFrkmnPcvEVM2CNpxlO85cREj1XGGck8uPpERyu4Oem7aghys2e9UF1eugO31QWBRLJ
cxwcn0AUmAklvHrxcv0+PkgCa181y2R60l4yWq6ewTN33yyLBW8bSPMxuall2aie5drOTt+PfzmX
+gDYSSltj+GUqTbGhyRtBRyQGVOYcU9t2Pa1HyLi3JK+dJ/mNzDIdgdi7PKkbQ/Vj6ekeivitPoH
Rx3GL5j0ATm4lpbwemf8eubbAy38X6+aD5SbmyYTKFa4b/imHuKj5k5+PDbl/7rHz/QzqRhr4q3G
19ZzrO35uFAItAQLqrIwScfPehJqTtMn/P7gcn2qkdIJrcQjC3UTuosjcWFSdJ52Aq+OeCPbft7G
0phX11iDSLHMGXi389S6rwT0S8gXNA5sJ3290lVv0gOyQnotvDnPulKA4cIlkiE1RiqqMkflrOZE
u7W0JzMS2eOeGsloHsHMTVZ9Z1eFmmkC2OqCIysa81t6DaZzUgzhN+rQElhRjB8U7ldN3Piiv/zh
ua2IbtPVRZMPSQoNaieJupHGQbfdfqMssq6ogCTb9rfYDeTCWIcWO87E8U1wFWc3+b6TcApBCiWl
GP90rYt0b6yFRQRSG848Z4hJUrMK8tdMtrvlOIlps14gRzVjWLVNl0//Qaz2AzYLlZQy4Huo33PJ
b9Cv+WWAzZT41bzqKmAW3INbeWf9ScRb0RHo6EejjvbB+r+w10kM1NSPtfE3JkMr88JUZCveSILH
4JZjNXzDYAX8O9LuTowTgi4KKQxvlB+2XbpPNYTZx5UlzKdSWo8YtSR3vZ/+1z6bTAn1oI1i/EbP
EpWA/F3dCo14FW8vwVPtOZfCy+xPvEPwYqR+NgccezbHcKRXOK4rVVxLNlhYo7OikaCdgEiqMG6R
/QlqPK+cQevMVSpBcqBWLZ7P8srPx+pTUd8Qt43/tyGyRjhoEIkrYP8+WRPvzkYABBjYq/oIGPZY
cNvJi3mWjGSgUyxBkkjUtuaFuwCXvOHuNV8zPU762iHUj7N17cytgXHpcQ7Gq2OFS09iEnDilTX9
JRLcyfAxWfPReOTdA/xK11Y05QwXGAjwKPmiegzK2kJfOrGi9Dve9aJD9wsET/lrzvfuklDErvq7
0aIArC57zxxcx0IE8kKs9EmaJNJFbtEKopr9VjQAk45wKaoKFgo2Wt1IVprWtShbh4dwIwcJsfM0
uRO8AKDOqgvUrGMPTyVLqLtY2QuJOVAzxFR2EBLi4uSgocdH5FoHNI/jJlieUqGAh2r6beVJwVIS
28fJkbnIDmK75TOZbUnVkMVNLqSdE07caEY0DVHat9NxgscLpO2TIncyfM3P9bRIbOl0DrVt7OdE
ksaF7vybb9rJ7KK9PDOgiTN+1uJ+gmFJhbmi+NaikkBfS0VcAj/VrQqR4esiHzkl8WImJtIuQ7px
00k1qlpJXeCcEFEjJRAdY7Fr7QL61VSS/owDw+45MmIzjD7IOIDgHlJVmYoyZMuGtnOIJZSfgEQc
HNqTwbC1zY4AZf1NlojQBZiBkqr1hopkUbOfbHG3cdcxZscoOAOlsg8rGR+D+UYI7bOzyakGxpPU
dGM9D/LZydXpJnrtoDFPU4Xsiush8nGcF+zN0TEkQ8c0zuIUxbgnD0DE3FjysTiXoqGMcNcaRpkr
Uw5wtBxw1NiLVrmqxqFRzbNPc8MXH/Ly5PvUkJU8IhYq19s2YxwL4+EkAVFooenwlHxaSHpWOKNl
KwTWaQjEAe+miR3xRyzzqQENCDPINDOBbizPbeRJ8D2OdMdY1UQ6JtrwlkvaBAoevYf7sKoN2y6s
ylc6x9So4WpOk8mFR6EHwQ6ni7PyIqNvfiC4JIoeT/i0oH8m7NLjhMSImn8ZpW8mxzPEGuIz9ZYw
Id2dTfA/iECMAoCVKkcqPzQEmYkJaddDNcjs1OYKq2YURCIn2TUTnvfx89bQJdmjhxHIXaNoFRWp
vq+V2k5ZIBXclIGSlKcDirSg6yeEYVYbzQcuial/7eNcGaU97Ue3yz05xwNzOB1Zk1YfR/6EYzvV
s5WFCz/Uvf2UOD2cRlFcfm/2vGwdsvXxY3iVmx1eWMJbDzgc4JM0GxHCeZUSrIqINnjJLOD7xn0C
ZhtfzlVWfGOb/1F6Y0wJZqEpPErrd5r85HW44n8pLnd4sNUbzeVds/mXZ3aMlGjXpF7nrkD2fJMR
F2R5JGyr2f1fOAcyXkjA3loOXr4iM+1AMvI7d3+L9WuhcRo2YyJV7HPcQAAj9lJ8VoRGUZcmBZuL
0PLeD97zsYMIcmj1iSZwinbZoxbIq/FM5NUtgrbIMLQtyiVaYah7CSTVStYjhFvKwAw4dpQK/eVM
Cuj0UrB/kqathGgLUeyyp1EjMYwlxLvrTilwJYSwg7lKD6Mp33OHaO24il/n1mFcCqSokOJCfihn
Ij4v5NSbpBKneEO7Or2ujqRgAbq4XKIoOpLiMAdXud6uhp9pRmdueKZLeLNCLzOqAy2wwHgTFSaU
HiPdK3gB+utfKAaCk2Zq7aKNkSAaVMMHV2fE3UTC/PVeVNf6s/TnDF05gNCq2EeXVrXcpRIc2HLW
V4/bZxyVKoDPoGP+cpTmU6Mc3ablktKNQFt08k/5JZxVttmCldlhFeHHk6OvMJhQ4hsHXzCsm3qk
9tWXzTDEJokZjEzHGuTag9ewkqxjmjbA77AClI5a9E1L0e5jgPKggQDY5em70hd4G4A6rexB4MSG
mzRGuCDqdyn5TXfokEqDBuie3C3EdgA9y80V3fhsbGpgo+zmyhLR6tjEvRnCT8i3Mh1DTsOZFngc
exXGpqxY2XXLoY0MbTIawJ7XLPmi6z5jvljSxC+nEnPas1lLOI5AkXB13RIVgvEJMFiKgZLU5Ork
VWtY1btLmcwc1CkYDMKniG1kaXAxVUqwP0tgXRQPst466GptSQ1MlkzWo0jG3hiXDl0Xu1kOyyg5
eQvLvE+BwNS5Q1xIYGzD/0EMCLL3c6SekFtJDRpiTBxIG24PEDfMlcXQK+EjchXp3wJwkE5BNKBW
ehE0WT4DpiEGmxifMo2eTHfIZYSZH0BJw0PIEbXBkRZNhqVDZgpzPIIFXyypcUXFYmhUpGR6YHAT
swZA+G6TTh9W/wFeYp7s6P2dALTF+FpEIXHlHLjSLznLZXzmYa3kO2x1ua7yRhN/OeHWD/8a7os7
VC7jm9Vfk/StYwMav9IRC+nLOqdaxlPx+GaQr6aWA969SokVMkHawdmK43t+CtOG2CqKejCw3e5e
BYhlLxBEvmhOy7PfKwkPGXOKdh6Zze42L6M62GqcHlr6sE9hT9xkT8DkwAJRvp6zReVF9pWccxqI
ur/U2EvyOWnZTeQveEnjx7sIw2VFIvb+B7KUdhuuVAhpwc9FtTY9vXKKl5kQuIsy1BgOfV3EFeXr
KNrnaHyBbn8gaOLYKopb/Dc3GbyD+LYVtY83SIYPkW66i2x0KUOOVOyMRvv3/C1HnZDRwiGMJHok
T2nOoKS1mEDUqSOB1qRPGNCXspZiOfgTAj1dpxOhL2qdmcbAPd5A43sejslp7phRtzxz6l71+WsC
9aNUQlB3elfm0IeTH1cz5bweQj9ASU8eF4KOPtFjvd9HReaM6SjDe/Dj9zsBg6XcRljoupN+wqRL
cGiNxlKV5Zf3FPSyk7FLwQp4gn/vHRTjDvluL1YKg+xRT8JrDXIWMW9ZEWNFf4Hwj6EWu4dCoG3D
jTDvDJoNEaJivRNJ70bk+rYavSQfMBezihtxwLomoCzNwdRuwZHMYAorStzqlxg8DyBSbOYK4QS7
V+T8he+ABW9x4lMIIjPnKLOs76SihANU5TOCiA65I7QUCJEBO4bHJsCZXuyQ6+70Gs/JsPNp988u
J9p0TieCgAS3kJDQnf5QqvkgDL+u2oHeffxVlx6A+eaHK7aST/9dmHmvMbFYTelvSLMzFYICzg1O
PiLHDZRFlFvNvqApTZqDj+htQ4XuNlFOeD8pV+KPagldzausjFmYDzrbs9lG6kLBuW3bde0HFN3b
fZRWfY2xNvXT1e7QIsJABsgWIW3yOzxwbj/B2uezEgISHSp5Jfz4FI/0P+H90k9kIl1Q16HrxaZ+
zUmLK0gzArYd/7WzKBVQsc8uo3K7kYh2AmOKekxlLo1guPqHqWoVoZ9NzZm3ltGOaSTEBkljC1O8
GKJIFWLC2HAFP8gGkqYdcN9EwxN2Bwxuj+qpKQ0TG3uvKKaLajIIh8amQ3b59Zm/KA7NQPddDeZP
ClT9aueO0lhGfEr3PwNEKYJWBazEYcNlhsvpVSTXmbRtXDEmYtLBPbj0o1qJu2of3ebigennY42B
9XCJeNRdrgmtT3jBPKHKKR4N8vOAlGGT2pQCJMRrxzvtMkkzgZ/3egudCzh2xaet8gIe6fMgOo4o
WCqdpPXt06XxVYCfCzVVw/o8voChiVieDaYw3vIbJA39eNDB84qvjGe/ymdPx+exYSOfgjBzOnIY
lNLz2FMCNMvE/yt1LLLyfEsmGNo6S1clRFBWY9PVuBMwT9ODQGpOzrIcmMLKYMeJ/RF1z3q9wsWq
b5WLcPASYN1d35r4tpPWZOhwp6+0n9R68Sj3fBvhJfLoEhhnagawtczeOyPWSEMXf1aRtJAtDxGm
TFac1em36XCbLHw6kIlKthwTdNoDj2NrwgodaJUFXintfOcYuAmBpWTI4xV+/oHGm71W8nhr2ZB0
w2FmVlnwt5C/wY9jNx9PGFmkuY+lLaIlNmxZbMM9ZNYYTNTc9kgsrdpo4BgMmuh7YpIjkn+UzwoN
RdGnEfQaZlBwvyH2PYVSpR5CQ42SQp6OTYlhggkSW5yUGMCzbxujC2YwazUHqWsigBfWsPGLMM+V
5CwKiMpwFjRp5MjzUNu0VHcQ0Ps7ADJIC1WDcURXpZbGvp3y72LATC0wtn7EAAu++hLSR+s0M4N7
XUTnt20gKsNjXjYqtN7EI3mEqBoGfORYgXbOEnY055gVCcPTjrPdpeh4B1U0G6ab76p9cz721YsZ
vriW3qcsiiuLPrEw7Hb9wjRUKUJtIMtXE/Q0YRVhazkg0pLTHDn8l9k1CmYPpCKXNHCN71iv+R/n
jNJvmU/86G3tnGoJO4OQY5O/SVDtzqP3q+VCnCc4pN/piubKEJscYesC8Y7KzeKEGdXLYrPOc74F
+KZyn9XtBAK9j/gip0NJmigTT+HXUlXrqF5dz2NaNEjbkht7DtCBsASISuicKxV5h8/QbHFwCADp
aMzbSC4HmKF8hC/BcJMAk6oqCmhmjpjfiIdtXDAB6kDQXlfAndvX3dWnzhDd9hlonaNd1ukbuTl9
sOqwKQEIaNIdFI3D5nstjD/zzoUBEAlmbVIWMiYsL1hmeVjyHMFtWbIAhGKdhUcW1ySHIamnBi/l
/qXhKs8Dy1ddfuMVJI5MmK+b2mMYWA+7AJbnYY+VMZL1pBOFB1S6cFaIUaLj+9skkKUHnJOuhMjy
hD8edMj0D7J8kwPFdS0mXp5dik+oadW+l/0BcHsPrchJqGR8MpF36ZGM/U4u/97sY6LvfkpZtfRx
4S3UrVjCNYIMiypru2uPn1SiolwqFunt6Xk5ntXDrCb0j4W1MufLKawtZWafNEwIJUxPzdx3rJb+
/rFfnUHowqieBeHfuEmvyTRQKcoVMkpFap7wnwtcBWXTu54mCW5TS1EKVGNS08C+mkmlHi82f80h
CTwwgLu6KsMudhUA5h5ZYYhLkJOD1M6ZgkZSr9FskiYmAze8XK9CPxs2Wy8a7Ehinu7yUIZw9zR7
Z6He/qumeKMNUga3S5ofXIzNawRZpkXXvRcIJEJfS3SaHgGKie7NjUB9YOKakLIEvEsZukg7I74T
o6W0PlOyVXsLpKtKcp9H237MJaVoi3kbAf5gmEXzkRxJ1/1guIM/EIK2SNrx4aXWyRIi4vuGG1bB
p+41Wnmaj6ukvcx/Grzkbu82j6DbIGRu9y/amLFjZ7A+JOKvGUIw36CX6K8mC4g3/PLElaASO4ug
Ej4wNKqCZZ8zSinrT9v8xzGZ54F7NQRGnOmj6/NlSSVZRer8aoe35/eaah845XsH2JOX7AuFEN+e
G4J/r2w+chtCSaaxM2P3qdcNbuc0n4de9Ep/kHhSvVqRrfHY+gdBAT9d0M1Z6xgPTrDjQ9tpNR/t
r9r+ctPKczH89U215MG7AS/uzDcpSqy/Hj0FKojCHlLcO/aQGFaha1EpaoYJWK48ss6oxsOrJ82T
QViknwcIdt1LI+B34pIX+yLckX0pPrNq5EBjo/S/mGA4JA0X5xlQF/AseDeh6+9tCzJMp7eND7zU
5J1IHF8l7udni7hLjFW6DI7ELZeQB4DqzySAba5Bth4GbQL7AbhRkixfXp/N9Bt12t8w9MO/4jdI
PbDmUKftgdUcusP1OI6w++ogj/vOHuGsJM2zsEImwIjJNn1MZe5g5jEzsn3a6cp6EjJLNMCazlNq
gT0X0Ng05VSDRjljW2m60u22rmyXTGmWcaUGtlKKJ2Gq6xcREsmw/p0sOF8HVmcO7uv+R4xQFR+k
zps/lJ5fTpMxJq8GW+oyeNbHSEnSoUy4p/14eyxkGd5+Z0bNRJSawfTe2a3ATe5zkxRvVrCDNhzb
3j6HPWHFPlYeF9XlE377HmBGaY0oH00xnLVGkonDXvvuOD2blz+sKVgn9xfx5Zf17GLY6NR5vPBN
LUzineTrmyoPTIzYa3ZBNfW37ZdJO1SvhY/ksUnFWsJvJXbUSVEQW3i2bKVdoD3q/OMsqWeAFOwU
91nlF/nTbeJUYtbbOZqrfDrAkzx1ORJN+3tBBUO+TpbfKqlC6VAR1wxwIweN1mpsq4t0eKK/SBtT
liAtHYWkyhLOH1i7IgmOWbeA7TVTZZXuogzwjGICVEY78zJnudD5lEUNa8Y9FxPyNT5YFErZe1gX
ZUUesjNe9Z4Xd0GJlxWf2rypD10o29a6I46Ruz3fz5zfRy/fMmACkq17asTj5f1GY0Rr0E8uykm2
xO51mEV2xBuMT8BNmMjxU/+7q/LoOOz+VSRx6pr25SPPZcKFdOLr7HIlhYu3MY2K9DReFwVeeIMA
GIMjIT0YbPLy9lNXck+dtp8VRhnoZqqarqgr7tU1NjMcsopTGCCZUQYsbFZ+BwhRjZ9LJjbHcHrL
BCYzXYcasrz1qtL2sRTHtWI0w6ce6NWK8ph2bFv/xRZgpPwMS7yVvLKIPnDhiqM/OsWq1eyiRV7n
9DRzNx9T/p5YkmfHgh/66pi21V4uIgqk/dAswW/fEZhbdbtFXF2skhZjFECzdyvz0kNENoXe9fll
DeFZrhctPsHv9CvU5F77j+QQ5yKc1uRC7JGdl4fUQ6t8yWCr6te5znBXnsJs0Fuu5z71yTxIufNH
CTRoZlyZn4/ZEKY69MrpcJIPrevERJ9ROBPbM7Z5Tv7liZvkGjLbskHyPQhXTSBgiv6EPGoqTTCY
qItqtnEBCB4yWZ+e9Ouzot+6pyGcTFciAwutmRkeUBGySGQ3fE+v3kWJzhUAjJxKmCh4tqu+i4P/
zTfn/e1SkmQJUUmyk9wHXXtxQDffv1M+hDBjvKqSfyb5s2tk2xg1hkMY7f/PFCRYA7mQPesXNyUK
lYni6sg6ret86h5aoCNlo1WH33c+CZHqLFiy2f2Gdzw5CLpQB1rQ0V4DdebPd+65xB7DyhnTlNRq
+FZmrsWq5kOhHzoTwlg7tdbibhyAB83vVQtH62P+7idJWsYSrzrSpPy0nXokVyjhqLx0lbuJz+aD
S1Ivc0EZhD8XZ/JROgeqove+fDcnImHt0t5xZA1+YYakF0stCYv6YvcEroD6tub4KYk0bKhWGroH
1J9+ZfbpVF5HNbY7VWoYbqawA5yaIHmllNStYuubEQXQiyMmlJpi42fYHSlx7WPVwjEiUqAN9WCx
W/O6tuGKUlC9H+EpWhxkRwRfHDo8+b4Ofj0QWMyKh8uOgp5EyznsXS9B2msJ7w1IHCQOrKba3cUa
c5Or2w95D3JpaxYdy0KSImn89/GoLVjF69OQmys6rkuPFxl2COxvqip3gwR/EIz5uxxPQUaxG2Ij
bOc+LideOvWtR6R6MabSy3wmpAVrH2mo/eRK+msdLZlHFXeAqBD4giKFApEz9WY03v4Xcm9Bd65z
HYcQTUrrXDn3XrvNwIi/WO2fW2kMXC/65n3EZRq2seaqKvMZ1dr7AgR1hXYT1KsUr6U8Er2nTjtV
ibPdRhVL6zDICnu7lCIsxOjzAiFSpIALR/78tVxugPIT79Wv+nQieySrWAq5EvYLnET4x5tGEMk5
kudk7GMTQReUMTZvKnvGAH8LXRXCqWBIqIQ75HktzrPb+ChhTLrrxVtK2vM6/EMyehjH+e/kpQ4k
32lE7SjNxTkPHtJnNJ7DqahZLfefY0jbXC9Ua+979SLdszRib72nUaTeR65W9f7BnGIdu13tQksH
kF4bsZ6ArViKiHpw4RGNYOUTlH2F8fTJcMtXLLHWtd08JZR94e7QTzv1pkqoUKBlWzkxhq6RGc+h
ZeiZfUgUuhN3Xpk9lxc8K5KKF72CftfaVAWnqeHCL+VzFwHnjZieLAVvaxqfZHXpkf0FPp+iGdQb
JkMMeFlHRtHbVAvVdyr22v9UVXDZsGLlM4roQt2AQIfgfHfT1R8zXUb6VdAaq+SXajG8UU3A3we/
v4sn6pwevJYYRLe2IBSiKb56Vqz1bCxJyx1IoqR33WslqWrNMwVb6fM8MrgmzQTU2xnZlvqicljm
A9Lox2TAxmH1kIbQqNvt8qMrV8j20EFJNktwNLia3AwTvZWKEdwLpj+1Tk3u4muG8BWKLL0lxYiS
wbxZsusXd4ujyKUkMmiPTgO7y8lsEXgevHMwotPckYL1JY51JWguzMskDsfY1vcLgh6d6vErX9IK
TQJ56yKaz+RykgFFAsxeIvc44x9epmZxE14bFM2jVYziYi0PifRJ19cSimzhMiUwF1kmMR61t6xp
epEPgepRFC8HJUURbBny7AuYZndxdYA6giO/QkVLtj5+ML9xC76cswRJBpi/MWcEvPx6S00xfNtb
fxyg6n+UABpxRT3oOq0fKc6oEP/NymUcD/wIwZK1VBJWk7eS88Abi0H+k3MoP2ycJUeD+OREyOf1
hPdldtsI7yPyxn/rC49QWsMVT98rBSab48o4ASguCzovUdtiBXotVFAsti3UGhgr9WNW/WF0MHkW
KL2+hr4u8gzAmDSYp5r+8ZeMhxFfhM0VdURe6kFuN8H3kACtc7XwCe4Kx9aC+LO3af0HbdPh86Fx
6pxNxlzcH3pAP7t+0Rc4c9aqQ7zF8LmRnOAFvB3UVQz6N7w9Jgw2sNuIGclYtta9cWKHuVYlGRWK
jwktddnL+7G6wQFgo1JugSTf6O3goQx5hJcj0y/uhE3H3FeI3xzMwgDx0pptz6w/9r9kP2Ex26gw
kyeHlluXgNCaLvALw4LbN9hQVLMCorpd1L5Sgzhi/f4OI/GwPP2h/ajLQL+aJ7CQWO1Vn6CThghm
ArBaFXPkAaNtyFl8OP6jzy1q8hMk1LUCDqWjsby3K3CyCJFY4vv+wqSStS4OpPF6b2XebqGcbtYe
Na/IYIpy0v9UWMhMSI2G8hWrfMN8Xi3clXP6bZVaP5eArPXedEMqE3oiHbB+/1Pb6qfnPWA9Vr8k
pkB1NlW2CroDs0EjJ4k07x2+vMwBzzqeiRMMGWB4QvXJ+A5/L6MPZqei4PkK6/UjakCJ3O1jNYbF
vP8E9w7K39LF5nthq25oyNQS5JbBEfQeYmHFBef90fCW27is6m30TcQUjg2sM9PM9jJtr2ZUx+Lp
l765hj9EsihSCns0McKDnuZIufKCWbdIH02G6rtvofZBAEANmzCaQJMxQ3JGMGaeDNkqKyDP0lZE
cVY2YZruoxd631N87DJMB+w1SN7XN+i7s3Q4TW6avmah7WXZM6+yl74K2cvRzhv7pQ2Io01ZX9gr
ydwa3nOsFiNOWr14/Z/e1MUs0P4BLMtji/fQw7r18Y++0YMFNAyh+zhR/c0uBVualMYxGQ2zd+gl
M+YaV2D2jGY53uNiZMgLMKmVR2YK/1gwsVkYpGvaOhIHiibf7jKfDbeXgJfljbVxtgrQ4mces2+n
NZZVkjhpQPxjviEWA/w3OlfTm2X424WEGPnjFRIhJfEmvY3Nv8uziMULArX3AXxRbkrx8nAV57P2
uAh7SawXb1k22hnJB2VJ/pCc+ifHl81nmcc0EKyrHeo9sSCirVpHSNbsn0XSjwjDA35kNcfw5UPZ
z/HhCcIsxYlWTJe+rXCwvgkXL+NZVwFy2AxrggzbYjlrmK7jfEK26QdfW1HrhRoGiufUPaKdVNpH
Bfy3KQpCGn4lQjoWzhOKy8jFfQy5ZTiFumHsDX8CD4UkFVA2LxwrRprxKU1kPl6DPDNKyZFwTOa8
hdbdaRYXyksAQbOVnp6uO2fYdJJoHFfe3Ol/hxi/KHVi7V0CpTO3XlSkRXi1jTFBah8SI7xfTLZh
UIIcsjTwiBB40KFJlQ9D7WYwQt/ewPkoU7guFKDVv0KpeupyjqIcba7QGK0wROyyTDAOf7LxBSKt
sLh113TJ0BwRbSy4N88oDUMWMd+bJ/j3RJ9VJ0TOw8niRvHHIPDXY+nezQ3bmnJlHnXpZsMv0/Nk
pMQ69G16oUE19EALdcd23yzTWOcSiBg/Ul+Zi6tjgoOzZr4PwF3wybogJGGXF9U3O97QL83EP9wd
xxUtTibIFVi44lB5Z6M9W6gHHWqua2lBD2Toc1AmA6zkYOotKkaBGiEUv1bHqlyGhQHV/YFm65iT
jOzSkl4PKx+GO7J158e4WjFHnWJuLTQpORMlvfo66z/an6645bdydFtL2RjimkWvvEQI6pg2eTFc
9ez3SpovF9DJeWzHtPDpRoQ8Q2QWo2VauFVZV46PFb7oSDK2XJi8GV0rXVGFH6dpi7yiiTeLAYOp
q/MAoXO6k43+Hlb5/wqPLrbc3xp6XFkyPidRbb+UO22HV9lRqMKnTWsEwwXSL6ydS66fJwpda8d0
XtHnRWmahtWV8w0VnBLrZKmrLfMFwzWdft3kJNR/nQmR6myJLVNpXwstlvrQwxuntboSQacmwdBG
icMIklTQVrVoG58GmPkkVsxWy+JqKurNzEqDrdHyWHmDOMhPqv3j1hSk5zXqbnZf0J92O8BcPsN0
+IH1xqdER4n5UinsWS2rnX7Nk++v/9yJRN4LqmSoVTrk+xR2Yte5ycfubd0Ce3rfUsLe22TlD1hQ
9iBJa3VY33wLXOBkkCTaVkH12nmCdhaWgTHdWlQtDrWqeFV6SPfJLsO+IFdQhc3Z9yvMstF/f1ye
hlaan75cy/fapN3o1KlDaRbr7dTyqYJ3to8qO5Il8lbstxtijLzxKFsKZ07UeJlrQ3ohxnQoQksA
1uIFS9AUb+YsE4b/K2Ucnol7ts0VwysbRkUvpt33d1cwJ7ynV1/KVN86uh4uZTmiqyiGl/R6Gf21
n5qYpqFncZ380L15qB/crV/UyZxqgN6tD0J5Wl8WE1iPuCHUVAjfEhCjb14aMbQViNf1YLaaxCW2
UxbL5J+sCzaoZHz3RBkBK7oa+nEgd7VPdCGIeIHqnjHgj5lifQxUWHyDMRVYwx6LrDr+xKezG4S1
Z0uSlgPTasnZQ05aMuN5aQFwsjw6FFLJi0KXDKMvzIIaWvsLHx+sDmuFeVHt6W27eRGLtEe9Yckv
EvRXYtN+2WNW2RcwtatCjuWNAf/IhczqD4HgdTJ1QnPZseQgn5u95OTjUKG6r3pgJQBve+J06tbt
KAMwQnHgkWcEIdqdar6K1gt9h65f3LYXPSFKweYhwiaixuisLz6/KIaIhRTO3fBKcHuAHTCQJnoq
858UR2mu10kGUfWdbccN+8bcxGBsNDd61R3syxdQCanqGEAQhwU7mDVVjlWp29Yjv8AcbBadHD4A
tRSvmnMf8BhOGYpnZRCicZQDlC1+6cd9BtAUT+S66qn1TcX91UU0wBlDnJHflIhSnW1VrsG9sVXT
cI6LLfk1s6UCUHdHhorVBGASk4b8zgDbflimo91y8BXrvTU8zMMTQGLbmA3naBT1MbvFytAPVsLo
PTwhRJJEpdWI9nXHGGlHz8PrxoIrYBvctio0h+RyIDxAgJoPcNr42l2/s0G+GDJ0ni5/GfhQaV03
E2nMMbF6x8KfGH7OHWBMu+QMwCzy6zN2dmFZyfs+2wFAPFw5/Qlg2QI/GCe8t4dyKkBWUqJDxBXh
YUd7Y+XwYrrZfo+m5g6GYHweb5csam7I1km5jDUvqTp74NGzjs4P0dqlgzGHUhAqVxLSd4V7aTG1
/QWK8KzY/WysLIKYqSwep0LcYDfusWh2SX09LV7J+X5WGZEydj6tWXcBelpDxmio+4VNLVIOlJk3
CFIzvArY4SY4yGdJtyNcWSYOLSaUjbE0a6yuJjHNJ4JOjKnlGaf714+s0olMd6Io/u0ZX6wiMA2r
qAVmse226OpdML+eDkKZsv4UHJ6PL5H5ZEaZ7JH15SrsHkUieh1crdqykYuK7Mq3MtkthWUaRmcr
zrgvLMxxNKU7z4d6+siHRpwWkReLJNSXamR6eYijlrdQYFEiaPGBP0x9jUk5KWBZR7dbiqIXvhRn
0YJ1WIuqmRePqkNsc2Ftb902WqP/ML+k9nNmKYI9YXC4uCRt6s8Xo+Cp0rveP3ARjVrI7CqPJK5S
2OxJgEG8SPvbubXtA48CVnlgBqW5SJncR0HzOSMDD+u+5sHC4CdXSFqIGvklty7DvizMGlgq4ULV
7oBXpSkj4Ut7BqV//V6WZU57Ugpik2ME0zyIqx/C88B+
`protect end_protected
