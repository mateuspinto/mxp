XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[�R��"�Kr/�Y�*�����#��� ��#��֣M��&XI*���b�$G_��S��l^�Igs\�n��rT�a9@Q��3k���6��h�/ǿ 7�~�ۗ�u���h�y�����:�
B��|	�P�*����x��V��İ��P�����u�4�@s+H!:��"�P��u��l�H��!	jɞ���T︖�d}�����l�1�˻�?n�C���(f t��9��L�ݒ�u d�gg��2�}ֹ�%:F���{d�HEi�ΓPȌ2�cu��!��˔6�'	[y5ӝ�	�п�m��BL{��
{,D6��z���	�g�vm��t�b��j��p>�Uu&���(�$��q���Z��[��ֶ�{ހ|%i*�u��,�~�ʖ�u���5�>�����}O�;�'������>g�^8�U/�z��{20q����w�_ػ7�+5��0����ݵx��<=(&{U��"�vካS�
�%�Y�%V�YG�Jz"�5��Oa$�KJ����J7�	(�j;�^�͔ɺ��L�����STx��P	�m��N&�L��<?%�I�x�|�0����HW���T\��|6m��ad���J�:�����t���%�/$V5G�L�[	�(�(� ��ѕ�_�ƌ�Ix�,�G�;:�cؑ[�YB��<�V|8<v��Z�s빹�y�� �c�9Cڅ	�j��:���w20�[���v�R)R;�>�x�p��{b��(����z{o�g4]�XlxVHYEB     400     1f0�)��Po�����g�>�R:m^�Y-� �"�p]YY��n����xRfv�Id�P�D�0��ő����O�3����8�8G�q�P�sC0��Q=Ǵ��Zym@r��Y�h����^����Sɹj���}�\/�1��vۃ؝ڨC��Tq��OdB븥��$��db���U��jzf���9���
c�Cľ�|8%HjZ͵fI�T"��z��n/�XUx��� �\:g抲zf���jC�9.��Q��8Ԋ����<�]�&���(0<����h�*�kh� d$�j�uG9���R�gK�kc��[I)�܄� c��E��φ��|`�[u�T%æ���F��Q�Ĭ�83�8��/�d��>6M���v���X����Jؠ��c����5��Αs��!`gɎ���W/�핡 �1H�������a���ǀ=��v���V���r������s��VT�p+��;�4G�XlxVHYEB     400     1f0�w5��S��f��F�{���&`��H���(ԕDoD�s����u��/B��B�e�eLH��Qs;L��sg��������|���M#��@�暏<���`R�T�W�=�������W��V�4(0��vr&]�B*�BQ3QK��/�_�O�~]�6dM���H�:�$��t�Պ ��9��QJ��z�(�t�7뱒���lǲ���21V��;��P��M�u��U)nC���x!�����k 1w�]�t�����{�����!���7���X$Q A�2*��-\�r�h���}2H�:�g_�4b���m�~���;��mC����~)�@-��u�B�.���+5!g�O5g�<%pE-tf��_�&�2��{��5ʽ<p>�����f�*�iZ&�^}	S:-'���Q����ڙ�n)�|(�Ӧ�y�f?r0��Ff[⽈��ș�9�>�\Z�l�x�>G��z{�'�$��L���26xLrg���MWcXlxVHYEB     400     1c0}�!\���sL}<~Y澻������(�,����O�����pOئ.����&��ɿ�4���UA����[��rG�S�hk��=�@��vC{�u�g���~W&6�	(��m��8V�4*��A�ԁ��-D�Fx�k�[�m1)K�8�vs?_�aj$��!��O�.|탌�V�X�rF ^�y��ٔ�G��:��F�۷x�T�F�.
NRG�-�M�����'�G�n5U?�4�e�`0�˰@���/׊���mi٧�X�|�q�8��������6CQ����Ũ��˚�^�s�8֠j}�d� ��1�Xܚ�OB�
)�=��h�g�+�Q.N��I���7�R{��:�Š���s�~:�2�y_Ƹ�P�	>A�W�\:M�o5Cݹ4`�M`���<��ѴH�
�s?9)]�R&�еP3�Ry�QZI�i��Q�(�q�l�<[���nXlxVHYEB     400     1f0Zs7n��(b�{�L����u���W�3&ɢ�ㇹ�ʱ�@ؔ���r���+Q��%���q�5j��C~��h��1�A.}����TN�����^M��,��2�0{~�\�tcǳ�Ir�L�7�ϑ��������?��um�������'����;)I�c��=���O�h�|���̀��5���I�?����?��8��T@����}.פT(�%,y�%��6�\Y�d�� �>}ǐ3b1V�Aa��K-+o��J�ɳ�'����������"����Q��8S�;�Z��%5���xb'�V��[W�m��:�;=�7	�J qaѝ���Ze�n��B�rc��f��8U�:�zb�aJ�Wg1=(�|��i�ɐP�����aa ��,���l���*XҪ���xW����`�$��H�
��>|~���Hʘ�<Ï"Y ��4*�^�K���J�((3��	�7�o���<��d��32B����X��LM��nXlxVHYEB     400     200�I��9)߼�=�[�.����Uǿ0��^������F}̗�A�Dnc�l��;l@��+�9JG:1F�F��
�`.ps�g����hՄ�ⱷ��]s���!��JQTO��rH~g�PA ��_PL`8�������.<pπDq TU�+I��!�?ʹ~-��P �a�Ӛ.ҭU=��`���{r]P%fm��/�P���**������B-�%�aA��xD���%]�"1ex�
r��ƞ�-S��1��a/��@[��eX"���k��d.�=IiM��}�A)*�I�+���k��8�a���l�����պ�{��ԿA�E�6��A]c�_�[<A�I������)jߢ�:NA��_��͉�"��?��"cOiP���2+�ܵ��``�{,(m_�0���
3�v�O?�Ԕ[�8��'E�zM�
ʦW�9�{M�)կ�#��gۡ���R/�t�ʐT�'ymS�؆X~� �qg�-F1L��%rG����BV	����XlxVHYEB     400     160B��[k**O\ >�uƏ����0��u#
ǯ�^�ò,H敖CT~���&�H��0�c�wY�r�͙}t�q�ĕi����m�?�KE�Hxu}�ikSJe��t��X�s(�\;�uD��(�-�l>�5��ؘ���Oo���[�:c(� t� l͔��S(;r�V���pnlVCF9|�_0�ʩ�Z�j�����7��?�W�OQ����J9L�W�V=ɡ`�G�ciOJ>_�ؿ�30-�ԟ(���/�cs�O�kC�S:@����%�4CGt��-�h���S����0<�\�X#C�� ���`���Y/~�m�D���,FG�+]�}��������٬��FXlxVHYEB     400     160�����=^�Ӝt/�~�LL�]�>tܸE�ܛP~�\*F7v�}�3t'�ũg�"z����0Ӿk��j�
��cZ2��)	���-�4Rb�����F�҈}��()m���
{���;}����9J1�ut��%Q��S}|ڔ��:����e΅��~�q(�p)*�HI� � �t#��P����w���'w�(C(��{�V �M}�u3�%廰"���=�G��(��ʱ�Y�R�_z��Z.T%Nm��E{�ͮU�([�;������aK��&� n�Ny<f�����5�����z��z8��s�3oW��|�]�5�E��H+H70nXzw��5����~�F�a�'!suXlxVHYEB     400     1c0u%�A��U��.���Hk�G�x��U��ݓ<7��������59�qh
��z�R�=t�oR�!&oU�?��oi�����&�J>�����#&��;:�~�+X��+ z�[e;��^�n��E����o	5����z��;��;��B�����x��`"[���Ϣ��A�%�j��-�z�4̒��C�}�a��;T�DCXm�w�
�8��@b��GP|͵ř|K2of��9��́������V0�~��ok��&���L%�G�� ���j��n���WG�N7�Q�!9�,�KQ����$6��T��H5$��`��b��"s�Y4�&�~#��Ǝ��`��V��'�~5�;�cE~g�J �T|}͚����8+
��o��Z���V���2�_�6���WM9�s�gKӹ�T��9:�goH�����#�	5�"|QΖXlxVHYEB     400     1a0@(�J4��4P����Օv߇�~�)vyv���3a(�߃�Pspq���@E�E$~)#kc♊��&�0��v�������"LV̴q�
^ˤ�T���f��f·`�%UyM�[Y�k��s��ص��$������z�j��*�飮�w*�������������D�o�˽�v�sz�����e߲�za=6�:q
z�r���g�^����>Q4ѥ�|���-�\�y�V��o��*X��F��M���S16�r^S��v\w[�p��VzX#��$�t2[�ڞ��Rbn����l��Q��Ws����K�!0$�� �AQ=�zC �$���C�{�>z���V�V�sf2=r/��&����H�@`J�-��ր��ň�s�8vW��Ij��C�ɎX��Bm2n<
q��#��rL���k�L�w�ZXlxVHYEB     400     180;#vP�\9�aq�ȟ��y5��9��]�3�Uh��	��#5�H��t@ܱ��e�y��7������Bxϑad΀���z�RfE� XJ8ɓ���FI��垗t|�eB6QL�.��Y����=}�5}ԪZEflW�&~x�q�P6�J�Q��ct��(�/n �r�<{��=��S'8���Kr䮾������>M�B���>1-w�V삙m1�l��M�o3�Fe���e��u�n{B�g�>�j�WJ�O0"�޻ܠ��(0�?�p]4�M��6_@-꿺���,</^�����CQ�"����}c-4�P���d�R,@5�c�$��-,�يg���Z,���5����\�L9R2��b%T|�˷}�55���A%���XlxVHYEB     400     160|'w�M���Þ����Y���2�h�E^Qf���>ļ٧$՟��B�)K����K���f��f��`G���(J`۶&�����"�D����&�0Ӱ�������W��A���55A5���C\��D�$�T�F�uTw$�	q/Ob� �YQy�qg��x��a�G
��P�|��� 0U�롟���G��-B@ˤo�&r��=W�sME�1�Į��t�N�,[�V&�5��:�y����d���a���]Y�y~;ܢ<�K�1��(1�rF����!F|Nxai:��X��s) �>�y"�����1��hbбfI�Ȟw�^�ɳ�0�`h�>�`XlxVHYEB     400     160��m���=���ot$��Y2���/h,�'�ds�6θ�����fn��xB�Ҷ�7��\�����	�^/�W�����?{�<'̻��k�}��ͭTzD&�z;]����%��v��Jy�D�ȋt�C=��<�Kd�������FN��U=,����)�$����u�$������"�f�)�87?ʌP� s�^���i ���bi�Ɓ����<Gk����f#�Xk�v�q؍��yA���ժ����u ��ߞ��	�µé;U>-nߵ�ʲ;�؝��mZ��9��+@Y�#�%��k�T�&�
���+K�-9��t��{j簆�U���Ԧ�O���j����_<�X�_XlxVHYEB     400     1a0:�f�	M����F:�`�-��۩*�Ǆ��PS)�U��y�'gp�%��4�&�$��EL�+��
�A3��gެ�F5��p����ZObK�k��*Ў��S�KL������tl<R8}9W�f���xq��C��)2��#�����_ASyyK�A��U�V)��l^
���X������Y^��������vD�d�=;��3)4��nkT��E��2N�l�q�*���],�T�����6�)��'�P#�s1���nvl���m�T����u\C��+����.��w>O�G?g�;'�aw%ħ}�+VZ���z�;bg�R|���IlT��ܱŞ�.��(�R��[*iE`����.���b'�/)�=�"�#l^� �_��ѳ�o�g�~;�����C���XlxVHYEB     400     1b0���N���`B�*��ԻѾ�U��:�ƙ�j�u���������Q����>}�x�Ԟ��^��o��6٘b@]�#���<��������O��������w뎋���|��.��_��`�B�6T��U�����d^�"�r�\�S��U�3�ǂ�q����&a���#(���ɰ��^d����~:À<����[���v�����J++a۠�w0� �+!��:"�}],#%�H3�a��U����.��O;���/F�̹
��֎��7���H�{�@u�HO��v��;����dc$��0�S��fO�BH�\��y䓇���[y�g�F>�HS�]�~�_KFS�A3*ϒ'�����?����'��Q�[���M�2�w��UpcQ��X&��s�m���Q>B��}=k�)�wҟ�b�PXlxVHYEB     400     1603[��1�k����w��I�!����֫gމ�r�YI_b�����j���{�w~<��/&}wi[�1�����fx��� ����S�Q>� V[s��(� �>f�8a�ܶ����~[K��"�6���V�2'���!x�I8ړ��8�ػ�]�<j{��[����zB�Rg{c�k���a�b�$'�	,�ъJ���UMrw@+|���q�8��_e^_�q��rc�>�f跷���%ƜK��Kc�d��|^�����L���tJؚ�w�b��s��U�8��F�K�W��a�j1�e&
<f��� k�(�R _Y�d��v�����}��Ma}̑ӁXlxVHYEB     400     2104H�&����4��۳�CG}r@�v�hiɡ���.^^4|N�{���i[���BLce#BV�=�{7��t�IJl��Θ�P��+��Ї���6��"T (Pl<�3�f3D�}�ʑ�7�i�\�t�ոj�eL��$��4Zm��N��w�&��{��J�$&ď?ΜQ�oI��S&g[������$o���F�셭\��!���t��{�d'da��P؇�c�?��ς�	==�wx�]��4 ���v�M,(&o;E":G�p���m�]�f6�
��5����e��HGtx��U��4��k�����ђI��
��? �K�1����|�1},%ԝ�m��7�a+l�+�B2�?@�E�;�gH���v�i�ɶ�����NZ��N�*(J������7�fI�)��׎��5]ᣩ����O0�EN�R/�z���� u�Po� ��E�P�B�A5k�1�`�1)�3��${��/����B�sb�r��}�����L� �C:,���U�"����̇��R�j�v� �T\ba�XlxVHYEB     400     200H���d������5
s8	��NW-�.�'�w)���[Y�Na�Dd<�yޟ|���oمY��[h�������;Эܖ�Rܠ��x������f�	�ѱm�S}���H�L�?՜�HP��E �ɼţjd��Q�=.����##�_@��-�'k�-�"{�;p�������jL����^R+��T{`�/{5=2�*�+�j��&lG�1��ĈZ,E������ļy��c��/5��A�֓<��\�8��f��q��_q�u��O�]��t
���X\�D����>>e���BW�)�v���雟���.N:��vc�G��#����5ϙb�l� |4�w�;����;UÓ)`��[���*+��������AKju.5���hb A����F�� ����s�%��o��Y'�GeM$U?@b�V[A���mmU��uX�����6=KL�HLŒ`q����f����)�[��z������/4�z���y�i����^@��K���+�XXlxVHYEB     400     1b0� ���hM���#�<���@E,��Z�G��I��� މ~b�������ۀ���1H��Ên�Q���]�S�)�C��C�X���&�����"0Z��έ���j��������^\��(��im�����v�JW��G�$�<[�ua"*Ty�h�ў�������2C������^J��;O�v�4 1�i�d�P3�g�B�{)Qd����@/9dWi'|ُ,�R���C ��0����S(MZ�0t�+@Ͳ0Ћ���	��7��cy����������آ2]箿��
sl�t��F���$��ۤ�v��Z��Q���K�d�)���E$���Py^+�n�F�5�����2�w"�XQG�c"��w�KP/BQnj��:�����j�2=q�R��A��nBP,<u �ML��[�=���*��XlxVHYEB     400     170	�cz���yv��/��W���dv�a�h�u'P�V�N$S��-t�q��]�bS	���5�u��&A5����?�4�EP�}�h��n�+E�y�8`�L�[���2���Ŵ���i�Rzղ-(�G9� ��}O���
&4,2��x�\��r��e������_�(�$��S��մ�\������p����i�,]��HF<#�9��G�4��7S$�������Z�����1ȿ�	�y�D�������ĺ�����	���ζq�6�j��(y{M��&f_ܓ�&OZ3�&�b�fji��e\Y6|$��eYG����J��v��Q^��RP���R��c��~�h�����#�ª7�|q؇�Q�XlxVHYEB     400     120�HB���<rt�mj:8�<T�+���we���M�*r\2�m`v�gRB�2#R��2�1�#�Dk.p7<���B�R|/�ȞM	��{��M9K�p%�r�pF��(ʕӯv%h�ӽ\1a��i^�e������#�̅o�_Q�0���ݓa��v)m��#sF�CB�*�ǥu����΃��	[�c��(�0 �p��#�s�_'k-����ЪI�v;�����껑*��n}_t���麬��(wcW��X
Î
��#���3꽫�ef*Bά��-;]?n�u8(]�XlxVHYEB     400     110(�8'���Cr�����]q��ï���	gǕ݈�ΔG0Y����z[m�
��٨��ɣ��KRgT/\S���t�o�N���^a�qQ��>9�9Ί9�O�o�6��K�{u+�<���\�V�:�?�B���qɍbz���ў�����(�R�F�^dZ�� �~6��������(�,��ށ�~�=����*�6��a�U��p����2����8���<�L��[�k:Y��G��t]�˞S}���:��E�-��2��*��ֺiXlxVHYEB     400     1e0-�J�<���Sݦ�m��]�I|�J�=��������?�`�M�UdJ"�*�0t!�W��?i�f�Ep&l9��u.d��S�U8��°FuJ��K��0�3���'���v�<p�h�E,sTf��_�ppʟ����{[K`�w��SX�*�4��2�b���k�@d��l�i��݇Њ �@��1ް�M6����$~��/:�Rf\��ޑ!C��?d��K vA<i��XS���#���ͺًX�^�j��L���\^�*���MUp~�I��L��8�:O��F3�˶G!��`na"�V�{tl��U�:8�:���g3"*�����Z���b�$^��#�&�n'��~�'���AP��z�U�
ȁT�MՆ}�R,u�9D���N�)���h�)Y��=��n��)s�*�%��t1M�g�Q�����=e�5צ�:[&Զd�O�U�4/P�:V�#�-5H��"X�������77|XlxVHYEB     400     220�ܕH�1�O�O���;<����_į1�ş0�6y7�Sd���ʡ	�i�2�d��)�L	dov6J#C�'C���BLjVjA��)�@�6�Z[HyX����UX�<d�X�oa}{���&��b��H9�h��Z��D�a�n	r��;���s��gi�=���4A3�/�6p.{rITóq��X㑱�@%��t;1�E�2駡�A3[�5����Ʌ"Vԑʉ틓�{w��uw��h�� ��� G{^P�c�C��b��k�����C�e"�䅷
n����Z���~�z�%�5*~k2�����\�'��`��	��S[�s2�9[���7�n����sE�­�?�J�`�F�n{^�L�-y���e��E�@OO�)�ʦ~Dm*ξM��K:���{`���F�d�D�Js�i!&7�T<����\�+Z���F�]lP������[\{
��X1��E���O��ᄨ���R9��&�BZZ�!���S@#(#�R�5:-���G��H�)��B#���uXlxVHYEB     400     1a0�Ă���z�Y�����۞@f�E�=��<���b$�C纔<���P�C|э�u`��S������ �X�r���7^@�@���z|.ԣ�4tn���I�uD����7gۑ\��� x�~/�KVF!A��B��z"��:�i��|�[���y:�R�(���!K:�A�'��N�G
(+=�x75��gE�0�E�gq$��o�56��(ӕ���@bd�^N;��6��88xp���+�5č�� _ )�;�]�`[ۤ�4�דּ�.� �#e�O�`�︃���	
2�� jKcY�׽���v/;7�J��u��j��@��A[����	Q��D�j@Foې�*�k$d�k�+�����Q+�@�;_A�>�4��b��0�@����Ȗ"OU*��h=L�.�R�~�}&2��XlxVHYEB     26e     130f�M�#�טc������)�<>Ͼd(+��`56,<O�q~\c�
 0���I֖c�
�H(~��%�F)JkQp��~wO:�{�,0l��_�{r߱o]
��'o�k%s�ϵ?���	�N�{�$Ah�����t��!���靺�����T�
�D7�'�����.����6�G۳N)!�]�6�b8������;�lB��m$�lD�����==nƭV�M+��
�K_7O����C�d3�8Swܝ"둷0�I<��_i�'�CM������p\��6�RD ns�Gʯ�x�O