XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\��:��� ����3jݦ��Qk�L,@�༰��%#�f�6�'���O��	�-��V��a��MH"�C�.f�R'mpf�Z4m��Js�t�ր�`vA���S���_ǁ�����*��G_t�zXh� ɋ2��z�{����jA��՚'l�>J�G c&sE��(Z�'��䡟\p/���2���Yt6�(��.��ֵ�oL��m��W�н+ ��w�*\�����=���L��f�G�[y�L�@��_��yYG����p#K�H/&Jb��@�ӓNXX� ^j#%�^��Ay>5�A5���C��,��Q�د�>�珮j�b@ݲN���Ke'J�+&�-V�@��,2R> y�ՍU��xH*b`�M	sOр���z������iSf��z��dn'�����]5��Cd5�=��J��8�#(G3�[}m�E&^%A�;
������)���4F��vDX�? ���ĝ����5�8Q�K�+�_7��>Vߥ���d6q����lP�d:�W��o���nWn]��-���YQJ ��}$LZ�I�^��q�#���sD�Mh@2*׶�,��!�q�~nw���1��͑�����[j��S�(��R���������-����O��kNB��΁%�Np���[�
�����d\d��Y���.im�S@'�B4	}��{'�W�h2��=_���\<P�O�'�|l�l?q����qz�ZF�_p�m�֢82fxR|��[�?XlxVHYEB     400     1c0dv)�W̞��������ߊ"�t�i,�^<J��E@�T[�^ 3>Hu���G���f�	I."r;�[ݻ>�j�z�f�͢gV�e��C7T��}?�bL��ұ��1?�ݑ��miе`@���/�2�P2ЍƷ���r�0fl�j%�niM��4�2��Ɠ� �川_|��mo&�cH��e�^��J e���h/�5Lj��~�)?���!���w��>)c���5����&A%!��B�.*^�୿�q�l/��P[F�����{��$�ٰ]���f��/���o	���ҳbG�羫Ο�����5+ԯC�M�h�&11�zyB�-4����WWj,���e<�=~���������[������}�d~�Gw��wU��gͻ-�Zwr���۰�i�i�%f�Kݳ�G�.g=�0\�RE��@�E�Ƅ+2�T��x��^����PXlxVHYEB     400     180t��M�Y����y䗤�y���7k]��/k=4�6�k3�*��7`�\�-��Ow�zBvt�bE�p������5��2��E,,۴�eO5�`_.�vb�Z��({9Y�|��|瀄ǓA� ��bj��ю��$������Q���K,h�P�hH1�UT��u���r�d��e�M^Z��*c�����Hz����������)���[�&�n�6�oSS�ov{l�=�E5_҂$\�H|��l�xiz�;m���9�V�Ğ����9��%?p=z������g�
��&�����cj/�C����O�m����	>|��@틈#2��!^Yp0�=�Ļ�i�+��F���6
Σ�}�N/ԝKo�1�b�qPz@��GXlxVHYEB     400     150�x�$k8r}K�e\AX��/��0�M��x�;A���˥!����� AS� �x���h���cԼ�"�C��O�����$j�d����e�!���������% �p�i̚��&���/p?c)!������B�֢��|��>r�
h���,J(0�~�ÝzBֆvz�����"mav4�s����my=A�9%w��L�5f��R؏������{�<�?�Êq�CgG�D��`(��~��,��X�P�{�#���o	�܄SJo��]���ι�=�aY�����;]�D��"9�=]�e�v��7�4�5hK� �H��PW4��XlxVHYEB     400     1b0��%�F!ZJ��� f�b֣�)w^%w�o d+D#�҃E\wz��	(]�;����#�ҙ;�RxŴ�t}���w��B�|5��5HH����ߴ6����H��O���@(�$�Ԣ�R�;�oPsP��MZ��fv�vG'?c��4�}�cBgz
msɜ�g��J�yy�
٦�MH����2�Xث�C��ض����Q'b*���"T{��}��`�	��el^�g��"9��QN<�q�� ��dd����������x-�,莇��o;r�����_&���P80|��n�
R \�B{Ql���@�<�!$>!��*���t<��`'�z7+���5�7��s���+�Q��� ��y�
zub� nT�q#wV�<"�T���1��/�����ק��xc{�h"Z5�Rʖ��	�-��XlxVHYEB     400     100�6_�~
j��OWz�3��c9�@t�\c�����61��y�⢃�������w�5��&��P�l6C�b6|}*�UΈ�/���B����(��O��'rώ3�1r�i�Q5�>�dD��h�����e�'a���x<��1F��c�Չp.�(�:�V�%R�i�U�X�� �[",�DdT]dw����]�؀�,\+�����"�5�q���wI΋��}�[7�����|�ܶߡh�>(=��M{]9ss�XlxVHYEB     400     120���$N��<�Ѥ���zv�#� 1
�3�<F2s.�"�	���N)D�hF�[�\K>u�eH֝���}Sb�����w%l��ڿ.���6�j뽷n"��n;T
�rM�b/��p!N>9		���g�ݰh���T����Y�C:n��Gf��o��:�i��b�~}���6*^z�ϫ�1�"x4���'�y5��b��8i_p`�o� :u9,�om	�6��8h��p���jz��IcNƋ�&�b<ȥz�.�f�W��S�\X��[��1�*�̶�8XlxVHYEB     400     160b����p-��:3%w�4Hlu��� ���2P����G�����klq��~�����4ZCH��c�\���B�#e�f�9x�"���!U˨aa_�i6�,B�m�ubx*���Af/��/=�H~��,���}�βfz�)��7X�1|�g�n���m=����o����Є�=8��,��p�,��Ȍa�|L��$��j�-7��HO��:D:��DZ�įy��zk�R���a"��(��v��(��=>�6y�P7�Q��FY�N4a})f-���6)��d�W��3���k^�h�-v4����9<7��7�[�e��I��ª�Ŏ2�~ǜ�W"�|y�XlxVHYEB     400     110��6饍Z�-� �a1O�Ҫ��}'�r��y�|V���ǂہ f�'����0�$ ><�z��@!��0]|�O���B��-'W����؈ċj���X���q�@�˹��z�b�Y�B|
j�:&]�|p���k��QGPB��U[h87�Ƶi5�Z���>Ӓdµ�9��7��]���NC�)^��<;D���Y��o/����d�z��bK-w�s?i9��:n�\T�#�H�����S�z�������npC%��A���}XlxVHYEB     400     100^���L�AØ��y�:��{5��'�E-Ʈo�u�-z8bM��XW܆�6Fd�S�MzND��x~��&��35����]�������G���J������Ã����fP2fk��QOM��__T؎s�mK��=�E�j�IGy�t��I6.L�ܐ�-��ԇ���+��ӏ��V�Ă�p�щ�V9A�4<�8�@�V��Ͳ�$�/��� F�`ѳ�����x�*3x��C�Ab�s��j���6��XlxVHYEB     400      d0J)����#�<���ڳ`lQd͹�w������IM)!t%���,w�p�m}Q�O>e$���n�e@#���w����:K�h��F3�X�`h�.IF���u��0�Gė�Bd%�0�
C̭��|�A^π2
����Uj��O���P�x��i�wi�s�P%���9=�<A�J��p~�pp�=�C�p5�j�<�����6��,�&XlxVHYEB     400      d0�.'��2uO������};z��7�C�Ly�!�A�֦4�C}�dX��d_�d_Y1��ڴ�7ױ�S?�GY�h�"��	1/K��"c�U���K�g/�&�S��]�[00���s���u�� J��8��Z7Y	�f�t���
aS��П�35�
�~��4ټ�����t?�o�3�8�N�����+Y�#oX�p��C��t��-�XlxVHYEB     400     130��s̲�
���L�lj���Ha�b
iyt7�:�j*U���$�,Mu��|��U���}�m�l6�ow��J��B/@�,�:7�*6��z���j�Y��qC��̼ͬ�b-���6��?�t!�Z��q�5�7v��f�Fgj�,P�\�����'�3��F���VL��av|����Q RU�M�mw�;cb�,Au�������~�؜��n���֩��hn��D|��;4y���V����u��HI�M&��q��e�=m�5�D[��ήc�
�����'o/��S��YXlxVHYEB     400     150 �WuY��	W���i��%��,
��ɣ�t�ۑZኮ�Q��K�VT�x���8�i/T���[�O�/����w�c�q���[���R=�G��<�����$﩯_K�ಐj �3M��S�g�Cы���w�դ������.3�A���DDU���^d���V#ҡ#(v,"m�Ф $��2^����=Ydy-F���4>ߚ���>�/M"Q��wy&Wf^�d� g*��h�����O�$������fF9K���YN7���MRA���a�\����31�����C���4�M2�W�����Y���+��u��KSQ�Mtx�XlxVHYEB     400     170��B�-�v���
"����y�H���\>�b}1yg�FZh%Fei�m�Y�Ǿ���<f��ӣO!�#8�iW�mS�7Gb��1;K��s4�� z��Ut�m�[��'Jd#s�,(ڞ0:v�� ��q^�i]��/�.��[��D� ��z����bm�
��"I�Ƹ�D�Y�2?v,�B��?����,��'��M�DԶ��J�P��j*�BF��N���v�=0.���_8��-��;4�(��H�jUmV@E��$R������Ґz�D\�]{���>A|�-<���Z�Q7a�!7�7�qjvB�'"u��nƆ���c�$��y�P<�c"���n��C)npu����xۥ j �>!Z�.�̒�XlxVHYEB     400     190��H�U6W�8�"�O��B3��3LXW����v/�¨�5p�}.C8m���h�@)���
�r�A��UG����W\ �T�
��7G^�@B��>�,Èpb���H�7a�'
��q�0�;�)����Y)��h��;d��vGB[�r$�E b.�:�qN�p7I�>�����y=+��eD��Suz3��?~���X��Ja�Rfx��+��{!sT� ��}���>;P�� ������ �Z*$��?s�M܈�L90*LB߂~ּ����~��������8.��-��)-w�p(�d��������� j%γ�=��s ���-��l��`���`T�\���PZ�\����'����V.zt��;˦��S���5X*toqI ��{�|�7L�l#�XlxVHYEB     400     180��NOb�v��S(?M��f��=�u�r���p���#=K�ʯ�3��tN�d:��� �?�8c�C㋣�F1~j/e��JE��d��o�C=�	�HC�qG�9�4�X��P�N��5�"	����l�T]_
�*�	����]��9��f�݊�*s�tB������H�t�b=h��kIar{��<;!ɸ���|}��1��y	�ڬ.,6N��#�:�a81�V1M�������ni����̀�E�0uސI�މ�f����f�<�Lc�XEɦ/�����,I�3�=*_�f���U�nx϶~H��Y�? B���c�)R4: g�B�J��/;�[[(��+����Z%K����EyX�I�A�hG���6���a
XlxVHYEB     400     140�Q ��ԥu��Y��"	u�b����U؛.�]�].
�X��}�ސ�Ga�$��6�9'(�.�=����bU}��zKV^�Y��n̶i�rI�~a�[F^����Z�E���J�op��q[���^��@���4�/[�8�T�$N	���������(�7-���Cx�d"��3�1&x�2I�b�_jV�L����͹��H�ԯI7�������[[�Ş���/��!7;�� h*p��S�ߍ�5�лf��r^ ���Eg{iGG�_�e�x�*�!�!!l;��IN�����8z����)
��j6P�/t���XlxVHYEB     400     130�DQ!���{17���gM�6�"?|�|�۽وv,  �43Ftk6f/x�2�K�P	�J2ޡ���"\�]�7k�[e�3�+YĄO�v'l�����������m�G���>�F����On�Rf�蚅�ŷ�e<�f�t���q'C����]ܸgk��*{��� pD�3��+���<)�R5&>87է����f!enXT?�8�y�O�~-G�|;��<(�Z�U�I��笧���ә�X���md��Uuy�h�~Z
\/��1H�	}U�|�W�0;`7�Ɩ�o���F�+��J�κ]XlxVHYEB     400     170q95�8@9ኂ/�Z�փ�S����7w�z�q��n�e��]T�J�����F9���t[@����}՚�ynx^�ME��q���#��A��ǃc�C㥚D�P��"�@�ћq������m~}ȗ���;Ky��G�gR\6��˃��$�7���Zҩ�$�z�!CKU5�Dc��dYRo���dڠ�`�3tѭ���t�**�����|��l���%n~֐�'z��ٸ�<���h�s,͉�����/��䱈�J۩{�RU�3K�̻��Һ�Q��O@R�������*L����Ѥ�y���抏����TnQ�3۰+]��ס�#�CT�h��d�������sY>���avXlxVHYEB     400     120�)�W�E���F�~Z܅�5k�zf��W@�aG�ޣ2	0FHy�{��\���ir��p��rz�9��A1��J����Bכ�w�mt����1�~GJ�J++l�9�$���-O��L�(������q?&OIw�B���f��g~A+�u�Q�>�B��szU�!��={�����y�ů|q���ŶZ>'�ҥ� �G�#��4d��W�����}w�ʙv,chEK���!�#8e����r��������s}9ŏ1��/O�z��N3����a�{�ͩw��$�XlxVHYEB     400     130t�qH2hy��G�ʲ���C� ߔȻ����ƙ��[��PP)"���Vv�i?$�⡨Q ���Q@��"N��
z�WTGP�%;��������bl�Pt����SC�D����E_���$H.�
��ٕ���PVgKW����
f���������RwM�{�N:� \XW��(�z��O�wQ$����$]�=������������*L���	�y�"[�����#�K=�k,�|��┍��ڐ�������ǫj6~�O�N�y�=���&(@�f�]�������i΄�9�������4XlxVHYEB     400     140|��Ʀ*��%nn>-�#��В@�Luj���o����"�������|�ֽ���(�-~�l1�:�ᆑ����R��޶o�r����u𐎲������Lű3��}��a�mV@���O�B� ��nb�����5 �e��4=����}�s�5����nV�G9�Cc����mٟ���������_��gLS�6+�ڒN�p��v>U�>��G,-hQcO�uU�Hk.�ڲ������>�&�Ow��8_����ᕣA�H4��4嵙��O�ݷd�!���.�O�F�>��p�Pr`�y�۵��XlxVHYEB     400     1a0��ȳ��B���H���˄voW�n�m��D�mە���"�˳��亥���*Ҍ� W�W���U��o����rE�l���ua���+[�JzUQ����(_p_�D�"�Ȟz< ����ߢU`$�P{[�������ܮ�tȬ]�1]/+��&��j���Rs:�F�r�i���o�m�O�\VU��PN����P����e!϶X�'�P�/PC�5�f��_��q>�)d<�$�LA�5b2��{�+ �A0�&�˧�VP
nY�1�8�T~���f_8J>����7Q��O*��5[�CϦ׻���;��'uЛ��)M�L�RD�k�N$�� S�?p��娪�;�[����g���Xc�b��4a�	>��Y*�v5,Gh�X^�*�Yx~&�k7�\� �mAM���/޶8�iXlxVHYEB     400     180�k�u���C��ԡQ�B�<�i������Jn�6ACwp��$��B�]�G�8X�ۺ��n��<���X�[8b6�C��I.��=<G���MH,�wi�A|�x���U0kq���.e�}Z�����3���(���:�$Y�{+���:6f"zÜ�ݍ5Ƹ'�� Sϴ�Mu�r�M�$�p����Y�2A���V�Zz�|�c�p���8��5S�l߼��:��C�~3��¢U^IΓs��WIi"��R�Z�v~��{D�+.�s�#�$�w�pLuI��.��ѷC�D�p5�U]��Q����򩝇<a ���އ,f�%���nU�ՅC��.�M�'�-m���q[�i� 4+�^�����^e���>��ڕ�XlxVHYEB     400     170.r3<p�(i�yp�7����(վ��_�F�+Yy�1^ȕG-
��hu= �d�	g��^�a;������ o���,�����qԙO���&���l�|����~9�	1N
����Q{�~���Q5�$��D�������RyPw2i�+�y��҇pZv��ל�K��O�"9m|O��'�^�d'%�s*IZ������W,~��J�\:�;P��a �f�| �PK����y�ߤ���2�^#c%+]���)9����2��4^x����d�݌V�}sr�1;�{P��
�n�m��$���)�3�����)�[$�3�������s���zhGq��fl��T�t�C�̕���:�U�XlxVHYEB     400     1e0�9�)ՏK:G$p������Cp����!?��U�<��S2��GfK�;P���D�P��`�Ҍ¡Zu{�7��(���G��l�uJ�y�B�xK�^e�1z \�@l�+�Ȅ[�Ft�J�Mg����@�H_�-��.��������r^�_�f�]r�Ѕ!�/�����2!gt�TC��P���U�s��Z�#GY2�~N.�*JVvK��g�Mz$�W�dZ|��� O��T�b�����h�|}ʡ��W��Jx ����z���Xi~�m��(/iD�	Xf�.{�SEL�ls�����W$`9�X��5y/�@N��O��-�r�W�hϐ���3|є���4d�y#����3i����H~=�`�wȅ��HL#2܊8/ᴯ��M���R��� �S�/mƾY��Fx4\��L��A�2�G%������@R�R��l��N>��u�J���j�����N�7�l�؞�I^���MPXXlxVHYEB     400     1b0A�g<Ő#A��Ÿ,�킞�7B���S(�����e�ƤY�$#�z}���LrJ�5Qկ��W�$�qߩĚ*SM8�����豑Mt�[��y{��g�.�;V��Z=��4[ˌG͵��v�p���x��
��'"3��?��vd��多���m�?F��.�j�L�UV���x�y'�#r4���9��q�*�� =��7�(��_��;A�X7�:!ס�XJ<.2���-\me���0�>Ȯg�Y��z@?C��� �{�}]�'W�6ͣD*m�{�'G۾]l�g��¿m����P�;F]1zA��wɛZ��FY;�Җ�Vx�գ��A�}�BQR�t����*=(�N뉵�?�p:o |��8�Ć����Z�0��؅��w|��3��q_`��hB\�0��IX��x�*�.s�XlxVHYEB     400     160
XXF�1�9܈�8B���5�[\�j�"��5a��'j(�ն8�nkSAHFJ�Pi�_��x ?��I�bx�43�s��Ꙣ)=��[o�?Ĉ#�LZJ��l(���M.�'�@���U4#i�J�	"e9�J�0�bE��O@�'�B��=�o����-�K�g���4p��1밐Bw �j�³�n�ʌ�k��a�נ���0ʘ�<ER��T�����<Hք"C��P8asË�
N�jq�w���GR��ۗFp����������bo6��k����'�gj��V����e���ls�Պ�쀔���Բ%�8]��ɉ�%��f��e�S�~�&)���Na^�^XlxVHYEB     400     150E�X��l3�꺯�G�al���4�Z��Q� aū4���%��m�\�a���(�����A�a�Ʃ}�q"�ޖ7�ۚ�����ҌA�^���0tt�cJ��O:T������ʰ���k�A3X�w�=&�k�$��@=8Օ���W6��ܢf��Ȍ�a\�d�@atF����.�`�7? I��f�j����-ycq�ޮ���A���W�}xІ� P��ߘ�����4��q�KX��r��(����q��ިa���y�B�j�d�{�#UD��q��2	��,�q��k[S�4�$8%%v���M:�YFWJw��{�DK�;8�� ��j�a�~�XlxVHYEB     400     1a0ف5i�_�%1x9�R�ƞe�/F�v�Hd����*����3gø!����X�y���'帵Wy����\���lW�:4�M�S����f.�kz$T��T^rb8��E�\���ƍ�2���$��w��ϥ��C�r�2�R�g��aX�F5�~��ݩ�ݜ�̄���7.���r��{��u��q���V'�ZY�˲[4�<�b���[ƶ?+��L���*��Ts*_���(m��H�P�՟KK^Z��j����}�`"d@�>�ԇa<�㎫���u#��n)��J���^c��lls�
��gl��U��yѴ��C6�"�xs>J�5+�����k��W�I���D��bCӕ���q�z�������$h<�3$
�h"����&���G�&���`XlxVHYEB     400     150�ɟIT��e�6�c-����-`1�� [��3�������{��n*:��;h��@sޠ�\ �Z��𽱳�^#�a�X���S�+r�:�:1�4��F:��Uen��h�-���ą�t=G����t�r��&lN�!�.�V9�!��/Q(�����I]^�R�,��_2�Ɣ}bQW�?-����.�%�@H�.�қ���x����ݙ��#�E���2]��xZٌX4h�����g�B�ƫ�֞vgs�s�P���K/ɚ�ASw8e��5���E�}�_:m�����lYe�A�O^d=�������>v�e��.i[/r=��JnXlxVHYEB     400      e0/ks������`}:1#:�`E^��FV�>����<z��:��Z�Cs����ʵ����MUN�i
O���QSA(#�dl�5+��f+�EP�/�tS��z9��&9(�)l)��}5��Dw��HZ!�Ð��9���P�
�`�9G��_��>���-!�i$6�l�l��!�,�1����2w�y~ŀ����7Bp��@�|��B0%Ihl��XlxVHYEB     400      e0��[�Si�����;��Rd�r\ㅕZ�����w��Y�'U���;m�6_�mW��d�Qlm0� �v�9�)0�]Yy�Vc��A2C轍�,j|�A������5}��u=���i'�lk��%��"�[ޅ�>-̜��JYN^q^O\ݪ��a� �]��dǳ��Uλ�_"���IWZ��JÑ�>��j	�q�l�)$f/$/{�qMzOYk&�RvXlxVHYEB     400      f0=��,��k-�:��bz�?�G2wW� @��-E*��C�˿T�;���k�al�ai�Y�4k���g��Z<?09�,̇�pX�D6A�K����;4i����v���]l�#k���k��T�נ�3�� E�U-'�H�4D��lw	q�D-�nt��,I�j��OA'm��K`W����K�㥠m�;Lơ���]8@f-��#��[�	��M������W|e�B\H�C��XlxVHYEB     400      f0����Dh�i6���
-l<�����R��@JP�仰����ƕMC�����Z%�n����6��:���n��=�C�0]P@~�3�e�~7!
��%!����&2�κ��Z�cp<3�
l~ol�2Z�)�T��B�2�1�a��ή
�o�fAm�+pXk��g�w�.�nʄ��,��3�G7�6�RM�V�[�5��;7Ao�P�����E6�;����h�j��9�LalՓtXlxVHYEB     400     110���	BZ^	�'�#��V��?�3!��:HrH�jE�iK(���{�fJ�
f���ۊ��k�[v��:j�!qY�>�Ȱ=|4�K�䦄��9�P�A9�s�y�ϡ-x����F�]��dâ����ŝJ)Z�:�EV`�㧹����Ԩ�*������]��z�������O%\$\��K����驂��)����o��߭1 �8F&l�PQ����.
���R�WP9������M��Pj+�3�U�����/S���`K��.Ń.*D8���d�{��XlxVHYEB     400     1b0��A'�k?��N��h]�y~��oF�hxGg��D��-��l�����A�!/������"�`�yu�/���u*xp�܄��z��"�]�GCY0@,�*�ԇa�Tc���B�D�Z�:O\��G :̿H�c C�f 7�S!abŘ6.\���V�W� b�p�Ҧ�+F����*6Hͭ�҃��{�.HJ�����j�4HDy�iƑ'��5O�D��U���_!��mD`'�l�%�`�e�NZ�u��+�V��߇<����~my��T6�${+w�}�r���-�B�
��%����;產�"�Bܥ��_`�aV	�M�ʠ3���0�>��2�����#0O�.O�Gg��3nC_���E1k���NG�u�"�2Z�U뼀�+}}� v}\:�|�]q��w}���+�Ә&�`,��sL�XlxVHYEB     400     140�����-$EyQ~w���-�A�ߊ}4�,/Ƿ+�Cb�!eO+��Ub���Xy��R:A(��P�����G}�ax�}̚��>aA[��PO��	Z_-~R�)��Չ�w8F����v��od���Md���!�;
!\���lY�rT���O���睂,�T�Ÿ�S�h�_���`A6\`�ИcgۻD�8π��$�0�.a���A�&�6��E��ap�&�X�̄DSG���z�l��}��ג,EM׮C9�$!��Jl_1�ҏ���p��Sp�� C6�<�����$��/E��|^V��bS�����xt�s�p8��[�XlxVHYEB     400     160~�Qx����oCᙡ/e��3���y}kn�w��A��꽿S>�`���Q�v�\vA�%Y2� ���&��:�M/�|&Y<uEo�bf��.*�x��U+�}6�>��C�K�>���9Ħ!k_x��_ݲ|�@�~�����R�˸}�:���=Mp�	ۭ��֥C��.7]��u���c �-b�M��ū��\wx ��t&[�v��f�I���1%�>=	�<�h��t�X��f����H���{�^���T1�&|FvQ��2|r�f!F-�r1�n[k���-����mH��$J�@,PSّy�.֋p�J��+A<�����le���TɃ��Mچ
	������x��XlxVHYEB     400     140�5�A��'�O���4��B� g���F	m���{0D/���%S���@�TNt���
���bw�+lW� !ٮ��n�\mm�����G���Z��Bё*w��i��`���zo��1Ҟ/�231��$"\Fi�d���i0.�[E0Ҷ�҆� {`����qB��Jx'�	���dUp�����v�ě�X|iIb��\��l�;$k"�����N����#MjIWr��<�g%���k��N����P��.���^��Z�m�.�����N[��ބ'̽ۜ1�&/`�Gu�b�=�ǭ}q1�&��t�XlxVHYEB     400     180�b�	�5:��F�R���ՄGs� ��~K�{�	>�*f$v47�~��{�T��g��}!<����u>L��|[�G��M��`6o��6A����������:��U�%@G`/u4��킄��5S�$���;	i���i�0�G��pPc�,���~[�I���T��E2Ϸzɥ��^U�a&�����{��	�FQ�$�Sj�2���Pr�5!���*��,��y��w���t��X�>�Ҙ>��4&�����&�%p�kS�
�6�c�(����D��+ih�wt@o��ܒL�x�bfņ�ːE�a.d�1�t3��-iƊ6��SѿYA �J���oJ�oC��Uy���j�pC�޺�b���XlxVHYEB     400     190���L�֬�'qKt#�Cv2lQy����iVV��<�u�׮9_��0 6F�V��e�e��[�2���:m]����b�Ƹ�j������^���2���C��5{�n�p����~:��K{��|ƛ��Ka�qx���#q�ifu�x�mBd��pY+&���`ϙ�#����~ˠ�� غ��2<4�'>�'�w�i���5I[�ER�g��fn���2�X���!,��(��c#��� m��(�������|�0����jpn�/5"�Uz�h5�Ň��7½���uT/jĨyPX�
�HK���z��*w�#��N[�>&�]�S����6����+��}a:�rGG�0&��P
h¦.'�!�����$��WS��XZo�K�u�T:m~@�p6�1XlxVHYEB     400     150t��H��V�)�	{[��ʄʑ�w|}�����[{����I�!-�g��y�o�S�~���NQ�h;�cH���{q����`=�K���n�G��/����7@�ӕ"��b\�Ķ��1،�Ru�
|ؾԠ����Փ}�f��-y��{'�D���5K��IFj��PP9t.��p����L ��߰ޭ��*y�"oA��x�IN���� ��	��bIc%6m� �j��nچbk��2���Cp�e�b�hR�L����X�rjdr����Sq_7��"+=/4�,���g���Z�{��f�ڽ~����I#�"Aӭݭt{}�~�8݌8~�~�CeXlxVHYEB     400     1a0���A����#�@����޼c�3^��)(�@_���g�$��lC��7P�'�0 {b�����I��`�~t�Zi��C���U�p��'#Nm�>��A��̻�8+�	�@�ܺ�7ֳ��q���&#Q\�z��E�=%��g�Lr�}F%V��Yw_e�G��ʕ�O�U�[�P]�^�o����@3��"eb�i�U�vE-+��_������=�&^�-W�b ۳��U�\�ǌRH%���m'(p$��R���M��
�Nfc33m)C���=�Z��cF����KT��;��=��vQ5fx�{�?("�f��d~��ˠ�)}}�`lV@b+�7g֨M	�e2�0����jEus��/�Z�J�:�D;�l%3 ��R
'���Ғn��7���C�����OC�;XlxVHYEB     400      f0���EC��q6c<�y�`��BҐ$�o|YqW����4�n���9v�1�ND�e���Q�:q��;0�B�ˉ���Gi���^��^�ԚQ���s���E�H�c�0�nSD褃c��r�[#I�c���f\�G��k��գ��#D��a�����{��,s�U�h���R�6h�>��#밢��F�O.08� a��r���S5�ҜOٔn\}�V2��/E*A��ɱZ�?d�v�XlxVHYEB     400     100�U^M�	�	K��S�(8�Y@��浃�{�R�$b;����@�2k�svG�\��Ŏ�6���kr!��~L1|J��yh!���i7m�lE8�$A�+�B�o/(��&�i����	��:�$�Z�2��F�1�VG�K�@��2[|��\D������ɻ6`�ǌ�v^$��Ȱ�ex@TZ�(U���q�/�=����xvS^�E�J���@';	�����nzs�=g�n�����D�����[���XlxVHYEB     400      f0����J��
v�Rq�U�ǲ�qan�$�D���lZo�{��7��Ɍ3�׀��lbV��k���^G��։ͅQ�m}^*:BG�8\=ߨ�\/�٭Nqh�%���P�s�'^�}gS1�.�n/��א� Π�i�`�g'�A�'8|�f�Ŵ�](��׫I@*Vc�wu?�&j������i�Y��ޝ�7��=�.y$5�Q���<C�q��\��*�{6g���\R�Z{XlxVHYEB     400     120��.	9��+�4G��}�f�
ڷ#�]k�,��d���~�m{#{	�hX�a���RC}>�&�b�/�4%���D���w3�����g]'A�/Oa��[�9�0k�gxKW�i�D�䫹$�It���c�le}@��؞Tﰤk�0%$�Џ��]�ys�����@d��8 ��k�s*�m��0��=�i��6trF_��l�P\5 !�d�_���Y�#��Q�wB�H�	�?�����D���XQ�0�L���4� ��̥J�Ȩ��A�]�pr��P���v�5hXlxVHYEB     400      c0��4O��)4�1�`HZ����a�/��ZY��� ��7��҃�uK�t��0�E���4t����G���}�h�5�2��;� ����܌�Q��Έ"���Bʌ�W�ԋ�C E�Gq#�^6�s�U����n���bК��q׶�u���rY������(����E%��.�0Tnn���+$y�XlxVHYEB     400     150zQ)��D������G�����J^ʍơd}����7_B���a:�����H[�ˮ`uN��H^�T�a?O���Ǧ�������M�(^�ɧY�j��
�Mrk�����k!)����W���.!*k�U��~;���i�. q��T�j?J�������Nj.���om�9u�(��n[8���A�*Ƕh� ?�õ�f�ev�6�qȭ-ءG��	ۗ)�u��Z����@� ��7��&���mM��=6�PA�����M��+�U�R�8��k�9<^Oð��ǋ`èDe�?��iӕ`�\+k��5w��!M?d"��~I�	����`XlxVHYEB     400     130�ױ�I���8|�����\�������3���q8�1����E7�^Q�Ѝ�iwS�Y���w�J��+�c|��\7H�{���;�\�`����ţE�s�����S�1N��Z*P֯؞��ۨ���̬|��@3l䒥l�7��Ӟ��@���7�?I�`�6��D@�g����+1q����?��H����G���1 �f���7�&́�ώ��B�&2���o�)$6mb�p�!ZJ���eH��?s�ʂ��$&:΃ΒTY�����`��_�55-�>�w|��XlxVHYEB     353     160�jY��Ř	c����]C�����^���0�Y/�����j0�g9�G�V~�V o�Zv�F�Xz��(��Y����<*�~`��Xj���Z�Y9����bSR��k��Y��uı-��Rx�w�ÊB���)!CO>
�3 M_���f�z;��+�c�Fz�9)�1`��@�t���$�\<�j��1޸ ��~Y�e��=���%��8�\�R;X�C��,�k�?F|EOH��$�Tt��](g��᮳�.&�_%�7ˬL�?�0���������Cv�� �Xh����UV]����1�'����D^T�����۟Y~U�Pi��7sq�k��+��8�}�#�5@�F��