`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
YealRjfN54m1ls+yAme904JYQtgPowGv8J4HMNu0s1w8vlbw4mmG1mbCT+ptDbmk0nZU9+KKdmGk
eLw59D0+2AFFmkc7MSQ3GpZO6Hd/IMTBCU2U9z9CqhxVvp6IY6UO5vfLgKEtWVuWUwcR6cwXv5wC
9hmuS7I7Vp4fgQRxf7C+8zhMCcnKyXGq0dkQs6/wWrmBe6efmZ2xRb7aOCUYaPvYlluXANEsQPBb
YI3W0cWGJmHGfvx6wKZsaxHJAlAXmMFQLBxknnBk+GT5BafoubGMvvTLbBFVbUyklWFcFeWx0TOW
575ChcKn30/OW+wv3XWokORj8vtanfUdH79uLZptCqryzws2VuPFALLZbkJBnAmhprhEwZ/S/FOi
xJsLdrthH6LS9+JZo1eNWhtPOeYHa/Nnq83bB06xTdCV47hEbPAKanyOWmdm+Fl7jV16QsvOyIyF
hqiBWS/5+mnOE2KnV74fnYjm5G8nI4E6tBqDd2rDFuub5u54DtMybLPEzy2wEZ/LrdF37rXCOz4x
nXFfWKVX3Yt65uv4hWfI0tE5kjVVP87Bfuwo0cwLlEELZ8ogF+tomwQ/Fia/cGRQUqKBbH3wo0s9
e4sshg1mpBzClZgI/sOkcgN1Ew87qp8L2ZvVW9vfIJlYZSY9t3e9E5WlBiE0Xzeav5PaWj5gfxTE
OBfFyxSSBjNklSOqauk0kDIStw3w+CCKtZwhZ1YSkAIMjmwy4Qi76llKKeoLTQ3ImCO/CBDl6RY4
9a6eez8GuMpMfAyYSEhYTCTK2wZT/rwQqA1pFM5IWblT7nB4bcYITeoIDkuNiSD8HpNMMEZdjweJ
hG5hRgr0UBGngtwp0MSG9LdTd5DT3/DL6ZxIu3hloXlCaBCIBX2RsWx6ERkDTVPU/+4H9GDTCLG/
aZIkpLjoWweDo9SbkPCReFhkHKukfOC0AUGgIc1dhLZCPC7KTUuvWDPWyaubWXWAMUlnJfqxM8xl
4VaLKnYa27YVdtDf23txUpGjNYoVrI+aa1tA1ahOtDYTqX9pmPMR0Wy3rXLAqQ/0q9rGIaYBFt3L
ZdNnUvR9fjZo8yAY6tsGkgz7Sx+eR+iZvQco4e2MVc/li7bM9lURRi25xwrQ3GXE9O9Ygrd0oqPL
h6FoEHu5v4tpQJXRijeuPLQw2iFdz1kxll1jT+2ZidFQ3lxOLvas7liDnNzwZZWEIKUv/Gjg4f3C
z928Du0R5JPBnGGEhfFrrx79KARISXixo9R2VxFXFYTcaC3enwcJSet3eHGHbLnMEtzSXjvoRjGF
+Y/6SBkmUuelypwkv+uP83XDhw8pHUN/oex8N3LztGNDdQQifidwH3s2rKOqBU0m94h9RYnZc8a9
79WVxehxs3JyHy2n9yg9eaQxSD6wzbge2mNNZnYthcGr8ZAGp1wygDoiE0D5/JH/u7+88eysfcT0
Cd7DXsuLj7ASS5cIqjw9utUOpf8RoeXR9FMZ3Vkr1nRRF+iP/oWC7gNVmr/G4peF24teBIPDy6E1
cml4Z1tsMzCS8XZT+jeo4HusTnFEAq+h438P5aaE4umd+jEF25dqBHMOS35j3qewz0XGVpBmt3dI
QM8T8bpdhFkywzTYcm/MvIx1lAmc5/ZydHn8XapaOBWI7L+k6CrteTS6pA0669EgDmCMC748ELWC
+QYJ7xyluUk6+efKwRl65jMuXdrtEOV+MuxU2gZ72vc6H7Lct5oq3QeYMiDYp0QdRYx+q+zrI8VY
02WRotaVfaGIVF8x6M7CK5JO0/HIcqoGDuABMUkZcj2omdTdw7p4W1azWxYeXqdifM1sPZEQBt1f
+FjZA1scakOzApgNRl0aK6zXOVLdmcClSzvgGyM9Xx+P2ZMwdQ5E913L1pbV8DS4+yzVzKZuu26O
QAkdNEcJbTPhDQ5nBVJ7DcpXqFg3c7yi9+fSAdtXI/e6XX4RNsCfm2px4zLG533aI6ncGDmZq47n
6+eZMlg1xuBAoXqgwwYNQbzqviIUERfRVa08fnC2Z0xiE8+akLKgN8Ucso+JgNzrIK6wL6L+eSn+
20I3QNFrphdhuSMW7lHLu7i5FOWq3HQFlkg8vEkf7AZcClv9XYEnshufrVejQiE3ikjsvKK6fPR8
GVj5TCSq7gmPPGFR8q2FYu+nVZSnz0OopEgbP+NDOzuj9AptVbw7nNcRyyEuKNzaCEdhnmLuCzoY
flrY5xI8JCv2jLnNmas58BocWN8jVCpXPGDjQThsj5MSOha5nGOpxmB7awu5Xa2KKIjyc+CE0xWa
eIlvS4aD3jVLsWQFGEhaGQisQww8E0moRRA1MkJx9bghAsNtl0dA2v+9wHNJ8y84LERBbPPx0yS9
i+UjGflhloeiDO72fhOOPATacny+Il7LA7CZwICQ4QNxTPh0Ha/zAJ5JT2P/+JhaIUQ0XtwzJ3qL
yzix8wzLyAHQ8RZvwg4Jjs5+QETI9ih3Tl3oBFfRZl9e2WfTegMEGRV3Tnq/uIIIS8EyEeSyfkAr
21tJYmlIwfwmXVxTe3vmchd2/tYoaIHh45I4pwWjl6jE2AibUoKSiijpSwZ5+Ee8FVGc0/0Laokh
kAANTrnX14v3Wr3NhDuwgdOtkKnRHdbhMYfloh6zZUbnu4WeT4aCnXuJByeDDWF5oQmYCYBrxyTh
71W1zFhv4UlmSLiVX0TJ7TafVlelmWPlMlmKISR1kzBetmyviQpUDt3s7mTchfUbFeOoIq5dc79B
tkE8BlTIRlYgT7T1pQVwDIfakUhAY5wN713N7vjbHOY2CNqKMHO4r0YqxtpPcef8zl5Sk/0pByaO
BFmYgDZRMaBwsU0zHFNMSIVjZVqy1DrYQla2ImsPmakW0sgYF/8ex5UUpB9XaNs4S3tIkskXtxZX
J5tpy0FiX7Lk22rvHQgODtzjD9J5M+nuFeAcZsW7cknIgF8H5uT6R7LOtxVJjRluLpbg4qEUbAds
eWOLa1EBmM4uuOCFW0++gUbIUZH6et+EUH8uTy4Sc0UL+M3++gpLNUb+G07YQw9edCpwW/jX1Me4
VPJ+JMuCjSopqa297cxCHOpK812+p/R2NsRuNHNmCd1QRyOnXw9T6A3PnQW9TZ1x69Lo1CecJKlH
zTQz61W1jaDhDwO+KQs8pt1Qw3ass0tEqAROmvoG8UJzjEih4ckzILaaZuErA/m6fXozGBrsLVmM
JS2IVU7B2aNZvlb0Ay5wLvKkEYLqK585mXmiV4G+6sQjmp7dNeIHq8lWEiA79dLyJ8dmQw3u1EgD
QXQ6h8c784TjZvcsE4wOyagcnYRmUjVIdb7t1W+nXWyZVsMfPAZxC7csE0+uqDLPYmsk71SADSjG
4hJ3U9s4zBMR1Xw+3qSaHhfYeBLRxeUCREyHa021NFes+pU22t3DiYlkOlLp5rcEr43RFD+u3Fuv
Ht9HAEY2u4DfKQJLEPwlVVMsiBO0lRZa89tRrlQEONLbNq6fI3jzrVIKlyifysOX9gmFlyu9h9HV
N2wQFj/HJZdiS8+JuvEAneJM1vW0uJviEg+LW/RhLCzGFZBLJ2GmHKuPlyQdFiGAYesXtvDHt+7s
6IUAf2AXrrIhan/RQqMy1f8eG35PBqO5mFHvy7sa/2NX2ASNsH2ZIPF4PDBfCj/gs/eQDzY/BHHk
/HzJhDQ8zlmUK2etONT2XLLcOp6BSPxqLmFfXsnlR3DFWEQiFi9/gQBVbd2b2njcS5MHJWvc/HV0
EyA7fNSHWg/k6BEHeu4NF9tVs8gwlSh8NrdH0X+DKrbXxtNI1Rqnk58PcKSWWldXe+ZjBPXGHUMX
hxMJG3g6t/TCs+qUzLsxnDls3A+Qvl7y5Zsw2rNTgrNXwc04KDlCM/0JEo781nyxMnDKce1NUJIz
jdlPyzSFHlGdQhSWryB1S8yz6mLr63xaOW4lOlMtDj0Z6SLdMBdmTQ77UZ2u2jQ7jti6okDNQQP9
FV1zcVriBwTuyqIW245OAWOHe7YMFPwnwU/F6ChFQ48ehx2wtI/qAxZ1LF9Idp/4std/eUOkzWst
XDzbfTCSz1N65MpAix+w0Nr9WofiS/rQIi0H16dyvjAMbmtt7GYt8CuhOamV1PI11dyggp77ifzw
Z4qWiO0A2ovkNuetEgSt65tNtwKZQTmOpAFmDvYRDcdRYw1R5hJfW/4dGcXC3i/qcgzA9ptTqpek
dmygCuso8j17jAji40QLKRgasqvZfOsoznhfHDu4/8o3NJowF51VGDQZcsBLnbLoDIrwyT/CI2WU
AzCxAxLHtxDT3TvFK5bZth8QmlbGkAVXApa7wlrdNo007qF8uZ2ad7fZddfGg9jb1ubIL44xhZr0
1SbYi9rZ8RX5L9BdH4ejFOb9ck8mViIDv/nkuWl0pA6V/d887H5RgqPrLlUIB6+r1BmkVu1h3DMS
Y5PuW6pdsHzq3PND8uoFbfle8CkrmpUQWJ75UuMxm0ENkvYISJMC5mwVb0kbFivKs/lPLXVKohYt
CWjqgKOMaIaHJ/Nadil27HxPeAvBZazm0E89U00eU/QYCb7PEUI074uCI1byKvUJwWivmMIwKdqn
brHqp+Sd6NWNI6hW+7JYuBs1L16NknU407+VQf4U9Ndf5q0Rurwph6EqAaAoVAJm4EPqAeH4wo26
NbGkrPeDHTMQ/51tkSBGgiztCB8tFpTFGSfK7S0oKA+SoekhbifwE+yKj62GDb0l3l5kwViaNaAp
mA9X7gTv3nUHiEQgzbZIEY7Smra3453rerMK6aHfrd1hGKbI8jrBmxnYXEA2IW4xRw4hpBwY/QNI
ipt3brh3FHytZJXvbNX4JtMoUZspDnMhYq1gzEsWLur+XJXwFQS2yeUXX4zM64bbermIsY9H+PFZ
Ltw7RC97eQLCHZrg+n0U7NnJGeKpTxDgBpnWKYpFgD4lPj+BNKUfM2y5vggsm3ec9WCzPciOjVNf
vhdwP2rfYQ7m3ilkWB2CET5s7gY1PKwOU6eIkfJBGEKd7Xl2wqwyJMiXFoGkP5VyDPiQrL5rfqXi
r1z4t4I09NSLyGz5nnJI7w2JUBtOAx/J90Vimvc5mP6Epo2R4e6/PEw7jni2FcsiuIpogPFIeSFb
g70D+r2YzcEVz2H25RZ246xwewiTMaXCuGjK67Won8S/PNtVltOJ/l4Qh4vrvF3tIQAtvtVERKu6
+dkZgoQ7fNo/HKx14nPz9wI/erKRyb2npesTem2Iw1Zu1bSxm2hZWw3DBgsfnQbO0XrMlo+B8Ua4
IZjIWr7RCtllgDcZYWciBxK5gkk6RzmkE59yNGsoGHWgkWebzJGrww0i4K57eEj9nO2jpYnEI6vT
fz+MsbAZyDYrTDidc3JTneNqVC8P9oH00Sk4iFpwqji0lV9etqew9f3msTPIe8f3mAwl9ZgCyKdh
b5m6IR3njwplrc5obesm5d8IwV09zS2HmQS4Vsfwod6xbpbW3OgJfclOphFJDd+wLxhYEP4t2dx4
uM8fT/uJb/hg+0HK/zZZftEozDRx8yu8nr3LhtdBBI/X8bzGLFLN2cXmYX/gRal18htOrdNwlJLO
kCZfP2qEtMazbUywdUesLW9gpSZiWSmwmBElwfAYx6jUf6qLrfWugQ3U8wuy0vyOpP7Ox8KJByi/
gl8fZFVp3idCE4VO0iO/X10PLH5ZUwGUMkKGKIaCoNZADjEeOi2ENZy8SqB8cPCkrJ6ieWekVklL
BmE6RXold1y5CetoPGbELQiku9/eUXSnMg0V9JtBEY67Orw7w5CWX5aErJoOYAnddasgUs7BqDXQ
PJNzj7ZbLPmQW7fYokWFvpe0tbzTt+GWqxxe2MMxPWS9jUR9GTgj6FVDUWlLeCNVEtH2PETgtS99
+W+2/IyKV/7ZWyTjaXPIH7MkBpgf2wrfhKq2t/NEgL9JYJqQHn8Hf+g8yx67Ppwitk5EW9FLLzNP
19k7cxcbgSniE+quDW5RrIp2rZziXqgVom2sfMk2IwsmTHD+zwFf1/WzQ/yAB0D0rb3Y2kWGwrFR
Mp8rYQAgFbXdTpZ5OleLEvhb6wEcXfuFMtLtwLcUGHKS4XZQkFqMLCULRx0iUjoKnNY8WGj9Tcav
0yrXZoEdBZPAsurGKqliAC3PFXXg1G2qmztcK9lDrgaQmi5f/fifBgX1YHWBa7yMtezVI3tvYg+a
+cBt7uHjUgubDiDjwJ0G+peAyeU2HSpBDriQ6avKrib5UjCneqNVPwxqvMrECCzIxBJSralKUMXy
viCQjF/Nr+4ZhrsprcoN1jiXM5dJn93d2J6Q3DGWVF2rJR7frNk+Gv/wVR2IeHlL9CRY2gZvwj5S
dYdPpjemG5JCYxgQaSogtinQq90CA1V+Jb2STnnq9MaZVjioCzZ59y/rSx84ZGpCDM9Kzua8v+IG
BHm/MptRJZxDHtTd1Tq7nJgLoj25FjGPa9qPik9pfs7LPaxG7uiqrfs0eiUm5wbpTKLPAHWEInLF
HT9gy3Q1oUfqH808AzeOM05xd0M9IIOxXH4lTzn9AR+kX6C9ZfgGVO2j/n5bDsFPk5akXOe9UYlZ
rMvr36yytTLQEtjGfMUTlhJxmWTqD7/Icdty0qf++J76DEK2SbmfX/OPmn2jGJOmGcDnwjF6YDZ4
3i4YVSrLXMRbuJClzWhpceGa9/afmaeb3iiv1p2SLY9iK3cIMm7mz+KCmfsJsQMuxcy4xKHgqm+w
U+MgiJJxp8ha2GHMu2NXcRBq0K3Edpe9veFfi/oesTIEd1R/Ktk9oPmGNCZjb3fq5V2QEPopEU2G
eh/OUm7dTJtJIOM7wvIsIFzZFsH1Un71jWYzZY9E2ztSU/BNABd+5oLEX2a2+sT64PqTnPbNDE1h
zqWUMHSSc3WJFmjlryWJ5qjwO65JpKBh0HFy0H72XGeTNEHqCVqi8kPvjIahheERBbcAwv98OaKP
hjhctWH0FM1zi6Yc4X2IRte33uz/BAhBmIaEb9l7mWyncsiSvuXp6k8XztyDI+QL38vBv/AIjT3r
+B/+3l6BpjVpnfiTqoRrZzAtA1FfNpU+J8szZ1ywG2rXgB2YWOzva6l74hdcKNGwy+7Cjn07ri72
F1l/gMbjaP+k+duakiE1+/OxwkKeYcTZeMqku3yUIyvapuT0qDJQJD3/28p/XX5/4h2px4qTExJ6
53bM8k/2JT1RlA9D9RsZqL4tLxAd39QKGIs9HN0Vq3InsHW6XhMQUdsj+6NDebJ9vtRVzbf9PIi+
dFAchqKKsf9INA/mv38RfD6+6yZLuZnpiJcU6a95AQFTQqQvErKxUmrc7MMHLIc2Z1yGGdEAr2A8
spAi5ckruOrLpum7oYRMlP7wtSVoJwDRGb9bpwltHNLXN2sWrTk3W9Lj0m5Z7rkLgVsJA/VzNe5C
Oi1snl7AUfpNJ3yr3cbuUwC045jKBo5iDRJdH1o4bxEXhgo1ia2n5Tah1z202L9jNZ5a56aDWm8i
ODSQQTRyrbwlyiR8KmIj4xUQYwoqKkkb5k8PrIxWUIQjd2I22wbuYg3uDAQDHPnPjoFy0ifv6MWh
1HHNgkFrzmRCoLStEcVISZXsG4MwjavrHPuhzn1gCSchE+hdKAU88oGnRyha5O0HolldKO55BW3c
dkinBRVr357WB6o6xbWQDejev4bDkIgG9tJDx3c+fS8eB2xk01B4mR9v1TZAk39CQ0kdU7jFbNze
lAob03whu0EU2l4ikTgjYVurPfDiTrlH8eMqdSWD3Mfbd3sXZDXkIBIp0FrebLmVEjtskB+kEC0Q
soUyVo22lscJ3DVfVz/JH57z1bl5Jtrhkkw5zOc5FbANAx6HthuGv37EgvYjd8UTFX0ZQFTHH5mY
N9JtitofvYbgIzldfk744RUXZZ/lIX+m7v61xDGpe+e5LOUx07lLGtbmTg3NERCtN5OiKUnD9eXE
EVjli7mkAd7Lha0XlnSyA4wA2D1syXflLsFm5C+AnG25JQo7B9jIy6lNvYVfxs1UuaVZIYLqtBeE
7u6f3yk5TcZDan1idutPxKbt/6pN16Ph3GVeLh1N4LrMUC43vulxrEq4jbgjJSqyLHly/Yv42Kep
KJ2rPhTWZb6wkuxJypG4Vi7Wq2KzAWDSrySQnsZHAc/x3EX7WtjyBW6RXsc20uQJAaQpQVZVVFux
ySwBoarSBnejW6qZ5k0AvVfEC/wHDdS0HnFFcJuJ+bIOOvt029J9MPhDBlbLhlH8XqMd0hB8e2gi
sjZwPhSfspbjBtVU2ic/19Se1MSTkKRzHxWUW3kBPVO/JJtj0pWbRY+z/v12z7uL1eq+C46NonMU
rTSyz0iSKeOAxp3DPJk5unLroJ+10UY1iFSeRclAosDP2iv4JBWUu1ZFbTha81VobA8Rq8UOPEj8
mOh870B6K0H9D5UTBqvpcq7+CJ7Ky0EHQcOKP3oddZdJxOnqvQ6XRCHDGgaF2df7czADnRp9pjXv
2gi+NCx4/vDl8Imbj40GuWAA0viR8SVmNILzG66ldxnfGBNw1Zcn1jhc7QOsb2bwMpqTXDzajAyz
DznF3TyTl18C+1EA7sjqclO+2aGYmlMiVij81dDbLoxgOyk8/T8nF6CNJpXVHubDWvZHGuyS0Gzk
4eebMJQpBP+WJKdB4zTsMcoEDGR4rq1TE9iRtxshwbe5AVhvONFUvGEi/DhtQ/sPwRYYhqG8/mrL
DM+JdvEE9RiSxRaUp6u6V10KEgEqgUSLPRuLbtvEKRfilsjtiRh7wHe39XXO3d/SF+EOmohVhDpO
xs+pBCIfnqM+P0m9tD43O5nimkypfC5l3DxXDida0L3/Rw0LN5VS1cT22u6CjUhG8RjGrcqJoY21
gbzhc+vbyxNYOccZyqTlx/Hj/eby3le8Q3+dBba4hLoJGyLiX1L2ZPDBejP0mlJtjcUxxjOCMRbt
nHah+EbnWZqWk0lDD+m1bLglz1QwLeZER1WDLFNNKlxvCvtjujkFTOlM2cQXq4/koztbtLx9ljpY
2tkxcOr/2/oY5qfYA3tWrowilAOinYkBsXypnNOFGgbyUlDMo+UJc54xTbySRVoFAKQE1PBy7qgH
i+WWQJliJNdwQsuwVDyt/YhInrYrhl/Jp8ooAnIXVUyQ4bP6sZdK8jXOWRH6NVxpzhiYeDfvxwxv
to6STTR/D9FNSAUQvebt1MfmuAjZrKXW9o8DZf+yu3VM+iM+rHYf0VxwfNte3MVbMyTy3Zj+Ozot
jfZu7VJ0CXctv88QaxnvCmChl7eAHPbJcVEur5LOLN1Oc/iJeFz8nBbe0SINUDOh7OejnHOX6vs/
Wdp4Qqd8L85/Sk2c0/lIiIXLml5utJEyVi5fQMQWG0EcDQ65VJWnXn4EBtrHnQhEPF6gS0acbBf1
vYIl2yYrWXrNTFAEFXXhlLJEwgo7pzT/wA9OhbjitpFKTOsp43tVrQWiXvEf9g07RKfYGjRBib0T
MvXDM+7IKW44peBylEaYGDKStyEasrSf/dLxQFnl/DjUbxj0CdAcz7eFxGRaClt1ZJ+7arJVY+3J
HRfBFO+528boBUtLQ4UFUS0NmvrTK8dDZbwKkkRwpHAHz7Cg5XmuyY3XEa0UWfug2iWZUdfaaxaQ
10/GgWCliWvYDrzRYt6eOy91gZYH+g1FvY/lGYrqjhxG8WUNjS8sNjyQnvchadRLGGRKTJcsbpYE
J2NwOqnu1hrZ8DVhgO+7mxNRXR9Q4UYZ4vZjs5Shb1c2slXbK27AcL335/5JK7mTgSfnnFN9AbAB
l4nKeYIh7xgqXm2EApfuqmszXnBopMMOw5HdrujGIWn4reHsAXQqvNUcv2mW23S9L55kB6FjPP2P
QDpthbEs8Tzg2NjsJvfPnrylWJyCr4/A828yrV6KRFkT/syAWVkotkSuSxke40n1LmONrxK6xsRZ
77SxHPHoVtFz0jRS8mbNMppuekIY1nySheB+tTO+i64qsrcq/taHH1BJWoJrmu7I+hXqF5QAL/4m
o8FOBzUZRqhmJY7sIy1dPM8i+hNLOVCN9ty0gSbfxkXFdkNwe9EvXPhmc0DSR5HJAmmhKeZJfe2D
NkA+QsuAQDPfh9w4DxTIaOATXc91r4LnjLDCSx5g6jq6EhpPtVRaCKw/quHAyNEPePNxWXhB1KUQ
RRfzyORt1st4F0gm6ZGNT4XHQzj1qxNrm8ITwA7AnOZtZyWJtL3Tcie049x8JynQygwS+u3xa2in
W/Jra8N7qeTazlGT0+DhpLaMavK0Jp1u0dc7RNY3VC5XbkPpUeQfT4JThvAag+c73m1kUhSDlaLz
PM03Le8KoD53xIZ3vHXc+Vllpe++BHRvreaVWPHUnjRi3s/lRKj0QdRUvCV09RW34wUCyo3c4EPH
bwkVAtf8qSKGB3f77xqycgdfJGhR5ncH27MyEEkLBXZ2WX2jCdM7cYcvRP25se8ciTi27+7Rfo54
kzBX9BEuUP5aCKfL3dsignkWIWByEBVDB74jkzcZgFu8078iPNy5qSM90f787sypmrPa+vbYHKaA
Bfp6Cv4T49f+G2N+KL6nv9FKFhD4ol/F48RQY5OWJxTGDY6XHU/06qV7Ur2g331hiimEMT3eWHEG
/AyY/I49uedIk4P4Mqhwlf93NHqy6/06qX54pz5FvvtsHOaG2R9MW9QQdfGqhu032wirTiUJc9XQ
sGGcDf22m0u82WBlRX+DZvDY1GCLhJdkEUZKM7Wm/jSi8FbrvwM7TWm+Qex7J2v4ypX0+aT1SBE6
ihl/DNInPrKdmfPmlGg8qiS+1LDqAdd8UHqab5AZ2VYnk0a+ongZLRirwqNbc6Zh+0ZWNhOcvraa
qVpivUnVs2dazyneu6xyX7KEB99rDiu1mKY3hSpk3YYj7Lu9CtBByIbHs82Zn/lUYKpAkPayVE4o
sgH9hKbRnRA9hlv37sRJFs/0W/uMHLCJm2Qb3MLWANrWDdepl5XgdlfyP5kN1cZ/5TpHJRBKNejs
7kegLU5RpEFfncpTEKMxnj9DgE249/WB+WgIQ1VoEJd8enIWKGsb1OLZm3Y17IAy3yN7wPgMdr7R
obhRxPpHgOFiAaxdSywRa/jZ/EAX/rCXoT0jiongSh7RxfCcq0c/+wq6ViHkAGDa/dVP36VB3l3X
FyfdsB3etciIe6AQWhfAYm0j8+fkwH3ZUbIc61orPz4s54BQpHMZFyVjgM0NjF/g25pZIs8DImNV
s9cKi44YEmlBYgQPVfXtWDbz57WhqLmHIOrt7ZxuiGTZOnmLNa2E7dSqpxjt2YJS61Cqisg4WvAe
Ku9iDsqArQ+sdht2oZUwchPdunN7mpaJFggqw6E4S0NOG0nhdCwUIEoUP6N4Hg3fC7uCmkI8+4z0
ZJ9/bqqFOaCrQaTg+NQtBIzlwD/dXCEBZDXu7kx71506XiNG0depYy224wcKSNUHLQcwIvpV48k1
mtuQoWJhS6VRPdaBch91+h8nRvBAr8evAqNGq8CBYvY7uSbL8/y/emi8BwQdd46WGwo3tljkG43o
fP76375ceGaac4/1f3/9Oi+oEuo6HH48O5jR6fGXhzhuAG3hWfehA4pj0S23gqvjiOKL2Ad0IJUX
KpqWJ/VDSIOqmjnyAPE7HOeJz0qrljIAFocvC98++YQRIb2ikHPKVFhTpPGNIuQQY1bVbb4dYPHm
b++2cJpRF3sCLlDWIM7RhsYoOLcZYAPRK0OMnVya1/XDSlgtxqQePj7GT4R1E0fH4CW+jZLtj1tI
nlli4dLJtdLQOPdCeLbuInirTfl6YIe+zdlQEXNfTLCPEiLZZWfs/PtVfXUyFzthl0X31e5jVcIU
bduj7lnJ0NIqPf0rU8AMGVsEWmKbnCbEEmIGSXmpSv6Z9B8TmFy9HFd5Zl9PCvVBFXOJ7cLefBmT
afsMaIQr4ytq/pkVuJ8Id/12/UxzHJmb6SJJSewOEJmxWDbuZF2GBVCpneLE7flbw14jB2TPVZM9
L6S6S8/uukOLeSjLTZL3VnB4qhEBV+AIe/yQhbeqL2s/b0bWWXwt8GRk/8Qt92F1HOKRojWvv/mR
k85Ej5DuicMQZOdB7sx8NKnePX930ugI0xvSJsx5pD2Q/nMoEAfthe/3e8rm47ybgwRfyu+V4uv0
e3u6VcW0uU6zC0FwlXrgHTIjT6MPNRvGmO72/0Wx3RGS/ZOxdKdCQBYnUJWSVIrxq5iw4QG4vlWI
tLEDaA57tgPpy5HOb36764P0uJ3/LPOQro/nstILzcmcwqibfthCxJzb2q9afoF7q51RhrUL5DLM
/IDExrDaJIuaQtPf3wnC2j/8HQjY3mrVi09HC6pjUtcGJhq1+oPTcsFZ1YkpIUd9ckIm6evQBLL0
zry2AX7XSEE1/51srATdOWKKR1OJ5aUqAk+j9Cw+lwGrEMgoL4X8QOeGMEc3ORW7HyKJIKQGj2tB
5Jr5GeTluxYV/g+znJBPymiffpmRuqN1ybq5flIOYCAEvxtlen5pH9D9GpxkroOIMnRN319nbCLT
u2NaZFUQ4aaD2sz/pcQ2c+EzUdNy4jIjiI7pfPbuCYvT9iSTzyLQhmIEYBvcL0AcWLEmyVnkB3bI
B8IYj2k2w9nxrh5TPR3RC5rPwvN7s98gWu8EqsaGoHeXwQd/6yvFdU8axKkBR4FnHJOzPBC1tWjJ
Hswxp/xa3HyYFmD2y0PgZyPHqNE1Xp9uHevlSHjhfq7gzo7R8Gu36tqT+Gy4L8KJLwANhq7ofCSq
I6bYp9Vz+s5emXC/u+QNFO2+dEPSxXEnuW/7hiG3moX6myQkkTouCudNW+rHhJhVNofjSyLQOeHr
4nmCs26ym6nkcWPqZ682sbCdcHcHzoN3TbVyXjeyIw8uo5V5ARIU6ajU/ZZW1Zk1kMbe+MB9wd0j
1JVJyL78eOV6+qnRUVmtuPFygVcroSN8Ix/rVEoIpRbUoCEGMajHPXIv9k/yI/cJlObVGUCjzQV2
7afAbKi75q3YaZk91Zb7E+2c2TzC72m+ynlFhbeC+i8Ym10YkvBN/6yQPAXKWCaNEcbFmn6Y0ZlU
QJ9Y6cqtfg+D7kb4CZbFRW6UIre5JVAvLyvBr2Iaf9HDjgybPS/SjvPleUVYtX1Ku9akuST13YlJ
EuIjSogxByLCHmQO0+8pssLd0zg7RYPkXbkkUGF3Q62eJfdLhR+dWu0XuY1oDJ2hysA/BEZl7rJq
jAVKekBRz2SVIgCNlbpJyIqYRWpnRomDlK12dCLoQdrDy4bq6QfN/DuMMmWHqhRWLe+/3lxzh/cL
+pDYmYM6Bog4t8EkgIObcCqxBcuUfljkjh0aJ7+5WSANGvWeFhnNekcPzA4vRVoiFL9qJiPtLysS
xZXLmvBfQImkkL0O1DVMRzvBUcxwBK7LDxb598/ZS8Btkscl1qbo8GYgtg+NB1r5Axdpp6xglp3e
5IloAqv+tSItu1QOUD24jltaBZUQ+Ml9DTl/X63zQ5UcdJBRzzyVUvqQ/8AcByxmTWhEiu4PQob2
D+wePnvD6J23viMHGf7JvNcjGtNqbsI2Lpce+7fSd+TOVKIe1S+gsbZvqaskIjDdlVxtHf4hmvwv
kWS7QlzRRd0W1uQhLiruqxM5AuaIKGqEvYam6tg1G15uUqeTCWJM5la/opTDcvYf/SQOqE/ldkUL
jX6tAvt4Peokl+10ml5W1YAMfeNWyQedvyj7Sz92tB10vR9zp1qTqiQ6o4iRzLcx1vqJqI/ysjFx
DXQsDD7GffPMNjSB9jXkBkIE61pkUr0n7RnDMoEGwixo1D9INiFdehEmEpqwfBhe9aGbQbDImB6T
cvwGXZZIZu7aRNbnUA3OQSmpKpDITxL2OpiGQ62CZTrCxQwAScPpCfjZSr2OgJTOkZ6ddrZhhcqp
ePvZTCF7Z/9bNUHpiHW3R/CnAJCUeJpbDnP6ekh/Eo1X8ybaCuFl3uUmsWdB9160hsSLnPNOMd+n
4l/Yt91mYSO4Ld7mm2avbnaDxz2GZwX3TCf9nMbawqYqfe3O7Erqbzti6wjHzwXAqVeukUISTMiT
MYXRK3L9UcvWzi6MrUaQnax/7jTMDD0D2JEodK2VZMHgnK36MveYj3cPuf6YJ4dExz72mvAPG2iD
arFFD0Ch7vZdOX1MK3uCGvwMzik2R2dP3MoSo44BQKsK9mw/UsYnDqQs/kZ9Qhbhj8zvBQio/juu
LB3paXrq3tzGrBGS7QzRtC2UwQ5bSO2v34dWYhUErwHk4ArZzH3XpnxCYfFJYyH5anJ/dfSq4EjX
AH2rjaR6a2MYm8jdemxKN2qoEXz+v5RXI+o1JblPJG8kpyQG1WBP7FB57LIlEzrwGg00Bpy2ca2d
zuNetbvc4EI3/nlgdeMMuf8TR/dQnfQmN8bmCWw5f9DKmBI6NH5jjZk9XrT64Z0wvgBEJDWVU/75
f7CcYxxzf1jsZRWxnDp4cHGfz0/8cBMsxaLcqX9nwBpf2X7Ai4D6Lv2dCoQ8dnCP5Y2iDwpURt8F
JdGjzIpPR/7j6XvxF0rxQgKEQ9ZG/NCgEcgVS96uBeeMVVnDIFkMZyKImqK9Y+waPeFPdME/XZ0m
lpxszzMXllmnucWX2FlqKj2MUGAifTNw7yhM/cj+iLOfVlDKp5jk0uSbXqGlM7QilZHBZm0ZgT15
LU0Hnrug1QObFTBYmw/dUi2w2/jkViuqCDnRZNxlt//j+nGL2ZfVSgnTzc3A5PmYC+kjswNVKjtG
Fe5HkJqMyHqFvEx1y5RaUBI2vR9lRlQUhCoe+FaIJLpafCbGFZSOJQHyUNZTNbW+jq9lhwOjEkRu
fl41nIlKi9luYEMtX89+fdKOkdilffHWrZgaq7vFPV+NsiseEcBz4M2q4LB2n04/SBwZUMrS3yKz
fj37O56/Y0RUmelceZ75bwUXGgUVr1awtNpvINUCDclHpLAUcWhx7vNnFLxZid48e5yp/46TuOzj
v448cSYqkc9bDzcsds6KW3cTCGf0wxGf85RFKGEl4rWFzFDf2fqyAuRs43OudHcF3Z4KNgDsH351
iSK5DEZWhZJGkTtga2q8t+K66yIG4rvH+qmsXeF3kI+hZKvqWesnoyUpj+AXPsDhWm5OkU40NhkP
rzucuvVrNC7sptG5QsO++2EBTJMStTiFFFMwgrnGbOpPtBzeosqvw9LVTiFFNlRuHAwzHVGPeeFy
SChEiosFqAUeUCeGB/PXV7OXU3hcfYmorpG/9VxU7q8qVCazChYjBOEQhXitYguCdh8ODmfrL5kM
wl3vU2VE5hTNBeHTD+cdqz2WS5BBVHA+Nhxmg7JS5jE+dx3PdiM4rQbjP6pjO2YfstqODUYyhmcl
CJeup34ce0k/eSYNpCa36oAgmkKz6ErWVmIXL3e5wnSpKKDZJjeJx7zRaMl/PxDaZveEtZcgffvl
HlRUbpNjHMX4JWwBbz4Ks4YSr+M35Vy7crN44/7T8hmpS0dnkOAhF9IkrB/JTDJkfhigbxgFYBju
Eox1iWb7MIEWN1pznSAvld/VWSSMcY38xAGUIwSbgdAItoBI3LvTCutoHWvJl1Bgxk/XW4d2aUkZ
Q5pFOYfGMRF8N13Thpdbg+3zIpyiVaXy6mRSSTFfPd9XvjMivBPxf6TkUsGh2tuW7CUvAWRDkjlx
kms3YVSSjLyn/oSfTS515FjVnsmAeWNi7uegy9ubefmPtKApoGenRWfJ+v//9mFR/c6CwQb3XWwE
63oHEVSu92F+HoUFVQjRoAf8V5EorbCbMPRqXAbuhRbc9Zj6zV0j7pse+s5Dvl+EhPE78c2iBoex
yhvAHmV+QLM1oHCT9kMM5qa9JZyMofMdvixNdtJ8CmmgiPHwdyvuce08U3Ivl5aiIOAabAb0ipCa
KtflbSia2QeEbY7JCY92S+7nF8jpfVIc8Ic4EOZkQL7VFBsX+RuRqHeRUU8isQ8q0RLJadamZUAV
sX4lfCqXFftoUHtCnh6ocUhaRXMiBbYtpM445jPMvsmhgk1QHgOficss22H0xUKwsDE8ntQvFS+O
tR8r4tFAkMBNqAhE0sRVPkZb6TsCyLSzHVfKuJeXNMTHplWv0Ae7ZsHsDKLbeg==
`protect end_protected
