`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
E2p9gl0dgx+3a4n8siInwdNVZ6k9f+cnHmsrUTFS0aaZylR8s/L5Hk0yJSbtfEBQPfCSl4q86oIw
uxZMoNAcH7JIoR5r1WzgWW/bDuqPXSuQkWfCX4RcaLt6JIxTINM2RzUS+wuh7rBOhiHUjZd3RlfP
BwZUh6QvZKPuc5ZMatGm5X3VPE+SuQ4c10mwNieUATT8N9RUZAyrWqFcOrQ/w3Ja6gxYg2/RZzjI
E5K1xKzWBreSRRqwkOhGUKR6OwIxpd5u39+9vNc2z1sbBqrRG/y9ZCOm0xso6Q/3XJOCuiA0kHPa
QgBmTTghu1YbF+VoUeJD4F1WKWgg4J2tNlu3Uw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="iro6JjmbNoNvwDHwTHk5yRrDvIAoVFdjtHJTW4T7PCA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7216)
`protect data_block
2cI+p5typ07UHO7ZW3KK5bhZOSbRH9sqY3OFIRFGKKAE7q5W77AhsZcsqPCwupeX5F3nKmYtdlpE
Ih6YtgopX7Me6rUQmI7nJB/4QktnjIJCfAVydWx8kMhkB15Ghijhe5CgzG8axZvw/J78YH25Sv3k
xHpIPKHqHJGlyMSPrIWIabneOWtcOy/DiUHxdpsGXrYcEmYaQpbY3N5oC8WXt9OWfIim30I+EpDE
AVYYcJgonCuWIMsFzrckdwiPeo1vt8aMllgJGmwvmjDQ4YaHVjUjOjzGgCYyqQ2qAd8EeI/LLy3Q
KodPuTD9zVy5ly+0Fe1FSZY61yQRFNtPWE9w2IkScpsZ1fiI7zSIRE6VLeOJAmpreQeD/sVpGCsM
rIGMpjbxxDvV+kHY55zTGlnTIawcRtYd8l3J8Q3zvcFye/5iSkwxEzUFC/r5dVBq0Fun0HkZM+JV
NJhibPgiPA7Gnnr5h/9H2Xms/ZvT+Yvt37VEoJvj/pdbM8cX9hKpBN138ezYrnheDnmSXp8kVXVO
zLrKvCYjVMX9XJlITy/PlnC8SALen3pWzo1klC6Erbj2rijBdLY+NqrjthFrQnHSyElSP+eO8puO
L4v7i7J/ZrANlYhGuTg5xS8RhBaut3D2sImWAAuXlST9onkFjdYHTZekFZK0/+ir+W90qUr60Cua
QmvxVxssi2BAfqVrxFvVrVpTTkVha2FXrZPxuYa5gokQvcGMBH2wOkx+/CB8DxUUtePfdBAP+uKW
wjhvcxw7Zy1nMlu0bfvSQXuLx3VXljKea7wSpFmFZUi5KAkoDoTxelAhqFbskHZn/EBPUGGUXWt2
e14HWpS/E+BEnwMRyp4ywduiue/LUwQ2G3JhCKlPSXRr7MwMPWFEzFCfXGo/87xniie0Ykg2SuLA
j++CWOjUvVaCMJgVioZRry8klFtSgDUKltuFDWREZwHs79sdXily3WEu6b+AhS/JDsViGW39XN4k
UZCS5wKR3hfpz4KR6/PjqEc43RzZZ17Depol3/0kF8abx3Gq467OMcyRP6XCOlvWKmvRmGm9KInO
FON1z7DxydoODWUY2fH9hMlDN2tDeWcPgIWIDZqqnzhZmp8eLm2VYyrzWgiNLnuPjBsmTcgJARqx
FZEUXUcoC4fFZFFyQ3y1vlMJxdcsiBKBRcMgUlVK8TDiYWYWEfG9NedVAYswaboAubkZ0NMdskIr
xwv4aPmIpQVmwOq5E4fmbPuT3t7KShrDjYwtRtvFuOph7/NVFgBawXBzF52ObbyeB17HQIdvVAvm
3RWDGvvh35KGLjh+e6ShSMVhZCeubiAxXKDkJOkYKj7vsfOG50dfcSAen8Sx05QpOxmzxiTUBUnY
VqUaWYDTzrvYFMG183DroGk3Ju9anoWjGnlULU6agJIKVx41cijlR5056I5qaP63dca/6B9r90m6
JaI9dnQ19dPBDb/A327q3YVfJjd3Typ56HdMDEgel2m3RYK6brB6EsDvrX4GxZsFZQMR6NErXUNC
agU8HiM6OYDLQXBfOb5fQp70KkGi8YX9I+kS4siNZlfjWObctd8a3+r13ozT/JsBTHofoH/0B3lL
f0rHnvjrTK7DSntoMwPqfaK56xw2yhkRrzQqaemJy4HFtnZDfIBnnsdYIhIu1/w4RBsyYBQJJGSV
/6L4DkoTyWHKnq2Y3EjzoTJ9zmVJ3MmZpAmUrMQthtxsU896a1SjSE5kg2kFybPELwHNe1XHuZ63
4Rirs7BibHErI5EEUrauesBjDbvaZFKOyo0i4tlT93FqOjUNZksbKEYqq2QhiRyppYecXNZHBDk8
X1x4y+vxNAfPHgeX4cbHy4r02gC/wHn8RyOPf6x1jnsJIDKWTbQqYdw/kfr7FYYp0kFG9Ey0rgNE
nDe3P2U42avujbyNWTkX6HfCNtpmMAYSxA4lcvkDIc9U1KrdV/+pxYLc0ylJGnLmHOOCAuomRRgh
Fzn8swhFRrLItrB5kjYNJiT0KS6dN9SXRutuobAYzpI+nUL+hwv4i4bf/vAbEY+9r9a6mILxAQEW
hWNYoB19fJ8PznmJlghMbROLePAk0eWmSVeoEK0oTlLbNPq7UGklXJA+f4cWYBX26TxHfQjV1uwE
porfjAvOaExFvrEdknPWAo1SXtLwHr9NYm5ERTtL1sf/41GrLXTR3j62OvydGOh3L1OCpJUmMpiQ
McnZaPyIK/06lX58Mxobbtxq9ngEaaGdx5P58jF/OyspfqT2UEyAQAqa7BLtJL2mJVs1oZTimEWw
02pgegn2n3mNg76eTDqXiL5M4v/M8K85WP9hVb4IB03FH+9pbfRoL29EhWNPM3VTc3KYj6QOT9cX
gPpZM2uih5l3lrPYDjivxdqbnuShcSpj7D4FepJPVUrpvgRl/iRkh7CkfQw0akekQkfYFRfeX4wW
6Xo9dPVQCqxS0D4NQneZrqGPjHbjNL1vhiIsVuHYydzL6Dx+1Ygza5Rbmdqy1KeZTYSUsQL0TzvV
uHCsGM2cnUUNKxz+Pj03CSJ7eYEKfc0z0f8oPklz/TBrLZvFM283JtiBmLrBhOxKIwUOg1nYTOR2
3+KTRblUvRdiTthy2c6KgepDLV+kBRkjF0e1wmA0KBKjg5g5y1/hOOfD8QM60XKbdT570Bfx7RTi
ZdZc235DdydLoSh0dEnVQk4upAZcaDMXequEEBh3u+fN2xnggsxzyhiCGdbX90w0GbFZvgV4Ecfu
h6CApjhbg5XGhW5Dl5AJ7Ruq/u4h3d5tTgbjMEeL4wNn9diPk/PHzUSHztxi4YjlNiMJI+UGOBUZ
YLEXBZE1FIVbQq12Yq1iKkq8PhAMWJHEEovc0KSMZAnpVKBfOsoBawHHHhUlC4tLxexmla9MsQxp
+hQ27xUj/LTscpOdUCGokvjXqQ4tj9EZcqKALTA1E5Fp+FB+cvBu9DoiDgFSM+CN9zoSfNzPIsKN
1/wy7o/9jYk0qIYQl/WsUGyQGSXLDyi+gJteR827gXHPGDPzF3mPtU7AZaRUMXYw+8+K9Ki3y8Rq
ns5gDh2y5fSMv5/7cnTTCH3SkZ7xaRlvJgCDCdjg7JuQzcpoCb37hts2MfRXLWZWRpWw0lQWpAYx
YNj5RKy8IRuGtwpNmH864E8YlEb7rmNn3nZ5ySDF5iJc7T4jk/+JYSENFjl4eOWWYBuGRbVxQ1Qi
HpKP/vmT9tiEu49QcIySBS42w5ixAPp2D5aj80u7/eW6yEaP561Eb0YzFSwfSiKTfSxltN+GVRcm
CpKRGrIkgMT98tIjWsd80o+3Gc3SpHQs7b501HamJ6PR4GgZRtXZlUv50uTi1llJfUnn/yzyyiLT
9YRffAcLc0509vSR9hD2zSUfWdGZ88a0ke+oZ5G40pTsh1Q0Wk00ljaNKAQHLvf4t1L5cRqDGIyK
OTJeL9YI6AYieWJo6g+aysKaspiSMoTEs3H5vpj556sop0JYVhBu57eqlHSKKJVRHXbSgxTfFF0A
lwjACK8Ev5+By61p1AvGmSiSzbUJFp4TJvetvUKW87ZOtv76VKWJG1+yWVxeRHn5nhVMppFwDfxA
XngnWedf3E7eZqy7mNAtwGHyANyb7SC9WP4dwvmcifnaxEeOiePY6OogmZLMULycr4Ca7yAymuH1
vEXJoRuD1sOwq8r9XYDP9lFXZhfIcmvnEQ9iAx1CfSRhmikDMH6vo4XlA3LC8j01LCm2+xrZ+Z9I
N2OxcKQcIjmOyAdses4+H2FGL9NcYnWdWjOeqNTc3ybUP6E9BypDhs8cSyCgz9uP+WWLd5YHCvmZ
9QBT8XSUIdJ7f+I3iOHLS/mjkUjtA+NzxUYi/Tmp88rm2+wL6VlAxy0OeVu38UW3bEsqWmxUcE4O
73lEgJ2fSVdkqnvbdZ/SxRhwyixDInmKz9aO6tnt5tnWD30ogh3zccHWGrYW68rTlk9kk6r5P6TR
kkqP7UtwG7xj+mk+Fy44s0aKEaDL3Ygfg7NSW+dgPkJmapCzcnwdvPuiA67Bh4dLu/WlNldr9Yne
RHvwtUPQqWuQAgUc3ETHoOaJ7ySjwQW2IV6XX90dpckIlXTb/KGhmgRanlKcDxURCkA4JfwbcDZ1
CHp+MDuuh4PTH64dcWvg5SFJ5+vG+8iUOZkL9oZa45ckGTDt1GS8r9L6yZu8+ltP2sp5FsCqCgZn
YvZLw7FAElB6I4C3EasyP8rSYb3KFwqt6bm1qOuFdZbk0WetPxQje04iab7w6qAgB6mOvwR4fU49
veVnNUpbKHWzGs1PCcS4Cmsa+9biNSBi3JqqtX2ECs9mmZgZg85zMpfhouYHqu4FTpytOKqL+BLZ
IsEc5MREgVO3LnBjR3FoVLiyj9cU6Lx57jxIPK1rqXfhnEArLC9/HRLUgvyRtkmMkrVtsjrMGZA9
0HRJYB/9In6LJVUjuQ4+bSgXy5LiF6bOFnX5Xsj7JYLVNi3z4UKxGnpC+lQ6rSEi3HhSjF7qh7zC
fHQbXR6tdnKmzZHwOdcGEYy4bAMQHEB/M9K7UhFws2gTwvC6BSjXJqbavofjSCLxFVKMN1lT6DIM
fd/wkafYr7IkpLIihpEwyt6Wt44QcIUB6NZgCATYdxb2u251LejOM2u1EYe7TMY0yreE9bVKYUNJ
jDTlU1gmyW6Ts35/10yWdwG4zqoAm/QbFNgUgew0SgcwOaeVPG+Ar+tVKIeJUipM+AbL5DOQnqr/
H79FUdFfvUPxAInzWxziX/qGM2aWww2+DdDuekpXUeQqlSzSjylI7RPrBwKesfPdho+sj/pd+WPK
bdZaTPmx6a7/8duryzzTZQbNMwsAlgt8I1JxGnFhxmgiJby6kS0wm2zlx31aCxW/OnYD8i+Iqpkv
CoEGUkbmnUGYi97ftPZu9D1whcFtdDDD5q+wHRf8p1bZPB4fLjsTFSy2M8YgGLEl/wf07lCxaEka
kPwofXmxpjMFxmlqtEIKtNUx+4nALyoOfrTsR9+4TY6BBdunjdo7TM0ppgrSOx5FIr1TFTIQTDJw
ZUWZonkxPWayAprpzUrS8LqDZkX77QCjIFkekgZZ+pBCajw22X7GroQr+yM263/g5aDE1YIeWB+o
lcPTjkM8VjMcH0ADov1YpkcSzocYfEE+5o0ghFf/mm3EvlndlNpBu2jvbYP7Ix3a8vLKMA0urFai
AtgDF17IyHiXrt+v321nM9AZdPC89467zLYf8Z3VRa1Ww9fJdsHSEnv0wiJ1wkjsUQ+4Ye+weaxs
kQFxvM0/syCQ+ps02dbfMHO4spdxaJar7oJ19JuHTSl1av39i5BE6ED++1lTQrcGutHLWAt7tvNJ
J83YtHHM3udXeg4DdCtFUB3l0t0hUgDGvZYYyipbYaAXJCvvkidlBz+D5eb7d3kkAJY52TPDgA+4
jQGIbUjOaPaJw85UzsPGeDduEEpUvTLWGXqqqbyYeNKpgtaz0o7CiRs2XMxuXn9x6MR5NW95wwVA
aCwYGZvdmDrIxbwl1WF5BUDmS2NpgYURScPUrDvqiguKblWZAbtJhe+xMMHd5ddg+MjbHtcOqktV
qXl5nnXwRGygvdAy6s89WkRJTNlLGfVQfo25wyY4ZeTOZIQioF5VID8GiztH6UkiVDbSzONSPylA
2Fon4vtd1gyM7JsGLci7/REsJWdHr+R6lWVDsQtLAnJFudVHPt+Bsh+JUjtyP1w3SA+Z6KR88aZt
6jMQ1lLYX7ujcoY4kdQxmBLIOxjwFe/tvZGhUD7RbNvOAV/rLskXRMUGcnyvfgaUA2tc/d1wZG7W
2H4qaGmWEcrQSPh+zoBquGG//wfaauJ6fOhRq+5c64oSc4qNNzp4V9OcE0VPmoEUEARriSdgN9hL
m5Ve2yvfEelSXxBBkJ1n+BzJZhJWcPuj8PwMX+oqE+HqZryQEZNIqnphB0MJuXlY6SmN6gWd/SjW
ElhrskMimxbbPcVlntjTC0NrrG4LB5TyexhEbPZstgWWllykJEQfkib8ad4y2tE+B6I/Q91T/dwX
3sbfQyKftDgWHrEMKnRNSWr6kMtHt1Cqnfhc/XgqsQmLHo+pZIUjoOy1MhdXKl+qjuhd6FMPLMbA
F/kddF+Hc2Ebn9leocjL4hER4gOduMuVBbLPYcnbCcKC/h8JXdDZ1srLF/yAQvzO65YJjhJsiSk3
GNz4TnpgKIT5EipDum/2xN5YvXRF7kIYp/f6FYZsMPa+pJgZ789+lst7iHoEfw47/XrCT7/1JNYD
bnZ3J30pzdjEjJuxOLndoFVGfNLk5NuGcX5duJQSGxIr2MO7WKeIZlh/0SzUpVooOdLCVek3Q9nc
Mqz7ZbgUzPEII9ylcHoFJhIFdoCRNqU7Tw8RDrOJVBhVnAwPhcz6jwlMS6f/dYSrCq0z2No5j/p0
bg6MbYcxItP1U4RkCS5nF9/fGHiSNyiIbFYJ+ZLK3qyOIXXXq4z4FYPBwZ6IOyHQ8X0wprKG36az
28tCHq53B4MkRFqX1xwx0r+U7Fwx4byQzElzuR3hMNf2imUVOl2igpCaMy13YPgdoDq/0bd81Adi
nlS8eX0LeEq1CYmgKtcrHLQphDJLdHAgwFhF7Wy/Cb2vccgbzj0KbqIXtCgUaauJLKIHmX8hsXAZ
wt982uo0WZ/9ZSMnXa/hUuCR0e4A+KbVKEMyKRW3z4980CJHUQzgwaTkiRlLZtPLeL9W2DFoTxWQ
bhh9OU6Eq+iIgNCsitpVZh8+JvmFFVkUXQP1k09cwVnQAFaX1BWEqLr1L4N4RZRdK7KFym6R3MYI
wSmg/lxWCdQKia/lcsxPgXtXmMqvXYRmVaRyh9/6ILc9pJdnKPHYK16Dokwpr8wGd0mua3doXSwb
KsBHS61ZiyuXGEYkiYV991pxSxoerfYdUOVCOK9hZFgl1ELN4xtWRJhfsYvJnSVCyfUzRU/OIqDG
xHuZo1PV+/PSIjPtBvg5nyvB5dt/Kx8IiVWfnMbYnHAM1/CAmScmW+s4wojHdv6/iXdLJuZCJ5ZH
gNsZE9ckO+QXGk+3dsxxNPZl33qnbEyIM6EcFUL+Y4Q6MKz5TBLrsd7ILsDDmJaN0uYD+ogAfUhm
M/lU6Lj/ZIdQ2vrE3L+kbGbpkn4pZ7PqvkWlRXKzPTSMcdkmAbPnObMjLwwTvTfdkh7MXRtK8C9W
ueUawNECC0OQCAUXnwFHcZnzROHq9W0chOxqV+L9hmNZSagJPjPdRE7zYhRMxCkCFA2bBUkR5M8/
JI4T6Aj+DlnHggawdxWOJi1we6v9J8w/LEA+1IngGXlnwfevd9JYLbet2t/Z4rkqVj/+liu5PmEF
ecEhFQnTMhku1Dil6X2CoElJUSuKZrlxgyF+M+TWGTzS6PL0dm1EMAJK5pUXjlN4DIGCM8UA2XhT
/5Io6OCEvgRBaBRdvVYQekioTYo81PY46JGQDl9F0EIxWBhtrHTEnFWW/BBb4I/uMOCi5J5YLBUc
a+ftsc1lihLx43Wj48+m2jnb6CYuFt5BykM6yCyZxjbh7gr0dD6VrGhh4H61kdlLbW8sM3rcg/cx
Cw5zEBIVbEUBr4pjTdLeoNNgZ3Y8V/ZfMiWWV9sFVS8jCx7LCNPnBFzpUhD8FaeXbDw/xwPEApQd
3EY3wrVPfDE0kL+P3o3/XJ6zzwjaPYEyP8bdj5ywA7HpQCMRJAOAA5q3zLgJDyvQxvYIPKMx3rCW
7Tw+sOX1P5OVGXb1uiNBHWhJ6CDMKFDM4Q5PbzvQgQHwFoiMA2gx7aIjSfTnPrrGWubMVnefXMW+
MGFoCa44L18iVYa3DzmAALMLJiGxcUtpcy3iqk2FIUGUOPBMugsi8s0RK6ovCxrTO7pT8ah3/DnN
ukHyEjSjCVpdzW5VztO6WdU+1X4htMARAvI+Y8twnz2vak7Paf0X1UWpLG/AGJuUWqUEitHuVyE+
aPDLBuDZBCw+2VdlmwR9JXoY5+OxpLIEfarFt65h07ucs3A4xXOECLhLSNk1U99RQl5jZmVlpTpI
PwXVdz5G1dcTl+FnLwUB/sfUKpxajhS95+wrYsuzpmyA/wfwGWsmHLuZoDDl/Om/Rtw6T4YjUok5
ofg5E4/C2UtpSLGzEubBijnd3w33Ue+rfhX4J4pb14aH7LpaB63CXfS9FJI8ADObblNDkhPZcSPG
eKK29MLVf6xW9jveziF0ABtV0UkApLqiNx+rMCn2HcbPi9/3ywH3yFS8BN8arlEeLxS7gkJYRan8
CCOOB5v/HOMsyCErR6VgsJfq2uy1HK/5gtb1zFTMlCXcpoQdAB8neUyD082kgfL6Dch7AxeM1k0g
7RGCZ76SBfzjfeeJa9HXO2lu5S7fJgsyaZDCRDzP11psZQRrIm62ACgwRD7Js/r5oaqdSxTCdhcb
QJ5EGyRb84s2b8dYuE+M7datg4T7sc+ggiiZuhWl6FFUqaYwvivnVl2t4OCqkK3YnWe+lO5+pxPr
YcKR9UatZBVAFHff3B06HU0pIaAKAgxbdrjzEW3XP4oWHc4BXjKvy3D3vlXMLc8gtZfa9/IHcaYL
3+F+HA2vpUY9fa5OpsGOnHVt/++T/gxTdXc9oCZ1Fo3yupTpMddOPSOH0EUIVlzBkVbWb57MrIDH
A+snvAqhKiDxTNTb8P88DafNzjhXljCzSV28FADSAazxzuEOJjblg36nc0MjbwlWd+LBrctk3T8q
WDXALYTBYNfFjPhCyVpu56MG06at9Dap01ZVPPMfgf8JxRamUKR2A75ohrmR/0gxsOW90FPppRhK
Ptk9KO9RBeHmc6vE8II1TAAt7MS924Y5Ilxeomb0MjFQjqY952gnOFO11afrlR4+/K//z1AGxrNx
0WRRVh08amlhzV/hy0hVnr0eMJp3aglnhC/JFiRp5MYHDLlIhxYUOGwQWNAevrd7/+V2jbgmbgvx
52SxHIQNR/igKkX0lteLBsyQ0/1UDtV1anWlNFUuaQceDJO6EL/Ordx3TGUDjz7fTa5naChrARFp
MPmuSZ8yuRlD79saVRXmEVL/+rq0QgDJyapcM8QJ6kY4AJpCxRlp0COKnm9rXSQT2I30eTlZ3gJy
vF5anBCiahK+oPoMlHJh+3JoXuzLoCggskFXjeiKEViCv7evdHwPUxuYgbWmsT89UIT41fgm9d5D
Qqvmov/SJFaSMkbKfHxCFhekJYJyiCd36wLCDTHI98qBVlbMx1jDlKloZDe2P1WVpm9Z0wSF0KtJ
W41cWQ/VTJWF3MoWmToULEGAiwuqUi7sdvOJ+JESKYyvvODpjAwcSd0OFoZMrUUeyNVqFmxbwWyY
ZPDqbdk7Wn2I27km2S0orBrd+qRPCstJnPSkc7M/Tl2DeFccokBqFb/5UGBqN2kR/+SGGdA7R20B
rVIv96/FFGNnl/1X8VZAjNveY4Id+LGHBKxygFYPSfAK/iyjvTsS3R5+Fde5fOVJdnLfIjVk6RHD
Oj++YtCDCpUDGhRgTY7Bb5uYKUFgmjQb7frhJSTgz9fXB3ZD3p1Xw7ByZ72MPkk9FtO61hngqWzR
Ywnni8r+W9R+GXatmP7G7AOECmUFdKOtIyZxbCVKfByaebm1JfGVm3DucTVisLKnPqKFsIyL5vPm
/EIMr77H1B0AY4Tot6xPZ3eDhBL6MySi96jI/ctGL6Qg9w==
`protect end_protected
