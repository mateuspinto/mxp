`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mhRXhGziPpWTDXQXXUm6VBrE0jdI9E2SqtH/J3NmXesyxgRCKojycfsSaYbGGwowj4/0jKkmxlEd
Mt86j/HmLQoFddFk6LBfjYaUD5JAbw3LCqMZ+kzv9uLNaGjPr6XjQi9f9PhHKq3ejPQ+r1XlLzyp
4/qq6UWmuD7BvwNzykAwOTfLHJiqXQOQKlCSM2o08+upRmzVQJ6e6CKrvXZMnNVQBsjed5Ldc1+0
0ElnuEqvXpO8SyaGcvDhHG3Wf7ccUem3cQu8ea+1nJMnU94efz7DTjYIOy+iU29VDL9hgRVKPVjg
/JDR0bO//YEazZ+F5ytKDejL4vSunPeryoR5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
IraYeYVMFV4GyOOIT6vfEEzfe5Z1+FAcQ2VjQgXWD3z4wSiLhzcOWZWT/Sog/nWLXgPxlpaTkGOz
XHJuwrlCjGR6U5lDSKmMoHfrR30ne1z152ACztdXKM6yIDyJnHTIWeheRPYepgTGODdnozE6wZoj
sRrpEkTbz5KOMY81z/yYY/IuTxF4zyDexv3jmq1XxuUc2u9THO0HV+vnc3syVFeuay/poW+Cdb17
bCqOu/oFBMDUmXNNZgFPg40php3bnH35UxsSuJyGE4gtYZWQXoFaJww6alh9gCv3kif/EjC5VWoM
lkxa4uic/feUZ/TuELWCAKvvZnVhi/jZq1cpIhzLSwzzK/As0MQ29gSTa+a2GQ4J2Xu4q0o8gWx4
NWNmlCOhVfMNi9NDS7RyLWFhv9YsZBckbq4CW3mYbi3XWav0eGgH6PmJ8BPcvfmG3SGnBfNvqHk4
lBgyEdlNw8aMSVB/4T3m9ATPgbFQPRMc4AZ3/roDjwKUdQycfS1I05prGfOPGF5oGYOPiyhkwDww
YWUdq4qqw2DQJhwp3D8QoY9LMsTapzErB5f61kIp/MmAtGIlPciJ4gj3CQKfh6ihD5qjk3ydPR6p
l5GBmTwsBHNIq5V/z2TImpayosSDMvY142cWxes1mXg0crNbl1PidTxkt2GJrEFtqpwlTO7bRAk7
Y9MoeWb16sCEsxXqP+FsYBiNHjAlLhpnu0+9tmv+aQqlwa4EvxZbUwJUoh6DQy4F4kr0b9yBlWkb
Keppz4k4VCAnyKt/oYObKW+2JVLsmLwxzItWoPdOwyWcJtZwMlm5J+ZukhewmIUdMx6M3j4Y7K64
P+8jrh6bC/oS++OcE2XUz2c2l/wlR8VsrH7UCQr0ZxNzhZqJbj+dBnh4PTXy3dDWljdVo11l23tG
CSBoXRcT3z3zSD6drZcISxhbtt/lz/Jxd4nnd2wG4p8cBdNqzvlisoqxnlxvPbPaCHDPWzjAtPYo
zy+REHtHOjKg3M0Q23upK4Fcr8xH9Y2nG8unFGNHEVkluGeaOm0hUtDoww0o4zxaKJxFI9SLQ+V1
kuUNVQZ/2s9f47QFI6nku79CBlVSzywENzxriHvrYYSIcZgLQv+bW9wenljSmXTiw1lkpin664Wc
gWp8YCF/+kL7RgsR6RZlFyxx9QBMrcndCXXNUd5eaPC9cyH+D4ZKdFfif4BkoEOUyd9Orsk9OYR0
Uk3HtFd3c34695Ix29aov/Hc1/PIDsFwqaaEkYvC6E3m1At85B4HY2yRL6+Z95P+K+fpnjv9DQWH
jjfhUcA8XXia8Y4+c+AHUJyD6TFCVeEXUh3WgOEk2/g0+n65kO3L74krm+XkxwLyEIdh6LCvRbR7
LF0lG1Eu6qfPDcW6amgnTYSfMdSQQZlWZbdo6ufDlIIQo5st2uRZo/1P/U0+8Xm4kWo64hm3Jd+O
8khhPIaph4BfVm4tA1vlZL5li4Oc2U8b/F7JSTXZJ0QzyTRDoUIJjiWRHmXajbWEpjZUHXumxPTu
n69mvFMp//IkMlOpmtJsI7Ugjc0UMMCZJ/0aZ7JigxYC9gB0tpJy10VZzHy54UOU8hG6Mo60nKOj
ciBzDcugZ5oEoa63yoAHVBFNnqs9AZdUyBpF0wNg80mZ8gv+tLrQkw/d+1BWj9VEjLEeo5/ng02u
RW6cjCPl++G0aAjdocjB+Q7uBLbk2NF2p7hK/ixkJiyrjGm9ryxvRpFy5kTuhfx8FmGR/D4ghRTq
DGpqtSNFPbOi0vkkvfeNNY9ebxt2lNOji1euqSmUyet2q4+KwT4kb3Pb08sdsUYRkssXliRj7o2b
B0zorw1iY3zmVGtSlcvSBBhqL8X5xmLmdVkpZ3zvsuZcAbmyG3zl6TuXKmrOFoCmwWzFMP0njzyN
hsXZ86ToTUW4y4ofYz98pSMy/jW9yB8eM+Z8wwv6KcBGUJtnSoQ5c5LJce2QqcympOq5lkTyNdO9
4VI/ipIAelSYT23u76SNggaZJRpq50dI2IeLJ/YWuZ5ylMSk1X2qZNq7rGe6Ddsq5qdh1PXK7WqJ
I2ot4ct8cWHrSqbVuCVGcTVNVVzKCtwKSKjJG0tdaqF7vzLPKKxegr1JKILv8dXYgCO+hkrGH5UB
EC+8Snl5NyJZN57gKKuCYkUeLkGKYFpML5EAErKShy1Zvik93j4o2saXzKmBbcoyq/QB1HpLn7Kp
rlsv87WNjxP3y1D7F5hF4p9fxuf/0i0G+1/c0+cyIAkyVwHsOEeGHKkJSra8bOk2wpcxl665ZtdN
J0L8jn+0qpTpqfZtVxkGeWt1k2SozXS4xoKdyITZ3tT1aHGx9+hrwATyVQsF5x4tVufhXbRgqBkh
Y7Z71in1q6ixkAesz0gfMBXGbflgwmXFnokTYcZqjS41xZoa6sl6lqZFWrljUaCQv3Xoxk3fIpcB
PDpSy1jQ5jCHrezVw5FQ1lHT4C+F0ACaNUfp9O/mb5qGLKtv4YKY0nyV3/3r3bszKSzJbLuLlQJn
G4AiZhJkCGzU/LUcprnqn/jKV0VeYYLz8j+bhu7X9zABzKM+O5d01J5WYVhRIb6v1g8k7fmx2ccf
RKmadoIp5fE8J4TRVb51/bwviL7O5NXPkFXowfbg9pGuXIWe5AEgJtZKsm+QPMWlvYqmxE4fEqPY
WgatEHftUFzRk633SBpnoBZRsf5lQpZ4sLTYk8qlGy7LgsSWaaq9Jug5IgfgivJRliEfWkdUv96w
/BzxwGb1FtAVRBT+QNwSb1X23MZtjmYMrR0E2XMHyMjhq2NmceqG0X6Vam+GoXzuDhugWMp3O6J8
MUnVXIuv0OrBV5Fl8OHaI3Zj/PLCMv6/85hvxnnjhObbtTXTMGhmOrVaxhEwQ8jG8d5FNU0OGfgw
ct7QPkPWbp+vtIOEePE8oTa1U+L/gNNKpC6bSyrW42J+1UNZXzXAbscsJw20noUIsqZuQIkbSOw8
GZabi/vc2IWbspZ3pJL/v9I9YVN1A76pOABGwRYZyjpSCbA8qwRC32rFFtHY7NGxiYmPz9yWqrcc
82dOcmrcp+gHKAw5OU4ub86xIhuItJxROFHGUhRdkHLKMiJmlqM0gujnscseIx8sNc5KYSw1IYNP
G6lfm4150NWnGyQjQjx3c9scj1aSDipQmFHXCR/VNpef7vjEkTAvPNyDOR/2UqQPBQW/r8+vehBT
cfM964oLQCn+j35d9EmzcZdluWeuwisy5WsgxhDC69nXDDpNBEDJwE1aF6TB9DLmme55e4N8LpvJ
IkAYGXCAUABMqCMbZbiWSxNs6u8rtmpobPCtv+ebEgCOGZC+9n/f9QmlOlDhtmysCg8KfvHKVyHj
njvUdxnRCSTSTz1MZWh9V3NN0NLd8UOfz9quscMxJIB+FgInOPtbhGTZuYoCt8T0jejx08wBm8/b
2tBD1E8GtdSHATJn7Rx5V5uq0D+H/Xy6q0rjI4Gsxzje2Fs59H8fUgT4BtAKX4ipASeLUvbHibJr
JeR/dUv/mNOuxV+ZI+DeT45nQAKwYeZnXvUN9vmuuI6S/Q1qlXWT/hF0WazOlT0yFGrM43NEE2RJ
Sxq1Mbm7EJevXi4Nmox5abnsD4Kt34u/tlsjuqbMzwzdi3c1YMfgA0oodl0hrK3DG45iqYc5necm
tVPdfKf1GIuOYFulJPbmGw9W2MryIarrx42W5fOUHZ3ZJZCOSqSn2xz3rPgjEXGqod7uMUBOXUz1
gTcb1C0rdlrT/ZUGdR1RtnoVVPuvxHSnZYyP2IGQM33IZr13R9WhWZOHe1FiFsDidPzcgH5eP5Ah
smlp5CgU4deARyvaOZLemO9t+iSP42xQeO3c+JMkwliDTiWeq+fZszps0RYsGeyM0vQWiUmkT7kL
0g7Zt3TCnrT9Kchcjv7WBPoNgTLp3vnLnNDD8Y+17PqeT0rGZxJ8ruvVGkJhdVWVEWJgLhG0v0pm
bLIVFYwTHHpgxAVDUkblpU5Dy0GxIXhr/Oxr7DVZeTJK54fmCtCAsAo94WyIwkHwrYKIOpOHqqxp
Wt+1PSWxjRZd7kGXr8OfUiDbVgsdKsOdyuM6v6PMrpAgbAIKcXtiFzRPzgQB22J0vHTiSE1SIrgz
U0gRXFDLfgHJdA/MGPeHioMVtcBCqjWiRWOCzcy84/Q7P+e+SwJdFYZDfHCrglr6P44ks7mmjLFP
hofHY82w6m2c2J4G1IhJ01UL0+9qtAR49EMRgTEmj9duWbck73RySbLK0nmhNcibyWX61SO9xO0l
ErAn80FUykW9kOxluoDR6Walj68dikBXjkXDEqpAVNz05poWP7WSXa8zL4n4OY4RKakMRQu9DGUj
iNJAFtp7J6juuMEwq6SVk/pqukxhoZdwk+yg7E+UU1sGTmJuNGCELIios4XTIzo561RjFEt6zqDr
dvTfykKdM2bzDIzeBE9nKE15dUHF4EdDRMmVUGFRJEnAuWt/idwrJeiE7Tps9JIZKvkwyGmDjvJ8
fL6pO0d6MwJCBvwPbGt2Qx35G0INUa4QJGsJ+K+ZK5oWw41Krh4eGGCCnbyFz3EaHHgiyMMbppzE
4K7LiJugii+n5KcHaLqG6ONQ6ryFOUe6YeKBOoYWKO9V1wmlOp/7Yni6uI+YacZ8118X6gRO/ceT
Hnui5OlHc0di0H9uyXZMyKmVI0faCOHyd26RLUwHKVPVqq7Th6Ohy35mmrox6t+h6zy+BJVFchiE
D0P4ADMFuy8vjPOIdNOJ0Lh/wCJOidelSn8Jyp5vNcbJFqS+CT1otDk5XOwevHrwmWztSfoV2fEt
sXdTtTIGQjbF/MvEPo0hsjxpUzEZGqMBw5hkWnGOG/wkQnEmZsWOL9WebLuKgPk4yjTJxN/LBt7u
zAC5hB74tDPGeW+XX1fuRxr1Rh7EDT4rXF04CPtUOyWq36jcyG0ziAV0GSl98gnZRvZwj8r7BXLf
vW0vfWbLinf7Lp5QGXQh1rasIMHqiu+IQMJgb24f9ox4rZ+ARYr1pVmKZCzIvKB/PwaALI4b5CwS
MUP44IVba51heC3Q3KNoBrTso8X0MnFdp+FIxiZArBwHCaSzJFUloxyC/t8ELPl6z6DIIzfgE2JX
gOfyNGpAtz9lKp8c9XOtfJeu+WFVj2PJ+YtZB0aaYMSkFoHmSSEj1sYDJDUT68hkiZlqxog9jVot
legPTszMGUys/05R+Y/gu58pH89WghumCVViTioqThYfT9SoG1RrwfjBZ9ZUsRTzqnCzIrCmJ9wt
9gmKA7naciqAY9a2VLql6FyTt5orC+Nt6tc9bJl3Rycl8M312Tsk9mh08YAYqCAklC7LKFerM/Gb
xrTRfz5Pnp0YzYyeT9/n8diSqV7JRO0yasgJLXBoKcBkZluNCBRo5EX/qZPd8On49XktnBMySZaD
neF+9Tfcs07qVg7gYQWkQmWg+fp2sBC43g5hmsGEMDSACZSnL/Klhcea1WWzX8Y7qTtOt3PGlcUt
vGZ2maO0C0mAoKX2jh+d3cggYQ2fWmnxjSGyiDi1io0AEXhnxyN6bvEnDdy+Q0HbaiST0UHGwzPi
+vfBq25zRNPdRGsvzZ2TSOeI6ZkZPw9ukwgal4gufuWtJECMrL5qpW21seOOJ1d2IpuZqlnaBCkR
4bQTzvGk7EkAL82eXtHl0rOCdKcjWIM+cXmrZKxOWwk9v3Zo42VIuIcrZ4R9Aub+/eA9NU3DF+5L
Vwp5yiUAXk1DANlTPkbu6agbxGPk7tPGbGtLcRusyfDvYccC5YdrXhsVklheUlzs+RdnONxO+awR
GEPOrcE/3rLBKmH1pq6FU2REwq0T5zLVaUoBqzQ+wwgDwXYCiPns/RygOiiNZ7Ou2ftBi1X4TF8B
otbDUMHMTn74sLGWxd1Lv32zLXD9Q4HlExklygj7CzDg8TEFSCUc3KPM2wVWNqIfrMJ/IJlhUSv/
53bE4CvaLeLt90noV931gtTUQqPvNvokWx1p1eXaHa0lbzYyekEIn47cAMnG0a50cyxsAAgMDx1h
bJAhtZMIUuDfAfBdemUtdy4PC5kBoWZo4ovIyPn/LtyHjC0ocytMGo+xYQgXzXhcrlXW1M7QEfOm
v2SIVAZPVnVjJYQzsjPagFeV9EXl3rDrRe1HTg4hxLvR4R+1/uzhfzitKm36cIWVW6raEraCP56t
ICGQy0Gc5tDKA9oSN4fDbO0vG6etA3oXpWvhi4RYQI01ZD3wisTmRml9/4Wdp6dGPR6km2w74bM+
K0Z4iG0tB5g52JCeXb7iW691/mfEuw8tUNkA35K6CR5yOr8VSc6cPMjlYturKgSyS6rd/LdXN8hw
d6m2BdFdJfex49n0fx95ffEDqhP4huGhjEmrgdoxeDBghY0RUuUWwpyhSkLCNVjBvyeGi3Tug+vI
VAEnfhM2TLweUNbDLopDOnsToVuIP8etZl2cULLfsUQzaW3wgbbKA6U1TeZFlmhaTfvb6OXXSzHY
L+6Nh9F24xdkYFpFgbSYaokI7H3OZpLLPtMUTZ0Jk44nXjmx1kpRwXy4CDE0cE7/vQD96tZyd1a0
nCB5hBOmcphUduOKKM+mdIYRgd/GNtJ8SQGixUmeOHApwZdo9yKiJ2PJ1wAV2EUoxQJjlBhtuqQh
wBqAwyG55PQ3EkBAoBmhw5W8wV6mHqY/PotsE9uvkcG3kQEfnVIMbGhQdF3UguPlXrHxxx+PB6C6
I71+PC7GK/4ggO82y+CzGMhu/vcF5dtgWhEzxzowVn/9WJ8ZPFSGLngYqwOQKu47MIMMVApcsMOK
kEtfY3sDSlhbEtvMj8wtvwl33fvia5qLyMfL/qKAUwopVrDhDPEiDg/Nf2cbLS7DhAoWL4SWPmHN
ivE90Ps1dTezPMXAhQfp1YuskkEAOUsX98oHS7nwsoGtGRH4QC6Q18EfwZUXxcMculcCH8Vah0N9
I/hYnyB1aQl6tAre8XUbMUQVo593QDKV2fg78wTolY3tcjl1A4bPpnuB0AYpY1B7gpETCcJh8H6B
7Wa/mkZfssDw7LctqPe8ZVt3aUgW0zcTCd8Jb4OXswPcIR7TweZHb5CyKnfe45TYzhczmvkdwWOt
+Tf99vBjgX3TkWM2uYCyigAOL0bmz1HtSUcZvMKojSJoF1eA2a9JR1PpgDEZEpvXJI7IB0+bLmGv
8RJqBWBbjm6Uu2IhqsgtFW4O0/gPqoFHTrcU4vzkAJai0IVHpNmQ1YS3Uvfvd1ZqwVgaAul31wt8
6ACU4c7GQTQ5lOknzAhCredNQkVkOk1VhFcQBdmAvZz3m8vZeBFhTAdh6iRp/YHYC1jEABfcF4Ob
RVf7on6tUsnqe/heVxR2r/pNjmEEM4cbxyZlBAbJvFytFQm/TEQgruYQess84AKYHIPNJQzMd/cq
8wFWdvFj3N5Acfx1xWyCzn51B7mq7vED05WlESmNaxTm8uC0snbfIbJFWo9V4m2z8TOBQgbtanY7
7lIY5x5EcKMcFnt1cX3lw0xLI4wexN2OmJwnI78ARCLwUMFeBbfBIjGlOCTqIA87hX79q4xdSRv2
Od6X2ttHhv/x3RiNGnqABlvsgmy8WI7a5DiRVAhXiU2NA/qkGzozxPX/nKdZGwZ/hDTd67jqSdQ8
97CVXLczdJaiWXIDXRVeY3RicqpgOZTjG0T4rJ6mhVL7zdmww7/nE+H3MfRfngAONC5S6hQApZhx
/TmXUYUdv/KyWj3z+VAzPTHoRdPPB94VOZy0fpj40yRwAlr94ChSUqmtL1f9Vsi0BAqeiTx4oicG
yA1O1N5www9D0rTXNjbnuAoH9PoG3iOUam2DL5PRP6NFakZmyLGp5ud4lLd+U6379NzxdS+8UnkQ
FvURowjulEGdOCacvrM0bOuX5F4rqBXSiYe6TGLBM2jlLWfYzILtePKcAYvCSkFuGcsAONfO18wM
TG4iHKBINXE4AGw+yzVh7wnJuQ24d3PGfdzxes0VNriWpl3b26aFT1SvHLzYJoOQbF5CDmGr9jap
2ywEBzVi6dl9t3DbVtqqjR3gv2Up4qUlrxQp9w84M4Jdgpcbj6G6dpNgilKpxwvwc0twJR/v4csg
G6Gu58uWQpONEL/1soXjIY159iYRcURV9rUfWIDehvP5JHedZjZ+oEnTnnX4GSLNx0NB3FjV+NRK
2vyaRCDY5+NS6ZS2NSWY0vi36mP3tSeNnW/7LT0ct1nDdWufS5bgTe1LzX8YoA5K45Cp4zZK6bl6
zDZ7q8wD3wbTdeiz62RxByzk04U9iQ/TRT5kP/HLcMI+SELlBbYEFyG0LjCg1MCpFypM6X8cEyka
KYJQq+hICfFK822iasg340cu1K2bgUHZRXpMEMT5tUDn8urNhFsApBcKkZDS34xdvExq6GdC6D3O
P2rBdaXyxq8MkpsgPxMgqMRMDl6V7nrM1O7zVQC/gzjOMnm/etYJ07eb3RRy5B9N34RGy6+ZNMju
89fuo8U4MfGmXiFlBdqP8J6xYL9NUCjYU7Nfb5uXZcTgr4FalnZrt/3Pnwt4bdoTmNsYAhwTaZuv
BPUHMVNShmchZI/5uMK0z+0w7AhK7UbeVlhzEjI5fmnVfgGR7AM2jZa4yINkai9Q3c+dSAVy5w5P
1qXpv9vghcWk4j+SqAzQUUq0S71xlDIl+Nbw8JxaOHYGQbsIbrchbH38YTTKfybxzt5joq7piuKe
1fGF7/zCEEbqLBD2BGPNwR5nbSXLBb+Byz7WsmUOFyEXoKz6SXfutRW2lJs8IhLq2HeRSTXFEVbp
Ookanp2qOUxSjWD8DzckcY/X2hBvZJEQnhI0FwSasCZpXg3MvRTOfDWWakdx5CYHjGFBAh1aEJYG
GbMFplNPKIrTAABLE3cv+aR195Lt2nMPJdCnLlqE2yYoSnEdDu3A6T/MP7l96NemAaJWkZj2CVR2
pDyvYBTmmmURMBhQ+a6vcHuDwEyDoS9ENchTQkZ0vmw80gDDZlJBL4yZZld0oMocp/BJBxUEVP+n
/C/36xgNwtd1QRPX3ETPh6z+tXrYn5Rgxm8svVBG5V08FlfJHRh7O4vsMKu5BE8ZLmf3uWLy5gty
BDuy/p7pt8uAc/kgwzqNwwL6Poypf5M/VLWr6RJvQ9I+rLuboyHfts7FOWljvW7BEZfskiQQpsTj
1Q8gtO0YDrsjCFPjrxoyHhlZw/WKb586cmnBwmHRNmjl1rUIYRjT7ir31ibdickiN8jBqy79ESk8
4c5d2fL5T3Oy5HqVgdeT2eq1OTzr6wKtVKUU7cyAPx310QT44tdiLa6JGgQ+QbOsj1Ese7XfUTBS
Zg+T5U3ejek+JYqojBAGovgun/bgcLYVPjBrIJ+wGzNamYw/s89zOszMA/lhzb1IWzPMSJRwnQYn
OQEjiFB9YYWt8kVTytZn0JqniuIsBJZbKqklpmAC8DP17Pv75oXT1xU+jEwChHQfN3zsyXG6GR5q
mUkhJxXimiGLK2iZpiZ38Kk3SfPB3gr8dNdfdJJzm0FofVD/6K+Z/3oSUXdA8+9rGGRRhwfE8O+s
xJzTI5lQyyPI2AzErzQ9U+exjgdbb9GfVZKT1QJdgrOPk/EdOZgC2t0RnI6ohRgKQh8qPyoUyAuP
kk9EoNVU6SHMW9d8/T5zAtNNZ9X3UgZ9JF6t+DxbuUX9VIiZSvYIvL9IWjMlBFYsfyrjNSukzHEx
fiuyAFxP5xpvkimAck4oVzz/hndyvE/+aoife9E7FaAAjDO+6mgeH0h8jwHXGGRV16fuI6LnO/Kv
f4pkHc8KpvCDGgVFYgkbi2hbi09J8FnEZG/uufYq9YXVsknBYG48vdODaJ0V0mY+lGS3/7DTU24M
V6mOyaLQnWH2YbwEq4jWzkfUtL9xZjOSETuq1z0sKIes+JXlLgrBtt6gbvHl3okEuCa/uTM4bujN
3Q9WZ8no/uCWrvR/FDpHTt2UdjTgQqo55MEFk2y8SGQng+QR51TrIefxEnhGPGaAJhCalV+tMhIv
pFqfNeJPNE3srtGbrEcCMbbKBA5y16LxlpoksC+SN9atIkUO42Gq1L8TJV0Ka2QCye0tf75qnZD3
wPIyeQgJPHa31JvKfMqd7+r47ZED3Z4S4LV12cHaT3oeFq0p8FsLnRkMp6WfWUWUpHHHNDLrgOth
K1D6oTZn5INhFf9ufn5k9jxxgOsoGLl4gs5LheRwIcIzpL2pfKgJu2QSXv71/E2uAN6LbV7aMDiT
nwEO0o1VcxEjZbyUpmQpUwa1imY78HxEXY4OG1BRoJ5DMuNc0hwzzP19Sk3NKKNs6yK+8Va8CZze
pnXSSHFnvtUe4TfXUOlkwCKXJFCzw0C449YB/AjnIfxAWyG/GlQQ/RaWl5xU3kkJCmQEabu/WT//
W3lGPqA3+a678CH3Rv3ifdptVMkUiPhazS7ZhAObvoERmwzKLbdhMTseypp6Nb8/CG32KkyMMlLh
blx9wlHp18EVt+NVb21c3g3yD3qQ7Ym09SWm/KkYVL/rhINfI+f7QOz9EOBCfviJOMZE7r49q7Jn
GsmZnBf8jQqfsBOSJwmFTfjGvYeBzozOKa9/pM1NqQenRZZh3A7nbAOcuiXCWlGSoxijP2EmavEY
XMH1A5LcEWDJ+gteacG+edwM9SccpWGf07yX4UK+HPoIUpG8UJHDJR5FpGAijbIWT6J1ifhXJo/E
3rJHEJdi0u9e2xvOVkvmymPcvJg1JhjGUBAfWHZAAfdJFD33HpBsm0NMrnQSj12Dz1ABafaa2XQH
Csai04DqlTxI4KpgPtBWtmwuLouEQ3scQf3c/F8tf/1A3oz+hTsObVZHxazhVJAj3jtUxppP8Xsy
HNX76nHp8PcBsJOWVUMYectemLaV8TliuDp4vw2EAj9xCdGjCAJ1Xm5QOzgBRnfr3DtKwtlCUaPJ
HOE4u+ljQP9Joqay2dd/u2V8bS3SZpkDzbgrMuYjT9S9RmhtRVafXD1UUo8z3eNn+ry8etDqt/jI
FHkZeqWxdtshrLseyq4EwKWd+ebZNiINtklo/7dnKXyyaWE/KPp6nRv/BGDHOBD2fdQ3r6hCD6/l
aOVRehw2MTRuFk734YoyPZbc5evt2fiK2D5yEBFlQ0vHYK4UUKlwPCEnmtZk5hHIwvORo5OWacpV
pIcj/+3hjmxrNlH2omMQ7ZDUnzYKlDP3Btea93skMw3wWTfjARuOEDaxEA1MsBnOYTDkyTnpXC06
uCHyu08zmp51U4w7uxAvCF2RpHtz
`protect end_protected
