XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���SP��;5j�x�9��r�k�N4��%���_���U���&X�R$J
��}�.��r���&�P����e��|ͨ�궆�T�3-%���:�T�	���ށ��xJZ�Ag��񍫵,ow"���Q��ۼQM֖z��?�C��'�+�o�Z��C�ր8����� M�{�4���9,3�)9<�����,��]K�h�Z�Vn�C�^Qdw#�h� 	��`>�^�O�oŸi�)��*��.M��:�q��0�Օx��k&��'b9��ܞ��;�kP\r?0�9�N��.cR����Կ�9�!�}���=t�ޟd4.G�~�!ȉum�SLqv0�EU�P|�e����k�	���6��Cn�T��B�hZ`ZD�m�
��.f�c��p�\�{�}D�@��w�3��:6��S�IM��*���׆��8��:.�*\'p�qvs֝�Y����#��C�뇝7�����D�Y.My�	^8��N`]ޱT�.���#P�~m�A����1da�x�0��{,��h���R��Pp�}O4�h��h��B�A��ݪοy�|Ƕ (\cߴ�q��{�њxi9����MX���n4Y��Đ�{�Gw��[2a����oTz��w�(��?K߻����h#�N��.R3�c6I�=�&�_.����-7	�7�;c 5ӞC�Y'�@����ӗ���|�}���P	*t��y���l2K1AJ�$�cm3p+�S�r��)��aKK�|����ˡ�7�XlxVHYEB     400     1d0�����&mJ�Ǣ���|7����p��ƚ���H��c�P�����X%�r��)��VC�0r2�'�~AA�*�bz����hx�����!|����
T"G��:�}^ڟ
�s.���q٬?����¡E�ǣ��ؔ�����!#��*t���@L\ŝ�D�W�"i��w�/�_�e����K��꾒����<d	�td�7�B��8�?�UM�P����
�A*����CP��j ��v�|�i�GG6�G?5��3`N����0���'������8�4K�0�Wv8���>J�#��[�;�����,j�@8
��\kP�i1��{ЈJ���Dr)Ư�����G��߇؀P1*n��-�s�8c�ðnw��("�X/��������z�W�O<I�Y)�`��E�����57�y	�,{�>l���^�|� 	q�%U�Ӧj/���g�l!�=39Q3����XlxVHYEB     400     110ؖe�E���kx�����N����"�F���;Z�wa��Z� q��[�D��.�dv�Y;���u��,��*1&Jμ
���K���+��ae�PoރF�~���aw����r���L���cC]�qC��7ua��,���[��%0�k�:jN����w���B�Y�A#�,/�d�&i��23��~^��|���s��٥8L�����}YH�ζ�#�;%
c���sȔ/f��t�-@&��m:l2n8���m��OA���T�W���V�;VP�XlxVHYEB     400      f0;����S1ӷ�u�X��=FV�|���~�qR>�ȵ�}!����C�-A��*�-�	�}b����#.Vˢ�Z�-$U��������쇁��ʘ ��i&�L��R�*�U���w�?����j��O��BB���a�n��8egP�����Z���m|E�'Sz�(Ncυ_�Y���^�S�5Z�@�Q[/��h=a�K(���"?�"v�yfT�Д�w�N�n�\ϫ�8���w������� ۖXlxVHYEB     400      b0�&�R�J��c�|Qz��f2V�����NP�t�Tq�?r��(]�I�mw��Iv;�y�kӫ�fo��dC������0�F�&kw���U;����?(<��?�h��4ikl�+HNDV,��Q��h��pn^�1�f�,d�[��� �?�xh:�':�sS;��w�ҽ�E�C�XlxVHYEB     400      d08�	�����n��Q�l�����eߥ�C��E��4����r���oZ�{���MM�?�����GO}��̛y1ӆ�!Ko���έڶK��+p(�ay��'�|�[�ra���� ��v$|XA;!�٪Ī0�?���?2_t�/���P���0��5^Y���(�V����e�XW2��Oŷ�*MӦWz�֯��`��x��fXlxVHYEB     400      d0���m������$���Qى*�Y���Q�cT��9r���̄�10�YP�#��1�p��EgGC����MPբ���л~R��t���VAT%�_\h�Z�7QvXL���Ql���g�r��I1���+Ia��S������>N��W�e�TOްN�w��C�Rĥ�0��0/���n��4���� ���I�Ih�B�гXlxVHYEB     400     120�N�8S�V>-*�)0�Y�E���Ծ{� ~Z���|�ˁG�:Cۀ#���gjrbE�}���e5=_:����і��ZuFޝ;�G��rf�F\��GJmR�3���3�'1�zb�rS�\eGD�=JP�����O�\��2J��g+O�ƭKdC+��[_ćS>��F�=A�� ul�Z��a:QI�.�t�R(��9Ȃd��L�*��9�7`��(��xO��];���>���VfU�L;�T<X]� c*�s��F#�u2���{� X�Ԣm� ��;�ƞI��M�XlxVHYEB     400      b0�{'��$�I�p��]����&��o���*~��U0��fP�{�7D�Xz]Nu��-�ǭp�i�*��:i�H.KK��P/��9CgF ]��VT�3�����r�~�k�'N�i�Psz��I;���=�A�0�?�Y2O|ǆ�k�,��_\�/�\���8Q�\(�S�vpXlxVHYEB     400      a0;Q~��8M�q��������!��=<��_�e{�Z�uaL��
($��(Ȏ$z �ݍ�%�
t���Վ5���G��Y!>��1>�xjT "�7�H�a^�ۍ0$ko2ԓ�r��Ϗ��(@7�y�<�}Wjla5�E*��kԶ��˥��SȄ�XlxVHYEB     400      d0�<�4����)�2$&��'K��^�z�w�����eٮN�O܆�w%O����p�tL{�<���[�f����C"�e��TOR�������tē.:,���/�Rҷ�V5���ݗ�T�?���W�O���2���Fh�1(��D��}�����"kgh�Z,S#�C���W>�����p`��c���	�Mx.��XlxVHYEB     400     180ƒ��̌�q�W�sؿG���:�j��-���,t�l`��qo7~VKc�8��ت_o u�E jsC\�����/�+�2S
�j�< �i=�?@o�x�'3M�߱��p����'�k���y�]��0���w�H�� Z/��o�'5\<���J���g-.W#�ޠ�ԩ�	�XN��"�D�T�����ovE3�@�=n��L�Tjo�V5��=8,�If�Y�#Kzm/e��]��s|��ph x�/�8�iP	ڗ��$�NOP��-Wgو.��6n���.���O�%j)/�Qt+-FP;�L
��ld�I=3�!sqn�GR���6K�,ڌ�Uԭ򌗻_�1��%j��8�L�L�P�z8�x����8G�s��z
F��s�XlxVHYEB     400     130vfy���oX�=����e6���^x*F���hAi��ʙ(��G*��R�Q��L�+M�U������M �Q�#.H�s��]l �!��U����Hb-��M��4s[�a��ں�EHK%lm�E�,	c���^�����M�����O��."P�q��F�R��- \t�p�ø��i�x a��G*�}���;�&����m[�e ���[r�ݒ n{��θ� ����Y��*F=�W�+��_6���˿�O���D��ܠ������:�)°>X~O?rFv�2AwYh#MӏF��B����t4HXlxVHYEB     400     110��y7�hE���lG`*!�
�[=�����������+�S����Q|�_�"��w���K�p�o?��B��o���ORK�Buw�$��w*�G�-��~�L_��
/�=}\����^gc<F��0P��0h��AX��~����G^+	׈+=Fu�x%�!�`�C~�	�0�j��M��l���{�]��J�e*�u�Q.��n�U��h0N���&<�o�EF3�����K�H��`wՀ�H�fkYC�ѿ�P�	Ͷ��U'���+!����:�XlxVHYEB     400     190$���'�|�8k8���`'U*$>4�gB���X��T��V��(a�1���j ��_��ăL�C+|l`̗I���4ЍhU�r~�^��V��T�]D �Nl9׌��մ����1��U7��T��G��%c\�Zڸbv,��}�\��	u�	-vT��a$����{�C2�ɔ}SZ���q�ɢ���D�!�ቈ�ۙ�I��w,)ճ<��a�8��{4;������I��j�8����͞��t�Gx�dP�����
\��|h7YV��_���ʸW����׀� �o����r��6Q�{�k�TxԵ]�E�ߣ���\e�xB$���A~�]� �Q��>��-k�"������!��'�T)X�`�ڗ1q_z��m�U��_�̭��o���rum:�t
XlxVHYEB     400     110oxo�Gi�)�!���vdBU�^].~�lB�Ѐ�.�w�'ǵ�F��ƫY��u���B}]F%���[�s��JN��xm�t;�Q�~ވK{f�I��N׳N�{v�����ӓt�Ӂ��Nl�R���co�zz<Cr�y��KWY��� AU�+�nQ�~�wd�ї���Q�2�"`l}��ٲA�Zq�c� �nR�|踅9�@�h(M�˲h6��0�NU(;���Na��1j&�)H�)+�'5�VC.�"�ꁙY�GM�XlxVHYEB     400     110�q�j����^R^Q������	��LMO� ���'�f�}/�tͷ��y4��ogO�fԂ��60�j2i�2=%��L�LD�Y�ƣ��b^L䁧�=T����ŭG��W����2izeJ��0�+���Ö��y���`Rg5��~
���"���͟�U�uw ��6μ�M�;����������'��� �g��FR�0�Wgt{dX��'��@.��#)��D�Z\��� ;��T��lPKK���r{}��bXlxVHYEB     400     110u�r�u��Ӿ�g�?�9<M��V�����:�M�	M��	]j/�O��E*��C��t.��� F�H֣n?B���_�wp[���!��ܱ$1�����W����Jy���P"q��6���FfG���N?
g�W]YY�UQ7����,@إ\p�l����l�%��0��ٜ,�8ߠ@n�+*6'�qE��uM�4� 3��}�XuiY�I��;����D5�^R_k8�JW
2�j�)Hs����u��mP����4=e)HG"D�����XlxVHYEB     400     100� w���' η�n���Q�:N�h�t�U��e�˨'�g�l���ά(ӊ��/nI����i���5A)NW2�&`�h��s��I(�r5�͘�X�|�o@�50v�h}&?�J��bUΙ�H^�nX��n��հ�Š�B�Ьh]t�E&����Wq����ݥ�P���������<�d}��������|�g�V�!�~ޡ�Kx�8GM4[��UE�[#̸�RA�p�X.tgyޕ��#����7���Ń[U�4��(�RXlxVHYEB     400      d05�-Ht5�4+�:*UE��k9]�E%s�{#�{��ؕT彚��!)c:#�<��5/�U��|�{� �����M��=����d��.���FN���\/��a�́���Ѹɩ��wk�o�P4�;=�|��"X�O�,�!D�c^�$տ��-/aN�^e�JY�S��+PF�S,-`j4�\#�*� �qG�<��2C�2XlxVHYEB     400      d0�q�g��rl��J�51D!檛�B\q�·�����Q�[�����WT9�j+$��x��C�JFFڼ�O�!x ��L&�߱]b�7�'�7����o|�ī�=��H&�^{�N�<�;}Egp`S�R�u�Qgÿ/��4/z?��*�_��R򦄎N@4Ф�56i3͌<9~h���F�a�	�ލ����N��0;5�H�\O�� ��R�XlxVHYEB     400      f0��>�Z}�;�\#�WpH�u��\���[��k��&��l����U�@���w�MQ�HP�,�ΐ��{� c
�8<�P������e�U�ښ6Ь�-� �����r���E���Y�QT�������}}{v2�x<�ۤy�ބ�d��=8������Z���&��YFdы�|�T9� ��OD ��/�;h�P��h��iv���K�����.I�^�#bS=�� ua��`��/ ���X����XlxVHYEB     400     160�WB}�zq!���'�<��t;R�~�]�1ك. ZJ����|�׎�;���o��g�{΃�'��T�d\��&�`���%Ř@8����4���Y�!��,8�A
rgaF/����2�]��x�����#2 8��C�uj�!��鸿�K�B;�;�S�?��r8�R�jO�տ�C�Q�i-���/�Ѳ\C��D��Z/�!���qv)�3H��$�� *%V�j�6vd�տ=�Q
��<�w=S��E^�G�{ H� �����M�����i/�����W�%;�R��W�l`��*0�@���_k�JȺh��||b�6!.��"R�G>�B��QJb�i����XlxVHYEB     400     150���N�$�A�[��".�y%v �6n
��v���rN�K޶��ߘ�N��r��\�z�7n�����ɑz��7&��D���z=DpH���Nu��f]��|�_u��bU�H���W�T���a(�9�ʴ�pN �N
��D��_������:�'X�9�Ą�u{]F��p�`�� >y�9�`/p��ȚS?�0�b��jA�$������[��5���7��@k�`����
A�Ő]n{�Ng�>JA_����&ѻ�҆���5r�VyʥSl�o�=FnMk�jϯ�-%i�Q?%��lm&�|��ﺱ��O�3�Ǉg����QXlxVHYEB     400     100�(	���&w��)RQ�ҕ���c[גx��)� �|5���z \w@4���DC�4^[+�
�$*�e�����}a�r�v�xmd�����A���8�2�0��2�w�\�܀
S�Yx��fDѓ���b�@\�nu�/�R-6����P�O4���GE��E�zй���Bv���ٽ�B�7!�#�(:c@F��5����	�Q����ԍ{�ީ�S12��kg2ƿ��6�+�a�6� ��Qǟ̞G>���XlxVHYEB     400     140HwK��� ҭ��boP7$X%�h�bV�ڸ��d�R�¡�[���L��"H�)��?��ԝX�w˦�����	�K9V����;�G40�Ӫ���w�,��tHRtD;��ߩs���wJ�K��u��A�lV�#��5 �����nc:�8O��U���,"}~,��YL�>�j/���vc�jZ����R�(��`��7�).���O�u�o��eO@���,u��G9|ЇvnE����m����֥��b"̘�����X?�})%RBV�ѩFZn-�Xf`K����.טmd��(I� D�T�X9ӑi$Mf´�XlxVHYEB     400     140yc/p>S��{��aQ|��OO����&��Y�ϗ�j�]u�\��o�M'�mR*�,�m \I�=�hI{�Ov x�:#Bwƃ\�0�E9 )�g5�Ǩ�$��E�B�N�ϴ�a\>�*��e��G§���c��Xj���c��5��3l��l�x�#e#e�N���a����b,�U�Q�8�g�DΪ�Y
/a�x̨$!����tt�_c�x����<q9�b�ߡ����������)��9���>��B�r"/'��C)&�b�unN�ϔA-yI#��n�m`A8��k	 �h�T���q �T䢓%�͊�1C�Ouoߋ�XlxVHYEB     400     130��KP��4�Қֺ:���?4�]
3�e�������"���j�]�Nإ/��=._vE�(\I!����ڂ�V׊�Ɍ�U���,OVNA]�{fgK�L;{T.d��X�&�l뭍�W>��y�K����Z�}DZ���vzh���`�;x��])���f��e��B>����-T�|�4HJt{�	h�d��|ă����uƥ���Z�b9N�~�o< �#!e�'cX�'H�+��D���b�;�L�����T�lb
r��SelXo�ݑ��xxQS@�B��?]1��	G�VUZU�XlxVHYEB     400     120�h9�l������ښ"~����F��Ehѻ����-p�T�J�'���w����0�pC~��CCv�E��WE�/�P��l%ڰ�\/�P �O�o���|�ws%0g`���n\����_��C;6�&�/7�q)�V��X��#2H�٨^��)�Qб�J�o����H2����>rp00�,"�)ઉkh0��B��Zs�S�G>�+�g�P<��N�(��i�(&ϝ/>�����0�^߼�SUb֤oJr����������J����T��E���VWY
�xXlxVHYEB     400      c0�%C=�<���r���բW|��35�/�Ҟ��-bGi��LÐ�@��Y�^�"�ΆL���J�8���|��v}���7�k�\��7��K)��n����Ň}�gR� qE��5
�LҬ**3��B�H�a�6��dG%;���J����Tn�7���X�'��r\��C����E	��˩i�s�i�XlxVHYEB     400     120���""|�
|�5}���O����q��ߢ��̼�����< ǳ��F>&�����d?�T"v�1Y��65g��'bS�n�����U(�DӉ�-��bԍM�;<�ݖ�9�t�Z%��g��Ȟ	ȣ�nKKW��z?�v=���0�g<w��Ynan��1�������f�֡ڠz���,l�rN`��"�d鴏�j�T��!>���k:�>�*I)�������lg�����ea5irG�*���kbݍ��G�$U̙s�Ϸ�Z,XK�c��RS��XlxVHYEB     400     120�����K���ےw��^��ք�!�Q!(T�J�mM��Y{�N�K�b�?!�4�>�7�/�������F);�)�a������=nƟy��;�NZ�|8u<�����G|p������}vDd�~��K s�j팮��V$��`v}Rh�.�vޖ��&y��g��Q��'��-����ԋy��)���߭>pb���A�����H��዗;B�,����ܸ����h�_�Q��9��Н�"m�g�C�ʕ�.��;P ���N�Z����G��$N�D$ӘXlxVHYEB     400      c0�3#���ٰ���uҳF�;�����Ǘ��ȶ�#��c�b�~�|��5��(?tM�B�����]��j�T��"�����Dy�;>Ě���F𿘎4���	��N���eX�8l�ӕ��\�*m�:���J9�X�2H�M/�s0;^T����X�w�{����}���s ��PK�W��r��^�����W��{���XlxVHYEB     400     120��o�N�O�X��8��٤�fu�n�0gd�����Vl�_�R����Ri�`��L#��	fݼѯT[��oOw�,��������)�>���<����LI�K$Va��	Vebp�A�,�g6�@!��-�V�����d˦��H����U���T�w�Ӣ;��-��,��P����&*ܽ��gϿ$:�a���h!zĮQ1x-ԥ5q�*|�9fFs���v�вR��NR�/�����Q�����"�fꗳ�A�i���ͩ�7WGx#ZUs��X����mXlxVHYEB     400      f0���]OZ�l�w*�V��\��	~��ݏYb�O��F&Q��5S]�=�Z��݉�ko���Q����
|W�B~���}Q�[�ٲk�`<9����yɷ�phk�,q� �v��G��0d�o����Y��2K���(_$">����h�1Zf��3"b�v�uL@��HX�A�F}(�Gظ� |��Y�j�������!�w.���<Ca��*�UK	<��E`Ytr�YQy
��s�<�K�XlxVHYEB     400     110Al~g�k���I�sB���Ս�嵿�G��ֺK�!~�e��	V��m`��g�0g�`��Lڐ�H!�\)J��2*
���P�w��#�8� ������4�!�߱����~	0������B{�J�W>�Ѫ ��(�F���,����C��o��l �e�nA�
堦Q��4�.<L�E(ݤ�����E�<µ�mh�JQL��&{^�I2��Rx�G kԮ��R䄱I���tx�}�k�]�|�SN���#4&���'�:�p%�-���`XlxVHYEB     400     120>�t�i(rk�o�JOk)t�b������ਤ��d��h�We��
v��f������8��� n�n�/�?���NKj����1��������n��a�˥%��Ϳp��H�ʊ�6�Y�5@픪];>����P0�ϥ��MC8)�NR}�|��qK�Uޓ�s��sC+LpIX��hh>�h؁ �Z��Bp��'8����P�a�X/VwR�~I���OMY�݇���yɷ��:�*���J��#'���tT.�Hzx�D���{�s�� ǂt�K�E]KC#���XlxVHYEB     400     120�v��~3xUy]J�wE��r���^��ځIY�}H��!Ԯ8�Iqڔ��'܌G�:*�Ye����v�B�ǊW�q&��%R��X����a0�b��L�:7D'��$i��hޞG�Z�8�Ǭ��ᝈO����?��o�G�#uC�L��"K��`�v�<��q *c��C��æ�Vi0*����7N��Ӎ����[g��8�s�J�����8Rm�+�:�ß��	��Dp�4wa	�pq�f�j�Eڤ_1�+8��Hܰ��i`��h�>#XlxVHYEB     400      f0��VzV�����CM�>�dp2�*k8��`5.�^8�m0"��e���RJs�
��&��D�(�0����#yQ&F�=�u`A�y��o*�@|��}�lv���������>�h*��%�{Uc/�d������2T�T�ԜE�t�W6A ���e�����jf"PIB��֫
( ha*��Q0�~keC������{��!�	��TY:b'~�� ?��-��{5D�F#���n3k\XlxVHYEB     400     130��b��
��#��(���L>yL��M�[����q`p��㌡�GG�{��)v����á��U/`�v�
C���M>��|���{�5�#oO�at,F��Q{�X���ץ%��!��n��M���nL�!C��[���0�,^M��L�3%��JZ"o�Q�����NCv�<�Y�G"z*"��wb������[��M��_�����t�y���|�I�����={�AZ���>F����>���AI̿��
k�0�� �2+��S�7�v	,Jڤ_�[ 3c���̗g���b�gg[�U�
~�	"r���XlxVHYEB     400      f0tTq��ke�Y�����{���r�Bw<2�s��Y�	��#�CV]V ���6��$eހ����p�9���U��ZP[������&���Jj0F�b*bvE�F�o���e^i�Tp�쌊�
��K��"յ�-��{@?�^l;�pQ@�:0��:[��I��W26 ����-�Ѱy���{ ��������^̐|ѦvF|���i�!~��go�Xӆ!m� 쳰bp�HPDo�A�ʵy�XlxVHYEB     400     150��A-�Ĝʨ �j���[��nf���A����r��.��`��	�3Џʜ��I<��r�A�����c="c>��~�̫v$���L��7@�8+�������y�B�/��cIJ*�PW��ܶi�0#0���5 ~�xy���Ϗ1�o���>"S@�ݛ��ҧƼp�ߗ��Ur�]��W{�n�k=�����r�V�ɍ��(�v�⟑����H����O1���\�K�[ǒ+Mؕ�IH��쾞]R�f
֕ma�P7��g�h�8X�c�iڵQY�<%y�M�rGj���v����|x��(���.�7��i�~��1$��b��(�XaXlxVHYEB     400      c0q�;�o��F����u#��rd���bL�Ia�x�Ш���\�;������Och�tc4t�q:�Vjz?�Vl'8����4Xz��/�&���*`O��:Z.��FJ+��ʌ7�^,c��	RB��M���u�y/�hO�.��תP��b�7Lّ1�]�醣o�����H����2y�8ͽ߯v�XlxVHYEB     400     150��L$�*~���:JM��p�l�2ͼ����q�	ohu-D���ʈ��D���F߀�334$Tr$��k��M�E�_�ify!�!�h�R�2b28��y��E��P���j(|�����X��rl�њsâ�o�#�H��\y*{�R����j��3�X���s��Oq�i���C�����{w�3���d=���7�?RHo���B�[I�!�XSY��?��-���h:�	�F��T{���T��F�	1L,�����z��1@�e�?R"ri��s�%,n�%H�1Y�aiWf�� ���7���c��kt4o���L�e�0�)�XlxVHYEB     400     140�?i͒�<�n)p�!t{`���N��4�|՘��z�)z�����.��>#b�`�F���j����0?��<w0� ��E-U�S��
1n����!J�\qݲ]�J�y{�?����d3��xnS��SgaW�/D,��~�!�b�qķG-�G�������DّHw�x�P�� ����W�?{
���+�,ޱ���3�Q�챦ֳ,�w�H��A�LpB������uT�J�5�f����]N70� �P ��VUS�g�Z�!����vU� ZÐ�]�MD��#;�n��wG29:CJ��/HK!�m��[<�k�XlxVHYEB     400     100�4�u+�W��q����̇��R��Ss��׍G� eȠ�bK?��	�K���p�{0R�C�߰e�*<��qq3� Mf��}5�̿��CI�|�2�sD�/��mn}�Q�Ɨ�d:���Vz*? 6H���N��DzO6�~H{�Z�Q~�{�oq����h?C}�]|�7%����P��s�&��^�1����i��X����	�:�UGW6�n��헭����\�Uã_L�uͬa����+?đ?���mjN�2XlxVHYEB     400      c0�F��o8^��
Y����R�"#���rD ��2%�&|��?�����ͻ���Zs�&6��̃Znz�r�����d�Jj��Q���-3]��a���8N�q��;R��Sk�l�ޜ���c8 ��oLv���q�q�i<6����җ��LJ�6�J�s�ބF?Ω�������α>ภ'�M�XlxVHYEB     400     100�Zk��O��i?��xGTt	�cC$ҫCj�f�/g�E�e������;�@"�]O�L�o�m�e�ޔ8r㿯:���~�\�f,-��s�w|#���9�� �Q���u�m�Vv�Z�r��%�FJ+j*봧���/p8z�P�d�j����A�-Me߃9J��;���r'���fa�U�%%OD����РD�l�f��ְ�h��]r�tQA��X�.f��)� #J�	���H#a�[��Alf�
���!T+E|�ߣ1�g�c#XlxVHYEB     400     110R3si���v�����Y	�,0����+\}�ed�y�����k	�&=�.����m���^��QvF��R��w��ֽ�l7i{�c���Y�2�`�s�Lt}�ץ6W#�ܼ�srůz�� �L��x�G03b:����6m}:�T��v|_��?�d5��>?/BKt\M���# �+���Q.Ml(��w�A:�F,ZÌzJ�z�J��ޖ�k6�W8Ch	4�#�����Ck�4f�6�]$���r�� �p>�Q�~� ��=�{��HPգ�XlxVHYEB     400      a0�i�`]Y9�/��E���*
�6r�d���n�i����a�]u��%F�]��bD@G,��Y��-�: �P�z3�����{G�.OYK�%|N�g��D޻n�Z%^�UM2�@����?���� �u�^��ȕ*�.t�<����3�/@2�d���&=LP�R��HXlxVHYEB     400      e07���?�����o��1(M~�*���	����O������v��#XLȃ�w�,v�X��6?)p����ki�J^��J@|N"El�x>�X�7�h�2��qYw�X�M�[ ��8�����A.�"���\����V$y+-.��ҏ�q<"���0 ��r
Ӟ�؎�4��CG���<�Xs��,&��o)�V��ƞl����%y'���V���C�Ϥ�Z�n�XlxVHYEB     400     1a0T,��I���D��Ѥ�q�����C",�n��'�3SF5w�[�1��x�[�r�g�O880�w��c��hG#�9�Y������Ã/B�"��x��Lq \Jb��?�y�]
x�l(/�n��J}��[��f����hw��e���`�ǔ�ѡ�س�ڋ��k�C��Lv[E��U�V��N���l���s�XĆvY�9���_��`�c��C�f��_m���/�R�S��3^��*���쟩�wy�М(N�[�b`T�yh�A4di�{�ֹw�����D�)$�l��s�+8�>�pv�jwZ<�ͧ�(�ә������m�$ȗO��ؓ�s��Fy�'�����ŵ�b�3����_�[CUW�_z:&�n=�X�"��<T��~˥ZO��?pI�&�0�l_�R�{�<���v�]rzcXlxVHYEB     400     150,@�Y�"Q�k�� ����e]�OÖ���'�d=JR�=Cv,��~���G�����U=a,���,�tT�N �3�7�P�aO��JB�4�F�y������8���6�6�~+S��֮3펎�}���ծ�%���� �q$MA7z�<4�Iw�H5�p���Ʀ"�@�2�ԇk@����-ߪ���g~ޘ���Vcӳ��1��,�<��y�s+L��0����Uq-�k�o�6>�G�?��}C�z��ϖ6�%��e��H�QKyxe�=Q�m����� B;��`Q�&��l�@@�|o��:�n�?��V�=*��t�XlxVHYEB     400     120��3�7g�=�a�yÌ�BW�Y���:��KI5P�����k��uy~G��U�j7b�8riV�L��È}����0�HJ/q��fҀj4�[�!w���d��EE�U��Ső���1��ݡ�eIPb��q��)7�%'�1xx/Ȳ\8��#>�e�ŃaU�vN�`��ˮ��|ں3��g���[T�O�9�	̊��&�
�BkU�f��)�׃U/,���O�^��ws�`E���s�s�%�_��S�,oۻ�u�W�oƋ�� 󗍧4u�aV�\XlxVHYEB     400     1d0�y��58J��N�/�9�ᪿ�INlL���Z.�XHr&ɩ�MW�Ѐ���^�u��i�����]�] �Z��b��� }����0@�(@Č���b�P�� ^C�Z[z�����R�8e92�W�".�>ȓ� G�����!}�8 �c�*�b�yp��-p��(�`��v�i�c����0g�t�.���3�&�H���ә8X'1}kr��}���X �ܻ���I�\�bn'���Z��)6킼d�,�)��1й���]�?%zG�J�q~��R�&0��������V��fԎ������a���#[P�_���w5l+�z�ZT�W����;�7bC�F�ڗ�2x�W��賄%�e�0����5�wkD6��y���2O+L*��T˄�8�n a��!>���)���z��y��p��Ϻ�Y���?NY!m�g��Z�jj������PXlxVHYEB     400     120�v__/vF�3����*��<��3��]$(؆H(E �6�i�V���8G���h���6������6乤Tf�#���~eaX/�ΥE��z��Bf��F�H��� ��~���$H������߱t���-��>a�����k!�<b�\C������SV"
�?#��Y�=��*4r���Y����S�Gr�i�%�*��O �n��� a`[�5��r
[5�H�K�oԛ�2��FsL�:�ԁ`��'���0�i��Q�2�x�w'�-��XF��Y�XlxVHYEB     400     100ڐ�Ɖ�8躣�F���iQq�`hSw�=�O=�e�p���1_]j�6�x"����|:�ʛ�D#j�	m�l3.�A���/�=O�?����7���3X�E���U��<�CW�y�?�N��gҍ�Nm^(�ʶI���%XW�!'��(�[0�Pxx����5�ਊ��2�r��3���pgOO.�V�H�'�)6�]2�uؔ��D:�b�l�݋��	ω9��r�);O_�T�#A�L�[+Z.��B ���.cXlxVHYEB     400     110�+�r��M<K�GV-�!;n�v�9�D�	�	j�J�	_�_����ml�$̐d��Lim��Tz�"]X���^nZ�(��n�@F��ϑWW�P��}aR�N�;q�ņ��{)���Φ0s�s���ި���Y ���t����^��mÝ�(ߕ�k�����j�����3ø�ق����Ia|�+�[��N��B1�-ͦc��Z�a&Rݲ�!��;:F�kuG���-�YĈO�T�+7a��=�U+��D��_��j�c�[b��|�K��og<XlxVHYEB     400      d0;|+�Y�&%2�* 02�Pܕ|õ(�d}�T����#�iSP\l��nx}_xmY���8 Na���&*�]C�5b�A*��E��.p��+�](:	�/-B� x7��w]��b%��xo�Vdv�����C�|�R�l{?�I��?�ld�2����L���K�Qq�]yN ��^B�պ�R�\��;�:,��D���w*G��H�*XlxVHYEB     400     100�N`�3D��0�ULlߏھ�K��f�.�S��&�7#��W��g|���G�"�3�R7�=���W�FP�['[�<,E�r��'Q�B45"373(r\���qa�6�����;����5-QH�P�� �!��<�r{�󱢨�Np3�9qTυ.b��\��T7��q�%���qv��@�@HR+P��a� ����S��w�%=��Q�)�g�L�Y��)���J$��[+O�x���h���S ������m��^�XlxVHYEB     400     130%�_������<���V�)Q{m���#�i}�)�9V¯����,���6�<|�! F�����AnrOW�p����R�x�g=��x�,ϰ�ᰌ~��?�6�j|���Ĭ?B�]�#�z�٭�P�w;i����Ā��{A�xr�u(f�y�FߨG��+rM9[�+)x��5	V�ur�������o�H!�n��J���MGy&��0t)����m�p�~�2�vKde~wty�,��Y3WՍɆ���ѩx�΁ȳ��O���R�4���L�]2�.�`��49�=��Q���Y��O��pXlxVHYEB     400     120h��.[�%���~բ��[wh�~��^	E��<�1�eYj,Dq�q��y�$��
r��܉�l�>,��E�O��(r,�8����~<W9<>�+�0��+W%Ʈ�(�<��	�f�;o+8�/݀i$�+w�&@C��}Y�k]c�1�"T
��5pU/���U�E:�O��_�"���:�v��s0�(�T63w7-'�=����߾���O&�Η�|B�V�����ѩ��Z.v�݈��6��!/6:"ГC��Ùfd~)F�`b��UuU#��9�3,gXlxVHYEB     400     150#���'� �>nx�cx���E��E<��#�8)t�ɒb���}��I��e�J�{l��͗�"�nS�cC�ڹ�*���:)�Y�p�"s@'��n�����OR)+�7�}�}�n�4&<���O`8������Y����y<Û�D���xW��h���)I��ȁJ����	�!0T��	�f^���a;"�L���@��]s���;<}/\�E��s����f��L���őԗQb��q3C����� +�j�f
�@ћ�)E�{�x»Uy��������1o��n+��֤�!n�gs������b\o��J�3�3?��)�YXlxVHYEB     400     110�#	ÒVfm��j����R����Hm*�L3�h�I^\�g~��9�'�S��" ]j4u�J)�q:3Ձz����`7���4�S%B��}��o�r2���u
:b�.=)������\UZ��tե�g�}�����F��6Q�K�L\<�7�q�h>�x_D�T��2��d2�3�c��J�X��7�6�kcY�� 3��{�_*�`��XĞ�,R*q��ΐ��8�k���`V'�ZN�tsv�C�/K�39o6��C⢻`RSG��0o� &�XlxVHYEB     400     110d��H�7:_����q��˒�~��7&Ku_���m
�<|�ꟼdS0�uPQӶ�k"7*�wͽ�>�[���ű`����ע?y����7����vi,�+�\�$�� }��}b��ݽ �E�����|�Q�@Y^EK���R�N�^}���ۆּ��2����[��2��n끮dy��e��l��QQsCo4�f'�4�(�����w�	�#������M�T���mn�)U,���?ʞk�7[9���Bg�YZ��Rtk�ȃ��0�2;vXlxVHYEB     400     120�`�UG	1[����s�ꓻD��:��E�\^l�w K��
���N�Ʊ����b���3tQyd�t;a����1H´��/�;����d&���0$�g��A�x� I�M���M�/�ė0���S�b���Q���>T�o,�V��������lI��� ��b��YUlf!s"�mǍ7療-��~/�'��o�Zu|�"����[=4�A�
�)7�@���(�Z*c�m͞o�Y ��n ;��`'!y;�ȶ\�\����Y��=L��XLbg�	�o�� }�*�j�XlxVHYEB     400     100����QYvW�Egk?�|�����^1�ǹq>�D���[Ǖ ��u=zu7H]��d�+W}.�p{cO��4���l�!~��Z�2|F���3���
��C��($]�f��g����ƽ8E\T��ȗԧ�����-)���0������[m�HGF�2Ǻ��Iut��8�Rn��X��y�Ed9*C4E9�P��}}�^�݆24B&�~׈1j}���c�\�]�n�����t�a�>ř,W߄��:216XlxVHYEB     400      f0�%�L�'f�J�� zr.���(o�T��������V��яtGn����#6DK�>��:|�����:�W���� �0?GU���e�����1�@��%�x�P�%(r�b��U�fJ@���o��z�
:���:�~�|�
�)����@V�y<�z$�sMe:ΥnI�^�N�+�)��̒�\���;��3��D�`��X�����+'��N*��Y��\X��:m��@��j����h,Y�XlxVHYEB     400     120{�g�MW ��!+2����#�1/1�:l�悞v4�$lЮ�X�)U؆w>MHt8�C��`y=͊���L�qƉk�`P9�(�UQZ��o��ʯ�WF�#uM�%�^�����)e˗��\mz��iUD%���^Y�+��N���5�f�F*����������Bm�@��&�tA��&�Sc�uP�m3� C箟�C1���l܊3�V81F芺�+����¦[?Q�@�@%��F�:�e�N���Z��}iw[�/`ڂ�7J�b�X
{��Y�Y�63W�hQ�I? �2�5�
.XlxVHYEB     400     110��D������Е��C����)�j3��2���'v�ߊt��$�7�#+�/o�RL�� ��w��&ቃ�2��եk
)�2X�ΰL{�8�Ӣ�3 Qܪ���x�h�n��(�bu��]���G*��H3��%���R(��l�MI���].�)5p,���ۆ����d;K�TU��ۈ&x�V� � �'��?ß cc�h�!��Zlܰ�P	F��F��q�R*�Ҷ�D�'q�Ů_��鸞v�L|�g!�z_��;ϥ[�s
uXlxVHYEB     400     120����5�>3\u'R_>Zݔ�zLߠ"""��̀�[UV2�E$Mp��"�Ċn���3I8�%k�J"\;��6�t���X����ӗ��K?[R|	�V�C��/���H�v�^ޠ?��̐i}�Q�'�s�@0��n��� �H)�t$b��S	���rc%Q�rS�)È�|e$bĎ����hdYЈ�㚒�d�$L��^^�w�6z���.o��@,�F�tFT�a�~��ب�mےf٩5�	���|v$y~W�x���DB�Z����SJ��Mnd�̱�:B��Q��u�}	XlxVHYEB     400     140��!�Cٻ�]
&.ag��'k Q���6
1�/@�����s�ryyƺŶ�rm��Y?�[�����@�U#i�RA��qLj����R"w����i������)�׸�\2R�N2��	\0�㣲��=e��1���%��PRdr��sK�G§�B�A���މ"��悗�u&�>�����v�^`��F׮���c9����=�����P%=-�Q3I���JOu��c~6��)�ڷO��|kS�-r���C�xeK�ܰ�^H�~%W��+��Qi�����Vv7�a4����a��dFຈ��L����XlxVHYEB     400     140�}b�<^G�%�Axwb����oq�a�_�(�~a�[4���x�xU���L6�JK�T�?MA���XQ;B���0t6�j�Em& L�h���;��sZ6�.5F	�=�#B����q�Ub){�f.G�>��2Oj��h�q�/9����']̂�3TK����ݜ9s2,�tP)�k�D��*�t6�#�d�T�㓠�Gܷ�fE<�U}T������ot�h�`\k
���������P�kڷG�jJT�%�oI0�[���hJR$�.���L "$�+١�3�,ڡ�RU�Y��u��O�Ö���U�h��d}R�*XlxVHYEB     400      e0���4X��L%�g��\���Vr��3a�N���!����$l#����ɂ���LAP��5��c���eըKB��;?��)�ޜ���2�u+d���DW	��$w
+�mp]�L�\LV�/=q?Y!A �U�N�y�$	I�uU}Zͮ�`FQq�a*
w��අ4؇b#ј㎰JR&
�����R�)U��mf����z|�����6'���0�E
��ڝ�J��rXlxVHYEB     400     140�4T&yI?�{�ɑ�0�n�q1�9n A-
�sKlMy�,O�Re3��d���=?�7�K�>�M�y5qٳ�&�&od-TJ�ZMo�Ř��+��E������밳sfЦݘYY<����O&ƙ��=\xgJX��$>
YrX�G��1Y��nJl��1Ϲ�),^�	�8�ߧ��lߑ��'�����E�
�S�'�Ao#�l�����ʈ5k�D�[�������E�	�m5�u��9H'r;��]�[z@$���;L�&:]M�2� qR���y��q�h�F�>�N�~�~�	\5MGX�CH��z���AXlxVHYEB     400      e0���H=�$�
�#��$n��8'}%�Uc|M��9j/��J�^�XF%�kTK�����l��2�]��$�䫽���-;l�΄�d�vb��N�c`t@�S\{�;����s��4#L�:���qK�l}j��<�JX�yU�-����]�"��� ���*~����z~U�c���c}�C��=�xZ�=�����`⑔lbA{픵�Sj�� &��*ԽL�XlxVHYEB     400     190l'�m�旴�u��캌�N�▤��Ҳ�X���3ɰ�g����N7��_\��[�7#%���b�d�;��=�	r�^ؕV$V�$�#S�^r�R�du��Џ�g�g6�Q�q ���nQ`P���q��E_s��ߓ�xގʺ#�F<i�Oƚ�f*7ٔ*��M�l�.�#/�f���9|J�0��TC�LC��s�پ2͈SO"�r�:T��w�ܿYy��!�|&ٜ���/�qU
ʆ�A�+SE��䀵G��>+c�����]d!�� >�ؽ��c>�s���}BYg�0��������"�D��8.�cx�P�����j�7�b(���X_Bp�5�rDr�R�eJGp�O�Xfu��[�幭~�:��iU���l��dU�Ô/�.�������7F�36XlxVHYEB     400      f0�~�}\���:G�1��>1J�P���E�N:�a	����X.�̵$0*��-Ĕ:�V5�]��S�=�izw!�d,o��Il�#.wף ;h�`��v�nl�mu�q@C��2���_i� �<�eD�S���������;�$ �)�X�g6�9���]��� �k���R��
E*�F�����.�C���C�!}~��v�j����M`|��d'��]��Hc�l�P$�c����$��Q��XlxVHYEB     400     120f�z@� 6v�%`)����>3��W�v݇:j�� 頏��&�NҐ�
->��M�6ѯ��2�,*w���!^�#R�L�TΚH�aT�ڬS��DWn=��h��V���`x�mL�P�Gף��P>��~�����{l|5�Uv�����~�sG��|C#r����( H ���pd��#P0�?$�P��2�%�|@��Z�����q�]�N�o�0���cYu����{27
\N	Ɂ��z�7�T�y7��ψ;�,˩�v�3D����r�W]�a�XlxVHYEB     400      d0ɶbRe0`�k1,�c��źz�rN���7>��"w ̯���+Q�{���Y_����>���F�)��q��	8�<��|���\�7Ïdo5D����V�h�Sa���͵F.~�c������%���8V4�iHؙ$L�K�Af��P�F�m���=��Nd9\�������V��]b�h���,��?E!e�eG�n���j��#?��N��XlxVHYEB     400     150��P�T^�mz�@��4W�&������
8�;���7�{Y��w}�X�&@���8�A���U�m }z������pqB.�����Ng�d�ƨ��~5!��K.�B��N^�S�4�[ЏCz���i8���\�o���NO�'�y�,3�>����@,�,��@.�&\��A�v&Ԋ"3��� ��\b�z��8|�W��H�A�f��2j�(tJn��혁8V9�#Yf9s��j�u���z�5{��;јIk�6�'���H����2�TIs����?g�~��|&MasD���k��8θ���ϼ��z`��h�7�N�B�\P|̆#��*�
�7��XlxVHYEB     400     180�3kxy�ޱvq; 3psF���.n��X%��!#�*6
���� �)Z��~
$U�h���0ްe\l���2�K)����D+������v鰾�*�Rn@���?}瘦�����r<�o���XO#�Bj���Vw��Iu>>�<!�.�ˑ�S:���FS����F*�*�y�������C]�󈬜eU&�����������D�S��r�4#7-W�^���X��G��ōu�E�y�"��e웸��U?5�dl����L�}ٷ��3Q��Ƚ�������Iv�Sm��)��in��K��a��Y����e����Œ�<�U�Gb��QMEi�d� )E1D`�����I�~[s��T�_��w^�QfV-�XlxVHYEB     400     120��㑀�?��?g���é�6��y6�@����<Nu,��c�F?�Ӳ�ֈ�+���3�p����C�������ʹ	���y�K`DBT$yb�����&ƿC����߈��bڍ] �a1�D��P@ N�f��]h�>���!�4�h�*јR�>{g�a+'�U��J�1/�>_��,��Ey����𭼥
ڊy�u�H���Ҟ���T%���ħ��]T' �������l���7�r$�8��k�qFpg�&��|���[�Aʱ7�|HR�]:mW�XlxVHYEB     400     180�Eƭ U�!��a�Ʌ¾�"��/O�X�Z9Zvv@:($������#ǆh7=��`�m7p+�8E���M^i����
@֟X1hı[���l�Y�p�"E�C�)3�Q=��Xu��>�!�/����b�G���\���1�em�E�eʨ�Щf� �����:q�F�D����1���?
o5����[��=��}�*����מ�BA&hG��m���!ԋZ���Eky�&E'�� l�����N���-ycGj_=8f�L�Ȅ�Y�ر��d%x��ay����ׁ���pzi%2f-��~*�V�}��b�p�x�z���(d.`p�^�o0\���ύ��V̙t \:�����I��2s3̃,D߬nL6�6S��ʶ�>kXlxVHYEB     400     120*)�Q|z�$2�L��w��Q5җ��>�&H%'��[C�P'�ll��1����c����vo[6!XUs�SvꞤ�F�g �'������HJ��w(��3��u����ajF#�+ۗ��g�;�6>R�u��]�,�ի�eZ�@3� 
�?3"�����0�[N��묳�Ѩ�i�dĢ�)��bWv��D]��v��=�Y;�������i��Q��Q��<�.����Sz�z�&0g]E��C����P6��/�;L$�_��:>����v�XlxVHYEB     400      f0�Lx�zFO;��+��:��'$i�������s�H]�l�� L�q��}5�e%�'�й$��]��S���'�i?G v��,3(2?�U��Z��T���D)[yͺ�;iTJ����Ѭ����|���$v�"�G��ԗ���E>46�BHM!7����R��m�+�N)��㒛���tP7p67�M.�! +?��p�R3�)� >[}� �������[�
��d��Py���XlxVHYEB     400     130�iUa	q���/�KY�*ѐx�|�3��Ӌ����t�k�0D��+��m_)
�YT [6�[�fLρ����z^�;��M.Y�?_9��<3׈�YXP왩`�GA�)]�j�V��е�� �[)=��t��V5��{d?>�Qo.��x�Eʠ�b�T|U�[]�@̝fRe��NJ��+���@�GM��a�X��)	�qV�kK� �z�F؂7YkN
�x�F�S.�<:e.�B�Х� Ie��Ϯ�\f/2�d4@�`��Y;Ȏ͆�~?r�x�����9�W]F2��U��XF�����4��XlxVHYEB     400     140ܻw�q�c�@���WY@5a�>�q�[����^������U�C}����Ktm2��&�	"H~!*�Y��]��~zu���Jy6 �([�_7ߓ1�c��Qr�FlkM�-V�,Rm��n,�[�,��A�ړ9�޵p���0�V�Ӧ�*l�r�D6*b"�hƽ�T�}�>˦`�sx�P�v�-!K�^q���lT�,��d	�ƭ�W���t��A t���05I�ż0���G�,r"ގ�ٵ�膱O�9>^�~*�l�n:�!6T�}Z��I�F���v��l��K��یR䵈�e�·������� tXlxVHYEB     400     140���x���1Eqy���1|����r�����z��.��tk���M�zx��{."����.�pYD�s@y'�FswP/��yox)�v6WH�y�[Q�/̘-N[�f���1Ǫt�7�M�N���j������Ò���P�W帊'_ܘ0nh�Ha����8A�E����������%XC�����}��3��B�xVp6�Gy�����(Rh�4
ʲ�E�1[��*gi�k��
Ÿ���QMo��Ø�3՚#��m1k��}5��.�{��l��M�n�CD|%=N�3���)���]d�8dҨ2�zXlxVHYEB     400      f0vf?�m.i�o�������Т)m��R�.B7ލ^9=�W[�Gn�if;�{嬹1��*�K�i�
� Th��bu|�<p/2�r&o�dk�wl^^ӴT�zY��)x�B.8�L�c^M��	1Vo��߿�l>��ۇ����R�'d�҉�pV7���N�4���I�U +�rFU������i+h�r�3�x!LR���"��֔q�;��.4i�3`B�����-��jا�O��r&XlxVHYEB     400     140��{J蒃H5��u0�!Z&r�qٷI7�.F�@��8 ��!��� �el2A�ْ23[��ƣН�
-��}��p������d�q}�]}V��&����!�N���QO�����eݩD��[�<e�.�(�֨�|6���R5;7�TF�3\����1~^�z<~���jd��������5p��P~�c#l�"���y�����-B�*���8����}Hm¼��OKm���Bh���8��%d�ѻ6iXq��� ��IM'�k�cGV�����	�#�R"�!!��c ��Ёa�|H��� ���7>F�i {󌼫,�XlxVHYEB     400     120A?ѱۆ�x�Ƒ��1���)��b���"-�g�j�+Oe�ޭ�7�����	Kʣr�V>kg�M�hz��+ߟF=������t�l��V�B5Kihʩ�zF��sΏ�?���,�)�R�����	�w�����?��8xx�[+�\}ӝ���|�9s�Q���V��Q"��%�ϗ"���I�ȥz�=?�A���h�P����ųq�����~��2k>M�*=�W��4V�����������z�/�K\�YdB�j�	�A ��lf�l��3o�Q�����H�>��A7?�����/�XlxVHYEB     400     120_r�[�%oNl�^��׬B�'�i��U�DD\>�%�� ����#;��QQl\��˨e�Գ#��Y��Ii.�� �q��;�ra����7I�/�����Yg^3��#��"�W�s���S��y%cZc��#��'���u�`���"['�X:Jb�x����섂P@v�[H�6W��o!*�ca,4�~�'i�,#�'��� W|�X��S(� l���Ӊ��|��_ٟ0���K���vw�ޝ)�je~�IF����l�����G�l_$�vN����?����SW�=�G��XlxVHYEB     400     110LȻ�ê�Գ���A�a����^�^F :N�U��h͂�:f���f��eaS �*�\;�<��(�N+�@nJ�훊1�q�j?'��<H��,W��U
�t��P���l��H��<^�>V��M�r����V���gL˅և�IQ�*i߾�D2�8�FzMIi���^��w�9fc���,�{����[�x�d��ЈЛ�!��F�X|�Y%���%�6\�xY�{��)0�mJ�s��݂>�CTK�?��#�'��L�e Y�"XlxVHYEB     400     160�L���r�:	]��A�cu�3üQ)][J�>���������jnWk��z�yicL����󢯋b$ҹ�Y>w����<'�
NN6ܔ��º�&��&�8�П� �=ԅ���h�)BDF��^[d�A��O~(8��ca�JFy�"���d많���K��M�rw���-����=ۻ�|�5P�o��gG�M�� �L,��|y9 "
��S����;���1&�T�fO�M%*���f4Ek��BޚO����U%iWM���Ya٢��?6��u��N��[(���8��9N@?ʣ���4-�Y8 0O�������$���=4;�+�I��� -k�}k�M]XXlxVHYEB     400     130��v��'���������<�>wߏ�+�1���#q�MN㽼�����?��V�-<��k�F��M�0k����+��Z�a�owDY��!�߷�Ք?-����])k�P����;��Q�ҙ�SUK�xzB�(�d��w,�U���Yn�䍆��u.�hp�͊P �4�lltbEZ���l��sW���A����яj�QQ)�4���a,=w&�'ٟ�3��f�D��c��1!R|��g<��E���U��.m��e�1K��KJ��7A+��W ���02���R��_Y�Qj�xH8UV�,��b~XlxVHYEB     400      c0��XB�M�GM��F*�l[��`j�ݦ1Ȣ����<��X^�k�2�E���Z�O�8.:��<$<8E� _�Ǟf��zgm4��FI�����:=�?�h�܏��Ժ_'f��83_v)�����~X�������K���� �CL�!�`�l�v�̎9آ,�k#�����ve�od�t7h�-�=T����XlxVHYEB     400     140j�c��KW���1�eŋ%"z�R��ĕ��eW;�]��� l(8m)¡�C���tQS�ҵ%�;.��:���=�xy�%�ՙ#j�Gi�j�6f�sy�}?�& հ�G������w�:���CBF�˪�D��![�׍md�<�6�?&]6�Y�DW�vt�u�M=���+0���д+�(p���s��VᏧ�2���	����JP��L�JQZy��4�iRP�3p���3$�*���[νЊs��4JIr4r�����t�lJ� ��($c\�)�1�
��X�;���f��+����g��8��xaSXlxVHYEB     338     100��g����^$wށ�&��޽7@��A�Hܭ�����M���v�JjQ$��Ẻ�8����*�57bjJNAGɆ���!���X�V��uc����*��ֿ��Ep�;g ӽ�}��}b?�ױ��|*�{x沪���Ns�z1컚5+����śJ��L�桗�<gL�k态�"�4K�����5)�qo�LM��xW�<xsx�W�Xp�����y�At���]H����	��,��{a�\��͹�͘_�
|��C!