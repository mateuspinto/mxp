`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
LHRvrnRls+bxY4C7Z8iEt7TMBhoJFEjhraBvfv/ONQMBF3+p4XMdMcT2Ow+S68jOZeyLXD71ff20
cSlFjcjvz4n5ji0F9CjYZWss/42ASBX3MTeSO1Ygv/E1V9AdJ/H2BeM1NjXN+X7jt86Z2CzYjGmO
fP0/VPt1IUP/M3d16wDLKjNGW2dRbjlUokBhVORQCRgiAN+PBCb2vHFM039a8QLOh6dlXJ9oCEQN
H+YNjJvsiPPfL/ILg7JG+q34ub/magGEwnPjhXghlPmbcRWDpegLL141aPJ+J3piV2QoH/NWkfGm
RAvyirqcptjdt37Gv1KFo2KqnQlCyTWxAiYQ1dK/qiUoEiL71err5PEv+/Qn70fj7H0P9cB6XD8y
asxgXEWT8xgvQUnBGe1W0z0gz8pgNSv7yW5UaFte2yq+4ij6wj8rOrRq0kTKkBQai3xEYLZxvFbI
pSy2CuRT8+7Wk2XXbaPuZfjucyA2BXv8UxgyOPKh3gNECRcc3PpO+nFMC/6iNOtl7CWjrhEgcQwf
TLvA5Sr6DoCEaXjyJC/XdI+IZuKr9c/Gm2kZWD4Sx/Vtfi5S+LUAXeXhsAfqofkssCnBoQPinfic
hqD6A1reIh91h0jTyZCTh3i3sTNZ3ovO02XRfDzkq1C40FCJ/75bfJaLUUO5ZpjEJE2t6MqBl5fx
TNYPAOYPKfaFxSfQxGyi7NuThx2d2wesLD73e9YOFZoHgBTwjUpwrgXRnHS4GA8SK2IBTZqzTNTB
P95WKT5ZOcYcIdgrxxOiAWcqFq8PaTWJAttCdyZ2/rcE0ldSwLu8GS5JTTrcNbCUxk8aXlb5IdHG
smqMU8WjOiGRmmSmxQxpQXn6DldhYNLKZYpt4lMz3E9QSz0fjRZ7rfQqZ69Ad/2afWN3AI0lR8zL
lB7jhBIeND047xmA1sPxvxWU7dBbrYVoFsIfIQ379A2tlcS4DXa38pBmMT+52RCej85AByYsdYDk
rTC372vwCkt17XaQ/ge15BHJbt7+/oThUY+cp5ZGMwtLF5LVp3Kwni1LKASCx8kN5uw/4+lKp/4H
dUzcehQ+m3pWYvCjlOzO0p55LPpI/eJVkn2hK4xx04Z3JpXwY+xy1IN0u+CfGGsUeSQjHXgBbInh
hqALX8/hmNFZCV7ZerUQ3Jtnq6xnSZZxYZ78N6Anfo66rWVbRtpIMjfd0yPiKGNaOvDNhY2cKCJ3
rSCQp4CfFTfjMbWahIo81ort/DGMsdgm2ZeoVN9kta52GHqJArv9uTBvmusyHxxp+JP2fCOMJ1+i
BQ8B1WY7V8dRksUChCrP3lS4A1HeZqb5DjYqd2HBMuM1RsJFuhjrcmE2weuDPbwWlDg6mKH5rPzK
8qKVBD0+54Ox4xJs/msPG6X8kUtD42E3C2J59a4QJOWMrtEVpt+Nr7ND3x640QGdEY80QCM47saI
GZUuVupAmu4/u2oRyLJMfU4Y1h0FOqdP1f1Z8wxgs4lBDrztkLHGlFxtNuFPcAyzE2x4RVLjT+vj
t6CDmhPXsz8ilvkc79wckvkXxYUpnNKAkXS6lmZoFPE+CidpojIhqwmjlCfyMlMlBc5KzaZXnXWJ
Ax3UoB6Rll5KinAz0TtuVEwO3kOnAJ5LuJL/dAOJvj+dX3hF5JuB0E0A2xqmDsiSLOgrzHHhAHLv
Baycj1uhi4v2Qw2FxrQ7PQLsNCsCDw9lJ7xO/S+HIj+5NWu1cTImYJ6hfxNl+1FmcyFngYO/JNK/
djOwPDw7jNqgoGyUf0JHQfNxf0rPzdsBFehYfTknkU8BDcKCPApi/qUGB4MP4MKdthn008TWPuJO
bUUqQtU/jMGke8srni1fMHnzhQZAp3zBGroq1YkTSUJ5OdVeeihnVMFlLIrDzkfoxVrvVgPR913B
jRADXMimGyZX8/qAPRtIY0fXpIEHspNBNAVJOvBzqLxtpec+p27LFKJ/n3Hu/ua0zgGNqw5KlYOx
jiwsLUemejO7Al/NtIZ6Jq+617QMcLSXn8YGCekOXgTeoL9EV8QiyhHxa6Sr/chLTERTU4Nxd52w
M05q+0B1Z2YMeZ5deY6qAqFDKfPHBKcn+e972jLwp/uLEu5aFYqX0lUR4TFwoE3RnphPuqHFs3KE
fDSRAynPJR3PkVLPOJ2Deo+XoGIPl4N3C+thEYMmlFHOV6izaDH1SGslX5f032p9/3xt0sQf56XZ
6AS3X5uihJZCRUerEhB7VIt+r/7fTDKsgSiE3ZotS3y4+WZtTPTo5EPpSun8UzazTIIAFRm9LGaL
hE8aaPtaIG25IXjy54Qy4TlMlBMbHFRqqxpB7Wh4H3l+kl5A20UXUSQs9vlt7CPfuYFeFk/zouSU
Gd2f5r6+IXjKGsx5G6oJyFE4UQacIiVUgTmQ/s1m5+PccbZphmIAQlXJV0tdGYAXODH3R0wDBmhV
WgfSiTNMqAaGZpmHp1tU97+YxArcvUnuIyYuIPb+E2rVakoCJp3IM07i2Z+PQUjBiERLaPj2B+at
r5RU3t8sqODcrYU/J92cYEvQdc7B4TnLcB7pebvrWqo48LGoDDdLxHs4rRQP8XIniY/ftSTCgD9h
NxKOIK6vnpTMb6VmCFEL3hGg7tERZOG8CFhgaORg+1+ftx3EDOVIU2+Pc1lgEMg6QgCy2gmFxGhW
mS42COMFZfmnMSX5wTsF4dbo/6q/TQUt7bXSi/5froD9iVug272rNeL908GV1jXHvx2fAM/6HZSf
zPiA9MfZU0fPERb+RrnFFwTtuez+DcIBGr4hRHaOtNZKd9XbzYqjmqYUOfdlSXhLbOMsOGlYTXP7
DjVlGPkGmdWyfOlXTogYNLRTH1QvmUBEAes9US0rnomCJ5EALLVEA20OSqz3HiuXNflVAaGT3cTc
wYd5BI5DrkGxysLvAuqWpX5dTnUKJ1nVq6j4+A+mTK6Z2Qsyyi4oVfignIjSKEBFrUizsBo3ysUq
zF0kn6oQjYokKhSTMFwszWcfJO4b0CdUsAHaL9H+fYUMOSpSi5BRwKBUVJtIQV3IeKq8wnjWBV4s
DevcXV0C4kO90fvUccdpu2vtLLU4heTsSTVBUmhHGoR2+A74XIvfya8LHolR5cOjQ0STku8oe+O9
CyF+g0DKu48WT7UANhV4UnLoe5rlhsOTJAGdMQhJgCB49ew2PJAe/QG5AuPx5FTk1Ih9Yo15a+j7
xvoZnxVJns20NRpyY4i7AZDhwwI6GH9TINa19/M0iU8GxYadY4fZ2Rv3kkgvCUXQgcCZFkGeL5Ej
EWVrfqbyLvwwIcPMWFgZhI9x6AdwRn49ZA8kAnEd9p0NeGG7AGxsCYgk7mZ2tlv6GDWeUOd0S4YQ
eOrA06eyh5yocM+r5KI0OTvvl7DyGL0oj/KQckjgWCHlSTQ6IuJxqKUnrvrpfkfL6m9PkeXylIkN
AJNaLKgk43iakXai1WKvLn13BjNBLU3c2kb+jKSNssEyzadhLReYN1nTRNN1f9qaz92Z7GVNJj2e
4OMpdtLHyjAnflXUsLbbX5o2rYnAuCKkTucChARLn1EJi8Bmi/VmlrA0jhdAHXr1p/4zXC1O6tqK
5+lLSG8kB5VzxJ0ggHHKdE2dQNd12r4lb8C1dmKc0MDCrZb0fmVZD9De1Wva7uQTjLGpnmaPp/TQ
79Gya9OK6Fh6j3tBEN8gV8w90tMvx188wTagyhYprzVUd3IlDT1eksLaZiEJU1POiA7Pv+1q1874
QNgO2mF/wE7uTgzDaVcHlnCiGy0VX7YIJ6EDdGCEfn4pi4Qw4u7COFbkt7UdnZSoxlg4RG72rRGR
rdwXkyfscjND5nAGiVI20dLgtkvqaUtrV658b6xf5bqQHRbzjYwsvj5PPl6Z37zp3zSW0git9LG6
TnmqGZyPpjAib9wuJ01Hrgu20Fv5uXnPeXAEC18DSW6nSMexMYymJm1IT/zeWbCAe0dWqncDhA5M
pAgk3STWz5n8K0pfR7BoUHCrzwFjtuBMxwEWY2I+X6yS9AmfZQlAaN8GbYuXtUZClw7xXBAllc/O
OM5cCv8gqmKytYhMUKCq49+ut/Rz4yZcfj/qQr7cn7aJ2ZG/qAhl1kXZVlv908OWDutP2OW/S33e
SK8iP8EhqBalhdycDI2DXkmxvd5gqMX8IKZ4mu6cAuZ279LZf50uzCyOuFMzBnMczXVxMO6HCupZ
g0Wq24Q2lvq4JHtrjxk2Mbz2aPah4YPYsvjEkvoGUENxl2agEhUo+GDs0VkX1d4DHGq70SFptHD1
esYoxhbcdjSjsFiR9jQnmhUaUrtgLEHyUIVBjotJ9rDwwqjh/jaBqobWAZ9cWrywNR1hReAM4m6k
IaYQvK/0gbZpijLLPHBntyYRpOo9Izq54mPbrB3RUyxGw02wh1n1v31Al7P6320biDEBnTCJE6Oq
2svY4BzL5+1oKyObdrUpu+hAQ8nANc8ap0mC1WEaYDTHIAumgUK8hKTb1xNoiZI9HClUdTejHWma
HUPkbNf5B8fWo+wsqTGJsBtT/OPHGJSJAm+2oQZ6mkuep0UjZW0eqqOvwEmo1F2F0YFSimiyGqK1
OgDgnIxJkde4hwcTsNd4l0N8IiV7ZhiSJQ4/IvhYQj5nFn/jwgfuyaodudl3bAPZ54P0LG9x1VnU
tMuCG79XesLsfQiO02elbHBzKQIegy8IUGxVNPZCwDGcpE+Ezm26c7oOtPUOUSYqIMbQSNGIFCWU
cUCHwU5uc6Sempwn/YKsQfoAVSnwCcUvDQ6BI4W5L2Ls9DlVwkZYbRJztqcePRuxRGqJHaMmbfFK
PPULMvueramfux4mh3Cx5+hILWqpfBgf4pIiXVezyKLnW9Tu3t4kmwlHfXNd1FKOh3i52s0vwc1U
pOwR0RWFb8pnrtFCATJ2FlfTo2AqQC8un7hKXEBvlEHW1w0IxRxgJ5rPiCmubEK4LadpPBADWGDC
7O2lN60D2qrIhC/WqR9ldPI5DMWMGhXll4W/PXV/HNnwylw7/8cM01YT+5GurDJjArAKmdne5SQy
+ZqIITBkkzDyFqrlLcTb6VL8ckedvoRrF4bMAaffoeBBnBwSMQ9JsPZo2Lix+praJ7SjGmA7B1Qn
7sVruNlZw1kScqQPwnA7vIVYAhsW0LdN0amCGMe32Q2CnZ2vekGdcQB2fvWzK0ccIQbpiKxCddoW
Qe3FNN+fuQNVb07UubmqcDNOYrj4frLBI5cVhQ506K1yOjLSgDR/7M/9/CYYRLF02dobXoQnvWU4
mMHC+2Sjw4NxIWsAykH21pGqsmFNhFcaxMH9KxUduVC/7mMMFq8ktA51xKvo2Ti31VNApMnNJ4RJ
xFcdBIdvLafOJRibYBcHugiTtHfnitm1luhA/aozlvforjsaGFtWz1/FP9QjVFxjTTovUx2KhsMk
nFBX14tzxryYvSp1rTzOYuTNc4Q2mVrBTw4z3wI+JRZdZlDHoInD4Ba+GD+DTndi/6t9DLUpcoW8
zezbVCkTr7KwDTZJ/X20m+VpPUUcGy0fbr/lXlZleOw5OObnZrUyVVrmdN5EOgmvf5ElYXe+3jok
iNQiF4mw1FDnVkTOQLCvIx+yZFJlEeHafcPbz6Mul23aw5vPx9oJgDHZujs3QLp6MQ5kYRfNs/PL
K9KZNeDlCoELNwCwRqP9lcbfwMLS0nk/3HQ17DsR4nyd7PIyVLoNCnRJkOsPz83ge2E7ge+3qxoh
DlEV9HC81DrX7GPK8f0c2b7FKXkwk8mJgigmTZvVJgUVE3DmTJ0Rv8j/rcw4sCDjVX8Uu/jcqRca
7hu3348HDdy8vQxHKJ/2WUSv5mrJ4MAsIQKhGBqHRJALSiJIg6OTkUNm7HCSfTtOasvkNE5i6aNB
xaloND73PS8us2BNaywSyfl5WT37Q88mb+hN+0wr8lVHnF9QtyPw6sXeF7UevGAyOJLCIued/f5O
A2WNPhEsEt6Ptm6ckHs/kHwGHAzLc1aRAk7InJMZDmXFaQIqIDD/WVnsqP36xdC7arO3+0NJht6+
WvKfeC4Vo5AffYogNi0zYExKdHdFlQ4pxQl/B74Iaj1cvDNMIYK53z7eOnYNU1LGHYJqK8ankBCl
Bm01v42N+Qg/S0hJwPzdWZA4ASW6JdFWf2ruZ612xe/BNSZFAjhLgDiSV+iaBDtgbEeDTC7UeAJf
CdRW6e/WcgsTMyH4A8U/VjmZdEGdF0vPJCj97sG4rmHko8zgMu9ieQNOKm+yryxlWeyTegkXfubu
0XDafNN3W3L0FE4Y7rnAZo3yEqsl6egKNwbbXQKOuEU4/y3SPTR+0pWDVVy+s/kOjcni1zvTgYA7
Cht4TspOIWe9/3LTFLAH5TSxyvTV6dzMRxyowBK23o+DXcF8zPj5yOwfNwTWLPP5rNET18fulzkX
a9U8IyqDyXEwTDNAkPk6qYsPmRXAIzTVQ/9WvFRmLkcNPG1Kk8Dn2Ngg9BP+cvu6JxUbvq1qbthI
O1ZN4y8ed635g9DBEgCxTrrpkCGiFYqevbeMXrIMEUUw1NIsTIm+abCvr9ksfkibcec7nCuJz/Yc
VFTG/6lAx2rjBn0en7Rm1MAGG2Q83k04vmIg/ZqeJurmQv/cWNIHoJsd2ET+nHyurAVlKzBtI+oU
DDXLu/YF+Q7aBudmWwzfMK4AONPyAXtkZR/Y3jh7jXJK2FIukc7eoNDI9bdoGB7JLhJqqtRPwxbX
t0oB8Kq4KDgGsIF91j7bqpCQxMQ6DQUHaHUjBGl6QxkSGl8BwynSohUeKrHXEeH3vj7OgrvJG+TK
ap5i2nOi91GsgtqS/uX6O2qQW/kahymP/q9j7bHeqV98aNfMitkAj1RxaXtfh7Bqi7UPET8yCpUN
+pBgxcOTaAYimL7SoaupM8ke08C32RNTSO5yEuHkd45Nej2IwPQ5XMOjjhhXbMwejrgaeAD+ol/i
3TS2MJPZYvZ2BRy/NU+eAmo4MvBRc8mn1sPOgmuJClndxihjTMERpO/3C16KvULT1R9Fzl3boptr
G5d6BunL+VcZa2UTuBgfTyTuWK6NdovgtkjOQ0ljt7nQsFpeJgqk+fwTzVvlTsfBqFrZIpv78dI/
B+/fVyZY8VrCn7jOTqxvQspo8xgHqE3VuTVLs1NcyppQtul5iFU3BFy6Oa2GhapRz4Rup1+RSFbW
Z0pCQKch5T7wEfRTpo1Lj/9Xnd5ZvWXYOGez4FqLgIeZvAuQ9cBBddI4uWA7uc4FM3acj6o7BMPh
pGMYJltmGuYFvxjLUBL1pCu5nxol2eazAewyUY1OlGf65Es0DmIFY7+xxfpcDi3u7XjEafF9G2tM
TdRU0z0rddaiv9fZOqNcer2B7laihOSdBRtsJSCRywrmcvE6mulVz7/hJjd/GbHChOag9rdMDMGk
/roKgEN7VU1LLzUCDoB8ctwmE/P+k6eslahAQKsfDjPM+4IwfUEPa/DBY7+8VeNErQpsNQmlqLpD
lFqpTp0zapr4jgAHLZE+39SzlgnzK2YuwGenJv9rLQzZnbscsgu0DBoa7Kchwr9ab7FrjfabBExt
aewFaJ2xKlynPRpNStRMHPAspnANhaH2QUJDiB9xTGMpvOzBJUyKOINCE87Os2p6dC4K5k76cGE7
IDUA/haIuhVZwg7dYXQu7NXbaAIFwk4DbhQZqJ4jmPQD7osQ/Vc2XK7UOO1rtApUQVI6Zj3GACEs
EMXwQ8k3rOxXROuM6ABHGmOC3+Dj5OOxFpX5YBgeWKnCHkMbtsG7Ez+dWz7niUv0nz7LCB2vAxXF
ug77haiDLfiYSsb0iTra8bOU9zoyu7AD7JxTwgHWoVaDHmA2e/u4rlqE9odS7PWg0M8x68NKsRc3
a9V/rXGwfZXGRtzJuruD+T+YNITOABrbW7uJVF2iKCsKM1baMFJ3Ulpd2lUuItMQszgkUYDpJ+OE
jpQN72GLGQXrYVmt0IL3tWbGuH57zjt0+3cfifntfNZLDGZx7iTASNy0W8oxOh0y9Yr1qG7Vb/RI
ut8zEhVOYkUK65x76kzGDfdCmv3JeXz21OhJGcB+kOKqHhX74/UF45KaeoKsxoV6Q+pBBH+srqXn
StR3rZjUXwPf/k25vYacWcnzY1ICzS2OH9KZenOXnd/wEteUfmdTUuXHZ9/Zu7iJtxcCGLFZbj7l
AM3eewKI01PQmjkYUU6BZBN0CTZBsBvFb7FsIN5blpJ4Wt7j668IPmklxOPmqeWJmkXZuUKH9t2Z
nRS4DqRERvb3DMPLSS5FhavJfbgK55UuHuSXvh/oysmj5xn3VMtT2nn1DIHgBm7Fk/89fFI2wD64
vTq+PdCcjyO0OWbBLcJExE6TsGbhzLOkWQ/IEzcTVHnQD6ZmEXM3mEPClEWA9wHHkYtl9ZB6AoaL
sdJuijmIt8wqXEK3yh/N/hNRg8G8fy3isX+ksEQ/Nb8MiREmaa2vHOdvm1Elaph5/EbDmT2sFu4B
2LqDm9G5V4wrdr56qApiiPoRcfrFjYiVR4/IdjDtTfdQFhe4lI6XdjlddCQmZiUIz8LLwZqoJeRy
AmbptP/mkTqitPRGIFDuPA==
`protect end_protected
