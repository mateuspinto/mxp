`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
CZQmuUxiEVTNl+nnbPo6e24dxGTQWReGynZWWZLBNmf66eOgnb/J/pDVc2yp5iUq97xPOfJBTe6x
627nKec3JEp3osn8n8z0R8H5ziQnOea6/UlkjsJWqfdTUMHuYTH/ZApQLkscP6Xl/caacSQyJAcB
uecfdQPnyCj2Yh1AULqHXlCrfMtItYFuHenuqnn5yP32bYL69UzAQY06HynPJa2NiCrdMptJDNHu
cqk58ppN3lqkq6JsQBMz+XrHgC3d5B5JBahmsyg6EfkSCcrPaM7ryPM0cV5PucqgJ2nY/ibv9XxQ
OtcBUGsKDCYae5uOus2F1krmJB8lfnIdpR51FA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="XoQU8PXZz0qBGpJytnLy4DYTRyp4Cjak6RAxUQvtK/U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
UdONN2pFGmKq9GT1ZcDz9aNh3QIcItjCY6xh3/GfunkwFHmPcGst2Fs8a7KsMrfzkbbd9ckmdYMe
4yVZ0+AJSZ47kj8BDW5UD7tQsiLkS6Ho//Ar0EVIuFSqWJzjAfbpS83YXutSaOZc3ho3mR+SO7Au
m7E6QTtBduJn9ApsYBvEDqXLFaHhwCbMczVvjX500a1eyOg8F7a/0o4P1ufc2qlLjHoMc8GzrGXE
D8C/abNFG3P2CZ805K33oXGTAX+yy60mrl3xsrKhDkYfab7ojuN6lsXlWOONMnIpsDcFMtIccHK+
fs+fOBx2PpOswtPHVPD9BPTDaTjO2DuyJihyuvU5xYskLCbK9gW5y2QYAwbnZMj9nlWaqiL6eNKz
rNm3MpdqIlMCfap90HgVU28f5g3AaDZSa5JbZd23Lm2I6byWFI3MOM+S1lI0RiCeLwK72T/PwcUE
wdpnxHkejVFldLhFmz50MaKBqsRhz+nWJ9vqFfOJmYTI3/cS/3geDgTp/wRy24fHWaLmBAT8HyNE
wqerhRsbIlvb5mldwI4iOALBZ2hyylPy1nWZTMPv0Pp7fyI7/cwM8Ezp0tsx1lcR2h9dQXNxznql
ASDM/UM5WLoo5b71Xyvjx358tNKekRMRIZrCshC0QJTyB7jFk+CelJE0+CbRtbUY3nEIVp7DkbgE
KhfbQml/PG3vtaXJzUSsHqyitIfHJrUNxOQEGwRhR3FqYWSwQbNs+PAriFT/OUrw/myal2vbeOqW
6qjRCkq+6nSg1sl3UcSch6rHc9ErsHt/OQUsze66qer2sCeVzjxKQzrUlZtR3idhmI9SRvwPbrxu
4L1TtVAShEWZ+N5G+1gsity6oixpVy81J07qruPXVWkOEuiHXeLWyufKOdCbwSNwVY8m8BTSI1od
kbt5RZOv+VRmWvte9jda0xiIo5jE5g3Pc6crBoGowdStmrKwakf36Ep6ntieLulN3dfLCp9t4pzL
X96+3GEpWnxbOYNDy8ho5g7yzUv4RqNljTzxLFsFZPAGDTBGxqm+1BxDSwDw0SFJ2QVgZwJizWjb
w85PMkX+cREazEQDo4n7Uc3ToIy8fvHta4fMYteqSxIgUyqWP+zL/CaWmvvo6D0wyB6d2C7XzTRV
BJhMhG5LBKNPFg14wBpOhgZN7e4KjgXPDj19Wl3IO5sBv8GBc7fO5C7pMYH9iYR0fLasd8K6RKeU
0gNalEBjLZzhL2QwlsQ5CujN99npo2nYSjXKDCbsE29h+xXa5OKCx+vMAJS3GZiTqD16LOz/10Gq
y/xVO6YryJ7wOm/Txb57/JTwwfq2LVzPGJA4nm5wlN1b+5J3lqTMNRFD5zpIJIMY1Lg1Lam7L+9B
aorZ6xdId5EI60AOddz3V7xVYtEgXDVJEhWehMJ6IYQfgSH4apIoInqS/9LXnaGtgRYT2+Nzj1pR
nc9+zU9U31OdHh/O2rDVTtNHDcAlmiKJdPR+2vaUzbaC1mgVgstf5td6NJ5HGz2s5AQImSd+4bG3
BvzF3Y3302zCABDZ26GZw29k2+Lr7NviK/aQXsjYBICVKqUxKoYF1DJc7SFhwZPaqzhp6EPNicuV
TnNeq/6LAkCYPOfdne5waUMGd3yqXIqLcEFeEQztHrKU1T1s8aiJOZltrafXYkhxfbikpMHcuXZ1
Dc98MaedE9lIe7eghtP70iorltp3hRn004t9fHHh3GEIbapWhd9MQ/kr/K+dx7DPMHa/SHtpoOHt
7Z42cvkubNd8duLWxNXhurhJ47McAHscL8yCypt1ZrOZpP4KB9n5k903+irzwJ4yjjKlQ7m84rrK
tR+E0Ew5qW2ohpIohZ4itI0gUbBWU01nTuEntck7j+4F85xAItk50fWeASTNRSBhqgggcMwg7MMJ
ZJvDqH9urPRZ+Kts2CdAZz/rX9kKHqRLOZr3j5jlX6GMOyRU9ec73cribKzDVEOAfNQWSEWbJhVY
MuCVqZ/cOz8oULrXcQ5HANoVfBMHqN+5IafWeZjv4bFj5P69VzMJuPBP2aFwzmspWHzo/ckrTypa
mr7ty0FCznQPetgfnmdvGFbk67O1zwjLwMbUM7zWCEXQwTOXb3MWp/1jaG9GAB3DKgLZSuXWj3xi
d39SzJYGjxC2/I0IG3aSSYhAods/nTFxbSRFJM8YVdCRlBsELfLVOGAQHLM59qojB+V/NExb2IQi
Z+nyBvaxGAps3rFgrCO771cujSb3INEuva8D7q0tK5r3OMwG4P6IMFQz0+g5X9qccVu9DIcCidka
rHCfcqBpYcP3doLCa4boaEq1Yijr1M65O1Atxmbu6oHUBbog9DGiLgfjjRlOssUJECe8A9kRqI/t
A6jTPSn1g/bD6BBVxjtUOoAcqok6qXw+uDRsbmNAV+hOfvqQyQa7KA8gBJQMfmzNZw4oRhTBKxDe
7SylOWDw2IdKIjSTwQ5jzBnKYt81+2I783DP6KzVEUKA7ypfDywu4xynxgfGbqVpn7L5KC6PMsqI
N8TVYUA3aMRFkGF0YCTrBZKlTuz5IKEZaIzO/TLLZWtvi4PoTkaSNhrpgEyRBMrbOAyOwkZKLhr5
WtJ5wDhF+mctD7qWPop9socWWNXVs41RfxP/UyVpC1HR5t4tf9lFukdFLNtt1dZiym58svVlkoEx
9lKmZ5ZYlu5fjDD3bJbskzLJoyOY1urrKujgOKEDTVYeASkZkkNpXGU9CM9d8fbKJVB2B2qWT4yX
2iC/VucOMcQGJV0wV753iTm5fO9hSHRAQnTgoITRqTIgSMkfxw2AwvJBvRGwBQcDFi4nZoejfuRL
iqkRUHdUYMwM9W7+6Cm36Y13ZkABYAASKxLd4hA4mrVyYh/lCs6A21sIBHr6O+qVi8D0JpsFlMBb
cvBdHGuyV6qhkaaUFJfjrbDXjlfEWq3SDbmYRHi8IVX1pHJtxj3xd0Vsyyh0069GQplEjNyldpaQ
8X+dEqgeRArOLNiDlBV1lpWDHpCYVykxKuhjt9GDFgm4Uo01qNxSm3QzCPt3n6yAID+usaZwwuvn
oUotW+g6OL8VYuIxx1H44UJ+0qPxGdJqhHjHp2blbfbw8Vralz73XiJbjD5J/O/vQcBN6kteAchV
8VlSMEhXFJp77qYeVCN/zgWerq3kE1Lk0xZq38oT6A==
`protect end_protected
