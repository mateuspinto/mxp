XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V�gH𚯾) �{�;H"l �%����ꑱ�㝯�#e��K���c)�bc�Z���nE��Y�M"�Q����S+��u�$p�<��jR�Ý[>*��%z�Z��/'j�ġR
��n�o��s�:R�B�L޸cyR�ݦ�z���җ�������C�X���������'uf4�7��T%͌5�4�����uUyʃU���|�K�]'�;5P��*Fe������u��Q�_"��)H�qԹl�u���uh�nCjh~_��]�Aq�nA�n�?�M(ɮj��!z{]5�ѿMh�v����q���:��b/�h���!OD*�$+|�4��Ή�K�� �ٱ%���j��g�6�Q��n��V�"T�l����ʀ�_T�o�Cݏ�g�����֭��������N-A����hB$p����&s���\��JFv�kb���6���?;��Yφͱ_�>��=�_(ِ?^Y���΋������]��;�����І�ѻe��袩�S/x`wZK!"�ªU������x���f&���j<mxp�C�;xÎq�l�T�X����
J�Y���i�
����Wh��I<a�y�A��j	I\\zx�2t��E$F<#��Ѫ���V�\�zr���H���2��|u����8�3�L8�ה�"L�1���LE $}�kI]�ڻ嗑9�V_rxe������vzc������Q�T� Z��(|�R]%74w��U-j҂N����l.�C��q�XlxVHYEB     400     1a0;�O��$c��wC��k���q��'G,&)d&,�E��9Q�+W��������װ�Y .Tk�V��P�}�U�`���]�y��L�.�R�.��0��8.�̕w��ZHdiV�mz�q��y+���v�.P;4l1��5
���4ָ��wl_f�s��EPa8�?�TNl�7��\_$\���M�9�-
��j�oI0,��iA�"G�U;A���U��w��4!�1�&ŗJ+5^����04 T�� �FE�H4�>�ySJBa��ן����R�S�o����ԉ=�_�?�d4,^=�����Y[��ˈ��BB���훾rL��J	��S����	A�?���x�	�c��:�<k6u^Lj��u�'R�\73/��Wd���Xz����cKB��J�2�(��u��i,�� ��stXlxVHYEB     400     150 dل��z,b ��[:t��v�)'لZ�����b0�@k܍���.�_&�2�u���}p2�na��{��4(GsY~�]\ ��j�U�$�U���~�m��_�����j�A��Q9�� ���iqp�ӊ�����׈���>iz��qC{us:�c���Z4��j`Xτ���U�^��e,-�/�@�AY��>���?P��1n�J���$E�X�Vk�{��Ӥ�|��3� gLRG�3�.�f�+���O� !��_Ѡ2�+x��<Q��H�=�|H�)wxGI�;	Cg�LP��V�ǈ���g'9�_=��<���\WXlxVHYEB     400     190Z7k6Hx��"�����A�|�+���5�1��<�pJ��Flh�I�� �Zd���<�&`��w�8@�;�^0Gw-_YW'��ћLB��u����*�oQ͍ ��D��[�Ѥ����/�1�XY�a>�0k]�U�4�-B��������ؐ���髗� ��5s(�$���i&���{ݟ.֜�UO5*R���(��Q���u0�B�B�-x�
��#��/2i�{&����ËW�P��a}��>O��^#�d����#���FfZ�+I(��LʏOm�0�@B�����H���Q��B}X��dݬ6�U�4)C����T��ig�����	'k�C�0V)�!�x�Z�dr��KbN*w1 ���^�.��Qά/�c�*�>�Bf��*��=tˮ'XlxVHYEB     400      f0}o'��UJb���T��^�r�"�Ŏd��W�C��췠8m��+$+��b�C���
�$=υ�&�V<���h��Il�5�/��<'`
&۟�l�:jc'�V=��k'B�������*b��c��.�KQe�S���a_��]_f���^|o���|ˏ�\�Xt����&�㒜Ϸ�^rM���Ԗ.����h���ZCxF|��k,!��7�ᘕ5H�qa;Í�$�#�,��ec�TXlxVHYEB     400     120�7Z/�dhbKv�ze�]ʍ'�rvw�#�q>7Wg��S__�'�����O�4�G�� �P�dj��)�=�%��5���"����.K^6w�s�4�6��1%���o�ܽ�p�E���<{��񦍴�m�E��$h��i#�hk�L#���s/���\�����D"�@O�6mb̓����n��A�מUW̍~����1�A�L-Ng����x=dx���,�,���4޶���A��T�5d��hٜ��^q6\��S�$���/Ef��P����g������H�XlxVHYEB     400     150���#�}q@�Z�O\��t l�v	��P���Ɂ�U�5&��5�ux�*\,�?4o���]��'��0L�f�Y�q�
�O8RC%T&�q֤��j��-���$�ؖ0$�GI��U��`$�ϋB�����ԹH�����ώ���PE�J�6ل�A��1���*�S���ER0r��]gSG?�(�������fu2��ԅ�~K�8���q�z�|yl��~�}��8����m^RI_�Y�(B!�2#x��DkL�S@�0&p3 3h����:�d�r�%�����#߫�Lt������𘣛�;"�O"7�9\e�5J�+�2\?E�4�f<���v���&)'JXlxVHYEB      ee      70�sIؾ8�I��5wҫ��������#�ҭv� 8{]��a}��*��������g1�S�t|?�|�ݢz�<E�{���6U��Oy��6��
�*Ъ��ʸ[��  ��{�W