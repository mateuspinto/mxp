`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49312)
`protect data_block
0USWSUGxovGsyBJteYpEoZ2WVliAMUPKxPEpzQ45dt0t+cFshbb/mg0GxwMi9Ec0HmPJeWVt5tQZ
vTDRwdPzb0QxrXeVjxweZoj6TLyGhFlLGwiFUlGYg0L0t4wZ/M4Om4hNkxu+eoZifwOf2cHTbbko
zkXDqmhK4vYLbRnhRyHa7NsMulu1sSsw1svCmELKqbwkcattdFaRGyGg/lGNKx+QV3JhvToSIEGv
7vAj04/0tNkT4H0YmInSNsA2YRpy3Y+PlvLC9Lxpba7qCH6rnKbq+Sxh1GAa1q8U06+ccHFRmO4N
xQES2VwI683Yz4VbWFq3iVzOVuOxKMqA98tkMlX2CtILpLX21rOhf2rqjYOWPCd1TcQLReqU6q3B
e4TE+syo4ACfnfdgCLVTkNQehgMGfgZ8JKxtsn8zG3/Wiq/ODQ2q3Tmt1QCjz2bKZa1/FQC/VRmP
Y59z6idQuE5ona1Y/UHJ6ios4CTD5eLRQZWpTCCP8JvlpznQzsUkDEAoQioIK+ZD7Q51fVMQFrXT
0BcY5rmPd/E3w+SZ88y3s7P7mCE1KiN7P44ntDrtN3N47ZQ9WfJupPIY0eM4rZL90SNwxBEsJK3D
/JNsdSoN1dQisvfo1itvTs7yrUwk0VyIHHN4yo5slGOg6mc78Lp8GhmYqXMxi0IBcnEIV4Se2dwa
xC/N025Ir0tqwhL6UUqDBw/3WQALOkjIvcN4aVumaF1w9Qbv9OHPgdy7aUk9k3DPrM6B7s8d6PFk
3gQLSy0h8172ubV00uDGAYgK0N2FfJk5JNx4MN4feQFG0CKf6fbzyA6peDQNL77tXGWZGd4o7DlZ
btl42WVBljG9ACi31uIeRKMnvIh2TQF/8hekFbOOi3g8DJ63hZmpM3Qq5Yc9c95gBIdOmr0YYiRk
auk+K9QdAhkGvoNvvN8nSszUVTaGL5XYpvhAirGqGGWJJxdtMrBoRRcH3iojwIRePfuI059TvXzb
Fr9ayOKAUBzCDEoIYrzeG6Nal9ysQyizgXC0Hxk3HP1XldyKT0zskWdbLI+X0hwjLsyoTMN4rWjQ
hGfc0ItCNqm5or9u+rXNsYk5I7WYvKs40VBT2BopboBNJwGxG9wXElTf/2Qijt+CFgHOK9V8AWOl
tk+hZUZ4HQQhN3vgXuhuWWdup15f+bnFB0S73egVbhS9Iz0S492fgTRu44hX8TlTqj7jDIgdZ5JV
6+JM+rs4BgJDWNeFFzSU17ZF5qaH44nJHEM3OB/2SEzrzNI0/ToUWJcZ1vUiqFtPvMDVnCXHHuDr
WId3uUTZOF74ctBc0u2Dg/6HqDecddxxLPNVG9QxK7RSGfKS4s0GXBUYJR9WyPNMIS8BrbgC7+rD
8e8AoVg05d3RKzcUfrgei+bjAVlkoBEJfhlcsuxiMxpa4OyhD+rzgJAeO8ng74I5iGH9rax834gC
Pu1iBijMYAUz1KRd+l5lEjOcgyIgzyhOcsfy8LOiQFEkJOa4BzeMMQnIfIe3Y01dyJTkETpXa/KI
d7clreLq+xe/VVnZfFUvgtkxPx1et6Xj3akvgflU9+LTeQpW8rekiQHvFvkSHPWR+SAx0KSBDIr0
PzoAmN1x4QKUD3T0omxoRYN5PDLHwpEMPnSrk/8c5+gD3UI1S5lzT1M4SqzSszN6CTS4Pzo1doal
DDscYBjGniXN+FpoqIzFODbY1Y6zeR5N7EJOdl/XvuG+rzW+IuqSopS49xQ+v2orKsVps/iUr6gy
XFyCDRrNGvwmhQKZp0vtev7JP1ES4OQQbzyE8g72bgJqKS0svbuizqYEoG6KrzXYj5cN0pt2gn1U
J3phlDIcBsx3Rhdcinhihu5YDt4u/8Ug2P6za/WNyhlUNXIXQKzdG7x76JciwoysUhja28iYMFTB
L++ljX3I1QdLkI6jGqgVPmuU0Ra7E+9zljvso/LAmb1usB/rII2ZOedrzSSAmvsJt3b7vft+cRVv
l6l3gl2CZ6uGRwEHMIZ/XwEVcEhd2etMMOMq0oSkW2UiKuWeAyBhpJSd57z1gQ/Y6FdOMnYVa4jJ
YURbX6XEpX4HO1hKvTzpNTrsFuX6ulSVXy4k3ubOBzmaPG/TlFViZFZkLc88ikZzqb5Pfy/vZIEH
w0nnKebLdtublYY12uDJLaxNloDDBd9rLOyf+fTbkeUA0Byh/iZ5NtzzZ6HA5rQMDcYKlM/odB2+
XbNPVt+Np7Jce6c9Z5b+tKb75DNcMk9cR9fSYu8HQwd309hxzROdQXvO7z40rhtvZwCau1Pp66Wt
HMZXxwXLdfDaQ5356/Qw/jfgy4dgikmXJ9aVPIMG7sxzAhgEZCpNP4vGGyWShUI+XJcBO9jWu2AQ
6grqhmlI3leX2MoFD5S6caHdn75sk0O749+M7clp80fdUP/DfblLCSMw0zdcbRPyWEWrlKfOWkzn
5MMP8C+C3u0XHOOTuHpK3T+dwcQOdlV3coy1O/YtY+bfEUroju2C9NV9lt0ar1UwmITmhKhcbDmc
nfvb+mXMQ2+Y96WMJ0NkeAV4SaH18xVGsW7inL8o9wdZLiMWXRquH3bQrrVoCCY1zpkFwJoSTR4X
aWm0jyCGOD0bVcMGjIHtaM4AQvTXvW65p1cMYaDPXkyZelhOc8tpi4uIvkejWfm/zzDDaO8wm8RQ
Vdz2WFKp50evvRyY4x5VaxjKB1g6Wjycgj39HGu3tHIoc/G4qfiWuSd6q8rUSLKpDmMsROYi8viJ
IZ5wLIaJGmtDoJ18I3i0Vrx679WbFON8WoadOhhGB3jvTMeeNQ0Phjdy7GyQ6MjnAQ4g5zH3EWye
0Uw3IBSptDm5qoxLI4WVpc5+ol9799XwHKY4ZQYDkGD2iycJzaJ1Hxr7OSPpmEC7OEjFeDbfrUAT
eOCKlSvRQ1TgOOhMqzT8HISso24w9gk6g3o3ALiWC0x7JEzG7LA1DBUQxxntCDpRNd7ATetJe6xC
hkPZjk0zcLllmTRltiHNCdlteG8GBtSGzg34ZdZQSTrPRoVLOTPpNMeswQZ1yqt6Yer6BFeMDr79
HSpfr1rFlGBrRmZzfO9AfBwlHWzc88S0b71XAd6noWobbxdjCN9QkwB5aAxG8OtRO6f4iE9WK7Eo
KBqwZoa4tJcZd79mHlG2oBfR1ppHnU4dd2bHsLKndpgRYYthLmmMTDKTvI1o9/paB3m8/j0x8BV9
soWTkmHV0Bcjw6USEhkVyM/A0Kkn5eKd+b3RjukdRfcgNoIMlRFCxPu9NRR8dAiA9FkXmR+UkyYk
FR+2V8nmert2CBvWMOWHXIxXMLDeNz+n3ilzcwNfag7CNup/lZ60KTPQISjTyO/HVRp45josY6lh
o4HiHVSYf6OIUYyy+p/oyO4aqNdVlxp4OZ4lQlTU0iSdCqj96j6RPlT1tjmzwFw8xC1jIimSGAW+
6Vp6/Df69dKqzvRG2tUfkc1ls62Br4iV4zTZlqMPXbxKX898uPJrHJFM4ft4OJtUXGFyd5xDGBLi
nJAdu5uIijhRT7fnN1EkC+E6SXjyT3wbmYuGzHTCB1F2yC8IKChrfrYxC5hWFHcUcldmFtXXTTSM
oWgwhzyEPLkerdXqIEEue6I+Opp1yGuC+6r8Es4i2giDnwK+0X7NPlbULxmJJMNrdDvFp6mqBuk0
HEd1eWC6NYbKmBcM27tfm2TpGZWpdXXDtrZ4RZhEt0MXWUeA9HzcQ2zil0AV8mdRGtTgCWQehkru
wgB18yaSDDVTZ3M1yIgecTex9u7MR6MAmlj9DdnZeKuoOiwBxPG7gwdlwR3gZHZ4NVbEfSLs18Bt
/Gdy1+pWsWtFeioXS0vQTPHGbdicada3Xc6X6JoZ91QzNyFDiIEG8IAfLNeLraHTEiMTiErvK8sy
GVA9mZTY0WKa/p9/0/Ip/AerfmlzQx36+j3U23LZOBEAtbvBwah2LHOCES7VY+4NAUrMfV8kPniz
lGG6nE2Nbzuw5Z1MfcUpCR9sRXbUQ15lXRVF60BAUsXlt+bnaPTAubsOEKywBMuu3urVdUhqzymZ
brBW7UFXsRpohcI1CD6wW+r5NDr/zVwyS0VWzbXuUhEcx4cSxbZAFnURj+cB5BPma9jth67F1a26
8PTH6LBz4pClY/ZDc195bo1DNYXRapizz5+v+vKUzfo8gq5H4Bm0NrvsW3YpOLU7H3qBO52UPUiF
DBqxfWP/eIG9gcKWARiJdGx+J+T4kYFFGONTpfcDD2tYciUo78pCgQlAdqIH63UJYiMoZhCt5fXl
u0w30p1s82RLCjkItsLRkZFu+aDVc+VAXN3xdbfjl9LwbY7jMBPo30ap3WIShNLOkeYwJMyaMTGZ
3561KB83g11tIb52ZOMtcfTYsWDPF65mVV1vRqaKAs+viq9g5lWoODvSOLL4Cz60rsPw+59U+G4T
gCZaw3MjCMtsJWU5N2sHHLSpRY1iOrZSZAtoCI/CA46ywKm7hGFYJipchFizlguVFA0L+jVq8zM+
640te6mzf5Hvwwheg8qY1VFXfVhZU0XBTJHgJtGPlv1sDtgXueVUulgv8/UIe8Vek4bmFtbGHZTp
7t/+2LR6sFw0fCTrrWIc1y6tDvD2IKIoUClpkdX8ASGozB7/wiNJEDEUi3PYBV/3wE1sFxINPOzH
nLwW04tcNYi82/5BLVBv2YD6nXuIkN+fK8mv+VFuuinGXR0NO7STUSFSCpUhsMeM6MhltFh+zlhi
HuHFX3kW4MhEUu9N7NCOeMVRVaLg32+p8mKdit99XFfBQTIjCfaGL8N35vrEUd47TlRoHSiSouRG
PqT27q1gkCkFBATnIXrmCLVtj9bP0WZJvldt/cbBwrGE/6ZMbq9KQjIwzPLoQT1HJDcmWcm5fPNM
EHIp53TIp4NJzqd4JbUDljZdZugeLDcLltwFgNWHIY0IxhWVe0IuBqv8TXPyEeoxZ47hswN1n5A3
KzJbKl8FD2hknThy9F2I8T9ixdy5klE2vz9UHwWnpWMlJs1NCnH1gMLSPC8383kbXSB3ksAkuxTC
oU+bFb1E8Y9T1l3oGjhfjSEs7GuSHhZpQWGqzVgwJG8BnHmfUndey4tWqxNIqwCK0xAgW8jNsU0q
md7BNXioUwEdKYHhDPZI1YwM4lglpvT2MgJBWY290nTrvNL1shypinPptM14vD409wP46jT36mH6
/GKnsSoJ+IPbWP+L4BqECvhiUsJ56CKvWUrMDJTWgoT82GWLTNQ5PB0QfndMltytyRO/it+GwG1P
PnDFqYqfK3LGkyfzunvIaPC5h69vCvc25NG4imNPYGORTP+FFG1psSMZfjFHd2hAgVTr+JqIvwxN
3h3Tp+WU4HdiJCwjdGu86QFbmeXTWobI5mPihhkOeUwp4T2vD4a7wapnN2JvOYtA7RAHi6FILC66
IkyGdDk3yYszdh4LWyJ3FnOYq3U36SD9Uyvm/7Snrd9u64Ajsz/gS4hTHd+dsw/fox4FeKflf2BB
o/YyaWC94py7pgREP05ofPb7jWVyhprvpOaRwv4eA9kv7w9HS8b95PuC8zfourmInCHOFDw39DYj
KMyHILlW32SRf2jDLf/11g4R8az/3LbcaNJTl+/Th7gfVYJSCNloa1IWDKOgDRrAr7Xea4RiCZAE
HzDO0r+FbbO8MwB+QjfIsMjfV0sKi+dy7No5VZelwSBaAf4eCyhUep0X8+HNJVA436fUvr3Qki/g
DsH1VMDnaOkFDcbBW/53BopsSd1LePKPiVwWeU686pgXgVH+/ic1I63SKq9WIGhRtYpFDPnZy3al
WqetHKg0jqs45KMyaaM3VEYEsdUi/TTFLuHzHwq/KbCm87hjGdz343rh6SWPcYLLhVdSJBkJ/i+x
9KqkYuRGRdpD9NinbbNRZJ5/laoZZLsXmEuz31Ao+Lh62U5s4DOtLrgPaKrc1YFrqBaqH2uvYAML
+ec7mX72je2U/eVPbXjghGWs+IFXxww4sJ8Edu3fM2L8L8QjozmNaIrrLrOoulF5ga8DqCQ5bJwg
4aMQEDP2Pysko+ILCUNWtNPk7qhM7lFXpZgfUNcNVvOyLcHZpvhe3HUIfBq88dkdd+sYo2S7pE8M
PrMgG+9qteZa+UwcDH5geuVwuImrYPFIYqWzQRrIMCTMXsUiq7NOAAost4QPPnCDJ47HHwvzImXl
j9dH20fynwc+mhDJsb5z+R4X56NvZu301NmfrMR3Cu3KMvqCBY5qLU1cXvzWXcakqnp29XvG+Rpi
s69gu61mcXwFdxKyyxoIHpPGVBASsKa4O5VZ1o76QvhUr3cdy73iFhj9iXdl+HUI8GdC08/sfwdn
oI4HQddJT0WNiwms0e2xeO28mot0T9ER/lcfl+JQRhMYZ1nbBEEDb6IdxWZSgknWusPBY1fz83tw
J8qtBPFozdrRAJNmWzVl8Cknl9lICdVEMYP3Hu5BujRKcozodAmHVK3eIp4L42bcZNTXfLreSTxY
MpMGDfUIqxHN7ueWzKKkJKoTZLMfYkLTe1IrLiVqeP2CPP2Dvinp4PHGXyl5YvgZLkKGvHoRpxiF
ny5w93VJlpe218agnDoRBRlEE0+hfd5CybHkY9Sia38I1/ttNf+KL0/A5v07O2M6ANUVvQ0Ecle2
ii/y1SCJtmv/Y4eMBLObSmVRYniDcZsKoGvVkWkGhZV/bLpOE7+IyVrZQkTT3Fs7sfMV8Nk6sIkb
LTTLgR/QzSMbRy+JoMErRLjU/Vvy8Pq7CCKgSwzqsNSb4t5H77YUpFdBk9QJdN6BJagVZAk+laOG
l/dOREliScjCPSf8c8x+SDgwiWktvLkG4Zjn7cwtXFWktGCjC0T+MhOBwnMLZdbGFp7FsSfsMBZB
AGC3AQ2VyD77rSs+yuz8t9YvpcNnNn0qnX+lW2GrEG6MOlZYNjqHB18i7BiYc5bBwvHUO8hxYSHv
F2lf0BLg2sziKqW4KAYFs8csfjlER8f822Is0M/p25aZYRBK8+VUbEW479SK0V+a04kcf6BZ87Bq
5JSzWjO4eyzAakIobEgmTKn7kVTbNLpXtaQvrjXqWbQVkUpqihXeUZi0ICkSJeOSUQOafRcDst49
BMtCdvo0GWvrRJ578+6KzjSYYNQlX5IUu3F6tr8dlS1gKkjLVIxMzphJM65kYDzfDJ4FoAi5pf30
IQVkPqxwC3uqT8LW+vYay6EeTCklPe8lSIMPAj0Vh7LSobuz1YfV93n8SdPWWAqEUHKAgspqXK8a
j58M1NdQjGyV//bwZEt74DMaMG9NttVgOmRzbX4rXV4TF6oDeWiDqt4wq2uniPs1Fh/9VPZ+IF4c
KcdxX6wvUcFzDuW9MBqn+Jgqcze3F3rtEKwQSsh/2T8MBCxH307AVsGXxXh3jhHq6SAG9ks51rSM
OrmO6youYgnqx5wZXbE1qgQ9tqux+O4E56TuCwizXBkLtD3bbxW99FABr42roj+lbuwkCfUbGMW4
MlY2wlNWJ731smIneBuNdeizQ/f7gjF1ahnMhjqeSXEVLEQ1aaN2qo3kHVXVtxl4SMo4AJL9bPlm
/MnBeZkHoH7xd8OTZ4ok7IEJz1hONLLX2OoCPr+yfdtLE1MvPbtWz7Jz64Cwd2s1z0Ohsp7hIhlT
wtVPyIuh1m24/F2QVOH1heT6VK3wJvznR7u5+xgYN8SRoJ0nqye8jwYKekJfl2BjzmZc706Egw/U
VD1xN5l2NtUQjIGjTbAZOBJJjR9X6NmFzH4iy3RfMCK0KQsX8vdj22wjjUVAzt0PnYudSJHupGDi
o3+pQMO78xTGYc+YgAh7ADW4b3+YvjR1Z7+X25a4o1nNcMkplYE55C/uzeVDmyFfrNzvNWmnjnyn
GBdTwWbMg3lQfznZxxLA8+fiauDacm2OZmF4xXJR+cuOJrxL0DvcrTXjjJmLQEhx4OvJoDKMvnGa
akGbeZialGOC+2Wsyik/qSgytOb81KC1MFL0WdqrcXE1EzM0AYgSudQ5X+EGQi9uYA7zrqK3iHWx
xS+TLn9BShLAi6uDLMg4iijbpOe2rGrAWZAoMEqIIfPNl4r2X5ZtGEwIowHZ2m4qjOlCENlGt2T1
pYwPENA35CQjGhL1SDww7ke3prYPgN3dVEUlT/NHVyneI0JIo/XsSUf8WGh4YSqdRXVNhGnNZEro
pYHShha7l0AEfBVokU7e8XFHGdFWbw24V9fFstJHjlQMmZNkrV4LmfQ7FzOMylexHfk/efvn3rn9
EH5B7YwvmrqslVDTAXEVmpuZPI/znmc2ufp9qkxF2mxTTs2QSssHhf/Oy0SwvXVGmFNxpSC3dofF
PNjSunK62VfjpwaTAgT2sw9zsJXmo0M4E+FYwPpz8aPwrbxR5BoE11yezBXe4+G7aXjS2tiG1usO
izh/Hobw7cfNQHa6KvvbyIjnnrsCHiesvaO79fn+zUPsD4YCUX5kRW1nEg+GLg9gSrvsVwsU6rNZ
/S3JDSHgfnydpVmbOI8wFlM41lwUNfe7RYUu/Zqz5iiovrwfL+6sEcPn2f7iZTBVgqMnVmPTqhKJ
S2bOiaa+eZFI5ryFUi+XkGR3wXqpR/9gwBLHm3g8CPaRcG3HBJaxbOYWXCCI+7saHAzNO3qscUoR
ToUJ8IX9nEFBlRY41/eHXL+WLa7UiwTQjgJsBmKMslZHgM0k6EePCz8Q36N5Na1352s4yxcpvimi
OqqYw/Qc6YFMK3gIaA2EWUB+F4VfC8b8QHAOjnpC/MiY4VwOfgaRn+oSrI8LOwAsa3XrXBoQgoZb
nWpWN2N2xm/ojJ1oPPHtzbHXm4sMjA+XGvLLgPeuUFCoIxSiAR374puN8WtWWHSOvrxj0p1eILBN
V2wlGpKey3kiz1IlRs4WQTzzk39/EqMMo3VUSf4oTNmABYGwo5GzBMDJYNjQMC0O0cnXxNpH8oB+
u+S4BHQ8qfQGUJ6K5zCi9WYRHNlwf2MAXHqA7uPDiWfS7gjws4RCmMJgYb1HxBT4J3FO0b5Ov352
cMCUGUnMQj271OTpPZ2se7FrrjaKIE/G8w6uV+hQ0AEV5EWUQNvX6YfttsIbm5bJbO2QeDR8Bclb
8Ye9TOGGqC8Z7XQd0LVrFbVJ6rDKj8MDPREpaWL4HIpq9ahUKoVIZMEYNxOXkC85EZrvhtRGzklD
9iS9QZ1aUr2rlNoyXfiLcej7++osbL8Xhit0fzvhcow59TUSIqyM4oYDztG1LNOF7Jiolv/xadfY
J0LIUtbJ5yAb33Rxvf7zpwpswO5dEbXvAVcFu4R8qKhBkki+ppj+PizvjqFbEQSpWhC90E0hPiDM
aHlmihNYjI8/IkdFQnCzNX1E2EgiiFbDF2vQS7Fs+M187xfHXMq1tZ8jyIqt6AF2SwuuCAerekb1
PTVdUp0/h0YeOKr42utAb9ynZu7V31En3NnhDmJjHbh8nXQ9+IqqJUmRE0uMipyx35R7oSdeFo5L
ShdwPtxZ/a0FYO4DS2GShG1AbKfHOOlrABtxvclhjwj8hUOFjbcxiVnVMPZUSdnnCV1bE0uWare/
P1rowhrh4kZCqM/shGmT34uWed2LuaJJP6o7ducACHqcTSOeqL+AiDtH7STR67PgN8vuaJZaSOcD
8gCytTCWkEPFAJ+4Y5dODTgcKGUxJk4Pp0jB5FEonxDZegeBi8GeIbvI7suhH/FbmCHr+jDeKfZw
HdXOongahN2GupukHd+gLtwOaUB0fOFLghGnR8wUpJSYpBXCyR5c/XbG9FgdPD17qgIL4cLQsz7R
qTCGhxt5O2ygSB8qUEZYAllVRx+KCIE0lOU+g0YaxLzgQRL88PwchBlKXHDwAFNizs+vYO4sG8xD
Ion2kR18+zuAGewUeqtPdgc974GYfChbhAGxZ+GndKAxyIM3HV71eGb+DKfC/krpepZswukxgTZg
/EZOGsoZuNYqxG7ch5adhrpa3YuOD37J8bn2lJcLMI80OQGWbxPk2RA5/wZo6BAyhY6rrOBdocW4
K5Dd+gojGxUG2trYxuwndjyR+l+xqUG234YDdnQOsOFlZ2kWUDK6HdXWV/i1BvyNGvhIgrYDmUSn
BIre4NfyWg59N5CnH2nNYC8brmlqNGWLOZoLbJnKSVSHLf/WtS5jrucWU+qzD4O1SUoz2QQ3ClfU
W7YVJIbLsyvmwr6F0S/NAlNPzcj9tq7CTEd0g2ruXCVFibGDn40lrNCMfuCaV2J8cFMz5vpg0XHY
K1d9ufE5nAtDgRuY1sf61mY+hrjyzMH7fpNZTmrvyP1pECRKOVHnoq31CLgfDf7dnnbdIhNk/33n
2rtYGE2jup8YL4SVNG3+JUgCyWFxDi+rrkKmXu7s+YUd+9O+YA/Dzw73cKFEZGhyIXu0VQw3Xux6
qDr8YDVi8N+e54u1E/NPSoWTmMGos+Hb/ByZzRpvj9AcFjdjchV2+h1V6n5QuVi+mFOnoMFW2Lkn
0BB1UyJ4s0kT4U75Tl6ggdbs8XoQbkX7PM3VVJPp9+QIsNSuZ4WfdwJQ7qBbEbzzHFRR6IUsYUwT
w7LCP+lnOr/8qEnadVNjtCGM47RPJwhTxFw/JSgA+eD86BEtXeu7qjHKkupgx/P3RqVKTLrdnUtq
qmNivqfbRM0cqy+dkJSyMv+JDbDIusEGbshtatHIoPPwGUSuhij3D3LwmMI5nwtC/1hD54oXqF6s
S1jTlaC/aUBQQi55NdR9c///mHqCQI4Fo5+b8hg2molKYGUZC2vfu0u/PHERtiSVU9nY/DqvNtT/
hgKJJ3fPRpo89M3tBF+B0avAs4ZgjVhwWRhtUhjH2T/cqnSBDPuiyE/a9/RsaFVyyo92mT3x5OEY
GC+soXVEMiznkHlxU/Nv637zFh7dNyZopjQx0+gn7VvGtTnw+KG+Lf4WgmDTHWKArzbrj63aYiLi
0hFjWRmdkEu62kbLUDnCxcgpStKuQifwkcnUGbxK8Jb154nDAWLHh7DhG6hh7CIzXVFK03LDSs27
/UK/rMhRy1YDQQrZvGTzD3Un0qEvLhV9HJnA8pC6mvIDd5YmFQO/iPvd1jyzKMII1HWFrB8FOYmM
+BnwV/2v+pvNCu1mo+/wKSGUc5Xn1IgjrKw1AhDiW+YtBDCVPgYfcvu3xvhYxMyDqv8plb/twDvs
KYrtARW4DOCCwfbRiCM5K5FNOmtF/tuCtmEUKLDO6kuApTIJDBdhrjGYnlGUIcmFZXS81OzFSPdW
98tt8iRqoOkCuUxEmp82WPsL/tKVOXp//dBGkg03HNGfxJ3Lx9mzJF9KuzIISt+Uyz7BxAJQLPic
MOSpJf1ZU8g2g6XIz44E3zaQzo4KD9wFxqRVg0LjpTsCWaPkKYpsrCFjSVCqCa2TdBctn0BA8U3S
ebgPWOXY2ZaWKcMk04+HxNCER9d3GxLukYqKCZrVfDP0ARqfz49qb0pPwK4TR1iGfMvwghnXFdzK
mmHMkS8+EJeWbnR3bOE6FRB7lcgVZkk3AbBTt5WDpzhIxTpZ0z64tYKDgXCSNv6DYWt4q8CGTcsg
TEc/wB8Y+pHeICCJiskqN25dums6noB4Qj8sx5n6sasZdGy5T+1c/kgYg4K8bbGCfXaMn5YzCF8P
IcrNiHpjffV9+2YZMm3tPxatauDXMLnlX+3U24q9FyDG15OxHpqNcbsncBuCSurrh805dXb9kNVB
Ra/eJ/kpZegx5F7ehYQ/b0eG855vUCWm/EEDSL6KlBzXkbTdlNbvBbmcRcJkL3zHLOToCT9MA6/T
kVZ6Xx3hmXhaVn3DDAtjOUjy+G3F71Y+XZ1duQ+VWvMXDFNsIX4M4xjpxBXhtUpz3cDeb1Qxr+UU
L13Wp1+zU0bnNujsTzzKEJM0ZT33qZoZ7WFLHcd2ZaHK9bCE37w3glpj8w747SU3hTJgORwUC9X9
ueaYdEVQm+C6cQZ/UVHLP4XoCCHluhdKET16+7MjknUB7qN3sL7MdX1yAaJCfKskmADbncUceC1v
//tXiAABebnZ815EgR1UVAd/E2SPjg3tC7pMuKms0iJqIKkw8KfXSf9JtpvWzg5TFYVLSU6/koXH
flviUW/BO8A3nefFYJ/zLoQ2MDe0D6QHD+Yb1xNTLFtTX9aqhjsYYf0lW45bRKMjOMio/wAuTvEW
L1MB55H2jT9Ouy6EQ+W3tjkY7gjB512CUAQAu0yUeoe6GMvozjBTfDoC9X4n3KH489Ec+FyrQSFo
uw2Na7y6+P0tRUlyhxWbo9lQWSOh5nj6m1Qn5GpW+NcQZSeiQAH/JsX0Q+RALc36glJieu4NezKN
gbz08pOakPRGvCKIhTM3qqCURsw/42sraDYrzPlwrIrQlTuIAy5UmEB5zZzYaOZ5xMafUihlp15M
ZEdM5sSrTh7M/DB4+WJaOIGjV3t3P9K75Hn/2VyUgp6MFIhuxZJQRl4acmTOsUzYOlEsIL3QNGSH
Zg9H6Gw8VIcHn7jdQpyuFRAeJ0GNieu6rW0wOhEAgt6RyWTqCLnxlrS31r3fxo5+NQZ46Ntwd7m1
Sl6+JvdrWEX17GGQghHJeuknMY2ge8DXNOjApJmN7fl0g6rSQEvNROJV5XqngJT6CnhbDOb0W4xA
1/hbcxlTt1jyzhFGw84UzKLJ65j9fSmroYQGbGMRWMueNO36jFXee42sHRn7cCX1YJHR0d+aaDBe
x06l7GazA/cteTFTkRDkKPF4Bn3625xu2wSpSqhivaX7Aaa82ZP/TIiM8dNc9uBOVcytX5gsisi5
euMPU84NIaXD5//KwZn+54PIEMsC6QiF41Qpz66RYwlxafONzCvn+OB0lYQVlqlKeMCFk9I/Oz3L
5zEsxn5jgKRmvuHrM2xi7rTmD7XLf1Wz+J4FpNCapnywxWU4Q8ek50tpHXbwkR/5yj4N8QWQXR3H
gV+J1zWOqeVIlWMd7IBGgwSxm5BIhNb8hYMyOFZy7ZFRWlr7hoDDgyzUh0K5Zawjk4MWOASxgh58
2PHxL+VXX1oMo+0ubQTTKTyvkpdVtDNvPTOoKhRCvzEbYs5BKrKF8sGO0h/cTc6zw+bTNmkm6G06
+0iQ0nLjL1dHtiERpUHaKgg0IS6GztlBkeyu0ytQvb1ZuD8q6SYHAUrkc0MvSKacnHXV9cPuW/pC
1uZspA24be/qDV4k3CqLEMK5pzZQmbZ6EVa8n38a/C14Bm0gKSrvzQujlbiY8FGpTbB9mPXJRRtq
zek+aWzU5LxxRPnwjWyFDUm8XD0go/TB/eYpkOspk0gey3+8MWm53uRMnzQk6CI4okIN4c1dXAP6
duQ/4nhuSqzOww1ZeSqd0JKYPfNPMYYpkhJvkCaPlN+v2/S4cvJRm6idzVn7Qd7tkWRKFt8GjF8I
7GwCny6eTc9HcujgLIj5KoE3f1MZO0t5wV9WIrxuee7a9zfCeQR1OtJyWRoYIj8985WfWGzaCEvY
+fFtrRXUAKXf/F3sB6wCdQq3WWpYZb0ub9Z3BS8aYds1+5qAds7Bcv3W1ZEs+cReuSisPzSbMQwa
7PIWnIZviKH50n6zjZg5lgMSd2OX9y1BxLRmtxTma5q1NTH1dAVBdVXke+uiHGc/TElJw/u+sgmB
e8NlQ1JCmw0eDT0fxRtJVgNt21rjWzmzxzRdRxKlQWv1v4O06vlgqzNCuk7lOxaTJhNQ06uGalH2
5QYQLPThbbpOYQpA1Bq0i/sDrLfwFuP59GTXoLWjxXkllRpuO5nkpIeib15GpCYnYP84xE9wilec
MCGi1Nk3SU+UnhndO1lUrzyqfChi4Z+coXBVw3y0lmxOhgFrHaqhu+DP81D8Tj+cOILAnlW4K7Uf
H0wXBCDP4rNVurQAKJSo9ZWg7wU1CfnnS7VG0Bkmar/2Z+oLbnVtBMCdsiuc9dvyQ9bP5f4b67lj
4s5I+wVc/ycTwIteWAxJTwSxVkbBGwIV22OFCRrub6xFyINVdb719huTylF59XqpurNSZvQMdDl1
5kr2kGW+9c/z7fNQp7k7vRBqu1sAdjEhuZTjCr6mfV/c4vt5iPU07hBG/GW6gX8Gq5eK7GvST4c5
CyIEa2SEVsYTGxh9axBQdNzPoYGdcqhVrzlIDZCHK0hqnxEn+AsY3yUno10QtkfPpniCVrWIIT2u
5Uu8I7qcg4kP9Fh6lAEFWSMeKKsCMDW4wmJ3pWpCVEIjF6UtvGBUDDdd//ga9qss4Q4QjBdXwMdp
t+16mxAXbg/lUqlEWoPgnUyhoVdc0esdH8ALpY3C7Fc8Olhfdb/xJ5Xj1gxXvoP2HemaH62cFIjM
N01JasvT14odvpwrmN9xQVIZIZPMeapYAic6NTUSocNehOHNSqP2bcNtmbSyzmdmO7/TnNg4r4zt
DypS/22tJM524r0vvEmxcBekDKbIlj/SJs7c9V7KiEfgNCHBOX7O8y0nSDghisXG5B9YRo5hlX9D
9pd8YH0ElHxFY7/2lD7Fnh3Y6eP2aqAq98rSCKtrIYiDdvvS7iaAnR3qTgReX/yBywwn7bluEN4F
Nw6TT89G06iBfkay32aTuMOne5Q+OtzYOcgbBJ21/KeV92Fu5Hcoj7iQ0qZ7QiLZhg8gC8Ed88X1
DSAC/5nS2E6mrs4wLYTYpCAMk0NoiE/67Pc3T++ks0dOJ2rvkJcjjJk3o5EbdX2wTKDd1lAQqbK1
b4lj+LElchcIjsDND+Dc/K1ny8apEAJJSw9qu/bcQFZeYKN/oRCaKcWrJRRP7NJQvyLYgcD5TI10
0uDxbrtUU2PIh6EzWpi9SrUrCmTLf/CdmQJR6e8H5nvxFWfntAWj+uxE0y3YRMy7AbDBmiDb4F/p
pawPLv4znQmFB86prYxYDNczBlrPOI8VHxWWOSASLKE8e8PgCzn0QnmDgtgTw8/bKr6BP0WErV4T
NNaC3GlnVgAg4NnL9wSb2hLHrAxiA+wUENTHmpaKPqtdRqKyn8xz6cSlpyrDBuXaQUSgwlLr+Qr6
MxvICH+lZYKNlY/x467O8xjRVtlNZsekPOuAAw6TRsm/4GTvG68s6mDaBI7OkbU2vJz+c2Ts3Vl4
DVa/ukmiVLddhk/6UewIBaMot3z6OwKC1UgXjGL+8WqbwOUYi/2QUIl7UHd0X1d2dYWRcOMv8zmS
QrwhO4f9VGa3dx3gU6R1ryuI5nD4KDbMKp0mnP3SlNQADrH8kqzZt8rfT8iWVD8xcid0dWzITQIQ
370JY5gkz7Sum8DGAYVkrfj8LXe+IpKox/a/4qPkpCAoSJ4cRcjWcbpCOBR0xSy8sKsthfPr81rn
XDa+a07ZCNPCQZsGQYn4I5ll6ske+1F/Tebn/oKr8skFtGffuo6A8j9jXwfHlJgB6rxtbT1VXkHu
w21HRS+rdsD3a/6jL91PLgTkLBO9eTbu9IrOKT88t7QhCeIMdbDgauGwsABpT6q3uy7gydPTO2Pq
uAD3m4woixyM+hfk7VYUD9Hgayi4jZp5EsZNgZ7GR//kYKYbFLFWRs3h0plfwG0XZJsXVZ12ca69
iKZ0ReHjdlVSR4wMKl2Lq091dq8mAojp2FMkNjnD8a2H958A+Gu41EQ9eZ4wUhdmYO2di6OF/YQG
Galjmp/x5ZhBJ//A2BEl8zhgRXSgjYH5Fpy4j9aKJ81FDakT9Ru6xNPmra7LrCC8lnCDi3ZCmIfE
u9jPhEuY5ACep9+bkckA6OJQy6SpoyDeEtgR843hYkRpaZfN0nc/giZxktaXS0EBF2i11OFa0sVI
lXdUuc2A8Pat6veFa7/1Y+ctBbyCyWlyEJHcUkHUcfAZfzN56fGRUElOTia7NPTQUxvUeYKPyG9N
H5DmWmJEp/hnEiOJ+3SRt34zquqhMSVvBzQ0MTVrBuaEmfqtmzxhFLXXMPT9X3kb40UrXahxqyAR
ltUFQ8bq0bYbJc8Jbqrj31TQbvaguA9s2Ni4ohrIoexMMDpGg5uQ+LEpbrE4JmwY+lFggrU1/V28
2JeJVjPRjkc4epLkMTHSWu1NFuSQfTDj/xFvf5LZfvSNOXxGY26ymU2IA/A4zR/sg/ii7P7nTPWv
2VNboP1NIz9CVHlxnTsDoYg0F03bSG+gpf4cX2JnIxVV9YWtFDj1mo3yIhDHSyZoZzH4Ij3pSUyQ
B/JZEBQ0tyIR9UDpTgDETTTaq3Ihs9hg0W/+6/yjokIXGr5RJ8D6z7T2JLlli7cDnI3MKdZMo9VZ
2c8M8O1Adn+9jIbo/nrSovePu19pK+yI0qQihaL9Ko5ZNQ8FYWDCox/OURipOnSbuZ4m7jsFbJcL
EwsYIjzE0N+s/DHovayGotCOGwWEH5Bhcy9FQlKuzYATbLNaP/sP86kOezPLRNiKOEZCkcRhHXgT
+AgF/XSHAENfO6W3jOvgm527ktCwOtcTr14bpmKbZULrys8pdYUrtnhq/11i2cZbxXDGP1WJ8dRH
6MkLQpGlbGMI+Vj04Y3dltUJKKIpfQ/JT8M9pQqj3CFSb1YHsuSKoNipZXUFmPJZzYAcLMtqi5ww
cBKM97SODa94WDP4MTsCP4wCh/Y6nYDA4gbuIV5/QSjCA0Ar9h9CtM9rigmdqQZGjedltf1f0faL
V9D764Vr503svQvN6plIAiSrMhHUwVhLDv6VIFoKFxNRB9sLMPs8tPVkPtHvhb31tksWTmh0gvJ3
n8zaKp1NQYhRSEX/VLl2L4sWL7vQGvIKrO62BfbPd4KMf0csMa0BeI4rEsCmV6/lNo3WT2rDouzD
NJaMTb+KvLj+iS1lpgUM0/wJAM19aJcTylJ5YuefaDF224YlrgdtVn24H0S0KDFPL302D7WuOv0T
GNoXC8inJsrGZgQBgOUTdbISX5r23zZo/Or/MLaElz/sqhf3x/Al07AhoNmWr/ZipAb45qL6DSO9
ms7qQEOgjI74zgmCwQFR7Xj+7JvJWiGtyrzcHy0UxqGwCzCh0/vuGmO+JCLBzJHX7xUjPAo4LU03
3MuvwPBSoWy4zaMtZUT6dpReJ/CldT6Lk86y6plQ7Fn/0TuKDstYWP121tsvKhwJQI85l0bSsp0y
qaedsV0DnxjtHskcYcoTme5Db4wveue3OjoSGYPYX889vJFSpNvwTF6AM7zVjYe72oJgj+1jsBND
fzy9XXR+mYNBB1+MM4ovNnRxcUvDF71r78w65vTRkq6pDnGsCHK/MQpkq326/hZck29Nh2ZVvOqG
a8YE61hl62eom+nd1q9Eu+G+S6blGJue/jEgL0s+bxwfKrwKdJM4YwHx/hFqMuB0MZULdEpsel9u
AaFZpi9cvTrItoFCOBudwzSJBXWFH121whdoDbO1zrwnE8i+KjNXqMtXM+KibsI66YHPTFB+mNSN
W46DKIwix+G0Rpq6BTOLlOcwVp6WRLBibl7qyIl1qPKzDBtehuW24FJ/tp+/RI9ptrRuFB4YfM2C
wrGlTu3sYTlcjpVH7QZ0+I+DwjEoC0hPFe9v1Odzb+g6ycUS3x9VzN+PWhC5/D3MTxCNx3myVOTa
dVFyCGvC8bmhNPZrUCqBc6F/fKu8n4J4zRwWUOb2M5IEP+0PAaebJ5b6OR38rWCA6D1en2CgFq+j
lJbcfgNNMjKXvm+qDl/iNGfkf0AdH2q9Kelh6uuQp4wuIi4HFYkT6oxcXFdV4pxtNjDpwHfflCtv
34ouqugjaPsjo0OT136XhYxWGT06iKGNReb+cmGuLmj7gCUYGrP9tVwo1RM9bzrtesUm+9ZDZDT7
n60zQDVWDfh9csqR7PR0V9YHMvZwSN1AfdBgWQJ2nYL1wW1xc67gAxW4183uekumbGf7Xjx7QlIm
gH/0jl8E0hFALawXgTr/TLUfv60GZ/grkEtB3utw+tKheRuhmT3IULT8u7mmOXeDb/8vMZZKDGq+
73QNlHGBQ7MlFgET9p3gIfSWtMqlEoSg79G15VLEYn9Xon5wMQ8hOmeJ0GZa9GB7V+coUHqTznS6
NFTSoSv/jIw07zkPRgJI6vy4bEkN5PyYfFSydNtZQDZ0EXTweiVS+0iJXzaCY8r+fbePst+glX8x
K9GBSNR/ZTbXf6tQh/2raueCQu5eB+50cVx52RQ4z+Iqgl7vPq0ZHSxkdBO9YJ0J7hVd1o/nSPbX
4L3XEwAlbRKQbkTgKIe8uv99T9Hend50qcXMCIYf4dxMz4uJJcQ7hMFci3sbr53JuTQIAn951XTu
rp6qeK1IPWt0hAT0TgZLw2A4ZkFDNvB8/pl1W4fX3svJwj04Zurpdi4PqK77Ids73tdmO2gtdGiH
YH7t823lYb4dyZxCae+9N3CfOSyt1ctJz72mWJqGAJoF8ihKYJ1zUr8V+BmSFqNhJx2x7kPNUNmz
yBiJlH0BRuUQ2C/xo//kzoab+c3IrDe8COAB1Jqi1stsTYN+Rql9LYLipvi3y51QtBUojJjToyTT
u6Pffu+1ysd8fk+UkamTHSEWPHfUhS9p0r1nWzxhaOjfUWqEI6Bxe1srDwfnuiGP5dZ/BxZFDXMb
C1WEo8JS+0Y3bwK/8aedaYuFjDL9PB6MC+TVWXW59fXBYKe4fXlK9CmeCSX84pVtNkd1DZwA0z6P
qfQ8n4LQbcIFVVMd+uTzsLFsayNExl38NfdJAqIVfp22fGpcu1xiYe9/bv7xnX7Xm8B37wL6iH8b
MP34Zo2DyfTTsSZ+n3YipAqv/phogN1uyecnbw3Oq/RRUV94ZG0bBd1gTDmFwijvnOPP7o8jIynB
ZXJ8w/JpFeR94xUKbdcdxRR8YlTZJuNvNYo+WCVimePhmWLuzwIBy8XOlZ5SVj7s1+zrQ1trmPFs
Ef2vOP9KTFfhfahlT2rFpU0IXmGFk7eHBzmTSJWOeT8fDr3QeE4tC0nMybpUbfWJxLlGgbLGg8V2
XXmIznByQjkyCIQ/PNkh8cm4Zt50DVFTv/NJ4APkp7JariSpCYTrwVRpELfYAWfiZySzJ6cUpCKp
bZnBU+JQHPPJblUoQZBlfDebNLn48id1rW3myqfya4zSHBJBH9fqUkvLCH4e13GwgKvCUh1Yhm7J
mF9ZiJoLkYaSclk4Juye06qSdoEU32hnmB36cpcbCib+FadAePB2UviR1vsTXzutKutjgOTkbCEC
d6IcPOqwYmQI/1zZdzI7Mu1vE+bLqm0HCl2wu7kPLCxjaeBVmdPNSXkgtB/OYyhWIKnh4GlX2PFD
+TOrehnMOKOCtraksnINHwS6OebP3i9TFdcPRT3EdkRyMBtjKS4EOe2JyyPwj5smIKOMjaZlh0PU
FAryuCNsvyPhdeyp9YIdIQBQmE3d08MEEr63W2jYx3bjTd7QC78lhw661KQ1kkg9RggXk3Gpp4Pn
yEFPc2qii4ThzZssZ3dnb1NzS6zWD+IcHTGiCGkShFMct0JIJppNWNf2nlLeBZD78Q7pmFLmo1FC
19//3/87l1a3InkuvAJain3FVy/9cVGRgV6nB9CJXjLPuotqAud5dfDqwlv7+MlGdm/uyiFsisLk
zvdDZaeXwi7EWX7RmoZIk2+Uev2t8Zk1sHCfW5W+X6hR/R7eK3vdfF6wlRJomdJsr53WVeH8R4hg
4PbNr9y0YDZVRWpXFw/jY18dQkQ4A3KT8BK7LUdTEh0IkP6b9YT52P+l5/mxOiDeOHDf3MOrXk9+
Ah413aEkZbXFkChfHdvqwYaFBx6uxwvP+JSQU7IHctO4dWLsPNIJJW/KjuKcs9M64Dfu5OmRWp4r
IpYJ+qpCAghrYbedSi8L0Dv8uNv+vTkqILWADZhWkbdYvm8TrdbG/Pcp/KSdbarpZA/iN3CxRa19
in0S79Mc+PuYWaZTenLr6d6XgPi0RV21QZJGAfgn08oz6VewteUj64Zj8O/uC6KcXL2iNE6C05Cq
jh3he7dxwubKzDNqhg8IKeeKgVohMsBIBbnc4NuWrtZ1zazs6YpPYGsvloELkaeignDtBrcUrN9B
IcXaExKY03Lw50Ut+6iWMJYSuDEINxxc+cV7+6eUPDOY/oVWyrK8307fjL6pZ3VwozRZaTeTGXUP
8lCNRN6Bz1AIXjYi2+8wDvgcoXGJcXniiOeV2hqFyWT5mjMnKP+MamLPGuZkvrfd/yPgeVh8D0dX
YV9BYfHpwrFYfokEuJcUac8aaltM2yNJ+sivCVrYmbcR6wGFtzZLzUMRXsJGZ5tbVFBbISx6BZt9
nvazQRjfSJIfDN68tQ++7NwqLfB5yH2HGBB5mdbPI3MwpEwZXVNarwDElBtawYq5bJ0TOt6BUeOh
9FccDTR6Q1VPl+mWNW3W+r+mKNGNLIAFqXuVwxy8vGH/Bdr4eHshGuNMdLxqox0poiPLp5Y2Sg9f
1bDoP7R9vhiBZjEbFgwz56WMJC2GpckKdlAuk//goL6I+DOEa8pfU9jU2qB64tQf9xxmxYpoziQu
52HWXju1Bfz2BRzWDGjcaja3SB95Du1jA4NJZ1KMdjXjMif+rvuFEBI63J9V+ctYbX1lbdB34sHk
xQEh01Agx47bAJi/lcbw1DB7xlsMzHt7StyHHKk+or9K9A58XvDVFbKFy3J4GYY8Q7UVbBPNjeu0
s+x+xsb1zniVRS2HN562z+dc7XNroTO8W4LxezOdAo6uTdKENLI90NOLZIvURWylzXEfbs4XpIfC
zlvzozHPkh5YlR6L/Ectm59Q3JsDK8S3vAd/Djc70Jsw5HEjDcnfCU3JwF97b0EuKm+uRJK+yPlU
LYEkHDlYhC99qau+wJZOT8tZS02Lo+ZVmbyTDYGzmKejjb19eZNuumlqbT3stbhcpZ6+QggO38ZB
zYXtOqiOpBIvHMZC0Cyh2K/LWxyECjzBN3IivEsGLc9uv5GWb9XCB2vpLUNU2wMExSi4vsHRt3Mj
eGnH6DLTdpbyUPG85xTvKgI5X3sKSNV4zZ0ui3cB7UIJb0pTo//YpqIY96SD1IZ+5LWyhdeE9hRp
NDCrqrDo1+ah+lc24Ka/DWzsm94G3EIlsOlJKzOl+6j3e2iozyZI6TBNsYF9RhBZY3xahq8+gqCW
ker2sAsB8/65YlG6KAstWWl6pEj0qtBDblajpQN8d8VQ8ela6hkc/kkpEdeCWAU4A1gThm42g9ho
mh24HAq9aLAPNBXvOIGq/75GIhURHl8BCFGdcpjgvbX4CL2N3krCe4Cz2gcArpgCxGgcjnGu+7gy
j8BBjzIIW3YpN5XGV0QPEcfbraLEFXMVD7tPXP6TXbGCh5DprE+TingFlSxG3Mp2nPRIV6b1re9o
PvnxdjpFVk967awgJGWrOFM4mW7GzvZN6rdW+yc036hRtI15zUzq893NQPa9le0wo5mDDgr6RQkT
jp30lNdjfIgQyMo80hullsWX+ErFQAp4udoTg4K5Jlk5AaeE4+ZVTZuGc0M4qCeX8ESdl6s/t87r
duFJcabDWOgBvVkrYXC72UWDJbDrSoNmntTa3qM8qgwfXjglbpY+5Fo435tAbvs04QRlqr6sTMiy
F+vx0cAcl4Ryd3BLJ0bIBzk5AG4tdEvObSSxjejb/Ced5u5g2KssZ7v7KOti4VFGe3o/UVOyLC9e
n3gbc9nMWLttkk+yEHHlb/MoxIlJWV7rsyuvDgwKy0T2kpu6C7H17SrzgWmF031f4rpC6y1BmVOZ
xdMyW88efoTAkYl43ItwXhMzxfEZIXYsCHg63AgOoT/DpmzRjAsz2+zhgLnKkhSdSnIiis+7aS/6
38IAOEwHiokeN9jLYTsLb5SApf7q1eAvqGtuUrZlf/zWnJI4guizp34FmjqpthLPZUM73ed7VfHj
X6e8wRk09YaN2ByIPvj3gtFHj9wGVx77y2ISwn8LkEfeYYmV2JH4wg987xAUI89S6hFxhcv2cxaz
3cdG8HX69JswjxXsglOZdOHh6yGfJb/yEyLKS94wQ8X93BG/fAgKUgouMu/ryommFE2rbwvhJZ1S
EiyJKjPIMvfPfS1w6x4fXpn7/mME0tn/0zpcG1zCD9kbJPRymNYDn1O0m3tm+Idtbv7IeUA9a/35
n9QeTeElgSkIv48AiIBavnNjMU9F5jPuYk0vNyiuFbATuPEgt2SHY77Kb8kF1rx8ZR+EwqSSElX7
h7lsTPNu+PNWS0da5Rn7GKgbkY9p1ij3flgX4HqVv0gWle25Kvr0etK2rEDImCx+cwKhE3la6zdL
9VRxIrlSyfjtsbVgco+4lWW6yBxjS3qfUvUFpTC9hs2a3c/UsAZ+dQsvkWB2d2f1D9FLTUy7y9OA
hXuyVKOfvvXX/hXbqrLvkFB8mfx6aZbiubJ7VtjsDSIipFLmw06tlnwTwUu5WfvK9s9OrkIF543P
AFtWuPoUDNWfSiz+8MonQE8qyy6iZjbZ5LupV2Iko98WC27awa/p1I9oDixgKn+ekCQGdrhMt89p
9dupcnmZqEmQB3FKKUeMo0vFNoUybLFt5Hw3WYWjTHygzRAHbwPndVt8tXL3qYkqJTnwjuv+4r2U
UMEdux+05/qKfUj7ZwDoWFR4O0ms5caP/s3prxUB4pbAlg9iooQzG8xOoDmFLUDPWCcJL7nkqzLk
dydiB8pJz4nYlcy5Ga89AHbmvJw8B994bIEufwBsFP8d4AKFhiDw2sxOfO8OmHly4wB7dMedCtAm
+zyZjtE1gjiFYlobrB8sJsCp5W7U43gEdYLloT/ePsSw5uZYQW6ASK8R5d3yIv2S3MEh6eLGaSNv
F8usZmd36LUN2/XnWitWauikWfA971AEYTwW6YAbMqNRUe07kZceqT2VJAJNwIoLiXMhXU4u0TPL
OsmsSRmgXK6lhUfIyzTFfohsCU1j7pHuLk3YAxUwWSZcQAfDteyZr+8rYkWp4MkEbZCR8TWuCM/d
5AodzPbp6iiP1OfZS31cRzlvm/9TiAerImCUUxXb7ZYmWyYRPR3yILddliP5hEIdPXTHJCkiYL5+
ObXCDI+6WEnYeVWSgIK6tOVqJYnWSFLGnmOcrLJPKhsqDlyJAEvQpBJf0y688ZwFp5jzpxKQ1pb0
abJOZf6RzAic/rBhn69bP3ga4+9ZPhH1bNhoreON28xxGbbeg8ZMVzy/okzkBntHOMnJV14Udu27
aT0iS8RUhOvJO2bJvWtC5bgHCFHTTTYM7+lvBlG+1TO3moMzhxj2nkrysP8E1BhF5sCgioUw5jbL
wh64pt4Sr/6BH13Pix77XS45cqv/3qfkepkMLNDO94Xnp4uowzO9X5GbXM9U+bz8iOz8KmCX/FNc
zlTWGjGPEoqjnXJ+PxtESNSyQ4UVN7IWUW5jFA7Ka/tIMmUQEfutUfcrZFbSIGQkl9eS2sBxDNGy
20yrl1VYvhpNyUP4XG95dozEx8mUmFFNWDYTaQeDa8/iaIfUeBtT54HzF7/kHEYb6bc8ajvBQM90
lREU0g6mJskzTaGOuinMiPNMVdrYSaIvYS9UKxSsjad/bK+spUzeJKY877n7bcIUV7B/y0708qar
FUSPlGvwh4hKo4E1c2pUtvSB+wVzBfIgT6x8ClHxPBZRWM3rXQ0ypDfSFePL4aMbi25VmOoJhlxr
f/w6sFGZeaTjF/M+l1RteRfitysHImxg4ec9IDKJtjxC7an0TR90d54qABYZk2KBiGs8iI/7mUiF
kj/XH3ow8lOnvTbG9r1mH8lDW5oRKLZNd/1n2faS9RLdsRHROHni2u+hk9YfRGyPsbpzVMBay1AA
TwvYSuOAJWoj6EJFXMyMsu9fq5Pcs6dxHvo82OmzURj1/i5DSy4WLbtqVf3DekpAZL7A/J0KtFse
cX5FJ6IeLEeilLL946Z8N2Jv5UZtwkCM6eWwNgUQZ6Tm04NiOATJs1JMxzLlStSTng+7P/isAJMt
26kuXq5TBcBT3/7l3YJYkCjOFr6NeNi96Sk9AkYQ0hUwxVH1Nwy4ZG4W252xwtsGb+gOb/KTpv59
tNDhn2sZnzhtxNkGyQDrfAzkDgB+JFMPTBVqhg35ZBJp8VLh5wGJMwBlRMS11xgZgDVtJqRLorjW
mfws3lBWSOZ5NbwAsERas3kv/QWU9yvKPl15JUntTyqrYOGzLwaPYq9RoTsWe3SKp08L3jrYkEYb
8aAc/zXXemoQdt5Xg5yL05dQ395YrRnJodweZs9TgNd6f7E6I94GEdf/W4htelb3pa7ldPY3Q8mk
6mIN7QiVyJv9aUu1xeTWZMZxrObhMOrS3/AtFlLv3fkPUCCZQ8EKtfrhS1kGv5DGeNkiWD+ozPs+
aurIgDf7FKS+cB9KHvpYfKhPVcAHyDQPU30gRNaw/hNAwtmvJ/lk8mcrtE/KZtUxm4xaLjK+Te14
ELhr38BvLqwDXWiGG4WXa/sC7+5/rMzG8f0XUZMkA47FBSA7cB1aHSFeCHbrvGMCCWIFJcw1oM2V
n8InRsQPmZQJXHEovUP4cCnpm+3o95BN4WJH+qenfLlD/vBmrnLxPZg08C/Z0oCevsGJYfQh2hvh
co4uqeZdFv8qd95+X6McEMK2aapZ07rztwt5efwnzgoOMPBp+hPKXsygvh0oCQ0P+rfBm+mpOr7z
p/IpqUvvCwCr3fzBVjUtP4ahHekkAMxyCttiRl5UBrvOPCDefhztN9Cjrfl1JwXTfWUnA//Zkp19
0R9iG6dzo1rQf+yrj9DfWfTBI5We66AtHHY+L48av44x/6Tl7eb8q5QLYegaUR3LJzS6tMXnMowL
0ghtH4KPuG9XKWGIH4ugUOk8KB0qH/DT+ra16K1SeSp48xJ/B+vQdLNg/xqA6CV3VJMMVWR46E5V
CFJ4ZVqS3sAWaLuGrIgux2hgtxOaTEXy+ZZhvexMFmGzu5Ri7r71mvfiN4cNEv4XVpK+7CJDb8JW
dmGxlQqM1Q/uqR/RQPNkz/VVhQ3uwRttZ201twFXb/ugY1GhB40e3nSkRZQCbJ23ZA0TgSWEgJgf
DIYJt40V/JXlN3L/D63OexRU3fnac10sUBASao32s2WwZSwrJJ0Wrd/a13dhOfoHq9t4B72ELes8
kwsIR6fUySxHWP7BwIBGYe1YCYvMqmvtArXE0Z/zAuHFG+gPOmotd4iypMitjjmUdI8J0myfE0vt
HL4a8KNASwvCGC8ThgLPkfv2y+YkKemqF3KePrgxrkdJ9BhzeMIzT2K+1S23H9h8Wo4Vbe9QAcSK
Ui4bgKl2Afd03aAUBjYrj+FdmbLAfGR75g840UdTybYduQ9pBR1P5DL+5+0oaseyEIir4PbmsJT7
86spcbxr2KKM72w0/WrjbGhhQCRk8e8Bm/O66ZXliR7Ss5vjOkb2y+yxH30gtJECo1CPP29K041B
eZQ9cTh0IAdRPskk39JeFSf1pbHE/Fy+3OT9+iEO3ZROf8+ITmflllQ25VtbLlnJRdcmUeltnaxn
aUSBFtKY95lAwPW7IXSUCwVulWHxNlWyFEW6782eWxhdp4tDuXrpS3RV4niOOTNJB02hn1cM+0jv
CmpLrpyIG934+8JQddwd5iLTE4CYiqz+54DCaoR9KcXjEOV2pPQtYEaYLdlNO+LabZhODT4ZkBLl
KIDZu2YPvo3iHehnbYIVEPDoRtf99RMZkTGT0QbQ5RFbWw/7M1BuE5HCC3pmNKPdfGKRy9N5ugEj
GVwAoKfkz+Dk48WwCd74/IyWnnitZ04B1Yybf0DocPj0tyw/Qxh0Y2fxAIs38wsYr5oV+lbJWGD+
Xoc9ZG9MnTjXgCSpGE0/NKLSLpn6Zpu66Yqr/NMW17bgw4WDFKfh2NGCxi2BWtHkmexdzlGeT0NO
tswiROGOxwy7CJ9TT1Hxs8ljLjykhOBJ55TLDDhlJ0SELIjj1GmhJfqZ7NqsGCkqXfL2ectIK2u8
TfxJgo3FgWrERxCmy53gG6kzAtln+gc7NF7zNb9TpRYi50K/W/LKJK58cdfeOSJqdk2CFg9jdd7s
CterstiJ0UGO9gSfIbXiJcQAzkZYdawIVJVpsPSxj17TPpp0HIKIJ/s9ICw2wLirvpJhNjqVipEq
BuSGxuDkhm9dcEFNgNmHQ72LlXT9RbQIkas5Al0pzogbvS8C+EgdVAIVyZR/kpT3DekaF/Gu+bCw
AiPXIS/5p5Z9acGHJijJLogyz4dOII7717co5QzroyeHkGBv7kTEskRz0uXDBptlSo/FzWhc88ra
to95XtSDnnRrJ+tH1fuZUgwROagUnvUvQNqELsX5v20F+iMBzSvuxhNCRRxKpMmef9IfTR0PJ2CG
CuBT2Ij5EM3AF/dTWNi3d87rInvv8pm7LkrdH4ebcWu7baV2Uhb2wGyKg7l+OYOFeHtJyNKYmuxO
uJ06VvDD2JBLeQ4HcEovK2tPrrcVErpnlZbLT706nMA3ikn57nQLjr5HlUE/ZLjDsnNtQGiPXkBt
ZfKxViroaWoiiExugdlw35AG4d9f6nhUL/JzLsMzXRfUZdIr9oWZs/vAh6V8WoOCZpp2R8RgUYfD
VnS7dGfQWemp5+1FRVib26SrP8N8K55YFRfiEH4wUugAZYOBYXFQGBE2xLo46K/PiryE2tznYu/B
e4UshObMeFcHCPTxF4BuG4mkWLQfpzUBpEUrfaeAoOwaQNthtJlaX3hM1XmdJwV8rvIlGvLW7RTR
QqwSRR0Q/QISNWEFErE8XaMfCTOKRHz1llQ4KEFmSqmUkQbuda/dcwohmyAfiQaAAg7HmH/3CwTh
cO0MDtEzDp1A5Gc2hqfP6XSyBczdLD9BYZEa04eSyCin+tkWd+a8mS57hq6Yv/2wEoERUv+NsaFh
sfvDPrRMSUTWc5/anjGSRUIKtEviCXls9PtNjKzpl9t5y/Pld8hsDvxagBkYVBfXvfWcw39T+EUU
nHlVShxd97vSmgSskKiN/MPv0C16usQVBX6FYnzhDBphVN/W4f5i2gqb2CfylBNlOqjvRETZRnzz
yau321B/W80q//00mN4A8P53A8J+HjIloIEUrzHgbmpHbabbkXVJpKrJv8yRnMFrOOPCfc6MkkFa
/iXm/0poVVD0LE5op6XXCgQSyp6KoS0Js/jicdwWgPDtw2vkYJCbeUI/ZWsjd5qm3imwyJmgvvb4
pWc7EiTb1ehOqiV7kU+tpif/rbb8Gp1H4igdwYdodlYkVOWWvZWEbKIyJs0yUeN+O5Vwyy6QHLCN
jifPlqAddD33beiXCNwD3JNzKtjxE4yowVR91D7JGb4xzlPcloBlxlmXGhR/uBDW7LL77nwHrrkY
U7h2KdH8LHmp8mvOBYjDHuGJTR3G0OTOnFWIF4UnHlKVB5roMgtllgKpIIw5NrgKF83eaSOIxzPM
q5Iv5Bv0lTUM5wUe8PdbzeH/IMWt5kqDhq6GxiIQoztnBLrbZ4p8+MU4ACmBWV/e+G9D4PKiIrfQ
+sFy4y4dgcUB+Tdrh+LHEcnBIz3AObQlGqpGGwAt1iYCecGekUBXcRE8cmCo/mJ3/Gzut4f4wlRA
UANwyEFTMf2sDd613DJrbzj1he9famP7/1jwOjKb/3Vuq++KGP5su7tFN54EaBDP57tUir0Ja7bO
eQw3UsCE03F7hHOUT0rceBZifkQXL2uuWhK8BXdfC8treGgfe4s5wTlqswf5TYkrqZxc/8G91O8O
RZdqs8vQEoHHHveNSYCCXSN/GBpK8gp5pPvTY1F5ykuwyec5DDMSCK8LLOdcj8Y3bYhyioO41/b6
OEmTMxrp7GJCB7aw0PwWlB2djrpKNCoGaFc9kB1AaG1d1ikei8C5/zkE0aqv4OYMMAgY0g6uTGxo
38uwDLA+z3Sa4U9LjQnpS3VmqSr/5+iQrCR+n724F55P7kU7hH85OGG3eD6djXFtxHPVs2onu9zu
hbiazYQdXvA++d3pqskJpvkQYixGHCkRhxY/w3p5JflrfgqKpRuqrQMb6TzQT5MwLqn0q4RKcdPY
/qc9j0hfF6R6LMRMtIUrPdrwgX0UwP3HNosHtGRFJUgq0IDYc4/Jv77XwQDzjJVso+Z8kahQXPXu
7WPqHloBWuoOo5ZVWSAgzmzP7J9BeLtUYmwcW37z1AedRPRVxVcVlJ5VF7GPXgDj+O/j4bjHsTiM
IzIHymvDgfz2FAI2EGtGTldT2yLXkYzEOyTTW2gzKBHBTzgds8NSYKals6zLocCNkUZkNwFM9Wsj
jMQeainAkEGM1qJtWKNXWFq7jZCvEwsrN6K5e0ST573LOU/hsz7BtfgjIgcMVJ/PrqT9wnX6VXqP
++oQ7n/q0zUbzo4wNhbKe6HZ5AsnHwrONIpknDZHfuM355iF2izCIjhwqDpim7Aa036MGC25XPQJ
joklBMFeBtZihXISkQDAbCtpv6at+/KIRL6VDCbSFssQ/NaUM65WZRSv4+vMD/IjDqOM3lEaz4V+
ZzXf16TUNq5Y1hsy0R5p9CSfCK1qtRvIu2+HTtqCAeZbewuYFAmisFZRFezpOllROvgjCADu/jXZ
D8pRfQd7aVRpWBP8hQdPVFI8lf7CPL+WgeHO0SshjVrTa4Mb3aWSG+dngXSgAk5f8rh0CIl/A9NS
5+motuFvgn0ernNYSG4KodYTNieRS7y1eT4NzB4wsqeThNrAq+bbH26q+TcBYThO/AZGFrblDCYA
e4NM5Af42iL4hSUR3cZ7jS5OzBFOY/5/LeB5OjQMm90/eWSSHo0eVnJHjGjrhYGmNX+el8j93VbV
0y/j8qknPZUM5xIy5H7kzNIenOI9fR188eDycpKxDkNVHoc4gKd9bv3JFLexUSlzhPM0j0DwKldM
2m6zpGiZFy2Uw4AaEScZpItBX5KQM9UVe0iA+GCFHu+20Pnuza/SWF9f2msC7ta84++WrcMFZpl4
ne3Xz8jLp8NSQmzjknSeD1RxH3KqRDxuOuRkyw0B9TindEPmfmmI3yq9zZB+FjzR+AAYEIYhDXqF
VDGwvEte95dZfbxOHTPsTxFiCfrS+Xx883WM7hXIj6QzEzOdGrjvjLUTMb85PtLJU/C8FHvDFs2V
N+8rLmrJVZECkxYJD7q+qonhomqUx3F44PXEd+6o9tUqmErffzHqXATYTNhwhr8AVIKh+0OI8O4G
naM6NvlKH3hgW9WKfr6K4pc2bYCF9B3SThKTU92aXzn16ZTBqS6vyA6od6ACEdaQ73PzlFwj2A+s
wtqKtjeQPgCmp0yQa4xMNz2/Yu2A6YOdrIdHDxMj/0ZLtDFLSVMF4Vc9IB8g4xNK3+EVs+A3z4+6
5xAI/mKwnTle7rgXDIrQUB6hHwLjZJ/fawP+DbATkCsdD2nr0ucuk1YOJaCHvrpuQ9my7y5dm8yO
D/u9mf1EospPw/zyJZJ445JahAJGwizCmkvS2QRNyjWIidqF+PNea33U8xsui7jjAp2tjl9m2pv6
IMD3+zbV6GjHDAXR86N0+Bf6R0ucQ/uFFxQ5zn0ylcX2qcP6NcU3PaOrw1hXsHTpctlwsHEMneZt
SnGTKqTYoON1eXzm3wRjueu+GqOTQtYef5RE/K6wCHIAMTLdDGxecwo/+20tU5vB9M+nsfYO56LO
LjDOSfefR/bpjeGuj6JqFmlpNhm9MZsFCVOrw0P9/vWpfBWCYHrIPIO5FGMUMOa18NugybbcQ0oD
Yr5S8slbMD4uPUmTMJgz7dMKzfhp3sLLDVquU+yHsYQrn/PN8W7JkKcDo+cBLWw28EeMSr+J6GSt
TA8xcKZuA97znlBdo46iUFi04yUy3EM9SooBzuPMlG3VB17T5/OxwbR5B1OPt02Q86AYicJJaypB
oqkcwfnuCCwQUwcuR7KW5DszquqIJnurQL7HpzPdtzIPxj3N+WlIRo2/I8G8qDnTc2yqOJcMWzDv
ste4K56/m4UqzxdUsbZgPUH6d2g2NTGKRVp2xC68Z5eIiCiNst4tQ3aGPlPf96TgDOH1v8ATG8SC
dAvP1sJs0oB9EIO4Nxw9le6adOIuXAt1SR9w9VtEkhg2vY+VvFMpT5uhoiEaEF3ypzVjTxI+Pj3C
WClVW7wfhht44e45jcowv6mJ6aL6Tk3AVxsxb5j2J2lJFGjunJ3H73Xys5ngklhye1yKjatcGHtX
ZQJ7QFSXr0AXt5gr6qHHqJWoU/E3nNPfp7PQFxJBa7rj9JwmvhtrZpx071DVokKr5swqv2FN4f2U
qBvcPP4FQYAkyzjH6STpAnQJArfG/W2hkUbCpKtJAXIJfw4yzOY81juugKd9hgBC4ocKebEEpkSA
+xc5BcsGhsMx6WVufwibMdKw3NAgFz3DBAhrqDM7KkwKh4vIJm9Vl7OaFzX0M64bXoKhJlWUdVzX
4nFfXE8h2ZGj1lUIxV6Su6WQwCQYbCLpe7tQshT6bop8vcQNR7LSAwBHZKl/44OVsRga6jYwyTRp
TgaXDiJDz6VF2PiCKXj7XXJY0qE2xCZssVPwPXXPrJ3x8KBzevzq6S03NWJS+rJ8AcHkwjU6tGxb
SDzOrkx2QtfuF9Yln7WHY9IqfvQDCKKLruEqynLSwkC7u1xUkLflAeGFNvHpj+X2N1MLHuiJwXkz
ybjowtiQLHBPvg6rQEWR74SZbo1FIsLmFQKaQ79cqaREj1t7vbpwyoZp4n/7JIbdbRaplKuMgyW5
EZEfRzcrvbLsGBOsnp+92uPGSs5WgRwFqmNc4z9PHiZv2BnpJuL7c5Kgy0ftjM4lDRf1k8di7/Zq
+KXv0tReQvM8xb2i8PV2KIyG0HI2gUJO/gyxPcAxPUmswECEo2NaYz2gmycBBanCV+EAM4q14ewI
NslgST3FnSM7DuJ4Cl/GyhAb547xGfBhBhKIe9v8d5TyTqTa/0jAS9d+nYyvPb6DEB4hODxGoupg
bkO7ngD2uIXOEjB1OatC3R9Usjaxr3GSi652ajc9YUu2Kkk8QhjSZcAvzZ1g8cz+rfxd7XkzkPJd
FhqXkxnAaJf6SvVfKgTcyMOVI8C6ZHiJYNy2vApWEU8MlCTnl+1eyDmtpERnCNzfhuta4L82SpLP
+sj8FSO1hbLrxv0Jx5muyQuUGDIVXNjR+T0Ka5Uj7/5zh3qucJCBIOO7y9EeF3kxV9VEzFzHtXQM
wARBwQDeMF+DckGTI4X8YIZbHcSeOtwTdNYOqEknSX6IvUc+JnGgY5+W6QYCKn3UrUbAXfIpKBKs
a+zT+vWWMRw49evmAiGCL/EFNh77eLhpumHkj4vMywCVJ2psU5xhsLURwuk6IQUMdaVh8Dz+P/Pa
s36mb+xD/pLy2gYRkhGaj9dCZLVN6AmHHGI3EESVFOLRxSK5n0Upyefh5wU1/UZr5aJGrhA1PTvn
SK0rYYEXVy8LjcOKa5K233u1xRBn2folyyTpricqqm/dzSHZWhQoPiRwUN5VHCuVG6P+OBQ46zTY
veBlcvd98a72YTokpMuR9ZYem7DKmWe3uMOb651vBMRw8i2RJLIh2TcXWFaeOG4hRVE+VWMcCS1t
x1sVl7YTMZOUqWGagAm1gYixFcObcxe75QgrH6TDE0ZUy7Lq6X3pJPbMDtU5D/lU1pJqnoZdBWaf
Pr6wbBVmNf0aai8ngSJHrcTuuLAUAncKlzAOSbM39U0Yqn+md8eHgwfkh5zeSy2bIV7/JNdzUMKN
X1vzSeJA3aMosrqgivjP7veycy/OqZ2Xom34foZB+o73ygtqY445lyBeJtQkTY9lrwnfHx9Ih9rH
aw406GZVAbAwpFrROCChTEYGZUKdMUguGrTfYV7VWyo/LK4wSmRDrQtpXvT4AIf1t1KUyVhnWyYv
0piavUJbe7Fu2VSFZah9LRwOna3lGz/jl+zBxFYBxu+8Lrith2RUvVRJqkklP6iniCHNVTXdvaKM
dAPWpeOMr+46w7GjYKuqBDNUOBzQHjSotKIWRXfD9wO/kBQW7d/VcIuY1ehmo241fjrGGqiJLDca
p1HmhMkC8VoLLU57InZ/6i6K1lvoosBXaa3GphJRWuaJsyVx0V+RsHsdQS0vlQ983KPwhIdHpwjb
KWhcZsOPwjyfgITdVJjS8/wEuCcYdir3gaiF27uhWxbP3EY8Y7vXbqyyMW2KpysOmP3/0MDGaDt8
xuAh1odBxl0g82KS5U66mYcfquJ9DS+mNticfOS32XIyGbEi90QOBoVoQbrBnzMsq44o7+PMDV2J
t22Zs3+ouFObsNAZXrHWzwPxRJle+akUM2sBThum6Yn4wNTlhrVwY1yCIp0uTQaCMjCrr4ZoVrAA
Vwpy1alq0g0s8PPo4n4/JN1G0wFG0rnqOThjidkWLseQqrJS2vi34XP0Pu5vPSrbpnVweCoyz949
mhqYNZEDT5cJ9F1fQeevXuhzMGPg2gBHIBaZmyKUKo1dmCjlkSvnJx7n0oTf/br8YH3p7sI9rAfT
0MK9cr+/oG4e3+UQe1xHBFuws9Z0/QLKfMgZl3LZBt07rnUzz1AQsuKxe2x2au+6dMpVKwZ+q2v0
JtsK7zuzTAkHV5suRqUyNXXBDm7uPx3OHorouf51Ni7rd4vt//iIbZ4A/xathj/033IU31lc59+H
IwSM5sYthUw+u2Snx6154oUobccsNa0x2URbnPL6hYPyPfzvQmsYWCIJORXoigyZodHiVkyUmCj2
pL/gyns0BlySvP24Wi3lqNN3PFdIL9dt97cQGVd5sdnVi1lN2tvj5FpnVvkkGN3nFDq7gzRtPfFo
MKVP3VkIZbUJh8yP/3V1dvR16puzbvfCyU7jB8rCcJO/5Yw5qa7nUxZwy88Wqhbnwt6FBImrc+n8
+izOXvHWpLZkkRG0RdLIG9oKYbSNCMBLddTmf1+vFEct8KhNs+KdNOfPp1lK1DSDEe7CQmQP2CId
vmgm2IQsTYgQsKQcS2hPTq3qoBfMWEmK5348Vq6M0cH44jr+3kBkPuWZpfHMIoHZs2qOcWMUzj0o
v6qe7jWXWenzr9usslDVWritS9eAEBGT4GghS/ZygOCKkke7ANwBiyAtKY0b/PPeL6pvFgZWLcBl
fZ/7D539iO7zpRjMP9BQb+z89IPQr/VEFh0RpEQDgF25vaf2H7VmY33QHiHfxH/gj8qjvcupjdS6
N032aRVDIudbiw/wBBHol0Fywl+Wlr8qKPreR8IiiiTdripYYz4P7SKtt0pZwN8NMP2HVZ6w/clR
aX4NRUAiDkcIdTLKxkISTXH7rJDt754m7JRAaBzE9NUNQ7DqJwe1Cs58uHT0aaR661M7cb3mBKtf
qPcM+9JrNFg2rOGE1R+1gHrgUfP9EOVutTTGBxytdFRylNXcJK33dGq5UuEAnnPkUe7GzhDKDwoR
96RPwqBduO8q9YTOOggXzovFeyNB9W9GlS4pJJiGtjBjyzcMX1UCaBlWrJ9q3mvdgVmFbvOD54nA
LUS8p7fTEOueafIX76krz6srY3kv8z/Oaj6MhSLvzRbmAgJnsDHB7VZbHCku82b4x4XkeUjeXSJs
NHM93i/vWa8IigDpc1PVQr+Hg+CIEa0q8M2xwWkbaa0i37ZBzFOHXmbEcXt8sRNIx83OGclmy1LQ
nUk2CFeSqZPDpMRYxekO+r+YaW+KmCXZAzrwnRGffkUAwwULDalssKqJtN/AlRcKTQskvHmBpT7U
CrOTB09232cWXFGXmlbojPgYj5YdLr/IKjE0HSzj5Hg2o5lM0wZT07caUTWVP/umMi/lbF+Vidq4
eXMfjPs5gV5WPWzmBZ46Af2ZcvDgfE/gOwOkgl0evlQe8yp/zvV71Od1wg4YH566I0pSq1vJiTt6
vgWLVVGLjPvTVbCHNLfOePG7pt1dGUJQPU3CIkpkiAuHgjT3mFuh8MD6c3WUbMQRxWyqsDdsMpk1
oZ80233qS9ONJ+qMbf7itpwTyWQaxGdm3f/jd+W0oUkRDe+t6RJnyHEPUzUgRT/UF0rYWEx2XlRb
PoszT5wzlP1TZas1Js0lKqvolKZEz3/ysaUKvv7aM/ffclLjnVky4Xs7qI+c6rDjCmQR14UkhTYJ
OldSV1xxMq8RPZEBowjWe6jVXGFHyFpfvbUf2T7Wo9MZqiMFiGyRlGtHZI4fzTqrtpVTF3tfUrmP
ZXLF0qw+4C4F3369TOaajFlrddldZZ/U0NPsZEAfxK3aVAUkuEWeQ5za8LRbXeQUeBGnO0pwHqrG
fbRd/C12YMiCTOqErKPXGYP+Zw02RfstKpsLTMu7aD5NlRjlZugLXVk/+qv1dxjz8WZN/K8Vk2SY
aOComHrmpGNYDLKJhFAalc0BGzBWV01xrkw3DAw1LSwgaaMcsmWhUUGbUI4qTUcpCSC+ckabsR/W
ycZsIMb94hQ4MeH+MzzHq0aTxjW3sXzzNPDRCkeyFtfSM2HI5p75vxNiBMbJA3XHk6qXvHRnw9Ua
lESpeGdVDvHF4WhEwMXrk+MlMad4+J3OtCdqTwnIO/uiH4yzJTg4lUFyC+6QHlh/SOnzuWtLUEyr
ONBArbGhRKUJ/pkGXAavQXoUmOUkFqVl0Z3NVPlfgYpgRG03rYYWo+yXqvmtovkNKFHh2Yr2veHE
zaeSE593cMR47jOvmaMn1yDkXipfVabUA/w3KMyeX1KwqQwRRFDtm9//4JnOorKikg9+taE5EL+0
6MAH5eyp8aiGi2H0OjTuPTp6IBbcssMCz6YMTXh5XOLpj9//vza8cr1F+uoOphfgzUreg/5YQB6Y
ug0xsBd1+yDdRa3X6E7LTL/flYo0WJTq91Mc/amSgUa1tqDVwBhPaw6+YhxcMC2iV9Jx/lpXlQRV
PzpbPqKiv6t4JH6mdE7VZkv+rb8888OIjy+oczVka0vlnPrW8P/D1hyI8G5kXXgIlyExN3lZmsEk
vgtEyTsSr6/5MG2ZYe1JSTP58fDa3fX27lt87W/los3+jFrWlMRcpSQdyJeeq3JHnz8h43IwPk5T
7CCqyxPJqE9XpZkyHpoZDjmas0BHcqqm/pF/lZyxb/zr2fhCeaay68jnCZLxf4x0HyrlzG7SL2wM
NVQpw6/oOrSngXdSU/yVcqsXKDJTM5Cp1qflkVLLOsY6bBONg5k2XrmT11dTc9nk6VS29y0iOydJ
WPk4m7wV/L9zgC4jwiLf5YJciOk2JuyDCep1HgxNhASAFyQZlUHh6S6xTLZ2QgngFCUdanApNnwW
kQFPXXylZPKx/DDcRir7hQZLAsAzlNOyPOhmXqy+vctdyeEw0ZYln+VBn/bnqJhH9p1TyFtzLoSM
jc5gqcZpexI4jpstT7dbaRudkyVq6Djerf3hSMdiwHc2Z3LupcPgm2o1CNC9trQSPBHb+WbLrgfn
a91F9xYtzlw5wA6Zg1r+xgTsfXZb7IfPk1//1FHsCP63C6ScTiOoCkCCHtalqHZL/jHqrAQBdos5
tyha20lNRMw13oncWCEfpdRafhliBqTn9pAf/Z/VknD9Zm55RRJwtvPX6DM+lY22shGusZC9xWey
D3Xz/dYa7Fm1yK2nMYlOspAF9yOCN30K9jGCZBd8Jay4qEDbyIqt1PwUKqWoByPTiGy7BYF0rFDH
91wqyaV9RtgxcQxIh3YunwSGTcVA7oJ2F17FGkuGwRIWvZfagmIWIi/9e/8Wdu1hReXb+Cj+29AV
kXt2qoqkn0vpCF2bvTOQ1kpEpAh00d1Urbpvn9phUyXFdmbip9wQhNdBdSpk5O0/XR5LRuTdLd10
ZzNp6w1UfOC6ePzMRQaacVWOP+S+rbSxD+4l7PIq6JNXjr5luJ19Pu+Vh93T/wgQ0DbQzwq5JeSg
IJgjo8g/yJc7rjM84RsMF58OVGhCb6zcxN4ThxYh2D2XaJQBDY5NZYrqSv/yWSyK/aiER9bMzYOQ
0ffXMoFAW9S7mbPeLWZCPB9/trmww17M2X9WTMciDWR+E5PMCPr5jAPymeYHRrDp59C8XSkwKvGu
0X/Mqs7iykZGCdWfdRXurP+MBJxdT3CF5dcH2v0SbMdLS3huII7c9n4Rjc/1p5ef3M86xiU2B192
/TqyZe33Xp3JoWFxFT5GVbcUonB222SnmIsaxkTELYezUU1D+iY+mksHPQC8W8x0wCucaSUbGvEY
4lOKVPsNUBfSDrXEMUd9T74XhdcEvngJj5G+dM/ln2D3xM8cd2e82nvFzPpPcIYBPtcbes47CUBx
dCwHo7y2nIWOBOGTJR/Gd2YrF3mjzSCMTtBspmS9HMIZBujIiC4HGMeldDXmnD4Iy+Euhned0cP+
C/HmIDipHiLVYD6NI5aftNNQdcHKriDJZMFuP4pSqeYaMpwx5PcarV7SDYzleRlErhrN2fLRV8VS
oyAxY5b6Hv/h7j24LpMOMRrvWne2StS5aG7jJB5RmZAsXPQDPIqr2ocCbVNxO5JM9oAri3WM/M0g
wPMh+p+Pbma9zIWiZIth6boVqNHe100/koEQdvrZBNpD3MkDYWAlP6svCdaRIXaiEru4yLtWkwAK
dPrMAInIARjeX/+QNSFLumu2/PoEAWzf/NrJ3C+QgPENawI2/gt6J0ZVsJ07lNzo8bT/z6ycalQ4
P6Ytq/pXpWLSNvlbUYedOenvHl+yraT3WsnutiVd64Og3g4oNepCqwe/k3XvCt6+qfIvQ6iLbjnc
xpwavYy4WhfrVFgrZ0cAA1c06y+lK75UVkDQViEUJSb3X3r76pw9sDkeq6cBsB0EXPBj/NZdRnzy
u0YXTaTX5brXxu+Ib49ckfIyV8gnyTQEqobKBcPecvQiH02XqrCn53yd8Y7OjCVGdh5cdjYSM8vD
DczCmS5BPbpqB3oDhPLkGC/wFlatG7hUbsXs8PPuAUK6iXN5XwtWxOqV6cCRvD95HX6PwWxlHd2g
auRE4iCLHbUsaRlx/pmhmKm94cIEvRotiAo8QeP1R3HtiS371MgCo3a7qB4TEC1EU7poJCS2p9ym
B0Bjjyt/pnvVD9UxQdnxoMrfFiOuhF+BN8Ct6jl+8YCYxufvlLD+UMc2iHmUkv+15f0aTVHcnUCU
6Rz0wKw9n0du8RfcVakZg5VPvGk3qh4K8SXqPH/uzgL5QeL5W4CMA9mRPXNI7GPnrXPHmvew9aJG
X/6x6BUX1ic7/a4XFi1ZW+QYEyu2I64/mMjjzztJ5Jn9MRIVpTN3DSesXkOH0/ieYJj8HBMBppSI
uIvGjpr+dz74dU/yUE/W6wLkjMboUeYG9t5KI4jId0r14SyzuAd23k+3TRNzTyin3iPyk4rgzWZW
KG/E7HdjmbFM0z0hcCBP9oOwbNGkRNahtcoCM74NIoQhirvyVsGwbjz2Fve1Hf6lMh9rTnwZbfUD
2QtcCbvxUQkX1LBXGCuQml8g8agPHokLEVOlYt3Grs7ZqJGwxKuD2tOO57QGcrKohsFUMk8QYaCU
w/kzdNOiuerqx1YdwX8iSb2LFXYWirG0sIH9Szok3p0WrvU+XzembsT0Oo/8qiv/f1AlNCFBUJ+9
BAHO1YrINoEUQmw3wwcjlQR9ycTHwPTaPk1tlnuvKnPJRsILXgfG+cODIqeXbwghwCEoG7hWGa/1
b8no0YvbJRDnAH5rKDaQqpmYFiMYMyBpNtgNpmfvo53J9EjrlZxiDFuHqaUQa+G6Kjj8xrPpy+h5
GRF/8q5zjdSA+TKiq1RccSudc3iQSOcM+KZjY0sqq1QXd8Enuq/2Aim/jeedUHqn+UfdlbqrITXY
6FZFP28Gc0+UJWZC1s8tkrc6lTjaOT1VYuAnhTORUnjTplRdHoPoyX8AW+p9/8S+YN54iepD9IKy
ED/WsV2EVTElIo8mqwjqeRTtjBrbwNh38aByI7lBRVkzJLrvFkiwgXgJRJeCGl5LC0zDTAzFGz5A
KyPdehdLqs6swWkVhl1n7KUPGl0v2GriQQnrkgS+khTuzLBhJgPZGWWGP9v4ZZeWH++6Gw2qn/zL
NTOfuLdOt7Rs9aA3kmxBLfe/vvSoHbAWJVBkz4poW1It0iK7Xkk3+7EnVc9lQzWutCPA3ZLjpTgL
f9HaQK8fn4Lbc6c0fdW1eyEKiwpGdtSGovaUWgrW+kVYwHNRT/Si3d5coPglMLIer0wmOF8vfH5s
JGTJ1j7go9ovSFTFl80ztUfGSOD+OmtD5kXO5kOCQ9/jSLRNnnf54gj46ICa6zloMBD/6EcHjrHP
cew5amPXpIc7xkv28FXzzplZDQwB+hX0BjHFsK9qbpM4rFn05BygwdpJAbc/1SkxclPcD1bZ3nd4
CZkDfgAc4kiyx5fS3SchzI2r6BpWbYaPf0Cp2UcwLk6qcpbtuMw/g2qqznbqWTNbfRcpuGlGl3IY
VngvnH6KmU0LEEjOwS/bRwEfXryeloURJ8XcjG0u+bCUxAlDXiw7mI0901W66wtqOZCqK9iBUs3F
UPqay/i6JQP7nu5M+Jy65T/0zxl+Tmj8Wj20mY7rPQKYMxAFiy9ySxJ2Tph0BC3ExEgeUTkZtRU3
ubLSAGpazzxLNfxYdvHhc2zNv/19FxQfaVP8WtDHJ3mdmAY2uEvFv42TCHcjRsijBHPW7403hju7
naWoBqTqITk1O4VGbm6Aq6+01CsbX0ZL9ElpfHUgR7Onj/w0FXB/D2LevLZEAvMoaHhk/W+Zedl1
Pkj1l+5W210QQt5xAgDDa2gm52uNbNM9lEnU6R5IxVJCbIUe6LPpgcdUTxhwPWvGCRT+K1zpzYum
Au9Ye3Q8NUlWmaBrk/b5Gtx+ZQ4avh5kUXTXL5Eb2J7MVc4QfFFNhr6fFHwnHpzDkkiWhIIXBx1u
5b0VT43NDlZzop+HKeiGHnzDpcy8yZ+W4xowjnK8eWANfuZ5CdEgZbuqU2u3RQHTW/01K4/6eZxs
jyL4P14aLgMd9JIgKmx0EEw6yI9eYjI11XxWAsuxoTCY0gCfROBtFNAjft61WbTxQNKTiCOixM0A
0G+GvixoMabqi2lObZOm3DH9bO+r7myvsYe9qTES7jpmpnZGyo3rYG5/QK7EUTpuH40isZubga15
dgNsTrbmkefyJbbjw+tRDMIP4aTj9kpM2ag9Xdfuz89y4VgMguCJ2HIHaQ70jhsveVUuRSi4Lxu4
ZR3K+AMHvg2Q0ErP1qxr7K31C9qJH8aKnrFUYBU2gUgBgQLBhik4HTTduD6/x9YLGGU8OVj+jRWE
aTM+ULCJB/Sj38Sc8BhhQus4jJNSkWMoQjc33Y78wzbJH4P9GkNtrKgXx8Q/OvyRDCZla8vOvBJK
ZgUam88+0ioplBx6UVY0gnpzRU0QiAw0uPRoPqN5tl/NJ1JkWXmBCQkK1vLDsX1PTOUgUQiF133e
AkTO/mY3baFCO/oYnvR2E7z7GJRpjWxBlZx5Gm3Aulb9Oxf8kNKimpW4enz3AfDSw01hITUDhl4A
dcDNyGxquz7ZMLBKCtAkP4hMV8EWttoRo+Hy2IbtPTUGGgUFUEuyVu0HoHwLDpFDqYksyDLYIaOE
CD0KVLCEIsPWNfiQgqb0bLRh38lZKTo+96/aFzqAT2CWgE1jBRn4IZ/yjVoF1BXixAO1SRradAal
+32SbJzCKVi77iQKk0xnCOC9ovGCB6Csw5AddGuOw64DvbcLCw7Qi27NcH3TBGr2xdLc9EZbeVM+
2xy//SvDNiriTyE/Psb3ryDiUHTFn8HX+sXccV1TM6QoNj8lWeJLsjwUC9mIlw/dhp6GdwtBK/UZ
cmZTFfb8mFClnkM1Qiqe8Lndz7ukaRuRvfrowFHWSGLE0DgUoUX2YiuLlf4SeDA0lEh4sHmUreZK
ae8PP0HYVWzutM6Xlv9Qc8G8OjHHtNPMTcWeqAVrzdoEyWg5+HSuRw3n+5TXHAIt1tSYBc7Byu0F
KxxwO12WGu/TLwvV996fjXpsR+jOPZaoMiNzNcUfDHp7i/OiEDuQVLUvtxBAGwdAeYGc4pV9fRw4
a7irtkvYKM0HjUzZ65ymZgIwd6ZnEIaM070KwxS3Icj/QqhZRkxgw3gUOP8ddboHRB/kJiqslUP3
Bq/yjid0ZieXbZwq9jHq9NCy/SsBOUTovc9jmszZ6zQ1uKb/F/c8oZiDlOwRwc2WcBfXRVXd4Cq/
0ocPYfLRNPMjS9ZK9/N5+kS4dsaAzb2XNiCFTtinGzIncFfh7OU1jAFA2a8p7qEQS1KcYJzkVMJz
MQKK3O3j6aptIOBXMrvnIWV7mbBJC7lWBHg2LVyIucj4rQxmGUZYFC68vo4nkBmHXgf2aN5R0sjI
gJazVvhhDe57dLvFWqC8WlVLVvHFvd30FVcfcAwCSTpgi2ZOa8hRpB0tnAdn/y1NY+zxHySfZ0vA
Hy1X+VyinrqFOhczmuFGJXwysF4vaJSTImVbNRRL0O1Z03a5d53UO1iu+pi0Omg3qTOYJZBmD80J
B5v66hHpmnOGA1CR0HiDYq1fJSdINr6AtYTo7bp3c68/wzQNvJy/LxPLn44OifGRfMuolJ6/iaUj
hfdx8dU0L2w7l8nc98DMrq8hmHG3lexI556OonGjKpTO414IjnfiWSNdAvS3pg90DwdoJGygBbw/
ehLPBY06FVp4CWJ4q52qvzxgw03w2ef8cCJ7pm4Bm34gOHXrbnk/5CBU42va7BGfk5LUZfteH2BH
bUbmsXkbCY4eH/drD6t7MytjHod1Rd9xZ/ssuyXpV6VrSSoALtFBPVmkKuhdWbR9CJUEocuyFX65
P3d0vDbwe0aeLyv3TgaLluBvzyF4DqPmHstLkc42QyChBveO4CyCZO3InuRW0jFg3mBfDK1lVlye
6cBhYjZsMSDajUNk2/TaUzj2JP6jtKENnE4TZNnt/IH8RlcrS5gbdnC6vFUaQazG/hTgsSlWmwQm
jflDGg582LxXEwwpkcv6bqQbRK8QGq43Liqi6JR6PZ0teMFxGGd8sFs29/HrWPc937zEAcXRd7vt
yOK0fLH9qKdN73b2k9YVUSj1qV1L57cxEakefwEhHnhDpxrRablBTuINirm8cTR6wRSXNbiNNXVA
4uFhOjvTVw6MhTP7lJ5HppflRlHtSwPipnzHx9F5evPvoIwdfHZCKI2oLud+7Q35VyrX8rxxroDb
iwREFaGwZeEichqX0M+cB3lpHYHaBBFK9I6I55nXShnqSclKgVL3bhQSCXqIixb78xVuvn25w4Tk
p6hbdR5ikUYqgf1yYppXhZbSz/VaMgstniCodP8nzXir1De6muMqYWPbkONIggW9QuQpSGFrpGsL
m66cgogZwHCzhMkZh7z4FkY0gWKBB1YlWBHlh0YTckYxL17QUZ26gAB5CQXjwC/k6Z1F18YlxBoA
mHW9N/CUViyYwVP2Onux7h1oWcaMCDSJkocbIdpUdVtov+nqRGLFIC79OG/Evi04e+/A5l0PJ10r
X/98aZoeyZ8p8wJEzswUHncsXsKDz+c+MieMD/+E4AWSnWkwD7lB2c6S3Wks/A8lKNB4n6US76ar
1x64WvwNLtnBdexa+cgLOEwO9dn5K7PRfXU07licyYHmJvjT7WDQ6HyTJC3JmfGS0cpVI1ifUupx
YF18xwVm/s2QW8i1l5YPpPy+r9T680PoUtNc5+XWoQTXoPJKyNyNjXrdqRWjLZ5DCcZH6Vi6y4ho
18insPUo2tiBQyurkFL+Ta5rqEARE7Ix03vR5y7Die3nexaudewuEIdxXuYhZt8MIqpPC+IVBmBE
NVvDx67rBZw3IeHgsKUcnhKyYA+/ZFfsPFsa4bh8WOLWotV1FT4c1yMWhcQ58wfdOZWZX4rXTDwQ
bxPDJLpBclAinJvuA99FEm6+2bcDY7S/2TIuzTxZ2XMV+RZ0XtkaVMpaHt+WnsNpXghYTtXMMs3b
Ufe810DIg3hi61vyw5TvBAQJe2OXt5Yn0CXQGCWHisNKkI4Izy5qLRyuqkC5Qt4ZV23KjnEREwZX
ScJeoLlL+Tg3+PSYdAmae/p+x0WCLcW6dLitRidejZTvpu/q7VU3CvZucoe0GE32r8GWjXzGsK62
s38nHxmc3OpgQSrQ0THdjgpTGcCXrsDrK0dQhAVr08V9VOXvA5aaF0czoT3nU3RBLpbzXo1x36eT
AAJwoidglpX7lN3Sk8T89a+5zmrG+cpo231TZrJsGtlccUIIcT19SpjAhaNPnr9oE5FqKet1r5Q4
5IVnnMMPuNb2YE45/qK4/+u1OUVfg1to6Hh/dfJOKMbXGgSAX7cLw9M7QeBxI+3Vznel8vL8Wfxh
7nbUKyTU1vItHxuhp3CsXRQNocivQ9MBRqqihsE1zBD7J8sUXkkFFdSncjlGaj0XxERCkWG2a6G6
+K4uM9rgEcQhPRIoBJY0q/GB5P7xfx6L/GClchRZ0akBlMx15aKGSyIOagfFL9/DABIlsU3EYYPi
lbOJ6J4sdNnlr4vKKs9AtGP0LBc6qZSgtrstblfc1js5FAHojzn3Kfbfw/XFQ2yil9MRbXyNBfQu
WIX3dx0vfVU1j0Aofk3PX2u5rst+MkwPZd0ubTOLdSJN8DCXRNlrYn72douXl1tY7ya2FDCq5bjZ
T9zwRw9YFHAreNQha6IjAE3F1ZCnyoNB4MJqswGa+ANDp+TOEEQ2DFOVk8Iz5HZO4jsNiXOSzx74
SkyDvklovtHyNGC2wOoDsLcLQXKGeWewok78kp2j4kEtgzboaw/T6Ggz5UK9oAhI6S01zrK3jWQ9
42TgpRo28JQ/qfZ1Phv53T+fvO5Xe71zMFpJccfW41RdbIPu7BFd6pl8rJtML8AygMcA1d3/e4cZ
mpV6LTEZk6iY+jPo5KYFLNzqLY54RgA3p9QW5q/qt/yu9Gn6xEm0jvLAsC6gOSe2PCdyZQe1giWv
+SiqsPMIhIxZEkfTab0UN8iupwcWCNQMNnQWoD+LEKoMlsa0KSTl86nTUZp5JDr1EDxmaWg+3L3y
ZndzZmnZFE7IwDBcpSvf7T+AJNY7JTfqDToNrrg+CB16n5biwfrU9YZ5HSI2NjSW/Thxu5BFNfWA
wk8sa1bl/lwDnXQZUu/8sXPCkq45Ic7edVhBvnQDoU/B9LrogukBe3cSA3ZzWCHH4Njv+Ovm519r
fCm6gMVCiGsVghw6AHG1x7OcrbCDFLAOU8BnpnXyG3sLmgLIh/7f83Xi6A6K3/L5lhOA/a3ugNuo
cWQiPZ/uZ891CY1uraEvK6droC7Cc0ZTMOwQuqSdjCL/sCbS+D4m5jlXWeBHkOXgFw0RLi6DqWtm
6/QzWknwDo+zrMjULGwLiPi8tfct5UUFlJlxUAa1sHvto2TvmjiwKFBNc801YWGvDyoM6Wl08TQo
3xCEcAqMNGTE/X6PM2XEBliwYYM8TMccWjtO6Jxge/tE0QYs8WD6YlpOuhfggxxK3VwEmVwYxqMq
X35aN7WzeDvZjQRGdORmLDm6+PIljLs5Jjb9yyD3jlBvI1zWkJKdvhjj5/9kcsru3JMNHssadR9s
UP8JWW/Phz80WvVfBeWHa5N/lu5C/1p8PpXCa1Q4K70vyW71mRt3obGmfCI607kF3FQoI/a/xCzN
JyDdxJu1UoiYQgbattj0vbITY/HbQQoiXW7kOXdDvzntHDeQqXV/+kEm9WcsgTrjRlWT3PGlnlKm
pXiFQeLkDlSRq4Ovt7GwjtEqWCnrnVqAmkxRq8PyWGylHOHN1niYSYd79Fu2oEr9dHCbjIk1S+dF
R6jNu73/YgEUYKptkyhuCH3OT1+hQa/fr30vsxoCTvukwyS9YM9SNlWLi9hGelpB+uFhI8pcxhW6
yaUocAjdEzGcM5dU7XKaH+wq1zSrJBGrknyTXY2HNujCXeC3/PUH/sX/YU1VL8BX5IwyWfLOLADs
EQNrJHG8fHlJk0zL7lOlWjTN0KBD3OdDS/waIDhG5FBr3f3VmiT7BOWLsJ1qcozSqhpvYSBttOs5
wlCf6HkO2i3cdx+zaMEhH9AMGZJ3qUhf5NMlVLy7DVJYcM9Quhq17DFEmBBKpqYOJk7gFr4ppSYe
WorUVNRbOr+JtY65YyCV1mBv/yX8M9GF5Bpbpn35vdvpaOKNWSpk6vr4iN6qCZZgYuTKRT5BHgQJ
Oi5IbdxahWLehonC/tWrs7F4z5ZV+V9obSooymbQpWdeLS+KOlAG158Kf4K6wF3/SwUOSr9/vLAR
CxxTbm1VSEJZDLUQMsNPlO8Gdqisib8LNTx9pgybtIzfFkTU6ZdY1WCMV0qcTqLYWGkNnNzpINhZ
qFyAGR6ya8UbuFnzbxO3nALfk3WicU/IdSHZfGydGBZmDS9jyM0aNPm1qVfc0oXcVpeG0VN8LoxW
ZeMBzBlGCih3K+Uhzg0kbOtCqOdQFjyJMYZle6q2idFjAtztxHK+FLUeSL+8wHhWXj0aSCNj0j7f
0bCJE6zSrpnVdQJbZuDJqazmqPPIUl+qYB4DsOhJlzvdxLia4mQkU3xjC7n2BMMCG8qArNHJ/U4b
e+iW+hRBbR9+lkstSR5D3aP0P8p6ltJ9BHxlgPjIhjXp4wUFhzcASi5T7s3urZDxX+T+v8dJl4W1
n5kOeoH8W6UNBF28ookZ5iq2AhqJ4MSegN/nYsyin7y2+eGGpLOOIxH9yInmBoG5ezxy+aTDkM3L
GU3SW4E3+6PIzuybVv8VBwiP2ua2qx2haqa6zaac9AEusIFn0pFQSawTvbMWFaWp/b5Wl0h8XTy1
dfe8QSVSG04h0aeOh57fibSH5Sv4pvNPkMz/Z0UVHhyqXpCLJXckWodfHpDe028ZKr3EvFixDI+B
oWyIikWi0sXA+L3OhXEO73FEABKSWUK4GVKUl9HMw8UpWF6xGi4D936JXbYX4FsGyPqewyLsfG9+
QDB2l45CsT+8dw6d/heAGJr2KNGe9rRsIsg9+1xjNnwG0yg1ZLuxtZ0UltffXxvPFlM+vIHJCiHQ
aAfxu7xfBbl60IlbgGft2UN9+lfX2lZtYbRHaVz2V0E0In9T3aT08h/sPKZlAAYJ9bc/MOR9qCKV
rAFP2ZNpO82+iaLj2586A49tTBFuj9fE/tdwqE0cWNzZ5hC0h6gXUoHCefCpTA9dVi+clogN3LkP
jx7kcZF0SwUy/UnRFVxTe3Ul8gmitzukn1bsd88zi+3Evunbz4ngFNF4HQ7/KKfONU2upthH+pui
A/g5cI0tuvW7kciCVbyWGlxIWP0YHvM4e6+Q06x196T3gEhgSB5HFTcOux37mGFpvXFWuL2LSMxR
suxqFxeqXwqbyuC9+025NBFINJTqOGTc43BIdb7C/g2Di0mpGorJlMAYOqI4f5ZC1oxFxUPYD6iP
ClnbYftOA39gvXyHSfd9bw1Sfpxcu6FXOOXNtdS5xPMprfUDguuRVLzbOmtTd3lhGS/KNDBYpj5D
Eg5XCFP5q3WLcRn4FZ1SAnEiOKi7Y51EFc9xRQh4jOys96/PYSrwD1X11zTYbr5jYEHtJNLEpjlb
FmIX/jFop4cj4bJ0iIP2zngiNShCwwhWaCIfbqJIVNCE1vYhrGtwW+2KSi12z7hoo2GRhPlFULcC
BjtbyHPF1bBEQLfbdHEufD9gONWrcFjlt2RKB0bU1pET0Eo3J1496oTdgrEVDfhr6oVtngvMtUYv
isTqOS3V7mwZbO6PKrnve3X2m8Y82TZ0Apvhsmh8cF+qo6bDExQmiSJs95qNnxsXHolUXRZZdZZg
x/sdvL6u8vbk8SERJaJ9zDOGy0vX5TowL82RlZ4TTMzeEZcFDaVXoWn5nD/hI3QcmjEsbdyed+ja
Fou873XhKQyRcTTt2LApSixxYCtIHPSbisy0W47tDOs3oOVj0nm7DgtP0ES8AR7afe/zXzKdCBIB
sG/Zv+eDAksrDcTFbzC52l8dOm2P1X0qySmdjmY6/eEHPGXL23Eg0qJLPvjzERWbL2pPN+zUsGf+
oO7O0uHt0ndzWBGmgsdFYGz2836FjWlaQ4W54sb5lph0CMEB0xUU0YH+ln2ZXlHGOx6Qae3W2cy2
2HesZpptWCNR/bnxcSUYp52E0iwdXcI4WsjLkO4HEVa1cfJ5Fs9AA4ECdZ9JTYZBb/IuQ9j7ZYJ5
XM3SlgJ8S0lirv82A8dqRrFt8ljLYI+9JhwYewYVoZMYOF77eWxSvNdxm4aHeXO0MQ2P+NGvtle3
hZ3s3+1lq3EVjmacBu5GgAz4QoEf7coxhTpX0PJ5VOdKnBPvtzmAIAj4RD/yz5uF+UTbL2FyuIWT
kcL27t/mXx4g1a/kdRW/L8v2xsytoRTOLR/4Xrh2fgMwJtsVo9nTsQn/CkcvXitDWWpijUtPxeUg
S2KaS7eZ90iLo14TtkhA/YhDdZI8OzFDRCfy7DqhlrHiaEkJtNosWusZKSNCohC30P/7eMC3Y2/d
Rh4antosS6sySK34bEDLGbBLO1hle/3DThTNWTK3LFnBbSA1GOVLuSZVb3jxc28Kk0H9DQyT4U9q
k1vTdmvB8TIXkku+O7uegcPZCAH2uawFrRaPcJ9dOMc0LtbYtR0H+Sn1nZHLdy8DvjKWNBlaOcz0
TG2ltzbkjwvsxiTdntxNSsmwps3QsrbP8YEaAbzWz827l5qDUzGemZMquidbDm3ZWnPESNJP9sVL
WBqP+yBCXiViA7FZWh9D1NeVcDm4yagxAQA8rZsmCBmJoaxr+2exjY6eBLK/hipYg8SNKQFT+BkI
ZDNEUcfsDvbkZgECv0bh5eZoKmBi8at9UAuIc67uDUQg6cqt/g7PqqbMwZh75t/oPUakmHLMJ5gC
/89mpwPTssg9ZDha2nWvMmeVFm8Q/WY9dggQT4DAjtXbgU50rRD75LFC/2/PTrH03jOWhQp1JOpJ
jMzMUXlt/V9f63Ew2kt4DL9fEvYeH5cAZcK5No7+znJqtBsF2yPksqx6CmwqmbPfnyinFAnbdbhv
vdOSRdYvmW5+xie0gwD2zsAUWt/KDrxEcqSRKjCusJJqLTdxLahZJFTg6Yb1Rr/vHQE1M6RDwPv/
Xm/n4IN126ysrFYoV8/+2Y/pDzkOBQGzTB+5tvBsLOAjWgq2WDwxzYrg0lPe/Tis0AXPryQ4jc42
IbqXhfgAS9xJvD30mcY9BzVCcIIlKyrLJD5/GMmfSngOP/iqUasP4Yoizhuw2Tu5Zxik4GRPt1CD
o1j4Nc3eDrQHDGS7MkSpU/bZJOPs9iYUQR3B5hMyo2jzgU64ExcjB7uY7TVe07SOewiAxVmXXqwl
q0pe6oXTCsAfWWRxaW1dIbeVeuikS+q0dwpYG/4xUDX0SPsKKCEGch+wqDNRhD8ovque7ZWPGV4e
nCBd6kI/vs5P6SHnlSkdGvDiTjCLTge+DkhA7uFcB80cdsOJB1sOI7LAkTi/zEy9mnJF9M5Zru5R
BmxbgLC6z1KYLKURSsohQKmSPdQmG40J9XsF1rFK0TavcK0B/aBjNMc+OpofxMQEvaASqP3oaear
jI+Rabfmsp4OrC3PNiccBVTZ7rox0bOY4s6IGb4Hdya3a4sAaBnXuuVwnnVflOJTYSiNKZnjl7zO
fh3UapL5DfYZVLfNJhCpuFTBycy2Zv2m6CXKeBTm48tI5R/IdpE2EFJ11sZSNM2qKuDC19brA/pZ
wRlN4v3ZgrdHoBi4CFGqAcXWpYhsX1N1e6ZnTvg+h6sn46nh1pPSOxjEm9pni3BH6Rqb4MDH8/vY
yK8ouo1obRsAZcKHgUcnzgUNAWFaiNTegzIR0JEe6WNytL7uZh2Brr3fCjpstKdpsc36Fa2VRAz9
wHaba0O61l+n5OkPPMRnzvC/SNs5ixCe1M2st8qD98uHC5SZy9JviWTPki6KhLCBge2McBTYergn
tWGHNbLvR9Q3FT0bpktxjztJ8f9/10FK9gSZZu4byGTKMWZhYfqN8+mOrM7JSqRkq/sSd77SF8cp
FteItimZ3haPmul+/NN116/JldUfHKKPohx7iYPeAZZn4j94ge3kCXH2/gsoVB/59vaF4Pez/rus
Sr1gxh51jXf0LYYWvn3OwAIlvx2InxAFxv98MBvHlA6FPfEoBu5NrLBAS67GNMd9Hu+KY5QObavh
NlBTGktdwcZ7jgPC9lrlW8f9LSji2l0anrKzplK2F7iSu12N+LnMEf/QO2dH1IDdZKGUAMNpGzLI
NvzLvfZXxlaM5ENXHejufeNtzFEd5fd/sLs8uqQR9CAvtTbLOdwMAOMErbr9hJBdnZi6gk4qbLQc
/BSy3l4GqYISJN99Xs0mg3m1G86rsUm3UQvgD8RFQcib9NurgFIMb5vHMavpg0Kt67COXFusGA9x
CS2oa4rp2VyzNhbVHe3wTsCNkvcolV98TT1rl6bte1gKSWSLJvKwbysA+WnzQKWJanJDTmTL4EhN
W/zxTP08t5wTiPqJbPqLRi1+dJlfyFy/81vNMebCgWIpeLNvsbqDlSjwcV20xASwHCBr4og3HTHO
V9J6RvaczwuNng7IQCFEeQhTp4y+SwZ+8Z0Yvk3bWymkPNhqooXZBYll5JNlasVhn23PMF/ywT9W
eL1BCToqvcbTNIMasm2DMuwZQU6D7s5efqARrKb78evaHq8xCewyVUk8+TrQF+woG6Qad3S4jOaj
gRExNbGDTaAKUlslKdRturTUWAcbWs1cT262o23aCmyUnn2RseBs7aVZHZ6I/e1+V9nhJJqhChG8
XjOUBcz0hRuA7z9Q7+OT+aA+paxhBGA37GOOn4SCV07Ex5Zkpi3EHps4jCBuDqL67XgSn6ttz8S8
wE2DNYB1F+s1GGwsD+BF0zhiQruMQqW/KYARJzCYZo0GDGaPPhZ0RLwNkoBSKSirLDiO70My8Iv9
cHqDqdGwrcmlGab/5eADO9gtw7C039NsJKzkI68GRN1XdALaHbtCfThRMkQulmBfv0cp3jp+oxQp
nTKV2Sy+Si+78gIW9JilF5nlul+UJiBVlaVXzgzf5/1A49wpAsFsbRUJhAGt0R9yhbApWaL4XT2j
rSdjVLJ8pLgzoCRs891XlAU/36gfkQwXeq152H0w5JVkliqk3xpNWaAM/vmgfTVk4x9BR4kCjN6f
E/HuRCPQMzruFCh8w+tCL3UYBmvotUpVO/vaQ3lHUBpSHZYV8dE2l9YNqUzTmork86r8iUm5tFrJ
yN97S27U2xG8KnbKlGxAIqo3fEzIUOZ+rKJwNIE/CyafrhPr68XDDCKVR44AXE9U20tr3V7Hjf1z
7xZ1IRJZLEBS8ISkS8wiZkyDjNhqy8g7g7O/uRpR9PWsm6YV+icjOXe+IynsIM5PL4d+jGmCRSem
5sSjcoKbuCF+oVuQzO6UmXEq0FgXTIGbOGOMOegi0CSU/eZzHdv8NjhU0yotTxwxVwywITAIBROh
iu/JatQjl/Lj61JSSvpJqCO6dgZSGRDh05vysdTKzgJmlaxlnrQkEJGoBw88IW7VvYtEg7bmKsIy
rKjQJ5Kx9Uw+Zc38iYZygYMtLkzWEYYBa37c4QKfNb8J1lKjSnrr9fkR4GrMrTSvqhuFYnyU/6Rv
EBrkojSKqr1dr8KQhu8g/lbYgXf1PxxCnlIDhy6ky/owMY8EHBAFeKq5QFVHFIzasibKNOGj2Ss/
an2FRJ/Oxcu/bv3Txej5jYiv1qxiAJn4RXXBM8l5LajW4/6gH8Z1eJ32+dAGCvPSlbg9sasLwVSd
73XWlt6GMoAaX8qOqQM38jhB9z0KOs1++QqH7SGD7VgfO6cQy96pscdhkvjlToNKn+Ej8hxYaY/H
YHR8Qz2zThjplqg3GGuDf+bHQxVGKQwmNwoKyzLXZzKMqqlL3V5F/C9GBO/0kXs8esSxg8GW8Rnn
wcUNFpTcFcmSGSVM75l1dOpsydDuTwWpyD36PruCNkiHxF5FaW0MOTkGGUD3Gv8X5cbIkm+ZTRjK
h6chCPZcqAdnMgXMSwhTU4Izfuy2p20EV3gIFM6r/JF9z+jOy6BdooOtkN2mI5v3z2IsVlSotvs+
z1H3b2cBQrUZMnNOdP/rRU8ONm398sMRaJj1YgkGFPz6KNpb1bu+Y2EgPvwJyLzvoWLimd6Atovp
ImH37lDBvtyJIE+y/96mraNoXd7uAKl329MnJOwQ0PeYxuDMIuRb39JjgYeMPbAmIF0dQbHaOxO0
32f9tD7uBZyhB0i0NtM2m4NDSnZoe5Q5GIljcj9Kkd0DjWsldiIRXBHIEnib3PPgv9TDbRD9DnRD
XHCIMkjB9qEqOy8ke1lGOksLt7hB4CvNP6XqIKlszv/StawtRDjcMK09d1KAHwV4wwpn5QdCPAXY
UyuTP4myoUzSdOYzMQCIyp87P4r30Kr/peDut1c9OHVMxdADjtc9KDxfN36FUaxbfieVMOJOfzBf
nP6kdZ8HeqdHGK53Z69ZfeXNWxw8HcMALJzw+4a4fvM9Vi3v7ScKvmrFLHi34VO7u5D7pd/8Mt0o
oh76khhNQ/IiJml9G4HbtUg4Y3lQKVsxDt+6mVBi2ucZYmoM4x6XxowpJDcUcnth6g6SJ+Nlq6cY
w8QOXbk11DD0TpxrqurRX4b62g/aBXW0Y/NZAujZsDVsHLILL/LniSq/1FrILQEHeZeRVGoDe6cB
aWcXYV+5GZANaPYELluDGvcwuVlR5DzE0RzIavKvO0j31SfYJ+/IXlDRdYjyZxdf943dGYiZ7pIu
p5sOvQv/BxyHDTwOrCx8y1/cYkx61epWugvVkL0/w52uuderSk26/jo5mA4Q+GuV08sK1p99qKhK
OAuQSKUa7W1TPn1vcLJkobyGrAER15cTarpopRkNP2OPDTV1+90+JIs4RPrtJntAY3jXwM2AxFMU
BR9xq/fEgols3pXquDkSFOiZ493ZNU/iTG7y/XT/9Hkq0a/AYpCySLFugYefj3EdF4aE8Vms5wFt
TQi8gbXoLrulPJ42tsNtvLq72SNdzP5JyYk9pxeuDKYt3Ez3jirgMPrfAY1gpEX4VVkZB5V/WlKZ
+M2ibUZdK5WVHFE8ajMeUYtg2rn8gu4/uRMNIuWWx1wpETT3R0KTX5E61+4daf/hWu2S64HTQ2OQ
goRxQcJipmLxqh76jbU1jN6cHuuo/4r8Ym0fQN8QdB4snjvgdwdyTIeTK9dbJ6Y+5Q8ofyV/fB8d
OwMw4NPdVaEdTGopU14hXdw36LxPxR1d5zvSwWqJKxu91dxGUZLjkt8vBffcoReNtDruJbAfV6vL
wJjvpoR5Q5PaCD+8NUJP7nGKhuwCC5QUubYjvvKkTTXijVpZ85lj9K2VO3Dhwl4zz/n3a++Qzlmi
hSvslBciNrDXQVhxaGb/3hxi4fnIjnWNeVU4WWhtx9baLLQXA/eLwpnWIyW4R2RW9ek7Egh9d6nQ
tpuHt3hJIkzi8VWF0w3+lOhMWnX1K5L9xqtoUKaT0xWhIxvbNR4j+bIMsMq1VU31ZwoAtYGGAovS
2XPil7Y/Ra/Zv17TnGIdwRF6TYtuJrpp+LJUsRXQoZQF8sVW49JjrGsl6EX6bW6kMeh9Mp0OBCya
S3nbxfjoUajG75sPQ4s67gSodaH8g+jGwE1DOYaNRsnSmgHn57qXT4qAPDEHaIlSyBF0aSX1xp/q
Rnz0/CIyA3XpAl3PrN3PALe7Pllo7osLn8pBRPy4+YJIU8kzLN384nkXUMeD/WYDUm+I6knDe6MD
WOxwERNXBz+16CHfQPaBAazBW+0t80b0NIxuSSO68e81nhqHHUKlBb+kqbZq9iEMFQ4hyvMaoSbS
czLSvfh0GxrZ8JhcNKrhkZP5xBdhRsnsD3FqwHGKA4Y84zOCAWnrlOjdtM7CcZ+/qdUuLeexlkYB
ZmPqGSJOFxJuvgtPw2NgeHq1CdaugVLxbO9iWsHQDk51Ydq0zUpUA8o29HnQlGfoSNLNTi+bEtOd
b/PLQ3pzlwWV1JMNP1q1INCby6RUdplpY3MbcGB+Wy1Bu8sjvMysp+4xadkwo6P8GcT3+UkWkPqO
2op88CLAFmeTiKLlfYSUf4bhCLeLB59FXesz/Z45wy4sFXaUZtBfpIgULOCd1Fusn0jujV0ghRgJ
Yl8PaeNnpR7oYJiCfys8f2bAnKCVLF9WU2kqsnFcgEd9dUP07bW0cr8xMhHKR7rcqSzJG9eb8UQc
CA8heqpTxodV7kMx/JmkGnnoTGxRblDyTsrQmYXOdTXMnpnfZ2LQ5vphdKi9idP//i07hEMXfa6f
6pUfrJk5rLZRcPqqKvYGQvO7H/Da+w8CNSnc4zu30lg7IhTyLduH0efN55lyKaczD8tiS3njPrp0
JeRiVWJ2D+MpzY6BV9N8nKfx61/LxcSA3Z1ClZ2LYt4cHHmAmAaUy+PocxDANpvUSvDfDxuhfEg1
uxPKq1ksOXxIKtZuSa9ifGB23QN2lxu6k7Sw0zSxsfLwB5WV/g3XldD9YeTTzXVYzsRHbKsm9Y8O
c8Uk45jaBlNK3ttN4jgQXy2zkgDYRfnQZuDlGr0bymKPQXdEETa/smQrtfV/9SgfGL1yB8JEBduD
VfaHZtdLv5lhRXFHbhFLRIfL+3e2Y8opFYmt+5/TaECCBOLc4+6chR9YOetZYLydTC0FE7TVyx08
eJ0dnzkXGAW5UhMwtukG953djxQehHAwUr0QH6BFwEkk6xgw+SoxTFQrADXNiAXLyGlF68qpwaFD
qsSg/+fudjiEhwo1o8i6Op5GNBlCQVGuPGrQbrp33WY+4yx8VXHPV7JeDsak6GYv3iu19JVO2Qzt
VH9qH+A0yBafskWPMTZ8BuYi9Pod9CKeBlkfkraBkn8oiqFuqQhnpr2n/obIcQJgEO51i/ZRROOQ
04PHtCiBtkqgs15LTpxEVXCYvSg+bUDHTUGUAswXEXSz527LGkI/lKusVI3AxvQ/EaEz9rUcXJSA
o7Hp+fgbaZ6yIX6n3PEgdBNveUnJ63SKbI0hSyjdsteZTgJYkjgg2yUDo2GP5RYlMDGIpdmlkvIh
coAba9IJ6/kP41eP3zT8NvMw5z30o4gIOIty9sKtsI3Rhf1OW2OGyBvq0HoEbhTbLO8D8qUZ/gSy
pUslIGE/H9j1AKJcEQ9bCPCKEU6o2QOmPppYPvzT0xdocszqi5VtwK9oxroFyMnJgkCgNhd3ZPHn
BglXGOISQLzVyYyGAAilbhnaI8EKue2B8gTUsbAHlzor/H4+fJhp/uZlYIg7KjyEDW/ZdQwaqHju
D0v6hnz+Fui6mDsEKRo0FRJYYo4UvnSAjkZ9YVL6AWpXyOU3guej1sdRJo7lFnptLVydDEFzwCf7
xatK0rejSWPY2JlTXQTojPkCHWcIQIFr6j8+A27pBdj0a8Ek8ioJ2FizMk91qPMZSjPI/ZebgRIK
kZeW/RvlLfPEMD7nl6OZK2o4iCyfzIDUoHgMFv/QxuSs26LQGk/E5nyAw+u7Uvw26ZRKreEdadQr
W5CYaDnvHTrRWBt1tMgzQH+OWu9uCG5cVOVOcjs3eKNPhIMb96JjsK/x3YFqIfCOyIrbD45F6+rC
YAvSVJk9bn5yxqSKKVc/hxMnNU0wpxq/j3Nd+Su8FTddXvJHHm2K2UGI+b1gElX0vlalfaBVIFmu
tjrocKN9911dNZ9uQ0VfDRACr3gysTeJDNNiNZzcK7oVctG684Z7Q7CqRsz12xrUvshPCsvz1a2+
OQ3EBrgHiWHjfN2COMuEUEYT/DxjcAVCdSYfIAJsHR8RxoBfJGWp+XnHzIsBZK1QEBB8ozoF/4kn
GQNUQslKR0do4hJoN/HhfmeZ22zIZy5YfIz8rfdH58t8LdOqXvE0xbGxlBD4+lmvIDddWd+jOSkv
doeM3tJtZJVOVprEbW0/3TI9VpmDf6JG1Lzl0EkSdFCk3LA7w7cH9mXsUxGDb/lZMrCO5ZXagMTY
OrYnPrmyhFyuKIOloF5hfn4XBxXHJEcjL1Z0dWdv/6Qu8uU+59Scq3/p2pk61PA4y00IfoBpLpoi
WKBROx6wNEkYhFR0KHtiIzmsCGmJlLgEqIKuzqjppbBNlnjUTPjj7jBhcYS04WVTxecpunKheMCq
O/eMvcJUvFs/0Y9YdsyoIrKO6Q/P29mfNAlpC/afegQzwyoNhr5T7ekAtT+EqvdUn0+ISjRVQj1p
dnTFaAXWBwv6ZJRQQAWvX00g1dLrdYrdmxSB6OgHzlhaqFnLm/LAY1MxDnZj39PGtKD3NulnMUQQ
IZhet8p6K+LoxrspC4QcHXLjHaiUna/ek5+6e1nlopdcOF9S/+xKeJvGRXwIgMTbpHx3cERgWjwP
cbVCUxpptLE1/z52lsvJqnGnhQPvr4+5F4Up5QVrU9fA++/UrLPPjId012RYGaidcUKQCoYx1IVt
GDZIboERkndbJdNL3uBFu8cB0dZ+TrFXKIpmfk9Trw01IzEqqCBJbOQQez5uGNzfVgyJN6FpPJYl
Rz0lckalA3gygNP37kXzNSKsgN84LKYs8HdwZqbMfioMY6inBOn3rY3VXhlofGbK1GzWNMtveiji
oFxunzeQkLi2jdSnW8Mheb2a9/+zmyt44Ea+c02++DxmgloorPZs+rUZ7L+V8VPjG/xTXK/POJHY
4tPVqFmP84HNlqmslpVqAzZMZO1nwTqWiFH3aQl8NdPsniIlU+DKY1O9mQOqRVETbmOAcAPtRJF+
wNNjmacx6j+c8E3VRayPIqzJ2pTiLKHUg2JfbEJZqDAHYehg3y8vdYiqhu3FoTa7qiz66CpSd5Y5
9ZT8movB4USfOnb51RxXvoKThrqMDi2jt39QVcCWGslP/eDuzLDmbv+7Lz/4iswUH7J4FZjtTP/C
8fMJGSKw4XSHUVQFANBgAqV/D81TiCca+CRqIlPzGx/4mVvRGdCIHyFe7d8pUNB7PdAeS0Ov4GrB
RjaZqDtAqWRxzrCBYeCBhOkjAQW6gm4EKrqXsAIAoDLoquHKpo5AbAcr09aiVFx0BUThAK7Y2065
P2z/sB4z4Q72wlUPu2doas9jI61QSOvumuke7Z8udkYqfM0Xox6z2HnBxnZr0AGocI/cE0ID0zcU
Bgc4B+vaW0Res++L8plZnXAeiCRGZ4f9A/4C7w2TM+BEIyDOlZt4GqrcBLeiNILoDBkuY5Q738tC
3WVGgmfyfaijnRUVoQJgT0hDNbMUCVTR1p0Rkw6L7RTBgs4EnZcqaDoIChk89HjZYIRbhqSJ1YNA
nySjjUYVY0iofrYx44HNXAG+2q2xBpTJRcPmregu63x5N/2jY9+W1zNclNHZeNpaQi1f6qzv4D18
XM7JDJM2YkZuWYAmRv7XKbkILQW6l680rZ2iQP8BcYcVhge7S8Fqd+741/kMdJXgIDnfx3MbvwEo
VunRN2GWZh3Y0VXpb3sU/k+DMfZLKgk0t7/y/ZBWOKNvW9sEdgw5PGnlYwOOhD8uKrzoL5y5Wh38
DnCEFKGgmEL4ZqdhwKsQ50yWFWCj9jWt3Y1dwpuf+f9FE/F7jVku9baY7bVYBUzHQbc38gtVmUU/
e1kItvvli41BsKIS/jrvG0X7xnAalbPTnAguY7XIFwwaWbdqdsprocvBwDUt99FULbv5RAHdgqIS
YF4EcC6qCs77dj6ac7tIWsAF8FtB6jKXIykTDE4NhYa2ZUJk220lm0uk55+G25mUGS1kCz/yiagc
WJjaRPQDSsbxZJQg99OtWJW9C21s/dqUzonBHQ6G6L0/rcz3Uyo4YN9F9FuAiDd5R4vM06YKYjOY
5a3FDAqj3YuN7gWcuhzhn28XlSpNuwxgyItOL8Hel0+hS3W12GgOer1i96JnYg3VjVMK1/ketl5C
lmrFdm+mbCNuoNPSH6PeND2O7lxIQJXeIVC0XZvH6G53vtWD9E7wmRt4khkdKvyA1cG5U9h7mY/Q
xU8Vu0uyqdk3pT8u85jwlJ1K3+bDQUpSigWx4/CpoyI70RMYgpzkZ7E//OzzkH4r0MehbsDgwcG7
W+C1GdnkSA1bDzKnrVFGr6a8MXOAe0tKfHUfohXJoFvAjlwnrDgrlj1iUK1uBJpb3UZjhoMmu2g6
LFYi5FWZYuvyrZjQ69lWNp7um9sm+R/iDE4IRouA+XNqMc7T+KJikHR8H5zxzuG3HWtDzr2LfU9p
0npnxZD+f9ImrOoxnnMXwZ+uOtyqg+nSaGjdxYIeFTbfoCXZGp60TrxljUYKxS8z/6/XuzKQFmpY
Sp9ECXij3X7fGxBNVEvAFMrLgZPZVkGH3NLeX7O8u3iRkkuPY6FEFOUqazps2lzqyfgD/E98YeWo
fcQqcaEGP/A8k53HggLJ5+hEhduqnKY2zNJZwrysDqJrXnIya4Z6Y9AqQfPFjKV4eYsXZMizTt2g
0Lu3Czlom9Ute1mRM4oiHIgUu+sSkywpCYULGwv9f4vk1rjfnT96z2PXLCvluIHcX3y1+nQHkeA6
mF9zFGvlNf4dJKEw6ymL8bt0PqXxBlzoIzacxyajZyyaWawvfwqYdc2bJU1REO5Xf5yGEbZwEkjW
9mhVyZYy6OMDgUJVRAwJq6aEPKZAKj9+fMsudW2AbNrqt2Gw7JSQ+9nEMWwJHPRX7fUMSu/viMLM
5YFon2cJkfVBC6NRpnVcYnq7ZdFf4pYgDz3rxZIZAhAyW6njG6tsr14A57JHUvW31+z5SSixtkqe
XnSWSJsiG/mQ9QtwJkHg3GiJvCtKDrd0YBTOZfPNXPK8y5VpOaZqVh2OQMMRZ4spEkeEBBS5XjT8
XbAu2wFXGYXJJusurfzTFxzFeZFgZH/CPaCPwo+lsxHl6AJsTNDa40wE6Wsp/v2NfdIKxKq7O7gz
pJRKdANAZfVxSGeen5nZ1BVY2u1LxW4SgHyPWfOWmm3wRTRmD39Kbj7HieIZujrMc7CsWlLd6qjG
0SIEAnyMz2TPAN5yAAKMiwNvvomxDRu3UMCYB+kT1hyl1jYWrDpO+kEGK3pKnFdEz9hyq9BPRunY
hGLn0GUQtfiYYIyFO+MzH/l77Yr5CHrz/hPoH9yVEz3cy++WWcBQhBrwvgerZzchTCEKnFluSiQO
HPm6pM//yUMW/3ERQjahhYD/P/Tkqnx9aSCEWm+qKCPsnKT7OY05aA7LKyX54eyyPyTGuZwFMaru
4EbNHeVCfcJXv5kCz2KAcDFz7/2A1hq/F2yE/kWRZdKcXvJmaq4bG4tMLVe7rXL3G1++3auuVCr+
WEuH3pYS7avJX6QCRaI48Z27rJZdhd8kXf8o6nJogTaZPVniQkQtAtAvyFjJCOQnTD8gHQ4ZncEn
/T7yZ00pMII78rbalk9iOE+rflAGuJ5+Txgy5nFoqvtTnXHU0c3edj1D9opIV+XU4Y2FKZ4XHcEj
jRbcVh32p6R8wLMoEZNqtrDHTbJdRyTaHdn+UuSil0Xdir6sxAz2dL/ATkeVp09xu2OL0rZM+wR9
UT7GfoAywZ/28PFOpNz1DVtO/xziSBgadx0UIQ/WseJ+R7iVzgeJZUFEd8KfKtsnNwkqLIDufg9N
P2lY3oQyC3LajifpQh2ZUCKOq639ypSz/nJtEw90Ex9r0sLQWi7UBo3ktjlU4u9KP88t+dLdOtMb
Kpl/1qT1+kZwNwgX8vBFNLhEcQXe5UxT+vGZ6V9mO3yN6udoOFHQhEAYSzxEPMLwx/UlOBFXbKVu
r5U58u0o974Rlp8gwgMspcFOOz6sAOrH7r1/Yh33GQqwDX6dT8xNVztzvicuTUbiNPNt7yVXX7Nt
GC15vdClbEdO4LCgrmHT/D4VISgyEwAYKnQY471qz/ncSi8TOnEeqDePW+dS1H0fJkkWZV98ozyT
z/1w7d2REsD2jVeMG+BoptSbQjyE1RHSF/9RQjBjrm1MJykB63gKiXPB7SykQ+RYJsqgjI3WZplQ
YHtxXL0FnMr3AMwLHCUgGkv6QXEEQCv8W6KWrD8yWp5IA/1IUGUhCjsquUetB61kjsMXMm81sWgG
nu5HXV4yazIGtOpMVKIQFfytxqedHkix/sLFHRKj8/NB7vsw/tksLqd+ztUdQUAChVqlkYvMunes
l4r798R/ZQqstzPH/E7g11UFq20MO5SA3uvXYmi0Ow9LS4toBr6ZfcnpyCTqv1WdYTZsnSuWkZrF
nNRhoOw/XMTMSkCDA4+0SOezWP9y6bkr92+/a1Jk3swudBPb+f7g1qvMTUdn7tUjZxn7ltG0cbYO
ewEG3qjwsG55Y6cRV/MT3/nHfetQd0m1GQxEU3Di56BGqoPVEBMfiTcnr4DBkCW03/mWItDxFziF
1g3kxo/bwq/s+497Kv4AsBu06Wv2pSt/gQoLjRy8PRncMCMBgxpoVvG49prcgVKU7vutBnl4xgio
A4tns5kxvM9KbAZ2DVDEnnc0e5SKhFqXncW79qaTBRsyClorl2Ufem2H+aq1KIw8USFCf9WT0jfn
u7zVgdo9xzX2gsYwnBIVYjxNDGjTPVtHWEG6l2AsCS4y69dieg6G2dw/KWcg0UvUCaV+s0lV07sH
vTooBRoAaxy+IHO+FdGZoTscvCr5oy1yKhp9L2WG5DJPaAj1Fh3Qx8TPRJIsEtsBOCiL/CtMFLv9
hhrFUvVtW0l0oUBs+ECw3y8eQJgaRuNRcAkcdlRnE9C4XGqYvIiNNrnF8X8hRYDulMj10iet2+K9
hjjkQp+CNYXSUqPLprztBlBb6DEmgvmUvvU4Omd+jBYoQhD4TEZbsWp4c7V4ierSjeescVRePb+P
2TtB7vG5ZwJtb2fNh0eVLhnsP2U1l2pakZ/UViQz+ujP8H5hWX5Rth+6pgUqtAdfLlk42YSsH2sP
vweUeDimTSN/UtJvRLMurHQTVt5tm+SMV9QpdNqSrofkzERkdCGap+RDgypCb91ekAeOYo7OpVll
WGgVd1tN+xwEbaq4j9m5KW/D1mbk1pH1btXyYnP5TO+AcG9as2uSDTFg9qCN+D/pvlDhrRU862f8
lHSE6Didi1d8Ge0FqeePl/Gcs5GfVw26HKmypLWJ4YOulBuqa0Vz47RClVDZQOVGe4Coi/JbB04Y
G5sqNzCrAtMf8U0PeJGHap/FQgBW9Zwn9MrhX0z8dKN0Ha9JM8KMTqUhDFxAZj/EmhI1vjZtMH0+
tUs+NDxpxfyYprHYOco3agurs7p5mJQTDZHJIDeqzkuC1yM5grJp4yT9AJwDVnGE+UwVAT0t6+LL
yCxuaOsKJvZe/gxzJb71E62eFmtUWch3qBn2uxBoDYe4elU+yrUggAZzzDSFs1/EYMh6cR2NR1Bq
53a0pcQCc4HzHxRYVdLsx43PuqS6rH9j11ccuImMxSSCWgWLLlN4WvHvyJMyEqQ1q1izpcKYzLF5
p3oXPx2Zupa2zzJa725ss6wlkvhgHjB0lUNzvhZ8uHDbNQ2SMK4ZnIqIynKB6YP1vXa/OwYwydzo
FDsQHV0wcICJWfH2fO74uPPKuEOwSd9f3Y/2mLVOhbxDNWrdgJIdhfM/HKc6bj8tdlGuZwBThgtw
XJ5nc2SgZF8dVRKmmmXNgZloHN9sg40PRb/s67rrIQmUBClsK+w8Zv4zTGwcXaTY3QMGC3HxEf04
cZzWNXhd3dLCgFtipzv1LZhmhkMvGY6UYU3jYQy6wciYblQPK5uZmFaTKrnu9rd7trYtbHZT+vwI
X4ReEBRQsIfI4tMFFrRtgSkkMywy2OYi0GtMXi36ksLL6AxbFjNPprJ58MrQRbDUJg1Nkd4P+s1Y
HHbvlRfOb6Kf0V9R2JXCO/awO35+pS2LrtLLUYcYk1F7vpw55aMjg8mE9ZkQP/6DP57+jVuT6W8e
6sSVYjy9C9hChbFhHDheMeGtPIF02ODBfQgRzB04xI4iqMip63JVLKja71TI/q8firw3561UXimd
r6QZcfQHGfQjjSM8Y7pc+U886ccFrR9895IQau54nxRra0H0+EjasYa4QEQiHK8Okj2m7bwMsisu
cIrALK+H8NmYPOhonCZmbKmj/vFtZLpoQ5OFyFUl6AjqIFcmoh6hPqwJPJqmCWJZQQCESrNMOEgX
WYJOep3Nt0PJFTjr9Jvh0xBI5owxyDkd8DIB0WWPRFi2tu8Bet5Nr5YaZqPXZciXhc6gLKDY0OjK
EOvxHFUkLj3uzcgV+xgaXEUOz4KBTS7dPPt7vw/huUp7RxARxiMlNa2NoYYf93OqpFx+vpkPjZl6
XSoFu3anMVYSsBKFjJvrE0ek/9SIQX+BbL83g4P5QtUDFkEOPG8CmAfbqZwhK/9puKXaSW9wPQ+F
l21p1o0AqYooTzktWA8PjQw8vVcK8/IbB/BESGa+ydjrUm+H+8ZYLdjU6g3Dy4VUEdy97FR0KbpL
tuefjK3y4QF/hMgeT7T4zsKona4g0fJJE09MTjkCWiTNNqrsX/oukDFSDHSaOiacs28d3jg4drfe
E+PYCi8+cdXH+xni9dbeCcusjkuZsJ9jmGCU0dg7tjDzgPxCpHNTYadW462+qZnH/6+zy51xqalE
e6EpCQXXZ+4fHuygnkG3wzKiXQ1bP8vq3cTe8io4+fvFVzgowkHT5twYhJaXYnMgRaYufrzFRVFd
6iVwrG6MBPLBpZkmMQzFAJhyklljaeGb5mLPrV4Cltf3UP68NXtPYziWEUmHVm+wQnRU8N53oyvM
LEGt2bM0/CS7jj/wBJk190gGa7fpoALIINoqAa3P0zfLKiw8gqLa7p49s9wxNoGwha2KR9f2+VOW
r/vJHNhV0KDbVU7HqAg7Ieyg8udqmBG7qxRGIQimUcEYFHVHOsMykgwoymc1inC0eBWiVUu8YAal
v5vjzcGMSk18mzhQEErZY+qksmhmy6eDMKP4ZQSjw+V73x8R3U12uJElsu4ECZ9cLYJXJwKEnoM7
YtF0DedGrHxBrqXC5ReFVDPyPQu+cpRwo0LQdUMvkU6mzzcJkH6tZjpJwrE4U+yymYOVpOrsq9Hi
W115v3+mxD93gOI055pzw762khjP14GBjbO9GyDMZNyUK8lJjv2Rq/OvWdTS0xqn2RO1qpn+/Czm
jhItG6CD7JKNdZfVlvUNZXa/Ur4TzYM6srA1IcSMgpktRVk/NfnLabxi90yY21CQjVi5jaeu+RDo
RSBeEPHBEFs/8oluMJPLvu3Rxq4GgTIU2lxX6fWyf3ERkwXULhUi6sEyEs1YfjkpqhPeMjB8WRhj
4vnig6i2/krPmXiddQRlJ2q213485NO7GTVlmpqh6FMBk6W2IOSYZTUHDfTZwo1ZNDzEOu4Xxoby
69/H6aXhEwhMJ23VUERghJbj7FaJTYSvvRw9loIL3V43evIdsw25YTXsnMLf1hv7RDRceyugoUC0
h61Kj1kC07+Xh96gCjZLIUk9VJWmcPktz6QxMj5Dwi2EzOMG4/n+AZMG4ZoHNOXW3ua0qZQMzQ5C
4HuzpF642UiKKiBahcZBkVeQ2NBCVuy9DLdgcmO2m+EX0JWskGrFWgRIoVtWsLtgjY2TYWOFZWgR
WVD2hFs6LqBW64fWj+HLHHLuZ/pFjDTVfIDDIfcqsKeqe1P4ZYXFeYzksZDWgZx+oPo/4gOQCGrZ
QF0tvJjbzoTdrfSigRxViJd4/p/rxMFVS22L/vHGN174adZmIEKUhgTZoaIrA74rngkAOuzuidfX
Ilr3XagtZuiGie/aTSWYWBgSS/HLrDtfEw2puAIqUAMg7JuhMIKTBTWmcE2ow8xRylmQ3IhVR3T7
+FaCoMo/rfkBWm8zOogjUAo1bG2rQtGhjdHJp1KrnSHi4vk5RqLUw5/fd5eWFP+HOshcbuvNgS2l
cYaHCzVez3bgYy69Q8SGhD441COo9KgeVoOrug1noFgr2y9EdNu1putxk7+3aQRCSciUvlY9Punb
V34mhBvQ24wJVBq4+fWfiDmKdNVXLYR/eCo4dfD4XBjXC/q/ttrTaKNWRct7T8IIiuv53DMG+9oL
exEhVVXFm9zSdaox9rUMP5P/KSffizFAQ7i1LF34we7Ns1h9sRC9FlwyqBB5cuA1P+z8IeE/2UYk
Mn7svg5jJeGf5sDEfHqd9s1lL61j/f0dtlTjEB3dX6/QIHGH9lxW5kIDNu2aF4ln1yevvHNBVjfO
eu0mMOcBIQZjWpjZheRAYA/WgloQ2shE25o4xd1IZXEWFtD+hJOGjfK5xl7XjwET51GfvvCC8ZYY
nqckZuHU5x7x5DkYEaMQclA58GhTF1z0sGzp2WxSkmUFmr1g4khTcWLbfPyHV356jTeYzFtBaicX
G/M09mSGe7JnAmWb6WNdPltyyEGhsBj7sllPAcaTEPLqkSZuxXnZqsp6+IHymkGqKF7oSIZOxZaW
poejdcMgyje0ddE6A9vXgfiahPCLIEzcBm5XFx64C9uVGBWs6TLHz6YOF5EXPy2E6sRTjY2u02Tf
zwthcPtzHSIWsSwHzvvSlJnOwaLWmPRfPdjBYnm63xBiL8JLWFzqg6rs0dJCwKP5sAU78eV8YkHv
l0uI90KZd7IzMxXybE3PdbXx0ypSFgub6aCf9a6Duzv0KshMc/erjDg/4n5PsAit2D0vFODZmSis
CyxlQLz/1MqhESJom487FV2smM2rN5gsqT+TJLVdJWEx0zwn/NS6HO0Qp+lG3KUSFrBPMFCOueTS
4x0kc2mgf22eWFtuaMyzu5z4lk0pgGuyRPQyomI9wo+bLmSpLYOnJfcuiYe+UQixMGQqSARcfMsI
lt3FjQktTp5MGjFkTj5EUwvNMSvkAPJUVBRYe6LAmH9SMK/xKnWt7v6QmL1/WDFeXDbs/vjPlozE
u7dHvJoObDzRml4ZpFXiGapHU/q/exu/CseIoiyOt6If7HyKUZtOg0vAkx9MJkSGR0+meMQucoEf
uRPQRzHoxVKu/oALM6DKL9VMBj1+LQJ244Sv+OOvVHdyPFTYm8bzV2vXu3u0cU8YYK+PofRyK0eh
b9F9Aw5X3rQDVWz6B1+xQHsYZtw75FC2AUanAy24pFrqtE4c/0lZ4jJvL6Emd1pRIoEu2ZbeNty1
sjPXhPnWhgOQVI3bENF4A5xAaH5bTxJ+EqdRVjMIxK0Y6lym3/n/CjGBNRknY83Lto35AaMCSgEO
IU1D3BWmaY/wRC1KqoIYFeONohvgTFvjvLtdK+z/Si9YSWv4XGbk6tNjWdK9VD2cyKTGkpJbWs8j
8J4iGp+Ln3HsFe9kjPwusOhHLWP/WGTQULWSyRACTTaF+JJO7YhCXXTyg4cmH0IL29AI5yXrRwzv
K35TujDof2sNMvJQ2p04JYYWCaAq39w0EOt+SQLjwJXZmXdlCSTKfT2B2kMxHiQfG8uL7enPMk6G
CY8q0cs8HD3d9483XmUpc5x54VxPTfGSMdkMyBABSDOY5aVl6Al/COECAsJfb2IcGBBnJuPIYFm0
T+E4Lt79qS3Xk8QBkDyj8nVFS33P2daFIZLGtxTXKf0VkPgu8MPyCyklMyqYEH/OVaykA5kH5Toz
bCNffVzxsjIpRaP5q+lhdhSS7cqJuyyJER9O6MJ7dK8uat1X2CbRBsb1hHuhZlAR2xdYyn+7C9FZ
PxAPbZEJ25DUxc3YMhttQ7oXuY2vTnpFNj1IburZZtCEGsdbIsQAXJYUit/c8GagizErdOOl4Nvn
9rjy0/Q9rEXodMsziP3DhbJfFQSD7TC8zgm4k8oI3qe39qHFDXScgu+gI3hEGWMzttZvmofsToKC
rBuXmwhzHvEvYOBYCoEpRZpnOodISXr7VJ/sD8rr7P21WaU0NVgyZ8EaV4M6kwNugDmNJS4o2NIy
LrTUilPL0dMZjBdz+XLrQEwZe7IGzT1/CHWQjEppYi1/tn3CDhCOSu3saxlvXkag2TFweSVaZu2d
/uhDz+9LfhL7TPnCNx2VMYgGqBNCXyKumSpBy2nCQnLCosjiBbS0SjUUxKxzLzY5paq55AHrSC6M
SwgcEYunsyo948JWR94+b9mqYKezhcxQDYLi/YHcj4rKwVdSNm15cz1tjDFsEzImMSxW4N0Hy9Mn
dudcSCZl+2tmdyASeJ/yHKA/+ignZpBb+XJocbn1wbor3AOXdTQgB+GZosABSPDTWltkZffPOBd6
joScyaBGe8xRGDTv4y9070SF/z7xB1VbI8w+RRrbhiLaNsIxQ4deqNGCwduUEXtBU6JOJNHXVrf9
E+y/FcNISOxiYAV20XMdINdZbxNfpU2IJwfs2RbnntgDynfBXUXdw4U5+bAOt20MjIxU4DiaXxQR
nYIK/Lk66/RHjQR0oAT+LMePDzoeArKKU/i9MY4T3MImaZmiNTjy3J9SV6bcRcbEzfT6ARIUz3yd
zDy0SUkAaXZGDvYrE1JYBO3tmAr5bousPclhx5Lh1FGG5kI+Mx17pKXaz6KIkOU+jUOvGl9B56eH
e7WL4UTU9a7/YQ+BrDNyE+G3iyOjrORau4EEbLOFQpecrDmHmStAw4qge8OQZn82H2zMfJ9zMbAx
usSGJ/o61O846HK0I35q8Dj1CQ7WAMlFPDfUEud+cd2zRez85rjznJnmBcsRy1bgg/8iOIVC1r4L
81Tf47hFoz252XRVTIMds/1kJCfNAsrZjK62SGxOk+vffj43t0TrWvrZW41bKOm3AhFYYKvHGGHD
xLZOmeSS72IHpy7t02e2lMUvQPK7GwFyoqYTA0lfMzOcgPpGEP+f1qEer0URjCSWoUxepDwSTEjk
I4k065fIhCCrBhLSygnWaxGiZmyDqCQjUd5wc5oBeD3boVMXhRENv+t7IGJl4knwRTI3N5m7CTph
Lx3IKxPzRyaZZvC0KJSfWmhRwHCRJLLIyDjchwN2ja1kpxk8N42bEiVePov2zV4IKWcFmaZSQFXE
16n9BnhaBBIE5qtSZmiKHN5f1DtuxgkAP0PUw821wTmyZFf8duqcPpiGsRfQS9BaFUxNSw12Ed5G
bNjeOESZsg4o9anZH/wtXt/ZXsd2brJZ3Uu3lVlJf5Yzmeohbggg9JIkKcJGT7zgwG1JqMBz/r69
I+S/TWOer5uQ46ljFrJ78CqiCiSv+uKqf6e6a9vOeLnPD8PrfYo89zrwJ14r2CgUoXTmZm/PUVl2
JgxGbA6fqSIWmATuXho63fwjrrkt489XrgwEM5TqYC9vAITtRTjxwXWUvKL16vZio7Z0PgtBhJzo
oourANGPuLruOeeMICyL8JQa4ULP2xY99oY2JGP7ZRpvlHIpcDzkMVt1ttKfbfOl4uExvgQYx3sq
/Lu+vviPlwoitnF6uWmAgk07XFug99R22LyoG4p5MnmFXjg6STzQFSup1bF+OPzpLBp8n5qq4O9i
JuHqsHAXvvM4J3nYQnuXAxyKcHVhCN8DXgf4LzsjZx8B/0HpXEjcjV/HbFwV3NC2E4hppqOgmj1L
iGLSRBqgrO+TKLVpRSNyJB22nZ3gZV1H6JF6PxxxmgP3UbqF3ACATRV2d8T9TlXjHdXBjOFb/Bnf
q64Psvfj4uB56K8ptiMaOPwQjAYNdGcxsyu9Ho4z9M0iKIeksEjG/7mtOoGz1PdXo3iQc/vu8Wv2
qJM/NPTvV/65DaakGqVVivWuGBNHliB3DPZ2ivy8f28obiUQp8efFNURnlFfpZsNYO9+oT16qb/y
tBYzyPG63hi95XatVSU2+Ft16bIibC8VqOLp6BoTH05SamnB5ORDRLXulgBdIP5GRcBIWWXMl1Ar
qSj93J5eYNr/V9Vqnj2Qz2qLkEY9cFh1CGRIxvEj7Xzv8iuwZCbGXFkkF93VW6pze7jUs2KLGmp+
o3hzVgOrkIgJSI9ewWrtep0XfLzzP29nh2dxRd16GCOxK+DlRf8UeL4cBQA1O9v2qsfP11YHyete
a9w/O7VRrFYQQ+h6VGF2TPN9swW1xtOEeKuipK2jBCC1xtbik7bgynrt63Bg98psAcAbvfix/bhk
WFIgfRf8OplPtm9aE2Wz4HupZvhmzVuIMOHnaowCQrvLUuorLQzx8tDrMt1NgP+HM9fpNlCeFDab
FbHIkSCQ3FinlP2kDvH58nMaCLhrqpOAbZiwVHnoUA6vmSHeB5nI0qfn0EqvVq1QtFleUuJyV6Xx
tkKBRJehu+GQLQlrp6k9WqowngTIBruK/OXLtDUgHMYUWhWxND5vd5bgR5r+1hSh6qsc4xe5FnXY
HApyUQd5YcswQVu/IeAQNw3Zqb8o9z0ey+yMXL0r+UCHukpsycyTlDk92aSZg1PmKcsTniCxjFKN
wVhqIeBVvQ1Gsls1qrs6QFovtK9L6Jn3suGscKj9Wuhh5U5aOcUpEC/GH+N+h3Cbdn3/oYM7q7Wi
b34Zre2pAg==
`protect end_protected
