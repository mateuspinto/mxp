��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���]X�FwC^�ݘ��j/�B��h;�7��dǑ�X)�����&��P��l<uR#��lBo`~xh%����U!�qP�<�%Z2bM�]6�1��ԋ����҆�����u�ɑ���'`"�G��S��t��悒���)�d
�P��B�]١���mf�yu��ro�o=ʏ��J�"F����P{�B���đ���q�ľ����=y'q��<���~`�W�P�ͩ��B�;,SY��bd�-��m\�o�	��ە�F4݆7bZw�N�d�j$bjb�� r}�/yx���Z�0�<S2�^�(�P��#��j��3T���ԭ���HD�'O;3T��yEy�u��n摝p�=t���+�:E�ʙ��E���1Q��9������ٴ&?Xꞅȅ�S~�~��=*�Z[����O��h�ˤ����{Xj �������m�K�~�I� �ʜ���r@��<�d�"��Vk��W�@���!�Ya���� ����E������v-K�:fCK;�#�����&�WN/��TzP�7 C��I^z`ɤ���p#/.�Ơ&dӜ�K��ig!r�N^ �$����>�vOh[3�"L�����������s���/���{3���ő�;�幎�f���3����PG���>��0g�v���RE������D�w�w���:��FVZ6�9ou!%lBt��D�u'�x�N)��JV����V�I�m�����dn�V'/�[lYX��s	[�}��Тc�YK~}��]+��G�>���ܾ�az���Z�\�X/=\���c@_��h䡅*����MhTkٕ�C������^�\�@��b����'�ߜ�B9,���~5���U�p��Gb���a��?��qOwVNfQ:��Z*�]�!>�;�C���"9������=K�G�_7o�*v{-��>��"i�ɸ�ٿVX5�^]�֧\ٍ�ݱ��Ƴ��W��gp��A�������˯��e�t�c^������W��"U�2���a�N+A5Z#����>�u4l&�s��	�a������G���U/?L�lj�g(|�f���p�#�W��U�����f�"!R��؛������*~�|A�L�:�]P��e�E�mL�N����`����}o��5׎�W���'���g�T����U<A��.U�[c_�����>�ݿ������YyO�M]2�0�Sg�{� ֢�a�A�}	�
�j���l`b��l�Qux��Ӱn���Q���r��la�5����-U�\��ζ���^��g�W�`�}J�%G?@��, �(���,�:}�B~�?訬��`0���Ƀ�t����zy6��E�`1z`�拦|�t��c�X�}��Nr�}tT��?k\�G�%b�%z�.M�{���`7]u<Y�hw ��FN��RN�L!����$5l���-�c�i�k��	L|��F�	�,���䁯� ��
\����y�G[Y���2�j iq���A��~>x�,"U�R���3LG��x��-�Cq]���m�Z�xu�n��������FI����<�궹�R�_�lk(�K󴹡ET�E媚N4zS?6=#3�������}�f���I�.68b�-ک�w�ݧ7|��qSNG�mF����}e`./�j�E�ŉlȠ�h-��m�,M�mڐIa"������I�zS����E�x�_Y���)=5�����m̅Ur�m��7�Z�)�N$�h�#�bL�_�I\
}�I���;��K/с�����E݊�'���mÓ?���+�XN�u�6\+a��_^�$X&�p��W�%RU��f!D�f��#I��哣��$wχC��J�~\�F��!�r��D�,h��gt�=ך��0�U��'�1���KC�Z��V�l&M�z(����1鮂�(�����<Η�R¦��9�5����"qq��^:F�I����K�\\فk��C_���uH:�0_u'L��(���޿�7i#���|-hY@!�����_.r�X:�[#�� ݷp�#��ĵ1�e�Wo�?҃�$�����L^��ߌh��A|�=My�����\[�(��\@3��g����.+W�Qf��Q��鹔k)#��=�o�#�v�)̗��2?L�.����MĔb{�����>�s+�®C�jj�y ��m=�}����c[]轻6��\(T�)Q��+���넨?���+ m�l����Q�Z2�i��Ƞ7*w�`�-�1���s�|V5�U7���.E7�B%fK�|��S�R8di��z�z���d_���L�O�B��W����@�<���}�c�_��F0�����d���~�!<��l��8�C��v�����ue��[�I�ʜ��S�X��^ ����b|�{ �2j�j84�#�"�L-���\�ܠH�a
�����T~.$X,�s�,;��6�缦9�VJF����To�.�Rf�W3��bG3�����J���mg}��t����s��7v1�����A[��)�o~�����rA������4�>Q
v@)4���:��e!Dt��gAFIv 0�:��=��?:��c�c��\9��֔i7#���m]I��f�֖'X$� ��cn�|U(��2����2��-{3�����`r|Tl����>��a�"��z�_ѿ�q����*��JD#lR�����������z+���>�~S3|ͱ�{7?Y�$�Å�����q,%�KQ�m�?v��;Q��eo������]��)������Q�)�I���3�R�L6��w��{���׍����J�i�lv�f�F6:3�d�l��k�x*h4�ߒ���-���d7�3w��5̒VI�y�����H��g��ڠ4�TV���^j�V������F&�_�rL��_�'/l�&X0�}�ڇ8k�u*(�b^�ø�#�:��n�x����ʂ�+_������ö'D�i�!d,ژ{.�<��'����(t]J)�:����tx�`ѯ����x��<�F���F��7�[ZD��MYk�׏��������9��Ȟ:�C3$���B�t���>�v���c�/I�[�D��f�V�4e��¦wJ��1�.����aV��'�)���0ꘑ�c�B���j+׸�K�bJ+v���8`�k �k�aNX��w�3?ې)�F�Jo�.�(@,�3�I��+%���m���!�'#�cD���������A+a�{ r���벲k�k]gw0A���{ۺ��m0��%�$�d���(��9� �M��$���V%�å�� �yKil�o�aܲ)T 7f�c��tA?�.��8:�ߤ��
j�-����E	��������ˬg���6gV��N$1D�)<l��K���9=*`��b7����vl��T�<�� �,��5 u>���Є���a M��c�s���@%���$V� &��W� ��f�����3m�$��e�2�ˡtK��e��qA1&g�	\��1͗f~��I������'Aה q�1MއuA-�<��������:�sH�a�@;�:�9���JI ��/ֻ~����ǂ^��Ì��r�3��q/�X}�:��=�*��'c�-�M���d�92Nã�r�a������6t]	�)+}�)�6�nH�' /�4�B���Z^��Q=u�E���l���l��jUs��s^Gj�'.s��:'C(�"d���~��'�O�U����"kw����Im��'[
�3�1�k���ƛ�X�,O=����^Nh�_�֗>Q������RR�G�(��� (��$�e�4"sc^o�~���un���/�@\9��3���)Œ`n$���B�Z[9r��=A��9�ú�F���ˬ�B�W����ot�������k�Y��$�G��	��Լ��L⮵wp��GHIV{"3�[�V�a��m�{��闦TF>k1�ֲ�#����w=Rp�G.��=�Ky�GK�.��~]Tl�j��v��Q�3�*��؎�fsD�i���_�{M�-*��a�<� ��+�gyj��
Tq��Y����:���"��X����H������`�
%O�]:-2�<@����k<�D��K�B!8 &����Rh�/H���
6��i|�|��7�j\�L�ch���.'��Ipu��9�Y3�>:M�%���݆��W�sp~���qB�7��-̣�/��n0�u?�t�,�����B��k�&�J���&$Mhi����G{�trN�]�`*�,����W��qH�[��Df2B���gi��1��K��x�ク��|�8����g�)��Zc�a��ӯ{�4��pƽL��i����y�����*,��	�1|�850��h����H$��:��Pf��ߏe��(L�kdw����ݭ����ؘ�	NP��-���n�)���}{*����>�(��-�����J�j���@��bӠ��4�%���� ���y�9?���]g̣���:6"pa�.C}h�d��\s��c�I��HpA��6��Z��DΓ����(��ը�	UήJ�{K>��l9V��>��w'�oN	>i����:����_��:�z %AQ��7��Q��W)���up�G4}���p��g�����RK6��v��b�h�k�#L�>�h���,���AD���|�w�S���ò̻��{�"��R_2��Vǝ�س�a.���T�ʟѫK,椮0C�4�%o ��Si�$��@4�D�Y��=������O(����.ԏ�P�����I0p�l5xS����������N v���z��s��8�<6�w)��I#��6��*�)��`���^(�-��ou�vz�_��Uj=gr���:"k�4��z�����R�ܚ5@D����<�g�xqj��g��:-'MI:���B���\&����}A-��C%�\�b[�b�eة}�̮����c���?�'�,x�����t���a��<�)+�����G��T�;՞��OybϦ� $ {[�PB�	\u(߆(I}��oZ\}��Ţn ��P(z�������G}�|$yTD7��sO��0X����R9հL
P���_�!�p,?O$���&�'z�/�[V����,���x=���{�9	^�K���j�Ֆ\���}1�2��O�Ζ�>&#R�C���Gn7��1ht^����1�GVU´'Ty��H�^ Ĭ�Ҟ�L �gm�M��m�!idR��aT��m��'�w� ��cM������S�����C:��{�π��+�]nf�<��|��?B:�v��$I�RÕ
o�۳���n�3\��%�<��{Q*|����3\���c��(�h��\�;?��(��ٟD!(ɍׁmp�@���,u�9n�5�[�X9�j��U�,}���q	ܐ�w�R�]���V�
dO���zӞ8j,��>�� x�ӂ����+㭂��G�b2u��4��*�d��Q&�.��$(?� ���rM��y&-�)�D���L�I,�Pr��<{Bx�]���sW};�J1�if��L2B�D���b��M��U^�G���ݤqf�,��Q�®ݚ�Y�ؓae]��Q��K��t�)z8m���<�3��gZ($^cF>�y�U��%D��R�q9;�yN_	ӊP��w�B��[I�Xo%���`9;3����h���&9Zs�p��w=�t�?���R׈�f_��æ�<Ղ�X�ɬ0 \!>m�%^���HF�b7�ti�@��{��n��ɶ#�T%�<0�+�u�`Q#%��,���֗���ή߀�8pY�lICG�$oH��C��aT'څ�ys��\0�C�㥛��tL
7�z����n�mu�(�<��a<!%���m�r!���,�5"L%-�,`0�=�����`J�w�jji��#nP���`���k��֯JVGɋ���6�������}F~(� >�0%"4,�����?�d�/�/�F�� ��6��������Ǭs�(�Sw�+ܓ��yi%��y�J4�l�|!�p{��s��l�"�>��5�PN��ϑ��cT#6竽�/sv��?+ �v^s�����ۃ&ݙ�5�w5�B<tꩡ�Ù�r	��9��+Ǥ=��}s�JK)QY�.`G�@��ǿ(�,Ҿ�\y�<$�X�vW�� ��Y��b�tC�b&�e��%����	�Y��8/pD�������c�ƒ �~�>�ф;�сÀK��/�v&�wO-�%�	J�@�/ƿ��..V��{�������%�	]�co����l8�c�������k�h��߄T�o��%>��٭)�����k����S�XȲ[\� 3���̯�aJY���J	p���/�e,�e@m�����$Y���������10�+E��7�Z+��? ?e�=��:>JvD+���`|0[T��"+u�t8-��?�kx�YW#�,R�F`�ԫ<p�Zz�iZN�BŊ����\&CLA��ۂ8���ֵ;��2К��V�H�S�_�C�իng�,2�qP���AT��M�T93�`6�G��d���ov�D���Њ��W]1��9Z�u��RH3��9�rz(~��@3*�8�
S�"x�B����aJ��8���I+�ȴ�i�hr2�.���P�H�߸i�B`3R�w�n����Aɷ�詃�����*>ؼ0�|W�&�3s��SX��r�mi�=�����|ƺ:�{�-���� �X^�r�_[�} Z������� ����:�y;`J]��?�r���Urc�����&	������W�·v{�v�1��<������!z1i3��V4 i��azޭ,`uA��!�0%�ڿ,Љ��HP�)xdY�R���)!��"�D���ww$���|.8���N�+=X̘8*�KF���_�ƨ4u-�rő��!�w��x	��A�9��w� ��I\�J����Ȥ�1��������a��QnL��9�#\m�9HM˕�hԾ�,%���M6����5,�=���r�-�σ�H1�'�G��egތ���Ѐk�{���r��L���T�`��j�7Nl��~�"��ü��E� �kꩬ>Kda}E��"U��S���m1����m&���S��0N�|OKa=�d���32̒�n�	���[�x��cH�m|�߮I���	PC��߷�G��%P�E�����ZE�e:s,kh�@:�Ţ�Ǫ(��pޖo�B��c����C�{o�@�c��l��o�K���X*ğ3��`� �6?��Xns��A�k�<�J.A �~` �;m�yu>;8���;aD_�J�!}$��hn���I��i�	�<�/�n!�0E�ah�����//����Q=y7�3��fT1�m�5�<�Y�6d��L(��[y�gޕ��O�SE��㛑���Z@G��cS��"A�t(�f��\�����_��R�IT�=βĔ�nX��f�.w��O� M����d>}9U�Cp��6����_�
�h{rP8:fs�_ 0sr�3��R�(T/�nç�9�[3kmh�	;��{�f�K��.k�>���D�,�Mر�BNL�4�Tۺ�R;������M���ޚz��Z�Cx�=BI��Ӎ�kS�;P�/���I��F��*��W.ֶt�-0�ɶ3�E[W��Ě�a��yL�4����9�iq�|����!=�*n�y�J�A�#�3�Yn�|l/��Hض8�wm��ȂY����R갏D���u-T����Q�E����N�f�z��R,��QL�)%�3'z7e��|�pA\m�`��o_gt����Nؗ<��d��#���/Da�1� ��n����1�!f�r���C�+?v�Ś�0jW�r�^���i����iv�}Ո�T���9�\oqc[UL&�t0_P��+A�>1�2<���K��T_�Vt�i
N=���>t_ψ�&��-�͚n����V�QP����e|�u�������./�a��\\g��|�+��8�l���U���H�t�8r�<����۴I��4����۟%�?�#��:e������d�+H:^7ߠ��	�3��r	��ZQc�v+/���FC>� ����2������� ���8�
Ԣ����豅��:n纐.�����dJB�Ȭ��-e��ILf��vP�r���Z���x�շ¶���g}��&Q:_�SQ��R-#���R�ſ`���$�b)��_�%AhR0�m�hsR��h�CW`qQm���䀒~�oq����_f�vݴ�6jˌ�TK�~�ݵv�&�^�*�����q��&��OܵV��{��b��g�fV�Ci���R�����$��
a�#��n���?;r���耜Y��t|: xg-7�MiJ]�S�R&<���,�pU�Zn	%�6I�t�' �����,%[{-L{=?M4�X�Qu�A��t�\������$7 �Rc�-*XXVS4:�s.���-��E��[��Z���#
�\ʹ�����~1B����#�њ���ql-�+��}[����Fs�ZZ������A��[��J��A`'�q#�}U�W��ć�U��h��m�^�bՄ"9��Гvۻό"jӧm)�ᑧ�����ޟ�bwQ��_���k`���m���,t�lGf�	�,�^��
/��QHJ!cgP��C�Ǆ��]�-������6�^��-.��T̋9U�,�T�uBe��^T��u?]�zv�N�p��N2��'M����������_ۓ�y��|������\w1��d"��d����&���=�_z|��z�$�<o3�[��6�(@
���@
6YKd5��^Vd�������l.$����QRt@�(��;����3���Qw/��Z�6*��c�5ǻKf��rO�����C(C�:8�mʺԛn ��pv�{����@��:���S��Lk���ǊgJ��'��IFý���#�m����g����_\&�+`G��5�d��xZ~?��2�ҵ*�q�k�M-���W�\�a�n�Q�H-��;�)V*���l,�vtl7�Yg�+�9�^c�jDi���b?�I�$�W��O>������:J9��V^暩���n��A�=�7c`����Z̴�o	�*��a�/������w�˴�d,�F&&�V�K�M���֔x�D]q�
��@�?v��l#�ý%N�ʡ�����}�&A��e�Z-{ám9.��-~���-�
&���	Q�0��u���pUKq���7�G�ߟ��1����s	�i���-�+%�0�GDjtqi3����Eaej%����K�����%�[v�?0���wK��� @%t����ć���I13r3��ܳ
�q8?�p��q�摠/V���[�@ަMG��9���"!J*�&ѱ��ĀX�o�h*���-����.=�}n|�Yx�K��r���P� ��8�rW�
4�C���.��5�������r�v6�������<-kn�BgS�ߔ��D�lKЧ��]ML�1pT�_�AKL��������uZeI���^@N+E���?���[��v����J�>�s�?�E8����"{
6��~V3��C[f��&�z-H�<"���~�D�pn�f�i���%�Gk���,>���Rn��M������J�Oyǻ�R`��ݝzr�E������E*�D=�Zs��ѡ�����`ݵ�h�T:�eĎT�>���6k"2��]�����g���çIL�&�!?��7k`Kt�Wx��<�q
Qz&T���g��&v�\�e�g�"T�=���?�4�?ɏִ��~�s��������m,,=��尣��Ym�~QX�č\l>H�1X�Yy �>�謐j1�������AB��?�;��b��u��&lv&�D���d�'>l��.�H��KI�������_B�Z�h�o>�#�9��W�f��w�h�9ݷ��K�J�m�vmӼ�6�lI+5�����������bG���mE�J�א� �wqYG��X��e���3�����/ލ�_��˽�ǒqA��R�P
�Q���N�F	(�U¼;8H�,vK�{�����am�h�eb�Cdpԗ"-�c$�)Cv�� ��\t�6G,&Y"�[��w�o�tul�jz��Imy�03簵�����Z�8J�u�y�5���tV(*T?q�x���fi��0�T�b�h��L��^�]�-O5a6u)	�?�R��I�%��˜G��-L�HL8����*�V(nAM��P}xh�PJ6!�
��v��N��-,������.�2�wzD�����ş�g�RV60����^!�ݏ��	��njI@�?؜/�+~S������y��|1O)>O/�u|b����fT�#�0@��?��U��@������r���3�D�縊�S��u�G�>���G5�FAN���O��n*Fښ������8�E��cd�v$�KTD��"=��q��K��h����}Wm7B
������"��Y�RX�P֤ǔb�%9���wy֊�6�܉TйQ2r�����=�yb�\6=�=^Rr�}�s���u�cއ�G$�}�?�M}N�ny�����i+3�V��i;��nOE��#��)'K�����6bU��t;Tl�l0x<d������$.H1WN1����I9�A;E�F5O��$��p)�U�i�opJ2��&8�q%ڀ��U0"����qO�Z[Ǻ����g3f�,�xA�܏K�QUi��'����юr>p��%=�1Zk ܘ�jQN)�;��kI�$�P�p�Ni���l��2hX�I*�l�/�$��0h&
�tW�l�M���=�����%�\l����c?A,��g��!� .�GS�VzG`���_Z�v���T��,����@2�߶c+�i��d�=����(ȁ`J�'�����,U���!	��m~@�}i��$>`��ST}+*�o��V�2 ߻��>�����zТ:.\)uK�5�F�u�MѢ�	���y�T��Vw9g�P�4��S�,�g�d����|���W�Lr�N	��9)������pl�Cyi�5p!�y���mT�V~.�9����xM��x�㋏�G����*ax0����Wo��M���q�P��u���O����@h	���K�dcκ���� +(��h�_����=d`+n��S��RȖI���>�"�٘��� ,��9d�+��M���b�>Q]پ-��_��^���x�W�J��	�*oI�詙3{��8Q�w��ȹ�d��	��|��xʃp��ͽ�������ݿ���qY�7��6V��!�Ў�N��j{=.������nр�h�e%~o�����+  �B�Hha*��(�x������� �i�Z(zT��*'�o[W
G2tRw�p���k�� 1*���YnK;O���!�%Zq�Hڛ`��$����?��|��}��`�2Hu[�]�y@X�Oԑ4�ۻ�*��
M��C��gl;e�i���\����R����$q˟��:����n���]ߏ��������J����5U��
BW��`Haж<���?�w`����<[�_�G���� �H$�`y_֖Wv2v�pC�v�!Ѱ�����uD�=m�\���(�!u2�1瑑��'*�r����(A��������0o1!��K������8H��ð��E�.��F멭��X	�J�}��N�1���ڎ��Y �^���u�0�߫�ں��~eL@� K;�����`M�H8���������wϨ���Ǣ��m�ͳz�v���1�5�i&���eiI��( >-�������5#	C�3["�瑛ڮ/DH2cN�Ǡ��,�>e37jA8��*̵�?��Xs�wSpH�ZӹH���W[���u�zw}4�VՆ_�sj�k/�0���#�D��!��QT������=J�4��%��ze�,� ^	�I�����ډ����'<e=�zj�8�Wi�0>d ���;� }W��&��g�(�4�v�5��
�_2��LmAj�k�oW�δ.�-NHӵUD���v�"�Q��M����79{?F��2�������P�`�8�L�m��~]�8�t^�#���aC�m�T|aʧ��Y3���U�[
��/fS���e��17�㑏���oӇG�em��Ǣ�۠ۼM�H�8�0�Fv�hw�9��l��DN�.�2þ��	�9� U��s�{�>�����=}�p|�D���ZW�N<��2.�r���uy�)��E8�f6��?���o�&���NL�~�Lo3��:^�0�%�)<�L߁�wG_�9)��4�iwA^�ay�����V�f>��Ԣ�r)���I���>Rs,Z��¹��H�ʎ�����'�bl���y�߇&a���-�O�%�d�����c�6�/e�`6]~�pm���x�pV�P�u�Z/xj����%sh������%8���i������wb[��A��6K�:��y�ʁ���ᾡ�r+Փ�oO)|א���I��i<}�	6��u�M�����p��x�"6V�(C67+ֆ��r��Z�@[�Rw��GF��H��a�4���~�|�
�H�>rQk�֖D�w��]�q�j����y���|}lJI5Z��<F�Jכ���-���_�м1<H%͹l
�n�u�C�yh�x�_~IT�&�-䃠or�x�
6bhTR����{G��E{Za�yQ�r�}��Jn��GQU*�t���v���\�&סU���@=#š�sZ6n�^G��=#��J��������+�!��y(�����Ն�A�R�4YD{cOC��Gv�O$�ܮ���+��'ͺaz(X�Щ�>����Fm�7�����R���82��❘�.�f��N�oo/�>�d���o]�C��w�3���G�ͷ�A�}�սA�Ķ2�G���@/G��S@pe�=1�W��5�Y��q1ݤ����[�U�_�Ј�ih#?}-ِd����Gk����U��>�'������M ̱���t�u����n���76Џ¤<�*����?(%YI���N���1brB�y� �h�(��}����}�"E�M����<��ЬO kP���GEҏ7s�� �]���nvz<�&_E�`�;��%r����O���������#�.�(T2_
���"�:��#�����SLي�3�zcv�q�n�rp��x��g��ku�b"�k������o�4�h�D��%ce�@��j��} 8��?,�r m!��"��Q8;���	D�b��]����EK� ��1����kR�A�.`SXhw6��"��sWL������pL����-{��q�K!��}�׬�H��`">-����^��o����ZH7���@�g�u'���zÌ��6�GE�Isg��W���ֵ�z�x=�@���Z���+w3�z
xѹ��0b�� q �΢)N�=�Ҿ���1K�j�:A4'�Ê����8�:$��Zw]�>�OO�O�dWq��^�.C�Gu�ґ	��5SXC�Ҷ^b�.Ao�/� _�إ< ��l��4Fg�)x׃�^5��� ��wXJd��֑bq���38�����63�D\ �lU��	b��\_�S��V���7���;�!"Ene�����A2��Qt2�&a���[<2r����m�{����~!�^�Zb�M���V�e�;wI��
#���2Hb`�Qv����/hLXy�GW�LK���ě��x��;a�:��q�Wnz�5 ��|�ǹQ�?ޣ�pڙ�dAA��=��?R#��o' �޿���Dҝ�����F���r����M�����������VS@�31��������r�n�9uH"� k4m_�5�v�<�T@�\SdƼ��/���5��h�{��2S	3w�v|$3�Ou��&�ujm8�����5�����K�2�汍�Q�!��A-fwT>�2�^�ּ+�?����}(q��k�Mk��yW��M��a��RE��Y��[���V;�T����v���o���
������J���~}��mnH)KQ$�;�F�.��aɐ@G/�3I;,�͡R|jy�����n���N4 �UA�Y<c����! /f�q裁^�;�R�qz�I_Z-&d&���kI��jb (v�;��{[�i�]�w��r��`-�KGN�6�xzs�\���UR�$������%G�@�}��W�0`�Dꃲ��e��{�m�(yw��/�i4��ٶY�.���?�f�)`}0�Y<�]���D	��6v��JZw�J�-}��ǋU�j�s�k�h��p��d3kT�l�M�վ�J�U�(��3�2q��i�T�zx~�΁	!H�5���\VD\!ܿ�� �y���ĳ��µk��&;S�%e���