`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
bR/vpw5zCwi4hftw5LDSegAoBbs0zGxExrjYhpBbFVmI6A2My1X3AiehwQ9ww/eYIYIlQOvw2Jph
5nJlKPbxszoqX9ZmznKQ0T4DFxQ+tI+IfwkDkmbPKc8TJiPJXK9n5fPKydIjq4HpEO3f9DYNBlwz
SVq8vKDusNxcsGhpEblbK+vbTF/zj3MQGUvkDQoAu8p5n6K5XLo2OXstHfWZUt1Be8NU5AqoC8Oc
PDPiyxPYDFVFjwjwrjLZvG2nw/Ch6AAnhvq4wwTUV5NG/ByaEVhnjHKyH0pQd0pgbrvXupTGIoeA
tg7AtWJWWu1BJqPGf/giN1eQQ4C8qHDYjmsggQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="0dVlJy3Z76Qh5Agw2shhmaV+lgMjkgAabzb7N3eTyo0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18000)
`protect data_block
AA1hAZgkEB0Yk7yv88kk8c7mtIMrKRmselVvlEjjfiI+PnpdCLfpyWAMuYj9DJmRsIrMi6qMRdWR
7hWVKKx1GZQGRAOIUFvbJEOtzOSyTZra9nyJRPof3yZhMwj19f7UAxzMLHod128Q1RCh9MmGkw4d
O4vjJnYm8rsUnPL55eCsmcr4ZBAl5VRBjaC0hKHLtomeie4KdfojDj13ssr/PXT0B8oJfy/d4PD3
jZsIqa60gyks0QCGfXZ4T74R2y55WedHHNxiAf0HXGlAtKI90bhB6PkkMk7Oovjnsu4jtj3uOH46
uHE7Vfc6eL1LjkD29PsBP+/oLsRx4gFLodK/nirdZUoQHOER2cMtGsk6Xc7SsGaaRATjvrLCP0s2
u8I9K0OAKoNUk3jJzfKmnUQpxkaT1+b7gJAIkurpHytHd7H5icd0z1gDZZFGlN6G4Es7oDS1AdqW
gnC7wZJ58a7NMjn40eOZYgjkUwN44903Jjqr0ln7CvLWsPxxQcrP79sVd0EP9OtJFy1PimvOWv5t
N3BO/jbi9a8n6pKg+TESJJ7hbWWWsBsurmQBwY7GmJ643+b8Rpn/VygzMRpyeREKd5PhyqXNHXf0
x3jSlHlbc8w0kvZVYJ9DKD3WCvaEgOEdJbuNopB8ofVGqBc5TxQp4yT2InSc8no5wsKm/HC6m3ey
w+F83suN5uz+h0hjl6S0ygIu7lNtKKgHroMQO/YBdqhkQEeAgh0WOEiMeCq2dc4w+Ln5zxBnWEBd
kiBlQx8v+YrLjflyDpwVAsrVMefRKerg+foeXoJwsXTYEAb15nwGnD97eUdb9kFnxc5ZCecCUA5k
DmHhzet+Hl1+a3ou3UAOMZo4G6ICse/QzG1cs2aT2nQuboMtzkAkbnRKtJmDA7joXb1Es1btzaDq
V8QjlAfOfT+oPCb7ASNn4VTR7iso32yIwnbY3WTFXtTTF96B++5WJ65bFPHlFzL56fBrqpnHCQEO
ujf6Wu+wxZOB9S+Hgk2J03J2wrpq/BeLbMYFrgvpdVoXwSi4XbFIKyroG9lqE2OOiE+oUQNmBcXD
n9hWjkaiWB5cRthVGUNJECnv5xYF4jEnsLBV+Gaf2sBFEkheZ/PLE4Htvym221xPJO1vi33XiRt5
yTBESlxcjghJKaiX3diPdcdi6wr9mStWwKWbhHFkoBIW0fytZYSrtvfKtuO6E2dp2V9h141oQ1TR
HUhGWS3eObQVMRUxegOHbbBj4tiOSxab2DpOFKsvmbY+BnA85563rkxlQ9qqcMZeR7JeciFSN759
gOorapN6f8+5X+WlHtdRrBsLM5hP+PW8D7iZHewpQMSoGv6V+AyUi1d0saAyPYg4bDOJM06NxnwY
eEHLiZ6blK2HLcwjNdLP8CVyRllA0V2EC3Nq6evGoqf+k2uetXWwNjw70Tl5k4WNRyea+hYSzGhp
n03z33novMTRFyIXqev7LQ7zVqfUUt60MWdRLKxzBGznltS7mF0RA79jhCSJx/jWO5KnjWEk5/m+
0Yz9v8Az0rA/b5UMB5c+WRGg3PaRV8T2V6dv++Nwj7TWDLMvC3u7qJ1KiH5zucekw578Ar/pfwYH
t85OZR8gGDzesHoyqIWJxSGcBNRrU4I/Q5Scpps2jOSidL9Bc8dPBb0NaM1NDnehNH34TBONcnMs
eZ4hlilUTuID72JicbHVMXI5r5qIk/Cz7Lndrusyn2ce09CnKsOHtD0p0DrKhnmgX5yVrjTkzIKw
dVtpaospnxzG+LRaH5yGEg1AV0x2KnnyPWVEmXGcOu+BKVKzqSz5YDubjgUszp/fHd7AWn3BZc0g
/LE8gsNjxf8QlpPXvF4PPURrZgnekkCGulXSsAyDW9b2kJtpx/N8RKsQoYCH5PhjqLqSCxh/yABT
cXuCgSthJGqHNNgPAH4LTFYumB6AAYEbeAZYpfWAbMFxe382S9wwBV0Ng3CUBjiLothSH+GvMgMZ
LsmCRESmlVbg6KsJyyaqUoDlSsuz5HI4WsuU4cttnRjMW8k4A5YpIwm3J8h1boRzbmg5zw06Hn9o
Sd2qbMp4KP1qMMeE3OHB9R2tp1F0zPrAY4NeIPBAVtIEm3EJTov7t9b2h7/jGwLvrjC9oQ2J/j/g
KgLJLunDScSy3l7ojjhJvCliGfInAVZHUU0Rp208dP3gTxaU3LAJm2nBKa2UVc7DzVydvF8GIeN9
siNSb5Yw3HuINj/NeqVVAjl7v8RruWFN5vWo5w1T64EwDWfTi++dy9ye+JD5N47fMXgRiZYYooo3
5Kj3f+eudZA1Hr6qtTOU2FuLPqtRjlR/yLcJw2Fqi4vJTOfFBAmFZocMQWWBk3LfT2MQcT6gPVa7
tCcql8TnhKKCNDtr/0BW1kdLrEqD/cauIA3KXuOB5g17581gnggTg8WIreYT1F37/+dDIWhVDFIm
gwLxTGVyULX2GOrdmOh59aQiVRPX0UG/vQHg5YiEsVWpcqhnbLUpJc9WusWDooARQxrhNFcwzAjQ
TRMUSNN9fPAQz3iljnWa8thfe9ZdmObE0tMQ4hUJvl2LdH5XakHTK22dtKtX+on+erycFHwQupfZ
bWVUPSH0gNCPbl67T5UlLT6kvhJkqgTWHqNQixwHZiaWWNUleX/nv1iLG0V/Tm0p2xC4mIuKpL9U
oup4bRPkomx/PCG9/G9wzY5MWWB9zBoHYz+rhdOcYIhVVEKwgkk1DXmU1vHk3vQY2BVBDYMPe+MD
eyLQ2jgf17IHpTkMa2bZIi1IBlAwTmBG5NcLQxyi0WkCHkppYZNtezgfvbo/q8OguN9StmpdOzLF
rRSlBLw1codOTLBEP6OHe/w3UUZtzDwm5jK2xLaUdPyBUWDGw5g1D0dR3f3DDPuaSbOYxHhz1R4Q
FJOMoiFFL8rNdmd6MzmMnQn1VHaDHrkXCTPT9k5Ow9CCRMW1yruaXa2NiqDp60AX7V1e0jOMe2ty
Q34/eMB0XWL1Iu8ezdIn8nlF27pQioxrZ+MzHxt3sLff90+NGWZ1AUFwxXSE1Mj0+Ox501lwAAFd
/dYZ8iQY4HDrr44tcsLOPzKynA4uuOIc+5bF2hGlnVdzl6wm8fB2y1e97O6kz7GK43cEmGDR+MzM
Vl9gwMNTUuRmWCMbsOvxGY0u8u3pkokKM3ERVtutYUJscZMqbt4enZcJQbGKt9ggJHf4diIOi0Nq
ycGJiI/YmE9+mnIOXOsC740GtPsTknEsmpMfqO+uTg5rnhv51FpmLz+KTV9F3E7tNuAwWlepZ5lC
EBO/0jzWgX6fziGsD9Ddevbj40zr7tXIUbo/pOv7eAJvySk0TD3MS6WcDvzoXMdjyEMmSm1oy7Y9
wH45+9nf5XTvFkaDGX55xo7gknvg1TSbbuv60iU1OkVQys1kOeYf1ghptfSgN8hniF2ohC+2SI+m
Lsddlvqevipfj+aRq0yRjGEt2i4xnPleZC9Hh7Wp0UJrLHAo3+gEitZmc9YNPWRP5F8+XhVMiOk7
MMql3uFKe2Yymxh3+MtNmhcf5qGkJm1etJiALhEhZCn/PyH8oqHbsVnTu/pIJx5dYdVkjxrEfwwG
KXza+bW8o+6lAbR9PEN6PU+o+PO0tzvwIItdwT5pOb/LahG4bSmPW57FJ/ugla6UX5sq0Git7yql
4yGqmGBHAhJTZQnMNftjlM0YMwzLPpPAOHUovcvEHvM0I1TNURb8tj2D0eCbIqWBV09nYh73VTW0
gVwbqkRLDxUsjx9JySVLAJMP0bMUCyhFGLAW9LrNa8O/0YowSQ5dYqh4MW67dTAEu653uUyG7aoj
op6eJAxmA20WY1cTFFJ/bvGRmZsWV6TPiYd8UF1qZ0BmcF4qAkNvf70UrUjDwPRPeybQRFKGd/rk
LOnkdVN6aI/oqbjRNgBzrjL3Rq8aqTlTg/TjoPr0+pblAGvDeHSlWSt7uJIl7hmyfVcqGkXqPktc
5TgNSn6JDNDOQJEVm5DNcH4r0MOR4xiwmvzzMuBHDMS5vGaOxcpUvGZM5lmaaCtPXtQu+1izz1We
fGMuOFru8dgNn2NBnHFX/dyk/bTmlLtsn9zSRhNRU32Q+MgfXIDtH/Ez8RxWDKAdEzC03jgP3yS7
6En0YsYhgas+oDc4dkvS5+yWIgP8oddKyBawqXu/tmmEMuBI2998BqO7Fc8uMtzpYU8hTM1OGGXu
sIQO13nGSzwlgyIsWVoFR+W3VyDyBiW9p9lQmPc1YEAhBl307sOR5TiixBXGyIUcvv6tzIQS4K3C
XPxc1DVg+HgSh/NDBYoHLQKzRAwgPELor7Hw+l/kRfe03LE9UJDwGn5bUi8O0gcm2BKqP+wICzP0
8RArSNsx/nJpknWvtpVlgbWlYnNVJU9i3BNHhQ/2NmpJJMqVjUCcVHOmd6sHbYWgqUvndaMuj+zu
OnRFLt/Trs/UsKRmb1IRBqnfCPfIt42QSVy//P2k74U1BUL3whWhDr/PFklM51lDMK6YHBGlMFLy
kQZppnnrCvotUwLiuW4YlLGY8c7bVWqgNbUmtz1rv4+20O4PEaUSzglEwIsUFE8pGLmfhRoSVCb1
Gnk0wAf/7vkTSzroRyR3rouqVCMSNg2ypEF3OzBEdFzjyPpEHMG+omiqEjB34RinkI4qdhjRtRs2
0TFSiAiyf/2+vMt6dq2VpqJgjkFlAE1U0WFCl7tsEApB57wNJ5CYfP2I2TZtH6qrOR9FgghUIguY
qJfxGuWG1P1Exr330fEip0SQukGEFIvB9pz2PBGec/Peuj4bK1oRAlgBkcc5hTU1pkani3ZSg8IO
VHoeaZotNEPUCVq6LN30GYzhqsVLWaU4Nw7HbjK+oWrPV7/Mol1qu5+51pYj7yR7UPmTW6peorln
PhLrRICz2A6Nm1GDKdtNPOggUhqP14xyRQKp4RtDft6H2o4PsNGhGTSohhJex+Tq+Q3pGzXAEWo2
xho/qGc5EvAJVR0UIeo1mCD5UAev5yfZ3EViRJoZ0Dp8eceVyMJPQCspe7lcsibZRYgNsCGZ/gO1
i12rAZQvzzWHnm6H/I6T/lSFy8nO6CUE0CWnVPDehACbzaozjtWvmA46KxP1Um+QLJLNO7+lad57
6VX5pvYCEZ19ZRCl9lYY4lE1rxyxEcp+Xm47BZ/cqzR0eMuC1HzLJqgDzaepbjkscgWpvk2lIYAt
KtMCyRPAMyUoZLKBFlDdrItzYW5zL4nPCa/EHbFtNAJOBW8OvcOhzFl/aLHBa2VJePI4JCVBZbxs
T5k0X9kxnGJPUEikemutvF0JBa88uckw+Wcoo9OEcn1WAhJRlTBnIQ5nVtQhEqM4RLM+YqE/TfJU
4LG/Zl7eTDPlwfy9BlYPoYIgyRBLEyGQ1yN++gECr4QFLhxUS04mHlZdtegQmtH1V22N94T1oq6w
G1BRYMTaDmmyNBio3+wc0qjcFjsHKB1CLKU5tfTMm7vccnwVKvIuDLfdeCjERhtMpVyhwP9LSd0y
Slm5zxeFMH1J4jzv4C8F/TlUkROiOYkVR8Ek+4BZ3CwfHVpRRa0KyQXqNnUPf6qQKtyOyPfhtAuD
H6wgSWm7aMEbxbH7wJ9KJMvUCZGGJ/xXMD1PmPYYkSYtM8NthizRdL6W0w8dC/Fabr+972mIVUx4
ucwRLG9OYViNpwcje2S+JQS/wgFWOlnqagP6HwOw57Yp04sRJ3pJ6IBod2tH9L/3ImTrgOtcSrj/
o26EXte3+BHRINyKpadk9SKzi26E3lO7v1hIygGqbjibtyDhpqIpScewCuA/yIXdfKhPnckKU5so
p9yBtvSaKM+dD642jRkBswbOu6OKvvk9b6p1B4918QxwgvpRHprGART1x0aIO20Nxb5MQJD38BDU
iB5KPEvP5TrmY0tHBO/CYClKu0qQbIlbnd5eFIZMSfFEv5QkOn+BJeltFULN+6+eFacFM8SRbdiw
+bNsolnqO55U/FCsr/JkHaeUC0UBQ9AshK0CbdkJkMoq+ucAk/NPKKOv2hthgO6S4QReSJ7RS/Lz
qaIOiqOJNaiBj8dBQ+yvQG+qNYfUIwNdeBCHIGMUGotHfhDjnjuM8MOeW2lChxlWeTXzZhRmNfcP
lEdE3mJVj5D3kK941mSGZyVtDW6fQDx0CxYEjsh25PrRIOFytYjJj7vnWmJa94VWu0gLAsjRsn57
im20xd1OgUsymZzmIJkmJdGFz+RA9uuG8uDZ5t02BaVvmlzqhLFG5xekmi0WM+Rtqqn2SsyMgtVd
rOUirJ91YVdOEZoV/rod6Bl612zyXjVmj/m8Jl+V8ksdnDqwz7vs/EN/FIt3YYoDMHr45QH2ynJo
hlG+FMhN04cZbkagzkQB135hHqJm2EZBBEISECtgEE24eNoNhFKnMj6XvrsXLE5EFs/f+CnaLngG
EwYrljA8UsYqkSPym97lfQ6Wdq7TatLPdNg9U9+lR/EInzFpdfVmT+mygBY2PVjIAGazac7JBvPp
xmfmOCBtpcKtUbWwFdWeOKu31AL3HtWjEI2K7LaiaK2KZopqKum6go9ApQK3P88fYuYNRClNvpPw
ge1kamxiHQHb0f2DjqenZYTMf0NlDOsEkDYTl0V7iVaUyvzAEuERj+CxF0krgiBUuwgHQBqBskMe
IAKoeYc1Dyx/ViYkPfQq4t6rUaKFBbeBsvVqxWza4mOrD82+JiH7CxcxTg8xq+/AQw2fMeA5LQ0X
n+RUichzrBgX81Sg4XWrspwIZnacEkjv40fkM68Joc4hUeqGusKfMXX1MHE94w9l95LXRsrLvMjk
NRxlnBwUKibM/Scgn7ik64TU31TBgM4OmEGb9MjMOeFaWIyQG83LNGjWkEnDuvrPPEo8H3T53Y/w
IfpDD6b0sgqUZ4Q5r9XYg5kiaVSzRCB4Oka6AAodqJ7hLfdCte0i9ujHUoV8MQ0KKLDgXbnZjKAn
Q1g2ZdX2/k/sNGaKP1vTNqXULGomA5E9ox/zDS4aQ5JwHJWcKDLO1rJTnm8vWDsyrxSwzTWXS/hH
NnBbCXgTnEx/2qESz62ffuBSO6y8ZWts/dhc5S6/IcOMoZuqa0ojJxqLEx121EhDyeDfXLFZPS1a
UanXE8WLNyokiXEaky2BGaVdKOBcvRKb5zE2HrWhmK1eqYVpjjJpp4E6q06F3Srb+QORDlSaM9hj
vTZSQQyji+37aJKvQrah+GJxWvLWcBs94gw2cpFhAWGGakkjRPVab39tcs/q5hcL/+HvuW+MoDIi
bMfCkqFaLvWlxySEJDHXemKQMAf5at0Yr1ea7MOa/A6nqszRxSKh2xkLkmg1IudJkuIt0LNuka2V
wciHvEToT4hckkC6+z1yzAO5oj8PK2mu+R84zPtBPklllxjHyJpPXLG77muI6cEH5LTIRxAeiTaS
ce7JKnFPE05N2P1J7BgmkDSfBz2g0J4Spy2V5n2MUULYt8R1lNk5XyjzkVuQnQj9LqwWHwwyYOy1
d/ZWj6/MKfgsc0581VN/Sbs+gWPHATFU010hcmf2A6L1AiRJW7h35anjaFU3MJEereLvqW4Vea+3
E9LRLG1wutn8AVKDkvwdhwyHzYKbtcH4LLwL5AB/1LZZOia4VVqUnlNZVcs1+7Qh0KUJX/m1pvu2
qQwz3APbhVFgrloBMZe7CFm7+SmHAQLLsiF5FHADbGlcm3HTxAigDP6wXJB09sUuPWngrZFsKNB2
MiqJOFegSk9bBwLVwjDpeYpM4RIysCg477Noh4pAottG/sN5rGVx3AG2BmxBoQd+c2IHAjm+7il5
ZzKNm7X0hcHz0sklLMqEttQMuWluAQF2qjf/EyinfTFQHwG80NhmaTejvJbt6tsmx43ggbdGErbg
uuGGr28WIB5LhsfjijNmXwkk/GTeHsL+u1r7TAZLJuBNBmAjUv2rDJrrjK5g4oBkySq9yDY1iwb5
8uhpSso/LGMn/k3idoEP13/G7E1PV0mx2NX/DFLYLZVykAjnx4Z5H/xg1thchDpSAGDZlXN7a8mV
0UMSMP+4aAW5X4U7upArbcIs+nT0Jz83zoY6lCMvEp/ixIiBBaexhW8RKdEJzrU7c5tiTV5LBoxr
8sDKRbqcr/0yAKCIj2HzS8m7cOejCzfgFInDpqUK9jHBMBL7ah18gV4dCMRPXygb50N0oMJ0iA38
nt2ahhUafC/wWqXd675suGjYLrvl+O9OKjdMRkoyg98sVIKjUbvTMwgVXOlKpmASlTG5HsqnOSG4
hBYmKyXdQX//EHvKncbWoSWFxYFwimhpPkQcSp4KJ0Rq/3vOiU3Ir0+H4f7Kw36BEpbEKLgMhU5g
rKq0pZZoVDgjHk/V1bxUYOl/vGzr/+DV29dBB+O+gs40xH2PbfuVq3Xpw0rtospPyaGT6W88juMd
c1lX5XkC9inny9+uaUJ8q40K9Gib2zu3nwK1zxYywpKOBSglYb9MUpJpKGkHhDhpS2IQfD4ivrww
DtJUSxWHUDkEKANX9r+9TiAoq14OtAC9n1ysDSg/bdzXdt6tQjto4H4TOW44vDgdyi2r8VcYUISV
+C2JDAN4+cR9yKcLvHJ0KTSjKnU4SvXm8hvNGYl1M2Ep5Hc/CHaDfDW4gf8Z8yYV7Lm7AQdZrk2t
0iTgMaYU+0ZgPdoncXM0RITvkACmsJbhFOzKWDKilapPyICnnXL1DuhKGioyXI3SIpSEQoAXRlZg
kYXnDGXWjtMqDRPSENgRji88Z3+pa9AAK988u51CsUu8SGHVYqTcGjGzlce2Cc/ychSOSWK0z6E0
UIR5sX2MPLk3Hm9t5HeovyFJvx3e8Zk2uU9kKuKicx6BAs9BAtk4ARXCBAb5FySu6bWB5Vl+6P+E
fPgXk4SsB51FXH4mYsPQqwaeQypF2XHeYbkkWbZ8z5g2kvYcwQUx/ikODIzFC8U4NmLJ7U9nwZIS
dSYPjE/FwiemgLcje1F7Sn2h/e9iH+htO1ac6Oc0iXI4fpzRNj8TZlS/+5hiiWToNNkVENB4hZLg
LV6niSNXx5VyxJKWHZQIuSwqS8MGqqZEbPJYffdVnFm61SKV2NAxy/zEPsKN+bqhx5RG/iSDCKCY
Hc9bSakZRBiVEg3d35w0BrbLH152Jqeis4I6gxWqwWUp6cJf/Ch8xfzGWPXqg2/iY/Zwj5rka1vJ
8aWsbc9O9j9Hx/GiAg6xjy5BoMji4OKKSn7Lw9DqwU8OWIbog0+RFC5zreI7s5TO9ciDxsb7O0/x
u7z6n054RDs6fIvm63hX8b8mP/4LsG2RgIS7HGGvW7motV3R9zAEvF8KA41s7frTPstWmP+fqfVD
SAI3d3JEcp0J3wqiSn8k9V5mQKw6RyAyyx0S2+6zwT1JCXLEaYhXo4HG3M0Je4o3PNwMrv3lIdAY
XPpuYczJBoYO+CqZ+JhCgc2n1e7zptd64IcsOEZvqPflFHMtCfzzl4W6pZCQrmEMfrNsPoYAaGMI
OrwnUwp/FLNrYRzF1j6akRzy5wSrGBQBIoQzfswdF66MfcN+rBtaoYnW3AzBSmp+4EI8ALZguSgR
7omCdpCCcZxNaC0Kw4AuAxJLHxy2Fn48QCNewNLhWzcXUxhrah+iVFiChOooIy+uu8YNSSd/Y5Az
AvRbRuV9oLngJzMqMumJr0Mv3N+lryMld6gmrvYsFQM0Ar8cLqgZX1vDzMJfY/1RJg8OgBJ75ZFR
RGA8qCOUiqRYCLAP+XgCie0NEwxbf8bRPWZ63lpESRat8/jMjSKHS6DH+zo6AnI1KEbQqMKLAcKB
SfAmKtlRkQfI6X07Pltl1FMvI+8JuC/KXJWaXo2bnwm1etIOCLWLEG7hFDPvNqHZDpKJA0LSJ26S
TFX7ybm3tmhmnbZDg1i6uWCuEj2AZ+ftT1o5e9E3aMjzdKD61xgTFqJIrkp+KPSDKJhEL6H5V7/R
BMS+2lmtrWJDuhFlnw9hiQC6EbGpjta1pzFR2Uce8JhAXiXFgrxqe7rjd6nyD7wL9bO17i84g/k8
y0BmJc6XXOKyUd6fKLe1IrmqL+PWyFRxX5SzCyhT0EJAKd0XX1tvz4rFD9or/vLR3W6UUo9ezngC
/MXqRohQP3a/+OwbwXUPAw6WR4IGuLaAaxo2vtqUFEA/ncs+mzeQzJH8O5LVL0XuEK/nWlxZoms4
wfLySA76nLL5AQLPaAFiam7Yh5sTBtbSSwzpshSrR01OuB+wmjqFSe6wJmvIs+JcI4kFRTprnoI0
mcxaV3W6/M3A3VyoQDP3W6BM2oIi+NLTagVD9IS9wWS3hDV6GgVAmxmPl+PafLtPw4IcowBmZRX8
deAYvBGIi0CS5qgoonN0gumqdPmxnMbWnmnvGBtOSchJRCqydqHaYqjvmS2T7ylwGRZ3y1HT2ILe
3s37P8Pxe7U2Z5Y16TvTL+qimDNQC2fqnNlAfNGSOugASEUfkcAiortwjGN2Fc0RibkWHLA8qXzs
0UGQWdkDYMiw/2X66GidEkJSzobEVdya6UrL9FcdDoMLCkSYLdzv2KVVqAn3a4iAKTHnS9JS7scH
zhyaQ1MD954wAkNYX095u1gmTVBAmrstEC+Cai448xiNvGrSXW0arZHt2OWoNo7KZej9ILSoQ5/u
zfYz1qFsXuhSU+jjs1IvqzpekrJcM+7tsP0jdj+j+JqqpKhvp66qr6CPyJll3bpND7z/p8feTYfM
ZVDvgyjCAy9GKcmOLxONOZwXmPPwKr3bAPSA1pTjyUmfdq8gBsC+ZLBa/B6CLjv+vlJkJwAh6kC7
Z6YQ5oaVN1tMDQ5h9/9KErabbhXXkW1yAMBFx/AAmdItLtJEWpVUHZ9ZoxdyJXVrBN8bqNEY1Rrd
oGeIUo5uObl4oFXKEOcTuPzQRox+STm2zGCJ3vLeCfCG8ipr0lRyVCW5u9mMTizNnWhe5sQUzVL7
Q3xBQBQCRxuJtkTv883Uiqa7Nrp6ykDusPn5dt+sjeJzDP19cvm8rq+y0Xe2u2Zo9Rvl0cadGuRO
6nHGCaKxOkqDgXsBcL5lT1Vm0eUWwJXRWmDdb05mAeg6usODsM6NBlJ4/YPfPPyE/kov+HzWV/24
NEm6sLLsIfRuNfuffV4s3QDG2yHQh70ZzU4hRjfRlyVJfCKBq9T2ei/7c7V2y8wBwkKn8hssXTHS
SH3l78CozvmBaviM7uymcd9ySELcV8Gn/H7u4eiSh9DC+BiXT5QL/wKSTKQazJAeppua9vZVhgWi
fqZGQTil9f6yw6wMX4UOyvPEPFOqpvhAtp4ovteQmwqM3tN8d0V1ASlzXI/tpEsEoc4V3TxItf4Y
IrI6iBIs6FplscIstiQSax+mign8jpfhK7ZowCAbl/i2/xexJvhiBQSIh5guGtvIb+eQ2sq7GVBa
gkYQWysv2TqO6eYbCODSDIUMJV8lCKZdQZSKtvVjcD5KCjobyBfhQzFSW0PkFUNXSnICbTftkF/a
tCTrtl6ELkvRGZcwzNRBWJ3UNqmua8Bd2i1tpnxSdU3F/++iStcNSZVBe9I3vaJFNYyke1N4fP4F
04xnMVqYMcrHMM3pNck2T0oYltcC8C2EnIXDqeFsaKfwneor2MbRYDgo2voAasTMCFTsPZb0T4FF
R6+rvniaDTBzD89QRfYjJRW1lQ32FI923BRBOpFzKYoamy9SKvRtjTcUdaHionifGRbbpdKjpq+9
Ox0IjN1hUSL8VwOsh3MPhEV1jnaGXc75qd+WdhYObKfHTx0cFIkiAEO1smAIkSOdwES8lvQrEB4F
UhSUB8o6gvIMBaWimFz4sDQgcnU6cES62ciKTlmco06Lw4k4DQYVMlaTHetRmS+d7FOk6LnP1ERD
MBKkic/xpuE//u49hFb/44XcD9QIJDdJzgPZSOqFAW62+7u2RZIQbTtf/46BNQ8/DVbGv6qbwv44
XdRit2nuQfPp8IY8MlcB62XO9Jf+5CV+nSs6WVWRmR/xlmSiCeXCaRo6e64kXVXFQSORjFit/xJo
H8/ef4ITRtQX32C8hxrQiWTD/mdIqnFeTBSII0ud51Evhk+qVQj+5k9O80xUqUyZ4jT71susI6vI
Z6EgsxdQRciTy3f8p7ZiVYVsQwHYJd25WYIjpSyZsUeTuN5QI9xWKAedG41M8Ws1c/PkZdQmW0UV
nehSP3dvXismOLKrep7XTLB7kdiFrEiYTGpoTC1G87dAPupn6AYSBqxWVF6q6Rg7OdKpboV63mHc
VblRkfCAae67q8w42ehnchXGZ5fla/TkMIMuNtxollyhH7E+80SkZ/gZUSpqk6kqdLk291s0K52J
9VkQsqqLQKYsZcV2VIUF4+vlYtRsLYgGScNI1xvRhJcQQ0d/Tkxc81Fq1HZ/i+J3Y8BytfXLvlEa
nqVV82VZVLGPSTRUOa1KnuVkT9J6/CrovUf7N9+KA9jr/ToYMNJ1+sGp8cN3x0cdtyJVZnBhTgps
+QWT4L0SbaTn4POgbVoQpSNBsuBnPgF2jmGspZgMBJ1OYaBY7QJIctEGvjW6kmCl1vDDFCSie4m0
OJ6otigpZNSHBaszfbAWtE9hJjPd4wicmohLC87nK8dW5WofUrXr89JXQLmCq7MkthyMqlB5/uds
huBo2NtuiwxL+M8aFI5aBERGvgORacMLyz4kyBDsbvsc9A1gH09dDteJqT3h21TeimC4jy9EkO/P
ngpPdaX9zvpMsMTpfkQ2qn4ky7BkBCgWfeObbIpxZSzKfzNE3P6I4JDyDsPcgJk5vYezIuEdbW78
yfyjSafPHWnByVrfwXo57pa/FId6MHGuVnUne85HomXb31HeYPKJO/qmZ1yJxKKXX95Ulv+RGtqj
6SxMiZ3X1XfshxOb/gm1mh/7cbniNf4PIekauWc6/UzY+mNsuYpzHo6lro10p9Q+kf3KkBOqMqu4
2DfcM0ycbkIxI650vecGXyYu31DcIFz5JcbEP63YM4l78v6S4erOxYZ7PJEiuj/817xQT4SyOxqE
5xMECcGcz3XTet3iE0IQ0TCfeQvkFe3Gxy/gUwGvfe/rttpu59W0vgITIBsEPx+DXz2b+WEzR21M
LGIAKZ8uxvSyUmDv7AdOH/DTs3Mii0f5h5y+3ErjsspQisYCkHte5Yc0rZU3XjyNSWNqBkqzxbpQ
usZIjj5crn9UYNwFd3GubnhB+uFKEHIn6B+wA1U18o780o3Hxrkxwkkfsp/lwXHLmQpJ1XirDU/T
HFbDSmHHZS+k0YjoWpz35Qr94zESgemN/hdwG7CkFXm3dcJcNP9K2lV9my3xATxFx4TbEfvG/tcR
hPqSWNDYH/duUv2rn0qlYWD8G6uNkXBmCfzYmueR8xa+1FwW2jeJCjpfY99QkP55cuGTRTTQpuw8
rkosrQpSwAFk3GhnbjxJ/NO43bTqyxHqFDMbJRxfBZJhhHh8lUnz6RG/UzdW7ziF3eO3FnhUEdly
B6UZd8jU8Z8c4O9XBSnlJ6Qc/+aUS8VZZ3WPLfSyib+Yo7ejuNQL7tg1SwG6yeJZg9H19xSUW7sH
9Kv/ICFMkfCpi1VaQdKFip+F8RlahnRaRGwoCakv2rwcyhTgtEQhh4WEYu9KfKohNd4yUTKgbXbL
qTiyElDo8NPUcQc68/ZAteBQWpGFdrV2pT/6+iOjlWNqeE5Wv0KmJbe1iUospw5F2B5m+DRB9DoS
md+xftfvoukpXia/ls9hM39wA23o7Nw27pdcCdtxYysSN31J0nrH9k3BGjfOExPSdIcRnULrTu+O
cCtmgq9QIVRMDPMc9S6uN0a2U902EnY1D2aDk042ng2LhHmBalIVMsKBvHpaygCgS3d/q3ziZiz9
6BHYpyJ2wY/0lK4X+fV9HfMmfxJ5jwA9oBCOCrdCuYm7odlU53I9PlqDsjwn0ZrE5UrbPYtTveL8
YOBpsqb26J0ISkfmMn6CTEgh3sRH4V1vY+skRSJbX3kQvD0mfHcKioPoGK/hS8IuolSzYY5ITtv0
CIJtZP2cpXVL2msz9aBd8dUdidfqs5RmrcDMxMOS1ijDSOKaY0wkCNxOrl3c6N2T3kET3j36pR8z
IcoKb1S4jIw/IiSyM7CH8TMFzFlajOjDNqdbvWWqDZ73LaEX3TfoAQEXODs7FAflnypb1m4E0zG9
FlOEDQqir+4sxt81Mloo9YOl1EL+O3wCnNcMugsBgEPkarO7GqPAWXppatNRubS6mdQp1VXBjOf9
mCgwEHojO8RMZCDJ+rTRf6J4w9IZIR+lMN2yEQZ1CmgRDpBxOkqnOb9pZnCVi6U5+hYEijCthHlL
2dTXLpBWFp2SodcYSBwT41PimBgpodjskWkAMSQqo7yLCxdFsPVwWf0H1NQQTklSuGhueOdlFhpd
lJFalZLE6uGy+BtjMC8nLttxJMRb+rMjf8dHMRAtxly+dKSwYA2aKykXIgU/94IrKunDfdKY7lxc
WO1MTemHCnb4CEp/c+V/O/gR04K8T8011GojTYty6VqVBduWc+AHtY0nipFofqlPNc5+XVTcqdlw
J09OxenzK6lUKTU0ujHrDP5q7zUVp8qaYqJc68Ewq1FqxIPmO3D6vqr88olZSDl/X1qmOhTFs0fy
RmQYO0/trRPs6RU13tjsMSp8NWfsn/uu7sqd3IYMwJwM21dXi4kxKTmercq0QVjjh1dbL/XFoVTS
Yr0yCxvOEVQGCaL8tQOhVvbFURc73nf75sX3QcpiKWctZhUo7XT7yszUZrJWiFKAFkDVWMZNfuzk
vu+2aTrbXnosyGmdCMSfYKJz4Er+zpyjeqgqcRCR64mz25ZkGnZFAbvX82xQtwyKJMzXtsjGqieM
RQV28wzVPPWtJI+CMyX3GEqm5oonqru3T8xMwcNURxprX8pkSV9QogWGrczAaCjohy+eZmJatweu
s1aJcPSKwZkRVdPzBs7YOK2GR8vb7fEU8nCABohg6QC8wWT5LdQSgqBPi2Tjrf1Jeg+t0abidAVS
rjK+lkjarPJJ2VwLXqL+ynXU9Z7Tp0A3TXECN+pFX8J2Up95emoA+k1Jx3wOvpXJ9y1O6s787sOF
8fmJ3S6Gzyn+ykZUkCokoRbQxADDAm3G1nWmoSooBl+0693iDEMj37CyNpO5R9gqKZgkR+q3i6se
zHalgK7/z38gQ6FqHs+jYqN5B9/y/zPGf04PkXA5gvmyKbCJSqmX39iofEZrwt+p2YDUr4pZTbcg
8Wq2zBoHt7feYFkP6ANlCQ7SSjnGjImFbuxeNtQHKkTOOVhDQVRHWdJsAq9tssuMVcbf97IbVAXP
lWvchlE0bHH5HjoiuorOZJVIuyA8czEiox6ZypNxovQQWJFuD6eVunPllSfAy4P7XSSUbQe5hBie
xyvQIzhyIQPivOkHV1uLvCCbR3oNf8HnZBM+6hpqerXbtUgVkL/GPjtxo2963UEZ3801zl08SSFc
UnbBfET2xSyx6vSqsR3j+z2U00wFX+tXajenL1hZGSEcq5Du6cvkV8DFfsTGjRXdwbIEqMRedAx0
1mgMaII1nqzYB928ToF40i0uKDdm2fIf/aSqhRylBDfZdIv0BJ1oRX9x4wt/zC//gN/whA46Fv+h
jCC19ge0DfYTDsgkJdPAvPG0ihaoRdzHb84QB/nW33NmxbhqFa9xLDfw8MXglSCy5EjxbxNFpNHJ
rAoV8eXNADEwjpx91UIpt8bZmuZhGHu9hX7R2BT5/HFtOgieVsSEkHGEFb8544OOEuwS12UHYIa6
vhwauvZ2WUPRFTjjTjeCxy/52N3L/dudWBvB7V2B91+V8QtwtmTm6hM3cRmZ2QGJRL+6ZczOTJuN
RC+RHSLxkm5MO0+Fn7MG2yxhFh+WsdDP2ZelQwqMcBBODkBKE+bAhlA8oBfyLFr4eR3sKg0XykYI
Uo3UNb3/BRgMRxKCcoA8Kq8hTXOrh0H7BRysNw/XeB3BvPAvADlPeCmwUQ2VmC+/BiKVC3U/+t2V
aEp7hsJhjKApXIEzV4L9lVD79fpVxMj1HiNy6TcXEx+UO/G0UgD9rY/iJ/3eBJBo4I43kwIUHZRa
eK0x8L5vV2GoQttVJFvPPr+xJK4ezEPryhs5hXoQdmBtMrE8YxSGAz2sMHGbC5yyvJNGsN87DFro
RtQYQA9iphL2OE3i22365TTqr2tPONCy0jAtsEvdDM5xk0LBVHCko3hcKv7ODr9ZwtaKNgb9fDXS
w2AMqUOzqGjOe/pR42fVmgqWlz7T/kOqulfQqaEYIkRiH7qAIkYajf9cgbRS8ZYGaPD0zz16hrpj
DpNn5dzJfoKeo9r5cwlonGm4lgcfmWADoqnetNLod+odN+lnn51VsoVJB8HgbgCI2kRs8A4amtzR
PQdP840qdGhYj/DzMLd3zmoMztrYzfJ6jR2CPtLBeqmTDSGce3mNBhdKbe9lY/EPuvW0taQRy+Kt
VkKj6YMJauoAQWoAp1f1KFv3vADrIKLKo1IZ4iYIzgtEIZxmPbgV3sVvTBqLYWOBFPMbXhAh7TLz
4g57hWQGSPba8x7/z5+h/mJ9datuWd2tN/ar07kS6nWUWhEyZmvD3G3oRoUk3CbQJitXNnSI+cFQ
bwkL77crRz1vSUH2sok8x6UA67VW/fDUz9Kw5VpYdoHc4L5zze64/I9G+Ve/TLUQOb1azgjIGaqj
kHtBAJkXjYQ8LkVMCCW0Jlidg/mAHjEViTVJb1QXjb5fW71AyNlwFZh8lcfKZGoXBjX7hcM9DhmG
pZhnOtk1gZoqywx5OWnanJZz0tgLSYaQgzBFsbNtP7mo2014dFKkcWz3pmNk5mBPESB3/hiH97lF
o9pWwmaojXNE+EN5GPk4PAgbZqIUrKB4YsFZJNnn05AQms4JycCeRyHlkloHdWCrPz1L+/RyTTNa
GJuA22YfBluxStTxZI0UKPZbIcNsW4At8ghT4ytRSJXVECcebzwxnDSzv4C84YgYWcylFWLSmW25
mW1Kwc9G+aEGu2P79Dkxm6t4ASILxk67Qf0tLIx2qltPESgjK9fnRtntcSaZaakJcBkeYMWsEBo1
ctMbbZUlUR3avDcHiafGCgMLi1FzKbEITRix6UyCtsC1lGoCy8ibx5tDIg80gLxO9OrRt3wX+AEf
J2n90+SUL/FWbURHAQqHIAoKx/4jPVozgy/a6QNnLpisAdAKu+sGhQZjqqFM2B87+ao6MQmEM0PE
J5WNot1+8Vnqd5XiomGfIPwQbHxOpoG9vMm/k3bidNoRY6s8AVqZHVWdYi+8kDcgFImYayGFDHWP
gJRg8VGy0MSX3p30ZeUM3BBORdfIcFy3fH6l6Q6RGEGJnEqOqBEAKLfWORB+8qM9TbKAqramhCp1
Ba45ZV4bSlwgDwcf4an0IVkk3VQH6e59iMPV5oLeNZx9XH3qn6kJ/pOb4ToMBlHD3etSHlK/EGS5
P/dDnHDhBrYKObDInVA2RXYDhvSVpY8SxvsFCaokEBXPEV0He6TF6XT+Z3Cjixk/Pqt1nNr5Jt3F
0GZD0jwrVzeikwSQsptv0Ca/ekPEOefHuYiC4+sMH7SYEbQdAAm1tLTWgqsqu0v4jyC03yX/pK3K
4GYLrKAmOcpMSVRUViAdwBMxZ4UuP8zDFE02NuGpsIAyW9JlHz3qHryVXSmpV+JWtwkdXB/WXhf6
5y+4GKeFijfVtWd3DN1iRnk0xa4Mbhl+016eAprAYa5X7zpqvPk8hoEJP9a2aveu5anTfflNs2Lr
tTk4H36cDLpWNpyrtr0UEviGwLvsn+A/dlE3xstG3ASIHkQ8eYp9p7eJLeRWy3bqZ6CcMCewlZQq
omNOzi4SItCit6jWYmLVE9aUGcZKaDUjhOHLGwCeJe/jzZQBfH6jJTvj9ggUky4jo5CSsI/yjxXH
NXnRePMS1hcB+mFVDT32dmYJ3SV5xM1xXzyfZcKN3QpQESG9PeX86HAq41u3QVfk8WhR6E+1F/Il
dTqDlAC+CUTPZBFeT582wTmgKQF5I0tjwrMrtNf4yfAcSWr6Rw+W5BzcbCFL3ALWvEkkyTJrPOUG
0TkGSflvHpoB/Bahiii1I1+z35Gln1vntgjRbbIOREfOPXrLYyWF3gInbT8Hw8BxR48X4xCDKGCd
oFeuIrlDDkDaWHwCLgiR7QzlOooe3+OgQDqQdpr/gxblLT8GTJywUbanXqSTQec00i78V07gAeTs
Nj2gbgD8etsCmUhRIS+ioxJ3xQvTpS+nlEKLQLD5kox5cvGz5XAHSXVy2QDwV8rKG3d0ba4vXvVI
rj3UVsvrAHqExkBOIDlj0YoqfmeNmkNr/ppf7rYIebsKdYEoQ5kW0+v50PSX5nL1Y834j1aSVKNY
zp2a7XKPoioLjKW4zECV5eV2mtdm1qc9MI9Fn/zDvrMgOZoqnCibSLIuSJ0UvjFbHObBUipXUA8q
vNyJU0tBxQezvrT1vKCfGv3cjlktAR2vUCP27FwBDWOd+pbgS/O5NZiszi+s5sdFsYQonwaHoePz
/UYFazQmgMn+a4g7Z/nJiccG7olIye5IJXN8J813S2xKHOHx58T+KvUzKo9jlnZODZnRvxWz7Diq
9PdDeyzmFZd5f85Bm7yAO1id9Yzia4dttn4u4/XnYYtUKSxnprxY9sBFU+P2O1yTPu2uKJkHBx8+
dS3xIrL7fmryFPcy1Wpiwo6lDX/YtnnK+dE9gS/pfdHvW1OfdWOE1xLx6kSy1MDLf1FMSLqUlt8g
O/Y2vSWJ4rc2IXs6OMjMJ5BpW7NqJX5znFL8cedxHaRD+a02/uOUtK4SMfBXip/wz81fr7oegTeC
XiOcWXqKKPUqoMbPTQfTYoETdZ4fwIcPLv7/vE+E0IlvnRNm9QzyLMm1FtApyrIh+UeQ6iOLzOpc
4vUqqJPYeAIn3/QigmQn4y35Q+W3YkroD+JKygSfjoNCA/ZIIOzRod2EVPvKllqJLnPCx2cvrVTf
KXL7SXTGJIIFCGAKgKm4VJc++KP1iWCzOXCTzgFjoL6IM468joljbuJK4yUen9Kqer/XMCa9dfjd
Ha4SBmxuyFSgeSC0VJ4zSEXfuQDTG8KyIGHjMJrUz46/XVc3Gn4WzEjVrel/xo4FE+04GZD3hwKA
QU8HJ4jNKAHc72tRC8nRpqiliHm+AUTJKAnxyxJznmwL1nMgi4E4icYnQUoBZUZjoQG7H4zf0W3c
FKvaPPjtaw0HCzi6n8Pa2rgdXKb6jImKBP9niiQ54tK73gCGfIAHvP9nghueZ79GNriF5ub8DXWw
wG+uvf7B2BZFZ2Mpbni+2ljnII//9XrYWSrevGGOUzmrkzct5CMhzV4f8Zzwisfoc4kH47YmJ9Ai
bNvnmta6GrAaj5p6o7TnzXIYh3BpYEFiZAi4YTxv1ynTMiImCoILDzIR0J6Jr8k1C2PT2kLwSyIM
D6oYlBIYJ6NzG1u2EzSBexLH7GCTpadb3Rm6qjc0GrBZHtApxm3GF8/y8Z84AMlgXF6qDCoVcaWl
CcCRHlQrimGbloANtJbQFSl07cyL8f4O+ypYzBtaBMv9hVzH8aL7/SJrIRpiXc9kEBifF4ZlyZyU
E3m9sf26SporjuBMoNP3ebjK5QGraTuDJYhuDmTotyvENyLI5FDz4LMPKjhN8NcVpFOWxxNNSdAr
7wl5M2OUx6OUAOnW7Hr7CtTUp2sSIUshE3oWDeyNTE7rJzAl3eV7znp/Yc5EN5abIJ0nvWgCZR9I
NzGxrahVprQ5kgJOAkrC9u3t9CMUftq1WT2qRbspij2t17Zsr1CgYM93nVM4P8hlf4cgD/T/Pag9
ym9PVXL0qAGZB5K7Zhb9t/3C+5XfrkKhMaBSJnu4uEnnj3xNy2+/QIpvLHI4PeF+Wxm2FmaG5J6Q
xat97dngLLFGxnw1tU1aYE8WkQtL7OjnM9NB9EkaE1+j66mV8ioSh8AXV6Rz5tRrHv8n6haZ+fp0
ERHzZAiOLnLjUCe1vMHdPX+K0+MKyuS9vxsgO8bEHKgeEg/Zs3Bat1Nw3guA5GJSmX0ACznBBhnL
9i+TL8et4n2/tLxAhiE1sHg59qkwGuGXXfqZJw2YCo2kRZF0hSZNyQ9aRYw89XuYfy0U7Jt1hPm5
DwTb3fAfkw3vTPmaCxos6LlAOjBVHEZW1vahi/rLZMBeUUL6EN7mlM+NjBcCqGjiuGvvmGTjXaNi
QiITkaCbzZMbxiGnOuP+gDbGV16GKRDRh9MzbCwZ4WjLDhCp/5iEnkQhjvVoaEZnnrxk4hToeioh
CxshK9ZiTnrBeXyuZ+puI46b4LVXm3YVNpmV1ZxcOE/BZwcvZP7BPoKXDh8FwoLBmfSSTAuF30fS
Qv+KgDt1dbgwWUxF53Sfapv8yDryd8hEKLXzuaIBhTJBHhzwQKCV6NGYe08LEsWLG+W5Tyu6D0RT
9H9TnRP4dngaIBEHxT10g+Qf6tTaxxJ96RdfXLk5cOYLYorzg3fInlZwRkxKM7veuUzoqH0k51L5
Hho8XGmuFegZM0BHthTmoAexCMhvvzGDS2w4FH81ZRi8ewP1XS/jHQA8HSI+WucH6fbB3b25wK6I
8+SXPaffiVpoAhqX5Ymm+5ptr97GrYoM4XLG+N3FGrhHdu1Fe34RjmCJ/dA2qYQgvPrNs0jGLbI2
CbOUM8c+DaAhcIv+YCw6ufnFacHBIe6XgJSXN0P2lcTDF4D3KIfMpBEf1ewJYvmdwAA4Nb7/sOKA
aTsCOoUXm+4CzxIRksR6hJSi2MkxneoMFqdS94de8TA7KnLMw9t6EDPYrZ59z9n3c2rmP2phu16U
rjNDUudqGl7+D+XjAPG6+gOOd/ed+dKcymdK2ChX6R/+F7wkMWp+3iHA/zbyVruyGAR0E7ze99Nu
59hMISK7Naz6/IuXmuw1Lao/9Qn4MvqWlJE9SAjRd7harCg2EurxDuIU2A5WqwpqQ3nkLOEtMI/a
GkLwli/wN9s3prJfwCY6u5y5/sSrUcyQFegm6brLIqOcSDKhT40qt7W8K5LqZaN4lVQy2Y/VF8NR
j8hNBXKvp2cW82TXJ8fZ0VfN3vK7sHA1vYVGNgpik9RHTzN9cjiNSwNhNJaioyoMZEXad7lzLg/M
Pgk5HW7457pnSNNRu4I+mcAvUE7+mSuxhXTonIf7UO0ZceZl471cQOePfbSvOXokb5qL3FRJohDg
M9IiC2+9+UcMLLapedoVjIUA0U13IPg5RvQf01OfsoWms777qvlpsdx7pYf/JqB1j9BYM0qAf7oR
WI8OvakxsYoIJDK40mFvQJnt0uPvb/jVosOGLtlde/B38q3qkDP+c1A0WOWvhJ1iDtppPO4dIj3a
XR8csq2sNz915Qa11NoUJcx7tkDIS3eMFnuHc/2JWxIiduFReT4Oxgv/LARkqZHyYJ+f2u97jr4l
u/IFcwk9QK5/NDVkV7X2Lx8FYACeznt44KBCo0xvoVpSmlZ45RzDTueMyVIqZQ22JJ/ZX06M4gX1
03LdkVrP0P5W6fh6Dfjb3DGfpKsBmnGmkSeacSWZUm2Hi8O9qgdC7N2gTKoBHegRWkwUzB5OBtHx
8HTOSBK0zuQR+EsXP1e0ZnMuWZ4ZURIJYtcD6PJzkpI8FeQnkw+j9pVJaVfxdEDv5E9TMUlxA0W8
fk9uypw+Fh5PKUWBNcXpXw0rbwSanK9cijf/JpS8ruCjZVnJHk32NpRkYzCfS98bhlKm9dxRihBa
GUv7bBlCGwAc5aU77u6+6umCaTerzQfg7VC8GZJyRn4O7vMw3igUKoSVKGwTSmEAHoKJJCYFrgkw
95u6BniHDbMx4Km/zGfcc2glpoQ0v6ZOuDh0EtFgzgU3Z9bpqM00yXovGD5qJYUdtFRKBAmlCSNh
R8iqOZEe9FI3HIDnxBt+BOJioteobezw/YMOqI/pTYFsn+ETY394xQgbsC7ZEZFk50OpILiUHIFI
UcyQvQrSTf0cytX3Gwq9sGFEoeZIU9hVs7TxAkamQgXuw6I+Af6Gcwt1vodmGmn+QSUY196+0F7d
tLbAzTXDBtbNYTHSd/UVn2vmOEJI/Ix/znOpFOmNR0EI6YKxFtR3meYuJMRXmRyXhSD4NtLHK/UO
8C3IJ1QlTr/ErrbB84SVZn70KVyNeZSUiN2rr0Q3ikGUZh18JVDmaKEHFH4Ev1PUGSJFANHU/Dlx
wqmpMt5E+jYgtR5p9b5gA1chCY2QYw6V4n9S7x/s15GuJaVE0Z05G7/FjBlpFAmBejVzFHN/Ne73
+F/wGpGuC+DCnBXI3pk6PBKskRW5dJlruhKIP4eGEmDjJ+F79KifBIOoGhm8sDP0sIL36RC7TIsi
HO4eS45Qn0pPOnw3hc/hBM/t0DJzta0V26NqBrfiBNQUKF+Sjm+r+BRj8M/HCtodarWemf9/h9XN
C9x50xuxPHs1bAC48ychkO+sQDwmVGKviYgCyV/oZI/hfAprYn42lufBn41QhFiLmBI+GwmfDIOV
dB0NdB9s+J1OlXbKMAZefACkxh7YEn5+55veL90asQ40aUxWC/BACPNsQM/SClRqBvqh59YWQYln
XcFqVwvadh3Vn6Pu3tJbosW1zUjK9hp41x8L6+k/PqBM9CwuOIYKbzrhpsQSql6R7Kf+5Mil6w6y
RNbZ8g6zDnVzww+bHS1Ct84dZfSZG61TZDM4w0hYqXpbFCt3hrcQERySA2idfEyO16Q2CqcKz/0s
vE1fu0z1Of90oiPc9EMvGkHu6r0yWwKaw46LiVVy6kXjuW75FB3mpUBj+fLtVRYhlwEJiAjANVZi
W6pGDk3GDx/goBv27a5sxMfwUO7kEKmzLukY1pCGWyYFQWEmwM1XOFeXhA09x4coMCCaEAUlTycv
6pYGUiZ4IFY4srQWW4FMYIfLg9sP37w4IFG5kc+aJrOm6Cyg+W4u2cj38fuNDsOQPoF8xwgM5Mw0
5McyI4AJtTfmNr/7Zta1syT70MWyg6ywYzizlDyjInFLgJE7xPyWHgb0q0sLfq5eL5rs5hLe1xzY
GVngaqWX5yulTQxC2WKyP/36MZp4Aj0MYgUySgmlpZYTJ5hNOGi+lqo9FmPQXfLpOxwczPifUdGJ
xwOlYPLBpBWl6ZIURK+hh7VIaMSPml1WF5xN4tSkdHJ07Ro/LLU/U22H2H074x0WYKD6eQ7zzkiN
Vncd78RABew0baITFb6wE153yQL1/R5Gs3397mK/PURefWmenV6rn52mUmhWVRaW9W2hPbFitNbQ
lT/2qgC8lnugUW47Pjkxk28QJSF9/ATRs/mEyuGZMKWaTK/B97QQIvupzKuaFX87FNxVw0Ass539
8SKsglMtfMSv+UOb0kZrwzuqBtMEGLI0EPCNSiIwjK/n7xgWqnaHrYHx9fwGRBZnW3Bvp80F6EkZ
B5ucQXqDzP3tsInsR/uKHaJ98wIkG6Up5xmt6TKpfQK+m1hi8CXWok7BloZIqpkyMqmr1IjeT/ba
V2kLRl7vJ0tCDrKr5kmUyvu+8e4wtvESByIG7b9/yTacneDees/jExzD5dobiWcgvLnG9h6wPje+
jJSafqSIiwmXd04/w5T53alsbVG5U93q42GEnpPxENBbUkTGx0NtLkEux9FLUdcQ+FQH320TPdPq
pP/O07DiVJ9h41wAhZ05xBK4o2AqrV58Ujs0UR0K5Dya6PLS5Y4UC1cctwnIfn5Guu/WAu2tXpRg
RCQ4aOSV4p6mN2WsldBxuYurNIsi7GQKFH6Db+b8w18UbstbVkPLtVPSgLp39vatXQ6LE3A5ny+W
zt1BRtXkEvHj9w5BCJ268FVa9to5FSKTAh9kE3HmnAky+G2z5/gZboo1dsf8or4aSoSnmWGiEi9+
txT1GqWGH9jZ418jAAXw7OzhbwrZQbMbkIy1w01nCEI0bqH62YT/3qN0/tj4qoRb1kFxNr5cWwBy
IpnCiMPiUlF+WXVha9UFbo+IHDznQrp6yLU6KvRvfVaDFrj46i3t9KxYaLkJSuagL72xpMp1WS9z
VBXJTqIm2zACrMNlIOfwBag7P+Brd1EyoRRSIJXpn0OeV5GP5h7eH90b7VsBAjo15x3dSaMyUvYj
yuoSnOK1vwogRDxCGGuK/BhIqm9zIkh1NnGkdJlzt6UHdq69uP9fy4QrWnU8
`protect end_protected
