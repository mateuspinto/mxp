��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���{C�%�P�*�S��_7@8�Jٵ+��Y\�����m<(��!)1��°�g$J�m�	��8���9�U"�����loq���9��Rl<� ����l3� &0�F���g���&�+�Y�z���Y�ZZ|)��~�~:[��}�����c{�	�~W[z�r��Y��1k������]n��ڏ+��,Q:� Q�-g���qOl6����>bs���t?
�|�� D�Y/�5נyb`2�u�E���d��Yz�{�J�[3D�^Hۑ�
��F�6)��'hᓰ�����������:F�+]��`
�|��q �Zo���4��t�Ɣ�tg��MA���ԍ@wu+-$Tx0� +��*[�~*��'W��YB~V>����
L�C]8����H]j�oɋN�2�t�HŇ2wZ���WH/q�
X�Éݽ��'v�� a�l��9�9��6n}�UH�j�u�{=_E���79�����jx�E���j+� ��,d���y��;1�G�("u-\���e��zH���Q*�q����f��1z�d�0OuB_�k���-n�o��VK��{�OE�}��S�� �O!An��H|�W?�:3��dd���EtL3,p<�E��w��D��i�"�"S? ��Y��7����Z��#j|� \�3/�w�0%`*��Yg5��g��� ��-R�\�X~?#@�����R���{�G���ZӰ���8_'-���0��.,D��0&(a�����>&�QK�����y����(!j3����d��&8(cWZ)���R�"�� �&mȥA�1���;ozj2��FSف��a\��!t���'#}��dh������Oo�ȋ�!�0�.�l��"q�P�-���~�Տ���������Z�{�3����D��zn���K�^��)5?���2�SŤ� b
������@�ɛ��vW���2��B^
�oPK��
�=<���B]��J����Z�E͹���X==�|��,�\�NI�ȿ@�onU��lHa8�,�	�;(�-oĩG",�"V���+$� S�@X̩�,�AO����ݔ���񀁫>�<w槓��Ԭ�Wf �����~���
���d���%[^�j��=�q��L�T����w2k�;� F����5��G�R�Fҙ�洤r�(�/9��9&Q�c-2Ţt��?T���s��݁�����6F�u���\pe�ĉD8��:����ґ@�����Y^�3@�sm�m�ݩ�����P�H|Pn�&�����6($iJo1�I-i%t'�	[���p�6�����ʧ-A�X�O�vc!�K�bêD�F��J��~o�.�ܝ��O%�����?��,�i�
.�RķӸ��m�^f�K�Qpi9�-��Ǉ&������1�'%W��#ׇ�'�tq7���i�2�F�� ��(��[��T�7% ����(�衵"��/���[ �e��zM,�o�a�W�a ��:RB�z�<b��8^S�Q�Ӊ��/˶��āf�͚�)�b!��}��ݯࠉ�'�8�7���� ��P�����R��;�,!=Q)�|���`I���,.�>��1MQ)bc⋕sє�/����gYfr�6�uy��_�i���G]t�����~v�.^��0G#k��b`f=���H��hP�)h}*+2����udO�N����Gۯ��:�X�cY�.����\REe��3�&~�1j�]�)C5L�Ѡ�%�����Æ77��_/{���p�4;o�,�d��Ш�\Œ���2^@|��y�k�4,���FF8>3���nN{h �2�	?�R���w�c���UP1B_$9���p}�9�����d�H˄�?��I�z��<Q�a+�g��8(a�;�[x��0I�]v���\XU�8��E)w����Ud�Ѽ��n�r�O{��c�$�	�3*#��G��QW��.c_�c�``�j������{��OCk2����6:�9�	VD�V�C �N.�i��Pf3C�{��8���!��,�v\��|�z�n�#�ؘXY{Iኚ4�L�q�5Ѳ��h���
���0�x�9C�J�A���Vt�����|?Ȇ����z�l(+QL�Z��r�'e�MWDc�&�>%(�E����|^X����~g
��]��	��w��P��
��ro���I�,IW��קSU��l�3�� �2QL���N��ޖ��+�t�Uq�0�\G (���7��
!v���^�8ۮ�5�5H���5n�_8o�(JQ�����)w��ml��=(�z)�_R�Ii�Ǭ��%|�}:��9 � ?�(πEw�O�[�yU؝��$g��<i�<����b��!m|��?'x�(��]"=m�ڤ��JŊ�*)S9�θp�Ft�M@o%�m��`�ߚ�9]�^qQ��s�`��%Ɠ���{�.�ѹ���&n7b���D�Hxؚ��{ 	��!;�p&Z�2ax<����� �<������)��%/��01z�X:����ܲ�p;k.'%d�q��~x�m.h�x�50���V6�1A���k���3&�)�y4�4n�>��'(p��YDM#�&0a�j,/��Jۣ;Q2�#�ݞx�"2��[FhԹ-�!�,-=�I�B7��<T�����P�!��~��@'�Qrx���<����_2����.�2f�9����|�ޗ��@>Ml4C�X�㖸��²��+�f���;s-���G�V�9��yG�(���b��ȭ̀��!�� ʠعdL��E2�>�٬aQF�~�E��&<5]�A4݄���;\ '�󧟏��!�ȶe�(27|����)��;%�7������J:tۙ���j^��l6����Kf��Ȗ�a�y�g�[����a���V�GE���ag=V��	@��<��z��ŗ��j�D��8e�K3p��9�[����p�f� 2Z<�� �ka1�(3N�į��AKf��
�(���{��c�K���,��nbON�6�W*�,{
H�fJ��P�{V !R����7���F������2�m��B^��mQ7�4�2Dl�%��D�k5��
7����T����EE�Q৖�I�$�,]c�`�7��xX��^���_�%�e�[D.�N�3*�D{��Ѐ�RM�lB`*(<)�	+���J8?���d����·5%'Ma�v7ga���]!_[H���R4*�����+��H�dE���zI��ω"QiwL�PO���u����< �!u�\�3��N�r�㵚wv��2=����6�
PaEZcru(S�����}ѫ�݆] .~N�Ԧ���e�jE7.ᰲ�D�0��Z4��@�)Sǥ���a`$%IZ�E�/ml&�d�r�f`�SI��P�[�~��m'ВJo�C�Z��F۲A�������%L7�Y���/����{�-g��&]k�Ĉ.�T^�M�?�g�;���3�/�����)#0H�qQQ|��-r�\�Sc݈�}Ƀ�r�e�9��V������R�(��ڊ�H<��#�:�[��=%ޞ�<�z�o�"�h�Wi$h��6@��p� ���T�59�*����\����+�p�4{4�6E˕a�J�4b/��QT�_�ڴҿ�sٮ`����#o~3c�Pk��яϔ�;�g���@7>d�+�k��zJ�����Oy��ZX�/� F��ӿ�p/+(�p,��,�h¼I9��E�X�[��a��M*�?+V�f>�g� �K�-ɱ��V𦿙D'��.5� zl��S�Tʰ�s%& ��|��s2���҂�+�� ��r?}�g�w�]7�.���@���̘w�����#��B�؅ﴎ����C� C6�ǮF�[2�7�g��&&��g�o�����%�M%�����-5�����e��*�9���	��v�E\�������Mݪ�Cw�O�妱 *dwo���T����j�>iqw��E����",���-�XްU�l����Z�ܴP_��=�5�_�=���x\�����sS��TS����c�r<	4Y��l̐m�p���*����C5�YW�f�T$��\�KL�b��C��,�z�u���-*7z���2f㮀� 
O�@T��#��K"��Hc�r{�Y��"��,�0X[�a0YM�-b��� �p�|�����7V�VQ	���V��bw�0�>�����
}Re�CJ�[��yu#�i7{��I��ی
�uB�ai��O(�-��]eCR]��-�����G��H���\�Wa��T��M:��-����%#
(_؋:�����pa��sx��Ȯ��j�I^�u27�?��3K��%�Ǆ�{mQ�N|�"Mo���a��9C%�c��y�~�%�ݶA�����$H��T��n/�>z0f��%�jL(�����:����K|�:7�t4wۋ�DC׻��f0�~[ۣ�^�(���D���D�'�mS0��D<��dͮ5`M�*U�D���m�s��.�q���f�-?����������yå��F�QeW��y���1W����.\6O�\޵�`v�)���1��V�-T���$�FW�L�~x��F��=�l�{b����Znډi����ȩ3�Xm�4�b/c�pqZ�S�Jh� Gۨ�����q��)�[`�[���l�R���-1��Ǒ���Y1=��vJ4~��k[H��A�@}��v���������t4V���Z�>FJ�4��$��\�ƁR �nz=o-�W�n�'E�e�������쨷c�B5E"��n�$+�?�!��"�!�Th�H}m5��}��FUp�V�gD�7:`O�3���U��=��ӓ�Q���*	�

�V�t)7�����Ob��H;l�~i����D��7,*�Pgr~\��E}�}��2�5��.��>�2b�)p��,E����Q'[.�S�+�*��Ҡ|-!k�#!�����ˤ�l�ɋ5g7��&N�P��l�Zt�Y�K��Ì��?a:��/ųϙ˦l=�ZA|��S�Dq��������#�;��2���'�;�j�`Z���r�����2�h��x6�>�[Rce�ܙb+��"��M�'��Lp�ň������b�RF
�Wz��p��9����hbw�1Bs�p�)��m���Lbt�G����A.\l�vm,{�@�ʐ�>{�I�ZV�ޒ�~�o9F��%�eŤĤJj�y��\>N�r�����fwx�ua���Ӧ�f�'w<��� GU���zdg�[�[���&=��\JL��/�o?����Cʕ#�o����'��
j��R���H��+%�K[\6v�׺�vj��A�()�����9�����m~h��km�R��B��e��X%a�I0�^#=#�ȴLp]���A��'^�tE&�Qp0ɬ$'s�nW)�N�x�'R�L�;iF$_�&k��(���&=,�������5�y�Tt��FC��{�PT���(݌ ƛX�(h�>d���9ɣ��0�#��Y�����),�����u:B�򀔾�#X	Р���ن��*�zz��ICRew�Z� o�%���E��ڴ���rS���{������%�]�a�*
e�[�w�m��D%M�G��}�Q/+ȓؠbl��κ�@iP硫GJ�p����1:k��;U��,��D�ny���
��饷�n<3�-���g�ϠtM6[Qxh&�p!|�"�րY�7TC	����-�/vz���$8��"�r��Ջ��@�܎���d��}��-�.%E(Z�T�m]��?��_�5��9��v0|��	4��z:�7n�ŭ=�=��E�~�C�K��&i3�Fب�j�����D�Qd�M��-3�H�{���IN!E������^�p�#d,��$&q�:��[��� }g�
��;mi�IK��P!�<����B���4.Ӡ���z*�adH1�a58ܞ��a#�/]~�lJ�a�jlnB�M���M������4�)�:�{��EB��Yt"	�}�i~ܡ�X�k��|��K%~�W�_�o�.�su@^^(�!jkj�ٕK�K��J�%Wo��K�cq�g�&���Vl;�Uq�Ǹ�r���$�����-�"�aok�Cms���b�lǷ~�5Zz����GMx���WY��c�����-��
q��b�m]�����C�kAIc�}=X���`�����F.�G���O@ I���&΍g�ug�)Ba���z��q_�uC҃�V�X��:.=m��%j�I���C �-;����"�qU��='��D]��{bx��&=;Ųt0Rf��#U���X���N+���ۯ[Ų���'�#��fB����[��jv�A��<5ڰg���G�UӖo����Լa\������G��-Iհ�����N�Hf���_�t�ӓ�*�.�72?�0��-�h{��%'�A󼇉p�.8[H>��3�؅2�����p�^D���JK��Lk�����;
3I���Ey()�Q��� =JU���fؤĲ����|��0ېZocŁ{|���W�ra�Vc:u0�B�	�[�fPi_�H���~�	`�;�DH},�#U��sZ)N_�#ݏ��7��=�R�||��#k�F�0gE~�4÷��㜸��dW�l�~8IDr���0";;�����m(lE�Pr�4�s6�~(["F�e ��2��o<W���w��+�Ъ� ���pV'�Hv��F�=�2�u���qd��E�8��vYfsKY7zD%�2��.������ǦYG�P���O��
�a�K���t�q���C ��.������k"�z�[�8�y	 2�qx[� + �QT��k�9��r͆�ͥ����:�+"�i1����M���2�Ҭ���"��%�s����������}��&s�4e4�2s����z
�Dde�+Y��QD�8�Ԁ2�׍�J\@�[�;������NU�AV֩�9�+$�B��#�t�-���%�Ezx���� C��VH�7<h�Y��q:��H��������VM{��Bd��@L9��=�X\��i�IQ�S�q,����2|	߯�Ee{@��C^�{P
0���+>7��F���N�m2�m���<Q԰�y.��r-FD¸���H��s��{:sW��Z5
�t����fE�E�?���|�'I�d�;� �jZ�j�����s_N2�Ɍk�t�&�@���s���Y��Mu&	I�$�"�G���3�F����	�~�|ědF}�������
L[�w�L'�!t~� l�O��q�)��C	R�-��{��c�@b�k��p�u	���X��:�B�Gw�`����jD���C�-h0���V�)��r�ު�ܕ,�t��z�����9��@�g]ې|���m��@�>"x��R`ӳ��i��z L];vei�����V�a�n�|��S2�?���+���2�w�[�ܟ% !��4�)_Y~Q�S��F��V�P�q�J<��?@��	������H��I�\�*�p�>�Īw%�h���y��T���$�S�D�yN��;���>������B�X~$^P��k\�tq&|�'A/YԸM*?A���Y)<h�ev�\)������L�l��>�%ȚD�=b[�|GA��5�9��lͿ�S��*�����ˆE�m�z歧)��q%�2����0��K��#�Zu�TL�%�u�t' '��n����.ҍ.�HHLt�<C�VG�Ɨf]�Ͽ��z��HP��|?υ�{���z�����3��Y˄���0Tu�c%f%����s �E�?��+1�%��>�%GPQ^sq���v�J$�c�R |��tak��cg5�:5�*�� 6@��հ���r�7���s��ŧlg�!y�D�����B-եb�W����D,�RKA&�pY��檾�A�����&��E	j�y�k��P�g��*�拣Uȹ;k�' a�A��=��l�P�~��Yw� ��x��U`SX���R�}5��Y�Z��M�� �_w�<^Qqn1F���a�� ��\4�1N��� ��4����ӆ���F��*��\|��a���"���S��d�-�3����^�.Wi}��yg)�lL%5���O�vյ��Y]&8�Y���[P��!(d����l�9��W�S3JO�WH��QX����¥�e�?�i6`|Yua��M2^�����EJ4�%M�~.�UT�x��C��*��9�=�b�sȏ�1�y�U��+\7R�]E}��{o�p�^(,��S-7��{�%�p�i��-��~���)�bh*�KՐ�S�5:���}��%�R	�ѧdЬ�޻>.��s4G�m}:W]B���S���i�a�:;Oe8Q��\̽��&^*��I��v����籁�j�±cq��J�PdI,kV��<�#��,�V!i\�}msO4i����/A��ٓ%7i������N�����������V/;N�AX���YqԌ`[��������0{�?�x +�	�:<8��U�5��jn�[èkY:�89HS~��J�K&{b�|!-~j�^u�����O����lZƪM�Y*j�ӷ�)uN-��*p�v�r1]ͥ�H�j>�t	�(� {:,�qo�g�Άw9>�[v�n�m�mN�����-�EH�� ���x��X�n�Y
bq��D�?5�^�ˢj�Oر9)�xL���w9�.����d�S�qa�;�y�k��Zq�����?�z�
ٙ{��ڞ6ٗ�<���$1�5�}��	5��鎸���9)�^\/�k���'Ux"����\���u�J�������<="��ݺǩ%�찤RȮz/�m�W�鋦T���j~hn� ��D'�Unk��̶�;��47	BE]���^��1ڸ�v��(�2l"<����A3BH�K��nu*�k(��z��$���?���ݗ�*9v��7���F�^�#zx��/e��GR��i␿�t�h<U�N�Ɍ���M*ѰӰ̄�:�H�&�Ն}�c���=�cr�g)�+,��ɥi+�4ns���ܙY����I�@W舸�YU����V�²�/��G8�c��n�_��(*)X3�|��IzҼ�&��3��-9��~gA�<%�QE5x%1���
�4g��<^��į�0o�C��+�^�A�r6�k|{�����\!�d9:�