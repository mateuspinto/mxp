XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���XH�n<l��ږ�?vVF���x�tlU���Z��sC�����jj]��f� �z'%��2v)&�uk([�$�(��n�!� �)#�J�쪽��fb�[�]� ���p5����k/(`l[�����}�;GU7Q�E������~ws|-��7��檠�`��o�FH�:	LSHm*a�7������B�3��E:('�~@��^t��'IW��}bĝ^�D�;��J0��u��x����6�QH� "!V�S�w9�8��͙��a�<RS��|IFy�Ӭ�>��L�xk�ƴ�`5�N։C�&��(W�y�/i��%��A_TeI	�F�w6'|��3.1[�U��v��>N~��R2��TU���LE��$��X��;��H��������#\��r���^��;H]�"�m���AAl��ð�&�OΆqg�Z�y˜nm�د�-w���l�ϣ���";��nȜ�j�˹��#�o9E֦���%�g�W���`��i$�������8b�(R�۪�������P�1x�7�	$��o^�7�����Y8���TM!U�dj{�n�觌�ċ��K忚����O%8,�&��qHս%l�ZnabL��c��^�,��<я�?@��Ss�F7��r�UU�م�y�&I:��i�eIo��&e��~1�"'o4���Zgt��dI� �5O�Ľ��``���m��ͳ���?af�J�����d��k��-��_c3�� 7�ً�g������A�XlxVHYEB     400     1d0ur�9ULY<�@��1��1d�r���w&�����&��"m�P"�Ih`�@_z7(l��#`��
�}]�dPCy�R��9b0��]#�.�ʓ�G��*��x }v!"���=X8�t���7��i�H\��ͫ�1w՞��Ox�E���m�4�l;�O�q�s���{|z�����1���< �]=oP�=�Ef,�6����T!_�߬cx������7x�>�':�V��:��,��LL�A7������~*>���pc��k�x���/��ᷨ���E��ĢK|�nVFG�|�mx��%lpW�CB��ƅ���Ӯ�"�f9��d��U��º�&������?l(9rߊq�@2Ie�ʎC#����S�! �1q�2KZ�p�$�" Kˤ��>os��1J�*�T_SV��t^b����!�!�)��B�w⵽J=�}��lm�u!=�\{h�5�l�wn�C�XlxVHYEB     400     160M�d*��c��":�_�g���\��!:�'�?C5�ߍ�b)�ԭs�2���R�v1�D�d��\�B��L��QD���7�H�7o�囌p�M�����qɀ���r� B|�V�$�$v.�JE�q�a�Ϣ@��N�{P} 0�I�S^r�e>��$��������9���b�Wf�1�?_2jm{�+��ec!v'�K���o����o6�&{������h&�dx3�uU�((_�T�xZAi�_����K��I�;)�}�ԔHI�����N�
[�x��Mf��i�S��
�"�~.;׿S���ڼ���{���u��N�-�ë,@� ӗ\���;�k��q�`�Y���l�XlxVHYEB     400     110t
V�u5����ul&T�/}V���*d�o����!L���H�
���r4�R�
��&\�I��:�k!�=�I�07;�&_G�]Ub��i�Ș*ֺB�V���#���m��#�N|�'	9yz����'�"u�y�k�A~�Ք%�N��c<�d�@^&PKZ��dX�^�]2/}Pv
^�oa��5Q��}��Cݸ�Tk"���Ji_�k�=��@�/q�3�P!e��,��O�(��a� 	��'����� I]f�;��y�䡀�o���'Cg��u�jXlxVHYEB     400     110���7��=yU.�^y*A�@i
ɤ��(I
Vm}��^m�뾚'�o�z��A>�o��]�q��]�i�
�($
�%�W�J�'��}�<$�%�g1�!��=�<�"8��Z�S�a�*� ���������`�+�r���X���t�VP��_r��������S\������4�ںÝ?�8@�Q��%�hĿ�\��F��kF���r�����
��8�I�#�
(s[��x�ω�`�N�Q����-���Ls�8a(ZޣP̃B:XlxVHYEB     400     150����4��т���e��=W�u��,ӎ_2emël"3��a�{�"( v`�۹ �z�'��M�u	tڰm�`R��u��X<��I��6�_eb�
	N\�'f�@D݉b�C�/:4�3M���%������;P99qT�#=n�����ی�ZѪ����C>��sQ���5��e�F��͌#g�^ܚ�@+Z��K���@�Us�ԉ����7W@V�ga�8-���!o����(����4�4�l�ߪ��P�"Պ��]��G��Sp{��P*�C�*�9:@�G�C�;����!5�⦗!��֝�#`ޔ�l��Bve�s�]���k_XlxVHYEB     400     190��.�-��c׺S�$!!�Ha�ag���I�YmP��8i��i�HuM��Y����������9sl���/ȉ�i#/�f.Ny��n���Q��ͣ��D���"��Fd�	/� $qٜlQ���Q��7_�DWl��M�D]�\/���!��Kj�h��Ve@�5պb�iՅ�z�m��3v2�D�NA�zG %ل�P�V,�]r ����hլ\�������W�	C�y_��rT�r<�D	�P�H/y��0B(�@�iH��Dl�����͹��r.�;i�H��б��O�أ�Tr>���o�>E5����|ZN&<ha6��4�A���K>��p�Y?럴��2C�Mr�p�#�)7���4#ĹX,�ڈ���9XlxVHYEB     400     150k�T"ً��ǆΐ2N�N�X�E�+�r�u���b�Cd�Af�e�7��Р��+�!�� (}A�����D\��!+T�@]��ޛX�g���5	�g[C�o �������\*��:��Cz�:�OB�%H� �̫�	�&������t�V�4��x��@ ���=B�r��C�ypjl��g��^�3����D�e��z����r~�% ���ԫ�.����L�>C�P�E��m4'ϋ��.����d�_�r��sT���u¾'|���S�
R �)W͔jRd�����8�M�� _)�d{:���>�GUW�T�.e�a���sCyp�o� <Or9'�1��XlxVHYEB     400     160��'�MO��"��Ïٳ_y���H��(������Byj�j�Gj]�s��ܷ���ˮy�Ғk�p|f塞=����
������@�z�Ex�Qɖ��ھf�o���������n�#�fY��C��*������Z>�c�Ł�����;ո�n�3S�Z�\C�N�o%t��W�8�#@\I���-���}�h6���)@_RP�i |���7#�`�U�AFZ�A����W�"U�\b!��HԒ��n��3�^�̥�Q���F�d*�N�� &��X�zk{�q�S��c��}��4��D�6�w;}%�R�ɹ���$ts �(���r�,�c����E��.�:���XlxVHYEB     400     120��_Ō6F~K�f�FZ�ۃ��+[ܧ��k�ztpU��7%�3q��p_��Ǧ��9d�+@�i6Ou�xrzi{�%�iJ�A�LxD@�W?f�'���#h�A��#_n:��O������X��%�	�F�l���@�� 0o��]Cʰ��'5n�TW��Ck��,�+��B�ԕ���eB�g��"?°��V*�y2Eפ}�D��\�$�Y�ԈF�}��e���r6q�:�@����J�M�H������d.�l#��a	���-��͠�
�N{�xXlxVHYEB     400     1b0M��.1�E��~�U��J� P�2�T��{1�;wk�Ķ&Ԣ�p��G\vJ"�R�tÈ=����:�2�RQ��:�����H��VCN�r=K|''wDV�����fG�J���{ӯN�[��:��
Ww#L2܀Q�^�5�qTq����I9E��Dp�f�]C�ҡ�
T�N����_��!p%�/u��^ʵ+V}]m���Œ�BL��'�نmw�L�&c!(�z�?.:�䃚�a�7K^�.I�P�|�u'����>�g&�S��$�N��A���s��,i6�����"e�[0���iŻ�t#8Uо��n�]��Fl�����M�i���P�*U9蓏	�iDP�-c@'�L��AӚ�+ա����1��M'\���>�t�ۗ}�L��?�f/x����h�Kcd��g��XlxVHYEB     400     1b0���������K�gn�5���'��Y��;\^� �+��8��54-
ݔB���� �$���v���28dT7�~�Q��A"LJyĺ��x1X�W$��JW�P+�'��R%�`O��;/��V}��"�j��$ƩC��"o5.�h<���;��v@��������|���v�z~܉���U��I �~O�T$���%<�19������5�r(Ho�&~*^,ӄ�˩I^0���*`���YTΕqJc7Mk͜_���E�^�,ܙ�z ��?Y!$��͠F�����G;�F� 3�IO<�?K����85:��'��%fz:����3x��n� |\ԢD��J� ���O��}�+Y�� ̷R��ǥ�h�/lO\`a\��b�]�
#vX,�\�}�vh�d� ��E��>(�-XlxVHYEB     400     180n=�X�Zӆ�KHM�����:O�잳WG(n�C8���TqC�{�:j��&���E�߲|a�L÷{�:��֋0-�7
?�<1�����\���e��tDM[�w���0��/5�`��1��s	h���	�Y
��G���{��חV�'��d5� ��w	��2���\0�W�Ʀ|�� ��F4[�B���âJq��Sۚ��q:�$�.^�*���eZ�8>gf~��I���0��,K�.7<�OP]��G~��C&����km\���q� �!R$\j��*$���+,�ko� �6D �xA�QP=`7�=���ծO<��mX��<FSP�E�S%=K�x̶]U9]PG����i��bqZ��O�l<�T-y�ꯟXlxVHYEB     400     1709r���~�󅜐�b<�V�@F��$Z\ �{ک�������ђ�?��f��jmpI����s���k�pt�	��[(�F_$4�^?����!�����Ж�1=Gh��P�C�t��=��1��^�\�/#o<�@l$J��|g3Sa
k��.����ͅ�o�G$�q}{�J�c;�؍�2�Ř�&��A{Ո����\HҦ�cC��Ɔ�.Y��"��"JyC������d��чo���[9G*C�z���&h�We'���X��=`DƐ�Z���Pa� 8�rL�"��CF@&��+:�/2�w�_Q����[�G��g{���]���j��2W��չ�����8�\PmU�G[���zK�%�h�XlxVHYEB     243     100�Œp�;;�jp&�5L���wY����y#)(�r٫LF�p��/�Ϻ�XTc�|�A����.M��G�m!,��vR�W���0�7Q������y�Џ���5����Ӟ�����=���+K>I�Up��a�;����x�Q:fҷ-�vY/��R?��a�&Xȷ녋r��4�s�QH�xH)0ď��ZāY��4[WD0qW��^@A��hA���4�x����s�����>�I(:�iv7�r�ȳ"�MX