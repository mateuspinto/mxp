`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
eIA1B4CN+clfh/RUFip37oCjXehxNyR7+UwFe4avaWUm85lmCb6T8OCBj+zUd94QoFadXX+QMtb2
2a7KlkxM4I21Nvkaqd7xKvH7GZ+rn+hO4V/bAFvDrlWDuiPcryutgd3hRC75pogIy+b6X1J/SYJf
37aqIzE9FgUk68ECI1YkVEfE8BhLtLgCkj2m5PEFAfu/KC9kyfmWczZYZM84Nk7feqKyMWxkPvoW
wZfWkznLeoUlhauaE0BEa1W6UBLvc9O62Ln2nsjMDiC5Qvgx5S4nSf+U/FqlwbeQ++9ahiQ0CR3o
GYhYFxzk1MX5xSNyii5asezkW44fsip8Zf37Zw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="1wYkgWUy9ePrHYtyb3ZVTN7HAYB/6ZG93sIqcSMJn5Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3600)
`protect data_block
NMNbqw6732kNzqh/UIGq4YzQUHPDDi87A9XsQtzFj7Zvq3HvtaZSy+FkOT0QMlatdd8v5zOXnzft
TYGscemCHCQp4tCBi6JutPgYGtbqrScVFRNXeubcTRYpJgv+cUMmzhov6hHoEqpIK0NvVnrXwRPc
F4VjaCy+TLF71w/BvD5FPq+5/qGZmw9mXUy4SQ9uFUD40H228v8hcy5ZYYqyNhl2M7G21DJuQlSv
GVaZhoHarBRiaqxzarQ6VlcUV3I9CWMZmra+u7bs91DYr5Ch8fVaTYbEpH8voUGKIcjvrEiQh532
hM8J4yiqPbzOnv/WdWdIBi4iLHXVkgSi7c/QY/rc9uPOl+ubQfZuVYqE8E0ZmMQ06szNmjEcQw0Q
QknAWIS8Vu47Zxj3juJOM0NECSuJfajc2rgnIWb+SjV7c90BVgHiq0uDhVDNoS96pHeJ2If1M5LM
0+N/lBE4xf2ZBq7Rs/YlQlIe8tFEF+42b0B89ReVRPWo69pO8N0G5nxNGQGcYl7OokcTKWCtAhJ3
bLhHOiH7gR8awrCotIcVgipQoNvrNifBc9mAfKBg4Nu9c+w8BEA2NyQuMq5FjAyJWkZ9s+hS/o1k
sRiHLDon+NNKK7+UZ+bd/ZBuTHl9LyC1OQilIqD9bnpRx7BusGdkL2+ltPmoYB+q7HZqmHyQ3pWv
Sz29TCw7xSNAzhvvys6Tc2cQJZfLHYCJ/3qDvzaUIaJ9LLl+pxkTiuufYTBrcYgPOCx57Gbs4eN8
kcPVe5X4MRMPQV+9ZPxpEBEYqMeS6l2xMqQmqGd736+kgZN8kT4FdNoeeU99tu+runAZDj7TwW/N
VkWF6QtI/7JYV2XQ2PnUfmaUy6kahfGGKQYBhkcxobpLkYaJ+s2rz1SFvNE6MpcJFM41gQOlyZf5
WTFMRLFgIQz+FMvtD/X5q0uS0HSMmXHWLv2gKT5AsoQ1fwfZaC7UEbSEj0wmAoI1SJ8xh2+9+vRZ
qRuN7N9yIq2J+eUIMZQ1PgkqxutLwA54odHL5l5VbD+mUU88oSfRppe1M7JBR0h/UfH4lEqBzLlj
tRzdp3GXVPWfGeoHKfe16Iv8k+kBWVCdv+QBnia75dAXwFw3eo2tg6FOeBj7quYtfIHqlo421NdZ
g+HaY2Eyn4d1r7XWwUybHwqcw/9xXTknFVbi7SozbBUnapxYK0BkTNKaYA0Ctib7Eiv7PQFBsvyj
7+H+TekQYSLj+IwWA5J1tNsMJumoLc7GxlwowmJBqAVWu3L2uo6K422UCpIk/pg+9bODjjWvMRN0
3jVrn8On/oREbQy/Ty+JlnWwhqAE3YCzySoetfabnJwwUsxH/yxIvqkQQ6R9+IaU3YS7QwJC8749
zbLg/WCElsM1n5h8vLOqCY2dOnueGMnWKHmEcrVuh4mFYty89Vau4bQa4Dt2VNyN8CtIzBrEdjy1
tNtQKmEysmj3CaKtw5PtbvZ224W4ZMzWhMfKTOI49z6pmYumrlLjry8Maxpz6MFg2EDYguo7/XLB
wOo+tqtUDUH8fB+6o4svH7PvqgOPh9W0wBcSwmZ8OC1xYOyBsBW1OFQ5ftMwY4hb5eCa+aNg9Zfq
8ETs1IDPFG7qW/IUOovir04UjfYWfAn3bqSyuLL2rMjH7zjHwZVV7cPrpvn2tIOy1nm+obiIW6du
sHK47UO992INRZNd/2jIntYDztSJsYUzNwyp1oBcoPofFqmMmzCQf2cr6ECdkVMcNTYugnLICKfk
9Hxidwz3gZpRGZ01fM4G+eAJ+fuU/PK+Op+0WGCYnIqXVAd+CERvY10uz8rS/E6PtgG9eZ2k6Pz8
j5XDru/4g9sgJANubVZt8WzsQZ3dur3ysa1zbiqOEg/Eh9hpVKb2s4qeVikQYlWMb8DSSgR+pwfi
QKjGF2LjsD/NPx/9zRYQXSgKm6apZ3mYTZr40kClFFsEkpA7S9DDhlkYvj6A6UUSaTPNK80pbDWJ
oW5J67MbTVSVa+AUt8DedbdB6f5P3uuN6lWxQXpLGl/AIYim4gs5itRLj+3tzg/uVDlno+vUqF0R
Ca+/fdeI9b20cXhBfLSDpjwDRGn03BLsQWp61qFlSdxKFNhziw7V4wWHgvXwk5STI5iK0BFMdRbF
xT+QHs/+AmRRMT/xK/90rRqX7BCuwuPCNgDBJZuYrMtOLQI9kQAMUy4nyjGbZXO4ovAhpQezlJQF
ATg17NTtmmVEZ9KfbKBbrIkSNph5cyPIsr5aoIScabzshqFhH4nIfrBeiOYNWg5B5i6ClXTQAv/I
vF4icbPnC49kWYuSPCndHQAf5G7tEm3aYXqkFWbuhmc4VtCKbk7waVYu6Mvsgipfamc3XkGKxlf0
GAButt0pDg9E0qgmfkR5y3UBd8JHPsidTyF9EP2na/dAov5K03I4QDi+MFPF+RueI4sI4SS0VMg7
nv43IewWkqM5VcVPok6lKUGp2a9h/MWn3S469VF4+VhMjVKgH8piY/wblUwTggIZv8PlrA0rLmo6
cMdOJ5H3/GnFv8GAr7Yg7y293aAXBKlwRyDADy4PB+m9mB2IDVbA1HhWDYcq3Pqbhql+QKzOJMUr
T15dyrCh8YAYRmRCqonH/uO6bbLAqII73B8r3nRdeT8q+r+wd0CJHM5UnRJGYdtAmMMqj0oQWUHC
eNrozIgKf4NGOSK6sYdokE6MjlLyUEmQwK5o9A6TROcaEF+vVKLMf7D3AmxkiCIa6yeRk3eOqeSd
SiOdedUfwjR6j9cn5c5JUdqF/1vldqBxRS8WY4T7zmjIx3d3jmbhtFHfHKbxaes3Ai8ZKXNvN+jO
NB8UAqcLK7q8npbHi67AxAlcqfMa4mvTfOZQe2V/VRujGrnDAsOE5yZHGdWL3useIv7sKMqFX6yH
2BJ4DQOnAYlFfHhqxMvlmtXzqzCNSG2zJZJeTZ7otLzPuyJaa0JpxjNpPSrhzipdPqbDz0E9z/sV
aZlqQE5H77qI5AKGq3W/z2+LZUiF+sQBWAkA9jWd3v7oE9YmdymybRejg3fJMj7z4m/1qCp8EZn9
JH7IdRKN/8mwcxZ6kgNZjBPtfK2zQ2pH44HP1ClRq5ANVz9QSUs2QiGfu2VsLRrMkSzD8kCVQAvU
WkPOvvjm/Ew8B2Tx+8WAdnfrEO+eXQvxnaR4rR5DwWjfItIZpV1i2uGJz9/Z20Zgu2dc+UaTvXRz
6Ahl98Bni4BAG6yEZ5MSY4GTKxOKLPohGemfmqfGIIwMjZK3Ncm+ceyIfHyfIEQLUvkG4wGB7W5X
K2h0VpqrSukzG6s7z+sUzyr/VAimUsFZ15vv4qKZsreR1RuizAF+lTh32v4Fqe3yqGHUX8F+rcTN
9Qbqo0L8P3LTqYjlkMkvcCxGXUNhBgV7WRVMXQtFk2oqxBk2MMb7HtfQQT9ciZOmqoxENLQVLfvK
yn12D1Ng/Wl2JLiJbCl9hkrwwxCoGzyLJvmBcUTHR990lXUqMAb3FtuUn04GKF2DuGooglY83k+j
4lvjh+cFFWjxRtoCIB/Kfdk5c1cwSsyVLKnPCiVBTUljOhrzbYW5Y07hr6xTBFvT3KroikAqPkxV
Fp/T09WwDveEaRB+O1e9NmxG0Lc1UqQxynMrVOTtMrQwD52UwM56GSe1nPcOAHupXIm+Z2jGQJRd
Mpi3PwmbxQWDEysrlAItU0kUYwu8iuE2dbOgAjulL7EgtelaPFt1P6o4ZvM3tmA6EaVqcU+fal+z
NUR0Cz31N5ItULBgHk3osfCKoM5qMMJw3cASNSASf9wlfReD+aDEtUtvlqicbwBiW9JwUsU6UMSq
g71h83LOJV5fv3RgzWp2giqBunTuoNXqv/HpVFsF09TgnWEELZCsECgZ46ux3TiZK8+BdKxk7Rpr
HCQ+Ev2+eAYvbS7bjX7tT0em8cZEXk8n7iL/fBAfP+3l7R8Er4j2cb60domRxeqGr5XKyoO72F0O
hd7IkQNUJsD6FP/+YFWHuicZq1MsrS84t29b8pW1zvUo9GLmtZJUSJktDRWg9Cgbh7L5atySNsH2
mBFfqWGGbag5V/cNCnfQQkJNG4er1Xv4HU8612qeUaKxMkjpoSNcIqRid29vLIHrY57F3doA++0J
K7U9/mLms0idMV6bs/OdLdy+SxUzShtrpefNOXqpd5PKW5CEE2tPuHjHb+TYg4zfXyLgBLsu22tt
H0c0KPiwfIhIDfn/oN/zVLGFAt/gfO+wsg+DpLXkkWkdATu8T5uckuYsizURCI6WqgQ06/zSXp/+
cGG9bs+E5CowjiQnRcDnO7ZIlq8GIgD1ZhAU/2TZ2RHU0oKhJzuoEFAvt+74chhyNZQnzb8Dx4rx
+uaQs6A3VS5miYp2RemC5ry5zLCCmPtFMQ2Nl1gKVsFh4oxurQ/hXg31hcs5bi1QmQ8H88xp/84f
G/beD3RtAbGJrP84w4t/Z8F68+cKNbpX/BWZhz9Sxjubest0r6t7RebZn1DUwwy4m6yjKVdKly1u
jTphrGb2mlEwzRxWmj7wgafUSYg0qgt4P5M0ETfzYbuXzCtotoBtH+WkKZyIOeO2F23AUji1zcuy
V32jhtIPJOELdeAiorlpLXRF155O0pkRHQF4gQyvb/cUDqnDNypuZtgHKLvzkhyPyTVBPRLOyCxD
3ZFskIaMiEnbygy1P57lzlI02QZ788AbS7wAtKrKy0H6ZPMmV6r+PKO37jdDsJTIT9W+6ajYUVSO
+j1cl1a1fSxC7traUEvs6bB7wTxZu35gN/MG0T1qZMASOln2sFb42FbW2OOv8WFgnPV/9MzKoKIV
1Xb4fUCDsO3v
`protect end_protected
