`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
BsaurmIdPbkGAju+2GkaTIplk/0MZqC4NaDfrCQAqovwbBZsxPZ/Js78HCmgI5rkEg7NJ+PWM6XT
5qvCIaC/vQAVu+y0etsDJgv8vikgXRlUd0rFyw49g5XV2ZxYa73i6rVRgjxSfws8k/JfA//8ITwY
TwZ++8a/bislAXajhccLkXHCUlFuOZPJPQpMgu+QS3ABWhavDYu7aIIEiBN/eEFTVxgv9V4NiC8S
hlkvibfnKPqkfNIQGNjpuwWcu4oChY2xDZb7uaUDtC4Rj4Xoc1jYBV74+wpjHbscRe/LAUj28uF0
lXKsmjkBuJfuLAyE+cdEoHP4yO9ut8YW4XHkVQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="MCtjyLyyy1mol279M94auNcfclUBJtJ9prfWk81Vma8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5792)
`protect data_block
/2pytTIazvkJtTZva8fKtV/Pkwp3xaEIJfehYzCg8OHgi1/rq37yXv8botXvKCrAKtYCqSqwr/MW
vk8SxdEYqYcjQ45wO+xzk75qyTbzGkPuLATD+IytKm0ty9s//Aw3gmwc40k87w0roHmrhShAmGQa
Eox1qyeCCOkFckgSYz/GSYXtZ90abKkeazIoU7tj3pzyishZJ4aG+bVxCUQOte67SqbW9qmBLjHn
BhHl7qGvPsH1598+IhbrIxtJOz2EuUw5y266liDWJXfxFX0qAA0WwBQVa4mRlc5BC6NeSifc4SYz
nXWj6mIMcfMVNA4ccmOpQILUgAb2kVjF26OEoN3s0Ue0bf3BDaxrDekAamJTUaYhm6HaHJ8a3a+g
m8uNVJKjGNdJx/fV+MI4xJHvnUulusD3zK5XtPvQ2x22CVw5b4/5dkxQ6tmRaOiw8aEPBQz6jf3c
v7zX/oiNwYAuFLjiZ6uxWCNtncRdpsEgGtp+IWWSWug6+ioT+HDamN1fjHFuSheGCPOV74QVGuWm
RzOl+YziJx1THfJKhJofSYwV71oY7QW3Ub7ADmeheJxJ/QUHLT2iiyQXSN+/XEfMuxMOSwj2q+mQ
RQMdePwAm6dlXMcoayL/kRFFLWXcZSmS0OBRVovn4dVEXY5H4rJDkAtYVfVXNFDB/N2nzs1tbCZS
4UAD/pA5ac3sgtFnOT9+pTrgwCqKjw2//kRExqr/cAuDth2gnWJu7it3oKGTnIL2BY9wmWJl/fRU
MqxVM1cbwIHMsXju0jgEZaFS51Lkf4Hsn9WtyvSCc4fkUgEamsm6tcLdqpTI7ktJ6eBoTwfcrhm7
qiK25NN64fqTG4Y/ysCRV0kfKZP6/rlIkc4+lfqbUHH3D/d2zd5AKxhKfllG3bFUFJHaN225TUWE
TPoSAmuuDaPdNuOOJKI0SCqgS4eHZCx8l7hYm8HdzVi0kGM0WeUilvGbKzw3Kee0zEV3UA9blrY4
QEhAnbYEAaoJWOLai6JHCxSvPpUYcMbjSfrmeVDvp0fvWnQ7bVU1AWOGXJnKRW6Xz6a+THs+Adz7
bbwLkoy0L31guAU156VYiMC0jCaSCNE1zMo6fRoiwSVGHD8WtKw0PHmfCRLmx3+d0msDYqIZeiWd
zuhWvXuLWYBlzh3qUw6edriMMKUpgQY7/H9LFF5vb94WHUbRrx1jY/sIr2Y5qCYOV4bajrp2ozUR
rTnn5KTC1pbjpDSx3VeSyDBeYLSdVXlENZwaLUWBUkhIq8Xuo8AET9nZdz8lHQECsqrl29z1wF5l
FUL+l3ITBDW1ys2WC21kg2C9Zdbf36xlU/ynI2Lz9EEO/59iPPMUeeycGkWUvARkmQt2L4IMuaib
iiAgKlw20oAdNBQBB/DZndhKsUOh0eoo3NZmXlNBcpMDUDCq++jrc7oU2qnYchAjR/zxL+W+lFrQ
6znBxKkOQcXFa+ecb+JVXvYubyMqeSzItwbWxnLl4v6ohjkv9K3uwkA6sVx7prNa2FZT9yBcnPZH
8wjB+2MvOBPpLT+7tUuDEVFaHrsBV9yaS+raS1diXFuLA+K/rVNIfgYZo4OVSFoEm4Zhmv6Ktgoh
5Jwz0sRzCNbNIFsV6LJoroFtJM7geAF6ai+u4iuIW94d6dinq0mxwcXwlcLp3m/ozNJ+GrO7t7t6
bhk5HJehJCQmPxNptTY1oQ84mIzYo/zrKkNyPRF4ngRTl1hGYYA3jlbOb+rxqBPzGSWkzSU7IlbL
AzVUsGa5LgQuwZ23tOaLCvOHH16cYnywMt86DY4iFO5uSab+JesUG+9NjbP1mlLKFzk1rujCowUG
wgg1eyGA1b8+gW1lz49NGgFDXXBnvdbHsGxBZboUC+GelGEsH0FIM2J41wNhDbsC4LBiFPuSlBWZ
BmU1yOkzwKqU70KbEfwHRrzPlCgrqqf1z1ahIYTUubSVE3+lIZqvvvuCga0AExxZyzUHJayfChSh
0ZDkpCde7hdLVPq4pL8UGpjyVksuLIUvRf8N2ZKpx768oVoZA6xM7IHQmgOcvx8RnKsKfJFUu+eq
l8UJV+vt3PmyCUyfmkrGHsk+PkEUutIG/+RignJbx7WtI+Ufhg0BheyLNtyZHjSNne11X1xfFZ2R
+uMrj5R45uDq6kIWtFNc59jlra+NdpmmVMrzmongptCc6A6Xl0Nz9mwU4wwNODOk5tmoBJcs/okf
Jw9355dOOGrTbNHVXBz/XWJegHNkgO9ViNfh/MJbqrz/6sq26ImZLvqyxfryUfbvbfl831OoaDfi
q1/4PG+VLbqd5MoNHwC0SCAvUBpvrKvNBT4tsud/FFyryRXdnZ4q+7WpnrtHPCbiQxx3hUrW6TdL
hqZUbZZx1v4+oAeltU/UnZIWL5XG75mLZvO23ysFbUbvPudPdXOUT49i9+Wp36Pf2JwBNCquXBSE
rgAkH0VA+1UAK9VTU1UImaPh7AaAv/uGgvdtIkpCXSwppICeQ7ltBXSIB1Pa87zM+s7oOmSzAIeG
8ralJrnuqgywJ9rMTCdzMMdUwM+N3amWVInMTOG0xp2mMmbVw71eUzhrEuTwrduIHSgkIpOfGoJp
qmd8G0GVGKkpfkbIT58xg5C8Ggm8dZ/N9XgNCxCIf26K8g6PbAXYKVU4rdjoae5Q65cnPyGdH/xY
wY/KshZIOHvKpg+AjwM3PuizLecSAk1WrDQ+mmzDzb9Fw3G0iqX3q8wjf1srclsbiIPjROVoOIIT
3Zr11RB/ApqMo86TyU8ihvkGKeqPEhot1Q13gXAwZGNzQ6pMd+k8/GBxcwaLuAvtfGyxniXKy8Af
ixr8Hve3gl65cajjEGBaWkWyf2lvPvECt8Hwdxd0Us7bvyz3wq+EHT0to8G4E8iNWhoVDqGo/jzd
awm1sT6upUMoJgPGFJd1x1pMTLGAcVcW7Gj0Z0NsJONIiZ48yT0TV4t/XWMffW4UHBPu7b19zIIa
uNcbLAR9Oj/PVF/2R+8YyPsaPpO8eCjLoarQrqN7Q8b/68dRYoFOPuCQxojBohE+nfGkWO/gJ0f7
kWAJPZ/slCZ7Ec3ZGw3BPt4RPrEB0NUS5o+Ems/ZdyqzXacp0nrPwMU62757pHZphn8srG4rkS+s
YR+MItJB3akVBzxUiU4ZdGqeSDK75WVWJponORenw1HjzpJqjzGx0MWxrzB3AIWMfYbai3dMf/Fa
O/+iwmj0pAhYPCVCFtiTQUKa1/H6QiT+t616b3YK0scOVABjEaDICW/m9431g9s2vezFVi6gv0P9
2C0jztfTOqm1pO0MD4Ud7u0AAy7m/tM1++Oo9j0x3v5ncbeOFJGhU782d/+SsgWNq60CtoUsK2W4
XA+Gntusd3+4O4vnl/1kzqH6QSA+Xr2VojAHc0HG7dYi2czO/e6E8oauMUK625Srt74HomONZtEd
LVpW2S1uHnIOdIDJLqwyUqlDPpcO9/IiKwHWz0aiQ3NS7ZnW/Pb7ZHxx3JBjt5uQ7geZJKh+AK96
gpLriWqoJwaUzGCNzcIsxeFxjwFbCdAJH2DSbnjT/F8IDBI/HGUjcLvJat1VuJQSEJcX+JylKrsS
nSnEVa3KdTCby5PkfvAnm+ST/YqRr6SRiWOEoy0tBMwoD+wzoknEQV1TofA8zCZP2x+oi7hiCXvc
MlK1sBKelV3QE8J3c8uBJsVu5iZLj61idhxndoOOA/JLmTu7DcRC/b/sDY5D9muvFQjZq2nRfbwQ
H9ujbZuF+8ww2CT//rh2bXgNAxXqJtDRgQmsmCXuej6i1x6/eyet27l5DsBMN/Gysv1IMBnWEpbB
cnbmw22CZOp8GHDtIGTYM9vfc6a9Zkm5zzcjNT0fT3CcslYX09NhFb8VEQ0HQ20Cuz81ihHWZ9Rh
zw54xa49uObiHv/5UosPfwYhPU5BXmsbZTGYPsYUCwYWOsuDhDpcLayN/u+XfT0A5O5Eout8F74h
5V2b40zokd32sRUXyUuvpnXfI+EfzqH97dHZhOkyUvOOMH2tbbKIGllgy53oqM3Py0c5ByekG7eZ
QfYVxZqaxk8QsqSjbc1C3w+SX3YiG2qrQmo6k6q0aPfJDpOuvLpGmrT0RDB9K35dd5phBLLJbAsd
MBdw6uy/wtsN+YcIJooFr5JWtPGKaCPLV4cRvBovYO9vq80GzlokVNJAWH32B+JI214X5Js5gPEr
jCS1XlEcGv1olBAkQHSu8iSjl92avMHY0Q47VUElk6jh/6IXpI5SY8aoay8WNStlJ6iQ72rBc78Y
KE2KQ5D0RAK3ahxXPUUfgwe8oVwrXpj/CigjElxXQa5oTug1As8DswxgmS7CMAZXC637k9AJAs1K
URES4H9UgeFAGJ3csTowBQbPqjrwEI07QNV3EzXQ5FxlUzHcT3MJMKfnc4nYc2nwbTsLZbHxnUqe
pJTZOst2JZuUQ3dZj1rQvU0GPW41T9UBQZH98u9YeX4TPbRzgLB6eqbNyAG7Rvq9zXpD7duz460s
T3D5PX7oVrP6inJ0F6R5cZhlPtonviOEM6Fb0juf60Nl+QGYWQgi2PHoa0F8tO7VS70a+GC3ERdW
lw8YX5FVQruRYcDS1ZjzXsM1S/T5pmZIHA+ouVc39e1L59ESt7nTjCNsiKFRUzmVtsehfLp5gBg4
u/NISbLQQZQFw+wOoqo7tUpKad00xlKOMY/Ck+/ENpI0laXYaCiyut/d/al8zug3CXY3f/41c4eq
Z5FVBEnoh6Nsd7/whe7kewG+INgkzHdwZyP3z3O6TNmLfiG9wOSZfR8cc/75gVkGd0TzG3fczWkg
L1unaGsFGM0FCEqb6WcXCO0nD9ZI7n6DwS/zZvW/Bu6EMVPQtqRItVPaBgF32aPCEvi6yr1TUTkx
0zLZlupHfH5QCOBBMkDb5/Ei1hDFmS5cN0mmQXZPyQvATlbKdnPiDmKLB4m1UJ8Ew0n5LeiTIoaH
5tEV6ft/R+Aa1bpMjxjm7/W4B16gjPsvxl0/Rz3vJqnjnVMfx7rD7MDghOYrKS1CAx4JmuOedYDg
ijVf+G8G+Mcxku7Rcw9rY9AfljLTuL6etTRsJw+TQk63YW8NPLauG2HGTnjAo/I1YdVp/NCeyBgF
qvZAHxCygEiz6HMkNN3Ja7XpdMBIKs+Xgzn4tOzWZHY7L9gh2PVKb5WWVs0gLRVNTS1WDZxyQ4SM
CFT7/PNVOIfP3FAixyMwOGKVmBcWwIhwW9EjSwhvU/Q9jxFFcyyp/WZTgm3/0AOc6ZXPuHiTbdcT
pgbgJB1MEQ54OLnvVOBPQFk8waAKTzo22yifQlzEw/XfAyJ77ky2oXHgrTOrld1L6vFg/aeHj3Z3
4PqDiwlMsDPwcmDjUxXxU1UrDP5MV+1TKz1VVl9C4JfPN/e4CDuVyYL08iH4tfrlD44SbBK2Tkdm
9gmpHFqPZbXQBtIZdyAVfO8fHHYMYcXvIiFb/MpnLHJ0zPjXfL+H1iWxV8hTAqrb/2od6R/KzfDQ
3/G3JzNbhSflLTbGdajuQHYyP3Evv7FxA186yqwp0S1sqvoWhWjehxCwnRZQGwFxbzS/eODAOSJT
ehXkAaRqYhVQfo+SuLGtviNZx+eZxBf/VYQ8uVRcQ+pxzIJharWlFKAex9OxK4wCjqqjtoShTI4i
opIlGVXtSaEVCZmRkEOVkTm96qfCks1vkrR5IvTtpmkGvilI85Y2NVZUhE9if1oriRI8QW5JVqoY
wSXGh+Ey/zcrGNRhPytCLbZFTJ4yeRZI3ug5H2rrd/xl8oRNbs9Bqh7icJvlcrJaPBFquGMb6jAJ
7gr0TLS8NbXkMo7LY6FmM0ngsKmrOTDTR+aff47vf1DFiLsv5fw4Z3Bv4bDW2+6fy2TIr+bAmwjV
S6v43jrUMgc6eQn9sZExzEdA55PCOhp/7yxAjGeKxkP3WTs/+MWr6Q0hiwIDp9BwpUq/gR7TU6yZ
7v8evPGsnrFJ9VISuZ70K9JppNRqhQWlhXWMnWtzNlNTwJg5M5jAhQ8IzI8p0YlEjGSHpw6fLUGH
vIK1RXyc3MNdmZKxI++sr1gjOewPQZK/onP9uWg+Bt0ywPZ1LOmXK/md2QAWAKdLfdAfP9+cVktw
FdiRrzQ6204IWwdTJ2WENpKACbkh/iz4KUnB4JdOwlCo5sfqf4tCkDv6d9+5ekuxqWwSbXlHTqTO
F0zY/SQcIWVtgyPbmgrkKeEdjkv2w5G5sNiKfvFnerfH3Z4obxajcFZcFNowv5pqODXoGIxAHfMD
ivxGDE/3egkSWu6L+gbcVj7oy3FJoS8DOYYQUiqE7b1XJu/ETSyVwPpcJR1X0vOaFwGzOAYejhD2
oX47JgMww99zkzgsdc9FOoK086Z4VagegxONGRDa7brxRI+itfMdgD8F54I6fA3eb+3Uklli29ZG
92F1Nvn2T/J+LBafmtDCWsetNo97tnAH+iqQSl1qevMnQHcgw1D9csB3xmwhdrxl2OmJEvZECwZG
ndY/7UOChgbdrt7NGURt84VQyzTxx8T7AIFhDlGVzVamZITkLWxcyFDhsR5eYfI9PClXDQ+pQFuR
FeV1U1Fn101kU3TTDh2e5I0hODoUxjOrWnCwTYg8cPHVtx/XrXIYtGx+G5L1hPEJXuST3acfKdV6
GBcYwoCJTyuo5ez3cb1LIfM86Q6xUCv7+G58COsJ4OfbaM0vZhpNU5JSCLyh8qxLVZttL21AWGMe
B2IsqK2H1h7HotR70StwiAzh4Vbl+gC3we8IzJP16jq24UUhlNwPSFd95HlLytNr212LF+skDVTC
n2PugO0O5fwDDq7cntNRBHSLykVzZSFPs9TVLYuJmULpnSmrA0FNSwY9VTUz0HGgzpD9jPJmu0Ej
fkMJtEhayfSE9FAeCrJGOIgceMi7arfXnCxS+PI8tpvVvUPaLo6ls69B2PwQ4BtY3Fi/KJC2hqKn
p+noYkTRdRCH7OKWurtevgk5Xj+FcLsjIjv/hGjzOJuEJWGnYk17Qmu1twygTBmgXKPZ30oRFm0M
ZuELxm0rMVUz0z1KGU3hic4+2Qzoo2kCuwFyjtfavwAQHtfYl4XIRjkmJxlPN8G5OQ5q95dsXKTV
psgqtjiXTuvJgr2EsZ+a99+NcXgnDws5wKNJ0KVSPfP3u0osomZvsHSFvKBCUeDLT+aXyDVpXRwE
luJr1wfmi4HkNVp9m0kqGyTjDsrYW+0aSxlbWfIzUuQ3sVOtr4yOmJyzayQg6nIQRfBxu0zIdXzW
H3mLnhoWXPEVTTW7+zU0saaR5FnMbXmPbZ+myLV73UV02Q4d3Zn2is1NuAgagigyODv1vQ7nyaHJ
4t/T6quRuM76Pg8llKU1gRSSSSn/Hxg0MvZQnHW552DpIVEN6oA56V406Cx1ppb4cm+d3KFo0eTt
QfFkhQ3af+AzEWZqDA+Nq5vzdvuJ7EQRI1OJRyim2dNvbm6E+8YKlVTL0kTK1ixU3PS+QrfOWByx
DFSsPshSuwXxV9ory06Gclh50KHR0CQHgVJi7ra2rgxsRXFkP6dzJTET4IGLJoMndCtmeSJYQiLl
gHbZjTVl27U74piRybitV97kvnzgm53PBTtSk634Rc896Gw+0wkWpk6s8apFXJ9j+0ERJhHkhuY3
oNGwnGox3W4A5AEoVWGtfTimGbJ8yKm73AhbmhiNVnVQlVlaqiRglXz3vYN/J1m5t1z3PIaoQ+Sv
Nhrx8GB8iE0hl7Ii9ObqfPEk2/jxH/FGcajKrsecO+nzbnQ=
`protect end_protected
