XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�Qw� ��:�&N�~��NLQ>1�4 ��+r#'��\�!l�mT��\�cIAj7�'�9Ͽ�}k<�,���Vj�^2~��}�!z��4���$�XRC��YI��1ו���8� ~�TaM	�4���SPC,O������t���V����H�9�7�
��V6��w>�ٶ��{�.�M*���1����cw���r�@UB�tܭa� ��Mf^��[�u�)1�q&޾�	!<��
���2�L� GY�~�� z�\���z� ���w�f�QBާ�X2� �+L1�K8��/��]5�����m�D�,L{Ϗf:ȀKKx���z�{��r�Ad�|k	 y�NO�v���{ݥ|/FB����]VC��Db��]A�5���L���:�UI��T��ޛ_w��H�O���t����o;�*K�,7�4?\�B`��$��������+ў6^ڥNWK�{��3���?$`vW�#��Q�R���=�D�E�����L�{A�GI[\��L�����^�=����!|YY��f����%�P��(�`�d�@�4s��4������t��P�JX���L��ó����!��~rh+S��;��cܩ��u#���3b})�*͢�wҙ�]�}>�FP&���q$�`��l�s�/�bn����o��u�ѷ׌1L]�lp��f���$ߘW�(��>(b���4N�I[f��,Ui��
��xR�>Ļ���F�0�J^���W8�P]���M��0@|�����m�XlxVHYEB     400     1e0��Y�3��@�HU��(�D���I:�6_`'�7��3!��ֺA ��'�#IN�#�N!Trn{F�3�N�Iw�{��Վ�_��k�\;]�қ��Ψ6ˋ��Cn�PCqCM��]V9"�/yT����t�f^A��}v��TP�*�J"�(Aw���y m�g�����!\k�_1_O�'�v� JD_����X���U�(��7�Wl�<��iwZ�ᮩ$��x�5�U�����������k�G�\��)P�bdXVs�@������jU)�ӪyJ�5Е��e��N�PZ$S^�0δ)t�oAJ$�+��g&t4dNR	�X������
���d%F�efn6�M����hs��x��X�`�HH���e]��lg�a�BƮ>�U����iB֠���,�������}tnф�B���A�g-g��P�x�0)��7 �H�"`w"Ӏ����O���:h�D�(\|'�_j�H]�t����n<	XlxVHYEB     400     1f0]�;�j����Mⷅ�XG���+�c@��{E!Y�w�̌i�6�a��CNL��dg�����8�Q��̂���� '��~1�.��r�f�[�5���-ga�`����_7{��S�bQ�%��� }�d!-��	��9a�A���Jo���{y`|��)H�t����n	Y4R"��޷�猾�Hr�t���1� �ΰ �0�r�������+X��g>�Wv�B�֤�W|� *.�V������DtoY�XS�LNa���b�k�b�Gf�g|�����F<s�4��]p�?	�n��"P�%˺����o�aa,�B�4"w��I��M��B���*_���f����j/Y�q?U���[K���*u
v����U�%3�K9в�~�
�z�O�5����,��`G�M���jn+��f`蜑�NنQ��h�w�t��dѢul�H��+��Mp\~���IA+��/�HOc����f���XlxVHYEB     400     1c0��!,�*�w4f�^T��xg�<ש�����D�r��K�M�M�6g��A0��.-öu�,Id�G㍷I�/�b��8��g7�)�\��4U_���aR�*��fH/���� eG������p��c�Gּ�']��B0�ō��x=R�bF���gY���Keڢ�M��K¹�n�G����nMܾ~*�<����p�O����F�t�H���#1�Ihr-qF�L[<L��~6;�H;�>Y��� S|�z^� ��]�x�䝑B�����͉2M|-Ӂ��9+q�i�/j�T� �q���0�+��]�'��$HUm3R	%�š�|�!�b��k��~	(Ͼ��"��y	�H�O{j�r�� �P:��'�%���x�(���b��V)v����o\���&��c�����ǁ~��I#@iB��XlxVHYEB     400     1d0�M@L�P�����ưA{ѧN�|i�귻p�L�=����/����Z�X�E��I�SJ��Z�{���ڮ1� �h�)�]y�!�G�Ow��� ���.�7�;�Fi?�`]F��Ի�@Y�H�j���SB�~�|���!R�����n��H�5/�姶�� nm��l*O4����8��&�CQa�
��n$�Bj�PW������L+�a�J�Sn��p�����a�U�����?�Ĝ�1}���$H�J[���E|��.���,%q��6�A�č��8v�K�~9��C�J	���@��~r�Ņ��އ�ai��a�$���α��Z����p����;��S&h��mt�%���l��Gn�i���e{�E�wh��ïwb�%�~X��?��}�F��@�i�8�iؙ��&���M�D�]kH$��P�s$�@=J	ا����8���̴�B
�ە�ʥ��fXlxVHYEB     400     200��O^^rg@���CX@a⳯8���DC[m��j���<QƦ���~RhB�s�k�Wu����5#��c�Y;d��y��	�u(� ��Γ�[��3�6�D�+���¹R� �O��3���_���d'?*�ɥ\PME�V�t���?���������ks���2���o'�J\�Ur�G=�r���:�v��M�°.����{)ƹ��*)z������ᚷ��s��?w$�9��S�d���yp�2�\1��I��b�G�Ɨ��۾��?��`D�B[��m��#��X@79ӱA�q�"�wv1')'�ǽ;�&��I� ��)�d:0�(�ʤ�m�_S����d���I�L����7M�|ʲ�mU���g�&��$t���PNuﭹ��%��Q��&�5=�9��� g��U���S}��&-*�Q�,*|�2���w2^�����w)�/v)�w�L8��.m���*��m�t���O��O���=]�Q���3������瀊:�XlxVHYEB     400     150�ik���U��.�4�.�`����x�l�T�O����+�w��Y�W��Ҍ�jb�6��U)��n+�[e�T�f�͹�������e<3߁�i^�Z��n�D��@���~ސ�\�3�TL����β=]j)���5ǹbl����Q|�Br��G��p��p�;�zu/>�@Me��_�>��t>�	i��(��By�x�M�'z(��'lSM�J�Z�-`�z�#L��!#��F������������4sy:�L��.Q90g�]��Dע���D�S����<��8�!@��a��-I)���^��i�� �^nuƪ5)}���������C��sXlxVHYEB     400     170@��X�q=ZM��˻x�y?��򩬯�B���{�}��Ս]��	4I�a��o�H�ʈ;5ֆ
wX��:�1�E�bq3�C~f�CO;!|��}���r�!/���G�s_S�}B�n�GV��X���Ɩ,��<yˇ�4T0�YB��q�1�0��2[Oml�(0i� eKl>���I�Қ�
�"�1!�|{��@S��
va/�,�L��ҬQ���~�ӄG<R���f�ߋ�\v�#X�o�C��av�RPyj���� ����yL�.�8�Z�s?��U�i�J8а�)�[��]���ˡ�o�6'�"^�d�/?�e���w ��Yb���7	�n ���(���	�\�!��+���xC�h|�EXlxVHYEB     400     1d0�)������E�g���eh��uQ�줩g�ֶ�z���:���Ik�)�A>7����tZ�o��0�̮R�O)�v�h����6K*��bKp�2��.�T������w᪮d����l�,j���(�����Ow�I+��[�r��Ph��F�.y0�Ŋ�y�<�l�G�0n�;YvZ��}����7�G0��LV@�+N�f⓾
��x�T��hNsC��h����E��V����Yq<v�H<t����w �����٣�Y��� ŲR5����xDT�S���`N�dSq�9�j�{�}�q��+��U���X�K9z4��mL���CO���������/�h�x�_ί���}=��).*b��ھ�
��\'�#0++����>;V<�J5���l���b"asXG��^ң�`>�o����.��1-=�R�I4�#Wɏ�[Z��	/����	XlxVHYEB     400     190<��3��Qa0���R�$C?�x��B�}Z�ҡ�*�z���}��:-%�YA���*�iL�p�vj��U=z����ᵩ^�#l���V�&*�����|��/QQ=��UP�N"E��Wmfy�[���kl���Eݿ��#}V)R!Wuzw2�\ȧ�#�nJ��$^���uϑK�Y����܅�W���e��I7�4=�+]d(��Wdu2�b�.چLeXskO��t\&�jv���D&�f��|��H���ۮ$T���Ҍ�̼����u1t
�J��?�����j	�J�9�͆��~n,xl�����7r��%���As�J�ו�}��L��v���T��$��'gCG]�l
H�$۱����uC�k&�>�㎌ﱈXlxVHYEB     400     190����r7O�x\��Þ�P�'�[���PE����u�>" I?`�(6��"����;��"���8��]�Ӈ�:A�t[��"G�y��|�1�d4-6�s�{��9�5D�)��Y�(�ĭV�JtK��C��[�/̚��m0l���D�q�����d@%�mO21�eJvUn
GYt	�M�Sn��3�x��W'�<�n�a=���ak
�;�xqDM�)O�(;�^�)��ZCK���L���Z����"�
�^�r+���!jHX��>)	��$�����N�A��As)�=p+�����q&Y򳀥�Z���"�K-K��I|�7�Ю">�c�L_�{]��]��ט�U��hܩ*�{K=rzɋ��NԼj~<]��&�Ú06w�1�7\J�*�<=�1C�%�0XlxVHYEB     400     150��t���,��P�Y�Y�]΢��,nr����]���s<�'��b.��X�ɥZst�&�yuA���~7�'�����c�V�'�m��L�Q�BK��Ƶg�Hvw�C����m3O>�x9���J}m���־�,]B}���� O��Q��e>ѯ����7Z�Ni�w�"#��l�c��q�َ���:#���qY���B�,��a[a��1�g�M���#��kS���B쒮
��D�n��S)F=OL��/i�Ί�~΂�k��1�+�!cS��D��Ƃׄ���Q�]~}��cH�E�>��\���x���F��d�@��t�8
�_�Q�XlxVHYEB     400     150�g���\w���Y:b�oǤKn!1ȒK7�-��.�;�>Ow�~Ɓ&*�����&��xFo�A�8�'�� �	w�'��,��k�Ui����\�ea��w	W��ܬ��[cr?I��E��z�Z��W�tj�,�����W����*�����<[��g�G��F��5xXwD@
H�C{���ޘ:n�m�l��܇���Ozcf}�4܏Z���	N+�aO��' �^+�:�|\�@J��͖�eә��8��D�O����⅞?��l	2��Q�넘�X�qmO�gHDl��^3[�q��M�t�zQd��IB���V'A�&�z���"=XlxVHYEB     400     1c0�m��@c�*��6#��.�P#��դK������Z��)XjUYt��s��dz���F,��iOv����Y�"5aTlc���]�0�n���ȑ�G �
�0|3¡�^?�X+mgط)C�ڑ$�{?�4�2^
���o�n4HPC���Z����J�e����Ytǉ�n�x9�On̙��������V��t24��_?�MU�8���j0���tl�	��#�k��9|�X��&	�F-n�3����}��R�;��o����*O�ɑ��_�UqX�#7q(T�ྻ��F�Ł����V6�AGK����a4�"����ˁU��b���]�[��*�������]���Sb���U����4��}�7y�X���J-�m1�*F�r��(��n�!=H[�<�v�ͪ�L�G���ݙco���B$z�s��qp m�U��XlxVHYEB     400     1c0��?6I��j�q�B6eH�S�G��^ŔLFdx�LD��Dcg��̡u+��G�[���Z엞MTT�rM�ڞ�a���`���)N�ȈG��	�h�>�X�v!�@L�=]�r���ư*�*31�@ f��(yg�KN�콊N��ì\�`NR����b;�e���r�J828QG�^���G
��_&r���B��J;�kZ�ZÐ�jz钕��\c�F�^��<Dx�DM�Wk�e����:�|%��:/�� ��GIK5��h��!�횲��Tϖ���
��i�d0�'7�X�^��ǰ��"�aR �Z�W���;��hV��K��y� ���|Pp���;���w�0�� �'�!#C�	���]��*�c\E��<�~���_)Ks ;~��n�V_!�\�#�W%��h/$`>��8�=�NxQ+Z���AXlxVHYEB     400     170����,�݃�-=ږ��zh�����דB����+�\���NY���A�97���j^��Wf	nY
Y�K1��*�C�����>�5:Ƽ#٬-Ņ�w!Z�����)�z�����i���K��:�#8okrއ<8ݗk9�ٖ��m���RW�v�M���7�oIp�.C�Sȃ��bѰ���<[��A�O0����弖�3U�<��F$A���+b{<���y_��E���0���y'����e��ڬM�.���+�I줉��Rv��uU㫬!T���I1�����&o�1��n�Ӈ�Uǧ�&�mt�E� 5��M���K{���@��<,(��-N���g�Dsvt���&�Ce�XlxVHYEB     400     200�iԱ� �y ����*�P#L�<f=���Bi�� ����ke�_;�[�|Җ]�v ip�^��S�d�$xcB��DXIT�Vm�x��w�&yV��k�#�uvo��k�[��͡��c����Y��ǘ��'B}c��&��{֛G���A�D��透>}C]�j��Q�K�F-��^U�\WK�zG#��i�Gc����= ߫!���Xv`+�^5��j�Tj\f�S�?��@,��|�f·g���f��%q�sѫ�b���Y�,"��W�Z\��Ȗs���Q�B�qm�3� Tw����_���d����I����~�_q��Ƞ5]<����cfR߹��Sj�'L��%�?4�Ն��ߺK�{�˵>ۘ��i!�;��<ܷV����:��T���JY�9�9"`ng�7K�GJ	�ا�C����?]4;M=xh��6����h���Hx
ǖǚj�]����V��7�X5��:�l�Ϛu.�:zh������ڲ�MVO�j!��7�J�8��uHXlxVHYEB     400     210ܡ��{�����G��%%aP�ZoS��\�tf��K�SB��Ml�A;,�1�4���GCڤъ�j�!�E��?`jc:��U��Pv�mjo�jxoȢ�5�֍ա�T��^�y�.U��*�6��U��~[���&�ON�R�1�����W��^*�ʪ��) &�:m-V S�����G��;�qϠzQ�	�)XOȏ��*l�e}l�"S�8�+櫶��ځ$��`;��^���1c t��Ux�"�j7�Mԙ�_�g�6����Y���$c��=��@io԰� %�	@L����S��頙�j���6RW�Ubx��V��v?:�]I�f�C	���|zo�6�c9��W��h|h���9
.k:X���(��z1�X�n�E��W�P��X)���Ȋ7y�<4�rD�����>��L��c*���������u�>���@m�� �$H��h�vl'�Efe�AU�ݎ�w2�!�'l��F�n����6��*����&��������N|�ED��oSt=XlxVHYEB     400     1c0�eȚ3 [��^צ�`X{��ih�'v�g�E�Ϲ*�Ԙ����b�V��h�e�~jE�ǈՃ��#B?C��MjD9�.�$�YdLE$ݖ 
���k7EX���:
�'�'g�?�A���%��k�n����[�4�� =@$�k绂���(��/���֛p�"�� 6m'��3�	\T۳i��f��TJ����5#鼻uBO���x4�.�8Ǻ̋w����)���Ŝ�R�<9/g���������V������}�Эo�X#�;���Y�]��T9�WypJ��-B�OW�X�V�z��U�Xrxs�y��,�c�(���׬8M��A����q��͇�|��[�_՚Q��2�qpf�P�" ��>iKޜ���Y�_��gK�%����	m2�[��i�3�gy�ʂc	���1�a��}�I�	�B�%��˷xi�R�XlxVHYEB     400     160�ЕtF��{v� ���(巀��g ��U�G1�D�,5^���{!��W�⸁�������[�-�$j��C�MFUY��y�U��jF �*PM�I�Ȭ�
���{�!��<��^Y3%�Ĥ,�����<��Z��Ǵ�)�G�//10��H���gC�L���M5o�aw`K0�I'����~�U>]�cү�{�4Ǡ��ݩlu�##O�ڍ�3~Q܉���r���d2G8����4��(��]�?�R"�wڥ��]|�+o{"�5_6�\����p6�xx9 p�S�(|[d�
y}9��d%Uw��x�0,�p��c��MIi��yg�/(�����XlxVHYEB     400     120��@�?Ոǳ��Ac�l�6�/F>�� �(����t%���L�
qFפ���x���H��Y�s!ɢD���UUn��A��xL�/������NZ�킲��G~��3��v� ���o?Z�ύF������$	5�_��ƍ���C�S'�aj�ݬ��g�qdT�W�2�d@���� �����D>��Q�� y4t�+s�X~p���wV�!|X�B��1|�I�V�� �n�\X~��M9����I�{w��TI��q^��b6 �/����_��ۉT<�XlxVHYEB     400     160�e׌%�Q�M��q�>�p�*�k8���j%�-�ux�ɀ ��c�!�����.Q���!�&��
�B督���"7G�עqK�I��T��VӃ�k���y?�+�Z�x@.GY��*q��>O��8\�<��x�oܺ�f��+ye��ߋ�c
G�Y]nl�|��;�U���l��H���`5������e�6�9���<�����VPBu���u�F�͙��d3���)tƪ׶��Q��y6���6f��)~�Z����	�N�	�"�èL�~�Az�}�AX�w�Q�ms���ҵ�tʨLQWJ�zn��"ba��r`��`x������f�ں�#���(p���XlxVHYEB     400     160x������.�{�Fo;�n��zpMB�d�3z"0�.gY�D9��Xx�%�L�x�G�W<� ���Y��R��ًjG�Dj9�kv[�M���A~�� ���+�:�L
�`Oi���s�t:�����U&�L���v�ǅ��~�Q�oc$�Vq�pưAa�e'*��T���&dyM�'�
��/���3ݵ�|B�)A�֜1&V&(�g?�]�S�)մ����̜^ŠN��X
E�))�	�*| �^#�������d>��[^(�j��Se�[z/��u=صL��7�֓-+9�.����PAh���Dht�9��FC�?`w�Xۏ�ڮ{�{8��(��t�@�Y˚F��XlxVHYEB     400     200��yek��ݤ��-h�+1Y��a�_f�`�_H���H �/�Й1ahyr0y�5���w�>^�
M�C�Yp�"@܆/����
���nȴ�g5�_����LMP���,D���^3���G"1�������\�u� e��4�Y|����`�Xw�B@�P]����\���}rޤ��*����w]K�Gח��ԃ�%\�����]�/Q^�
K&�m#W�"��aru��8($\�&�O�N�٪'��&��8ݼ6�~[Q�I��H�נ�%�M�4��p�%�$h!�*��{+�x�i��St��nu��Bd."��9�t�)���_��ͨ�Q����u�B�u��\<�j
l\�mT��|����EX����¾sR�Ո���&���".p0���	��zBy�@<����qV"o��ťf@��Jz��l���;t����U#o*�r�jw�L����zDf����c'�7��JT�V1FH;+
{~(S'�z`��2�J}���WOG�� �L�XlxVHYEB     400     1d0�ʜ͝0�[��ņ�9m���� ��d+��x�.~���'j��}($�x�fڇO��KAd'O�*�T}�B��x�0� �	��6"*}2&͞�]�:�	���<P�����yP��eH%N��J �sZ�?&xH����l#@]��;�C�:��4Ld�W�N8���k�%��K˙���	{%����,����Z�ćo�T��F_�R��+>߯�� �;`3kN�����L�,W0z��U���@zYG���E]�4�s��{���-��͞(˯%]�i���@9v�-Lt�0U�ޏx��|�U�{����X]��(V��0T�q�9�
}+R�����d)��6��˔Τ�B^�κ,�Qj���b1Y�l�~��(��=�T=�@�Σ���
Z�*��d3�J?�����6�Y�tr+ܾU�������X�� M��Ѭ[[K*��~��N�v5s}�XlxVHYEB     400     1c0�ͭ�'�:>��2�7�io6����BMэ����������@D$������J�T����[��8��V�!ұi��P< ��U����;�X�,�yՔ�!ae�@V�=�[C��PO�?��ܭ:��t��;پtl8�ĐHS� u����D�^=�����6%�V��7>�!�$�G0��HV���-"��ơty�w!�M�G��U�?��p9��*�%E[T��VFk��G����.��&c�'�s��Ӥ7�(�������e�$z#?�����xQS�m�bY0���6�.pH`J_���0�1@{,�ms��x��_�t�E_��4R�w��s�O'�X?*�]c��4�A�p��
ނ���������)\N\>��	+H0�����_�Au	��n����Dw��W�CVw��9pvg���/�k�5?T�,����H����.XlxVHYEB      42      50���דM�}����o�D��ĝT꺂 �~�RB/��o��P?�F���u�*�L��\�r����F�� �ȯXǃ�+d��