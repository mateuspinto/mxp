`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9456)
`protect data_block
0USWSUGxovGsyBJteYpEodNjdpmsWVpNStONQj5zxQQt3qEj5HKpzimTfYj1ybcKQp7BEilkv7UX
Lq1S1TrAgUZsPG700ABVV/uSGne+BZtEqctw/oPlcKCitvt56eP0RwMn2GgTo2RmjUHpoTUDdzO7
uMu6CXW3vlonxzeTFIdAZvdvU7QyTZfwhZMdP3MROjQ5ZVbWUD+X5OucuFuZr0EkPCsbTnoQnGct
9fzNtJKHq228uqLH3258bks5dyoLtx+rt31nRvEvKRC4ParrYJNP2u2cP0b0hk06HIdfbDEVkr9G
/sNAedcUImcsXctjgeomOFjTXOkCLS6In0FX2GCUelbzh7sBfokqe9rxRVt71SpVbWQAvKg8H2Us
eM9n79q+dg2mnAI0lH8HSvELxmyJHY8IgYNvMO8tLMHs3Uz0CDPuHu3j0vHVqGmiPYEwqxku8zQP
o0hUokfh9YpgX8x+lUQdSTrkQNCRYcwin7AoS8kCI0ejqlAyM4meDq/QI7grLjAN6+z3vcH8o3vR
QGjbEsNGNf8XpsefnR3oniF5i1OLUSsVm9xKiivbxb4eQ0nOwcrFdzbKRzprw/8mxk0lhnpVDP2k
9OAkUPZLgUt1cP4UBoPkfob6sv5ftFCgpLuHZtCA9DzNWH24Ksao0Bn6lcuywbVRgemRzecdu0UF
lPHS2y/mEPO/XtFmrIppZT877OlEGI5djjn+8+Qz+FKTpOxKezDh/aO8/3voyzfnyWdSkGR1N4md
rHDFg2P/UGewi0oPQ5HPCjv6BsJPHt2DiCGctSYXi4OJooaFBYvAQB7rafsooDo0Fw1Ub+kgMn4X
6RSdodsV6WWQ9QTpDLzx7Y/xp79Ae01SM+HOme/8t15P/ddYyf/lTISH0DDsSLSmLdyzwrSNr9K8
MjkIO/B9SItBQD2lPKfi/D0R+Ykkdlz+OmmA7wve68L21UxqSO0K8fk2lFyjFl6Hv6mplXH+kzJZ
WkdamTliO+zzfvdzKKiRu7kOtnmUeovGnkU//7/GY05S3JHRSKEFMcWb1ZWhVwAjKp15LEOluG3V
NJ0SUNrtC/Cc4u7O10vjTbc9EFC8hwJ5ANueN+cHQwQvxRqcgeSNl9CO6VGlckJsmQsczLgjHlFo
N3Q6ReTxbOGHy/H52VxbqON9gj9AWqf7FZ4LujE4jInn9ljBb9SAEM4diT7Znmo5PyEMvPEx21Dm
z3nK9Ci0Zl98zxNmefnjHGyoljlPjyVBFSWvqNSE0G+5xzRNiEpvT6pgsGQ5Gzu83XPwCLZ1+xrm
3bCXCTl+tqdR1YQ5biWl1DyWdiGjEHo4LnV1qWpjibStjQ4ebVL/GjL4bjGnDR58JZZzfyR5/HHp
b3nOQMIrPriQnf58sP3ovDrs8jA7Xtp/itgycAdJKSo/DHlvrrOeWjCFqpAFZCVhgfykEr0LUWo9
NZYouHlh2KkPHJujkE6HIqhF5B+RAfiHsqHBmH75Zjc7fCz6Z8vo8/IbdZIgEgPDHHqq7mmJrtJs
ehbQyWoatRWu8PLWtiPFkqu+uVRpevv5XvIYRIOe9u4g4/i7kJa6zk8poq5SbmPFizRiFLRdzQR5
mIoCt0CfGuJh1dqC6uQbfN0TL4VUYD/8PoBpUqj4U+cEIG0f4/I353AS6JpegiepYOmrBu+2M5KY
uEYGSOJieYTrTYXjdEHLw/RdLN/+Wwbi8RUKeIQYEpiyDMdYUnl6erIpsHFyOUjiJBz9NaHmV6AP
WPxbtKNADH/Vu8btOGWzHSmnFcb5ctgSWC9KyE4GZeNRIFLfsoiWKhUkWvrd32s0j0yhNUl6psnA
th4YzM7Q8FNsj66va8NFqGbhTrAHYsfoXoIyQyvV8DhDt3LxXEswnaiRoMeUyMSWnOF67LAILm1I
oX9QCKgMRdMmP3rzD7IqEqXI33WmOc9My/PzdUf8o5lfvfQzAUEJc/K2eDqYBBdexabcWOe5zU5e
E1Ina8z8ZiNUuOOFoGmtW2JvVwSf8sI6tbxZi02kCb5oXKL3VqWbc8EdLYGwI8B+7MHz/WYuzXbp
EEO+GasrDy43vMjg1bMJGkJdJtsVHqkE/Q07Jmjl0si/pLUbY5oP1ZfnQ2t0lSW1vDo0sKLV7vkq
cgrJpTgKZTGeAo5uwPD7OHUlSbgfxEXI3JBzhLOSsoTTG1TYG/taS8i2JpE+e+XdeG0WFG5YLtkL
lbWrShyzI0Y77DUJON9H6bFzADMNneORjZHNj+r6PnQ+jlDdRwmLPP/ANVSp1jOfFi8GpeS0Mqi6
8t+petYRfctyNuS1q2RwzV3cpIzwn/38wHmbGAOdDTsCqfunxs0smklPJvvHqSYg/dmqMBmvQPsE
nGxMX0eznFxO9OJPt8eQA42iLpSrFq5Z/ZPxzCnLoRje4w8nxO7rkVbfJFtqcuE3Xzuv+Lxf4412
k0+EiPPtqlh9FwdSEJnl8xz7kqP0raL3xJgUw9WOEtXStHjl+4NNO6j0EVwljD8JhUnRPUdvAWdF
yAg9fB0+dmuv0pbho9ho7t3paYYwyPsMRLZv62qwO358YdGxxb5tL/drslltjDZxgq5SLRzrFMdG
rEa+Jo/DilMQM6Xr1/KGewEepDFAhmm2DGA0yiI3hn9AQfIkghAHwedFXm82cMF4GrL0XFpr21ul
IlBed2DtpvUWZdalTzncJyKPs/dHql248G9Skv5FMA4cvQoZJFBriY95jJO0Ss5fCybSeTZ99kAB
a7DdJ2kujC8Tc5w3o9svjUDyXmbJuohlIHyaPc+dx6pbpOIYhmz6bAWha/Et8HrbfMaqLf63OLFj
cPIg2yMJcla8HGVuYIlZUHnxhbV6Z6ov2+sbX9Ys6ZvfDhE3598RDxjYitQ0p/OyZ/ntNO7Pn+bg
bkwRwc1uFPH7GOm30PyCP56nkgJbxjHKubi9XmtkG18BGXFug8kilR9ECAkLs8bIF8SCe7MJ1trC
ZE5eR6TzjcXpMIHoZ0BAh4VSSRvR2rwCzUYbtjLUK2Rnoxq6AMJkbbRa8MPtgVV8KnVY9g3GGq5Z
6z6plBVpkssPpMSbKSrF1V2MWR0gwvGibh5/Nf69N2vs1U3voEajyOxUqw8LfnIKRZn7HWVsbUBL
QLyCQCtRZWBAm2UNspaZ8wPVuOfOhBKLcViIYFSi0f+IEOjpjFnuntNQh2KSluaX7ixS3DaBcYEa
sCpr3T1JhfpoVyz6o5rgkJVmxp7TuKpzOHA69JD8CcolN+ED0tvAUFQVtKxVcE2J3mazhjRnOWTz
HLmzGdr1Kvskb5IGba9IbqwYUxkuWfm5enhvDn1BwgWdn5nhAWbZwBr8bXjI62G4tnYlgYu9PwRf
MPN3cBtdrdfNozrxhZL6YUJsRBKCY4BDbPnq9o39scXzNdP7XMP3MYunOxCx02IBqWaU54AgWoU8
SZkbH+4c2T8dKLwvKVgrfVq84D0Pt8FVtlMPVpAMJ5o1R3oOmxcz5DxtROxVJxryHIiTGqKv2Cls
CF2mP1XJxkx3SXKAFSviAwaCcr20ai9JvThMnnqnwfWZxtqK0NRzFpnL0EBAJq+6jebWkvOGVvWy
uJGTY6vKKslbMKF0byjmrVvj+Cxx9+mV6DRoC1ra4ey2gbqKR7H3XOmjwS42bxVD/MfiRGEk7pKx
WU8GawEzr6GMFgzmm23htInfZZP/SDceemyp7w/JWLWyVI85u+cjDwBniVp7io4474l6ZUO1EWjv
33oSrcGkl+FJk5oz9T4P8xwNWzY4C6rxesFbyoisfg/0B2r+obLJsiYyFKmwFAuTLp4KqQ56gFoA
cOPakuHd0/0nIjDY+UrjSRpjnb8PU233W/ZRpNJLcVdGFsIb3ApQtKpbxqJnD2SV9SxpavVoSn0P
7M1VIngs0pnp1E8XB3AAZrS/9bR2c+usYtcrdQ9PH5cGyVFagg1xfSlfV+wXsLUFEJ67RUJZitg7
imrpFC0p1b6nYIZMFNDJV5OqUC8hMXgz0xwsVq58jdUIMs24lCPIfN33jvlhHlvc8kmIY2v8ULzr
DZ3/WxywjfJROz8uzgRIxoaQcYWXKix9+DwrlgHh2qANxDEWMK3QP+FH1P1qYthtelFSLp92JEGu
85xXLqu+ClbTBhnlXiah1UBvg2QMkA8J+Hlz0i6Ybyr0XagdHFg/ADoBEj0Su+29avGNGb+xD9/X
ZD7jZaK9rfDLkT1C7v45qGO7FZzrLOsxcHA2cN8l909cLOisvFtf7/krMGst8Jqk2eE9wFW396M6
+I/5s9nSH/OTPOvz4RIqlraPe8VZ/VCT/lCkhxhtOvcnECv8Fa2mm+5VFdoUXikUFhkSp54hmeAP
jK5y0krtEYkxYVA7gExQv7KdqLbBPHyzfGAQOBfrR/vfJr7ZflwF+i7Y1BLRvCYOmK4ddHsCeub3
qEzzV/9/LAZ0DNCAY/8wOL0z8htJMrEFK6zC70fAHzp1VHvdoz/3G3TRNUq6coSoQtp6FDj3IfwV
EyU3Nrxg8otD4JrKr3xCWy3/UFwQ36st7VecOEGA5l1iJA9VAdkVhYK07U3vzIilU66teNBpCsbb
zTRjhlE7FZ0cMlc+9ET148C9MoTd2zi8az2lMN2CXrtS5+II6Q+rC7VSb+kMycpU/0HUzoGoJMip
tyx6c5il5JeptZavX1gHa6RZNMbHe6cb+1nOG0OwRXHC+/YO6K5NZy+oGv+eybQlBht+VJtaegiO
CeeCYSvugU4B6F1q4FhqWKTnB40gKsxN6Ez2qHQXOQ2C0qY1IDDE+L3aD6m2eF4tIq2MKeCJwaAU
xoUcYDc90fxCF8kxJ76c3QPmo0zapWM/Z+jBkXiZra2ZxoX4p2XyMnsgID1SJjDFRt7qY0ZwtzsF
iT965pERJIm/7/ZUJ+hd/pl5ksnMzVz7pINHkjvLckXM2RuH0gW6i7GLk3eYCmbuiyK+/1Cn9hZi
4EfMxfE4V8Xv14EbJpWVD3DBKc6k13i5H7cFq+tO+YF3se4Gl6H2pFk6W9bn63Ze+JTA0Letk26Q
bGLpaKYZhTWFiFtVNdWnjEtviMzoF3nsZv6qaxeJMoq9qNQrWlh+PsYewaQoxqH+Bpkk4eoqiqFy
FZdLYCnCB94GIUKaHZ5VuGZkwxJylUVOt/bC3KNOJZgynpKDHmfcGdiDw8JEQ2wGnQgyRDisqWQF
FrJ7/xyhIM6sBmdEPBNy1KtsHNinFDi2MP58EGT7pdopyVeUVCdBI0Ms4nQee4XeKte8ITOs/Goz
/9Z5C1vsRcC8sris4umf+gg13/GDejS1H0pZY/U6F+XpcaOQ0IKGIvkxBMlRKzfVLq5OaFLwwkEi
vw153x/aknMV+sY/GBJQLajBII4alseLBFbTY0Wb8HhIoSQ+tgN3EVrvEU0HMzASYNl5vgGHhPmA
yTSgzI/aS5po6wAhIXGYE1VXbODFX3kflY52vrO1igLaplyLDS5hEnT/5T4NQ6F68lZrFjagKCiM
InlMk1pKnij4K2efFZyjnDkXCW28TOwrESa18USM+b8yDscjY8LANivcOWyihEv5huzr9M89AMLd
tbCcMwUKSRz3tyGcwQcQpsQuwfok8TJ9u5uYqHMEVQHGb+OuDqpZz2sKZo4kA7tGiXwxyafAlWXq
Grb+nyPYKjcspTAU9Hl9ntE2iGpLg1h6CdaQa5tJCddsOlm1Ont9O6VABA0XYkv2K3xB9do/jwPy
iDay47Dvy20EwXa+0g82tLHU8aJgiTBhkwBjso1NaQ8XlGPP1bSUXO7Wu8F0yf7M/OGL7ZM4aH2i
nlfw32mGCEQY2spnkT40BStFW30qiZOmzKEXszKZaA9pmhBz249SU1WhtPu7Xu22Z4wnppyF3LTG
iOmMhOodMj6RDB8UMNxOZGISnGvVcaBqu78CFxJtx5YXr+WG3zDzslpCdqE42nrd/fA7uBH9j3Z4
yTMqdD2ZK3bVebthr+Lq5KR58fbTxrJ3qyQTYXVP5aQBobh/BBU67gANPfVAPQAsqo3Z2sWuG5fz
02gd9QtOP3n3nnLpB8rmlKRQggRgcs0yFaE8jTTCsGmR0AdbIPgSv6M7RPxasTct74bIPZdYrkBn
bg1jEs9N9IxhD/aLsX5Dl7ru0kfZKYpXZ8AAQv5fnDJ9gZkE39+Vw91qQteS1iTEcm8KXlVszGXd
BDnWFOWoR0wrktJO5c39ma0lyF0VjXOxIe/oCBbd1cTL3TXOxBhvBd23LG9WQRKeNII2e/k1wRUu
Hh5UZNA4OSoULZC9Om5oqx76NoruF0TOZ3uxXd0+RMTfbj3pgS1vgv4+H/Nl1hLaKLDv4FgggMdU
6GU9foZY9JOIdPECAjNoOrm623+1LevOVCaoo55QIOEvN5SpZB+tqTgQwspHuVeAxkH5DK4uIQ1G
Xfp7pW1MSvygtE18T1S+L+9DFOu+nDyAvcY4TTpJU65VlbEmAHRugCIELDCfEKJzofokPsyk6tKx
10zU13m0loHOebWNM8JDMX5f0if9G/w1aiiMuZccRwA1+kjMh1Xowh/1yJ3Ju1kBXPAr2DrlGgYK
CJgqOBZ4HeIK1Od9btTLNOFH7YP9wl18Tgif5FlE6uLvqO8tKOYK9PG16Fc9Xiib912BuOynJ1jt
Sx8tE5VC03LE1BynuuNg7Vm/08LCgmBh0W1ZfgWnyG83wT9TFM0p5gOMANlCdE0jLa1PFo3WaN0C
kYYZx0IOIi1U1t0ZAeaHDWhKAHBMvfEBm57n8TeTA81WmhceviEm5THKVu/n8roiiRDwoDYqPJAy
OynCka0/6KvM/uJd5R6FmhP50mev1u1WzcKj6EUIZAPLPTncVJI8BelJuiEF1U7Xj3PSnHgsYKgW
MSjWYIpVTQI8XNjnCwxorX/LFCIAkVIHgH45nLqnbNtbSml66UXCPvqUZAGJtLvM/nY0t6oeZ1yl
CQxdsmv454Y46hQuP/jIb8oCKIIgilgNJN860+wrlDHseDCz+g+txMipCC5s14Yik36zJj/zxklX
KbmExOsYaxEwd7bQuLkESQ0K/cIJ66ahNvCX/kEUl3eAbcdds54hSxDx172tnhAKIY8xMQPaUfNS
wRlBvgL46ooOvtYJ9NZIecYcpCfCbmTQ1EmZgfJqTs9ka8IPWpr0Z8G0PGC0brIJ+UDwZcIqn8Rd
A+zQIoXtVgohdpc57UKd76RsLn9RYhJPeFEI0taJ45r/2+1C+yR8wM7lU/M8yWMTF2Av6fxYZnWk
lVLstOL5C6rZXoGQKcSuozeDcO4iAp1bOf8ceeTuSdfVEj17zTgzVf+4EVlq7G8s35MX1ervoc1l
cNZrLNfqYJiAuImiztlhIiZb609yqBP+cTASD6wVSZQCTMmBp3R4FQQ3gUoO/tf5FpKAkjBGerKU
2655E+V5CUXe29dpyC+Q2E4OmC8GtgQ5ZKf3O18FddB8yJXNB1Ew4xa+TK9EZf6WsVsZ0fyUBdPF
+l1Wt4Dnacr2t9pVG9tsRlDgEDDc36cdlME3WyPJIJVavGD6RkTeBgqj/5Oz45QtsrkWbr48+3TM
+4u6EWDUYZuxZlbr3DFGbb1eERJqrkBsd7HMRAQhY6wzIvdpZjmfuPWI+HDBRIhzxO1t5tPgKppE
oA0nQcwKwaMlFgDkdXg31RWHRGiUHlrgW9xkYFr3EG4vNXZFxY+rrdJdetcFBIH/66nMNyEUVDD0
2fbZgewjeWU4qMaS7fXDkqw1hJyMVv2EXlgNp8Zl6yojNIBkUVhE7likWr2YJW1Lp/0XoRNQCj6l
+QsfTd8Od/ENMAfu7jaQt2fVcDs/lZIRfUyvy7WIrqQAQzzkxYDYFdk+ThQCYKnvjsSie8ccRvaL
MtR2qFUP9Kvbqx56Pd6MuQolDLjj0osR0cXu+cuyZxJ2y5BIB3w+LZGLcsEOAznt1i5ZrSXVwNHD
FCnfckZxMpwgQhb7yuRRBJ1iZN4eI0DToZRtImbm9RX5pUWqEydO3CPypjLYtqsXDGv8OcoKYjV4
gH1Pg+11+YCseUEj5yOCUFu7ovSD355r1xZbgoGn0XCYhf38ZhNiQ6TrnPY3xOqJu+9qoCyloFmw
Xr6xOiGc72p5m7qyDmCQ9q52x+05ud0Fpk47HDy/t2l/xkMdUl7ynv5LWDMeYtx+8VCQTB9vHACs
OvaFOwbMu6A1m5VQcWio0nNvo+Mm8DzZ0h/CU4CdoXq77zkBYWbZ+r84+NtGf2tI8Er1SXXUq8N9
iJXmvYstsZudxRD5+y4+FRBk57KOPmbcXpaUhn/kGkPbcVTqGNSQLXgfX0r5AGT4L+SA6RBly33O
oXqLZt7ACsaXYZamKG9wl7PboWrb3az8krPFw9VEHeVkGWjoMBl0EAFq/5T9bUhslq+HeYpKbhrX
wwV3e+MLJo1m4VvrgXP/Nw3UqMKb3XPsrMjiRBSFiEeJoI22XimfHWjWDrbgK+DhKdlIOfEAtVd5
gfrF9JfL/dGUQTReuV2kW6fo2lsw/fb7/3Z1PwRZt3SqoLf65mm1CCVw05QA6r4Lt6MRjJuGKu4w
sAvVUdcQ3MneYFKY/Bevp1XdXaA96wFxAeDm41NVASI/jyEk9/cJLH67fLcMUMsC93Q+lamMKcvn
xVEmm8OAtyQ1eSxi01l7FkigLpLJ0pV74JwXdRer9HzBmprkyMecVLFjbkzh9wbRgg+rmmzDzKJG
YYdG1SRvoc3fz0CSVi+5juKojH7aN4S8uSR++u2O7MIUw/wPK2nCPHUfkoCQ3i4E01Q5LAqi1XaI
3CzNwjzYxMlkunAi/Iy256UBMaX98ISMByUnWoaNRS2Mf3jamoh0zZHWoDmGfmLjDd08FPz3xlVj
uNaIUCRylK8IjB+l4eoXsHFJ0hVNKfv/Gu+fzN1bjgcQ1DWqN4aGb+wpsl3j95qE3rdiP5/Ojm7F
FQs2Bua1GplPXV0J/j/8nA5eNusieS3DW4py7pEis12/LZpPwoo5sleBQhKnfFiL88RXA9zjpF3T
ZWSE3eDfzuTVHeBzEQbUwThvRI9J6iOshT+E7wruP3mJecPl6hFvInA7eFwUax0udWn3k7USLyXT
3mAtc/bBP/CTsxdbPMv+jH7T/VavP5Xgnoavgkv6AyGfKVFU1JiLE6FOk/i0oyoDoPqj4DlUj2+H
AawLmC0GRipNVr9M1z7VBglqJPeRU6ZEbNx1pmU6KSHFocIbPstpkWd6+42LjioVnIw8siArVvOx
J7z6snHONHS5GSnJK06LYm/kiSaWvUJXLBGClr7eGYYYPXDqYF9zPqrMFtJX5spieAFqME09XpEm
hD3eqoSDjmY+SAleOplhTnRv9OWUc1O+qzpUvaovA2BMaKcjT59nxHZG6urEaJQGeZ3yZQv+1yCw
F4Rvx+5k77ladjVh3d4dvTMvvyotOMWpwIb/qeiz7LOw3AFIXr+spB90pFau2Rz+nw+Kd6/I7+Od
k//EHCzVixoVI1rl3kWxoCZ6D819wAvzEOoX3Peu3yQzq44yQWpelkvh0xBdhbR8V4f0YyXrSCBO
cKJFMxRc1vTRnMN0dC1OEGC3HNIh6OMr8F3SqKzYWgXYTQ60naxQenZ1qnCRjnjFu8vRgM2C/AWX
KdsaK6qSanI/2S3/730L4SQgxaOgJSmkuWP7NxvzyM3b8cChRLRRUZ9iYEqOrgaGko3mmIDRHjxr
dbpMQ+JC4dgfxJhfdKFbeqoNgCXbTud0c7IKomkRQn7wZRILNxVvoMM1+cMjNmBBarU9WoOSN/y9
WX7eEsuH1qQtES4I0ArbvwRUOKalk325zgdVTlUSz1mxTEVsRjp19xwJBdYPfaxGVu6dJDTiltjL
ebgvdxc9oMOKIT9NaRDnzM5u/AYImgJdht79vQW6QeT+Mi/ir7kcrzx5jcuFPjvFhkUV0riROrnS
73wWW2nb491VkKv2Z54uhpl6cakXfoedYAnnqjE0467ZwWG6HmKZjNvUfoQ5cZNXCBuZLsSXtrz4
7WD8OWDsJY8u9na33dDVLspw6O2dKxeGOK+Agub3Gpa/eUjPfPd7lOSvYHlPv0RVOAZ0x9m791r+
4wscw8PETIN4yRd7K/R5NDoDL0OjCos30PbYfnA8J+UtY+bmGqGSHhN4zVgdFgPJk+R0qbw2A6jo
PcPbD52pC7NbRCpvQIvQbk9cSmzCFMDs1+5VKNCMxfRT7nz3e+2V4Y1u2KC+vnXmPCO/xngxtJ9G
J6OLfi+482IkKjfYwpAUKXBZJEpkQhoAyvKyVjuPEGAYvTOM4PA13vWHU6MGy5zaXqRdS/y5iPu0
fWI3+En4vwan9w83iY+IC6Y9gXs8PCb4oZJCTmDRlm2NA6VgjhDkpXPdNFOAqrXM1IaPadTZMJwF
sFzefvHz6uC4AXhEsV23V0glFqy6izM61tV4cm0KKm0m0UTJR8Fuxdt/Lk4eof+8QbFVI5+ocrNn
cGPUULtAdr4Lpb31jdrLNevh9UZCT5icw2mwk4ddt7D5iY+6sEguua+Dk+flh/rdPilrhPGPMNdP
sNrCR5W3UdmKU/YzY2a3Yl8uh2unefOwz3kXuPBrRGbVWoIO72/lhJkHhjxxVCJlk+0AxfN1SgO3
8HyKKb3Yf2UQ3Bt7YjzDwscsPOxRXYw5DLzMLWq5jYomAt7Cx19LUlbUB3/ttyXYAtO6j00m80sT
ed9lLfJItFVPswyn3jX40799i7rO30ebN68xYVjvb3XMRM1eT4stalrP5/Q1iswY3qhmsKKUW/L6
9jAWT2U01rP3+1vgziGT3XA+a9SRADU1b4pAAK69okbuuldvWjPmRy5AqubcYhxpZG/P/9jLw8AV
quT/KGvA1fyRiD2HhhuEo7Gx9WbA3ZmLnjZQZFETpsgwuDerdZA66TgFXJx1q5S4hYLzuRai9D2P
Y8+Tx4qX8P5oe+s7VG+jDdC9pfeEDmQZQ6mV9nGs/x2Ok6jRSoXE5bFEpuHesv+HJANxwahtHjz2
Ji60lyTMRmS8G92feQozFdBvRgs7vRhwG86K281HhnwXGv0rNQhljvSKrsj8Ofxs6iBDo3w5RNkp
rQfeE1s3RTcvGsJO4wVfp7FadfIsyzQqpLBKCzo7mr0zdE0WmtoRwRKS7LVg6swAguv+9+Dtiy7z
7/rVN85rj6Kg/AYrbX33IgzzTBrrQWxAmwOmkaGNT2LvhuxcU0fNvHpNrBIX+tm9Qk5hZEJY8N5F
/Vm9+z0jLBSEEj/CiD+wyR/4iqDTM9xp9Bk+P3DeLsa0gsiKjTMRCTb6zYgSu1BJhXuGMIEHH1+d
ILDLwZQ2bp/eTQpy/yWsJ0GdjTPV88V5N8BeLaLkbSBzKQzmzynZHWq3hxo2VIQsdnJ/2Q+fyF0I
1mG/jcwAVYC9Emn6tOVn6hZmDbc9u6zy4jyf3LOKTCjGTW/upZmLWKKTzvGYqQJbeBoYrjZ+KXWU
qTtWVuldCJAXPJ6tMASPAu6cKMAejh30Ep9i4qjcWkbfNXzomuOdFOQKBKCSDO4iPYrrj9lhXEWh
SLWpDoTP+kwSsLroY6l6cDlfokM86mGz0ar+g6u+hAgNLqIbqlgloq1V5TIAWegzoIpwmJV3uKQ+
NxZYuXidu+g4AAmyTm/7qieg+O3Em/5wVLbBrbiw/eFs2mLsTOdt8iZYZo2iREKtfyELdwkKmC5D
7Quy1WAi7+i0sn1G7HKW4K4v58UKV5YxAV63YcFBiwVKAj9imNhlfH/xL/SsF+S6JKdSHWzE8orf
LgXlVZ9GIcniQicKtUQKEZuBZLlJVIQ4vWI+kZuACTwuCwdJ3p7h1IZgbKzEufaWOxVY9j8hgaB9
H8Rcmo1LUQL/dYUwsiKJuUCPN/N45C8RXi9PtdNULNYUPoan9xk+EGydJUwAOj9hycj41nVa3FkN
/0K88jxJanb5J8aAlt/vHPRjRmeUD/PonMsQVd60j604NSQ6HrpnT87uKfDQquH0cVcIb4ug8XBD
67mZGP3iFOTwNM6mQRkzn9uORgZXQhptmEmEEReWvfu9EwZcbGDM8eu7KtCs0XAtw6milm1kDyEz
DpuGdLxegXNTlA0wD9rBXc4IOdfhC/z0llh80AmwcevFozQKDCJPLGbaQhmvpWwEZFLphgpzXEaY
yDljz/OkE498lv0N3OueHHAoVN+rL7D5/CXC9MsM4O/2djD3Zg72PhB6ecML/Qucjpd4UJgQndvI
MmOeoPPI7j2s6xCjsOhpCrzftGA3w4zT0VcwG0Wtt/+IqdWY3R/kjk4C2DOo4rnLBny0wucJWlDx
b34vaTWaXuJ+K3gegHtdQbpCYeUD3UsuOiInIak/UMio/A37VR/YfE59zUnMgEtAu0CwfnheteCm
3KMj17HA9HM5YeKIFfZ9yDx4TmzyQccmnU8Z+jbbMDm7cvCla+rLkTRvrpLRbx0/3LBEgGOuUVge
zuQ7Rnbhlq6o7DwE6j/7RH72zCwS8Qwo3t6SrXF5ODnBjwFQ4DUUcqTYQw8IMs2/WxLXrn6bS8tg
ObIgmQ49dJ3Y0bzWIoyzt06i4tq+8pMi3ohAWTdRenBPIP/2t0C1OrHsUK3OxRFGvrOppIL0A5c2
PqjtCp8xWmzMbILttWiTXioVxO2TF4VWWGx54ViMZBHUspSEh5uv7E2QD6nMZKNR1aup
`protect end_protected
