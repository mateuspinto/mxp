XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)�DXt�=H�����u:��-JN_�}kW����߆P�t��L� 2�P?S�F0d[nſִD8�8����Cs�60Wu�1͂�V|L��E�D��"*�s# Y�H�p�;�ϴ=�E<�Jrj��@0Z���L]�C+�a����Y|4麖���ӵ���/��N|+��r�8
 �]
��{'��8!l�xiJ)�n�e�X��Zʞ��sQd��~ �4�bŝ\�� d!y����;�KG[$?��L���1�'^��J%"��R��&����Ͽzn��(P�ʬ��vk $�z��K���Ea��x�e_��}2���T��x�h\<S��'�Q�����V7��F�\�1��a[ġ��Ϛh�*+��E�9���k ����z�p�"��@�j����x��;3���lH����(h�j��K��My`�����^�&B�;�Z���p��=�Ŀ ��0�D���TY�BZ0���a�kl�h|�Z���+6yUC�φ���F�!���y]�J�qG���Ά�������w~����=���dù�������z���y,0$?�e�s�~T����t��G�b�BQg�z��2����J{����;���y�Ns[UT[i�#/�GN�}v����j�[}8�5�7|ߛ�����!�}������N��ȈV�;��$pX"�!���>]lx�IC��]���Z�R���)��\uG��߈���/O���+���)�^�������*XXlxVHYEB     400     1d0��j��)#���˶/�mR�; A��x|k���*�:���U�ۧ �v��a_����gCYSR�7��i�cmg�F�T��R��e�b�����+�J��
���Op�f{#���Ð��:a%ձ���ҡ#b�!�6U���f�܃����l�3�n�>�פ�-4V��	`pg��u	�@���ޞC࿓��}�jͶ��St�{��0Y>z䈲ݢ@�ك��-ʏ�PN(���9,�J��n�	g�5��?�c����D��=W�d9xt8���m���K���@���K�Թ �N5A�F�xY}&�̄��pO�L)Tl-2�}�O�c��:�\�Q"���;���Hot� w}f�A1ȖЧi�!�yP���|�����[!�� �&#�M��a����%����! 3@�;�N��˗pF�Q�9wN�-�f^��p������Ҩ���!j�:
�����XlxVHYEB     400     160�l.�ŉ[�F�2�ƶfݰ���0�pGV�4�Kr�ǆG�e"l���*[`t�~H���lh� ����]_>�As�+x��Et�@�zp��k�5��Z#��Ay¼Ǉ) ���J����0�	�M�Xف��^�yݡ�H��-U�/V��cE�Mq*����i~|�����pȞ�^�"���e$��'0�v�`��Ķ�l�?�Y��d1>)�M��h�1o�z2*3~/���@h�<���zĪ�Db�[5�m��_�~���R,��rf�u�A��W,�!�kj�)ly+e��RZ4=@�D�f���+���$�W�a�¯D�䛾��w��}-=�a�ѣ
�[�%~(;���ԧXlxVHYEB     400     110z�ؓ�6����������5%���Y�-
4-oͳ�!�="�f�x��:q������l22�CZ)�ݑ��դ���vT]����,l`j�!A!�cNk��^�ָ�;>��@Z�ZG,3��x�������BA=��@�Y\T7��	��Xh�=
]�t<�h%�.b��+g�Ń�հ�4z�e�����/�:Zy*4裮��*^x�p�u/1;\\j��^����@9愥���9y��1��i!��u3LbU��R������:om��2�XlxVHYEB     400     1109G���]��.p'z��F�,��,T�9�A3lBb���UA�d�z����(=F�0�zia���]��G���f�C0�'Er/3Ⱦ��q�=��wb���P.x�J�*15L�@Z.*ܱo8���#���%U܁�NY��6	�ү��}q�A8Ӡ����(��߸D��ZL�t�i2�B �Y�� �t�P��������u27�j5�*Y���F�dV${��FX�u��c�%W����˧ۨa(��E����1ݿ�>C�G�]��WXlxVHYEB     400     150��إ� ��l�>�7|�u�u
�n{�?��<:� ����C'$N6���N_թ�J���SBK�H3@�R���	�������JC�������b��Y����3�B8��@Γ\�a���i��o�݀Q����d�a�vcj�p�pKp��𢍗\�M��ɒ�/')*��LK�+�c=�ސV��4t�彐'��[V�����?��l�08�@f����j��ݝ٭�M'C���P�r���j���K�x�8x�؛ �Jq��,�8�"|̀@�J�u�C;⣎��E�(�9� �&���P"����tS�!�{����u�j��O��ڜ�+	��JXlxVHYEB     400     190tڠ?��ʴ$��/��ۣ��J�$�?��w����B̭-�����B��G��dl 
�0�c����+��wlO��L���P]��M�̆0M��8��l-���v���ƞ�G�%{'��憂�Gh��+.�%��J�Ӵ��R��~��QAQ�|^�{�����tN����RR��]���D�����u������He�N#�v������0��ܞ�Q![2�mO��fƙ���O����'9Ӝ����:W�>����K�)T���de����7=�k=tZջY�!���<
�'��9r}e��t獵�m�qK$���aͼ�n#)3�gI�=�K�����������Vi8����' �L����O�*�:q�fz� -ߩ�/p��1ywuFu�u�՛���&��XlxVHYEB     400     150#�p^��e@�^7�P9�,�%L��P8�D�{�� ���aQ��T��2NO��
%�I�qDG�B�h�a�m�Sf*�����@PnR�<U�*��*��M
1w����ݒ�94�J5�7�.�T��9W&$�R�0��0w�	2�aĉ�p;j�P`W�Q���������:�SL� ��d~|�~8ҭhU��O�gs��AW�%�:8��;/�����C&5S�kD[��R��~���әλ��itx�]�ѐh�)�'I7@z�~MH/�ۙ�U���:)���8Ykr�6Rf���0�A �6����_O8�oZu2�s�P��i>C,xXlxVHYEB     400     160��[@�Ruߺ!Q�Q�u�KFW��G�rGJ}�0�H��^��j���i�al��?��O(���TmZ�m]_��`R��,���+5f��A;��v���dѳ����[���ڝe2U��z��N��a�v(�}��P�R�"�B*p����W�hE�#y]+������'EC��T����%�
���98��0��_�!-%)����!��x[�f�ۍ��b�X�ى����Ϊ�����/P�٥X4�sU#8BT~3+hK��iU�R�
S���L+fƠǸP	��)Ns6 ����;ZD��*sb��)M���jqV�m���CJ�D(���ᘬǄ���sIeIXlxVHYEB     400     120��=YB��W! Ug�L�~�M�&]T��}�}|TJV·	O����c~S����XJ*DhZ�"w����ͬ.ҡ�W��m��_�q��h�Dޫ�Y�b�@�X�`��Ly�y��)Lhȃ�J�V/Յ)]�ʖe�ܑ��&�Wt�|��}�V�w�;��53J#�.{o3nI�U�ݺIh��Z ��cD�ݹ���d��>��\�V�o>t^R$�[s��f�Gih\UF�����a��Ǳ	��	LEo?�C]�����U�;~J��O_��g���XlxVHYEB     400     1b0�5��|����N5��3�����h�A�]|/	�\H�2B����O)�2�fv�r���Xp��)�3]��v�#��{���=��tP��j�i�nޢ�+�x^d͗���]�iB��B�=8��`�ˀ��0��@��q_�@���o-�˓��C� ���<ߍ
 0���݄7OM�qЂ�	&h#���Ns(�����n9���E�o��	��T���mY� >�m��ln�-\V��@M|�>6���F�GwTU��u[>W=$H����C4���e�8��� ��(�0ؿF�����2���k���ZBt�ZA�	���}����/;2�&��^��^�Ce��:8+�<V�V��m��>��s�J/*���Y��v�9�~��T����>����q:�<�]�[1�ivV"WZ��!!m�<�u����XlxVHYEB     400     1b0��+���l��<[�,�I�z�؝��_�m�\Q�}�=���4�/��	�k��[�6�En�d[���{|�=��r���a� �T�W ��)jPO�P*;���Ҷ|��D��%Z�Q'Ydx�hwr�,�N��Y��A1t+�f�����$�F��ַ���>󰅐Pְ=���&;:�4}ʨJ{��:������Bܨd��1��=)�8�嫥���ȵ����ؒK���N�q�l�����9_�Wk0a���P�|]���92�?'����ՉT���"V!Lw#�e������\*ʐ�Hc���6��{Q�Lٞ�O�U��JH��LVr�a�JB�tA5~��d��(1�疟���m��#B��A�$��[�>������ B���w �n5-[��6-m�(�u=f}i�3'�%��XlxVHYEB     400     180i�HF9��
`��ףuנ��,O�k�Uh Ñh*q�TY�S�e���PC�|v�ӟ�K��!�(�Z�`	PVA w [�Pp ����y\���?��;���	k��
���iC
�yޓ���:9T���1?P�ѨQqg�"tG����&�9D�f���؀GF@�Rl��-����O�bV��;NMt ��&��SЛ�܍x+��˂�z��j��]���ze�@3|��j�؟t�:_�/v��/���ve[L�*<hG��������L���K�Rk�1׺A�^<k���Յ�֫�{O�vn��.�t)H��bf�'����6h��m�\95E3A�F�?FU�2� 1RgB.{
�[2=����x�mbXlxVHYEB     400     170M�	R��W/��>��`{���zk]��z9˾LR�+��GE�[n1"E.���}7�E`��y' l��`O^�5�\����Q� �M�b.W{����1H����:ָ_��,s����(��5����,a֊|��H��eg��rx�V^�徻���A$����8�<!~%}d�5,�d����/�n~Meۊ�����(�!�p��~�;B�ݹVa�	k�s
�W+��(!��.�V�--A�9�͍���,�k����H�e���W܂����@���,�y�M��(���:�qFz%[_&��~z��� T^[�g�݆A慑��Z}��s X�vB�*v�ۉ�3�m&����Ѭ�%I5�0��XlxVHYEB     243     100�rp��T�J���/����ݚ!+����y6���	�Qݠa���[�ڇ{AZ��`�>&�@����G�KD�����V��X"Jb`�CrL���D�2}p�4���}UB�K(�U8U���sҝq�s���o�����d�(����X	�*)��B�ų��vs�`c��UA�cv�p>y�	�{ x��'L�@�#jr�We9q������K���;S�]f�7}��(َ���X�^�U�e!���t�h&