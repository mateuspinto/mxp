`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
3NqBMsWMAYew4sXZRAH8KuirJ809Z7le1cV94OUOsQ1WNIg3X38KNA255vtuKmEdxYk98liqKyIM
CLa8fptIa7K7AZr8dAnzH5GgtqynNxHqQiGnDRNIE2TyVPFybbOusCsMDa+DZjqvxPWfP2z4aSCQ
GZBM/CgBlIamqWSJeG/M+JvO1dixQHMsu0FoxxI9xL4tZeG0z8Hcfz7YaOndaQ4rjMIq63risjoc
cbDrwlme2qtP2UF++ksX2IsimYexksDe5D67myYS+vv+U/8kcDGRuqFDaD+UQdpz7SiFdPknftcL
gLDU9d5twl96/jGEVOHrJZl0wZxl89o+smFS/CducHR5dpSt31mtAYsVXXwlkJQwvs90KYgrMVRI
z3U14+IxpxvkOgvigQJVF4ICD0OhjNFxLyh8prJly1awlMK3OI1ll/ckR+lZgPMygy6ONO0kU9PS
rPOP/3XCQZwGPhAWIgc/j9WamprPh0Ka01TrDOAd6d+lS08v0rYmg2w4X3znhQPaGnThM0Va9mgG
MhLN98bvcqFhsNzoJrnkvKVYq2cVOuZOKTTv2D3vgrC9FKzAhFF9xeQ8vznZS6KmZTLGAcA7AH6B
nVR9dwEw9Dr4VsrI6qvUSDL9u4w+6bWpkQ5uLyeDFLoufwhhRN37gTLX8WioN2TvH8Wh11l+Crbd
LLSaNwnYuiT3JlXNZTcXT6u93Okv2yVCNqVkCWHDZtnMmj40WZypks8Wr4wMQLfmdtW+vgdLlRZS
k3bvq9XUIIL1Dgdy22RvzDaM1i9CMeVzyiJw47CveiwGqZB3jfan3+NLvnI261ocfXz3BobaTgaD
G5+/dqCiKw14siVJRuCiZpigK40oCuJpG8uNZBdygMkOP96jRX/UBiC73u8IKnF8GqxI1Mjz8IFI
eYSXS5GhmyIZphQCJpbioY4Me5g9UafY/2Ejib48mewcmLFylXQ/8TEkCrDfnHNlPViHAhIUrVMF
WMMXCoNkzb1CtBelj6KIFeLDNkPZnujp4yZRaYvJ46FsAqmM+RG/znoM4D3In0Zs3DCQxpoclpf9
bgNd8yFxPZ2yj+ixUv32rLBcUFnjtL7RBwJsIHdzYQoBJ6dnLkIaKruKq0XtKNgAhIUycy1XGukn
srvffNUFRnqoqoa2CtzuE/Gikc+gwJI4vZFMBDEO2dwPt0yF2nV/PWL4dH5ziXtfwdeZEK19froC
s3A6oiMBVXs8jA9S1qSdcNk6O3WnlveykNjpTd/QTKwSlKEyIIr2x/OGNFgar/tOd29gH1VFjDAq
/2OnQpgkG9GaTWfD67hrplxV7H8HT3WUAmcYtmJ8TxeiGiskOYFMQkVS4HpaSAPTJhTPlRXvZ4AV
f2cdyHZjMJlhFSr2EGivWpy8uFUuoPzR9/V4dF4aCUEiuizYNTHMSn8Ratwghetnv9W9USmpJaPI
hxN3AhnVE2gL6wwwjM6/zc/6WyBqCD1hWbzfxywpi2SY6C+fE7If+u5Zce77BANEwUa+5VQf91ho
bv5NIEttpJtSNsk1G0apUXo840LKwSxBVuUyjNI9IIhNk3jc5w4TnLnsClgb2D7lZxWj8/d2qC8C
/yeWmqIshFXQleca85zeQqUrlKAvVHW+ngEvnTrLAMj+upoJwpxiuz96Ok6YWksmigGiDOijpOS5
9A2DeSXzBYJi224d+u4sJ8iH7nb/20C+lA6gfhr3rTzr8TybinUurevbe1GnQRDHoKgJcKEfgHXQ
wM9pPItdwUKW+CYPhOpDeRFi2ExSnx1zCltWzF5SccDzXnoh+qlpOxm3SZyRrwXwC0IY2TO956WB
wjDpH0+EAOfW8D4db7un3PFOI9k7P3uhrMEMuiIp175hopXYcL69CTw3PvrVWi2ElUaLa1bZqqu6
/P5yNSV2s0wjqOICxS6zdPDjz+mJLIMXFQ9ztkflYzkFe8WK3685wvneaf1MnSnJeKSvyIJrvWjF
75pmhuR/IEkp03kFYBLtAo50OzYuUJRNWdRGSrUYDRB10XeC9uyZEJzNIubaM7Zrn3TSh6YhlZBM
zRx7q93AIQllEYMMAnUM50lVOCnJTuIxiY0L7JCXGP550omXCfL6lZg385Evt2+CdT4gIQMZl4xj
DdQdnQ2s0W2iaQqCmmfeTs/sCO/0kE13/ffklSTKHEqrOS2TO7VxKTmt4GBrLjHRAQmlUWsPuGMa
yKDdIa6pMuLUQY6qUhe/ZOeQJsRsAL5gg7dQujJnh0YBp1QNMTJTOMP2C116i7RMgYwpzcFX62sv
06oTjWXKO7b5R53POREJNjsJ2fnGH7JO1LZtLbt+m2zZW2AVJZKVlMJbpovwuMdKuGKzO4YNznAk
96rSTPFQDRvqGu+YdQfhcP7AUHpu3rgMhOazG7PDrDIJTIE6Qt0L8tiurjf8uNdCf+IMPloEHcO7
xz9705sxm5/lQteah9jb6oxSQzdYOhaD8LkF76eCTG6euR5L5ypp33rBYnbcBqF0PbBeC+1ZJTU+
48c4+TUzDxW6Hd6btkREBUcRf6na+gWh1DQ6QO+KEW2bxqj0hTEGB4X74JEnkMaVfjJAfwWU+jXu
RhSI95JAaWN86sCGPOZ1yYPZ7M8NkZOk7LuRtJ10kGdeFHmhHTtZpEM2ZOIoeJt82yPGDeXcpkcv
ZFgFN4q2kXdSJAqFdPz0SOuMC42tmix+7EApPj/GyiKARxxDvzks9nL+++5BVwWtVxEkaZ4Q9nbx
5EFiMiIUmZFPvmoYtQRyZpi1f1I76hoPypeTdKVPOThUOvCOgLS3tfKfLcW4YAv5W1lgF7a50t7O
DiwiyeB/ml2o1n59KVYDhBfyJfPMxyg7+jv1FvB99awTlQGxBog/mzzv4j0cP1qhTkzC3LyAN00A
XIaIDSkmGeNPnp99j4DSA1N0b6h8DWj3jMfJ14R84jV4q6FsGLWrFWqYES+o+YZjTI0BpI9Zx83D
Y6ZdPSqc5dEbfsI/tfy16HnYhgZz3LmLwU8qudH7KMOdOv8l8StOVwGRvQH5IfD0PeKSyagMSVl4
Qefo2wDGdELAaQDPkS4NbShBgbGoJ3BsDL1ZQf/qrxlGxALsvNCQ25OoxmaBMqwAzoEUdPv4Bpbv
B56ApyVNQUc4LomT8Hsj2WeES1NneQLxsPyhRHiMtsH9qaes8HJD+3LHrn6TpQJVIhwOLILEWUTZ
Gg9AxBz8/oOoNBq4hctpYP6GIKa4KEfzKnYsBC0fn8vHfk08hvj1ZucLJ/Z2Y0+FeCg/txOkUDih
dUVm1TVA1bAlcMpCx+wHtll/QX1eoKUM9E3MDkgi3mcXXm6VP73STxDaSVu4iqqDPcFDxp1kfCAD
fmJXuzk+BJ9hd0qIjUfHjIj+hS8201ZXvMACbP3bWbB89KMJUd/fkPZ8pS3rTHUHf/CpPflmgBk4
8f6jRkjgOB37pj6T9ySzUDFhFClhXy3vF3KioMA3mTUf6Ldj4WhsgpUKJ/UQ6Fob6CbRgob4gFfQ
CNRAmAzJvEk3EPengXv0pdxtt1bsCKNmL3jHed9LLwFKxyXJWhfVuV4j8GAzkGIZytLiiUnnVSLQ
sCbqAknF81CJVL+tD/QZ8pSitqwlsq5j/T9wK/p9hsvla40PmCOCUomZtL9xStiK7QuEgSF2a782
UfqPvSuiP3145rnBlEn1OV5+VumDclv7q2vm79m1fky1ogG3ND/zZ54VXl4z0a/GBIiAgmr61TfM
aAaXN/UyJfbpsumYUcG1bsd5i0F72lkfkMAzV7ZyZuM7xF9lZgTgmE3AjUVjtLuoEv6IcRrm6W4I
iY60n+TXcwKuyostykNhKOOek0x4K0Hc4Uw/oVQknziw7hREJe9+B357Nk+eF2LRgxy2BcvOqPmX
+oNSYKpz2Rnk+Cv6+h1Rf+He8FVLnEAO4QLLwYPJTr88lz/U0+wsIH1E504g/ahLbuc90pX1/IjQ
hMozwLDufEbgakIRQWXUQAYOIDFiyxs4gJnhY2szvFnQJhjW5omUZ9O0pxck/VYhETwRSyolLnUh
jEMgkcK89xtxI3tpro2EOkreCi6uZzpXHKgvVgmr2+9jICQKg63CSbIbOmzXSZcHBZbjbT3GYThl
75joxSU+W/v1yKnWhLmHyPSa/S30/MszLF+LHSvly4HWBe1ZYxwgkaVDU+r7r0R1goy9ATzty922
QRfGRcetNwHHU17jNHjaVwHoIeQFhs6EJ3U1/tk++/6kmDyTQKj84gw0Xm7ecf0ulpvDrGWP17lF
xkLv9HVfIFT3o1EheedUmOlZbtwWAcv85QY3bZvilnOxooopREPLSff1zar2Ngvi38/FcfRBEBvC
MXTcC7q6ZqXdsKTkRSSjIV2Ww7n0CMF9E4Moas/k4rzExQeVvQev3P1zeyC/NSzFHq16aP9NVnOO
kBddH749IQIxlcmdBM3Kxzw+QbNTyf/ldMv5Jh3xSLc5nhusIiEb6tjzh1vlwIi8U+PIX6vfLPbb
eIQMZOC/DHTyMI/7+tOdsUjfprqvAy+zwdDAbrqBz0Jh1Q8DpAHHzPHfapr7Cmgawo6dFHpf13Kn
VXl58vnZjp4J5zJQrsYebNowIYEkuv2vgRp+8dak3DGpCxynuuuCRbQwcM4WInpm72mMLGsxfopH
Qa7mRfxJk0yJd7Fn19BXDPOimDPNH21P6v5w4sTcmU1LYKv7WPnHhjEyd9/7hBvKxucnGWyaFgwG
OWVgblKma/2x9nCqD4UuIjr93ijzXZflQC7P7vWkxSNfeZtP297sCXH/4z4zNpZjkfywOW3SNlvW
uOzUvEJtZDynhBDFpteLr55zRsrPMLixt+VEt2pRFilh++iKqCxW5nlz3CD1ayE7ka85Oq7PUo0L
M/MNSIEe5THakyaBARxqFCWVZNaAWmeySuuT6FlhmcRrzdcgsA98o/ATAED1xHsCdYOB6yawvU92
7MERzIZbK8A34or1o5NvaMLyUDxCT9CIglj6DR0WS22Nc7GOFasR5tJvntEmMhmq4Juz7IbvS14p
akh5hojxJshTUsFgensQel8WIDnLl+y2iXVfmzrOQ3fwvAq3Doporrvw4XwvDXoZLtxAyQLdeVdy
oHqcbrtGz6v/AHE9jf+jQQfI2ocSO75DI2qJOyCG/cJv6+v7LqQso55Uzmr6SZ7elwgno2SnVbr9
a25dq9vxNVx0gwRaw+3E+erb4WmG/2WYo5d9g+EPmsd/iizTpClCmecAYDIywOXkH3P8DUd2Zxq6
3sXDNhNbnHlB9SL+YoZKj49ue0DLu7K3mJxam+ArkfRxBoF3w4xHVQ5RhtHufnRL60aYyGn87lJK
zD4SigrLtuZtDsqldZ+eKT7Tkyy9MasSZnv9DfJ2ENHA9FK0VUN1+wIZuUQpYtx/eg8orx8CHgLJ
aXyPmXsdIA9UlLp/dKcJYHgcTqYF5AQ/CXH9PoRGJRkbVitI7MBSn/tzsGuf5f6IOW8k+rNT1CW2
baTDdCK4b+rGHwEBq5WX6LFYcW+0XeVAf1OGf/bEbSWGawhcbhJlX8KRJZLfpm5va9xVXgLCoHKl
XCQlWicdsEszLT8a5wOJERBq4kP1rB7w/YQftqteEQfzK0XwhIYzLbIP/vSp+doG+V0CbZOLNtay
P9q7fqq/uzjli5e6sQjtnC01KibRHc2KGdUQ/DtAPuAQmzdbg+P3KzXbE5bCdRAelYcuUxXROQtl
PvjI78yvQFL5AO/G1VzYL0hQ7JSgGPKrq/LPWFVmEN22yui2juahfAOaqbK63RIcSkIn2v6SSobX
adRdyEm0rKCCr9S/T09UNc0ElXGg8L7dFqRFSeVZaVWu6Iw5dD3V3A7Ss0CStiw059fdUtc7K2JG
5sY9EPPR9dEIEVyXk/zfJtUEp5oiE3Cp3q+G1jpI6furNvE8BCgWpOPnymgwxTQYuQhS8Agf8aWA
T3KrNjLkv5G43JtTik+pCzZyCJKHQc82hIH9jW9VM15zu5HUSuu+LP6Zysp1vi8ETwTaoBbIa8yl
dcZ76KbCOPF4vlkawN9icGvxKC3kF2iJ9G7BANyF544BzrgkltRz8ITN3ukjrW2cESPjNSExx0W5
AwVS90maJmKikBTwb6JEkBVqAJW158aORosvEHpfSYpUqEBeNaWEIkkqUMGQqT+TEsIg8sj3ZiIj
4Ury26qKunfITHXtgv1XNiC/QmcELlEJGIC5ZCYWIRjlvAHHF3ulUD4JHJvoawuqZUoMcli+GSpy
kQ98u+YcCrVChNLyAtWawdZQdW3Iaqq/VyBj4M9b0xH77LujHuMBd/ew49JHfDGhgzwhxp7w4OOA
WxvqGUhftXibp1QtFnm99ZVA3bP+lK29+7pFkuhQgN9e68CofN24KRbspgPscLnu0VQlocOF8Mm8
sKA4tj28f2Nh6RQh8bsVBNLgNY3pZwVbO/cpic8uqkK85nc3h2fgeyfQUIurG8YbI1dPQGZ4K3Nj
HZGgTPhlYyAJ9/iTHQsN0+7MiuU+YuTt1inUPdHd/zjnzn5COtVUouuqYJCXJyATRu+F35H5MiCP
VFIL0TW+N67vd2xHhvIT0BBdiZyh5UcfP4fR/7ATIqqLdu4ZQjvVqwlJcrX7EiCvpCqU56xO4R7T
Rw7+en22denWRMintLJc+lN3wp+o0XN/ozRUFiarTed25gaCJBVN+FGymQ+ywE55HcJ8Su4LLZLA
bM7rW5B+qG6Wul3rBT/fR+0hNinX1HJ+zbgmC5Kwl/uGkHqw7SBJWSXUZqh0uN2B2oUVxuc0Ea1D
Cy3QvcIqiazjJb+v1/toqzCDqtPHfO4U7fCl48J0yjoSS5FkEg6L4j2/bEXl9QBf/Xd99Yvb6+6L
BZMz2YEfAiq8c+VMghB8R/u7iLz2r2ZV2VuHZj1YQSKLJqKlnGvnoO6DMEjT3iJgWXGuPZpJs9xQ
Y+TLCc1IH23NcWRVcmbsqGlPWlR2uw+rxc4zi+jdENO//R0fmJ/jmqQvyy9t8XHtw3ZVg81jvV07
CsJghgMeUxqu2nebtFaPAujrDNLPwR3UBeQJskEZU82NurGZtSoA+wsnXAGGJAJFIIn0u44toTLO
NVewCbp7mzFQMXYB52ksMqGfvgZPvbQF5VFl5oBxpa0+lgwTz0kG036mOWHvbjObX0t+k48WKQGP
h7Wb8/5uz9/TKPQIfnFLC/xGD9MgB73C9uIaylkQZjWRrCNwJFBaANkZ+WDpBUj//sUq8fJraMYU
ktU89QbSVZI7rBlkjSJ9VYVmUNqTx6QgUI6zCHQtM3bFMWVxeB5plQetNQzOpgQlk7dXX+o37qpV
Hvifuvxa5/I+VyrsO/++WhK546yIEkj7sVCEoxKrRKCP6gWxLCW3lmw4ORVAIv4LMz3UAf3dzgLo
hlK2wakR5BTRkhZt7Ge8XwZf99kH91Mu2FoZtqs6J5uFvAQM6jq60GZHJhpdjvQUii5Kzm63xfQI
mVBcRy/DAHImrYAuTb1au8/VwjZKEvfBHrsQT0cB4PIZveS/RF7cBuRYFvqrDzy9co2yT4ZQoREi
lJsgi52iR6n1AwcAExyLuIMCsgXGI92w0CrlZ5P/BwyNjLxZLIiX7dUt+1FMr2LPxiQxR6MdWpO8
gjXc+3jxt0+mRIn09m/c0xAGobMK3jpI86WI8aPTxu/udYjrppYQHPSgLX3xSaMMroukdJ8pFqVk
bHhS1E1VOj7ZRiod7BtyPX7WRZfofoyuDByCNVCFPMyBByTHFw/WGlUkWydceaAoT9ZZqzYTAWvb
t2+A9PNtIClPKs0IOfdeAJait0qAAHLJ2wA6UcSxxS73v5nZHOTJ8JGTNBKRQ290G8gof6zCNtWl
pkwOZ2aynbAb3Ec9w3I7J2rQ03w/9/qZBueNz1MkTNYaREGRKe/IcXdM6D0VUr5MQhoVyM7zn95N
q0AOyB0Mx3uTcsZYkkNgyZMJVLYX988YyhAs0S/r42auL94w2sdX2XMOm1AzhLVr1gVIV3g+Cr3w
mGqZRehdv5kwkITDi1OgQpAr50n2/v/DJH4lEq6gGiw7PofEqbUP8OkLhtJrPETFuMHKK3E3rEx/
dglTPnsrord8sZJ1a0/94HuHDmXFWJGmEOiPcE1Uoel9jzlQhX47KmfZQI5iAFEJ+QZm0o922RtD
/ETGC9b6RVq/x7XU9ciXUh1aITBnkujlGmlvfGf5hJ1ifRTyXa08ee3hjjIDEHtr9ts+LZFNv78H
HXvL4blRR1TXV8EAFsB3z22BPh8T6GQ4p6Ffhx6jHb4HAbF7t61qlWbt/rkcj38EBSQ/KPh0hvTH
KMdQBwr5m22N2wHc9/v5uQg+o+zTjAvUQhc/OYQfp4zJi6l/gStmyw4aBr4wWcQhQJqh9OqKS2t6
H09lM9lxtRDyfJJCYQPFOLN5wgnxWjTt8P12U6WC2s3MoL4Q3H4AioUuuiZWePFr8fHOeEHy+Rx3
WT2nky4HFUASvRikTtKFdHlKIlQ5t8QJpmxY/qguHioLoD+c98go1leofdzUo9PR+4QXs9nEU5w6
o2RZHnXMaAcsPc7RcUvTjNy0Xg0MtKyuUWqj2bNRR2GgN0haVc/cRZ3Q1G152Vto8budpAfXVBIw
KNOSjC5AjPxYPWWftpJa9VT80jYRNa87GiLht9RpSzrYQy2DfOwxJ8bFinOC/mF4G61Y1OTr9nrh
l+3IFKmAFRbaPawpLBYhBx6Fo4hkok1O4OZbAEAyLlnkjd7wwG3GEfp/5Re9r8lFMV75RdRz8dXw
Nr9tibI+QuhRVxWsJUeyYB5YL8h56cOjHLXuKayU/gIPRYhq3FHci8b7nvoFp2YY1h7/meVw2jz+
bKlSBGrk+M0dslbFluuE0g5E5ccBh5NMQ0YbdoRv+gz6FlifDlTnVBfiIxls1NHudPSpafyu8PH6
GEd6xmmF7Sd2jwwZQ9H2bzOaB+d8vhKK2p1djFAvEohOu2YYBg4S7lrCUEQE1Sz7m/rJUPOK7kr3
O17eycydsalzhsOA2wS7FLubC+So8Vm70CeT+KT4SEt9c7J4OnXZIpnD2GddWNhLso8MPolupeQA
j1F0suN7CuoC3HGL9uaHq+ACKlMby5NKOaUp0WkLQWYwo47kNP2ktbeKLtriu6y+G55NV55jjshu
0mvGT3WrbLsnAfQnMhqX2VbRPsrxW3K4iBmIchK5BZ3cronEJyvqmLZYammfzEWCTLVCS4vUayRi
6xLzg9O5v8Ax/bim2nc7sFocnhwnrmrlVpVVmrFnmIOzSVm2rQVHAxA9CHCqzkz1KZjuFaHs1oOw
qGWYUuQfk08lXG9zjHNAZAD2eG6wZKlGrdpSI1f9hu+VUsfN8dPg3bnr5VIFH0s1rwrjifwtdlIU
jy07O59xpeNunYdgZXRLxBi65DdzkMOfSMoMkTo/jh1ZIUc5FzUWus7CHO+0q2PO62O9swN8Mm6h
CDSPM8cjH2VeMM/yKpnKVU6bYHFY/91bRzuPsvRg/ubMx51tA9t+IssS6OA0uk4VKCcjbNCLblZi
vigQguu6AFbOwLE4zX2ZXmez/uvkh8mS0N+kcShK7wtVhioJ+mcLYrV1l9hRGfRVp/u5TOk6TjXC
pKy65c/KQGsUgVEUsIWs9sO8E/2BW1tOe7mWDbilAIETm1u3yB0tPOI+Iah8AvT08pmFx0AqD89U
0M2Rs6r9gdQqp6zP0mLw2tr6PqcU4mh1JrCa/YzooZiY5JbaCqbsgCS0EoOt9Q496/lo77ag5D32
yHuVXiShEDCjwMTQLQzUFdOKXCboJB9ASNPOZ1H0W+wdoS12ZJUTPAbzL/I4OfQNuMICd++12n5E
eC5p+gBTYHdRVFKDTAyUSZTjr8DICtwyVjCESiKVRWc4V9+vyPEGXZ1i3DAURNEQNlyMZzry0yzW
w7XXPXDKFZVaMx2s4CW5eA2vUFk/FiH2fl1OrLu4cvFaBtviJtm0oKJZ05XC3SFEhJeS7fL8isQy
4FD+usaGsAaLw6El0AHFUooXDSBlvuzHeaaZCRAsBLM0H6fRvHM9yy8Z+nzzYVf7XgxmDKIfUrf0
4hWGMoKafdtRIn9nZH8X0L38heQ/2sHGnOXrbADMGzXHaJHg2l6mUmzCc6ceZNtDBkP1egWgPf/T
O7iZVA5G+p60Mr/Ys5QyUyiwXOl1EVT80RPF/qLYMZby822hrRJX7vt/qs1RRqNa51drOXlKTky3
Lubne6sxCkaUawX0CzeY3fInvofY47IayaDp2QzsH7RbXaZbVZefH7yhhrIio/+TrzatiZkNhPiB
gHFeiDqwL1H0cg8wsbtSDtkVFeFcC8+PBs9Vq779NDCVBVtBPYnOZ6yQrDXxEW+mdvgHTytTBfrF
ppk2qdeNbafHxEXLzFf2l0Pjwxa8W7vkyQeWDhOhC718Q6CrIRWnsuTdl7r6wXgPK6qCAcu1AGyC
6nORpn0MGnukO016GkuQ4wPLHJS4dBjWT87ko9wadHjmeeFyJ2M8K3V1Brel8WO3yCZIYi311dsY
8kk7zymvYfQFIgFJOqHnt3GCnHUgIA6wMPsGjP/ieNEbFuVEKH9tD3TDNr9uQE8CfJTyMzs3Np7/
GoejIVoZqTGfv8kKdLeDeTnGK2LDyOzZe7pCaaVW1xiIGOpreIsUEhNVq0VK6OYZpVOvoxO59r7Z
sMk27xjUa7MXqtQ9bhQGvtgZKE8TnNAr/quVui45krNlHY1rvQucnHfxXQjt9W+CsYce3ZnJCaLc
8RWgBHRhKUQU6VlPhfLDPUVRD/8T9AzupzEX+TyAd9y8qLIHUqgc3eoDW9OBYgm91RJuI+qqRxdc
FDFrDURGXNAluFiK4RexsoNtKtbEPI6uzms+wNhjZ+syYQZGAUStzCeV75ALvIux70CGy78WMX1P
LAe0p14Sr5rgxDwYV9OlhvqbJFO450tAWwWf5VtpydVwn/1NKFmFJ3HmKhMFIqek2GpL1G5fF4/1
IPLMhCuzE+wlqsceNmkJ3cm0L/PipHT+XXZ4iDdQUUdurHfxgMRFhu1RcamVakMw9a9XKwA/P1ac
sE9mTrNZ9ggpaW+TXTxfiQ1P7m1GAD6m5RxILAbqxlJQOUwk0VTQTw7SA9qKjQb4qRfSF7wIwLkx
73KOkOxxRBVYz5q5lRdlmGefGmcjOSwkATJvB54lhTXea3TfBodj6f7ItSXXFQqfioM1AZHvkq3f
aux9Fb8PXPTAJcYQj6utvIONGENQ0/4dJH0A9EhNdxMl6FUY8b3JQDGaHh/jeqzGDyigf5qoucWe
TMa2xzh6zh3aoJ/M/OVZeeMt2T7M7o16v8Bo/O7coazw7km9nwUiBjkRFX5EphJMUw0qJypkdkkF
Ep0HBnVEYMPQ/5b/3f1d9PS2SPDsobWcFxCIeXwTjfa6EuiC58/8SBJsr84UlN7PqEEmptMNMSO8
tPQ8XErIaoLZGxMxJ8OIVjol01sciJzVRyxN+OxTH682hPd3cNJ6xMXieZA3rpZL6Me9CnXCWirJ
hNMu6PmHjPYsPqsfxhClnu0szpPEnGA6RURDW1n9FywApVUmQBEYvPJAJhmlnC31J531iO0J+HDz
wJIib6Z+10dErCTvg0zOzIcjWoJ331mnw5hTffHW6pWHBWP804Ln4at5XucJSaIz1RQKW0QvNQUM
Xe7vglgmnzTcnD9aOymoBkExs7YGN8Kh8OuVsWV4XvyA+kPMGjg/1tRxzgJOMXfecf8KlkFWzMaV
1sf8wUr2q7xGR9yWeP3YH7HYr7X8XFjqxJ8FOsgDrcyz0+gI/GoZiX1V6TdV+JUkeZN3r4ksxBuF
1Gd/VyYu8qNjOZVbzL0zXIoS7UA0MoIANJZS3EU3QEQNtGMvdw/Ytx/4wlboscQF0WRM1TX0Vwv7
cvgjsP2bkcwC0iR2ZyW6tSZl1bya9JceLRmIvs8CXGSsOnCyYgFbT7+r6P4BdY/2sQfrk+Wx9hoK
MRxUvnBxNT2CSc7HYlzEWNPc1PJBu6TqoDtjyxHqRnZuQFCkWu0YhkkLYMnTOnEuodYmbi++vMF1
5JpacSntD9ktmmwlppEFuZyDYZcNt1y/AN8Qd4eGU3otR/9XQAYKgxxWJcp9IHOkBd9Yw8cwegZz
EWF/tjUFAauJEnHFYOIEe6t4rlVJiLPbiSZjQ4Xz1yXimaA2AnST0Bzj0Nsa5J3fkiDDNhKG5ehI
PnrWRsH5x91FNzjugcygfbkG07hZFDlM+fGWD9i9urdDl6nFJYh1xscYmOJIq9Y9WlYiEFAnO93W
njPJlInFAR56IVsQlQVhGDQZBQdijgwR4YNeszpkpd6yIz7dbPw96RVajGSfIkoJOd/p/FI+Q/qa
n7GIg1v2TFtw/+O/lnFwCCjZ+rd7mT8b9aykm9xNpXSi/o2h9M+aAFMAmg1+ozKWn3goZXPMp1+7
Ur1XI8m+LI9+5w3HBzuqzbgMJ86Jg/eugb//WWcC2lDMMMCHDPQPuPVfRVlzDXaJKtiz9QWKDKh8
96oiOXQPiBFMFkg2RkYfbqaeiL1l1OMScZ1qCwsAm7mtqLZ6xO9q4xQqlCDn+DQ9O86S1ooNWIXj
4FgD5aNs4JutaO4K0ZeWYLVUaS3bAaEL8ieNWi0kLkygU19CCMPo8E3OxMEjJV5taylp3XTr3L2U
vh48xj4rYuZbujo+c2uXfQsX7q8jGTfrFjJqrYo3ev7prJqZSJmUXzp/d8uCvlIe9FgAxWyBlnA9
AZS6yDKXOJVzhqyDzE0aHSu+3F2lsi3G8gOj9gVqoqdDLMazpW5JNOUu3oFEtqaHMk7aNrGonPw7
5P9lrnhPdQwjfqNj5m90gN4ypv3d8VNeCwYvBFeYDmlRsk05IhYMgXAo5YpOAaCvJpbhs1i07+/M
kIzYs9Kpcb1GyFaWh7nACYNmUibdcq8J1laG4F5KKUUWqdlsGwfFxIiXdgukazhqRjkS9bHYpInq
PsGjSjtW/MyRzcRkKlqXsnZuy/FbhhzV8lC5p2pz8eUcFr/N08fIdcyXDbNAwrB8qxwtymAsEeMS
7el9CQOzUGO47K9K9xtaZnqpi5sDHYmL7mGyrWtCpolBcWZUMVzxDhUF7FsxTJV6ShIq4c/Az1Lh
0zwiPCi3HpyL4+jkvCZBuAuA12C4lp2dfnVfk/nRYnFZV9xirnVUH66GwLh+5QU7TyC3HQwjtzco
TfF12tTQ/Rlz8TNg+LZ9QyCiageKlOeqUg90Pp59e1l8theDC9Wb+VG9p437C2RfUPu8H64sBrP9
xr8rlGSBIzOax5N/corbbqam3sK0Ts//pO92y33XTTHOfB8rgmoujs4c3tSY0576d9f5q+K0YxI5
2U04mYf9UFb8v5K7+8OtN0Pom+mZ6CXI4Q==
`protect end_protected
