`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v2YSda9JslsnIPZcTMsx5KeySKJlJOU0EgXKmKI4Dv+qfxUzpN0X0FlGOI+9lx6YuNMnf9PtzNkR
ekcDjxbGAxaaTCpo5aA8ibltdBdSgftU2Kfv6LathBDPQZA5A+1oTRFAVxwFrveIvnxHxrrMfQXO
tS9ro66KcAXSQy1YMh9pz5Ygl/71Dtf6SG5g93ybzFnI+HKGrntLCs3690duSiC6zFMEeZRO/kyJ
irGm2UkI8qCy2hGzMzBmI3ZMXajXxLxtDWkh7BIAbYWeksB3OJrJ2nu8Li0otPpX5LIc/RVcpDIl
sE/JRlIs4JtOBHMmqE3Br0X89f78AqtRbZbb/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
DZ3xiwCbYJ1A/RMoWHamhC/FIAkIeMIZ/ur5XyYU37NpmvYHZ82O6PYJXHFLeN1NCNWy7hHjUL7j
sXZqlQt9d65QAte/LANNvqWCXfuxo2svQstZXrMAbg88OdSlqRU+YE15KaY0PmXz2JztLBU813r4
J15gq2qtGgPoMSRGjn4Zq8nlAkSnkgEDyQFRNlbwUPuuja2zZA2P7tCj8ZN6n7XgV3DPYxOSBgu+
KZ5GvDrAdDhmbbfNhmcwEOeIuH/CClFlrBnXi2EERZiyjIti+NPf5mV2x++GqovIjzRZtyMQp5G9
5URc7M8PAPubo+9UZy3nQKKUcIiQxJykO5i1DhMuO6E45joT5hbMU18DYzqvgo5d0e7ISis6pIIu
GnNkJTlR6uwCQcLMDh8iJqcgoHp2ffI8MNRMdQIHbFlHQEgHcjXJcSxueUUepjO67E1sWA1kiEvt
ktYjA80kLWhgJ38FVwax+o+BxWVlJ7THUIYnu/Y8evtGf3dibi1rCan3Ig/PBXJ7DicG/Cm1Y4cV
JX0RYAQyNBArHs+LOJH/rfgQTzktcTXngJadjckaJbRGDqvgolmMPPn3zg3Pglz5e9FJoOm0yrUB
oFScXuV2g+2Z2NtZXOyeCpP2gfShYlB2SJr65gfJvZGJHmvUzTFhBNgA1ZilKM8xs6+yxcYkcJXJ
gkSGhW3m78d7DXFhLqQ1006jnYmhgLIzDu8kSKwKGA66IOzRBP6xj0F6Gdk0AVaWPvX3sSM9x2ze
g0dBJl/n+DVlAEDup9iElLra5iPSfOZuabqdLTr/wZWdeJN0a7f/3Maa1sqzQOCqAwqGLwX+9c4T
pq0mUk1E204MZibst8LKRMiRfh25PmNMiHZqKzF48VK0uenqKLAPwCpqR2M4p+zMHzLefnefhCe+
um6nsqdF+5S+Xie02mw0qfjg+T7tGkH9549mZHZZlBoTIAcVYdivdeFzEbEfchkND7aFkBlKaJDM
IXDycD+72aFSXQyJAlt+km7bwSHbJI6/0OB5W7OLUqt/dW2UdnfInntR4xzef35riIpv1fQRBHgt
ZHiRa21DwuK1BauXzw9ljGGtsJTrdmGgUWoU8YBYFJDNiHoZy9dW3w/WUvBq6L6yXpgK5pSuXpYI
cVoLt35soiFf0QOz2evLI+hzXhlIAaZCwmQDLIl2w+5Bjmm1/BBa4BLR4e9CJhTxNHJhA/pafu4Z
OxqDMD+53VFdtcGpG4NY2YDJHXO3QUPopM6Wtte+QN7xGHhn7QeOXblzfUB4kG2bTDIaCUw0S7Ow
YsUsuCJhUGr+X48zRau1iBBVQI+5RqbuUfquSQsSyT48Bzo2D7T8bdbwFKN9RQdWLZbrQB744J3h
OH9NBmerzxjBX5pbBaRoLpL9/hNCVBv/QespuFlLF/cpptI9zCIiWf9o6/dwKO6KMlOyTaASFee5
0BqoDhDJoZjR1cucaYVpHGvZAtqEwZjX3T3j/yezXRyFHbEIWu/LeIVIoDZqqGKwCLR3hmAoOIRE
0BpNvzWZQ27JTks1+udGBb14F940zlQVBU63hGJvN2sNMI1TML6sqq8OD/9clLZbZHWDcK5RW+pE
B2tHt/3zhvsG5y6zViLz8YdYWHbaeo7ULFhAiXST9fbVmmqCJurbfPshNlRihs5W7MkB1jVihwT0
H1SZi8X3H0tKAAy1F3bwc/jzbYDf/YWXmPQEDopgMAur2ZqgUNKQ7QvfQ0dPN9MV896Pe/+VMqV8
VlNA0BIYzNNisDtuI6IjwkhOPDLfkdkdCJxHpFOVitBvEIZLkXyk+dSjjYe3OO9+y6JBUY0UPXGx
9T+gRTQgK8b/LrdjYhRbWGd+6LOFjXbLkPetlP0NMufefoiVPe+REutcAmtRNiRrj5EmD6zE2unX
eusNkdye5IsKpCXISOzXA5lRvkRTxbdhSbf+Nw3yJC9g37jrj+WREMZhbisqSTgIUES6Xo/DcG8d
ZsPYE309mLT2SDaJ8mfca2SdycFS0CoCWuc59XPJAAE01lFAZu2esrJvya7Kz+L0mLjgoDmo+AeZ
SCgplZyWxIPALuUk4kob2nxQUpawT3FUwCzZ6aKNyrh6/47scEDhLWHeMumUyBsUDmhH4sSYPUFz
8syeeQrbtmV8siz6PNdGT1iQiRANcPhjPcmlVN/0U/+eN8oryqaZz7Dnf/Hbgs4p37oqqbG19kSD
yQcagMuNSsTztcd97sm5CUa7pJOmUv2k0PtouuBa3h3wk6h+z/q9E2GkOkINQ0vO6HtOpcACxuOC
ZiGeYVCcsR3B2kWKi9ozFXuqqbBVYrekdfKMyQOBFE+MsEDtr81pqOklH8bviVcSxGOJ3zuXHwj4
R3veaoq48gJq1NOac9/Q9Cf9mHLOREweIajiXlsN3pys+k7obV0ulaVXfhvXQ3vfXslGdX6QnK3a
8akSOjBYB4Jbffq4f+z+wx8FQgIbyZ0mb90baZV++PP+rEXEIZuysTkfxaLYaZ/WYvMs+UD7VsYP
7BLOOuh1n2GuLVGFn60Il99CbaTlkFDj/VWvjj+GKf2XKsBOVp59WgrtC2G0QjQGnyrsT2HyvP9b
R6MWq3Wzy46HAJOrOkW2coO5yay6bM5ErBDDnVDFJZHnyBL21zMfGF235/LsRknbBZzNkDgUY/HY
vBvgZ38wvawOLB2bMtjMdd2gd7xRSQOxMp2BRF6L+NA9UelxI359KuSO4/DPBVUOSbT+EGE+UKXD
vIGV339GxRCDpUkTvPLncQu6gE/DZNChfwwX2+FuB4pgxszpdfHI0kRzFP1Ay0WZxExYNzUN0UQS
YjLAhTLc6fqK/W+Eln6olI8PMvPi5BO78HyVZQoez7Tujih5E1xLCZosn9ydW406AE9AK8Y+7MQM
WSoXBwa1Sds4Yp8i9FStrQSWN7pQG9Gij41KBr08YC5jEnflZWyPW6JB3VidmMi4NzIn7KDtI8p5
+D6a4xTgsdeo9/AW3bhB8eq9Fj0Rl67bUK93C5PLSu2BQBFXgCz2iA+rUPvx9Bm/VzWSWeoKd28o
5Ocq+XfwbEL7ZhhvQ6m9+h2w+oiXNrXKnZd1Wb97vV7cT/MOAoa86Ax9p/NZ9aGDpJhGweG6S6Yx
9sONrIdYuhMAyxrAz2X/u/65BoiSYe9Q+JL0dZiUB8DT1unVuFC8k8kZaFZPVF2WWpXpbIRUsCsO
YihmfR0qr4Q81NbagSKijRdzsNRPP+dEIJnBct10CcUIsUOjx2kJY1loFsUXIy8F0ZOMpNqGqRd6
wkhljXDw/1bUWQuzX60ikk4VzCZmXOeLIrO/bRqTYF8qguLPRDwbbfgXkNe193vPB8TUCbv8kLxp
yd5OSBS1W0TwcDWVjLS0ZjcBn91+SrCEjmkXlMEQhgkdsFxBAY5p83XAQsOzSHsLP0P4qxamfu29
c0PuVAxry/rKFSvJgr6dPY+PWAwfNx3v41c3TvbEKWthm/krz+zO+mVIk5iW3KpbwucIwMOyEuhQ
JX7ycDarGN2DlIaqRuy2SN9eiyig1SxyPEFRZ9VYv5fw4iFj3YlU3Ut7FxyuJEWJFTfovyCvxnDV
0suq+pbxeRM13mBYeTXQj5lpll7vM/MOLIZRMwbTOl9e6RuXUtSAMKmnYvM25BQpNcoOb1Efe3mV
1P9xTU1knPpUDjir70B50AeL1iT3As/Vaw4v83MQm9Qe60pj+d0VzmZ5DcJfsobcnAo4T2XCK6Sm
X6R82NVIRQfsEFaen4bCfIXgd8ciGiuBvhF2+1GxKJkHIMTNBBUtOSWQIFTeSiFjqbyvT3nD3Wc5
oUVmq0XsJB8q7Nz/opzHfhzU+TtQZFJr+Y2rnTDPsu6Le+7N+zVj7mcFSj92FTUD62DHMVQe5BEp
tP5d00YyeTOtWszrWmsVUMzhZHr+1UNSZ31V28Z7vHjUgEUHNVCYZlB7fZYgtFBvPcJ4/QYGxekh
kTJlcUUMksbZ41NFSlveZzV2APcFvCmiWcNmJ4EgwfAYL/GM5LtCQcuhU5r31ntxPgoDDDAr9LqA
Qhq5ILpqr5rLm13kqZzNJBCAzSoQMm0K6YQftPjNKiosnB3D7P0KLW1x1AwJWEm29HBOpH9AQbmO
K+SN5ELzL92d7q9pavZdOqlWQ8qNvSR8CY7Hjj+oGjSKzvJw4GCZIpVhVeugnpW806KWy2ZcyBT4
bFPNdRf4W5QCmY0h5+dbGc92caSKpKLoBj9j706senCYv2bhRE6KG0ux2vgVH+aZ8JbdBRQM1GkD
X6+NyGg6BsBhIiaAdvIS+1ln0+CM0HxJggX4linqpaPgUWWuEp14Zwfolao+MmpiA0VIetiST8ud
Zs17eoM4a6NnVjaKoDIvN1q0BN/Q5XV+sc+VwKCHW+Kz6ek6tan0QIA8YmhYFCE+JD4APnTgdyvu
i5EpGTT9nWC3SP3M4z1PsdVwG0Fnca4VBIzs/ZvakOIbwMElpH/Y4bZBi1rkUGBnUzQW6Yfg9vkB
G32v/WBJrvlgYJJdochiAbooTWc6tt+EQZ5LZZbj01Pv2oh5VWeKl88XoLRqehtP1FYoogUmmbUO
JqP46MQptv/4TxSJKkLnhmNjdLB75AgJ91m96O9e0Rkp0VwqEXtMGDQSO1HBa9WpS1ohKLYOu0pq
h8TTnzxjQbcd8PMwI8q3jf9AgTaKQ15/SOHTJGfG+IjX+1Uq1lXpgbBdiqEN3rjJhYQTQwk/aC1f
XTKQTMu6vOGOzorozTWbzmS+8IjqpdNdd3bRcF4GlgtOiiAt3Hkah6vzAbjAXe9JuPY+lgRTAo1c
Oi42A3XOLKiU5lFN6KMBnJevkxmdLeUIPhdZq1cgTZCheHvzm0TnCOZrlwhUXgqr9hDPmDnRhn4u
ack/sPuZQJTcGlW+sFsET1Bg/krXhlHPBSCbEPCxtQFLfs6DH447V3oXkVxp+WwDlAfJ8aDDjh6n
DfkNky8WRfJFJ06+xzYLo2cVUZQSlUwLcHF+XE9HJx6SHlqkLyH6hlMxd9CK5ZfN0GqjDxZJJN1g
fukLN6hdjEw2EdaR9sfTt8XtDV0gpxcb51mKAskpL8cvLadgBfnKTIVs3mUZ13cEVwHhTahQTkp4
AesLM0cXiZYMGYmGGF/gyKDpHMVw6tU8g4O5KgWZBwOtpSGzA7mbdLKRrh21Xsh1nWtwM8TiHHX3
DKLtoMpXkjDfKv7c51XJ7u1Ge2SP/HX98Hok98MpFBfhVz9XZOtOHrzaoFHAgPN2Ex1U4UBaW6VB
Y2ozg6uGRUWSXbTIMS+ZFIyy+nIEEqJz94GcXpblR1bonjRogBwa2hlWp0t7lEAQAWWElRzhS0ys
puuSuZOLOT6QzSJuwIISMBWkpYXEHsURo3Txuen9uCgfj0pnrsrzyHTUdJ6px/LmLJUEsozmZa1C
D+tTQl9WyOMg+n1yybndKwf8TNymBFq1AAhOkFSqGcfhZmRtCsYsB+WnqESU7mAA5bIb9BHwM6n8
zAkc3gLcy1+Kk8X0LXOwY09IJ5K+igIXaEto9cFG7X3tHgdAxitOZsHiVRXqKlkx9lt1e8aA6md5
igQOKeJv5nT8EOTn61EmerapDPvlC69M5gLE2DgAJSHkwzB46lS5vPwoNJsFZMfvGRcJukW5ixuD
OEgYpfznpPs6/llHrLkUrDxk7ADOfp8zLYKO5Tr7IwblQjIZxyVEbA/t8vQxULR3j8rPzkt9h21T
xQ0Kspm6F8putPWrjKkMRvcDvlNvNA6agLV3KmtNv0TdmVOEyEyW/XAVla30Fyj5fPz8PskV5RQ7
DsDv8f2jXoTIsZrbdfuCUcPoUUs/75476ylyR5/RO0tARgKvWIPERD9NH6zDhWoLkhWnYiEB1TAt
J4NVw9nUILtcLFdtvCZwpVnnwB59GrSzRiN9ro6BwU7kgZcDkqrXFu7U0dicZpE92/Q90UPyMZcE
/qbWR9dvpNUwpf43ay/MNflG04035dlixNFhTXahF0+aOTI3spXhUIpH23JdX3rtGVc7DMtZRt6B
OsjXqVjFo+9LZskYt3WSDyzGrDONIjL7io1o0Px0YBNuVxVjvtyp8UYv7imPowahyDLAYAIJBkx6
e5qONlnbldYCExnQzokWcyg/JZoBsPxzHNaiwcf5aKcwlbcR8JTc7ldF9qI4vLSBYEkHfoOrqcJ2
Xl5Rz6MShyaX/mvVJARCeni9nzMAY9H4mhnh3sTQei6cLaL2fX75JPixln3lZrWq3cFbRgXnC630
pX1rysvCjyGJlQgP0Js0xgUVl1nVYZJrLZnjdB9h1GVIAWrI8siHn5dBFix/NvrPDdCoUn8MVWFm
2m067ch1BBhwwa4UcF1zfa9WTeMD003JmoSi7S63cd9/P37rtodeMhpt6CrzXUc6XJCSTp15ZBK9
hRzvlLb1tsR9gpmqVCY+a6f+Jpva0BMCGUl9BaDkrKAWvAYHlPqWmhnnkW51gIt364QdXB1G1FSj
rCnVzLSTRuWDkRH/5oF8ry7HY8nvo9cCUPc2TuZp9iYyZZ1YQf9vWnXMUiStl93vXu77Fi0XSps2
C3GTk8Pg2VUFgPns421LGnMHKD6eOVkDdnmceZEQI1Xq0kcOASri/vpu11xMlicVEkqvhHu7uqWF
X0WVoE6/iTap0XUVOtdHG/mSOeDQXgbiusaUzeCjG9LE45UQXuEWS05kLYrlLFwVRXwpIhj21Ij6
gnsF+/iIY4J65uQ+/r6jtgU5sm4vneEs7+FcBAFuvebfNYMXQ/55oQGghuqKej71RwdmIIlmwLWW
fojFyMqNlLQnljQyj5kf4sbm4AmUhc2/5hjj6UNsLuEMUWwZbAfD3F0CZzZdRCtLfV7zBECYN7um
QRwYNE/oFCGtKFvoHQdRveV/ISUGJFtW16+N1aMdQfyWLw3ptwComlbFw7xhLteCpHVl5urf4fCM
mLT2IWYgVKYADBDfloi2WcgyZX3QO7G6Dms0RZdlw+XDlK/h3lrP0WXXa5LauT8nTreM1bqLqKG0
ZJIw0U1yfqR3ZnZuZ2uv7m7oD8f3MkjimVjATVN/MVbP4ZUj6b6S0mIkq/8DmPD6fkbZsV/uqmIk
wxVArxCNhq8ttRBWYdor5g875bwT/Wjnb/dMbY0UnixFSVwL2NLkB4XqkRlOgZYEFW0fddfrceR8
NJ+2amYHwDI8QlfxQQdVluA8vWDmEtkzqUz+O9/pEOxgGttVdYxs25XzCW+PfUxyBLxKBoJKMfjm
PZ21vauywsisiiHHbHeUU2n0jUX8tQEqvN+WJhjAkxq9xAelkHDs1cpKcC0LLmfXpnZFJrxunV8F
+NNfyNf6d3KpQX968p3/QsBbisXi74Bd9eLEhrhZFiI7tfni8FTHCHrog7BcHE7jzBuKOwzdsofj
3xLTorx7rowANrkgCNL2bp2qYSVUse2xlAYCqxmH64Ig0RgzoewF+mQn6Go9SqzBfB27keOW7HY4
o7G0V3PPIrFe2zw3J7QMox95VsE01BIrQFHXELnH1ZtTH2Y2U7HiDKEU9u1NcB0VpHnbrm6OVwpK
wQ2ZikrHWcpnmEtdKheh/RvKOwYqvCjfnIH0eWDdzBBz3Lnho9vfz9eo2uuQGD1rmnjWT9UriOrH
TTwGBw/tAPbO2/7Fu0XSJFhHSXke1E5fI6wRiO+wW7NM7dIKIL+VyCHeqLOhJCSGQ/LR5ndvn7cl
pRDNcWaH2K3hR+wnoNxH8NCMuC5AjIc5QodSd/lf4RfPUHAXQ26ni7J24jQZOUwKcNOwIaT3fJje
ct8x22ht+xBBANnAfhSBnPRmPZPFFqNZGM5LjY4CnA59hZPj3492PYs1q2L427JkI7C7u0Vpo1Pd
QQGnOoC7sOIGKEGoOAou2fj9fd3/hNfrtxUE0ZVDq+txWqFpcLphW8u/ng4P6PEx2t0v42+ondM3
eqAtYD/hhukUwWcmqdLSsLvGeBrG6JZDxBZ11NVjmVgrWNE07XJhboo8TZe/iArj9p23sY0m+D9F
Y5P6b0RgBlMXi8fEMU8hyG2R8mo15FD715LXS+w9YsGqgXScaAeCwuQuPDjuia1Pg9O+5n9JZZfu
4HI0v5U/ocNLsHQB5g7kQtRCLMSi1suC1HfBxIjl7gFGOijF64Y3Z9SxRitOj0HA+tINltaiTigT
4IZPXHlGrWGpDVeuZSwsEdxMnbieifJUn7PRtEEKQYVjqNLKWHPmSKRdhz7ie+LktDyurdcF34hd
NpB6NS/FfIeWWH61BuEQv1F7p1yWBQWcLP1RHY6EP8rhS69L8kdkQtiL/cnkV/lXpEI8sf2GIQHX
7hi6carq2XCtMmtPavezE3htOAI96q2HZbKKrVY/mCUYrPsCujwv7wfHnDKoIwcL/n79ji3jxFDt
OlmnOf7Z7iF4bqnJOWT7scSUghrlQJQwxtD/GH3vAmRih+RrrmGn6Yk9K+HDwxw8h2LUZSRyJkPB
YyHj5pvdcU7IK6VqujwnIDFVndy0lC7U+Y5I4Yaup8qztb10djwhU4Kq3ISMEOA47dwxF6COKbdR
frS+IHyf71Ir2Q3ErXBPniyxGLYvp8sq5BiSWyA+tZ8LE5srH515AA6rQU3r/1Hvw7wG1PF2BbOx
ce06YvlGocBSrFbL7+qkNOrx3PNg54FRSdto4NBRt8+utgS0gUfqjHeSlJ1EYXl0BLII/RhLvK2N
K9wIgX+xjEhBVIODABi7/ZGEgbIDTdDKc6oevhGslf3bEwMZL55D/TFGZlq67m5YYi+eZ3yXd+k8
p1KzJAd8QcMGnLuZx/iq3trbnWhIiyJozQfNPSwNeUnY8VRUlLA2LOQS4c/drsCwtlg4IMQ4geTQ
5dNoqPTMdr8wx6wJR2rvtnikEEUV36chhISMz49LkdGKCbKf2Gqd6KgT1YAowFXX53xpTqwgXisj
XUfrzGBqDADvB1O5B7DdMtcd/zOqCHKwP9khzR1PLnnymosumAu41VED4RKLfhFG5fTWL2S8dI61
6E42cVzlIzs02GBsPhIgCa4CDeSGSTzurqsWvVITauym6uu4nKhvNjl+MrY5isMwMxRMmTgI8GWQ
U0lihhA9v0L6Z6zSsKagDZ6KVYwvRYVdYg1FtxnCoFuNM8mNkFPQ9a5SQacFTVs0VGAXJkFZLD4n
CsTF3G+KCtOStzCd58MubVaCSvABuEZ3NTdazBUCMXMolJGEWpQYWFpZ7aUwWT0f7IEi+p1Q5QW3
lu+vBytD0vu0ZwD+oGEWsfJ8cwT9v9jADLreWA8dEEUEuHQTRt93goD5gmhA4MtXiFPIez41VPN/
kXbDkxZkBa6TwddMkunzPzXgw7J4PxAwDFDZMoaRF365DIyU4z9NCBR54IAiKR4fY/JBWE+sJbfS
w6n6rXur9ILByigOKgb6PZaHmnff75hqbHFoYR+vEt/OYT8wDREhuV43iqLqavdZUim6s08QplK2
iMWX5RGXUKwagmK1atqs2PIs2sBy9hatWKCF+2/Bx+hUb7JpoFuyHgzzeesVqNQdsBOBZ+pGHrHw
xWzSFFh6Wy8xob9J6AV1nAgeIdx3e1eYPnjT3H0Cr+8oj1gEqKXDq7tXIue+P1Wi9j1ZiVz4GZvY
Q85/it1D3iBJ42BVm/v3EhIay1yiLF8EyjU78PeQUEt34vwiPWTAZg2qVUqYulS9tSvP7nkdq1Qq
nI0JI5BBRxlPSDGWtLbOkd1KOzr77h5gpbbkj7eITiGxgLGBBIHwLKu8B9IyBNmfiO94L4aP/p/Z
mOliQbrfx/vYMn1VfwhT4S+hkr2PnjfwlGzhZ88gKUW8B6K2j9cdKttpr6cIRKD8DHpplRIylZ1p
R4NtO7eKIJ8rMBmmlxAhoiWGV0HDngoWArs+gc6cpNu9Q3WPRIbUZhqr3uXGssrNsTx7oppOl+MY
NQ2zp4YNtwXV6nIbnIYxVxKjkZfqy3/ZGu8FH5ndti1H/8VttpoHVoF0YNlk6F709WWVZI/GZPST
5F92c8MY0IkmeOI8+p+fMjUg5YSma9CvjP10Z+8Ka/mYNNqW51cmzpkZE3uNkwQ9Pqi10yh8E+QE
73qqCGMliixMXCdMTqFUdH4eUvkS11nC00y8waFVbgXKzzWh1dyx+dqJudPEJ+69h8pStuZabLrR
Jl/FLX1EJ4tEpHSQURIoTP/3Es2EMlynPxey6bzSZ9k1uSlbeltZnd7sfz+evXChS9wIJFqDNaKL
VOpp6sHcCyhe7npzMRmmKVFlwl9FfZI5edHa2DLZDNSkVRXh+V5omfwogfc5S27eiLitXaQRTnEt
t6eGGV0riJ4318Rnvcrq9astCjbBFBpMtj37gqZnEL/EjgQOHF2HYQMOLEib9fTB96vHd+DEZqXy
sQ/3TxSmgYlJzyQsRFldT043fZwgTyY6Oa+IPbRNyg4SQBysf6YebPzCbOl4Nl8YbhnEuXdXQ/iS
lJQ9ehWgSNZhey1DP6StTWbEY9ZoXGWwHAn+7mDCSYVPXFmP6Dy9uuzHBj9cuTXsgZH4anwJljL1
UTG/l54E7K0/DwNL9B/U1LhBtPLfpszer11iuGsVK+MuI3hu4Y6/6JAmw6tG4Upb2rWHvmj7DvGk
2fAgPl7Juen46tNgVAaeCcnS22mmgQOwfP5YfZ9lcGuB8RiNO736m/pZL2G8qIcK4XAS1VfsVCuk
071vWjXNT8FgveJXXNEIIHgAM6rPQbNYWqidFhPuD5xi9p4DDLEfpmHivWvlG7cTHv0L7i0Yq6pv
QZqG24jwu2OyIASiyYDOaXZ4zBwKdN3NrHsg0Tj4vfP1rJBXAB6F/9eG2fkdaKfxMzAnZeqcowuC
sdQWRbnqsqv6Li3F+BBSADLw/+2tsWCEAfEnVlUIwXuUXnnoAsENfHhkbTCUFtlsu4cDGO6o34sJ
Gs3pAcM/uaGSqGboUUSiBkNlnZp+cNkH0CQLJZZDUkYSCiy6ee8M1neIm9c2KNH9iE2IfubcL2Fk
xdKEyEP59osRHewTVw76shr6ofVTi8EEmlBeqIKVpbRW4oxKV0yOFaMYPLPfGWa/L6w1WsDWaQIT
WoD8eHxelutSJYeWFV9ba0FYYH5KXd7jtD2RaMhjI3TM6vZr4PjLxjQmVcnVYLkdF0y9hlGCdKiW
A6vYbXaJ/D9MGSXoyRfL1ODieYWLzYfRlLbY5z7XSf6cnkC6D815sjEn2dOEtErzStgA4T7rNiLB
zQrzPyahLEj75r0z2c2c1y6vEx/PqdjLAsZUQj5RgWPiJccD/qFLaSa1fJ663hIAvrOU5OsPxRY2
88/XPxZLpSZVWrq0jfSsmrZfPequi53fh79H7bmj+BwoCwsrG4elyq6VepBFcvLYbRNeteB0Zg9x
P8d0+mHbQswBhU3vFxUrCGc4bfQ1ORlMIwNa6dKziRCEMH8+/vbSG4mMm0AK3WPdafBtSz9JZu7p
xpwSDeaKGvF8EnDDiZeq8lQgBLBzdgB50WHETipv/1yM4RKc1qFhtZEuVXsBlS3ZeqpbO5NxtPmi
Jln3FBKFXZmwf0IWLBXIyf/R262JCY+U22fcjB5npEfx7AkZii1EJnTvtMSmvdgGiMLEN2lLNinZ
egwJZE+cf2wEQWtSWbIh/H7d6HhUwHCyEi2urggpg/AOKPYrW6Su5WA2DX8md3wZDWxmgrue2jVC
P4kuIhCObjhwqOW9HuENPhQgA3LAQ90ARASG5EY54JYlmd5qauZ+MqpRR2xQjzjQnlyGfsp/Ze0H
C6/BpZpr1gHDW/sEJI2kLepNRnNz8PLaVUiSe37JjV4X1Zdz3VO8M4cUTWTwgHbgS5Xp5uddY1TM
xpOg3IVUEhtpD4WKsuhixeEI6a0utFsx9LuaoEPkYnwYf4DhT4VIpf6835W9velfvDngsvhw8tec
PEjM8qb8gKtp3gKvUYUhL8hgczaDKnHNiq5IBaMOlYu8vPhEExbe2MgE/rv/M9fB9ZyjrQkUPC+M
ZfGKN8CiSwDsq59t16z5JHBuhxwqXBhVeg/QWlR02Kn6gZCKCqpWEXF7EI4o1UFOh3CtEi0eMMYm
qwR2vlRpOzr2YVJnOs79usvf+rbj5THc72mUYLEX0tCD1Koy7xzUa2mwxhI1ne6zGtO5TuHrBQrD
+b2N6jdpXNuH+4Z6R//01mvuQwCINPuh6uFlPfDoIRgsEBIQATP6IchwyRJrw2nHoVP3vc6r9+Tn
/+2CNkGKH4WhZIJ4SxH5g628c7Lowt/8JrWF5o4xM+vJLhIVox1A7V+ZCmOiQFmhiMPlJLJ6YzvK
u3SAvFiKI5RNYoO4DoE4TBOL+KtptOFpthv1FU5CDR4e4CwiMpi5c0eGV+2PL2f2A90LCjCk9Ui9
EaXNMVk8BoJNIZhWxFJFFqrt1m1xnQAtsF83yRKCFuipTHKp/rIyQPy4fxicf/vs1sAFfkYIsidb
x7lf/4JmkRe1S589O8+S5pxDatFcIigx6puNcHH+RNHVsofZmrL3r5qghCC/1ZV34e1RNlywo24/
xD3hXzD14ci/aPaZX+HzqzktKu8NadXQJK1FFKWhbgqkBpouYqBT0/bTzESqxR4INN1D6i+tD/Dt
RBnNNRzkeZ7aruVnU7NPFXO14HscAyBbgjJJru0sfeqR1O7Wr/0FdgkdxhOgeNJ+ZSHJ5s0kVsah
R+iCRwXsZLYcZDUVx8H4cBb90rdTOsphIE/Xl6gM09+7TuWFI5O6VI5HF7jhlHrlfuZTKMJGkura
FORdFgMxCLMmkbCY9hTLF1iJynXggpUq50WDMEgJt69v/VJmPxTZWtlywkQZ7o3bT2acVWW1YiKU
vCI3To9hYd0E/NxSyc2yb1ahYtTaQRUUtEKpbSoD/rNiow5naqbEHccCbMt3MPlGXr4IwSWzoNyg
VCjd4KnY/mmwpRZML9EaT2jCuAr5cwaaHEjxd2xEnh50iR5X4OHIn9NPeKX5TruI5i+DIH18BjIc
cM/8e7FifBV6XFA+LKULfgrn1u37Bx5sHu+FXqv/6kIAwHIgEy6maqmNsLgiH2b6lY5oNCEl3mMs
ZRFZZpaUb59vGcdMeEwoh7W2x2bfkZjZdFhk36I5PyfYSIWe2PdTp4XEjNFN+3RZ9nlM+eggLFMq
095gYzoQuMYQdHpkwBuOrKGpVvnpLFcQ2+tfXME9rMbxsyqJ0+pgomhbs27E05wCRoOWc/xATnQ/
NpBeVwYkWsabYr8D4+LiqZWrWJ4yYUPaPQ+68HSXKOVb9JSNTNWiXE5gwEaFIf5C8+uImvl3oVT6
CDy5/7R82JJvgd2OQifGdU1ldbX9/+jBZj0asNpIrCgl0CNACP2BTTkoTnYdwVMm99AabwP05p9w
06CG+GkDMuTOGrLpDelmEudhpSk3yScxUtNrXHvS6pVerGf4xGYS1EXKMyBh8Vrnms67zceqyasA
Sw3KjX5r4hQ0g7bTQHRSzAERbsl9Kt17VLBSj/87lCewjLgnnYZ9bmSPRhqLEv3lGWpPdEZ++MOn
P413xC2wc9b1RZweTQ1KaP5hxFJOeAS+SU1caefNcMAWJ16svCQ/K6JK7M+9ks+87hxA89NrnPON
QIPc9dtnZqZ3AskBXnGNemFeYh5prCak5aALdjk2DD5dWDfFSAXxn4Itnaj3/DNgnFTs/4PHpPIP
LDiM2hi4EDUp+MlRt3jk/a71u3TS/2WOKaFQGGs67+jUdGHbbpWDYJ3/v5UR9a47J81bczC9xfMj
67dBxn0o50UOqVVnxhxGE57WVMN4MK2U5Zs4KyMNi5mL+Z46zEvpt9rQ82y+Nc1vEsjcpZDnNRi1
ZmA2GyWzosKtQi9WNFiQ50RW741p0qbWea67grJeVmaGQtLjrQ3YLRbEXXdk0EGPRgUArdUxNAL9
GQMmb35ngCJc2vC804RuYGE5LoPfMTXm8Af/4vyucuyRDhEMjFkQFRBw0I9p0qqWtRFr3gqKRPiF
qZWu6ga1IzdWPNlyW/9kghMTFzx1ZKmuYR7qDFcZTQV97m9sNg4rhG3EXboWUCJaIQSkfMKpq/d3
aCYW1OAsRmP3knjockGTM6ahx+w2ZB9BxQJb9q74zfXHnRtKARJX6xgn4GVtQV7PfaOSRjDfSHE2
5tOSNYP/ME2+CyUZVcRGYLVks3AXqUdvToKEsnsiKSSwEZVtkXA+k0CDZhczZh3sRck+QSylWAHZ
E9d2aNOh32e7FuOEhjZq0IrsxtzTQAPmOCODXjjO+47S187EnTJN+xWld3a16/S2utXmd2bKsnuZ
3e8GHifHIGJz1nhz+8ryH7Q/SQ+kauGvUF9zbcN19i1plZqZ5GvnCGgPiDRoZ3f0DzLNGyigsHuy
5NIkZQ1ERdjOo3F6PPZV4N5nyRPreMMwzD0Uj0VyPJLB4h/CueL4OfU+EaqyA56UucO2vUq9KbXZ
FtXCTP0SUcqMtf0U8hFTE2LRxS0TDDQSFX9IMtmNaUu/WYcvAMvK62ZJIYWefLTRMRaeSO8UYBFi
G0Sh6hzs7iY0KdmOXjmg6nXOJVd4/pOZYQBtnxujTa3tBK/boIxKz8/mghM8tLd0IkOY4R/cocvD
9x2zT/GUtphOKvCd+L23IfD8C1/JWBbQGwOdHBeQZTe0Q2uQu+ChTWU9ozcsYYEE5HgLJIAhWLqI
ApaZD9cjQY4MfWYJ42JtjBP67ND0cP2fYpvvhUP1orW9XyIHcbVEBxdOGmsPkmsictPhZXIGZMf6
NV7d5QESKbSvH2kMF+kUPu1G0OdxdNt+bahzjdiUtjgO5X10VbMFOJgvRt0RiOuFKUqdISRCmbJH
iK1IjrSt4AKjU6KGwNMXfq0sgJYfMxoYLFofbl/M33XiidZljwH7ywL1JjupoGk1AwKTuG7Na1wq
HkK6+FaOkkMAYGSfyOsAmW/pY3Tr00bP59UGt2X3n82VrEgq8ip1UqSK81O6kcmNgH/YgXZgU3SM
bcP77mw3vOnfKsmrQvXL0YiCTAVM8plt3fe3MAWYgGUacgPCRRQVOaDrqy7A0CAMqA+4GXm8Ipgy
sriD1OGVz0SiCamHF0OpiVvd5Ef3U3tfVj05A1+PUaq4HGnoc8n019+OmBb1B2px+bXJaMltzbHc
N58RheaaGjHwn77zwKFNwMkkY/LVIj/arUHUe4yPi1M1WLWcQKkNoFX7XbTFv0zOcIp/9DZmqNSU
RRf8KUHXTnvx/bMF+OSpVQ0CbvP/GsQr4hInoUbfecGLPG0D+AAwt8ImSJzaWgGv9hukxgbQagE/
Bg353dlY3GvaOhkQBUugqLWcaA4d+DVuRnteeaupeR2L9FpoR7Xc5V6jJQ/AvJLOOVDZysTLDow/
e4MdM5N9kOnaSzmPNrhMITYaH2asLkRuPA7Vu1NehZrEvEPUdV7Y+O7gOE9Fl5lffnc4LZBPzaOb
RKcJaLBxQFugl3/HhJwR44eaa4MArGwdHd3HtGiGj9OIsb8pNL05/P0gFFCtYXLdk4EVpQWUjV0j
rosee19N+O61rWpNdCw1mO9SVvBbUnmJ6I5PCyOx/zB1SGiEBTHpdUv6lAJ33FaXfo9dlohJ+7oY
hnho2KQZaiOuZ6dT4dSTTZHQw3Xu3zTv20tgwQYVDFkUiSE3See/tSdlXduLR05fBs8WpL3IHY/b
BQU94JsthnikPIYIsPULiEqybfkH0t2Uz2u4I2xGKm54okbheFa5Z1xSXAVLMw55ukQSrX1VJ7mz
yfUwFi56qMxLmWq3rI1HereI4PbKXRXBnPLOdAtcswlR+M8XCkf49/hI2Y+812TTsqX9KmmICNWM
TAj7+I3qFH50Mf24daAwZ1JGhaRJJ/IHUlauLxOmwFYi0j5gE6myNYAfr8XZONPN70DebEzpMzm5
GglZBHdjc5BHgthPQwIJhZ8HU+/OKFV6sWAdbSoV99G1ZzrCnus44M3IrTSdaXzyKUdEBiTqI9jJ
Y4MlwyetJEWpjg7lRpkc7wX/ZgHrg74jiMLeuK8/YzfHSuIQSITqO9WRADExkmVhPF2EA57QQeQ7
DKq7w9ue+6fHQDa69GpS0pUil5/rgLI05lzLKo9ePYUN8+P6emQ4Y+XDs3+254fhHPGrsH2lw5fy
ppcqnVw1z7I9Oy0Esg7vXMhUApJjyg2lqshJKoJ2ULPRSWIkBxFEN9Nb++ubpRm9SRlEkGMS1atJ
4Y9jEvhdgU3zhPCV7dbvbA/0RHF6mSWtNM2r5qF4F917UrhIJ4RlCq7wrffdIfGQuv8YuWPVjds3
vdY1fWSJeoJKOCHyPuPKbhOaJJBRDrCT++sZyvv8u1G2VUyf7fY3DSIXU7DTqVKMdPGlCoyQ7tFH
A9NFFfBx8ctpjGqhrKHelZouXYV7v02u+RZexYHwSym7MM0+UseZ0XgzF4WKPbML/DKO2lB08SUm
zgPfw6Y5L+kjWhm6g/GgcCoX0Bs0ygDVwa2vCGIe65kTUDvUpaoSEgNAVss1h6glq//45IxJ9dy0
TaHy5O+HDAE7dvUbzczcrFAMRJIv+ZMDF1wWIi4Oem2y68wLazdy0YPpgPsZPScQNH77eAJ3tQha
PCFVgC4reJPrEkykKSpCbLLTjyhX2NKhMHl8x8+LBg5Av4ahQ1kZqi/2M0K91Notv/vXk2/vBgbr
lPssTumVKGZIVv65lAke5cEyoHzI9F5SjoGmBoqVWec+22AOwNpMzNjj14yHifKXWg+B5WKx9tYG
TYfCXe1McbS5FboFYpn1iaoXwpd2JQSSiYm97Y0gMZYmquNQPvdUNvN17X5c7aTEU09J00uLaIqP
5hRTOxln20hGAreTUhRgwKUwTeiUr2J7i8snT+ueHQ3Zf30MAJ0PC+8+aA8BaFt3OuwDPZv4UNar
UDbZME80HH91fKBAF3yTASzQbSkDTxsBzCNagRFCZSRQrJT9Tq+zpDkbm89cujUT5AZj2UUj69LY
rQtEE8WtS+bBI6ou0Rw/0YdTPRx95Wisy/ZQDYL0cxJ7ek3w6Aqw5iqKlZu5MFS3O+w/i9bwZICW
U1J1VeqhRlQx/hizdDqfZcycXYfdZi/m7BZ94zYpFfo6YFVEvG+334t4MisqVMeQ0nQCcBbsJljz
dAe8aabjRFQs8YBZNID6sm+D2fPBPAmH5XrYCGG/VJHtOD4x6OOJRgj3lAAFwC7nNV/GHVJTagF3
9k0cuLsq5AW0ZyuELzl54GphSsItzSQsPB7Jd5vVDjAtOQC/dDdDO6XQxFDJPS+bGnHFklClNPCN
fNhP1smAB5ZOPZgoh/iiOWlsPh1glqJCcgnuD/PvvQyO/TR7r35zH4lVUqPVVJqWcy/TPSbTWzXU
7x1H99iHP7ENeAzfysw9H6vxkUAFjO7tTRi6ni1WVeuoUOJ2syzms83lfnbcn0+dZmTAFSwy4mPy
SFCYgQt+Af26viID494BtViQCcEd7brpzGHn8+6qIVhOctTy2aMOAwuqHoQA3eVw8rpsegVT1M8b
qS1l+CqxAd8cu0BvIpFPSp6xGHOqzM1t+jTIPsDojqXBkGSPZmMeVTcUPWXHHErhZoud042FiRgk
R0mq1XQtam4s5rOAkxg4RbKBxp/BOSE1bzI8Omi7xpuQeCJGB279Y2ayPqAoDuG+DMEtNqRBOOBf
xIL5VdOQMSrneGDdSvsM3c4eiSu7d5DRff1zMU5wHqfKoDgn1ZXipWvDkjQFmiSuCvytijQl5NVn
8YCCGhTenzB9RAwJvp0wBh6j0013hWiRbzuX1qtaz3IJtVOGxRPmclhPpWaYQrni5rQDB7Q6QWcP
09YlaeWlJQcvaOrOmBasKwDU9tAHb0eDwyg+fJ4P1bPZI/z01pmAbhCxURjDL+2gFcVhAgC0prFB
lscG/IRvnCXd/+EIy/A/kylveG5yrkXQbSmEGWtfWsS9hO3fcdBKPFXO2QjQRx+qtu/TRrrXFPp/
sTPK+iF1Tex4GYyrxHmtkQSk42b5657HL1hj1a14yi4IeTDLZAIqio2jGhgV1CWy837SN+5KJj5a
K8udNavWHtInNX9nj5z2WgrQJQvlxiSqSSU9D0nTEIyUa4s+PqSAV3eZlUxK+RDqszEmfNiXlQQA
dPBmewbcZlHxcERkLvsi8MDc0XUAVQY6LtB+or1oVUI82SbvkzKSZqBM8BUx/NK/lL9rJuQcToY/
yPfU/PRPIj+r32r0CeJ9vvcK0tSYtIT+qclFinAi7dhMpaAH5V+Nnm2lt98VtzJ67I83wF2hSLik
HGHeC9td2BuBYJ/aCTSlNkWC6lUuw+8ggv2QuBok/BT3yzYAfzYVTqx24UxrmwRGCQk6B9BxXSZ7
kVMzV19Gvr2DcHP/cnqPRMTw5Du23evVd5TwWu9KWEQ25ed917MMKocakroW7++zV+XkdmX4rCag
FNyoJQAukoaonjITRLFGgiCHFFjRa19MvZWGILni6n9j0zDivbn4nawXz3hDOni/kQ57shBQ9jb7
w+OhrK/OpfUV4YKNgeWo/a7EHd0G76FwBGNtuiyAECdO2U6nNUZujlR3DomzhT6bN8lSC1v2qvwA
7VRv3hmUG2JIrsIEPLjI6iIi97g7O7N7wPSeq18zw8jLboqcXU8qv7Zfekh7Gl2evDyH7Vpbe0rh
6zREjOMMxuG13tyRx8da3BxWzZDdqs9aA47I+cyunk01wkRfT2XXCyhSg07+kzR2m9TcFmBBGbok
ili+9lSTPMEx3IqMxajoHF9cbHfadwprPS+mEckLnn4043f/gAUXwkGga5doPHBCNmLBlw0OHCXW
Ci9dfx86kEaKm+6O22kncNp00jjpulBvVdORmH2DidPpmBTtSDgUSEiWFLkd4aN4lMzUhJOt6I45
T12A8f+Usmi0Tc8BHd3cF4z1+WoABKaUVqcHlcmX6nCgDAogHsMTUnBDyi0TPC9EF3ckcKb01Tli
lies1Px3Uq1wJ2jhbezotzKNnNwGdpIR5sRPbx4v+hRIMEoBOC+fJdPAGDNjIgs7CVwBz79Jjf3S
rksfWT8HhuyfYfwCNj8D2zgA9ByHqIQrj4XHsJb9SzhvkxDFomlVAkcV+Wz39kpRWhCRxs6eXkjt
V4i2cWPQFJ/x9q0+649ZP9FigbveGo6QVpIxoKpnFva46JY6NUTc6sooRcad8WJQIPJbLt9tTT3b
Slz3wx8tsLYCPuNQlfGEPqhSVwlZAnVDFcoFCcZGIdch4GUjJdohTUZm5I/5tFiBwRHQHBMnzAoc
h1sdSviEpzeVyy/T+u6tUY2Whsy6FNFWMjIXFgmbE7zj2ylUDhaYl7HTnGTFLqVs1KyQCv7/l/7a
miwsPECBKVc564Yv3+3SjDoXKPRTPIGtwU3dcqBqSZ+Rq80n0foxqyki/UrfiJKi4Fz9jhyzfWd4
NL4HRjzW7KADv2s2hvmh6Q5Q9fBTmFpF//2uQKtdy+mdSq3WKyWkdc3/z6K/W4J9FtE24CIOTBIl
VdEtA+p1qOowsGhPE5kT6gPslFXk+0/g9SUl44hJ9alUbSesrJIE36azyeZ86RvDvx0DlikJ8OMP
suoRXcWooRP6GM+yi1jgpbhFwS/HfLqNvS5x6xhRUhnlqNKP3cTV+PKEwCpG774uKl5r28ZY8CYA
CmAfvVFgC+nbYoF2shu0+FhPwD43uROsjAuoZmWIsb4HBgTEWOYo6xCbEPDOL7w2oSPkTaYwr6QS
tF3IKqHNdvLa/fiJKEmPWRBWDvgsGUkmW6dUb7eSDJQB+XYrTjr6bjrA0HshsfacW1U88/NXdce+
zIpFaT2tFlakPrgbM5qkiYxr3ny5N7r6rG9OVSI5vP6tv/QZaNxvq1+swwiRI6ChBRtnLS2yIxr9
k4X/zeQKOtmbZcvLlb5Jg8sCsIyZcAR29eanZraqz00pV9zmihtHjzYG9HqKvGvTzB1yIoEwHm0K
UtMqI1Qc7fsr3kwqwogwDgPkOW7dmd9ZcC6LkrHkATck3O72z+/NyQe1OblAG83opjReHHcYHczf
lcitVVVQlVs0pqbg9EYOC2/xAoXjZ/inrAoUGrOYoX0Xv6mTSwbgYztnjHn5n7R1FbF04jrBoT4M
bkH5nEIh/owFZKfGde+FFWHpWcKgE8tKnH4i64f8cQsTIX2lk6L7dkcAknb48vNkJ/yyTMNeYYM/
rVF6ihfmZ3Wav9Kh9zpvhfkoloks6aaKR1mkx4VhQqM436KbnRMczpB0NG1m8doPX4GXQifuvsk5
trpv4er9VlOZ3/CbFa9gkJmHYPCJ/ytCNktEyqDnxD8SLa37yXAepCRWNDyE+DUMIXNyfl4rR7Do
Q+BxMH5CxSeMzBKtRnJj5YoHMtg+JAeN95Jt5veKR9TBqdgN5PN3gGNRrXazNz9sSHrcyk2gbWN6
fOy/HYHZVaLsxX6khoVEibNYEch7Dz5NLYo9OeQIjonqwx6V2gDi3dqhNgnMT2OKNw8ydqwfq2Xt
Z5bD+MZ3/b7btB4b9Xvf6pCnSqCrWDiv7ogD5zwvGlSQTCXG9tqlyarxv7aVeDAW5v9ckyG8dEb+
NPm8O0NvhrbPmNsE6J/re0AhbXUtuFt7X+k1gcZOEZKXZQESzF+rwFCsIUl6562S2fv/D+Nz9pr0
xpofef47QBZJEcn0HV0ewoFguhCd9jTBtsvFn5j1ipmYToKr248wg4THsJzgzwO2kz9KlewPUhvQ
tnaKBj2jQWp6HCuTq9Rq+zG7ElDCvmd0hXUR/SbiEhH3an7vJQEY65uikzfT2mi1wR0F3iLEfbxF
Z/Gd82nYTeApzPUmsBAC/AsrVRUwDCHVmogG/40WVe6XfLu4bOR80b67iDDI/i5VSgMKBGS0Ozam
QYpVOrbF8Iw7UphGQoiJ2QFnfJUsnvLSMqRQSx8cpWmuvzuruIq7pan/QeUKfRXuKOwWkbiPT7Ta
yRkQca6XxVxj0RjregrMeuT8DNRIOEJ+do//T4FrOBAr+6octlJBctsGW9KyDse7IuukQaTmFeiW
A4SlUBFScoTUVjEHOKPuvr26ZQ9BpNz0Ycrt2SYmPh5HQwVin5ioqvjTFw+HRQIFTbgjKQhs3FNp
6hwrfIm+NSD6rAPeiWvgCbeUvR2IG9JrlHDhdubhGGKnRUPZAbAwHDZAT8b0npFMhYPtlv1Y1rhy
sNspMwkDjTN0Gdga0H6KxsMvxm65xS1e2EcWS87BqP88dRCM1vQkgMxMvWqQx6d6cz8TERZmxKDr
87/oqfDlunEOdc1yoYKzWsKDp/qlzIGPavuit8WjzXNIbrfy4rPGTniFzVXOqe4gbujweHTTCAKA
jIh59i2tasGnjzyiLc5cPCjlHV/nEih5vuSt1ZiVBVPqcopJ+Ktx3CatGbuwvH6OnQNFT3fAdaT9
EDTBdxTwbkqihTaXZFxib0q/tbSGiEGsqWKs7zBtgIdCEVBm3IWIEAFxAat/+yiqYlwCGfz30ptX
Rv+PSqlQeBtzQbm+0iaPtmacbaUnPcvPL9K7UDttXJrOe3vIG556czifZtTFqhpTUsxzybQTt/8W
89NH/TtDrvXkDSj59GcFI6eN2mCdpJ7A8FQ751QotKCcnpkomzazPp4B1Ny0d2zTsYqUfBxCk4LN
K0BU8o6Uh7KITqibiO3QMRr24rV93UICp4iPSlC16cCTzZPifSom+csp3+8H5twvNx1AU6TxPWff
H4DZp3UDYlffkPoGnpET+v/e2brHK5lDmKBtGFDU1kWpNH0L2IP6Fls6ZdeRRNPlEpg9waaDo4Lt
b7ye1hK81axP6fyXIbuWEc/KBFAxCa4LAdbFyZZUOkFGMbtl3JS0gAV8a8lwnBA1C64NJuYnga2V
qKB8sDqg7IwHFZ0CixaOIpPCKCjdHoN9VQjggQfzh19pOlXGQlc0r7/QPoglARYiKG0BT72Jfvsn
TE05tf5VXW7YNNyjmMbI08RBzH6detKxM+//wUkksCD3cOztfvrLB6y4rU2Zy451hOirtvKMzzHE
YXD3febA11XyLU8hk09XH1U5lwyuCE6YL6L7krdnNSxadZpbmAMK/NkDvFSQ+kGCxngPkOa3ADC8
58wVAUDrOAjG50VTBJZdFByAYtS3UN4Hw7yzD4pVXANAr42j1V1+XSN9WbgtqiZCyLxctTgkXAXa
3xC1DS01rRN+FQoqrt4DN4Hhb+5/43nv7tUrXi+scv0Z9VDCJe+cDiWQcp/zk+iAzFxRVSLj5BFj
CwtMTKvIb4JDfnpTA/mmruio92G7jm7Z+OcpBVX9pixLo4La9FqeMRgKckDrKkh5VTCMXGyHjtms
qcjgrNZZ+UlfTSOx1TfGKXyw6bekJedDNlqyRpIUjddXqpilIf7VKeNf2zruoNsCzo9qqGdYsRps
CRdleM12PwdA+SClIriz72P//JmqGQ0cEU/qaejioz/t1x26YwpujPu37rMI6vgopzJUwERfiSCA
lhbPdRc6/OPBaD/gscmUpJdK9UezyIN5Xcoav/zAQdTF2RE2colq4M7QiJAr1fqh4MI3Gv+rvdbR
GvESg+toUIVUQWBIpPYu0jzNtq3QOEp9nMVeQ4JB3VMlYhVxZdUWe7bNt/R6yqTEr6NpvKBIByvt
lETOoKO+ZN2qgEfzlOfU/WfRbpXcQ2C+TYzlukgbr0uXUMO2KwTKNuYLb+MGmfkaMHOcCddNY2HA
L5CiWx6Z3tzmc1LZc7F6umdHD+9Ws08vKGvUNyoggeun6nHnVknVi/hTNlbLLYhdYI+uOxVv8Emg
nAuca8kGdZ4NeWkE5BRmZZeo/Sxa+96jhM0rnwuxT3GXr1TbSL1tnCzBqNRIeJtkyLqqHVqR31Q8
scvhQ/mgTwBuVhH1Wi6az8FYWjFqK6YyI70yhOfA8iUBM2LR2+iQxdCigoQdnQ73KCRS/uMB2h/k
eMvrxikSPwKm5hOe4YZyB7LqCE1AgKajjGcaOK1aF2xURExLRUAjwdGkrTLcfU2Fb4tv1zeXl4S/
yEOP/KE4gQR6OobdycFAnNbqU3IA01GNQnvV2zdwLoUTd561pu0gjdsycHZx3OW318F4pzRq2U7l
59a/Eqs7l+j8sMk0OCv3J5jsr/Fg0OT6QABoCLeURwOHLHyx/zQcn3mv6zUozu131Q62N6mkuai1
CI/olKmeaF9cvYBpJRUxSLwOPmknJMIDhOBn83inpTtiQUvoKuOf0qzwHTZRXj1dBVpHo+jegAVj
Vi6e0Dp+gNaa7HrYbcLVIaBOgvb3rak7UBv7he8ollfIN17MEfXb1PCKofLcsByYLaIMRQLhthEs
imz/w2vCIqIC4VWxu2YZv6Z0cw9H1yL7ZKTPhQhpSiKoye5PACoEPevStx+KOv/x6IwKIoy0xByj
HZbFD/1uvrs+STIx2AOZzFAXUQy45Ok4Rk7gtXiGG054oUAEhZBYenhYOIWHfLWnPW/hJfzPCYJC
7XkBXBbildOKEr5Xdqox3qgq9GiM3ENSXhasW6TheW6Kry60rwDF34iKeRyiVQ44VOnsCEvJcTFp
c8FMrS4aPAajPk6J9Q3VvB22q8KeN5m9vw0UiVE6ePQJZHoXXlI8INEva35e11PlWy1MhylNemNz
t98+ugXmL8rkndTFu91HibauRgeyCWS+GhnzD33YQuYOqJ4H0fZ1ITpNqPj7g5EGGs8xXNhxcPiS
+rOsB/J3R64R5M25Q+1/9BJtPG0mdVOouUvfpc7Ilrl/U0g92ZBz83P4narW79JxHCPq/9p5UbZn
MBG1W0QKIolxMLzkPU8OF4w/7oF2+JEYFncjj6+sXk65g/dU11fA8/4f54J1tW++0UVKcQo6wslE
XwxBmWOjV17GQKy1AZGcHUWMVcugfOgT7MKQgKT1OCpA1pTf9o7lmzxtu0ceRwWR+ArdgKTcAU/I
iUsF1qP0D5mKHTKNb/w3jERYCBFTrkn6txAvf8Q06av83UNvMU/+vWg9NJEhdw2CeABYyD95Z/sI
IaW4CpR7Q4fjxI5OZjJQOGIld54Fgs6kc9fiMzODtOusM8tNqbKRchL5awzVNXVAoUuECDTGorWz
xHKj+CPfjyLm4MFjLcqQSm6otCLGJbPXmJTbRtRlQZizAEQ5tzhfPzGCvsrH2XmrAMbiERW7gPfp
NCR9DLH10R70q8yVli8PG7GSygapoyod2gT2GWvi3ZKUOHSU6OqAq5Gd9EJLY5/rbBoLKUk+TAO+
au5J70iMqD5IO23XxhouQA5qT3sUMGGY16ivAkQuGIBXsnLsSfiRQIeyHFiJ8GGxVW/SCommB/FG
Dht2U5h1fDlh0gJgJOr47VE5340sC8/dHt0UFQgHc2CgGD0z4H4l++g9DXO8fp6Xwj4/YhJluYUc
V55M8lDJ8ZuOBnUkfzyMFwfHGe3URaMRDZIfAtybrqo1lpXfFjO4pUZUL6/NNYCV52vyUDBUjsOM
gOKjaWGKDtFJ82CrhI5zuLGi8/qJnSSNVfvYnXqPihK9z68KHBWjmt7s8imwRTdtAwRa1PCKyZ8/
/It76p8iFm3Jkl6TbxTZkPPpFJ16cBJ/5LOG9z5/N/1+YD9qB4Fw2328KJlXWwdcuS+mhW+2usJb
FlLh/DIuxj8UL3Sh0EZ46SCzDK5TaK7+7kXP4kQL70OmCt/eESU+2djFD3JC3mEX6b+o7TojtF09
4t4yeyxujfVjunh9esBd9sZPV6y5WClCttc+Z1LPG1TvmXipvYzrXT7OafbSXiZHsEeDd3rG+nIE
+l+3NEvdYRkbH5+SNbxIR/Um17hUQNjqNZ0GC13cB+LQvVQHmhL4bw85qqT6uIrbNM5Dcz1GXlzY
igs7AHyaGRw8QCd+mCVusaZd/cXecFVUAtZqF9fFdiYD5MY0VulmqRyTQQEejjeZ67jfXmPWWJWd
54Dt7wnellvrFmqb33dH9kLr6NR0GAFwxn2Uko4lkQqPWitW9kXrllIiWDE4QkVM8E5D4dC0EFk4
9OWt1mSIm8xj35N2nryHvRMw8MzSEBeOw3uasvbyOitpEXKHqh1Wnb/3AZnKJYvxUr5zWvTvmVGN
2krjYRGyYAcJRBB5+YulRRcGKoGKaRZQwfbgkhgTe5RPAJziRrLkTbqf+K7A0zm8MOal5oZ4Vlxm
3KPyKLR/enBM1Qnf27D89trEDD12Rc2ll3uxroQR9kbo05PI6K1GIGUt02pAiN35QVcnqwWYgdY0
A09rKXX9AF5PPbivxnW9C0hqGVPA4w1639s2Vuz2dsK0IkUlhTMmQ99a0FHy7j9ylavXD7sUenUT
7czgPn+M6XaXhcyk4/+6R4WvJjboI2WuWh/kA93EcAAdY8JVqRzKpvBsEj5dzeznQ6UU+wKuRIPv
6IwvFX/3hQTwWlbV2mk5ajBDlgcYB/o3PaPk+s6HraXJbT9bpES3ceIWMc5MN/Wza1vnyKxW3Sek
HUXtn4qpApCQOhvP/DnA1hluy5uGcz4w9pf8/TkcQNzJeK1DWe6EbcfgWyfJLTnPLMeZGLQ0UskQ
7RyQsryBY9xPzV6k34HHbLOqXL78fLFlYd4gHFBvjUTWkKCXAwJ1rjkaeGbP60PySe4gxR1NvWVd
zleqjczqeC35Bfii2NKrqfd/skILjgJuclb4eQtKtv5VigD6DkNRn51Y5kNwKtIRDEsFPmgBzg3K
XfNbUyEaWcICeUo9mCrQxR5XMnUGtBf/d7I8ytZQd4SksSnT61/8o+vsNDIU0saRUoDTcQx1Zlih
aChT5UMkCxqbk8KPjdJYlGDuBwTH0lKj+5Jt9s5vXyiF2uy8DfgF+4LyPnYOPxGo47wP3Nq8rU1L
tWqPq9blQDqNaFmtUpmVSMYF8C0Q4pzqBz7MzPrFfPL9opiwarti1gzSuYKZhFoqJOY7W3Idebpq
PZ46+V6FEB2ww4OJmW1Eg8Y8CU6Gpm/coyMUvoOFO7xsmgG6ePpfz6O+lKxiRiq/cpWzdHcgn5n5
rdSxolrjLtqDVH+f1Xxf2ngdIWBnOqftEMe+axe7z1zGZAQDOVOLqozAdJTzt7dn2oodDinXQqcV
2o3Er4CYu1FtynpjNtKiAAg3/2KjkBOiPAcRF0p4ceX8qCnDLI7EXqCbaLdUpwaN6dORUN594+4B
scjyv7iMbXu+sH3pJ8YPgKCwahmjZiNc7/d8J2vVxzw7K3hKbhKEsmbf17YIOgassc0Z6zmhSTHQ
2/ERxlCFOdMmzQAYnXd+Krz8VnG0G2/49Z0kpAToaaTd8Wsi+jm2mcVCwtR6/Us9qGb4j3eDarSz
VTbhx0Q1B8tHu7mrouJkQT7hRD5OR7HBVEnRwTqpXWJOBdwWSLo0iCwvfcAyoj9KTGTxmQfsKACd
dLlqKNKHyL2vOym2RQkU3WfwO/4StYYoYqCLWvIcFbQG0CGNYKPPwSmClldl+HgBB5YTQt5tOJhD
45lI5PeaDnJ4DCKT5KvHwh71ZplilO/l8kyQVpETaTG4TMrBuZmhmWVXjOssTzQdA/9r/8R0hT2q
a6mXXEZM8AMeYNCVSWqN358WnXIxuAl0hqLVv3v3j0UNNDYLFFXg5xBAzMP+6CCE0Mr7b1c6OP7E
QoIDf0P5ydGcmFWSGBWuuYUeGH00iGTeu7wuO6bby8gYfWn0+ZaHNcII2WePkOF2UDKyx/WNWMXC
U4Du4oXV3kJ8voKr2LLKsGuuFSinSipgGZCVTLVu2hrNb8vK/OqRhYq340NlI/HOwndcQ7hUdn0q
1DLUKBvuJLD0HsqF4a+XMjSM9FKXoXRNIzazVsoobI3Ii9/2wtFi/8p21Mme2ziAEDjd3ThGyf+d
xy2UInnfpSVFmVp5TB3tiRcm8B0f7n5/c4CEvXvfUya3gdzzAhmlGHw8sYK+lh+l4Snxx+hVLtIW
IBlKIJheyWBV9t+lYxefgBYX2fWTH3E9yKx4UIYZ3q47wxFfdlBIcMVq/SD69dMOdov7wsUV+I7f
cCIbwwo1Ml74CoezouRZY1wxHe8w/I2Uk/6cSgkQgMjKUs+tNCVQE6MY/+xSXqjB6k6RQfXM6JNy
5LXPtpIdGlibwTrmwCLd2vPeV2IsjybLwUBoobHWD/Aa9JR2oCj7fytQvt87Vx6/n/7Z7ej72nmE
IDhW4pS7XU/47qeJBminlBonpU3rbmANeDjOoUHeiAyuU2TrA/4AlYI9TVypbXpR9gBEUI0JLyBl
d2ovUNIIJb9SC4ekdnzXvRFVxFCnh8GObaTdQ+i+qD/N+mosQsUM5xXlqLPTJx1lOIsjT20dJWEc
YxKLW43UqgCAHY3PsjPIguaQLwulRT7jsxUwCDN5G7MTOGvjkK/pHdTMYILaEVmez2QhVFBQ4inG
9PK8NNxfU8bsr0foqIAhHBBm8qIawAC5AY31ea2QNnMBM/a8FWh3pCnmeZipL/8/6N4OYJQjPUDd
qkn/mjMcBlX4x7bA4mhM8HdUqotKkgvZjaAmjWSsvG47+Fy7Kf6GGKgm+4EOc/vaMcuD5z8g91gs
RZuGPMn+V0VFOcFs7kW9De4B4U8qQe73ybdHU9tVPHECDdbUxUBtlMeALjfGELxT19YOiQS+Xkqr
EqWuyTFuIiMpXf5aiJVKbUNtR68LtMSq+qcSrptw7Zi7amMKe10pnuWmbRU6+BMyrDwu/d82/Gck
TCF+iYKIW/iLzd39zbx+XHfRY4e2gVOgz7KgWzx4LrFQ/wgGUN72gGNMzZeDl3U2BOsPsaBIyK3p
BIFwFigYwLYMdXuhQUkhZaUf8cMSy7auvof4XVlJf83YvKXXaj8unoO2hS/ij8YQExHEkI3aiqnJ
o10liXk5n+139J4IYBGpMzgk6g/uVkTP0/BhD8Xg9vVRiEG+ZOqS9khMViqgqmeI4v+KYWTHTXte
PTUoUhOZoFTZAaggO6LYqPHd0emn3X+ORgABjneuilogAePSpxtoAK3u4XLHAAWBLWJMlVzBpSed
S6ViJKMt4NpRcJuNR0AE6jQXD3RuqK9hITsqndP9jT9ZvVYMOU6imXDMPfCNFBYU2vuwBVDPBoJd
skSHLLZ5EF6ayLxlioPg4ZRYBvjA7t7RNt9e7QT+Ohd1kXBKdxUeyfbnTL66T5hsRsWT0BN0k4/i
fg1o/Ax2Vx9qbiz370F1CtGd9rjmD3fUFA+/JNIJxbOzfMs0zz99GtrI354S5YIjjf6srvMZLjU9
C9HkTRu1NcTya4Q8aF+c3Gjj9s0jWeRSQRd9uDV0QeXdfcJiP8oKowHqKC12gyYcmyxS8OGS3vFx
+gKOG2Iz+mlsof9heyVcpMolgQ24+mdr6F9VBzt0cpoah+bbCS7jBJogsjyPtoJI2f6N+0A5KoCt
HBZ4LaReuleqn3LkR4jZaLLEER+AZoK7B+QiI+xmhdAgB5WQGCuLuVbf18RRYmfUz87JEKedf+G4
o/PvNKQ9A2T0WLPJ5f+s/dx8reSx0eSeCmfI9l3k6/7K064am9UPKpFc3UWP56XronMRJQIAyVpj
yQpSU4nutpFZwC+jCmg6SdCuQCU69e+XPYhwe6KY7VnxBG0y5vGy+Js2vqfTa+JVv7HXC1vmeodp
QzZ0pXMDWoKeiYpfDfTg+CYCV29w+h9Q8OdIR4z04DC4VIIaXIXLUKd+hdN/it/UeweBH8MXY7bZ
uSlgCN//6UE/hadcBZc67uxJWdH6O0vMfZsNOX8KC+ifUiOZz92o+CnHqt2+IcXQVJfi/ZYXaTT1
JTjzwYBUVb23p/s+2SDFG1/kBUT1pipvLTvppHC/jrm/Ng6CvujVK/c2UlF+faEgQS6YgZAjulUX
6kfNvwizLzIzX24b9RaB7Zgs1LK0qN0r2aTsJpY8bLP6vA0XaulKdXZnn/4eM1YqptSV2pT75dKM
7gMqwZ3ohSyIMa4r0QM2tsjd4Mith91xv4yB+EWryNZ3oCyDNwrZlrqsDtI33aB6vTQYYbChGtff
XaDXFmvjtEXeZacauKmMR2+XE+vzzu6Vo6NjlmgFbB/mL94Ton7NpuvO05xvnI3GwG00egGVz0d9
HNe7mqyvxmGT0IzuRa9Mv/oOMYqWIIDjdgYFxCdcLoxWUUFd2ViphyTa+YGJ+uijAb/ruY3YsWE+
DC3TgnsCcY6c2EM86RiMl/rRc4df8rCp2RUn7dSVq+dPWhYmoSU5sxfiEpzqviM7iHEJXdf8N9gF
6CQlsEn2B2N3PJzWo9MU2V/l8Pg6639VIMJH67KI4cjvCboyfQNEu3MqrwHSDsKxwcn95CrJbeGc
GLDKQhjdDHXvDdh+UULvPYSpSAjyiPNdciroitMbNVjivmEBM7HmvbCTC1SljkdO6RF3bsG4bBYO
mTXIBnUsrRu36FgNcuplDWFb6C0+rP0lWUiwahkbTcvqjsz4k/kKKIIzOVvHyY+tQcaRxEpVO2RC
ZC7DBVOzyTFTbWiSUd1YGX8LmedWHazgG2I3yCxr4+gyK9KXLhtDEzIw8r/1lh7Hdv3jD2hAJ8+o
+K+HL857t6e8o1M2cLTkSitZwHKeL80BVzWaQLUAst/0NT/gn7AhdKMex+SiZNG/u0f4fclC69oA
wHRRJGLicXPRpnzM152TOT1+yt7Jco7BDuLpu8Pn62a5ccIV+JZVcm6Fa5NsOSqC5PaPzSkvO6P5
CjJKbLrwHOgwlm3rHMUi0TyOXwfOxF8iSTFGBxypbq+0sDl+B32r5EjiRqldvZdqxk0+45A3+/cK
MVQcMxMXtfvNJRabaOfhHHWwZ73d3PSzEOQW82wTzme9Vq1qpSPU470FKUSnhG/QYTyp1uQXc5cz
tmzxn9zBVvRmjssKOYCQRvXHJInKN1h9JiAv/hGMrK54+y+JIL9/PtSw0o6lzA1bBh3vkSZk6FJD
M/ZqFBdcyYomVq6pFxQgAxr8EbQ/uzCratvOF94FPzUCYo4N9kvh91X+Dcz4iNoThvtnlHYlT1qW
cW25mWz+3lU6p9ulcuj7fN0qeuAlulyfLgAqmOE4SxqgIuL6YFnLylAUwIO3SxlOxUhxjl+WqKPT
WEf3ZiJokYvDexH1cS1YzEbLwhwiXi077sGaAHMqVFcYU+G2m8vIK0KnbfItW9qRpNRGYeiq4zWl
M5OWZ7jVjg71FHfoAS2Fka1R0NeUNF9IGsQGJmwMKdUHvnLsYGAPW04qdEN0w8uFdKUuUkDBxD9D
q5Ny9M33TXcthZejCC6Mu3/I6JmfrZKgdQV8IZmcTcMGjkR3468bKx92dCMaHfTQWFoo7lOfZitP
X/2S0quf/s2CQmt266ifhBwD2+veQbbsgLiOpnkVAWdWk3Sm7E/fpcq3a/3ycuG+qVIdrTSVUAr6
gVY3oduF9bR9baIhIvE5eRPl9xD6i1qszbN790BbRxn9y7SuNPi311gjFCEcHQ8Hd90YVcz29em7
kJEUYaEn3fkOa0Olyz5gv1TuSQbKKzza2UHuP6f0lFihfMVQ3RXvnj+u0hLjiCgmM34Ba0Cp7ae9
WPcQ/D5xg8urQ1oVVsIrR+MKNFGsz+zQbzj8dVHlH6t6V1ovr6/OK4/mAbvG5uuf7TORvLqLf93a
NvrorfBjT1OQk1i98PpLagE6C85OzjDsbVYWKuUli8rGwEZOwNsalR1vbt6Z1UNrHDPn0M/nVJvq
o++5sFQ94Y2tp+g/cHV9VQagJvN+hny8cWz/34IzO4yVvPzFxsjYWeHZoqIbIUIv40faU7e5MBMo
FjSp2PisyDO0BDBmb5q4s5CTWtSi9Rv2RuKYfEiL+KaPX1nnzz2ts5I71QdNL6mxslxNEj243oz/
IMQr1+qAbLWrMYLOGYVqxSOVwvWgXuDUY+GrPbhJaegIeHPOdcfDwvz9RHClaGWIPWTGkroCQR5/
iBz/AG5+Ao5jlwp+DSFV+NWmghUsZBOLZd785kDdY6zqrMWgcQFar4+KJZ+hufGl6imyVPGOlOMB
DLAX57aMAU+HJwSGwoeXpknazkOSsO9He0acp0sFsn3x3OdF6A1xMMeVR+nCrqOzYTXWiHgtpCCV
us5df130aZA5jIPmMgXlta0YQAugeIXBQp8Oni+OzT+x7KvlMEzi5oVMUjj0y3kvM13pp5PuHSD7
HE4R3+W9xje4yg8n5dCqIsDothuoKU0eBQ2lAkqnLX/5XjHFdhRjPZvB+jsfoWp2w3YtxDcLXfsD
LT8ob976v2JBbfH7KyRy0o5zyLRXYzD6v7/bcZXouQMnjT704Mmp8NFfmOSNI4FGda2Q4EnoKtP7
lTfUyaaMRO3E3Zo1oiHHXz3LCy76ae6ucPuPTedHdzu6653YPuL91o/Xud3FRhcqmV3tLsNip6et
a6bVfYZCE2h+gQvXReSVfEXe+LDJNv9EJsxn7lD+x+xRvCh0/oBoXJKFd2u6hOasEqd3oH0Ae7t9
rInvtgGh5Z9G0VWIYt/ieTyKv7hN4v7hz7WmbIg0k74N45wR6p2ktTW+9QU1Bo8MvBVX1435F7aS
9o02+lkPJ2VMer+VEJ1sjfB5fciBQ7WtQ08nuVqnZZ7GMQCLkCBN4BeWcsERkR5KyOFVhfh9SLMb
3BqGGKPz3M/1XQnF71EmOk65951Joqh+0iAGgeP3wyqLPKp0YI/JTlShT4146+yQJJenYxZwEsif
UOOOjx4rp4gLRHWfvX6n3Ora6K8PXwuciUEce6RpLBFc26+1Aiu1v/HRPQbTMYIg+6zsQAc9WQrA
D6oVe9qSlUrqgpqdPVthL28BkB72eAIPJlbq9Y20TLL3DvLvtSFK24Se3DmH3Qua/PkprCdh6prK
uC5M0BfKZmkfqMkRymOwlKmiPO5Ur7RT/E3z+zMSSKHAlDAOr4yotJg7fdJRlLJU/4CNUURVvdoN
BMjCPPaZ8UqgP0Lx4lG4V8Vgr0DXXFAj1jzP//cIV1vunrez07LyVrpnmJRqxjbLqIQs7zoVsj4g
+Uj42jnwKYniKh/ic8Y9YgtesIgqlj8W3x9cvkOYDZFojb0tqsJVIcYNX5juB3KRtEZCHGWPjf9y
Wsc+Fo1qRDkgHEu34gxXx2Q+jnvhqarIdzxXEclMdzI16m1mH7PtkoYdSuAUuJPVLVpdf98vMEs0
j4SJOlT7HG7DVzD3eLi/j7J60iUbRIcdk5RI1D8hM5aTtCHgn5PUkb+fKvVHoaILd0009xBJNA22
lQ4l2B4N27nNfdZVjnAHNkbwjTYnTvVi9CZDLqn4yJU03K+DDLLtHb57/OtxTwVBNjMdKpSh4rMG
wM7S1LMmfRTc3gTspOCLq1hFgTL+kCBRxAgvq/Gc2AJ+935tlhLqYefnFvUUbdYljOOc0wsl8SOg
Y0btDtSEFEY156U9xpW5jKZ5GX4C7/HEM+hG8n1yDFzEhGjgAEBGnTQJzgJFh00C19uChfIU+I0v
2u8m4MDu1QxiFpIcmS0X48soUW8u5VBcwbtsh8r0ykMOw+JMsKf921vCiB97J5fyWz5047ov7DCX
uPR1j67LtiaSZ/tChBfW/AtwNu/UuL4F2uOZVfokTTVYh92tnY5QsLY4JF/iDl3vlI5K6UUrMa9r
+HLhJyUQBobgmM+9NrDo+zVjbGifdSkZrp+1groBoTQuPyFOesaWjnhyLaJ2bFTef8LeExG9thAc
xfPXwrej7yYZ4UUC49lCnHOj/wNZmBcUaIHzvhNFwm6r0DmwdQUx+aM3zfVBdR9FEI13szxzmMLC
96UVVcrdmJtZDkVeBPHnMWSEntVWDcDc7aBxmsfqaO5O7RkKJ4SZlUfIATXTho6r8+/IeFoIaJHJ
ebAvuulXvT+XmxhNYutPbq5Kcdbv2H60bFEDCtIdUe5Ko0yOGr4VD/6hgoRJGbfABdZdFTkoIsR/
O0SxcmrDnsqkrWxZdcqZotZFe9G1CacmPCDd6/JzERxcom3us5zNGEF5Sd2b11poSg7Y//Zmsg4r
v17AdZKPSnSZN6Zd6bFObuQjr7Hwkcpd8Bx2oxWt/2aHRrD+iS5MuIc0mrvaHfB19w4xz8Ugtwh/
bxUOuBuoRQqpFu7zYBSWah/9ah1SavbVLuxGK1TFSbUnIxoNeZ5uVM9jTIdMhy1Q74gOsq9UIUiB
MnF2gaVy5YkCWYvtvINsU5z+EGTxlC2bZLxratTslwV2O7YBTI5R9LqYKMGgdq1g+BJaYHO4zQ9X
X1Ue7l47loZyZN4nJOdBnS/Dpz7Mxw7ybl+6ONX948oaollKVt8Yt/XI861IW05Ip5+j2TEzUhQc
8CuxV7JhdUHZcgzScMeyvQC4YflFlVTHBkfJCszr7PCTi56YYYGL6RBAuqP/NYFZY5GayoSFO3cM
TGXz/khlAW/FQk7wnSNuiXTGriocIvOQfjHc6vjbZFH5b8Ne6lHgWbBITUh0R/Yf/Nd4IrwwqYmx
0wNoLjFfgnOizUwk1RLsNMoLMAdbZpjmhy3fiU4b6EqoSR58tXnOiQ88bfKnd+YreogrJSr5Fa2q
BUsF2oUxfm+7rlsfxQOYK/ar343BVabrhrk4thr4BNSA3A2KiiaS+GXRadXsWYVDYUs8zXTkhn4Q
uOEaFcTOcU6bwKZDhXSVeICR6tmucxrwu4/bgTpW7+G8BdWlb+f+zvzKEvhh0zsgIQtHDVH95wuo
cjQMwmvHpQJx5T2qf9e7uj7aPIA2sB+UUEs0spqi2TwnRAkmHJh/6HDBi/f24QvaNUPTyZpx/NbC
PUbdZV6E4la0TzZzaV2z/zsubJKqSvTdE1Zd+Kmo3FJmzsLQTpFlGl2LZkv80KGnfP/QGcu++YB5
UVhGev2BOhRenc/5qx055iw+WMz3Lux23lK1w8ttsorMTlFFiAG/L1y699rjbt0juHkoaQvhUNxN
DLLlmXJuDI7abPXOGyluZE6ufufrNuKlX4nPkPkJ7jfY/go/jcRuu9fAzMVefkFaSAM7Dkl4cjVG
7K8D8UgdGmzp/ryAEvW7MpYRpJFNRqj/Sg+wThRB7tuMchfPSx7UoY2hyXhZ3gar/+DzzwrAV6aT
SlgluzODid9EYko2nOGl5dWSfddb61l4qVC1aLi2s7WvEVEgPdLgpRGIyOMdhXFpwqOrF4STB7rP
+A9Dwz7qkcGwoBJjHBVd3RGKxzrjq0e6At8SH/wECjAgGLw4BX8HI4SRdvGNQJ8+DKUfunFMd1Fn
2sVoukGpzhVC5j+zLcQMRhmwT18MpXYy9/5LEhUUgZPCIxXF/A9xTZ1QV4uwWNygjP7Sc0WLXvSh
QZUOIqXDRIJ0gU+18AgDpZjSYBAUCD+evWfR03FspkoWVptIkmMleYzvtKVQ8tPmmZdhF3MMJhy9
4gyqx+HLg1Zg72MFcoEPJRh6uHSbAk7jjcCjFBACRwqKRNFyzd6dUwn4txkhuhjpMu4unoPnu6pY
sIDVRuJjFz7wHNFC61yPQHBRilhWsahufPDwO5zzfwS5CAD8laT8bkAHqDQKnFG7HBT/SUMxgDbG
H/zaoSPXJo4q/gEy/ix1ZwBYFh4yKdgJdsDHhz+6e7PURRxXFrH2cyeWTifQ5n3ANtc9MNCeW/3F
K6JeOGcj0uh0LbNVFyKz8bIQFI3ZHAGZAt19IlngHEeJqsLN4ffy9h2UIJmnUFirvg55HgNXTNqF
tRH4Img/tm/NcUD2IDxuoB7GG6/WONT+P88gnFxDA1MImBDdB/Lel77cQqbJxVryNiKSVEZ6H9YC
hY3nn4bUHpN+Vf9rAlDppf9rSE3aAGjjF4/YTO3jfub8K/tuBI8DmGikgvUtpf9S6TWf+LJ/RG6M
nBkciN7dzRNLMJW9fo7T+yRxZPJJtLyzd48Mc+V9nGIyiHYXxwGNbgQsxDfb/kdYmrQsCkVFF1cK
FKnUexAXBZIdXX6vN4Q+Eb3uOTincpMv8J7Tk2QtiVTRRTjriWWrfREgQ/VpfxrgYcn9NIUx/J12
PxNnG5bb3ZAJmXfxjg899gBUp1eovIdSP/ND6BACziYOziRrj2e5yBgec1p1S3xxuE2evdRM4tEK
wlpBqLFGEWpgaJlJX92wA16m3UnIYtyxCNfh9Yhub/WhgtQQsPzFFP8CcWVljZbmGYQNxb6VaOWL
nkqJr5KGMTXTuzVdQybjRTGRc/B1ESaJXJefhF8GhkigJAlWZGG02rLzjZrvjASv/yYYzRc++/lz
vVWtZSVqhilD5VHbQCBXocIZ4syL6ttqqKO5MX1OH3/xw960mKslgSsiliUmmu+30O+8SEjve/yx
N67vNouH6jFFVuS04XLhgCTWnMowIdaoamp4PgcvnzlrrDvYZIoBrdPImRWR67akY/PquQeLhklh
b1tJ3lnKZaONr7CnEAVLnpTBj8wDzgx220iL/RtKIxPYn26XgQd+YLYgDXUdvBLTkNU7qi0r1Aym
Ku43PzejYHqIJPTKrDoYzWvs9CoOFg2rtv4N1wuQNxPl2LcT8nun6d9PEwguEZxa/uB1Yu18AmeJ
HJJkFFVNB5ohCPsl570B8LcWgnjTM6FWo7syuBO8NKguaTs6rgRW9vuhKQRgZ+xH8j5Bl+wi4StM
xr0FnJ6Jgv2/G47k79jWVvFfOJXo/yDCJMg6RcgOcNTlGWhLrz0tUowv+g2DIxIUv5uMhek8B2Pk
ZAVDDwmbpzk41qCUOeKyl4QAR4tQo6yo2oW35hBdSfERBpxNRFqjtjfOmXen9DoGHpEiIdE8WjMY
tAtauXPU6ql+L5DfuP9xpBCxLzWTYRTD68HD7mfrogUleOt4MznTCvbTC388RQcm57vu0qvmx9DR
5HhIRhpN2GS/sq8EZP4a7zgdZFed6dUq50Xh0x0XWGOD2IQJPys+oSkhEcU0qYd2l1KytvDi1iQW
zoXliyf+xJKGYijdYZLZHvlsBOvz4hTMo33m3NtJJ71J6Z/yYVnRpEw0Vpfvj6cy7OmS/a/xvF1Y
+e+Co/V+spR7bwucsfZ2x6MYpib5TQFpeqYHsUdBoHlp3F679bsM4lYPxteiBm79hUb+i7geTO7q
/XD2EN0crlx5nX1hZsO6gUFBA+7bb+Wncpu0h9j1NckkPXeU3T+1JhDB4Rb4Ig3Bk0fjHBAeSgAT
CYK5l7ahViwgr1zMv9GNbXDBi/HKJTxNU44liGDKOhrjJfUU82LzqVLCmk/HuKTN0TzE3YrMRV6P
ePcoZr5sz5QZsHY81ZdH7nf+6UUAHJR8c7cA+vYwztLiWc9OL5RZppjBpqyr4g9gDTSGupUeG07I
YbIazbS+CpuqaR9oW+oqA1cbv7b5IH+jXBz3BNzxUMrT5qwHRj3m+AkPTgrYWFY2H2tvgaYyNFq9
o9OHFxN9LHWyrd14KfFFkCBDAkZ00OQ9apfzy2IkrOQmoyNTLNxCbQSAO9T5IH77yCvsHIFnN3P4
o1VLcQ85Tmm2vbdCEeFQiv6bcNtHO7n8QoQqu23vicdjPyoKDhFxQBVikocqVXTWXb2sFxklDdhb
g030mCE63clMOyPkNBSrwCRww1N04ZRUIPnlTGYGb386kiKfEPzUSyRNHFOQqcNkADsHWdv1rj/h
tsuQ8cqE0dFMZA8GxThuyHEBqRZudLG1u1NggPoNZ3hEe/zFrhCQaq2SAYM6YL1z9cvz2tSp8TjH
C+kPOOfl2/Acl3J7V7MNEzlLDPAjCOjZaX8XOmSMVDYqbrR24XpX1YPrlBKMLNjn6rCvHmWpP2cB
wk8yb1D4n4c27ZmOAth2X5z8OdhUUNfdFFh+CxZIgRTy75S7ueo5ns9PpYjzUICXPxp1teQhERPr
wfbtZUpWWwo7YfhIaLcNb6DDkAPX8Oeo/JPIC7ZRzn6A34klSc2qjRlxPADNx36slOh7AXPM4Cwc
/rb42YkVR+qF0vlcjy9BWiD+gQ+ZudcFQCE6EyIG5Np408P9aJ+fYH8JxE69H571I++FcJmUxKgp
a8s24g6/VGjTghrniQX8jQaWQNrgUDzzj6SaHf8BddckHKvI97812uXCzfqumslg9t7ngYwER9V1
nqVSp6tFdx9rQGrK6BxG5HS63IzT4wlo/pHL3P+g46mYnuG0Mt0AppgYwvkEyHYJCdPctW6QXIe4
3psmbX4e5mO0mRkQwZjU40FW4AitYo9iOi+HVcUrLnE9Az7hA3kfqiBhEXv/tRX7Lpluj8H/l90I
NYNxp7Mcc74ckddUokpETa4EfuebMs6eDB8ceCI9jL2k7TD2otqEoCEFr+qK48dezRiGGw8cuWFo
WkejGIr4h8mydrzMM+AgJSRnyTUrz6LWwjEM2RPWQsXq7jRJarsFIU56MZosha/EK8s6N861sZeV
lZaeWx7M9Bv8LmNsXNHcdRYHWwxnREn1/xlF6sP1UCQAuFVYTD7BTyPWGTAtAmAuocUbEv77qf4B
VVdHbmuD5tvLYsQ3lCf7Rn8S3KfVPWoekR9BCGOj9sqNgN3jc1Nhfk8wTDItlEkOFtdGbSY7aG2m
VcDV434cSn7zYn5RPLnMLDXyJwCw2dPK+Owdh4+jR6fUEEKTa+7turtroC/opyFleEqVSEs+OXqM
QQrxHJoLx2yvqOypQeALIpOUsW+8cnX0g4vizxeeQu0ftCP2fHr7RZmgRly54CO+UE5i4+zL0Z/7
v05Y0Yv0KBoqPU+Yg5CGjx2/qUTw8Bxg9RZYO/AR0/HhLuGk5UPlfoWyeUM/LCPNrIhuZkbG2rua
9kiwmAI/gw74Lk19wp+1sL7OcdoG3g1t7dSsjeDfStQ8t2IQrheEf0CskbUdwQtEW0GcQDwRqwnk
/ALtX7iC2Tbmjetbatjv82NUWVsJapzd2J7wYVYoiP0ivfDRBclKYvXtXiRGwtO4QgTaHp7I7S7t
cxHt+pmAsgLJtbDN4AYBpI9n6TajAx0v6wJPrqSXjmEOrh8miFrfvQfE5YzLOyEtbJBcs6leeTjO
RtTIlWuDif6HsoXim2yehr0NKF8fotPxs5lmgIb2eVfJ2laIyCv7vzIIJN7wJ5NC+JF5CBPXkX2G
LH5b/mxcGXI+2ydBnZ1Qqk/mqQhZ6xg94XgPBUKPXVGeFMlzNsErWnXtiVGFr9uQLfNBg/iOMtmU
ja4Xgwx9IaSrUMWjx7jHWbqppesDVsthi8gpQMfnCIAPKBJXK9F2S0kV9Xge35u6PfmcCUkd5OQw
l70ykcigB1tAXHYJEeQ6yXZ9gCnS4mIM0OagsZYQzs4uFVkFzMAGUX8XJ7n/w8PxRsqHDAbIxIFV
MmLG1aWBos/CK5V/roilQAzFaqPiVW68eo24vnzcK+PNPXaq9hVGMOkt/omc6oropTUD++9kKQBo
AeKmPnYyJM0D9XprKJ31l2fRjl5mbp8TlOZmS/RYGzaS70hDMTD5vnuFjg4rUehJ//IGFK5UinLk
/ySKTcHGrO3xDPE9uQxrTnfmT/9/1VztkI11FLrI/YLUoA5Scki4tQuAD8k9y9swL0ZlBxjZJoVM
NZw1ZX9FFanU6SscQVvWufQ/LoFGLRVsOXN067DD7lAObvgrEySoyUkysEbPobraZSeujJFRYPEM
ooV/cgOjAGCfRYkacbzsCKLdNG1lfl3Jt1um8SlbaJmXlSimyeYXe5YR3bqP908UHLilLXd+QyVi
eAPfCrrg6B47v2XuQjOJN5CcKn7sfnu71B05YgoBE2vzTZR4FUNVoQ44qm4bvLCxyX8HA0hS3M+R
RLlq5l0IkL/kudnJOfFh8Sk0YVq+P/XYZTcaGb611OGtB56F8mV6nP2f/c1M1Ajgm8QT4bl6brcl
WYefHqULlHrfa3paC5BbaJbHg170oAut8/U5aPT+eTjk2eMx3dLkdkX0x96QmcIjfk4cOo5WIVKV
RKmUB7Hh1hWb3wOTIS8Ecmv0WboGjlebQPVpehBUSiUMYsBzPalZ/S5SKrxvXAFlm2nUB3L2dvbE
Dp+APmeWSzkFMPDRT9SyzSwzso8ElRJYQyd4FZe7pznaLqLIpf6H3LUAa8/j68otAeNYkUBm/XdT
zK8ZM+qo++K2SjB+D8Ltd13pr6ZGoDXWB4Ze0l9z9Hn9RiZGB9a9DubaTVwGqTjj+utAlWlPha7C
iefcd9emqtGGd/6KhJlbLYZmBOSb7td8alzabl6AgWTLHCpwZGMW6MLcu7/7869/IBPjs2aoi/Li
jWXCD/GjcADWmd7EN9EzAujDEf69kkI7zKsVbgClROAQQ00llAGrSaodPaKOew28VGuGPYsOlUXs
znv9cHzpcE057sZIMSHM8eJDYF1RzFSQywUAP4vJ5hNd0ZXTnTwJaNzNaoW0WFnRygRjYgX6K9PT
Ta0vaWBu3tMThzGQ0R7ooGHx6lBBEgXY/nzW8NqFoa4a8DtFxTfKMMRXkyg0EMmTctcdRXyHbAhL
Mf9MWc+28LfD5IR3tDQjztFd6mo6lYQukvQc/WjO08h/lhjV3bBaTs3ImYKsnPQdZIK5DsnLuWhn
ZYnrrJ0KQQ3gtMBybq/MPSP8jATVWUWwZYbg6kViXca1brRevYMVn9ZU9YrD700V2VO3b7XUqyHn
RfpSQGZNSP2oYfyKS8Ji4YByffkVrei4FI5pxYzwlOvclMmAIYcg36zOFheO01+7lO5wPsaWfw5D
d6we9gJRt9xHfupbSAnQ7xjffwOqrDLb3+we+/jI2gVcSAbwBJGXvembVY6AQcsKV4oblucLOVI0
jJvIC8fSqQo6cnjHN+6hsjYAyaKfJyw2MA5dxUaX/qjau62HNTYBY9ZOKaeyLVpcPbkWxBcneUf8
GkzDFDa1DAPwgMWB18WVCIpK1kpTEwTfMw25wonrBSclcEnjNVWltPnsEhVYIvqJxVGJ9fpmpYbQ
mLQRCPqsRFIxlnCh5SFw0qmmKxsOR+BtUqSrEfUuw98BbNXT5cdGNHoYCu1LOa8PVOOlFRyat4qB
fjTW7xUIaCpw+Em1lw1eKqbOSFuWm2t1sOS7nN8+kwrehJLXv3HrZtyCbguZpoRjPAIm6pBl5sRy
3iT+V8/GZ11DwNHMDPao1qL8X4AMASOLS6DjsPkpwQAX8MxMf0CwKiDxsL6kJ90sSvlKGTIUE2Qj
umsqwm53BDQuOpOrgnnnXueN9bOZx0RCK8vSsRx4Kie9zmuCAKq6f7w/GLn+2fbTrBOyDeIlZeO5
rfhVeNDmzQymzIqcV2EXunVhZ5ZTFzATObbyKD4CtMnmqJKhRAFV/6ikzLvXuhl52l+/lh8ohdKb
qjfODpBATgoDD2rAVzHHVpPAKkJXAvRx/xOsd7FEg2bPFRX4DNGvQJs9iTbkuuLGqep7tDCqgI4o
UmR9/yURBt40BNOxYISm0rh5KNJQAJc+D6UEnb4Q+MG/pFwx3864cmsZVvquDLRcPbOKlvuigZjB
1/d5qej1YtttssmLR1tGifRyTvH6vrxRWOOojqj0boOPadMeGP0OoqXR8qQ69tr1Wpw4xrCpgeYV
cBpEG44Xjx6vM5Hf34SGU1cnnZmLcGz2X04fVWKmMgbrzy39RH0A6do7vUJnf529rU2Khl0BOKdf
EphvIFHK2L+YMK0AwFiqz2HuGQLtdOq2VcgiZTq3toqGY+QDCxWL7CPUFCQpDsFQBmUl0uhDuBOb
bcgSemJivaqOlL7zsxW+WSUudnFGhONgJgP2NvifpCx0uvr0tODBgIYVBueNL9xNj6plNm7n+SGe
DnxpX4vlswlDrQDjn1YLOQcgjXGESdNia2V2qvWoovjhy/GcdiANqEE365S8zEISA8mGAwSZfg8+
N4RYjXiW1mIqCH7SnyhReSAdCOoX1rTiKDRjVDwDLBXPoJXjACS49PRDbYEoqX+FmLsmxohqNzsM
qqrVMQDvK4OGcxJw3Z/nfDAhBDEBQDV4yI1nx1rqxjuLCxQ176C6LtvGm/AIscN11MSOplom6Lvv
QpQdnFApr0nAV3ZWBZs5W60DKmcCeyx1exB647S0sV6q3NDRzg7B2ov6EBwMt9oaH7cLPFIg/CgF
q62DLauv2ZhmBMZdF4cOUBGXFPEZjEPY/yifjRMMERc6T02VcErbM71QGSBwVFGXKsPdyrSKe0I+
kGYLB/qQww9F1oBcIlIu6QYG6V4DArJE/508Fm9fzaGKjcQbss4jXytPpE+8kPwawhUMrvuO4053
S1rmmdjVd12tvqrOAOe8N95s3a4g33sH/FCbeSZ8qM9YI+hL2ZrPFRJQtU/zZBhU15KODgG8Lkb5
bxY1i52KLqK6V0CAWKBZ1pFzhLjKNCUMdVZs3LEoCmg6qyk3R6IgNso/knF1B/ZRqwfhfWXXHaib
yX9tee0D7MiDs/SJ9osDaLBkgsPiQxGHl4qJdLAuLZOJeWD+h+6mw4g4h1qwBffcfhQ9TBpHFP1m
n3hl3FSvIaayRyiAo3muFxTUB0KR1hz7qUaX2ci5f/WTEqNW+vJUZkb9oOttLqBMV0/rZM0vwWLW
2UsxkWXRTV2Oz6HpeBP2p4Njt3IFr2yH+9UKCNrCvAT27tQTboYUnj633x8vBVPZ6OSulW09Cyjf
hQIme9Sy30C6tu/Ny2AdFkLbpRNaz9ur/wrvK8EdffRGVx8YDJcyWyPJa/q39JGsjitsYNMqihpr
l46U0HlYwS5Bo076B5HrDGD+FOns4YklX6291AUcSLyjnerSZl8NEjRhXeFo/b8oNBKzY3JrHnIq
rxmP9TSw0c2qUzf5corkjehtWLOkViqXCXcilgsfgv3S2Eq/q1DkL3NtftROpDdqqIM3DjaUVZFx
giJaYAzZEQfz1kZFebLyH3lt/H5/i/RvPzGOvfR77MDYqvxJc0sFMr28lItplYkWBhr2HaMryXBv
ROKLUnKkjOAE87TVyH3/NeGTehMFjZ23Fl0FpP1NOu1E1X9rnEC5sRnjaSb0rG3lPT8rRo2bEmZ4
sOke4ETi+eVWF5gy+qEOtTVSVvmphKQhIIIKiX9cxhs5ykYLvU4CYjfB0osn6tyaRAiGHsZxwDo0
My1q3gvfqTkYXqsOO+pE0gFAtRHoh/y2xr9bBXDt46EH1oMGXxSCQ0GF+I6rFGyrHWwi+mSKOPn4
F7scPgUR+LATi85BlQOQoz4pyOpctq6q+gQkWn6iSXFuRLVxpympeL/mRX5Fpq4bkaRc2NeYE+IQ
KqLwfMVVQLHMtUQ9rR/l0K6Yjj825CyuKY8gHpxAB+dzIhs1ILsQvDxY48xRi7tQi3BJq8wDgQdO
VvMvcpewYD9am7IgZ/IL9e6ZJ3afbXzT/TcjkUtDQ8R3+FVJd/LjqGx1aQrwlR17SpVloPt4IpCD
Kqzdx4StcFtgzOt0g43RSIt1uY/iaQpIWxge3nAG36uHg7rMP+raa9Q2dEJ40LydHELleEwcWT/g
YUkG6ZxiqjmmgMA5maqyRO8HI5SWwwwUFkD2gsrB6ftXd0q52jfa5MLKpi3ngnfc0pNIn1aBG+in
i/p0f71QS1cyELQYlLTt0MTLa3m8IvRDuA1uYn97+4O90R0ajpJGqFunKpTWJfQ36/HzZtU1HNh0
Af1Xium/iEgJhpvksSizrWorOtJv6MmXM8Qkih6vVT2iwfANcA0UNfqoWHP7Gwf3nkByOS7P+MOA
v7ZQE1XV0nv3Knxx1gtNbP68X7Yq1xQgjOARcUOAU9D4ZDGDQfzei9RJ+GTq9juSsEnRtscRzLsn
UJvYcDqS9Mq5U1j8bNd7SaWCYZjpw0vhpdSCw5UhThTCN87+LtmYX+gGtwdEExWuwXbpXrOE9F0u
NZny2L5tk2I1UqzbeZksKJyo3U71LUQxd16P8qYqlm1K+fDghx14IOZ2kusJ0mWvNLar8XIphlJS
e5iXR/8krHt1m/9tlNG2b4oM1I5QVU0WzMvXrwYE0dD7GeqiY3lJydx2ak4qUoy1QGJteuh9ScMU
Q3Du4jI8hMJz/nZtfe1AKYexElxuX/Cv/14popGixAyttXCn78G8WUHcsC0v5x4Ip0nWlk3M2QBa
HYs0mp4toG4xIAHuFKjrwvhZiAR3XebMhTPzDuI3efsAXPzl9g82guavhuT8sTivuQtUm1odg40P
NvVkrd0wPmOt/RqkU1iOg1bX71gb+TBPT9I+upPRuc3m4Rnrd78A8MT3TJTEXjqnbvxn3spitGTZ
w5UYR5eA/epd4s27TkjdXcnyiDn+oKNKfxDmLnhHWjQ9GJCYA/GyoUekWSzOCaUBGm3+B1Xf1iH1
v6Kh9KUriIi4t+FEy6AK7/pQ6ezVcDo+8p8ixGlNR8653dHRmsHLKMC1T0GzNg7cH7+2EngXPv/q
NjvZEw6q0AkMGdeus/gMcLAb5tTEMDd+i4U9vCiQFQ6VFA1XtsaTDNbi9V22CxqUucx4Nd68mU5w
pKDukVnvUrsXQga+lGhulpiJ/6sNJvQE6et/TB5A0XyPQFanNEutq86eEQqcdTdQNb3ZGY+UIbEQ
iSH15lgxd5ih95Yx8LkaEQoJZ6PFBhKpRKvokxkZf1+sMQ2EolR30BTGY9PKrSjNdtAJcKrqmxok
lDGZ9ThUPUE/QGNByKKPquPrMPqx3rAf7isAHUUNILO/obq0gdgZGnqtryDb4nOdiZxiDA/4GEwJ
GcqU50S3YebFiuHrD61Bu35CEq3ePCtQCMPFXwryIVvJpgZBw78hSZEAjT9gJEg4yXpLnhF4u40U
NsP5T7HDhsdRfTm+XZvOffBiG5hgMbqaYbzzQTlKqrLf5XibysYef/bNxV9urerlm59RuX6gqMe6
tEe/OxP1/G728xUnYAGil4Lf2yv+gplFJ8d1xL5T0kKLkpw6PDsxDq59kZl05cqc05Jf6XkRRx+n
5/udm6zis8l/Z/wHBzizG7px9oD9XI/i7qEkb3Bg7i79U3oDVV59XeJEzlyrIr6exp30I7ziaVkI
OlIFNkORk4UuXtgX/ZaLFQsw4cs7cu6/67gEX9rjEmVeY/OVwrEM20+qThtmRwahyyVhFZ+y6P27
nmOUr+6KA7e6OJz5L0EaQj/hBBNNlJGM2pchr4QvKKJcszJWUPPKXbYnXZtCtNEpzdZaignov2XR
fp+i8njP+8gWtlLZwULPW+KeJ/GAvXTapDrslPma0aIy2IyBOcvB0JEvuSnED3ggtJTahaspY1GY
PqNAQXFBV5a3SzEqOElafgzcrKwGW/KB0NHrD8c2P67/m6qW4H3/oni2o4rvgyQS4cYbyrekr0Vt
EblYaLjuer0Yu9LIGdM366GZm+kFg1zdl+ac6ZyvqLIq0MUt1Ut/soyZmgXrBzQs8Arbg/sywv7e
35goSytvSeM4AEdQT6Re1ZjhLu+B2U4uswK9WTVeCx5ThZud+A1nJoWb3jmCxVxxBMIr4+Y3BTHQ
6ZgBAOSrCAKZl1t6bU57kcTfda/mh+0Rh4eXxSUqSZ6AXBA4AomRc2NzIE0yVlsBRZFuj7Zrx/aU
sHez8PVaAM1n4H7yA9FvrbqTIA/kLx7rRwQDRcLNQiUnopY0E3VnHDjRI7S/j+wYVWpiV8gR61rp
IUtkgy6SjwMU6F4Hl/8rrcnq5OX8/5b9WATDFS02MmXzB4C/uKLBMzm42mAfNhXbXSqOfkq3hDa3
vHmvzTzV6sk/iRQF1V953khvRgGF3CDlEKJdmnEFRFhLL2VoW3LJw73UsxP1GCSvx7ZwfxIG2Uy1
wY7bDNKh3+SbSrDRiH1iZFS66/2fkdc6HThd8MArOBn0smk9H2aZtktacYzqMwmGvSeWfQ8JGe5N
8qNP73rnFRk2Z/e07re6Y+VkqhT+Vf1KwlD+Zj4i0H+4RWM69yO9xW+PP2E4CWVXdqnPUzTJM8oX
QUzpn3uavOOZt+N3LO+xs2v7WtOOq4h+0eiDYf7+A/itECXaLWv0yHD/RqmFw7qAGBZ8vn1DxTLt
69ERSIRajxr1t/qa7G5izjQ2uN9MXUF+X8jWZtuV1fvkppeOfZ0oXD+RLaFmhXq0lw2RQ0ZoQRwu
FJyPWEaj9qgbFHiMGCxG7fiGSqlJBa0y/KgWSBfUXAZNk3+BYkzbgh34FdRrH9IRq618cR1nnf2D
C4X4k8Sx4m7HKwHyf8m6SqMccmMXjcye0l6dA7+vr1e6IjhTXjvZFHJaexXiBuIiwakmsebZJzxb
pXqP2xgd+yjaFj4ur7HBRq3dcYFUwGLt6gp7aub5Jv8iSkQ38jxvwHXHBioSLJxabV52iqp58VPS
lcdaJtwzal1XEpt/Rc9yybcjZbbrVm7LItjTu65iVsUi6YdksuDtniHPk9BdEtA6cdvcUbr637+E
CulR7Bz489ZzXfF7P5bMDLTDEuNunHfc0q52ADXnZW/4eWigDlcvuDgVaodCNW+WvhJQiijNZI9D
1b8512R+pE6R8Mq2CPigPW+4NAre62rsrrhjUnph4h1QkN5d6bX/SodPE6fsGB3uhigzNoSD8XaA
K4LtNb27t3HAdx15200X0FYWkEMRoZ3ImWFD+ZQJrjCDXv0YN2Zwg+TnqZfmZcr8WM39+mbBf0Jy
DXHgbvei/PxhnTRRK/xMLbMH6sXiZXo3SB5zVvLvLGH7d/xFp0AOb39IpAvfBO1H4AC8myoKh1wW
LjzN72wIClG9TaXpNERuTIVMS3Rk2vppJ8Sz1dsZ4XYRC/qZspbwnmHcNk/xxK+OKEkUXb63ENuC
QkNZ8bs6rOX3o2d4/sV3t9MGHWswqMP5PDidOvU56xgBp4/w9tS9rtQjKGDLIRevG7cXoUFh4dDw
4f+h5hzFQQKRtMFKf3KqHm9VXQOKgKvc8I4TFV1ZFRzKCqXE570qdIYfSOL00gixwNzONH6FQhTA
MzZXyVAYg3sG/oKPY8AVAmOVN3HvdB1pewNiHaPIKp29jouCVpp5JVmjOiG3bt7QwLRDwmiJm9Fl
V5yVmntO/bQqEyrhlOhj43XdgwxY5Y3XWKzHs7jbo63zUffcq51oaDya88BoxYkW2smgX5xkCTKy
l+5x9Bx6uRQHjq8CgqJw/ut0i2XUebZBiR6zqwo540uB57ShVGe6LA6al2OZk3WkRXOHlXfLyA3j
3nU9OjAYKMRce5F93sNLn6H423LZaz+y98oZf0LtH0Ae6oJzc/YkORb5WxxD9vOtLfY8AAqDUkU6
eYutY4JRe5ayQnCi/JOSnVtGLPpl4NaEzF9EhVI8tRPTv6+S/ueEuPUF/J6mxUH9Jor/0cXsjTcD
d+Y3Tpp1ZqyU076xQntScxNU+Wbx4pTS5XwVPfOydRI4peWreHBY7wIfgSX0Pggf5KcJAzwwNN9P
bpiR7m+D54MYQWWxnwNtoCE4+JYO2pbj043nQWLkEjLfQAkH9AySJ6cXTGK682LlaGKyIMb1fVBX
kYA8XPK1t8HmKylE1P2w35SYvrLVdEQ3QOkdhAL2xjlukZvYkQj5FHypd+6GVgx5gVTyfvfG4svg
R+0s9GPLGMvMYZ/MzmyZ8anihaT0DcZ3c1+I8XsvwnRVk0Vi70Q0EBocFszOc1vE2Bk25TvqWN9E
NdkTP7q9oMa7b6G328jTc54iStc0sw5fLfweH0rnDJlsKDV+No414KbT/1wA0axQX3j86l6+irJA
b41PjYzZDWKWypxk5TE29Dx4UbhaSYvswheis1qXcW45TvmodYOq94Y6N0j2+qZo/bHtLo64Oxxe
wSZTZcFwHDKJghZE/oKytGuCAwTYiQpCY5AapO829OKBrghORopDuuiK4KLZg+39verCNDy+0EM0
Ynpt/nUNvnzl6451ux8ZBjPGAL6wAWT+DyuWKaocw3tYyUxLstPSF8uzzbURuOrEP1hxsMnrXDVM
KQKK4/o9rvJH3R0mdtZTqhcjDK/ENK8+UxffElNunXs62JDM/nX016W8PKrrpcmVNTeFHZvQ6O/B
vh66jNV7JtYUxVeCvzOB4BBxWdfKo0zh4ttYLdgU2er+9ty3j9EH3VkE4UkrAwatpzvJAjiCrNJK
kBI65CyxMx0UkTuwdXAUSxTympnZkl9zAr/DZ6bBK3LbSELGTEEssj4wChQQwC6yNPisowHnxSAz
8UgbUejdXp50y3gTRzhyHNwAteKrlWFIJuS1XQLugOIq7znD4d2qwn2sNcp+kMMNAl5bP1Uup4AR
Y0v1Uj67cD4iDjX/JfjpOVPKmWSjLJQU2Gda9ZOVcF3TPMpkSmJwLe3R2TvVt8jckwsCYX4VEZ+1
hUcEjykxYMCaMtgxrnWx6Vj/IR+dDPkUkeFJbW/on4E+5R1XGNbLe0O2ON74XMYP0olhoyrfm8tm
WrY4/O6LzPdHCxhzq/T9x804JPCbBx3WXvRguh69hJIJkcMNCIpmC3VX/aJwIfzfUkMv9/5IEd5X
WG0Dcd5uZvlo3DmtSchphMg+YB/bcFgGYnVdEOGxY7KHsYHVzkHx1dANyVyevM1Y044iuoSONTzB
soPmbazOUAuhK404z8jjZQJaP8+FlZ3uEvGZjzFy24DNfsDAOVN/vUN6KuFAu1w0Jy3GLslZo+jZ
I2ttnR9omp+/1KKYGTZiOkWtaE+AAU88dfwHdjbtS4IMKjnnN16d8O9SIHt/gz81Jt8pk1IX2FOx
FYdeA4hGse4OI1RinXPTyoZYvdRy5oT7QC+J48uq5vfdHzJk8Tl24zUMfM2kcsw3gkvNT86TE3UC
pogRZ27shgvPoC4EcYr+NCVt6B6XgnfAKI7GBmeVwhyyAkJruQZ5P2s7I0O9A+YoNvppSgh+6n8/
7kxJIeY9aEqNqQ8Bm5Ka7eqn9BTEV3GXh/k7sCQmYohScbza8MVMd03bMytwF6g9Ah/XVmfHZ54L
m/NJuZBoQY2qhgS3OKZARqybKQPqL+/bW/jSEbWbrVQAjZ5uJ0RpN6b0nWXGtHEB4e7TTLvRjIHe
4lKqGCkL13EfaHzRrgN0dbtKrse8ZdN8DuDMqlEPeSdrwpYVVORjh++ifHq1qCVgzXsm68Yau2+k
D5yZ/5KIRLGPGLX/al6QA6bkEgtOif2AczdvxksFQFRuB5yN7WXt26BiWB8qGCQwIZnJNUm+wyZi
oTvOnB2TXqGpn1NuRYVtLXeg3azbc6zLMzOY0MgA+UGYcpOdj5FTOHHeZAa5J3Njv+sIMPrv+0pQ
uS3mmq1uHhWEZ+rQrNsnK24YNCe2b4rO1b+G1cRZnjPjusZTHwcnaTwHdZc94tYpRYCuxY4UBwe+
1RV0Ets6NWSAH4BbF/hs19aW6SClPfc9wiiZ9eWg5bpeznG8WUZ90S9v3LnhWyRZ+AJCxvHE1Lwq
hzwjf+PTgSSZUPKCrw2JNeUH0n7dehOs/ee46Xb1TyVpBQ1v1eLgBTllYCMmqhAvC0fs/tU5iuts
TlQojuI18xMgBgvUDFNE3n1PATg3DZD8q7jCOCZhMc3yyYm8DgZLSR9o42Nr+xQ4kf9wJeVAPXqI
DjXD4LXuAz3cpCYxG7QkC2V81QJRxffW2K6nmBRlHfEcRQTbMEJDOg7SeQ/uM0sXdnteAFAPWN+U
L9agG8bEQIAbNk2diDUu36EmgplvDkuIpT8+44CxmnTJZ9VgmHN3/7Lh2SVdUs5sm57T42BZ5TR2
J6itflzlJO8P7DIWZZMWW2yZEHIC8vieLS65p9JaBSmkd/c1y+OpUcrSfSZUGcfBOhSHOArLHW3i
q/ua7xB/5PIskdg3an6ULW2W4lSv0o7bxCnSfGMrfBmdiy+9GFSUgFowJWYM6SU5orpLWdJCQtcJ
IxPNvQhgc9h4Kcx5xTfUBF48O5RRq303cJbmfRvKcOtYDqo9W/z6CBQSkWjbSp+pYg0Tzo5gnlj8
LXa8Uxbe/0Utj4suhY+B8otrP3QVCM1b465rBylR+CF4PphZMQfzFrKWYh0eKKhBLGiEbqCiP1O4
I1ZVqAVkj25lfEi5jRjg+2wnEOYyKZF9URLVnABCbx3jfBHgnRpaSwUFPqjoOM2RTPLpcDQhJuWk
WrYTJcF8l9Fr0ULS8EFvMyYm01doY/RCScmR6G44L3n4ttGujza+TjdRYpmc9RfqaBuuqrf8nyvG
e8E8ukkwMwc+yAKLUwqN1dSVGi2p6Zsmd6vk2bbyfy2qb7XbXX6DSX2LDisTOzR4eWjlmi1fjVF8
rOcnipOgBUvnzl/27zHAeFaQv32rP7NwZp7jWhleirKFujB5jXstVoZdwKZWW7i4ZHKPrVqqHCoA
HSs5Sqxrw/hki4Ahfs25f3NHM1TbrZ7CsES4O4VqLbE+gA2mjTybskNIpPYvYntl1uYibraXWQRG
keY7kREwoDuAb8nI+mlImj8slzw+gQX3LDBQZ9ehAHYEphzf13XeFh4luy6wJbEauvYMqaGaqAG1
dTpbCC8XLOPpuZI4+rr5ccF0ZfZxLp2Z+huhkE37t+nIgUaKriCLjRvsUiwzXAQL8nsRg1BMtN4K
HXgo0/fieC0hK1IQcOgWec76zyFGd8iryjHMYTvY+IVn/3AHsT8sqJ4HS7rct6NT8ae/7OZVJDrz
Q68G2x5etEx6OCa5ZWIRi9aYpwBiy/o8Nhmmn1+NbKNzd0HFvWkYfNEzg75SBY7ITcGY6GfdYtkm
zwhnRnwkyyIIIDo6Kgyb8gSdkFUeE+ZLbOrjG4iLEQfxJ3ZO4taYvx8M9rgc8Rvh8TbRkUF2MqZE
XOH2bbMNmextZNTTKS6at0AOwd8Y4CKDanB5MFMjotA3whTdNRZKoTO1Saq5KSxqE1QN1ne+w3H1
N4JkTkaMEonLs0PMrcZhCwLbmw9+2oaFU7YHAtw9FqvGYU0sVnwlCht57u9Fesp7tZZ3S8XZMsVl
5b58tCIR7Epiu7VDJo1W9bI1sGlgQ6KUichA4L9RdgUf1MOnYs8iw5XxWiMgD5v889n+5KtJ7KXr
PlX+2MUqOaPNVbfmU8rBdKlIzpbrL8IDMtmXcn7m3gn4HCMClXyZiGuBS3j446Rp0K4VITkG7z4E
GbB8/aEs4YJuxZ6vXPvnyGjrt0jbh8+jJBO0SPbLPqiej8MbHR4PHL+1iOVjgmTFn2c/eIi3ASev
Vy35sXNerE48gzqAFcn06C1kCOaofJe6wymO3Ic9o5MwBSK4d2i4RJTq4Nm88uNyUVDizWOwmUoE
NJtGyE9gcQU4VsmGtxghKtXvLw55VC97N8TfmwX6zJHKgbtpoN5aiUKu1DcGV+h7xLlu18gXymLs
klx805Wg0QCuDt/h1fm7pOIHavT1NHquFcKlBG3H+hC7abAZUct+FlSZeJgXSMYy9/llG92W0uI9
N3bXQ5PJ0lpri9f/uGvQauFKBFy0Ksh7Pb3JAc0bMBIb1mXuDuD5L41hrrrnwIN7ra5VCvw9Mnya
vLel+R9roo1peaebrYE66TRaErl+JRA4dcc3ta56Cnwl95Dz5JPnpqiZ+hCPL5FRIcTepmn8iY+9
2dzJHdHJTaQzXdyN5J6IQB5xgAsNmkl7kkeoQrgDxQSutz2bBB1dUc+P7LbiZxivxc0v8Tte+q1i
I6IWqiDq8EvIFhO5B2UfLlg4oXjzdIB+1jDSvyHAc0YqsZW7out7ZZf4LIecLMzkllSTflEHedTM
wGzZaOswUcICm/s2TtWzdtHZ5ieClGAGbkRIzm/rL1cPX9I25RW5M5hZIpKqfPVJBLG9usjvyxAa
4Sj97lgrnXPS1xZFei1r/N8NIHcpNvNFT8cn8Tn9QOYfjI/pzVFO9farkkqbIam36kWyrG4JnNg1
GkRAvEuY8OALozpjz7wW8NOl3yZEOCCJdr7nwdD/FyiZeeE+ij+aLtY5p5spaqwpL/bbr8J3hs1e
fftTirCF5TWF7RxGiPRSY+bdcR1lumFJYOeLfrimwqT8n1aVdTbOugMjLmNWWGdU+GI9Q/HPPQkw
Ut53A2w/SES2hT+dgITFxwhf6BSlHyCbZBLnZWGbvLB8ph4ZPRybaLLelrf+WPfXund9oHi3cKpK
t/lvPaJhGwjZFKhv9wxoMQy5n1QO0z634XT+vHxNvAsUaffWGyM6CLtg/MlPBUPOUTJPti11doV+
KqAGwadvwUQHZzcUR1k5+rQYxGsdP7LXPObySCzgMy2CdLxIxFHflKJOOxLwTmc9ujBSoXodUw+3
93e4mkPwlKWA03jeZ5z7KEUE56/ccrE18x0nq9MuYRh4LpQYZ6hgUFcZ86MmQjLC95NxrObaoZsn
+dNhRxwKoUGAcXN28I6Z4LGlT5uu4piixltksqV7ooPvmyA/3g78zwiI1CAoUM5DtLtcG5Fjg9s2
zwMxyjua42yCAlDwt8u5rMFl/YCugbiKoAkhLV3VxKNLCX1GCJW616RBSAA0tP2XZ+jPuQUX5aJ3
EKgouo1WJ2mivBNNig5fbxW/mwKRdWZRllqZ2Ty74vlYfHQbkUGXwHAsryxbTJqwtA5/X4tU+xMH
3QCyvT6qHhrKL38esCKQcM11oQ9FXEsR4Reb3FEgNCn24Joab9JNCn5BJPnjYIdbDVrr83o8FOCH
wPj7JFwtzgFzr9aPqtocrZgoiCSXFnT6k5tp0xucdKiXdfJ26LDM61la6+qtIjbGyC8APjUZYj+O
H2ZkvUsMqIlPaQW2cNf7E/ULQGlajvhIk2fOsoElksVwlEOS/KLtw0/ET+1HHzbwxQlONzm6RzSs
cHT3jRtSmsNOu1mQAyD/TAZFBS0AmY5qLpIlp7JFQ0jL9BXcG11pTCmJ/afutp1B7JKdfR9ZZHIQ
smo8ym8kncOXWKNederil3OELwY41/3n4Nu0M2Xs/0w9hkruCzVa3k5iPP97c+dwPZ4LiboUEksl
i6b1zrZJfgtKG33PxXWtN+EMlTjAK/+q1Zv0QgABh6HMCbBc12C01dVGsPLWZaEZtkrzjM4ObT34
ywcb1Q4ebDhf8XnZqmD2AxZJIPqx28BbUZaE0ZU8wjefhGjkivvJx/5WuqR78l6Mt6w88IgqVKTu
CgipbDKQu+5st9I/KQIc7sDd1fIS/zDuf/Jp04KsCgZlgEnZueziVLi196AQcM08bvbHMSppJ+YI
G8fxmAEeOIPI5sOCp6uIecgvBPFf/VUWutuOQoZJWZzd+61VPFs0OAwEChS4qtQBo3yCUtHXYtX0
4DnELwysKg/eEaTAxLGNY5sxWFXnZdfe1aPS5gIzSmMvvlRr3wujODrdqTiHnIJNIY43cezLqlTm
2Nxwnf2y+b1ejNAEGauS4P3wqQ2VgPygCUjBU+ot6A170g7HEPy6h3Az5znygxdWjqA5AzbIApfJ
R1Qus6povAgQjx69xXQi4O/NDFR3Ro18c9VhYbRHfZMKfED8HCdjVSfCJAKIw2FuluKYvxgf/dKp
6KIIP9jC2m40iBLflPVPV2QzOuDxR6rxR1kLcOccMXm7SyPmoH6RekTF+al+vgBcPUHnRoLv8YJo
uRsuuVXbdCoPamhC1vsl4N55aUawWWr6V69PVHo75km9yVBCInSDL1GC/BWauqxUt2qwrIvDE3nZ
oed4WsoZFDNpnQZ58qL4JqixQWvp5Rjp3EBddp4xkgck+PQERhQqSkes6hkDdPHw3j5nsqfZWF0W
uUDtHzvIs4l3Z3LjnRMMnSurn+U5oTWv5nH02gkqL9fVGD3Q9TFBmG+NW4YvzpmtfE4MLlUHG6Ao
AFvSF2nvGnY3M+Jwfb8eCZ86Y9W+zwbKqKebONxhzWAatCBCCedt1FPCkgNq4CKKzuxyZjQmYwM8
36UHlfTFPIKZB+i8XWPEEh3GF5GuhZdajTAk1VgZZbzsVKz5ThP6+u/Bfi7gL6GZBchvueAAviqx
wxNsbryki9NIysXRrb7khVCpTx/jUtkkHyk/RugEPj02QDoX2KQPSAiGcX8wK2YQZP5pZp9r8FBa
cPPEl9thwlxNHDrb8yLAKUpCecOCmq2gDdMcg5uhWcR2/kbirYYNiyS3JKz3JWR6Magk4zQ/HoGg
YxRbFnKDuwwUjF3hUOkx+uJVSIhJb62MV39nxS3gRR9yOB7P/LPan4cij1ve+BhqKjizR1hq0oma
/8dEE3XUkyXtSHgT3yc98HlOlZ8fExFZvPtvTAwdKD7zirHuv4vYeyC1uiVSXcl2CNGfiuLmmjv2
LlEf1FadUOr1CRKqMOeStPVhFM778R8sFjI4tvqG5I9DFmXlIdRuxvMIqKATfxdQTgQcV4xbe71L
A4GsyevQawmTYccD+8ZUBEdDHi4Fjv9IQhr6svKAApdnMvybIind6YaaHr1cjPdgfgkrR9EuW03Y
3q5SX+yCGbC0OGSkgKsUBpfiCRiAbNyqTWRASGV7a5bsUcRAmeCA+/dd2PSTHyEmuMJNPvOhAHzL
rtc5JxsEFGeKTdlsn/cDKFyxIlOOqlRgNkRqb8fghFqV6Bu7XpddmtrwRp6wyO2EMrfmuGBDGW6o
yEmzkwxPoTdoEtsg/oQmZkuwOoOYQFTOQdPn7hGzwLpZ7XndToyuUeLBSkw7Qwt0GZOWvnjjdRDu
vvUzbs3QEh95KkdDie9dfgecWVV/txLbWGIR97jFWki2Bn1tiEFBHixJmAW6IrLumvnvHkXm8FPw
EwgnGJpKBDs4/MzYMN5T6a/mfJNke6WUmziujxmWUqQ3GJRoyjKY7kddZS161BhaJhwKTBbOCa92
GL2DkUDGruw2bbgllP8yYC6/Q/U3LHKeAMxVb/HNINGg2Fkiu3qRKFWfXk+Yp5rjnSfaxODe0Sqj
wcbBBnc6yedktSiwSJlDAwilZlz9TZiUH7RXPGT7AbAlCPL8fZlMaZKycOv1UJBqh3JHa4c5on6z
vkYWAvXpijI0QkiXgxBW3dqGa4INqmxQGoSgCJ31K8/KDhvDFknLczoArW46+BItgpYLDgFbKRmJ
ukSSeQvPjn16YAxR256QUNH9f7TYOi6H2I0tOHgnkw+sxG4z9bFdy3KeKHnrjoaKMRxBrV24h9q8
kIUy9E6/qGYrTH6RdsdVWahCSZ0qhjIFjdP3aAArYxUDJrBbEwxUJfgnWi8qkdfcD7LeFwcdmlJK
lusj/Qz2pPHymDhRlq+yy/pEk6mlKPkfQ3WGmUkAMjHgjQfK5tm7eB73VPvWEu/kdImsG0LxjmrV
dOqjqzw+v4CRpu8jWlRekwcfG9z6/oNWfelWCzvbvy0zYXCcc0CX7zBpJzKCxmutgL0o2YoCHU8Y
JBbtst2sViQkHq6mqsHm8eLVw/ZEXRUN2ojXOsO8+7hqCypSm9sp/pUS4Ywn7ZzLt/VeT52jKeYA
r40RbrkK3JqcaDCkiBY1egUrz8cdW9o5fEyTZpiZb33/QH53HO6BBghzIzgkOkp8B23NNE+j2clL
XxCGzI/8t0ajUsE8VtYWRPqHn3wl3ChKZK/7HJJ9F3fSvwBMdX80QjWLoiHrDGCyKTH4kcCL5Z3v
6USPJgZUCfHPRAqAvQMPyRGWFdN2cRYgz8+YMcAg7E3QTxQmDClYTf7RBQHsId/kRoqXSjU3CNO3
QlNZxJUW0jaF/tdnYOkKOjqN2eIXARjtQkmcXHu/FP506V/oJi6bEgEAwfa2D/k5cMZlDUGdFNy6
jAnUBZC3E/afkdiWqGPboLcxuAl9uMmbQr+ravJ03FyxILRmR9tdeYR3Nc1/Ani6f84GN/2h1eCT
QwPar4haGW0UvmJO65du3OsBrPgLvw1uUcRvqkqgOuA0fd51wXWSaLCrmj35xagNXZt2G4ga8Xmn
wvslJFb1SloOJxzAd+JJlRp1zaJgBZNxiMyI/ToS216tDYD6V2ZpwqTQQA6Y7D6saBar5kGKVoEy
TYbudXgJNs32EFm783x6Kj2h/PNSjI0D2aPWdr5SiBTf/07SyN7+T96pkTLxm6ob4lWDXK6VTq/n
I3Pv/1xHP8cnimae2Wm70NQw1FC5Qi45+KxhR3Fb21FCdhHveKj7SFVNkezBldGGuP6ytA4cNIwd
NKGOco8LLVSXFvwKVsM87alPkKPL65ICcgnlNhmiqXzAVOEcqt3R/gbZwI4WCc7OmzoZ1wf/25Hs
mWTOQFJcWHtqQCeVDB9PdfyXSzk6kbJZzLzWZNhM8UgWlj4gqzmyFu4xak/ibwz8jx0dhnIkzHZb
T7zFYRZjFmKYyVZcmJy7eja/+SftXgDyBmRbqvVTHTICUyJFuo+TuqpdyQ+YA1lWiU9A1a3TCN5J
RkuHsojSMNk19vfv2lR62VnhNlumH62t+TVXRY7+yVpxWQMcmbQCH0043lflAK3H2FQ6MGYwmGx+
0xoe/qeZahK5ZBkRcgsLfYgwE66VkAAublumhBIj0ztOZ1uYCj3j8V/8lrrSxIRdx/CVv+VrD65p
mLzxbN9QXeIscjGZQ1YEJfpjz4jL9iWno6SJG6LiJlSmH2725/dJ+6t50duqeERRKYfvxlLVt9dR
L10ZgXSlSAMRdL6ZJFg2dXKuSsUk9NSb+1GCiayvE4edf3RAr07WtxyVRIDzRuhjI6iFTsnuNKlH
Aa67TqqO8unT8PKMbQBBYVvv+bH5y7dDoNdJINXfUdZhVscuwf+q4nL23IDL3pdXoPorzwAlLGe+
740YPNzB0ejZTsfI6/iVgW1xlqt3CY4uHjRDDgs04+yHpwqwhM22A3vrkTlJrGrqZAq9LPtmW8d1
cWDHfBFkdbANh7FgoTQrD6kuG90wvXEtVEzxl54AfkwI65mqZVcU80jayYlub+sq5Yc/PKHqtNXx
FZjozbpTD5+cUKh7yaSzZJSiWwTiGnuPCO8h9y/7onfcTjxoUoeyKOtQZzue/Was6UkBZJZ01+ot
0BIZ9aVz+NQSFtlBldiRDdDCO3F4ttwVgJ6M5yKMgby8PuKUrEjDv/dHP1dm1aFDxmytlX9RmQWe
HKqZa+4QDULkN02hwFr0vj2T+JDHyxyB9cqLo2NHcN08c2vHK9zyPdeJP3GFVzNzvauyIW38+/4b
pjAWYKhvORVyzpEsJuRz4Gdjcc4Cv6eoLdOL6Z7CKE21Ki/42hVwSQYMv5vjgnG/gFyVjVDAgeFl
uOR0M5UurKGbXB7yM6A1g0SrotrjklH3acDuTlJv7eS8hvYpn25tN2a1OHQFAEtE5fY2nTHswnoG
NhDKkqrwILApIPjWMiU61RQ2f7In/1jZiysPJlQ8XpHmvVgppd//+P+C3QSxmQ8al8TREHCcAuje
mANfnXHN0fVK2iKdOItTzmR9TukcAAgrOcbtqpkSbG6DZhLFBMLKCciVU+x28zruiP42toeEGGrL
11K5qF4ERRlhXFcZq24epV7G3rqTdXrmfrZkOSLpbNESlq/1cLEBJHeluLs8Vkc8OhHwUaygAjUC
FTpb462TrnhWtMcpPnvrWPzg2cnW5GlGZ+BeIvhBsw9JoihQKhOd6Br2uFkfqLESth+LMsKaHQRn
q3BeqEj7qihosZWQmUN2J3hlPeJD7xtGfev6z6MolWhVFSGvgy07vib/R5ysT9UuxbJAPsKSxlrI
onmc+ohyJYielPPU5JPEThyvhYlizWIdcCXWTm3fWXBVMnHeUT5aC6dywvNUBRcExBc1O/gDUCoc
SbYN0cUK9YnJ3HvwSCbDVvq6O2A8ioMX4UYvahxzOYRkz52qeqv0pYXunX11QlPfaPkzvz3w/JCv
xAuyrsAknp9pr5cAX1moAZg0+N6LfataL6z7PZznwrqprmzIfQHWFTnbb/3IBZ7U8E9tg/IlEnb1
OiFlt+02x2U/eodiBkQOlE6qVoAYI1/yXB1+1v3qk30fdr76gHbFOx0j7Xg+PfFuPdWUlWoG8TlE
KwDuafW/dtLG/FW6JFmSwW/FKjSv4KY/vQnnVX3T+udvm14FkS95tFRdvtlHbzuzYkCfG+V9sD04
+LmnT2GUC/iJgeg7M+misco/QAmJJZHrjkNfeRVxRsWz1Wr/74P+OOGJ5D6UlEcuvBurBCrKszmX
/4P14DtUhWzNwmwvyMUIGpw/POwFzR1pMSKeXnGlejiglS8i6Ek7gyt/ftUI7c4nFMLZgmBd0Uqa
1nAG8ZzYjzOskNvZAp9kfLHhFqS65NEPxcU7Yv5uBF1XYE2d/39iNC3LLET2zZkIuKDuFUUpmYkt
RKvLRB7dOAuUWmI6mZ2lFgyl9Bpb8LLxOI+hOqu5x5/V5OqyOPp/zsFH+FsG/aJSxpfUhz+nkMm8
m7UbpeQl2RtDEV7F2cKzyJYPGM81hKnWsx9zylXMLwwRxQqqPrOe4W1f9M9nLPIHMGkf/TErc2nD
S6B26YRge645sJfENXSD4outprY56oGvx+CcWJW/alqr+vG0vDmKpCiYMDx30E+Q3Xr7TPw9+5Q1
F3WgqoyCSQwz3RGhoZCQ4GN2MfCnBlhrF2zWHHld/V8ONH0DDkxPw8jhmCQV+COXfFfiXaBgyS5C
Ugyqb1e3hI2zUIhTAMkcSiTcrAhibvCd7dIZM5zDlf+UGTTHY7gdIggoykZZurTaSMGaBX1uC8JG
p4cObwjDDUBCte9WOxR95qKezKFsudn536nAKZTasQXexWubMRX/KP+DtqOXPCBiL864ffBTIjc2
atP2B6LC3+3ajq7A/tE/pbxbdnDUnxsxEemxAyxV/UHmwts35O3dOMQK6KJEPStPS0BIs0ZH+5Ha
AA16fgxQIrq3V2cnPSO8DIHJc59GpN3rIcF+9jeq9fyWGv2/VH+ARRgkC/Lqd4aKK03pAOW45LuG
K0t++viMgr7UX7ZOQaFM+wB/WLB+pON9a5FyVfd/Oz/7TED5D8a4Q1mPaIGfNKOPf3xrJAE9ivtU
yiKQJzTJAChVxNiPpi28M6f05quN96FDjGFUm7iNHBmtR35eKqC9S9+Xy5o1Ycv2uI1UFPfD1uAi
J3SBp2t5urODp/ToX4NEAgprww2kNrYUp0ewUlZJQCkfwDaaY4cbxKeyAcOjLM4YeIvnYhr5IFAp
luDTYjvS/FqU5bC38I3lO3Eep6wuuF3H0Dm/6azd8DKnXxzGsgUwtRS4EMopu8G7oLk7y+F9xOCQ
Xv4JwJZwRuFw8a/Q1hRC4jgqIAHwWjrs+PaBA8jBZE7JqYuM/LY8DlEchKiLKzgk+6CDK79GChm5
mgNYAuF8+E4q4sgwANlgVPbpvTs6mYFMC7yarGt9/cw0H//gWUZYDQrYYxAQ8W+ESRUoUDVW8KHJ
ov78iPQSGQZElOz3xpnrpXGuZ1yned+TEoQZ+4wj9LZXWnv8nuJGGlZyTKLKOFUzQEFFHIiyFDEr
NVt1v9aFdZXF5eDVAt/0WTiSW8yrmo0gd9C92VOIagGE5QQnQr+xtLXcmZ2hKqfia52sQjl6ZfXD
xbAu/lb2K2p0SXn97jwJLF1GFoHsgQ48LdAAEyn52IA/t41lPAfI523orncXs04RkdTsFUb6ujNT
Cyw5PTR0m1MfDTqhAij2SeZ30plLkY4dnKwA5KAUfDgfmavvd7zdzcalESsnu9XMBFVLC5z8EbWX
6kIMeY6zExEZAYF8gx4kQzLen9vMW/2GkENaIbHF6U8t6kpkfdy01yY5sj3PiI/hOiYdMjYesqRK
TxYzIgdft23UpOK5jOpSIlIYypdJixHF6kM0hghBJTbuuy9rdDIo6PRQseMONO4xa0SR3hUA/hZ4
VeYXeYfsMETO9wkUZvypBlhqNOebnoaNuavHs/K1vGJgILH0Pf9MKYPct5XSjkecjdU31VMO043x
BCpN5/YSMdxYwFmLO2x84JtH9YE8NN+I3v28gbtQNb36PkX492x/uBl7dMySMYFLjpb+xiP+058T
KAz49QNp8HQdklUZALZ/tZbgsnHrleegkdu/EtAnykD9t6g3CThnXCcwXOLjfEhJSurorGYAamzO
WZwF+iEouBTLJzCow9uSFNn3+uxkJwDbnCtMKGcpHkrYhQK4zQVXlFAXcwrm7L7Z3lAa5RSqFSJH
uak8KfAn+jcpt1W+s4CiFvAguM7KjjRVfu/gu53miN2r15aVl0AVXVSgbDJDUvltHQTgoKWCJD5k
vWiX6Po0gUo1/uFwmg9iEnG/0CwayPuD8TDh69jtVmLXV6cus2APpp6aq8UQvuD7zaGkNAADup38
4dSXJp3wvAZcOg8Sq3wFF1xmnIL/IKxfmM0SSKDe/8T8+oUhlfcSvG5EXfQCgImmtGKS2FmSJ7yx
6LgAB7z2gINueEex3S49/e/BOl7nrIH+ytNBfqQXtAmphVJk+g1ohkXBq5tGyzWSJgAvfucaSObC
23Hs7CS/A6+zUbhUhPrxIZjeGV3Fjp9qs78Tunf2fQ2LBHKWJnhLAn9ifdNjoro4PiQQxbPvnZn8
VE0pNsMGBpois0YNQWPFC2jAY5edDyFGMQpO+6JvcE6opeGb+ViTnUVBK0dAO/PCzroE5EY6zbo7
1gXDpvcHeUMpYtVEyuVYu/jr1yw8Q3Nt4qFA5T6CMz4Bik39n4pKln49E73S+p5mlaLmujOSq+LB
WQOD6zcCij/a+PFHDOlYozu6ke6HjNa+OdKDaxT6jxBNxyXlhmXnGfcxrslZ7eqCGzM9/gf6SmoE
pRjbs2TWGWLhff+vH1fmdborFJOyZjhYs0Tr5j0Q0W9LNPR+zFZkfKenZAE8ljKVsTnjQXQho6wi
epRKPkBBECTkaNUHoJljKhsTMIS4n25ZNZFK5i/HV4p/h25yLUZNsUQkImOjPrBhoCNt+EoNlSsy
6sz6kZoH5cIWg5j6YGYVMecCBWE137BXMaF530yiJLTJuPf1Z866TITe+zPR9cufz1XKzk6+0H92
WLarpo26oaiNoigoInI8wJMv5FkiRDj+FsTQneEG/Qi8ObvqsLB31yi9Q0/kBUbHS8nrDD+WS7s6
2fPiKQiJ5dnIdTbEanWAFeShgSPFMOdwG84aqtd+SSKB1I/nNPkNrbb0EWL+JmpRQjuj+yp23G+3
VAOk5dYVHQwZTXamcd3Hng7kFaptRiHzeMIjpLiq9xcvw+VlZBt3z7xKSW9LiOkGSP/w6tNWFfcf
tggCHZx4EACsDSMbi4TeN5VLuX0/ibHYuY1P66sPRuo8ly3TVR/hupEB0HU5ajDdTzz3SPa0rQR0
HRjXYxEW+cEDIlXZI5vt910WYriI1S8gw4Xr6bbrvBleOFdtJnaYmR6V7SLbyQO64zSyqP/Fi2KZ
j0JIUbgoYdpl1zJf/Tt+Ei54rwk4CJTQjq00lQpnqJqCWB8daDzLWw/3tiSfYdUnHfEeWZA/9uy+
5ICy9RxTwrPis/1V5Iar56YjezamH9p6sg7xyUSHJcpKxL+boDwh1eTSpnR25gNS+rVz5qkz48fb
pxB8yZIVWIik2ApVvPYp34qW1pR94O7yunSkdfLfHu3T7rxEv5zShgorHkhIwJTDN3lxD8KxJA+L
zNiEXM0yG2Jrq4L22CHfDzpWKD0touAQIgr+z+bCyQHYR+sEHPlhE0d1eh7xs/qPNYo2SflGGCO6
Ybtu5/xSv6oiFnOP+7y4i4Wpv3PVCeRcZjJnFSl0rtdDMl0gVtzcDnCe0yVh3tbfjYHdCzPCPGzQ
8s0U0Zf9/x48Pf5eirC/vvbAal7iXuxpJnwi2KnFxmHa9p/jdKudXilBH9Sq9NYvj2+15pEmJcy9
Sc9LaKIoh+9FVhuUOfrn7XFD88VUnjmEOqcMyiIluxjPrpiFTWTKBIpL05ENuXybMVOWPfxeN9ex
Y5MuaYiOr7e3EVxV8RPsDdf1rRUxKYz7DYR4Bg19pPu1AXMNjMMhxM5dm+Xht//QAyDidLTcJ8ID
NVYH2XC/EFK/iq/lBatgqZ8ykQMqw/JPGR4+OcBcRYY+v7mMXqtxp6Vzou1RkDwbFSpfGptHJ3cf
UL7NNnwNjifN4U1FJyD+tF5MiyOX7gtiweYWvIkEYqAFmVN22Oa89quQ51k/RwVqvAn2i0yfHods
3on3Y0AZA79GsYMBe/YSVKloxOIARmnIz0HK49+3/znmck/q3090vdV+ah9kj7kkEAoCKUaLCkDW
Fiq8ue7GZGdYxN1yRuyJC/QmHACRBOa+yticTobYGbBPfiLaoT3jBALQtcjXXGeeeSBbZdJW96kR
YpoCQzkT7bn/5MsHci1I3jHGhxm11dXikAgmp3WAqMHb0i6IyEZk3mVvg+cXe4DE/e+tzu2lW4kG
IMX4OUv8n4wP6GBE/NIk8sO26YN8sUznQ6UNOfLqYxOL9Bgykh08tde/fPCeN2/Dgge/QGgfTSFr
nzokNhhZucCWUKlu7CYt2wsBkT6ZbTmMEiSdFn9bzBhVe0tjAEsTgzQdtiXvzDs6JnOiPAoz0HKY
azSR4GVN6gXnr+j+I6WEdaG2laNlTfZamp3BPJtyG6gdFCj7CeH33IWnFI1oEsruzp3/odJbQTkR
zkAvLFG9XnNkxEazCWg0jLBtx6JiWyxIBagrGWPcewJkXgVYe1qSdatDt4TdL3He8lwZ53jKu2BP
iuRYxRJEg9tSOJhpqzitnLsYDkWLGSBIRM9/ixZK0YJCQkRe5n2ZCma55yRF7pNPfrtkDdD7hCt5
TkOkC2Xcq1rS6HiUCuARNFrGLZmoTSx87rNR2c8nHg619r/z9YbYjud69hmMZu4AZWW5DDzTUzwk
1bWYe3p88tMs4aLhsKJyM3h+c1B28n2rIt9P+f/eqpeztr0XwSrhrTptHSLuPtO8Pr9p96LyK8EC
mahwPnbA+lOihrf8Pt2YOclzFBcZoZMucfwqKoXwoZzKOjLNvgaXBMmjEKlDj8w0xSoTYZ75eW4+
jA/CpEYtZn12rs6YaNAOvdVmtebgOWykurfueqwatvn5Adw5X/jWPsx4JnddIjQDFm77EhJQcLR7
09P+d4bqjHYWE3drar/m2RFBRHnwAXHKvYD6q94CwbSCnKDGnASW+sfe7ezEq/suwEYfB6DD2T4h
+RvU+Ji0v/wXo0So9QRvB4l7EQpJJ+85cdC9bwhqVW8TdgOzzE/XWHz63BXWj20+yFQYTQtCJcHi
rPxJgDSZ3zCNX66x9PrhlpGizWigEUSyWzOvhMzoqVte9DW0V0SbecbKAq+z36Jl+llb5f/0ieb/
gtDPm9t6DIb7sTnuF28cu/FmcI3wuKryN6Py+nNLVIyVVpAxn6fRG2Ef6nOET0sBt+Vk3MJulWzr
mTAMwV5VJ8MPOuRzhmRAn5mwxi081V+nAhYJvb10xIO6Zd8a0V4KdPrGArpfZY0yCG8YkxiNYeks
2HlPUt1SsrExdKuNfFm3dmIo6hLo+TWgpL/QyHxsJ9gZHpWWRpknnkwCMOnLCXjBur/J8ZXzjyuO
Ek1nqD97YwpWAmPBdrjWZj7nAgTd+p+XKQB+2SF03lAYTwtUQLXYR69ykI4+ogw7+uImZuAro/1G
wL9DM39vIz3Wbj6k3SXoU+TZHd1ipT0qBiWpj3l0BaV41/NHODodvQSHco21n5Jz5jHdSoiqu/p1
GXrhGXXxFvPRl7AhetyfmVGyMBXDo8HZH7W0OCQso/3KpHKFSWCQDbytQwB3ntF/g4gvTfvXmPBU
IXtDm4zG5W5v91Vn7j1M8OkkwKDPmFPabFEQdqO6iw7bxqaKlH+Yzdo7PWWjCEST1m4qratKTFFw
WJSEHE1HcgshVj8xTB/KY5bY8YISwUls5dyvLOHjrav2mdvFhyYsu7Z2dMt45ldtXw2VkhEQfeiD
Yf4cn39imREyKkMxk9n/zJs+hKyDvUCH8D3diUSES6ZOVK8Fbundr+FXqy+lrT+q2ngDBHtwViMj
kXtPzm0xy0FrIJ4dxrXY1xFg38buXq/96ZyGaJfQh+HMu+C2YBuSR4c4U7J3UqyvWuqVJot55p1I
6K3mzKNRSkpARSbtdvjur1neuFR1PJazDl39xHfbiJ7qvtoi7OfSZmHoZsc1PndoJKSHIxkGxVfs
EuvcVa9/7xtD9v6BHnVkfP5DoN9tULCi5M4GVnE/9R3AuiWugMATi8vJkqMinEc0IS1OuuKissR3
lZ9J4tudT3W9X/NAX0h6wYE3jOdllZKnoV9PKk2XNNsy0sWUBdUi01u3Yp+TJaTz308l6ZwrcFOW
el6EtJTYbGl52Nz7vc/+l2NEEtf0xgyYu4sb4mbmHhlVCb0A2+kGqkPOkm0yRSqszDsJxaGcJG+a
pTYxieqJNmuC4ZtHsbxMsXSWnu9qQ15blTssaAKdQZoxCrgxgkg0LjD/Ujzzu2EhHdmIIwvh2SYf
xS7xKjwMY5y1o0ZiYIgLyXTOFwNRJNjNV0OeTzlj8eEZiAmRcaklruR+0Ps1EoW1P6EXVG3ptdyv
zZCO/nlQAEbOo0hfIM2MHxGC1DwVDOQ5yJVJswcNz+yADFemdMmCOXl+oKjm7od7KYp4qT3qj6Si
hK3dufM/VvmIkEYfw0YsCL2uvUYI6Rxu6gHHTnN8UEf1kwqx4g2nrHejiajUjnmPwcmIzf+bQv/X
bJ8TcY1b9jYSng82Y3pHulnZWoDSAD6LMkonNO10ZI1LwUuUljcI9VDXlWDlCULGBXsT+oMIz+Ia
yolLBPhSV+KHeTRGC8+9RBONg2h2Erp/eVUkifqCpCwjyqBksZy6p2eRMl/uNQv2g8LaZlaEel54
QZRngeI4Mn8NZrQaFJzZ2kda7VV/tmGrSG58iL+J83xMvnUjVNkDLbs5zM+EMdHti9AImRmxPVg6
I+L4W9CYdIAwGk0abWPqvZKTRUo2U4NEoDsAGjZkhAEv8CiOwguHHSFUxZaqlH9ujM012E0znxbp
Aht1OjLmkAwEAWkg8qJsPQOCSnzdR7FKJs4coVILlMNEq2Z9wc+zrFkjbHO0yNuN/FJWTMuoORyE
CExRz4Ne5CLhAps9iDDQB1Z0SeiKAgoJin/cpOh1Dck1l+q5oob+BSnkzcRhXZY7VvEVMrLHjBVZ
Pc5cqgjIS3RaEvY3RiRzu+UqlfyrYFLm0TRDtDzNwgsDnUrve0qcwuXHQTXqrD/DX5b/IOKD5RtA
4TWNKDLw40j1wroVlUExA0FnFZqVUpxCwQS6XjxMoVATclnAPGcOyTXT566H3LSoQxoBfy0tFMPN
VlXoPocSkEMlDmvVVo+kllbPwZfy8z17rPGAWyAYHQ7OdiFaGo+KIoNq6S3TG3e8x7CA3gJAJSSK
cluwdqcjR+6dd2TzRDze2wMAHowkuKqofGQhnV3j8fggccyOvE3DjFkYvzW8oOyQ+5oc6rmZvn5U
4+xBIgu81drJ7mBqKsR3XSCkwrd1vyhfrfSnr0ikQDv/o60xIIWs2jgb/bz2WPTheI4VNvtlCx8h
wIs2lMrfh/RJUTTvA/SHM5dcIO+gkWG+5MrzWCjJX0ndvxOySM18qsjcZpEra2btx3+afg8EMqMk
hW0sEjZ74sDc3ESSSnY7licm0RCFiiuXLR8QKw3R+NxCnKym1asZ3KUl+jsOS9+2gNI4SpQazFip
copDhig32G0reALiW6wPgVPCvcBBxIEbK9sAA8Dlkd11tqVWIfamD5prsFGyG63jvBzb5RCRPMzw
Hd3mo2KoQ0xCUYvov5FyvK6UIOAwMUg1aw8SGEnp5iSbeYBbz9I5VrKB+9SEt0n1IeRnlXhY7uHj
pY3twRK1TCay18shwuwBqjbd99qt+VAVjpSLII74Kt2va/1XCyJ9/ENjJa6PlssmDC/B0cr0Mutj
FNZyacE3nwehnGBigmYKLEpPuf0PssK/ja0+wWOPGD4+6OKCpLY5rTFS8/G0ttlQrL4K3nNIYou7
CHYlz+I4S6ZrQQwjkygtsfMBcLD8SxNU7ex92c1/1qiW2MFDcAOhJ3U7zrrDeYj+R6XRQcZRYFND
Dw3kSW0CfKkC3aapVBY+KdUhAgFb+OfAn8nLSfmfbEIWyFMy8pYekraWJVDSMSIAwHkSP6EuXwv6
7BbUnG9K2MWbZIcp0dGZzhQ2x4jrQ/PcSJ6GAZgteOFuwpavaJAzqvE2/4/kw5DoDr3ssOdbqxXR
ap8fQdHse61GL6wCRHBhxx5y2Y+obb3pNRYn+i91QT2el01iP6fiulQiVF6yDTNXikiD51WsTii8
jijCdaigs+L/GzHCL0YmokugduqcHz29g8d/0vmfQO4m+sZDJya60irl9zLnr9nDGyiz8p4kARVL
JJ7PbTZYT04oVYICQba1fKPVqAnCoJHk8F1gW/Ii5jiyVxH9QYJJ4N1/989+TsHIynz57BwOCKIw
CO9iUNKAcN9VbsUUJqLDAIT9OBzBx8FxrNwTtShGUGApC0NW2LbRst124z4tqLGb3gVBFT8fdG0w
DCglcQ3zNOZaQJvAv1kJ8p7u9djsrvGIZBGehkSZt4n5+avNxHRAgvawEtUgNEu1QTEkLjbq4eVh
vPIdsSqA3j0iq/UgW8TMDNO1YUnZO/lY3kzzwAm1563Jz9uoKAKeGCXTiIER2j0y3peQbzpTyEH7
aaXNiavt/i33LOjd15+DbVhpbKFHUZjcIBqsiJFzhZYagLxUedkWb55Y8MJUltAciTwgcdGECx8o
DB0TTHyv84sSX1gdTHvU+H+fXF1bZcwT9wHAtE9Ij2j9OU8ec2pG/2LkLmR/qvN2mFI/ts2Csgok
aJy46Q5lTllc7IhZ/3AszjhexPeQzESPywr94cfPPu/ARWKb4mLhjcpG4i9SRl+ZQEtN0RnrT0L+
ZgiWAyRD+lfQcDh21H2Nqn9dKfXDURXKf5ejm71strOp1b3sNP0uMSGZh72Nb1exlk97qPuGOf3+
00iGVtzJl38rsOYwKt6Sujdoaqy8N+ddgp2AsmIKLSMBhtuv5Xa5PAy1uw/wBYCiRT2P0wIQEaTX
ghaf82RH+zdzNziw4FwgZt9336zR56JPZ4m5yIVveF/CyXzGhu9jT6b4W5MoFmKkS1TXeg/Fh6+M
OBLAWr0X8Q104a1RbIIUe+Sf8pu2D+vZ0LybFPhkT81SiLDfgb+wLcqjeBZlfg0FSRzjzeA8Wz47
Q2wd8j8/mXnlojZH+VqlS5SvpUP1ukKeAP4W215uFZhxhez15OE/S3RjzG4gwHFcGkDJ/jEv195q
e3tUsIEEAT+B5gWPYhCS8w+NQWBfAFxZFj+20t7v2nLj9fMRxWiz33PPqxIcA0y3RDqCXEmRYHUG
eS7KyCW8bOMMlujvsWRoeN5WWown/sPMI3PFv8BFBcNZCidK5R3Au3xAO8erQQ2YBrNv9pzpIRdk
mDf8ictvieljW1UuPX9mVji5vDMbY88yicSO2YvLagWkWWcpm3YtmlLTtq/+VT/9a717Eub4YOHt
AdHPX+kK602MCbvg1VZm6+X31/MFE6WwHzMzc8Q3setqrDmMw7grBzu/Jbk+pmIJHZ7QAOT4CIPl
4TTsJi51+iZy/ekhfhlus9iRDDIN6G0nyU2w/pHJasSyUX1JUyI7O+XCRcPubmdIeIwV8n9od78I
4dYsuwHxJxQMfD1x6wH7mjYQIF1aHbn25IDIPoEo7kyrHgQskDG3zEYH1Su13WLRYfKqZr+TuFQE
kO0vkbsmh5dCZ1ZLmBGP4PK1TRmFiu7Dw87dXLuu73vjIfSvDK6MhMQtnANxykJK1+0nGPc2c+pL
4OOoUS71tfK0J3jlTNqTP9JF9AT4BrSjX4TuJ0u7fLLuW6XokqVfpMFg0QIg+Ao9Huos9vCZbRbL
/i+fZjl2ba4Jf1q0gzWwaG1XMQis/rLvgwu6nKj8jS2EMzQGeplPCYUi29k2mz19uIYnZB30kzwX
Wj1VQqwhZZvhQEUEAsrUCswY5frGAsZbdA6EdZCME30hSImmftiuDIQs9eh0l6m8uLgCyiD52do/
JvgzgQOcMvV7CUbfLD4nzgJMSjdiHt/TTKfQ5/cJDOY8sO+o3mWsNgHx4cc0y060UhCN1ACXuwWC
gp44NBr2dUfE5CNrs/i6hfkCJSjUtYsXcytNELlZvPo1ueA2kkOuQiWOPtpmCh4Sp8kxgFC7f8O3
1ZP4hQ0nVVo7varBm02f5QfGG2sn6kYYyZx3eO6zV8BBCbGE9XRpPf5jxvjxn4Q5qOdDbiLZvSx4
7tGkYd4HcSZRslZ4OprQVbBFcwQI9a7yc1AYn0SYJKwXZaqCyoL+VdowrUuJlV/sNQZ/Lm2jVD2u
y5u8blDwDMNI8WSrw9JqS6imSz/3Mv6ns1DaMjuWdptjutQt7pft+lxLESe4FaTXP+JqIWJfDHss
IzfE+k4qdtrGSBg6JpUSHFKlYSMS4nTE9kXRBeqAB2yyhlZYW//AtNBIcX81iqEjoLd6DUgxoCyb
MWp8uqZ/wCpjKxfJ3e0WFu3mGVQTaCHo/4Dhdqah7Bb/yBSVAax5vxe2xFdrn/vxqRxut6CVmFc6
4wDKpS+X4sdnG2AU/yDQ9ERO4H72iorv+7+DvSXMcTaJKMkaZgN/4ePZvWUqc8w5N8kyBbgUOXQA
Tg2QPzSrtv4ij9hiTTne2BN04IFI3Q/z3H5uP6ldp0mQECN5ExUPMUB6LIweWpgY4xHjc+E3Bcky
FcWanImL8lo3Uoy0F0zuGJmItlaAUiN2Tj1rdf25U3wwZIDlii9+3WJQeyzwHXoSL9hlJCbXz1tF
GIZDQ1xfoXgJeO4BVfXPjPpxFUkyfks4tYHro28sM93cz0ZRwK02WJZobZs9C6jdBdnLSGKQ+cRD
r+VFK2VYqhluyFroaInEfnJgtYzfYubaTBvzR0lkLE9T6vYdEw7UumyLE4NGfDprhzS/uzw6VjJW
numhCkHoOarDHXAx2MB0G0r8heEV1iAGjHp3N4nd8SDIIV0wXWU+IlhsK1sLEAkD4yhDLTrTDBQ0
+iXpPBnkk9zfOejU2p0kMLZDSzLVlxpq0l8AP7sll8tvCMqvHxUseySvZcPX+I1q3XqLbokai8B3
4xHiH5EJyIb5DU9MO6Nd4U7/pF9WJGHfbMIa4kVkluuOv0NmPYzfRgkrsZA9i2L3Xx3MehWNqZne
L2WrJZ1jajE4c6fa3uHjhdSaJ/Hj+yAOsmggz4Z/2O0T8Eoa9tywaeSeCTmZ6UAK9HkCee5lqjkD
EI1FAc9wMi7lg5jGbPn8a84+BDGE+e4Qp0kULvIkkZ8kuz4ETMgEAnLx/w1cqifboiPC8aebev2A
eNUJTUXjVIMntMs7zKxPSXuGv2fthlhsg2awNhZrA+40aDOD533IeMjXj7nQ9v88Tcz2EGLj0hKI
1jsSe8c78AH4hLcMir+ar/bxYLz+dLF6FAFAoG3Jtfk1QXjViyJUTxmVp3yFA/lkng3vkojD7igF
/IPY2x5ddX+oeKTfDzGvyjzeK+921mpfOcw9fgxPVx+cD+abWiXlQ/WRHf1kenC6PyhUSHg3vX85
lWTqRfbBOgD0WeqH+HeeXp+5MMggbgHkQrA/IgBvAAPj2Tyn2RewCunUAx56NjCy+SqcLSx8Z+lw
JgZtq1svDvgBgI240lettXrTaAXb+MVKFb4L7Zerue0MymT2dEtJNr31awo87YJE5Z94cGGPFAxX
6umOWYewZDy55Z2iApmlgH05zerjXYS5k24Y0z12oD48swNq9EHjI+sAT24szNx9YTG0TeQy6ern
W4zVD8bQLLCjlvAlc3gjPbi+0ffu8yWJ50V6ri8jNhnEx9r11cbYI2e0SZ9G3pi++CMIi2vFlatV
DhsCGk0TZEzcECWDrR/swEOwfelguRVvPxLwwGOkGPPGrJWGDhzvI8w6tky9jV1ds8fPtnyU41I8
9l5rzJm/ICD1er2v7VI5SiTzlXgkjy/0Ssuk/D5y96CJThsZiA42XbkmnIgIoS2xwff8jaO1qjWM
5PiLyJliitl61bUQxMOqkTwDjis19B8mTPq1IquZe+EGy9JeaveGO8350oWcfWxxU6XW2AHH2LwE
/LasDooCfwPVgP6cfyKHodzfYGZqZ8LpPKOkcVNUZfv8XNe+3z6FlNurM9BsXGfdmkZBu6LmyDY5
gPxZHAEB4aS9YgvNMatCmq0Tx6S5MyqaJ4kAaQWRZkZD8usiRy3WQJkYlrkEvsN9XXQSy4v+u8oV
54o6ujTGduJkuVUQRiFDyiO1I1qsRlXPm5Hfey9AnlIbf9XSXQdG6SrjovHe/Kpgm79qighcndrZ
IX+7SPcV+W59JOaq/SCVrkCfZUNT03RnERJx8LlqLM6AJGmx1m04+XlAOKmCGNC1ERs6DjLhjxB/
L17YlnFdFSJ7DqTDPh726f90PdRY3Az4nD1QXhpSsl+BmxO2lpw8cS/I4lASkHPxbUbI0zohRhYi
aDbPoWYkR543fJEvGHgL2vY4qTWRsWrANdJ9fsORQSj+rXgFgjRZEpdEl6rfOLapQ2m04lIJKvhx
gGrQ2tUPUBBOWefTmDA9T1cqYWXdZdgp99RpWEBYPWSLUk1VhC61n12gT+BBwaTvtvPxQyVjehpu
qF/FEzRrCP4kPG72vEaopj2Oz3mlMKmT0dQqUxleRaww/VlqgrCEkxiFFaEvKLp53dG+qhywyafJ
zdK3p82h4DxpL7GJmDyjJcSNaYSUt0vvkwuLsYWnII/3wd/4mc4kfzEBg4AZT+OZurmgcwc06QCM
xDxLBUJTDU/DdguS2t58a528vP0JBJUWXhEgMMPKMRsH70wLywWILg6fGPOpsYxhZGIh51JlR0mh
osyU/iDkNwKejOHfKtzSnFnocB7sotCL3ke/gyLAMV5lORc3POZtLUPSwQkhEl0XqJI+WJehH9Jz
nTA+kVoRxlwRq503pD7GBdEmjSqOIV0+wNiS7UeuBwnuWe1RkWeOX4rK508ltPfERuhiSFpIjafh
1PAbbSyYYYGu0+0w0DYueVT3lzQbsny8uyWle24rg1pQ/c2yu0HEG2V+K1rg4MbmcCooLtoVFjUN
hno2zYgZL0kxkSDi6m0SM1cHlOtwZhkojyEn3Sj9V3+iRIH+xWxWN75QNZgyJxNZE/6Bx6+P16Fa
g7lPGLToCICNCMXglUaYlwT3nYLNKsGDlYkEpasrobp0KVUKQJWcXn7gAv0hXyyO0Vkmsi8V72Ef
kT3bBblZysxgQVwu3wQjK3mlaJtzHzOuYZrrt949JO4X44AtVWgXsQ00IJXi3rxlaZJRVDjSwtrN
3cGqjnLHJohWohVQgSlaJmKeWebAyivo58XWXAMS/ctKRQP2qHAmy0hO47K/CnOCkKQSm7SivF42
i9mLuzUo6GGEz+YqSW8KNEzc/f9S8Z6uGpQrgWKso25dFEFhfs30gHt0QWjUpPn2fb1KJtLUoGmj
Jeg83ylOKvShPERnXzEGFpBWC9HGnXtteGBT8X8V9pAnjBg0wFJ9ZR6EDD7AIDpJbqPkGvIRgmm9
tOplCpbykhu183PLN7teG/6OhYUHTSSOJGHd6/+2XcZKPjxWqSZDib00ypzlu0Wh6uhCZ0RjU2ps
eOneEBbvLIfH/M+QOVAQ9hnAS8z+V21dSNDT/peP7we+931AsjHh5Dy72bqAJTILfflB1dmOjXEU
juPluDUKEKJpOiteAlklGTNmBlozJZRAfknLStNMuOI0+Q9UX6wGzgBZktUMaySj0HtYyWTy3+uZ
m92a5B6zeXfNTq2Om0WBTfM5BDkuqpZBznjD/oD3Ab9Jt6GKUDnJzgVdSyhaHpRwIflaoD8uCmE5
DzJ7zlEPeb+rXo2d0bJ4QOwqPEmX5fQWML/SqSl/y4PdlEw0e4+lkNYJslQ9miktB35ERtyB84sl
9GPuTgdpVSjNmbVs+dDwfUmkNmIvft/e7rPTcx/3p0zKKXKJQo0hOW0fnt+iAC7ZdxewtDSLuHqg
7A9TPOQ7150K0cnSUuOebmrlOsu1WBA6/QWecS6QmZhc+fCXJelWBlQWeZP85yVwH4OzNqpyZU2H
+vqSNnPi8xkTxoxzL6S69FJvRiSN4sIjrdsoh0tKm/GNuSZPmdRtbhrXtAxY2ukgLkBIw3rhaMpH
YL2iik0MgAh5lfE1pGIqrodv3l04idIarQR3Rt4N/3sVOxOwhy43KyrnUoRqUsWdtbrvSF3h1rlS
SjRaiPgAqPrajt5cERy7hF4jneFC/eLZrZ1+B/K3xnIaVzfCRuijkP6Ernv4a85t/q/rcbUMW/Ah
id9oYz5w47xO4s/T6J03msRL5h81qrChAKwDk4PwB1m0580mkGn7pwvcXU50XMT/TXUk4bNaivEl
TbGB05mimnuuOUHawi8IWR1qNhrIpSYsTokrlX4l2RmQg1MAMubmUZ2t8T2OhVeDJg6PmgqkHNH0
Mrk/XkPMjze0fRFCm5mi28/LAKTjF8ufkafJ0QasvavwSR+DDg==
`protect end_protected
