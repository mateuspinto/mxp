XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��˄���}�n4�w�^���cl���n{���U�<½\�ъW�����:��9[������O��ٶ)s�滠Z~�	bWVeq>��M��擽�����Q~����e� Vuѓ��1!��@�nQ%.�2�20s�hH8��P�v�����.��AX�������L�k�ԍ%'���
���љ�V��!]E���N�%V�A�9�TG��~J�M%��J�{��]��4B!�cĺ�X��m'��}k�ў�Ċ��TFRPj$z�c�Î�7�Á]���Y>�\�������]avl�=\�;EYp�j̰��Pܳ�o�@L��C~n�/z�kmV�������郮U�&�3
\f�]��@��y��튭b�$��{���g?���8���qNȄ�Z��ed
�P��nqU��HN�����~�ͯ��=�D��V�shOhB/��(
����j�z�:�މ[�\��H����Ov?������5/�#������w�|eAk)�
�>��.4  #Gz+�"�)�LA��f������c � �8��u؋3��ڼK�c�N���X���:�Y��"HH�����'.�f��w��h>�Dk���z �Q�v+k�����@U?U@U�]p�h�*)���O�ܮ�jeI��XºA��L^�n�l�6jQE��3 ����x�T�c ��I�{+	�<����{�12+��i�2~�,*��L��j���D�UTS�+���/,�W�#yC݊�G��^����XlxVHYEB     400     190
�x@?y�D�P���#��s�����P�ƮԻj���{��4ů��N����h���v�s�剪��μ�N4ۓ���ID��_�>5��Dl����6��`��א��K�9�+%LSF��)_%��;<�Fq�E�I�Z�4���/��-�>��_���L��A�K�s�B�=i���:��z	{v�L����[y���V|����� �2��!c}_�����K��՚CƦ_o�0�������o���ڷ4�qPs�8<�iA5�>���:��~Mt����+�[�!5yw��R�6[v��F�3R�M;���KP��ѿΪ\s�92*LV:�n��B �⮭�A�egjMe[�Nfl������&I�%hb$��k5�=Be��XlxVHYEB      3f      506�d�8b/��j跦��sc��K��DJ�bc��@\���^:��zj�]p@)7�ȶ�#�������o�,y�o�?��