`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g03D4rMsDT6JfeI1+A0W4/BrCqOJgiFPieh8DdQJdSi2z8RsbZ67HiKhCBUE86vdgPK6/RxhM8Vm
KtKAZOVBgUF9GcwaHdBAIhShTP/HNfTKRXc4eNK4SvxV13nnSQ4WDi4E4oeiQfzx+hW1FEqDt7gu
aLndMXdAlUv3w8OEfjRmDNQDGvLvbDQgnPVGfpLep6KGZKdsctCwbC6O4hqF5AoRpfMEmJ43eWqz
PjBhgGTCLznyV7shuIQMIf0ZvDbnzyioWgxuGIZ2piHDHVvLmf6eTjlkhBBKCJyazPB/8G9ZY6cw
hCDz2Y+jb31v4lvPlwSaRNID2/zcaG7sNesEjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
0USWSUGxovGsyBJteYpEoetM8dBXIBYjwIIJqt3PQwU22X1/g08lEhuOtgxYLr9N+4bWHOT58XnY
whRr0UGUUvYM6/e6gn8Vm6ux+0L2bz9l+OXHkjSJXmODieceLef+mTb7qjzWAXuecutxY+ZYPSUs
V8TWiAt4Hw+1SlXsmxjusu2x/2zuYefMYM8WlNOUDs1TLipnXGfoDmB30YglSUwZNrtoM2+uXqL7
A5v9f8CrXmZxrLFCljVUWvYtor0NxYlq+wxXGGdayHx4YsKftCVUU/p73dBnqQtQ92PmH4516tyx
f9RrxP2/WmhkMvmA12Mg7tFTTEmV7TeJr5UkwUEkm1CqI323CpFWQwKHIGMmBTGHKoEHvC0fVEbB
dMG8mmhnWCxhQ2jWsHbe5VuvWXQV5Ou/g7E9vsve5zOE5B5QB/Lqq8sAagdFzXyx4pyu0lhU2M+z
HmpTP+dIPUjUchDUC3uNu5/F/CLLVPMf8rNEvooXFcOhksR11fhiXNpsDVSKL+InymRCl9y1tIOq
ON5B7pEKD7yKLc+YClj15VKLpUpOC0EZtBV+ORcs7Q7qxQqBfpVNCcuz4igWttjOyP6q5zfKdKEH
1WDmdqONZMS5fRg4T04j1hQMT5lKWMJGFyol9ng44dZnRU6N9PvRNISOHR1ACC7aRHCxICfxo+kR
YqvfHbaAG/oKVryd2iyBPUZEV0QU3Dv8ifKnuq0N9PwZUD3zW3oUnKYbkHEL1YnMSgKaTjYBtXGN
Ku0Jy64nbPqFg2MzllH+ozHA2J0lQu86qQjSJbCh+UUQBxlm1dDgbHhJbWizSoRb0OlXCRLS5o56
3Z4jDyo485aEMzHTMHIIBYBU+zWxyhZoDRJCaaV+CYhANdMDu9Yes/9BaiSS4R/NjcmskYqFg0Kd
70BDtjJeLxeMExRSKeZgNLGdWYAh4qZ3i5OUhL2RCPMss/gW5z2mYloa2q29zlj2MmpMiQyZhEKI
+KxIRbTePNgJE0oT2G3spSlC1uJoBG8Nd5jK61+IX/FC4HHWOmaZ2uAgjB3KtrhwozowJavdRSWG
iiH/irDkJgRZajOQsyHcwxMGWvnjOxONGeVtRgRrdbDDCjdkT06m7P20dSfUwh+GTypbp8qN95+q
SRR+pOsSLDx1IgTD/LMH9Ux5qPVBdNsa3kn6w82b8gKYQ2vMl/Qb+h1R7GpUW9tPGdLTPbcPgyRz
B6xUYx44fZaKxV4UusWM0acNY1ZNhgjoxcqpo5pHc2wZqSjvv0sjXgtA2Z80iCR5Ybc/ofsdom1P
tfPH00UwnktB9wiHWBKjiAoJEp84uJBTHDNsD3QuYEOQywuVXQ7kwhP93chbCq3R0btGRNONZ3e5
pxmKi/o8fQlIISdpSDclln9frbiGl+SbpN8ozt/K+3ICl3LpFvj/gsyLDtTcRRsszNw63GrwBNM2
pD3TARLYyUJxR54XwNLVuUGyEbkGitdLLhVf2UWEyFRcZ+bzBxAhhfXJMiKqbex4+J9kbZqjaXd7
EVKrJIuumuc7NqzWWMMJBZ+C9qNcxsFBczxVolfHNNaDGlnCP/HfSVyHefNccQJe9z6lXqoO1bMT
6dEGwwZrvaS0yH6sFlplytEFTfBSNklenB0kdEUJiL+VF/7GEm0k830xhLHQjCZjvpQ7R+C22pzc
oEP49jQ3fgRZv2jBfUk9mQxkYLzUOqGpMqVtrtLluIBvZ6lx9B+f1jHc37IHgGAd+8LrqWepYpGk
PcClpQgq0NmJnwvMRyUPfk0RWEJ0vOZXfKqndkzC7OvuwJqTvkICRFUCdcfqD22h19xsbOwm+nse
ufY1nWwXD+JP9OEbr7sVV71MAjmTlistnzATcbe5n7B6g6T2a+0/7FwciEyODTYci1ZDmzWqm0t1
d1kuFzqaorpgpWBYm3JUye2oC/ytEDsOWc5MK2i1SR+QC2XF7u0P0TfECS2jzQu+hvXiNQE2YwyI
iT7ZOoZCCR8fB5hBFNCAkUP9tfNcI/vKY0xiSxG0z+n1eANKhs7kKiM0UOl9MBcOhEBj9SXTHDP1
Z263sC3UOB1TQQzQGU6cmUPDcLWGqSRajvaACw38A0nsA+YUmPaEH60p1xe+axKESxjvPtlyNFCb
CV8yT12MCRCeiD+sgnpAdhlmA2WJDzmAao+Uwj0z+V48k8H7MXE9bOzTvUFPRCkl1do+QHHSSsEH
VMsmHKOs53NC2+fZIuihs91/BE48RUI65OMZv8Wt5N5U8+FzRLjeZR/hoVOdLhODw6ECpBhj6OjN
LWLjbrsYNW7ahDZKxYZqJvWv1W+CPCRXrc0Nu7DopngCxVz475ccu2MtUuqJuMmpdmxTsS0oc64i
/0fCn7CFDiIYZUlOpvToN426TU30mY4Yuo3haPXHjgfNPi4HYKatusrsz4Zjsaqhvbdm8K6MUnSc
fSyWS7ylpJ6K+n6Im5dnFOEDxrUAaHSGMUsiTZOfvVUq4FT9G/ERNX95ssDNo1pdg9K2VJY7MuLj
/CKQloAPjWcZ0xm1MAidy/n7LHSESLywNi/qNZDaUTUsKJxiFo5BxP+2WguYtp4HH2mnceEBODI1
IL7UMeKns7XVoFqFde+nV0mCH3R8MdHfawOs2+PuNeWvMSHJeABmJtR0DQOXayx7JNdYq4K8r961
sNOkCNGVUrdluqd2vauFDkwdybNaoB/M4/WBjYLSH8De2QfvxwP+JN59/Y2yM5nWez0WnQkVjE3J
skdSQ+7o07wNI6RS3rTNLqDGcihqagQKjSmA2nwa0UHITWBTsY0BEptohVPCJaxZSu0qbTqc7BdX
HuwnhK8w0xwCrKYdO/QKiLxfrBwOxm65nlnaVsCp/VwyFV9shH/rX/f1vdy7cUxdOlQcu65A3D3W
q3p4QKQmD43WN9htbtnX9LtgHLp9/3hikoqbVgpXlc9j2mKrxD9nfRbt7CRmM7UymTTxJzq1HifR
1Ty3aQUKXMn2yFg8iKc0DNECRg3zkokr6Bt7BqoiwV8UedMcDUqYxLxDUusNHnWZ0sQiuCuIS9E+
n1sf/5kftFgOdwz810vxjw5sFPwWjAOOycQPWVbVI5tra4oub81ncwkgGP04bQhAI0Ttx4kjS7WX
Fgx+WAwP3A62fx508GLmkf2/02v68olFZPQyMmbl4D7fqvommmUQ+mGTQf9EpypfoLEEQC1+r8IG
SbE3Cw72xOfZXrzejbtAH6422UHIcL0X1VcZlWb9UvvuMd+7Rfept1jJUOxKvS60RSrznFOt71oR
Nmsa8vhzy4r6AuAjL9kSMU3fw5i0/G8Lc6pSqgHzzPz7sOICI57Xq2QpZCMbKTNunGytgko1q1Nx
Fq18X7NRzAJmXR8VoKT4F5k4hI0zpA0WxdnSb8HAFir8i0jweTesTE6pg0/TAPmoaK9d4ED8dZNM
GPGQWnbKyZ2/0CxuW0/RKHjgDbdI7OWagHRZgWFzKuLREk9BpWiu3DPd2zoXTtX+Ht2T30YI1Vy0
HI75/9C1O+RMNjqCtnDHV2XX9KXsyBqE6PmFo4mLmwV7r3YOwFAQdNtNMz6DJAImsBe7KUwZxEX1
osurzRoEQ5qxqJYzXgPyVRLSEDeAb9HpAMrQ2AzB0w16V5Qt6z/kaI81x/kZDXkEDIq4wZVt2wFn
6iycQ/We9IeWiUQjT2E5IRtFE5ZCBDNdQJxNgxqWC5TLQUlzkcEPLJTE1EJffa98pU4S1p1chFlz
uqwijtjAuv4Evlkx7Oyo89m3KnZr90Zv1l2EzhDDOy+jhQQC3d3V4TBDGAIlrYhvQDvmzEqpApuV
LaM1qIt6ZGbWx4bRGHdZnlbRRsaKKbHfSLzeS6yX0ZPdUgyTN1ndlwI4v8ZCMSKOnjxFL63gmovI
0KUSFsKfj0lJW33w7zn9F+Rw0q61RzV9VhpGNAauXNel/0MyjQQ9icrKHes6bJUml5NlvvVdKwUC
w2jjgi2IgOVHUtlfANB4gHNFbn+ZSfj2Gc6r5HOx/A7UzFl8+WGUP7oBycf5SgP9ls43TcSuwjAs
EC9WBk6mpLvj+GHzGcBJIwyZebLPUXSAKZpqeee8CcQh3huLKrawSvUVR3y8I1x5hwfWvqqx6ax2
CgnSwl+T/KRRILA1iRmbEI8CXCWcot8AkN0lQlZgVlUHSeCJmhcPvOx3s2dISIbHmUgoi/2yTz1A
Z4iv1USBPyyB4c1VTJ6iBGaL3wWwFjamAiNj4riTUyZCo1ShDNWpI9QF2Gjlw6ZFYoS5iS8Zfr6t
2AX1gvYPqMGTS7GRvjsAGvIt87tBybfg/WErm3025/odLx7UES3ON+xMHG62/3mZ5p+ij19miYMD
CSBum0nxhTeC983KFnxb0dbAnwu0xRTwCI6Nxng+SNLB7Y4YHl3idIBWyrDydY4SxKab9VKZBSG5
1VdwJGlAwFKVhClAw+jWB5XolK1azBzH9kmuGFQoTBwkswV2ckVN904j7pZxwFWUozaLbGFEoXqR
aevRW/Sg7+T468/iJEz/lWp7EwsNaq8djmgArF0zihRKwAEa2Lj7jvxeHBAva5AgA2dBEP2qBB2A
BQlQPpqJVo+9DZt93nau9Nj49QdbEI3P9A4CEAqaPx3T7VaLJM80GCLaLaGmQAAnew4RAvE/f8oi
mt9nfK5h8Lx9lzRxdZdSE1HPLhm+q2fwnlPJdztyxYcK1vsQw3P4Czs3fRgUTeTyfGfye3HR5jSh
1frwvku7QEck9/LgssQpJ+5NDqHRwow4ZHagTM7LtIYy55i4KIb4v1ytgzxZadarWqEcmEn4GCFQ
JaTd80IyuvgbAs3PTITZMpKRW/pXvbvMfgdqVZZC/tx2LUkYzH6d6CEFz3FMp+3+sCi2hlHGF40k
Zo0XhNqmaW9LfbXuYUR/yRNkjszj1M2fSAKUl/CpiJE+IIq4xQzwK7S1J16bfEdPJ6ctM5TFx7UG
B9Xnq7TIDtHHRLwMdWNrzb2BOuSBr7s1kv4HF2Fv5vSTQxNtWU8RJHQt+sdbwczsL0FrcABXTkFD
4ZAL3/YUw4Z+f1Mj9V/Ei5cQRMADxQAuKJ8yssC8o5uDGjh2mjzOC1TMS2RDOYkhjOVH0+er2hpL
2ybLVmDnSg4qj0xU8oN9SLqhqfFAVi8yi9HlREmShkxl3mxu6V8c86BKbRlS8tQpnk3FUfYkhbD2
odcjAh14T34+TOHvL3+8Seko3d/aEU/9HnUiOxquiMjheHN/cuwhnSuco9pD/rC/LpbBVvzF4kyZ
PC0cuU30mPOKWNl57vsl7ZjJAFS6IbL1liy3DyEERW6tkINh6RNGd2ZCH6AMINCuUNjlD5O+Sj+M
3c/hKWLgFLilx5skkhQDLZXPn4Is6wjkXku2Z3F7DjG7uk+YeTCgRQ3ZAc/gcIOnfIRQiHlJel2z
4TTbvEcIP1dNclQEp7Urk5BGfNquYWE1ducMBuXbYVuJW0iHcsnpIzEWLohRn3fCpsk3k+7h8jiQ
OzJQk2jw83JHfQ+oGWbrQSb1n3qw/uIUfVQvcG1iZmHCut1XzJepNnRc6RrZqgWw1cKEH4VTMXb8
SFWI9VFz6s0r9KXlqLEso9MHfZ5lHaQ65Ze7KHNot648e1PKITHlgi2a1bk6K4YDpQ22imebaPP/
UJmgZQLPPzXVKKOwwNl1RJ9L+GOWSzn71jnatY7DErbA8XXAy90it9KVcuIj5OdZUo/HBl4HtbIu
0ge4w3XDf3OQcBXs9JjgLzb0NBzkz4ZllZBbcqcKTCEza1FbmWIgAHrqhgw3e16tCINA2DX1dr/2
l9xVT9bOnKoyyAhW9tHjCe69i/egGcsnSNri0WmdJAaegGTI46Tneh2hOpQHIeNp4yYXVQ5xcvLS
zZOJJeTU+4S8uXrNvqI6xOHXmbnjFuTCQo9H7/hQauA952Q7oLA7qtnq3ccoCSlI997KxGTk013i
0y58xdRlhJ9cxKwfnPQgqXi/KHabfU8X331uRgd+B0Deew0f0j7gOxgAQZ75g3CqiQEKfUAcpVm4
cP63xJzI6yHRf16T6+OZozfHmWjVdIPghGHs7+OF2GK108YVLI9TDW6Mc6witv1urm93DZeG6AG0
eNHwxf5VKYmuti/GXKmiGxwtdk7lrB9tXQtPNtTzxc+/wRuDZ0FHd+XmmJ1FXPZyRHuNVl1R8eBN
rfrLYyTmkAAAlL0G/SuBkutU/Cncb9RxahFoUBWXaR9uKQow2qaRDkKReZcnIGFv3kmpN11IxFfj
RlQLuL8XzAjaIViHJEdrXxDU++pJ10v0hLO+6j8YQ2t99ySc/wu9Z0iemvAQiF8cGG+oUVRMadvJ
G8xpIl7yaA+xFiNbiZ5Zv8AoRYTZb1xeI8UebXzn7bVrHEU2/j5T3MYiQmw8voevVUNttH78Qig0
eNeXROicQvxduNCwVXfiRg5CLAPxw6l5dXoSje4FThIhMRk67cQoN2wMTpaTcv9OGa/Qd13KNB2t
jyaHSJwhLVEY+u0Bx9h/5AKIgzspl3nNC+RkTKiI1n6UIwFRuVlVGgGOUK93kFFDuiofCJ6+nNc7
Vv/PA2hVYX3QswULPmYgbLu4DJ2NE2+FO/+MpWwhEpxpkyTARXgrOtRIrdElGZwjrLLV9WV5hLVw
68+0/Fkjf/Dr79dPDKkISfa+0DPhOHX3nNUiqTFmVzU7I0RcLQnLNCNonRZ55YYgw9kCPDqKBlbS
HGoe/UZCvzVD80OZo3QtBwStoySXmjqgpS7g2kD5Yz9dtZVx9gKTr3WRhPSMVKy4bzz+qKzFCkze
TjX1VviTjrFpYG3xWedZ0gJ5TSWOBoJX9gm9vDa4Of33wGRWOn1i/rFOiggsRtTu6gO+Bz2/GQf3
DXEHFoJS+qnavRxU7Zu2dg5MQTLTfgedBR5J4QMwHj2lZ1ccLLfv53j+KNMwrgA6EZIg9xuLKsuX
hWsAYYBvlJ4nhGS+slb5BxvRDXr0SEKe75EgiYyQWEH/gG02hSq3l5rY+ruzBWQue9qnca3nkQ8k
s1bwb6S+72MJdVbdY29Dr+/oIgz8lNWARJTnlIuRKIvaqfC1pdcRRaHJD+7RVybWvx33MrHoqqfV
8E4GqTDvXPDgBuuavrLxcnaSRit0YXmoVcdMeogQYu6yzi8D45BK9TWpC8dDuKocU7OvHYgjQpcH
r+lArA1/XQSQLPgeSZR8q7irX0dcMIt5AN9DsutMaAGi2uKlecEJ7Vw0MZMTtZwcSjtdkEe8XXyQ
cgAUsz+U/KXGy0ugmDQtAn6nN4sv8q3oUMRwIWu3yC74cU94PkRck1+t57t75YsFLwLl8QnNMYdi
YBALqcb4a0d5vupllckouy8n/hzXm1aWe0LS8oONUvtOs8XoRsniYXe7eCbMLwsAQvrMg6P28w49
gx0aOf+eTlykLsilmVJnVHzSTtoWMewKklOdBGg52Ju9oRDv6KGLGPi8tCEJj6U9qu2ybDtbT3iN
t+gWJXNNF0HFQLvAjlNkiAb/K9PobnoPPKGVCzuCOIxV6u8zNv2K/ixoulkR4UoN4N0kphD3nRwR
aiFs6X4wEUG53ZdFgssdR23qskMUiZLs0WsCyY7tK+M5j4OO9z/v3qbbJfdw+G3BRxsr6GkDegpY
qUgQ6G0hRCz5gBqTTGm3CQKquj+KFamO1lc+jv9CJkX8DlNMLio6nFcKWnyyBJrV2QAICd0U7yE4
zX0y1AFfMY77EFJHwa2823/idfG6zmGjQociI33pbqX3/Qfyc5wMD9h2w3w2LvOoLReeS9R9hTo0
UlBzqKzaD9jFSY9txptUC7XIrtkWxNabaWT7tVxKs9t3i5SwqvciHJKWBmQ/fDYJ0f4hrLgnp3K9
z0Nw9jmVdgMu313ymJdnr3eOnm4XUuF0qy0447VU6YLLobXh/2LJSazIk/tNg5M33aZHJFM/JIk4
4VHY2NU6+5Z/nFev15zi5ONPKYzrSZlAiKlHk1eSozNm13WZtjNzcmiMrjlX1hQL8HzLfVSwuGQV
PH8xxlWZ6+1F7TDHjeBq0I4uSp6Nwn6alfS64p20bvtqnoKAtbth/XC6kxK0tSTcroPAbIy9yUWP
+5pl4SY6szvHPpqThR8XdmUylOfkLK9P2vwML/2fza4N68a27jM6AQg3hMbn0c2fMmDMYCZbuyef
JwtUdWqqe8ozdZRSifsP14cVkVJomuH8C7SczquJLrSFG+hT7P0MZRdq87IIe5Ld/Q9edRmADuco
rf+WYkmemAybPwlkLTIWOV2TY8tPddHALz53VFzdeOaZDaTLamCL9OMQCbOkq73Xp41i0AsQohkY
EDcy8aGZFEGYUAmFvAoSh6/iij5m2cZZ/RdtLIH52WRVyVf46Zw9ZfYy5tlF/qoqNrw4dZgbw6kO
HLDYd2Mm8Hugoft4yHhGOqQF6Qv/pt/MoFFSqEtFGKRuOmGJkyRHKPRtS0N6Rt6Xyp/RT7kGNxn9
OAZuA5my1uCxkzcXHereqWowMPY8SLS4TehJf5N3MWAK7Chr+wcsI2uUb2miF5mO8itJxM6D4MGN
nSlbYAhygdjlGrVHkWlbze6046+TCIoBJKBrx00rlORaXYyWWF3nM4A9n9/L+FA73KQkZGdTOqvY
wn/YXLoE7ahgUgkHbzv8uZc39C1PHapFRg5S1FC1IdqqjyXAirfxwod9Rj9d9wntJDjyPkRwdKth
O5pGu9qR6QjmKFjhl+4x/bPktV7kSEQQdAM/3F++YLAEiwvwwK+WIlP/I9GLmuj2YWRyeq/YHtTL
qfoJyviQ73ikqzyTT7iAYVtK02C9c4CfwJkNqw4/j4mbVw4rz8N/TRvptoT9X6M6vK07dGGktz/s
KhUAlfXZSsn9mZjHO/NhokrIQQpE3Ckm0KB3HXtXdkBo/Yh/WpZfhCyBKW7bXL+oyLWFspR7kNp2
VoF6nF9c6xDCwWUgKZYQDwPcZ2Mutdy9w9QoGQakpDh4Q4DPVPNuK+Hg9qb+09kl1IlXY0iSqNx5
o+eDfjUraoBzrLrVF29MqTZGGuN54qzL6EQqibB50mkgmNqeMZjxqrdeUu9l3Me/iZ7zNFYd5Ije
mrVQ6VY5XKnHEPvp2QRT0cqEv3XSnjyNTmQqyyVWSw49wHjRojbFmtksWFIrDi0mv30BrtajozEX
Tctl4ep6vb6wwtORb1jh5cEU6VDQZByybtO03Yudh6FWkKNlj3b1eKpzecQ6ICNIwKVVuMdkfADr
JcHTDhWI3uYHn6JsrrutWqj8eJXN8puUe/RsluAYUmM/a6RIQuPuHT7A/ZxvQqQDRvY4GsS6hQwg
dzBt2oh/aKfPoQ++CGlhDQKFqD+Xk7yCEobra72+vc75+BdpbVplYADXX1grgZQMDTH4PFx6qj4P
jBXdvJ06aXSi5YKImSkj9BSEw9rj4xHy1/eI8OGAolYgFCzmSlt1YOajrS7JrU9z347tfFGdvZOV
EhTIA7+z5d56Ty3wB3fuWSddHi1KlvdtORrMvE83hwsCSKJ4444ps8oHgLl9rNoSwpVoxaYiTk5P
Gz8LJAVGDgTemKNuISmKGAr7xYC92Yv7tnJZEGQHWA0DGonIfWum+HUZ16YUs+ykeV83KyZ/38dk
K6dQzdo+CAK4KaGyoxJGjvnIRy1n/yoqwXB/MbSwS0QxhkMLrDqxWeF+2ZpRiJAwN3VWy3O5wr7v
qs1weWBG4A366iZxEAyQq2syCu7aiqO+SX7kRhIIHk3iSu8RdAFlNb0ZmQbSHtwoHG6tWrb/ObjU
9/Luj9BLPXbEIPuWIOhMPgdBk6TSW/n7P3AM9JixOu5ryxlITFCmSDd/cnmLrPGepsOhZQEY8P3k
GXVjHGcG7AdChQ+fHG0A5WqwR1U6z+6rGC2/J3nohHJOtpmME2/ZmaaYzjGl7RqXyyWazvtdVejQ
3lpl1FhFvh2l/XrTwRQlig+RBSmNDpFXpbpKEmNz2LElC/rPyxg8+ynzPQ97Ly9Tb+dqQluuDyzP
hMBPlSZtHcRpBVmDjMXd4UfJ5vuii0cezEvd+5sqSRA7nF8iyWOV1iUNOT42+wQmD/lyDTpvX84Z
CiUsLFZZo8EUNgPFGNH+Qbw+yMvXA2XMHXtNfSMa3yhjgiPCrjGGDPzS1yINGeqVEjBk36CPAjdy
4NjHKT36kQZ4jH07rn99+Q/rO9pTIzBTEiajFiXiT4V9T5CwtBTHbD+lrYC8zVZv/Y5fALdV9tS3
A/vWJfqrWB1GiOUBOWYvT0VUGAyQz5BCc1Mdokkzow4jMsCgdRvEY3jglBOI+spxYYhXMj5OWwTc
UaLtIiB+o+7IJwVyPfbY4+l103QpixKcrzUckWmQtJkzWnyN7FP4/p7ncNpBfMerAksfzGLqdSVC
IrxodKNWs0oNrRwhyzftt0m8i+DN0SuAUZnF+wlLHtqQBD+61WuSSK/Z8QmxVzsXC0WT6sJ3p2xy
2CeiKPiv6Dt1zIm6i1WhS5hwMI5j83wUAGq1cfw2tumfz8mDCgy+WPfFUfVLgDVCia2aPaEXYUxt
eVd9nqb68TU7d/ms/sO1exreiauFwfUE91+9IbMxDTxWWbBaJ7Ctyb9TbF5GHbIU6uUKv68gVLoy
eEb51Co4OUyQ0rZn5VHE/eTnlORciFbi9gS5DpmFo1nlS5w9BiuICp+96V+dgk6BR2wOlk8gFfJy
XoR6KlbgHR/VvTl6iSqgNXnQHs/MvBsnS1/wpNVRrL2wSABU5IxE9N0q3SgPS6IOVU2PUk9CxXNE
9qw6SS7ixgG9rdFugl3Sh3jeIW3cmPcY00htvu46GlRFhzQgFJ8awPdNgcBsl6yCFUJt+DYJUst7
0ekH8Y/sUJqmEO0dR+aKuYfLzDpVn6COW0+P7rY4tNlDhXGlF1lX6iEQtauo+BjoQIFSWpBLV1tV
NvBikOrEq8RUVJ6hNZW/qSoTezXEnJb94pLxnfO2Wcgr7w+bQtj6pG970PevU8RAqGHGYgl3WjVD
/kI35hzgNKQuAirXbF3PLc1o58HMPo6opEiK7RpEKXj4/r6IJiG7rjTitwcucD7fdEN+OCTt7/Wt
Df0QNicWDbAalO4AeSX5VG4yLPyt2gJedh5aYj8E1AyRk6zZm+gsxRmJ81T2xZEOlpLArRGlwLPm
PwPcTllsyc57NZCP1e9DwBrNjrAcn403nvD+KIAJoXFachzwXiRogwJHbcUZ7PXWCrODuMcirLyY
n485cH8lqsiYda9hf39VRNm/MFTMD5L1ce/wZ7J2glkB8MtRlygSDWiiyGifRSh8VQTZP3iu/bsh
PwI9nPm/IMu8XAB6kMd60ITRC6ZzXuUw/p1GcvoNpYUSjPPF4uAdpx5/yx+rOzP+X7brAoExopLe
irASXR2zQjJbsnmvRHV50SUL76N2AixxWchra9Xf3VgJd44ANzqGzdWOaiZkwXs22YaNcb00mgTs
Prxt6OtvsIkHLWKiPwlYo1zHGRerJlW6kzGQnyNXualHpF6cCvbheDLusfGdTgiP5FnVv/ch6WVy
eLwGvD6Ux5Yr8iqt/LhyIWCHL4MzBpwr0ca9QY6Kn6neGSjODhdxRbIh2/KXSR3IX3XBkJj3g5ou
VVFPLAL7X/VraTajiBowKnyzBp708cpnAXlBK9N9I0+RTkemEzoUYk8VZLlCU91FsreXcVK86x86
UUoY/i+xqVN4i4FZLP25ezcVxz4p2l9nXV5TGzNSsfGMAnHFA0HKTq0gIzA0/qN+EK6bvEIP/5by
nDY61JF0OdUqkF/+iNzD4Z2wsX1MNUAUEQJIJtPaRTK0DXUFELMccm3QEkF15PpYGUh9HSQcyXN/
HpVa7mLfLFFLgW/QiGKQRnCm8WsCKtArGAW57HdMO+INRKfrN5/Dnat3fSCNBYMqgpx0ucpKZhW+
q7QZkaV0V0EmHUn2XStbm0EVQXIVfU01v79D/bt77xIld4lrKBqspZ7MuQcIStizrU7lEnH2T3oA
YNbl9h1oSQspcT/Cn310NoE4GKg1D2u2+szavWA11494YmDM3OfQefJpzJ31Ai3ateqQ7pOxpdDV
I+ohMPkoQyPAKwDSTpPDO+F58U+0Y195mNwlEj2NmzFTxVqg+c1o3cmfPZbuiXT5kq3IS3HlSi8l
Scx/CgSYR6Cf/YV8Vt1fFrfUlmLQOsrOOfVOCeHF0ZwVC7mvfyPql0Ccj/uJHDpjAv6X5ydgU8I7
WYXnnYREQzhKBZdrHvR9g6EVt6ptuyuey/YutKDvWbFx3xY3E45XhuTvOZzQ/mzbn4uuJb70gGwB
IJ9KZoHrbD9I9WaSTcDXZ6Zii/8Ab1vGydEbAxKAcnFlQNEf6hSCI8tunqPgLXXzlkdo+wv6fU2T
ylnH6X5slPX9oI9siBnPWIz/voGqyDnhPnfBvgSzlzQ45i9UtxnNZacq6LLtzd9zIYOGKk3a6q5I
oe0GyiNfEvRh+w3xOpyX+eODGA9on+5dNIsFIbkzMXmmPsTfHmNdMQP6KBdA/jnxjRMPfxLZS845
H6LxeDMcTZXQQ6zzJwGTisICz/rWayeEfFeknn9Koau/Wh3x5kUFfZQpHbxmsv1brm8tldCzQToJ
vO79s5hbfpZ4MKqViAEMqBko+r1vm/3PqysuSwwuaha9NDnOxEB+aOByPcMAyBE8Jr0qNUPa32d1
XYS0hS9YArDSMw95Es9WGqvhSCvBzcNppod3QcJ/5o6apAgVOR53NRfQ7HzY1fp92Lgy3/2hYDQV
/oukfN1a234pKLLGdlgvp35fDIhgBCn0sZBiBNwKPK77n/2cIEuA1kIDKS09do1EMPQc0W4gjYiS
RXHpYa6IPN15ZPtsSMEemwlYk4YPG5+9OuJc5rupgxtrv3jVh/1yy5eL2o8dzLi9CPLLDIIPHxUD
GpvntCs3qJrXnfZVyyHORi4qLKWDpFxUnfs/DoIpz0gzKtl7ettS4lvpM3c1Ukdp5BLZkDkYf5pt
6ZsupzXLM07yR0BW/X7O90r6yf68I4ztbn50X+FaJw3Qij1rpdmPklxuclbBb4lrMhGUuXOQIY6o
YrnoOeTxJnFAja+Sdw2eNwqziMYAOHoUdkyk8f4siR1Wzh72lktgJJB6iC6JoEUbe5It73CknsKQ
B+mxqV/oEKMbWsTtPrnu6Y2aFLbJrmm2Tn2O+IRH5pXlI+qHScj/3h00zB6CBrAQ40QLZJeIdq1j
+7lEFxUE+uz289PJT/hDBu1VFe6efMNut/8kGxKQ5qom3Tt9ptrNpk6eWZat46H+nUhoHjyFXbT1
w0xRY1JCT0/Qwh8ftUsYM7Pd+kg8xR8ajpfZB4ljoXSo/+wCbJRU4GfKaxoWlkIjcZ+AnP35P4DE
V6xkicRleZ2+5C95OS8VIAMjv9Su2PVLWRThkPujVLHLn8ajyKH6JTgk5NLzo5fjR9ot/jGYm1ck
01ARy9pI/mT9BUctv75M58Nat1xKPYRkYIbM7zO3xWkbcYqIMCgOhs2hWLbU6p87bCar/JLfOlsq
lM47O+H+dPlK0mARH0hJV1q+feXb8WrCERpiP68qO06d1y35BPisw6NgqkVlQofBLKdBxVaTBtKh
qIytR49J5S64Yx+6CG9AqiXBYlfwMyKM5gdCAVj3/faEk5OByLR6ps8SNS2+BilSIoB8RxA7MZW4
6xQKM2jbMb9P/TXme6o0XQwZIgeToVKM4u+/GVs/UYOwl/5lNiehV6mP2myJpIptQXz8YyZbSDKV
1g8d0wu5cHeZk8bDDknAW93sxad922OxPdVc7LyGJ8pVHRtQX2juousDiSb9SdlTnZgna92JAWTa
24Z8SYsKDEeNXAnK22R/uJg1+yd6A5KAzwqLd1GUH954FdG3ZiLOW9YEZLEKFq621EPbeTqTkuGQ
ZC2umtHd52rj1q7jhLwayCf+OC+BOi2i1Xl3z+UlakU/kq6v9ksmdvxctpuPB/doyEFysLqALxDD
JaSHJ8qlkppHIIv83ueMBb+VwitzZijuJ3R1O6lJuSjWMYOUqKsb1ciFNrydkufkZE0NcPv/HYql
CiWIyT/GHMDBDWta5rq0wBIhHbM+JsYxbvWMoAuf4zJegnlRJeSsnMasYAqqj0HCgnyvRCJ1Btz/
GdpIF0M0iaNGxxsqeBC+HJai1BChyB705SsEj09vH//uKGfKLJgXqxj2lAwQ9Gwui2dvVLX4fxc5
Q1C07oREVTnbmW2dCYun3E/5lm1pIN/PvelQlrrER5QyvBMI1c5/RD+jNy/vhu4hSMwKAF1wbIoI
BVM/W32xY/Fi5iWHv/A1f390ye0kOpGuy1vKZMpmXUYkCrvi2c5Sye5iGWA0DjLpJreJS5DmAAmr
jOgyqHdhC81LtOZ5uS0oPuANmHgaL+ZHlZWYy+xZYOHYpKzaCO/xJhykv5TPM48fDdmijG1pfQJX
hCttraSadRlXtLvanNB9VPUTaiDt48KuK8/SPx4QNbYSKO7DDIzKPPIbdIGqfrFQn9RAWqEJXHrV
Fuf21KZTg/isrDVHDxOlthcMK2vcIkCJQhP/ye6ygaBCN96zXLgBZguk36dbCbumFvgEMJ1r1uvW
wQywNerXJ0JVls+VZUxyhtj5NkjhlF1001TbTYXoQeh9pi3wItqSY2YJ7osu/KeFuOxZDLH0ELQh
NfYCQ2zfWK009IseaCmIVWgQOQtbXe8t954VD/qqRiwh4nxLkTyy0QsXzl6XmHZqKzH1D1zCHAcn
n9RQMIvG0fc4EwtLc/BBTzQ4VsHxdQpbq6DX9Xm4so3ge5hXRh9sDHYocn/y0hsk6OcbVMkHkdax
lhCf+SgqVuaMl0qYKOVAZiDORyFQSK6fanObwkDnsq3/QAY8IyAAKweSKxqBr/SUen1COS8WBdAc
pJLecmuJdE514kwfWLts22hA1KtPL4hiVCi6tyHIpHuBFll9DJxdt35n0G+2TKJLVFJrO0flSot2
+w0pTuAjWTaXtq+Ve4ZZrnbBtqfSVdZvLY9YOhFBZdx1bOF0GJHR/SQb031aF+Xpi/ncPloxwfjz
lBfuZuZTVDOZxhQTpzjkvf1OnU20WENgTPvK/ps019TdAGUBZk1SR5DEEIhqtJjv91DqGIRVsJ2p
H2YmnHFILpVwv5eDjw3MdpBqfzXBVLKW6KgeOKK6UFTGFmNoC7f4oNYenUtpzdJV1v4qmXgbXcqF
1bcyQ6FacnshWSQL90x0INe8B3uENkLnku2oMF9uy5P5+iFe0gc9GyYNTlpBaMJ89jQlzSZWVmBz
YTAbKxUWtyr+f+VEetcp6zHkQW6z8aigz1VrrrNsmzvIvviKVSl4guyf7T4FMTOQGN/Vn0E1wvHl
4qRN1F77tFwthoJzKBuGdigg0BOXowLGA1rrqvj8gnSvXYOILt5x0XsumEL72a3qp19t0PCEDTxt
CxsG3XRT8F1bxYtohOFMeswWq/ONryTi1qb+cAvYubh2tQ/WAdUXRfaITnSNNnLSp36Tpsdmt96t
hinBYGj9wUR/ge9riAR6fF94g2/IKWYi26NE+qprEHWH0OAAK6zsMhLmc9jVYb2oPaNg/zpnBzta
IGZqFT8gra9wW9mG0z+qb1now/5LkhflPBFd8NAIQwJNorWyv40ohKGHp622cE+vn34WZIz4AKSi
J54rX7vqBQw4EOrxY9lUS6ib8KBQ4teo5jJxcNEYPmOg2JO6N/7ODmcywcwKLfhz8ClrKuBKNTlv
An654dRG7wlplZyDU8e5NwnslXBvxjD6EohrTXX4f3TG4sOc7sluLp1jiJUHl5jZmvYF86O8cq33
p9DnKTnctNqlFueKKHe3Zu6s3xmrTzofqA9h5lYRvl6qf2tVlIWoB0UwdIA0kzwxGby+Hk/4z7kL
j9ClbzM3fFUnX0tfEzhrI77QgIWqldXcUVNYH5UcO3W6TPEFVL0RDAYeG/tesCkXVKKffaBbQULW
ftu707VD+2aOpe727OiMsWyZcIBEgeIX6n/2Nq2pGg6/U8YVUeoE8VEGOSHN8Ot4y6ItiVSSt1F/
rQhazRR/Ki3F0bJvlEVVgDo6y36DbPcS1vLWno+ITBseJvPhwHIg3/8JhfukJKkpBwWoe7VIl1kL
nB+ig0l/u0EjMxp+rc8SJI7kzadiTtxix94utw6Dgu+AUoL1gt2+7v7VS/HE1SXvwX0Mruux/fwf
hrP4RLnFYGA8r+Tmqtp6hNO0UbC2Ngq3bfp9t62E4tmSt+FS1+lxYouGheoWuPkNuAYIaHEj35Qf
gTnlbIdCkoSYGYST2JF3MkFZ3D73xt6KUqs4AzUOFHTSqe4F/WZ8FG6SOYkGnJm0bIyRu8ZQIrI1
57aJwT+alakI7W75tc8MAa58mzLFkBW9rDI9TF97liUFA2z4OwzkHQgVROErrO+/USuRTGaLJ+m5
1JRH7dg5/hJfwVu+snGyLhgEvCtpdLf/lmf0AssBssgVWmgHoFoo0kIjo5kAy+kK4UmBO4P3UHP5
MkVLplGilcvHWrKYzq/XFuDWhnjz7ZbS863WmhMaJcYufqIS0jwLSx4Nn5YqDYh1Q17ZzHW3cFgr
a7ZzuBZhGBo+oVnxeAUm6Ao5fhHx8gI1z1rY7zXL8lsDNvHoc9UY6FhRdg4ZajfYVXwb1XTd9GLf
P8BVvFQaVEhXsVd+dma4AM9oL12ODjVyShQhYcs1taKtJN9kZZ4tmxxptQX2DQHScqYUtE3m3YnF
51dPf00hqWd2Wo6tLGg8Rvi/wNlhp98fL81RLdeToZcAT1f91T3ZBEbE5z6YDp8fB999PGrHwOM0
mtL4SVZWu5bKrY6b5BR1QY2KWb3E9xHx2NWlQJ7lAv4M8hsCEs1G2bLMBupf4cpWD065Dfo1l+4i
urLsSUAxAKrGGbo4dFs8AnOElM4bXY/W/KGjA26OukLy94FeHQiyG51IZB06lbNZa0J6WRvNrCko
ma/zP5RkLjfiD/vsYjMbPLbKUcrLDMmHkB1dW15kSAg8unyw9c3LjjbeR49dAzvUx55iFNacFqH5
TpLG9XIPDnSB0QU45KnrWljFaj5vzqG3AIU+gj+HoTV4btExUnOXUC0H1kKnuOJoBi8aNL5U+q7w
IEytNfHjQMs/D5xTB7GnkjXdTtuuIs9hFhqyfWsoyZVuA13VNopbKZB1kDdGACr/1RKBG3DLmMPL
6nN/+TDPWZrZfjG7wKfPeHBv3FmBEYL5+T6W4h5yTrx8QFfgcoi65YYeodxGD6sle80k2yiWVdel
ECoHPIeYhI/yPFAX/1rQXOUUw8A9USZT5nDm+MP/3qWP12cvSheAu0uGEtfRwOxA9ZVZjKJJNUXb
r+IqFK2FdpCKPwIc3KVQOAOz3I4PF87URldioytKGWtDxVuIFP7ow+5KFu/5ZXI8XARcLMgC7oSB
8cfFhd4eI8/iq4fp+IXpAakb1V6MMwX23UZ5uon6hjb2UOiHoSMNVyyT3GdSHnG4Ba3TOhXhKg/W
8WxDOmbaPn75ih5XLqKDm51h2ACt6W21NL0RZQXpDHRueBEc7reZL5gg3ACXpuS4fJA3oIHE7aSz
Kq7kUXsEiOn3OtS3uiaYt4y0kOps4dre7XEYpnlEpyG+muPXPkqLcg/3TEgoiCKvA93QCLwiIY84
rFYOatc7Xw+/gtcqIAcyzJ87KVDegZQxIZPXZH6rNVsNppJxN2E8Pf/+LRCb4QoqtS7jVL1riJbO
03uR52S19uGF5Bbe0anIAoPKT0A/fcGEkR6av25CvyiXWY7KAQA8c+GjUA1AxoU1aU3JykwiC3je
O6yDK6Xm2cKZSUBRjGThy3PeH0rWF9M3YDCCubMzi0Q+H/3AY1rVkLaK0wVOlqm4ggTKvptLfeli
uAk0b+DZ9ijTJNJ/pAPUOwNvY0O68bLXyJ7We4N+p+sW5QrtNUzUbX+tlhLt+TGVonO7yH7ncAPw
Sbsxqv1lIP5wx21dNvr/rHswDpIZWRndxLeAt3dvb6A0Q5XgQsQs5EedZXaddvhNLw691RDLrFmq
HLBq1fJW4YwMvRKADHUUR47L+73NqbkiCSYWolO4HRxUDOWF48zLiSWut5EYHWGDV6jDmzop5Lb0
l5VvC/iEG2yRRHWyGxR4N/DpsiLmNOKSqXibDFhRDQNWIXZDgyPbyi6rZwhcBY3GTeRssOOY9c8Z
NqbW7uO3Fr3M9agPgdTVV79D60c4pTz8Kz4FQLFi8CnhD3OKaclh2iubvFaIzCTLuanBfcIWyrar
s1aX+e9WMloaMJfa6tS4jnfYUDLVvD+1FiFIvIg6BCzOXzqeZr+cyEwVPfDW3ji21GGtKsq+6G6W
PmaoHI9zwVzpkQgmyqgqT7HescAcyIQbLExGvcCh2D1XrJARNwzRTTPaq72huDRpRBgyv1QUWpnd
tXr25KitCcCUj3Ar664oKrEK3u+lr+6/C1f8MhMTVoWPayv1XtDOws/OSJVsV2OTBGGkCZWAyb6A
8WTf3CXZugx9g2HStvqo/uMgbSwrewa+W5Mu6efL6tjwjEf9I+ABpoUNsfBL4U6/hSRMZNEm/RA2
qt32L4dJClGvDBAA8tEyTc2ke0CQ3GisKLP1wQiqkDYtNunQZbk1/Q7VjesAVXa9XniB01iFhkRr
kUeD/7RIEQn8YCi5OB9hYV7OyZ2y58sYEYaaA1Vrig+H3WjllTFmKOmUbYW762SBpkZ4i1LnRp+n
gUbUt2zzNvyt0Ewq2gZ6rOUFumNaPWdsnsB6XbE/zJSfzgvF3TCM7yis9ugXUiNaxyzcyjpaUzPI
+FgA3yytZ5s5iS/LYEqP+pXIvtE0DkYPs25RqKUZKFfnFOwpV2sM14JqrjE0GvQMoY2CPhDkkP42
4q0IMoHGhK8HdQ7RZSv+jKPxKqdsPyZJ4l6o3pc6ggcYb2Vt9QRwqgzw08h3nHE3xUQuqIeYwWom
S5dLVBRlxyEDRfZTH37KqqoUC9IGulN1MOuoEuT4/mbsVA2C2XlxwKuJfvmODBpAwSqbZpiok0pI
Oop8Dy9hqJePwDZoq+bS1xfQHoBBLODCsNlTMJt+pVahLiicneLQMM4mVIrtRfAL1jtuAxcS4v1O
8OQVNtfpl5m13YiOWgABxHnd21Ing50Qt/wOtBUvpDKxaXFhZemUDq6q82xppxXhFj4X6K5Tt1s7
Qlw2XW1t//Ox7RSTp5EkCGGJdn9qbISAeAYfeU06kJmEfhe3iLJ0i6G8wf4VPggOHHT3VezS9uFM
LgJp2f721DWn+iqhRQU9B62NuwIt6IzBR2cjv4uugjjhXkY/3O2LrAwKBqj4hfAbBkuGr4iqI0Oc
RvWcQg8cTXNEZBivYutvGrW+u1c7Mnp2On8sMTiXUFI9KrD0hL7yPkhLlMH3ArerA4fLrYFx4wgX
7lBeOu874nMJdOlPT0kREtLHp0mQ8RE50WQ3o2UR7t2uC4DIadBwv5KydIZ1Mepsg+/MlbQG6rQY
4Rm5RbrCuNUlS0O2uWKzIWyz3SQr8YufzGgGZZMRBPbtOyKQu518ikkcetj6Ia96JtsW9+PObY8Y
mdrfE7zb1Mh+yVgw2LHlxS6avXS/lHFe4PpMYgJirCDUa7axKC6vd+epd9W17ZSKVerycD/CrUMR
UMviZcQ2LCY3omvUGtKvGB+9/uap2gYFyKdU5hbrprRhdYCIQHxzrZcwQ6jg6YK9UkAqPdNq0nDX
DpBuuTC0gW80uEk5M56tRsLZZdf/o7Uhe9BDpYFY1UR4o4lFgykPWvEHysiDkImR069O/qKFvn9F
+10mW3IA1aXNnpsaxolC96UUt+2gpMG8/BMWZ9nrLfRfMDwYuxPIY7Ikm4lQc2SB+QQy5ZoU/YcM
r4qIEzeRwkIt0F9jYGyluoFP8Wn+0ItlnuPnsshUcJvLbmEtQdChYz/r3RF9FfUr0aGX/XWnqzfC
RQEAjtuzDNii37mvXh4uO32a6vhsrWVYIQ6DMUZVHp8SZQ7mLCMwhrzUGkjKRiLV++R5H3YTB6Rt
HW0kbK1PwGmDHMhSficaaIvdr4uvxo2bdMwL7WTkibf6TY349QRYEt1NMlN57Qm+D/zmDBmDbb+0
0M828JrOf7afdUdzSsL4ZlcXOMNJy6ma0lZHtIpTLJp3J1Z9lj1BJxm+M/26u12nXeraLB7UdojL
JbyDU1KyWtF1CNJN0CI96Z1goMWKP57BiqtScTwA3GekxTbU/LWfUQkBE9WNuu8afbU0tyHaENiX
YkmJDnJKiWnG/YLnzhz2zzpA8tzEu7B6KJ5Ut5zw8QqDswBHfcZtU3f/nr9EY6FIKFfE4NjRrWla
+hiuU4dkacoxQ9a3ODEds/wRT5rXlM6hvCRUpkqba7/SjBYmC664VmJYVVC8YwEu0Ru1pCYJ1g+l
IAOc0q3PIvbbM7Xyt6fDcXnL/ZaiNQ+H1kZdLvstzFWTjFrAhVPCFkRpKTm+Yi3dQyWVDYQ28g6e
ccIsQ6YxAAz5vUplRKlvlMYInrfm7myse/ofgU+R7fWU/HHdhPx4mkihAThCSCxePnqMw0Ko13rs
ncOKa7g4jlZY2QmeTGcIoC6ec3e+Kc897+o7ECTXunjMwgxjatOakcbEIGzXWg3qraNlILMuVB8i
s79QwweKyzioTTsOLCQDXMaHQrwI+3rH1OQXW8IZQbDzwaS5RKA+Nw9DCVBcV+JxjKEXAgnSM4ap
iPjN6F8CxVV/BMrec4teCAGmw1yaN3VkDsGGvo+pLXlw13WREDXVxVMRfryVsIn9XBsk/Pchs+1S
yxiFFnfMJCN+zQsj8btD+ss+AHpC6F2AL0TP3nDJb4dQFScCejkYjlERP/UOPI/Myu18tWtpawVp
lwtt4mcG/xXpvTK2Pq9BiP9u9m3Km+mAwEeNVF4sQd3wAV9l4niN/gU0MKJKLtkmdzOKh83boyLV
J2VglLOf5fEpI6eWUj/P0Kijc0+WrBdEYI7y7yxA9fRtGi2pfXcfPZx+OD1CdzCWs8asNeVE2P4o
PFP0pxBDwZaA1zs1dFFa875D6aFNpIhXdp4chnM0haBTZ0rXDY/piKSMD325UHIuTMf/NM3j8dMF
UsJ4iEn9JlRB/GiAUMbGol7sZ2u+g0HUGHoy7x2wNNg6NCUC7gDcwHHIMOQqiVuoLncAab17z9sQ
gGofabegfZuNSy3hsAOHQvk0qqsxBv+cP0Z5F6GI+CJwfv8pRIpUs+l/6Y5MAWGkkb/DlyfNo3Xt
p70VnTndQE+M5IAUflCEOzD0Sb8nDdvT0Odk1rbg2EBVfRI0CkRKdRC2UM7wp133jOLUcNJuOPdQ
VN/ttdKpkej24JmzgysHLvzW0ZtXbPa1jKyzItEpT8QyCioz6Ov6UIUoxgIJUTtki6ldBdxcY4yB
/mpKoxI+4SfSxaWzc3lff/D+cHoWMr+dfBuk8pMG8FapfwOx5cqq9CqOheGBQgcRVg++klar9pwm
qU+ftsszsunxfALQwd10Y8snozstt/B2f6xCXAIQS2aiXbJBMrYKk4XMzDl92RVnyN8tDFXIsoPj
TQ+P7J7O+2DLua6ta/0CihN2Q98oYFaRQx8iYZXt/lTt/crmH1R9O9gPBfUoZs1SFVdrpupj/yth
cglk8wsauet3qu20PmdJ7msqqSJUvI7nJ2M7USmssDZTXh8CokndPPVyAB7qiDZ1ClBYwWW/p644
RkuF7ouvmxJMU/+6AZXy6GV/Rf8/u3GTnY2z7BapahI4xzu5+ZHbVzgIuhOWZS3U0gliRtvDDHYV
8PVdo6PxfvBvumFndbFko53R8jdUvV8AnYO2tYwDz0ukVA/WP8YwYehEKFIAUNPLy7VKTqfWjaSs
cdNl/B2TTEPw1UAOGBbotXkJ0PruXEFZD2aN9f2UhGivbnon32FbDkDsM1sFoZPlm5cSalK/c3q/
JFt4Dj/xAmIxkArijJCXm8V1znEcQY/okqf6LN1XMrY6GuFqMrmLBYjf9Mcq9a40DI8kOTEL2Jl4
17pZl2CmmuggpWGzj12XuhklrvdwnHDFMNb5qB3f14cyzcI+ZLF/e263OHeJkOub2rKM7nYVW8xX
POOWH4wBqUbSSKjKt5rkQ/dm2a4FY5JL8CrSrfwIVWTw5p+Jr4csoRrkdSnnO6Fij6DFip0laTNl
18tgJZ6kRGkk2esTKFAB6XwRYMlGo8L25wwHC9yO/VMgp7Fkdl5MqWllWPzcfrPkTgR7BqgkHu5x
KBk84oSaV9zAfs5xzQv1Wf9Wc12ZKSoqP4iqnAf7oumqcmQfGb5qyY48vHwesjZtUxM9foh5PyBA
hAs+pI6icB2WbNAsZH+8yN56sU7PPqHXlJqOy3ZPwEZkVy1114qJFKSq0AWqpbwrEL0PiczbIV8J
nUaxHGq+KLDG/zmZnVMuOPpa2S+Cf8bMg3g5BB1qnnwJ2/e1i31rOD/92k9J9KIYYbKb3IwIEFnz
yARaksnRjHqxqvYH+huiYtlM/vc2TyrQPIwKq5IYlhyU2/hpiHsIpiKzaQT1fw6LOtj0lmZ7nR5K
wQm4i7uGLYshsWwwDQUZR264M5dQc4VdC/YlbxWDSe6Ficg9GbvWUJkWoBUEVXCFiET3PZukCzhe
tA3bjTTR5MEnn88jPlynRhBjYdpx/2OQv4YjSUUW75MYHV6XRTyX4j/1guIF+QhobA4CM5o3Gmah
TyzyuuUK/RzUA5lK6+ad2a9COGnw4IpagmKfrj30PH1bPKXdVQEKdI44xFqFikZNVKNCM6iwRXpv
D6DxRfSWCQH2dDUXR4ufLYlRcHJVN73oV1/Bp/ChUPHAoDYvV5k8ueOI40PZ3hz4YcQXV34QpSJi
X8J2X/KAc8pPeLHgZIjF6OsLopnIb1DR17zDS5f2wAG/O3LWe/Q7hs7jTpH48zoE1QAZ4LkvooQE
b4qx5ZXUUG+XbOLI+gEMplK1GdKR1YZE2LhVkdY8ypqd49+AqR0+ScObMBPg5ofb71W3MOIPQQq9
qiFf2H0YycGiMzfTWRIhL+f/Q5OJGoRePioVpu7qKN3h54f8huAlI1mBJ40lfWTM6fK2C1+Yb46T
lFgaoTMLVT0wXZwdeIt+qY/RKnleuslI2q0eo3wDhqhecYpvfWyQ1NoH6sZKS0UnT4AVNhpQDemX
/odaucdHf/xobN0jR0Nz0wl+EvQcbDBlDU7+YPoj/EpfQxeiiz24QXmNHT68nQQlTi/Wevo2QFXw
6WSSdxYBMJYX3TBTbmSb3r/+ILmY9fRYIMXZaREJsLeJKuvjQslHKkNq1X7hFxtsAVkPYVbn338s
NCi0SVY3GHt/d9eZigaQZldUBPwpl7D+30FQMQWAuGwAwq47uwDlqCZedDlnytJV2+4FmEeSMEEi
C3BjA5Q+9fec3nsYqwDzoULp2wO716yUxLYPAFMRqWM0oHfVeIgngw+s786FU+LLwTew7rU8BryT
i+TJ0zZnHfdF7sH8uwIf9IlN5nxD+qfK28/ns9wIg5dC+EW1kEuIbbA5rwhiXqSaVH8+zPSIpdiY
STpt6qN2kPzmZGDCILlNvUdWGaFNmVWYlen2cho0h9iX0Dc5VmGUztHUT8gOPvWUC0lV45efwYJ0
iiS83rxKmkB6YX2IbmWFsWx6ZopW4MEAbl+OId9YdbLvD/udwlDiwvcTdLNKCrZF4ixBvxTKjQT0
QGI9SaRuwV8SwSTcnto6RyBs7PFz0Po0H6ZAxDY22vAQmJJgwHUr1k/Msrmjd9nVQjVQ6cciTsHa
5eymUXgoh309xXkPVR3WnSJ4vjFJYcFFfFptcSEN8Uls8xRg4fOzzakLWq1WeWjdQeTaZBdACzMz
F6xugWwa28w658gb510ej4DilUAzfWZbVIiQ5lC7fjDaqum08J9J7iKg/xi2kaNPUbF6jaQ/6eYy
uxNoN7eWy2vgdah/W4C2SGkRxuaRHhDvelfye/affRJQoGTGUNTHfcDwFWc9M974xLZd1v9DV6Hx
8ZeIsuBWFfyGMHqgjT0Y2CSKy4jdAyOQxig2qux3Ndef5PJ/P/rBCvAqMOFAqle/1vduMUsXQpfs
xMGJ+J7w0EduCqg52DYbntr3ofib67PAdD2cDuFU3+2CcX5TJcGVIRl4MlkIGXGlahEVDqCocXmz
9g80qKZHRmd8e9ua+WDdCwAit12IWWHzPRW7IPu+J86lY7fz8mBnLWQfbCFjhWUWzgNcL2TQk3qy
o1R+Ddh1nCpGm6LmYKnMqYiuQlgOPkzlbL2Hcan0KHk6va7i09DAbSAgcyUpp+YY1K5Mr2RKmJ5l
sKNgNV2FL0I+pjOAdgz3y187eju9aD1A2O5ThkL7vqTOZU7JTn351qjStqMLGMDhA3Mx9/+d6dXT
75pC/mc+d9SUsDT8qF4EZvmh8h54wwBEzB8O2P6LMkVddHYBJ4ZMmzRzzKZQZ6qdb3ccbNy22STC
nh+b9NI9+augXkRfobUnluTg/WBU4pwfoNk5q4FlYYXEG7oMIFTrntMNVVJxiSR0vQ2CoR2vSXii
lOQw885NoTtp0FirJFilrz7Khm0UvEeoG9RwDdV1o9wGFoBUAHOyxhWM738KoIxfciCkr+JkPJAZ
kG4fcxsR5+qJ1eT16Vx+IiXb5b/El7zl1wHL4YnY+vOljTXQ5sXMAEF8arSFkCtEf2EZrkncPkTc
hyyzTRwnmrROp+he7PscpxVs4Gn6Z9Bri0DxXXzDjlN2OxNZmRPOzxaqvmjicJdY5b9YdAxYTQxs
75sAG8qrDJCJxkx3qUqwS5F8P7AM2ibDetf4NgGohYbKAjn0d+KYlIE01SVfpT7feHrq7juYZ6T7
2hVqhsWVvEUhF6M0F+adSk7vHCWOHrNapyU3rXVFw4UoCa7k6vdhH46kzntu48C4XyzJFX2Ihil7
HOl7ff39/D0Iw40ZnymPbywtS15qoS84MCWGWI0lKpshkKXaBYJdUKm6/xWMIIaR409Ce/MpRqkK
dWXP3z1E7+Fn+dp6GOUtyHoLsjO8rVskG2fBSn5WL5Q4b4E+MCXOHgbmpkJ+ln/vrQ2U9E/RsMKo
jkyHkxgvPreJgYMvwtT774K81pzogWMe+cEDMHLl+cehfTpwR8o+kfY8fmtFOlGPcCrueV1y6g6m
rcgeXuz/XQsw/IFhrHdFekPYu7EzwM8fJ94tuWAnFf3aKd6f4wuWhkwVkYc8eGDuYL8b4vDfI+gp
aGcJ/gqlmDbvTpIQaNxgNw2AJLcMlECJ8CdNAc98lXhQ2TmIwGmDN+4wpZ+Imm6hPR62EphdYVJC
6hI+C7X9ZtgGuNY28ZvhVaGSATasv7k+fpE7fYGGSRaL3kp1mES9aE0XoZDXyVAhIffftZWzrn+i
OR/tsEXpt1mG/mviRLkGaTbitQLj5Fgq1IQbnoybUDCX22krb1oxID2U22UFmCj536vayxEyPskn
O0c+DSLjNTrBfgQ39j09EDWKZgVhW79jBTiWZQ6MJf4pY6DzcZxlEIs3rLwmh4vYycV7scXYl0Ga
sSy4XpVH0XrB79GO3q4Vf3WP6C9YDwlh3Y4G58JNZzryuNWNInc261OjMQ/bmbUFCXi7X/fzY/YD
vbip1RR7KXPhyKEvIMifDDJF+8oTzW9CIxTUYVdSmjCkeN5PptiJg6Dg93v0leSvjXf3c7CTmy8L
rAWDfUYpvHF77yyTANfQuttznKfpoO5FQGItMJoxqrKLbyA6tjrdUwdjHrJezqyC4nixOkTMWZlC
kopyXAaEKbCQBHsr9iMnsLpxlKdG63pf4vrJlVebkP3FO/dyYaUjfSfW+bLGZn8Fcf1b+jf5VAeD
KJWzSzFeR2+zkJklFbZ0B1det90ebz+jC9JnF7KI8i74fxsREvqnjQpB019b+xebOOzqg2n1tqhS
MA3Cfm0Jz6GcTGkDUAMYh/Bq5+yfznvLzVaT5GKdCaR4WiOPp07uwuv+Ciyfcy7Y+oMNjkdOxAKT
rPWrN+oFMmwePc3YEQwrsJDuB1oMnaUD/iSq9o0YdWnQOaZDTePQ0e7bs1VsaBI+cqFp6GZxNber
m58miDr3+FKW2lBX2AQIJR37yLf8q0C2CEY+sFvTrYprc/bHjNgqKKDlLaDfuMwn26yQW72YIDVv
4wCBx6mdYtKIXnNL3n5K4CpqRiDuJBbVbKla+7WKTcxqjSNO8fpd2+w3fTU/rkN0jWqxoMCxup7p
XQsrZjM2W4SgmyuNNLM+npcrgBj21TfWs/eL7ghuSNGim9Q1k8qKk/tFSoj/Zov4xnfRCSkyHCvD
JvMV6Mx2MUJ6r92PnQ4DDrBgK6EWYaRLiQSEmg2Kg/ImJplcjyQIaM2W6jIX5ODinVvhb5Xy/0SE
9edqRNQL7w+zN+wtrLL39AmyyEF5kf6/9P4R7DAP7ZllwtmBqylX9tifUU4/Aix6g7xePUMsIcMo
KnvDUtW7fCfMTN3hGy6vIyqfsYqi1lLjgiZzQKDCO3fiVzu1hnjB+oKT4Q1i8CN+c95yT7DtOfcR
ye8F3Sa+pfY8814xLNtfBOHIwiur4pX+9wVaBz+d25ARmtHIUkn68qXRbNHGCpo3zAm1scTlZY72
BaJmkOrp5kxIx0VQl4gSLP9AM4Eb2ceaaXzkSfjORw7USsv4WPwz/Jd0YQpaVYvIRzKpmvUxVnUy
8pB8UOtlvHZCV0Xj8i/9S3MOGZFy7iQ6VvkzKbpUuywTayTPook9zFhONWEyinN6ewBgFl7AZWDu
8FfMRykLwGP2LHuzeOavvcebcWsG7ou54jTRKk4MJzHrisZylv34EH4LtVQkFq34WsVgRirroW9m
CxpkUw2F6rjiqGFhyCKHYZhuAARToA043QU8P52iZGvGFKY9O6qQT0XVQidF627vIxnyc6hJ/4as
l1lrT8CE8dQxLTgLENv6JpQ8BfKPhQ4K4i6eKcr5jA6xI0854ndtm7dS0yVLRx1AiyuhAuzQ/Oxp
8zox5c2pIHX01oSbCiBmLoV6dUmXY6leY12o0LZVQDia5YbysQuwmcZLKVbG7pUEYcx+s32BboYn
Rxb8vDm6e3WcbyeiYp7nOm8vMcSL1XobpapFvzYMOXBm2dGuRAzTyhpS4MG6W9wc3RbjDI9UvGiJ
WFIhSKoR8JW6oYJZFpkT/WhlWZXZVnZGZuXpoMlF/UXhkW5Pjmcc2l21vJ1YvgrxyKbyOdj3a2gE
H/GkAx0dykwk56fRMjlVTyCV/a/hHJRiE/CjlPpZdD9IXXV8GSPeQjxU4BxxQ2puOZiFhFfU0Fnn
olEsqBg9vqkWoYDeLbHLxo5vZ/GR+agArOYcIj6P4C937DdlLLjVbf7Ks8lj8v/ni7TekBRBpNWg
a1BO09dUq3isQfuHO+xMqY9p2QpHJb6XzahBb/EDmTtCL7j0hV2JB1V3ICWtu1iE8xrdhjo1QIzJ
hcldLHkjgOBKabxVT7qj3F60w+QJYeSC2lUZv58G3FJ53Vh7thPu3Qwj6K8ivN5LBErYd8NOKwOV
rjnlWEw7ExIvze4rJdrRUxq4JK0mo4StI4Kzy6sHoWm+duj4lTrqtr0YAe8IN9BlCOvyD8dNGmo7
AefqDe8A3IExEwWN4z/kuOH7C0MkWVv3PRcs9AHOln03iVMnZmR9mb27+3lBwU+mdmYPa8Bpxm5I
+0+wm4AaVSxtvzsBkMykOuh0IEdw8OEnEBKZbyRYD8oqXn5rwO2llwWYzhyTZNbDWnwRQNUeHVUH
iZ+O+47/GFOKu9URqbmQjLxxzGDfln89fNEWRSvtmQStUb5+n1mj89aX83g6pQ7ODDAjnnx3xZYU
RGFU2fTQpHJqRluzu1GaFJIF36IogtJ4CyofzjGX/ETjZpW4c+oIdlM7fUEDaFQXgLCR0h506EuE
fjdYMAv3JgMIFsuyNCo5t+NWTDx/4DTKTKXtuOBQMy1eKdeZYwv9KbxvfM0/Rpgv4W7iTqQ2JBjk
PNiQSGjRERf9zg7HNUJ8YvfP+1ivJc0v+eL6rv2NFGsxbThBWUxKYDDmzh6uCI1Lh+Usf8A60vEP
nSsF/87Z35O73qX7KevcnNrToRk2LfXEfBSGEjiMo/LYEuWB/NuZPsH65S7TmSc8PeKWxKLUdduQ
ZtVXHeRN3YG/ZKTbuBUkpGnvVfOsh3YZJeebif6eaa6okP19otqJadIRzgMIwLeH2CmvlQXFZ6I4
oQLMh8Gm4GmOL0TgGMVLCcq27yqQdvVGW576PHWncNtl5VthyBle9lJMSIQTTCLEYUPbFnqyLkby
zVYfxFcfKQWsj+44ZZ10VjSMHBm6y3Fy597cZ60DW1U5Ci6X04VsP2J1rhiQXib3FIiC5ZTUjEnT
1pano4v25LOFIBXEzLIiNahh+l61IfnHStLg9UgPpi0V0i2AysQyMhNe6qinf2Af7FexDt1RxnI1
siNlUhOdC6jTS4y9dY53KEGj6pWcyHUKkgdQivo+td+8HXTjlU1N67oIRmE6GUkaE2Nn7263obF/
GOPJnXmrFTutw9rx1p7DmpZqMYuhhlW4LpI0/JfY7ge4m8pFABPQt3FlwcWzuzZVG52VrOhP9ipP
rGCzR3cgltbXcc+AQb5wdof65wFC8k01b3ueIJakyii2VSr2ICBxCSkS4O7yWUMXIb6wU5E3n1HE
sLwaNnKICnxEyMcxB31QSnCrdSUeC796wNZGlKD5YV98N5LE+TYKifcOwi/1ap0TwjUGlfewJmJl
Ab/2JsN9hIPWpq7f1sLco3CNjERtWaJnT4C199fNPe9JeRDYeQIQsMliu8LBq3LFNJqtJwdDYAHl
denVP9Hsq2sqqOY7J9C+J1sWmwrq0zH/XFkFOhZUdJFAOEZ3E5rmWZVr3SEtYhDy6EjBq+bquyp6
86GUM2uvgxEPAjF7vf7IWVvAEN4UI5OBkFqVWfrqx7x4sAA6YLf1WbJtEo1g8zOXSAhypYDG/zZN
jdYbBhSG0+iXC6Foe9JSFW3b4XsAfJxO1zD/4CdFPBFgIdGcrDmZIxzhDk3jnFf6ufM/BNzygOZM
KUUw+YXEVKJ780rqutAWDAMXWeMSaof4h7goJ4ldSfSm7ksFE77S/0xZHUGvaRAYP/GQe3j8UGw+
s0hLFDsFJgEcwFhz4IQSgIgxAKRhtr5voPIxfGaeH2A8g81K59ZCimvpPRGpBXlPDFLK6Eq5SVPq
Da4+dPLnSKyiYYW1OPXXxbiMM1MMNM04SMO7nPs+T3DA8rIz3tGbeGb7ggMAtJWIzupsyz2fbLxV
kZg8h/ABHSIDsfnzES5Z4qt7GywpvklGIzmXPz94+6wiN2uIsLmBXNTrXBeZdDicjT8xFBATxyqK
xE0JIMdw/d8zBGFCCP9GQ3FBf0JC08eGniYgBCCIgYx19ThqO+dV+WMWoQwuzdWONXbKozBqDOrA
Ns7k5WSutkfUw3ZLNs8IupMsphGcfxXMthB9pdQuQveNXDoCcMipsNTMNAax1GDvFzgygsz1/5Lf
WgRCBFg7rIdFXJ0uLczywbcZjwzl+3d+nsce7gO8oC9/MUk4f/uYALdD6t9Lp7/Q3cUu51/Zeqpi
xqr8mRpgjtLPKGjjH/3ehMgMUZ0aD03PTrsbztxIWbg8ZF9zLeNoUl6sti/LQKayzhm1r3yWRniq
Po8uQqiVzgfXhAloQLAEK0G9ihHyWGTmR+1j5XFqxz3UROWTOTkfiOV/sk4UQ5Tt3J8UeZNksujd
75MT5wxkJlLLmCgggn2ihEqMT1hVOwwKIM1IF0WLlUCN1dvkLRB87XdwrCdABW/gBlVZZjI0TBhV
CF1FJfoyWFL6WV7KrtZbQomrNiNlmST6jasKbrPT/nKMb1MdtrLDPnNVPtbqmBRV9eI5NkfxbQtd
38MJztf+RpPEdubtjfcN5EcXKoV2FYoFsrqx8PGBKcwsARcG2smpgD1Dd/9R+h2zAmpo4w1zsQvh
RULtG0RHDKRZfRh0NzXQ9pJ+wyPlCknirrIJ30IMhRI75nxyXN5ApNUzx1g+w2/Nd7Bg6dxXqK3w
kg9O9cQ3SCbM5ch8doSwADcnsEAW5Fo0WG/d2iUOfZSd0m1IlGqB+ziiia+dcmMq9u/U0fmKOVvE
Q8q3i/CFD5gfG3C2XWnTE0kV6xgxC9G00w4J7bggbdOh+K5W41QOFhzLsukUdjCJKYhGvpqMn8jv
lLzAHZBePii9jJ8DhpmNuYUqjFLqWRsZJO11SlKcHxfw85BY60z9BwEJhD2Z9BSfFS3creb49fmY
OPeuTLtuWyXrppQBjvpyrDYRnc+aqQBzzWHn5CfFC+BrKYFpdl3knqTPyIiZ0GtbC9BPT0FDqQLo
0ICqYTHvP3PZ/XErJVt9LbdTCWYTNqAXxpmA+2ltXaw0ZK4uja+rQrInu4y83JD0OJe21Wzg3+VE
hoteega+RxiSUKvPeJAeFV0QZzHUVMTiM1v/yY1gfkIXk1vYaE9PsYKjh6HM0fCm/Iv6KRtyTfBD
B8P1ollwjnwegNHTpC21vw9gTGLNnabvla8wFeNwbZi1Z4Vqbkr8bWP8tc5KbvQcfe8uiVCnOkQr
dOmoVZQarh75o/E29X4uXrC2pawwUzDUMVvnNQnp8zbCvLpNVa8Igb3ZPVYEtS4amQvgOLrNGtoK
Gq7X8uMqGPPN/CyditPirgTYT7o96sFP8bdkiwpupXzd/q0IMJaqbsEeuB0i3MOfxcA2WiP1lVVV
5p0Cc90std+CrdS7gEHvlN9oGqN7KFVAuyiUmy25B6hBDnnIKiiq/ja9H1PwabBfKBgY5jndAPjD
vEEz6suUs4JBBTe4lzrkKsG+Ta1rankBMyHClRZGOSxC98p5L+TfbPMMQdmm9IkxnE7FSUPW1P2e
r5tIfqJt0kiuX1jOW83DSVy524l2GxHPscyt/sN6hfeyrXQuqaeneNT6UcYYBwF6iUo7CMJXT3MY
u74RQn1G03DQKPmQmKAPQkyM50DCHksvtxLYZU4wlT8ltOOR8t74/TfWXZdeWq7Bpm9fuoujhbZT
IHDOnjj45qy02UuHCHsFBeU3MLZ85Zz5Igh1c8mtjd7wT169eQbHnG399SfSWvOPopc5rBe6YM/c
kkTV/9eW6zKrpAjYv4GVP+afPozJ1Fshu8XmTvKMw53KS79vyvqiQ5NNInTl6XtPhmQl1ljhPG0R
Uk7WOohoMpvxmawBj6X2F96uUv4uklguYoTSMPorp8M8/UqU0j92y1rIXOHDNo3wfIfJ5vgYEuSM
LT0cgdHLP+JG3QUMEU4ia9K3krjAyVIPbFK9IIPeDkub7NylvmvaGwRw/yTWajDPgljprPeTNjhp
mUSwnSIh43nZxVkxBUUDVONrQF7uYyD4ycn5mcpeI7lgbMyOHj/j/D5RssmjcKEVCbgCTl0jiZuI
KvTTzidoKhfrpXwfSWKsrDN0oxm26Kg2tGWQ5AsOzmdXQSL+hZsRKn3/3v6b07kcHSLk/zDrq9cF
v+b2HKhlVVe+b7iAH9aa74B8hb8MvqH/8eI9QnushwNmECx7HgE/PJuad7UcHm5HvlmVtG6+p7BE
4wyaRmYK0+b1DGSEaeIZkSntlKwt0KO0dlmLzUZId89BMyjC6YQI+u6l9E2cyvHJ38obnxYHP0W7
Z/nuC2zdgqaqSD+3RL9fCAa9a7vyB/F8vZyZi/f7dFaoY4bCGND/jf2K6g8Mssl62UuZ+YVZoIjv
LiKYkjtG1YA1dySFtJKLzjt7xz/17G15BHU5p4g1dLymc/kMq+yMwxfBP3lxHdtD7L3kbhcGodYd
RrYaDsofxIW3FHhg+Lkji1IOnb6Z/CDG4RdmTTeWRHc4axdvAOYY8p+D/YNVlab9He4zgVkl3ipo
cBpZ4b23CYWMfF4KoUhEKdarPsRgfYKMBHMss4vh++lPgrYUDhBjZE5UfRh8EHLKpBxvAD/MXdQX
N7w6Xc5lMAfavJx7juDtHABOgJwAgKrn7fw3yL+GNNLK9l7wt2Os7sBJBDK+Pv2/jt2EVySEjHY3
34NO2Qg0HUbGKxe5wXJD03rrSIoST7qy326/DoT2DIQddxm8tdrHSkNaiTbPNwp0ZgQE+LzhNlcj
KN8aSiCuCDoO0RDmdDLFfq8cIOn9N/nHOoY0LdeOJCgZXsPOq4EbAIVig0siuIvkdLuUtFab9t9R
Od8zBpkF22vcuMW1YcnRZ7II2WC31N7Vjv8zocrgXBxM/EfczOMEGd0VFG+6W9hGKrSETWbN6tQb
Qe/PHIqm0veF/vBzAF7UVa6AWOLtd1v0zA/hwsJs/B5Tn1UhwZJFp+csw/8OK2EIV5P02LyoEVQT
za8XLpez1/n4xoHNSuuM92lCzFJc6K/tmNLTPWKqGTcAYCVmT+uItz8S9/NWzWIFcMEPyGiJBfA0
sDwY7EKXkuuuVmhiqlKpeqHBeyxs9D+uKT4fxBm/YqhKDJKE/j0tByymdqgyJJeENEbvspMyGVVq
1mmP4t1uUSB22eJn+O71mIhSMmZ2E344Rh0bRsx4i1348LVvniFvcftL5qTLIkWCUgezPajczygJ
izVvha4mgiW+VsA7l/pet4IfdZDpCiLLbJwEiNQ7csMGQ10iuOBUu/JNjUjNp54504vZXJukc3sV
TX2r8sks4OgQeFyK3YRWEksmeqark/9ZHit89GvvSXNSUkfFFZ47Sb+xvU4Y2eNPGggksPNCaXs8
NUQ6YWcDA8VuY9S//O5pBnfFMZ+nJhNut1HZGqwTc8euaWYURlOvMO1jCw7ECT11NQJ0qG4Z89H4
S0YS7N2TTCs0b28YgshntQDRNR2Imzf0bl5tyUkH2/x/YVxPMOE10NKoMGMj/a0oaW6KwMNO6jLU
TRRx4iMg5dA8qldJkwUvGyD3V0vfMwOq8x2JyZov6aKB7y94mKhFFFpyyACcsJfJlzh9q7mu2YdK
KKr/vaq0KnwqOeNGDEHXsZHI3SXrsIGY5hgKGv5nxjqwLuoJSv9UfQsTL3kDUZeX2nfxEpUsD93C
MIGV8a5reBRsgUSgJBgu86wAYjhYgOhu0eFgA8qvLM/VNaLko6C2yHWZV9UPj0sRcQEvjuhj/ALo
TVyhvp3qxSQ8HaPde9hNXgRkMA1W5U7wMOHzqGCeB50TY+4TzqO+QNhd0fncCP6ztcTUNlm1kRsO
AQqU2L93F71Q042dFpdvINb6IVNCP+BUUDqZK0gzCwswY0uLFYM6SAGmrkGxkKkU3/K/xrWjpRnW
SsgOaxFk3ngRl9IWihf+19HMgreK0JLV255CPPDZ7mrHk4/3qnD75Y+pRYefNalB4RRIJzaTEIAs
E49/yEfjs5Q39nnt/GXZzPiwpXvcmNA1pyOsMiF0cHOHGWoU2j018cEJRX4XB1R7k4MIWvYkRNXd
CIpKBTCXx/NPr+kuCGw/NbbU4Rn6Lo49qaHCXgaMbQ7Zl5nnn2L9FsKfZHsYVEAU6IPlSkftJl2e
vZmalnmXY7VlTwIg1fRu8nc6cc3Uy51C1T0WlwBxsc2USL0taFh7aRkpYblX3E3c4gDrlRXyKA6F
LSXn1Eyk+VYUmDw+xiP/9SudMTv1HWjLmInua7qdcRsuVMpKr+SFeXk/rQi57TXf/cLoegw4PHVQ
LWavuTsDiKqYpzz/GVLnVu/mPdCa2AatEVfAJDC5AavSgrDyDd7/SbVtQXE8zO01xngA9Yyx6lEP
ky+ajCPiyVR1izuYQjhdht3a6Jut6yOsa2LiU5VGciXj4zDXC1FPCoTiULNdvZbqg4dW9M6xkLYR
S05m7UuGDJTQ/bHOZaJQgxbaTzWhgDOk9hrBNy46u/y6pdK9eVO9zItfu48BAt2Zo8UlHbtr869H
YskXSJHbE1/4aYoV/ArSTrOFZY5ZW0R4JdoyXICS2s17da5DQVrzemgzfluCwLSETcNFm5RprLax
RV0OjSHgxqVixeHmC2LhkazO0y4TSlLWd7iOAfrabKMyb+dG/WHX618LrPruOoAg48bX7/HS11OX
3pHaE557lgBV1H5JlzMp/M+COGEeHvw6yX48Wo+H+CWKRu/puFU6EG0anlosQ0ZVomaa8G6lWh6C
8A//tzsSDAMyrs4acuunxfPtwHVsZ6OeDMBcGI6USLRtbHuCO8HUyV5k4MgXdk/ThaPZ6PjTtVe/
LWLliS54VeSB7ksF6kNu3L20FoRMLCZlY77rHUmD2gnF35fxKFwVI+OvnjlpXmR31J5ZoZ6SzIT7
VVoTmPZd6hYwvdXcuvQZrc+QLXOom9SpBWfxe7lWy1hF2jj5uHL/6FUMalKGIMXWhbKaRrT6pXs1
BRvfAuHo2Udw2ZOiBB/fhL1XdVXC0nR5/y9YAJ8qh3jNCr/QiLA9uMoXTCtzGkl8NVfQd3Y1lu5g
aPGU+icMUIzLnMpeRF65MmLUrHQRSJC9acJRvpysWNoYFpg3rQlMOZdEzNZBA7JMG8EZIyWt2xUZ
lqrS8jCAzbOryFDb4iKuztUdw+icGSOfP5R9d0b+Zk+CUS1hKGbYZAEorGM1KdDRVDO+BXip4A7D
hKVRgzgAqUIiTx7nSubcwXq/ItfxpjsLhdVQZ6vpOF01ftz6EKmbouzNMuB8DFpppAgp6Qqdn5vw
HClI+dGVKgzdGHopThPnCrBUJXhPyhtWCdBdR5XtXGTT97vTT9EnOHR3dWB7w4fTANGgWoxJEhcU
nYp1e5YfDWJX5nFbkmIHwh1+UiXR3kmZ1v1t5znUUEUt0QpcX9zuCgV/kmS5K91aaMRv7doWlXEU
nYaaHQjDmwAmqMJJUzQ613PObY0tSqYxfuVHS6QC/Ygurk2uEJfRBwy2KjaFfddG+V+BWnlIvbDS
+AEvQwrv9XojahKzHFR3lf4TiodP3d3/kB4GprJXIJxY60Ta0PDEPBf9VHji8pM1ezp35b6kBpQx
AeA03lEDsqJxvBTjDmm1ntWw5ZM2fivdDxM1i5WLe8j2tOK/vsF5PGxOf0H2wbOrki+LAOXuf005
CY6xhqpWmWWNRwld1GT1Km2Tdy5tT54F0pxpwQJQ/6R/FpeYNSso3MKDBO2XStO0OlHPRhllEfv6
3o4NowixoPRMO9vwo0PVKjrZwD//UPO89zzL2QBYqMtaFk1YdYHe2XSqsMpmLzmced90QYCo2e76
TvDjOhBAzhqqIpeSY3lHKYWgm76h3FXIzzRKGQgwq/APdyS5/dIqM7GVAlUgF7a84VTnPE5pr1A4
pCbrEsfF45ktLi/QdWa4Ry8L0PpBuhp3tEVBYyG9d+cCfaHw0WtGREkQiuUOILcYp6uzzilU2Wkk
yAEAxfSzPrsottps+5wb9v516gVZEyQ+107oXfU+aZztowW623vm9WenUQG9332WwSYPv/TPp3W8
S6g9saGH8UNm1mnfsxDBzaxscvEkFDAXYfaCLXnQQYjoFeD15/EafwDX19uban1Bn5C5p/I0bS+p
RVk8lEc3idAjbOC4ynhB81yb1R+PxhJW3faHbngRFPSqVTpBrQVL76tOlIW3ehbw+28hczINF2Gp
Cyybf71b27MI1SGpdHsSd6pRz40SI7rpVpfHcv5YACofFMWOcDTx08R3tpPdhh3YjqRlE1PR9HNG
TChmTt5UxG/I3ZRFkMuJjELUXxf1B7Y5JItGjYvZblVwgeKZuizI6lWS5rqLMusIXpDnZOfDP/Au
FwqMFl2ng0W7nmWH2wao7OKU/jFFKqO9ELMEaTDnRwIZ96J4kKLUmQGABEikVT0ajgtT8hrEIytg
IgkxWyUKMsuNEetV4aL7UsY9QqWQa9v7cFEWafg+F0OLMwfd4OL3Kdp+sv05kdRos2vo+W3N7T5J
bz8l8OTIOgGvGwxM2iNCckMuswy6rbm/qoQxvbORHkpIoRjTtP6TFdTZTSeIRB1+hN52kUeVb5eg
qf/O3Wk1l4OzHGVm+mYDBtSWau4iMwDrV4RioyqMVbwuypKsVgjkA2BnnLMfeeFZvZ/+7NxrqnW4
UsNUJ5tKThWdKKOF4MfVvdqFGXoKRLbU8H8cVm1XYh+CgNycasQn3b4x7xe6WoldH9do+Dv/4N1x
qJCrfvH1WfrB4EY1Z2L04bjNtf8DLHxrBfq0tj0cJuWlhTFKcLzEEvjvju0tA4zZDrunFybRT31N
h6yQvJyo0CqWXjudSaG1Jq9nmDmutUkNJ5B5FKBAib4wz05r43mqm1yB0MrQMOszTRQMe0PyPyMP
qwqWWgjhve8XZLPRnBtsucmmawm5JDh6cdxBgEK91UOXF8iYDGYbCXZ5oOaWyhL5+N3PAdQUPYm4
JNr+0Awtc07aK1HfPS6e0k80x9FV4o99IiMtmNBtpPGKg6vly/qVJG2vCefylMvqaerxw2muUenf
ouSM+Q98JkGDYzac87gMoF4/h/eI2yF9LZ9DJxNwD8R27VQY/wAtgqGoXDFxbM6wEwSuoRVytjXX
a9S0IQpZytMl9pFriwY7RJOLcWAQDMnrmoesdGavTBsW/mu3LHSvwnKhBaBcjRg4FhWjHJART2/J
Ntq7NQZcPz23+dYJLh6thF7lRZedg6fp6hSyl+2lliH8EDLa09AYjkNu8HNmd0lzpaVPGU7oXTlC
7slKHwxuLxfi8gmprUOQi8VzSqR5nVvnALdWSLoydM4ttZtBPd1rAri/4rf2i8nzBYoj7zT0ONYH
XpKDuY/oTghymTivqWEwI1ZCHZNF248YvRWYIAQNT3P4tKG+Kr7hsYCxWd+diZT8n8xE8cLO7pmj
yQ7Nj5u3FoakyJ6iocvzXlg4+puRwJTspjD1zG0RJDICFEYW9kO9L2J6KMbZokfQ6mc1hzxCiuwd
5FZT5pxh0ri2X1H+uashFnBV0fAsP0r7cvwvn5O7o24RNDMNDCAX2Cr9m9DPcIeWZmTvQ0AyJ502
EX7sQK7VYlAOJ2j+TxfCGto+1eDQrkCkkAAIoJGmb4oQ1ItHx9B04EQBiuqhPB7d4T+xqK01LYxi
WPocpC3LSbJ/62ZTgEW11mKsqc88PPHW4JkWn92NXM7WiggvY2lt2DjFajQMXTZyf7oea9Fnu7Bc
UXlpw4MLKtGpad2+DhLe7WaHWqUeb913zfUqeyMVeGw19Nmz9fEVF6+UuzT6V2pth0clvFEr40aU
RtqPJG6Z8fC+4Xm0049ZpYNQ+RDz0hyKmhfcJprheBQe0XUqz8z4DIDBlehl/m30xuubmZtcxHtU
glLl0u1TFtu/u5olGmE9gHRlVYUCyXWKLbDKaJ10019oJUiaxv7wvO1yGmiyQgJB+1LohPtv5+nJ
L2SfuvexTgk9S6WTjMnRGN1Fjpj+pXksdU4yo+g1/3bQRmkVjEz6uBYN/Z6y3ffzMAg59M3J3qnB
V3zLlpSRPNzQcY1VmBj9JeitSnb4uJ0h+QoK0GjSfjM2m2Mel3rwDOpls4fJL+jylRWPrJ3SmKxr
u0D5tnIkDXejqfd0KPCCZKU8juoA0QMiATMdZdVb3RLFEtTZk4ccKV1kS4Bfx5NRpy5J86Bs2TsU
deXJi+n3KuxqEU5JOexRKqThhl4pAYRj2/C8pfQ2QEXIcs4zNtj4Vwa8fZn799yJNPbubSMdWF7W
cXRFXcxn920zYmbJObVNqyIU0qWRsPkNiKOqNfg1LiSCwwFAZfh1kUGKzJs74HhBJGibm2L2fENl
cYM6gF8cHvstDjHcbQERXB0S0lIr48KF0zGHRUh6/NNXdd98YSSyowVSBl3og1buHAbn07WMMRrG
4WKDEwgVsOR/DmskkRPfar/tcRoM5Neez0DRASZjQ0vUJzDG8+E7LRcXljunUgWychqUQhGpWp4r
uctBi2X2zZWIDfkhz1QT5+pvIso+fekb59GnMakUB28oOtb76Z3Lma5DVnHL+wTuzWXK65zu5d4U
KbPjQX5YSPjE1b5O0wygq9JozZQ2dWQArdL5hxdV++wHtXN3QbFTiFXXVQZvkFcjS7Yfh4WzWzpz
gp/En+9yk4uufbAW1nZVUpeT8ZaW31VVyCUDI12lmamoVhtqyrWG4M/0AEysmyxObw+T8MjN8iTH
O1FLJv2i86yl7Kkdaq8W1icWMHfOjgEX4I0CORlqu6h5JKrX8hB3d08KnIP6UjeuuTVbbKnhnJ9X
MJ+WGsFEJR2G7lr8/tD48TiFQD+fX5TDP5NmmKprBCOnHMwZx95YsS8XIQh+Cb+6zNIsJ1h8ujPV
q9M7DxW86vrXqi64GddoGw1IRdVoTVSocOuYOAIq13/HxjlFbH00t09dtlNzjEnKhaHlOmvSmMxF
dPTdAy/PDaddu0DSFZ6Vzfx6ggnCmz50waJZzRCcnvjUMecwy9GbXU6AmKYo4pcMt30uYoWOlNLB
YPzEEu8+FQGOVWMIMPHouPySPRRNjiXCltrg+TmamR7bR7pi3TN1skjUWMyA7d1I5V/MwqZMBaGv
P4Wkw779ZWPNSZNhVmftRw9nTjgOhYN7l2ntds6eHjkMHPxdx0nwCgq6gRC5uAxDuJC1MVVUmG2N
RuEmmNh42/CgJFjpcRiXGSYHCDUws7oZR/Rh14nJ0jH1lpztWZn+d7yO1hkACFkauKZiiIEVuR7A
doQLDy1clCM8fN0RywBjUoAcFw9ukUNOU02ZCMgKpkb0rG0k5drOiZaEe+NiWLdmwqKTt8fxXFra
Z4mRqTrOU5zHGsdeNPi7sm9kBkvoQkHOrD23MNiz8w3IRh3qY8Z4R2AEx4D8zKaS96Z2JDZYRDVW
9KnbkhxgVBGj24q8OgUHUl5i3+XQqTktE5GrXPBUxsPRzo4nzmXCAnu6tS/quTJGawOXjnyb0jqS
VhFl2YomxSXXxtnUtIbF3DwDdSsmvSX6KTr9+1POaNJ67bmiTCY85DJ9wFaboLKGH9grEGEP9Woy
iuG1QNjKhYCazls2ulf84+OAp/ZofP6bd2syzK2YJhWyn0yc09qcz79FY9zNLxqwEPOpkaY3hrur
2kJs6ebytBGpoaL4Eq5AdrFeByqmsncNlxyp7IAnZthKDUX54Hq54gC1dFAGT6KWiIbo9V+ZSGgK
Rp19WuDGB2VwWe1g6dRipLI3DSKR7pZNscw5RFHipuFKwQT3mLTNVfH0VyIMlr/ybNhBPP27ylTR
x0M7PEUg25C+T6umDeZ8ceNXrRm7z9j5SNqHT04VfKGqbcFw/ahtJwN/tSeaa4U/sBTN9dZHoYZI
xrszhFArFX5pcwM9LCYNzs/uxjJzb+p5y0lUQyHxwbvXjouaPZpHcG4wxtJNgIbZa044H3EFm3Lz
Z1R6gu4yDoN8lfdVCncZ4EdxCOwbqLEf3SGXZvDIM0heVFHp59erPfqTh5iYwoeOcsYh+Mbt9M60
qusnkL869MyOjWV0p6gme6lJ/Za4MBo/LSVGiSCyyI1PFTEzaq9wXc7Ktz7vU8iTLbJrGyoH0QfN
PANHoREgY6fJNmKRvqTElbl4683OKDr4PnAxFh9nxFfu/RnfQPPUdxkBDGpSGhi0r5PNvuevlu59
6f//+5AlCNiUYX7qiHkx5AvAzXGuf3lZwheXe4DCHZRTbQj6b1op85rwDXgdveqnrVIsG/EoQ+vp
pXSy7d6y6RNx5LXFqr44fizo6iA4/DWdzW8IRrxVIgUqDh8gkQnZNOYYP1SeY36ZHbe2yDiom6E/
VBOXuGcM3A7qOdGbW1Qh+5rd/ioveuK8JQ6eDQCvgtsO9amcYDBbpBcx8Q58WLDPW35t6wO0bpB4
xAk3bVb7KRKXTo05XXfbT0YrXmUdeS8E6kz3aVmv+Bc+6zm7BTFjJhlnqMg28sA/WnEDltkvMjyG
fPhMKfizuzNX/jUQlwuvck/nFgToYT1j7oDPr9kxIQB9xXIp4xrD3K81H1oZ7DAyhfjVIpktsDdP
BDMmsNFm52zELLXuAuCeWxhbAZNLO/lT25fRJnacUOd1bmF9AUKwsplFwOXeeNQh6pSmXImg+zzi
eXr8omTyvNrmpAeMYnVw+lqruU8vLzr5kDSiCc0dMUCKbu4hGqKXn1cX0puwZjOsxCELwsv8lZPc
wj6DXc0ORH/iqt9f/WT+YVW9llTX4P3CdG3vVxdNLMyWmgMQEdPiOTrg1mZK6Nm97cijqvKocu1W
MGZstFhSqK+AFgSqgn2MHj3WD1ClLoG7TtyJACnsfOTP0rIBwZoFrbgWhvAb/xPZmjUDXKN2rutU
Oouf1ua+KS6S1JjF5dRfgkuIkl9WpxpMovaxZmwMAclW1kWDdzNMSMTvFBXLj5uHnAEYk8HiOjRW
NsutTQz7cGOEOVqxtU87aDV0aNyJKomyNFbGoJ5rYyh2VkZVwyhx8DhPDzuJ3O7yt8D7d9RRlj9d
AyVagzO2oKDD1DfsCaURqStVBS17RIjDWYgw0WUp1Z4ndfvLBzu+ci91EN6bBeGj/OP5HZIX17R0
LjvfX/eE1OjTzfOwVenxEpQCC2hzGKsrYbqdRTgt/dJ4mTP6NJlCtC3GOpqFj4AWeu1Mcb+0+M8d
9dhviHp60nQ/mVvHqx2ynBcO7FnLXiGgJSwnl1SxUj9BJeEEsromk/ItllcVED0U/ND2fKHATpTm
hX02Jr1HhDEHXGxJI9P/lQWg9zNzLMy9350vTd5OcX6WMie3HZM0GeFGlj8iiHaURaa3jEH0ZmOe
kt/rri4qX6ZWHkLsV9uua+LGkSYn1nZ/yhYCuxcRgf68OI0eu0cRzTKphygjvL5yLe/TMi+Mf1C7
SnnpIZx1UIohMhMJw6j5WNAjtjYE6F+GMLAo2J8Ee+tyyd1NvVQKXI0IhTCtSGQ5Fia50MS4D3Lb
Gjbatr9mzH7XP0BXtKMrjqJdOIoTQYhDQXiRBdGDaQZUiszop2ZsSADaW3Yux3BWaNUZJrYNCjlt
3hizTdH2U4d1m2ChR3FjsJ9jkTeOTIikWqQ1kP3fQfzxUx4ToYY97KQ2wj1NyuYhdvTKW6VDBYgi
LikpP21CXfi7BGEb0riaakXUKut5SmzAFQer+O9ZXbjZEA6e2KYEBCTmWOEIXJ1vATanaDysKeTl
NB+RofyOlDo8wcs4WfLe4NyThOyLDkD1JiBrZeEmTqMrzo9AWv+7JAibQUXNYB/7DqrjRVsZe5xa
uOgAS2lQsXtSgdzpHlcd4o6Gvbf+L6T/JcU8doyJMHAC8Lj8GmFCW6i/eUPYCtZJiVis+UaIzgqH
EjOvgqj1NGKaZDB/RfqLYryj9UwkbtWYH1G1uclRvzV1y+fFbOFGvIQW54qO5BLanjUqY+Umlfnw
a6/XS2rTumcZDWRSmO3SfsXkAZ9DJubHMiQ3EV24nJMuIgUpu2dqSoHd3aKL2bl03IJoi9egfHiw
LN0dBfzLMFvo8vjouKCKZbwQbvvbFovPdJPv0NMnXMHBXC4InUYZdCsHHGMLnQkrDeGos1S9Y5Ax
WIDFfaCZwEJNsbC7efkjbpj0lA1zHSkqBe/UpkqagAw/+Fc8abJkKq5YQ/qL0i97/w8kQ1J/qgaA
oHKcjaf9zmwNaVViiH3Aefsr/tpC7BAGoE/hVBSblO5gcnfLLin5dCmp/9c/nLch3iCNESJtHmcS
PqHRxBzGQLzDrnp7YICcyodugflkoRlBvhRr9TaySHTYlXuhq7CH7ZKUogjDr7NIhafBRUZRbLhL
q8j+6XLQk5ZGE85rwusoUUPE/iPq6VT/ynFgwpfYqruoC4n0vLzaFyhiJvwKMznzqLUfjIj0RYkJ
4OGoNh2O7/H7mndXTAqLKvLLo9dG6MB5Wptf3sLbr2ZhCgW9lTM0oWi3BdfRhLpCDtQClq8EWyB2
uuwIAG1pPljn9CA97tmF7aPrywetuD52yv06r4PPxozWVf8CBkDn46Ng62B/Py9U5DUsRiHocMzd
LdkkkxViV1H45nKa86fvzm8D6vZtVtsiGHFKKl3bwVT5VFnByqqEOQwxrXPF8Gb9CxpCuXkYhvXx
GI2yKhkVsTVcMMX5z2LUtBltB2OnBPhunr6Znoh2U3XY4iNdUWDcZVVwO0MIBz0jTfsXLm3zwuoE
yLfWWgPDUcGFTY1Lw/9VB3h0fro2qDPwmiaPR64n51x9gd/dAtFDDqz83wN/yipyX1vGrOaayB9O
ZtBTDalSzooEBYw1qj1BfJuTvqr86+9wQMH+VhqBYhEVF2pCMtkntjLIHT2d8jhlbopln7GQwCjZ
QvA3mIRRkciZqsrFyVc7jZv50aKsUfAkbnvX+QIhgrni3YFZConZLHo230fM/kM5wSYGovNwU32A
j0Kzbkbc8Ey80CWb0JybRenjSLJUjeo3WHa6NiAMh4tYtdINkatsPbNejs+0K7Q7wUl5/j8OKSoI
q7FyG2ZuqfnUra+m7QeXDG2Y8GX9WyeOFRYaEQbHptnfchWkjakvLrKpG1NRhtqXV+HA6wVMh+HR
rjz51Zd+Ngjn3D01IDghhD3oZS1A7djhqqKW9n88DLbBUhmNTrNwzrJnI8HVL62b5tXH+/pos2xb
WXKy1GIw/ybbad7guArG4zPxClyQk5jIJde6myGepBLFrkZDfJpIEv71x2g8dyejYapFUxxl0ekT
V58fZiM82UcOIjtFii9wmFGuEo1EONUfiYZecru2aQxWpOXZmljYP80fXWtXUBKxfZ+RgcMKtimF
ZrvUGbpEYMl/VRmpfdrfi/POMS3n+YG73b1wrRk8AAh6Cqh4s6Mgpzu8B8jY3pyFcsFf3M9ClS84
jt8zNtReRCGXV48Swa2RY1tE8vXQzoaDaGHCZuxdLbU51I4ybXEcO4YblxeUj4Ttza8DkRpFcWkd
6rl+R+yjw2mU4uD33FMo8BlOypzewjLZuq1CAu+EPb3j28S78555fRGwTn1IOJkres44ib8TudtU
jt8PTJKFYSM0QxLSs6CyID5dSXM6qTkhRPBL7Z3+nZwW8m09yXiz2YRvtaLhYlKv6uuZnu638pK1
x9ujqffs9tbF7PI1dyhgaV6DkKqLhtFLzwVf8nF+bK/RhO/MlVMBPuIgDAZkX2QrcB0rasnKdtck
tUsyeW5lj+mxJgZ+L94Ivxobe/K0lcN/Vi/ubxlEYgK+MCye9EW3Wl+BzdQ3i2PV8stHCnZ7MCsU
MpDalaoUn9Qn1WzI5EjVWA7rQ/Zbxvrt2bCNWeZ1/sUwYxWjhbkCB3JQ4LUGfHFhMgIk4QSYAkQo
bpzfOeK0E4X7H5pqqr4ZJCwEuJveKGtCq9U4lfU/ioivQx52h1JqHCRrwZFySDq3NyR4myWo2UH3
FX/3xldEOhWSV5KKTsDQjVvjmg75Un822BUP2yu3l80iKJeXFvYd0Na/qyonVGoP94Onp1kouWtE
SzoL44i+82skSoFzRqcUvJEZlch+d69kdriUeEcoiCR7LkPhb7hi0r3qFHiWtYw4IbZiyQd5GAC5
8Ns907Wx/tMyWUrTxA5yPqjqCETpcDLRIk6FufJ0dr2g3fuGCA302GpPjZJ26c4Eirv5A5RkziLZ
LhG83S+fsKtm6qNacxUGGQHdewIc2skfsRMmOzHhmxhlFMXN9UPfhKARbai//oNBRLV8HEwng7/i
3KApAsg+lax3rvDWNJB41tqEfytMgAQ+3OYYDw08cjDsLrPUSZmJGoLiBj63axZ1orBs0ROuttHe
rcgd5Kcm6CER0fgzMujiKBO8d6jU5prKWb/S5w+NK0DZdzAljO3rB7Xx7yFp1eislehwxqtv+mz/
stjv05skbzHdkYr/XJNcm7IuEud0aYarvVvZYFKDxlVe/ZyNGg4jzk0nhKn6RqVekt2f/r1MXLBy
LiPigaYD6EizrkgVZMR5x6s/h85MsMDbfKh1/1ssHNpnekL8ZfVGWkS5ApoqkhlkmKxt8TP4df1e
1j827LF5ewDaf4RRt6PXtCwpIiKdJfOj/L0YGy0hTDuCtjnO/lTKgLjb/NrKCNVOAZgqBlVV7MH4
v6f1plQcZPFdA9I1WEgFxDYKQKzki+ccoANr+G8OwOhJaKAiaWvKC/Ji+avAxQd7GPK1PcGzhKhY
hdQutdYQtFE8kqSaRELTLPvoG67VwCkyYJVJ5pK9QRA+krAgSyYf6D8FBg2xiSk4eeTbxILg+TKk
cXin3WVxzuJfSiMtWI+u0ZIV9iqVZhafKiwY680sGC08Qyme6b8fWIgGczGlAAUyjO6YL3/PPc9y
uepGTSeWUvXHCPYZHQbc33qAHAyMuSO0q0KZVLp9EJuRrjw6bk+FSn0cJPoztrJE/a8s6hnJDXYe
9jkpPRDtkouU6y7Nt2RCl1zCGyuZU3wXop+j39h+WkmJsLn7txxHEhfg53LyJ/cmgv6ehJWJaX8P
nXvVKt2NQTUivzZTYnGaK/L52zqFPxrJ09lnvE4tOsn6Q/AfCH4sTAJ7+URgdFyp85ty34eSdBnv
s2hK7Vyji6DPiiVcBgizf6g6nbC4Cwlo/WRzn87ozuUx9Wmjm/VUX/F75z/n/jq2WioRsNGIJikw
09pCsydrzwHltBxMHssNfKOK8r5GLlJC7jqg7Ajuy7g9F6aS/+ACgGbeciMOZhC4v5AX7pQwLNfG
2kHzn4UoxgZwXaaHV38hKIfmL3oUlK/g6hSkST+oFDW5kDHKr2atY2igz/38+adOWyf0kZZWO1wO
lHZW3ggFwHLleCEsYMNezJhx9MDMqMWPswNYO7OCqyKQCW8C1d4Xswwls3D8UL81/2uQbyCVYtpR
E2JnV0YtnKR2TOnPfrMD3Q1D6ZTzeZ7VrKO9prTdlG614y/MSvm0owfC3juelDVdkIaJE13l9ZQR
u/+gaVqDn4tBZPRNZrjI6MKS7oJ6WEMlhC670myDIVhU6FmrEVfygXQ5us983FJSvPFubqK/xzQg
JKDLvg0wrHAb9qR8Cmp8exvxZJKKiDvScMtaAr3CUbyyHi4HIz0TBsRSY1aWuTaElPZx/Y+KEuYz
ZUZa7qgeiEukeH5KMhCzehCdAP9roubft5t2S9at6b1+TbN+pZ/VVhYduOf3mJSLb16UMmGIkXKp
TvIDKRbFwje3kuXZSUZNcxJAnGPKQVNetmx4fDQLYHJA0GE9oX4LquTdCxILE3tzqmrTDYyXDDfu
hCMH+G5Zkn8nRMFPQeX50RwKzFdr5J31e8hFBWLaNSo9mGysNCwRpIpixxI1uSjGZjagO7YHUpyr
YNT59hB+imGBbR8LQlB++iTCqcaq6bZnwoW9+jKxmzc6V/6Ng0CbIpAEkVOw4mDfJvAWaDoTPoCO
/anb9LVoPfB0TIWb8+djOAO/TSoUEM76+hgoeoCZGyAnqDNs3S+96SdTTtaW6Xhyf23g4LeTwKiy
EXXjYcXrkTeFBZ9/9sEeeYOPeLbwrOrurD+nJrBS1bfOjztcpSkKy4hEbvnjUnm5tlDBnGfQjQSu
t02tGQ0dY+TG/u9yAqAuTGBGyBZ1tLzeO0lgT25obcVkxyeI+a1BNyfLNkRvHztRxFAjYTq6zDQb
CZy34W3R+5k3+BXm9Cp37Cqdgxb+1mQWstzmbB1+EeiYdH6/EGEOg5JB7qpZOAV/2eW76R/WQBmQ
80NmCPhA0uvb3fbeT5qLXDPd+/E/t1xgQ/rKNhLMeMFjHah/DDSvsCU258QbVb8QHcG/E+35xFQO
2t8mInm9hz8exH7dShbQQrI5QZdm9m1tfdAQ8iBX4e5AH04Jx74sZtOQqOsEDhqejFMiT5CDR3NH
RUDGaR6u46G3dXvSxuthuYHB//G4CMeyRlsA64Yp/B605EUjOOAFQN4AWgvc9GyONpFALRjeEZO5
0L5FEFsysqN2dNIHTmYqOjuLx7KBMdG3Dcl2A+maQN/Zx/Z6AcBuK2z983zPSCromfVckUc95eoF
gPhYf8uI/YO8Pkh+3H4hUJUFRQzCnrb0RU6M4SDt/KctB0ynhGCiN7FqrHntDHnZ+ovjdEoWquFd
b0p8nDF1LxxNnJcr8NO7ijjgbhKPpcj9D/6eWfECPK6de3+Gb/9SHp/8xImyTt8K59jaUlY1c6e/
MtNs70akUQevbVb5sJk5DT6fZ6lwuRn29qVyygjU2oqtQIGFh8AeBAM1MBsGfFCyyRg/ypYOmb0j
DzGNoQfjY6gQZ9f/iY+3RnQn28Bpdp0ux9LkdBGd/gaBudNZDVCrigf7dByPq5gVIJM/TC5FsEXQ
00mFjG2hh+7/S7Xgh+iuSVYXPnXLRMlQB7/EecF16Ry1Ej15ZPZ3aOOFrhvtEfwtNcc+tAeiDiTa
GF3GdoOcExm7GecUGSBwi7zmzIKbuTrNLQf+6VnL8DwLhXfRwVusYdj7hO8mTy75nyh9RCd+AvtR
SmBijtZ6sIEqJD6y4v9yNQHMdm0ceP2xoVgMlszQc7WQx7v51k+rwLsZWIyHTLQYxrqAgehj3Vxi
mj+x2iyY5woBIWAbwYiNjP2aUkzwd3DsmTGeSS2h7Ltx7zN4wN8RFbX9nPVHVkfcKimoGIP/ZxTO
eyC5fQwNXOz36b7FQpBkew+gH8frgxv9kMT/YNdOwLpiCkVeZNotR+SoOjnZnRWhCnQlKh5Lt/Lt
ymnihORYC4wdZwvvzGoJ8TP0GmNmrV4t5RuOCs9uRykiQR4u2dGRTr5qseaQGQJz2D1ZiQPWMaVS
v8PpzFHpJJqyar4KH1XwcLVciify0E2hPvR3Wvz8vn3LGJeSA3SqAYJZLOuupZv9LIJdveCxiQgV
kb8YzdP0C4wMW0lnIi2M/l19mQvUBz+npKacn96lE5WQX6p0btst2tzngHuAUWuuqCOiLJCarWQV
S6KnpJthY/Nc5w5/HgMvGOuPouRiXVX2eeG0UeXoif+G1WFtrdXi/1Js2MguCWsa7lOH+/uuw6jj
qoZqp5uA4SpFIzPJ7S5PQDCWg/kERupyruJ9GI5EOzGb3e6qdJ5gjy82MnBG/GIkOS1aRn/qv4j6
WXpOnclyJUf6Vc4l584/ezhZOa2kANJsuT/78mYVi5k1djP1PxUVAnUZrUSeI+KvxxVUURC2REku
nygdFSEitAnmup+GsfQYKx7OqCd5jHi4Te+iLY8EuJL7deDk6+QjnhICZhcmoGgsgjeW+K+RxxYd
SHc75cK8k1tyOl33BEow4q/AiAQXUZ0pZYZ0wlH0/+b1lYQhhEXVRPs/xKdphTT0ikSRW9Tv+3t3
2d0+F49BV6C1Xst7W86DVbx+dAsnhApNL/VUFiAexdlxQ2A4/l+djoMcjQoluIkIIkuNIj7qzczq
XsryGqs6dUC0AGB89pBdOzGpmoRDrhtudTu9rEd8Teg5HVSz31ocGiFdEAWD60tGfqGHI6sCEZpo
9ei5JW5ya2erNWEhXlDdydQXJNC8QIZrFUfu4oplJOIdJTjD+SvMZiWEGKJiW3Qdxy7gzERD+HsI
VLmQFubgZq5Ag1UbS5BY4OwjtZAtnlkRJxhCXfTt5necK2a1Bj1cV/jPgIzJXCqGw4HUOEWP+wAP
0PgKDrwvp2cmty74tJsTK5xx0SPtsOVj6BiMGMvLjUiPTj+IOdVBXZjr3ELGya4w32Qbq7CSfdti
tJaazZ+bzntA/Flzz7e0LuEdg0lNTTS6C6D2dpKEVqOUf5WZg6pQdjJwC6XhIocNyN9iV8+BMU03
t1SwydOU1D5vBui+I71LvcB6DCRQ1uCnKIToybaIoUkjlF27TeO7/wJDXALzhvhEG0dVfVKyrYlU
aYyngkpb47PkgNIrOD9mwptPOSsO/RyG49DaEPmCWo0F+CEqgQb4sLC4W+pK1jyCz+YExLMmTOH3
mSrCDA2C//TaZv93dL217Gizop4jum1OAeOQj1yu0GBfbP4wY0RCeY36yHRt7noTwSBf6cGlR/Ga
BOL0ZtmHvv8n30+ExpX7t+OV0LqnNtvRg1iWXhXIeZ62fwyVGo2C0sufxT37IJx49fLUpNcavQBG
+OpgaOY/ibhd67OqcknbvP6y4/BsFWaZz/2Cb1a94pWb5M+spR2Jh7DK+VXaDn8sCdWDKBXPeip0
bwY+qvhXe/vmrOkXvYeAfgJwgtaoH9rVo6fugdJ71gtNebSFQ52EHUyrmbSSELcB/nngiZTWLVXU
RNfBgnt6dfjKpBMbXv7roBOzVF1K1i4EMpsmWHVT7WPCURpnNgCgv8CFawEvO8YQz0dsDEOFWJ+0
MRNJP03k1bTYluq9fwouFAlAaWBLohef/eXFG0LBzJJ2iRHaUsSnGsuEF0AfAL3AYdkL06EdEKai
WMMlYVlZWTzX4u+mCQcJyGRHbz98xKrpWs/+DJx+pWyDJVJ+hHnYKXcLRRb4ys41fCADuIW0Njxe
73ysdXF02JY91Zk+fZJLUEPOpT0SZBRhFSeKYg/H9BjTS/tdLjyJ3oydJmwrZ4Vp19G96jeS+lQu
fIyIUZLbgmNoDb7Vrtry7sbKgVx20RJGoga0fZUh2zAB5IwNLUJNnp3rRzFAJKVsZuZmXiCqBuNI
dxYBy4VeE5aCohm9s00c84c+YwBeP+6xGomPOT1ktdM+6XUOT//YlsUWC5ZxZddwaK6uEqJgTb8s
toiK20Kc2bmAiZOF0p96rcMwl2wem7cTREfX2xc5EXxbbynj6z0uwG6lsy3misZ9rCoAyUh10zIe
2QGiADoHJAWuVZL9KPST33o8c5KKvT6GONmnDk7K345VuipZBmkAzO5Tza5BqwOdNqYScvd1j/ud
q9XcQ8AbVvBHhdhxwIdK+ZuC3WYZ9We3q23BaOeoUf4W8rF01Ho/7RA196yh74H91eQvtr7gJ26Y
0UT6H7sbHr/4RFNSpYmC5YKnmHfnklIMFLPk+w4xB5VE45FgUJ0JOEEr2+v/ir902POxCC4et8Iy
i/cXMYaYZkGJ3rMuN1LdPcJgafRaBFyRyGQh4ls2aLV4ePMRejLCLQGFifSBhe183bKuIMLDpRq7
q8S3lgw1U7f81As6bQFIK22IvUaaR0uQnitiGMWuSAv7SJx+9rI0iapisEZQnwEo5CsnPtJYzNSF
QHW6hutPNMtRYkklBXmf63JYhS+GexjspksoMb2zBymawY5xpVEtJjpq9moYDuZIiKBpCkV6YZLL
ocIepZYX7ZuKKwjhtXQeCgNc8hw74LJN74D454aCHomyWR25YIsgEbMvfx/PuOfMggzenkfitEsV
3asg6vPzjDmkkV2kpUqY2BkHZ/zyf6rAZ8xMIZzkUinq0rBmJLpnb2tXEMh2VSuPLLneYqN9uAwi
1ExfX1h4M8ZT1TNwhhXDOr5+1gKwLfCf1eiQBzyC5WM3PKr5m6ekXQ/EaiaqKKL01ViYk4xy9kcg
ZBnG+dIIbWXUYg9mCaepsE38xti7O6FAO18XO++gs2vaTaMuMvcedo84wMLwGxezTsRoncU4HApm
gXugKiXLx5dJGH1OYMCAoilRA7iTt9TO14l/oKlBzyoHUqC3PAp0evF2qS1HU98QHkD98uHW4p9J
LqIMT9dgttRzYw8I+kuVn4Vlh6e2JGcHFhi9jFgCxdL9rEhQwW4KBY8Ppa63J4wZjcG0ZfmqmV6n
v3rCZHXph+nPyc1jfdI37AhsASmwFLz8zuT9FZkk5jqi3O6oBZts1dkQmg020DmOiImmzBtMsLjS
D3P9Eofha6pRsci488ECp5VK+e5+WHfhgek81SCuRiu2+XKyW/2yWskECrjXp1yBOKqnK6PCzBsp
UojlFTsafOtt/xtD75pLthRfeP8y2FGFoMb9QnST795zJuNg/4+lfSzn8ulsCZpR+GImLh5wKn6v
vyVWJP2z5Z1WmAiabRM6gphX+AoiAaIoK+Q+omEcH+UAKCuMeo4Ob+CBY8vQ5SVtkgTm48UA3GgH
Lrnr33963+CZ0slUyf5JgcEOql4uaO+zTHXncsvDQfzOrfylCBwcwcouQnE0f4Bec5ua/BZWCJ8s
4HnBk2pktbL+b1+W4jmjAkQQlORTmqhjzUMCsvyuIhss4TABE3zghTPWOrsL7mSXu42OCKO8ruAM
222zjV8rfEGoGhwpiaM2DxWq4L6s+zbT7VbO0K+10CXEG2mSnqPJ0TA8eucmctyc+GeLOAx+UMOG
PBQZzdIudLaGJlOHbp9y37OFp3pQF3ARsISSxgavnsrmMpf3lBoiCLmsz+oaCKtRrdx/kb5gpQBz
pKrOg5V6QzzSYz/9XiuMrTGGcwgbOJ22lfO6dwfchadPJ8LetwoFQ8T9DdXGJfefcW2nxT/QJ7T6
ijvE6tZfzH+v9hmNA5rk5tBfJR3mLujwffOa0LUVICrKKpmO26bspyy1XbsRz80xRtvpWGAyMPfP
a9lPgt+E57kBFZ4AIiY4J9ku8IUFxmcnvOKwZ5A+LJvjoCPzPnJaDbTam20CbZI4sdUXZ9hUN2sy
r1OmrJYMZdCSk8uOjy7n1+K8y66pi7q0Dt33jfnCTd3vgzySdmCB3sOClpmyOcydNsHc2P4G1kcU
LrtSIop8j7VpHFLAupwjK/lVoXfjYRq7HlBasUcWDqxffifouO0giAg+/eT7aSGZtCc74ruqS9PQ
c8SitfD8a/nlc/2sKGRoqkvwhisZgl6G5HupAwZwS/fIcXr24OeS8urh9zeuIEmW6OyW9W5xrJqX
76wuHCJFE5X7zdFUWwcb1iJhfq2qsBW52lqG0prfqFZqKEatKxH1+hNgTinDE+HxU+mAJ3Wnaj19
+9AwFDYE4ceYdJXun1XrbJYRgbp4aa+g4VOTygH6aQgYgZ6MZ+FxJzFwoNKNK+yt4tXoWCok39bN
qAOZjx8z6eJVQ6W9POmV7FXt376JoJbKf+iN9Fmrk+RlWY4FyhcxA8E+yVTYC738lUiSJkLWLgE3
Y15c4W73MtzOfKcpQkbMbIXSU5ise5ypzEVf3tZXWdEwj75VjDngeZKJJ/wQyxPX/ZIvmIIloJ2N
gUgoGgjKVvZyxJ7oyktt/f5AcxdeMJ3Frqnq4+qozVULwgoDkVZCCBPNpY1lA6gpGpPn1klu3Tia
IYOfHX4NBx5A3+cAsGkhsuo4KPGpR66lVH5+JQj8d84uh3XNC7/jgvaRcK+q9ZWdPCSKOvl/zDbG
ClHSXcPH+54sZtONgdMp+FkT60TmfS+wpCSFET+WCyI/ZhTmMFtZJ0lnyG+rVOmKvfVho8dTPFYp
wmFCpCRm9qw02Gn7j+zyuVl7w+5sE7BwhZD42wSzoVE51LdoR46db+1vwYf0A54DRIfzSc4FbkF0
G089jbKUUj6ojFfrTZ0bGZ8pNTJYIutxWBJLtchkFOE7vPWP5b8jnL2aoD6NYqtvAEivuctUA9rK
UpBsFjFiET7OYAyj4FLT7rOe8uQeql4MTwOOKmzVJsnqySJ/QvyotX3lwQOVq4uvgjHsSHpFu3kX
xFc786uzzTfYtbGr9F7YtwvBb5TUoaWEn6fhoa+QI7wt5QT/EgUTX244D71mYS3Bpm8OG3NM+Daj
kBupHyd2K0yDgJ84Z8L17DUEFDGdZylYpCX/pYaLHkvGikjal1yimGoNzxDRv2jIXDT3xxsxqckY
LRiEqiT0thrwaEjnSBe/rvmGWSa90supZk8v7kIN2llb7w9PR41zlz6PjlS/SwFkb7/MYIABjE4J
ZWGdiVCrZs44EXrqLyAnYpb6oxOLqWXuSSUWdsZ4KkUmr+jBoA/60/xDjovh+WFNQ6uX34LmbD4T
P0vhWP2jb4RSHcN3wnJvMXGPCBy8xD1r/BbZkdenLMQpvRXME2pfL/e6+xP97bIoJL9Qxjaj2yct
dOwvY3p4ZitDWsD+J0AGn5Pk7t1voDCKuDMZCLEeyI3vuYgET0XgwIH3WwA5O78QiTqcSTxZYfqq
npKPDe1X/+gf9fN0evPadnlEvU7vo9DpKcOhRjv9axYgBSR4u5R9jNGmvKfhM2mxIT3D46euDcd+
IUhi3HSayGrni4AN8Ki0OP/eaVloOruTbW7E4y70ZyiMz6WxV+Z4p16YDQuruAD63SMjKGsbXkPl
jZMtyj5MmU4CdDlQp7xFPjhEvVH+nwa6vDjf0n6Y0RSdyyWpFh14GJpOdAlVRcgP7yFKpai5ryn2
+uGndURSPwmBO4u6XOUVWS6skczY7NXe4nc1C7b8Z9ZZhgK4WM+ZAQAkMsh6h8azepboN+R7iphW
kgFswVNqdlnxFi6Sdw98Pl37S2F5TkJPuNTjfqlamRVa1idWftHpbTkiwt+YyaXNjtUJWnz1Y2c6
7PhZsZ0uEBxe9h6XY0SSU4U2M/WstaqOG3VWtsuucAnhXipLOopStdPwQehHQ9McM2ozUIM+nh8m
qS+1VjX20EPQRYvvDvRFknQb5EXNRZgXimqxUJ+HnGgux15mGmzE2KDTsdIW66C5ZcIu0coxIAAT
fHnrqhgZsrvmkmBhII2apeVybWFANsnYKdg/MSY1zEi+rdH6h1+1zQCI1lyTMM5yJeajhl1JtZok
wUbFUfkODUYeIbZMBqTEK5fwMryUDftj/I4zustE2ibaPlDuGBBJyMQkfOCQlnN3E9pHw/vI5drN
+PHV9tJyFQbboKnSEo5jHxfA/jIuLFobSkSMIym112VQ9UahbV+FWepZyQy5VHuBiuk4bVVG3DvW
0B9DtkSdfLtpCMTd15YaEMBzaclFr59O4zsQI0oRe1QRBEmqVExIThB1Y4kzypwmgc4GQN+EqRr3
QsqquXNGkXfObKstG2/VRzkr26WWivMiQlCRvwffIejYBMBMU/Hk/mR0SQGSQby4hFtqbJAJQPi4
TLJFx9CVmUepSxMecve0S76CubKp2JqyawB5T3sjWev50s8YO650+T5IAVQQnYM2i57Eyi9U8ieW
jX38BMAAsXSXncPf3X8Gh+1RaLFeIZzp38o+al27WXtN2vmRhNzk8qEP91KyEgBcPdQFSjEZzk/3
oOTsXeqILK93GqVlFu6Aq28PoXXKDM5MR8Sl0WmMFYvuW4DoVJqmKRQpC03BFnyK1WwsbxbawX1b
GDuvC5xSa8AZP65XgnSt2c3uky04/5A0W2PnGjGwqGGJq8vexUSj+9sirkUiqMoGpSIuvdSA3Zze
EJjWMVD1CXVN6YKAiwOBXGJB16KdyTgOYkbNDfEJ+XnWURSYZ4V4Rt/d0Z7V+Gv4iAtyHC8JgNAd
10/ypwhSvZpPnyGMWRZ0IXuODCmsHwX3WKCp42CFshE7hMkAjYuR2MCLSdt/7u6K73xJcpILIvyM
t3r9zh9oVpcj6kVOEX4yhsv4HBlhCJExTTQl/HB90Idfa+3cqzouGnHK+I11rNZwe/hGD3RvS/Dw
WfrU7Q1i6fkUvwlfsL8gFKYWMsiDheC1cGLdQ9B3Z9g7N8aaQCuLJUAIHtJ2cNTzhvoKLw0YinvF
Mgl2rhJjbwaOa6DleKVdLLWKRX/5hsDpY6gUvVeFctiER7+Pu6VYT7+fQuIFsTMtn2iv4iRGnWv3
WP+lEmfyIxe/ugbVzLCjvCSnxqUEYt+13i+KAMsdLc2pzzMwK6ecFjvIt4VZm0hPLlwc6uCcZGxM
KEt6dda9ZloMD5p5SiPHtIVCsUryfOPmuWuRVBeX81L+0lnPlkdW2/k8ENO8mV2shSt3LcK8qa/1
bTdFlD/oZq+ru+MMOGREzNUnIKQsngitxnDthywZWlfjSgekGZ07dKkEqCueinqMzsS8Rh3OWsmm
jhFhjboMt+rGEZ7zJ+6o5D2yRlko9mIWd8xMTsHtKxdbMDgihk4bYx/HeUDO4bFYU4DsncHO/qBM
v2GicH2AyteA8xdzjeCoOxnr5MDaNAo10MOSwNJpbqFicdSD0mw/ghZCXwbVToMHIjXshfRQoET6
hnFYdecbqNAmrApj4i8RBv06t+AjLSGCYoNfULAbuwcomuNIh07UzoJYoXCTGaaP8HQL5FiobLrd
QBZ0sRqk1zfYm7I6ioogddn8oUxmJXqRHZVvik1T1yuRNUG4Gw5UiDACHeh9DHGMzt69IaxLWTsj
cdrEv2Y9vskAp47TRz2v9uYaLjSGNWQGhYNSF5QRXmI2xUsxwzjBI+cxfM8CLoGpaliAozneyuFN
gBl8sVXzMvNEGi1dxKLX0cudiN1twwt6QEOlv1tRHOU5wxOKSB3Cl/9rbir/P6b6RaA1MqdvKSPj
jc+lz/HSD0LfJgXvM7R4K24D3cfLieSsSN7Rs0fpwNTNKP/4H9CxxAp/A4KB6R/eMhu6yNCSlDXw
l8Gnj3mO+V8hS1V5EvR9j0EbI9OqqzBETmanDJZ2vjfs2Ylm4oJbcM22wh6hCzyKCuAOVnpP2u1I
VaD235mOO8eWKjFKRBtckQu+YxIAOiKUtEKY/DtnOXNhWtSvSa5cuaS5w/o8nsg4hnegBsUShmJ5
e2DiDjh0zq+eCXZzITffuK3tnoEolc0kyRo0di/r/A3eGUkp/oa6u9/lflXAa0J3iKOZjeQ81txG
ZCbG5+g7L+EA2k7rdfEQcjEA24neTtdZwGKLQhVQ/GX/6mJcTDlc8no4mObLY/jDer6MpzYUosQk
72PzfQIf5pzyhhQbpiFg5CKUxxQ2mw5LfB3pnP9LOYAqyp3jqp+twrkIZawCnjLPN6WfcAjy0CRs
PECLfkoABxBR6op438QYor99BzEzYCqFdrohCsHYkfYOLdFmFbZC0Rp+I/4JXiZ8rBCkRDceum53
iQBSF+yU1QMavYZJEcBw5alLEZcI5klooMInYxRfgmvkvjnfSRfqqCFdQ1hDGngMYJwKPqWPDmAM
+bmQIfd2DaWT8HsS86o/e42PJ4JqbrzSHekmiG4cq5bvbyVch6umlBFABkkl+urENw116UhuR0/u
R/U33P5SaB9nQLK4f2m4dipbFqbgL08L/7ndYZZFAMiV4IcE+bl6P9bplD7j5uuOz8R/F230B/aP
ODsycq+YalNLgWVsN6bARD25Ckegr/jww1RNuho8NDn/6+jKAfFmJ6IjCx/r5i3XY+nMZ94ZzdH2
abWeFq6K/ytR7Kmp2NcUaHQL4G3gSrWq0kvUMaKWJzXWWI7tdEl3/acRd0sd8+1h1MOKKs0/1Ksd
PSq5PMGvdvCPnDeRwWpATJ4M7rPOxsKtxvGR4Aybg7/WNPrj4FDIkrtq63L2A+UI1PEwy5kNLwW5
GL0PDee2Kt2qOfFuHkfHgCbcRX53FIpv3Wf9MHy6hbwF7tg/g4U3O26bnJ10ijryk/NsalkWv23m
H5WlqCVsMz2Ug5HZFnrlmygmzmq2cwSvPw67+R61EQphj/ZS8hPoHBKmzIfGR5hlLCoXUolJYiiG
SfBeVvcr3YekA84G9gPt85SZo/9nqhrwiNGiBoT1ylDk4oViG9WBQlMNdXYSR+vQe5X34Zy/fPHF
v1bGHdSo540gzqxPaySvVYdZdiVuoveM/iSJeq8y5g7V2Y/jvgtrG06eDMM8XTO+iOrj4yvscSrA
TjoyR8qv7rIekzt5KGw6ckkuCYpHj//tISi60XoA6LYTEDD7uECRVW1T6JoXpwqg8Nht0Yewh3NA
1VZEhNWpKcdT8YsMuPE1JmF7mAS65VeUqzyLW7W4jKjoGbMiVy1v9I86Y12e0wPRNoEaQ9gADQ5f
SL/R9enHoo2LUF8KJ3bwEDrqIzmDw1gVygEpXwW76LLdEB1w240RhE/KTu0P8cL/BGLSV3bXTbty
poRWJ8TGTn84YWam04OvYP7K/VNBVLszM0DVbxj21Rh1cCHN5Mh+bmz2iJHj9FSful3yCD4zSOP6
agiITcKY2UL2JAtkEPGYuhOtHm8aPQNBzRrq4lPxxx0xUX5ssQ59co6p/CvHxe3swxQceJ/uiDMu
2mK+cFrIhRi2Vi3zWFpuYFKwPAPrDH5Yhray7uC+Zo3Ugh/iEe8ED/FBlvqh7RsW/pwRT4dH1ksP
7bwBjTKf6PU7ZuVH82XMTKeI5W4bwIID3dxLIGN1r6sRcO+GooheDTGHbR3pkrISSXeBrZyZCdtk
5Prs/onaQnu1rW5xeSO3P0KDu7GNj0JZo8Z+pgwhusXkYbQxGEFMsQScI9PHZ1uMgavkJcFwPoro
6w+LRgck8553u6IJCxv/Eo6eKA3JGaWwDjBrMBeqOzoCxA5TpS5qpGrVYYr4jE9OCytbYjOLeHVE
0MuG+CVu86pA+1wqibEC70Ja1DYAIpaRk+Z/rIDQQwD3n74Ta2lBvLxQ3LNEStGCSYWTbSxcbHvw
03aeJX3fhd28IvLdPRsiFeb3O2t7KxPEIJzn1VlZBTPbb8lqyUSe9KKt6n0lxLn/3arZhwuMmPTP
PpATswQMTzByiN51UhE8SmUOEk8CqmcjOeHTBNH3EJhIzudh1mcEWP+0uJVmmMVIeL4tlKPSvq+H
mA9srTcMRc1zDx+qGB8zEnEFprbumh9kCcYaGSaMg54hbu1LfJ4LRrNE8O1kzvU5oSXsIyoUFd0h
GTvUrp6NIVrEsbUBkQE4EnONCfscEm59Nq8ntHQTGi3H6YyeYGkCeIuuX1V+B+y6NgQ6YdqqeOiF
g7w8wngog+9faMgpfJeHM4XYfsAAmG8aMN1EmwvlEGw3H9XLoMpQFwP8x5OqGMRvHqWbobiNueck
uXnQXP4XYQMwfArV+DGGiwOOgZJ2pVg5bHcy5hZCSP0vw71JUeI/a23m7+raQYxDPJCNlcYAZKB0
8k+oqvKZv/j+Ckxu6ZcXw283S6LwiBm7USugQMH8Ygoxxu9QT1h0ZLP9/N2hTSxNRWtrUcUNRnX3
GJhEx5FWplkzW0eR0S8IhgV8NnOSkLD0+0D/pDfMg8shctVr0VUKLvwJKbqKR4I0Scp3q3EsKrg4
4TdGNaQF3mATz8tc1bLNEJziZD+D04327PxJF+JReH54JLW5Ia5bMUApjy5mmV0xmczzY7H/ykwG
5IOoIpKXIMGV+Lv3ALLz7zMilFn5hXpkO07QqpMUEvvhIuXK6wqk4fekSpipKsVAaV5GhYcK58oQ
sYII0aHIKGQMTNkf9+ufF/6mc9iavuGPSYAqypStqXIn6NVzANFxS1gohEtdn/pVdjcDIfEbBPn/
9TNjuH97NAX5KHH9z/g9AI/RBfWODEwG6v21mX9nbZ/qDsjMqxW7XD/VPQHgTg10OZ0aRK+mthJO
IhnQ+hBtWDACrJymyKtVScf62QjwqELDvLPYVVTE8G2dK/ZXAsnXkqqoXvGn/gRACJXlGF7KH+1u
LmMmyLK5IMTa9MG9rAqpst5OWiHwhOBjmMXvHg7JNlPFvSP32CpOaZN1K1LIn6P7LvZTeGu5/6hl
3vSzpvpI+zQAnANJcp/o6jWteaMASZslQ65N67ur99To+Y3eVMLIZhv8elV4U1j0MQIGsaaL9CkD
u197AcbZbwy6i0Dlvo+ucukssNVSBjDKEgh6YbTVTltWufs+DjICwsjYiyu0hnjGh4n6yX1Rb8pE
pG3FazzltSQDV6axt1nxLAxS8pOlqdswxCogFhAXz0DbzTC0HlplRg8ZUcSZFD8rJVIDoWHNDOgt
b5KFEUeA4+Zh0VWDxyW7/75XeQl2qj7TAG1k3g9bg2oLIsFGScbatfzylFWdFpDMgwxFnzBUmWN/
5uaWx+cF3PU8qjxD+FkmNBiYe5q6AAJmJCiiErhyc82Ou5Otx4F/wVp1WNEMHJEcgH8PnPD1QFEy
ZFhXdS1U2YrBpYnsAwSGnsEcs9QwykOEW3Ubm9pO4eQA58AcVDM5xe5KnxvNPO9X4aSjGhVMHLOY
zfd0VOEu9HivxXZ0PHsrupw1kugscpar6MIT6VF+7r+Ka9wQtquUgmSLe5aAScYrkvI3r83DhkuA
oziNFMfOQpOA6LPi0WcdqyuY5slp1BVAJEA6SxrmH+vBAmPSxyW0QoX6df4N0AXHy0YwMx6/1EC6
+9Sk513kG44OBButZyZtqQJGHCAqg5SMs7/a1FNGIco/doM+0iho/Qj+zWktbalxOvXzcwxW48rp
gtXRYV0fokZ+d1k8oyM5wTDmquw7Em8QPrqgQ6swSfsdw9JB+EBG/81RqNFcMixoGpwIFi/MStLK
CEWCVU+VA09Wpzt+bOKujGu2OZHKcnbtwA1JqsBWi28vVqjYW2xfbrwOiqcfQKJ1omhePsJlSpoD
4GQpblAzCM1cQFOI82R71y582R7g442OcyHKIrIS0oTqFVd7nsu7uyEksW0mUUXSXyC+zb4DxoDa
Fm5FqrQ6lBKGVM02MDxjKZwF2Px5BTBBPGTWttyR1945Ll8DveckXA53LQfE7VfqLlfc22EmpoO4
dVgQtlKviVK2pNqegDfqcdYPBGGuBDG8nzB5ODSpG/724YZj3Z7SUjSrdQMuC7YI46L0ovZzs5/X
7wcN3jmUfxVS5VjxpEvF1XkQBSB6XnE4BC2FLPyNL9wSn0/urWhjchInepGaHSHERvS1+yoqlkz8
ViX0D0yGUp9fsQkOw4FqyYyBmmJm/Ahyf2ARtl0f7wwuCMXbcAyNwCmVOurfmZkDZK0F3IWe8B/6
+zC+4x5WvhlqyGOr5t/RFFbFw/NmY68kLshAfUxU02P3guFOdoK12TSNkIhHyFpNL2YWfCWRV2sl
tkInoDv1sfyHPoUtLlXkC7sCv8eON7kxw955V841gzSBNlBOQ9j4MrVMMnU34PzVxbCPpSH3II9K
t5ET6eokMWvx6pa9I/aXI/6hvFazCaPuEMvXeDrnfvzagRx+xUutOJW486c4ZvjETI4rqryjTUMV
supi/WNVe8YzH98LjAp4JTDr53eva8qw2NW4NGkt5s5YSIw7hMqBv27UJYX/IWlgHu6zhHMyom7k
EpVZVnfACqVJ3dpdRECGpcvOI6/LEXbe/cVI2z38MIk9eslaRQvUltvW/seBKJGwxqmQn43ewXZT
+KqHxLW1O+92yvilbm2UKSBp84gcNjJLnXLyUpV6e11SXhqSHK+myrS4DdSmWlW1p4uLonPHS1Ik
sGOrAcDvPAcbrnwDnOi99r0N8ptrwHbYezIo8NLrFxGN7zi8A9p8t/qwq+20lUcRoNsGfj4mBVwd
s4CzCREpEAJCofTuasv50VO0MOJXzt30zwCPUKDbiGDceLgm+ZcQZ1KSo9NWAocSK94EZTsTkEDa
HunVE5pu/+L+Y0PVsFwPSeuRkIqSKV3+GNJRItpdWlhBbv5VYxfyIwGgvcUhM9AFHsJprTZIbLKZ
Lwb2TjvIwe9ww8qwI3TThqS8RHGDNI92Cd4E8mpG62P8qdyP9PzXTY3DtffFgtbXku2dXWM/3nJB
+6vsMuarlK7IdUqeEaOhaK3ANj+soUJ5xDAOlDIZ9Rb64/RU6kMLxmvbTWXTcw4VhPIwaWbHCK1m
Z+Q+v8dMET+2XVpVKCKfamWUoV9SSXOwyRFtJFU9XJM8Xt/VVMcU939JtsG9+JxTyNGGD3VbPT8W
vD8w8RiS5hviYA3EY3FgdiIUrat/6ELwmyx2MDpXHL+7gFHOuB/CkbKDCbtAtD3z5Lf00VbchFKl
7YoTzvFAWkrZz1Y0OE+NTVU3+Ap+vlx2W7BjAexZeadwvWUsV3pWN0Kp1OmsbHOmrx+QKObHpeqX
5YFmKNF5mV1TVUctEdtW5ftq7q0vDyrKE3YIs2kH4Qv3vTypoQ0hEpbCYNqQjM1L1SkgfbZr7fwA
sfidR+Rid2Y3r8lrhzy1083vQV+3Tnux6RZgZE3ok+b7LPsjaTuW2ksRfmnlFTkdvllxHxzOdaxy
G3IQMpfOB1vAMzPkx+8zOnJYt8jLs5iEzqBdKmD50qVav+Tby/SvZXFfDPvyX0SA3IeylcHhTrfL
f8QofAChNl79aUum4Tyrp470jAX5nBS7KcbIUw75BKH0d6R8PpjNmD1Zwv6cLp0Jaz4Kht8z45md
E5STAUpbnSVRcxeu8G62mOcWCGnUpUFgKNytMC+l0gWuzI74uDvctYGhyZTe1tIQzp8UQi1rrkly
V+9I4ZQHDwwJ65tpRaEAkbyLOSQyMzVjjoYyMADZgGh5Cdg+8LM9k46i0oyOm3Ch+4GlU3g1W8lP
DnhPqHv87Ll8ShHBxfPV5fiPUgt7GOzwOJPGgVfegVAPb389KS2B6ClFILFVJiczsCAWMRio5+C7
nBcLCjvPxDMSyj0ujlNVt22IbbPlCdmXjaohr6JbnSe38iRd+XjdRp4hZXHHwDC981P7ASdG79sO
/sMcb2thHE04ZTOd/NLQ6by0QmXaciyWGFvZP7Zdnl2GUgUdnIOpwsHt4N6nbc1WKX46FeeMltuI
ZejNJQdp8jzXrjD75mX6/bztMIxg4jM6BgInd2faG9fCH+GySjoqzWiHs+8L0CvwE2vDnrMvj2/X
n0sIS5p5KsZ2MZajMtQGSVUXxBhGtc7N+XMB5QC+2W0MigFA82Ab0kXJKemNcnwaUMlAjo/Occdl
TVQadiudlscC+KmcyXe8WvxZorm85PBWiBxZEhOjzJvm0dOsqHScNIhrOa4j4MPfLhACsBEc+Ag5
oP4pFgvtf+xfwyF6AF8jXZdZezSgyWirClcaeMFn4DZpWzZXAej+AgLrknHaPYpfgcXnN+VpOGPD
lYzrx6U9qfQAcd/RUQKEdNgBUl7bHQ/L98ajc7noZZDlZd24iWMgcFxw14nXpEAQwl/9jYfZBDwh
8V2lJvEd0npzKqLY+xqXPpgOZOxsMoYwmbtOMMW6aDGlJg+pTs5HU16fMPa9bb4VP67P5eH4uRgR
F3yQOsZCe73/1aMomi5A9F3ApR/uxJGNQcO9pz5s7rreL3RDk+f8llfhPB6mNdPtkEXsmqUJN9jG
HHnGow3PnY3XkbspYJlvNKeuwShCkP4xKbbzwmVGxlDuGrB+qE+RKS6Z9AxwkdQ2Rmjthe+FYZAi
jB4MVu5A0Zx71gqGI5twx2I+xTAXEzd4LM58ovJAi20+Y9hV2KrcfuMCcD//L6Dynoq5Om8hp3aG
l8UUhvH6B7BEkcecQgosya7HyiPl01SggK9UF2/J8qn/gTLn2Z51B0iOxzHy3PPOm1MK+9I4fSdP
p715DKEsxqWJkK8Fp6LGQeSQEHsFc/IW5eLOah0Tygn970sHs0wKpuPeC3sjzxYxJJwCUHsVQm34
tOe9ZLO5TjvFvgsuYE+IeA/dj7XCfYKjd3Jk46fvCK0M07Z9ORvuR3rA2WeGXgSJHgyZrWinyAVr
WoFMzNL4Tw1YkwJRVAZHrMsf0SLwnHZHaKOIYKTnrYZcQCTOYa9pjUS2VatEYVOHkDEhVrSDJLcu
jYJwfbJHKluuJ1+OWPHWOFI+gQgVIlrrFL3cBme//xP9UljqKa4YJOYvQrvOnFmhInqcVmax2R/F
492mEXBfxg6UMe9X2UREPBECs133vFIu3uAIDe4iVKF5ZMy3XujEV3/4aqNmg+z55eSfjRLKO/rj
YJU8OZKJNGU3iOAVacukvZ1enezXeY/lNooC33tBenkc1AhncpoAkHOsHCD28qLkhH/+dM4=
`protect end_protected
