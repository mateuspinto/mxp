`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
d9jwDDeh+l2mQx9oDZaKTQc+ZHiWBQNsl1NjbGvbtia4oEerscFFcsGBXqi1FED2bwhrEQDK9dY+
UyzIq7tX8VMF32LUndB49DJiuzdzTNdRLuQaj5VwbuQymSaQ7a34wkBUbRbt7WLB/isJiOyzSvRd
YGqdLQKu2DldgRmLs0V4+xe91Psr5QEYqKuOPIYvilwvGGfe8O2dLijJ7aaWh1hCVPctny15OVq/
NbkxRr4fXyzMSgjU4GRZ6+EjTnJEg+zaMf8zZb8UmiLoS9Fhv+kwZQoA4oCL50P3mSBuBJflH2H0
h3V+rHRPDYji9/Udy+5gqlNYjLBBruqsKZLWHw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="amx/td8bN8yF8xjpUjmMv9NyI5DsNDV4vOOd3/9oWu4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
XTQuOWYeDexnqBl27tdrHwK1r3blmUheF+gTh7NUviplSVo6sPALzGuPi4UVcc227CV3iI3Do5P0
fp3MDk7IRve/AEO4kAbb/Ow3OWcOn5ApVKmEYFD4WmDD8lsbDZUF3jqwIg8d/jxtSeDTLQHLB5XF
S9C2xpZuURX9255+D4spcq+cWpCybhiLMDp51SE/D7Kjeqy57AckLGYuCkgwPktdlOcm8T9zr+lM
yqDw0vrfUVXFbLQoJOtjtVNefxanmlnUvB45zh+gtdO+TcJAtsB4YEU7dXlkPBmAoKIpInIZbwdw
WUNkTIqD+9A3domnqzyUTknv8jbG0OsQeMZn5CH+F77EWHEUB81XvUURdkUWFtw9SKZ4hCIGC9O6
FrF8WmeY4/KF0yMPhDgEqw6mbJDnrB+B68BUexgIn43uNeOP/QWq1MbCLIpf5qEbwWFM8GXKEj9m
iKRzctQfz2Q1itkCBh5LF/2tmPwPS3B2mqdiXzG6Kig0ejACPHvm0EPiqN3r3aGw3F6Uhlu9SW/I
eimbBAC9yX9STG3KSVMO6nm+5tGvZWn2RSq5fK/NN80l/d2zAf9vplm7dizm+vVwSOFYh0zcMqkP
y4QtRS5FFSjPWLdovYhSfm+FxmqxkJQwfxkKjosNW0lQIrIKaHuXJbkPgp0ZRhMvFyFBxhh0YsKA
sM+KoB50vnUZS74MCSN5r67IkEPeQkAf4cROVMhrLble2f9D0bScv+yNKKcjbVUHmfQVomLGN7J4
u2kyJvZhZOVLSEchW3epmL2/y3eLRPG6bzXcjWjJXpDnJCNaYBdrAtaud1pcurlnKb5umlgYYVww
LYwwxcFYPLqjv5d2rsvLbnJ7ob56i2eNyvpAR1FKdhajgqjDdFEoXfQRI4Ob4Vs831NOkg72N7AK
Hzbxo/Z+s85uBrmga0Z/rhy5AhgsEA5+7ivm6OdMwBGBO6mG1/BW1n40ksqTHsPzoWPFxzj+Up8H
k2KvqnhZ4hIcczwh2x8acADPsT09uLY/UBJ00NQC4hNSdmEHMDzkrt1Z/MX6g65PHB9BqSFaB2hj
fYyYJMBZAJ1AxwOhcS4VkUVXdCJkckwLWsI86SFzQ3s9uxa2e4jHFEI7UhksCAx8NOe3OakfwU0B
pE5S8i8FA9M5v9qV4O1tCdfuw73Dn/mrHsyG0Pb/KDmQLIywo+x/55RDjyjrjeQoxXIpPALbY2TS
7nP0bRcg6Vh2ryH1m1M/QgC9ldjS0Q3G8djYbW1wl2pbl0ymyC8WiPZxt4G3HSx+P7qhDvDvfjxx
ZpgwXUEBf8w0wei/tuSqRT4V+UASmkYUh4VowLq9WHmKocKHCJObbTzUUAkFE6RijxS3zAqbptwS
8ZVc0oCmOsA3Mu0C7D5WpiYGM59osFA/5PMD7pCfinlxUqTNOiTgBNoFeEWux4/KL7KLyo5KNXig
eSfDiCwvDlb/YpgDxSy/IAUeAgvgXlux7IJVGRTWOrZ10G+LeOu22x1ljFPvK0Dyh4dintsQJ71l
8A2jdgP2J//vw7u+APNN3iUOiYGLsSVF92af54p8StMbbsfpRomO2FX1SooVGwXdKT8azrkmwBaF
F+HxJwJs9wegG/5tQ+7rE4ezj3g3N+tTDqEgITzj+iHjT3YAMMepbYRiS+OjHOqSQCB6vAU/gys0
SDkY3R5g0Eo2AUPn3yyauUE4/DmWXXSJz+m17my9VngJ3GW0sIBITZ7+9bONfC86C6C2CqnegZq0
V3apPIGBAe1f/H4C2YnrKQuF5unk/6FQtxxvXTI6OWiI+6D9NxHPCQCQR1ubqnDeT0mnDyM0jc7V
H1vuE3gNG5xz5Wk4hfCDao4NHNyRuSgz4eO4Ms1+PtLDPVq0eW5NbVQwQmB71BS1zfKrzJIO0iww
6fAhIsX+pOorh0RqsIfRT6Mn/QHDGEnD6+JCZ5UDl8TqqSZ/BJ+uUcZMcgiqr+M9RWhss7TTFqwZ
LA+6YgrlYwE3/DSzY7ntAPktcd52k5fbq+XE8es/aajuLGubD1clS3oVv9gjo6tY8lZJxn1WivTY
kb99dHLBsXuYpSgschAwUHUSwyqLpg/7CGKQOG4M3y6/V+Vs+/reC3YnpULoaPLdPbKpo4nqd+Wn
5VWtStWtDZfcX5ot7rYljMuTkmtWNRttFnR7n/C4Ykx6b6vPsbqw7mymMFGIfJHtKGhNKmGjhkuo
u/fqm+Nsz7q14vas8AjzASMMYr+eu0ZXdSPRiGCJVSzQ1iY31WnevmTmkm6yyuWSE3DAEk1f9F4x
E4J6/uv9zqaNo6Hl9Y5x5eUTgVrpq8q8U7LuoOz7j3Ax4SGH9Ta0Clm3M4MRsctdgvA0yYIsWtnm
YcC5Lkf0p4X/ZUemiTSKvzxLkwG8tcpPBuRRwLtuCljWT1oL7PVa7KcGfKL3WfJ4YQhZYM/Ml0Do
stTGIlP3Z0RPkKapthbHivaTNk6W2Ez4YfxSCZSO47DEws89NN5X3+HaFYTyD3tjosga9hDmpDwQ
zgCeXQLQRrEXYtUnYSdh4cOfIPh5qFW1UJ1AYETMmSVEm+Sj3qcfZ2ikOBBYex5xiqqKtr4Q8p5o
hUqPrLJ5RXlcsuTtfhHpS08r/TdqWHhqXxNOx/Rbu4qcrTBjX0nSjPdB57sHEhdLb5+ihl7NcTKt
aRobfsRtDn6U4/ern4KhyOruXHx+Bsl4dDHfC64ErhEadX6cV7yCcNsPqKC7g+8v6G56An0btQxJ
1gnlIayxnvyqdFHSPQtmfKUoGwla6dciXjhAgar0V6HmKRwPmofWSykTGjpgpa447OY+CA13/S8g
+V46aytz71DRm8g3UHzwa0cP8GU/J2RIOZc2DU6FLz1uUMhSU59vafMomhDKSLljEsnf9Qg1Dumi
AZLJ+r1X0SB0R2VDd5OWqHfesVmn3axND1eAuH2ul6H8/DoRpA7zW1ht4YRftExAaSx8sTPjNzC4
WZSx28lTl20saoFgpQ3fA1vTQ0voOldmCaAn9f9wAwF/PS7ri7QS9lBu0HShJHUjuGS9hgHNIdyo
3iKYHrkrg5PkM3jZjLcrd11TeNZveTcdf8Qn1NGnlSVMiBnevb68n1LvF5cYcIKgAPwfu2gNqAch
Y89vUVjiBxrCWFQV0yeN4mBhjDD/4E6fKnNkfXIo41iZxf8TALh/CB5taTjJ4dpMRaJtn+P6RBSj
ds5h9bJs7Ns9bfnKt6hcPL6JdcBfNMk82EnVL9yawxMyJrpNcDwcPv+Vm8K058/7Ihl5XkuldQRz
aiaLmHCLJRpVfxqnn7lFyr5jpWfpseqklW01tc9Tx81I73OgpCjZULkQD28LWot5CsDEB5mF0yCL
dTOqh5PHrxvt9vtzkTeNr1EOpHptOMyx4+g/Wxm7MvUKYCS9Iej248DNa3o/Pb933Ultj//IIw7J
CBU9BpyEcNr7uoBNXPuKRn8W1OVU84hoBBjJXrNJHc7iRZpb/KEYlxp/BS8JM1G9XcDFToD7wh2h
2up5c2UokpFjKl0oPJFVSom9i1QEd6niYYrdIT9S56Er2Mtjj/6sTwi/ynjNsqhFYzxkhPZKnxUS
4bdqmJoeDLGXPUCCyedpM+0hJCJWlcNzXbqTkRMCP2HY+NMTCAr4/hgs/xxps2a+Z+CC7wSaj9Zi
GSn7CC4e1go59M3FMM3sIOdHCqD5KJ7MgUtTZBvRCrKpB+wskVICqH0CFMVeZqDjWUI4GC9C9ocI
gjdLO1fBDTclNvCUJVwTwLMtFS9Ur7gdRfRI2zuw3r/8U5E/cRw2MMCwfDPfWXWMo/jT/SvtDeFX
DXWBUWtmKiLooWMbinovL83qQdqFtR3sDDHNlpPPQbAoZF4vniSU6+MMsX+u/8iSFhWbsusG/8OR
9NyMs8M/6+XAHerPOcFKMFi2kQzHl3p5SRD1BKVyqL08rJwAmJ/eosw7CCGrJUXrkvXqxiGOcLKz
HJltxQdtSJVFq4ghMaEgUa2hmXfmPaJRK7stQfhlyFjchheky+x6+6hujtsnM+dS0MpnbnMeDe4G
HvA4cY7BXNhKmI3J2xVrGQl66Zo4VEHImwip0Yb2MMm92VYP2g4O5SWHsc4d3nngDPoRrobPqGUN
HF3yv1MynY0ZQqK2wS1QQNr3My2USGDFCIcUvRUHIdU/E3GJQtpGFJ/7LPX7EUdKyIOXslXozQO/
aExOYyfvchrCwLo4aiDm+Op5sTnRoixXWul0wOPfZmJTqJOlqUHKitiMhoDnq0zt+DzVdND99+u6
0ccF2xJCnOyYpOM/+qE1gPexjKEEkoz+TN+cSJ34gsXGvGH4L42M/G0uhmR4ZHrOKZkslo/k4Wvx
/40WQDfDvPXCX3BLljb5dFUjzUG1miFTb/gPP4884oOasA7HATiQBuB7Ey47YJS2Q/inHaRNKYXe
rEufkx0kz4hKpvnabBEz0dRpfs2M/hqzjyH0YPvoDcc95HZBjtrMMOdnBYy60kNuu2kHOomzrplV
xxDMOynhI79RKmyhKctT4L6l3UPxZt0khlZZ7R0J8JHEjYtfthO2lR+F8/vtqAh28QpvTpzEZpUr
PtXP0k8JeYJkY2xLqn211ZVie+kuxqTBptfItkb1VW9yP3+R3HSPxMPrOdfsO9/Bft2SgLGXv/4Y
op4BYKa85K5xayH07T40U064BJ9grdzAqjdCF2V7OB27eiSA4iz3odWVqrPQFSpnt6vz9nE2gSTh
BoKxcSFIyzkt9lDL7vLdbWcOLqYrz5Qy0kULZatx50wUAQOtvTfQbYKDrQ1ORseEGn+EA11U9Tda
K2Dw2Y/us6WoBR0BrxD8eq2Wq69snnUsEzKZKPwpwPhxDVLhrPxhpEwTgiYZxiXvOZXGLXp7GRDo
JiRHfg0TRtWkjk0WuUZ+Hj8v7QnIFi/MCsWQ7SKrncMgvFASqwXV5XdOdiuf/FsVMOsPH1uSBjr6
7r1Xf0Zow7I+7VXrxP9w6G96lWFcWvdNv4dzOLSPh9oY41GXhu33VV726r3OggTPvh8fBB/O32XX
nyqt0GKvS/08hnLpYCZF/9Sv5PGXRNEZLjKGQoFHYor2uKzoxGsTTqpt4Mdsnw5Vx33j7QfvNEye
0PReui4RWXhly62MfQ4oMtpAIrlm7ILuihgEXO67s/4gBguETT0je6dpJK1WKnf4xLXi8iGX/kd6
7FhKBh2S2ZGNuY98YnAWBs8Y5Qz5LfrXdX87Pjn++jhFAdMKphyHRNyhHiMItSCmzjeQm/MM5fND
aOuHVf5p0q+EIhsM7Glhy11WDs0ANx8RZAxy9dlOZFOJmn9h7F13NjOG3lsbiTSIb7cNgarDIS+D
WxmF/F+xHeJn2YI1dkxSXVa7pg2cMdEx5P94eMuLcxT1PnWaI5/5/dZhO6Z2yDiS+q/l3bnxTzdb
p6Vj/bpNWgp3R5VOX6voc1Gno7oLtiaUS5g5nKqe05D5c2V8CPnaV53/V8JJy7uvvCORDBar/Dgj
xRWrJUMOgn2q6wgXWh5zmHJeuKujXOietAzGQq0zR2UKiw1czDVWazmrSHVQzywj1B8S0rh/OiTo
CP44+2dq6KvQ+4x/ZUSwh8gjlV9ZlfxHNQwOwdQqitQ8aF0KgsrHfRjH7vlTACCESpR6voB8BG42
vs9hS+Khb7vwy6ntujz7G9IudnmaMy3W1nOps7xqo4v1TdlVsmyeCYXv7Dmt2NvqHVZIPpkty57a
280Tr1heVKo0nU3IzDBb+Ejsb+gBgPXqQTNRl97VJmHDx33ZZNNj9vaCk9YSd05xvU0IJEOMnweD
gR/XqFDPmel4UOGWj7vSO+6AqR2NIah2oYo/BzN9kK8FzDXaZjgiNKrfM/xtcDAVBUFX0BBjC63u
9MH4UMoAfSEPQcWC5jRuwf3ph/K4tPFbubYq0N5zIXId+Pv8+mnNwSJJkhQUH6Hhcwp4v55e1knB
IJ6THya5KVUSw5jl8+aICOtA3EImJLO9qcDxnGpVk6+a8fcUE7afdBT3xYERICf4vhjHHy8WMpXF
kusfxhexseebLckz+v720TXyXB056C4Yf7oSk9jgftvGRmt33pcotF7a4+HTUQzQK9dflPEl9U0u
bCMjHGYhk06XUkEV/rA7MEbW8rSbIJ0l1JojXDSZT+SKbwpF3AIU5RnV2Tqp85O/184KJlAxB8o8
ZxQngfQ857UABWEDIcF8tV4F2g1sMSWGq7TEb/Ev51tbF8DB1Jqh23bx/Jmi6cQsTcr409u7I4cU
FvHtwcqCkW9q1YCEeXOQcAZtfXR/gnfAgubw+WRvm+VRKdDL3GuQIR8KXGvbse5HmRtqwyE1owOj
SGZlWJPnnzHxs1rjD7CoXIwF4UaEDrkGJ+iLiCVj2aHHNr0Uc6o2r3a5st/rP3uOwaZpL+XegtXB
YOrRf+JMmaee9uJn+kbZEY66IUBRt9ESXpYO3RxzdsQKypKGefFnLtSQ/yiEcdfLEaOPacGkvZwF
ISJCyPLkPw0RGVClsv+o3bth2w4sxp/GGQAE6tvKDNrjgO02l9EcfHv4qkwhBfPS3ZzsqfGJ4RyP
kxCAU5y4XiGgqlW52v76qKU1wwfUsxjlMMKE4noHkZreJFcoG1yNgFclcHsWda9RyV8uDpKI2Js4
4gropLnoKjSalNx6YPe59+TcJGcKk3/pLJ1D31eJhmjSHtcW89oEYCngIPTZdA+JRdHytHpr31k5
fvyGVzTRfOszOByTNKgXCY8ni9IUKPj7IXh8LpIvF1Z5391lkbYjE+RtHmM4cT51wZ4CoJigAbt2
FTZfnDpxpXcD5IDENdIuCOoMIgcf31ulsUms1LBrCuCH8t1E8/HZI4glbImMEvCTrX+5rJSEV7xH
JUHCwgFP7ZPBAlzY8dbIkIQDdA9t33ri2aqT+jM6G7EACYUL2/N5Y7gwyHizIDJfkaRpGx4B2U+r
xjDYrkMZSOJ52gKAKHJ8r2OphRtDVxGoyyqUIaBEss5ImL/Tla6kXwCt31wRRbUnKheEdMAeVPRi
XKyeacnrzP6uJhjPrsvJNvwzqHLll7gjDRdfxjBnwG0CjALmzrmP11GaaQ8lwtCDs+AiM0f/ofrC
xwyNb4/hDMUIOFYeBzfrv8PjppOHEuDavb90eI8IINZuJIe1ZUIjZuHcqsEYPJBZwH0k6xkBOO5L
/FQVJQely8vCyEUZ8kgCCoUXsIIqny1InIPEMcZcx6PyfOnuLSSjd3U5yCSf7hVYaG4ofQSjuJhq
pDow/o9WFsUapXmseCUkOrFjAyumKQF3aoLmJKcJpxK5pbuaNbQBtjGVkv8ER7TYINBBi0OLNx/T
7AttG2nBmAJrbFlWUtmugPJ1TzRAt5Tkne8+FWLw3ftCtRekSDvqjdDZSjHYo8vE51OUC1WubizS
BTgC2a6Q8TFeYGtZhjNnqiMOjSqhJHbIpd3PCmLGhv1DrNgdMDNFa9szhFrJnAzF1fxQsKVSSRaI
VmcA6FUjGFs2v95kR8I5DqXVFhBTi/1QMnuHzHJIuA+ppP9N5EHlfHCQItWZReTRT8V/mTmrv9gP
wIUvGbsALx09R87qaSvdHISbnBXndYQ2wzg1HIKob2Zbcs0U6m4RoqMY+G7Y6By/EnBqTpk65iQQ
3U9XFJ9OCMK4rjONDOKEOzGsDsCvMtW8zHxu0jQHVgzxaHPwehFwyYoOOOGqdOIUC9mPwb1bU8cQ
yFaD4nr36Bb0NJRjzzWv8akefNqIKC/fL38Bpabu647PUVnkZ9ny2R9BG9QlxCb8Dm156umSw/PX
oJjyicdp5XD+bAU30xMdc3KnjzKYmG8Tgpdv6O7Dud4ljZ4d6vFF/Itr6yXODJ/1lV0DjTyBwMQw
W/HqlAFRiFKuxBn8AVT5yu8WqherS/X3BQ96HqiuFlPB1rYy7ugVYS8EDJP5fjj5cDKTak3bFU4N
9bM2wPCAB9q44LZxtApvtLKo29rovI6LkY0CgOLKQNdKNZBg0cCa8cC5LAu5jciNuMbAvqPuEXev
NmU+C+6Q2TlyNHdtanYLWHCTldjwibEIl/t1zhGKJ6pzf5jZWkq92sRFc4V59ERyTipZ9V2puRYD
yEX7jRJU5SWFSL/eoF4jh9j3RrXClkEJXbPXtHl57mBrsfkfOqnmU8MShb2Zl3LguxT9e6vAOtto
SU+3DzCtxNe4A8qkMkvhQv3A8uKEL2UG1ci3vsGfQxRX/YQMMKQSn6HbMY0UxgQeMVS4YAFap8YD
iEsSTf75wTx5z+U7QCvijvY1ReDAZYFOPbBUk6c8RAlaUEXmzq9l3/mgTWnwKYHsJB8l+KFmj82n
jm06T8i2NdXPcUYQvrCaVIraNDrqdJPbb5qNCUl1o66/nE7Hc0ajC6TE/kA8ZL1+wy9Nzd9y6nT+
KXhHcZutTMC4qbwC3K7f08bgvwf7mfbv7ltIfHO8K1v6gZ87vew576sh/qACkO6qFb5CuRiUmSxV
1jP3qxOEiDFPAKNDYTRY9uTJmSWz6WJEwxaL3kxZsKhzilk0YjBYNsU2GTz1Qq/6Ab7X6QxUuf+P
dXaQeVHq2nrelP5jL7PHM0ufhyqTJEtI5wAd/Xpfv/2YqxXArlZikNOu1zmRqkd6WRaX7ktl6kbz
tLrwinmA3DlCigYwqpQlQ9j2NSBbcHOT6RukcbiFsqcycAi6ptMtHVQlcsY2FYBlHW/eN0zaMpC0
LQ2GRAtk1FdNwdbPdUMpERVdJnYxXQXBoAIfwKYgBOiRSiiWa4SZLms0Skc0aCwatfmrFQbYO8Fa
17PrSd+XbP1s2BGxolvSVFHoOCFRPHJrimIoIH6WOg7usgFfPG6gjVaoYRLFAWyCUyESceIw/PvS
x0g3gS9hcWM/VJfIAdyzO7UDWLBH71a3jNjNSI2rHTV4OlvCm6S+h82ceYmmoVLY4ZRiyUN+y7De
GxtI5sozbWEIDsDYDn/DIdqleXBxX0qOzuT16mpcOcSIODDc8a2iPMq1XpdVr9qO2oAGJZqOGrXY
Q/9TZJUFjnoOcV6Oes2supq3JIkA3XdCEAOyrqEh8AxaR1Of/BexshQnNmZZCRS5+xr4DfYMOciy
9kphAmkzlrbrNhWOR9OOqgfbLhzLXhyHFD8Gg+gnPzUX4wrmvT9yAUmDm7fwOfQm8KuDhXgEMlp1
eTBufYDVJNdYEjeBFrMik8llf3LFcSmMx35V/XV/ZRmyzYopBqNEpovWe6TzyBVEZIzHzbtOiYJ8
nx0MDG3p4ISLLvZcWpzslYf83CwOelGJOQbzJFxa7NX+WpXxIggAEOsIRmZhnBTdChOku5C8Um0J
arB9TNu8fvGUZ9DQXkAr83W5gfdIA+n8AyFLf/6p3NS0j59FW0sAPHjNmDt9dlwUQBIzuoDppLxs
d9AHiKfpmk9Kgfa90oOq4WMGdiQKWIl09s3n8adUWnI1EKWHw/2/F1IWwl04ZpzIr7TLBYNZzzJQ
5xo3I7S3RVeSiOwlj1sKWXHtw7VWZ8vmg/LQI/LqVffgcyekMdbI3PW0MXLfE0byD+/RQkXtnsV4
+V2qsXlNbF+CTHvl6PTl5qi+n8z3myGgMuT0U3zB+no4FCM0Ak1uiRHMlJRpSvSQZ+lXL5e/aAJ5
uLuWXMmpMhIaQt4k2JIZuh9DRlq1LVfr3o6PJt4Bu6/zYH5ci8IrKLTclqOpEtxUtd+Q8yNjpVFU
mkLMC4dBqUUubOZlhAwOoSGQy9/8iYRBhPHVu7T4Vbt67IzMfD2mrOcDvT8DGK8kZC4F9u9zlTys
7Wvx5LAORiUaYIUnA+bjB06hH6qjmArSdyV84ck4MqcFhh8Sxp/J+aipn1rzSjWOmOnAg/fb8+6k
E50mcXukj0vepWS60QRrsspngc05Qa8d5fxBoPa5LbxGC2zs437/001UkkCF3dXdlKyqIDLbs5zz
S0L2e7t652JhxhZ1Mm+VlP1RojB8BFzhS1lM9KkdCuDTrNMIchItksrA94dWcpiH9pADo2uue57K
BcWcKa4Qrj1zpq1QA7ZeXE2qlOR5Q4pjP72VlNERit/iVvI0G5YAA1onGSRw7rJJQJXDc8dlSPwQ
/ITWPIoumUIaMppRlBCH9zG2trxrtU59cn1z0UtsNtdm+FoTn2EK4wXc+k+1cEY2sWGI08jRJZ+h
Tmel+2fPAmZsxRVBILrjCv2kaTXr7DSFui/8cIVFZu2ZYoTDV0eL+ALU8q/DC7H5fnobYsQmmgut
ls+5YUNDLYgWGr84Ez5GWbvbT86sf+SVfCXIzJDVYEqzzw417HiqPXyUIokU0cat9wlel+iJbNT/
JLBBypdSuO9BzdO2VcZ2tVGnCULZOrb8rP7AYeAJ0CmZ6/2YW2XxYXFLQy45BSUc6u6+QITXfovg
hfwuTGQt2WzCfVYa0q4Pt0VkYzaaLpgCj/9ajotB16c7JdBrBpe+otFpYwexwq4fEz+QQ6D5CEUO
h3uKFGL6reqAV1g6wHcOE1ESSYIFGHc+OtWq0HQS5e4r2prAsvbYFK02LKKghHo1w+fDQC/xIik6
hE3GUzWOUUVi3rzkyNsrWhHSfiyKrFdjffbrzosp1egVFNzfuYed/w/0duCFCwyQB5rVSvW9XSar
hMmaodnlungTPO6y2RNNzIARx16hcmI3uPvLgX4gz2ufCzn30aHIon0lO72inq7qDLriLmUEytTH
w9pS7lB34t3bWpMFem/25xxp5N0pncWuwowkeT++aWS9aruHnVm/HtJao3jldMaPf0s/0k+j2AF1
o/Pwd22G8W+UBi+OOtysq8Ieo029RTTcPS7usrGQ6T9pyeV+lYmjPexhmySsEuwVEsef+iUfuxvQ
fFPGu946JxhTVRqT/gpN/dnGpHSxzdh91V7a7Rjkj9X1AC17weLB/Hpgp+tD6xRDa4q/bwizi40A
WXSEhWtqajg/c8E1/4kIZOGzqmop76ilO7sH+wzjAzMK5QgLV5etZmiOxKIIbVsh/xWNP17qaHnJ
36XKxndf7+hFF6gPYMW4xGcHWXOgAUglEm2YOLO0I2u/ZIgNROoMW6fN3zM6R0iU7k81Q7/ljBSh
UDLbLni4kxJ5dC1vKUxzEj6XJToDRDk2+FTzuunu/KAvGgvmXl/1CRiY+4i0ewD91samEwJnTVTD
Og71cRlm1gIXK00akZ/X0fryigtInis8TFK/O9VyAL/kVI89hiEUwksejnyUA6cDvUNeKclGpLzs
xB1S/tSY/mbpE7TyWi2aPYw8O2T1YdSrOC2ZiVIGwlQ9SoeTYFjsuPKKHWLxIAv+wI2h5fG/5o8t
l5d+l8M+cOB579Kx52/7Ihn/kF8DNeMLCJT24d/DSGRp3NmC7KwuSDqkgQSrtSebFsYNizvzm9bX
9mMdyJ+/9vR0DomYFejAwPCOoVnwLHkzzkzKzy50eeLYR8SinK4+Yk3MO6MH6wGRKGDZePCpH4n6
eKu/RG6ZlaGYboxLnZl/hTL4ZijMw9cKvI4Ndy66+TYU03SnogUnToWiji7/h31H8GSF6seNxFHi
47URTlSMHQ4E734QnQlobg18h3b82sfbuquqW3+M8sgXebV1jaE7H68TESJO4E6nq1kGIUzZhz9F
4DJU/sh6VH87x/LsMJQxRcpQc1cXa+wfl5hZ9K5lmlpxThlRVKjy2PtSGK2dsMwciS3QZOvDoge5
k82oO2vBSAr03iHMY9Bmd+3Z/xGvBcj/unGj3PWaz9QvjerCQWEsCGAF+jEv9Yse2w8BUmbK+GA5
+LcsbqX9p1Ugs3PJD+Y8tvvdiL95ByXQbHNJ7wTfd4vsppt10SB8J+g9UhrHGwBPNyKeaFuPzNJK
ZN13Jqftdin4sLeClWEZrT9uqVRUz9/zvW7fJFTOIzEBPMQIqj2DJhLLvl6ug6ChPHKOG94qck+W
zh0jIVpBeUe0EZu0dzXR3jzBLmtT8AU5V6cHXx9UZ1YRZyFfP+NCwvSC40UxcxZdXQWxb4wi8QRC
DSRbwOSg43+pq8OVVOrYFrNNzyKmCj0OVupNlZtWZr4htAeYVZwGRmx+BrdGnHNB4NH6+SjnHt4N
ruO3Ny8WtvpQtuWEDqOUWuJ5mykDJazf9P0pVr0KKizn0hkWGbt4ChiFzvdZ+gsIinb97Hylbjiq
bon2jvogoQiEHxV5FXp4irEcM6398/fNGxCvtvcMWx2gtQI9RkyCiRNRldtRGyJk3pL01+gibvTm
W3SMBtECEikupkQb6Z5wmx3j6iZtFyjLIT9ZlqTD6znfd+KVQCROt0QyENLMtNOZAFxoyebUqupq
ah+3BS1+w9TtdjJQamCDhFviyPtydXgQDcH5mWKioR06Va60b7gAbxtE2C7WZMnARQ+5gsQDL2bx
MITpVyRfmEvE/AKuAOWb6PZmKJ/Gwjh4ZtJyqSBtv46zqSPSI2YWv96op1GlcyiujHLBXjJuteWS
e86+zXRXbSxIoVKwhqSDY9rZFAWdn4dTNepWK3Ci8yjA4wNPbnPbHo3RAyfJd2+fJ5eZN8e0YjSu
CP0dBOsXTYBxTZFPXz/V4cKae/mPXPKrsSez1XSMNhlpuI0P2VEWTkGPi5LYRIxKSmcgH15lJQ01
9Morsqi3BnpHNw9wajRBsia53Q2U4gkAewpHGS05fedZ6gGQGPETM9YITh33PkRmmB11ljW/bOXL
W0M7wlyMU3bXKs4NQESPFKXPR2Fbz56j6AVl/Gj/dwWwVN19Ly2yp8AhCRVRmbetrQNiUIEqKr0k
jDDqGM2Xdh/72j04aKaMV0LGRekgJ9gRZrZMOHVvPLjobRrwLKe5CQubLENxieXZWvx+3/2xVZ17
lq1UboTIvV+2lBXKEcifyD8KQNp/gMFPv4RS/rvzgD0oPGSM7V7h2JVmf35AJLFI9t7syOeFQ3Ig
lsx0V5QuM4Hasp2bNUqc8qjfj9uNFuhh7Fh7lTB1KWHghFA+jGpkyEMBtLxnsnJB0LpcAum0D7GD
3x4mpskShQRK86RDhpMZSOsK48Y7W+xAtKOfTFPE9r3CSmGb89m04V0OdcH+O2QrrlsqwyWY3kjE
7qC4lwr2mfC48xxgUimcPjQM1t6tw2z8Yx+D0POarTG1Sb/do03ymRvtZLIKuG5ScH74ZTaS5kEk
6ugrcPlkp/Jg7USZC0dpuVKyzmwzMEn8JZV8A4JStfh2roto5SCA4B7nSe3SDumBsR95NG6TxcGW
HNowB02VJxq4qaeqBbYjKfsxngOQGIzP2Sw5EuFB7ru8rwX6H3jMIP/ZPesHh22AuL6nD9offJkx
iO7+GuBddVCW1vWTfRO2XvFHFVgdpMDhKMxNCLTFTElICLw2lT5q5GqMcX2lU6YOxgfxtQlcfbah
j646oIAXAu6Aa1QN4+d+Pp44Tl69ntEQIRWHIHr0GtboTtK1oBBzAhQ0scm58QXiZhf4DyJmmC32
hn7GQtQuvAth35c1hyAf1UZBSAgOMs+tE19+H351N9l+u46BRE/aqJEoKl0BvUVYy9uZOBki4Duy
4wPav6VLg/98J31O9gaK8ywSK942VX6kQ3YjfP8ovotWcksjdg1kZ8fu0tL+MAe3XvJ02pxkjsGM
48Zv1HzCi+ZAbBHffcRTuJyaKwVvoSAXkmXnf6xXmIo/oyBS80ZNbnnIAgN/PYL9+SPPRd6GrOmT
O+Hxv91f19ljetGIZA1DN14SH4yX+6oq0MsEWWPyonlnIfoqbFqmdBhZ+pQyCawOGx6C27SmNdQ4
OY0n2wOzVQWydTTEs5p5cG9r0aGsv0leHTLnLIAz06eqfOqN2Xfd2HNwHVqg8yATqNNuik4BISlA
8I2MhIOQyTK+Lyu54D8NRdkUYBAAWMI73OiqNLRF4NP80Rjp9Iz8m46//SVkDeBkSY2WVNBYQujx
chHhcEvUAj8f3asJOmccQWFn/K9KI2UUeajo9hL2GlBSo6h/kcQyhdCk4PqJQsZNYtisIiegpbwq
ZuInbBsqE8b2UMJHfLkAc//rKb2Z1AphhN/5X6ZqKLO7aJ4e6pt3FA+qeKe8vymIzwQT2L+Z6sB0
2d8mO9Bivn6xuZoAjBscL0xmE3gsqaNXZjpfnwEaq0sFyjFSYm660VxKf8BhelTRO0h+HHxxNDtY
i05skXxcnL8FUZV7RKv2pGhwft8REo2xlqhPeZWYa9cWzv9zksi9CBUllU88F8Dj0Q+YgRZR04m7
/xLtqWV1oD+qBjfh0akRA24VIIt5Ea799YdPqAyPcWGpdagHPAvw1VWPLt0X22anzZocUoAKV/mQ
BuIZDG/HVzf4ak0oSFyRBryEoNv1lE8kDbYjS44roQjl6u8ZR23tLFU2LyFEgeViilopjIidteNN
t9PYQGleaNasJRDNbJj2X5CjV/Q5izSN+MRkRDfdQR63zhUgVBZ9OHvwFohCk3BaZcaD23hIcXCs
jTYK+NdKt4iL3SKyzINh9qY18zmYqm+H54ZIxyDFtsLy4ir1DpGoHLLFk/hv5j/2ENFpEDk/8ar4
E8quYsWDlOktynkOSfjjvwcB8/geEGoaULP0Lf9IBg0agX9vt8eIcxjvf//aR6x8ic6HmM8tFGqA
1XC6LqKat4CC0LUzg0YpcMglMVOJWtrz+gJ+M4OkJWh56JhYjyOrKuZ2RE25dD65wyr0btAHt7Jh
B91sihDTLkH89+3cdywCA6aLvUkLoOadHvOk11O5rgUR/IDmsQGsAss9IqRZVrvBmNsBR+0Re2aa
VCSVFugt++omx8u5Jjv11rbMB15vlh9FTrFsWUEeIBtKWfA9nYUhVoDA8Lk3lW684nXaDkGjCbld
rZliX8oJ2OSNaz7s2QePbw3nFwTcYFB265yAdm0RqklPJjp2kewWq9QER081RJV6hEXUivV2BLj/
fwu8NCqrwch6RAkWxMJRDsXLSFnuAKhI0RLq3LEfdffQRTSKOzhpUub5UKgDN/xQhiDLYmzmzNWn
SF6prOKDjXaaE7ECrU3lFHWnzgyHoBRMBgIiXZZyaH1hTltcotxXGqfmVemLFeIlMrfHtnDXrJA1
M9uGsg30Icyigyp3PNL0wn+nTwCWZRfPYi2iAqnFPcw7CGfDnCGFpj8UfE4xSUokN2UNbq/GYVhW
DGTg8CQ0qOSUx3MxH/5HzpEec/55L/PbOgcXy4/rABQABhcGzJfqBJDoqyvjRstJEMdSIa9z5XEG
ueWwfaIfqz67IHQnG/9G6TS+/DfOprTww2JQ0JPXbnHQx91OJfXakxleAwmxkTx6b7LveH/2evoV
cSL5nogaqyNAmBk/bWrvQ+rM92kL2oUxdnx4D2qJ6NB1+qLPEQHkwQcP4ejRW1N3Y8Fzu7sc2LkB
CvlKENAeLq0CQ/q/ZAG0znsFlwLpcJWCjTevlX3aJxnu8fplb+wLBVlMIh32Hyw8eZuwvVe2SYZa
FugOV7UVMoNR9w5fN9OqazolGkUDQDku35c+5Nf1WwAmLoq2yOhpkn3rNwmWwC5XMjtmCPwbYLYH
CJDZ9ipCbzIin/rRV525tgwI576oNpWgMJSUAeDWrPcT5J6d//3KGyX5eMPAN8w83j0olH7cuYDq
QLdAmkf9j4Dq3OMp4eMKdER1CNbZDigZcwOFpyrDMUEEx3nWBIWs0SgmPf13BIqHGKzRt3A6zpia
i2nUiit1uDOIQ41maArAQMTHvp4QyCgkriVKGmroc+lPh79OH6G/IOP267Ug6S+lF6qrlFAkjkFB
j+DJsIMEJn6n5nCNzn+FmDJDoRwm8BLi5hU6RvkSdcshk++cVLMkQAGL0AXcNyAMjMcqrU5CmVZn
Msx2Oxr8z+NRX/hkgbPTsnoD2KgyD6MxlotcWRn+iFlZjhpSmzBQvtAGlFyOZrYI4I0pamTB56GL
g3NojwaaGu5ZatjWeI4IbRxbghn3v275cuKNv6Fnttun8hxAzWOLZ30MSJyMBACTVSiBQENNzVAG
G7q2zj1J1OlbNRP+8soaCKw0T3lwf3mU1jruuZ2kpR8LNrkIhyvv3qxiB9a2uEKE+GVTw0AUIM1r
0pezE0LcOO4CfwKXVwnyY14cDB4LRu4md1IlnuS16YzrOtNKO22B/Pyn9zVwEEC4EmMiE7ivUpBv
eWOwf54nD0LNUhETMglkGywBPia9Jaa3wvdtOYOpTVipFb52WOJv7oJTNPtCL4VDcV3d4QnhF6oR
/ZUS9JgYLO44+4DNJFYVYeL8U+bIhoKTgF2O2gRy2rfwjhGgsUqDoL04MGWIOR8v4M2jESqTpNRo
re822yqaLaonbEF/E4X9gaZOZ6uAt747EzH85WTyZO9alw9G6znQCYJuQiTLkdxoUAmzOulkgWK1
KtXHJiiXDzYGY602ek07dmyne0WXzLy7WzrrViJAtLrAkl7e1nsE7rULI++T0+YmnR9gtqY5IxB9
sArLEyt/sO1rd6pst47cJc0SZzSPBzZoojxt76azVu8j3jMrk/MtQ+kodknLZr9K12Dm5dvUOMpf
aPjpLHoVNfeqEyDALihSFbKtnnalSBjAb+Y1kGwQNLVItT18rk2vLfQJpAX6Y7sQ719xEYoScNzv
ybf7m8b1xKJNXxC0y3l57Ds1bvtjsnYCNCWZe5VXjd1jKi7/zWFC0ZiPP7piNI+w1v/F3OmoNPTT
UxvJvx8VuYYaNSu5jn+Fhech/Ms2JLaNE3a9KSDwKr1oUSmjCnk3y2NZZqPz+csNkCMmgd25Eg7g
BAMPFwsC5s4eB6XUMxGtYqlsay+sQ0sBdSeWT//iBzXoqBSpPxR0U4e2aEVPAD61euGTwiBkDObp
tcQpWyjQv37r469LZksC6YmBKRMEcUKDY/gYym3fYCHvqOAqiGCTrS53idnumsQF7BFL1eL9J6CU
tYkX9zTiMmostXO3wvyk95OZGFEpXIPqT8iH06e5aaufZxU7BVBNdEMZryNtESFlhlbnCAbhj1Cw
QoXW5T0j2lETAeJh/euwonleAZzyM2xzIPGi5cY8+m07M4vxg6o3DhBu1YHmrwy57kFGMJDZvPXh
4mxq+MpwVgg7K+PG0n1Z0Ck49NPv00s96Ik9wst7Oj8qgBLysD5xtjSWF8rjuSrCGEfhdpFC0ZV2
jkV9J56An1BE7OxRUlhjsUhpPkwHWO61KLU9LQrAOAlEim5QjNYkZ+F8sCBN34f8rziC3+T6HtJ/
l+h2v5wf1XbmRJULjVNFuF+Lj27Dptxta9N1DZ+XF4fTx9ZFdZgeQRhAq8FmoPw7pZUIpXfpMwu6
kVs1ddB2Bvq1gjNLjA2CpoAznB368Qd9VZ2be2fG+qfgvQTawL/AdqSHNZkiN4G0ubC5Jdou/aPo
c9zOi73KEH6Zqr15pbDINzcXsFpCvTQOzLbGiBGnUOXq0d7s/HsrHn6Fm0GKC04LndFz0TI3EIc8
WUiNZTLrDIivGrNR6XhM009S9gCyEgepBkuaqD/urceqRzP+GB6O5zekZIaSWj5Kxm1gAm+0nZwW
CDYy4wvv30181uDaQOsr38XP6SGQ3h4/ZjSMU1to8PnYuqC+Myp44KIgpBcbRT3c1zKD68VOza77
auFU3J3K8GcY6YrZSpKaW3SzaKvO1uiFFUHrFDQlcqp+yEuIl6nJ2yM7pCcmF8ncjjdK6oVhniaB
8wBYrNWAs0KZ099+Zr8WEvDK9cHYit1QFUcKiEOqC7LV2s0z8F62wTheHVfgN3G+zob9H+An3EiT
2maNJihoLuiqF8O6YJtvem7kkyBnp9Hv4RI1ufNq7JKzfzW/NmqiHudizFuAOdsIoMvEhnNJYQ5v
vRk4/YUsAM1R8lWV20nFmLJpHrvbzidj9wzzdQ/15dzSK4w85YkJd6ft+Ioyutww66BtGAFvezDo
OUW36nQmgV18M9rV0hck+bVngHVDgbCdZw2IW5G+x6t7rKOFxmJm9CIjeHtaE+hMwZ/75QBsIu7P
BhBtVo3XvJmgK3mlXdUNWiOvCgUu3Z+U6ZuVqnchaGIOTsY5yI/18/XqZR2zYwViZho4UgC+h5HS
PvzuZokHFea+k6z26wD1bq8R4OG4LRJ2eItoIh36EUVhqCkgYQYJyhp4ktR30P46JyhWK+6wsAra
7W4riWzXErZNQrO/kRAAjBofgrPFlXgJgiVwjOyUcAyThhov95M0R96lK/BqRwFeE9a8vmxaOn8K
seLodB4nEgBoVqQOd5mFoDFUQG+6pG/YVj4HJjt1X6eXEMEg00EPr6zgsEo+P8apOh6vEH+41EeO
EoLGF0+J2sVUv/+1dgV5FUape1Zm/3J3zGVnKcX0JrAZPPmRymEZq2QH3yw6YKC3Jy0HsptoXJhB
xPCArtPtb0/8mkNU3O8AVJmmXJRcSlDn4DFTmzklTW9OrOTy1PZXuZGv4QtcLuzZRRPiUxsKKfW8
AFHxNnHYmsw+5mIfYDa3bFpslO9lkEledhaaU4W6uITtqAKeBic8kE/niyskYD8WU0p651H7PLns
ce36u4piRRU7DgUKBB5qeb/WO9L0kg1zC1jzdgnoGwmRhdpoPJBRkOT+6VpdVGEGiaQR4UMdUch3
WaIBdw2sCb5kInkL15bBIPdgOiuRZl4UnNTMg4WuvCJDZChQD2s5tmhJsewkTygnBXezvcxdVGDJ
CD/3a5q/vuGJDwrALA2JrrjB5BX/gx/N4y2HYt54XvbEE2ua7UtoiCNKB+iv9bavWdDU+pfTa//f
AVfaYErtmWgrYie3aQQAVwFXhP5UrjUCE7t4y2QwwioDznYYZlueD37m5O5sqpiGona8iNt7FPmQ
DuzxqseHLv2AIvOWjL5dxnir8sbxA45VZ2KokOCNjWoOFhKrX6AgY6bP5YvMROEy8/Phi/ww5ZO0
5jPVyhfwUwU6TEHBormccDpQdL/FVh3FDXN3hIan6bCJPmJ6yP2VvkNZfqCReeCPe+bBY1hiAvoZ
sQ5JfS5jIpS5afUBjriYwykjs2h0kq+Cabsx8lbn2brmq/TdkHR3HQ6ljHWNyC8dGQMkEoBg43Yi
a6nvnHq0GJ/JqL8KkI28s+wuALXhYa0ivgaKteXnpXVQ7WJK8Sl3OClu4eXB4Eevbyiyg1E3/D+J
qMpPA76rxMjDk/UrjiYW5hSQnMcgrcyWGzNJe7FnxRFPHGnGnMloutQHwSVPnkGAYMYfIyHP7ypK
0KDsooJ2W034ew/65QuUqtd+uaA10Deb6YMzWuuplZSU4vf5pcZMoPw9RoispKuzdbFTyO28py+X
AvUsmDP60CbfQ86CTxWQUzJCIn2oaFnj/DX3TN7Q/Ueb5ogDyj6X8WcHUqM5iIWrSnfxt6k4tWG0
5DEY33+ULi+EypmNxRidVHAeOECQFWa1Qg/LUixOtefH3UvBKnLmiafklWSvPjIO8142aTsWKbIm
+2a8PW6jQALDtsAb+fN7dzcZLxEeH5cQs69d6nISuQ6pFf+m9OJKnwO5C0q9A1TJP6vPDYATpZ6T
jIONE45u31YaM99st230Ci76XRoU8d7y5ONBgwGrXUL0o9iwDLMjAkxZ78T06927zW0ecPLIDofU
1Zd7upZ0BRXmqsyI49BUryvmwcxsEwU3DZBJknCm/1cSD5KV0Fzgmh+vAjk4h2m3lGAA1oZnj7D7
0SNwqHMyXh1XiZj63WE4yAPhKkoebBNwA5eCAy5BBAIbsxuyyk+2rHzO/Nze4SOCEgB8ihFijoUD
EBge1minCKkqCST1MWNV+Gnilslo3WJbL/fXgKIgYPDjmy7x0QEn/cPGYlcUjzG6SueIfqfKy4sC
DQntEGgRHzj4RfhVaqKYxJLlgE7gjtq8RULOu8KHxXVHIPEyLonO5WI9Je9lWROrq5TteLPnGP72
cWCI8v77YJn9FWASvKsGQhkHRBEXiZluRHsau1aYxMgKeBh2ghTRmhJbioVJfIWVrgDL2IFDegyw
2KfdjPqglck0eydCaOL24iYIUkRnfivyhs7+E5F3saso4vJUpB7bqVHSa91sAyZiSc1xWKPFPlUS
QsVi1ymQ7YntFtXzR9rCvsNXY41KJUuVBbgZrLDMG6/zJYCwJsUnYg9WUh653dgSUtlWEmAPUXxM
JWWPfhyrNux1e6eFOSdGjlUhiIEfLbYv8btaLwjZqxWi2/tp1+++qzb+qGee0QodYGVOXJvyA0uJ
YsRtsGASt+WTaPIaNdXlzU1IIdgFT3xjzrdHr2FhQYtc9J3kJGq3oT6o2AGFj6xBBhOzy4oGxbMn
DWdyKphN0Zp+XCRAk77mFrCbdF9pZds3oT1tHr0YxQYXld85rBJ7JBqYKOJ39Si4zYa3iEPK7HH8
LwL7qM4nJ8uAfu4KApvNMtU8eU25KQKN+O125O+C0riiwDTan0DbaSCqbQxB8NwRoiyks+2wOSNk
cF4AMfuX4X6lj+awDCI5L+4oCJlHFmWS+ZfYbZzBphkS4rtrqnuQF6lQuGXRMoZL96tM8czHFKiu
mJjKBFyzC60XmRUeUHZfqBbwb3AxDqX7a5ugkaJEdabSDdblwKWq1Qhtq0OywfQ/SAfWpo7bn5Mp
x/1h4uHcmOIe8DqhSSqOS/aMCu0HxrGlety0EbiXs6fxdUyJYhbk03jBfNoEM9Gh/aYmzDau4vfF
cFa5HZvV4uquqw6Lz6BysB4PBsm2zZo6D0Gy2250qwvcBpi1TnHiT4WCbVQEljQLkwV//o/UO5iu
A9wFHU+85NFKprsUwtFamuKmqmyHGYUeRex8y7J5HYNMq1swV5+vB9IEx6EgO6Slbu9PEONigaGs
ulfrTVXV4ltS7p2e4ucx/7oHCcqzb22vuXcyUZmbNDHv73edNs6qUaztZ+qziZRIDrmre+1lwJQg
xSHvE5kcljN6w4ALwSFGARlc5M6t/fmgBK7eE9JSTst7NdsFGvfxcJg5OCrD7jTTPqePbKT/C0Nq
u91+ifX4Jyf/nGomETYzNCE0+f9OEiV4Dc6ihRKEET+6kaLngvmjsi34+OVEa1LXKlTbdMvCcUem
kvrWEVxOpI1LlMu7sHHOXFLoQbvWJj8SV12tmp3jFR3T3CtwJ5EiD094lHXNiwHW0PW4FR1Fyrbk
yP3jq5MlFI2nqgVlmF5b0fzmf/kwhzRIsNpD8IQ0r4AN/gl7mEHfWKIWNTkzIOUfJMy1DtP44hlM
xHKR4U+IvN/I0j6zWspQFFJi7ZQ0RCRhiJeY7rUL9THUIVGAtsNrzkG03J540r2KwkBK40do7/md
mbfxZZYhmRV6GfIV91CFI1Zm32GxkO6WqMuIVC2XWLtHzqtmfTKGw1dTS2HnaDIp8tgABrD3EI0N
VvdA8VnVm2AOGF1jsel33LCHJBKZ6/prCaMMW+GQQK63QtrAb2kuhMGGka2iIItNj2WmkYLF6f1F
jrv5bKqx6hYDuxr7dLubpNb7Ig3h4a3gPwmTXbsIgepJILf+bov3iURl1cjdeUbaG8HUOKnliadZ
KGWkfwH995HGnMKRXqU2WyW3EnQqSVdJx7m0Be81qbEctxIQhtE7PFRcFB9qfgBdXnaHiFe97Y9M
iV5d1yCsizK2Vo1Vym+G9IX73KTztDyrLqAdA3hmmWKC7zUraOn4lnsa5h7QYTP6iOPKs9x+eB3a
tKQqO5bf9PM2rEBgLXPhshwMcl+j2kL+IOHIyL40Lomb7OQirCuJEKArFASNQOZm/bc6bcsu/0vv
tA0iR4zwT2IV7KwVWSsUf3gMgYEidGcIkxlj4Vf5oeS53la+DnVCRa2+XQJdhMza+JyuNQ9ZlbZV
a584IM2MQIBF7Mrr0OTEfeIfO09nUlEtC6pRjpKaW0HsetD8dWSNM6uqM4VTa0mOlK0vCxBT7EXT
5A16ZL3rCX31uYyPZB3NSdJdDas+QN7Hf6WZD0I4wuk1rOtPElmUWMwyQP1CCz7XFkl3VUWvTVth
Vttg+dzAqheXji3MJXE2y9Vbpy9rzvhlfGWlA8qsvGw4+oC9FEVgnekFsgfWGAkPhuHSFXZ1TTwL
QTfak9zdUAB/OUBX76gO1HDPPeSxKofR2r+Ihejd2grITuM9eSkBCf1w5Z95laD0QDnWvqVoiizz
quWqY1GRMORnlwixKkj+O0QIAtx66UTJhcsLkQ6wc2uM+RXPV9hBss0Sr6RztxJGTbQliAu76DDT
tIg4LWD0ytN+CbS+/UCyopWCfbBZ3Ww2qjddrF72JfcFzl74TAXrDtamavGVuLWMLzkuj0JDLiAt
5Ex01x/byQBiWasrYG6zLsVyVDsqs3gt3fRoHaKC6o55ytk1IYbV5v8oBjvwRk8dtmj4dsvst8J5
3my3ATonRkj160gIsUXfrDKaC5anH2va3mWR3yU5Snk6g8J2zbn0EiHP667URnv54zGOdp1QCn+7
XZ/trW73vSqsfh3upc3QCYri9eb6FL+daVrlKdgWJncXUoW5CfiYKUZJ4P0BIs3hMvrDXkljp/bl
J9EIzJtzBACRk/IZziuVyeKOCwBsxxOMFCvPyM3D2WTe6Letsx2IQEDSnwprGy8qYnULjcjSmUpH
FY8CMAijerdsYb+vwYPntb+4pCOZg87SB9kyZ9DQKcODacFQf+BueueFEZaSRJxKtS0kiAbg719G
OrAXW8SaiUHSPsRQphfL58S5Hc+YFLnuzn9Ldkxy9Ww5BIhLlRtpjbUJKZ44qaGtEmoEQFnY5HYS
PMKQbgU9IIx/wxoszeH5cRU+bp3o1QvcrjZ+eULAKv7ZhC0vTNcEsuv8+k1cSfF3/Ve4SW2sYqud
YZiHUfvNeKnkfG0whbi3G3W1a/WSuRwu5R/O0zp+AquyIybw/fBOYf4JRzpvIjStWE/JPr4E7Q5D
nHkAjGrtYCO18QrzUIZ/6tlTlvjRlg339rrvzMfMv1FLAW4dvf+CgBKNxelm+OC0ZKHUwBw4V/Ud
IypZ7myR4g+bmluAQfQWW/DT6Q6n4Mp/mCYymVT5y7w6CQ6zsyc0C5S6BumVTGcpRLxUpue86h4u
8tfPxTqkAjL+zjk6g0+4He7hGk//bD+4mQY4u0mTBFv8t3G7FfTZaOdX3OlX5H7F+zzcaN0mtkq2
4JfKNHWZ/Wi2p9K76DKfz6EETi2FTWWL0Y/v+kB5sGfJq8wHzYTMzWHey5PxXTLZdeEO4tE12e7h
cdcVdAcqFuwyhbzjoA52XAFMRPi0hZ0ya7wmNCwTJUR9H66Yknmi59qsHVfRfGU4dJahvlYYzMLa
NxFmsLGYUKOYKSdUfeM37+rRoVb8U64GVdRrJF2jEeo4t1mk5L6Dqj+3A0LaVpo/L1V6iaCvTQE0
OkJtLU8rI8k1n2bGt+FscbPPJjayJdaRZqiAOHv7elr2hlvXYZPPaMMhzphwk/77GMKoowrz/PDa
4Bipne6BCLl/jwxITWx0Zha3V1juKlYI6oGA0DFpxotJJRfAqjvH3vVKG5B/HsX09ufrpxD5ODY7
9xoVP7U2mCkTdkXjMFmwc7hmB4wpR97X6iEP0Xx1H8WXOctqoWlxVvFDx/ODximcJztdlmDTJEpC
MZLdmYrW+5tuiKDWYJmLnVajUSjfBmN3YQkelxG6iEiE96sGQsIQFf+jEuuAKCHxbNblXLmvXik2
KVaqGfhWt6Ek/IrM8+VdlaPIHccjpncRTb/49D0BxOYehBKVzugKdriVWcCRZP4PN46gRI9Uz32j
t1Q9yu14/jsqn22zArZZZulDJmtucz5xZx/KUHui4D4WZ8+Phv2fJ/IVaL2DWWnKvqD+22yz3g+X
wbDqP+v8BXOidAR0byAutKWBs+B+VeCiDic50S5/g0xvX6ca/zMCj88912UQ9wUU27c2Boz3QWhN
oBGRb3pK0R8m0KslygcSftyks1mQd+UGCoUmVJsqbdqyvNQfpovnmNZ0i7wQtQDA4h4sCe9IReCD
/YoPBpJwjev8fhOgWqVU5n6vDohruJ+4dvr3aOT/e1t7lLbTD3iPdR/0Pi/0JS2+U4fpMe78vUi6
Wf8e40/FwMOwe+32a2eqRLNJH6ARoOcu4MlKmEO7s+FekRVHzmR7yYSIhlzxoV4h2q2z5i5e5VS/
iSdzvnaHoX2fIjv4NgkssqY775yBoo6Wy0reTkDddQo7QcDkxwsj7MX5v4xHW/quY3l/FxdliWVB
tppulxqTvYMBKK8FvgN+QZ62CRPAOURQjZyCv+Y742RIKKCFZfIq994bNP7mSgTS/2wQroNbTl6W
oCT2XQpua0/v9MwWFq930kmS2ki2IiLPCV1w5qMkzZpdA3MvOmACZCxRep/uA+eFcT/vi2/diVnw
FUE28124Gh+4hKcgNHhucM7vlbqZwc6ei5bTis6P5T8e7vFeyQzFuu0rdm33VHmeS7qZYT+swJUf
dPrWLWg5OFbUO+hyLI86P7jjpkT9vQ3Eol/xbdw/M+9cXNUFG1+SA6OwhOhL9RVFc8ecDTxtkz/W
kKGwD5saef9pfCjU8i6uIcxHlEMvLxtYiTSK2Qa+DHGV2YjL6UMnP8eap8uMQ0REL0Ye9O5sy8Dk
6Qkr6P/8onouqfN5Qs+vEK6xWVzG8oMzE+X/j2rejxukxgA1xXYrsIBGW3GfzgRVw5h+EeEQ4YfE
aEEx/z8lXo52xW90OKZQWgmzBPy1Oo3CI6HA/Uxxo7aaIv5qA9bkMq413n6RW58AAOrRGppk8zwI
A2MbsJI05N+ayEWB3Tk8ldCUWkzT+O27bzsnqjMN1u58fdUXUtZ2Fcr3CQkmRhfTeXB5EBTjA9SV
yhXHQRC4bgnILXv+Y3y6JDZrYJ+9Pc4zhPr4oqPoRGg5ZbgX4gzRTYJS3/bd6eAPAiiuUtQtkDQS
zUKvZxx2uYdm30TUFFdYm+yoXwnAKn/vrbdVBG/7kZr0OOmSGWyCAuc6SEKJvCX6wolt+RaYomCc
wCvaO+xNmVJQtSQavy1TrwXKA5QLx5lY3H8YLZym6GrAayY+NEU9PHO9SrX4fPd2AWEbIrqaOP+F
z6IA6IlE1TGD5UqBZo2cV/aRpF2P3t4jN1OJqe6xxhILrqkyKqfJJTJDU7hx0aBcz73DGdz59m/E
B3AI3P+AEr+Ai+6HSdh+SHiTN7IZ6S3+9Xd9ORlb7XUQOcXMBnmx2FE733CLvw9Q7TUMfNM/GE+B
khgUcuMS5IrtyTUSVkgmH7H8pJTGM+9Ldc2SQTo8BDhRn5asxfU4VzSx4kGYcolPlNcwMfpDzhgR
isugKo0Q6dMuVyQvaCEQpseQMH3S4ewcQopI4qtuV+wl2BluYOIUJ2oEu1zPKfCX0RLcnTUnDkSK
pIdE4bmkoQKI6ohJLimR84c3mfAdEERFTQwE4yItEvbVKXghfzYQ9ATToD8n6GsYZog4cY9J0I4W
AFjkCwDXR95zIpIjDdnVA5Z2ILHXkaQmNnf4t69fAaufWE34RX6yYWavU2y3geniXOCvUs2kiYXM
uPi/iNat3MVdHll1Te53BV7EVxdzgIVBst/oB5OSYPJOp4V6um+ZrT6gHiY55hEaRRU3KXaDud4I
+WeLlQktrG4jhywbjlyu7GNK1EIcA3pQojsjbFml5MBcaY8OaKhwLyReyOtN1gJLaQvMLJCS4Ga/
jpakK+ihOIH7LqE6y1yoUmUT+/SteWwhb3XdryzN73BKEN2fdsqxaAHd0OpjbB8SOoI7uE9rRM8B
EHhGwnxUXIIgdw3nMTJAfFrTBxwuye77xdM4DzypqgQcGljq27Tr1wNdK1ead1BzJqn+ObZukeOa
2cWM7se01X1W6rAofPylFNXekaivvOPS2qL4S28KsnIHq8e7VT7vlzIePo/ILEASzko1+JS/H0Wn
a1bpDjxMYub5//owXnodPRo5+c8JHUyJ13FDo5/iFWnG3UX76tmxJfh81Ob0jfRe2akkb3tiBzqH
WRSBB+sjhIu6wuh9g0kbW0uRbnMQRjgYbeP4jwzrv/39F3v67W/4Ny9AwjEpbkLGPKaUrlS89Pz4
z9SWuaodeXl54fAVF9GFBwte/u88l17bkTtF1u718woWa2Q6f7/7PzSHBGftf99n82rvur9J8lrs
ozO7cRFBUb+/xDjBaH+B+7Qw7J5xYja14+Z5nQ3ixQFlUsZb4A3OEIXgNgKDUe5uCwAnmsBsx5Kl
uScL2q3S58KnoybPxxmvqstzxkYrQCB43ukCgG+Gf1aHOTrRoTQR8p6ady5Ni3fZUNGX2HY1IO8g
U8g5YIb4OGXO0PN+JnYNUKGdkSmoMR/7E51xL3xsorDirbwaJdpykVLZ+TRbQqOixQKiLlGc+MsT
330l/BzWG4DhEt9fwzJDhWBYeCBALYdykqi7oo/TJqggL5PdVng9TXq8kv/7XqlwlGE+wbUMd0VQ
5Hl1h1nnu/IGx+j6T+ydpfM/kSDJg2q20Mb0lX0w6+A4j9jsMwCF6gbV05pcqKkFnyytWaEUner5
VCN6bjrWJS4aeh/5DZVbgPtrRDLLI0aKUhKgusJyBIVFcWw321drhWlGcRjna/VmpQczNMl7cfrA
n1t7S5kBDBHmH6/zhlvvU/pIvsFjnql01ic0CuxEWyCo6WoT+vSqcOF3QUjOL8zj4ijDWj2qNTli
72ry7lBPBybSVrK2GJaaDDeSB/t9DT2nJkNY8UUB+c5VMOsCcLkExPI3/QPaXIBU0Pkm7uyJLa2h
o6u5bhvNu/uANAxLnZpQA/Jlf/Die7RPRHQujI2IvMcqI1ahMwxGI3VAmFf4fAsEqnLJjsdrnwFV
5ogOOwSlSX7GBMayMUn5IqV9ejELo0++v9mtzngQormJQppfJ+v/M2A/mEM32g36nWApl9uKkjlU
45fTGbOxMYZn3Fsn0l1ekWjSTsV7+NG7bVAnEY66qEbjKuTX6UzZETY+6uSXDaW6muGc1mvllS1v
xWXoroC8qUV2IHZi6fKTqqCV3e2o69IeKG2JSntHMsf6JCuDr6kBt0gTyzmx2KBlXDqGwssM+0Je
Dry2zQEdAUT9hIBLTLLAq5/TfQLSkXfj4N4e/EB3p8NNuJc2Su/NkotogsOGyiejFxA+oxKGmNOb
cB25TbegvRZ9JOzK3P+3gU+aKlI+InOKlUKh+yguAE0EXl3YGYLO9uRwmr7tSvaMLdLn6bAU0eRj
CMK/Y7R4qBdVCFRdkApfxVzOHsMPG7AeHFVQHyaed8I9fpcGSxt0hyl6CPT7Lr0ORLBdxdAgiCQw
IZEgMUpcHixK+FnOoRIEtRp46FykaVKQeD9Z/gW88ZP0qxx3RRexROdr0KhDd7ohXaLOe+S0O/SS
6OTC1KzAoujBU0vUmN/i6CsWccIkTl05S91d/05MDTVT/HJYXiLTE+FHXMVgz+j+JqVBtzJvqTa+
yuDY90XSK767XzluGfMeub9cCZ0MXqDtr5d9+tTjvFfIOsotUh7CsQJPH311GKMpqzAh6h75/mvf
JmmDz4mUbpahAWP+v8fwxfTksU6QfeOclqnxGTEn8tDCSHfRIgTWMZO9nZo27vnUYLRwovknUlmm
rADaz+3b2i58ZOCNEeAhQJSPa6KlG2OpYLF4fY5Ef3djVokLW1Lt/dEthSf+6BvNOhuk+okLqJ19
L7rckIsStNrvB0npwT5xNYt+qsH7OoaE9tMc152hlvWUE2LRGVsObGy2KOX859GSVwenlYieibe8
3BPn2IzpFzTy3yI/9j8C3e0cnqMK46hj7gTycRzuwKGJYTqAtRr0rIZxaPTGnJVHJ2TyjHu01NIG
w8J61482QmjKc4OKLCumT5UXx91i/YonmGqjjvDL3g8ClZf1ejIFK46GDAUuqqU7YXFRzIZ16w2H
BwH/8TtGlT3tjTzccL66ikyDJBTAFxMLO5a1CMyItLmKFJu6wWjUpH0ED3wtbXFVdL//75DxhXsu
Rc31nCeEd6mZFwf2dOmkauMTg5da6NcP3+Iag+JvZT4ha01NfWekH3C5QIZ7QFXNVDv5UoAlcCnJ
UkGVqXFAdBKlSVPwtp/89kiiGwtmcCh4IBn9laJaiLIaivpo+gIisXxv/pL+ODBvx5mAEZRLNCZ8
Yi8warmtpF2ncCY7bW78c8BJxGDz4c3tbqN5+zjYMQ3hMZEImptoc566pc3TLScF+aE95paMPPxX
8+pMSbn2lzjXy/NpD6fsgwGpO2861I0jEiOgaLmC+z8l9Y1KKIJCg3SR+wZDw5xZwborjw1z/aWv
2I2S+fTRR2Ls4Asti+3ouJw0tExrOxD5cQaXzDBD/R8UuSgdl6n4k/0P+PW99t0adIy6izhXPhil
ysYrWR+9x8cg0sFp0PFgcOvQ7AQGp1UM0bkvVjOLZhI3iDg3NlppaqRhUhQ8E1HzQzCBgl4l6rQp
6chlxQyyKDE/hdmTa1viWPqrNO4l1A6G8pVt+TlAzQVegbdFcWmU1sJA0VWvsOaBMsWAX61titDu
RCTkH23bYSvHrZlBhhaMK+ILsdASaXKSQfFTu7DmNaMo8ALTNVv2ZNqBnpR2uwzOOSpKvVNCYTwR
4QUFN0WR4KPz49qYtKchsIZpw2ZG+qbm5QqiL/W6Z8xbdBSyQuT4J8vGjduRpTNI4pPOscpBRChf
zg/cuWyNBoPnaKH7rONoZFWRzW2ZyDmcvGEKetSqb8INRJ2tk0Vb/xIwVdXEeXSnFxxMEJsp7DeL
Nx5kE4nV0TWVQ0mlcLznpnayLvpRoZqfGTdKE0NLTqhtyZlfTJ3KUmcPQekZnw2A+5K8JRZwVMxt
bECljTdAD1pV37aB3sbvXWRGvLJnUoeGPIci7IPm3XNzk62QhXnxE5PPMimkdgYigePJm6PaJCo6
FucTjWqPwBtyt+WyFVLSqYPvnDl8c3AnxzkLCNTLg/nC/f0wldEx9K9GUHrJWlQm+qyjcpRqr4Y1
/xH1gmXy5o2BcWwDl/Xq29KTKwFgH/uAmDkvjRl73RgkvNS2XW0Uo68r4U+JB8TVVUa7sCZKPGht
b8lA7Q+DWzzQ7vTjHOX7soYyX8Bt5mS+cEL0sdD7dyFR/dd/S7su5Up+4J7iS6yys40UoRKjzfsO
YXa6+IBOW/BzbQIgTzAMlvxVngnRDUBm2+HN3uy6olanbsofbAczxNFuWlId/qsO01MkHwurMNyF
c2nSeIvkaVuHxf9Wl3/oND7vyQaRJsastMt4//rhnQY5oBGfgNhlt7wWlAZa0Yg0V/XXkWM5itOQ
JCAMecPFB3T9QwtCkXxzuQ94Vrj83r0gGkV0baoULy0jT+iYv/IGL4Kc1RQrNu08yuQVLjhvpek9
gS3BRCEQ3mD0V7gtFBI+HbGoh1/VeCAasKanfAsID7L7dJZPfjGfSJsNLgkWOqKCLKauGCZTbM71
r0YXQUiH8Hd0Ij1KTi4aMMr0g7n0HKXIXlT3JQ2Nw49pxZ2IAEZkzOFY8hXsuKgNhM0lk8xYnfbX
scZce5UkXr4cYUX5NuFezzXSQp0+cAyRFVnTYiHWEEmDiPAoQ5RLdtByfydSeBd7lFsROKXU7guh
KxB8KZbqIeEqMVSEHT5m07R0kPzI3+wYA04PEG1a9usN2V1oABvzLAxn1cU4lmtT6c/o6iakycxb
kNApjDFhI2uIgGtyqrJ+9hewkkdKl/xJan0dydJUMFNurq0T2j2Veki9+EOGipuGw26r/YDz8hvA
7miR4rMGtyR6ZIne5J06D+0rbq3OwP3SRXFAWEUhPW5uFAJ601Cwhz7z868z8TJ86PiJ1XVy0qA/
MKVaXwOJz+G8+oTr2ZjAMiijOB1TkOMvqYeQg3eQnw0mMOfS/ZTgKjqUcNaAIG4Q2kSCIJilTrzT
YlEqlVlTfZ+P7tNogi46IfHq9CFwUID95DhJCGgzy1C7ZC1RjocTVp/2kpP6zNPAdFDFTat66182
YqRHXt66JltwZZLL53wZEDsYS0W1qh4B3mGBRo7w+52O6UGKi500J/NYmYbAhO86IyR1YUVNyCID
IZNvp1yUqn35qlfGuhqKxc/Xv8k86azAJh1Dx6G5tJYji+a7yvKnK8Yt9hCIcPLM8az8uF8ziRqX
aZjwX8z/Fc3ZCegC7P0Z9SRgjSKrNtSllD9sYuD3Ry1G8pJxCoGgO+okkFUPePuS0paE7arrz3Ct
7RgyXRJiPkTk3xDnqc0PWcClnrPMmnkq2MCIhWeo4mSNVEb5xUbOF7QRAlL/JiWhIhcS9Ruuy0df
WkXhJ5ZASGgiOSsXbtCGoEzOkGpaQ/v2fVP6TPF+Sn061jsY8V2bO9jBlhPuRMmkpHRz1sjH4Urr
aBKpgzCFFS8XYA965Og85N0tNAPWJG03xDQakO/ISG8GeJeiTrHqhRz1m5s0/702OKK8EoiMcuqc
x6LRbkFravrTiIl/OUUBvY7dZRc36JHwZ8XIQR/byIva1JOxJY9fsDmf8D6Djwf7WnEunILM+Nmt
LNrNhiyhjOFcCcH0wUTOWjui0WTcWr81taTXJDzu6Q7vsdeobHRSuBfeyjn92/uZtZrVJYn6eNnq
lZ1woLyFnrG/6kmx02XuXRNApl5ybnlDKuDQZSX2aq8LNIU6ODlixl3Q5EepKftRgm5uu5SqkETE
cjBxvWMx8BNeYvSnpa1Ul9JtZ3oa6Oef2aLK7zBZoUNnzZPkjSBV1CoZWsCstSZ45hFvK6IkiLpU
GeTt6w/tEbm9ZldhmFsPugiCxQq1lKV0qqCkjWRSOIhjz8FZj+MMGjwI0Zp3CROVCWdqif3rEG8f
Nnv/W0VBL2JFBrDJCcwgpE9NSlB55BBXV8FjtTgwLmBgJ115dgIDp1I1aCggdu26qYofwXkjIblr
5Yzj068pofsQG0gBJ9wGtYpLwus1pakij3e7tKeOop3R0xajPe1+KcOV5Kx8laXUUOPN3EMtnu7T
J/E5bnVJOcvGe6UHW102TJNbOyR0KXx2wrbEqCzCrDYK2FPOvouCeVWvZYEeppsSpkjo/a8w8QKV
f1PmmkF9Ad2qf4fkxb1nskh8oFVVzJWCOieyiLOWZpKt6Thohkke+clOrJjJl9RQQeVzJPCJepsr
AI6RIr2y4ZV5utnPMcyrP9Ok13k4HbBggebV13nS9E1DWpz/hAJRWJV1lcU3aPmFYl0CgIzvTlsl
USPUB40lOoAK3YkXR2g9U+GSkIst0X7v+uZIm0nusgqDeUSdwVVySOaocm7vGpWqEZ8+Wlo5ECV6
rrl6KvoVB739qxMDYpUzVOa/XPUtAdB/tNBEbwQG0YW7fVaLN+gco+UZiWrf+qDoNjx8FOYirEni
MDvMgJi0Ret0KOhIUx/RFr6zEoYJqloOi9Yi9/bUWb4RLPQyIqiCISBADUzaCUM8/+d+HR6WS+Sm
9D/OlEkXkZW3XKbu1YOf1ZMEy+tgeshtnLxiyytY20jydxKmYNkTpalW5ixLQjQxPzJcoM/5Rr2H
0bmqOz9NENrNSkFkkjX2MEqzsqiJaohKLBfuzGsn5ecNDM+nhugK3yWBfpIkTuj8w0R0o7pm8m3P
PPOVT1/4rL4+EHGjOJqJL8fRvknm/ZHmbCN/VVw5Q3AvplQ40At33Yn6t4VLyJyqFwva2XmfFZ38
G8mfWjB4JhSnSMF0ddZrfgsBXmX7rdb1mJrxJ6u77q+G0Gu4p0oTffBg0PMxEJVVH1DDm9MfC+nE
I8iUjK6XxK2YNjIDZs0y51Q58CBT+LPqqdTWnfZp+DavDpmWOE0ZZXK7YbWr0Cg5XLJvga4F/6L8
EYnsZmkR3kCHB4hvS3WCtaW3Vhi7LUseza3k36qGvXTWvwwCEmsR2e9rIg12SHDYvb7rd17u3chq
sUHlflgZnKhknlZv51ZKeZyaW4keBLk3gOM0LOOOWZumkjDcONErAUfomzJNX9wBuBuj17i0q054
SCkIWRw8Qb/x637XNwRknbpIDocTVrE5I2HBO1cYHbmVZjdc7QrlzmSL5Eptzm8aoeT3jD0jHIF/
wVXuXqF6d4IkzUIn2gQjHEbp2iKQI2VVBvqTAMFEPybq+PnaXTe5AnA8A9EXlmtQaQyfN8UnxBxx
ARR+jfuyd2A8RqIG4JVAgofgc5qyea+QKYbpobq0OeiLpgg94wRfKq5M56LiwjFsxkPsKDj6q2Jh
A2gfPHDOjdRVurLrVcNh0gbY5qpYzPm3zgMppTlgmTxVmjfPxIBUkjSe72L1ES/r8MusIq3Af3rh
PL9eLRWi9FcyjOskxeJcHy0h3C2f1RhdKcpTOFaL1TSoPWnkx5NxTYsmtlfVcL6DsyeajDpgOKMK
I/SmiyKzGo02SGfrhI8MVisI59uAciLt7y08eNQF34gEpyUzzAKhm8Nf0wE7qIyRo48hKLSfxTVW
S5nmGhrQOiz5A6yPrvSMOEI2hexdLJw2p0ALiT3c24rA9WSVs+P+986NcxGE4sTBgBug6l5amik1
t1BRX8eK8dGndm66ES5KjEg3BmvU9mapVlw3DmyScgHnr0VFw3Ot6IGQJrqk7T7qZViRrhJm1HcJ
fAPAMo9AI4phthkOI7xIrBxt/d33o1+QpKJtR0Ut4z3lDqBYREcJK8SRedYKHbgVEu2LPaDfKkiE
8/P+tMlOiNu0S5dPSIs5l7ppvlO+Q/JOt+/QbYqAJkeurpNebiornWmtVAkaGUH2OjRDfMr/Q2O6
Ai3oU29cudfzS2tb5ZwXxbN8CagWd2toy8S9Frojp0RfKJMS3ULniZrHv+F5/T7SMRWzytNR8CpD
BXynmWqGBaQ4je6u16hQPyquWnWrysS/iN9DAaVL+f9dalHHYofBxPPOkmcad75iUk+1Lc5Y4/WR
WQiOA8Fmco3vL1SD8yudWjLoft0MKnufLT4bsQ6eTVjlgWcT9hzQ7ZPpU43AgfXlzmlZQAX/fkyM
ukrX4dWea1NsUbzoLxWCo6ZlnIQ6PCcgyNdiRhBARRokh42NjDR7vRHAX/O9Y9p5ZVtfSS3BpJRs
g4QMcge2Im+FcpNW9syM5Xl4vMt6hTU9HLThRHd9/CeKZl+zw7iFqL+JMfljsWUiidN7hQXVxPne
aBkZgvmXUsHTMw6LmZWbh2b53OWYKAbSyVM9Nq4xvc+4hdV/CxOyjtA5Dp8vz0Tefc5qWiL9O8Z6
yFxwhpE0bJxBGlgKPjVG5U/3MHoYJvq714EDvfzlqmH9HVVrR+7JOKx5U0F/5JtWz69XLMfutIns
1MiGqmsKMJSlEHAfDpjpTXxTX64L2ur0aziF4LPJb2kar0fALArGSq7JqHWYR9Z3iz/nviQqUK2n
0IN5UPk1SDCMdr+bx3JVTISVStAOrjRl3+LF4ESXZ9coMKzvKCgAzI0v6a3lq+MyHAdSvbS7TaPe
RxtE3qN2YmYtmGc2zbg3cP1tJB6+wQwedRxJbtuZibF/XC0OHDSBYYWOA2BIpalbpK4W8PzQxx7R
mQD+MbSYcNXsQ+o6ChBTJBvnuUCQmQrsw5WF77cUK4s2cg2k9W400/i/3ZyLn3L1mSOQOaq1kDz4
p+gmzmns2njlxHsK9bmuNz9eNb4X4o7CLBtZQqNY8PjfPLxNwoujwLk4LrMX5I0AjTLjxfk1PkLG
wQ/AYCY7k/0HKBR4cG8WYFjMBESPWSnTovBAPvmpb5P6odLoSBbcPeBZuPOM4vp9NOdLCJG/7SdF
hoaSxo0Bi9KD6IokRy6/OtduZFgNloNcSpp+1euKDeRmFBFaAzMncCVCutfE6zqVFTVnGjWmijs9
1RAXp0v20Yl0jk6pfmE0g99DJraM0eyqNWbLNRHaCJr9bnjziGdKAL6yC2DHU7wdoZ/AYr9Jg1qo
wxBBUQwyTUC2JEB1RZdZWRhEPFhJzVS4FtDI8kYSE0POGfPMJhtH4NCh5IZ+a9E/1vU64nH6Sh1B
hI7AnPjLvpdW1sEHyubgjd/FOig7MSrhRy/IioocvMWb0MlVJ2sUXl5A4mcvpYDtwbQW+yQSvLor
84JzfVC1XWTcmbCTrA+Y2GjdH0JGrGK52ZuBHMnc1jUrLVRkfELJmtW3o4JJSAYdZy/eE2tpvB9O
3ZNAR/3fnLbw49MF+XnrcGQpznbxfk/mcAP8J9kxpVr6R/EBqykvuAQeX5P8C59rfrtFUwQzqV0C
wZkCbr17e22ed/rYXCSHwUz9OlRqhQDs7Qpb/Z1hkgvFq5boBqj0jAMobHVldMkkcpBtoL5OVg8B
oqLbQOyec2GPcXUSGTCPkzAKeD7RP3/TTMeYjFaSEMxHdPlCnhsYrWpoQtfLM9mSJBCBXgQjJVmz
xGm6h+uff6J8vUSPE5HDge61Nf+S8k9awS3PFhBUxo1T2uBS34t82w/0BsFNZ9sUmoXxPekmXTta
uSNxcKgeDrS/q9UcJIRw8D6CQxglsYcDUNEqNEk1sfTPrT7bjwb88hY780OrE2D/Nth820qOEsPi
ODrCvIxoWnAiE76n0SCCsRZkO1KUmzCKqWuogveXlOUhJygZoJDW2s33IdbEMXSXeV7hPtx4IeTt
xQgnu5PDgM7bKJT15z82sLvUVfYu4RrOX6nQKtjL6WRumaOgrjvX0u/hWNwizVqUbxbsF67xmj5x
R++dAnMDQ/QUu7nEsQEdW99vehnlYVMqU4XeUjB6gCSkagGT5JDrcjVL6Y3hOG3eoRpFOjzp1CwA
T9u5LHVRkB86gQ7vgnsLkzo8+rVDx9z2ozh8wUicZ5sJb7Dp5vE0ivk6HRpY89j7cPU0IK1Rj/zq
xj47kWwcu634X2B7Vfn9xSWe+Y4ge7HD/F3Oo7CIf9X51ASEpbcrDJNMnqy3NuRcrR+C/32cq7Ot
53jBRMEQWvaqTubhpK2nQfWNa+PkoHkEgB9uf+yFcMa7m1A+ZdIZXYu7jCFgn0dDPJnrrfGWYnmb
oscSJFOoW4CMd/ICv+KRpCCtYluB1F2d8VMMzA6UGraRdGTUohRsCodEQZtsuzKCs6Gy+7vlQNWh
f2W/DmB6cboVyEW4vW6DFZ4FgbR7poTa6fpIWAGMoAMYvTZrWDkxgCNzpWR5wgTkn3tenwSr8Zey
me9ldAXPsBTgzFHXOy6Fu2EaJhr3ZNvf9EV9eRHdE1H3mDcEC1Db0DIGcnHGJkEq+VOFqrPZUQZo
pmJTq/mRtywmRgGbSlZpiZLYS4RPZCeFrGFyORwYQxNnWqOfy5WnMVGgW4Z1FA7nHdRQU0NppBFn
XiZhoOyCFp19efmwhKaK+FAgHyAWuiarM2CXiBaQdi7dw8XAnMP9jriLJ6SxkUNdLaeWNAMq04qs
mcCELt7akBJMRP15BagcNvtTTNLVHbfyP6cfTqIh+3P4mzYFWRSnGlUvMRCjJq+4qPjgsVUOYr3E
q7uyWYqLtV3zOXztKsYkDJ3qFY/ZHmpwpvXQNsqL1t1Wv517n1qZRywaey8Oq+o5ZWB0hawU9fjB
leNk5k9SkhYg1pRh2F6nbDn0WMSFN6kNvZ21e4Ns/c4oLs9mNZOmcwXKYm8NvBupEfwrcfqTEQii
G8khXJJXLWzJYd8TPUa2eEitgCLdZ5QhP8+do/VLR3pTHkSbo54isiaS0rVZd8IlwFd9Ww7WwpW8
8B+qi4VJYWEH6Vn8GECXpQlZWzGAxKFU08L66X5KuPvasY2hv/k020GeU/DWnhvFGMOyEgVajuGF
HQMPaRfXX1PzTgFi/d3xb+t7TBU2Caz1MaPPu89aoF53yWy0wm1NGPn316zN/SSFyf4FNmSfiBnS
1ita0FNSmKUhi6ksMPN7whxn7u0yNSqHQpN1DW5Cl3eB4emUU04XxvnMKRMkZ5hbEt9GEfBDJhg/
AsHdDzvY3NpUThLQymwafN953sQwBw2sDp8TdgBw+r7Ub99KqeIe+CK3Ea1BjWdjyVe51B+/Z1aH
HuBl+9PyIlTw4HbHa6n8XOov0yvebQuArYmcFoLe8t1XPlognN5lvH8jxQFR2FqgrPRU/yuf6vwC
MR2iv761U71XKG+V91vw9AKw5A+zgrfC4qINFmuK81HlYN7E5/PYfkFQWp3CqL/cyeYDXMSry1TC
6NOYj0GWLmZZjSfgUgO9hYezrTjkbaxJ+G+DmfeN3SIm+LL+bevu9n9UfIyR9bV+Vh6yyEdG4iZw
J1SVS2TkcpjUfYXaWy0D06rOTbph8annkMdQwkdnyGOwfF7MkJ9h/W3LGz+yUF1kGEsToLcVMkD5
LvHxXZhF9Th5MmyPgA4LNiaZmSAvQV2f5A6oYn7AP0dCxlmhKM5BvIInpX1DyzNBVt9uwHUjaT75
Kdy4xTyPU5cNohGfhTJKTMMr/f6GtcPRRP8itNRWSM9TuoGJ5XsoG4P5uzER/uNhL8Iy3GbPaj6H
qBrFBR187Bnr7F2JxMZn9N3+pYIBA6qLej0nv9xctj7ke+YtKx7MflCC2i0gfuKwDDe8KQUMskWT
weKd0e6jjNm69hwHachrLlP6DsErgoTs53xS4dtYrdr/pcYx9Bp2z7ehNeVqz1937Y03oZGq5sjk
qyMkKkB01iBSyaSk8oHWT7QlL46a4fD2cicok5cWKsuSYlQ0UV/Pde98ySAz6h4uOB5yPjRr4e0l
uxxQW6BdK7Do+UdtRbDWKawssOMQoCJk/4rysVl5WS+I71UEYEoiyUEofE1X0sZxefOUuG8Mp0Vk
yWSB1GqQTVTtc7bwmbrMv4xVbGoF8jrBI+oub+qUbCntFOXJFLtlJXNEvsCmTCcMKWp1jh6mcX0H
zbzkBvpvJydsddKXYtAEE35BO7chA5r14xxiDhiYNuVsotfIJCsKh926AnPOuk90rYzY3ic34Oa9
6aDsL1aTQg2DFLJhDx7Hw0yBSEk6D1zZOaF9BozKl20Z0A8BbCbloQlrSMmGtqzrx8SRms9BjHmV
WAaN+KW5IS276b4ib5zYMD3lB4sqMDnqfAuBmHY9wCK/OwqQHavUuJS1t+aROOOfkCDqTrOqshzf
/gkay15yvPDKA1Fx+DdLtanO1Qzs3ALia8UAIyoOKl9Vqmw44g/bIUWABqDntUM7lFpxOdtkTOFj
xls1B656tL6jV6S2wGuCsEtSzzZTY8elcYJS5qaraOp3YAC6+JXs9AQawM4vsxerkq5l73fjzYZV
6JxUM5MQuR4RnIb2Lm+8WzyUM+cU4nBsCkVHr/5/DctlhkCdmoTnyzTfN6UPO9y5dI/Md6T2yf3g
FQ930l0I9hA2GZLBjOJXVFH4ZQ9TBNrehJV0mbT/F+tFxCe9VnuxeI0KlMBNy3NEEXilkrWdj2l5
NvAg5W6ekns4Tbm6jtEPOM4S27St85Qs/FyU5k5Qej17AeBGBleQRYCcT7gJOVH+dUjbbpG9jD5y
DPSUIrQlR8ZKwUBjUbMwauZtXWA409aeZbjwji25C8LSw7raq+efLhtYenmcK+s5s6HmC0+jIQM8
igSYkQtbLFdI5kOlceQif6GXdTLsAgfMpG3TnGKjcnN/BKX+MMq/Plk6aUiZXHziAXd8CS1gcfIb
8RrnDN8M+RO4EQfYDnnAM1FKLH1ABa9BJw1FrXmkY52JnT/2t+0VBaxhL43Azch1r7RmqSl9hEws
i7DN2ObNJ5QL8TNWKncZI+kzTCxusJsO/0uonLYPOpRPNSpbd38a15E0Oc4d7mGfCvaHD/Ei7AO4
YJc9JVbocjDtBR6DsfaHyNfsD8YakqGZlbAkgIsuFZ4QCCKw8LIGhn8Ui0jnwIzNsk5E1G+K/8e5
CGcCKGoDFnfLHH42vCpktkEI6gR2FKpXVtOAS59h4c4MxARfpSKc6ZzhO4DDT8d/IvWJgpSQ8PsT
la+P1llDKTZqIEQ/p68l8qVivviGgxy7FrTUDbP4J7WtYU132p2WGiORi2CAh8qce+sGLTkiU6ki
udvFu8BZPmS1E/vjWugfsmuDdcooGlZTrg/j9XkDzD1oJ+94Wjp1WeWMjbURlM2Ki2/aIfZmxACB
JWh/Lsyi4yWbA3+hkigyD4vIxQyAkXo4Kcqk+X3TEgqdA18L6SW5kDXtTdgfXoptlZKWZPV5pD7T
+L+aPgq0h1Q4/LoIcErrKBi9Z099aCODo2xNzGfEEVWCkTl1cWVfVcyBTnMlU2CrOTcFsN4x4V2b
31TZUQkqRCzQpqR+oJvh3YIiSuEyo0+r/u8qwrIPO2BM2YM9kJixqT5f7Z0OIMZQIMWGD5w4vgsK
qQTqF66FGFYbNQgrVf4a8rPauLcXW3Mt67Rq4PC+zgWbVzfulKDLr/85KSyIWBzOzgtk1/b8Q792
o73bRZlaEIeAGbo3eNeHCPO4OMe5nraj3oLJe0u50jkIPh2nkJmzDg6ze/mBsl03ztEgVzvTo01Z
BA7XQXzIO85LyF+cPu0MBGl78gsMP23P2Fs/5iwKn1XFTyytJRFuTjbDwvSS6NVcy5I4w0Lxsgn6
hOb3JC58JSGlNJfboS37XERphlH2jnOE0QnhTS0jleeu5w1PY15Oh9b09V2zSA/rB8mpsTymHe70
dAA0gScZBFc6CqfI0y9kcTomVAvfHaYSy+54zwUgm2vYnyftTTz7wyP3ayMoFIBxgV9VCihhQz45
W6jTUyTfk78kLWV9wNnyDdOCFWAJM0IEagVikqBQA5ZkH4ty4BUXA7s+4tn7XqqgnD1hg2PdKIqg
ouY9b/MQbdt+p2eflEiJW1crqasb92FFhuLbCMcBlwc5wtN/H3TAkbHSfgdsJpqyDuEPB0zxrQ7g
YFvP2+fL48caXbk9gMaxwF7Q4fBqcukYSMZcH7MOTJyBnyNvBZGW/M77u94VvYDHGdAABX41JecK
D7SS6upbhpJDKwyXsoIwIdZbRycWi9A40J5Ax4diewo3keCT/fi/Rh9P7nN2O4YBvq8cZl4QlQ0/
0clzVVlX100z42PuSuBPdcV0djgo9cPgemootALCgxM2uDjT2VXXE8TdS5rDTbTiCU/3JBMp9kFh
98N89ErxGiGcDwH3POo95aZfhLMkBQsKdGpnfuerhs+OV1bgetmWsqyqJp7dXvrE9XhP0hIsEBst
nzfPqMJPie0qoYNkZ0TSRZ3MO7xd9GDZ1ZeAIX9jj0VZkBfCFSSbsC65OMhYXHviLhEEA3px+xWG
REXfL2QbCpCpjKYhCg58y0scG7Yewc+cDyxWVmdR1IamzQb/KzzG9vnFrIXn5W8NqRood2ITzoI0
wT+z7/Ra9Gxnlhci+4NdJC4BrCyiqYvFl+jg95JzuOk181zVJlI+srt53Gjnjh31bB+LliUyUboU
29TMJhRLvk/AI4BigWzlVj2sXFMXYLJ13sigo77AzlTqCkloo1PnDBXsQ5w7PwsFiUWpoU+DU0X0
m6GJRIa31cg2BG0Q/M7VTykHVOA5uw4HzBfqnTMYV1emKbH/haI13E1jGWpy96AeGSfn/KIJZQ/w
zAQf4zqIEa3641AgLB2gPho53Pl4q61BpYlvFvh6DD/8i/XSJYAbmY5thFe2uKFCO2312GMfMut6
AyJ6nrGaQf4DFM+ubZrZJTgh1qJKj31VYRfpqnsf7AaT1AXVhWNP/kauDgBjyQwyOA4qIsI+qWlM
6mHS+gggdZcVI1wRNPhI0C7xEKWk3H3E48bZ106iR/ELWOuJf9K1Ji6BSRSDfWXC5vF41FvYgcHa
AVIPGVH6dGAD7LnqFf4F69uIMmo2lz3sw2THdallH/ozWdLU1djZXlWbKi7eI1zJpx+A2ptRm8kC
QXoVj9gOAwFvhC0L7Bmxt+CRenNQIoSqsT/AEMIegMifQJTQ5cqzBNI378aP+IOboW5oQtzqIhM3
2IMKCVL3uCkZTRWf6stR2/N/bBWwGiWofJzqPhp00D4wqY19q3XtyyfIAsxfBM37LIh4SuRtXqAB
WABCkRDuc9IZejflP4cx9YNNvIEbnE4tldVf0QYYqbNuQa9voBPrM65saEPnAD0fN9rCFroBJ3I/
FqbR+B7/bm8olfeVJyAUbRwYobLuTRmkIGfyWjMoJaXDu44fPUXORS3Wupixthw9rOr5/9nOY48t
wrCHIse6tnInWzh8lCFQv/ohMB7kQPurhISPNZ1XDiSajh+T0aop023UoLll1oJnr/RpqoKLpH99
LDlQ2QtKt4RjdtEs7kH1amV3Lp9pWDhsu1PxjVm+K+/qToYkGWMJHx0B7vOxlcOyZ2QXhrt1u5za
KVaVp2pso8hGLrUE7kpaOmp+vm6dCGz2daE7yxJUBClH4owtrvUwoAhL/mnS8Z/q351pb3byzuF1
iakL9St2P6JwVQO3LzPfrpMN5YIsc3UeJ3eIXVqz86qMsMMCpiJiSKAw+3c48qxlartFqQn8MHx9
9TbH+2b04KeViDL7HpDkRmr7HtSc0iNhNNDW443yfls06abkumsFI2CmPgpH8bwE5LSoVmsC4ZT6
vluLZaP1rXIdzIHhLZ6K9XRn0yQBCj/wKedaCww6t9gA8CgLVQwTPPq8gogP+OsqrxViwShQMn26
ZjblZKIk+j9IiIyDAZhifaTj2hXiAm7YIW1pOWrSLrF/MDpkm+u2KJu8l/h7vrYKpGbPIU+kzKrV
0Tsu1s/bKMbxbaVh6H0ZVHVaxf6hhjAX7MWoCSW7W2miVeBGIWGPN9bdEBqhX3ZZBDXqBU5qSSb9
KlewY/UFmhfSj8xtcUPP2zgWnoglrL3zQktmJlX+P1wDAIqvSnwUf6FYqXo0xhSk8TFmgJHeqhtQ
tM11Kb4JIEa3cFzOnMIbXenRrKr86ON3arZBJIul7f1wG49gbCEE+r4qtQMG33dJN4AW5Ijv9hfJ
trN4pEhT1UsdWyT1KDsEaR8izbcq4TLcNfEQ1B7TBLOqlttGPJsZC4zO1u1dWnV2+jbVkfUiBbHM
UDHX/O3UYjl0QAi0QN3rOUay2D3ZnArhmR1da3NxBavGzt7G9WdhhDxN1CER4VynuyWkY9Vv1c0u
LsLgmfWGdE6vgdhuQG3NT4+wylf4gAxvHTth4JwxLsmgPcDVXqDdlBKQCeMFBzQUn8ZHYd61rkiV
XhWK6FEShC52DWoExbJhe8hJtXl4oUfyuZ4rN4Eaw55fMBj2JX5Z5QOKgsNjsEjiaiiexTIf5Llq
+g1skGhiBp4vRaq5gReTv3xt6mHPmjf1NeWX/eTJAjP8IPeks3WoSoJtm125PN2p/W4pEGO2+jsd
qzDoLa3wOikb82pMDNrF1ZMtX/rv6iSGU9LIIipXjVsoKdHSfUK1g13X1QRSBbQPpn48vV6KVDRr
QC07T4Bcb5HrUik58JRLAKuEgcz+Mtfo4essV7y+wlr1ubNTmYgmoO24wXjjDlP/c0zTZGT9BDdh
cImaak+yjPlb1eJK0VREkykuYfpmeW7mPwvKFYK4HKM5FDw0Pvwkdm451Zxc/lnbR01w3TCEX56q
3WRld3gNe99cWGAuHO34F311bWNodyiWcM1no82W2b0N41QJqf3F0fMKqfdZodJhakqBhhVXcBeS
/m7zTE37NxenZGTlLTSSxj8GcAdEuMvSfcMd90hM3pVWRftBo267I8qRgN209lbk49JjkPa+qA9w
4LuHuk52U3nfbSGBVVcwhLKRCQMXI3vxcJ2CYgcF5J7tXLflFs+Ftz9o0L7w9LCUgC+qfWkUCLYj
gf+kWeLb5oN3+Sspj9suemz9Dwp3QRlXQXIeQBiVPO0jp8qnACe904NggLNuJnSGTOUdMes0M4ti
fU9FbwjBqk91GJhVCSgeFo0xT4pUKa6YIQxOrtkPw9ugxkxqpigJucqSPSW0NZ4wL54MVs6jzmMu
N6dABwK8zywlZ4SWe4pZLR6whYOTWjlsD/XzXMXfw1yqKSaEZRphvR9YdrbXuVwWEfVyqGhAUyJ8
qw/3DgZ8EfByXW9EMQl44Smq3mQw6SAzKKTaj4eK3t1eLz8fF0HI6Jlkd/7828EyJfS2LINaktdw
c1yezcluiyQsGdFv8w2C1uE3gBP7SZGFlsioSsrOx9Wk3mJPrjnAh9YIapxbRqT6QEpvHqcj/klq
x0l3Z5Du3ozo4J1uAsM5L/dTbMULRZJAtagNjWtte2wwGTPnVTz5lGBbbl48hnql2MYRRrTzNBIu
TtPL/8PvKViIoygy2swUH6yDiC2sgjhBcxN4EwXoqT2XvjnbYJ6xn9FdbnAmVMqNrHtEgVjYWvtx
v6pdiXdCNeMGSCuuqdkFtK83lg1GGb47kpH5IF4MfbtR46I9OZN17Y7sGV8E+56A0GdTId758RYh
bVbO2S52OMj/D1Fv1Icwf91FqKdTAZv2SS8u/yH1kbSxLeGQZWjAyxnHdRDYAGDARmfLTZ1Lrp7j
NOmUh/Ruy5CDRuvhtsDVPIvc0ZmAqV28+M9ZoTde5fSLZBn4VG3D9+/PCJQq8rjIllEiLcYxeQR5
sJtMsGsKmyO+Y/18FzUQ2XVwV9vUkSVnZmGlH4v+CLQlfBUilPBWEPsO/VmQ36LBGbdAFIFTLUVj
T0n3BHQ1WUR50c/s1wHn6Tz3rHbi33uGqL6BNcANLQyGvAFgRdiYd/grhXmTPOffD6ot/RiCGm3g
LcMTNB2O6f79AZb0Su1PHWKZCKBtvSQJa1sKA3dWNjQdUpnsyjgfAA3awh6UlwzARSdOUZfnHz/s
CyFm1XCumtD/+mzt2sT8BQ1aN5v3CUgfkZocyui4/8d4zcqcaeRbJ1gBz3sKlG7JzIWgIXcj3Cur
J9AIDnd1OPg0iu1b5rcmjmdXt6rQ95KgfpllL3TaZ56G++IfCwdsvqpkcQfNLSRjG2+yDhuSb8k1
mbPZ8KBdzI0qGVby2T2aHIZ2XU1jRTwgrxw4p30qE6kjbgCR78Vtk87VI4mj/gLGc4VuPg8ylsUL
9f1A2kjKgt86e3S0FpIG6uGRq8VJ+sZZVprWB89P5T/w2cBF1Oqt1SKVZ/NhTFhfvEav2EUCENKa
bhP6AM+zFFEtoQuY3PRMfbK2JAphaae0/1b0PqspaWTvsggCQZ8hBVtwqGbGItCGO/5hIv1xBTKW
fvjJJwIlScEQf+GdIeH39RYXgU9Dsn45HM/3H9NRa3MXzYWsUszxDGqTpxJJHnX44Kja0vaLXh6L
rj0u++yZLNJEVpXmGYiRR2x55lAKQjALC6J3zdJejZ+w7Te9AO21OhaoMWZ7UIKlF6JF/TlXk+b8
tdsAwCbagJp/b1HU1cbUNT37DVgBMtJ0U/aL8Gu43vbxaP9pOpUKZAPFg2Av0jtxqYwrxv90E6QF
DytYyFLB+r++5Uee33WN7tF3TCjvs+oLKYCmyY9bQKNnK4QErNyhcE2tm7gXMTpn2eUar7vvn+HU
URMxIypPiREKimNpQ6dcd1rp5TskX6gc5fcS4kTwaauFSf/mRQfLO2iY38tx0QeQjZONKNXqFjAg
qhqWFQs0BYJo/M5mZKJo0zFzkqpy+7ygB5SQW3RY/ZpFVAJbl7SNtH1eSeCff/M7na971TWzvgZC
F4X6kuXD8iqbwHkEnhGhtOLaqluFgGtQWDA1efUyhOUIoUu7tiwWEJsJy174rzUTWfeZOev8obMy
qlXXyH1zf49KhLOPTx4AmWeJRroajRa6hsw528zicZa5w43p9eV1rXT+WiKMG9UaxH+AIXmxTjxM
NRiCsCUsMXXGrzw8X8+VgkRBMKY+9FBYxfJihXcgxfWT8cwEzrokBGSlWXOC6EEXp4pEPr+dU7uz
tOhn3veeyb0K8IhaWYVWMou1gNLQEHV06ovCidjYNOGojp+RL1xgoLw/LTxzKkDH1bJlmdBnQHtI
HPr+ETLLThbqO4TwZm4YHkXf1yKc+DCpnDDkG8gFl9T0BFH1NCSXSoYu6yruxFwK30DVtdiVE7RH
dt+sHNn6YEYOsi6YastSUxXWChUyEfVzU9DG8wB8jDxShugJbCxI3zsNrTCDAtQcSQd5hKxYDwpV
HqRI8yT9/CxU8jdG2MYLSUoRDHlWiV+nDHGRhO8eVix31fntFZfmZqqaImrf5ff+ss6icFvpzCVG
Se2hD4rF5hL2QXZTVjh9CMXTtr7dzr6CKYf1oc/xvhNDYSW0S/9QhflNy90MCyUlGSjFpaiDvd4j
mmtrSCQkQbvzOH98J1lyk6FFtBa4Ik6vSDzUciuNY+5KbTbCOo2A7MY7C6NmeUxIPBtWr22it4SR
V+zuiA/bbqjxb9UJe8i2W0DVOk8d6rLxTsaKLnAZ5vPfp1R+cmAzbE/00QeS6lOfSCb69Ly2iLRd
CnShNnnapYWbt/8wtiNLWD0mQqjEO2aauWloCg6ix34yP2fo0xPuaY4vHuPP+Bk/l9Wyu7xGEcdP
ixqT7i2gyLZTqV1/BZcd0an3540f3cTznPQDLOwACxt6y17K2cGoMQLRh93ABhzB2uRHX5ZNSEIO
ZwEqyJ3u38MGLZRzFLrXPqJm1h7mBiZ5z3+UxZI6E7gDhnrLmJdpdi0K+WP/UJUYiR8DJ0lnGpPD
jsBdr8fdc83Oc4MoIlEcvTHc9nCvnThaYJ4XywZTKcqXxbeEzQkT7riSGftnta7CoB+oWzPOsmbF
eMfLTEvtzHk5h7I6y7h6FxdcnICTGW+h5Clu+mL8yPTzrBgxXfAWz0jgMQvU45ZPFP9w78bXSXZP
aw64myd8M718invHFpxa5y09rZEPrfy5Wt3VmEQ5lxDFT1DuAQu3CzhArhsO7z/0e259XDK2HMOt
vqCxnmNfpJlr46ehjNiA5fNVvmVD5u6d0rvwQcRKw8sTAYMEapQh+FQnutokuIyC4JpE16h4xiqy
6NIEuthQ4tOkao9jx39OiL22Dx37LJOqVn8t9MKzAX1qPmJX2gIvurNdJ5IO2h+A961BuO2KmYHk
4C62JyyBjhFohEClXEtr5j5HAr72gxfQCdc09W3M1u8enlB4pSWJU7ZYc9pmI1oydT7ZQy7nAVo5
DOg1AOF8Znw+yVrHFWwSFqFkn5+deUlLqzPmzVBPwOUIqvPPSayq+bphRUdxyFT01I2uBNW/DRf1
W6ksixKcGJ7M1/Z3iqAAnkxATCwd0CiRROidsr/Q0mvvSeNQxEKc1IZEqmRaPS9uLQHxJOKTV4WB
MRapvWJBf1GFJ6hQdnkcOt7LiwrV+FpWflFWT9ygmQeuy3AGVb0jYAyMIX2GmVb0ET6OXXHESpow
mxAzRgSLt4dKaD8L8rVwXYs01SVgfZYU+689rDjZqvZjGICtnemTeXYCHRg18o2/WIn5tpYv6bQ5
pyYcxGIqoQwEuWkJpcBvaMyggs9uwIHPt82JGtVht5Q1MG68b4531P19var/KkkCpkXYQJdexpPb
KhBkvAmFqSTfssKoqKC7oVT6atAbj2wMKRLtHk3vvPxmbqIcRrZmIDnMuM7ayQDxdHmOR4zNQLNZ
kK5Iwnse+FBqeMBqi5+Jci+B0mwgOKchw/i9O+UBtquMKAf9pQsgJMhAhrgXZFFPUtJEQPjKKk/l
A1Lo7Bgb8S7ZhGASqycdykDsS2c0Ie1Aq9mZdxMInVEKlFaXXxLTkm3/ndnWNm2qhPR6IQpRE7WO
URJOstlhKIe0H6t7c1pAPVl+HNs2Xyle5vBrWwSBNZRtwlffUAbE1slG5feo4jMJ88cshqPh5Xwq
TSofZ6abBi//28dedQxTm49opxZdZYbIea9bEU2goR40Y4PdjgtEjUgZHRjeKNDIn7/iU+KlqTRc
7tJyoTa2d0Dn/t7aTZnMt3q5j0mVeb/1tmWGHvbYUqkC4fV2NW7YnNg3CtofbJbuzixjUvjT3zuq
sAemu+A/Wxa02mfTF4gkWyK5V/VrfuinC7Z4A4L1C6NdgpIbRStaTEICNlf+6HnH0jKFzL7kYEOP
MW+vK9IYrRUlhjGBGWz3JTVMoNiJamYI8MBQMXJ+AVh2eMlZB3to9hfEKVRaTtr1gO/GnuLUm1KL
RPV2/toFEqMreCPU6Nhpnm9BNPSh6UygFsLVqR8m1qPDTigUnRxKYP1VgcDcf5uAYDb5BTXTF6sP
eXx3x0pJERXm9hqpLZTklyw7LW5nNCW2R/pH8/1HUmVs5qdXDbBEEsyYdRqssX0NtUgh3U5dhY+R
Jvibe+H2/rGD1NhLtVSuIwvAxWyZs7X3tmy0KoAz8a+IpdzJfOOWZvA1RgHqA0c5CgEVk1NL5hyg
zAq7G6q6u1Z2fRP+vm10DtXMXN7qI2CXf3nKKaflFEU7qky+0bkdoYo4YNBhOkuAaZw+YKSw1qqS
IFk+jiX2c1asWKyC3RqMXipsoZwZiYUAabICPy7CkIe5uwpBA/w3GdhxyPUCoST4qJ8nQl3Mgids
dR8GXS3EBuHmzYBeDCZ8oHVoBvnjgpQyqvWGCs+5jRLGPNa/A3lCA+xNsJ+KmysQuvfqyly7vmLv
OpLhqgbCdBEgr5vStiRo5oBdI5UvTG9RLmaBhAvB8ddusgKEp/lqNI8UmRhznoVoNyS1K7HApM4h
LESlhrmJ9O7o5HeXi3DHwotM4zxSsLFsybY47b2C8mSpdvaq8qYDAgb6uLydY/4nbVfQfrdiDM6p
aFI92Ibt9LsJg+QykNUydcswCWFDhb0gXSGaFVWF9hlSH+zgad0OYCjhCIvIo/WrUyJI9z0GqE4q
TwhUtikRbRbXqReMt1uOofP9T6h4NJ7dxeB7p+K8iTDdjOD4Cs1cCJw/DTbxHaMjH3i0ula3ntTv
6gbwMTU/74sc15F1Sx/B7G2de1XpXOPhZw+lI1z/WyzQI0QXDKWyKSEtRsqGlJXt4+1KuzcFCNff
3ve5+phtMsVaPpBTns+ihMQJS1jo7LdnvugT6JfnrsbD1QasRAembsYtGvMRsf/0v5KcKkXU/q+0
lKCbT4iMJWm5jo/6d1ZUcfRcKiGGXsd54DZhOy3VEGqmYmXd9B0axePu3Ryg3J+U6MQlIqLiyyRl
+HxJtWLTDrOG2V2l5OA8BAJQidf0sRK/qt6mLrZAgD6lJNGgwCIw3+k6eHaHS02gVPOGcMFWPQr1
wfkN8fUfRHxBoDhMhI8V69NURqYG/ZH0sjaYMarOg5IURbSb7JvH/WHvkL5EhyE40b1k3aQmgy/x
7OXAr4kiJDgbt/cu5UTzQ04tmOsiynegTShZrp3x5JeU1/efvzDmGKEv/PFeNyBN4sIGwY/6KGCN
UKECkU/2MNUNJ/D74gQhzCZ7npbEQWVM9tkw8v3Wjck3L3WmIaGY8O4H1do+4vIwoGVjV+T1cE7S
LbF72WdCKmTPtoMKRlWReARJKcq/F4rqqtaU3LNJjrOU2XOy8ALtqY4wVWI01f7NDFuCvFJLLXCX
pCP8NBw2NMErl2XrSWXCpdIcubUp0/1wWXhqdeV2U0lqDcjlcCrXxq1i7WoZ7WmV6vckEB/5nRdg
PZZ1KQJUYiR9FQ7XlGN1vJ3pwaVghTQAmqw47pvYv+Lz+otUIOPr7iq4uCnImS73PhimMrJBa5q+
e4v3y6d+br4ra4PBh46GD2y0qf61/i83u5yqnQqtxfIheyP3r8TckbJYkVyVAZWzhFF0oFTPxusT
S+jHu1LgsnuisB+BQSDRWzG9wISPLJ75ktz97ZrjcBerkZZGJ2xMdQdRovwIQSIIhTfN7cULz25T
12kDes6HDyRFXSHVQLmdY4utVFj1Fh5n/tKNgFq+Lk7n+n59yjQPpQHN3UGbN/kNcOcc35S5zvMj
payA4Ict5LDZOA8CCDdbqCrCVxjXNJMv1Vz5R/dk6wgSTDTjDQLLWs8m0k95sEkVVpUljsW097Uq
9eXT7wI0bweTyA5rE9+mjJMaGl4RDhsX47QbhxsyZ3wWSdOA/Mnd8oVD3qvnmtQpz3SdTZpYdhqa
avVBe/79hiImzIfRDYgNyujBhadWk1zZ578tFD4wGJDJDTHyjW7fkye+h+lG0MXHohMO+0+EKoW2
FuGUGIJ36AC3eyN4AlW/5PO6dMwrK6Wwfban/13Lag8QIXMA15pzRs2IGgM5SM0daixV3OEfu+7F
u3kQa5JxNj7IJBgiwjBCXK22+Tn00LU/vSBZvCoIfCuwVtKBhjyMGHAiDAjXmO5BGPETSuHd4h+m
NLpT3Vriwj+HbNOgWGw0liwkbhci0N0HMHHxXNKDeG/SfKsjvxPIR27h3qBl66f4hBMjD2N5fxNJ
AH6AoI6iw1zwdkCViwuDvAjFNeOrSnI1SQlwQ+ohZe8vRYfcaYdothetqDRClVyfzsp+TvLl9VvM
sxwOXjXUM0d7Cp+6/xZ8CIyPDXEJ/EnEaKjxj16mdFeLTkIyE7HEPnhtTRgZxnLIJ+9ACEi1uiDx
+TxuXa6lcsekPuab/ORhehmKtJ1MO9ifhZOvQwGD8RGJlMXT3au20MV9tQRtY/vvILfCExLr7/26
9xwtvzLIoL/bS5FKIc88gPCuw10CVCXeT14OapsqS6Ar5HpmCx/XZgcYBCmYxZAkuteIOS6y3jkQ
geHGtXLdiG4XdqG5QsM73glBtsggoSEE/S2v6r8CEWBu8v5xi1sZsAxFUqfGprEEMIH6PnoiGnxr
fPbOpk8WCaOmFnHElHDONnHAETbLbrDSRUkJ0kzZIAA/NmStgV1SAiGbCB5SxSFR+0NSx9K2XSXG
qY2Q6KLLGqczWWTH857FHJSphRvZWR/Wv6H2FvL6Lhc+1W1yXwDr/K0cYQTc0ZMWrr8Uiwwt6BGr
1h+zchn6onH9KpiX2UIO17Zu7FlUqni1OgP7aTwBoLysIXcg3yFuPDfzK0Z3R4RPzN6oT+UZwuJZ
O//18Zp/lA5jMPuhrsa3ZKgnB/RqQNbu4bmMlVuzCTwLbzLW/EW3P0bfK1K8dP8m09FaRpXC6tgV
yD5RCnzETXkkJt9Y2JaGfOlSwJ9dn/UgJUMtMyyIVJmfezFvDwsfG/VBhEMutednNuUI2NUScmnL
YEqllukiozvr1Rp7/v8cTyoH+3YfendflPavlQT1vGvkT2bpLyxhPj9BzXl8GdCoAqJLBSIYhnA2
/q5hZ0uAnXrcfrP0/8fvakLK1dOYR7GHHiOMvfYIYucnbgG+o8accZjr8d5MJnf9fiHVZ7DTeSs7
+i9vHbR+YkFBgIvFxYXDg+OPr23vBziwirFMnIWfYHZYTDw7KhautDlCX3infYCRt6XUZJ+fTcvo
wrZGAgnPiyX2Ism00mTkh4+PLSvrTLpaF9DGbxpaRxnsklEOToABW9xvTYFDxRRaMrq3QIR/e/DP
PCSD1b79CdJuSQLUnep6iTfQ+tc2bssYtrfklfW31nLJKGScFNJWC1XChOuflkfnc4pjXefGP+NR
xLWB3S7OAdZ4yDsAfwYY7BxoritAWBTz4MDZiZSJsQqstRh4vgtDibj2B15zdBeSIdAoeJw+rdPW
DCN7vWdChCFk/8VP0EByplizDuwYVsOW7TQJEF81FqBX739LLoZe06CDquwo5hV3HjdCKzxQuCID
DV6SB0YUt3mZ1xMgB+wdsQAbNMnPC8kO8I1q5U/bv0xFB0UHylJTDKQZq4gUrlG+CrG193QWOXgA
QlTtgjE8ZRvw60GGwlueRYssUbgduYRgnXJWRN6NyMibcNlvZ/IqTOoHACcdZrHPB6EBEZzBD0pA
kXFeWkz6xULkzSaVx9ewt2MMDgzYnVeLxbZR16H/8ZyNJ0mAVsO0HrBklWIxfGn7K34I3hBD8tHd
VnsW8kXzu40k5NVGWXIYWhNWDtNi3pLJC5vKfui3zTg1CXwxhDqbm5J/X9ahLRaf+aNyIxfwFJXY
mXkc3wzj1fde0//E9z7wKn8iJATNDZtdInXEx5hsAmHqT62yBBtT6k0+WfSNi64n/7JAAKfLJrxE
QryHVH1WLh5kuwKAKk3ZNhIE2/yi5umvYh61mBM9WI4lAG18vBPXCyIvY25K4GFXH8AYIsOzLxiW
jBmU5zs1tfqEL8ZZRPpd98Ls5vXWcWDiU33lt65Y/E+ZNCQYEVI/LdchZjSG2bBErr5JGVM3OpBS
pk5uo/ToCQdUZLsIbUPKDUlzsHNc+rDCgE0HdBb1eu9Twvb3HMW1aFGoJJS5KwfWnDUauW8zHj/b
4fUmRNXxWdZBmOHWgBJqMFqqDMbb605GirRsaSpz83P8PMVibx5OL103Vp6Oxo91pGsxp52MrH59
0g/gCU05bKD6B7DREwzC7VKc2z+5H1XCD/lgeBbIbpxb6UQvA2xzbnuwrjzdFRmUKn0AGYM7uCVM
lPy8k5uqI+TH6iruA8Ufu/GaEAtnnH9vY5pRfEucFfAi0kr/uIL3p/dr1vskrJ5TdOXyHZZAjgJk
Vghgs8Vf2dzmfRFU85ZZV5RPtgMcXlkLkixyYCoPR+EyRfSnWEv6boopg4Vq1LB7OcOlD2rUi7UW
2RP/2EfQaeb0BICbLbNXrv3+/jp4YT92D9ztxJnnQIBAOloruGCnJfcEVwmocTIj2eUlXRpyPXNd
gOpv+WZDR+HncQZ1jaRIHhTRZvQqTjNH+fB4gElSHAb9b6RZKhSD084ASsMumgZ2383zu3yMn1d3
au1arthuDwEISkYscuComwI4DZ8l+sDLQRfnEyYamioGKKGvSE9LFzStW011P5XSODGHZqaBSwyH
xK9ofSF57FgRJYxHHofSAY1fwXZh4zvJyrzaQJBI0j6F/XMOzNTPjahBGE/4z3NZs2oGaX5nTR2B
sHxEXZqi9GKzH4KLsvnFM/0qqTugWBM2xUwCvoh1TsrVsxsas+FmcuSTNjWYcA/E0bK2bMNIyxfR
T9PHWgaM9ZRX+Kz3a1BDApDfXk27S2iA2BnhkJJBOvlOVEiWspU6YcPQ6k7uzamrmAD8XkNB29zB
zIJgZgOgPBO0sMwWR4DuJ/5hMt85hNHjdig6npRe1V09xSPdgRfKIjkOp3WiuAX82YrV5FVgz6GJ
r5uI7AgZdapPVnVxRaS+9w9l3uFGUa8MM4eudVUcPJV9YOpp511NS7+MtHSsiu5H8/SuuQQlLXkS
+0End/xNslY1WjPklSpUFgsyfbxMpjHCZx2Sw/OvbPGTLxmWrJskzl5Tv1hGLh2+wTC4oGCwjSi6
NzgTkUcSRdCFivsuvge01XJswxvxe6KNaU/IgjGhtNjVXhQEZKq8k3pb+0UHIMZaJCUOdiy813H5
RjHTHvt3ZznvR3o2BLtvjTd7liIJqwxt7B5Cv4CeVBBmD34cuHZ4/W1Dyo3C56jUjB93snkspRLo
pjF/I8sIwRGu8b7jyNWLoPwlYsSnnYj5ELehHUadN7XtQQGW+b4G9ePWs7zA9U2hyLHGm7i3jzFw
RdFGufc6oZHG3Ifg7DL2kpecLvqKIJJh6KnE0UBNHvkRAwcU2AgT+rVS4rPEH9T6+NoWUG66Bh+7
D2wYWAd66lEuF3J12/a7yOL9POnyTPdoNRHgOewzbn+uD4tdRXfOgW37yxXBT1LOlP6aGntnTjBl
UVvBGLOYodHeyopcvSuia45bAYvZTVsQ79iMGVzVuLXjmw+bFuqmn8x4KD0blgLFoJxtkEzPhODZ
gob0gaClZHxfhE4E7FNRELREtAtQl6PloS84zkcKHxOdMxTUfb+QUaGNcKjb49R/iW1Z7bZiNX5n
266X28mLni2Zhmmynnbqx73gocZaNqlfVmzNy9MSV006hGwmts2YLYcbj3k5kKRyDXnNUujfJ1BX
JG4ZCtZBOca5fw6YaeUknCNbCylh8vRHf6TocVumIV9G+h7p8udZ9x03pqgpU+wmBVek/JSKUXxi
IlYvQfgaaExcn0FfROFVDIOWyyYYZzkyE+5GmoFrxykCNDHNenbCh1rrZakxQb+dDVK6i08nSlcJ
203cJdUShF62D8NJbBEjKllV4X19YOe9ry8p3WWbHwFUC+4eAD6EFJXxFwrCLB16EfgWU+yVPd2E
7LqiX9znTATHnjterMvYQ03+LDxCeXaeNUcLoY4px1nFG/hdy6bENYbBhYOiqMPEtaZGdfeGOLdW
ob7G8Me2SziNypvEDI5lXphD1Et/IddeHdPUQzsLNBtFb0d9MeSoA9znbjDUpPHx9WZEIrSXq7v3
uZYOf6U/edn3BAonVSZrruw/61YDL3S5nNedr7cDK6taa81FS9rFGkhQPh4ou7cIP6CkNX1wjjlb
xwLzwjoyI6NB/HOrZPu2jDgUQznRhhn8ptC46wniz0BiC6QNcJ0NBwrcVQK9FYRzGFuqlIbc9Qxv
uKJreTNewD1Plx/c7wwfXIhSYGTUwAqquqi/BU4jQrBrObV1u17yOb/kqmnN01XcBPlxnj7Tu6aT
0SgLAiFHdOpCVktrcv5oss9Cx1ssz86jke+sKU5z+/yOexZ5cPzkpdW07x9SIb7e1NEdqJrdfQrd
MxclkpnqeqzLXscSo70+NuBqqDPL4DNDk5PhJJ2CzVxcECRe3RouuDLxl50bKT/9+XDvX+wvaBMj
nqNZNfV3o2LmNCRLs2pocaxxiTLth2CnBXZWieXUk5l1ht3ttijVmLwzGrQoB4CUVLv/vWfwLlnS
8XsLMuUrez/akhRks6xyEIGShLnwm91OpimtIG5gjJbuH64MllmD9NjkzHPCp0CyipqsLPEQ9Afy
FKWroSs+NvKdZYeZ2Nx66g7hbapuewPvxiP2kZAYW3sK79RkdBtxfLEx+JzOR4LEsifwOTKfbfwu
0vQoMjRqMlIvlzm2CjKEfpfbCEhbJKdOx54b4wEO1JFVM2Td8jUjLekCqHT+RSzd8htEJi0e7xot
i73XxCDDiU5CNR3UI3OmyKWkrk9NpHmDBObpj53pBn/dhIHXOu3YLtTGWGJnsoUQS2ORIbnCcQbE
Vmc0iAJNq8rGZ47okHe2W5Wjqye3MC4D7/1sD+1jvHmv5B/efM8VObAOAExt5ZZrUZFniDP42nvr
+HfM/zWyYg69fq6VSDrmome8tmXY0Maih9oDoy4nWnxIt5/0X7h8JW075ANYnP3sqQ4HasTp7xkl
FBJCOaAP+gKayQRZ0uM8lXXn+gcuxY/8vF0gouDo0lrnDMiWqDbyDaI0k2YavFpknJMq/0zkGc2E
9Pf83flINunFyllOIYF5AmwYnpsrrp/qBJo+A65TZkoNliqQdm5ZyJbsSMCuVIKHi0ZTwTREsAMp
cqwseTYqpCBNRjAC9zvyEpdqrW4kWHvnz9x487J4NOhgIJFwoS28TFhBOj81r0LmVv8xqhyrBx8N
sSz0Gi2FNNswF57UxnA8wLSL3w/97iIM+4a+wu5Pq6t2xCJ+zsWbAA/Dya6PnuFgzQ7sTr38bSLX
OAGDvxWUbqUZCFBEbYH/++SbePDEUj2NHTYMd9TWU3icWy7K3LGi+QdZMUvTl5XFMYTpAkcSUyEq
X+tF3G5bCnrWtYQkJA+5cXICnLG+2yOyzXcJoKflRwwPH9PsPozUfdNyFd+pqq6kCN7Gw0EPxJ8Y
61+c1HeFiwTRV4PsJiTrN/jIEWPEwp9cZjA73dOJqTsck5v+m2cqKrvlWMa6e/HvH9vTMFBK5xV5
VMLNvMiJIvkzo/oI8yLinxi6NY8DRRWpjP/hW5A4Rq/fYw6HSwt/bvYhl+HyUWMwbHE7IBJC/2qH
34FYn6gokkI0bMA2OqyPwGFn5OYpG+wD46CX9cdnRiz/cpol1m0yIqQjUEqVZsBI7RzUuKpVYFD7
kF9y7OxZkjwiE6QZhLVCP5fCQAW+v1lH+/hWCUBQ+THrloJVVijqYy38YkKZt0sL0y4nBcRV12QJ
IZcNjpl3Wnuuzcl6JdpgapsU4cScQ+yjRtVyu11bn3jXdvu+On9IPCxFoeLkVvUh9S4LOC4qbhaz
WVYJSQfuzL45BhgW0PnjD/NjLyGE+KMARppI1LM2FEfXOPxWC5GhkRXopvqLcdTInR3aAnkUxp6A
eaV2O1bAEuRrWvia5JMv8YfqgYrbi5pMeUhbWhZu8TgXADfid+wwNLCc3u7P6m6Gmu+eeikZ0HDW
DFHTXA7awvgs6HlyBdRlkYvmlDMwiZQEjz8ABuX7wCL5pFU1ekabkU2XYBKxvlJqmmTI43XzvAs9
bfyBmTAeFiaDyQ1RMS0/FcmHJrRb4clwsPzAWJaQX17XUzlhS+iEbBp74d8YHqgcpiYRDbnU4p+9
gK76iJvqI9R02/HxYk+ClJf1Xtl7vM/NymLF5HNZfib7woDwVSfSwb0SYQen86+J8yTSzmK8CriO
KNtxQRjilEG27pp+QKE97/A3XkgH/NOS3M8odj5jX5M5fGuFh0Z/LP/xyew6E3ZTPjUdCT457GqE
LeIa4eKp2GOf3QXTGrlzPpwh6X3uAydfpoIQ3gUbnNi7sp7k6spSIyqtV6AmMqZK8lhtbPbk09n+
XaonxdQX300wyImigrCOufjGg/AG7jhf1E0NSoh4disFsJsJK8SpOG+z4xLpjiZ6eDQO7nm83nml
k2R4aE+Vqk2zdogAWplE8Wefoiy6D/q6dz/ORyAsos/fBmGhK2IT/I1VLpxv7KHWkVEk0rTXaMpF
Lc0Zr0ZAog53kd4P8u93q+za5vbCUEdtTuHBLXw5dH/VYwQfPOoNGW1MW9E/VHmf0lou8xpT73GV
GW50m9Y4oNkAEvMnoM9RCkC0CG9uaRyd91h3wc71Vkdj075a81w4gtB78TzavaWQdYshiF5S8TAD
QrX22iMv6OzqdiVh7u9ILkFi4LDajC/emyuAIPDD4QOWQe0TX8bpkKvotr+55O/UmfqgIpYNyj7R
LfPayMeozyPDdATUzzROc8buwwKvzb1l0sg6e6UibHi91Tvf6l46PQAfF5FVOm5rUd6COeNp9TSh
i6NMEDPXIYw48HycCXsFIzl5zbXXFAzuRmTHiF2gpzYHHxm+PtW1GGCADyu3pARyzwhEN6z9z4e6
aNCMgka/hE1B4giqOkkI3OvgxI7jQff7jDwTep4wfaUc+A3AkfVbG2XyiyfFCjDWIumpPhFkcj4H
J3co53MacuD/4lFxEZurLIjFy8m3M4gKqotdV5uvQpghXTGt/y0uQFY/FZ/C7EOsgAYxImu+Xg/z
+9oYN1YYv2HcOfXQi/EqPk1uUM+VhNF0zAlGzJ7BSdLqUnNKaHhFhCgcdVibMDhHgc6gLNIUdtfi
c4JXQoZH0ZIpPaGfWmypK3t2GXyOE4UXZKP54UJ7+3QGraRGFhsIbUPxqL6sz1Fan5XVQu9FHn/F
nDMk9cyu9gKNUtMdogtup8XOAdDqgDN7rs6XUDzQnIebkrjhJgUGMUyweuPNq8xVb31UAdIf+tu2
5a28DBDWKWQPvMP7OJwuKutCa6cqA56i8pQSxODjQgnOaao63nkQSXaElxcsHNxWLRij1Pvafde7
SDot8XEUPdwqZF6BbJ5xFY7dIclMuuJIoiQ0U65vVRxJyjcrrRpWZ+aHahZ/JSPfFsCgmqVKLRpf
ZtZWhzIIxeEnhy9uU1mRxw3d8SrijJNrTdAS4IJduSIb5urF6XdKn7y+IoE8TvQmPjChNyg4GMwu
Jl24Xh699AJ3LmagKamghs3viFG+H3JsXJA/oHx3q4hpyaB/TsIYrSKSoxSrZrSbEXuQOA9BVE8u
itOJ4rztoICOrV67hFlDT2qouOgQKY9sRQAz529HvvFkwHbZKsqoqs5cFcJCTru1hrGOFhipurvk
un+GR8eDbaXD+rcy3KuQmgD7Hzn1VjNknvtx26hws+hP4SqSUIm4c3tq7I4YHYSgdJYKLIjBpzCY
HPJ3CZeSeEOoVtpTGOav/rS+G0nBGRzKpeumZK3JNvYAuJDqDlkOM6O8Vdq1Xi/Ptke/QrWrJcRz
LHOza7MVTicpnX+C9XwoCrZLAuJxQ6iUndKevQI2KZC82t70ajNe/de58PQgdizm9HJwELqWdHai
mce3lkzdTjZi73aEG5CfoJU9tIW5xXuXJH5kKG2B0usfhrohAJMloGEJ6vsX8NZYoHhKrhaH6luJ
oD0I32M+7aKxU8YFv6vBEB2jlNVtrBj7tIs8aT2sV7uxQ63JypOF8z1XX9UXpX4TVTZc1RbYo2IH
iy5ug09qVMSDdxX17D4natFY274bhxCN3vAt/cGobZE5SI90+mpOmTAIPDd37htuIcsj90FdoLVN
IySTq8ALeLj7BmlEUXp0mInWXGiVgQOhd/up3zI4tuVFniEgXcKzRe+Jxl0UaBUTFjQrmzN5NrvJ
vVhvy90Dao//go7Lc4Zqk008XM2/BKGu2Qpi9jUEk5eTTG6wWHJ+3NA60L7p0FtUSa7OI+vNWWKG
CS2egYb2h6v2Cm12doPr8vXzg+fOrDniuZ1rDCSa96QnOZ20TGvPKE0oJ159lHtP68CwDxglW+KZ
0zD3nFbN+S4BVVTT1wVu/1iuvgJby1E2PxWEPJ/f7vGuHtmQjssZ66iHT4NrB6Pm7Aui9I8JrIaD
DqRUhvHQ0N+qRV12c3ZcWq5MsXQiUw1qGBRrwRteY2MDeCkfHf0aibiSveR48N/SQNljlqZ9rQL2
lVm29xMAKUzRtiTc5xl55JjGtsMKYtWFQQQdzsTCAmhfTRv1E5Zsij2ZqQnZ+Cv2qekIktO2fLnk
vrHaxP2OuKJxrCi2JS1duDdxfl9KyYHQWnzZqBe1EHjwzNEOsvQwaXld6v4tnwYbDxu35BIjgTBn
XyUGg1rf5Sz++jf37/VTDz2eZrGNDLRsMcc6tWngpWvoxADj9GUdwNUWkgfRftxQqRkrn8BJHU9Y
MDkNvDHJpNUvBJdycV8+f9Vp0YyhAnt9IfgaGJK/3ykK8LT1wnm4s3eOm2TKjMnOX2qW0/vwzCu7
1JwVtGLrOCliDcOS984pQcvutcLy6efP9l0tkLzghjzlOaNki5BK8Qgx3PJ4GI8B+njR8au55xOv
abSicL3Gvh7uH55E2icVoiTfJbt3A3tKsPmsr0qvU3PdJfefBubLN8tWV8BM4m/mDjT6pcVCx6uy
dU5RzUZ6G+sNLgEHHlwMtFd+WSVRlhxzpTckA1Gjr4WVvKcCx7svB3vr4eKQstmaj54drzosJ+qp
aUNX6H77CQvqyGQ1+MSi6nR3M8zZ3k5BG8otpWFeTnF/4VpH7gDim88yTgr+fRXb5oEPZlntM7AB
ROg1vh56ZWxuvApxYeBAA1DD50+Tkg+2nZcP2DZ4SXPyMAEARmSQ2f0meACY9P4SttxGN0PJAo7n
2Ohqlwbk3XfrAvgynSxRf9px/jbhKQ/rPM0rwHTvrbM9yx++03qLzyAGJrTdkSutgvwWwdaP4VFs
xAijxc32q2l/whv5GN55mv+JWUSZBHHxIIWvnxqiGiLjw+qZHJxDDrlSqYhwtoTcij7sQ4FVSgId
FbiYxYwBb8f/Sh8uX1+knwFu5BKvQeWWtJtAINzIzpGXSo45Ngs0nC4sdpXAFlqqNZOCW5rdbKl7
Txmv0yoqZ9DgNlR8QTzOkEkIBA/DxC5aCfS+OMvYbFxahh7DxxzBUDNsd/+lfWQ/EWdqb3BABO15
lCoDAAUGgWNtGUdv4QeyKArAhKM9QK06J60O0oipXAiG4F76cuRlHHEBsKZtJIV9MbmRJYukwtaI
CybGwj0UAgo3hVh3vaBvjfAjqBpjdihLoXdiJU8Z8/NcPjsphOEQPXScDseVCECDJV3lVpQ+N1R/
Otm0rTSMk2/V74LS+lyB37e2ACf2sCrrXXIr4SJ9e79+vL8lT4jxMJ5ep2Vp7Y3JEP/93Jrga2Im
CPWOpWAs226zOjzvI0U3Q2b9DtTVULAi2irFIV2Gp24zSsLJNSf7G2TwK501+i3SKf627oF3DrR3
xA4c2u4FDqTm6g0546OpxJC6zH56Kcr1dy5mYaWLnmmHSBsnISmTOPS54DaSGzIboifgN4ykbX4R
vL/QS2kngdOysaxn4iORfqps9FAUwHNgcKJwkSYgV+0OlsCdNmJjkz1ItXOrM3RzKTVtBmjyEqk6
0QJimWYdN2lqkfqQsh1k1Rmjpsp/odNgW9higPCEqTyu9bij9/pHKaTQ0REv4ENFAKRwwTTylmh+
SiBSGu8EjuztpLbWCtCTcs42r08b/jGGJiFti3vtTsu+glO/6JaNdCXnCj85ow+vqrssJIMZbqEB
VxGPxfpL2gA1vnc3OUBYseOs/vT2Ci1O0uiVI4rrDDawbPYINyIOcYzCFufLYvepEGyrEHor1nbj
9Gv1G0K/L8YHI2E38Xg1NrJhMj1INc1TK/fvLOCz7I/oYrkhcfEgbARgEWzf9EK1TOxAJVgdJ3C1
YqV9Z8W1osSfGEBxbzYIg57xx/fnDVZgg3rIarV9MTf1INMHJ3Ny8+eBWnjI2E3zjw2nT/QPpwkl
UcxCiKCX7nZSnyHePmFvwMut/SiPQgSjylEVTym+tgNspVzxlAFGnFV4ByXkEu8LO2r+1QSmIdma
erWXbqIkL/mkUI5vH30122NZl4vpV/pXHyW1HR8pV3rFRfgBDgkRuU0b0WJ5wFxdLEWVMyPt7FxK
1R7b3F4kRkwj4QBU6BJfLvThBlzptCtMbDpu26mwD7Y5IUkQ0djy6jo/UmfX1ndlYcnGOHhG7Ak5
d1QCve/HB9fP7ytAE4skpshPQs6WufSacfzEfUo/K+VTO2uZ+o4TRFXsa4TYfzzzEY4HkOAC0Iqz
gmJ40MnH5pQIBiyem+e0GaNXerb/1cuzTnvAj0AJ8BAQ/m1RxfKxeCBrhKSR2CTDKRvI0ugugEJE
KM8oxyrhqtGFvxP338FR0NrXHqoWGvO552Jcs0L6MGz85fiSB+RtiEZn52hxCD30h9nTn7BxaVOX
q1DgpKBEDa26fOROvwBQZew1PjWaP8uZN5o71FioQANSxsF6slHQm9s6YbI2ZR52vWucysBrzn7R
+ILwRql/e3loOn3tREHSQIU7Y6bHMROwir2sqgefW65RloYhqH+VWqOY69rKiRYhTV44VRJwyDCM
4+zTz+mMz751g7lIs52DIZcRIvEyStLl+AA9BqjiiLZDlSQeboBu0o6cGovPmieF7lJfU2hf8u3G
SN7F+wR1zeaWpDmv4GPYZLbKLdHTicMaEGoG3xYNc2/ZFoKdktiwSbKVPT4i2dpP90jLyJb4xISv
KNR25brJx7A+87DTIvJB2TMrC4clAEnPr9xDJ1WeRSb2FcKiwjLWKBdsHBdbc5Z1jIxldV0GGXra
UUYT1cBvzdA9WOaYuRg6B9i+G6RhaPVQw90J4jyXW1uoa+zlXuNKA2+HGqqWQInQgKKB1r812Hqd
d6RQPXwRWL8N8o+ea/ytwXjsN599KV9EUSBHpUW/koFA0sfzQ5pq6JfirqkNxFil3JdA+I2VxLjg
oK0iNsW+q9MMRgXxwlGOFYF4CfNRgHqwEIz0ts3PDERA1UylEpEJHsTuBZhoa1LJhWvXSJqIk4tH
ITAVdf1Lyx/C5mj+bpKpeQvNk7SoaGt2t9Wfeh4lD3r4zLJQTawExZiC8zcyC8M76/LzLCs+QqbU
nrCDVKzGZZPDrz/q2Sth+jW9DsZ7ivHT8jYSMzVLeDJ47yHfI+aiATBWjits0c9Y+sB4/ZQUubOP
BoaoAYiAd7vgJdQXBnLACAbWf8tWD2ugBIZjokgk27IYB2WESfyd2Y9RDZ8MzXb4pLbvTDJYrGai
BOJiGAYlvD5AZVUk8+pa26MVvkefDy43D4O7tc7pbLXxmzpu/X/RaHbVng0Sj9dzoX8X3pzBVza/
mgLvh+JcThiW4RrPBdP2fhMXsPl9lPwpI5hmbj72CYZ12Ln2e82ZXpRJttpquUERIb5I04SHTIo8
uZ0+IsNVlVnYMdbAkEtTXMbX5qBgK4jX6RSNQD1bjyx/kUaCGgnLyLZubNTEDXQTv+i2nKKF5On5
OBjyFSb9sugU7oIvsPuO7gltZmTdhEfgRJ0dw8WSh0pQQ1D1PqeosnX0rlja/Aa7+Aydzqm2scHO
5HxL59iXza2skG8CWnz2pola/ALHbP0WSYDzDsH1eyiBK3e+wT5Lgznwdmku3aEP+nTn9e3nAd9n
qaQqRRSOt1sg72aavCFuT2HMIqNuj1bZUStxM2/bR4KF6mVYFRGrjhugyF4Hs6tNJUOFci988CK/
pgxvjjixebLqoRquHYLZId3xy/hPvePEj0Q/xqzW+FWYf2Z0PJMDlhxMm4jU4Wr3HEvBIjSfj+Qi
W/rrmzsKttmb8mYcZmrtjEyU83yAWtOiPjWFQ0GiasugvsahNhrFXj7ScSBJmjyy6w3oP3qLKYol
40jo+u2ql8RzjhZsa0uugFTHiD6PkwhlY0AFY+px4dw27xtR+Ts2fTHBfuyHmI2v+PrSTMkaF2ri
ihSUIskT4TFo0900DBM2mo92GNlP7lduGugdki77PXE/PkViR7/Yux9xPtIB671Hr3QzBBXM7+Hh
MBXzXwYQl+f9tMUwcz8/SR05Kiv+BGBnLhNv8bQMlKno1z0EBGtCLgLWQl7uBV2dMt97WAtea7J1
J681f8yZIP8zKMc2zYuOzx3OaF5bOB2jfJTtTHC0K050I8pgwq6XvBP1+Qfdw7ZpiP4SVxuHbR2l
4J6Iawj5QtYnR79lPQFhJdYENDUnBjkzftKVYvf+u94d60KO7QO0QJDRY4hac9Bs4pmrPAx2nugx
TJ1z4ZEd2rgADi02O53/CV5QJ2uALM5vl83U2fNC4E+mK0KR3TJW8vWhfEBcBTKgVtfY3HPzVdrZ
h7tJpAt1uCm67uuwgut+JU+FUckvHSDVzN4PiSu502IJ1zI+MWOezLKm8K5mhPxgGVoa0IP4RaFP
zcjx12uOj9n4k8Qn96dVbyKn2s+fEMI4jp4O3QxOtlRbacSPXuJ6foFP6+QhVzPHZ8vubQ6X6g4A
QCjHg2kHeGSJnQNt1TIwia5w4GX0/wZFrfnwd+hhsJffipxCZQ5pXJuDGDNIPoCRG7I3CT9fssHj
hpu8hWUA/Z7vmI0A/93Wyp72ZYfa6mI68pzt9Q33ghN1aKgnpFoN1juG9HYBW49dMqc+5hhA9bYF
EzuCvkJbP1HBnKkLsuSvlNJkarOFZ0SgUCs8z1cuMuS9+5pWwlwwvtCE/LVDB0Y5zmo/gEC0xb7A
6bC7I/RLLqg8nRAmLeyBmi5GtsXMaUp0tvP7DQ28YRLp2ezKawoEnFHJW52bBJkJoRwpQYE2I/pn
mZQ6L0DfZFdpFLiZCzqTglk318cqjoOV3J8j72twPjQXP7swQM2svdVPwpcPsjaz3PC9hzJvT2Aw
5AaBX0AvUksUdxuC9Gg4wG8lDw3MCrxnSAi3TLXB6FmFjqS08HVPKpgcSa/EsU+cenGxTDumgEQw
kS8Xmd1YNfanpZOoVAlcQyX8Q6AJ89jsYDm+nFTzuhIkmB9FTs86LIA0BPSMuLpj8Ps4TKzPmruM
kYoDV6oDDNYg+2lJIGsMhla9XazGpoEeFOZ06S+6fELFOnsLmexHezlpkaynHGgZfpLi6rrhQ9qY
6nRbrh8OLHY9feYp/og3/W9V0x5Iv7bxX5GddOpKBdXwwUY8+NM2d0J8zRqT+roYUSCAPgTn2GHR
29Xl9teWyZ+b+GKSrxPhUNw14sfMAZ6uGQSzh/JN1Rq05wUEi5FGOrdJsY0TB0bT02/y7j195KX6
WEZdxbbo9CmjEB2UgzN0wust0CX6o33s/+e3x++GHuoMKGnWil6i7KX1UDdQb8ypqd04sOCZRqz6
mwFPVK5RqpwX7nFOfvywLdN35zqihKjc60KuLaMPGIoYpE+ZIFugZ5Ou/ALTrCnY45lS72+al6dt
K2dIm3l8iB3G3Bh9BHSQsFK8g9AGfT6B4sf3RA3LDDZJ0YbA4jyvb/0Xm1hAphxcLvBRV3m5ZOgu
FepVjTYylA3rtDnKIQaMFzrYh/kRrXfbSO53HgNNB6el+OLMINxKlDuwjtdNBbczuJ0Kw1SzO1TP
xPLp+8CImVUPIhMKSdn5bhD6WKK8Ml49lBtl0odb/GyQ1i7TkFKwale4WfoSQTL5A24mNMvsSya0
YRZx9Y4o5S5S8Xs7eMw+iJYttjdT0/KXuJW+4nzKB1pNBbHs3UL7fjnc5TcFvAcFiZMxUrSezXFi
c2UXbSNAdV8DOiwSGVqNRevVpg8PwVByW6BLmMiOKrVGh9Sh8pyajhIxxkw6gRuVD/bFyw2UBTSZ
CENvNlx4bo3yOsoze4ZcyHVnIemIZqFuFbJsJ0ASe7NnI1uA627ZTVMsY3i4pXS4RDa9C0q8JYOu
Rm3tszZQv7ggMpzPuY0fE9G2HR9ZHYmNWs6wRleP0sNmjSwe9Ry142XFl6OfmK2Ju+5Pb9DjcMWf
Sq6AH7aEmDGq2kWChCLrwjtr4DYY7/3DSK14PmYn7Bb3zccQsHDL3v192u0jc3WSQkBUPtQsORJA
L9+VvAC5tjeAJURLbwwG1TBZ5nrTzQg+ZnDHis/pcxoKg1g6IZgapUhVbONLH3WaX44sAPVGItpl
FgG+i3RhZlSeNLobYC5AfvoaFf+onI8luGmDEg/3WeCGcNPjGu15GZwsDXgOaexyta6LAZkIpMLr
CJjpoMeqJOZvdFZ9ZSoeqgbarBAcEJYkxTHX1iPLLp603lOgVbGxeLYspKejdyIjfUZnNgIEQf7n
kTKjB4gZcs1u0K9weUMwyS87zrcDI2ManJ30EJXxM2kUMDcurDAvkRNg+r05MQz4aPvtAye4H1Gn
gu+fUSy/ThnAZyheVbt0cajoFyfBaVbPvSC4YQ2gAqf9Q2E1lEVw9IO7UgAvLtj4Hdv7GGKdJUX8
848kExpOgsAGz7wwNYaXlVJswqYpzsTWLvXcmsE0Ycy7k63uIYV40u9YSCbG2iBcczUnZbtkGWn9
8lbk6CVqtaYJIbuLdG3wV33zqNrT1JWf9sWm1mUwOmHxEMoqMOehpQoKF7QP0o2fdJkrO0tS1HwC
3uwoFAzacRajrYs99PEMVSBAk/1UFSz1g/n8SDJqzvQvnTzOqfmmDRBLTrAvyBTrt99ZvFImETaR
Hq/vZ+Bvx8s3T4oPY/GXUie2fJoLe70gNcfkIMelZXU6wUypRsoMbnk053AgTRPffoBUrmHW5Gqp
SwLT0RxyiYe2yPLi7blASO5pe3trC7NACdb9kq9CheENfZAxZMFVED/rnKqkjgXk4Dbq486lFQjs
2U1HugbLWhs6+vCqe9Isyk6oK902/mVwgiGH5yGvawDEXzExLEwNbwgMz1cItmVJRNpSKMeLYKZu
w32zh5+IBvPfrHHlvTWO5QLPQlXg0Qcypc+R6e7Z9A8OOVByzbdifjRGfPxJ6lA9JSYBbWaI+9f8
7zMEeHbYHof5J2EHiGDesKYYn6Xmt4+8dKRGcr7dk7Ax9dRO5VQyx9H6g2INBk4JFoEHtRY3fK/z
mZRJe5dpB/3nrJYC7oSG7YbJsFFnSYa/X2MO2WxFgCOtF0H7VsBSKpUurgVp6N9Jxyis27nlYpXG
ibQSnG2dJq2lzJQpX4k96we/ALLJXOnc/Za9LBWhcEkdrfHxhOX3eQAOJUOiWvguVrWVKOHI8Nyi
O16ggdiu6qJ7yyrOjakNkoLdWwpcFWYSuT+nRQJVElPtzzRlAGQ0zfBlbOLtIeycCDmDMtssQwyn
jMWjnhwZLAza9a4iW3Lbarg+atU9z87fJ6a0xwwTAAAsEYiLkYxheQ8KQhlMxlN+XukU5bTZq8EC
qmjg6WuV3lbmnEDwvsbGJdiO6R67MaSdagwjljYVjqXt3WO8/rP8agJGoV+3QLQzV+UC351iupau
Yo64xNJNdNEfz37RSGyNKoibuLOAT1MTGDzYuwLJuUmasUEljsEy1nIkekOPbF5agSJtGQCit1ic
Rf4dNW9S6pICXnFYRkQhD2CMJewHUlLe3hI7vZZRDO5jg7DYsBP5tgCfou3ReNCtSbl2bXaXpmo/
Bg436n2w8IQrWk7zwaWYGpBEA+RsDAj0P45oMy5yRig9GZVePV2eldLfMSOayrjeXaL6jx/mQRrm
+t2UhyP1BkCWm0uP9Jq1bqWBObLU1IIIZh0M0RYNkk2WfE433et4g4jXhuWqAKBsyXD0LvifcD31
AQjdSxYylfYRLnjz5l+6DGMFFrTM4EmEh8G3FWtGQuHmHgkNEopIX6nuB9T2AgijwdRcMrK0d3J3
32PemGrrnvNSHw/MGPLL9C2TtTrH8gSERP04YqcRY1vB4a+T5WIV9DUZtFlcFTYsubwiiKfYAZAr
iafK+YOktrJVoUWIP8kY1WgTt2WsfXBp2lLsKDA54A29EJC2SY6sIUp74zsGkz09tj3NUa7oSrOe
QG4ni0a6anVsXZTqE0RRuXe++gQ0y2Bn09s+8yw6V6HFTSC048MhRtEypi76szYeDd2GQ9+iiyHS
OWECeW4gJxwSxYTncWie426eNCrpKp0+mg+jd1vhu9CqMTFIp093DJzzLnbI9Lado71pQz6OG9Wu
IBmNuFIWlMSGq5+Sj15JhC0EUYtVYkcUgDxAg8hlK/ob24jnEs5SSpSOlGHcHl2Deazc31PDVswN
3QmEjTPcGWMpjgeUZA55XxYG4MmXZmusjETScWghL3CKxqAq+6T1u9T4uamkEJtvoKiphO/nUkWp
d8BFHLe8d7DlQnxGK+N9AxtW9CGPdHUU7U+38IR3Faisuy4hDmrE5VU8xMOXVhcW5k7dM5/ygnCx
HOISCXC7GD9u6epk2tjK78gaK0hgcT10gBcPb+pPojvSPM1sq1fXhaLfT6ag10C7DM3XGnAPgBpq
4xT/uJMCmUAI8X9aUY7TW0ZPSu8FEmyXFZyIKzKthlKWHWgpsbiH5BlW76KTW98hKZ/GpJWR7G6s
qJIZY54FTEHOpNgR5QhM9Hy1Kfjp2pJDWiOJKo5jqVppVXbAgEcdUo9fK/rxxluNFUSkIfS3yjhM
UblC14koGyAvSV5pMKp1svlOTU22aoAgUXV3Hrx4sd+Fm2G0dga97j5R1zcKs2n9yu5xMlhJqcxD
uwzXEsGWSiXjDSpk58WNL5vp3R4SzE98Tdm57hIa4NaztZSMWeDH5/7tU0g8dGM48az59WnweQwQ
GHCjFhZLsSiZGLFwrHTZjJCP+HYX1VtgI3i1rD7/3R+NDxrLCvxGsylHZoDhT/LmqH0p4qk9TQJ+
h2ZnhFsZborDoCO5rR6siP0j5efSlL8bABYu0RzBqthcIiVkdLaQ/KJF4OnjITYeQmGz+tcqVUap
nGVDjNuTGH43FNpCtw0HLXDXvOepExrzmrq6w3sCafCCSDu5qbnNax4RBC45CCvAABexz0scTJu2
Hqj9Cfz/ZfGeCrpffYLAjfpl2jSG2l9EECAdzOnUvbRIShcqDUpuWPXHy3yB3tCey9yWZ0BY2hP6
OIM1u7j3rJcINShN590STB7Q8qffZ8OLSBzGCKYx23A6eSQ8qVQq3ZNiqkuru1fqiRI8K7mFpdEC
loMC5QKYfe2Y0IUqh5ISJxbsd3lIOtn8SdpfRN7tvjZ8jfEPhPp7kRdhWbfJ0L8jzBCQfdui0Gmy
uiqi/7K2qMVys2fKMf3LGnsk8gwyhqDbHWBGz5SbHqMvqnsbGPRUB72M1qdrlF/vJH7N2OEpDnaj
NyV9Cxoe9ZptCS3M8XBnWeC/Hrxz9ljF+KQNrbhKHYX59Ubdeua6Hf+Thb5wFbta4L1IxtsGFUZh
1sPOuBBcLSiF3u1CQZYpYHju3gbUTL8xfvUwSnj3KH3jVqAFhesC3r9/bqsJWEzvTaMKUFzePKMR
9LHyIGhJB8Crpk+//KQPIWZeFOshNmIl+t3pG1a6i8twvPHELmmu2mvj7dGRJPEOnB6k4HTk8yqh
CjXUoAjiYy8ukKy2mW9zajApMPO/vGIjGFJWsJ42acbsX4Cz9722f43GhVaPStQ99r49mo33C0kO
w+rdUFqGGA6cYi+RRf8t4mjE72mpPa6hkDtPBwisg9yF6+KB/QA0IMwZDF9xJT7JNU9G+Je9fwYY
l47PS7i+pXMtALRJX78uSDrga6MoEt9PImyQBrZ3ABqzNzuuvb8EGgZ5MNAR+K6TJkDxxo6q+g7G
EAYvkzML/xLgigfUzhQ9WiB+3xlBKdNowRqTkBFLutCJJGgVjhWdOiCzxi7D4iTn1EPaC11hdauA
38W/pIITayhd2fvBV3vYOPHIgZY8XK7lxtp6/+II+Mfn8t4BWVj1u7RmdHH4RQqIAWlT+ks7SCOA
vrlbyuAlX4xoC8qdMa0EqCXYSGp5+rElbpnz88rraEkDaa4YS8KXFoGB4OBnCPzxn3FMDf09CwRK
INp162v/oo+4LN3kRGggf0JMvljC8DFtDzCa3tVGx7S+YRAGcoabuAV3atATeQGg0NgQq0JME3Tv
3BZNR2Eg3RMYwS1ne4Q+zwdYciCQGynDT2nUS52olqBXNd4hGhVnXbfUxwLvyPidbqy/bQm9FkP9
88a85996YvamV3FSFq99lZbC7QN5latmp5LcQkI//WS75z64bDNaATzAmhhlj7vS2apMCT1S9XZH
kXR1lOfjS+PSKKCvwit7gRpOGwUUlVzBlEObLyWxnBuBo6Qilw0gx8PgN/TW1TDqEbUxVNEX4Y+b
GFkt1Wu+WrNNZxmX+fJbwPnAOGSTuFdeiqiy4iFzG0pxrtUWjK/szHq3ZkhxLxLTeprMdT9eunAx
rQzKk3JlT5VUy0RKpK3cRUFLo/068fFiGUMHWtMTJvI7MFPRgDqYGrDDzFICK0jWHiq7aEGNVPm4
dZ88kGJwLi9ZeGyDDnfd6uPFzFfAefRbwaPJkvMLUYAGK2OovpEao+hgvBsI9GyRGoQIHjRRg/nW
Uu+MQjVDUs0aV4sdZMRHW7Y01vZlJWVhL71S+0l+2NORy2vnsj5ISnTviqkWaYgS61bhzTrK3XHn
o2u2mVr/v2siLyP1MgLpGgyrvnoBz0L/9l9mla9blxIauJ1bLcFRCtw+vcvdvpMQAOLjAR09wI7Y
gei3S9L1MjJWU7lhLympbb3a37DACjE4ZmQVTfA5kgHlP9lnuXZxPiMh2YGPPcqiTF/wNpr/BwK4
n5SylsIDQfd2Utgs269UHU/y9dvHr+vxY55FjqFPWvJLOH5KdgjL3hN+G1VXd7gfmHahMh9chol+
2MZKe8YosufPMIaobKGuJ3GE+sfZtUsZPhMqFDN3Ask85wdx0vxhLDwqs/xrTt6rWzdi6cgGDMG6
65Ct5U6s9YMB41kiiIl3IP0whMewNatRWjsQfvgxcxiumQjbiT4oQvqC5ZVeFjKBeGlwLF8vHmTg
KZiSY66obY7p6+6hDN4Rr+k0rBtUQP29FzhXy3c/FVu4Tf5ciWVLfMY8CxgZonEno/FwNiT0u4cu
dPO5Il8WGLASxrNUTR785ZwR2rxI/liQdtqDdVOKVTSfGa0sbVzbkF4TrqjdnqzNXSPZIq8O8HMD
W7u0I/J50Kkf4De8QyXWHW192PCDAApb8zEbhkuoNmYwVzaEmr0NnbFzo6Z0bgbqv5yapCY69E0J
yHcb4M7jzgh1uxW08kwvsbCjCh3eNSmb4FPl0EFXKMlO5Zz6hB6cvpxAnHD6bGFTxcdZxTZgexxA
uWWc5I2RidnSbOiClTJKykVsbBSm7jt4mo1Uso5DwxgKs1S9mGZ6yNopWJSBIQcGTMc4H5GP91+Y
Ttn6cQOwy1/IskImbgmYQDwBpY7bMhQsVVkI9HBWWUUbqdIgiUBM2bx3p83+HMnF29wZvt0hkQJR
eY0AxPsovMnFhRqUi7Nc91qguhEgLBhNnWcxTT/zxOsM/TAw1nCvZXRuYB5ukibRTDYiw+/mJ3oZ
4o/ri7w5cjkX2vPBb7m7V3LwJcjyZqEETz3fF1i+r27L4R8RCra0vgl+fbTR47+KmrTNyjS7UBvU
+DKCX3y5BsqHSEKoLnWahEGJAT6w3SEcZ7pxxbANSuT0tjY7vUs79s2fzTuF09kgnK3UJVWucGS5
zh3eEJ2yGDdB+hobYPn/2Pw7z+Bl/u4mWNOqZLMjvhggGSydhNEfJlSnNLkrZ7NWsLtKO2O+KYND
ZwnfYKY9bz0Ikh+zfy9iDnXbKg2XjDBjz3no/CjDlGXXwlTi1enuKMnVpkx5jWes5ivVG8ToFPcP
XN0BpdYYHYQeNf0wHId6YlFq1v27lNKP5R0orWzmQbxQhJUFnGTYD6yQqqQuTQ1bMkRJWjUkzMsK
K6R8r7VDEFsCQUSSrJWEyhRcfJhD7BMbAK8g84lCnR16qKk7k4BU8rHKATdEOMD07f5ly36KKd53
rjT7VSpHWCEcSeJbbXifhvcnEy2LdsXCQjsq9GzhGfxFt6SacFXCkgk2eUS+1RBfk4qUDxGspe6E
87VDczXdyJ1BDL6lGIt2kEWutIE4uz9dHcB/pxbgwUNU6T5cIuyUfxqfoQ5E/IWz3SkX9hPa77q0
TFMeEGQca0EyU0gEh1s6+mP5e0XBZX21HPG2UDQ6UkOcIj2LWeKn/H3j/rdN2Q5EM8B11NrSBrZe
J8YEuLw3/Zg8a4LVQaSlKynhwVCd6OZUWiZYRRydF9Y/Vz7uNdFr0ma5kBz2DEAMv1Uk2WBzKdlz
wF4LyMgdjvBNsq3fHT1HRN2grnGMHQG1Uyv/CjfyT/ENjCSmawFdj9biwI6MvYgEAePi2gmS4i/J
weUM1KTs1y89ubbKdibiZTLieleW8bpMzLgSRqvg9T2MJ2fljNbIv+jTNpxUi9HtVVC6Bk/X4dRs
y5bqwE0l3SO//lzDWKu9kV8//fBs62Hmef1oX2rmE0DxtuJyDOEhLC5MCSkUp/le+z6HrJ6CngPa
IVCXXRcY3P4z/YU9nHu3z7NjwHiqWBKdXboNLP4fD+euZTUuRCm56Pm0tvDpWiAgDHBMeDoYTOQj
cpvzma1UDOYVjBh17SGuy3XtvCG+GQTIgbR3zBbgfI8x2+9KeBrDdJI8sE8JpxoP2eMRUqrwIH/2
p9sVm4ulFRfj5E44TIrbGJ032ZfiDpUaST0WLfSXuTynALhmt/fGL9M8ItPoDDCMRdrOBP+x/yNS
DKgh/4Z/UFOZe2KUYS8u0cAXLK7chwNbth6uhxG8/udjfCPdm3u6+d4KHrgsX84V3GFN4Ws87Cmb
CfakBg/0l/Wa6xgHVQOwE/520Eu/z5Uew/YCZvYHWZBGPSCOeq7kCl2E9ZrLXnUY+1gU9R0isHeN
bfldCVdu5j/VJrg2/msNRVsVHvrgqYfie4xsiINCqfenuWJsD1MFjby4jebNcP9g20M9slVwxkP0
joxqTnlr6Aim0Vv784lN4de7z2gt/KwBB801Kw5XbO3pWj5uwPEOnPgT/kJHTbezxSDF5xkadKS+
gcDxFn285O1cL/PhB6EICZTawwr1ePUXv4BYWrlLn81kVEnSAGpIzolE8nd3jRlyItOAcbJw9616
cZn9Rgfu7jcTNmR6o48ziTicr2x+YBgFEESIDCH02Yo5jF3KI53KefFb4w4JaTiqikVQenfK1FKv
ZIYMnvCaGrObxn4lBnsks9jvn0OSa8OA15dqlgiOttpf8ktl3zlt9kuHsPvOgLfLKzuMF6lPIvuV
HFpSKxfoyIR1NDuoKBwLIHZS9XdSU8T3rIhypHZEQhvUelw/ZD7skyqM+T8bNCjzN7AcgHiDqStO
nU3f+Eg1qzoSAMyp1hg4ScaLojvoLQBtBpBSjiawnG8usC5hrWxVfPJsIGVDb7GmXNkgEqgezBT+
Q31xNfVV8CVWzLRv/oTtX84unRYfNLPFCyGnJfFl3rxrWZtl5mZw8bgUfWFMNm75OHl+rfmV4zJz
0MjUvE1Y816PFMzwgezpJcOmr8aR6fUTD+6dA8FczEBCnb1/7T8zQ2Zn4AAxHFeYiYBUthZ4J5dP
V7KeMZyUTby/ZY+6D5VsTYrM3FozSFx1fV4bQ3Rl6w4iO6JaPOPnMcToYm0arP+R4xNfE3oUx/te
uEZxsdcFdSuu3h3K/alcFH9gSGqEV/DhdB12XSsobRqaSDoGoxTTTUEbpTDPKx79nlERS1/u2T5N
iJ+ltUvfDmNh2Xsx8LaxHxA+Y1jTp9aQLPJOmvSdb5VlTcfyjTMt3PPXqLMPeX9FJdQnsR07eLgM
0l2xjzMpIkboJqAywCL+E0RWHtqmOWdfmb6TbZ+uYPX3V8sQFdr9nw+iJjlNQ7YZwUWnT0QKZ5qU
opXG30H8VT9YQD4sbrmwCR/XmuV7ViMityRbCUAM0bZOjNiyBVLJr7fmH1Oyb3nZdxHVTyX5S67h
1CYYUnd8YQgT7jvcRMawSvzONTc0fe3+d6pj60muotpKk2w1Hru5gcGSJG30jvxYzYFXTWKqTmJb
IRUgWOqiHbLbx8qo/M7Nz1i6gDM7x1nqzFAD7R3uiijJVAarJBcqUNkeDVvQAGB+C/g+GV2bpNb1
MSW5p0tj5Bqx9MSb+4zQi/opW7WOEFlybeZVG7BhVGdilaCnIH1gBwBlNPrTQhedLdQ2WmljleB0
X0/S7qEWiih3tS3bp9iGpGzZcoimWwT0iUoEutIbD3L7nTMgZyhdjFKQ/DFxh4JhLt45fI5OXb2q
ALGwAt+hFrZCA5h8BAMNe0utFpR1f9Ka3lI12cqe19LBEvxeAyYcTaN48V0YseghaIJbZCJVucIq
I8hTQgZ7FU63p5emUi7d1TEloDLsQJuEgjqQYlboiHye0+eJm8ARz6FdoWEOA8e9n8Wdam6sVfWc
qznZZe2MrOTzWLV5zISCUz8iPsXbnBm3I5zs0lHLFZKNwV+cUcY/2M91Yjl1NHLs17QPbmMvFjlF
qHFlcYM89P/AvjrQOK+OVxqN7arNrqA9O34kIHeNdX6pnYRTz49DPhYLBDE5oQQZobJnx244YKYK
3qGzqARoehmUzdUt6NhNwQ8QJQmH0eaYpPtieHGEs8lmwCiyKqYXToc5p3hWXOT3V1Wy60e7Toey
PQDg3Ij20EZhglmxx7K0lJHWi/NE+kN02zo2scpZk11W4JTOLmRRWGr2o6Z/7gwxk8Ac61fwytBO
bL1ojAyxl1tvKYga/jlPGwXRUxPWIma9JYiyXs29a804+r4pv2tiw3Iz9yjZYi3j1pATlqsqQ39w
qA4IWSKMG3KDTidOjW0H4kiu94L/Jsm7qxaZ8DVssYn0Cjrez0NiEhYUGoL/TZTPkBNoxsRrqFAM
dgbJyWqGSWr3zrpYFr37Se89oMN2gW3NdjZNJ7Mbcu/SFL9z6b8OgqJZeXNU3qaT66OrKYG9Kqlv
WnxZ3kKNeoXUbl7owqE9U/T5OCG9k2rKP/YjSBfmTPoAhl0GGh2S9U7/3YiCHotsKSQtiWem3p/s
ZvkizhOHfZgjNGaYxqVxfRhiKYXqVLc/EzjPc2XaMIYDB3gZ3RGZs6Kv5zKWNKjxLTYwfvdFCNgR
5yFusKSckYwpUoDcsxhUMBRUURkZ8GP+4QeF5hI/lL0jzFDv40Fxm/RXxCJDxRFqZZqmbvWgh1Wb
dwEVvICjaD2UtRYrHeTIKMK9v6e5rEvz+EtwDaIKJ2Kns/J5hJsv9gff7LWrHWVLxJAE3T1wgLzD
4dthfjpNHNUy+Q1F0jhX0rXjt7zfOew8cfvl7ZL/GHutQDM7yFk8REreqbdJ/memAFmTFwbL07I0
E3r4QhAJiIKEd25EvbGUc6uMtWlPX/wHMMOAdcJM7bxHX1+EU0l3OUAsSuOGmYg5yXZ+XEVOjiQJ
8mi7H5ugDMqkkQMabCzxot1sUDA6fxnWPT9yZpyKsTmraRSvEN0QCvRc/EbrhiyKoMX/g7q7Je4u
WR47MFbsxKuI5xmZ3XBc1J0QMkRpiOUXjRMvYh++zKSYeVKriPPbzsunpiWkCphuxP2oACsGKABL
hk6mlDFKhKY+TSs4pqusNYwxvjhzqEQGdGWZPmt2TFRz1J7KUkXZg6NQEaZzJCVGegcjEYRY8VbA
bczvD/xaTWrSbLvDQZxPtM97DAACYkZ8UTIgA9vPj0ctUs2gw2yI5b3l/e5z/V1gI3tN2jWbik1B
tQf736zR7vBNX3z+/qL4cAuiWaL83fShm1DCasVqzmSpZstpOEGFlbYdnm2H2sQmReRjsmTX6dWh
XEO+HKN35K48gXUS63GUo+IBof1OE98+S4F4rtk9jskfxEQDcN3+CBxRwUQnv3HvMlwf1l1ERFe6
Mb80I20vWQrOgU8c80O/GRUWjp8YgPZ2cmxDpo3dY/yl6af9GLMTXczUipv5ZardjBs38xgiOvY/
vq6NubOraLhd0ltZ1lVVRtT35o/fpWkiuZS5m6FivX5usl9jl16Kvptf7Rp3aFIcVZzF0xdC6/J+
DWuLiSG06dn6+NsG1ilaoPdu+34SYFHC+nORChHG3hjA00xT/8F6VpsmQ/FGDpQFaEF/44ghWZ8p
kaxZv5BiXjpqJOFvytyqQ/DNNo4Q0VMAjQxMblpQQNdXBxWVlT5rgz5+Q2EGR/J7zLM1I5DCULnu
V/zNhKqN5GlNQz8To2GuyTzBA4a36ikp9foriJJZ0ofGkhZ2/wuxhcrFniXabFngferCKHwcpdOk
gCIYSnKVsnDACeYA0IrRUduLn82IbmNagzM2AG8AWxpVqGxJXWBItFW3SNjA4e6In9Nads/eDIoT
kakgZAuqxLkgcpB43AsB5H5LfpctnKxspd0d5zh4ESTF6Ka8LwUoIKz0iGe0Ka5XRY8UNhXvGTrW
BzkAy/t/qY19pGFwnk7y+1SIdmiI8J43j80yIvvfkVcKcYVY4tk1QyC+9nr3MqNWzX0rITdslaZK
9VtW5dTTpq4E0c395ISoyn+FEwHeM/nXjqSD0R1zCtmIXSHGnEPlUhrCwD19OxABAQm62JrV3CCx
Hxp1MuF8HyYczhje5i6xtAeOcUwt03mpuL4UcE9M4IarDU7VaNWxU3JAEweLX9h1uj+pYnTSxzQX
1YphJraTq2belMo6vGQHSi931vtj0CHNSgqts3AWoM+0PL/F8yfReqo/xfB3NV2dVdVvBwvdCq5C
1O/N6kRtl3vguDmj7sg9hI+hc3owYDGUpJNpWYrWmNcpJ2H6xFhF1SjL8nPl3IPhN5d2QeAYOjh2
U6SJEw8OMauuVGV9I4On3XVAH1nM+RepjsQBABLX6E0AdQdO0aNwNaaJfmtr8oITifxACxrO8tB6
IOkBecilkrtpkSLEgSCBfq2YLpdDdCZZdgQXZivHyNZSJqRK7TxrzvUJxz9GDFsIbYGKVYNb8JLw
5N90YtW6UT52KuIxtQz8bncUUh7kmlkEN+qbteCswyz8nE6bYl0/Pa8fayFOBsqoI5EVxG9Yqpys
ykkr9Oc3jG6FBhdsWpr6aSCsDl2GMjWsLlrTvIj9NeYjS1tV6hMzZvAcbAJT9Fl71417IiOtGDIN
4Nl85h0pgp0zImpXdtaiCEJUBhfF6H3acTU/eWC5QaJWx4DS8aJhoPcCmrDQq/z5IgqSNKRLjrjR
TOuRuxqNTxfN4XqSty8Im7O46vD9Mz7okAysAH2Ziwp8H0+5Rl/rkL812Q5i10nI7fZeIN7ZJfCP
bZLf/mlcLrDYiT9nAKdfGt6gkIii4S1QE+IDC/i3AoFnbBIOr73Qphzqr6Vx17/YroS+EAodbzuO
VNMxHOfgXLdIvW+ohNUiynhyxBUZrdKB9W5wPDbFUNblZxIqzBO/cjZB7ub3kgVIN1BJ8GYwbDxk
deCwSO/FGP/JpLPO7U+f6wt4B+U+MXXSX0/axCoGWnnS7PeRi7zp+GAyYZ0JmrXpviyVhzrkIVdy
jo2lFvAZd3mCocmLURQuVRhTEKA9lZiZlLTHVAbPArDBrce6RHToO1rF/XZePlQeBpG0cZSNpNzg
WLajrFwX7jVCPK3trBo7Z2vGDxPvb1h9DpB4uATzLmXcN6qS3CDZDtxoqWxuyOgJDn9Xu6Aaa/82
nA4DelGzI776yW5mdum1wZZa0S6X0yXu3E6MibQ1GUfircHCxo5320KdB18lKnYlRlYGFn95wuc8
MUd0tkSXm6jOS8qFIXhwKaCgu2KZUO4Y6rm/7xwdl0dkXjl/QaVRLIws2nOu3DW91n3T/AtsWOTH
g1YVQ1djDNwoBLpC9riG/dcH3pYGTi/n+TwFYu+ZnTRftV/F26HVf0PASPZ3kiDMC/awKPV0Ex4H
5mk49w9YW4etLAgWEDhaFWse0Wefgp4AMpQlIMdBh+Rr4iagiie6pvS7RFC7yHjP5WEwnP8DUBVh
F4KYSgDX4tnpOnI2HmgBdZEc/fVooCGMksTTIsZVbpcpDsk9jyN1GNkknmcMC5kd0095KusiRj0J
URZk3rSbYiqR/clktwJllx1u1m9ydUEROGyLneKGs/RnFrGibYJ48TXa3JQyLmTOTrk7l/IsceEk
f3+BwmxhKCHzbX466xGkRvxKnvk+Qy85lp1IDsOzKy0T9eyaaqRxdTU76j7gGM56PknWJncgcfLw
8XQATEz/ezBasuU7wGaTilyZkNZfwoUypDdV6oygMEnZf8M91p6+mfCiwppRjTSGm2CW+rGfxD3z
hzOCkBCTABlj4l/xypHJXQDJh6kapB62UdQ2SLWcxdvxa2OISRzBSf+iLqSumNaVd0l79s6HdgXa
I07Dbz2VEaI8vxqDXjo3yOslkNn6TjeUW1PARxCVLjlG+1cn3CUHAGeHgNPnDL/ScZqD3G53r8W1
uDfEflPwIdyalsyJPgN7oRMh17h4pw/EvgWuQbfa9w/rJxmtCjuFKMyKnXOutNZKWBVyROAPwCHQ
dBGPwTUd9lWte/OfWy6fJU3U+aboEW8qcvlNUPm7VqvFkSRjAx2Z8uEd9vLesqzPsFYsyu93ymvR
DERIqENrXQG+VsdqPss6WTpqrxSbfEcxc1PvfK67cb8InzJoDcrSWyMLpumsJk3NTRvsYAPeIabW
SqJYRCH290S5Wa4LzeCOYEnaNTT5aPtFSWfR0ut2VnoVEr/W+XwJpkxA+aV+b8wt+lNxgFNLo89V
TNTLcLZcxoD/qburTQQDVMzmzT+TEVIf9X7FnfjuMYfYfznqtkXB/1hfEr/n96k0UPTBrM5kZI2R
+yF8zZEjalumD7+tdpaf/zyKXv/97CC4veO5ogldvBko06/T3Qy9FtCRcHg3p/KLVM37oG4WJkL/
8AFvGj7AImzFg7RdSEp1VuGHn0+yyB+e1czqwefS8eN6zNuF/shnAkahzVh+lMzYd9ajXI7K6Zfn
i+vBQHZ82RIjtqKny5NJ7nUpkYM1GEuoGNTBB+kCtSNs8FKv7d6uObaP0M9AUe2hYzhviCaSZ4Fy
zm9p3GOo4uorKR29CMzRLGGAt77TtlXBJwgYOdBZ4VfHKsfGfHpe9X2kM+PUG9pwI2/DtIaFYKUB
RpLWKh365xRdwt6y8YxJynYjKhZUFkd+JGccxGpR91SyxMBiwnIxsfqpqqpIVeuO8Af7dyFUIl+V
pijTAMav/WosVVBQrmzBYZpUe/GU2zgvmlxFzzxme/KZcRE7AHNl6mBqVZQnMVzsem4mmMWlhGw/
hBN7l/e9vyQUj8ISFsJxVn7a0qBlnab/F3SbSO3YMGI7LlTcFv6BgrkdLbyFhM5svsjObEFxsD79
NufHEKlUiCNrhcvo2gMFNS1KU810WczS/GP36JSE5bQ6WcnmMuokEhMvkM4EI9DetX0lgIp2BWmk
8BB3boytIoYO8YaPxtJzBIFqMdafo8t+20fIaZTS9WikwSJBPMmureLZ2acROZjdsH0zdT7t+NBC
hpHPinLrtCYaDyh/TPoh++UtszvDb4gMHValQZk+38vFbzVVWhcjjwRJJ1K+TFqOqkDgkHntbrYm
kRVuwTEqcaZa11rSZbH3ZcZ+v19i93C4lzqXl7ZkDukpmF3f5C6B+NJrIA2OAy+VNyunEdg37VzX
OozOuCsHJ96kXU8OweyuQOLvc2rXUgyd7CDbwUvuQ+wn8zLnaNUa0stPEXhSKjmOYQf0zXMKeZzo
YMsiOEAk7sNaF5e71KFnhDpU33mLCylsNSTSVdl8LmUeVVjqHgji/iDDO3nkB33/EmA0qEyHGrQc
ghgU/xk1oFg/fJYpV2tUHUomxXkFHkdOVeGnj0tHsI+2CjDXAc7irGZsAPV8iBO1doZ7FvMB+bNy
+5ZX8skWjV5+m5tV7I4b/wRhzzmRcL2OD0GnbxebSD1pk0H+YfQP+t01BrZnVruU+h7/EuNPEJcc
OQD+hHu3VHQq7SqVSpAkKN7WHpq6Q7YiGE5bXtCtvXDEA6NGCt186wcZphmHLfFCKg8epWKmNYHb
xtxYemS0GuJMobOIdmWZ3wynkofvP99XzhR4607KtJxUSVsS8JjqLXfiUqdYNyosDUJxUJh4ZXQS
76YxuqzDpt/IY5qmcvV4HJtVq/h3U5USsh9+QurFX7E38sfIX3dxvsVquJeuh3G8Wsr5RAW/f7hM
0VuZZSobw/v9XfsGo7BzBv7P3CT+PbuQjiO8qfT1dylx7d4ojCkGoDYS+Xxz04gqTQ/GnEnkfD1A
c7Wo68PrdW+JVtrPZJW18oiGC/e3eNiJn4kHv8obpTca5dbPxGuo6wGU+aZ1BqR3NtutcttGIp4n
QE8fHGkmwXzRg6O5OLhio/emFpbQG7GJ2SmHauZmG9f6Y0EwgAynhwL6pVuZ1NViuHSuu8IZKPQW
/Ae+u39SAu5do4Ixkgik8HwNcBNPyRTAhRh4GwlRnuaH11DNV05bNSOBd18yyQ6SuBpYoMqBfiId
Qtii1z2Tg/77ZIQUg29bhfe6Hh8egNSaMuve9rVLSbrjaoURhGB2OjJlpNCCGD1AWkc5TOz7TUK7
W6DpLe8pyWldDuM5PYgKP+xdzAdJAKjPWKcjTOGKDYakqOX2q/FULHXpxTPM0ExS+fjc16oQTf3b
0PVTXV3acbQRc1V/LnDHXZlPfO2Ig6ewvAwjjt7c2/Uxx6jgT1ucmszrVfesXFyHc5RVJ7sH1KY1
AQHhRc5vfwliKqVdSPx8jsiJqlMQLQExHziarDWkPKSWUEATUm/aTGOQREttmOzZUZQrVyE9k+dZ
w9qEtrY9+Z/JRsMy5oVVsDqSFvgFc8KMB0GRw5eBEZu59EDxE36jkyO8o5wHwNFr36QxXA4mohdK
zv7vJzWrqxJeOJ67CJLYc++S0hgXzDbiiTlwpxKN3HFfGnZsqmlJshXQo2jw5khIEf3sO9+5M1D0
mPyVCgDkEG0JUV/s4WjzjpZL3ukGBUfOcZL6HPpXpR3VpQzTr3VOkbpl7NYy8eyqZnjp4B9EyjSW
2ZZChLQN4PEdAEF6D/WTZc6gFz98AkmHInczaNHU1p3tbCV37WYOQFPNbBOyadEFpMviSF/PKadA
hSHyVWTK5Q2P3QBvkTqx4Sb8JCs4Q/FIH5maduqRY+6JQUWPqUg/uDDHIWgUO3a1wE3NUIUc6Lme
JRzXuBn8nfmhhD4vMrjSVRGI7JDQzRB3BUxDC9ME2+QSF9wE1j564QvgEjXhmIEjYY9zgV94RAQ/
MK3er/w46A/BuWFAe/hKhKsyBi3fNbcpFeQeMcFw7OLB9veQXy+DnL2y9IqfDntXKc3IiKhM2bHr
Ru30EwOeXWf4xLcqyFLj1zUzPXIuL/hneMZgrqFsCiVmYvlPIbUb1rSunwIzWioEAJpPspLtPoRf
VR1IaeUP0JkUSDZlyXN2+mxMBlFfiiG6RuLtU/qxEheHbUXCh0kgbB097QF/SmBY3Bs05IXLdU62
nRMFAQaJg6csb49n75qR+u/mjgcEaRZGu+fWhgYpvZImhrpkVgdSxuK/HCMtL7MBWLzUd2MANt94
arQO0jH1L1jvY/uAZoPEsGdwbTXTxmVuzg3v5B3UnszpkDSix4eWw26O18NrJG/vatRX8lCWsMsO
Tn7F6tnh/xgP/wymZ8qJ4RffVxmwTe1E9R9pfYB9O/N4AtVSHzXHNBXisA8vqqSYVZG9M7Sr8448
WlDDCe9y24LfomnFERcjQQjZD3xZt3WMwRtb+93LHS5KhqOGCpnUrKRL4Fh55k4mt9nOd6gWiC4Q
SgarQ4Ga7gGXhwe74SfQFuKZqmEQyjNQa+cy6HFA8HhWr99tQRe/Q+chF3MwmNtn4EeqKw7XKhMh
3ZVLwkx0JsftDpOD3agW43a14xkDIXcDi26YeF7EBFgvdGwquja1bw6rgQQr8V9EkDWAWDoTkQ97
rjKkhnH6JOFE6y9lopTFbe30he+sC4lCU6gwcLi6qovckTvreVpyPY9kNpgflKO+BmNu/3zuUT0u
nKMkaID30YOBLqJkkzwguQUZByr+IYYZJFUYNldVqiIsg9wG8kn2FDfJ+xJlEXWOS1fFYyppSKHW
JT0yL/Sk04zluUyp5V/f1Jgb2lyCmASW/sdeyMaKwty7tT87rC3kNS3aZx/RzKa5DUdSaQ2sfRtH
qdVl1Eazee1e1nHYWWNZFrpW6GsTeKlJGeaMHBkT8c+JBus/yVKRQCk5wW9CAz6xYCfYQPBxZQoW
QZHteEirlfmutJ/TVQfQaq5bH1DuglL22E3Gbr8XjU0L0V7/+nY5zgrBb6EUbftZNVVqib6/7ID+
/vlsglvQzh4v56JHDR6PPhVH0aOkV4tHeivrV0X5RZfpRnh6/lE9EceuPE5nPMzAq3ko1uYW8F+O
OJmnOYsODix1Y/DT7R5mJg8eHYwq0FVGsyXN3fvQ26NtX4rT3Qr1s3b5S+EOTRqad8UOJJ9Ko6zo
yycP0Zp5MXKWXwL/N0Ldj6qjhwCu4yxnURFk1j8OSf0mHhXuvxD/UrOVC+tJkqXFJjgDM2Os4jt1
QQJlI5oJy5NIZsgruKRNkmZlg1kj6+mF7RoQc+RmtvrkEDaQ0s/ohzZuu5PdvJ/f9SF3oOCE6hLl
HeeKFE8UGypJf1wEjzqR2Z302ZOqPws3BTnWY0ns6nTd1oqnDW9DgSfRxvRkPlxCXQ4VXGtqNvyg
xtE3tRfeTtQrYGmkqap5HcvrwK6FQXcgvzaelrLloTL8eCC4LNzx8AWQX0u4uKt8CdBbQk8rNit2
t8L6qbtTOBTemlq1uO9uGAFwWlEFT1uoe/02qxIuIqvfYoPfli9fhFwZ2BXMNq3LyYS7xEudUMDq
ZZ1v+VlGOr9YAZ3BOlv1V57szjf3+83Av0dweVas8rSLZj4RLfykYchsLFOYpHdWlcDjAAgV05tB
J6m0cSy29eimeiU7mylOLDfvHwtBxRL4UbaHoQ2VyNFOzl6YYn9/d5Vc5quFL1ltNN6zxNt/GCKO
cfGSO0NZYV4nVCNByO7p/7RqNrdbKLTpe3XzZUCZRwzwnkBKp4CkPYTifrHZZ6q2Sn8jo8hS542d
E0sUcm/u/MhHiuU2Gdkaf0g0F2IBWYOD+gsExj/hfInPbTpeqe/OXaX9BXziGClMCHxUu/DVjy9p
uzMAVcpuEyLnICuzCN8Nay61EOBMYnbz78AIpnhOLR4NwddBbnRONCwIaMdwASHa+RCkJBeozO+w
lSL8wNFN0w2voNk/z0A35Ks+0SqpsnHedH5Ljv2sr83y+V1aIJygZTGYDikYfV5osXKD0dpv2Ojo
4T0+qhtJ/vL0bdRTPTbU00XZ+XTpLDBHB/97eIWDYqNPByZZ3jcVk7fcOCH7xn1QohS93kF+yLnh
pQR9auUSbTTSd209q9RY+JO/X0cEfRv6+HbevTHWj4jALJ7uB1XjN1XFODyfoZxH50sr4NPwRfCp
T0vpjkpNY8GojNfAcvYksz9EmZ1Hv+iK5p9br8Q6TwinXlmR3Ql9CA/jH2hu6/xv5SjNpQAL5yCC
4ixbgOElug+3/9AOfGMOUkZdJMz5ETUQQDr3GgdMmNOL8klVk4MEjuS93NDKPbwHGTaqfFGmH56C
aDzUIVm9/FYOSs+Btu3qmsS7/VpmPhAntW91g++VG0edR565ukh8Q+xmFnhKNh/azj9ZDFy8WuAx
uH4JFG4nN7M/N2DXPqFvwDlI8zF0iFY8pIY6/gRqUXe8IXcI9QjgbDN/fixK0QiJFtK/eXKRQD3P
8ZVle8SFjaDT7FcPUxC8geina8psFE7kTvg33dpV4SwCcMlYdMAzin0EmBU2Ju/63aijAz8ErKTU
FRzaN8QhXJO9oL+2Zn8XSFYmkkBVPWbRdA3PNfw7J1eoL7UJqa9CJETyBm8FknwcmIZB1J++2mrz
FvnJaapzuLSI/p3QOWBXLFC9yeqoHJGiSICiWw3y6UsAkuNUThn6eO0hRMMxk8zhJFHTzUy72otA
U6Wbus/oOoQbLGXRMcwGTKJC798WyEPlVMJAWhOzYnYsDDG5N09Vy3fFpt+EoIclNlCKPgc0YNc7
NcYxBx/PppOHvpuI4GJxYcl3S7/MVcEdwmnHqyLkOIJR6Vvj4q8NkVrA7LnCxOsFJ6CyiqQYF20L
cIiVHZIHvljJXO50Aii+o6oxRtKUZLn2zg54DDxGAED+JyACZkADOJ1lQKg2W1eLCZHC8MbbAM3L
pDZMNrKT5EYJSnGaA86SoBROGns3GoE9t0uFJCaTb7eknNgGPZDZ7SXT1h2kM5p3NnjqmRV0aM+9
Rws+5NrixTIFc6pTMi0LEwOBtfkx2qe6ps0+z7XI2uSqJLux2NlGmT8hlJedAAGuoejicnfHCiBI
VXPfd/p3YnlsMWNhCBtLzYcK0u8ikbyjbfyeMPlzv411i8YpnAIqHrCCIirOqMLgB2VHn96vx8WM
GOU8a5zndO7klm37PplIgEMhc7epp51n8ER1lRrK9w1Z+HO7GKPrQlsjtndoJVPppfpisdYLm2D0
obWR3p69gOi2s1ziZZiHTXuG4aVdT/lLa8YCxvR4HQbAV7i8ytI9wQEXVzQuuy7Ugva7tPohqjnA
zumMZPCeq2DiaIC9ffQozJkC7ujIiz1RShEODRj145ELb/nx140FTQP2kpWvLC/dBNqYTpMoMlEC
d7MeLEjK5AZ/rlPOoDNkxuy7sOBNQ2X6LQX9xzhLZDxYmtqgL6bWJPEPP38FF7kyy9Cjz1OVzvhM
vY+//iABotvX9dqekAD9XX0VjEA13K9audcE6BFYHzyKpNWaofE0kxpD3tGKgnNl0OPQPp6/i6cS
JSQLv5zT7qFvxKExtdXe9witPFgu0LJD34+i/1sq5z7SIs+7dmOU5QPvmedYXo73RXVlekJ6GeeA
lRvLNCt9ACrfZpJey56u8gJBUV6o4JPUbggv/7zqXe1qjqePk1U160Vh6VND7bRkNssCDSl73SjO
m/ImPGc3Qp0BTw71oaUxt9Fq7UCjMXHSMh2w1KAzFeQJH7zl4mIXVODumd6AbzmZYqD+M/fpzulq
+h3KKIylM+uxKctbNje4uuAfo6M/0Co2Y3QVRR0xUG7tiV443tdHdHiGFWtzhzXA/F6OnDbXbckT
EEPqI7i+azjsk0Hh+6vCDu0IfHhUewO8dDYZGSlCdK5xPn/ePB4wzQl/99RW44PQpA0pqX6qdspc
b0QzxBfFwvzUfoyNlzxF9k/BDDlCgbmnQAAMT/uXfvIJMt6yVzx+jZQIYAN4Cfq5aQqtDL9fW4yA
54oYmRKjdaQnLEW4rq0dfjMvq9MGccCaZt3UYGIPY84JZB0NspUQPV0N92i+I8mHAAyp+r4t5ck+
ZHDna9aR0zhOt22EUCqssw3meij36QYn2pHyPxUh+tE0ApJFrBMR0FDXkivVR+vIkLxVDRsrAObn
4LmegvdxLOPteRdYC4kv7MP6aep9+cv+zrOBCJGxB+mhG59zOrrH6rMdWKCQhy+CFoVB7NcxogZE
NQ+C4T3A8LQwdx2f+RW+AJDtBK/OyDJwXY2+Jed7QIqdYcr2L101t0Ofhzarwn0GYZjHFO+IRFgf
Wq+6rxSSx/V2K0htQ+wriM5i9NBus9uLQwKHhl2Csc2x436TpLFurwVxxSqMHBVqq2RwyWThyluS
V0GG8zAUzfJMvSjcvniX+gmbzC9FPTjhpC91S193wgJNV5P+rCRp1St0m7JrrGt49K+24MWvW1cP
Qc1sedqq2VYSZ3Zsed+s/OK5Jby2wdV06PaPEMScgsq1WT4LPx8GpehivbFV8ep98dEOFbE+3EDA
IZ8eRulh7wogdvcyX+S0F9OLaYYCy4XRaRnHb3dChTc2cHJm8JevdEq6qMw+aYiOGj0+HKohNP8J
rNekvo+aUP4alKyfxtSfLRqusqkZAeKALdxCrZHxT5Zf11lpFSgP6uZMz8DejCgshgq2XvC6x90J
6eE8taq+g5iaZH4Il7QR2/ux+9WBNiiowoWRKUdOzNS0Z7xdP0RMKS2WSbmLg0XvJuYfjsRRzra4
3IGrhWEJall1IYG8+XlVsfrY+vqJdSyWpoPyk6oWqxnXCXgt1fxsiK0KTVHZrycuOiSHw95cyrp+
kSSWft9baZnPvP1Hnf0lzxSX7aa+JNw/Kk4peW2YmWL1xGGJUXj9O8A5q7hWIjDQHCmLGwGKRKQw
m5zdyZwjZTm8vjKGKq1KUgibGKnI+uCS75bM0gg/aAFBMgFgWGsHnxtQboKd7cmXw54mc9QuN+eD
ACFu6LxKp4UqoCOzsrsqbMqYZNWw3d5G4g06CBZqvQLlLfLuCq59Bi16bVMOzp5dpqzJbBqHin2t
X+MkmQPU5B6EAu1uzGctZ2V9Burg9lui1qjp+Jzl5Y6YrZDeb+QKbuiCUHKvEq1UgQV/benJvASX
bpShwOvRMlXMw/WNfgiQv7HFbLDg7KdZN7jbSop50yn/cBmuqnHbRgAhI7H1F4V80pu7C6QiISz1
O69xspjntwbTcp7JizcUrObhOIGJcFoUTLEoOy0EN6v4YqttpG4szQGov8xbKaa2poLC38CixS3L
WdbXGWtwAcycxus0yldrGrq2RA/MBiNYqbKuTML+Vp/fRr+KZ556W4T6tYMcHgiwhBl6xl6IAi22
OxRMoEuZ6u1gixYB2Eoi+GDbLaaxiEazlu8gjuJRM4pRsLuO2KZAlUIm3cHtL3wnBkfQJ3ZHweCK
NjmZ+kEfoBvvnTHlMVYtGkdqdq6A7kk2zqJd7Qkz2/RIUfUNfaJdGc7iSaEdZo+g/wNtsmGCXODw
hxigzbsR3ZolK799WlkuSBMA18TtQEd2iVkNXZgFiUAXNn2FCWSUuleoIiIKfdgsqTR8uROBrHev
iyFnMjGxwZ7EpDLUqAR/4T9XdcPu4hUuUpTcBPIYXLCfA3k1MR4bGfPinYWlLc2hL3/N94uJzdZY
b1PbLnOXUD1+UHh22wDpBQynV9z7KZwX8PsowIR+mEMah0memYhPsGb5/fStdAKjznosHeyBn0Nf
uVvNbMey93ytTUxZiSWbip47V3uDKKAtAFq4kCb1gTA6bRwwualofjCDTtxX6I2YMK/cvBhx6+be
AFZR2xXXONaXW4xUcMM3ALDlwQMdkt7s184rAOovp8zyF2PJOrW8DgbJs2Q0OLqhVpc2r9SAe3kT
cysw51jaSPwktHmvLfXa5HTYwSOX7emsbQQKv0LxjCk1ncv3Bay8TOeBKdxJhYeU1c6qv1ADEyoL
RfNzx0Kqzkmulz0bqjaNO2kK5+RxF7RerIfPV3YGrNrxd66xYAdw4W+fI7q1jHoMp278+4haA39w
fNQjibGvHpLhhiLbujQZn7FqZofbZO1fJiqELa6o5F30Bkwxd7eazgCUQsH38eSjd4Cw98UmvZJl
DlF4rqFKN8rUAvXynGayaQprzDMjiX34CSSktBDeckhgsONF7GJPf+AobR8tCwMXeb4ianxQc36n
5HOluDUqhv6B+ZHqkoOGju0EO30ALlh0SvSfWJHhT6owy3jwokuu1uRbXhB96ZKuzirr0kxF/Bdd
0NRPKp7o53nqQ3W+Z4VcG2Vmoa/QnIB7nWE0JYoLBpG9JmMrwp6dgwlGJ3+4SKjhTjPlA++ZraWU
twDXWID8ssFkt1Di7A198vK6dz5DGJiGidtLgq66LblGUtALXMKEfnYHQA91QdX/Wsj5htMW6jck
QqH0/mAJPqbPSFHowel3CYT1/60+Iv71ZUz7e7mAPRoiqtj+PHbo7zSDQm+xENlbLSoj9Q2tsZsM
IzOscBZITUoF9BCjE2fq7noS6vnj8JbJtOgTT0kx4YsKstnnuVi6iAJ44tFtBmbRdLXr92Sd2O9e
+xA+s4U+VwqDyvESO6djj0hkanMsnwxiy07z+Vw1AtsTF4bwpmHvmXL38jQeiiQMlJMzN7+Xe5QA
iCC11h7HUik2qs/c0QkmLd7YFajzPPSo2tBxZKcb+b0X0IeaLr+CZafE7JpG3gxuGNjZbh4anQRr
bYxkaxvOOa2SRwOH2AyYBI6RMJ9OT92wgZgtcnZepf3syF/Ssa6yWQNY73zLvlvna1F/B0+j4k2b
e10Oh7JbAuUmUSxRkVorKcshHmImuy/aoMRzM2JiXh3cbJBLshkkcAN6pQR67HeiMigfCViJgR3e
pP6HfN3RXdYWxc23QJlW5bqWf1yo+Vq0CTAR71adqxIJLUUy3ubZ20c2i4tyqDgMOD00rydmrPYm
euSzz7Qp4GQUCka5Zvjp6XcIKVkJIoLwqDCj2e+Qy873sC2QGKS4klRk4hFMqzJvQ+Wz9gjZX7CH
kQblfGYCBJmREA8kfVkiREBf3tZRqKMNKaVUAxt0ZVkDJPCqJFh/7V5qS5hG6Qjer9t9Fk0OA9jz
ztLZyeM/FVobpIhP5IcCYLeNKRr1cOJ7fGHp09Q215HB5VBZMvwlVrUkc5wu9MXBzx42VfAw2YCb
WynO/ec5UovgiOMIQDrznlVcglzmpP1bcQRz6ygFJRHdPh1JZoNKouCXx1YVJ5seNc7OdyFUfQpB
j50y2IfAp+xXQEr0CN16Br9L73ukmwIzlfMtcqc/qQ+IvrMY9VKtWrMCNH7Thh2IFXCyuiUGdMWs
u7EiUBtvy5ic6hKe6mBFDpfyvFiftTz83PEVLT/kxemoUZMKi6MT/juSRRa6xhCalMHcgYsAqRdi
AOhyZnOStrngG7vEXFHEgXP/0SAGriCLidfJDImuFmPsBQWP82j8tX9ra9LhqBBcWMtYztwMYyIV
avygbybz+gK7Wpx+/Lnruebtg1zVh+v8kivvHNrvlkwCssSmK3xlqNXlxD9aTns5WbF2fjSH5PpJ
Cb1hwxplZN4uB4Sj+8CvFsOQhBmT9LNTQVYCUC3W4wlc+XV48UryIY4FvU2UbEb2aqF9ZugC1RLT
kjSdAYipVqM2hktv9adDg8gKSbfm0Oe/TJTpQ1Z73F9HlSEIQahaUxWg/Nc2ugAXpcNqjk4aT22a
nTlFTyR09rfEz7Ns0hF1F/L8JTSYVuuIilnTRutLso6AcVxvaF/z+TDWdnR/GZshBnqc8rpxgF1m
rM030c+zEIpAQdEcjmiEpj5tK0Gb/rD38VGypY/eKdFEaCRtiC5K8Id0hx/X6WdhYJgIn53ywthW
uhgvuHo+ggUnPIZ2SccwBuWh9nzYl6uhnuYhkUuUZn9ICO7KKTnj790zu1aJ/MllB/hpJParOcBD
VQ5J1erke/J7SxUvZW/4NzM0Kjx8i5ZTt1JqieqP+ng6KzsF8RmW6hTR3lzJ6blkhokL7NsHpETL
IRtZIVzy0C83D+eme3S3cBEKsGkclKEMjPeZNuwAmIx67sGVpDns58XYrIsl17nvJ3nzbKxjobFf
dEgmHWLfVoDGRxxXJpqy5lEm2GCticXPncaNymbhBB/UBUaZiM9AMdmqiLimfyO/9NvXe48g2SiE
eEly/Ss1ENkIBVeW9f7fUT4RW567kYaW8dB+mzX3zHstEBnplTj8OST59DC6PhoxdUzuB6WvJTAj
ZES86OwqaNcr3+CpPZJBoV2Np4qh3yNEUrINKRTHsgnoRow0ausbdZGzwthDOpa/NXcSufb8ep6P
DNBsLSaMiwCHWYLPs105SPAPUI5rJ7JjDIVD+Y2ifvP8e0EemIP9SGZyXq4405zOhZLiwUaAw3SN
x4PFYzOKZLj8fI6FRuySyz/eIJNAEfJFV0bhs+soyxjYzvdG9DpBCYb2jp7N+0EJGml75VeU0mu5
3z3E1tpovKlhHOA1Au98WYviDzTnPkDfNLwfCALsjcTJz6A4rwFMLsyRzWyO4sU9mQdLjmpJUUEY
KzNidpvuviHlk3cAYWTbivugkZD+c++Ers60gsc/qYKD+zBKnXdrda45rprz/yduzx0nZafirK9x
rYuqD0AdF02UFoX/rjK+OaKs91GETWbzCRanUmnZfnSWwCtFLxT5NXhy0rGn/1iQIfPbPZ+UQQ5F
w9DIacxLURXY7Z6o1ygITvyDTR7lgksvXurD19ngLgB1/r4AVpZyn7L1dnrU670BpGt0ZWLayP+1
ZidBN1jA3K9ZpTNjLJpjbtHbzSoQLMwnHaZX2cxd/3YsV/4KfXM8UqgH/Iuwvpg7E+sz17K8uP7T
5Dk24Dc8EV1q3jq9eGLKS/XKPQ8gv6huMXlMG344WDjU73LMXyWpiZxpzQFfnG1fZMxVB+9rkXTY
+pdJgK5sXUHJ1qR0OENwIpmhO0hdHOC8fX7wwCKtdgfyxfbIizxVCdM3x3+EVshtnyNclpW9NH8Z
F+nUu7BKtctlSTdPbIjCq62WkC7gAa+3eRYryA5ArggGkQXAH1cMrC2X7SCROGs3zFWTBxZf7DRS
/BF6FX5MKlSqfDxx3780JBmIJTJm5m+Dgx9bHbTTSqwSnCAMUteIeUIOnj+u2VZUoo5NQxVQu27B
uRyrJ53IebYR5z3iPeCP8kNpw5jK3GNWohj05SQkr7RzEbLDDIXK9tyEtsOcJMS9iVE3JCbkQ+nc
5ev08HQz2eIgL248+Em5TnIS+fa2bFm3Ofqnjgx9v9qsxKzXMMVZ1e7WpLjFPAarDzhlt5Olp5kn
w/rEIgF/9ivN1aUXE8Y4gQyxW0fQqqVFdUWpkZH5QLw54s304VmgTJsTCkzLgwBkbXeC5/u4Idzn
iOW/fCyTLPBXntXDN29I9IuOX3fu9Z53uhfOc2dsX2uDdwhAavdY128sR4ElJnvilUbakcrrJGC3
XyBcPeX2Vpvr9KOHCSWFtsPpvXR+Wf9B9IY+c3/XKCCK1pxDhXvhf03rHJcQM0BrJmC6GXU3SdvN
nr9fNqwDWj4NgdsZgHpJAjCyVJV3e5iqQ38ugGDOiDpMV0IQ2cyE8qohb3RMU2PZtK8QQGfJHf8U
YGGklyJ5Oq3C0y+8bazGX9v5cgGARE/9gmsGtBoKGkjXyFtw0HBEZd8a81w3ewFZ713zbxRi2ycZ
TQJE7Nht+KPpyutbBO1FsD2acBusgTbkEyySN1aHop2e7ExOELxu+7ul9BTRAiJt0n8pahY9ydZe
8uW02Pns/b1Syv6Utl0UQzPyldHyX5aXI2lFkM+uVFnlPBgwKQF/cGnAdU7PXruwobrG8gg/opWk
3RIdXIng1631pdcCtrhSeefVqJnImFwWWE7VCTVuJxq+o5d31K16g8UKN6BJA9MpPgKGaG+N5I4h
mgYLCUYdPMhfNMx2MLEQ8/6KIsfAhajuUUEHjAc90KEAxdjZ+topo5jrs1QieSNmvZGMvhFEltLc
zE/S8hmP6+1J3ANcYYNGMJdFdg1hZeXoqnRoBGB+S/qM+g34CHk5/jeY6hNZ/mxwWitfN68HVPz3
WVcS+yMwQ0989zTby7Q65NX+0VijjIvy+OZLdcWAPXVCd5xzOS1TgqB4yZE7FbIsoMkgSlUpVLP4
hKS7frrxQgPsTz6APdwfrVvUuSNkM66Ch++RzmxJVWL1OTtkphNmQpNKQzFwA9KJH9qfVW0ajM5s
PhdBUHd3/OXR4igfqwjFSe3k2CcJm/mgycUTLycfOuvIzdn4PY4JbeE5u4aEsO5GkPUKpLE0x4Ph
7bGsZsuOkwSfoWykRn5x+tWkbd+AxQ4BbwcNb/byA2vMsUdaNp1oNbJEkaINflinu3k9puwdNZLz
A8O2uxZRitn8a9dbSnUkh50DlLSTlelTCWal5mRHEQyPSiccrCuaBBN1PNGcFU8yz80HGK4ybWGa
J02WJqICKaWNTmyjltFTwMnDoYhsqPdY8Rn4+SPh4bRYE3adVqT09RzL06PiZkUezrQleY4HDHD3
imkT78cOfypkeDFVbebYv6TpPTuExL8/VXF4CS06nT/6IVQAnbqe+cstrFZCNPm2DLqNcLBuYVaJ
a9TosAObV3E/zPBz/OK4bYAn+09LCG3c+hE8pXcrBpGEdzBdbJGIEldFj8qEdcytS0IqlrKfsKdH
3B+b3lEVLeu46h6bQR67W8mrnTS3Gs9snx0Aher6JS2vcKiltLWlsOtcJZkHMN1FnWn64kf8KnwO
7HiMbp9x4U3drWUOgNUlQToIk+rkbOQl2ZdwgV2xUJhLBmjuPUVetU3odkd3YmIxc2D40I+76iPm
wcFUwW97WnGTrB52q1Wzm7SeNFHuAjAEZ4kiQw3pvThYLrwimT+e/h5q95bsvWW+6ZplDNZPn0Ev
WM8wYy8aEtHoA2BxeKYzXjt87LBuvTEIrQz4P2kgZabboVRQ1bm6EGBB2BoLRg4srUCNdiKKgh88
PXdse1pVBJzyHONvYChyvLM0dcbNovDncqyFUno5qJk25puRor76ns7IZxUIGiRAzoDa2Kngk48F
/1GoAGtF36qrx3HPsFWOHn1F6v3Pn5ZLh2puN8dCr+dBBbqoA/fR2LWvxIexRB6kMZt9HAbm66zi
luoE6NjrcpOOBgd/34DYBWQdmCElWrthAYWDNdtyQ2LfSt3DCu4aRxCa1DRuHVfrYeoW8cITfeQK
C00XLvWP7kq+SRe1HdN0/4PquI+tuuVvKOzRROvqUrP+7PZnP0IyLczgtlEb9MjTOTfxW1YBDxxL
/bdyvHk8Nq/vK1ACPNEMQqj6lgeKKw3cAVN2IPAlI50GFFour4btjBebSgmhMx3JVw3dPgBBwcDq
Fx/c6quSxPAfwcGACHjtI5s3QwZnT7Ahdz/SjwQ48MkwdhJ6e7T2x6D7MCAOKe8Zcv2ZNdN+monI
REwbZGtIoIe8zT/lMt3jWy2RtDkis77bwn4j4MgucLYG+h2cwuvLCPg047/YcaJNNrn1iEKQxymj
iWeVfqoVVnr18plCFIF4YhODaqPiYqPqYo7MZpkKEPqPagVQABKSWwj/0mmM9vQeVQisPixpi4Bn
eO3PfLsh4lNfuen8FM1h3Nbhop77ClXSFeaIe0hLo07+D39dmE8qUf/V/8Ojl90xZRiCQ7M2JSIi
mGrZATe5LM2p1C3mC7roEPZNRb6IrPrsGgofvx+A32D44ZJ2TNFd2SP+5RysP4o7pLjtF6h/K8px
8GBXEbNpeRCkVe6sI2xNODjtLoYL6dpo4kAIbn1KRWVs9A4+sr54HtYA2A0chdVsToQylzNMl63p
OIaPiYZumEgVR3hpKWvHzr20sjwzU0lDw3xBoECDaRS2qBbKiDGwujCN/IiPBh/oAlPrdb3eGKZl
J+E/9qAlGVMd8TwXOw69+/WbdxfTQ6pHaQO9DxCo3OvnhutZX/9jsRJX/G6KGobEt41QJ7gRKFFV
76xSAgeXzDgnw7xnv/FZiNRn1XZZt6BT53EEaMrSfPfulQYiebMaOtlqO7Jc00MUPgReG1GCzLpl
rZn8PaEyplbiJwbLq55/qjlqD1Lb0is6j0SJ8NybzQmso8itY2IEYZ+89jzLIdeckKhISBu3688H
2GynsWKvvRtRxKzve2qAlaZE5/Mn0pG18NrLTCkM1cQVFprDQpuw5TZOK4YRLT6FoRaWxesn5h3n
JqpyAuF5VBeS2+/31MDw8waPGmfpoQq22Z/BpPCf5lUI3LoSAt6Bm0TIIe6349iZ4wD/vq5XWu3D
7BYrPGhFrBDeDniiqGaLPIhCfeQKajdiHaPqxyk5dbIgoC1EKFEie+nYeXFOoLwBjRuC5HJiyxak
jH7ns178+/Rz0BjJp47mUxi4dMaNWv1VH/WWzJN7Poh2zHRu8a9ZALsyW+FX1kYL7jnNAF5k700L
fJ/O1DYr0dQOrzU6dwYd87T34VSs5yrU4yM3a9V6q1MijYUchQP42FMvrxHpjU/rXBlhXPuWfvOG
S8d50DgF87uZ8GWQBBhkbhCp/IgxEdPFQ3Qpcty2Gft/2u7JPZYA5JQ85wjtYrbIXDIrB7QWoc9D
5B7tNw+pXjHNJtMt7grcvvROJ0a8e/jv9dSfrs5hRfVQWwuDvjNI10l2pGahO8HVZh/uiHGSa/Mn
KszAWhkRf2Kap9HwvqtlSd9m9yQkxBMgHbfr1hwAt9t0n5H2OBfpYAnGfk7G4+aJYMwH96i9uCvP
0qXwhJckahymxGaN2WIusoUY6B5/rgA1qhxA4pmqqtgURjqESGrzJ5H/Wlh6IoA5aBw9EuyjR3Aq
tiL8UB+VlOzEtXgN5ZAbHLdJiY3vbLrPRMJa2//9kAWbf6MJ7m/7Orh0Q730w6paGcLeekBQjdI0
zzUm7be1P5jVCLWOTMgMP6RfZ5H9zrYLmYzSqz6smCkDNJryOK1UkMqrYxKfH6j7jApvjdoJ1Gyb
g2FyqVuwAxMIrG4ng2gCF5CumD39WF6ijMEhd38sjtFj8jRsqcQJrz2/BpSfAyKtJ8SWL+SawUje
P/r3IbmwyRTpUv4bz7eOqzrmL6UZ1LyRUIU2s4LtCj6ZiDYUFuXCwDGWi27IejH3pUTY7mYozaCj
FWE56unDx/wykqk0gSGdCP65xYBLaPVxI5K4BvXI5vy6J/wV2pJKo+jmAyswJW1IFeExTkLo5iGV
ACBKAZKBdm68G9L0TiL07Ufvaj6TT4cMSkp3pw/LD7NYhB/q56+Tz7cMqvfntggf7acIYD1+wkys
jTfVehXRQvTPEeQxjgzX443wf7/C/f6TqqSCHtaXwDS6wMDBkQWs9dllTio0NmTYH15eMEnQgdn+
DaqHa6IOLrlLr3DjAvyS/XM/BLKqFcDKm1GAuG3V7SXsEvwT/wW9I7sgcNni+LKqV+3eB8ZxCk83
/bgQBtJ2ukGqunQm972PRTPIAoIiUvBErMqzgjGJs5ehlLVAMPJrkgCyalCphhnOZ6Kmzh3gDLwe
AgVQBh1Et6THmc8QsZ8fNWmXuiyjRnqlv6jqy5LzONjNU5NYGBWNsXALvOK/OoNjerFu3vDnxSfp
t6Tud3NL3TcK5Xx6XhFnXyL/kXawwGOvFCIAxaX4zMsBOfDGe8NJRGdvqCPHWaRS8Ij7HNMkteb/
TEpPI/haOqsKq8+RU4rJqDOXP5zOWdKtjXG4VqLfvD3VVdhOBNCrQfHsmYqDZ09nUE98V93xOapW
n7JwVQAhmYWT+uwLvy3cTIpfp6wxLUTmArksuV8Pl0jiyU1QEFcp2zaL1wH3QgbrEKe8LE66IT0k
Jxgb4T6RM9P3EyJOlawhdsn8mknF+HU3D/LWJI+ce/u83KmhoACkRs2zdEJ3HLwU/X449W99zKR2
IFdwLlhKb5Ha62V+/gflRxWC8YnFOnl4N5CVUQFQ/Ue32RqnQee3OTPLN66kFDrkAFYL7JJAhMNP
ExajmWVQgeHpJ91YmCxcP11iye6xa6cXCAvms1Nd6Vy+KAEB0+ViX9A3bvRF97jq6VmrD7GGy5mA
eVqmSU55OBD62OitOknB5D7FbcXtW/aFMhLhYBkhR8akFbkYwUlPyTSRa1b1hePC8n3KL10WRwNI
vtrSMgjBLDvLw+aZXOfAf8CfIoLFEMSq0iqKhr1k1dw5kIL1+aXd8+ktZtmSDSMufeK6e8+z1ttI
AUcfMRe6upvxIIVw4jBhyWEC3gxcnYQHx8kdop7fDG6gBZEKrfuVuEi/cFJEqWerMW/Jw3cmGbXL
oCiQhRmn0nBljNTMecoNM6mepMRYKk6WZ4tQpHzHyKverwytlpPd9WiDaY1DTxpi3Oz2Hpe8Vz29
eG1nXVg9PCvO5s8imw7lYgvVPh3yxvVtHGBAWS/buvUa8VYwMBg+Sn8+BI1XSv8LOznrbVlZ27nA
e4ahqWUtG/63nFxjBR7JrS6Sk5cZjqFlny+friH4/bi5XQ7rqJpYFORXZQPeeuGUl6Gfbbbg/C1k
+jNkh4UMnljbCmeavggKrN1AthVR46qJH2jxQp9FYoVRST9JTpy0YPtbiZsRfpqzo1QSHkUIBkuO
ZtR0l/ZRLvct+lrSQpxqDCelbRana53PkRQkIjIaHxqkiVawzFd3nqZfuOAA9hxrpBAe+c1mHUfU
tkA0aqXv6pWOlY/660lhFFRkhBLGqB6LEyE7IWO2Ag1pzuSBFaiO/uCWGkPEVbCPbImRhyJ6CHsl
ErNvsGsililtR/EcDI7I1JukGOcn2qt+WKK+BXuJO6vI1OfBoilmU/H2sGJsyXkJ/YZags4wdpeQ
1tYAop3ZAQKheMe28zSYQXcanp6Md3ezDaMba7W950ThvXVlUre9N7VQzoR75is/TIJa2DwMscew
KNuEVOPevnsfe5y+9FifTneHcDXKgYLLEWzCynQls0t64csFU4gjopIuMc3nqGgEINjuTxuyz3Lv
/++7WGlbAAry1/9D5+ujC7/pxi18mbJ5NVB0PGpm9QpSWco8Vg4bS0AYEaAGcLr9fc79F58W65lu
2UuYVTK3AsdAVLa2s19bT4jKBe+oEyNnrEZ8yN/NFWOA4n7iDBKRkXJYkUxw5REv0vnYaRcGTi72
HyQ6SitBRLEMwKy08XMxReoPNdMT9xNUAHfIv4qfB65BpnvmtBRIjCM35hbrTI+lXyKXwyO6e3Yd
IlZoNFx1GPlDgyzJiTJAP0lr4FUE2biwxhnpOas7wBzlLAnSRUCjD1EmT24rDV4X8w4QAubkEyxQ
sPW/d6QIpc/188rh+UE21lMDkV6Ugl/mas7rCHPcQz0+0HdINYN+5wgyxv/ghu3pAlk+P5CVGwWn
fm17nXK3QZ0iMj3Et5jHSpYgpO6F3l081KnhXDosudn2h27DQGrXXzwTra1SrTIwNHN2X/AVUfTQ
plMsTMGnnwD2Msnd56kkErnoM/knMSdW718L7TylMUHPnQ01ZI6hXQ5EVGRfy2Z3RS9zRu7mJ4v8
JKY5M3UD/xMbsxiPNvdWWBgCoYjP70NTnH4AVI7n0Dk4fac1xtQFz6R6axttqQGqryukBguPHl9a
WCzhYXLwAsvBeaIqsA71PZIfmoNQasqCAeHDXb/FVG+17ejSNBgLqmL959IvptKkA/gv7UzAch0p
8YWvupdGAZnPILceM14KCH0ScdNhPKzwGBrfPlU/gfc/GTs98bS6IcAL7q52gzlqQNGnVtCtdvyy
7iXrA/Nm4mrfzBQHIRDxnJ7z+MIRusRr6Y0ZCXNTI0Qc8cek3V6YYw5YznPPID2KFiqQyJrVo4eo
6tL7Cgao2QGVy3LXweGE++MsrIiGkIIYGv7ggUZgN/cNb0IcuCDiG0Rm0KryLsghONWTsEo50YAQ
UFpZjUcXivhTURGm4CtC0Xj4Y+AKf1k7pGDVMsV0YJnNXRl8+TwL6mYo+kjBCBWydpSpqmVhnPfV
4OJ1V9ac2z5BQEFSaEoOpwgbZljAVe39unTMs32QqYmfIiBm97zhB5FNSab6kiG6JLagAP8worwi
zK33VkigND7E+MmlCiPGTege5UR6ua5SbEysn0trAPLLR0JWgk3PTKJRGu/cem1NXrDpUf7cWTki
V3wkdZDYXOVFVPykRB+deOnurGHqQCfEx3dqRCf47I95WqdrS5hTEx+mCIEA/ct30etyXIcOUQWa
X3nFmYJbJcPShMIkYtbpa+fQi4t0vacYr/aL1w+6drzS2615F3V3v5IEfOpAl39UpopCcjZbXLhT
pPwBn8VZyYkfm3jimlUXmgXRlI4a/DY74fbSUDfNmqpZ9p8FNgQq+BBGNaorjAeZUOfvS6rOG6oz
3aUpihk73m9wtEyM7lLaJMQdKb6qdfasakhW4D3kWque9rbJYr7dKU/aNVEart93vCAcPg1xmKcR
zKgFFggdMqIbJ2KSKNfFCqeyVYmGHOV0NpRbfUHkkwaImDEGUShUARvCTZJlSwu+YbMtNh9WzRjk
mQsOWtZPnXB0zmfSOKIcnamdHcDSGeNntnvJquj25SFECa25HaJ6JU+MCxOW179I/piXVCETPK9m
L0KJWMTqdYdMzUvE+V2VlvztbbISzRHiyI2+RNkEsPySRwIOWoTFYkG5i5cYLS++F526xe5RjF9u
BN2KGlHQc//1lcZRMP0k+lN4Ro2W+a3O/XF+MFnNG+MZPFJYTf6tUAFWa3XqdiuwwMBV4dXxwg9D
dZ0rRK39JOpyK+Gg3DP/GPByE8cF++BkoqVprb9T54qlsZB3+tN87lpFEq/IGet3S2h4r2+zV/Co
2w4ZyFqOQ9doB4X0y6Fp+TE0o5V+O+Yh24LySkR6x3tx8Fgfxh3OzTxCY4T0VQ8FVUTES8ZTiMiw
cU4V1k9jMidHSqyVsvUyIv7lb7wNCoXZmv9nm9gbxj1QA/3jHni1Z9F4Wkj9UKpHob8rfU86X5l1
62i6udeynptEWI7cYQbvKjJbBuCgecijmlzP7LsYLorT8tXQEOXSQP5R3uwSy25DxJNvSEchsxxA
2ejYzdB7u6k3aNYEUjQTZ4gAE06BGcNtabsPrMfvC0M1TUBidtig6hnDlMi7muP0mibX3v8ZgirI
cQPbJbs06esCJ9pDnvJPJwsKcSxuczPgn2eT9fPKD4/hM6ZDQ6fSLJPJowwsBgvvmo4m7ILR+fyP
0T+TEH9iym1XElKN/2xVq7T58yYRdc/HlRENicFjUa1+FTAMNT2KqKH0M3qyLn3zBcNz8dtbgmUp
TUwrOiOQsRvWfiPOu03TaqaXUHeL2fyihj+RW4hBmJNVorlwnHsdae2j+BioHPXJH8XlO+Hb2WLR
mxw5bDVMqvaNooa7wh+LpgKvslrgI/FKZvQJsqTvvqkS19Cz6Kxdj/NL20oqqc4w8CSvJX0HSH5p
A9BceVDS9TqufhpeaEeEuQe6LrtF4b3ndBdNXQlgP9t3jqB15+/pPae+oKKfgOlmBdJNv++0/4X8
lhGtg8r/bcypyCbxhwCwEHBr103Lw2/74Ghw7B6oYcOGSjzYxyQm731zIgemqAq8rnEy4jk3lzs5
NaeVONJE8KTEpcvN7I7HmGd08fBEVqPiUZeU1u0wpxhAhBUoKupKZGB1rmLtST/ux/Xu06JIwfKt
fpHq/jjByCKUkSaADuyiKZtfe2LdKsJU2FcmaAalSxLPu7Cl4Fu/bazYvZ+A1NdnzeonIMpx8W7Z
Pgmm7DVD6hnSAVrDgI7dEbdri93n+NaEmfazjwZeiy2eTmFZpJlqNDTm6ZHN174YPwpiRgO0nTAA
AjWhWXAKQVh7P1Ubr3s+8iQy5lG0wipSCbTN6hnQaW641MnGCkv1rPWfOX0iUK0jc4Z2xuyi/cRR
y6wpukdGRkAItuZhMO8IncXnWPsrPJdCluz9L5nKa46IN6vHzzzf6/9vTPatBWRgpN+1EjF0W3gb
vjShNeMJuNHfaCzXxd7M4xqZ2gotZnuuQOeBTxon/IqE+w+QGKfKHTWvmiAnWWsmv6D5VhIdTny2
LL9vH1/qqtu9HfpuptpXEGYGzA7HzHmWc+foICtpvNTZfzFjv26HwJRGr5gE+qcNHvrcyd7W2bFA
2J1HCGkTYeByfID6uDlbr+U+srVF2q2WLmJLEIP5/jJAcJuiNjfjUKchTAGtFGeyHXZqBHIC3eZz
Y/BFoeBv53AHsaQh6K5Z1WeuoIqaCcvwKldXWtGsy6Fs8xiEDEI7clsJuPZDD9goO2WvpOQtOayC
p/ELEqZ+nw0Ct96hmlSjmWJaPuzekco4CCXL/NdNr1C/mmlv2QjhDujK7Zucq+V7RESa8J1A3I/Q
NsegzZBcOGu9m10QuFjZRwnvMp8hfieFCR1hz4QjzPQ8dpOOux0fOyf8VeRCUxuhvJRTP77Z/Kg3
GsZVbNA+Qyp2/CuXITU0av8VcTYUuHHYvEwpxeHmrfwIBOHs0NVjtxVpw0Z3ZinVByG/5+LzGcTG
USre2jlHTWSPmbC88x37c46EyOyKtjOiJbCcZzISIy1wSlmDsl5SKXd6tWfkgltMov2XW1QN5T48
fCrWfSiBmmSRnNs7kS1cfDfOFbp4FLc2+3ovb54Uvz3CBNUNuuor8qO1F1hXXsHTm3Sxtt8/JODK
1bD1UQgCpz+IsPXHHZ/ah+H33rtx7eC6xCLa7uwCiydhnEAcqRNJ4MTcD14Bzd3zqRJHDRypw5vh
wtldXH3AVkcYasjrgqLE97IdLPIRwnn8D2XzuuGy03kI+gQRIFZjYoWq6jYKKgSPGcNaP1J6yRUX
Ud3W9b5mIX06BjdX+d/RoDH7Yz2/Ju9LOp/0YUq0ImOycicLG5x3aLqdx9OEFaTq3kqX5U7N1UQf
uX55+XkO69F2sqhE8edvqfEJ+BYqxUIgLlGoSOgyS44+fRTKyNCtdPWHI0PAyi2UIZNvb+KQ/G1w
BlSYlH4oEeKrdJiDf4hfgEBW8n/9qiyrFCt2YAXWOat/Bz1M6wF8bdVHnH+qVL9/oTZbIknIfsaH
aJ/ng2dlh2K1yI3bu7YT6qjyrDjASMIktzDlNY7mxBbm8kbRuEn+GbfKiJQ6atw7aZQXqFE+Nrnj
3slEFWKVdNwxfCFAoPhxoL5mgxeZQOqrPhAboq4POmtPc08laD5YqHOlnzaqZ+ZXqd1uxmQuFiis
tplTao810IgDP97gi9OPD4y88H5SPANkvL0Z66U3Gotfb5eJ69qQpZdJFlj4tijLLyP7BdWkXmAY
xUYICKj6FQI2c4qnYiWex/BxhXvSVec4VNYzXV5TxDAMY9TI097ilgAr5cGmmCs63Vq3fkfZv1m3
PSe6KpaFkhe7wbg4913dxmXlGg4Y66+8p0ku533wk7Kzi12HdUb79UH3vr0LMwZVv4ZIcWRrILC+
his/2UuNU3yOg4+CRLmGPGraNtuNPiioaRazAGwEIF/XArpY9rSOUza0PmBiDlqU8A7baSBPJdfj
Hd8/zThx5Rb6MYHrJTDNEDwwkFoN/i3qos8F5hsAeNw6mYX2nhkyWECQjeVwbzqAcDrVz900sFm+
RKr8eg4KFF8glFbWJmxm64YspIveOMrSl5Z2raCg53SoaOpuBzQmpV+3NgFDiXY3Ov35CefUowSZ
juzuvnYNC+U44uHO/o74PDESTaN+Yf+2ItOVzkBVI7NintLh0jnEOI90ltOt+5XyIOy65CJzmOho
BhJ9xSm0ZXtcAxmcqklWNU7atbt0W4i0M3DpOuRLHoINeZxClByQGBGx8rEatjpnbwlmKWROB/pR
yFMn0+RQKj24fCDrO17WacoX53MFJ1l2QfFWZeFJQjCR2Iw+D4g0rCvHIuNxWYaxhen+NCSK7kl1
kvBHbMIsp5+r5SFD5AKPjnvtzjoQzgzfu93eS0Xne2vgA/ysy+66WA5Ghrfobm90y4fG6GpFe7Xh
GRRHoRoWJgvG29oeaZjM0JNdGKA2zi1FcXC/PmiZDVFk+xcdg6gIcl828shguiHr3mq9OGnf+FHW
KDRsweabY2UfofN4+SJofJoBy1UJb4N2kf5doLAPBSz/t+DbRrMlZ5dvd1on77nA5/JYOKu5cZr4
UgMUC5zqQLTgtW+Oukft2JVIuAJVZQmp2OsVxb4xmVZ0fHbxfyyNEuH0NOYFf08FppvMJlCaRjD2
MMlDXg9oVNhCP6Yz+Hkdkrom0fTuDbpOy1RWm7+ebDv6pSiP0p0U/sCsZrgip8vd6tR5rp5EAXeS
rN1hEnSKin6arhBtoKNdPzoKbz8ahglYqYxmzjVm1pXEKmOEOhcRpuBq/L/x7kOtdWsBJRLBrBUZ
VWIgWHfH8Y6FOFFXnXjM2pz1NX5aw1cWbjQh327r1ROCyC+jFFwinOsZqi0OKCzksziowkKJFfg8
byvzZDQkKHZRQuZdFktTzlpSTok32K2FY9BV4fue3rSFHR7V3xB2edZKAWR96onM3eMjm3jTX1Mv
EL3k1No7GDSUDplQu2OrTQ60X+LfNAdZkq0st+HESFqRKhPUccT2t/lZDPfEYdCeaqgx3+dpc7rq
4Wiw22PW9uRu3gUDkMJgyZaZDFhPnIiIuw5zCVKSRL8NczgOcyttKNG4fx+kJtPjQDX/ex2OczDh
Jw1pMxgk4fJdQBGXhy+QeQuMDoeLRMdg3e3EG0+wpDNNHhdUm9UziMWA618YrmMkg5Y0fZo2etQm
eH1IIZXV3YSAXDhcjbEtJK3UMUbefZjdwpRw0SEffPxlUobihn449c747Bw/3yYuaT+V63OHbqow
DGvhI9fapXpy/ajNZ7ok8zPwEK+rDH/w0IgmRl2SRMWLgCEwAp0Z3HKtQ/Y2B3vyYgeUQff5UaQi
m2fZmdRsR0WrZjT4GQLpavHHDsxQ4cCDvO3v842qW3+Yeh1kxL87qumwk9mt2PibL3rCEyrDHud4
iv633pKRK364I0L+F3G7IInWMwrb0BfIY1CirExuaOnns0th/QrbEbua+/BolrAUZqCWvhrpi3i7
WPBwb80NpN1FB3Ot+jVIDpmD6bQWFeVCGgLtJIaQ1MB91BVK7BMWvcTD5YLGguKJZbX5i8k5A8HV
jpCy71JxcLmO9oE7KpgPpndu3urX35QePPbYRc5JQV1tRvz4KwLlH1JOQl2RBw+T8a5YGkZOxmJW
euZTUoz53LDUmQCgA+ZlhA4Q6yydUSeLZ86fsV3vfmwl+ks/HmW33OLUG4Wi8qdexIblo6ygnK5B
oWYYDpeWiReAe1QSYgGPxMRHU6s2NOXDYq2EJoCO7DvT05BZlAmU3XsyOwUtWZMz8L4B1f8QX6DY
AVoSH3lpNrezzrPkbyDT5fjP7iAM1rqVim7rrQwdt07H3Qh+xgPp9o0F4kp95oQLk2JtQ9KPJuTI
AZCOoyR3cVVbP8zMrJJQ4JcdoYqhe2nCvyiBmiWUu6WyGgFFGKuqhaX7dn0pbVNHccGmw9e6ss7A
10nqz4xyEtoTlx3O2p6aM3n3WbX45efeX3FbwjOVmtxU14JjC5BF5yK0iJAaOgHXt8CCwTcno3Ad
3y2mfBWv+W42nAfp9u/cOAA7KSfAmLuykaGi3pziuN0=
`protect end_protected
