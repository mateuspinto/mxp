��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���� ��8�F���GāV���sD2�Ysh��"�������f{f'0R`� 53���j���u���q��ZUh��)���B����e.O��}J�/� �\xn�ZP.mwl�B�k�-�%�2�� ���H0o�.�9w��!��j��'�8���H8q6����O��!�lf+����e�DD�s���U*}��m�:� [�F��N��K�,�� ����A�bMmGܹ��94̿�7�R}�g���^�煷#�4[��>�K�Lڿ ��l-��{��A�I*�	�(�rU��_���@�,i#x����@wH�+���čA�lP�.���,�(b�z�ho��u"�XԌ�!^ء/�7�v����rURem�ytG���vA��>$d��JA���o��h�(�y{����`�5��Bj�-��D��N�އ
�~�e���A��=��8s.�	�{sfE�[���zV����Z�"1�8��E�OZǙc[ ���|�[��O���?'�R~~��Է�	Ե%�Φ����yΓK���ok�0*5�v�v�/�\�`Y�e�eeXl�Jv�5Lr����f\��Go9�%|	�=*N��q����|!p>�LW��l��'J秦�^']�U�q�xОA��>Vvyڞ�Ճ!�r`�.߀�(����i){�N+>�<�D�a�&7-�l�x�I�l0E���w�I�Vr�q��}u��!�������V��ա�þ�}\��L-��V�b�ywT��k$�{Շ�m\l�f��
�v9� =;5��r��w�5��(�q�ʟ%"G�{.�.�p���$1�m��0d�q� ��G�����	_ �t�E�J��e+cUe��n����+���۽� x,W��A��G��3ú���7�'�g��X�t�"�,p0 ֕�_)8S+�g�l�;ȧ�̐4νm������~H{�����A�����#b ��#q���9{=y%-F�����+ڐ�ݬ�8��Z{�د��=�X���I�4P%�_�z�s߃��rC���G�dڧ��RDT��+]ы��q�"����$:S�&���+���ު����D��"�(��b˒k$�=4gt���uH0�g۠hZ���y����cWu�9�t�8;��<9�w;ś�m���r���w����8�o(���5����g��W7Us�Ÿ�M��ړ���V��ie%��a{f{�k�@1�y��n*�M��9x�����ôd�w2��t��Q��Q�ߧU��S�i/����גz�nZ��sK��o}e7l����h��o�S�6�VO��O�F}7I%��$R�U��5�.L�ɇK"��y���c�V+-lp�P�t�n�����xsm���
S�C+gL7 �Ώȷ��jʹ����bU�rf+�׻�t�KNi:��6���w�Az�<�6}�]#�9)Oj�/�e� �mx7*6��_����C���X0F[8tt���ȷ'!�е�ɘX!�*@	�-� ��q�K���%�1vO~��_-��bm�v��&FM�	�n�I�����]?o)bB�Ӻw}�j|�p�1����M�2�Q�>�g���X-�ݴ�E|�6<�N}�	=zy}�)?^G��.B�`��w7�<p�6�h��Y��|��|p*g�sU�u�^S[#��AB�Rlרt+e^���π��w�T�?W�����	`V�\��IQ-�����Jlw�wj�����BZY���Ik�^M���/[#~��#��T�#��@��ᩧ���G߅f�2G4)���oj�J� {��u�7ge�Fap�ʠ-�� I�=[/E��9%D�4�`��`�]�rǁ��s����+�I���5AJ;9"�d7�a��������A�C9L�C��n���NX�ɼ闀	��5&�|�t���-�����-�&�@\������/-�Z늄Z�m@M��*����y�`i�R72.T��0��L��cĠ٢c�F��z�<!9	1x\�v�,A*���s���Y�QH��@+��l�=į#�u?h��H��^���&h�������� �jX�m��>wr�󄏫HȜ��s��t��b슒�� �u#�Ew6Y�o�#��ɲYl��1��~��K�L��YpW�!i�T�e���(�V_j"�u�D�D�
�T�K���X��9,�u�
�C,���o�]�� ��;긕�T�, ub�)���>|��0��,a3�	����^�9�E���+��W�3��������J���ZOo�< iZ�ģ�������!��Tb������~0��8<�/m� ���휸#����9����l�B4��Z;�߫����đ+�G��\(,И���	�>k�"KG�C������rdh2�1���A�j.|�a�z@�6�}e.��Rl��S)��M_��&�GJ��k��+�$�M	��ӻ��Ng�֮k�v/:��3`�W��fN=ٝ��c��)��0 ����A`N�$C�g�b��@B��o���_M=n�t*���=�C�x����ɶ�jM��<4<���L�<
���"2?������x/�.�ї�6(�ۙ�L�+$m�!h��rj�e��mp��?��Ծ�������J$?���`h^�q�h��IQ����뤯ݵ>	�B�S��0���,%eF[�WN�I�h�����4K܈��w��Hю&�sꕄ7��|��2������)s�8��C^�ԍ�&M9�5c���M��VV���|�����ˊ�?�7M�5��	��G!�ތ����Xw),ζ�q�]/���O��OSQ��`�u\�&���*q
Q݅���q�S4��z�r`L!D���-u����4rƝ�C����
�S�'�Y��Ϻd�#@8	�(�.:��6��w����X�%��6�.|�� )���/�<�&���HIoR������ܢ�ٶ͊����/��_}�nWG��h�3u�ic��~�Þ�w ���B~����ͭ:4�L
5P�ԋQ�E�y2~��+���t�~�{��[lQ�_S�^׺�8���뫳�}��zy5� �O���<Gs�R�R=���~ˢ�}2}$`�-�b�R�@�a��	0)�������}1?_��?�1x�� x��"���ûg�4��w��P�|ҁ~���̖�����1i�]����9_����՛�^��at7���H�G	���qɴ�.�h���+xKh>��)w;�س?�����3�~bU#�"{	 �ݑZu��?��ֲ	@_U���콖i����q$F�05�2���0x��p���F���l����a3�}zf}��2��쮶�i-x��.��Mؠ���!8:p���4Ч%	�A�G�46�<�*��(�R�k�qv�)_�����a�&��_Q럻y��Wy�	�����/9���`A^�3��x:�\�`�7P��w��P��{Y�ͅ����x����"eW�����f ��r)Y�QU����*чX�e^3S=���jǌ�ߦh{x��͹��.���X~�,�o�N�z
��P�(۹��h�L��;P<B��i���gcC��zS�(�^��k���K�D(\q�~!�i2k����d���	��0��;���2v���I/����%��2+!j����T�;�[R>>�7�ߖ��ثrQƈΝ/�kcQ�k렛���x�frw�=��qٶ�Y�K� ��=.�ZG&��'����fĄ����>pH�pZ"�������f��N����=B���9p�ґ����16�P|�HNj� �����c&��o,
�nl�Jb��IY!�TY0��AM(� |u�j����H�䥽���(�B@ j�}�j�y>9�旳�3�G�6.x���芪rߊ@��IPS��w�ā��t�� ����#!�ix�a�D�{�x��-r����0�k�ˇ$@�O�g��&i'~�n:5h���s�ȧ1��%hZ�Q�:�'$qq7��A`[^aߨ����q:M�?��#�����6+eW����}	��u��{Z�v��1�a%�
@M���}g������e����8��nk����Gg�(��Գ�~��t|�}N����9xfv+y8]��\v��a��<W �d��"WM.M{��xg�;�V�~Yz�<�9�ˏ�i��W�����K�1�e>�d��#�l
y8��DtVюB�j�p�U��hSbf`Aʔ�FI��s�H��^\��1#�@��q�ֲ�.چ8W��s:t/�z�n
?��T8�vzx����{�h��� �9�$��ɍ�}�n�h�����0&�UL,�+@Q���f/�x��[k�?�1�BO��1B�����3���7�Am=�G�q=�:1Y &J���j�3/��:Z��[u(�{��K`D<a@��{R���w/{xr��]K?��,
��F��?i��y�DV��'EF����V�j�Gs-����#,VQv�^�\;s�'�ׁ�ïE�m#�سe��{c��F����4��$Ղ�$�F2�)�\'H·�.�$���]��|K�2�O�W �x��݆�@J�U�w�I-�eD[	�^,XmÜ �ϸ{�Y��t}$p��q�S%�d$Y�I#⸆M�@ g��?,�z]z��g>�,W�gI���g��/X@�Z���XR�ۿ�}8���=��B�4��O&t�R���iã	g���r¸�s�P��#��LA��V8_!~c}1p�b����'a���#�q���f��V���'�xO<y���.��̨�xH���5�i���o�>��1�LS�N�"�J~'�uK���t'ԯ��(���"��� s��)
�ӝ�/���F? ��l)U!�@�C4	Wa�xʫ;�����ԅ��Sƻ@`(���[p��S	�G�⛔L��%ϖ�RZ�B^���Kp���i�kI�|��Tm�.�66#��]Ƒ��;w�Li���%	 ���QXO&����Dt����3*�h��jӫ!�.(&�5��M�e��#���-��5�0�igC_,o^��\���k&�Y�JO�2���ZR���P.m��Wv��a����VT�8J_|OYh�����u��*,m��J&A�
=��Vၸ���~5��>Wr�o~����҉ ���t��c����Ih` .r G�(O!"�}��Q`T&1�[�ap_�����NbaF���!��ŝD�t!k�p�X���r����;\M�ec2k��Րb��qLy�{c.��b�����"�Å�k���eED��V�����'�����hxBEi;�}h&v���(cd�e&��2A-��+��y�h����Um,��=�6"�4a"�F>�)b�T�{_���vl}���q���=Bt����ס��E�8J�:ޛ�-1�G����﭅)b�� ^6Ie�Ð�H���X�~�d��Zi�l�v� ��6r��i��N�G`�����jZ��= ��A0:&WVbȖ�.��&�t�)	��ƟV���cʆ=E���������
��W��=�����V��T��|����B}���^;�ײ�K��z�T"j�W
Iyw�~�8��n*灖R`�Jq���gO�=f�F���J�+0T��Wq�,d첲����j�� ��V2�v�'���<�Ǫ�a�o��-'oQׅ�U�K0�4ad5�B)�ߧ4��9s�o����T��@ι�7B-yP0�o�͜�(�$\L�8n�TU��M���6�G �߉,֊�!s���^�����3��
�{xfx@(��/�tš��3��P��ЁG� a��vҬ;z����u�sJ��g��o�@������c�,Q�Z��C������`�8��Q��i84�*!9���+��c�ֻixK.��E��rz�@��w0BWNAM�~�h��IjW*TE�z���j��h6��RT�3b5x�b�����6��W+�l�Oʡ�]����کX>�H��
�
ā�;��i��ɜ��1���\@�Q��BW�
�|#������_���m�r5c��}�n��0�\���寣�s�x��dMP.Ӓ�L�4����f���\Y�R�bP"�t3�܎]�I�q/
�WLK3K����%�uf�3���.�׳�ma����W��|�d�V��H�O$�ǼB�#<߁�ܭ)G��%yV���1�b���#��e 4?/�r����GȀ�K�3��!Kp̫H���!�T�SH���6�ؖ���'&�v�z@ ���2�����N;������ܑ��5
w,!��3#�hr�@��Ϡ{6+u-5�4�� zO7�a���+g�ڣ`��&E��_�)���2֥�u�{[ܷ�������]64C��1�Ȳ,������u���K��յR92���K�e}�$��+G�@U˸�9��t�b�ݖ�g	�C���~�/j6I�Q�d��pOhYȞ��$�O�w!���S	m�d�q�A�}��4U��O�� ���7E�2Tn�K��������R-�0Ѩ�[������~�u�錅_�fΌ��\�T����m��3]�U(��=qƎ�@N�\�YKU�q���+[w��p���ߚ?�orJ�z]��!8��ה�֥H��[&w���:@tH�57�~�:��J$iRu�s�h���P�xN�ր9	&6ɭ��%�Ȍ�%��VV�40ܙt&�h~���&)�(�d�:���FgMz�6ӆ��)��攴��^�V��R�U�g��J�=GB�.����N�[�0;�o��:Ūx!�ԡ������eE��Yo	�6E"�f�5!��l9=`y�X�
�o�V�o|♪%����ʃ�ġ�Y���X��l(o�x+A�ª1J���*A �c�9��yQ)ŤJc�y/��f&�AZG�~γ7���,�F�.��IX[sֹp��>������6F����r�1K[z
U�5�Y^~(��dR^]�Z=>�e�Cv$B�Ϗ�9b����y!��>������-ۛ��C�̧>t���9���e�˧#x���U6���u�yj��d��)'o�(l
��[�^ޜQ�V~�]t�B�f3�&�lI��"�z�?����=��p ��1���:�%eY�twvJs��+������T����z���(ʉgQk�!��[�����2�>�5Y �[q?����e��+���?���B���gv[3�X�q	�ު1M!�uFW��FU��W��]��s\<���:��"!���Fk�K�vvG�p���X�1��xɔ��M�:���6���K@��"ObK�����r��_C܊�
DֱvR�~5QW�d����� ��t�C_V锷<`i��D�}�:w����7�#�#��w��{5"��\�	�|ͳy��!�=�;�5�ł��H�?[�<��FpΉ�f�#�L�­�F��vF���O�Vr�W����vE�r;V��ֶ��'j9d�Ee`�~0�����7���L|��@(��A�u�M!�N����r�L_�R���	��k"�X�Yh�DBa1�~�0��с�"��o��Ɓ�[���ǌ6�卹�,i'�=z�?���9A,���!ֵ���h�Oب���'=�&7��.�~�:O�E1�K�&�����Z̶�WD�`�q���Z���&Q���L&��-��;�MY6V9�.,��"�R�ű�ؑD��K�ǰ�B�E��[�e{�b�d}����p�Xr�3��}kӒ��S|���ܱ+m1��ce�Q�&q�Yuu6���ŕIN�b=�oo�#af��V̨Z�RdՃ�&���X�+QS+?hq�I) ����yO>B���u�)<�� �Xa���)ʍS(�A�S�5�bE����%V*��H1p�������:�۽_��c�����q�J1}�o��05mSWqF�}�X�S��ׁ��8vei0�@{�U`'�<�ܩ�(�r���٤Yj%..�n��+�<�ڎfy�E�q%WphU�Q��YG���ZM;=��8m�+I�l�s����U{D �d�͇�zp7��u���
�b��(ب3�h� �)rqH~����<�V�a��a]#���k����hz��]�[s�ߕYL��cr�h�t��U��C4�����T1� w��20��g�{�V���}6�S\�z���YG��Jm�ęK�&�O{Z�ra�l��m!h����� #�D{�'}�pi��Ǣ�,�5�u�X��M���ϒ8��9j�i�9�L�{��6X���
�6(�ʰ��hH'V+ZHL_�6Cڳ>�E?��=��=!;�]���A��-����.���W²�v{�q(��Ś��s���-� m�GÒ��}��K�K�vj0X�J�� ҵ�?0A��m>F���Y�߰<��I��l;".²$���Oc��Z��4 ,��!�w5��<���R���7�B%��y��t!��vD��7Tf`�Bo-}�9�(Ղ콳�#I��K�R; y��M@?	d��=��}�4�)���~�'Ԁ?9h�~�5e �&v�ĩX&�)uk�c4��ғ�,�lb�/x�����NtZ9�e���P�F�3^�ڪ�I�IbO2����y2N��J'����R4���_I[�~p8��Ĳڙ�Г��c�pS�����}���*�G܁E�~�������K���� �7n�A ��
��9_Ak���ro4���5;i�F�I&ְ��})�ڤ�n5:��8e���U{�P����@��o�ja���(|+x���ϵC�]$~�<�����߻��` ���&t�\'pF�u� %��va�Dx�1k���b��ܵ����u�*&|�2�m��@ƭr�31E?�8�u�0fbܴmp5�`+�V�
�#��8�;d�^��G�7^<z~��:���Qĕ)�3�#��7��.��裷L�!��rpY-�y��}m��F�2��]<Ã�ӛ��$�>�A�f�h�2�::1�rɚ���u�Snm�2�^ટ*j5�#|H�4���nv�xqe��uO�0�d}L�����(�zJ'r۫F��EN��>��Ե���(Q%����rbPdbe3�@�6H;tݟ�<���%����krKe[���_@��V�@���O`>1Fq��{��e�y�V��zRI_�
ٓ�6��+s�m�k:0&'�m8ɟ������A�v�^�ۖB0{����y��ʶ�Uܤ$�c��A���s��Q��Iiq�ɕ��)nTi�>~9/�T����=��?�A 7.VB �䬕dw��)d���&#���E�92-��ߦ�����
)Zd� c�NN��=�I�>M�����!�r�-�蚾"LD��#@��([}T��(bx^`pK`�';)o��J�(�ɹ�?����l>��'�]xK�,q�D��5���&��J,+.�a�o���5
�,����YN_��]7�	��?��AK��Q��$_	G_���T��,x��P��������Jـc����]�K��`?GU��o,u���"
"f��D�\ ������4LN��L��9j��3:h�Ê�Y��~X�2��ť��C�F���������.����j��	�����p��}���1ӕ�秨hF��(�7�� ⯀�'X%�����T��_i��&�^M4�Ͱ��`�	f�24?o����W���n� @���{�[�T���ce"�,f����>���C�'�f5�d�&X��b�*1l�'��Gzz����-t`ɱ�)�ʄ�i�K|�6#	x�|��[/v��a�H>NM�� b=�䧒{+yZH���_�"f[ ސ?O[��I�#�>�c�)fIB ��*���s���1��I�yYc��`]���&늰��4��Xݼ60$��T�/c�G+i��� ?zR.թ��IJ-R�T��y���w�EC�B{��<��ucq]+;�d#�HV��U�D�ls1v	�8(����x����%8����3"������C;Lŷ�y��uU��]��m��DQ��,�@?ڲ���e�˿ 2w����T3dhᓡѬM;|�;��+]���OW1]ލ��<�iH��Еn]W��7ל�ۓ�����n�5d*�����խ_pJ�	���ü'R ���R;���?�>�W���	���X��}�,����:0Ż!0s�t��96����l��y����!GL!GT)͝�4�U��O����J;��uvR|i�(�ZA����g�ը^Z�j�̦Sjc y8 �L�bo@����wv�2��cm�8�6��8��$#�PfjE��6�X�M~8}�2�:�T����1 �d<r�u�v�&Krl7�O`�����f��>�ͷ��t=Y?y1��Cf�s09X��0C;x_��?w
�q�:�}�t#���*8hD��a>�Z&�ɮ@5�L�c���EA1N`����}�����qٿR(��Q�?�G���xLKec@KX�S� 8uٲ�������JUP��l�Pnd�3��H���ӝMت<!:���z#�ʡ��>g��w������ȝd��e�[��� �	�j�p=�45�&���	77�AW���'�2�i����
Y���6��'�]��2�5j�'U2�JU�ƅ�u��p8��}��t߇e@�0���H9�;�����������S��= H�L�+�>�����^��N��h�N"�}x�~�df�^�����I����h�۶t��-�J�_�V~��b9�ZȗX��"p|f�'��p�&zX{R�zT��^z�X��L��R�%t*+P6�8���&.���p�C%��=W/�Y )6�#�0�9�e����i�h��-�,HW�3���j�F�%���ȵ侫�`"l�Y����W��Ga�%3��^�?y�{��&�9�[�~�� w���|�櫳U�tα���>�[+?Z/&�QY/xE��*<���w�Ĩg�D��e�h���k������$9ۣ�z�Vε�Z�$�6m��6%o�+�Z~�s�ԁ�ʅ(��HZ�ѵX����期g���z�B��q�Ҏ}��}(��(���=��������5�&6T#�"E��$[��3Ov� 8PA]�ę���e\.7�l�-��򭝮`
�	.:N�t�7�<�Q��&fDI�� <)��/D�mT������~xO	���Y#�Ch��2�<�آ�����ڭtX���ɵ�U��&��\��&y�}�:��,C���@dJ�m�>��Ԋ��XpS^��hG� .A}��{ߤ+��N9-��y�N�0�p�  ,�Hǭq� �����_)Pў���3�Y��	�D��ǁ�(�Şb��?{���|���Ll��A$�n�ѷoE�4��k�ߖ$�#84d<�b�]��"a��^�A.A�_O��ͳ1�?�d68o�.+5�]w7��Wk)K=����7��*\ �y-�]3��Z1T��h2��}�,if�?0P��2��'z+��r�`6[ai��9�[y/��OP��!k��s����<q�z3�H�`ne;���>�+U��
ِ��Nw��OO����"4�z1��B�V�RT����aD;(�������C�W*���4�����+���h�O�;��Sj�t;T7&*$�7��l���/�\>��)^�k��O=n��e�9�pq�B�_�L!1<:�r,5�kum�14s���#3��$3ۍЅʅ��g�3Y���Z`��xQ�_LQ9k#N�Y�r�?�'7�	$��v�S���CI���<ȖH��x,�Gj�9�a5|Q��V;�Dظ�w����HjE(�_X�h�
f�C�k���]G&Jΐ$�C��S�bt����W�(�Z?��N@M���5�G7+_�Li�r�/Z�W~�;PՊ�0;8���s&~ �н&��sڊ�B�:VFI*�����7F��Gi�kKxۢ�0/6�XՊ���A�)w��u��Z�+۫L����MQ��r�TH��! �_���0ި��o��8I}Ͼ���ɘV� {q�<�����t��Rp�z�P�&j�@`�����ԗ��<Zy���D_�����h�	J_]/�36����@�F��"���&n����)us���K]�G=,.�����k#KF*F�Hj�
r��zѝ2�C�x�:�r�y�t��	��60�B�F��w��������\���R}�S��h�ʃȯ�a5jˑ7�i���ǥ7��j�ĉ۟A�ä2~Df2�H���rI�r�����Kf�zN��c�6f&�J ��8�7���!G����^c���J�8��'a��c�����F��$f�pD���d�#5ϧ�D�`\��H�o��Z�<^�
�:m&�p U׏���7)�`R[[hԲJ��}c�}�hh�0��~PMr4�"F ��a����	tr�����-��Ϸ7��ۣU�1��3"˄���$�W��)��*����<a�t�ؚ{l$��t��b%)F���+|ttg�+cǕ���úG�H"��mq���;6ܿ<�Ҏ֙_|:���H������_�Tw`O%���C�r+m�?e�֗��aw�JA��F�ļ����f�ua�<W�e`#��ͬ� u0ϲo�(@x��(E�w�&��ّ��M�<g5X�\̫�h��H��҅ɼV������I�����5G��g���[�0޸YD1U�aʎ��8	}���돿�8R\�k�[�b�g�j5��<v��Q��&`���|��Ǥp\��%J��5�����n����*�p�#r9��b8�>ĻvtP����.��:C*���B�a��n�XTV)�d��{m5"�4���̙���������ns�^�������\���>y�ǵք��L��b���6�ٵ���C�.����[+��U
��h`�k�4��!�P�.��˚�O'�w�I��3�٨�x�>��N�ḵL1��ȁ�� q�u�
rP���v��A������"^߇_cբ&��H����X��@�r��=ʾ����~=��mVk����cƀ�<�5�΀���mK�^g��,�W�M�� �0U�������������T�@@\7R_Vp�t537�8����0[�vf���Ž�Yg8� ^s3��Smm��MmvGlo�b��'6�����;�0��v|T�){;���T���Kf��Jj5����!��Gߨ
Q�r2��7n>�[����K�RJ�~}�u���T�5��%���
�+�ïF���lh���%��m�w�'kn;�^��}��R��͒="���~�2�b'%�-X_A����0%.�_��f�` U�Q���2҇ɮ��x��vt��Qk	�/�E����F\��Lv�����˛� 5E��Pd.d$����+�[S��@S��B�T�EA��[@� ��nԁ,��G����fX�%�I��'�Y��ơ#i1n���m��3�QO([H1RM�Di�_�GM�2\b#���%����'