`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9QNpJbjoOi25V6tKbp0ux730bmrNBVBK6QiyCkTy+onhgEoAuwCTjUWFmcNiCZRARqx3hU7xkp2
uVLR4x/Z2V7h1H3q4c3cVkUDmPKpg0W7rN6elv2RUbUR904+2IKB4R27NTKkWazElpaIYJfdDwCA
ztRy0ubaXMO2cKTXp/EJ+r3f6KY2LFgFJsnQBTJa7lshAY2qaXjclPTQwrZNRj5dNz+WlCANDR9g
kfZd2N0B45TlRSZ8n92x3ETsHLpFz6mMbNUVvIbNhG4lPYvbqj3fGtnohL69h2P3SGyeWNaMT8dS
i1TPVOATH1LHWkhe7NiP1qb8d7HwkIN1xnGTNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
YPQPtyyLSZanGKUgU0nXyrjZN0SdgoqaIRs5kIBDuQBvHR6Dk+mLrep07bx8ML0tIp7n2s4TXlZw
EexIGDWH8eS7wdpSbcBNpvVnKalTcAVTDa/AAYdFTUqYOGrTSSn8q7anZSa1cKmCh3N9PUG0d0JI
/Uh2UC/UrxrvCk3uni6PFblIPlSVXZkQVeYVyjwJ4PMdriAS2fa8p3xS98EegFmWxsjy1EeyFbQw
6kHGpzx0WYJU7QswVopG9oUYo4wse5xLKsG63rAaHuR3Vf9mli+Ktma0Zf5LVXZfyXv1YOwzuAD3
StfwDoYe/k0ZxYRW4ESWJiZNWObMgw+nHsnvhB0lEzRRcLtFF/l0zuxuiiLQPvjeO0E5bfg5SYgI
JUG60SooZTcLBlb2cTSRcP+SZ3KhlC2sB01cp2Hk2lJxY74N9hpug107/o7x9x8wCqPP8hjupMSn
pH/QPjNpLw9MOHSlIjYIz4jY0pNZU6Ba9btHutkXYnzZOY6ces8OtmT+Z7WqH7/m5N/Yw5hZ/NOK
3jkNG/nWvKnLZsiEyj7E0JHR4Vjk+Dm5YWYZydNzZr6Oa9sa3QYdNpbezBzedAWdp8gYKET6+UMg
y99cRZoB/eRsBG3yQFW2xgNZUBgT+f4UE8m0O7H6awQoctazcN2uteZXwpq83Xn/5K/OZmPEBUHT
AqkoiZW8XOf1CjUxeDvws+6R7nf4OOBoVI3ZWWHimogCs95k7KryJrBQVNc/gTgn3vFxs4bsvkKV
B/cGkRWVPmlM4YS1dANg213pw4dg+KLA8oHDPubyW8uvyf86ViYf6GMm/nnxOZctLHPMucWDsw3L
oUGEbWtCL8PmbFnUP+VOAMRPNOcamE7yRxXkk45vo0Xaxurgs/BE5KMNRqZIfLQ7Eo1KtXNqVbxW
HNM7AdZSOEWCE2m8+JruZHvmYdzZMTmD3kpihIbQuxtNJ/Hp/injE5CVzBC/lM3CRUZSqLwLq0nC
8DBg9tMUH2OmMyYLwKIpydBMxbxgwHbqtTsQdHbOYvrTabXE1zZHhAIXeMHgyPAtLUaF5++p2d1u
lNlautZUPreFYJF2lBnFTO70n9rgR/TEdXfycD8ct+xLb7/xlcphC/zWdPZb6wJfUCfMAMldNBHu
PqJLkkLWXAZe+3rzVyrGPUlE8lW0HSuDIWOMqlY1PTpQSROvVsaSo9lj9yOnkY+ud08Lcvqrhzcd
DXOjvbqoAp8WLamrBgelvHf2V+8/fRdUk1OFhbQbDWC2/IkC84m2xIBt6KPQvZ/00M/sVLS/LE3F
un+9bHsCyfp7BkdcfYbSo5pFI6RMCXrldyMGEtKIM1m2ThYwp9/74ZQH6mjmi7+r30S76eoBxVKp
xIa1fZEEr5yxFpYr+IjVswj9uGe/Aw1+yDF4pwARm0PCZ9Vn8NTzAnuME7QjD36PnbdISwzL3B/H
n5WjMrXT2JUEzOf4bXTolZZIrgfiYM/or7Wyr6d1oLwtdXvFhVt1k4jsG+a4y1EMxwfiXKnVgiCB
RZz0qoFKm9rJnT4geeNDxlWvR/tz+ESZmLI1iXUhfS6kIrFCBYmJ4oAp38wGrF3fWa7qIyX//xra
KdtJ9yu70+ImCFYyP+YbQLf8RL9yAFMT7p/IPoeHwAfWD4vtbUdKd5GlnmzMm0/TYXWlboC67LZr
NYNlvfKQsuFg1EXKDNX6Xeb67k2i5ENesFaJQl6fr6HMbUoSU6fobz31P7Tj999zlEXUSQWVzZje
/oDa8XEeKjLwaHqctefhCnce39hbItYnldlUBvwAGFbfc67LoNUBTe7MvQ+c++k6SAFPMj7FJJgS
fu5PQ5ZogisE1CVdVFZ6VAdJZhuRWc2KymHk0VTsTxF1MAp52ztGeRbELHL6QciaapIMIbFZ5L7o
v7vnqQXg4jS+hhqB5qyUb8/JnD65lJ2LWXHAbUiMvPb9JVGmiN3bYAaQCfrMkYKu8elZzdSEweQ3
RIfSDropd4deSTATQzS0n/VXswm4giMRA86Q7GMMNZcpUCg4Ks71Rwr67NGUDBDT2ULwMUY5FzRD
Lhc4InlvwIkTXeMgQY4ZC5gSij7zRqExaDTtRkxawxG9aOIyWjxLyQ772KXvS1rG7/0fTAHyevbW
2gYG8c8XLaEf46uvHWnd7l/QKfAT/WqrezGWi3jy2E493yufjba7ZnLGAWu2dglZ+QC4qea0qLpM
hUiEI8WlnLRLS9w5Q59JHywZQWK3JpJa2L6veeRaUulktY43EEnJl7dbs0VCdFcm9vo5UQRMNYC4
Btl94uNHUnGp80IemI1qegRTkvgvtihsFumBckhenhxykKx/8GoXrlAvVzuOpAEnCOJYKHi51sDw
wnh7Gl+H1TNdyxA8352kZPmwhuGMw7S5hlLbBkJSS1T5ojq4sKgeFhmdrYv+92CfaZbjt/Nc59TL
L8acvYTlMdLFiCQy2A+M0I7/8xWngEqAtpnWYPwujBINjwLr9KOn6Xbx11vi8K3+78DevJtWyKxE
oC6rerdUTeP92r7Dad+wkwqielCaHpjf9QWb4jHJSIpbKrLjPD2og8mOBPPi/DN1zrJnDN1HbKZw
RnCVGmU39Xd8tREYnvlVdQrC5oX72MCQD2eXRBcClMCBEGS7SaglvxyNHD9weAxPV2jjaw97BZxG
w79lQrN0ahdCX8LTY2Gdoz0rrM8DruFfc+OIpNzTK7I3ILCz6mK2SuTVyre66TE+W6fvuAXLwI4T
ZbQEcqAgkJ2q/P6YKmVNAQGKxGj8Kmjlzbe/a4pvyQxyS8JA6QAPJQ/quXjHJXIuKelbeMqFp8f7
LuPBci62fE88WXvHdh9qnPZMk51JCNa2HR/J9BrrOmMjQ2YO9i9B5LQ9IKoxJcuCM6WOtMbXtusY
UoZJkJBY1AhSvVKdkEatHQ8EpJCmdLvnHCBhYIGlWJscynw0VgkWGH4RJixnKg636sgN/jtQsLCY
pHSDGZWiJle3OmLl2GDBqKXqyFg0DmvGkYWv0EtD1k2o0aNnbOJCvT9863RdXPJPkhf4yi7aUGNO
lpmhgx2fFPggFMuF+W176c1VU35EJd7kfR82ad1hPzW5syXct3EaAWrL1xN8KQCalBHtQ+xmYzMr
Zo693YqxlClTlf/eMf2PMh2VEBm65KSfg2uca8+kXIshipLYMAVCmuQWeeDAnHCLM25qrrk3Ns4c
EWS08+nQ9QNHs2HnHYsmsvSch23aaWVVkW62xtlmIFRli+d5/rgoQ8kWgl6LtQPK5DnnrBejZzSm
I1SVNHRLXr3HbZloIwt4zIFwD9s8O8//0yDQMyTrtBFIvoiHQdsMg+WcoePMNSA6CpsRKb093Q4S
4c6Qfq/IHyBFeb10IRrx+MlzZGP0nbvpH4mjLACroNnSAX1gOwYTOOEYPubpAuXiNjVUjr2ddNNy
L04tB/ci3yN+TegFxX4kubfp4Q7Sq/pp5yXJPn8vBvncW5B2GWJxpx4+qm/vhnZEfnYKs8LctXhN
clJa+vqvyjE4A5ry3sWXp+UqDl48x8EazZ7k5ruZDkFRE207xQwDpM6Mt2iHBNI6Y0TVlFcHEXnD
RY3qy3Z2BCCDU4sEszOn1904F9v+qbDQME5A/bjLbGqlQx+aF6fvxpovE3ryDHzc1ncnYb2Ux+I9
zgQIulUpge3TkQE1Dzgl6gwWe+XZ56wcDi9JHYd6/4j1dXmJAgBup7TrebZhT+rD/ju8gdrWmw0/
LdOCsPyzXYGaie5lSFZO4FnQp/HdsBdndPhgzJHv683RI/AKTi6EsXjaKrUYRAad3hQFnGCS96ub
9XIYBcRt6EAz5bg41HGWZrNUOASlkHzJNKLf4cBGsKrfP2PiSaIvSAJ0x30s7aBSOVjrRGOs5Gq3
5k/nnqNJP41NwNBGWtdQqdY7sTNpkpGuGsRglvJDL5ktIDrn9DjnVRAMI/6vBMaK2NXITEXPbRUZ
gCRF7fEOdjk1a0mllzBnDV4Ftqfp2+nxpCO+kMobEC5KDH+4fC1xBZbKInrfxlaYrnB/iuziWFH2
kIMxu4gSp9iEaBEPGhvmZNRzxOxUgGecyrZzy+iIIO5yfuRsca4sanyqNPBNfTzWmkKBQDmMBHMs
H9wzgw/XKU6XeIwU0JEXeDrrCeSS11twJUPSGXuMitZboz42uYbEnB2rQ7nCROri5b1mAGIdHN4q
DsJVs4DxSpKC5+o4lgwph5Qkh3cvEjfBbsx3tOYfsmz6YACzCpnfZJ2cmtS7aQptQ1oH1ljOMhty
d7+HDxpta/X1gcofTCujx0uVXsEyNdQinrmX2uvZM3FY6tnr40jeVTKOa4uQIjrdDS96vvt5hqKj
Detz1/3Jtgg2LxLcdfTAyrcqPkbGZ69DrKEG9uI9ECxcOJRskahIIaRlfBsAtf5NmBHq/RC7+q+f
vDDbkvDo8v5ggVspBTcMHo3yYiScaq720JmmrKKLl9DgC+zbp8LHka3Om6FozxZC/obGqplLS9zZ
C/C4qLDqdy5wCcunXKOIjCN/mwugUq9y8D4ShIe2sZsAaH0Hs4jFQXqaL2Er8TAdkKLefJJmoli+
JU7PiIur47MQ/O2POhreshKHpa4dAiWE/RlRTmLobVFvVYZM3F1/0ol9a+YEHU2i2N0LHXvKkDxM
yVbXjDYJ6PwvEy8ZHgfS22fHeApW8907v1oitFOueBvTHrF+O/UhDpYn6oYtlY+y/5OQ4hpzaiYj
r9ubZMSfHewmuJg5pO5NmLQv8dySUct32qrTILqTlgVh2AGxoPvrj3htBp1lNQOygzKseV5kpRQS
xkAU2uhUdP7ibzUI7US3N8kceRI634/94nrXN3wtxFEvv6w7LapJNVgRhycZKCZJz3eMnh2MGae4
G10MoJEVO0pbx2mi0kRPjHuABz3OpMR6wMQ2K91fl/rMqeTW7bGFQ0DcuNKAjazWerx08D0YS3jv
7Nv+5jMWQYA2cpZsEVMvYybreHJjy9KyjkrMNRKbPiJ0SPJpRDfSzGRApG1rXUS4QpjiAeTfcizN
VCVZkgheVLn+qnHIsvYOvfMpWzAphapT/zdecdJktswtLrd5JcwN3LMzkrovBsw3jVjJgu4kUz7S
2+l83ZloqUYXjzuNHtWU1sXpvmMv257GTpAWCZa5hpZUGMDFR+KWrVfl26zAuYZVEYDYtERiPC4H
gXqk0OheBmQyP1ak7a9OmBM5p/2zaoVWWmtayXFe1LgaHay/D8IlgOsa5hUMyN4u657xYzsn16gE
ek/5bCn+Emaov7e4QEUyAaUs8Ys2Y3C52owkjfenlDwMRw6Qu8WZewrDtmtJaehRG87LHXplRF6A
+30os2R45o9S8F5d9FS5CjsunTkynhSgJjAJkHtdNmq2vAStwcez+YyfRfG0Ry7P2dmAw29n88IW
TaUynb6wUMym3p98vpTrInkJ1dNJaOEohjKv6hs5D858gLkm/xF53X3l+BHVKc4HaEH9vMwV/A/S
4xI88c8tQQZ0Buknf4NYoX0Eq+tOdmbj1Py+GVbG4emOlRbhk5k5e4PZqpfDq02yHfra+5RihS/l
3L/eV93U8iQfdgmhAV1a8mSnItOTxtvs8B24cRUvzb/2Pp8ICHfE974Hb0i5EHRoo+wSCmSOiDSh
NObd2haFw4PCNzjcQ4u0SVNraXbRJaDgAq6qepd2RM8sjQwiP9r3Suwbkva1pRDkaV2ovjsLb0qe
UN/b4pTqXyrpBAAymHqFjiMg9w5wZPMF0n68fpDEVqV9q9tWJOmGjOKjmy2Q1l70/k3RDFXvQ7ji
GsdS0IxfABN0awQJqKyP8AtXWpCNKYVIHiEW+UxZPXbB+rbO8bZLPZBHL5+fS3xo0dEiRD5zeNVE
vxej10ir5sE2ltljuegyNUS7O+qZBx0sjk/dsVko5HapSMXmIgVNlAa/zkiNI8dCSMgX1H3hSaI+
G5TZAYLB0W2BfVWJofMK6fHu5ZwCZrvNXo4lkgTW0BaurUtssExjRXjKkAicbPHuWmV8sZQNDzT5
bgwDekbCJ6wuG3pvRSlKbtJ8YDmSVvNHni85KogpaWrI7XSJ+dv5XdwGElNdZWGShBJbroAUld/b
EFUQsav5jcgrQ4rDxEnusKWYtXoq0grvG82uUaQ2VG5p2ljWaiIPl6jOlNOsLZx0FNh0WEyw3kn5
SbjSeXxIOkBwZ1axlIjTqHwkFbj1MO5jY8gfaHr/khz+Hp1onc3fNqhnAC+zIGdHoEQNeI72LjIf
TY2sFkQyZLXH5zoWoYNZFxXXqV7Xdzt54ZxwPjnNOkDAcsD0Fv8dfsYwsrosW7Cx1IrWEiL9+iaD
t6/pcVMxdH0hfl5inuSBZeDtGQo+DR8nLx/4UndMwsqcBA2iw86IpQ5sMw5TRxdU6PL7TACYnYfW
ORZOeVH2kTI3k+U3FrGssgmsXrHyEIAQEoifIF/qCQ6S920Ya9U+XzAgjlYeZMTFw2dbnbZHMq8J
scdYj6d4Kp6VfmPiP/e7y3z8Um95mznSEt7t2i/R17WojLxJ7+BN/LIhbfcNhKPwHITRPeEjT17s
8Wu3lgVU/DuH0AQVPcAOrZfEJqe5TtmsdFxfbii8maFBTJaOfgJmJY3+aZaurNzu3yOx9dP3O176
1lU1iFirfMcKSis2NWV+SaaIQhsvJ4dX68j0WPS4A+tTx+LGHrD06CnXa02wFzWTb/9u1EjLxftZ
gP+RqkoC0kZnp1sxp5sFUb8g3f2i6oE3vxRseQfcux0yJmbO1EwGpMqM9y/RhnmjrY8xuY5p7F4x
VnAofux8FkOBlRQLsBFAyKKdzHC6pqcrYn3lR25pVcfyQxhRKYRPRIB7pDt07OUCY1DNN+i2Wwjt
Ib0pJGJ9IRH2uYdAy06G0d9clm2bXy35OPcHJDg0/EHC+Qe+JVQPyrwdCRSrlJosqzvpYqlKhiBC
iUo3vndA41OTIFHfU5woWYKj3IOopvy0siflRUrTbob803lc5xzcPTZVnq2nXSFzhbBhzBklRqko
57opfJQyiz5C0pAJzhKfMHW8cBZHHmRbt+GMzUV+Loh4IjXgz5l3ZXXUjqRiCEyHXyQNFzYLvFr3
1KUmcGW5nx2Knh4dtpamMz3/DtT/Yc4xx9ThDVihcmrnk8WbOy5P55FYRJ/Td4g3W326nYpCy8/e
6NrFkC8/HYxG7x3LKrb6Jf2r6v7iVg10wr9xuGS64IL+3eoskaPTPiO5OD4T/zINhFc5vn0KG2XI
vMJihARuKi+gSLUg9WDMcGejXnUlY5BQ3rdZudAoDaY0hw3HKvEceQfjhIy4PRb1XERWIZ5Pmh0j
jG/Z1aEA8GjPOYX4mMxiBRN5xWYEAIuQh6BRl56u3lcZWGdzpSoYEGnWwGShKLDTrgbzg/6pcHI3
CO5GOO+wbF8qFcphA2tkCGswSN7dUaGrMLuuPtiQKbyM1katPc5m9vNITjrkb3veK+iqczE6MPHm
HkpZvtxaTCF6QCZCJ/4mQtY6S/eZa2sCN3yLFmBvqWC4wjSfvAkXnnxri7NDSICizpKKtcfsgXgN
XhV+vgkQ2qCc8ELl70kbZF9jtSItcIAX2vycErKPJp6ZMUz9lJYaoJMmisd8jtNji+/dOeYX2eM0
Trcjf4PLx5xrjnXTNeO9Wd1PONyzAEwlJ7WEoezq+P1iF/pFxk/KKd+AuPWcLEC1t79VEHjXvp6W
glCarRn4aMMCNG1J2RE45X5f/GEgKIn5wy+dVxUqtMCgqoYtM0Qoz0q5eH884zU5Ef0Iaxp8CJbF
CkOSJGk4d4nDU7fx0PSVyap7JGbuJYI5ibNwyn6a1BmqT3tYFnHOjbuoWvqkFly5uAzIav8MAJ5X
rCsMLn5WWuNIcgYtsRFS1NRMSyWHeArHg8DCspdOFppU3Pm9TZ9tWumVwvPoZ83eEvMOTJ3GdRQD
sxTY/co9+/Jtha7rMz5GAf+WR6USxxatOVmbdcx1An+vPSJeYj5RxhS56lLhkjHcnAs2jVxS5t3E
IW+j2aC2kvbEDkUt92PNDvftU+0jKMYgDwvhphBaeFAw8j0Rd4g8lVTcPYopTeE7pnYQ+fbPzKqt
5eIgjT4WhyQFnlY+EKTVjQhcwJ6q47zGbjfKo6my7ewvJx6bcw5nUBz+4GGIfncqdRUggfwt9q3w
eU8EfuXOEIZUGPtlwp36gLGFF08ANZ6LnaPkTObfTYUC+BXekCKG8luXkwCV9qbbXFhDn7qoZsMd
yQeMqUQ5vLb8ScJkr4RwwOB40AraVcyTMrDzhIDJAGAl8HpFiBR/6tPT08p1wz766oc0MTmlEKM3
MWJl5HuvA+OHclTaJn2SZ1px2Y7HbPD0LeBxKo7X5l0gT8EyEmX6vRQqZaBp60YD86bv/vnhhr+C
6LNhyyg+O6yjNQCaVjZx7tCceef+xYcn26yeRwBvuZo9GYCKuipMkvtl5yOoGZnBKSzB5Zf73N6Z
IC4wNTO2S2yxMYYKPm50lEyMQ446hPaQofsNQzRi6oq1C8kf2TjouaxXZ3j57bRgOYTzWdDgK7PG
GDz8T0t80TVEF53kglgvYBOYV1falDpGtDRwq2KKuwMuntdAx2honWi7fxK1t9qePCdK7kqUvtWR
VyHWCfRqqae47n9spkClhlc/FgxSiL1k4hrM5SMeX9mw74+LU+ACxkEUBQe68bNUeT20UIIoXGrw
pEf7e2085Ee6KIneiwOBjO0GAZHNB6K3p/mYtm68uOmU1/6NqXXQ81stHXcEfa+Ee0H9cZSFgM1D
7sBQ//pnNB+biehDM9XkbSeL8Lgjt4QdGlc5MTjqHxKYB3kSvcFJjfe6Zeqti4EndyB+hzK/Fnd5
wBClomG3QfPK8MrB0zKfjuzlTQhkrShSVsJleyL517+WZlmFoW5bFpfPvFuDMNxMGC3ZauRBbACU
xBg83OD2Rror9ArewWKiwtql41A3OLruw8fHlIv06prwVXclkpFGQkS5abFWYpIsQIp+VMezhW/q
KxXMallIgz/VovcVpZyS8dXhjblo2NwZ5QXiwpyuobrvZuYbkeNqpYqZEici1RSs45LhL4HoBicN
N6zRX2ROH2AtmdZfQ/HfvXez7jbX/nWoB4w1g8nJlRmprqhDlVbvW6bSq9D9WRBeb9rUGtYSHqQC
Qnzo13ipxFJgD7zTiJeikjNjy+G6lzfFtQBj6aah9i3L/ixPSjYXWPZgCOSQKCl95cRq3yzuzf7A
B4nGSEw+OBBlwiCArurgv+DiSbZpZWPg/NmKPjGZ9Sf/mFyJVWiLJEtHJXd7b6tpgydjcnT8eSG1
qs6vWHZQIftG55htaGuY7Nhrfw4YoOAhVH2tU3H9tBOoSCFzy2OZGq4Jm3gLIzhl6cUPnIcqvLiw
Rj9c+YBWNTe2O3IwcvE9/l/p/cpsqrGn38SxtKAtpX4PkF+zqL+GIsfTAaDQpFDw+R8MWQfbE/7C
8w9t4S6cv3J3RLs4kJkAPc1v7nJXXFa9hRoD38TM7KTmlSPwBlF5NQdeXxyCzMffcnJfjLZjBA9Q
nXSQZZUJDj9pIAN+xJ+pHpSxNL56vCQmXXnD+0bcZQYuItJG0ivRlx893HX7gsPtdBioB2Hb6qfJ
D6yLjZLAKWagnppF9nd/WU2wYAaQs/DiaIUHCP3yfCo/FRVjDCca2p+apV663+IXd7hgDXmsUXqW
/ddOiaiPPdxg6GRfRIOBlGMwa0b/xV90YuYXKMTWO2bCRbEG8va6622q5pLOxOpYYsx2p5Vpmig3
E9ozuqCUlFtHneN12w728EFMKvCnYtwf85x+/jwW/o+xCuoKFIMdGSORS6mYReEipbYC6s11n58E
AODm+Hgj/iVQA/pRVFR1k33m+CAYr7ElVjfG8UNThqVvu/UUqsVdaauMNmFSVWOpLgTfmlmKNqld
GalyhlkO9opQdQ7rKNQmhEF1tT9KjB39FG1YmhYyjr1DigfHg6eyRlRqLPeJ4JEK2emMB3MXmG/w
5xenCVSSbUTP01v49Is+xzRqWntiSYtby/YZg2YgdofIiA5dxutLgnEYDmOWhXVOW59MKYiO9kwM
a6sxPxOIDdgPBAYcoqDqXmkErfm6cxbPNYmW5nZNa4p0u5k0ius/s2x9VT1S3uBsAG+iP6R8a+bo
qnuXg2y707Y3+rN7gkjacZO90qIya6tZleNZMjKtPRU6eZjJAFytWGkUXtTr+BSUfjmr57qJcyVc
vX7m5n91nwO6bDkUfyGzy6kvMRpCtf+X+t0s4gY3JVHO8x1bScJvgWktRbIkA/BuUrq21w9+vr5Q
vUovA2OYXc0tPILn7T1q1MGfAzsfky/9wSOLo+9FpzuarBiaL5PJTqVDk+QPF9chcCtPULIg0umI
gBkFqC6HUVzePCOuV8Fc/PMfC51tXb2GQLJ2UsFTe3BiQIsDpb1aNKEoeDyGUxT7ZVtCG2sre+a7
F9g3iU3QzUgtf4J7zc//nlq6nvebDQiDipGNXdi9m4YBWVkcK0KeXc8YA6UmROwOK4su9fVMmrpf
myl23gXYhR6BzB5Avl2nFKWSVRJe4PYrDxi16ji3OrIjVVuoy9lyKWI96Njz4SnnyrFjiSp8HBnZ
ZLXJhAObDf2iFTEmwNbxZo/KRmH80F1Bo+RkSZSrXZz7uXgRLNcEuIGZ5rvNLqtk4L6EfKPuL7NX
qmi/ZOwkPvqYiOfzQUGvNEl0hg0b41mR2b9H103WQ0+T9hy+v0SlYTs2KUckRUrH2VbllTVzn6MZ
VfFzIoq/Z8/PMXshhPjZOCb/cakD+wZI8LewD0yAQvbdjFwzcKO9l5eMvT0CPOrTdSqmIAU6dN4n
Q2vDIl1y2H/SK5mbYTpr3bf+AvzXOXcG9o83+47EaPdtspzaYOFZz0hEfX9z7V7Dlb6qg13VJ6VD
TBdFEvSbayk8hK9xQDS7dofuz8KuT+L8K0yHb7aHdFi93/b2HeovmFXlr+Lrozja7Ae/Ho+4vK7L
w7JN4B7ySVkPxxqBTdhbNsnQ4SorwvdnjVkxKtC1jT1Rjku2QXdes36ilqOWXRjWhTlgOBjTY+Mf
1fjMRvlqUwobzUiGazqoJxKIsxDNGrd6qQiGPDx61omQPgBSiJDNy4tprXd9bR/Yw+oSoUGpyZ06
Mn2iV7tYbumfpHyAThs56AzOL7UNqdglemQqx3KCjMYT6KitsvMPh5DJxSpKxNJbY5BcVaHnEEwm
L1tAKF0hRMs0/n9MoNYRRbcmQNZ4UC3HA+ttGE0lLIrpzKnA0BS+k+AKHhshg9NTqWsm0tI7xeTd
KHjFeW6Uxyi+4Z0o6UeDKyIpiF0TR1QU+iXGAqoRr1ME1kiilcDGwCDui+UqWhdrIHJSu5tagCmF
+CS/FR7Wxopp7WODNvj4Thtb7jypuF5xndOQzADGsjdQMDAe9LKEjIbiY245KYNc2CNARiuOJfYM
zpSj7R2TlWSN1Wx7KwfnUaK/9EPfmpHXilscgE7SvcezNuXi90BsPY0hfttS9jcAbF2+DRSWEyk5
4qYprp1wcmGcfkNbPmMsVB688dPMHWQI2NbzzdtzR0yuHGHME5i8rureyBjvYdTpqt3d0AflU6Qq
IAGIGJKtoxyByBA6QV3Pz+cd4pud26EndOupaFU1vRRSBqhlEOKFPMznp4WFjIjyAQ+m9YCKcAdQ
MEQZt8kaYQ7fbST8jV1SuOzgofjIX4rOsA3aNPYrnDg89lHcRLT8PYhfDw2Z4WoS7szSDmkAo4lG
2njqAqLy0DSreOLVmQ0GN/MZoM/iixWYufSpFGrK1WSUHQdgA5i4od49EVeOFRwFNKeLMf4/bKJq
E6kjHI0p8qL+f8iDlUE/hGyZAiide+3kgEMf5qZItnY1T0PHvLkvZ3iFPsNHbkPA9WA8vofnhlvC
mGsIH/qTedj3/PcYFig8JW+Shcp6FGpYoII8bpNfFVPMLCkx/nq0qmcyZrIhG8ohEOni/uiBZ8Os
sqrbbIrRo3ZNxkHqhAIzz6sW1PBb9Zxvf8QwNgQM1oK9oUqnQdqu1F6UQ8oYIPvfv430JQhHeeXc
DhqVHuGfhxZ4f2bw6LnnJrGeO1pN0DmC7kzJ7SFUqIp0IKnRCHqJ2icLhiR/PAqB06TTNrbEvQRJ
z20HsaxUkPTeb4yyhAQV2K4nV9e0ryJEn2ubxqeOPpRyxG86xXtiA3MKenhnvxffOX5GvYBm5enD
+pB+7WkoWtGMukKUPywiQE5OgsC7scXakYgLwF/GxWwNgdOomKF0Ij5G/k590kuDJ5HuVJzevc/A
J+4bbJMnfOiVj1KKc4cBXoq+xkvkyYUwOIn/pixBzTGRHWhS3d4ch5OsXgNjNpXltNPAKE5C2AkL
r5ggAAaqV7YD3xDEPg0fJe4KJOptu/EwmD2Cr07IeXI1zv8roA52i0k6wwircbWTmnz5scCwnwsm
CDprRE8NQ0TeGq5ggsoVqqpBA5gF1UXIlSLh4zjApBpNre3gu7mXoQ6EqeKNpKbIpvDofMBMqdKn
SYymY37AUlFqdEm4V8uWkarjwqCBryMHBkaExA3RFmYNBc6X+6kuAg3MU4FoFchRyQWEYgzqN97E
ILEZGAYoEjAhBoOI9SxaliuYXPBozqcxQajn8O2DEH29ydgZWKxIYegi1vZOR/E+pYqfo/oH7blg
sFB8j8FV7UMhMkbhh7wrHyFNSufYuhQCjbqvHOt9Uk1k70bYA3Aev7rt2UuOlLiF/XxprJTxEdXD
iArR/2Kt3owNp6/E6s8hyWYgpT34M3KHxcBJG6XoW9zRFiWaShVDatpng7E4hucEqu4VfWx/g69P
w1TP7AJlIem5cgrgH5D1MfPDQidQlbRK4IQvNuW8jWsof1PEFr9XahxbISX4NAMZL2Kq5ee3qwOH
1+GYAO4mZTTSSR7pRvkKRp/q+IEBTAt6sjE6hr/0SPEaokMmbsHSj5duXsKdtguJGTQBW+ZnKh3X
hgIa7o/wjFscKDibLIoT0fbaj5UKPJYjOXxeYDCpY4YQDF07EtANiloE5d2/T1IO6esm3gwPj9yV
iY/RwJP8Re2yJ5/hg2NIoOrn1/M0KxmZsDwcYKRt2/0q1O6NStZNyzlojWyuQAoxSGBC8Hha+kM1
0JmAaKF98BhhBiajW3JQt80gy0ObvNUInU6BU0K1618TlHQaiEdX2U8zoSFiRUj6HYAcONqLz178
y5pQm7Ug87GiaF3qh6wmPABa8nLaJXKA83JpvtBHqQJ7rFh8JBS4Ty3cBIhnVtkkbgrRBYmRedOp
v0CZX1KUhFwyS0PMU4p5NAcTTQaWnYDVzsSQHm5pNNE/CDPS2seNHNUPCAlGew5CudM3eRv7OuG6
B/RYY3Org1Oo6udbUyh7ypdDmiL9nkqoBqNeArB44C3uBL56MwXVK9DvFVmxCNo7LA3TOarL01Dr
SnXUHMUX4KASzm4g8a2gthN2QDTx19y+cWvv5oK6eCwK+0rmYB0qWyZK9p8PKTWdK5VRkcUSk4xQ
seGdxbnsxfuki01W3jJo/3xmO7t+6Ziu84XlI3FulMA9hjhQr40jemHkTEE32nGwq2/7cVmPFgNq
vRTtf2/uuF5WFFDKziXaAzQiKtvPJprP2SIbyeUsuDIOSajEkBo28kL/spwX/PDSBLSYz9e53b0+
ILMhmQINzRE0Ch+7HxCWbTxbdkw/DDdWImt/+sB3TrVJ+MGaUfrToF3kMQrfrtiMCpb0yHzUZYHN
WUM0KNdgVAuBySG3mGcOTkoNcJ+hUXfXGTdhCRGcDIor7PytNn5zM6ZROlq5DnKIJrrkbOgGie6O
e8fMgYkusm9kMrDyATZxaLzIazDrIXoP5HZG5jFNpPL8vWUdZHSquhdapL0b/GIM2Xw2c060ysV3
ZlFeMHPihjN4Gj/amHI9oUIU1cgtBo8lLb/IgEaKHfV+WyDxbW+9R0guHOGEcoOLEoSItC/zTTMK
tERJ6eISJtmN2QVYsSVHJZEcqb18/I3w1MIgSjT6Mo7LMhGisIKEnQI2bP9rQ98EZiq9/Ty1NFpa
ZIfT07tkuO25qHzru2YEk8J0cxyv422uqo25qAb9OYRBdca//uidorx9EB456z2vZNwpojw2kgaR
SWkpIFj/Uf6yDCUA+G7pUPvwmb2oOdS/5/bXtanYo/DGpoji5yb5T1L0x92bynBQdK8MiYfFOH/E
wp+7xmFwJP24lICexADlXLA0lzLE/dJMe4jDk/RiXB+NTwcp9R0E8KFmpeRqCN9zfLGWJOvzKQ1B
xZPmsKC3692ED6PTeBZFbV+AK9OMH8LuY1sMTVrhlu1tuBJ9iJo0eVEOuJR6JEXC0DhEjK8zsUdb
oSiak5PhZfA8EMlN+dTHT/HnFfiXQfopQS8FKTveJOzYuwEKRdABAbpgeVnPHKcPTNuaF6H+eVDz
HA0H5AcqBsSdFuH0xfvxv8dIS5sxyYYydpuYKktNl/jyugdIskbYe13Ssiz+XWPCChEAQz7yEtiF
E4XbzNr0BKqjCGk0WVKccuyDwoZ3np6kUkCbwkvToh+wQ1CnKEpGwO8OHCO5gKei/H5QS1bvbyps
Im9g2wRKFI4t/+fj4P4qAArKPszjbVXsEXWphu7wKrJbBDQOQ4VopIj86/CFKXCoMAebMysgke7T
UReZocAi6R8qmH4j0Og04jkCTpR4863be3v0dIdlKLcsKiozXZvsJH5HAn3tcISWeY7pCYW71oRc
OyWDDugJ1c1q/vtWwDo9AvKN4g5fORzH+GzWVGmHbCIMDdn31jKN97ytoDgD8oTCzvuprYUoIFSB
+jsXqG+AVT3BsCdqdFwIjBIV396e5N2xGPEENFEYp7hsBkI7Xf50swJgGEWr/SaEeMUCqclaHd0N
K9keDfzfuDaGUVC0dSq0vKGLZXoQTn7h5PCZ+ajMC0GTcpvX3dqBZBxz84qrZnW7+IYdjKTiJzs5
HbNjQGPUFrwn/Xm9jyUSLsM4No3aZI2Zmu86zEq62L1QKvSgUbxyFiK1lYZwlyOGrFrTBzCe07By
Ghus0TAcVBkkAipElmYXqghyr2pUD/2be/AiRGlFZm/dQONrI5zqVsXdREWgz2XZJt+sZ5PzaGhZ
2oXK+vHu3dMHUTnedJd1C7d9mOJelcxpZ4IYo8nOOt27ixPmoPlLrWd5mcEh9TRloKzcNQPWTxsd
8u8PBElpLhbvU0zItdc8ic5G6OB+M6o7qOO3B/Tif+pdeaMJ0ezV0BajZSMDwxQPyRpb7Z2lGl3W
lMdZL+xOKhuAiACF5FciCG2GlzCwJIqQJRnXehiny1v/3kOouywsIeJ9gYsOZk3NNv0Tog5UoKcW
TjonEEGLQBJQVnlHeh4Hxz3+qjtDJpbg+FfUY1lwuz0E5Vqm6Fsjl4qQC5Ui1hOWfyXG9D13q5MX
XABjKdj8TcFyUc+TOby1EdWTL6uWgZnzKd5Yta/6jbuOxiPgKDvGuguT8VQiwhZa/rX+JbmJ5vqM
s1fbaqYnQYZxwYJ0uaJiK19t65AfMsspj5qD7fq5squIEQOEwQhfQ9L3x0wT1xppw2dPp6BBTbBm
DJnr2MZFnukr61YCBYHzz+3JaILsYK9ZYqMDTgzWH8pXkc+1tvSfAvt6TssUUM8itLaggYexY3Fo
XXbArkWi8bZ6Bpp7/I9vGTYbG1SqdGjFpwoJL4vJ84iVu/zeXDUGp1j8Jy2CLigeLvBWpcPbx6eB
ifZj0ktMMnUfAIjQ3QwntmIFe+Qs9rqw9aOg/7HCroGPwozoqKGNGpeJnK+AA3obEkWCZcJyG9+u
2GuLjhz5v5hNVQyXAU9Dck5+gzjhQhM1+KzUwGVPr+/q4LPw0hO4fXPAiVoWQD6qmOA7FIHV4umY
rpJQ4PnOXS+LHZgP04BEZhMLbSuqxjYc1hN1VWsIz5+Vn3BBu4jPTZ9Cfrbjz/h1IchVlE1XH90a
yaoGvdEBhJ/1rFRf9FSBUSLeVCT/d2jISCMzuGwAzzmwzkxfap08ZjSZCovzjB6FMxYMzgjXwMk9
bL5864JPWu5MnCkrCBYh45oEcP2TWolTql7SZkdM6l1DYX2XH+ML8ybnayT/s8gTvq1IwEsgnovx
hpRxKGjldPX6l4CeA6KmV2a4mzo2aWcU0kKGGaUnsdQOyBAj0CMkd9lLPMqdft12WCjiOzgGZzBV
LeFrkOnmyXnuBbe8lGbBahx/NP5t1+UI68oaVIILP3bC8bKrZP13YDa9V2SChfUhuAEZk8QgKUI6
rsuXngy0xIX6nhtS47fUTmq6DhIfUagGXjxtko/OagNajgey3727uR6RGbDY3AsEXnG3
`protect end_protected
