XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G�4õ{�W>?u|p��+�Ea"���Q������K-�c���;K�ZϾ�����,�0垞��>|������c��pz�C�=8x��"S����X��9�k���/��%!d����t
���9 ��œ8�t m(�4��@ѯ�Оq��دSך�T�J���_�g�sAL�W�S"�y�E����1��ƀc���`�H�����3(S+U��ц�'�qF�B�f4 �`UYy	�7�^,ibU����>���(�v1!���?vr(�̀�V;zS�F򻭒348m��Hm7ꓰ��|$U�������4�`p�37j������HL��Y�6��=b}xS��.M�������!=H�Z��Ϛٗ��;]����p�R3#3�s��o���{&+'�:�IA��g��iA� Pŷ�y�.WX�<Hzx���~қޕ�V�09�R`ᕝk$�
3r�E�d42@������w���=C�]��o�L(��~��H�z���T�Y�c)�j�g���!�h�������B��輳�3|�jP���06I!!� 00'W��gި�|�]���@a.��eE?�,��Y��踑�ƖA�V$�u���9iS*���MS���� Go]�}��;���#��^(�i�G�%Vf&<�cBE;�!�VmbM�>�?����@�Lc���G�y�6����c����3%�jU"!os�@Y�����gz� `77p���A���čj\Hơ෶�XlxVHYEB     400     1d0>��2�9%̵���j����!��3ZU�5�.��=�-�T8�(��ZY2��� #�>
�F�˷�"��G�w�m�=�D�+�kD�Z}�V`A�5�%�^�;��.}�FK�VA��]d3�@yb}sN��GO
I, ��:�[L�s3x
F5
'�)���pg��I�e&P�6��)7�>�V��7�l���q��������1L������3���-�߼����T�o�V#1��b�䗕�Tj"s�b +zx�!��N�x�,)�i'|c�W��ɻb��J�=�eL�`��m�:�|��A�)徶�q���z<�^"q�=o�X�/���Ch�u��2@��jN��<݀zկ��3BXdV��V�G����Jgk?��f���+MU��-�.8�z���n-���nJ�������X��Xؔ�k���x�5ڤ\I->������͍���3���8��XlxVHYEB     400     1300�I8�j��e�M-�B��>�aUB�4!f���w�D=Vb�d/�6���_0����#��ȃ�67��7�Jk'~Yt4;/���ia���4J�A����pV�/��3f����&>՗��J�6�(�����G������Ep�!���|���2B�eztC�# 6t\鶓l�	2,�@ԯ½�<�!�Rnv���_o���eX�pyy,
Jc����10�I_�9�"@���$���y�8�S!�h#��*���K��]2
J�!��Ҭ��rInc���B�"T��^u�(v���A.XlxVHYEB     121      90����v����|�K!'Y�]�p(9���h��+s��GꞠ�
t�H�MLv�2�ch�%��Ⱥ�8�eRU�O"�e<u�G���:7�w�M0l��F�pݰ�kɼ@�N5Z�l*���\|�.��� bwb�����v�L