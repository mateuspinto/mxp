��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��вV��h�tɩ��P���Ơˮ<��K��],��Pt�[���xq��'��>�=,������0*)0���X��!9f�
?�!��AR;�e-�0}�۪�c��:+,8E�% у3� ��-��cR1�=$/�b%���X�f�K��!8��£U�|�X*�'{��`c��S��_�<�W"6�'bW u���NT�[%�}����?���c�H#��'ޑ��@����N(,�Q̝h��>�|?��A$T��G.��V��t�q���˕�yfO�]g�b��!�W���Ĵ6�uX���ߢE3�	%Iry��y�H�0�Cr�qz�6�<z�{��:/�Z'G i�����V�������hJ��~8=��8��Z�ə��@�j�eV��F�)lC��'�� ���z��M<����2�cP�A-���YH.u�]�;�4bT���#䶯���NKf�Y�N�3S7�1h���*�f�"N���q]f8��l����!��E:N��vQtF����0�X]���~ U�.�`����#�Q�?�`��c�G���ư�IS�\��0��ȼ�W����D�R��:���U��Z�8�`��f�$��y._:�ZYY���DR�:��Y@�AP� ��C��gRL�q3u��&���_����%F}Uk�����of�m��>\`^z�*i?�h���0�گbJ�s�l��G��#~�&�dN�j�R�h�	O��mM�X�G�쓰��.]?�>t�6x淋�R(u9xѤ��L�S�x�9������U z��X�/3Hi$���Q���i(8>�b2?3D�ڐ��H[�+��8 `-�&���6$t�i3��Pz��_=6���g�Ά���1���:Fj�Ժ�žKg���F��/L���0ۍz�ۅZ��uG�V�Ml޻a~$q�3ɪ�̸/���d�jM���:�q=��$�`(S���<�w���V�C�0�.��v���3�5k�$%�����w�<��b�Z6����s`H�߰ 穓�{�%�Rt��0[�/�	���]��8��G	����^}���r�x�JW��z��J&#{���?�J=V�a�q�H�?��P�L��fT�+W� e�9-1a0�;u��y�5����ǰKj$(�"Ѱ4{"��������&a4)�}đUK��߃qu�α�L���Ԋ%h�����=I8r�7�f���ߛj�KB�L�.�?5D��GG�Aڕ5��ԍa��`M���´���%��'�v��,���aI�n���Ȧˠ_{��YC�$&&R�xР~<N�B��sC���R����{z^�X�3`-�ibB�����<�ړi�[ m0f��ç�0JY�e=#�ļN��u�q�^�6i�\_��V��!��D�I�ϋ1�q�}�^:"l0$��*���6�C����/i�.�l�}a0�e�dL�e��gq��r����9WS?Ӄ\1����[�y����(�[Nc$\1�KuM	g9:�pJa�&�ɦh�Z["�vo���Yޡ:<'|�Q�Z�c!��\����~u��� ��=����ϭ!_����~�0��4ܡY+�s{�sP҉�RR��k4��:�9|DS�dټK������ D���8�D��tP�b8��'6���
{���w�Ρ�N�+@7u�⦎O|>��N�c-<1$���H{F����XxB�?q���X1�ݪ�@.u��t���ޞ��~�_�X���|��\@����4m(�z���U牀�P�I�rf+�n1�A�>�5�V��#ȿ�j��������f��p7]�k���Y�j�����c�}8�y9W0���&�6���8����`m��lv��M�6+����F7�O�X�F~m0��l,�X�.�7��uĕ�����t��6���lD��Q%d�����k�Ä����}��`�\�eX��D+�I�Q�?

Q=<��.���=�(cf*FXP�?�`agl8t8�$�]�u�67��N�x�rsr�Ր��R�qt?��=Cp�t�����v����g���%�����ǚ�`����N�H[t��#?I|��T�bB0���U�A~4ܺ�"����,�x�G�_��$9��|�JC_�V�i��p�xl��!(��s�h��hk�Z���0E}�x���k�͸����Z�ܠ�n�C�z�����u��H}!�Z�خ���7wQ��r,���:��m�v:���zƞ����%��=@$�?ձ��������t��	����SEH����b=�;�k��];�hCN�n�����2Jdq�#��?!�LG��~�Z��>=�����m�"��Vմo�d?���^:�9� 2�j������"�md*4�!C�}���ER/]+��U�����j��~�j�ڗV�YWY�k��#j��F^PRI0O@A�]��Jt���$=�����!vU*׿%�����$�}���y)���MB3�W�#TIf� ��yhQ/��I��m�2������pq(�x8�������d����M�T�R,����TC4�Ǭ8���;`�3��N��'۔d��Y�,�޵�=�=B�!�u��AM�F�w/��k�HS�'�N,�M���U�r��:���mp�lI>�������)H4f�P����ܱ8b�Qj�%����3��/M���j�<-�ytⴗ�;���6aj�Μ��Qҋ�05BPL5�4�s�N���O����IM�Igȅ|�A�[P.���ݶx5v��E��TEo��x���]#r�[�4&��O&�ۀM�Ө�%�'��uG���=+��I�dz�!�q�H�R)�G+-�X/�U�)Bv����𝩝���$.oV���Q���c<��`T�'�7�5�,��j�*E�Ȅ$�P�3�js:�H*��c3�BA�AǏ5�k�׶���EI���t.M,�����/ɸ�~tǔL�=��;�
�z�8.�H�b�.䧑fBSQ�>�.Q��,"��+��G�1��B����݈A���}����*�uT�Y�8��z�hhɍC'-v�+(����ܢ��0\�?E��я���8L���"�ߊ\a��,�ܩ��HKPA��o����5��P�YM3�[���+up��F2YT�Z,k�����ƂL�l�*Q��
���,v^+)1w�*M�q�����F����7�g��Z��|�k��:TX���	yYD�6^�UR�3��CM��'-�8,?_����{r�.8���� ƅ�T�?�H�HfV�40	��c�a;�^0�8���@���]�8�f���i�o�~2ss#Ҁt+�*G�.���Fk��\)\�9�d��ݢ�H)bpwxAGV�(�x��F!��Jpvg��[����&���6��67���@w��ZWM`�\+3 -�k��*��OVKH��1������K)�Ly��w��YHETX�K75Mh4��T�R,4�ȚTh����B(VtS�-�4t2�Z�<�E�iL����(������� ?�k���Sl}���T����W�u���RU`����AI��J�+�ᖘ�Nk��5�~�g�Q{DǺ.�M��t$� �Щ;}�ud�>����Ӱ����nMQ���U��V5ˊڭ:�R�̮���Q�y���K����t+Ǔ�Q_�����P�ꑓ\27��0Y'��3����ޠ�]���+��zʯ�>�-�/��\���4d�/9��v��T�H�)�����^�p�z��>2� u����n�&���o��k�D�ӭs��|Q���Wɥ���<5e+g���vԭ�u��3�"(�{�qg<�ò��^�����:��������ݤS�QV���P2���q��.��kv��ᙕ��on^�&�X3,�)�N�45�ܥQ��|����Z��� �E��a|z0Ȍ���T\��ץ(�
_�/ߗ9��a�o*'�I�-MzkWq�b|L|y�%�bK��[*:��=QN�w�U�"
ˍ��s�bc�G��:\����\����g�ޅ�t�{L�*Zm:]�$P��۷)\�S�A"�s�d*�&�X'V�<4�p��on�M�S%��;�Â7Xp��\D�Iط	�A���;�IՎ 6������{]�4<U�)�,�JS����mg�[��K"$o�tc���f�ɵP�V=�)j���<��P�"�L'�ծs�8T���3(��@˙-V`�7��0\�\ k
�܆�U����K�|.	Pp���(��j�\,֗� F�X�l�vY�KA�h���L'6'n}3&�Bǐ�{#w#{�1U�;Tc��F�?Mx�T�n�o���Fs=U���� � L���.��Uv����P��E���3�Ö�������˨S�V��'(�C3��u��v�>uŹPe"�-$˸'_/X��_��,j_5~���h��d�>D*�>����l�lp�wI�V����b:�q���qĬ�@*�*�M%��1 <6hNޓ��/�� �#m��Z�>I�(T�@�OB�4X��E�^�����`�_��h�~-� ����N>R�x�A%�eG�\��b�-e�R�HEν	G|����aL �F
��q�F�:�2���ݴd�6[Zً^t�ٹ�[�2�ޫ��PL1J!(-�:#YeWv�8�ɋ4�=�@~`W�b��*�\��`�1���l�s����Ԙ�c��]�o���AT,������� IY�S�j��^\���9�qt(o�I:�j�t��!Y:�lA'�E*y {���1����{�����%�"�WH��t/�1٘S�ʤ*�.?��NvM0u$�lv��0�A��R"~늡&�QG�&&��O������F�u�W����d��"�N�Gz�3:��������0]��^>b�k���U*�J�\����ڢ��ħ��s��=����:s�d����s�?:a�k4 ��g�f���p�D���i���̰�E��I����f�����i�[�Gzn_� �}i� ��p�F	4��8���3~�5׈��Kg۔��P��y?S��J���:"?����A5:|�K�'��
Z�0 0z{ڳ�C�A��yDf��?������"}9.#/6��8L�Nxi�hJң������$C���I��[����3������歇s5�����d�_��M`���(��j�0s�
�lې�-}8'a���._�ㅪ���ƤKI���+�J�Z�g�AԷcBD����u����d���(���&�;��ǔ���!nӫl;���cArh V����<�}�>)�kܝ7�u$�E���ʊ]�zX����|��?$&��Ou�vv�2�若����TE��c�F�d!�\��8�`�;jJ4>2.W>qj���D)���b;	�)޼�{���S��I,�|�*M¹ϐ��Gn�!�4�lB����X��?��M^w(\����<��f&���[��I�$۶��e�������
޵�r�L���\,���������s����������w8G���k�·�LJ���(�a7�C��
�.��'r#wR8�����Đu�,T��Ha%Yt �c3�y�a\��!փ���U�^몟�7��#��G���p����� �i�\ 6%h�m��^>S?��SE����t�8z���
A�Âlo^HVUЕ��zve%�7�j,�N�(��Bƙ�2���*��E���9�-����Y�2@Y���Ȱ `NZj�f(2��5���Y���t.�������a��V���ș�A�v3T0f}��f{sk͵�:�=Z�W%˫��+��' s�\��5��汒����`]�kx�땣������ӽ���g�[��,$��'��$0�	ȿ�P�����]���^�6!n�0j�#�8,�KO���}q x��u� ��t��^�ɿe��c�(�U��o��vc{Mpi��p/�B��J%Q�,����"
p��i �t�x�$~Ϭ/�E� z���Qoc�X,^�_�i���4E�����ۍ�{P��&VyNa�D߸�v���v�	6��I�{��*���V�i��y�]�/��B�Ñ�k�����MUo�k
��Ǥ`B��)�H=8�u��F�u�*�V.��?C5�Xz0�2u����?��ˉq1׆Q�A�tY�*%����5�[8⎅.���K�R�ع6h�0,��' �#Ib��6�#��ī�ioI@Y=F�K���w�mT%�b!H#=�ȼ��jO0��38n��ѷ���	�T�T3&�$����M�"��%�ʏ����}r�F�� ]��R�	�_������������xi�4���ο��,M 9��O�_�	x���*b����,9AG����]��dP��E�+"��-���uy��?�����R$FIk�6���oK�+�>*�!���jY��&ӥG���ӛk����]�٦4)�V�X"���su�O.*Z���E�e��󫤧8Q`�U��q��KW&JF"���'������E����9kv�u�����l��!�&L�!	��!M�V�9qC��u��.�M_E��9m��B��W���ˊG&��I`Z��p����T$��SԈ�������H+40I]*����9w/��=��U�[�On�z���A�1͆�n;����|�F���F N�m9��A�P���5��4�ݤE��'e|��� �*��5P�޿�[�$$�!B�@��P��fG��JR���W[�s�g��4�jT�zo��^9N��K�nz���l��\7��Z|{|]���h���."�V����W�Nm�÷�/�t��
�`���s]�o.,kɐ>�P쨽oǻx��gaN!�ْ���ǔ����L���`����?��3Մи[h�Z�B�� \>��0��)�q��{ҧ!#��U��+-�n.�Q�#-A��,N0�oRN���tu�]}���@a��tΓ�)d���,�P���3�"� >�q���5�_d���.�Q�%����ނ�п�w=-�W���漍tGRf�;1ݲܥ����
RF�r%�B����k�K���@�j�B��A�eb�HC;������2�G�n����Jԉ�e���Sx/�-#"O�B��ܡ�9�pvH��:��
a/_F-��,,�w�!窅��-�wA��a��n�! AB�:���D��3#���c3)�Mk�]�$0s�`�L .���i<��5��Q��r���L?�xfTiH���y�k^�9�{�.�B����X�S��s���w�^pk�6�>��˔jn�.T�5W�/�(1Ԥ��Ҫ�˵)������%T�Ѯ�0i��-������$�7jC���ص!�=�U�&�Zz���S�ǉ�ԧ�p��]�IԎ�e����
�KF��(+��,	 �:����A�5�kҩt��`�K4g�'U؎��a��H(��e$Rsy0]��`s�,�tؑRQ�i1���������:}�#�v���J_���#�eHmEs�u���@��Ƶ�	p��9X��r�-Ygo���c��˭*Oz� ��&�V\��L^�k�< a�t���B�2'I{q�m;
Ѓ3� ����Py��60)�5��)�9j�*��wZ�t��Kl�Z��a ��9�O���R_�tL�	�*!���d����}�T�a����>`ފ"j��C�%',�F�f}��Ü��`�v�'�q盉��6r��g-w�#P���#G t�17��v�v���ǫ�h�b��zl-;�]��9TE�Y��R���S����[��ܬ���l��?;��;�_I��C�28������U��m��r��������s���H��R���7ǯ��[�Ε��Z5we���,ֳ^M�~����!�#?d�[@�\�a~�gS?�f^���p1����	E�Β	0=��'��}Tֆ�x����hqz��`n[� \��6� �
��F&]�ᰗ@���%�M{�o�Ћ�'&D�,��(�ۓ���.�#ד���4�MGP���6CjPɵ�;�p�in��$gS1��_��1�ě�S�4��٠�����{��Fԏ)���kI?������s�N�p\n��M'_��ӯ`T�E�ZZ������̠�vM��:׾u����U�#Y�0le B�e��.�g`��Pm!%p̋\�$����s���<�؇q/����gI���f��1���Fb���[��.t�@V)+L���R�AÔ�/T~~Ve'�0#id�l&P�M~B��ѲV({8*eGRL8ݍ�c��؛.�ˡ�U�'���J�O�a���2kT���|��%�O��Ux:w��[��/�d7���hߩ#�I6��Y\�b����{�"c71>�^'���/�ڋ*H�D����	Q8��8	����o䎦)����vzD5�DG �63/��ҥ�D�lR�����M�>��p����eF~�J���H���{��X49����A-�@ý��S����S贆��"oň�p��[���X�=K��V�9x�۩e��x����Tͤ�=���-�7�"���#	���[׎��RX�M��H�/N�>E��*�FfwFJL(@M֍�t6���:�o�M�$���!���+��
 �C�<�h�	�`���nbO,^���}{�E�|��@?�#�M�1(�Q�L�O	�1()z#a� _��d~�i�� 	����"`�_��.'��ߠ�6I7�r�g�vv�C�S��^*����l��1�I���ioՊ8��fok����m�`��@4?�d$�I���]���6���
��ܯ�6g��%/�\J�#qO�VH>U��A�o�*��L3lM���e_��hݬ�J��C9���:����`�T]��o|.�U︿�f�Z��]1'�?;'��������2��^���Ä+��3�v�s1 k����N�eF���)��\��C��G�əƮ){�0�k:�ʈ�(Pp�\�2O1܉�������g{P �oFbu̝LL�$����89��%׫wo���mY 9���Uz}d��:fy5�i�|6���B��g��Z|$�(#AA.���C��-�Gtr�|����i���4$o*��h�͂D�׮��9��x�rWonZ(%Ԩ���<���{ǔ������AA���)EU�QG����.g��!�W
b���0�A?��7���x���܂N\����&���wO2f�4I�E�;����1�J��*�UYIvLW�|�u�G\!�� ����ZT�N�/�*�<�=NRv:y����
�Y̥�׵�}`��8�ٜ�g�"�����.�"��v��c�vJ�o��ݍk��4��P��k�!�����۾�=������h]wQ�	@�8޸������|�۶���+3x�p^g�+�bR� ������[����K�e��6�R(�C�i.���/��l/;uP���j&��y/x�H��[q_	��+ڮ!�R��,��a�5�y��;H��>V/9��T�ÌC�;�E�N/�A;����Y�G]A"�^%��PL5Hd=z�ZB.y�9�.?��z����2��˟I0<�{R�D��'���o���E�^k��Z-I�v �R]`�,�tJ��VagA:�k���hz���kc�����8BB n@`�7�'^Y�ِf������_l8�Γ�	򼖊]��e���U;����w��qqpUX1>��By��#�ߏIr�c���	���3�Π	�@����T��Qzӽn�i�PP�w��>[���9�Y�tr]�Qgh^�>�+����yWT�KH�p_��,A�m�dݦ�3,��M�C�g+t9*���G����_�	>V�*����w
P�qZ��-��T��Y�ZWU;<���q�[c�Ҍ����%r�W�J6#a[�{S�-�z�=dկ���:ՙm�v��6��������xDKR1NA��'\q�v� 4K���Ƞ�� ���ĩ&:qkb���8����o�HT�&}��־kM��X��DwH�s��H��Y�*�_����8����p!��WZ�AK�\6�dQO�����:���W�}�I3!t~V���.;�I�D:fcX�E�~�x�F�����tmӬ'����״�\��A�90�1<����UE�k3���R�Bd�<V$ƥ�qBCo�sR��aC60�f��.�{�t���"����}��˝��N|��O�zK���0��@�Ͼ��)�������:��9E���!rg���R��5��*&�-~�ğ�Ѯ�s6�;�&�?i�����~>�o�ʮ�W�t�q���$;|Y�V��nR7�y�$�T<���5e8� �$5v�xDk�A6�L\����9��F1���)�*��1yba؅�Bmr4?�W!n�=�İ*-r�Ap\�/�Ld��x� �q�H���$)ʹM�m2NaJ)u[a�+��4Kj+};�j�4}s�`�-���玑��G�������|/l��h����f�h�har[�d��l�"ԢbM�)bͰejI����
�n��U\*�"���`�:&��C1	A�<�q��q��3Q �0�3X�ŉ9/�@s�^r{����$�եk�9"M3����T�L�h��.��?�S�Y�Og�����J~�ƪk����|�Ёȍ��C�kR{p��S80��S��V�I���M��<�X;��^J�C��D�����8�e���N�T��ӝK,��+g��{���r��1
����\�(B��؝Ƣ~�� W�e�?G2�SxXN��mu���D���A˝�ȌT��y�&�T�`�~���G%����3��v�AGB��il���1{I�.d�x8��>�C�w�>	�脱9��ׅn�JAi;2&�|h�0�����6�l>@�2�D��Y���,��������t�?ܻ,F*�ͤ�(�D�ktIΔ�}�S�v,X<yj@��D��p���/���9�@��l3}޹�폲E]��4EOW��a�j���
<�F���d9b�ф昆�LxI�/?-ׇ55���骳�������B�N+��+0돹�a@;W��=���v�g��ÞR���D�s�X�B���h�	��*�k�EHnkTGy� ;���s=e؍</.�]��o�M����#����:����"�7���i�r`n�_���W��G3P.r���Vz+[1#мϱ`���|�qY,�o{dA]As�^P����=Rm6gq%�ˡ��Pr0��=2z,2ÉA}�����
�~��������M������B`�?1B�y�nbۿ�ӢN?얞y7����é;������Q%nGݲ��n�����BK�vT�eQ�s��Y�Qqj,��徼�1x��?A9��L�=�A=2$�f�r�����
T�};����d�������(��{�) �*�F+E�	Ԍ����]�}���L95Ҹ��ַ��]L��s6#g�ݳª�%iv��\<�`]5��!���_�7�I���[N�l�
�G�6�`ۺ�s^��qjЄ�\h#3BB�=�[7�bD�jS���Y←v5��:߄{f��6P���-4~����`,7�A���7�j\4���BL�	�A8�nFR0e��� �Ȉ ���*ǀja=�|�˶�*�1N�Մ�N��J8���,rϪ��x}�Kp�zn�