`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bRqgFPHy3CKSpQy1pNoxHjkQd41BqQYO9zoEqxfTgWXq5QJnJIKr6wHowqwXN5tCyhGG/UOv4eOp
sMImSPfCvhkv01vIc4P7/3QeJi/qDENrvb58VcAzBU02DB4z1u5bb0sspOUMDQIecEReDqE++pSq
xccU7Ir0wD03U6XjP3045f6qywyVrW4rM+ClDGAjX9oYmZgpScgCwARKJsZnjGOwO+7mBnMrsgtW
Scv4WymYB0mc3RLpAln0wyfFBAU36gMqxJ2MgAWnD2QAhT/2bS+2cjg6s3FCt4Gll9cWzUcS1Qqv
2cgXZ/t39n2TUShG2KLAFRAgD6QVQFGsg2xrbg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
3/78nZiwpBdfv++opJV79E9wDVBA06lQr6qCpc7nsq3bUeUnnYWWlG6c67nWCwf0tBwlx5HJczQV
HqQZ9JCTAviCh9tp6CmHxobxviApheM3l5r8VWd3mhg3/hjGP6oN5+AYmaJoRkY36fn0W8uRrVMs
OSr2ZVBzs/3wENjtRgrLqRkHzSDQXmmElaM1lFUvdSSL+ETTyYHsdD7lWw41CKX5shJloNTBi8iQ
5iuu7oBQg0/v2jKvWzQmzoyct0w0FbZ1xDosnJCzPdLudPoPYfYuYm4G8I80Cl1NvuweYHJptWG1
b+0D0zFxa2atLr3giXkqZUCSxVh9dy6dG25ZEus3H/3T5cj+DqaBX+BlVk6eINRNV/giufgJx8SI
b4bRA22anszSawQ3MKGa9uyb4Kr9lnKFOr0zIO75+XloveZIF7jvzfseAJ2SFX+J7HmM4DPLq04p
MK88kouHOh2XgP2OADHU2dXZvodq13rLigQn/MG67nW2wPevsua8CHc6ZC/Jp1EJBMHiaCNT6Ucq
/ck/mS5+UbFlD3uXuo8j6m4+7pyjvJy4qk9y7TU7xoj0PlfJ9GfhFvQ6u7/srq8UENjzondtnZ4M
SMF0eTJwFBWXQzFGe3fDnV/9L8sgHcId6tpy+TVLgxhR/zAKy/vf1fY02fu6QNoITqMIlaTGp1ur
vwp76iEaQH87VrFUJtD7F7KV4BUvwrnVfwk4NphiYJY5UzF0Y4y4is+PfLwuQgmWsETQb4Ewx5YI
oQyYDms6jX+u+UhYcdVyRnltNVJekAPE3EfvYYnYKT8/2FQLcTrBKFzdNerEDO873Wz6TG2L1ph1
ElPYyFC/ud9zorslfEPoT2F3pFPS1ZnFqMF3LQdi0myiN7GKYRUxYgtvDLCNwyDsHVMvy1eAZayY
mdXQ6JGuz6d7UbyaJXDV21P59cbKLywPB9rMmf+IEB/OkEYOBQVpFb3T+vVxdOs4nrVEsuybAqVo
cIxMdspbLMOlIhsH4exqmXCXYgGSxo9YSrvKBjVno4Q0iOv7gUBzLHM+eoQLHBxI2xrObx25rASi
A+H5/M7VYyjAnGgCl+debfzElA2Bha6xmqUrn7KCXErkRPmOenZPnD5/m3m92rZwU+ndF77WNXhW
p64Hc138sCdrPZ6OEKi/eUo1jONE1xC8SDmu9rn8oYoy8Pa2x756V+VW3n5KbzmOeNZ4zZWYhY4d
d8C0q6De9ICKZzGxtyAnvhisM3I5OsNFKcWC/dUP2Krk1Ih5iSAJIFqwZi3jZC0JBybQo+/lo135
8z89DQYEbDQy2OTzKULTCHOEAjJOtoMY9GzhqCtwDwaX9+ubvrj1DKm4k+ehuMPXhkqPtUhlbdtq
OKFpioDK3I8gW2sxbpW8bmnCzZVhdp+bPZTHNvrW4jdNQFnV3qaFVk3uOZ2hm+URwDhom+3LjREP
76xYhEJceeedzybBt08C4RrAf1h3l0ClAssyFxVmP2d0qhlgQHUfUFdThObTlzTqVl5Y7X7EIbov
E19nSf8SC0X1N3XcYMVmm7m8XWS2doyKxRcWApgqjPr6RF3EjQl4eCxKQQy49Kga9hCJ5SY1vY3V
wnNrJwQEXVMqp2OCFaz/m0vAgBy5O3af4yrvL5reR9aKKMJq81qjmmwIQHfBcHukEQEYdHYSYzaT
OzPmSJCfqbWQ6qBaxzJWTz/Qj7BH/6Qr1r7vjrHB3vYAeatJpbciEVmID5cNC1eKJ0RO9+JS5rHi
scYqAf7IwZVEUuulJexKVitDqF9JDPOSzw3Zp+EY0mJEmP65kH48VBJZfYNonF7TewpYoN1n7phm
mOxTimeTn89TWE3++AgVRMWKIZxSkiQevLdid3j3oCWKAM23MroCNJ74x8RFpQ/sDWTzfXJ5vhWB
JPisnKqtJbUjz3eNNVEWx7iYOd3Xye2U3kKWXcvSgRHFbdNv72uQebg+shHlxtl4Jm9yG4LrMrU1
nbWAyEWt52fPVXkOZ/xHSYFccoLAYQJDvphPc527Rgt4JnXc7PJdEJYHs4k2lfd17eKkbSonuZhm
MwvUrvGxENgvLs+AUzJ4v3VJcIPHoaqikuzZo6EKbOCyYhIn7CKadektOTHPrU1XonpkWRPE9tD4
ti8/Q2VwHKm/i1MwmcOSaUFzqpp8hQawNkvh5l1JuT0uFR5G+jD+P9lbH5sWgRomfToh9ft9cHpz
jVQYKdSyC0H3N1bt/eLfWd5kGP24Fh9L7PdFuKIsMkS6tGG+iG9m+UymBs0XvtGGEdDIO9XIQLDM
BnaMTWqVyOrbiiz2vW0WsgE91DlOMrkFI3LVqk2U6yFijZkIo86Ohe3ynUkZETuRWkhHEx5CLcUK
im+zDu5pob8/VMIjjcq/UffNVcdmclveKk+NKsrizE04LJKw+xQk97RaiEQdqoubZuBqe6XmHs7G
Q8f1/LLZJAvD9YfgLWZv+O1vZLRYx5Sh5U/44+fO9jL/Nxqi/Sad9qxqfd8JQO688lNw3OKTpSIC
oL7Rjtiu/8CMSnTxVRr2eyEw1Y1D18MasBLt5cHFBQbMnVYAjg6fGLBA/+PiJXRD/TRxyE682Pn+
OcZQVG5iZa/Bfaoey3aAUj8DRAyORxpo2TnNH30yzvsI/ux+gwhlxFz9tcULq+cQVC5OY8VL/Ux4
x/ihw3iUFgzZOpGbqTObl7GV/YwtyadtS4UFTSlW072RN1eplcL3fUXUIpatYVzojsCEzw318p+a
wF1QBcOhDxSkwrEaeP6q3gTXOIqvhFbz8acq3+NV36pVkUrKbP40qjfywcOrKLYuZYT0F6qCeaDi
gWrE37ha04ros1DYX4+Da93QFxbf7l4tD3Y/p6p79EpswIxnMUDcxFGBUSo996m0kNN358giyn5R
R66+QrXymcGCFLuWZsv4Guyuz+4ox+NmCzPfDWVhKNIoDey0UexfhoOM/s06RkUv+QiV3/Vw2P9p
6aL56AjHWFtub8B4bpbu/9oKVqdk/JatNJH3VcKzxLQD7ViQd0chxeTziJ1uWUX+c5DcyaYjcHSU
wG0xpslzOLB+VTzNlgF4y69QAPzeh/vRLoOIeiBebbInKI4SXFFyz1i3XtqmhBdwpzqLKkqrA3Uz
8jVUUlLTWZFys7xh4jbzpLNAtDDsbpSBun+PEt9CDY3sIZ+Ck/LJzYtXS6YrjLnCihKsVrHBa8O6
0xsOUlVtZmzpxtwY8Vq85CdlnOCpbOVWKhMU9ASsrzY+l80sJDlL24w0JaFJTZoE99Q/rRMQxxfE
xfLb/5Pzkptg3DZOwUIY9Lf7FuhjAGDKKDct+TOqhhvLHmopEq/6dLagkzXW38pjygQO9tyiFOCY
N7kthmVQdh44ToVNCQhgJNgnQUj/7+azgr6Znlc1FWBifna+X/a9tmk3bHiJU7bBTejz4rlwsvsv
wToWKGcWSNC1RwsdaIs0j7LQPTR4KEWK3ecotE0MzpiWOgw7h945BdzXHFplERFRH8rAnPt/626P
zVX3tD02AeoXvs+mYHUbV+cxUmCdiZcPlZ4dzKiYVJNrCqXVGhZe/c2pJy77gSFvyAQaP6jJAFFE
ZhoZ19wzi7OMrk3QxfmQacV9ROfakeTG+WIPRha/bVNgaRsWHHCEUxOl3joFpBC7efnu/wHrokmJ
5xC6cAVEVyADdvj2CfBERptDg63KWWxP4G75rG7zH/zKOG/fzAfbx6FjvLO3CC/WI5kHU1lCD+nV
ukLov5970avgwnLWLDZr1MPC/2woO48yxq0msm9BYeKqRCU/CQAJGntG3NyJIMkjI1il1CvzcG0/
OP8YxYscrn0J3dNAKqcm8dtJgmRlkM+1xcmd5U0KO5cs+oZMWNnR3Y2bsfXDDn+/sqeyi+vYNY65
/jL1emLTXDPDG7R8qaC6SVqxI7KcwzL/r6VJQvm61knQ7DtVVraz1jGZANWT4y+2oem9gY3CJjeO
YmY6TGZMK9pr0+Z2ssys3/UhFgS3DUj+u5/OXcOZzjohNh/irtIXVitZLM2nmcfJX/JWXJfLvq/i
tt7bqhNFGfnqMbjHrdcqxMznS3SqrQHndRa1HtPHLqymAkqTEAdTsWAuFreU0ZEZUyNLg8k95Fjb
jhd9a5lYNSYL/RenrDvOnE3Zsv5tG5yolfYOqNfsQEdU4V0wu7/1ZWA8KYBYn5nzORJ+s9guBK/f
b5dSupDnSKUbJaszULfLaKUxr37rR5FOOGoVD5Nv2vNynYhzYa84UL7L/swuUhU5oqb/OFurXsvE
hCetZ3gDZdyyKTsSNgnUByTKuUC/mfI4oJjpK8qRgY5SyPkAeppPBkqcwvIXKlOqgMGKZ/Br/YQ+
pm4MbJzvsvpcQHGPhCVDGD89Pu3pAhfZ0L/Xiz5fA7qdCPZzxSe0gyuMvjEnS4fM+WYWjiTCby8v
L3d/EC3dI+kUMjMjsGo/509fdkX63HxB57vM3jZle2pQMlu7WR+lIkyM20gKURjQLUcJ7rt2f7Wl
yDhzu8vTJKpnhUahuP4HGegKvml2XQ6vL80lUbwjdQI2/TXBN1LOnGdHyooELSywRPxzUuxWToYD
de8pqvFrdAxspJD/JEFt0KrWtCgZ1y9dc0YaNXMCPn83xIbd45sDqH4E7ww8g2djMdAuzbBr089f
rHnAMjp3ZssYS/K1VsVrFHLPQ5gS1T2Y5PmSTZDeOFAM4iInjSOMPRrCt4ITtQsvURuFxQCAVFuJ
WghPXKabEJ/wKYLhH5duzutsulaBObeEyU4G76NLHxraLKFYZ6761mtbKYaCBlngN9PwgP5rxAhG
9XnuxTIGeHzZQiv0MPpsKBRzcID9iphJRp3xdyRBRAGGJ/AYRwdRqKN/0o/oNDZeXWthYE5r0w6O
+JHYoY9dYXaRs4f7JqOsvN62d3D8pJVzp0jgEAQBLnLE+ZFh5poJA3cWgbWZL6LFpNB9OqlZvX/H
DUpyd9BlnVYzRRWF406D2fBO2sOaYQ0YdVkRvlik0klNHa1xMnkj5cLciIvZxFqBwbrB1Tfo1rL1
vcW7o1Lnpo4R3J6sE1SO55J9mmLpdNHU/QstXqQZMiCvjS/lW1u+btq28iOGKmcKi4B6AIkGpxky
DFL2zDSZtO0KarAHvfUTC6rqj9HRQA2WHw5IBCgPKBn9UmPJkt3CWGMKENgAuu/y24H+UBZi4LYa
ic4qgsEWYLTR0DS3BwXcJIrbS2qgRF7+cti8wXTgbhlp3ytWxKTwSNOUyecAaS/MRnVfhXrOJ0E1
tyAN3fkawmctc3iDLhJXPEJNMeMrf9GkeYGZfNiemdtp8hqjXuez0gnXEgiyddakwF77D/VatY26
c3xVBEC5BSDEseY70K/3V6HpbjuBaWbYQM91/s2mEbXLRrnrt4R27R/BFAQpTpHqKZAmFPn656M/
gS/YFnesx8xZf2eFlF6DUjOB8H+jBDVEyLJ9kH/D1JBR2899s4S7Bu5d5OIWlGfJHCrTh5zPQJFB
BtLgCvTjxBUgY/yYWNrlJfeFpc6sUNvJcchQon6KqX5pG+bcBmBiXkKdhknHpAkhy/lxA7ANsopx
AGktui7mL05aZ7CHfNgGt51qId29PXm4GSPnXwld9aw00EFXOaAjGph8YdpE06pMslHUi2f3w3YJ
5VV5txUFtez1e3yTckVUgDLWoRaOvl+dqfYUKY8Wllcau5Gs0rJjEKsuchEJyAFAFx+recymEUiG
qmhH+cZfHuqnrSMAdy7Lv81zP3He52YqzP2e1wxr7Ve1lnHdpW1D8tx94BsgrnHC1Ta9M/4Xkmm2
M42jmywP2z4rCR8p4wSk3TJyTS/i3iMP2aitgbpnRoEQ+c1z2N1NdZ9u5rQ2d9jgdJvEWex49EcS
PIwfsZS0mbE2mFGkj4zVbJ3XIsQe0oVWJgwpddDypXrFct2Gver8sRWxihlJMBdgUPqyPremxOa9
Y0hSLcBiU9XCpMy18XfefObFg/TVy2CH8Mh8XFvKSW/JJt4b2KU5CNCOthV7OaXXH7MRSgvTMel1
r7LDoZef52kLbQVr+jjOTspvNlbwnxro6t/2PcZ+DIFtZv3ZXeHZMKh70BhS9u187F0u9BNu4otE
XW30jhEB/yAZwgLHdW2DEWXKgudyjAK+GkmyecdMqRu5Hi3wZYR9CHheESDupvHzylHRsw5SClWS
eslE3vmDV/b8rU84rbeDf3kcxzDpJMv9qKRbD7yTnN1LcaIKbcs3Ub7Cpsk3WdirvpDgnzTh/5+a
ljCypMn3a3f/fvA01kgS23Si+WzOZ/316s/JW6JcBbJDqGfyUNMzQegO19KEN/8bPGQAme0ZMUR9
7At8HfItsTYjeGtoMtB02u2r6K+KYDvYpL2vI0aBNzRqtHcjyGWBZW+Eb7a2+pF10XlN7QKbmC/G
USFWeFTjXp2nzs+tYsoMzkLNxRLt3sysaIIqswLNDM1BWJ4LzOhx5hLk4OUSCUVfM8ZxU2DPR76N
42XLSmXI6dTlUO5mQ74UKQ7CrdshI6pWSbycPTVh/wirzUCaPB+WR9otQZ8moLpIO0DGyQNuWEQg
xIajxEcSTMIRZMLbNIMaZkkVEhW8bFhZciLnv2P3mvImtmNtgcf7Upm9mYt46LAa8Cps3DyqSRzO
jvOFIWWiid605IvCXNK2RJ4yQdKJyFqIRpHDIIRcu9LXxWjgg0DB2QhsEjD15L53uz9T8zFvrxEq
5sOMSm32wiZBLcGxiJQKgeDDPp6H+tkszs0nF13nINrk2BQBG74diXu2cB7HiV/H6p88c3ZCNReJ
KOjOQJ2gXPhw4/1CGTCtV+0QWkaFS1W/Q1sQHG7ktH5X5tOW2K7BJN/JX6in1ELIDqJXuuYoSCOX
szHHIwatMfQFE3PHGS3M/5PYMMoWA2dcf1RQZ8G4pxNMip9RHAJ9W52lOrvufc7Y4aqrBxR7Ru83
CflvMhWuESahqSTkEeQjsLCkXtx2YO+FZkmtP/JRs3H2++Yei3cJQU1ebmuVZxQK4WBqHgc2/Fqe
PFO1izMrSFKbzLACO+auxnRLJ1QSsEPHA+QZ3PY9OQW1j+0xk3CdlqJEP54vrwZ+HM360Q2hFGxa
372XPyHt7IyGie6TXQwFC4Jx9dmjKlJJ1WKVbaE6fmdvWGifXk6UyeF56/BvkX5DTzKxZ2Uh/xW5
MvSYNeS+qy4gLi3kmSJPFASf/kdSn3j9oIqJgIY8zXzE7jGpBZ41RCMcoeBp5QwagvmWsQAFU1WQ
hQegtMVnUufGXeUAQq7n634d4wLzXSC3ICcub8x/5Z/KyUeqxlqp03oryg4+sDoqPbP7bdDr3Gw3
O99+DK+gWV6q1FYV548FQSS7wdLvbsnjEiqhPLXy7ZJjZfV0RuPLq3tqyLvOBEvmVSMBimsF71lI
nJ8BnXp9PZUJYKCj43QZUZ7hsuZ6J1ugxpjJ+ll8ozeZktsoPpHi5w96KQfsI5RFXEo68T6/YppL
6tBHsYCnPplWIUe9cs5PGuLReFpXZcPv1sxCytF/DkZRMHOQRQEj6aSODzH2mbCm2xHCtSIsOSpx
/wwCPw8eVSRVNdk3XjBt4J6nnw8XU00gIW2Rcact3QVtT2noowkrEkfV52i5B9z1WBQgTXnPsYDX
PUTj9v5HL9zXu0NjwpJor6TVpkim8U2SgIeKBlnZBJK3rTMs2Ibv8nZX+ufMLhhD7LXI5HuTyFpY
mV8eG7QE/yf3PKK2eJcS7BO879cj/WhFPl89WkjfyQISzyTmRTCbnkxk2mA1px3eNjIxV365x9MX
6KRZpGIXkJpO7R02d+kZRT14z9hhSi6riVjyinUNe4Ij5akLB8/lVPWCOkLoOOfFVr6CcjfcRfZG
QEJ9BazYKWM9PN3VWBNmSPzRdRmP/+9oksWF/CPSr6xtkbwFXosbknjNyRZPuC4VQ63BCvNmxh36
tEDzj87uc3H8H4KdMLMgCuNCzgTcyqq2z3MPkWLzWBNV2omyM/FQ9F5YEyu9lV25tbmVhoVYgVeo
KiqGkv4jt9+16f8oB57DRsYCjpauFuzJmipV0u4LJbZzGN0bnzpfL6WDOql1Kaseid4q+DOY93+G
eGZO84nSOXh4hMbQDh8jL0Ay1Oo9PigtsKHkInziM43EL7WWLS9LAxaLaYY5M8XMla6zdRxZfDC7
ZmVZptFdowDHZI99Q6z6Qr4WlmIVXetxAMyiE/9rJCKes9tRAvdjqqmEibKSRoYaueHcAFh807V5
6ASMboSPI1A7SlreMfZb9w4toqnu7z9drpQsTvgGnj68AQvIxsyqBipZ+aL3YYjFu+RAcl0uZlfx
b0sz4nWo6Xlu+sVVbI9RAzcm6SMIGFElVsIE110zPYElu0U6NUN4j0V3FeFiT5wBbe2wO+Qeiysl
oGJjdUogHLxwdiCzVRFPjyNs+g7KwPyZZI7+F9oyDEsvFyfHA6vr897eue/tCmOwahCYK1nHcC6r
DQacl6l6OpPHdUlJs9zPEAhM/u4cOTySlZELZHYK4xDUZ/xUnXeWwAa0GO3ZOgQxeJ04/7VlpfmR
1JRpj83fp6VkEWkuXFJMst2VPArMUUC5/funJfMY5RYvX2MngLhVNemHZNAEdEfjeIzQ3RkW9nXV
yL5FuWN5P1pifmyAFblC+iKxSrHBXgeH5AzfpsI0C1gDalziuTclH0okxoyxmXxFc4FKtJVfRqeL
xIpy+ex6/o/x2/vv21sOd1//4eIBO4/5gfrBlYpU0UYidALuR1Lmm6ZK7L0xfVR46Ar/bn2x8fB6
Q2h1/VwkSmUIDuHB3DKHBrHssmDmoLPlWvMUr6rh83BYuutY7MNuRG/b/2k6sfozwE9yb70vEmPS
9QsMC4ut5W6VPftl1dz6iwLUWYEswyCpfmUKVTXdJEBo2ziwa/5CbeUST9z2GU3JPu9HpfaSboR4
kY4qM4T04LoOs6Xlv6ayhILfcO84xz94mbuGTlIXYGbmYanDITnc5KAsyMsJ1WM0E1jalkUxwCfT
l1J2IHZCI9JCOEUg2S1TLgTk0EjPxhMRJ+farApb1h0egvyNbzGavDFaozsv/gjTa65Ob20lB/am
eF+4o1qz9e3iW0hmux7gVOe//cucc2Uq4Nx3NuNp/jij0z/5GenuNWNPEAss0VDq1+1sHLv2qSld
B1hwcqTmp7Ph++u5rElD3es+7w1SO8iAqKzMfWxWOh9G5oa/itDnvUV0EqoaS6i16lxAFpwfMcZj
RfLSSuXx51BDBpfDLo9zapESC/AHDempoXHd/4zJJqF3wX/QUL7AUHZJlPh1p0txgrHVmLNRjDoH
oQj4NKErVfN21T9uiByCRDyOTBzFX+GcQd3gKI8h2dvKHymvAlr80i2N1MFKMxqsguXPQywN2Oeo
64UXOpDkFBqXs/5saFyDpV+iSzD+Rpw4+YSuPnmGTW/Zxwa6ogTi/9gYZJfeVVXS8+pd/oGZV/pM
PR2N1rYRiSUUmqmj9goGLMlcU1Qokc9CV+AD6h3fer6pq+nsc3mDlrqtg8ZrPgopC10m9L5MJbUy
DZSQEZXMu4EDE5UsHQr+9SCDFH/gooxiDzF4yspJCEYEuJM3qN9ILnAFjvRTK5eptsMNbcg6o1C7
ImH27PjA7qTxxkBQEX4p3VbU3rmiU69DRzEIrmWrQ0S+iKdauZZQ/oR2ZDthR1NnNNPlLDm6HqD3
SzveJ9uv1n7GnvqUxCxh4XZpDxhtWha6SC/7Rhb6JMGzW9iJR2UIMsIOrNHtlWGBLcNrT5LcKAQb
aVik51Eg1NaVh0SA+Qy2WJ1+YUJqVupT3tPQ6at11I1rt9nYQPWdEBMUWC5n9qbKBduuQ1V3+Nkz
vdIRSDoycq7JpYus6ufLvuaFXEN71hRZra2bVTcR63ErPNAeSX9Wr37cR0ZabpacS4m7pjo8KkQl
mmInYQE13fMACS6AD3il3KlCIfjJyhPV5RxTr5wy+4Ns/gABtykTr1wfkGZwKqIlZaqokZS58GrR
T5Kk8h4=
`protect end_protected
