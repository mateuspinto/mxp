XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��otpa����3V�v���2�+a�d��6� �Y	���b�E�ѷ�����N��?&���fϕ����;�˲ /P����-��}ޟ�]��f��R
�_��l݅�/��ަ&����H:;v�E�j��yLQ;�e>~e2��2�-AjHʨ9���3X���ń0X(��A&�����`���sx��l8����@���:
�ƃl�R$�	XvJG�"H�b
�|�p:o!���6|�}{�-�V2�Y����ha��%k�u{��k!����#*p'j#�[�������(�z�8$��`��r���==��o�.?tC��?�Ů��=?�Eת�<ջI��j�0�fQ���x�u�����: S����)n2���I	�%qx�<ִ�`��h����['��	��K͇�q^�
	����}����&���y�+���ä����X��|��ZAm�9��`gv�@G��P0|���n��BK�N}#��>�H�1ޭ:Ta�k�Z��~�r=
�U���3z�]�ꗗ��P�׿��j�q?Y�e��O� |;H^�W���s��;�X;��gx���wo��v���^м��̠��u�Pw,�i�^Fk����:��2���a�H�ȁS�r��u��Ν��4q�+>=��J�"{��]������@��s�O`;��E^�B(��^}��B���%"������'� 6s����{� �d*d���	F�׼�|%`�3o��P�R�8��q���)���XlxVHYEB     400     190�H�")��Z�����E�j�ȗ� ��^�mbmnJ��CR�w��h�� �XJ�C��
�#Yw�y "u���;�Y�.sVA[�2�&�UW�D�y�X�KN'\�4M�T՗.��t\���d�Qc�� �����������Z��)[{Ӱ��B���B5��f|���͸��n�JQ���� Pޙ�x:ZdAWM��W�5�Ǌ�/L&�K�"33���&ه��x��p���M����ڣG	F�n"��,W0�l��4����Ċ3�[�a�n�(ˀד]��)M*1΄���?� �HU��1��Q��}����ڙP��%	wu{��F?}x�����J{Q�SɉѦ�CAa��G%�&�T�Vvڡ��g&!���vJd �=Q!	�=%�XlxVHYEB     400     150P�j#�pUs�� q���ؒ�˶�β���;��	�5���I��Q&i��J��72��wk���ΓȊy�F���JڂW�λ���u��^Pw��������M��c]F�U�\���ވ��a��/�8yA,��gr��+P�����9 �-��$�+(-��'t��T� ��k�o�W,)�[�a���'�0-��Ft�;�,����>�:{�"�o}�!�k!���I�9 H����(�d�`�=)�����X�Λ�u�~�7�=��s�J�a�-�C���
('�݄JuܞV�<Z�_��Sw`Ԯ	�{������#�M��LGM�UXlxVHYEB     400     140i0�X��I��N�(͚_�YR�x'u�g�J��ǾE��s�\� �*H�����
gO��i~�@3�n�/���	��� Ϊ;��+��&r�kƉ#k�����p��bL�bs�J/�6������5��6��y���^᜺�<���m��x���Jdʂ�=Eg3�خ��@)�ZV��O��C*�<|9@C�W��ز��9��F4>0#�\���J��z�
����9]�p%hN��O.��`F; a��x:J�|fPd{��$�Z�&v?H���6x���/ګi&??�o_�`�`�].B�|=^��6XlxVHYEB     400     180���5s����%tS�p��YC�.vX�oG��p��bKp�P�:w�a��$"���?�D��������Jۯ��K���B��o7#��'X>'�7��z�"�o�z�������A�u��;�xte�"NE��^��d����`1"=������k���@������^/�KuS�Y�e2�1X/�=�_pd�⡄�W���Xd�Hxp�@"���^��K�1�F���6w�[�t����y7�hlLռ�WM��~��^{; �mH���ю�#��Ƒp�9�W�3���\�r맹��n��z��5}����hZ�gf
��[݈�@�w�,��K(+[��a*���"���� �Zo�&��]�>��nLu���׎�s��S�gqU�C�XlxVHYEB     400      f0�M`�dU���ћ��k�.G����b��2K|�%��,���hc�h��z�}����[�G�pTK}�,��I��T��x4���a������Ӷ�(��X�XX2:8��CQ�?z��C��eRI�E���%�H�@v{��T�f�7 �/��Y��N5<{y�`N?�4;ax�h>�9i�w���XY�L�l|ѹa0�����a��c��,��EsbI���j��һϴ�4���pXlxVHYEB     400     150_miS�K�w'xS�0j�v\���n�T��}m&�R�����"|vV}�S*����_��F�Ʃ����/Q4�6�Ý��)H_pp�
�!�QM�g��{GnB��4"�-�͈��l��o���ZjZ��x �b.f��t����'�ke�:�b��|Fs������:h�u~ׁ����i�L#Ȥz��^O3N���*��������(�)i��4��|[�a��8��]y8_��ɒS�R�E|DF7�&�QjsWxK����z���(��	ձ<�{����mt�xӯ]�c��8�O;�MiG%���Bay�8�KB����6E9U��0Rw�XlxVHYEB     400     150L���f^�~�!/�ΞN��r=�w�|lr}�Q\R���y�򘐪4�iH�v�+g�?q��)W��g�-2[�e�Y��Ln������Y,����n}�����P�� �Z��[��$ulןBZ@��%��tƘT�qH'�N���@��h�ɻ���)q[Gi��d����t���c����.d����,����HtuQ߁b{.�IE����q�7;��|-8�'���fVg�1I�O�z˛qg�*��]D�*;�QR���mz$�Dp[�u�Zw95�[��H�]���N`h��2�S:|�N˝��7/�[��f,6V^���B�=�WE��-S�XlxVHYEB     400      e0�]$����N���w�ܻ�c�&*(8���^��z��8������I�9�WD�:|�
pu���'����u�����6�j?�"�acY��f��	�\o���o�kن�Õ2_PlB��׻D�v�"��]_ �ެ�5͚,�LTN�1�l�y���ٶ-&$s�w;͇�J�#0Xf�{�D��7e$Z@\Cl.5^���s��~�7���0T��'XlxVHYEB     400     180�wQ	��*�����'�eG�렇����X��ŉy�tR��`^k�/N��b�x��G:	�0�@ 9"먵q�	K\L*�n���iw�N�����RJ���+���U�z(�xc��=XNs�M/c��eA7���M��Z����dƹ�k)D����RZ,�#��I�{��W��-��^���ǳ	���h�Ā�@Uip���]��h��Fxͺu�:���Zq<�����n'r��ǚ�#�K���	�K�;�;��^;,)�O�����q-��i�O�J������oţ��i��+���U�/ǼaEj��=�7Z���%ma���F�+K_ٱ�1���J���;lW��ߥ���=�6!��7T�ثR�cM�._��dv	_fBXlxVHYEB     2f4     100�c��J�-�wI�+B^�ۑ< ��
k\�eM��mC����r4�輈�� t��	`o��n0'�ͽw#����L-�[#dy�~x�o��@�&C�*\�Y��.~3?�KpK*�q·[���Fa�oΔzt�~ͽ���H�k�f���Ă|0�5@K��ԙ�������n�R��y���6�dd3���IC �N�����>�ϴu䴕�_�SqFR8��8� �Q�U~%��B�����:h^�m���eNČhE^�Px�f