`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
IkLjosT3sbPyA6ib6GLk/QVcKer62784zixqtNvliUVxHiHHf8s3w9BuEOnlSR2uNjMicWjhQtlI
Deos9XevD/mnt3878xpg8bPrtaE3DSlisIse3DUm5NoiCFfXnzAnmpDnk7+/IsgF42AJrDNU3Swt
sRgZK560wOquk39dEcks/tuu3CD3R6KKYpWVrcyCV7n+WxNfGnsVDbg6FBKne4jn9FGTSNrSkeG7
Z7khHSzrklgRsZp3JEXMmBaz4ysq/X398SFpELitGzzXH5Jx5z+Rsb7ERqmrU9eVglQq/kRCW0/n
xEPPOyYjOOSDSKLOIRbyhu2zJDXeYcHXLxwXuA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="LHqMUJoWDq8ItP8ysIaLPXYOpqc7vZJmILT42MQBDJM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
0Mu3bES38vYbJDI4FPpjVlY38VBdBV7SrXtAv3qXiapBzhq8rYK7SZsjEEKY0QAw8d/hrwjf0L/d
Qbfys8cvir+FuGs0KnqhKZapkqtq4K2bDn3IeXCnYGN7cscM3O+X/W/OJO/Uco+I0puyxT3GzED9
UHPKDbcizAw5DziT1QQ3ebN7oNjTgLarKVZorLDxWNHFs6Fv217Gf1viINFrY3Skl7+q5vDxbqJS
tUUpCIldsWnCs9yr+OGOUxa3EVAn7wPDYVNnHQS6LkMpd1AOkBCSWkuLNrNAzk6w1U/YrfcHdCIq
P8BRXUXDz3bgGZGh0Xv+XJvYVyDSj6YZZgiyYBepBvkp+DOp48E9L2TX9vb/dtphJpK2mXIRdKRU
Od1+hj3oVFDZZ14zsaI/1V2YENk8lRbPlK2Ic91lkv0Y56E/NwKWhtyLG82eltuf9eJRsx8kUURO
ZFCniR+5wPe4nZ6u36j+B64SRLWBIY26M+VFTtBAu3ybGzfzVgDnAcnMDx2vOiCVbMBqolmJQG9G
6oODH0yIoqsAmOrewQ2vToPjtj2TPgGZBDk8uUzZ3mU10oTQ9xxf2xgbYySA+xlTGrzxKXtb/f8L
u0h0HP6khELVIauLqL99aoIrM36cdqMN98ctGlJ8/Dl1K1NvDnSs8OATDSEGCHn1OwNgJtK+jOkE
fOXxRIM09d9I2yEby0Ieg76pg60s6b592V6Am71XuVy7pwUMH47F0qqYioMvxc/uCknOtlyIvuyP
4RYN0V/F4Vp89ox9n0zf3kfEyTutRazY2sLG2Zc4tBU23K8KjG8GyQjvJtPWYhJjYIyi4Q4VoSxZ
iOi+3xKRQfpO/N47jJ2pfR97NB5wf0R8a7FOaHf+lf0QSYCXI+gTDD56Qgzd2kgzfpsjTgQoRxIM
CHABGrdd+WozE7VT6RbOgspJlVppU9uYpuqoWDLvKx/QvWHEr0L7O5d7SDRSepcBra9eEKZq959Z
FXwyz5EkXOuuzoUO1Lo5H+5XJc8PbE5KBl141RmEzfLb2fpTwEyyzdb5QLUTPnC3OqFePCT692Vb
QhqjkOPmNt5zqlTsCXnTYZOBMVeSBfE8XibcU+XMPawyJaKHN45tTUG9dqH1uQDx27G3XpCrYXFO
sAPiD5doXY9cjrCyjCft2rJ21tqubvHNde3zNVuatlFvM3Gb5PK0i8g/giFKE4CEZtLFIEbnIE+h
uqjz9DrOSOpOCRAWgSLprw==
`protect end_protected
