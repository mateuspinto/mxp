`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption=(activity==simulation) ? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
KKS81l/IzyJt2RtsUzxYvm9WuGzTYfDu+aCCu9CVQQS0xFhk//sdIyNelRFl0VdCLmlzI72kaSXn
lRhLI6cyOtT4kVuuQdB0ei1JMVBSAKdsi7oRusZaM4hScT5zARfoQardWmdEMKgFkzCEL+OwuPzk
acZ+kVQy9twFkB4q7PXKeZqAxxPu22zSrEC9GPaxQfXOa+UOFEWe4EwIVpkCJujo60rxihHvaxt4
b6UdN8iw44Trrf/rFj+zBqCZnDtGkhvZDZ+OWhhMIOBYHf4nRfEITZEIOy+bFs8i9lZ6N5Z8TXZB
aEgiu2jx0iohNpNydRfVYd1OYmUos6hhWStc8w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "false"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`protect end_toolblock="kQcbK65L03LpIGm9MGjSufwI8iesksTA7V4n7yMWVCY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3872)
`protect data_block
DhtcORi6u8j7mvNuaKDkEFpdK9t47gI0x3U9Glh14LfYmqyR7VP5hxwLkwnRJOVuMpKXGZvZUibU
xXoLOKPTUxJcauALHcju6U/0/oDbKUix8JXyfiPsy3eD/lAlp32LoVxJ9X6oOCez075d3+3WXbi7
RafTcK0CPn2yNifPk5vvmyqLbTex1rihv8bxui/KuarHeaA8ZwFB7rBHJmIQei2coRqw0atBqRyG
hU49olXFnvkN2psbOVM35HahwcHL1gRlcMHXEY/zXX92zqMrxoCOaiPsPjTpPpLpS1+H5VooeQSD
7JUOSNrqpbg+HOhukPdmKa/Rio2Ti8OjWJ8EwKVB+YU2mkKyllAQG9IsT8XA/i4ikioczwzSrq+N
3l/tfXLQo6jkKu9geG8xgO0tMuNVvQAZf34a0t3P4YHFlptqyrrCiLxwwx2qbyB5IlEtwGqu7uQq
VV98xTa71k3k58L5007jNGls5atwqGcbiw5N/KdS8/gBw4xVuKG+1k8R1o08qM56gsQXJ3acR50d
RKiw7ZkpekjwoK3+87x6tq3/Z/O3Ysn9iJFFRC4axAMvU6/rlBucBDCtpMHvOLlsb6Z1RDmqIrcX
0+hdRNJUm8i4a3pDubFhG9LUIjUZ2Lu+EhaFz1yhklBKWrrj8r8dB5ZM4xikg50Aky6DKWQaagsW
ldxqCUDpJR74uHNa7M5F7OVHRIokYeuG0mKX1qm55xf3eY8tSVEzIxzQvj0eKaIYCOS4mjDKlJYA
0dhCbfDWQB0ehe1k91PhxfXVOWoSUBlUvz3hBAErF5fMH1I6fObgIWvIfDu2J0vjk0xlW75uI3PB
aoEffNaHGSdkdJ3EurFhT/+EiP9L4ZZgpYxz+e9qdUM1JHIBBPgfswDkmAEwDhdwhZBm/7U8DI9t
HkUgkehwv0JIDNJ2wu6th+IEdLQIPYiKcx/8so/3nv1k+be4/ehgf1xzFkfkE1HbMOFvVy6vcb8n
zvERn8XgPrpliocSESIdp+1uCf5ULu9J1KTReOP7OrDz0graEsj7kv4IfK+egRMzTQ/W86ypAPEu
GYaZSP7WMpmkSCKgEpcihAHokMT3S2Iudj11GeDwbPRO/7cM1teqwpM45quhxBfx0gUFEurLKLgm
sMq6CZsC3BOPrZTJIdGgR51pzVSDCvbRMmpCAPRFdY/hncUE7M0LHDVBuVZgcJc1ELa4zh+5Gr2j
71G9QD2bfUgQMf4cwhpvWF4facb6B0x/FWN4w/vvc2aJhaMj9rylS7X3hJzLWGEYc6+SF2sXkDKp
OCZXhDjcK51PJ9aVi5jYCW32Vsn7oAnPPpwVvt1U7bU8Oy3uzAW+aaYHxoyDnPxVeKo96UAUrtnH
lRshgXvhi6b/Qmcv28SUf7NddJRj6g1KvOlWU05ZlhFw2IVEuB4qCuw+sK3/EZbJbp73z8S9vsQb
J78D2C8aF5YxQgIuR7GUwgBkfY46KIdYoLZZxG1AJ4NgIJD8b4CtCju9IXfVkmSxwLbekjrZ5Opf
u7jWF0yDb2pUtZ05nthAisnzA+6LRdF0abA/E5ShqFn5mz6GRAnGPPllVO8GD2ce2iaun7S8UeqB
v8Cfv0q8oePvk5Hv87u8RxqX0p7HcHO3CdPJBjJX/slhA0B0Yb5/Pp+eDZH6Jy5bkvEpbCJushAg
6F6CrVstVZ5ivY7EeXVGE3sLtKtk0hhicc3q0rBPJr/KZNE+6/EGnY4ayu1DaqtVbS5Hu6EHvTHS
y28VbubpiKdhq0o5Qkqz0kGvtcffNBgDSPshjFhsTTrSSrQE8jvfsLqPX3YhqHdJqja+xOWGs87c
nigyDpwA2nCLBDNx1Y8WPpUeY0U21Nqw3dDpRrjuYrrFojFWfH6KTX3yUgZ+RZertnjmmbqREJwd
LtTEhFjrQwyU4MXErei3CPVDDl9RK0Bi94mO7qBfOiKGnXc95Muwqshx4OW704ro35leg7BYSp68
Hhm/VpTVSXBIpk/JcUkJfekgOzuN5jRFuJHlmTUT8DZ7Z9D9LVbhgKSfnmmccWB4scQstIr6YUIn
vIdOUDrkJF5qAbgir9TaqA8khZz7wM0RCQoLfIrDHztOPGGPH/Nxd037d7Oqv/B4RqmfEiho69Co
4Ww9KpWwrlLtdl4qBLKaK9n099oFXYeqqI2JeFLyQSKFTRa/W83x6I7AAZuB65rh5HDmVl/Fd+qH
tklCMT7g4YWh8ni46ZU8kJr5nzIrXChClH2/XW16LKkM5KS3uwb0g4GxExc3vZAjG0lWkJnLI73h
L2kjO9HMBL1z3+IncqlypDd8m5x3R1CaACRMZrmOVppjoA35T7X0tOVfSkyZQLWn0DBqAmSeD1aT
326gSAxiRBwIUz7gGx87rUDJh5gKJLkWvI5kQbWQLURHxRmmWWp4lqRZ5jh1sGt4uobnjOWGGiZs
xgeRr/n+Pf766kcAK7W3BNXPzMdceYRCWkTlIWmnF5Lt1WMGJTY2UhPE0CV9xaIoZiY/T/XtyX29
FiIvTGue2WvxrJQAseY+ipA5+kZNgOgiffd2+5PMXKn0ndVgocmZw9udvfai5BfuJEc/RsemDkmA
W5q3V4beTnpyVmkpJ1g9xZcsWySMwIBnxX99bnvQBMFb7Hfin7hveS4STPPOEBeNPLLMRzX2zN96
imu8Zkdck9GhvbAXm3HfQ1oRgxRo/iVgoA20JRouos/vHkByuS1du2ZDOqags2H6bJj7t68nIka/
nC0j/sUjPAzEoFWdHf/0fbvixWcILM98jrNzOxkJJgeuYufQLlxu1mqSz3SzPN/Tk30LhA4RVDzh
CA00SKdoivwtbmJYSxQPSiLBdxTkcRQUrrO7S1227gTCK/nO8rrWF18H3yWybFBafv01NrusRI6b
hbNVpclp2cKfl3RSWruuKNsdnnG0rs6ea9sJliWYJczeKYiRqgqzOsg8atZguQoNUI+IiSlSiE/E
VS7xEs6IO5nFZ9WAGqsP2Tss/Ae6eLWVJEkPEzxsy0tDuS4/4cL8DuHOI/jzYLqbYWk+fU420RWO
8U8kWbn5MFmUfEI1yymTohK89l1Ypod1A0mi/YLF88qdCXlspEKyBSJn2M6wjqi3Y0PmgvOg7Cnh
gJGjPRAe7kvyPmbbnz36K0+zyIPOIHn4XsX30D3drjlUI2rzJYulPOoGk/MQRGrNFnU2MvLGDieO
K1X/3PuRPGqpgTf/3nWGK2ru6/D9vqXKQYUgmByruJ+Aq/MYGmqdo1tKPVGZWQonymCtfk3krO+2
lMloabZBrG7+Ki+izJvbTr0U/2SurYj4ri6+53Y8hoHjzfPL3o3YvtOb0LeOQzxENkupfpRJTTB4
aNXoFaaOvXOM2X6LCIWd9Qln1Lg5v3re+5bY5ioQS/invSFqe7Y4nNHysPvvNoav/HebOAYotE0u
+YZhUqYg36oqxDn0DC4+5voaNYGsKTW1r79OBwkn68yYO56Ft8YG7qUJX3qXVCEBVCdC6zqwPeBL
U9eX+gHADZDO3w+mOC3Bdh3W/AfWEaZM+LeLNeUiEltC+ui9ykCTfW/vaoZbdCOjEdW95FSowS4K
jxdhWjRtcnWwSMz+LzPxwL9QaatKhawPVs8xUV1HUyx2WNHDZdIf6x/aF9WYw8dsGIcDEjxhEGx7
zXJVmugs+H8dNi8/L2uw56n9Hwa+cXBq1mgjR3ZjP2qyujReiGQ2TZYmJXtrTDP5HO2JoA3ftbcJ
YzSv6Y36wXSh/4ZOVwrilBgNz2c3wj5OI2CTKdGZFDqwYt3xF7C5RDpYdVyriMwRdC8xKsitdGQv
dt0DhDYMi1KLjQRVdOlhDsHZj/TuUy6zUYCfXRXWdqSlIMR16D20AdRbq2rWLmtqOLFpKUtrlDo5
ZNZOwp/ABnSBpBrL7zTRf3434TVMxio51dpjj0RO/qd5FzJQZgw0Z8Q2pYoepT1EcvXSUVcXQwAs
on6dEECxQHVtd7XA3TvkunNa2fHiOnGpJhfOjPWhemz0Jz9zUJsPucLqtG+ttqdI6YLC1qrfuilH
Z3WSM4n2IpRFR41cpO+Is+JgM+fOnTCG+XgILfR62iXVTL0jQ3osZTjGvhC1Y60Eg96fh1fAjW5s
PZ/z+jyJeMVoL4JO1KaH/CgMg6xvdPSbMYwZt4jNLeEn/On6DZ3OyRIGIV9UHP5dje8vSD7/Ind9
fe8KI1BvJQ4ydj9l5e2Wd1Op+RXNO/5IQUpbB5yNGC3DYh5P5KqEnlh2puffy7CPz3WMXO7DxupE
Ew91nstZ9mv0FP4VDagp4dW58i0UxErIF0grxFT7VBIIJVUgs85MHe3srfxx9ZgdtovkT7mBEoRy
zGmHQE5x6gAsmGwwdqRTUsr6V9om0BhaNlEf4+wpJfQENDgCU2eZW+MnkC4Yu5EoBhmP3Ks0JHh7
oNGYVJ1yRwF8hChCnSahC53iPcqqrC5P4z9nqcwHj9sr8JI2+qQkdQIksD3DJhmQ4fkHnlJosZHk
o8zyUlGMlaXfXgeliXSjj8YytYXpyVWFlHPklPhoCUb2e0dP38XpRfb8NIAJ2a0bPsxD2G+RmqQU
rC+0sLMt03aoraSgxNkuZHPG5vaekZt0sGmGlv3nOFvblygHCt1JecZjb8l3q2XeRlP3t8UAb9G0
jeCrnrw93DEcK39fFwRDvlrTFDCc7b7jgxaW4KHOI3EwWG77fGypzOJa+6MfK2ijdlzgFNgBjtIB
KQrQ9qtwcMZa5SmYZs37Ukxn19YRHVzyBc/dXeKoTovZiIpTRvzdORaI0VQOfw6jFIEbO1vbG0rQ
iSJEoeUNulimeSVXfXHM4owWg6vr6H6zXBfpwIZNTcoBAbY6Xc282FQ4EtBMsB5VqfYng4kP4pLU
gEAkou3sGeoL/YSaSVIQV8KiC7OzI7mqd3V9gdk3iqYzskuhpvbXo8NAtjlnWIEg64phmW/Mb4oh
z9bRvsKwJepEm0j3L9jtQ0PyZZlcoxvMVjc3E3bYSkJoiBlB298igkRdbisCbkF3A0eUYqEsGFZL
7NYH4JQVEOe9JjXObs712IFPe5gFr0SVUtaUyQbxV3schkxT7lDj5vifd7srDmQEj0NK8tX+cEh+
oUaKYhW8Z3WfKgI10K4+YhxFLP5IsZDyIbLFc6ZEva8WX04/Wh5r7pzLnz0Hsj1MiklUxNA=
`protect end_protected
