`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j8TT0L0MZmVcxSF6URU8dlcdkpOtmaBEgNc6JwBLtB9rT/VY/0M1+gqfIXhpArCPvRC9YBHVq7b5
0/4U9BcJ8GGh00OJzyYz+k+ZFqYgssB6zxgelhxYcJnQ9Qrydo1L3nhXcm9r0TDWE8bM0Bb1Eu/X
BMj4JXtXuDCklnRr4yCeQoCCcDSNnji+TD5PLtZBjUmqBRF9AN00++fZJ4UOdBIZwnlgGsmruHHq
/bAlWiKdn8XFsDJlZf7AJmPq3HZ2lCxmHn6dyK9ZqSK8nHhrcECB04DLE6YCRNqoH2aQ/Da3efDr
vqDdFOAMkThqvFVRBeg+WMSqQBgEwkGh/yF41w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
GP2lQyAO9SLLp/YCsuu6jXEih9Rn2WXBALErNL++yEbHTAsDRVGvYS4ZZRbILK7NCoFGIuDwYT3A
fmiIY1e8qF7TD7aIEYAeCsgU79mPdgwfgjgINRgN4XUNEvQyaW/2YKloJmcenzZHTuNOonnzkO9F
fth73C+mtXDd4/e+7eFc+s0iOq3rxk8l7vKNW4/HRatXJkhWVyogm61gz/TkdmDLLbVQ2HDF/8aw
Z7Mh7enCOxiqEUq8AeisPhIQT2cVsWcBIntluYksN/g4rbRZ1otxW6EOXUPLb86v0TLx2SN/l9sb
bbehKGcrql+FspATePk5eJVAW/MwgZYn36Mt7YJF9UdJ2eTBnvm7e3lVe1oh6MJalhqwyG6t947M
lIlUi2oVg/S7WxnaA8149Hiv7Zv2qBG9GQefgfU+BttIKyHGgj67LuelPLZPK9rqZPGUXKOyotqB
lHe5s32Gd61d7QHlNqle1fIrzV2hj+T0WLG4ccMa2R0iapxP41HPJze6tc4iHLxS82FBH6Kz842i
RIC9SLg9iiT24R9Oge8I9+e651Hz4ceifV5v2owQacLfMLSe93GoTXC0p0j58ZbLr76jp2UKwCsj
UgdsiKxqw8TlGS4rKEGBLOzHQWsdSR9L5YVdEt7aZ8QF8+buAahGvEHkieDSKm0otaOB4M0T0/Ms
bD3C3ZiKB9cUIY2InuoFa/nP/YGfJDx9xg1vv/NbCswtHrgkRx2lAWSyd1AbEvkq2DBDfYeHYTtu
4UEanTmYXA8AFSbRNlfStQ0kCfAMqujHtZ0/hyh0RbE9OdkY7dXsHK3hrCizRl6KAvMbklXZswqI
8iTl6Ie4ZvMPbZ0Kb2du/T4CGt867oNL/XedAMthZSD0fdlkcF6lWkIiF67Kl+RIuAFxmVIC0qak
9OjYoYyjYBUIhcn6Oy0x4Q9F0sXD0kTfP/GdAoPUenH8CA6a/dXwevu7ef3lquIpfCMFwncghkR9
ilGUqtque/LOjHxQfNcCRUGF1HU8LU06er2zldj+hhaXlYhVd8SmaEp5jafUBFl6exsLxtZjGWlb
wxSjh1GhCrKHU85Ow8E3eqUka0nA5146fJTUNt2HyXJdYOIzHtMAayEo3pBAkk90CarBzQexJ9Tn
7be8w44F+Akz9BKsJs3T2CReWYCkRWLPc2d3cwzHwau1QikfnwYF26oebbz905MiQmo/cvOqypIA
Cav+6wV+2s45vn/y8eXP3FqthA3LGa/PGKP4RwVctJyiXkQtPhoFduvjqw2+fKd749hEDkawEwwV
bpTlPxpc1JvycUOh1RyiBi9NBue/v4u/5q6Ndvx4jO3NY+EQkHTYIYCXpl+qIuwJMq0LL+2ySGnc
ySRaqHKXTqBJdq/9i4Y+EfWK6dOly1HRBmcdY1EmiMPG2Dlc77aVZ9BONau91HyXfSbJLXUsrOii
tMCbWXEOouVs9KsQSMCn4/JBItGfs4afoZY2XZ9gh+Iz6dD1xk2QnCqZw5c7ripZfuXdwqWW3Rxp
EgJ+40lmUcHTbzCTqlBkaAbItyVbhLuCOD3vUTv+QZXgvUUipKNr1acLMsiH2zLdr2rFeO4b5MeU
yJE64wICmYYlEL30oW4akJT1xbGNlpZOmqZZ2sn37vlp48g+Gi6BBRUjFm9CL3kXH8M0nQ68PiuD
Czuna5ZpEVKUaDNEOCIa+fGEjCAwqwSD3oxO7a04uG5uCp+TV5h8g5c6P1WWwQYLwxMk8HxLwAI4
/hVkMejLdV8Y4fSBPJ3dGjvXH6kHzy3LghZvPVj2S6U58B37OGSWW1xhOj2yr9ckg+M8qqCsI6MJ
913IrDJcxhpAQaIgmGFvw4X3un3PoTLOb/3jcXPbQwvIaFNuzC3GiPpNF5XkiqVBbfNn+kLgCBCi
6tL5HWF8xCojQ404szHuxj4U0MSfuQ1Miqf9NT8WOskvRF/IFb8uWNq3yqfmYEhtR71BOrbtQo2P
QskyqoLSQchIeLZR1vAQB5ngBc6MNU1Ej/iv/qSHV1++wlIrmCPQAdSf1NKoOQCZLDcLdI8kctun
xcf9u36HShYt8nNh7ZOWCglFg9+CCdb6tSJwmrylBS5S4N4kcSJZun0m8InI88dzARQ4eLrmwh1Y
f/EFrs3XJwlFnrNb/lcln/8prL09RohX+dG4wLdWi6pxO7PfbYI21qSa5NcKnTrxm1JVSJ7Qd6mc
Z3wDQrOoLIDuiPyIEYQFzkmGytAj7s/A/IjXg7Hxaxc6XxFFcpTyycBJkEPI05fCCda/eZqw3SBl
Lpe6zpuY4CN1RzFffs0rgvs4coyqW3fZ9tcgqEgUMy6xvGIYNV2OYNnma/o+qDiCE299H3O2yTw8
13MGFVgiJAL9Df5/CAwmWn100DzwKgHlglx9D9Qh2XNKF3StGqw2LjQMbBL2V4NmlVGiv044qSmT
IQWbaVk5WvV9prihHljTTRl7bntXG8+dCv9x8fW/eWJBfPM/8zaF6NJlcjFZ91UkCt0gehdKaZn7
Yly3gSnBa7vkRUono7HwjTUsmwSJijg2KGgk4OV3eKAvbCG93UBMs8t+PwiZEwVDc3f94m2gHDQA
Ho0FLpsB/JSUBmcH00q1EWyRyAHVdT6TDXCQtEFg+9j59EZJFmhQm6DesA9X4w0JNE5itRCNouS8
dehfufWf9eMlXeRbqaFTnw/LB9F9lk70yIkvw2++Tff0LJazF0/e7+aaWGrv7bdSlRBvrlD4MmUZ
MoSh5aWqRL9yda+j1oOAyiB3JLG8kjZS1g/tL0Ee4MOtfrG/kGdZ/4xTxW0nKKFVr5OJ4APFTAkC
ytrk7eaAlkS0HN6RfSa39oL/I4vhhXwba2pQL8wB/C288iHmgjjd3gxULs7qNHtaRzKDZ5EQeUsB
7AOmf0DAoOkoeHMWvTeH0AhbIFi5jvhpK2hwIYuGyeNDa5eQ361TrReAv6ZVgTWSZUZOCmIF7aOr
DbXBahl7AZxbA/SsJlbxKB23S/tz5vdVWbIxR+t/te7UOX53CAfM8XNh4G9BXNY1SXYh2XjRjmfA
DiNyrpC9TR2cjqup0Eq6duB0isRbTwXBjXo2yBZmoennHUJBEl2HtelewJ1WDcCrt2Nmki7+csO9
LHxjF88Q9bQr6c8TVIEPH3Ut35MahfSE2sDHpkaCsJpI3uFdohTawbrGJQtgWgqMXg1OFf0BPNji
poUuWAlxrERioS3RNwSWXP1K6y+8W/jc4UpaSLmRhRGda3p9eAx2U1XwJxIHA/TxRoExPYqaOoPP
AFzy3rSugF5IfIU45viUh03MvyfPYqW6b/MZ6oyqdzwSfGEhkwTwtwQ1ce61jRYmiVcdeHTfVaeU
vN+j3Ui1ZSVA4noemcRUxdCbJL/vutmGPVK8XEpzYJKeuY4I4AWMtyElprhsR7eb5GxJ+NUoV8BG
J1rPAaByHqSOKLdtk+vbCG1BuWnvb6oZOhajJ0tGxTlBw8rIlwRldOFggM/m+RpOIBrA5n5hflOb
tEBaZwdrbPkMMdhntHWXJELFcuNdfOS4vUZDywQQsei3nfoMoznthDsk0PY8nFM5o8zSMdxFO2na
NqBchsLox04zM79TLaE6XJDCJ1CiYr10U9f5zzyrmpRdsyqBn/r/CucJtMPeAfUiUwYR3JzVwZxK
IDlz7yp4ikdcCyRky5Mu9mf3kmucFfA98B0haWtu7meudpHii/YVNHX4QPgUiV12QflP3hffdmjg
vM7jJ4gFaKqZeQ7qDPIvb7mUaiIeAa3Di1a5X8HoCMv/h4VNLKb6D5pT9TDownBtRp06HPktdtOO
vqKnDDXY9sLBX2FyhpXvqjkskoRbyXiN3cxj0IzjvgNMn/IgrM+Ia3wZPcVFOHIqcqA68lq3tOW/
sq1o8CbscDLV6X9fPnecx8En0nXU1ijAvR0UQHRfeHDbXWp4NzHIFzUZ+DM/kdv+qb7yx/s+RUJk
aws5kLgulIvlNFfWAdx2PPZF8a62R4o4676dzhPxsqk3FOtI7hrsGuO2UCfcdMguzP/COeCaipDf
zzcBAnrDDxGn40FLwhLhmspwUJRZ7NsNohK+3vNjGSqcuMTZp7YFRIkxz19UtB5dLiTK+XI9czul
hZmjLNi9DvdonST0cBMc6YNhP5iW+lU91MdOjLrToULK68Ifw0ws4YFt7TFWRRQra0xNSlSwj7qK
SWdbSWg76yGi0Z7i4WialEdF6uKsKZv29V/17zmS3hgtdRrzSDLSaLHHbaWAkKASp1q+PJ4d5jOb
ibUr49nnOU4/E21P06PhnlKDX9k18b/rnsaTXlI3D8Xbk6kCqwmkUFnHRd4R/q/U05RXB792mSwq
d3sE9bV/FRlBXFbQjDtURWvBDjavMa7hajZCwFFSDTbEq42htPuDBvc0YIduc9OFmVbbfgKXVaCo
umWHErLBo8ktGuG4eLu2fu8w3X4EMTSqyfPy312Nq/zXjPWD/U6qp5JSAZrW9VYYBv6zWNZPAps1
Wgo797Ce6Bd5fHNLlz51VuU0YGMZwabWxT5XUi6ef14N5LRYx++HIbt9FvNx8paoW4ELFIqud8Ns
i/yTWjMp2xdtG8E+QQtRN67bWeF6IKOxTnxCG/Nvb61TaSvCV7M60mf7l87uwBGNXkfWkclCe+tW
xme/KcOSbSaVEl5lniWQk2qVZNJqN4ziOOJNpzpmXizRc+lLZ9S6R/gD+a2XochMjxB9n/GKcMT3
aciKFPqzGptNtPco/riSwFwzJ5WitcK6PWY0yq3ua5rjyW/Y6X9qpZ8BbctyPRPYbU48akPBw2qP
WiMU66HUEPAxCyt6K/rdN/eyFDodGA5BErFE3rA/EKM8yMU0oEAJDUt+bncgSu8NCPLiKhZflEwY
+mpS6TAjoihWqHUIeYwY1ESCEQqJkqKTxaKb2SgB1mkrGFPx+4anVFvcx7uRCxtYP66B2z+2rUq7
+W1ch/hHnPBxPn5qRutxbF01hPS7536dNqoWF7q7xvq9f11LRPizTqJzFehh2fQs+0vzS95Rr4Bd
EeGQ9n4wVhBMD4K+sNc41WmmuC37GMzNBTmTQole7TbxoKdXM1aGqY+eZWBCmyOdTsXuwyE9Eyne
lYnuiUYO45KPuLi7lCW1Dh3QwYkmt/0d/0gqCBxLc8UVIcW49nZbR3auhvLZ4ukhMLidjOUhO0sy
k2EweerJK2/3Hi5e+biVsl3k6vWkOET9NQ6Juevs4wSCRBULzQXld8n71GDIwoGBb29Ib53bvx8O
9mOkvQJ37L+WMTBQWBUldLIgEzBf+Lt4zzSMX3T1JYIapBGSLxUzx3IFZRyW4tRkz1taHcw4UKVA
AjZWSG6t/AMuGdN8PUHRHM0GTYBwryTyYVG7iqkkBR8382HO8TKGbSonn/VT/OKcBC3/+OOjpjXe
1a0GymmZxp/61QQg0UGUfudVKA9LW1DQpEW90reZHqhYOXytT4Uf3bis98IRFHQP5rWtpKRcN0/N
xOl3Jg2YNkBgGpyzb9Vg2XyNmUc9OAtHkeuFSV2n+tE5x09YASL3Rp5UTgA2CSrLWkKEuE7Jjtt3
kQ8YOFYa3PZJ7ydpvRFV2yAzxfGCUeJzsZrhRqPpeQu8pxjAEGEjbmNiVVlaRVdDYhLK5uGF2yN6
tTEsQPyO4Jce4dQSmlRLm+A01dhUVoNiDLCpzlqXXps2g4XWKhrMTH0AlQ5Jm5Ux0AVt0WHeo261
pz0yOpqx4bn7V/w5oUREDs2doxo+PZOx4MYilt7KP/dBxR0rQpKmH4isRNH8iUMDAOau5YX9ystx
cCn7kNHvkogq7XE+UWY+rcD8VtIYMDV53QVINq+S+pOY6U1XG35uKuAxexU2rusI5QJ/mdWEhQLs
sRCcz8DlyUIVEvU6Y1QJyvEKmzfHwo9HhnR3MrXI3suWes2ge85xB+Hxo5hFYIdURgI7+IfXAZaw
eqr/ApylEWjgyb3up5cg0w0moff2FfRgDpGd/qb2/DVxMJdhmnzgEiU02jKFcJJR6AwcPi/6aXeZ
VT/nBaBZV4e8dGJx2dt9i37i+DUWcepGeeAtRvSp+BNuweP2GuaVV3ueK++K+20eo4Vz/dWALur3
uXZwc3K/X0oGlTnSaPGzq+FB2aInZeOpdrGJepSCYPRIaIgRh6NgOMgY/Qk9ERto5ssM8hE7cFGB
RcXFUxq6z1V6QW1SSwWB7LhOLOYp8rZLObZA1oaBTvMA8ug8DPYUfxeu/XtvbJoniZEU8mmhWHjV
tmgHIeIW0pafIwkuIYo5WRJ0cbDazhhqc3wRtpx1IrpLBfV97auQ6CxBRAGwHADs2kf85DziBQAP
+Ai4qr6L6RvthgfnUEuCtxpemuf6KDjekQnv3RtWkl8uvfnZZ7X0mSToun+mw9iGxQmvRS958SFL
dJigf5YhCmQPDwhTx1muOrYaSRkNWoRwKYrB9ZUCudq4V7sIFLUkLUs62xe06GhyQiTOjGdYhzsQ
xhVvh/l1hXWOxlw4g6UehgnpGm26NO0Pt559DEsD6dGi6hdN9jaGEd871MBBKasI05JxQEn/NHfo
6K16P8IxCUQPCr/JlBY7ouyuZQRi8zEMVe1I66leFVQKGm3aBzoGL3p/N3vFxW/wS1+L3WYhBnue
iw0+P0T2xZCl8nbRLxNExiUE82OgRDk++g57fyajTOoZ33vBBwdSdz+azMHK9vEqdyn6jBWxh/AA
KIfVroUXK7SgRy344byHZejV3WUZAQ7oafShE8NArEZxFRsdjuqkXAS5VNC8Ljfos/XIU0cY5qYO
0JwsHWjehH/p7allFozkFjnsnf028luuA+WZ9qvZP2narTLEUKFiOZhcn/K2StQe3eOzi3TZoiIX
tzzZd7RIdpjtFdAnbVKfbjSQGe/pg5ZQML8YSwt4e9eLihmw70rtvtHPPke+BZQ7ztqh+8tUqTS8
zGRvY+8ybxV/iJl1PynqW202E9LSCUfOZPnw47QOPT/XDhm1NGTjRSSbMCL6Y79QmZ0t0Rv44do6
QLcN5ocY1qoZ5OTV09Bh47A+mpPbECNayWvbfcSdmU0ov82MMyk87+GpyrAvjyQQotl/OunYHe0t
8LSqFNgHoV43qYiJxjYh/1DpkdSCcsFbortqCgU0eLaT2a01BqTTQRAfvWr4fIJUSFGHiwtDyL85
NBTDmPdgMJEhsH+YTd5CXRg59N/3GQwzaHTNVLhIo9i/DbCfwTPemz1yHBd52D35bNwrSvONHlg8
VtFMitV85nX2iqvUddCSzOiDBtZwIDCKr5CJ7eKeS6NsDNa9QEEWSbyW9BU+ZgAo1AtU6Bj2f6yB
9iF0iBtgoqxm/5fdSagRrwQjXZgbPDZubwBOlbrQ3adypi1rVUaZ6sOImRu3xc2xeOU5Koqsvn18
IufCQyFXTQeek+vyTWg1F8r8QUh+3Za51pYNujTeldI8yV8POa5iWJYuO2J2AQPGvSuYM6/jaMij
PN583Bz78SZOltXi8rQnKNg0npg5f2cqAV87MuJfAXHa48Pip5GMXA0DVEVUnCH81WQQtFJC0ZZb
slT6lL59lbiu7Eba4m6IFhPrnF0MK1DUwZKtB2ttJPmf//+plwEk2YYd1hldqQBm6gi+Iqme8Dm3
yVlXKBlKVmoDPvs3l0GaP2duc7jtf42iHvHz8ilAuRGb263TmDcRMZdTapm0ostfz3IjWef3Z1dg
2YnK7+oAagZdCmBByzmHH/q3Jhax79crXl0TFUuP8sjNWP8aHUZipv7Y3UyLJ9WSYDsLjEByfr5s
hmnsCQ6wMc+b7bhkVw3zolcOUOVbNAh5HHujVNDsr8XCZdAyUz8UwxNd7LtEfsrCxeCgh2LWCZBz
TYbQLWzRKZUEArhl8IUWoVjnp7Xz8KMYqgB2gGIfx5G28QaEsrHX0xvbafQQkz5S3QGBnHxeCR3v
RlND2+g+urQ44iizIHCJYm/3YpRSJN0YmC8D4eevn+/bkv7MSsKZ9ZoUT9a7kkjP+7jyfzK7+gRF
Oo4/np6INRpo2++PzPWorG+iH5390G0fIlll57euth/QQNYOBgRzfCMESCCbYL1AC89QJaAkFfLa
dxdGeMXgBGjMWyXMPAPN/+FMvyXUpNadtmlq1VhfdaJ0PPFLMWc3qtRd1Xg1zRf1aO9Ww2r6A5st
5Iv7i7gFZZ952Vu+y6caV5xiABK4QQLrYAEjotTNgX+W4dGpHBIJV1sYYxuwhfm6qTbN24RO5fAd
H6+Sx1I9LOqniGaYnIFgpsNE9mezcwATgi22+9J7V06xZH1nb8iRSn/TMDVGFV6BpVXb65Yhjsnm
J2uCD9qHdKC2rZRry4R/ZGXk0o9Jn9ER5QGaPBdMVf8jN/M06/Rx4tHJWIL47wtoX0gt+TNZwXPy
xxndLp9IU93E3bm61r1Yaq7ZrzhKMnB1amBnkudOcOoY025J+mVRk9pEtCA3wwcs1QnZQpoDNOur
rHGVYe3yxuwnJ/gj5Js0I77ejc3U3uIdTNN21hPMhZB+gcPf0ZDUrEzI36cReN4noaPmoI3jUtLt
aqoupFOn8XWALYsAT701Rg==
`protect end_protected
