��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ЎW�����S�s���z��R���at����ΰ �y��Y��yR4�;�x��݂���d6g���@��fY�	Y,&�I~4�UN"M��@$7���e��?���MQw���+�^%w^3���q�Gͻ1�Y�0!�#6�a��V6�:w�j�F������A3:	�B�W��ݑ�{"��X��}��&���g�oL �H�H��,V��y�/&2B~��|/��tۋG�?���?�nU���˄F���޵�e�E:��#5~���س�_Ew�]�ПR�R��&�\ݧ�e�E���`�!�tOE�o�I<�HI3�gI�O�nԋ�}e�I1�@'D�,�#,N�ȝG}�FoL����0��[W,^95��"dZ'_������+�M�Vm��F�h���$ۢ0���c�;0g�C�UT�+�sM�A�:A�ۦc,7��D9�[�(��@��0M<�C$�t4���W�T>�d������dQ�IG�
�4��;��.d\�� �3zF��>t�%D���fͭ�5!�,;Ml�������D�=���d����9���9�q�&�7�Ղ������ �we?N�C������;��=IEZ ���4���N��Ϳ�R��\�q�h�?f[���s�a��(�n��N\2H��숾�՚��ct#& ���xudsO�|GM*A��*>�X->��R��>7~9����1�6l�����Zp��"N�y��*G�jC(�P��#"���׊�N���|w�E8����d�ۂs��L��),"�t%BR�16տR�l)i���:���@�D�|�|�R%���(�"oh�L$R<m9{�0����Q��A_�Y�E�Y#��k��F�&��>�;Հ!��~hWn�N�5�DR^�b����k�z���Ťe�y�~�����TFΗ�����vukB�f��XB�����Ӂ3�����������gF��%Wd3�H�~�h�:P�;��4�ɣ�%��և��kE��.���`����?s��m�T�,W�8��J�Q�nm�J���S�����s2���^5�ӕ;�P�ֵ7 ���;vFx�[u$��7;�hTd���#m�6|�L�9�������]!䔇���bq����u0��?�u� V�
tY��'�?�Ul�^N���}��z�P8��}�4���?(MV�ܪ�(�4���#P�fъ����L�t�J^�f���H�����!3�yi��X���V��v4�dN����=���PNR�o�����U�qC�G6�
�<F�1ʡO/atp�׭oJ*z��r�x�TPJe�r*<�u?��D��A� ���Y_�<�o�z�xSH���;]<�->����sB���̎0�F����*t�a/��z�6�Ne|�%Mw��^��{���)}ʭӨ�_CID����w�w"��t5p�1X�>�ʷǰ\�\�L��=�ʖ�]�6�*�O�%x�Z�,��1̿Pv�#���U���J�
/:���#jx��njD��E��
����3VϦ�.m蚖��-�k�a�s��N�o�eEW0�O��E]B�ǴE�"��mu����`��p����i�\�Z��?֔ō��	����fK^PQ�d�����Z8'C��i�������03�l��O�C�<6�8r���W��~���v#%넧 7I�c|�s�� *���~�y 	��\n�	V��u8��M��ר��b�~���@���{a"�vQ
�jPx��<���N�r
+��G6��J�ܭ��X��q%�5�NϹQ9"�y+�m���QpF{�3P��y�0N��{\�G~1E.Z���@%�*���3�^�p���w��F�9��3�g�{*C�,U��9z�p#�.���(*�⎽�8�l;�"�-ΰ�OBR�;���.�Y+hj�}Nz��)��fe?[D_��e����~q����ϭ2��ϟs�^A�s�1��M������zV�4��L���q&y���QF��X��]��\S�ֶ�}�r��Mݑ�ۮs�u�V����E��tp�s}N�E�7V&������>�ŭ�ff��N;�)��|4v�O���Bڗ�Rw+e��#���6/ɧ���d�6��k#�:��V�HL���ȧ���
=6C�qC>��y��R��S������������T�aDI��~����Y�t�y���Jj�p�@h{bC�C��ys�Ї��*�9}�
\I3��z�H�@�b�eAZ��p�y�)*��-��߭��<~��z�_���K�x�v���;]m~U|��$��iG%6f�/Ypa1��̌�X+i�ǌ�Lt�ot2j��K��K3��2:
є�e\Z� ^���:'�E}��[G}�{hR$���?%��,�Q
��C�6R���KX�ڼI/�4��!��Y�R�'?EpP�֩���R�)<�M�A�\o���cJsG��u�+WXOD/w�'��p{�ґ��2,�~�|����}F�#�v2�m?[�`����:����
[v���ִoB|�`��^�q���4�ǻ�߀b��O��t"�9�ri��9}ݮvHhZ�K��`OD2d�T�4厮�(%Fh����aB���N����w�\�˔eDՃ�HJ�����MyL�$�5����mm�gT���S�f��xX 6*(�͛=���i��d�z���a�9:y��l\¦�0�n��z��p �N�u*��-�o���4��z-F��]�[��Zd��%H��^��Ia�c�N�C51�4K��J��>�ݣyB�: jڙ����/3��d���[v���珒3�+�E5�� ��?�<^�T��#�?m�+��q(�;�ݹ�K���^�m&�P�	�7\�ꂶ0�:9�|�3Jͨm]���C��ݑ����O���<,��X�_���'�٥��B­%��Ŷ������A�g��׶Vr$l���e}����3��!Ͱv���x�yC�O����;O����E��aʎ�""BZV���{���]r����������DOүw��g6g3���/�,�Ձ:%�7
����2#W�}h�؄dP�	!ۿ#��M�NLd9���}RZ��7���Wƕ�#�`WA�a�>�'�'�t�]E����~��us���%��I�i�QJֻ�8�vz��k#�93��d�E6L0�)��U�4�GU>q���Er�Bn�ynaxW��K'UĿ~�!|��6���2�cL�1%��w�YN�����I|�+��.��
��һ9Ύp��Ƃo��ǣ1u'J��5�Q����kMr����)d�r琟ϒo����-U7B	�m��h��]�L�$=��"$����9G�-�O4.�JpXP�?�C,�s'L�����#�7�g���1�ܞ6�y��p�乻�d�*��ɡJX�ol'��Jĺ)�:X�Bm"툯k��w����v�����?:B���"�� *���*�&b���X� �v2�=�Ŀ���گ��I0�*Q��a���#:�@]���/׳�J?�����]B��V�)���0ÓW8���`d���d�=��w
ȿ�I~��?ߞϠ�W�.��qLV��"	L�V3�SP�z<�&�s�c`82�dj0څ������L�I�V���f��-[;���Ш���,��Ö�ԉJ���;K�T�g��.��0�Ɠ�[��vtч�E׷�u&�0sY8{�ܵtx�,��SD�\n��Σ����GN�L�S.�w�"��|ƈ��G^�8'r�S����d<�%>���� ��"Ά�K�$UT�Etܯ(�n"M�~��:�j0 \�.�7�: �]����<U0 /c��춟dȠMVE���n��/GdKJ;�O�T�������[ui�� z����.'��Q%o,�� qyK���*��D�T�xbp6v��݉��0<ǜ�u�R��kͻa�~�{�E���y�_rE�^��ZN..r�u��M���/toC�݉6Eg�O;箎kh�KZ�p��P�5Q0ހ�b�y(Ez5~�X��Oy��z.��1���U)�2|ͱL��X�\=����?>���^�����uV����)/ ���lx{��S�l��x+z+,�4X@���W��[bkew/���	{m}|�OI�q�f��կ�1����>\ ��D��|�j���!��[�[-���$�w�fI{�},"��㰒���l�n��2���|���$ϵ�g's��b��IS���8v�+�B�L�;]ż�P��p�Yl�j��|���6�5�w�1��)A}RV���������e�*=' ��A�Ծ�8����fE5xK�s���]>�Q|[�V���@h��f}���)��_�����-W(i�BX�=d�J8l�"���I�))�Hd�\��1'p����o]y��j�/�W�[N[z�5Ř1<MV���$OH�&������ʗ"Г��X+-�-�������,n�L����u�a	���6���=Y��A�S��(A��&n�1�>n܊. ��f%�S��ƎF���A�RQH�����I���Qĺ��k����2"]��k@Z�^>Dc v�L�ї�������7l���Al���̯�������^4%�p+���6	�Sz�iى�)8ʯA<#\tb���gRށY^�]OpGK����GZ}Ȣ^�F>k�75��l������f�Р���q�2�h\���T���C*rbV��\C{ӷ�V��RY�i׻_���,y:
c�^]V����
Q�K��Ő0$�sN�Q��J(W�����F:8�bȒ��+���sA�Lր;�sC�F��%SCyN<�f�|"q�e�;Obq��aNc�#��¨;�O��#��x��"���S��B�u�Ou�Ylm ���5R��I��D�|�]��F���@�ФUw0j㝶+��S�SA���(?}���Gp��\���uNP��+$5���>m'"[�Bq}I���K|bf&�54GX֓Y�j��5zrrks����ss��3Q.0,l���
��ݏZD��� ��G~yA-,���ѓ]��4���_�W�"֋s��h3={t�M.i_U1�#�]�����?�@��_!�A%ӂ@ۈ��yhj�ʹ{$[�N��Aq�#_��7��ʆ^�w���G2�nj�?h�2�f��J�̅��(7s�k97 z-	}:��V�d� ;�E�c��b�XYB�Y�Q#��Lhq&M�B}�5���jF�h��x�>���@� bxN�`�G��!�d!
y\i9�v�+3��ɸ����C 3:�r;���i��M�W�aR2wNI��
��>T�q�Z%9�J_��$nv���x�3h�=X�֜4�@w#�oFO��Jيu>���"}+G�޼�UsE��Wȷ�"�r�u �o�Dgm?����W^�dK��
�x��j�h��?XFb_��i�X�B�ƈ][ܔK}������U��CI�=��.��m���{&Pj� ����&��М����6i���q����ō�+)��4�ѐ�B=�K{�+>[x�)g�����Y2[�WSmX��#����|���7� !��C��<*(����F���.�Cm�9Si>���-�����6��d�����]��TUH*A�g��_����*n������̠����}��.s"���G�#UEĦ	[�Z��u��1>��rY��k��5�>���Q4@h��&�#�c� 2,iLC�͇º�8JL�5���$C�s���������e�@�y�H"o��u��~	�5� q���b?���y�]�lDR�f�٣RO-��j���ש���^��ֳ�`v�k��8��Yϲӯ�8��k��9D-��d��F~\�X	eT�jVX/��P�]T円9$��<������c���o��'��d�#{��>Q�_����\F$���|��n��;��w�X\Q`�2v}sYY��ؼ�)� [tQ�ENz[�UvE|�g���ǒ���6���4v�{N^�oر09-���l�������n_]C���	>3#"+���@Qz6��j}~{�l����f&��[-����i���A]�
`z��*�������h#��˶X��3�+ou#���!��N}+��^n�8��Ǚ648��t�ʁ�ST�p�~�'�F�=�c*�X�p ��"6��|
�p�
>�3Fz�l�������%�Sn�"��Χ�ܳ�묬���랲*���3��OE�ڳ�P��b�9����{x�~�b¬;0���qm��(��1�@i�;0�Q��>������y�GS�c˵��U����eg��/�:kD��Z)�F�?Ӹ��k��F{0�_c�G�� �G��J�W!���t}f�o�(p�)� �m�i��di)ڀ�������PA��A�r�]�{�}�66ŋ;���E�n���7����en}|'�p+��_�z���\�#W�D�L�ް�l�Ry��U��%�J��u��[//�]�CX� I#8�Z�N
� j�j�5�(V�OOt0k�~�e9�J�W���=�OqDk�:�+h���ځ��]�3�RH�����