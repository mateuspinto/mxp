`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q4PW3ONO8bbxtVPSvagXLNZPLIRpYo/6C3Ue0lVGKTHEP/dSuBVftXOZr/rsw/wxkpKWxOupXsx5
//x0p8sdLrvxT9sNXIdlyYEvie4UCOfnUCmb6KEjZjoYyKeDJLhXb+dJQ4e7yRtARRo+2QNXVigY
2cV8HhbyTRW+ybOLgBFmhBNLLPixOxYXAEn76R18szMhXWYTbSmgzHzF28kNwUUBVaJOvnSFHEu9
euVklcaR4P/saYdW8qV7p7snNuANKIQb2ek+HM/bktmFoSR++akMGamJgM1/PcPYFlDjxIToXuG+
KhmrGxDT8OrOkMBl1cliIm5f8ba1pBSJAl8xRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
s322cH+jhxrHSuyqg6Y+WvRA+p/A9IJyWX0cHfdfkhuhuRoe+KlkARhrq321qNkEKrsgNi3LT8OH
tHV25IyGAfUk7vfF2elsb2JkfHCoYh2meqWSvYXaeRT9ZTTrl4nFDXNFUYNmDqMkkuUPOZFylgTu
gS/dsFYUmtOse0T/iX7x6PJRZiCs12+pqONCBlLYh5kLQGoOuM5cvsGdVsnCMXkqS90DfWjL9miU
d0NBeOuHfibC0M0JOFLDw7sGbiK7ZhOvKJosTI3qxPP1VSuXv4Fn9vcAWWX4MqtR0IYvs6kigfSO
UCr87wdt/2d+W3Ga2uNNxJKUEw1BcXCZAFcqgRqPGfsZvSeNSF4p7ntJCxzpCcDtn+QrkauxIpLg
MQP5DIRhQeIlz4BnkoJEuFezqQKp6gLOP92Z9Ejji+xlWO9pHGfnl3V9TT7k368hsyy2zwktqxng
A1xICLzMAJpBNQH0dU+dmyL+zStLcu56OMIGlx81tTSCp+tRe/6kUNJ84MWj9vHb1L/mj5lfd/Ac
qXqhcexpxrdU0tbaHLkuGGCiIV8yFY0CArJx7lrNymAhgmopbepZ7an6KzEQ8jydgU7NaP+LAsXh
ZH4dOeM+CRp395DWsJIhmZGERWyXcMh5veBMICRl4JP6g7LIVBWxJF7iOHl0Nu6Njpnc8npQUkn8
5/ySutnfEvmP1yKeNW1nmEWwpaegXQ8DNZysF22M5cGzBO9dF1RUKQIPoWDWXswGP7Lka459MxN7
IlB2i/YsoRTrJk4UY7n1cPeXKsNQcuOC/xTQwEHgTC5gIt4YYNMyCTsKYd6zNni4FOkqXZHbMYlQ
C3t5nJcqYe8oZCRJ9dDtt5SrQfZpKcps9k2rH1G+lmzRJ34EwZajcaDSrm833pL+o4YJF6HXyENE
Diysmc0Ab2l3xFlfo2gfz6ZEtkAsA1ueRtJmdzPQ3L1oAh4SrlVoP8erVZ8fm8FkIW7DC+0XKnrq
AlCJAp1ktK9qxd8E0kO8r/lza53YCilyGnO6/BqAgHDB4q4Fwa7Ivup5wQ9uJt5aRYAQHswZtT/D
M0UwExUD865rnZ14Cs1dF1NHuSziXhpQjIjvSF674ONfe5tAxgrfRABXU+IAwdJMQLhEm02Ni2qk
rvscWt9A99LDXZh50JxmfP1UmTBAg5HZPehDpFo/DP9bxvLJODXqn8j62C4ZhOiaf7utbeaZes9O
/O1UJMra9QWIO7FYXDhr/zfysm14g5FGwr7C+DClrgC4k6FS+YBqKKjLTteO8vcBkcr9osS6Pntr
u9kUBUuSZlGvLOuZjWTUqFofaq33k+smerzT3klro4DDmS4sCW7g4XE10rrPZjgsgBOFSv9OiSPL
qGY8HQHvWRPC4ZEEnyycOatZaXmIylzzcZZKwISqbkLc+IBaxX3I2vv0EmVEA5OfdjLS44EhS4a7
NapxIQja5rOCpO4oUV+W4ERWQCM3MCYcPTvkuqHjCALc3rswMC4rxm/MmayxEJWFaqd+F9A/Qf0y
tg/MybqX8wJxcjcUwjwN0/bjfMU/wkZ9Bn3+y1KG55/Zbh9/yggAClCGtsTRSaGtmets00SGcRA2
8JGxdzb+kSLaTONHTRlFAxNlrAh5SW/tO8g+6Gew67NDWI48+XhDmYf41SWXCXHcumYmcGA8VhFq
amb4/4mzdt21MXBuFsSkEC8LHyOYBgGxczsg3LvfTOsOKaobwTTSoZccaba22YIh0d0ztUTN9csp
+H9vMZG9zp3CaCALe6gaef+FbXKAOKWJtX1KoVWZ2PbdWPZsST/M0swe4hdddMYFwaOzQpwbP9/+
LASPX+ivArzIIioucPnXFUzcgRT+YEGqUZlWhOqMzlu4FR7++Bq/RfxipucSpB0BVBgVp66Xfrb1
laDgAuIGJeptazAHj1U4EYp1ZKWlPivs+GYmuQZobLIKUUKEEVRirsIMLuTklPZdCGgeJIOIZdE1
6Ps5FTwpAN0BqUM/eIYXy9/KMeX/FY3t9BslC9DOyn/8+Pl2x9XH5O8Ij1W6CVClm8JDKwMgshW5
/JQEPvFcy3PpKnRMEFYKOZroigMeFn0a4EHznnhkWAiIN5WBDd6DnMgiomfWMPU2lkomW3pTsMHQ
LUbXl/3dHHgXig6Q+cacNXuiv3VePONEvlKzmdofKsyTEV3/KxtFqYZ5IY/MJN6a0ZS2cAnNca1H
k6lj1MX5j0LLIgrxopISIugCZbuzrNPAZWn1WKXUhV86+hcP1OAWvZpNE951goAr0pMlgovH1TLs
DrGkhsrdR9ym+qIRZ4CeBaI4j09JKyflWJ96upN3u4WGJpOtBYjDAs+DvNylGF/FKnxwNNpf7kdq
Bb7uUp2Oz30zkdzGmCMD1nlasMryz5BDLfz4JtxY5wwCH/09oBR69YdiRT6eXciiugvL595jwwNy
v6PIsmn3IKY1Pry3GOrolKRUCkmlspeVdX6gz5LJZdRs2G36uP55Ygx9g5XOKjDxtsyN5WOal8IO
Pqrz/GkJFDd+/uu8qeheaQJGrelo58st79rvxMPiq4snTKIdcuCEVlGHxVqNbOLcF447Sl5+xqMl
C+HHuH2FKqc+OQWAKibbh0iLwGYcJD5F3U9MfOQeeXv1lqNIVtgkMJ/UaDonwYWUvHM9B0k0F6LL
vnNth4Fv/nqibJEveV4uOAkZOcDWaBQH2Cvz/ASaUuGYbafytIi2mqEOvSaR/qNHTRUcbd9Duy+h
YVapBVDnoS9tqGpvRg2tRCJrTEy2DKOWO/yNPtkex8GnmE27MVfA+t9rsZzCzLRk/u2oXbRaONxB
0jzOquIBQ3qKYfJwqXJVjZfDrmRTuI1ZrIko/QPVF+TSg5WvXu/WSI4cthk5CmpGJSG0MbFCzQ8L
BSsKUQdMLDoQnw8lV38M+2V53ejxinlkr0dm+dUH7FZ0LZu5ArurGMRBnGldABgm5PEJ2F9Y2gJC
L3p/mOCg9D5N2e01sb0BqAMBdXV72acfNSKaf5M84qmTdH/e15NwtUGQdi6+qB4PdhHt74UIi0Oy
PkNS9hm2jqkzlR014BtjifRW79Vy1aCtvJsowQ2Ky7FWdu9C5zXKSxVCqGq0BN7qyDj0i4sSZl/s
gLjlKWDuDh316XCH6OVN5l9wDiT/8aD4DZocgDPzzP4Kf8cZJvWmhGzdb2vieTBjITJthy177rJL
rJhowaP7WBuekkxgm73RaYMD05gPTkVTR6xP40m8wP9NbMh8hfRbWGrMt4XhPTsSTR9qNd+J6ZE9
y8xp3JR6uI73KWMLKyfap/vfg+NqBDBGAbQwaoXPz7NoLkKE4XOx153JRo6UB2dZwEK0MTUZJNqo
f/v94O0V4S1OzKK2M1Do3IiGBLfQ0OW1L6/SaWm3Hua5qFVOAw4RKjXlU7hweoGX4SsQ3LqUzK3U
MeFM712n1QVrvxkZORH7/6fZme5Ox6b2tUDRzeE8MAbzh/p8uVrS6eP7otYGPUqe3S4MwynX4axf
TX7xCL4xd8jGniBqBKTfjFf+whwNpoDlrI6CMNgC+21tHC7lW4q0m8kWyQH1PPQX1IqRnKxvQY5q
MY93wL9hmsDI3iIyLOfpp/LQzuyAUYpX9si7TCZt36LkM/8MOE5sHhTbyhMNmTv8Gmx4rVADLHc5
iBZGW68qC/8u6Btm1t7//SUrNx60kQCsINY6tKDNLuVrhuVNV1PaXQdBtBtFUxlATTih89LTCp2O
aNONEuz3TXqYfNeItjq3mPWhlXcZvRQVIflcI9Win9SxnMUOGNvm01xcjV2g4bZD3qhbEsOFT5v0
ZtSXRWwSwRewAMAKwoeq942WqiwrgiNwVtRgVBwvBwBEWpV+Y2y2guzzrNp96G3DA72oHOjoZ4SL
GbpqkMlTPL1l+mQBPOs5juqSEugwb14+dZi9d3BQh1z+oj1zNPBVll9jrTYNdR3PUNneKx16c+V3
UxLcZqnK2aISuKJ1D7OTIPGbF/faLW08Hy4o0u34r68TiwDjuJufeAZNMdGUTGLIimjqW6Y/e477
2RhsOJaOmAJ+I7WSDiVssDgmtxZKw6aOiUcP5LA+7V10P78n9uljAhhAd8Ow31wp+OAMvYFmLyX8
XWawVQroY8aAdU+9eeYy1A9NGlQSgCr2aw33nebgSq788xSFWYYbcj/1l9Ed2fOMlnfcXBanNXaU
iRUyINlO1O0PZG8PkE503VP+87qcirNfRsgTRVrBpb/iDE2QBU+q+couC/bkn9/QtBnvK0HONp9H
skqEyV/xBquLd/6Pot+Wrjgc+Gas6Bk1yuEKcuPciUnlUFQKTm9IKgqqXbq/XopQX++iKgjRLsEG
gzdjQ3w4pIoHHjAtp8ow+bDByuA1lww1OVUAJFB12RdJ1pJctnmz7NsfgDBMWijY4C/J0iX4enqI
w8I22akJkDKqxlDHQryWh9habKKshaEPCK5tl1LWVme6JDrYvQIqQrVsZ3R+wCgxkuvMkCNZaSCY
agrONSKNwfDY/a/FOiOGTbk3ZIeZz1hoJZoCj2YkTC762b97QfhASYSJyx7R18F0PsTdDnszF7Wa
bkCwoR0DedNlSarMzoPtBC0yV1HcXx8YAA5nbZwH6ma6ieGGQxQCwM+9rLhZVk7CX0hdbjUCbBB/
axG6RbDaLt+5Hj0w12SLbyiArhNLA5WvtOcCSq1T3lrukoJldYRM4FS+4J61UYW9Yvv/NIJWWD+V
zkJD0JADdAVcSem9W2Cp8UmkIhkagNZaIGY2NYkoTEcMLenOiBm/4EuwMCmQk21nlClCtIapC7d9
IWdtlLaFvVxWVTvueKMdtCe8FDSU9jzLygoy03g4YumLZ/bnOSUI2Ml7jOeX+vj00rnTELh/LCIy
JiG+RZsf/a/pwfXUL8EJQNrNleYAnm5AfCgjDlvh5yqJLqjU84cUbmyE87ce/rOg74cSh/L0Fccn
Tw32v93bbrS/l5+YRMeKVM38ukVa9IWleNLdxT9c3uaZDnXF7TaUZ0cniwaUJWQwLhfFQ7LrBWGM
jxcVfDzFTjJcsVAoBxAllp4JcF5dVim2R/wNA0u/NLBo1bGM2BOFhsCAa1ERn5UpbccsESvK4Vd+
AgWpn30nWKy5Ohowj6fBdjlIw9f/UJsjWpgY2xW3bdZt4dhZ4RduT4DW9EACydaJqWACBL0hlOsz
/OYPoTKF39b2Z4uiQDd0uTiC//PWq48zJEUGkQALEWQ43kX5bNmzrwjuZkvjC/wSWLti5A8JvIni
lv23c/KRGuvtBLr7WVUrSsDPJff2kkcOXC2HJIqHoqkBlLJNYldr81C7/EnLzSzR7i0McajxFpXr
7mIE8hk47BjhFGesIkTNhe9yQQSNtbvZIjm3b2Zyz0n2//6nmFA+aazAbZHzSNGOVQm1+sczndyi
S0jn9LaUb1jb4MhZF+dZ+4P3oMdKVbHzTspa8/wfP4iMQxUP2nmmA5xQ/9SHaMibJIf0lAGkv7Is
iqALA+zuW9CJe5cNS3518gTsXW5YJRdVuH5SnLHVavSetNLVSc/SXmq7aqHYrj0y7/c05emWM92N
EV0m/cBqAqNBKBaP9gAxtqzHdHSHDWdbj99W+sPJFjYHOf43RIxmiCMHDfWsLwJy15AbYLPQHplj
Nfgi++HICGROcY0pzDnz/115Tv94TXIoUrHE1okhxbcrSCQ3O32t+eVJVqIuHYlEHlelVFpBnj7I
SO9pulP0HJc8AFcYFAijiqE8sNOustoflFvcrVPqg6i+wyoeLmLY4jdSQ8FGVspjlNK6FOSVAbh0
kSh9a7l6ge5UeS7GqPV4cd20oqiHHEYW7o7waUDR1EMQprQqfkUz60tVsPrWDFrkfHc1F4r1Nzxt
y5VwafRb5fwBCOSzUF3KY+OLj7Dj4AO7QO9DJeqpF2xb2GaLFXiBygtL/bza+yIK7K++cMrtVHQl
gRyqsCjoKdVh9XPRqKQcJFB539MpX6jrV6V4lMkH8iGTPyliJrvtIj+/6LFe1e/Ui2MVG1mZxp+7
YYzIR4FjXumHi5EY/CrsQztmpMhD0ogpkUa5din4Mh3WLgGUhULZaUKJLd6PyDhC5ADnBSWFFek1
6i2OfboOCTEtQtz4O44pKdK7brs7P/EH7bL7tbp7NH2sHx903+J1crpNB+Tk6nieO74Y3Ull7YRQ
TH3nxOPWaGt2BMyNGRFw5Rq/AWIDxr4o+axDlGBUl4f3Kv8rqF2Z+UHVhfANw7cJuAUtqE/ZGKdk
qxQPN8EZZOKFtCATvA3BGGcQzA9meyZw/WeECi8wawNtvYSzquudZ+nhsly+mqOe890iJT5lEg4O
ICr1385JkNYFrruHvJN4wmscixFRVgDMiqG+lKNOk2NU/1J4Oa/Uk7sDxPSvdsDe4N5xZ4zZGBaG
+NIbFFHdENIRhvMiRpQGQskTvEVBicg14JpPnLD1YzHFOUQYnze1HuurpbmPe9P4gashisKoHQ11
aWNIrc27rqMMfg4X2MHwHuX1xymeEFZMz17y3orMc9ULovS2keEwLqPkRM2BtYoFHEuJWdei74P3
xqvU5BCahWwdm0nsId65Huu2S5jOiWR5kjgbCpmfsWoJ8UCuyJ9vsUfnjrAntRT/qCJvQx4FLjYK
Or/d91e2ds8VBfbB3MiFoEgBZd7yRIpvHuLtUlQfdGEQykISJycEk+GxG9xi9zyJRY1SgJtIUM/w
cntGpzq6MaK/Zk6SNXWvHJt1xCbtMQ7ZdCuHqDHXCZhojkqqIPan3gxd5l7RVHp7rpIlUzjHWmke
9mGkz+hZTsHyjL7A5VQQR5HOkLa5sFmg9zt8ymYfPJIWfftyzfYs0IDZ5i+pnkUPFBzjK7j5wN17
DnhU14jENj4tlBJlcjHW3HOFH/QEIAJo2M1RX26rfEDiatXjfqjxG6ab5vWjuOGpe+NBl3zswkdn
SYvR93u1QGUePkTXtPxOpxkBbD9QvfXmnyA0c0dNkGkN2mMoOrsSq6AhWzT2X9o7wD1u7DYcPOVk
prpO5knlv4IyimltAquIO0YXOSLJtplN2Xd2vCXY6LsqGs73HHIdSFLOa4iRyN6FrdQ4sLAXkCwt
M9kWMEzEXD7sFdNAprUarzgrRQ66XZq0OMnarOO45kiw1nvM1b3lov4Qj0Csm5x8XQhLbDvpxczs
IFyMYdUoprl1nXjtxbgtSbV8vNCQm6DdVyEqs8eLqx9J55MZShYJIO1TRXXJZ//XcuCMnvyY0+1L
HaedjkGs+W4dVuYgXfERR5Gj9MUlhqoh1s5E2D4+fH8CrcT+hRGDszmb2Qyx/P4WAfbvLbtwVArR
aonf63YPeCuCm8aqRX+5yqcEPV2ejRssuMW8z8bgzd4efBRv1km1n4OQ2EWUu9DcPWW1mWjm+Chx
1XKHYVf2+bsk1e/kBoPC17pVNSoXuBf9V0iEb2jeSI3PGjxdXwwPenjcxJqSGqcDDX9d5hUhZo+9
ne8kGy5sa7b0V2XbGF29+OCoTq6/uu4LpGgca0C6xC/RPfVyBGYCoJ20lrfBK+ppuJXHgqykFmGY
lNiINMK/hSPa6P82DvCgW5V6ghPTvm8F0nG1zeNv4Q4QUkLFxyR6cO6Bb9LvSP1JFIzDMmVrNzTW
s7L9jPTCma97pAiVbIo0iwc8V1++kVHLC7BK3wLioNvd0dR+mig3YiPJHxZkgoewTrC6ahWmTWiP
PPb83/P0SvEBJhw0vi7VMygqkOdPjuqXVnzBLN6VKpLiqj7tvdOk6u6uNrXJ9aXi5RH/xGpmPbur
ryc3rpMGUIwzOkYE4RgXtw0bmc8kOjHb9nYqIrJEONBqU9LYo6FpjdEUClgHZZlzkFEn4RMPnhW+
+vrRPiCrmBAX8JdhUFyRWATc6iSWbgMfU1wP6gxOc95zpBCK57qmlIt9bG98nLfG79T2iRInOMmZ
Mj7lYoKDIee9JFpdOH6eoh6VjuVYi3WvQJ+9HepkWp8gEE9Aq9T58my+2+J2MnMyuk8AmyDKD74n
JS5FAOBbwRob9Oaf6kM3cP4iZu+Gh9KyeTjK+HqTQJ5/Xds3rKEfnhTgPVEr3dNHctGSpi1V12Vo
3QZRJi8AOgFexCJQVQ07eRp6ogvHYk3u0sQsIrzparZTkO/bU+kv8MhlXaBUW6Y7RDMEY+pwz6xH
gKmlzbSCOui6ttGV/0VP4R7QjgLnIzzgw/2H6KQHnIIbATj3apzdmfu1JTxbgDDT4sFFXReZY26W
u6h9ikb+iMBp/RCysqAsQWniFGjgoxy6QUuKVHBAL/Bx04Kdbc/r8rtWX/Ex5flC8Dk/cONstebZ
CZhm5DbR6H7dyKsHWQd2bgjOXg4XVxN6I6wIgCdR1fSNf0E8ou/NM52ObqzJrFYHTTEmVkFxc3uU
/8nglEwBcCRXid8yWA+ZuXnfwvdYJgFfE3nIW2vOVaJxn+5hX6Xz6aPq6tTmVCdqZuXNqDPyFQC8
GIQZICrdAUOtgcYGbpMopUxmdhKJhLj0SZChb/H5+gSAXfB8waX+5/wCp7KWXL8IXTGFrd5Dzz2S
5PNML+ZwGmCimccXWQNkyEdGyOp/bby/v5I2WQV86lzeJeVOI2tQ2/1vI8B9d//Yyoi3xJeR/e6q
tCAJoV0mdqvZYNk0hAXlxyYfxuS/VF7X9x3ZjUUhDxH7qMBWUT4mr12FVI0XRvWBoY/ZVo4jl9A5
8HAk6uYhrmUD12OaN4uyN3YfCIajiHPxkjkudstU2ZJDRp4pudNw9l8s0juM1jnx3GJD3vFe7S5a
jf9WQ69AdAWHi0AmcSK43c1WLdeMQ9+DAr2uxqUVjdQTR6uDV1iitQo4LEPy8+8ftKY3lsZjcKpy
MC9YMG4djqVh3B1360GyJ9405w9jAlBKtmVvC2MuTeqTXmEVTS+Hed68HIEKO4ERmW+HE/nQcXq9
qlHkLFSBs3H+oBuNffMsV8nlRU13qz2j9pjc6kqDdIGY0Ai1QaIFxNU8Kph1I9aFhObJ+NChtm2U
zMMegr0trnVDY8Xt4afDfqyES7aa+CipQbiyByk5GBnJWgUWfPqBEBoE0Qkd1IxTpX1OfGxPiuqy
hilAPQIcVc5wjqi5KfbbA1qvkMaNeFhKCgEy+w2Vjb7OWNrsyw15Aq6D1BxO8ZtVZfMUKm0x+h7N
geESAItGj2THqtwNCwsOiSW3RXxz+FkdiJfaww/zcwqd/Zw03acMNDsn2t0OiadCkdVgoiAb9t17
HdPbz7+z8tKIWxfJEmqs3OJCl7lkeyAaV2zGJXVJx3jPSdGXE9X5k/Q+90hhc43xbf49DH6gkRrL
SWg7VJeaXy1Yv3n8OTgy8sn3GMLwKBp2UsTPlXbvCUs70JuyfCIdR70xne8kUiWAnbxyHCzIp2ic
IYWi80Hm5AXkG4H3NrWfZGM5Ab08d8yMsRrrCt1QtYDHFw/8Usy4tC5PRYlsFURyoiUNgSlwrCDQ
iPjo8T9HqRC7KROWqJ4yeiq/FVQ6NHk77GpIzEmLY+m8HTgVtcZ8iw08ewNnWwNO/KWghi0iZz+b
JgbNQImhYjML7pK7588RAsOl15MVHUEBf2wrD/+x+JZKHUBInKpxKXYRLAU/kgrO70hFSmXQbcl0
Uc0py+11TcoNB5HSdBytkTwcdshhUcsNgOgeerNSrW/TVA96h5qesw0dzB3b7O1NdBcH3UoCtR1c
ARLBR5oeLb2f+FEyhMHVrxFeUW1A2enPiN81oIJqU/zdGerDhGB6M/XuxZ3IEECvG5TmJQM3Uz9p
GC8AdjsIPxYLWDxTew3wXT8WX37lEMd5gChv+gvb7jel02ptCPPQHMxBgCMdICpLqDTCENxCRtiN
D8WumOlLvC4VQRL8CWDKmqKdBNqpQ/KtD1lxlpFbS7P+JwmaDTBB2hkW/vcuZXXQCERQFv0P6F3K
v1Oz+IuIpSEoH8o5L4rSasIF5/qZC7UoCeust9sgHgszrnjrlcGVbsiYB0tukahli96YOsFUBXk7
dUlmHT5P6ilCgmEgbx+UcPXdK4QPVuv77sizSvgM1kPnTdPN8IhSAJIL8OhctRnmpWgvZZIJXnZz
ZFk06Hj31YcqkrXQRiK0pYXoylsAsgGgiD6crjhZZuzL+IG+yZXrCdjCA+lmlpCk9+xjJSutvble
J2zjP9ZWCEKeJhWkBqmZEGA3x7ImL7Lb9ZfBLONN5mkLwTiA9FM5j488tCxMm0ZIhVxgPd9dIA6P
CprgABDfJLIGpvLAwt9Nsdebpyh4oP+EeunALvnOIS3xcK5GZ6mXykv4UT41T0Xt11dsM0fYZz5y
Owgs4RU8+L27cAWt/MjjqFSEONYT6eGbbzbhA8WOR6VuHVnu0bick4RniMsGnWX9d3hilHdQZ75g
NCEf2aBA4F2JViPMBjSrR7CZGgVV/npofOhpcBug8+vM/w6QSRPRQWI/zIuewMlRPFwlzpMZ/UPj
KGMysGHHSv3LhpLMPL5jg+XjHnSrVZIQefyN4Rfndz92X/eQt72khMkx12r/vPB/hUp0jLzPHNUB
izWgH+Ejxd/H0H4lssEFSda2QnEFl7YmYtNPdg4ejmcTMu5C0GdtKvRSE4W6j92jnM5xcmS/jvmt
CBnBQ/qjqiG3+aLaYhIqjJior1nHQI8bgbFHbaL0Fy9b83XTfy6fkdLeJXTM1RCknaoJQ23sqDtP
mKoKtn+40Za8zBbcLIcZRDW0+x2PtmsMwvJGmoIcvXnxtZWGh2whYfGrlWKwleSI58q2X+TMofPF
m9lMOj6sWGSqGI+uSLpZ+GvsFrxLQEOsyNBBQ9baktC45uwE1O8uDzqPhvxcE6AgVcSkbDGK5u5J
bNpLRKXfDTZt3pWnMRoNEFsU77N9Rvs2FxGvrJBq/4WNL5snoMgEx+93vYjSpe2jnrOMT3LL94zP
BLZQFVauUJ2MmI0amuGVs0MEDTGZ9pQWJSpukR0d5C6/XE9DPubI0uZ59Otv/c8TWyTARb2sj/WS
aBhU8IE/4yoIaLusgktrW8NxcmyDvnjFeZcqFyzr/qVDKJWoailoLOu8dXjUebSLcgAxMRcLVYFD
ywUfCbITwKonbMI96NgZsUnLUWTpQ1OiulGcfC89vTKJfNm2QNzSRJ2MSVCCM8aJx4U59BI2UU0H
cB9mLMI/RFEeCPHSYXViBzDqxLBKJxXQrIfzy3WGD8VC/7iAKFObvl+I4ViBy+FUs9qo5I52swzp
I/V7m/p5mhlNC5KxcU0zF+w5LFrbQj5MCkndquhC0cpebNvDWRostinbCFf8R7G2yze8L+mY8bQA
hooZqwUJgGuxSYtql//OUnBLiX3r8QQIHhcBkL/GOrBI5ufEo1L0G86fA9fUNGxjbazB/J+uMhOk
KuDRAEZgTVowfqGka+mL/NRRnIRO5MZ6pQBIPBd4iUT31430DZz7E1TDOaxJols8lSkMI6J5RNJ7
wx9jsV43FsFJ3XXCmbFykrIOsUgf22E47cEt5x1DilHDi+qUBRCopWyy0FUjq0a/+7ELR53E/vso
HoJXTgCakwrKnauQ33axNqngK8IjF0JspFTLUhr1L1sBWueyIsjARgBPshmXz8k7GyayG6MjyFAL
Q4iBhFuJCl3BQNok7XUCx1QiAzVFMS0veJ9IvDuSjmWwRXYa/VUHkxQjNCLIrXxZG6JjVqSuVLy1
4QSDssx/RuLT2V9RlBjYnqvB3yHYiDaUu66IM5maUfoTNBJZkzn2HHkicafJ0cXWY7lu43VuOaLO
cRChnSsde+W97Vnbxur3tTjcSmxWJHj/NUtblWDXfSwfpHnUzyIvV2M1sRti69JW1clfJjnmAPDV
GNX02JiynkdFK+yCaEET5FtTBw4W8stOE0dBu0YIs9W5jZ37jcJdcuDQa+l0pDsy5SHoY92xvfHU
c8RlR3ibSJ7O+/KXE+NLlLAzc+zzpixtm6eKFk10EzHtAOlJwcLU012eQLPWkWa1fsRekuBAtOqE
ZNMNsmnuPTo6c8ni9lZm6vyt4XaiSyJTRxx3G6PFrLaGtfgZsWI/5JUJQvSnIY+qJl5jBTmPiTv/
8cpUDp9ci61rvK0TABmf2tf7IPKiN6S8spXC4ZUzQu160kmcWQZ5mgnQRCVEqA5++O+R6Lmw7rhi
UiXirIcvr8n9aqdfepVlJaMDCYyHVMy29BPUnNrMUrj7/eqJAACb9gECZ99+umXcitgN3wfGCXA0
qNlxRqbc/qlyCDS6CNM/757sdDfNjPw/QOodTOdPTbhm3tL8Jas9QPYcDZXS+LjpvUtcejjpfQHC
07i9s8gQk++apptP7ECMGSG0npjnnH2HVy6tyRjhzmw+nDm+QMmitbovLxMsANUMo/IlSAvQ3J03
x3nstwTzIEMPacpSsFlnMzpCsnx2fdFD0fE1vvK5bHjInf4Our8GzNEK/Q6rSs9siaFVbCGTCumc
wPJS3yI5QA6D7BvEx06CP9iES2vyQPE6O7gUUtCWuRVezpcOuaXYb74P9q/EIaLygBK19YJ4zTLK
6fLqNr7tgCSjPFMeZbwI07pkFD/oyao82EvE/NOhcM9NnCZ+2BG/CKS/8ieQ5On33eHpeJG4dRe3
vMpnRr5UzMmZcCNAlb3DqiWYrvhBiz4CY5RinD3cHxG5hu+RvgehNta2b98vIhBY14s2tGcnbD7M
4IK0REkLKxGgMYbCyWIwNXygu5UBDjumvpVdh03OF56gD6WWWfFlaFxa6C7JqCsnagjRLjpUbLHl
rgULI2T+xd7jw/aU6ZUdvY6ka7B/F9JhuvJ9/X96EJn4Uc1YNNaE9DsiZ0eMHb5pNERV28I6EE4z
Rvy6kX9KZ15Iwt06Z5+kM/FXu0G6cvImAoGoWTBvPGarlF3PhSDyiURwPnpAl3DzhIu3W90E5SCH
4n9UTsMANWkrDkWRkvPNgCXU1QULfvkHgqdDqj2qEAUrcMV+BXPNTcTE/h5RtfRJG40czwD53Izr
ERyuX/okF8fRQB/oHHRoZpTY4MjZ2nt29ar2B6vxUqmH4fwwDxR2kjvymRWVtDZZZCgXD1WR2Mfu
6DFpAZXf1YVtAE0BtnKHZlUME51ORK/875ca3QatkqCmOQ8HaAOZEYRQ8ydnNbEQgo4QQmfLkK+K
BYcLjOkiRJUPSzS7ZufsabPgoRrdxDNfpdR3IH4NYmp2xhVZ8cBBuZD0Bb/jvZf9JZx3U2nGlYq6
R8dXQjLGiJyem5Hn4p5KZtUxqvdy7ZkcDdfMPFiMveXGOJdr0bAVk2UIzBLKw+k/PlOa/XtlIWPa
Mhb7nZjqAzYzWlBS0phfPC2X6eo3STLrkHUiIEwgBXDgPaEiVd2/JfgOPRqprRRFzqnk8NZ41uau
WGTwj8F5DmnMGXVJT+PpGBvqATUC85Hvk/954pM1VjBvW7tCGR2VMc//Z1JOgMIbaTEy4lL9Mkjs
T04fzR0V4tCNHtRL3qtMSbPADaPkQvcSDBF6H+8McTtLqYwE4/V7xL+7zQ2YvW0GC8B0D+mpVIcn
gzTzl7pTWHN0rTJW4N8eVt2sJAmcHnXuZrOHIkLRUiOom/JU6TXqh/H1H6xFRRSsnyjUKAcgfLp6
itXiKU3UmbIxWlMFq8/owIYnTykNTABGR+ynZKXZ7oa9rAlJzK+K5FFELXZ7ENHg9UtWC4syx6rx
pxA0re2vXafwKmPYUdhimsMo7ZfjQOs6R+FXwYFubL8jLYmo6fYOQXAPuEIMPKUHO+L/HZ0SWyHR
MeOVqSYRyOYBVUcffdVIhcW8RE2juqZzTGrRGlnAbXxb3TXccpzWjsm3Yx0o0gFr1PNKJGBCx/Pg
87NeJtKffFwtkzwUNlVXBeYlEhzUPbuivXdF1IZ2ndLm9hMhsNJcmAw0TY65riXNpu0/uSHWGJX7
cLXfOBXaX3cZBFLHePBH5YYc7WmJ5PlX1cbdg0SfBQEnZpr7jftBxOhMjDRK85kSVHDamMaKO2nM
JGIczGnz3LQOKiQgmeP+iIH9N9r3abNrXz30RFG/CjSCyajgt65GQ0123twc9sa8cQkbblOzy6Sa
Gtki8CkC0ov/BAGm+pvwEurXhZz9boFlSTuHTPlrtxvTukAQ9dH3HBaqStADLPCTj2pZL7gm6l0K
wDXiuAuzIUIe/5OMoJxwZ838OTRyYK6If/PLQXYtsE9DRnxj1tv+iLxsi8sZp0naDd+XPuQdLbMn
pSDBEBQ3/C2/T/bn/6GlNh89zFhVO/jZQyugL5cvykY9DYGfZdcjPKGuc0e0nAfbi7IYBMzZpwnI
mUAMzxbPbEXYo1BWfNOi/dQ6NvrzHoQqs2jP9y196Oxn8gomLCdtbeIdnoSKepWXkPQbJYd8CAPZ
kSAUrKr1MTZk/stMV+hIH3mmFaePA9TOFNh/GZtXkV0xPPE/ToRWzIqH18nyjq2FpACEB193WA93
YAtBOojVQ5mnBuA2aw6NA2se4tPcbwD3U19wkW9TT3U4+OCA0ZOH7JCrLYxz27nGVgxx/Mgkr+Vp
jLfy9b/PW+llPRndh97Fs+z6ctMfQ4OhLNp9/tBK4UsIDZfhP5txmDBnK37YjTieYFkIBkpANtYq
sJWT+keiR2GjEai3bberOFWZu2jMch63iY6clsGJ2sLE2LZPsDkTK7xK6c1ZXhDhnUFh10P/JNw6
AQdawK67kQ9cBBQ8aT/uuYRdSbaWc8nmbNSYG+r05S7QVqvfdqhSsy1ifsD8r5dtrtbLaAzqjI87
LUsee9JTzNVPXV9dy+kgx6Ee7wdP0ovzaWJWa0T5GNNSCxDypYMq2a0t3dIODHQk4wg6t03mS7/0
oUlH0O8jv9+FJjS6umnH22PyIo5skZ2zCjKqX6OwWCP+XtJjsd1dbQZ0YQ/WYiEIPQtr+UV9+qN7
ct8ivGd1pD2wy2LU0WmHJ0mMwPc7wAPOCjvjJ8emMYPN6VF606LlgalKhgD/V9LMs9ONmOpTty8i
P92YATN52TgmCeImPUa1prgcOO2rxUH2ztLraP1zWVbTssrVrhqsJMfWJYdvROr4Itb4a7Tmn5aJ
7qptR7M+zzRKUky1qXhACU4BtpaArXazkI3wBdziyAfqiFx98ue5xaE8WLjNVnmi/aDclzxTae7A
F286Z4+hvl2vYy/37Vc3+Z5kt1coutOvadNa8nLJU+rXi0XI8J6N8AosgBBlTlOoB/orehMaih68
swCeHCEEYLdS+QDNHGW6y5akmgrv/X1yPB8FUp5htVsgY09Qhyt3XlGwn7+KVzSqJbSCdojdWUfr
9b7Dc73tIauM2DWajowrfyH2wedNCxb+e7u1FeDZXwBOIOMYgOWJayicvu+I+Ugl7g1aBrRkkkCt
4j6hhVnWKoqAx3XZGrhoPWZIO6UAaQ2iPeZExIVgKXFrYN45LHp9hW8PnC2Bq3n10tKFrPsn7cI0
lWPJflSM4rsE13loY1C3EFh2+/2v4ORDoj+RG3aZLTyZ3nV9cmige6pqEHUFd64v+pGZPDGuo0+Z
sdqkpUb47qxhOdQu8DT6jDvRRktFSz/qa8A4IKkvgHuHW40krh8ayKtmZUFw5/A1Ffc1RrMoBCFM
mOuW+chAVDmICcvB9yzxKjcOHiVih1dd6l0XhmwGC0E29fcRPZQcANaaQM+zcFKhfRtaOUztLgPz
84ISroLDn/tl0KgH4HN5bVZSCikNWw4pvpPqwh96OI54AdPNV2G1cZlgFkqtJcYWx92IbXbAkV4O
0sapi1Q8NwpQYO0kV81i0EJj+2QyCREwyqQWhNz00R9G66rgAoRLuFRuRNjqWz3m9NOCMeYpQop2
0K6GTw1cmpeWKti0LVir0iXSKF0T1Q1dm5G82Q8cL+qLuOzZeRGeuHz8AsgB1DQHs7zSiB73s+Lv
oAxso/tigPcSo8P/8iL8qqLQW76SHNV1o4mplFO/+JgzZvFeVO7ToTKsYgVTvnVz880TpnWQOpWY
zqDtplvoaJtam4HAPoAaWrAUJxlyobbb6yfeQdLvhlTZ3XCek/n57Oc4rsOo+4rXdLeUORZTnWQq
+6R1YxFkAC1hYg1jYi9ClvS2O+G+n8LavgsXXsUqB/sX6NAUWX8Yn0B94hJhUSPqKDd0CxpF8TPt
WJ7kSht/3vCRHMLgNKzWbaqxG7NcSCD6mEa+eUPE3/nPAlXiQabeqDRNdsRMo7cxXxBWczyGSBoz
2YvgTneGbhpCQvuOS2BJpg0j0jRR+sdKyAXS6eCqnLVUMDNtLABDWIhrAAL8oW30YhmmHGqTQzIr
ugK2bD+XpK9rk+6ea052ixbK7AOc/EMffmmyncfj6ChKbXD3XnNYYg3EotkNLqlc2g+73vgj2QgW
Ai6dkqmW4LeVupS49S5TJwj+xGSLwU5688SwCsVmRUzNt7EdIbcGs2uYKPcKBIi2sBzlQBq94tRi
o2xqiqQYLzZ2wo0Hgc5P5BxlyuNlg1xp1gmigaQpnUxO5NTURWPxhJccR1Trr7W3bVwdeGqYbSp/
eN97zna+5IvvxYztmxwt9xwqWzIfFo5Nor5SfHkA9/h0fWb3hvVJzcNsH/lQ72TcjNzTM6ZMYf90
ydE2MTc00SpzJsttcdA58TyfF2NHm+HdXXp/3AnXDe0wWuQ1sQqISKA0XqV8QkUH1DzpE+DW8h8D
wM6f43X1hx25CqXPnOwR8W9YE8MaYvngJtA04RH7bVMkVStAFZJ8jpNDt+6Dxx44LXRux7/+CQ9J
GqGs7jKxoetOJaEB1xataSSv0cGDfYi9MJrz4x+LhH7xBTDarH7DAfFXBbck7D/u8QbJkt8PUZuy
B2dfu0WIW/SfEsd+kGMTJIje2nGCUVodmVEoJKv650tNYYPYtxmQ+WFExGmszovnyG1KtZnIGedW
kcY5YdiOEbj8q9NjwQPok8vQYfe2bbMVLJ9xV6M/M0VRhB3REUZIxSVM+oqfexim2DWVH3edFQav
zjOmeY74P7arzVNAbJJVECadmMcwpKthhPqyZy0+QKbwPOHiCtRQAtJezy8y7iqQNlOxlJAzWUKZ
NA3HLTQaV+E/dcQsoaFtn4KGSNdQrYtMH9OPIBxfVfOZiiWqayE2PxXRhx0U5wveTqzxww0wL/37
CaZBmIXoMEgJmjBTM/5IR3un6zF09dFevcFjfkqukb55lxV1es3simxFsoyHx1ahd+tJLahjRB7M
7pI9sC7wU2MZ8lfPQ02aR2Q1fR+pvMVAtrO96c6ZCBCOqmJf793o21AYtv21sjk9rYCex7/NnOrN
l50TPdRpVL/TsRbBH6AIfN/ckVBidGnlC+R6zJHwDZq11fbJrN7+OU4b8l5RGon1EK2+jQ44mL3d
PLLgXulkHgCHIjrcki8TRX7b4h64dBo5yZLn6Vy2bC6v9pW0lpMynEHLotnYjJd8TqA/WFTsLEaN
rb5TZ1brGkqXMtwTVJzmg+m552rSW0HZ8s66fB/38XckSkAx7u4OzXyBUHo49PTevS+h+HrbJLUy
MwNXAKQ6WlWVcyLgF6HkMNqLLGnKRj0BpqxeR3ysJITkqZHKEg1n0900FtX2LsTQTCz0OpyzXhu3
iFUyj6SqZOtmZ3UmkJQI1gYM2DbaTWuQV5y+l/nYF2iOqSB82Y41LTU6+HgLe+DjUKt94leZVYVK
qfbQ0ntuEX/BbzB5z5gOAF6EDzDH+mhzcExSJpwit0c3syrAGRWyv0hL5aftWb0UbvksjDK+E8kU
Nne6iIanwlZu78Ntu7172JrQpPix8gu+VXPQoAclSO10fyVmztiMtBTGaOsQRHIBY+5IxqDDjUs2
iZgmJKPkCFfzSfgKQsgjSorAaeL0woNknyWPJIZyh+ji747y1ANJsjfR2sqoyZ/bxYDHXn++/Y15
9k1FtOU9wBL6r92McyTvb9XSJIud71vMXaSyQs2XYFta4BmH4phP2yOaEvI5zfN3rSCYvsQ4PCHw
yeyRkTXh8pKHh5il7qhR+ZMEF4cUd/Gp4xe51vMNtiTVOFaSr5e9sCgSEnXIaX++kmqr+6RgSIgy
4QerWQ2gymE3crKXaUL1PZScj42/tyQ/h7jNAMTW71zpK88vuOCbj4y0VzSdE3PzHHc+21PXnkf1
v1qGSpTJSAxl7nhef0YiEVbD/6ln8m3AD/NzU1lj3hh4erH6lPs2AvqV7JRt4mcQ4WkOgpLRjlgD
QnLXYImamAYRqQhPymLDil3PWmbbNn0uux3X8+PTLmOWG4K/vS92bFajYkDrbnAHxL205EVyIG3a
uCwYtuAxv3tlI4t+Pbop+Y7/W1uRlvHzrLtodWvMwpSy/d+pZusikomZR6Z4iTi3ixpX230TI5cL
kaihhZYUHVC+MAZu6aMSeUAREIrEvbVqiRcgEswo7jW/AwAQDFRUHZdSb74p6Y9nNAAKe+lnDdOf
OArxm+QAL2u4sJoL26X3LKd0CEnZ2iy5iCz/JWUPsERRTk8KhG8G/TE7xuTAldpWc3KRyD9IJ/aB
JK2QVgZ3vdiMofinw+5IbTSV8gXVu5RSRpg218S1WMP91nGeB0LQWXEFIK8klI7QaNRqxAgwR8DV
5VXGuKH6te1UJetn+AyH1C/DbL9X+4Slu6KkSYkFRt6EGfo0q7cK9vHZqNWSt8e0IpBEi/Aq2nIt
kfS1oRvyckZoFyg/44nJEoju6UVjQJiAbQr4nzKdY/E3LxY8mcwTIpkWGek6nJ1BSie8FZRsTFcj
Zfl1SIMDsHIBZzIHOp20GZmlbvTg3QJaKPBhK4bjQJX2CorUZSvPsyfBwS2tXM0VoLssXrw7uKk3
JzzFYnuWRv4rgMRbCKOLD1lzotQSIJJqPl7pcQ20dIqwt6WBmGXAi5+o8cY7NR3zDtXDaVZc0kxi
0SXcoGfP5podiPM1Wxlsg96n9nzfYDZ75W1TVvRSZY2QoQty33h3A4BpEzn0fIXBDsSgQO1A9VJD
FaJCSRsCcx+18U+kX/fUrMZLc50QOXxZ7jwxULDZ+F4og91LV3dCIsfs9JVPgRq6zq045XEKT3uy
ugzqj8nZ+9FCD0+FqcpmAapo4obJV1OdaJkSw6/owBcNSalXadgbh8oJPhSH1UdYYBzls58PZJ+d
Fb3Q9sfylRjzfxx4/ep0DGkTYE5A66rV7phDrEkst1tEAMdeoB3CVMYZhnqoDOhOhiyyBl/HB2pO
ypE19tYzZafwMWvwu8Bi0B3GXMsNYcCQOa9xT88DMukGtBDG7Yk0W+d7N1OJy1GbMY4vISbJ3300
ZlGReZvNJSoO2aKqQOGIgXx95Q1bwuhvtsu+7tWbAEg/+rWq7igprt2IpSD5tSQAumJugns2Pw2o
0NVs8Tlr4C/0Fco56CgEIKSogdfqoxB6ktpA0wVhHJkb1BLrUYjAibRMdiXNh5Tk8hI69fFnDzWg
gJX4Q0Dh9QD45wB3gAeciVP+alklrx2KfwQHE1TrSkb1i7M1AVTWT6OU9TvyMYHZbUS45WuhlUjr
tRSv42b8zFkMS5A/F3CshABhdFUvYdj7sCqzhd7zn5CoB+k5ne0e6NupYZ3t1Z2tMWRBEWj4lawy
Vg8wAJ1iJ7o4179plMmL36dD0/Nbp94PFf+r1Z4AHwFI5kefnuaPYzvaJhZU0tq4LKc+xClFbi7h
esVOPMJwxpd3dOE1js7LkdshMn2Ne9oaY4SmgiPUanUL0vTwJIvkn/EDp6AlNIi2cumLBG90hUtV
klFrfksPbh5IwI94uBqMr+dNrBZt9r6YKSrfe6rWPrTg6ZGVF4qE16IJ4wr/aopYxHpfHp09RwFt
hzRR4Kl0J246r4wjY1BvAW4zagxeq96ocK0K+80UgdpXzY6qeeQeOfm4E+GK7D2tMlyDC2xmOoQC
Xkuw7yKvPP5KVjJXTQjghEOof3PACAhL/LCqtgsp5IHqmx/7XI3fNhMGr2MQQ2aF78MVSblnIMn8
qUD65SgpHHKjg38i0cTdAr1pm+U//RAm7uMeh4RGal1Z6183LhA1PT5ChuAodg85qeF3HL1jtV7V
r51Hl/1ct+maTj96tjZA/2h1BxaVJX7RAobZtEYDarrJmZ+y0UGMveJz7uj3RZL83kmTZILhhvne
5TKcYEzYnvOEhtThqBsuxWMcmVFY4GifV7HmXbiqQKA3NnCZtgxulbeQG1+XyABWUApPAnLGualo
sJMU6WAEa93F6itLxIZ9GBKWHYieNkcpYNIoftk+PkYIqGf+nzW79yruSeSGnt9vBTXxhVp9TiFG
W8dWFIT2mDZxVdk480WriGGlv5oVC4XjIz9A18cj1i4xk3XcOJ+SLnr6zGMq11m1DqAhw9mOe5g2
zaUcEfbFIE+hvF0x3UlZf1eoORDPp1BG7s+E9hHw+MNHi+W/4V+cwtB0CnzxWhq1zlrTPG8XPx89
l8sQ9BJ/82WxNRuzs4jCFz5NKKZ8vQvYue2p9UpMFd7pn098kkuy8lEHv0WrHHVUQwgH5YZTzhWq
KXwBmXJ5jn2B9G1mzEPkvasMi4+AUrERQfiCcPdybESwQZrYppAIdRn8sC0X56iDZ4MgcUlI8DLB
MUJegCPmtVQOlc/o0OhWHm2LyD8sVCx3t//CgKAbuOXMcE+cnRBezVbG95LjH1xnyGKkkECNQY91
4LEr1btbEpaWeJU+Ctd4Y+kaT1PsR5/ERbaPJVRWJeA7ceYq+cKG+dA48hrmRmhW+XQf3541EL2P
jSuZsGN16U3Kxp54ATOBFempxu9FLpafOPhJyzflKiyMHwiM7P7OFUcDG/TJ7GZvRwzaXoQESrtl
TK6x6zznRsJonnpn7ry5FqTJzIUVqc3feoZgiqmGxoJKOp0GgXXQIn5yp65Dj1A1/+Y9oy8mc9Te
BR2Q5c6dOIoeeOhZ0nypY+N4+jrmg7+gZFvekALucnBNFqgdMwZGvS/wcW03rybAe0TzR6QFkIGo
t3PhdwYlnDM5Tch/6lryqkZca9CEkLwIfFdUfAyF+nBjUSh6fk/x9MQA9LBtEPasgemJ4Q12im5f
C31Q8vcd2PlohsAtUgEwHz0a0Qg3S92pWyG4lXnt6EOPtG9qXGiYHuo1FYaYBLG1VRTQ2ddS/lyE
HGnu3lN4w8bIGcn9RPdBaie1WroE99/H2hQDcfS4D72QxnUNb2BY798y7vaV+vZK818FBA/BVO+N
Dzlq8wyAcQ0He45oLqUvORD79J49Dudc6iYsSVoEXPdfU1MdQ4dt0Lyz1uQ2I8eraYBtgFm2N12y
UdctuJSisscsdOpPEGEnEcvcb93JHQh7FJZ6smEcXcCBI3rhufbffdFPfEBcywD50bJAtnZmcSi5
bkaiL7GFGeCGnqa/j4XkCPD2GjcGxV9f7Ai47HEggckCby9FDGic9z9H7goS/Ujd31KkddYrpp8o
gR+F0E4RBoA5yuV1KfF8kmgBSDI7RJXHStUEFdKRsbBEx1B3C4Hm2C4OqNuzIPS1sg1M1ffVZHdJ
wV9rzkILk6MbSFaS/qtksh+1HRvCCIMI3ScOmXDl0VxuuwlTkc4C7DoyWACeWSJsQHj+oN+ds+1C
5OX3ep8Dv9aNgz0bNzwLlNBWfUlRg7s9doQQDgALZqQwSef1qk1AK+pT9GfB94HVyOgp23e684x9
zXhzNIWN7acw2pVNnb6pt3I7SVmz22cwhYOco0EzZVYipqh+dlyZKc1ovopiAp39EvSLJkwKWwz5
plB9eaC3Sk/bxEsed8MMOoHGYdWo6wtEndX+aIt2bbPiIA0aTGiBu9y4cB1WLma4J6mp4PGaf5c4
wQyUXSv4R7TYkHFEn0+Uu9oS1nE4HuqLwjwGAiyStrJ7QABe8PoWU3lagDVh6xkopza+ENT9epPo
ugJm9mSbwH0ok2guvr1IYOsDc83MgM4ecu2ii2pKmTjw4p8UasyNO871Ol7e6BcvaqmO9o7Hd6zz
NT0BxwZjFD1vX+CVAD2rdfgI+84fVWv7llPsfS9CIPDS6WKOe0aCq0i/I09RlBcRSha/xUgk93gV
xOIeHNxfiL+yi8FMGT0tuiHNP1kra7hEed23qU1f+bdAzXXRefzQOmkaSBha7U1a3jPluX2WP50r
TmjC45ziqQ1Ge7ffcvWJ/VXaf5qeY44H1+lI4/doDB7BbL8OYd3M98WmVDYlzWpls2TUN3PqUPSJ
kpSyiEaoBENhQr2PZkPbNhkTane2FIZJmqiviwxPY8hhLPbhRyPzf2N6DM7lEKNlilDt1WbtVKBi
KDEMn4s3bHhzMIN/Mp+mgK7oQTda1yjk5SJfoOJC+fexREO/p1Q2IINruMTi/UovCOt4BjgTidMq
0kWJ4qsh30D/2qD2+5XTcztXemxj8nv3kSEYEH458tURXjwPbSeIuhd7gzp4CAc+RrkIub6hQRgZ
QLARAaSJm+2fFoR7Ljxo34CuEE9o/nV3ToKyz8GUopnAer8tfFE6AWT60yd5pwT8sqraoP/qbr9+
zNou5zSujSvlFd+0Ro6Ph4Yo59Qg5TXwKN+4C3KNHeGTWQjhPHHdAN7+10P1KnNQG3Kcf2P0YOy1
Sk+vfod9/Y4Jby/ZhG/7b0eT7v5lBztL8cALJ0OmVSXDyu1z8XUAj3e39JUq149qjKPukiQ5o8Xx
I7w1cg+kaYseDjsRPwM/1G6p4FRCfleQKuLkTlzhbiGmTfBQoI5BfnW7XAC8rNIj+i/wU498gKh4
bYBWjagXeyxLKF7tAQtOYhMEJhTknOWT3ERBlWm1CRjWR/OMVWFNvmk0Nf32D8SioQOPB9Lec3JW
V+ie9XLO/uaiHCt9tX8hLdd3CsSwuszTOBGT/mmKTqREn4aeFZUgsbEHZyQE5MOm2X2oYv7c9xm1
uPq3jtPZiYp1jBlkty49+aMKFS8Kk7PQ2vTsgbrop8Z38WYfgCltvSqvmU+oFrZLEziorft+OM17
9s4bYtcD+LKcVl++N/Rwd+Qd4yP+xRhVqvoyjGcj0gdu2H0Wcksk74yyfKrAF4q4PZ7byO7/aGv2
CJbFud86iUB8ftfxSrt3jwBC/zb+D+NVd6/0WOs9MhgKFWJmO1eMZeiU674u3O+3gJzOIXrdJdC9
4YNWy9Pxn/s8+DeywMTIyB+uVbHlldXd8SmyQFP00w0BzYvJoRiaNB76apU023Si/lr8Jq50QJC2
pywk3rMqeqVmO1Pyte0Ed5KI9TfIqWmkOCjP9XUKx57vfBQjTyZ9gkbBeVxn0ncoOe4/Wu7glDVb
VTHyJsbfL1gKkK14ysO9PyzcbRK7lHO/OKghskl9K10InqBGNktdjOimMe3P607SL2h2ZMaINBSa
rr+lMV+mhVg8oaOMMHKFD4CSm8lYEd7e9wIytpbvHzMGB7BQQSSpqjzDm2K4Hhol7nh/VREhVh1x
E4B/Zx5xegZFHexrXx42pnZbzeuPjy55je8i0yJi5IBpB4wKKRGyaY47a0EKE1MqSp8dOOHUSw1Y
4IUKSNartygWD6AU9gQA3e8qidnwnUI4sQBmJxu1TtnJH8aQMWadaSKukVvQfbkKsY2mXCqiyeoy
1PtxBfIDrL2S1r9QVn3eSuylaUff6U4NjhmaNxD/4ED4XpWQlHwWgz066i0kaXA/kpjG5QJG5S2R
iSjmX717WDgjdFoXDXCCzI9/vh/OZBySfNzRl73XOlTlUX+SO64T7BONf5xd/ORCYKM1UgR58f+f
7O0Pa+xpjDrB3O7VZ/tLqZwnrLaEcsorVfE51bZp1FIQIkPsA3ykZCodUA38eXBOiSDBpgsP9Yi/
OctewhZza0by6mYa86kI8gw2ZA/ovYZfHKyUGA56HiDWqg+5C+8zSuFem6auNDlrCQaA5ubXvUOF
6faOaxraLtIXRPo5N03+hdmNSHeTtU15Sb5g87DdSPZf58p6G47lmLqlaMLLCTkMd4Q35fzkA1Nw
J64eGDjRyE1U2grEEIA3tsUHbkcSxkvbCXNw3nJ9SaIafegU2YRkyMAmnieZqwV7QVk9YxnLuJhn
OcQWJLgP8ai2b0e/eEutXiXBzBOFTokyQlLOs0+pwW2LJN1O6eZIM441JVqg3YAO97/abi2DII5N
9jgCskIW9LMKfsTSF8HXmzGI2EIyRskmsDQaLTw=
`protect end_protected
